//
// Conformal-LEC Version 20.10-d132 (30-Jun-2020)
//
module top(RIde67cd8_3982,RIde68638_3981,RIde68f20_3980,RIe5319e0_6884,RIe549ef0_6842,RIe549770_6843,RIe548ff0_6844,RIea91330_6888,RIb79b4a0_271,
        RIb79b518_270,RIe5329d0_6883,RIeb72150_6905,RIb7b9608_246,RIe5c6738_6786,RIe4fc9e8_6393,RIb7b9590_247,RIe5c5bf8_6787,RIe4fbcc8_6394,RIb7b9518_248,
        RIe5c4fc8_6788,RIe4faf30_6395,RIb7b94a0_249,RIe5c4500_6789,RIe4fa198_6396,RIb7b9428_250,RIe5c3948_6790,RIe4f9388_6397,RIb7b93b0_251,RIe5c2e08_6791,
        RIe4f85f0_6398,RIb7af720_252,RIe5c22c8_6792,RIe4f7a38_6399,RIb7af6a8_253,RIe5c1710_6793,RIe4f6ef8_6400,RIb7af630_254,RIe5e09d0_6767,RIe4af828_6445,
        RIb7af5b8_255,RIe5e1330_6766,RIe519818_6368,RIb7af540_256,RIe5e1ba0_6765,RIe4b0200_6444,RIb7af4c8_257,RIe5e2488_6764,RIe51a2e0_6367,RIb7af450_258,
        RIe5e2d70_6763,RIe4bdce8_6441,RIb7af3d8_259,RIe5e3568_6762,RIe51acb8_6366,RIb7a5bf8_260,RIe588848_6840,RIe4bd310_6442,RIb7a0c48_261,RIe5e3e50_6761,
        RIe4b0a70_6443,RIeab80c0_6897,RIe5331c8_6882,RIe5339c0_6881,RIeab87c8_6898,RIe5341b8_6880,RIe5349b0_6879,RIea94af8_6890,RIe5351a8_6878,RIe5359a0_6877,
        RIeab78c8_6895,RIeab7d00_6896,RIeacfa18_6902,RIeab6518_6891,RIeb352c8_6904,RIe4340c0_5995,RIe26ce10_5604,RIe162368_5252,RIe0d89b0_4811,RIe00f6b0_4415,
        RIde415d8_4022,RIdd731d8_3637,RIdba6bb8_3248,RIdad7918_2858,RIda15da0_2441,RId95c8b0_2053,RId88c728_1664,RId7c3590_1267,RId6f73b0_878,RIe4333a0_5996,
        RIe26c000_5605,RIe1658d8_5248,RIe0d7d08_4812,RIe00e918_4416,RIde408b8_4023,RIdc72420_3638,RIdba5e98_3249,RIdad6b80_2859,RIda150f8_2442,RId95bcf8_2054,
        RId88bbe8_1665,RId7c2870_1268,RId6f68e8_879,RIe4326f8_5997,RIe26b2e0_5606,RIe164b40_5249,RIe0d6fe8_4813,RIe00db80_4417,RIde3fb20_4024,RIdc71610_3639,
        RIdba51f0_3250,RIdad5d70_2860,RIda143d8_2443,RId95b1b8_2055,RId88b030_1666,RId7c1b50_1269,RId6f5cb8_880,RIe431ac8_5998,RIe26a7a0_5607,RIe1615d0_5253,
        RIe0d62c8_4814,RIe00ce60_4418,RIde3ed88_4025,RIdc70800_3640,RIdba4548_3251,RIdaebc88_2833,RIda13640_2444,RId95a600_2056,RId88a478_1667,RId7c0e30_1270,
        RId6f5100_881,RIe430e20_5999,RIe269c60_5608,RIe163088_5251,RIe0d55a8_4815,RIe00c0c8_4419,RIde3df00_4026,RIdc6f9f0_3641,RIdba3828_3252,RIdaeb0d0_2834,
        RIda12920_2445,RId959a48_2057,RId889938_1668,RId7c0110_1271,RId6f4638_882,RIe4301f0_6000,RIe269120_5609,RIe160838_5254,RIe0d49f0_4816,RIe00b330_4420,
        RIde3d1e0_4027,RIdc6ed48_3642,RIdbb8138_3227,RIdaea590_2835,RIda11c00_2446,RId958f08_2058,RId888d80_1669,RId7bf4e0_1272,RId6f3a80_883,RIe42f4d0_6001,
        RIe268568_5610,RIe172718_5244,RIe0d3dc0_4817,RIe00a598_4421,RIde3c448_4028,RIdc6e280_3643,RIdbb7328_3228,RIdae97f8_2836,RIda10df0_2447,RId9582d8_2059,
        RId888240_1670,RId7be838_1273,RId7064a0_859,RIe42e8a0_6002,RIe2679b0_5611,RIe163e20_5250,RIe0d2e48_4818,RIe009710_4422,RIde3b728_4029,RIdc6d740_3644,
        RIdbb6518_3229,RIdae8a60_2837,RIda101c0_2448,RId957720_2060,RId89b638_1645,RId7d2338_1248,RId705780_860,RIe3f8a98_6047,RIe385d90_5583,RIe182a68_5243,
        RIe0f3008_4788,RIdfc11b8_4469,RIde5ad30_4003,RIdd93500_3608,RIdbcac48_3211,RIdaff2d8_2817,RIda2b970_2422,RId977f88_2027,RId8ab538_1631,RId7e5f28_1234,
        RId71bad0_843,RIe450d88_5972,RIe386678_5582,RIe1bcc68_5184,RIe088e38_4865,RIdfc07e0_4470,RIde5b618_4002,RIdd93ed8_3607,RIdb62338_3285,RIdaffda0_2816,
        RIda2c258_2421,RId978960_2026,RId8ae508_1629,RId7827c0_1310,RId71c2c8_842,RIe3f8048_6048,RIe386e70_5581,RIe1bd4d8_5183,RIe0af538_4863,RIe02a050_4392,
        RIde5be10_4001,RIdd94928_3606,RIdbcb530_3210,RIdb00bb0_2815,RId9cdfc8_2495,RId9791d0_2025,RId86cf28_1704,RId7e6798_1233,RId71cb38_841,RIe3e5628_6050,
        RIe3876e0_5580,RIe1bdd48_5182,RIe0aeb60_4864,RIe02a8c0_4391,RIde5c6f8_4000,RIdd95288_3605,RIdb8a760_3284,RIdabee68_2890,RIda2cbb8_2420,RId9799c8_2024,
        RId8aed00_1628,RId790848_1309,RId71d330_840,RIe3f9e48_6045,RIe387ed8_5579,RIe183440_5242,RIe0aff10_4862,RIdfcdc38_4468,RIde5cf68_3999,RIdd95b70_3604,
        RIdbcbe18_3209,RIdb01498_2814,RIda2d4a0_2419,RId97a238_2023,RId8af7c8_1627,RId7a41e0_1308,RId71dba0_839,RIe3f7760_6049,RIe3887c0_5578,RIe15c260_5259,
        RIe0f3878_4787,RIdfce700_4467,RIde5d760_3998,RIdd963e0_3603,RIdbcc7f0_3208,RIdb01d80_2813,RIda2def0_2418,RId97ab20_2022,RId8ac078_1630,RId7e6f90_1232,
        RId71e398_838,RIe451670_5971,RIe388fb8_5577,RIe1be5b8_5181,RIe0b0870_4861,RIdfcf2b8_4466,RIde5dfd0_3997,RIdd96cc8_3602,RIdbcd0d8_3207,RIdb02668_2812,
        RIda2e760_2417,RId97b318_2021,RId86c4d8_1705,RId7a4bb8_1307,RId71ec08_837,RIe3f9470_6046,RIe3898a0_5576,RIe15b900_5260,RIe0f4070_4786,RIdfcfc90_4465,
        RIde5e840_3996,RIdd97538_3601,RIdbcd9c0_3206,RIdb02f50_2811,RIda2f0c0_2416,RId97bc00_2020,RId8b0290_1626,RId7e7800_1231,RId71f400_836,RIde5fec0_3994,
        RIde4ec88_4006,RIb7b9680_245,RIb79b338_274,RIde60988_3993,RIde612e8_3992,RIde6ad98_3977,RIde6a2d0_3978,RIde69970_3979,RIde63250_3989,RIde62878_3990,
        RIde61e28_3991,RIea90778_6887,RIe546890_6849,RIe546098_6850,RIe545dc8_6851,RIe545648_6852,RIb839848_152,RIb839668_156,RIb8396e0_155,RIde5f3f8_3995,
        RIb79b3b0_273,RIde4c8e8_4009,RIb7b96f8_244,RIde4d6f8_4008,RIb7c20c8_243,RIde431f8_4020,RIb7c5728_242,RIde43f90_4019,RIb7c57a0_241,RIde44da0_4018,
        RIb7c5818_240,RIde45ac0_4017,RIb7c5890_239,RIde468d0_4016,RIb7c5908_238,RIde4fb10_4005,RIb7a09f0_266,RIde49300_4013,RIb7a0a68_265,RIde4a020_4012,
        RIb7a0ae0_264,RIde4ae30_4011,RIb7a0b58_263,RIde4bb50_4010,RIb7a0bd0_262,RIdbee210_3713,RIb87eb00_69,RIe667bb0_6885,RIe667f70_6886,RIb839b90_145,
        RIb7c5980_237,RIeab7058_6894,RIea91768_6889,RIdbecc08_3714,RIb87eb78_68,RIb7c59f8_236,RIdbebab0_3715,RIb87ebf0_67,RIb7c5a70_235,RIdbea4a8_3716,
        RIb882ca0_66,RIb7cade0_234,RIdbe9350_3717,RIb885310_65,RIb7cae58_233,RIdbe7d48_3718,RIb885388_64,RIb7caed0_232,RIdbe6bf0_3719,RIb885400_63,
        RIb7caf48_231,RIdbe5a98_3720,RIb885478_62,RIb7cafc0_230,RIdbe4490_3721,RIb8854f0_61,RIb7cb038_229,RIdbe3338_3722,RIb885568_60,RIb7cb0b0_228,
        RIdbe1d30_3723,RIb8855e0_59,RIb7cb128_227,RIdbe0bd8_3724,RIb885658_58,RIb7d00d8_226,RIdaab098_3725,RIb8856d0_57,RIb8263d8_225,RIdaaf0d0_3726,
        RIb885748_56,RIb826e28_224,RIdab2fa0_3727,RIb8857c0_55,RIb826ea0_223,RIdab8e50_3728,RIb885838_54,RIb826f18_222,RIdabcf00_3729,RIb8858b0_53,
        RIb826f90_221,RIdac3788_3730,RIb885928_52,RIb8293a8_220,RIdac8eb8_3731,RIb8859a0_51,RIb829420_219,RIdacf650_3732,RIb885a18_50,RIb829498_218,
        RIdad4fd8_3733,RIb885a90_49,RIb829510_217,RIdadaf00_3734,RIb885b08_48,RIb829588_216,RIdae2610_3735,RIb885b80_47,RIb829600_215,RIdae8268_3736,
        RIb885bf8_46,RIb829678_214,RIdaef720_3737,RIb885c70_45,RIb8296f0_213,RIdaf4e50_3738,RIb885ce8_44,RIb82dae8_212,RIdafa508_3739,RIb885d60_43,
        RIb82db60_211,RIdafe630_3740,RIb885dd8_42,RIb82dbd8_210,RIdb03b08_3741,RIb885e50_41,RIb82dc50_209,RIdb09d00_3742,RIb885ec8_40,RIb82dcc8_208,
        RIdb0e440_3743,RIb885f40_39,RIb82dd40_207,RIdb13468_3744,RIb885fb8_38,RIb82ddb8_206,RId9d7370_3745,RIb886030_37,RIb82de30_205,RId9d25a0_3746,
        RIb8860a8_36,RIb832228_204,RId9cd0c8_3747,RIb886120_35,RIb8322a0_203,RId9c86b8_3748,RIb886198_34,RIb832318_202,RIda940a0_3749,RIb886210_33,
        RIb832390_201,RIda91850_3750,RIb886288_32,RIb832408_200,RIda8dbd8_3751,RIb886300_31,RIb832480_199,RIda8a7d0_3752,RIb886378_30,RIb8324f8_198,
        RIda86978_3753,RIb8863f0_29,RIb832570_197,RIda835e8_3754,RIb886468_28,RIb8383a8_196,RIda80f00_3755,RIb8864e0_27,RIb838420_195,RIda7daf8_3756,
        RIb886558_26,RIb838498_194,RIda7a7e0_3757,RIb8865d0_25,RIb838510_193,RIda745e8_3758,RIb886648_24,RIb838588_192,RIda6e018_3759,RIb8866c0_23,
        RIb838600_191,RIda65e40_3760,RIb886738_22,RIb838678_190,RIda5f888_3761,RIb8867b0_21,RIb8386f0_189,RIda59780_3762,RIb886828_20,RIb838768_188,
        RIda510f8_3763,RIb8868a0_19,RIb8387e0_187,RIda4aff0_3764,RIb886918_18,RIb838858_186,RId927408_3765,RIb886990_17,RIb8388d0_185,RId943680_3766,
        RIb886a08_16,RIb838948_184,RId96ccd8_3767,RIb886a80_15,RIb8389c0_183,RId988b30_3768,RIb886af8_14,RIb838a38_182,RId90bb68_3769,RIb886b70_13,
        RIb838ab0_181,RId8f7438_3770,RIb886be8_12,RIb838b28_180,RId8d6dc8_3771,RIb886c60_11,RIb838ba0_179,RId6c4d70_3772,RIb886cd8_10,RIb838c18_178,
        RId6ae7c8_3773,RIb886d50_9,RIb838c90_177,RId835578_3774,RIb886dc8_8,RIb838d08_176,RId8a9d50_3775,RIb886e40_7,RIb838d80_175,RId862aa0_3776,
        RIb886eb8_6,RIb838df8_174,RId99e778_3777,RId9ac620_3778,RId9b8290_3779,RId9bdfd8_3780,RId90fe70_3781,RId918b10_3782,RIda42698_3783,RIda33a58_3784,
        RIda28b08_3785,RIda18aa0_3786,RIda0b288_3787,RId9f8d18_3788,RId9ec9a0_3789,RId9e3418_3790,RIdb156a0_3791,RIdb17f68_3792,RIdb1b640_3793,RIdb1df08_3794,
        RIdb215e0_3795,RIdb23ea8_3796,RIdb26c20_3797,RIdb29e48_3798,RIdb2cbc0_3799,RIdb2fde8_3800,RIdb32b60_3801,RIdb35d88_3802,RIdb38b00_3803,RIdb3b3c8_3804,
        RIdb3eaa0_3805,RIdb404e0_3806,RIdb422e0_3807,RIdb43ac8_3808,RIdb45850_3809,RIdb47128_3810,RIdb483e8_3811,RIdb49888_3812,RIdb4abc0_3813,RIdb4c330_3814,
        RIdb4d410_3815,RIdb4e5e0_3816,RIdb4fa08_3817,RIdb51100_3818,RIdb52c30_3819,RIdb541c0_3820,RIdb559a8_3821,RIdb56e48_3822,RIdb58900_3823,RIdb5a070_3824,
        RIdb5b588_3825,RIdb5d0b8_3826,RIdb5e3f0_3827,RIda95720_3828,RIda97598_3829,RIda99a28_3830,RIda9bd50_3831,RIda9df10_3832,RIda9f4a0_3833,RIdaa1228_3834,
        RIdaa2d58_3835,RIdaa4a68_3836,RIdaa6b38_3837,RIdaa89b0_3838,RIdbdf030_3839,RIdbdcd80_3840,RIdbdaff8_3841,RIdbd9540_3842,RIdbd6e58_3843,RIdbd4860_3844,
        RIdbd25b0_3845,RIdbd0030_3846,RIdbcdc18_3847,RIdbcb800_3848,RIdbc9730_3849,RIdbc7a20_3850,RIdbc5e78_3851,RIdbc40f0_3852,RIdbc1f30_3853,RIdbbf938_3854,
        RIdbbd4a8_3855,RIdbba910_3856,RIdbb8480_3857,RIdbb58e8_3858,RIdbb2648_3859,RIdbb0758_3860,RIdbad788_3861,RIdbaad58_3862,RIdba7d88_3863,RIdba55b0_3864,
        RIdba2ce8_3865,RIdb9fe80_3866,RIdb9d4c8_3867,RIdb9acf0_3868,RIdb98c20_3869,RIdb96178_3870,RIdb93ce8_3871,RIdb916f0_3872,RIdb8e2e8_3873,RIdb8b840_3874,
        RIdb890e0_3875,RIdb86cc8_3876,RIdb84ec8_3877,RIdb83410_3878,RIdb81700_3879,RIdb7fa68_3880,RIdb7db78_3881,RIdb7bb98_3882,RIdb79e10_3883,RIdb78268_3884,
        RIdb76828_3885,RIdb746e0_3886,RIdda9490_3887,RIdda9c88_3888,RIddaa480_3889,RIddaac78_3890,RIddab470_3891,RIddabc68_3892,RIddac460_3893,RIddacc58_3894,
        RIddad450_3895,RIddadc48_3896,RIddae440_3897,RIddaec38_3898,RIddaf430_3899,RIddafc28_3900,RIddb0420_3901,RIddb0c18_3902,RIddb1410_3903,RIddb1c08_3904,
        RIddb2400_3905,RIddb2bf8_3906,RIddb33f0_3907,RIddb3be8_3908,RIddb43e0_3909,RIddb4bd8_3910,RIddb53d0_3911,RIddb5bc8_3912,RIddb63c0_3913,RIddb6bb8_3914,
        RIddb73b0_3915,RIddb7ba8_3916,RIddb83a0_3917,RIddb8b98_3918,RIddb9390_3919,RIddb9b88_3920,RIddba380_3921,RIddbab78_3922,RIddbb370_3923,RIddbbb68_3924,
        RIddbc360_3925,RIddbcb58_3926,RIddbd350_3927,RIddbdb48_3928,RIddbe340_3929,RIddbeb38_3930,RIddbf330_3931,RIddbfb28_3932,RIddc0320_3933,RIddc0b18_3934,
        RIddc1310_3935,RIddc1b08_3936,RIddc2300_3937,RIddc2af8_3938,RIddc32f0_3939,RIddc3ae8_3940,RIddc42e0_3941,RIddc4ad8_3942,RIddc52d0_3943,RIddc5ac8_3944,
        RIddc62c0_3945,RIddc6ab8_3946,RIddc72b0_3947,RIddc7aa8_3948,RIddc82a0_3949,RIddc8a98_3950,RIddc9290_3951,RIddc9a88_3952,RIddca280_3953,RIddcaa78_3954,
        RIddcb270_3955,RIddcba68_3956,RIddcc260_3957,RIddcca58_3958,RIddcd250_3959,RIddcda48_3960,RIddce240_3961,RIddcea38_3962,RIddcf230_3963,RIddcfa28_3964,
        RIddd0220_3965,RIddd0a18_3966,RIddd1210_3967,RIddd1a08_3968,RIdc0fbb8_3681,RIb86fc68_77,RIdc0f0f0_3682,RIb86fce0_76,RIdc0e5b0_3683,RIb86fd58_75,
        RIdc0dae8_3684,RIb87e8a8_74,RIdc0cfa8_3685,RIb87e920_73,RIdc0c3f0_3686,RIb87e998_72,RIdc0b7c0_3687,RIb87ea10_71,RIdc0ac08_3688,RIb87ea88_70,
        RIdc09f60_3689,RIdc093a8_3690,RIdc08700_3691,RIdc07878_3692,RIdc06270_3693,RIdc05118_3694,RIdc03b10_3695,RIdc029b8_3696,RIdc013b0_3697,RIdc00258_3698,
        RIdbff100_3699,RIdbfdaf8_3700,RIdbfc9a0_3701,RIdbfb398_3702,RIdbfa240_3703,RIdbf8c38_3704,RIdbf7ae0_3705,RIdbf6988_3706,RIdbf5380_3707,RIdbf4228_3708,
        RIdbf2c20_3709,RIdbf1ac8_3710,RIdbf04c0_3711,RIdbef368_3712,RIb79b428_272,RIe5efc28_6741,RIe527288_6346,RIe45e528_5951,RIe395df8_5556,RIe1ca840_5161,
        RIe100460_4766,RIe036f80_4371,RIde6b9c8_3976,RIdda31a8_3581,RIdbd9c48_3186,RIdb0e968_2791,RIda3bc30_2396,RId987e10_2001,RId8bc950_1606,RId7f4028_1211,
        RId72b4a8_816,RIe5d6d40_6768,RIe5117a8_6369,RIe444fb0_5975,RIe37f9b8_5584,RIe1ac2a0_5191,RIe0e8ec8_4791,RIe022a30_4393,RIdd8ba30_3609,RIdbc4870_3212,
        RIdaf5f30_2820,RIda25c28_2423,RId96d278_2032,RId8aa728_1632,RId7dcb80_1235,RId710748_846,RIe3ac2b0_6083,RIe3aaca8_6084,RIe3a9b50_6085,RIe3a8548_6086,
        RIe3a73f0_6087,RIe3a6298_6088,RIe3a4c90_6089,RIe3a3b38_6090,RIe3a2530_6091,RIe3a13d8_6092,RIe39fdd0_6093,RIe39ec78_6094,RIe39db20_6095,RIe39c518_6096,
        RIe1694d8_6097,RIe16e398_6098,RIe173270_6099,RIe178388_6100,RIe17c780_6101,RIe1805d8_6102,RIe1877c0_6103,RIe18c9c8_6104,RIe192ff8_6105,RIe198cc8_6106,
        RIe1a05b8_6107,RIe1a6300_6108,RIe1ac318_6109,RIe1b2420_6110,RIe1b7970_6111,RIe1bce48_6112,RIe1c12b8_6113,RIe1c7960_6114,RIe1cc820_6115,RIe1d0fd8_6116,
        RIe094940_6117,RIe090368_6118,RIe08b700_6119,RIe087a10_6120,RIe14c9f0_6121,RIe1495e8_6122,RIe146348_6123,RIe143210_6124,RIe140a38_6125,RIe13d4c8_6126,
        RIe13a660_6127,RIe137168_6128,RIe133a18_6129,RIe12fda0_6130,RIe1280f0_6131,RIe121b38_6132,RIe1194b0_6133,RIe1133a8_6134,RIe10ad20_6135,RIdfd70d0_6136,
        RIdff52b0_6137,RIe01ea70_6138,RIe03a5e0_6139,RIdfb6cb8_6140,RIdfa46d0_6141,RIdf7c7e8_6142,RIdc22218_6143,RIda953d8_6144,RIddeaf80_6145,RIde58a80_6146,
        RIe03fa40_6147,RIe04e338_6148,RIe0629f0_6149,RIe06c608_6150,RIe0732e0_6151,RIe07d0d8_6152,RIe084158_6153,RIdfc61e0_6154,RIe106838_6155,RIe0f8198_6156,
        RIe0eed00_6157,RIe0e2b68_6158,RIe0d0b98_6159,RIe0c3998_6160,RIe0b0960_6161,RIe0a6988_6162,RIe099440_6163,RIe1d3c60_6164,RIe1d69d8_6165,RIe1d9c00_6166,
        RIe1dc978_6167,RIe1dfba0_6168,RIe1e2918_6169,RIe1e5b40_6170,RIe1e88b8_6171,RIe1eb180_6172,RIe1ee858_6173,RIe1f1120_6174,RIe1f47f8_6175,RIe1f70c0_6176,
        RIe1fa180_6177,RIe1fbad0_6178,RIe1fd330_6179,RIe1ff568_6180,RIe2012f0_6181,RIe203000_6182,RIe203f00_6183,RIe2053a0_6184,RIe2066d8_6185,RIe207920_6186,
        RIe208be0_6187,RIe209d38_6188,RIe20b958_6189,RIe20cf60_6190,RIe20e4f0_6191,RIe20f5d0_6192,RIe211178_6193,RIe212c30_6194,RIe214148_6195,RIe215c00_6196,
        RIe217460_6197,RIe218798_6198,RIe2199e0_6199,RIe14e868_6200,RIe151130_6201,RIe153020_6202,RIe154ad8_6203,RIe156518_6204,RIe158228_6205,RIe15a280_6206,
        RIe15c3c8_6207,RIe15ef60_6208,RIe1616c0_6209,RIe164168_6210,RIe166c10_6211,RIe39a100_6212,RIe3984e0_6213,RIe3967d0_6214,RIe3941d8_6215,RIe391c58_6216,
        RIe38f5e8_6217,RIe38d428_6218,RIe38ae30_6219,RIe389030_6220,RIe386fd8_6221,RIe384ff8_6222,RIe3832e8_6223,RIe381218_6224,RIe37f148_6225,RIe37ce20_6226,
        RIe37aeb8_6227,RIe378668_6228,RIe3755a8_6229,RIe372c68_6230,RIe2703f8_6231,RIe26d4a0_6232,RIe26aae8_6233,RIe2686d0_6234,RIe265ca0_6235,RIe264170_6236,
        RIe2616c8_6237,RIe25f238_6238,RIe25c6a0_6239,RIe259ec8_6240,RIe257240_6241,RIe254018_6242,RIe251408_6243,RIe24e8e8_6244,RIe24c110_6245,RIe248d08_6246,
        RIe246170_6247,RIe2435d8_6248,RIe2418c8_6249,RIe23fb40_6250,RIe23dcc8_6251,RIe23ba18_6252,RIe239948_6253,RIe2381d8_6254,RIe236720_6255,RIe2346c8_6256,
        RIe232a30_6257,RIe230bb8_6258,RIe465cb0_6259,RIe4664a8_6260,RIe466ca0_6261,RIe467498_6262,RIe467c90_6263,RIe468488_6264,RIe468c80_6265,RIe469478_6266,
        RIe469c70_6267,RIe46a468_6268,RIe46ac60_6269,RIe46b458_6270,RIe46bc50_6271,RIe46c448_6272,RIe46cc40_6273,RIe46d438_6274,RIe46dc30_6275,RIe46e428_6276,
        RIe46ec20_6277,RIe46f418_6278,RIe46fc10_6279,RIe470408_6280,RIe470c00_6281,RIe4713f8_6282,RIe471bf0_6283,RIe4723e8_6284,RIe472bf8_6285,RIe4733f0_6286,
        RIe473be8_6287,RIe4743e0_6288,RIe474bd8_6289,RIe4753d0_6290,RIe475bc8_6291,RIe4763c0_6292,RIe476bb8_6293,RIe4773b0_6294,RIe477ba8_6295,RIe4783a0_6296,
        RIe478b98_6297,RIe479390_6298,RIe479b88_6299,RIe47a380_6300,RIe47ab78_6301,RIe47b370_6302,RIe47bb68_6303,RIe47c360_6304,RIe47cb58_6305,RIe47d350_6306,
        RIe47db48_6307,RIe47e340_6308,RIe47eb38_6309,RIe47f330_6310,RIe47fb28_6311,RIe480320_6312,RIe480b18_6313,RIe481310_6314,RIe481b08_6315,RIe482300_6316,
        RIe482af8_6317,RIe4832f0_6318,RIe483ae8_6319,RIe4842e0_6320,RIe484ad8_6321,RIe4852d0_6322,RIe485ac8_6323,RIe4862c0_6324,RIe486ab8_6325,RIe4872b0_6326,
        RIe487aa8_6327,RIe4882a0_6328,RIe488a98_6329,RIe489290_6330,RIe489a88_6331,RIe48a280_6332,RIe48aa78_6333,RIe48b270_6334,RIe48ba68_6335,RIe48c260_6336,
        RIe48ca58_6337,RIe48d250_6338,RIe3cd190_6051,RIe3cc3f8_6052,RIe3cb750_6053,RIe3ca9b8_6054,RIe3c9e00_6055,RIe3c9248_6056,RIe3c8708_6057,RIe3c7bc8_6058,
        RIe3c7100_6059,RIe3c6638_6060,RIe3c5af8_6061,RIe3c4ec8_6062,RIe3c4130_6063,RIe3c31b8_6064,RIe3c1bb0_6065,RIe3c0a58_6066,RIe3bf900_6067,RIe3be2f8_6068,
        RIe3bd1a0_6069,RIe3bbb98_6070,RIe3baa40_6071,RIe3b9438_6072,RIe3b82e0_6073,RIe3b7188_6074,RIe3b5b80_6075,RIe3b4a28_6076,RIe3b3420_6077,RIe3b22c8_6078,
        RIe3b0cc0_6079,RIe3afb68_6080,RIe3aea10_6081,RIe3ad408_6082,RIe51b690_6365,RIe500d68_6388,RIe501998_6387,RIe5026b8_6386,RIe5032e8_6385,RIe503f90_6384,
        RIe504d28_6383,RIe505958_6382,RIe50ef58_6371,RIe50ac50_6376,RIe50b880_6375,RIe50c690_6374,RIe50d428_6373,RIe523688_6352,RIe524060_6351,RIe524948_6350,
        RIe51c158_6364,RIe51cc20_6363,RIe51d5f8_6362,RIe5267c0_6347,RIe525d70_6348,RIe525410_6349,RIe51f290_6359,RIe51e840_6360,RIe51dee0_6361,RIe1e2210_5688,
        RIe1e10b8_5689,RIe1dfab0_5690,RIe1de958_5691,RIe1dd350_5692,RIe1dc1f8_5693,RIe1dabf0_5694,RIe1d9a98_5695,RIe1d8940_5696,RIe1d7338_5697,RIe1d61e0_5698,
        RIe1d4bd8_5699,RIe1d3a80_5700,RIe1d2478_5701,RIe099530_5702,RIe09d298_5703,RIe0a2338_5704,RIe0a6fa0_5705,RIe0ac310_5706,RIe0b16f8_5707,RIe0b9240_5708,
        RIe0bf438_5709,RIe0c4730_5710,RIe0cb0a8_5711,RIe0d0df0_5712,RIe0d8aa0_5713,RIe0de608_5714,RIe0e5ca0_5715,RIe0eb358_5716,RIe0ef138_5717,RIe0f3bc0_5718,
        RIe0f8300_5719,RIe0ff380_5720,RIe103430_5721,RIdfce868_5722,RIdfc9fc0_5723,RIdfc6000_5724,RIdfc1410_5725,RIdfbcc58_5726,RIe082f10_5727,RIe0800a8_5728,
        RIe07bd28_5729,RIe078ec0_5730,RIe075ab8_5731,RIe071f18_5732,RIe06f308_5733,RIe06b0f0_5734,RIe067928_5735,RIe0608a8_5736,RIe05a2f0_5737,RIe0541e8_5738,
        RIe04bb60_5739,RIe045a58_5740,RIe03d3d0_5741,RIde1d908_5742,RIde4a200_5743,RIde62e18_5744,RIdc30d68_5745,RIdde3e10_5746,RIddce948_5747,RIdb96b50_5748,
        RIda0b300_5749,RIdc00960_5750,RIdb708e8_5751,RIdc692d0_5752,RIdf7e930_5753,RIdf8d6d8_5754,RIdf9f978_5755,RIdfa6f20_5756,RIdfaf968_5757,RIdfb74b0_5758,
        RIddf5a98_5759,RIde028d8_5760,RIe036620_5761,RIe027530_5762,RIe01deb8_5763,RIe00b3a8_5764,RIdffd938_5765,RIdfefb08_5766,RIdfe0838_5767,RIdfd6680_5768,
        RIe1084d0_5769,RIe10ad98_5770,RIe10e470_5771,RIe110d38_5772,RIe113ab0_5773,RIe116cd8_5774,RIe119a50_5775,RIe11cc78_5776,RIe11f9f0_5777,RIe122c18_5778,
        RIe125990_5779,RIe128258_5780,RIe12b930_5781,RIe12e1f8_5782,RIe1308e0_5783,RIe132398_5784,RIe134300_5785,RIe135ae8_5786,RIe137258_5787,RIe138608_5788,
        RIe139850_5789,RIe13ab88_5790,RIe13c028_5791,RIe13d5b8_5792,RIe13ead0_5793,RIe13fef8_5794,RIe141230_5795,RIe142568_5796,RIe1434e0_5797,RIe144638_5798,
        RIe145880_5799,RIe146ac8_5800,RIe1486e8_5801,RIe149f48_5802,RIe14b550_5803,RIe14c978_5804,RIe14e430_5805,RIe0865e8_5806,RIe087f38_5807,RIe089db0_5808,
        RIe08b7f0_5809,RIe08d578_5810,RIe08f120_5811,RIe091100_5812,RIe093248_5813,RIe0950c0_5814,RIe096998_5815,RIe0986a8_5816,RIe1cfd18_5817,RIe1ce080_5818,
        RIe1cc550_5819,RIe1ca048_5820,RIe1c78e8_5821,RIe1c4f30_5822,RIe1c26e0_5823,RIe1c0b38_5824,RIe1be9f0_5825,RIe1bcce0_5826,RIe1baf58_5827,RIe1b9158_5828,
        RIe1b6908_5829,RIe1b3b90_5830,RIe1b1d18_5831,RIe1aff90_5832,RIe1ae2f8_5833,RIe1ab940_5834,RIe1a8628_5835,RIe1a6030_5836,RIe1a2d90_5837,RIe1a0540_5838,
        RIe19da20_5839,RIe19a870_5840,RIe197cd8_5841,RIe195410_5842,RIe192e90_5843,RIe190460_5844,RIe18e0c0_5845,RIe18bc30_5846,RIe189098_5847,RIe186c08_5848,
        RIe1839e0_5849,RIe1817a8_5850,RIe17fb88_5851,RIe17def0_5852,RIe17c3c0_5853,RIe17a458_5854,RIe1781a8_5855,RIe176240_5856,RIe174530_5857,RIe172988_5858,
        RIe16fc70_5859,RIe16e140_5860,RIe16c1d8_5861,RIe16a5b8_5862,RIe168a88_5863,RIe167138_5864,RIe39c680_5865,RIe39ce78_5866,RIe39d670_5867,RIe39de68_5868,
        RIe39e660_5869,RIe39ee58_5870,RIe39f650_5871,RIe39fe48_5872,RIe3a0640_5873,RIe3a0e38_5874,RIe3a1630_5875,RIe3a1e28_5876,RIe3a2620_5877,RIe3a2e18_5878,
        RIe3a3610_5879,RIe3a3e08_5880,RIe3a4600_5881,RIe3a4df8_5882,RIe3a55f0_5883,RIe3a5de8_5884,RIe3a65e0_5885,RIe3a6dd8_5886,RIe3a75d0_5887,RIe3a7dc8_5888,
        RIe3a85c0_5889,RIe3a8db8_5890,RIe3a95b0_5891,RIe3a9da8_5892,RIe3aa5a0_5893,RIe3aad98_5894,RIe3ab590_5895,RIe3abd88_5896,RIe3ac580_5897,RIe3acd78_5898,
        RIe3ad570_5899,RIe3add68_5900,RIe3ae560_5901,RIe3aed58_5902,RIe3af550_5903,RIe3afd48_5904,RIe3b0540_5905,RIe3b0d38_5906,RIe3b1530_5907,RIe3b1d28_5908,
        RIe3b2520_5909,RIe3b2d18_5910,RIe3b3510_5911,RIe3b3d08_5912,RIe3b4500_5913,RIe3b4cf8_5914,RIe3b54f0_5915,RIe3b5ce8_5916,RIe3b64e0_5917,RIe3b6cd8_5918,
        RIe3b74d0_5919,RIe3b7cc8_5920,RIe3b84c0_5921,RIe3b8cb8_5922,RIe3b94b0_5923,RIe3b9ca8_5924,RIe3ba4a0_5925,RIe3bac98_5926,RIe3bb490_5927,RIe3bbc88_5928,
        RIe3bc480_5929,RIe3bcc78_5930,RIe3bd470_5931,RIe3bdc68_5932,RIe3be460_5933,RIe3bec58_5934,RIe3bf450_5935,RIe3bfc48_5936,RIe3c0440_5937,RIe3c0c38_5938,
        RIe3c1430_5939,RIe3c1c28_5940,RIe3c2420_5941,RIe3c2c18_5942,RIe3c3410_5943,RIe202f10_5656,RIe202448_5657,RIe201980_5658,RIe200e40_5659,RIe2000a8_5660,
        RIe1ff310_5661,RIe1fe668_5662,RIe1fd9c0_5663,RIe1fce80_5664,RIe1fc340_5665,RIe1fb878_5666,RIe1facc0_5667,RIe1fa090_5668,RIe1f9118_5669,RIe1f7fc0_5670,
        RIe1f69b8_5671,RIe1f5860_5672,RIe1f4258_5673,RIe1f3100_5674,RIe1f1fa8_5675,RIe1f09a0_5676,RIe1ef848_5677,RIe1ee240_5678,RIe1ed0e8_5679,RIe1ebae0_5680,
        RIe1ea988_5681,RIe1e9830_5682,RIe1e8228_5683,RIe1e70d0_5684,RIe1e5ac8_5685,RIe1e4970_5686,RIe1e3368_5687,RIe4520c0_5970,RIe438440_5990,RIe4390e8_5989,
        RIe439f70_5988,RIe43ad80_5987,RIe43ba28_5986,RIe43c7c0_5985,RIe43d5d0_5984,RIe445e38_5974,RIe441c98_5979,RIe4429b8_5978,RIe443750_5977,RIe437630_5991,
        RIe45a478_5957,RIe45aec8_5956,RIe45b8a0_5955,RIe452b88_5969,RIe4534e8_5968,RIe453fb0_5967,RIe45d880_5952,RIe45cdb8_5953,RIe45c278_5954,RIe455e28_5964,
        RIe4554c8_5965,RIe454988_5966,RIe116b70_5293,RIe115a18_5294,RIe114410_5295,RIe1132b8_5296,RIe111cb0_5297,RIe110b58_5298,RIe10f550_5299,RIe10e3f8_5300,
        RIe10d2a0_5301,RIe10bc98_5302,RIe10ab40_5303,RIe109538_5304,RIe1083e0_5305,RIe106dd8_5306,RIdfd3728_5307,RIdfd71c0_5308,RIdfdc8f0_5309,RIdfe0b80_5310,
        RIdfe6760_5311,RIdfeb788_5312,RIdff1f98_5313,RIdff7f38_5314,RIdffe400_5315,RIe005750_5316,RIe00b420_5317,RIe0132b0_5318,RIe0193b8_5319,RIe0202d0_5320,
        RIe023de0_5321,RIe027878_5322,RIe02ccd8_5323,RIe0322a0_5324,RIe038768_5325,RIe03c728_5326,RIde01258_5327,RIddfd748_5328,RIddf9788_5329,RIddf3d88_5330,
        RIdfba228_5331,RIdfb5e30_5332,RIdfb2aa0_5333,RIdfaec48_5334,RIdfabf48_5335,RIdfa97e8_5336,RIdfa5e40_5337,RIdfa2f60_5338,RIdf9e4d8_5339,RIdf99618_5340,
        RIdf90f90_5341,RIdf8ae88_5342,RIdf848d0_5343,RIdf7c248_5344,RIdf76140_5345,RIdc56298_5346,RIdd75f50_5347,RIdd9d6b8_5348,RIdb67180_5349,RIdc198c0_5350,
        RIdc008e8_5351,RIdacdc88_5352,RId8fd180_5353,RIdb353b0_5354,RIdbdbca0_5355,RIdb8b8b8_5356,RIddb1a28_5357,RIddc60e0_5358,RIddd3cb8_5359,RIdddeaa0_5360,
        RIdde50d0_5361,RIddeee50_5362,RIdc2bb60_5363,RIdc34788_5364,RIde6e7b8_5365,RIde62ad0_5366,RIde55510_5367,RIde4a188_5368,RIde36d90_5369,RIde29c80_5370,
        RIde1c210_5371,RIde0cb08_5372,RIe03d4c0_5373,RIe040b98_5374,RIe043460_5375,RIe046b38_5376,RIe049400_5377,RIe04c178_5378,RIe04f3a0_5379,RIe052118_5380,
        RIe055340_5381,RIe0580b8_5382,RIe05b2e0_5383,RIe05e058_5384,RIe060920_5385,RIe063ff8_5386,RIe0662a8_5387,RIe068288_5388,RIe069a70_5389,RIe06b870_5390,
        RIe06cf68_5391,RIe06e6d8_5392,RIe06fa10_5393,RIe070eb0_5394,RIe0721e8_5395,RIe073808_5396,RIe074960_5397,RIe0762b0_5398,RIe0779a8_5399,RIe079118_5400,
        RIe07a798_5401,RIe07bcb0_5402,RIe07d768_5403,RIe07f220_5404,RIe080cd8_5405,RIe082088_5406,RIe083078_5407,RIe0843b0_5408,RIdfbbbf0_5409,RIdfbd5b8_5410,
        RIdfbf3b8_5411,RIdfc15f0_5412,RIdfc30a8_5413,RIdfc4f20_5414,RIdfc6f00_5415,RIdfc85f8_5416,RIdfca3f8_5417,RIdfcc720_5418,RIdfce8e0_5419,RIe106478_5420,
        RIe104948_5421,RIe102b48_5422,RIe100f28_5423,RIe0fea20_5424,RIe0fcd10_5425,RIe0fa3d0_5426,RIe0f7838_5427,RIe0f5a38_5428,RIe0f3968_5429,RIe0f1b68_5430,
        RIe0f0290_5431,RIe0ee508_5432,RIe0ec690_5433,RIe0eaea8_5434,RIe0e8658_5435,RIe0e54a8_5436,RIe0e2988_5437,RIe0e0228_5438,RIe0dd7f8_5439,RIe0da828_5440,
        RIe0d7f60_5441,RIe0d4f18_5442,RIe0d3280_5443,RIe0d02b0_5444,RIe0cdad8_5445,RIe0cae50_5446,RIe0c8150_5447,RIe0c5d38_5448,RIe0c3290_5449,RIe0c0d88_5450,
        RIe0be628_5451,RIe0bbdd8_5452,RIe0b91c8_5453,RIe0b5f28_5454,RIe0b3318_5455,RIe0b02d0_5456,RIe0adeb8_5457,RIe0ac0b8_5458,RIe0aa330_5459,RIe0a83c8_5460,
        RIe0a6a00_5461,RIe0a40c0_5462,RIe0a2158_5463,RIe0a0010_5464,RIe09e378_5465,RIe09c668_5466,RIe09a8e0_5467,RIe099080_5468,RIe1d1cf8_5469,RIe1d24f0_5470,
        RIe1d2ce8_5471,RIe1d34e0_5472,RIe1d3cd8_5473,RIe1d44d0_5474,RIe1d4cc8_5475,RIe1d54c0_5476,RIe1d5cb8_5477,RIe1d64b0_5478,RIe1d6ca8_5479,RIe1d74a0_5480,
        RIe1d7c98_5481,RIe1d8490_5482,RIe1d8c88_5483,RIe1d9480_5484,RIe1d9c78_5485,RIe1da470_5486,RIe1dac68_5487,RIe1db460_5488,RIe1dbc58_5489,RIe1dc450_5490,
        RIe1dcc48_5491,RIe1dd440_5492,RIe1ddc38_5493,RIe1de430_5494,RIe1dec28_5495,RIe1df420_5496,RIe1dfc18_5497,RIe1e0410_5498,RIe1e0c08_5499,RIe1e1400_5500,
        RIe1e1bf8_5501,RIe1e23f0_5502,RIe1e2be8_5503,RIe1e33e0_5504,RIe1e3bd8_5505,RIe1e43d0_5506,RIe1e4bc8_5507,RIe1e53c0_5508,RIe1e5bb8_5509,RIe1e63b0_5510,
        RIe1e6ba8_5511,RIe1e73a0_5512,RIe1e7b98_5513,RIe1e8390_5514,RIe1e8b88_5515,RIe1e9380_5516,RIe1e9b78_5517,RIe1ea370_5518,RIe1eab68_5519,RIe1eb360_5520,
        RIe1ebb58_5521,RIe1ec350_5522,RIe1ecb48_5523,RIe1ed340_5524,RIe1edb38_5525,RIe1ee330_5526,RIe1eeb28_5527,RIe1ef320_5528,RIe1efb18_5529,RIe1f0310_5530,
        RIe1f0b08_5531,RIe1f1300_5532,RIe1f1af8_5533,RIe1f22f0_5534,RIe1f2ae8_5535,RIe1f32e0_5536,RIe1f3ad8_5537,RIe1f42d0_5538,RIe1f4ac8_5539,RIe1f52c0_5540,
        RIe1f5ab8_5541,RIe1f62b0_5542,RIe1f6aa8_5543,RIe1f72a0_5544,RIe1f7a98_5545,RIe1f8290_5546,RIe1f8a88_5547,RIe1f9280_5548,RIe137870_5261,RIe136da8_5262,
        RIe136358_5263,RIe135890_5264,RIe134d50_5265,RIe134288_5266,RIe1337c0_5267,RIe132c08_5268,RIe131fd8_5269,RIe1313a8_5270,RIe1307f0_5271,RIe12fbc0_5272,
        RIe12f080_5273,RIe12da78_5274,RIe12c920_5275,RIe12b318_5276,RIe12a1c0_5277,RIe128bb8_5278,RIe127a60_5279,RIe126908_5280,RIe125300_5281,RIe1241a8_5282,
        RIe122ba0_5283,RIe121a48_5284,RIe120440_5285,RIe11f2e8_5286,RIe11e190_5287,RIe11cb88_5288,RIe11ba30_5289,RIe11a428_5290,RIe1192d0_5291,RIe117cc8_5292,
        RIe38a110_5575,RIe378410_5590,RIe379220_5589,RIe379e50_5588,RIe26f4f8_5601,RIe270290_5600,RIe270ec0_5599,RIe271be0_5598,RIe37b908_5586,RIe375008_5594,
        RIe375da0_5593,RIe376a48_5592,RIe377768_5591,RIe3921f8_5562,RIe392b58_5561,RIe3934b8_5560,RIe38a908_5574,RIe38b1f0_5573,RIe38b9e8_5572,RIe3951c8_5557,
        RIe394868_5558,RIe393e90_5559,RIe38da40_5569,RIe38cf78_5570,RIe38c4b0_5571,RIe04cad8_4898,RIe04b980_4899,RIe04a378_4900,RIe049220_4901,RIe047c18_4902,
        RIe046ac0_4903,RIe045968_4904,RIe044360_4905,RIe043208_4906,RIe041c00_4907,RIe040aa8_4908,RIe03f4a0_4909,RIe03e348_4910,RIe03d1f0_4911,RIde08bc0_4912,
        RIde0d030_4913,RIde131b0_4914,RIde17968_4915,RIde1f528_4916,RIde24e38_4917,RIde29ed8_4918,RIde31390_4919,RIde36e08_4920,RIde3efe0_4921,RIde45070_4922,
        RIde4c9d8_4923,RIde51b68_4924,RIde553a8_4925,RIde59c50_4926,RIde5e390_4927,RIde65668_4928,RIde6a4b0_4929,RIde6f820_4930,RIdf73710_4931,RIdc38040_4932,
        RIdc32b68_4933,RIdc2ee78_4934,RIdc29bf8_4935,RIddf1628_4936,RIddee388_4937,RIddeaa58_4938,RIdde7a88_4939,RIdde35a0_4940,RIdde0cd8_4941,RIddddf60_4942,
        RIdddb710_4943,RIddd5e78_4944,RIddd2278_4945,RIddcc080_4946,RIddc39f8_4947,RIddbd8f0_4948,RIddb5268_4949,RIddaf160_4950,RIdb7c228_4951,RIdb96c40_4952,
        RIdbbbd38_4953,RIdbdcdf8_4954,RIdb5db80_4955,RIdb48190_4956,RIdb26ba8_4957,RId917aa8_4958,RId986da8_4959,RIda7eb60_4960,RIdaf90e0_4961,RIdab27a8_4962,
        RIdbf1ca8_4963,RIdc00a50_4964,RIdc0fe88_4965,RIdc16080_4966,RIdc1c098_4967,RIdc25080_4968,RIdb67810_4969,RIdda8518_4970,RIdd9d5c8_4971,RIdd8f270_4972,
        RIdd82fe8_4973,RIdd74150_4974,RIdc641b8_4975,RIdc54600_4976,RIdc46848_4977,RIdc3b970_4978,RIdf77220_4979,RIdf79f98_4980,RIdf7c860_4981,RIdf7ff38_4982,
        RIdf82800_4983,RIdf85ed8_4984,RIdf887a0_4985,RIdf8be78_4986,RIdf8e740_4987,RIdf91008_4988,RIdf946e0_4989,RIdf96fa8_4990,RIdf9a680_4991,RIdf9ccf0_4992,
        RIdf9ec58_4993,RIdfa04b8_4994,RIdfa1bb0_4995,RIdfa3b18_4996,RIdfa4dd8_4997,RIdfa6110_4998,RIdfa75b0_4999,RIdfa88e8_5000,RIdfa9d10_5001,RIdfab048_5002,
        RIdfac218_5003,RIdfad460_5004,RIdfaecc0_5005,RIdfb0610_5006,RIdfb1c90_5007,RIdfb3310_5008,RIdfb4828_5009,RIdfb5d40_5010,RIdfb77f8_5011,RIdfb92b0_5012,
        RIdfba9a8_5013,RIddf2ca8_5014,RIddf4580_5015,RIddf6308_5016,RIddf8270_5017,RIddf9e90_5018,RIddfbdf8_5019,RIddfdb08_5020,RIddff548_5021,RIde015a0_5022,
        RIde03508_5023,RIde04fc0_5024,RIe03bbe8_5025,RIe039cf8_5026,RIe038600_5027,RIe0363c8_5028,RIe033b78_5029,RIe031580_5030,RIe02ee98_5031,RIe02c4e0_5032,
        RIe02a488_5033,RIe028958_5034,RIe026b58_5035,RIe025460_5036,RIe023b88_5037,RIe021fe0_5038,RIe020168_5039,RIe01dcd8_5040,RIe01b758_5041,RIe018440_5042,
        RIe0157b8_5043,RIe012590_5044,RIe010628_5045,RIe00d298_5046,RIe00a778_5047,RIe007e38_5048,RIe004df0_5049,RIe0024b0_5050,RIdfff558_5051,RIdffcd08_5052,
        RIdffa260_5053,RIdff7b78_5054,RIdff4f68_5055,RIdff1ea8_5056,R_25610_96cc360,R_25642_95f0d48,R_25644_9598060,R_25646_95984f8,R_25614_953c348,R_25616_96251f8,
        R_25618_96ed6b0,R_2561a_95f00d0,R_2561c_95f0418,R_2561e_95f0760,R_25620_953c3f0,R_25622_953c690,R_25612_953c9d8,R_25624_95f08b0,R_25626_953ca80,R_25628_96253f0,
        R_2562a_9632be8,R_253fc_9d20ef0,R_25412_9530108,R_25428_95f75a0,R_2543e_95301b0,R_25454_95304f8,R_2546a_9533198,R_25474_95332e8,R_25476_96dee60,R_25478_95f7798,
        R_2547a_96def08,R_253fe_95f7990,R_25400_9d21190,R_25402_9d21388,R_25404_9589e90,R_25406_9d21430,R_25408_9533780,R_2540a_9533b70,R_2540c_9d216d0,R_2540e_958a5c8,
        R_25410_96defb0,R_25414_9d21778,R_25416_9d21cb8,R_25418_95f7ae0,R_2541a_9d21d60,R_2541c_96df100,R_2541e_9d221f8,R_25420_958ac58,R_25422_95f7b88,R_25424_9533c18,
        R_25426_958b630,R_2542a_9d222a0,R_2542c_9533d68,R_2542e_95f7c30,R_25430_9d22498,R_25432_9d22540,R_25434_9533f60,R_25436_96df1a8,R_25438_95f7f78,R_2543a_9534008,
        R_2543c_9534200,R_25440_95f80c8,R_25442_96df250,R_25444_9d22690,R_25446_95fa438,R_25448_95fa4e0,R_2544a_958bcc0,R_2544c_9d22738,R_2544e_9d227e0,R_25450_9d22888,
        R_25452_9d22930,R_25456_9d229d8,R_25458_95fa588,R_2545a_9534350,R_2545c_95fa828,R_2545e_9d22a80,R_25460_96df2f8,R_25462_96df3a0,R_25464_95343f8,R_25466_95fa8d0,
        R_25468_95faac8,R_2546c_958bd68,R_2546e_958be10,R_25470_95fab70,R_25472_9d22b28,R_2547c_958beb8,R_25492_9d22bd0,R_254a8_958bf60,R_254be_9d22c78,R_254d4_9d22dc8,
        R_254ea_9d22e70,R_254f4_958c0b0,R_254f6_9d22f18,R_254f8_958c158,R_254fa_9d22fc0,R_2547e_958c200,R_25480_9d23068,R_25482_9d231b8,R_25484_958c2a8,R_25486_958c350,
        R_25488_9d23458,R_2548a_958c4a0,R_2548c_9d235a8,R_2548e_9d236f8,R_25490_958c548,R_25494_958c5f0,R_25496_9d237a0,R_25498_958c698,R_2549a_958f728,R_2549c_9d23848,
        R_2549e_958f7d0,R_254a0_958f878,R_254a2_9d23998,R_254a4_9d23ae8,R_254a6_9d23c38,R_254aa_9d23d88,R_254ac_9d23e30,R_254ae_9d23f80,R_254b0_9d24028,R_254b2_9d240d0,
        R_254b4_9d24220,R_254b6_9d242c8,R_254b8_9590988,R_254ba_9590a30,R_254bc_9590cd0,R_254c0_9d24418,R_254c2_9590d78,R_254c4_9590f70,R_254c6_9591178,R_254c8_9d24568,
        R_254ca_9d24bf8,R_254cc_9d25090,R_254ce_95916b8,R_254d0_9591808,R_254d2_9d251e0,R_254d6_9d25f10,R_254d8_9d25fb8,R_254da_95918b0,R_254dc_9d265a0,R_254de_9591958,
        R_254e0_9d26990,R_254e2_9d26c30,R_254e4_9591a00,R_254e6_95347e8,R_254e8_9591b50,R_254ec_9591bf8,R_254ee_9d26d80,R_254f0_9d27368,R_254f2_9d27410,R_254fc_96df4f0,
        R_25512_9d276b0,R_25528_96df598,R_2553e_9534890,R_25554_9d27c98,R_2556a_96df640,R_25574_9d27de8,R_25576_96df6e8,R_25578_9534bd8,R_2557a_96df838,R_254fe_96dfad8,
        R_25500_9534d28,R_25502_9534dd0,R_25504_9534f20,R_25506_9d281d8,R_25508_96dfb80,R_2550a_9d28328,R_2550c_9d283d0,R_2550e_96dfc28,R_25510_9534fc8,R_25514_96dfcd0,
        R_25516_9d28520,R_25518_96dfe20,R_2551a_96dfec8,R_2551c_9535070,R_2551e_95351c0,R_25520_9535268,R_25522_96dff70,R_25524_96e0018,R_25526_96e00c0,R_2552a_9535310,
        R_2552c_96e0168,R_2552e_96e0210,R_25530_96e02b8,R_25532_96e0408,R_25534_96e0558,R_25536_96e0600,R_25538_9535658,R_2553a_9d289b8,R_2553c_96e06a8,R_25540_95358f8,
        R_25542_96e0750,R_25544_96e0b40,R_25546_96e0be8,R_25548_96e0c90,R_2554a_96e0d38,R_2554c_95359a0,R_2554e_9d28a60,R_25550_96e0e88,R_25552_9535a48,R_25556_96e0f30,
        R_25558_9535b98,R_2555a_9d28c58,R_2555c_96e0fd8,R_2555e_9d28d00,R_25560_9535c40,R_25562_95362d0,R_25564_9536810,R_25566_9536a08,R_25568_96e1080,R_2556c_96e1128,
        R_2556e_9d28ef8,R_25570_96e11d0,R_25572_96e1c50,R_2557c_9591d48,R_25592_9591df0,R_255a8_96e2e08,R_255be_9591e98,R_255d4_9591f40,R_255ea_96e3690,R_255f4_96e6918,
        R_255f6_96e69c0,R_255f8_9d29048,R_255fa_9d28718,R_2557e_9591fe8,R_25580_96e6fa8,R_25582_96e72f0,R_25584_9d287c0,R_25586_9592090,R_25588_9592138,R_2558a_96e7398,
        R_2558c_9d28868,R_2558e_9d290f0,R_25590_9d29240,R_25594_96e7cc8,R_25596_95921e0,R_25598_9592288,R_2559a_9592330,R_2559c_96e82b0,R_2559e_9d292e8,R_255a0_9d2dfb0,
        R_255a2_9592528,R_255a4_9592678,R_255a6_9d2e058,R_255aa_96e8358,R_255ac_9592918,R_255ae_96e86a0,R_255b0_9d2e988,R_255b2_9d29390,R_255b4_9d2ec28,R_255b6_9d294e0,
        R_255b8_9d2f360,R_255ba_9592a68,R_255bc_9592b10,R_255c0_9d30128,R_255c2_9592c60,R_255c4_96e8940,R_255c6_96e89e8,R_255c8_9d30278,R_255ca_96e8be0,R_255cc_9592f00,
        R_255ce_9d29588,R_255d0_9d296d8,R_255d2_9d30518,R_255d6_9d29828,R_255d8_96e9120,R_255da_96e93c0,R_255dc_96e9510,R_255de_9d307b8,R_255e0_9d29cc0,R_255e2_9592fa8,
        R_255e4_9593050,R_255e6_96e9858,R_255e8_96e9a50,R_255ec_95930f8,R_255ee_9d29eb8,R_255f0_96ea038,R_255f2_95931a0,R_253bc_96eacb0,R_253be_9593248,R_253c0_9d29f60,
        R_253c2_95932f0,R_253c4_96eae00,R_253c6_9536b58,R_253c8_9593398,R_253ca_9d2a350,R_253cc_b7dc210,R_253ce_b7dcd38,R_253d0_b7dcde0,R_253d2_9593590,R_253d4_96376b8,
        R_253d6_9d2a4a0,R_253d8_9596038,R_253da_b7dc2b8,R_253dc_96eb0a0,R_253de_9596578,R_253e0_9536f48,R_253e2_96eb298,R_253e4_9537098,R_253e6_96eb340,R_253e8_95373e0,
        R_253ea_9596a10,R_253ec_9d30860,R_253ee_9ef0090,R_253f0_9d30f98,R_253f2_9ef05d0,R_253f4_9d31040,R_253f6_9d31238,R_253f8_9d314d8,R_253fa_9d316d0,R_25666_96346d0,
        R_1a4_b821b50,R_1a3_b821aa8,R_23ca4_96329f0,R_23cba_9f596e0,R_23cd0_962b7c0,R_23ce6_955f268,R_23cfc_9f5c4d0,R_23d12_9d225e8,R_23d1c_962b910,R_23d1e_95a3470,
        R_23d20_9632c90,R_23d22_95a3710,R_23ca6_9ee76c0,R_23ca8_9ee7810,R_23caa_9ee78b8,R_23cac_9ee8140,R_23cae_962bbb0,R_23cb0_9ee8920,R_23cb2_9d22d20,R_23cb4_9ee8bc0,
        R_23cb6_9632d38,R_23cb8_9d23110,R_23cbc_962bc58,R_23cbe_9ee9ad8,R_23cc0_9d23260,R_23cc2_9632f30,R_23cc4_9eec430,R_23cc6_9d23308,R_23cc8_9eef4c0,R_23cca_9eefca0,
        R_23ccc_9d23650,R_23cce_9ef0678,R_23cd2_95a3908,R_23cd4_962bd00,R_23cd6_9632fd8,R_23cd8_962be50,R_23cda_96331d0,R_23cdc_962bef8,R_23cde_9d30ef0,R_23ce0_9d238f0,
        R_23ce2_9d23b90,R_23ce4_962bfa0,R_23ce8_962c048,R_23cea_95a3a58,R_23cec_9d23ed8,R_23cee_9ef09c0,R_23cf0_9ef4380,R_23cf2_95a3ba8,R_23cf4_9ef4a10,R_23cf6_962c0f0,
        R_23cf8_96c3060,R_23cfa_96c6d68,R_23cfe_9d310e8,R_23d00_96c72a8,R_23d02_962c390,R_23d04_96c74a0,R_23d06_962da88,R_23d08_9d24178,R_23d0a_962df20,R_23d0c_9633278,
        R_23d0e_9633320,R_23d10_95a3e48,R_23d14_95a4040,R_23d16_9d24370,R_23d18_96c7e78,R_23d1a_96333c8,R_23d24_9633470,R_23d3a_9633518,R_23d50_962dfc8,R_23d66_9629b88,
        R_23d7c_95547c8,R_23d92_96335c0,R_23d9c_96337b8,R_23d9e_9633908,R_23da0_9633a58,R_23da2_962e7a8,R_23d26_9554870,R_23d28_962a560,R_23d2a_962ee38,R_23d2c_962a8a8,
        R_23d2e_962f2d0,R_23d30_95549c0,R_23d32_9633cf8,R_23d34_962f4c8,R_23d36_9633da0,R_23d38_9633e48,R_23d3c_9633ef0,R_23d3e_962c4e0,R_23d40_9554bb8,R_23d42_9554d08,
        R_23d44_9634040,R_23d46_962f6c0,R_23d48_9554f00,R_23d4a_962c8d0,R_23d4c_9635000,R_23d4e_962fab0,R_23d52_95552f0,R_23d54_96350a8,R_23d56_96351f8,R_23d58_962fc00,
        R_23d5a_95554e8,R_23d5c_9555638,R_23d5e_9635540,R_23d60_96355e8,R_23d62_9635738,R_23d64_96359d8,R_23d68_962ca20,R_23d6a_9635f18,R_23d6c_962ff48,R_23d6e_9636068,
        R_23d70_96363b0,R_23d72_9636ae8,R_23d74_9637220,R_23d76_9637e98,R_23d78_9638b10,R_23d7a_962d4a0,R_23d7e_96305d8,R_23d80_9638bb8,R_23d82_9638fa8,R_23d84_962d548,
        R_23d86_9639398,R_23d88_95556e0,R_23d8a_9639440,R_23d8c_9d18d00,R_23d8e_9d19d68,R_23d90_9630a70,R_23d94_9d1a008,R_23d96_9d1a350,R_23d98_9d1a9e0,R_23d9a_96314f0,
        R_23da4_9634430,R_23dba_95558d8,R_23dd0_9555a28,R_23de6_9d1ac80,R_23dfc_962d9e0,R_23e12_9555b78,R_23e1c_96344d8,R_23e1e_9555e18,R_23e20_9d1b070,R_23e22_9d1b8f8,
        R_23da6_9634a18,R_23da8_9555f68,R_23daa_9635150,R_23dac_96352a0,R_23dae_9556010,R_23db0_9557078,R_23db2_96353f0,R_23db4_9d1ba48,R_23db6_962db30,R_23db8_96357e0,
        R_23dbc_9559730,R_23dbe_955bde8,R_23dc0_955dd68,R_23dc2_9d1baf0,R_23dc4_955e158,R_23dc6_9638db0,R_23dc8_9d1bb98,R_23dca_9639248,R_23dcc_9d1bce8,R_23dce_96c81c0,
        R_23dd2_955e4a0,R_23dd4_955ea88,R_23dd6_96392f0,R_23dd8_9d15d18,R_23dda_955ee78,R_23ddc_9d168e8,R_23dde_9d16ae0,R_23de0_962e310,R_23de2_9d16c30,R_23de4_9d16e28,
        R_23de8_9d170c8,R_23dea_955f1c0,R_23dec_96c87a8,R_23dee_955f310,R_23df0_9d1bee0,R_23df2_955f3b8,R_23df4_95a39b0,R_23df6_96c8af0,R_23df8_95a3b00,R_23dfa_95a40e8,
        R_23dfe_95a44d8,R_23e00_9d1bf88,R_23e02_95a4580,R_23e04_95a4c10,R_23e06_9d17218,R_23e08_95a5348,R_23e0a_962ec40,R_23e0c_9d17608,R_23e0e_95a57e0,R_23e10_95a5930,
        R_23e14_9d18910,R_23e16_9d19630,R_23e18_95a5c78,R_23e1a_95a6260,R_23e24_9d1c030,R_23e3a_95a4628,R_23e50_95a48c8,R_23e66_95a4b68,R_23e7c_95b1438,R_23e92_9d19780,
        R_23e9c_95a6d88,R_23e9e_95b1780,R_23ea0_95a7028,R_23ea2_95a70d0,R_23e26_95b1828,R_23e28_95a7220,R_23e2a_95b2bd8,R_23e2c_95b3310,R_23e2e_95818b0,R_23e30_9582138,
        R_23e32_9582288,R_23e34_95a7760,R_23e36_9582870,R_23e38_95a78b0,R_23e3c_9d1c0d8,R_23e3e_9582a68,R_23e40_9d1b118,R_23e42_9582e58,R_23e44_9582f00,R_23e46_95830f8,
        R_23e48_958cbd8,R_23e4a_958cc80,R_23e4c_95a7aa8,R_23e4e_958f5d8,R_23e52_958f920,R_23e54_9590058,R_23e56_95a7bf8,R_23e58_95a7ca0,R_23e5a_95901a8,R_23e5c_959fdb8,
        R_23e5e_95a0b80,R_23e60_9d1c4c8,R_23e62_9625b28,R_23e64_96261b8,R_23e68_9d1b268,R_23e6a_9d1c570,R_23e6c_95a7d48,R_23e6e_9626458,R_23e70_95a8090,R_23e72_9628330,
        R_23e74_9628480,R_23e76_9628528,R_23e78_95a8138,R_23e7a_96285d0,R_23e7e_9628720,R_23e80_9628bb8,R_23e82_962c198,R_23e84_9d1c618,R_23e86_95a8288,R_23e88_9634238,
        R_23e8a_9d1c6c0,R_23e8c_96342e0,R_23e8e_9634970,R_23e90_9d1c8b8,R_23e94_9639830,R_23e96_9d159d0,R_23e98_9d15e68,R_23e9a_95a83d8,R_23c64_96c9a08,R_23c66_9d1b658,
        R_23c68_96ca920,R_23c6a_9d244c0,R_23c6c_96cb4f0,R_23c6e_9d1b700,R_23c70_9d1ca08,R_23c72_96cb640,R_23c74_962f030,R_23c76_9d1cc00,R_23c78_9d1cd50,R_23c7a_9d1cdf8,
        R_23c7c_9d1b7a8,R_23c7e_9d1cf48,R_23c80_9d1d098,R_23c82_9d1d1e8,R_23c84_95a8528,R_23c86_9d1b9a0,R_23c88_95a8720,R_23c8a_9d1be38,R_23c8c_9d246b8,R_23c8e_96cb838,
        R_23c90_9d24760,R_23c92_9d1c2d0,R_23c94_9d1d3e0,R_23c96_95a87c8,R_23c98_9d19438,R_23c9a_9d1c378,R_23c9c_9d1c768,R_23c9e_9d1d488,R_23ca0_9d1c960,R_23ca2_9d1e8e0,
        R_23ebc_9667ae0,R_23ebe_965f6f8,R_23ec0_9667b88,R_23ec2_96688a8,R_23ec4_95ac230,R_23ec6_95ac428,R_23ec8_966a780,R_23eca_966a8d0,R_23eba_965f8f0,R_23ecc_95ac620,
        R_23ece_95ac770,R_23ed0_966a978,R_23ed2_966aa20,R_23eb8_966aac8,R_23eea_95b1588,R_23eec_9d1e448,R_23eee_9d1e790,R_23a0c_95b1630,R_23a22_95b1c18,R_23a38_966acc0,
        R_23a4e_95b1d68,R_23a64_966ad68,R_23a7a_95b2c80,R_23a84_9661a68,R_23a86_9d1d7d0,R_23a88_966ae10,R_23a8a_966b0b0,R_23a0e_962f420,R_23a10_966ba88,R_23a12_95b2fc8,
        R_23a14_9d1f6a8,R_23a16_952daf8,R_23a18_95b3268,R_23a1a_9581220,R_23a1c_9d1d878,R_23a1e_9663160,R_23a20_9d1e250,R_23a24_9d1fb40,R_23a26_95305a0,R_23a28_95812c8,
        R_23a2a_9530798,R_23a2c_95816b8,R_23a2e_9663550,R_23a30_9531e90,R_23a32_9531f38,R_23a34_9532130,R_23a36_9532280,R_23a3a_9532328,R_23a3c_9581760,R_23a3e_9581f40,
        R_23a40_95323d0,R_23a42_9532868,R_23a44_9582720,R_23a46_9532b08,R_23a48_9532c58,R_23a4a_9582918,R_23a4c_966a4e0,R_23a50_9532e50,R_23a52_9d24808,R_23a54_9533390,
        R_23a56_9d20668,R_23a58_9582db0,R_23a5a_9583050,R_23a5c_9533978,R_23a5e_9534158,R_23a60_9d20710,R_23a62_95349e0,R_23a66_9537290,R_23a68_9d1f750,R_23a6a_966a6d8,
        R_23a6c_966aeb8,R_23a6e_966b158,R_23a70_9537a70,R_23a72_9539f30,R_23a74_95831a0,R_23a76_9537c68,R_23a78_9d20a58,R_23a7c_9537d10,R_23a7e_9537e60,R_23a80_9538250,
        R_23a82_95382f8,R_23a8c_9d21e08,R_23aa2_9583440,R_23ab8_9d1f8a0,R_23ace_9d1ff30,R_23ae4_9d23ce0,R_23afa_95834e8,R_23b04_9583590,R_23b06_9d20860,R_23b08_9d24958,
        R_23b0a_9d24ca0,R_23a8e_95836e0,R_23a90_9583e18,R_23a92_9d25288,R_23a94_9d20908,R_23a96_9d25330,R_23a98_9d22348,R_23a9a_9d253d8,R_23a9c_9d233b0,R_23a9e_9d25528,
        R_23aa0_9d255d0,R_23aa4_9d23500,R_23aa6_9d25678,R_23aa8_9d23a40,R_23aaa_9d24610,R_23aac_9d25880,R_23aae_9d248b0,R_23ab0_9d26258,R_23ab2_9584898,R_23ab4_9d24a00,
        R_23ab6_9d26450,R_23aba_9d26648,R_23abc_9d26e28,R_23abe_9d270c8,R_23ac0_9584c88,R_23ac2_9d24aa8,R_23ac4_9d24d48,R_23ac6_9585270,R_23ac8_9585708,R_23aca_9d27bf0,
        R_23acc_9d28910,R_23ad0_9d29198,R_23ad2_9d29630,R_23ad4_9d24fe8,R_23ad6_95857b0,R_23ad8_9d2a0b0,R_23ada_9585900,R_23adc_9d2a200,R_23ade_9d2a3f8,R_23ae0_9d2a7e8,
        R_23ae2_9d25138,R_23ae6_9d2ad28,R_23ae8_95860e0,R_23aea_9d25480,R_23aec_9d25928,R_23aee_9d25bc8,R_23af0_95864d0,R_23af2_9d25e68,R_23af4_95866c8,R_23af6_9586770,
        R_23af8_9587688,R_23afc_9d26ed0,R_23afe_9587730,R_23b00_9d27aa0,R_23b02_9d2add0,R_23b0c_95877d8,R_23b22_95386e8,R_23b38_95388e0,R_23b4e_9588108,R_23b64_9538ad8,
        R_23b7a_9d2b118,R_23b84_95881b0,R_23b86_95899f8,R_23b88_9589aa0,R_23b8a_9d2b460,R_23b0e_958d268,R_23b10_95390c0,R_23b12_9539168,R_23b14_95394b0,R_23b16_95399f0,
        R_23b18_9539c90,R_23b1a_953ba18,R_23b1c_953bac0,R_23b1e_958d460,R_23b20_9d2b508,R_23b24_953bf58,R_23b26_953c0a8,R_23b28_953c1f8,R_23b2a_953c540,R_23b2c_9d2b5b0,
        R_23b2e_953c888,R_23b30_953cdc8,R_23b32_958da48,R_23b34_9d2b700,R_23b36_953cf18,R_23b3a_958de38,R_23b3c_958e180,R_23b3e_96ddca8,R_23b40_96dddf8,R_23b42_958e570,
        R_23b44_958e810,R_23b46_96de098,R_23b48_9d285c8,R_23b4a_96de3e0,R_23b4c_9d28b08,R_23b50_96de530,R_23b52_958ef48,R_23b54_9d24b50,R_23b56_9d25d18,R_23b58_958ff08,
        R_23b5a_96e6c60,R_23b5c_96e8160,R_23b5e_96ebc70,R_23b60_95903a0,R_23b62_95906e8,R_23b66_96ebdc0,R_23b68_95efb90,R_23b6a_9596d58,R_23b6c_9d2b7a8,R_23b6e_9598c30,
        R_23b70_95f0220,R_23b72_9598cd8,R_23b74_95f1918,R_23b76_9599170,R_23b78_9d28bb0,R_23b7c_95f37f0,R_23b7e_95f41c8,R_23b80_95f4318,R_23b82_95992c0,R_23b8c_9599608,
        R_23ba2_9599758,R_23bb8_9599800,R_23bce_9599950,R_23be4_962f570,R_23bfa_9599b48,R_23c04_959a088,R_23c06_959a130,R_23c08_959a1d8,R_23c0a_962f618,R_23b8e_959a5c8,
        R_23b90_959a9b8,R_23b92_959ac58,R_23b94_959aef8,R_23b96_962f8b8,R_23b98_959afa0,R_23b9a_959b048,R_23b9c_959b0f0,R_23b9e_959b198,R_23ba0_959b240,R_23ba4_959b6d8,
        R_23ba6_959b828,R_23ba8_959b8d0,R_23baa_959ba20,R_23bac_9d28da8,R_23bae_959bac8,R_23bb0_959d268,R_23bb2_959d508,R_23bb4_959dce8,R_23bb6_959e420,R_23bba_9d28fa0,
        R_23bbc_962f960,R_23bbe_9d298d0,R_23bc0_959e618,R_23bc2_959eea0,R_23bc4_959f098,R_23bc6_9d29978,R_23bc8_9d25dc0,R_23bca_959f9c8,R_23bcc_9d29a20,R_23bd0_95a0e20,
        R_23bd2_9d29b70,R_23bd4_962fb58,R_23bd6_95a0f70,R_23bd8_9d29c18,R_23bda_9619ae0,R_23bdc_9619b88,R_23bde_9619d80,R_23be0_9619e28,R_23be2_961a020,R_23be6_961a0c8,
        R_23be8_961a218,R_23bea_961a4b8,R_23bec_961a800,R_23bee_961a8a8,R_23bf0_961a950,R_23bf2_961ad40,R_23bf4_961ade8,R_23bf6_961ae90,R_23bf8_961af38,R_23bfc_9d26060,
        R_23bfe_961b088,R_23c00_9d29d68,R_23c02_961b1d8,R_239cc_95f4af8,R_239ce_962fd50,R_239d0_9558e00,R_239d2_9d261b0,R_239d4_95f52d8,R_239d6_9558ea8,R_239d8_961b670,
        R_239da_95f5620,R_239dc_961b910,R_239de_9d2b850,R_239e0_9d2b9a0,R_239e2_9d29e10,R_239e4_9d2a158,R_239e6_961bb08,R_239e8_961c978,R_239ea_961cd68,R_239ec_9d2baf0,
        R_239ee_95f5968,R_239f0_95f5ab8,R_239f2_9d2a2a8,R_239f4_961ce10,R_239f6_9634e08,R_239f8_9d2bb98,R_239fa_9d2bd90,R_239fc_962fdf8,R_239fe_962fea0,R_23a00_961d200,
        R_23a02_961d5f0,R_23a04_961d698,R_23a06_962fff0,R_23a08_961d740,R_23a0a_961d938,R_23c24_9d2a698,R_23c26_9d2c420,R_23c28_962ac98,R_23c2a_9d2c4c8,R_23c2c_9d2c570,
        R_23c2e_95f63e8,R_23c30_9d2a890,R_23c32_962ad40,R_23c22_9d2aa88,R_23c34_9d2c810,R_23c36_9d2ab30,R_23c38_9d2c8b8,R_23c3a_9d2cab0,R_23c20_9635e70,R_23c52_962b868,
        R_23c54_9d2af20,R_23c56_9d2b310,R_23774_9630098,R_2378a_962b9b8,R_237a0_9d2cd50,R_237b6_962bb08,R_237cc_9d2cff0,R_237e2_9d2d098,R_237ec_9d2d140,R_237ee_9d2d290,
        R_237f0_962c240,R_237f2_9559688,R_23776_96301e8,R_23778_9d2d7d0,R_2377a_962c2e8,R_2377c_9d2d878,R_2377e_962ce10,R_23780_9d2d920,R_23782_962d938,R_23784_962e5b0,
        R_23786_9d2d9c8,R_23788_9d2dc68,R_2378c_9d2dd10,R_2378e_9d2ddb8,R_23790_9d2e100,R_23792_9d2e1a8,R_23794_9d2f0c0,R_23796_9630290,R_23798_96303e0,R_2379a_9d2f210,
        R_2379c_9d2f7f8,R_2379e_9630728,R_237a2_96307d0,R_237a4_9d2fb40,R_237a6_9d301d0,R_237a8_9559bc8,R_237aa_9630140,R_237ac_96312f8,R_237ae_9d30710,R_237b0_9630b18,
        R_237b2_9630c68,R_237b4_9d309b0,R_237b8_9630d10,R_237ba_9630fb0,R_237bc_9631100,R_237be_9d30a58,R_237c0_9d30da0,R_237c2_96311a8,R_237c4_96313a0,R_237c6_96318e0,
        R_237c8_9631a30,R_237ca_9d30e48,R_237ce_9d31190,R_237d0_9631b80,R_237d2_9d31f58,R_237d4_9631448,R_237d6_9631790,R_237d8_9d323f0,R_237da_9631ad8,R_237dc_9d32540,
        R_237de_9632018,R_237e0_9631cd0,R_237e4_9632210,R_237e6_9d32690,R_237e8_96322b8,R_237ea_9d32888,R_237f4_9631e20,R_2380a_9d329d8,R_23820_9d32a80,R_23836_9d32f18,
        R_2384c_9d2b3b8,R_23862_9631ec8,R_2386c_9632360,R_2386e_9632a98,R_23870_9d32fc0,R_23872_9632408,R_237f6_9632600,R_237f8_9d33500,R_237fa_96326a8,R_237fc_9d33650,
        R_237fe_9d336f8,R_23800_9d33a40,R_23802_9632750,R_23804_96328a0,R_23806_9d340d0,R_23808_9632948,R_2380c_9d2b658,R_2380e_9d34418,R_23810_9d34760,R_23812_9d34fe8,
        R_23814_9632de0,R_23816_9632e88,R_23818_9d35720,R_2381a_9d2bc40,R_2381c_b805670,R_2381e_b805868,R_23822_9633080,R_23824_b8060f0,R_23826_9633128,R_23828_9633b00,
        R_2382a_9632b40,R_2382c_9634190,R_2382e_9638720,R_23830_9d2c180,R_23832_96389c0,R_23834_9638a68,R_23838_9d15880,R_2383a_b806198,R_2383c_9d2c768,R_2383e_9d16a38,
        R_23840_9d2ca08,R_23842_b806240,R_23844_9d17170,R_23846_9d17c98,R_23848_b8062e8,R_2384a_b806390,R_2384e_9d2cca8,R_23850_9d17fe0,R_23852_9d18328,R_23854_9d2d1e8,
        R_23856_9d1fd38,R_23858_b8064e0,R_2385a_9d2d3e0,R_2385c_9d220a8,R_2385e_9535d90,R_23860_b806588,R_23864_9d25720,R_23866_b8066d8,R_23868_b806780,R_2386a_9d2d530,
        R_23874_95f7840,R_2388a_95f7e28,R_238a0_9d28e50,R_238b6_95f8170,R_238cc_95fcd90,R_238e2_95fda08,R_238ec_95fdb58,R_238ee_95fdca8,R_238f0_95fdd50,R_238f2_9d2d728,
        R_23876_95ff6e8,R_23878_9535e38,R_2387a_9633668,R_2387c_9f4ddd0,R_2387e_9f51b80,R_23880_9f51e20,R_23882_9d29ac8,R_23884_9f53278,R_23886_9f53320,R_23888_9f54580,
        R_2388c_9f54778,R_2388e_9d2dbc0,R_23890_9d2e250,R_23892_9f548c8,R_23894_9f54970,R_23896_9f54c10,R_23898_9f55348,R_2389a_9f55498,R_2389c_9d2a740,R_2389e_9d2e3a0,
        R_238a2_9d2b070,R_238a4_9633710,R_238a6_9f55b28,R_238a8_9f56260,R_238aa_9f56500,R_238ac_9f5baf8,R_238ae_9ee9d78,R_238b0_9d2ba48,R_238b2_9d2bce8,R_238b4_9eea0c0,
        R_238b8_9eeb518,R_238ba_9eedf18,R_238bc_9eee6f8,R_238be_9ef2010,R_238c0_9537530,R_238c2_9ef2208,R_238c4_9ef3660,R_238c6_9ef3858,R_238c8_9633860,R_238ca_9ef3a50,
        R_238ce_9ef3af8,R_238d0_9ef3ba0,R_238d2_9ef3c48,R_238d4_9ef4620,R_238d6_9d2c2d0,R_238d8_9ef4770,R_238da_9d2cb58,R_238dc_9ef4ab8,R_238de_9ef4c08,R_238e0_9ef4ff8,
        R_238e4_9ef5148,R_238e6_9ef51f0,R_238e8_9d2cf48,R_238ea_9ef53e8,R_238f4_9d2e4f0,R_2390a_96339b0,R_23920_9633c50,R_23936_9d266f0,R_2394c_9d2e838,R_23962_9d2ecd0,
        R_2396c_9d2ed78,R_2396e_9d2f018,R_23970_9d2f168,R_23972_b8068d0,R_238f6_9d2f2b8,R_238f8_9d2f9f0,R_238fa_9d2fde0,R_238fc_9633f98,R_238fe_b806a20,R_23900_96340e8,
        R_23902_9d30320,R_23904_9634580,R_23906_9d305c0,R_23908_9634b68,R_2390c_9d30ba8,R_2390e_9d30c50,R_23910_b806ac8,R_23912_9d32000,R_23914_b806b70,R_23916_9d320a8,
        R_23918_9634c10,R_2391a_9d32150,R_2391c_9634cb8,R_2391e_9d32498,R_23922_9d32738,R_23924_9d327e0,R_23926_9d32b28,R_23928_9d32bd0,R_2392a_9635348,R_2392c_9635690,
        R_2392e_9d32c78,R_23930_9d32d20,R_23932_9635a80,R_23934_9d32dc8,R_23938_9d331b8,R_2393a_9d2d488,R_2393c_9d333b0,R_2393e_9d335a8,R_23940_9d337a0,R_23942_9635b28,
        R_23944_9d2d5d8,R_23946_9d338f0,R_23948_9635bd0,R_2394a_9d33998,R_2394e_9d33ae8,R_23950_9d33b90,R_23952_9636110,R_23954_9d33ce0,R_23956_b806c18,R_23958_9d33ed8,
        R_2395a_9d33f80,R_2395c_9636308,R_2395e_b806cc0,R_23960_9d34028,R_23964_9d34178,R_23966_9d2db18,R_23968_96365a8,R_2396a_9636848,R_23734_96368f0,R_23736_9636998,
        R_23738_9636a40,R_2373a_b7dc0c0,R_2373c_9636b90,R_2373e_9636c38,R_23740_b7dc168,R_23742_b806d68,R_23744_b806e10,R_23746_9636ed8,R_23748_b806eb8,R_2374a_9637028,
        R_2374c_b806f60,R_2374e_b8070b0,R_23750_9d33308,R_23752_b807158,R_23754_9ef5880,R_23756_9d26798,R_23758_9d342c8,R_2375a_9ef5928,R_2375c_96c2b20,R_2375e_9d31820,
        R_23760_9d31970,R_23762_9637178,R_23764_9d26840,R_23766_96372c8,R_23768_9d268e8,R_2376a_9d26a38,R_2376c_9d26ae0,R_2376e_9637370,R_23770_9d26b88,R_23772_9637418,
        R_2398c_96c2fb8,R_2398e_9559c70,R_23990_96c35a0,R_23992_96e8010,R_23994_955a300,R_23996_955a450,R_23998_9d34ca0,R_2399a_96c3840,R_2398a_9d34d48,R_2399c_96c3a38,
        R_2399e_96c3d80,R_239a0_955a840,R_239a2_96c59b8,R_23988_96eaf50,R_239ba_96ca728,R_239bc_955b8a8,R_239be_b7db6e8,R_234dc_b8085b0,R_234f2_b80b988,R_23508_b808658,
        R_2351e_b808700,R_23534_b8087a8,R_2354a_b8088f8,R_23554_b80ba30,R_23556_b80bb80,R_23558_b80bec8,R_2355a_b80bf70,R_234de_b8089a0,R_234e0_b808a48,R_234e2_b809768,
        R_234e4_b809df8,R_234e6_b80c2b8,R_234e8_b80e040,R_234ea_b80e580,R_234ec_b80c600,R_234ee_b80f0a8,R_234f0_b80fd20,R_234f4_b80c750,R_234f6_b80ffc0,R_234f8_b7ddf98,
        R_234fa_b80c7f8,R_234fc_b7de0e8,R_234fe_b7de388,R_23500_b7de430,R_23502_b80c9f0,R_23504_b7de580,R_23506_b80ca98,R_2350a_b7de820,R_2350c_b7dea18,R_2350e_b7dee08,
        R_23510_b80cc90,R_23512_b80cd38,R_23514_b7df1f8,R_23516_b80ce88,R_23518_b7df348,R_2351a_b7df540,R_2351c_b80cf30,R_23520_b7dfc78,R_23522_b80d080,R_23524_b80d278,
        R_23526_b7dff18,R_23528_b80d320,R_2352a_b7e0068,R_2352c_b80d5c0,R_2352e_b7e01b8,R_23530_b80d668,R_23532_b7e0458,R_23536_b7e05a8,R_23538_b80d7b8,R_2353a_b80de48,
        R_2353c_b7e0998,R_2353e_b7e0b90,R_23540_b7e1178,R_23542_b80e430,R_23544_b80e628,R_23546_b80e778,R_23548_b7e1568,R_2354c_b80e970,R_2354e_b7e16b8,R_23550_b80eb68,
        R_23552_b7e1808,R_2355c_b7e18b0,R_23572_b805c58,R_23588_b7e1958,R_2359e_b80ed60,R_235b4_95ad7d8,R_235ca_b806438,R_235d4_b7e1a00,R_235d6_b80f000,R_235d8_b7e1bf8,
        R_235da_b7e1ca0,R_2355e_b7e1e98,R_23560_95ad9d0,R_23562_b7e1f40,R_23564_95adb20,R_23566_b7e1fe8,R_23568_b80f3f0,R_2356a_b80f5e8,R_2356c_b806630,R_2356e_b7e2090,
        R_23570_b80f690,R_23574_b7e2138,R_23576_b7e21e0,R_23578_b7e23d8,R_2357a_b7e2720,R_2357c_b7e2870,R_2357e_b7e29c0,R_23580_b806828,R_23582_b7e2a68,R_23584_b7e2c60,
        R_23586_b7e2f00,R_2358a_b80f7e0,R_2358c_96cb8e0,R_2358e_b7e2fa8,R_23590_b7e30f8,R_23592_b806978,R_23594_b807008,R_23596_b7e32f0,R_23598_b80fb28,R_2359a_b7e3398,
        R_2359c_b807698,R_235a0_b7e34e8,R_235a2_96cbb80,R_235a4_b80fbd0,R_235a6_96cc018,R_235a8_95adf10,R_235aa_b7e36e0,R_235ac_b807890,R_235ae_b7e3788,R_235b0_b7e38d8,
        R_235b2_b7e3ad0,R_235b6_b7e3cc8,R_235b8_b7e3f68,R_235ba_b807f20,R_235bc_b807fc8,R_235be_b8101b8,R_235c0_b7e40b8,R_235c2_b7e4208,R_235c4_b8105a8,R_235c6_b810650,
        R_235c8_96cc210,R_235cc_b7e42b0,R_235ce_b7e4400,R_235d0_b7e4550,R_235d2_b7e45f8,R_235dc_b8106f8,R_235f2_b7e46a0,R_23608_b808118,R_2361e_b7e47f0,R_23634_b7e49e8,
        R_2364a_b7dd860,R_23654_95ae060,R_23656_b7dd908,R_23658_b7ddda0,R_2365a_b7dde48,R_235de_9637b50,R_235e0_95ae1b0,R_235e2_b7ddef0,R_235e4_b7de238,R_235e6_b7e4b38,
        R_235e8_9637fe8,R_235ea_b7de2e0,R_235ec_b808310,R_235ee_9638138,R_235f0_96381e0,R_235f4_b7e4d30,R_235f6_96383d8,R_235f8_b7de6d0,R_235fa_9638480,R_235fc_b7de8c8,
        R_235fe_9638528,R_23600_96385d0,R_23602_b7de970,R_23604_b7deac0,R_23606_9638678,R_2360a_96387c8);
input RIde67cd8_3982,RIde68638_3981,RIde68f20_3980,RIe5319e0_6884,RIe549ef0_6842,RIe549770_6843,RIe548ff0_6844,RIea91330_6888,RIb79b4a0_271,
        RIb79b518_270,RIe5329d0_6883,RIeb72150_6905,RIb7b9608_246,RIe5c6738_6786,RIe4fc9e8_6393,RIb7b9590_247,RIe5c5bf8_6787,RIe4fbcc8_6394,RIb7b9518_248,
        RIe5c4fc8_6788,RIe4faf30_6395,RIb7b94a0_249,RIe5c4500_6789,RIe4fa198_6396,RIb7b9428_250,RIe5c3948_6790,RIe4f9388_6397,RIb7b93b0_251,RIe5c2e08_6791,
        RIe4f85f0_6398,RIb7af720_252,RIe5c22c8_6792,RIe4f7a38_6399,RIb7af6a8_253,RIe5c1710_6793,RIe4f6ef8_6400,RIb7af630_254,RIe5e09d0_6767,RIe4af828_6445,
        RIb7af5b8_255,RIe5e1330_6766,RIe519818_6368,RIb7af540_256,RIe5e1ba0_6765,RIe4b0200_6444,RIb7af4c8_257,RIe5e2488_6764,RIe51a2e0_6367,RIb7af450_258,
        RIe5e2d70_6763,RIe4bdce8_6441,RIb7af3d8_259,RIe5e3568_6762,RIe51acb8_6366,RIb7a5bf8_260,RIe588848_6840,RIe4bd310_6442,RIb7a0c48_261,RIe5e3e50_6761,
        RIe4b0a70_6443,RIeab80c0_6897,RIe5331c8_6882,RIe5339c0_6881,RIeab87c8_6898,RIe5341b8_6880,RIe5349b0_6879,RIea94af8_6890,RIe5351a8_6878,RIe5359a0_6877,
        RIeab78c8_6895,RIeab7d00_6896,RIeacfa18_6902,RIeab6518_6891,RIeb352c8_6904,RIe4340c0_5995,RIe26ce10_5604,RIe162368_5252,RIe0d89b0_4811,RIe00f6b0_4415,
        RIde415d8_4022,RIdd731d8_3637,RIdba6bb8_3248,RIdad7918_2858,RIda15da0_2441,RId95c8b0_2053,RId88c728_1664,RId7c3590_1267,RId6f73b0_878,RIe4333a0_5996,
        RIe26c000_5605,RIe1658d8_5248,RIe0d7d08_4812,RIe00e918_4416,RIde408b8_4023,RIdc72420_3638,RIdba5e98_3249,RIdad6b80_2859,RIda150f8_2442,RId95bcf8_2054,
        RId88bbe8_1665,RId7c2870_1268,RId6f68e8_879,RIe4326f8_5997,RIe26b2e0_5606,RIe164b40_5249,RIe0d6fe8_4813,RIe00db80_4417,RIde3fb20_4024,RIdc71610_3639,
        RIdba51f0_3250,RIdad5d70_2860,RIda143d8_2443,RId95b1b8_2055,RId88b030_1666,RId7c1b50_1269,RId6f5cb8_880,RIe431ac8_5998,RIe26a7a0_5607,RIe1615d0_5253,
        RIe0d62c8_4814,RIe00ce60_4418,RIde3ed88_4025,RIdc70800_3640,RIdba4548_3251,RIdaebc88_2833,RIda13640_2444,RId95a600_2056,RId88a478_1667,RId7c0e30_1270,
        RId6f5100_881,RIe430e20_5999,RIe269c60_5608,RIe163088_5251,RIe0d55a8_4815,RIe00c0c8_4419,RIde3df00_4026,RIdc6f9f0_3641,RIdba3828_3252,RIdaeb0d0_2834,
        RIda12920_2445,RId959a48_2057,RId889938_1668,RId7c0110_1271,RId6f4638_882,RIe4301f0_6000,RIe269120_5609,RIe160838_5254,RIe0d49f0_4816,RIe00b330_4420,
        RIde3d1e0_4027,RIdc6ed48_3642,RIdbb8138_3227,RIdaea590_2835,RIda11c00_2446,RId958f08_2058,RId888d80_1669,RId7bf4e0_1272,RId6f3a80_883,RIe42f4d0_6001,
        RIe268568_5610,RIe172718_5244,RIe0d3dc0_4817,RIe00a598_4421,RIde3c448_4028,RIdc6e280_3643,RIdbb7328_3228,RIdae97f8_2836,RIda10df0_2447,RId9582d8_2059,
        RId888240_1670,RId7be838_1273,RId7064a0_859,RIe42e8a0_6002,RIe2679b0_5611,RIe163e20_5250,RIe0d2e48_4818,RIe009710_4422,RIde3b728_4029,RIdc6d740_3644,
        RIdbb6518_3229,RIdae8a60_2837,RIda101c0_2448,RId957720_2060,RId89b638_1645,RId7d2338_1248,RId705780_860,RIe3f8a98_6047,RIe385d90_5583,RIe182a68_5243,
        RIe0f3008_4788,RIdfc11b8_4469,RIde5ad30_4003,RIdd93500_3608,RIdbcac48_3211,RIdaff2d8_2817,RIda2b970_2422,RId977f88_2027,RId8ab538_1631,RId7e5f28_1234,
        RId71bad0_843,RIe450d88_5972,RIe386678_5582,RIe1bcc68_5184,RIe088e38_4865,RIdfc07e0_4470,RIde5b618_4002,RIdd93ed8_3607,RIdb62338_3285,RIdaffda0_2816,
        RIda2c258_2421,RId978960_2026,RId8ae508_1629,RId7827c0_1310,RId71c2c8_842,RIe3f8048_6048,RIe386e70_5581,RIe1bd4d8_5183,RIe0af538_4863,RIe02a050_4392,
        RIde5be10_4001,RIdd94928_3606,RIdbcb530_3210,RIdb00bb0_2815,RId9cdfc8_2495,RId9791d0_2025,RId86cf28_1704,RId7e6798_1233,RId71cb38_841,RIe3e5628_6050,
        RIe3876e0_5580,RIe1bdd48_5182,RIe0aeb60_4864,RIe02a8c0_4391,RIde5c6f8_4000,RIdd95288_3605,RIdb8a760_3284,RIdabee68_2890,RIda2cbb8_2420,RId9799c8_2024,
        RId8aed00_1628,RId790848_1309,RId71d330_840,RIe3f9e48_6045,RIe387ed8_5579,RIe183440_5242,RIe0aff10_4862,RIdfcdc38_4468,RIde5cf68_3999,RIdd95b70_3604,
        RIdbcbe18_3209,RIdb01498_2814,RIda2d4a0_2419,RId97a238_2023,RId8af7c8_1627,RId7a41e0_1308,RId71dba0_839,RIe3f7760_6049,RIe3887c0_5578,RIe15c260_5259,
        RIe0f3878_4787,RIdfce700_4467,RIde5d760_3998,RIdd963e0_3603,RIdbcc7f0_3208,RIdb01d80_2813,RIda2def0_2418,RId97ab20_2022,RId8ac078_1630,RId7e6f90_1232,
        RId71e398_838,RIe451670_5971,RIe388fb8_5577,RIe1be5b8_5181,RIe0b0870_4861,RIdfcf2b8_4466,RIde5dfd0_3997,RIdd96cc8_3602,RIdbcd0d8_3207,RIdb02668_2812,
        RIda2e760_2417,RId97b318_2021,RId86c4d8_1705,RId7a4bb8_1307,RId71ec08_837,RIe3f9470_6046,RIe3898a0_5576,RIe15b900_5260,RIe0f4070_4786,RIdfcfc90_4465,
        RIde5e840_3996,RIdd97538_3601,RIdbcd9c0_3206,RIdb02f50_2811,RIda2f0c0_2416,RId97bc00_2020,RId8b0290_1626,RId7e7800_1231,RId71f400_836,RIde5fec0_3994,
        RIde4ec88_4006,RIb7b9680_245,RIb79b338_274,RIde60988_3993,RIde612e8_3992,RIde6ad98_3977,RIde6a2d0_3978,RIde69970_3979,RIde63250_3989,RIde62878_3990,
        RIde61e28_3991,RIea90778_6887,RIe546890_6849,RIe546098_6850,RIe545dc8_6851,RIe545648_6852,RIb839848_152,RIb839668_156,RIb8396e0_155,RIde5f3f8_3995,
        RIb79b3b0_273,RIde4c8e8_4009,RIb7b96f8_244,RIde4d6f8_4008,RIb7c20c8_243,RIde431f8_4020,RIb7c5728_242,RIde43f90_4019,RIb7c57a0_241,RIde44da0_4018,
        RIb7c5818_240,RIde45ac0_4017,RIb7c5890_239,RIde468d0_4016,RIb7c5908_238,RIde4fb10_4005,RIb7a09f0_266,RIde49300_4013,RIb7a0a68_265,RIde4a020_4012,
        RIb7a0ae0_264,RIde4ae30_4011,RIb7a0b58_263,RIde4bb50_4010,RIb7a0bd0_262,RIdbee210_3713,RIb87eb00_69,RIe667bb0_6885,RIe667f70_6886,RIb839b90_145,
        RIb7c5980_237,RIeab7058_6894,RIea91768_6889,RIdbecc08_3714,RIb87eb78_68,RIb7c59f8_236,RIdbebab0_3715,RIb87ebf0_67,RIb7c5a70_235,RIdbea4a8_3716,
        RIb882ca0_66,RIb7cade0_234,RIdbe9350_3717,RIb885310_65,RIb7cae58_233,RIdbe7d48_3718,RIb885388_64,RIb7caed0_232,RIdbe6bf0_3719,RIb885400_63,
        RIb7caf48_231,RIdbe5a98_3720,RIb885478_62,RIb7cafc0_230,RIdbe4490_3721,RIb8854f0_61,RIb7cb038_229,RIdbe3338_3722,RIb885568_60,RIb7cb0b0_228,
        RIdbe1d30_3723,RIb8855e0_59,RIb7cb128_227,RIdbe0bd8_3724,RIb885658_58,RIb7d00d8_226,RIdaab098_3725,RIb8856d0_57,RIb8263d8_225,RIdaaf0d0_3726,
        RIb885748_56,RIb826e28_224,RIdab2fa0_3727,RIb8857c0_55,RIb826ea0_223,RIdab8e50_3728,RIb885838_54,RIb826f18_222,RIdabcf00_3729,RIb8858b0_53,
        RIb826f90_221,RIdac3788_3730,RIb885928_52,RIb8293a8_220,RIdac8eb8_3731,RIb8859a0_51,RIb829420_219,RIdacf650_3732,RIb885a18_50,RIb829498_218,
        RIdad4fd8_3733,RIb885a90_49,RIb829510_217,RIdadaf00_3734,RIb885b08_48,RIb829588_216,RIdae2610_3735,RIb885b80_47,RIb829600_215,RIdae8268_3736,
        RIb885bf8_46,RIb829678_214,RIdaef720_3737,RIb885c70_45,RIb8296f0_213,RIdaf4e50_3738,RIb885ce8_44,RIb82dae8_212,RIdafa508_3739,RIb885d60_43,
        RIb82db60_211,RIdafe630_3740,RIb885dd8_42,RIb82dbd8_210,RIdb03b08_3741,RIb885e50_41,RIb82dc50_209,RIdb09d00_3742,RIb885ec8_40,RIb82dcc8_208,
        RIdb0e440_3743,RIb885f40_39,RIb82dd40_207,RIdb13468_3744,RIb885fb8_38,RIb82ddb8_206,RId9d7370_3745,RIb886030_37,RIb82de30_205,RId9d25a0_3746,
        RIb8860a8_36,RIb832228_204,RId9cd0c8_3747,RIb886120_35,RIb8322a0_203,RId9c86b8_3748,RIb886198_34,RIb832318_202,RIda940a0_3749,RIb886210_33,
        RIb832390_201,RIda91850_3750,RIb886288_32,RIb832408_200,RIda8dbd8_3751,RIb886300_31,RIb832480_199,RIda8a7d0_3752,RIb886378_30,RIb8324f8_198,
        RIda86978_3753,RIb8863f0_29,RIb832570_197,RIda835e8_3754,RIb886468_28,RIb8383a8_196,RIda80f00_3755,RIb8864e0_27,RIb838420_195,RIda7daf8_3756,
        RIb886558_26,RIb838498_194,RIda7a7e0_3757,RIb8865d0_25,RIb838510_193,RIda745e8_3758,RIb886648_24,RIb838588_192,RIda6e018_3759,RIb8866c0_23,
        RIb838600_191,RIda65e40_3760,RIb886738_22,RIb838678_190,RIda5f888_3761,RIb8867b0_21,RIb8386f0_189,RIda59780_3762,RIb886828_20,RIb838768_188,
        RIda510f8_3763,RIb8868a0_19,RIb8387e0_187,RIda4aff0_3764,RIb886918_18,RIb838858_186,RId927408_3765,RIb886990_17,RIb8388d0_185,RId943680_3766,
        RIb886a08_16,RIb838948_184,RId96ccd8_3767,RIb886a80_15,RIb8389c0_183,RId988b30_3768,RIb886af8_14,RIb838a38_182,RId90bb68_3769,RIb886b70_13,
        RIb838ab0_181,RId8f7438_3770,RIb886be8_12,RIb838b28_180,RId8d6dc8_3771,RIb886c60_11,RIb838ba0_179,RId6c4d70_3772,RIb886cd8_10,RIb838c18_178,
        RId6ae7c8_3773,RIb886d50_9,RIb838c90_177,RId835578_3774,RIb886dc8_8,RIb838d08_176,RId8a9d50_3775,RIb886e40_7,RIb838d80_175,RId862aa0_3776,
        RIb886eb8_6,RIb838df8_174,RId99e778_3777,RId9ac620_3778,RId9b8290_3779,RId9bdfd8_3780,RId90fe70_3781,RId918b10_3782,RIda42698_3783,RIda33a58_3784,
        RIda28b08_3785,RIda18aa0_3786,RIda0b288_3787,RId9f8d18_3788,RId9ec9a0_3789,RId9e3418_3790,RIdb156a0_3791,RIdb17f68_3792,RIdb1b640_3793,RIdb1df08_3794,
        RIdb215e0_3795,RIdb23ea8_3796,RIdb26c20_3797,RIdb29e48_3798,RIdb2cbc0_3799,RIdb2fde8_3800,RIdb32b60_3801,RIdb35d88_3802,RIdb38b00_3803,RIdb3b3c8_3804,
        RIdb3eaa0_3805,RIdb404e0_3806,RIdb422e0_3807,RIdb43ac8_3808,RIdb45850_3809,RIdb47128_3810,RIdb483e8_3811,RIdb49888_3812,RIdb4abc0_3813,RIdb4c330_3814,
        RIdb4d410_3815,RIdb4e5e0_3816,RIdb4fa08_3817,RIdb51100_3818,RIdb52c30_3819,RIdb541c0_3820,RIdb559a8_3821,RIdb56e48_3822,RIdb58900_3823,RIdb5a070_3824,
        RIdb5b588_3825,RIdb5d0b8_3826,RIdb5e3f0_3827,RIda95720_3828,RIda97598_3829,RIda99a28_3830,RIda9bd50_3831,RIda9df10_3832,RIda9f4a0_3833,RIdaa1228_3834,
        RIdaa2d58_3835,RIdaa4a68_3836,RIdaa6b38_3837,RIdaa89b0_3838,RIdbdf030_3839,RIdbdcd80_3840,RIdbdaff8_3841,RIdbd9540_3842,RIdbd6e58_3843,RIdbd4860_3844,
        RIdbd25b0_3845,RIdbd0030_3846,RIdbcdc18_3847,RIdbcb800_3848,RIdbc9730_3849,RIdbc7a20_3850,RIdbc5e78_3851,RIdbc40f0_3852,RIdbc1f30_3853,RIdbbf938_3854,
        RIdbbd4a8_3855,RIdbba910_3856,RIdbb8480_3857,RIdbb58e8_3858,RIdbb2648_3859,RIdbb0758_3860,RIdbad788_3861,RIdbaad58_3862,RIdba7d88_3863,RIdba55b0_3864,
        RIdba2ce8_3865,RIdb9fe80_3866,RIdb9d4c8_3867,RIdb9acf0_3868,RIdb98c20_3869,RIdb96178_3870,RIdb93ce8_3871,RIdb916f0_3872,RIdb8e2e8_3873,RIdb8b840_3874,
        RIdb890e0_3875,RIdb86cc8_3876,RIdb84ec8_3877,RIdb83410_3878,RIdb81700_3879,RIdb7fa68_3880,RIdb7db78_3881,RIdb7bb98_3882,RIdb79e10_3883,RIdb78268_3884,
        RIdb76828_3885,RIdb746e0_3886,RIdda9490_3887,RIdda9c88_3888,RIddaa480_3889,RIddaac78_3890,RIddab470_3891,RIddabc68_3892,RIddac460_3893,RIddacc58_3894,
        RIddad450_3895,RIddadc48_3896,RIddae440_3897,RIddaec38_3898,RIddaf430_3899,RIddafc28_3900,RIddb0420_3901,RIddb0c18_3902,RIddb1410_3903,RIddb1c08_3904,
        RIddb2400_3905,RIddb2bf8_3906,RIddb33f0_3907,RIddb3be8_3908,RIddb43e0_3909,RIddb4bd8_3910,RIddb53d0_3911,RIddb5bc8_3912,RIddb63c0_3913,RIddb6bb8_3914,
        RIddb73b0_3915,RIddb7ba8_3916,RIddb83a0_3917,RIddb8b98_3918,RIddb9390_3919,RIddb9b88_3920,RIddba380_3921,RIddbab78_3922,RIddbb370_3923,RIddbbb68_3924,
        RIddbc360_3925,RIddbcb58_3926,RIddbd350_3927,RIddbdb48_3928,RIddbe340_3929,RIddbeb38_3930,RIddbf330_3931,RIddbfb28_3932,RIddc0320_3933,RIddc0b18_3934,
        RIddc1310_3935,RIddc1b08_3936,RIddc2300_3937,RIddc2af8_3938,RIddc32f0_3939,RIddc3ae8_3940,RIddc42e0_3941,RIddc4ad8_3942,RIddc52d0_3943,RIddc5ac8_3944,
        RIddc62c0_3945,RIddc6ab8_3946,RIddc72b0_3947,RIddc7aa8_3948,RIddc82a0_3949,RIddc8a98_3950,RIddc9290_3951,RIddc9a88_3952,RIddca280_3953,RIddcaa78_3954,
        RIddcb270_3955,RIddcba68_3956,RIddcc260_3957,RIddcca58_3958,RIddcd250_3959,RIddcda48_3960,RIddce240_3961,RIddcea38_3962,RIddcf230_3963,RIddcfa28_3964,
        RIddd0220_3965,RIddd0a18_3966,RIddd1210_3967,RIddd1a08_3968,RIdc0fbb8_3681,RIb86fc68_77,RIdc0f0f0_3682,RIb86fce0_76,RIdc0e5b0_3683,RIb86fd58_75,
        RIdc0dae8_3684,RIb87e8a8_74,RIdc0cfa8_3685,RIb87e920_73,RIdc0c3f0_3686,RIb87e998_72,RIdc0b7c0_3687,RIb87ea10_71,RIdc0ac08_3688,RIb87ea88_70,
        RIdc09f60_3689,RIdc093a8_3690,RIdc08700_3691,RIdc07878_3692,RIdc06270_3693,RIdc05118_3694,RIdc03b10_3695,RIdc029b8_3696,RIdc013b0_3697,RIdc00258_3698,
        RIdbff100_3699,RIdbfdaf8_3700,RIdbfc9a0_3701,RIdbfb398_3702,RIdbfa240_3703,RIdbf8c38_3704,RIdbf7ae0_3705,RIdbf6988_3706,RIdbf5380_3707,RIdbf4228_3708,
        RIdbf2c20_3709,RIdbf1ac8_3710,RIdbf04c0_3711,RIdbef368_3712,RIb79b428_272,RIe5efc28_6741,RIe527288_6346,RIe45e528_5951,RIe395df8_5556,RIe1ca840_5161,
        RIe100460_4766,RIe036f80_4371,RIde6b9c8_3976,RIdda31a8_3581,RIdbd9c48_3186,RIdb0e968_2791,RIda3bc30_2396,RId987e10_2001,RId8bc950_1606,RId7f4028_1211,
        RId72b4a8_816,RIe5d6d40_6768,RIe5117a8_6369,RIe444fb0_5975,RIe37f9b8_5584,RIe1ac2a0_5191,RIe0e8ec8_4791,RIe022a30_4393,RIdd8ba30_3609,RIdbc4870_3212,
        RIdaf5f30_2820,RIda25c28_2423,RId96d278_2032,RId8aa728_1632,RId7dcb80_1235,RId710748_846,RIe3ac2b0_6083,RIe3aaca8_6084,RIe3a9b50_6085,RIe3a8548_6086,
        RIe3a73f0_6087,RIe3a6298_6088,RIe3a4c90_6089,RIe3a3b38_6090,RIe3a2530_6091,RIe3a13d8_6092,RIe39fdd0_6093,RIe39ec78_6094,RIe39db20_6095,RIe39c518_6096,
        RIe1694d8_6097,RIe16e398_6098,RIe173270_6099,RIe178388_6100,RIe17c780_6101,RIe1805d8_6102,RIe1877c0_6103,RIe18c9c8_6104,RIe192ff8_6105,RIe198cc8_6106,
        RIe1a05b8_6107,RIe1a6300_6108,RIe1ac318_6109,RIe1b2420_6110,RIe1b7970_6111,RIe1bce48_6112,RIe1c12b8_6113,RIe1c7960_6114,RIe1cc820_6115,RIe1d0fd8_6116,
        RIe094940_6117,RIe090368_6118,RIe08b700_6119,RIe087a10_6120,RIe14c9f0_6121,RIe1495e8_6122,RIe146348_6123,RIe143210_6124,RIe140a38_6125,RIe13d4c8_6126,
        RIe13a660_6127,RIe137168_6128,RIe133a18_6129,RIe12fda0_6130,RIe1280f0_6131,RIe121b38_6132,RIe1194b0_6133,RIe1133a8_6134,RIe10ad20_6135,RIdfd70d0_6136,
        RIdff52b0_6137,RIe01ea70_6138,RIe03a5e0_6139,RIdfb6cb8_6140,RIdfa46d0_6141,RIdf7c7e8_6142,RIdc22218_6143,RIda953d8_6144,RIddeaf80_6145,RIde58a80_6146,
        RIe03fa40_6147,RIe04e338_6148,RIe0629f0_6149,RIe06c608_6150,RIe0732e0_6151,RIe07d0d8_6152,RIe084158_6153,RIdfc61e0_6154,RIe106838_6155,RIe0f8198_6156,
        RIe0eed00_6157,RIe0e2b68_6158,RIe0d0b98_6159,RIe0c3998_6160,RIe0b0960_6161,RIe0a6988_6162,RIe099440_6163,RIe1d3c60_6164,RIe1d69d8_6165,RIe1d9c00_6166,
        RIe1dc978_6167,RIe1dfba0_6168,RIe1e2918_6169,RIe1e5b40_6170,RIe1e88b8_6171,RIe1eb180_6172,RIe1ee858_6173,RIe1f1120_6174,RIe1f47f8_6175,RIe1f70c0_6176,
        RIe1fa180_6177,RIe1fbad0_6178,RIe1fd330_6179,RIe1ff568_6180,RIe2012f0_6181,RIe203000_6182,RIe203f00_6183,RIe2053a0_6184,RIe2066d8_6185,RIe207920_6186,
        RIe208be0_6187,RIe209d38_6188,RIe20b958_6189,RIe20cf60_6190,RIe20e4f0_6191,RIe20f5d0_6192,RIe211178_6193,RIe212c30_6194,RIe214148_6195,RIe215c00_6196,
        RIe217460_6197,RIe218798_6198,RIe2199e0_6199,RIe14e868_6200,RIe151130_6201,RIe153020_6202,RIe154ad8_6203,RIe156518_6204,RIe158228_6205,RIe15a280_6206,
        RIe15c3c8_6207,RIe15ef60_6208,RIe1616c0_6209,RIe164168_6210,RIe166c10_6211,RIe39a100_6212,RIe3984e0_6213,RIe3967d0_6214,RIe3941d8_6215,RIe391c58_6216,
        RIe38f5e8_6217,RIe38d428_6218,RIe38ae30_6219,RIe389030_6220,RIe386fd8_6221,RIe384ff8_6222,RIe3832e8_6223,RIe381218_6224,RIe37f148_6225,RIe37ce20_6226,
        RIe37aeb8_6227,RIe378668_6228,RIe3755a8_6229,RIe372c68_6230,RIe2703f8_6231,RIe26d4a0_6232,RIe26aae8_6233,RIe2686d0_6234,RIe265ca0_6235,RIe264170_6236,
        RIe2616c8_6237,RIe25f238_6238,RIe25c6a0_6239,RIe259ec8_6240,RIe257240_6241,RIe254018_6242,RIe251408_6243,RIe24e8e8_6244,RIe24c110_6245,RIe248d08_6246,
        RIe246170_6247,RIe2435d8_6248,RIe2418c8_6249,RIe23fb40_6250,RIe23dcc8_6251,RIe23ba18_6252,RIe239948_6253,RIe2381d8_6254,RIe236720_6255,RIe2346c8_6256,
        RIe232a30_6257,RIe230bb8_6258,RIe465cb0_6259,RIe4664a8_6260,RIe466ca0_6261,RIe467498_6262,RIe467c90_6263,RIe468488_6264,RIe468c80_6265,RIe469478_6266,
        RIe469c70_6267,RIe46a468_6268,RIe46ac60_6269,RIe46b458_6270,RIe46bc50_6271,RIe46c448_6272,RIe46cc40_6273,RIe46d438_6274,RIe46dc30_6275,RIe46e428_6276,
        RIe46ec20_6277,RIe46f418_6278,RIe46fc10_6279,RIe470408_6280,RIe470c00_6281,RIe4713f8_6282,RIe471bf0_6283,RIe4723e8_6284,RIe472bf8_6285,RIe4733f0_6286,
        RIe473be8_6287,RIe4743e0_6288,RIe474bd8_6289,RIe4753d0_6290,RIe475bc8_6291,RIe4763c0_6292,RIe476bb8_6293,RIe4773b0_6294,RIe477ba8_6295,RIe4783a0_6296,
        RIe478b98_6297,RIe479390_6298,RIe479b88_6299,RIe47a380_6300,RIe47ab78_6301,RIe47b370_6302,RIe47bb68_6303,RIe47c360_6304,RIe47cb58_6305,RIe47d350_6306,
        RIe47db48_6307,RIe47e340_6308,RIe47eb38_6309,RIe47f330_6310,RIe47fb28_6311,RIe480320_6312,RIe480b18_6313,RIe481310_6314,RIe481b08_6315,RIe482300_6316,
        RIe482af8_6317,RIe4832f0_6318,RIe483ae8_6319,RIe4842e0_6320,RIe484ad8_6321,RIe4852d0_6322,RIe485ac8_6323,RIe4862c0_6324,RIe486ab8_6325,RIe4872b0_6326,
        RIe487aa8_6327,RIe4882a0_6328,RIe488a98_6329,RIe489290_6330,RIe489a88_6331,RIe48a280_6332,RIe48aa78_6333,RIe48b270_6334,RIe48ba68_6335,RIe48c260_6336,
        RIe48ca58_6337,RIe48d250_6338,RIe3cd190_6051,RIe3cc3f8_6052,RIe3cb750_6053,RIe3ca9b8_6054,RIe3c9e00_6055,RIe3c9248_6056,RIe3c8708_6057,RIe3c7bc8_6058,
        RIe3c7100_6059,RIe3c6638_6060,RIe3c5af8_6061,RIe3c4ec8_6062,RIe3c4130_6063,RIe3c31b8_6064,RIe3c1bb0_6065,RIe3c0a58_6066,RIe3bf900_6067,RIe3be2f8_6068,
        RIe3bd1a0_6069,RIe3bbb98_6070,RIe3baa40_6071,RIe3b9438_6072,RIe3b82e0_6073,RIe3b7188_6074,RIe3b5b80_6075,RIe3b4a28_6076,RIe3b3420_6077,RIe3b22c8_6078,
        RIe3b0cc0_6079,RIe3afb68_6080,RIe3aea10_6081,RIe3ad408_6082,RIe51b690_6365,RIe500d68_6388,RIe501998_6387,RIe5026b8_6386,RIe5032e8_6385,RIe503f90_6384,
        RIe504d28_6383,RIe505958_6382,RIe50ef58_6371,RIe50ac50_6376,RIe50b880_6375,RIe50c690_6374,RIe50d428_6373,RIe523688_6352,RIe524060_6351,RIe524948_6350,
        RIe51c158_6364,RIe51cc20_6363,RIe51d5f8_6362,RIe5267c0_6347,RIe525d70_6348,RIe525410_6349,RIe51f290_6359,RIe51e840_6360,RIe51dee0_6361,RIe1e2210_5688,
        RIe1e10b8_5689,RIe1dfab0_5690,RIe1de958_5691,RIe1dd350_5692,RIe1dc1f8_5693,RIe1dabf0_5694,RIe1d9a98_5695,RIe1d8940_5696,RIe1d7338_5697,RIe1d61e0_5698,
        RIe1d4bd8_5699,RIe1d3a80_5700,RIe1d2478_5701,RIe099530_5702,RIe09d298_5703,RIe0a2338_5704,RIe0a6fa0_5705,RIe0ac310_5706,RIe0b16f8_5707,RIe0b9240_5708,
        RIe0bf438_5709,RIe0c4730_5710,RIe0cb0a8_5711,RIe0d0df0_5712,RIe0d8aa0_5713,RIe0de608_5714,RIe0e5ca0_5715,RIe0eb358_5716,RIe0ef138_5717,RIe0f3bc0_5718,
        RIe0f8300_5719,RIe0ff380_5720,RIe103430_5721,RIdfce868_5722,RIdfc9fc0_5723,RIdfc6000_5724,RIdfc1410_5725,RIdfbcc58_5726,RIe082f10_5727,RIe0800a8_5728,
        RIe07bd28_5729,RIe078ec0_5730,RIe075ab8_5731,RIe071f18_5732,RIe06f308_5733,RIe06b0f0_5734,RIe067928_5735,RIe0608a8_5736,RIe05a2f0_5737,RIe0541e8_5738,
        RIe04bb60_5739,RIe045a58_5740,RIe03d3d0_5741,RIde1d908_5742,RIde4a200_5743,RIde62e18_5744,RIdc30d68_5745,RIdde3e10_5746,RIddce948_5747,RIdb96b50_5748,
        RIda0b300_5749,RIdc00960_5750,RIdb708e8_5751,RIdc692d0_5752,RIdf7e930_5753,RIdf8d6d8_5754,RIdf9f978_5755,RIdfa6f20_5756,RIdfaf968_5757,RIdfb74b0_5758,
        RIddf5a98_5759,RIde028d8_5760,RIe036620_5761,RIe027530_5762,RIe01deb8_5763,RIe00b3a8_5764,RIdffd938_5765,RIdfefb08_5766,RIdfe0838_5767,RIdfd6680_5768,
        RIe1084d0_5769,RIe10ad98_5770,RIe10e470_5771,RIe110d38_5772,RIe113ab0_5773,RIe116cd8_5774,RIe119a50_5775,RIe11cc78_5776,RIe11f9f0_5777,RIe122c18_5778,
        RIe125990_5779,RIe128258_5780,RIe12b930_5781,RIe12e1f8_5782,RIe1308e0_5783,RIe132398_5784,RIe134300_5785,RIe135ae8_5786,RIe137258_5787,RIe138608_5788,
        RIe139850_5789,RIe13ab88_5790,RIe13c028_5791,RIe13d5b8_5792,RIe13ead0_5793,RIe13fef8_5794,RIe141230_5795,RIe142568_5796,RIe1434e0_5797,RIe144638_5798,
        RIe145880_5799,RIe146ac8_5800,RIe1486e8_5801,RIe149f48_5802,RIe14b550_5803,RIe14c978_5804,RIe14e430_5805,RIe0865e8_5806,RIe087f38_5807,RIe089db0_5808,
        RIe08b7f0_5809,RIe08d578_5810,RIe08f120_5811,RIe091100_5812,RIe093248_5813,RIe0950c0_5814,RIe096998_5815,RIe0986a8_5816,RIe1cfd18_5817,RIe1ce080_5818,
        RIe1cc550_5819,RIe1ca048_5820,RIe1c78e8_5821,RIe1c4f30_5822,RIe1c26e0_5823,RIe1c0b38_5824,RIe1be9f0_5825,RIe1bcce0_5826,RIe1baf58_5827,RIe1b9158_5828,
        RIe1b6908_5829,RIe1b3b90_5830,RIe1b1d18_5831,RIe1aff90_5832,RIe1ae2f8_5833,RIe1ab940_5834,RIe1a8628_5835,RIe1a6030_5836,RIe1a2d90_5837,RIe1a0540_5838,
        RIe19da20_5839,RIe19a870_5840,RIe197cd8_5841,RIe195410_5842,RIe192e90_5843,RIe190460_5844,RIe18e0c0_5845,RIe18bc30_5846,RIe189098_5847,RIe186c08_5848,
        RIe1839e0_5849,RIe1817a8_5850,RIe17fb88_5851,RIe17def0_5852,RIe17c3c0_5853,RIe17a458_5854,RIe1781a8_5855,RIe176240_5856,RIe174530_5857,RIe172988_5858,
        RIe16fc70_5859,RIe16e140_5860,RIe16c1d8_5861,RIe16a5b8_5862,RIe168a88_5863,RIe167138_5864,RIe39c680_5865,RIe39ce78_5866,RIe39d670_5867,RIe39de68_5868,
        RIe39e660_5869,RIe39ee58_5870,RIe39f650_5871,RIe39fe48_5872,RIe3a0640_5873,RIe3a0e38_5874,RIe3a1630_5875,RIe3a1e28_5876,RIe3a2620_5877,RIe3a2e18_5878,
        RIe3a3610_5879,RIe3a3e08_5880,RIe3a4600_5881,RIe3a4df8_5882,RIe3a55f0_5883,RIe3a5de8_5884,RIe3a65e0_5885,RIe3a6dd8_5886,RIe3a75d0_5887,RIe3a7dc8_5888,
        RIe3a85c0_5889,RIe3a8db8_5890,RIe3a95b0_5891,RIe3a9da8_5892,RIe3aa5a0_5893,RIe3aad98_5894,RIe3ab590_5895,RIe3abd88_5896,RIe3ac580_5897,RIe3acd78_5898,
        RIe3ad570_5899,RIe3add68_5900,RIe3ae560_5901,RIe3aed58_5902,RIe3af550_5903,RIe3afd48_5904,RIe3b0540_5905,RIe3b0d38_5906,RIe3b1530_5907,RIe3b1d28_5908,
        RIe3b2520_5909,RIe3b2d18_5910,RIe3b3510_5911,RIe3b3d08_5912,RIe3b4500_5913,RIe3b4cf8_5914,RIe3b54f0_5915,RIe3b5ce8_5916,RIe3b64e0_5917,RIe3b6cd8_5918,
        RIe3b74d0_5919,RIe3b7cc8_5920,RIe3b84c0_5921,RIe3b8cb8_5922,RIe3b94b0_5923,RIe3b9ca8_5924,RIe3ba4a0_5925,RIe3bac98_5926,RIe3bb490_5927,RIe3bbc88_5928,
        RIe3bc480_5929,RIe3bcc78_5930,RIe3bd470_5931,RIe3bdc68_5932,RIe3be460_5933,RIe3bec58_5934,RIe3bf450_5935,RIe3bfc48_5936,RIe3c0440_5937,RIe3c0c38_5938,
        RIe3c1430_5939,RIe3c1c28_5940,RIe3c2420_5941,RIe3c2c18_5942,RIe3c3410_5943,RIe202f10_5656,RIe202448_5657,RIe201980_5658,RIe200e40_5659,RIe2000a8_5660,
        RIe1ff310_5661,RIe1fe668_5662,RIe1fd9c0_5663,RIe1fce80_5664,RIe1fc340_5665,RIe1fb878_5666,RIe1facc0_5667,RIe1fa090_5668,RIe1f9118_5669,RIe1f7fc0_5670,
        RIe1f69b8_5671,RIe1f5860_5672,RIe1f4258_5673,RIe1f3100_5674,RIe1f1fa8_5675,RIe1f09a0_5676,RIe1ef848_5677,RIe1ee240_5678,RIe1ed0e8_5679,RIe1ebae0_5680,
        RIe1ea988_5681,RIe1e9830_5682,RIe1e8228_5683,RIe1e70d0_5684,RIe1e5ac8_5685,RIe1e4970_5686,RIe1e3368_5687,RIe4520c0_5970,RIe438440_5990,RIe4390e8_5989,
        RIe439f70_5988,RIe43ad80_5987,RIe43ba28_5986,RIe43c7c0_5985,RIe43d5d0_5984,RIe445e38_5974,RIe441c98_5979,RIe4429b8_5978,RIe443750_5977,RIe437630_5991,
        RIe45a478_5957,RIe45aec8_5956,RIe45b8a0_5955,RIe452b88_5969,RIe4534e8_5968,RIe453fb0_5967,RIe45d880_5952,RIe45cdb8_5953,RIe45c278_5954,RIe455e28_5964,
        RIe4554c8_5965,RIe454988_5966,RIe116b70_5293,RIe115a18_5294,RIe114410_5295,RIe1132b8_5296,RIe111cb0_5297,RIe110b58_5298,RIe10f550_5299,RIe10e3f8_5300,
        RIe10d2a0_5301,RIe10bc98_5302,RIe10ab40_5303,RIe109538_5304,RIe1083e0_5305,RIe106dd8_5306,RIdfd3728_5307,RIdfd71c0_5308,RIdfdc8f0_5309,RIdfe0b80_5310,
        RIdfe6760_5311,RIdfeb788_5312,RIdff1f98_5313,RIdff7f38_5314,RIdffe400_5315,RIe005750_5316,RIe00b420_5317,RIe0132b0_5318,RIe0193b8_5319,RIe0202d0_5320,
        RIe023de0_5321,RIe027878_5322,RIe02ccd8_5323,RIe0322a0_5324,RIe038768_5325,RIe03c728_5326,RIde01258_5327,RIddfd748_5328,RIddf9788_5329,RIddf3d88_5330,
        RIdfba228_5331,RIdfb5e30_5332,RIdfb2aa0_5333,RIdfaec48_5334,RIdfabf48_5335,RIdfa97e8_5336,RIdfa5e40_5337,RIdfa2f60_5338,RIdf9e4d8_5339,RIdf99618_5340,
        RIdf90f90_5341,RIdf8ae88_5342,RIdf848d0_5343,RIdf7c248_5344,RIdf76140_5345,RIdc56298_5346,RIdd75f50_5347,RIdd9d6b8_5348,RIdb67180_5349,RIdc198c0_5350,
        RIdc008e8_5351,RIdacdc88_5352,RId8fd180_5353,RIdb353b0_5354,RIdbdbca0_5355,RIdb8b8b8_5356,RIddb1a28_5357,RIddc60e0_5358,RIddd3cb8_5359,RIdddeaa0_5360,
        RIdde50d0_5361,RIddeee50_5362,RIdc2bb60_5363,RIdc34788_5364,RIde6e7b8_5365,RIde62ad0_5366,RIde55510_5367,RIde4a188_5368,RIde36d90_5369,RIde29c80_5370,
        RIde1c210_5371,RIde0cb08_5372,RIe03d4c0_5373,RIe040b98_5374,RIe043460_5375,RIe046b38_5376,RIe049400_5377,RIe04c178_5378,RIe04f3a0_5379,RIe052118_5380,
        RIe055340_5381,RIe0580b8_5382,RIe05b2e0_5383,RIe05e058_5384,RIe060920_5385,RIe063ff8_5386,RIe0662a8_5387,RIe068288_5388,RIe069a70_5389,RIe06b870_5390,
        RIe06cf68_5391,RIe06e6d8_5392,RIe06fa10_5393,RIe070eb0_5394,RIe0721e8_5395,RIe073808_5396,RIe074960_5397,RIe0762b0_5398,RIe0779a8_5399,RIe079118_5400,
        RIe07a798_5401,RIe07bcb0_5402,RIe07d768_5403,RIe07f220_5404,RIe080cd8_5405,RIe082088_5406,RIe083078_5407,RIe0843b0_5408,RIdfbbbf0_5409,RIdfbd5b8_5410,
        RIdfbf3b8_5411,RIdfc15f0_5412,RIdfc30a8_5413,RIdfc4f20_5414,RIdfc6f00_5415,RIdfc85f8_5416,RIdfca3f8_5417,RIdfcc720_5418,RIdfce8e0_5419,RIe106478_5420,
        RIe104948_5421,RIe102b48_5422,RIe100f28_5423,RIe0fea20_5424,RIe0fcd10_5425,RIe0fa3d0_5426,RIe0f7838_5427,RIe0f5a38_5428,RIe0f3968_5429,RIe0f1b68_5430,
        RIe0f0290_5431,RIe0ee508_5432,RIe0ec690_5433,RIe0eaea8_5434,RIe0e8658_5435,RIe0e54a8_5436,RIe0e2988_5437,RIe0e0228_5438,RIe0dd7f8_5439,RIe0da828_5440,
        RIe0d7f60_5441,RIe0d4f18_5442,RIe0d3280_5443,RIe0d02b0_5444,RIe0cdad8_5445,RIe0cae50_5446,RIe0c8150_5447,RIe0c5d38_5448,RIe0c3290_5449,RIe0c0d88_5450,
        RIe0be628_5451,RIe0bbdd8_5452,RIe0b91c8_5453,RIe0b5f28_5454,RIe0b3318_5455,RIe0b02d0_5456,RIe0adeb8_5457,RIe0ac0b8_5458,RIe0aa330_5459,RIe0a83c8_5460,
        RIe0a6a00_5461,RIe0a40c0_5462,RIe0a2158_5463,RIe0a0010_5464,RIe09e378_5465,RIe09c668_5466,RIe09a8e0_5467,RIe099080_5468,RIe1d1cf8_5469,RIe1d24f0_5470,
        RIe1d2ce8_5471,RIe1d34e0_5472,RIe1d3cd8_5473,RIe1d44d0_5474,RIe1d4cc8_5475,RIe1d54c0_5476,RIe1d5cb8_5477,RIe1d64b0_5478,RIe1d6ca8_5479,RIe1d74a0_5480,
        RIe1d7c98_5481,RIe1d8490_5482,RIe1d8c88_5483,RIe1d9480_5484,RIe1d9c78_5485,RIe1da470_5486,RIe1dac68_5487,RIe1db460_5488,RIe1dbc58_5489,RIe1dc450_5490,
        RIe1dcc48_5491,RIe1dd440_5492,RIe1ddc38_5493,RIe1de430_5494,RIe1dec28_5495,RIe1df420_5496,RIe1dfc18_5497,RIe1e0410_5498,RIe1e0c08_5499,RIe1e1400_5500,
        RIe1e1bf8_5501,RIe1e23f0_5502,RIe1e2be8_5503,RIe1e33e0_5504,RIe1e3bd8_5505,RIe1e43d0_5506,RIe1e4bc8_5507,RIe1e53c0_5508,RIe1e5bb8_5509,RIe1e63b0_5510,
        RIe1e6ba8_5511,RIe1e73a0_5512,RIe1e7b98_5513,RIe1e8390_5514,RIe1e8b88_5515,RIe1e9380_5516,RIe1e9b78_5517,RIe1ea370_5518,RIe1eab68_5519,RIe1eb360_5520,
        RIe1ebb58_5521,RIe1ec350_5522,RIe1ecb48_5523,RIe1ed340_5524,RIe1edb38_5525,RIe1ee330_5526,RIe1eeb28_5527,RIe1ef320_5528,RIe1efb18_5529,RIe1f0310_5530,
        RIe1f0b08_5531,RIe1f1300_5532,RIe1f1af8_5533,RIe1f22f0_5534,RIe1f2ae8_5535,RIe1f32e0_5536,RIe1f3ad8_5537,RIe1f42d0_5538,RIe1f4ac8_5539,RIe1f52c0_5540,
        RIe1f5ab8_5541,RIe1f62b0_5542,RIe1f6aa8_5543,RIe1f72a0_5544,RIe1f7a98_5545,RIe1f8290_5546,RIe1f8a88_5547,RIe1f9280_5548,RIe137870_5261,RIe136da8_5262,
        RIe136358_5263,RIe135890_5264,RIe134d50_5265,RIe134288_5266,RIe1337c0_5267,RIe132c08_5268,RIe131fd8_5269,RIe1313a8_5270,RIe1307f0_5271,RIe12fbc0_5272,
        RIe12f080_5273,RIe12da78_5274,RIe12c920_5275,RIe12b318_5276,RIe12a1c0_5277,RIe128bb8_5278,RIe127a60_5279,RIe126908_5280,RIe125300_5281,RIe1241a8_5282,
        RIe122ba0_5283,RIe121a48_5284,RIe120440_5285,RIe11f2e8_5286,RIe11e190_5287,RIe11cb88_5288,RIe11ba30_5289,RIe11a428_5290,RIe1192d0_5291,RIe117cc8_5292,
        RIe38a110_5575,RIe378410_5590,RIe379220_5589,RIe379e50_5588,RIe26f4f8_5601,RIe270290_5600,RIe270ec0_5599,RIe271be0_5598,RIe37b908_5586,RIe375008_5594,
        RIe375da0_5593,RIe376a48_5592,RIe377768_5591,RIe3921f8_5562,RIe392b58_5561,RIe3934b8_5560,RIe38a908_5574,RIe38b1f0_5573,RIe38b9e8_5572,RIe3951c8_5557,
        RIe394868_5558,RIe393e90_5559,RIe38da40_5569,RIe38cf78_5570,RIe38c4b0_5571,RIe04cad8_4898,RIe04b980_4899,RIe04a378_4900,RIe049220_4901,RIe047c18_4902,
        RIe046ac0_4903,RIe045968_4904,RIe044360_4905,RIe043208_4906,RIe041c00_4907,RIe040aa8_4908,RIe03f4a0_4909,RIe03e348_4910,RIe03d1f0_4911,RIde08bc0_4912,
        RIde0d030_4913,RIde131b0_4914,RIde17968_4915,RIde1f528_4916,RIde24e38_4917,RIde29ed8_4918,RIde31390_4919,RIde36e08_4920,RIde3efe0_4921,RIde45070_4922,
        RIde4c9d8_4923,RIde51b68_4924,RIde553a8_4925,RIde59c50_4926,RIde5e390_4927,RIde65668_4928,RIde6a4b0_4929,RIde6f820_4930,RIdf73710_4931,RIdc38040_4932,
        RIdc32b68_4933,RIdc2ee78_4934,RIdc29bf8_4935,RIddf1628_4936,RIddee388_4937,RIddeaa58_4938,RIdde7a88_4939,RIdde35a0_4940,RIdde0cd8_4941,RIddddf60_4942,
        RIdddb710_4943,RIddd5e78_4944,RIddd2278_4945,RIddcc080_4946,RIddc39f8_4947,RIddbd8f0_4948,RIddb5268_4949,RIddaf160_4950,RIdb7c228_4951,RIdb96c40_4952,
        RIdbbbd38_4953,RIdbdcdf8_4954,RIdb5db80_4955,RIdb48190_4956,RIdb26ba8_4957,RId917aa8_4958,RId986da8_4959,RIda7eb60_4960,RIdaf90e0_4961,RIdab27a8_4962,
        RIdbf1ca8_4963,RIdc00a50_4964,RIdc0fe88_4965,RIdc16080_4966,RIdc1c098_4967,RIdc25080_4968,RIdb67810_4969,RIdda8518_4970,RIdd9d5c8_4971,RIdd8f270_4972,
        RIdd82fe8_4973,RIdd74150_4974,RIdc641b8_4975,RIdc54600_4976,RIdc46848_4977,RIdc3b970_4978,RIdf77220_4979,RIdf79f98_4980,RIdf7c860_4981,RIdf7ff38_4982,
        RIdf82800_4983,RIdf85ed8_4984,RIdf887a0_4985,RIdf8be78_4986,RIdf8e740_4987,RIdf91008_4988,RIdf946e0_4989,RIdf96fa8_4990,RIdf9a680_4991,RIdf9ccf0_4992,
        RIdf9ec58_4993,RIdfa04b8_4994,RIdfa1bb0_4995,RIdfa3b18_4996,RIdfa4dd8_4997,RIdfa6110_4998,RIdfa75b0_4999,RIdfa88e8_5000,RIdfa9d10_5001,RIdfab048_5002,
        RIdfac218_5003,RIdfad460_5004,RIdfaecc0_5005,RIdfb0610_5006,RIdfb1c90_5007,RIdfb3310_5008,RIdfb4828_5009,RIdfb5d40_5010,RIdfb77f8_5011,RIdfb92b0_5012,
        RIdfba9a8_5013,RIddf2ca8_5014,RIddf4580_5015,RIddf6308_5016,RIddf8270_5017,RIddf9e90_5018,RIddfbdf8_5019,RIddfdb08_5020,RIddff548_5021,RIde015a0_5022,
        RIde03508_5023,RIde04fc0_5024,RIe03bbe8_5025,RIe039cf8_5026,RIe038600_5027,RIe0363c8_5028,RIe033b78_5029,RIe031580_5030,RIe02ee98_5031,RIe02c4e0_5032,
        RIe02a488_5033,RIe028958_5034,RIe026b58_5035,RIe025460_5036,RIe023b88_5037,RIe021fe0_5038,RIe020168_5039,RIe01dcd8_5040,RIe01b758_5041,RIe018440_5042,
        RIe0157b8_5043,RIe012590_5044,RIe010628_5045,RIe00d298_5046,RIe00a778_5047,RIe007e38_5048,RIe004df0_5049,RIe0024b0_5050,RIdfff558_5051,RIdffcd08_5052,
        RIdffa260_5053,RIdff7b78_5054,RIdff4f68_5055,RIdff1ea8_5056;
output R_25610_96cc360,R_25642_95f0d48,R_25644_9598060,R_25646_95984f8,R_25614_953c348,R_25616_96251f8,R_25618_96ed6b0,R_2561a_95f00d0,R_2561c_95f0418,
        R_2561e_95f0760,R_25620_953c3f0,R_25622_953c690,R_25612_953c9d8,R_25624_95f08b0,R_25626_953ca80,R_25628_96253f0,R_2562a_9632be8,R_253fc_9d20ef0,R_25412_9530108,
        R_25428_95f75a0,R_2543e_95301b0,R_25454_95304f8,R_2546a_9533198,R_25474_95332e8,R_25476_96dee60,R_25478_95f7798,R_2547a_96def08,R_253fe_95f7990,R_25400_9d21190,
        R_25402_9d21388,R_25404_9589e90,R_25406_9d21430,R_25408_9533780,R_2540a_9533b70,R_2540c_9d216d0,R_2540e_958a5c8,R_25410_96defb0,R_25414_9d21778,R_25416_9d21cb8,
        R_25418_95f7ae0,R_2541a_9d21d60,R_2541c_96df100,R_2541e_9d221f8,R_25420_958ac58,R_25422_95f7b88,R_25424_9533c18,R_25426_958b630,R_2542a_9d222a0,R_2542c_9533d68,
        R_2542e_95f7c30,R_25430_9d22498,R_25432_9d22540,R_25434_9533f60,R_25436_96df1a8,R_25438_95f7f78,R_2543a_9534008,R_2543c_9534200,R_25440_95f80c8,R_25442_96df250,
        R_25444_9d22690,R_25446_95fa438,R_25448_95fa4e0,R_2544a_958bcc0,R_2544c_9d22738,R_2544e_9d227e0,R_25450_9d22888,R_25452_9d22930,R_25456_9d229d8,R_25458_95fa588,
        R_2545a_9534350,R_2545c_95fa828,R_2545e_9d22a80,R_25460_96df2f8,R_25462_96df3a0,R_25464_95343f8,R_25466_95fa8d0,R_25468_95faac8,R_2546c_958bd68,R_2546e_958be10,
        R_25470_95fab70,R_25472_9d22b28,R_2547c_958beb8,R_25492_9d22bd0,R_254a8_958bf60,R_254be_9d22c78,R_254d4_9d22dc8,R_254ea_9d22e70,R_254f4_958c0b0,R_254f6_9d22f18,
        R_254f8_958c158,R_254fa_9d22fc0,R_2547e_958c200,R_25480_9d23068,R_25482_9d231b8,R_25484_958c2a8,R_25486_958c350,R_25488_9d23458,R_2548a_958c4a0,R_2548c_9d235a8,
        R_2548e_9d236f8,R_25490_958c548,R_25494_958c5f0,R_25496_9d237a0,R_25498_958c698,R_2549a_958f728,R_2549c_9d23848,R_2549e_958f7d0,R_254a0_958f878,R_254a2_9d23998,
        R_254a4_9d23ae8,R_254a6_9d23c38,R_254aa_9d23d88,R_254ac_9d23e30,R_254ae_9d23f80,R_254b0_9d24028,R_254b2_9d240d0,R_254b4_9d24220,R_254b6_9d242c8,R_254b8_9590988,
        R_254ba_9590a30,R_254bc_9590cd0,R_254c0_9d24418,R_254c2_9590d78,R_254c4_9590f70,R_254c6_9591178,R_254c8_9d24568,R_254ca_9d24bf8,R_254cc_9d25090,R_254ce_95916b8,
        R_254d0_9591808,R_254d2_9d251e0,R_254d6_9d25f10,R_254d8_9d25fb8,R_254da_95918b0,R_254dc_9d265a0,R_254de_9591958,R_254e0_9d26990,R_254e2_9d26c30,R_254e4_9591a00,
        R_254e6_95347e8,R_254e8_9591b50,R_254ec_9591bf8,R_254ee_9d26d80,R_254f0_9d27368,R_254f2_9d27410,R_254fc_96df4f0,R_25512_9d276b0,R_25528_96df598,R_2553e_9534890,
        R_25554_9d27c98,R_2556a_96df640,R_25574_9d27de8,R_25576_96df6e8,R_25578_9534bd8,R_2557a_96df838,R_254fe_96dfad8,R_25500_9534d28,R_25502_9534dd0,R_25504_9534f20,
        R_25506_9d281d8,R_25508_96dfb80,R_2550a_9d28328,R_2550c_9d283d0,R_2550e_96dfc28,R_25510_9534fc8,R_25514_96dfcd0,R_25516_9d28520,R_25518_96dfe20,R_2551a_96dfec8,
        R_2551c_9535070,R_2551e_95351c0,R_25520_9535268,R_25522_96dff70,R_25524_96e0018,R_25526_96e00c0,R_2552a_9535310,R_2552c_96e0168,R_2552e_96e0210,R_25530_96e02b8,
        R_25532_96e0408,R_25534_96e0558,R_25536_96e0600,R_25538_9535658,R_2553a_9d289b8,R_2553c_96e06a8,R_25540_95358f8,R_25542_96e0750,R_25544_96e0b40,R_25546_96e0be8,
        R_25548_96e0c90,R_2554a_96e0d38,R_2554c_95359a0,R_2554e_9d28a60,R_25550_96e0e88,R_25552_9535a48,R_25556_96e0f30,R_25558_9535b98,R_2555a_9d28c58,R_2555c_96e0fd8,
        R_2555e_9d28d00,R_25560_9535c40,R_25562_95362d0,R_25564_9536810,R_25566_9536a08,R_25568_96e1080,R_2556c_96e1128,R_2556e_9d28ef8,R_25570_96e11d0,R_25572_96e1c50,
        R_2557c_9591d48,R_25592_9591df0,R_255a8_96e2e08,R_255be_9591e98,R_255d4_9591f40,R_255ea_96e3690,R_255f4_96e6918,R_255f6_96e69c0,R_255f8_9d29048,R_255fa_9d28718,
        R_2557e_9591fe8,R_25580_96e6fa8,R_25582_96e72f0,R_25584_9d287c0,R_25586_9592090,R_25588_9592138,R_2558a_96e7398,R_2558c_9d28868,R_2558e_9d290f0,R_25590_9d29240,
        R_25594_96e7cc8,R_25596_95921e0,R_25598_9592288,R_2559a_9592330,R_2559c_96e82b0,R_2559e_9d292e8,R_255a0_9d2dfb0,R_255a2_9592528,R_255a4_9592678,R_255a6_9d2e058,
        R_255aa_96e8358,R_255ac_9592918,R_255ae_96e86a0,R_255b0_9d2e988,R_255b2_9d29390,R_255b4_9d2ec28,R_255b6_9d294e0,R_255b8_9d2f360,R_255ba_9592a68,R_255bc_9592b10,
        R_255c0_9d30128,R_255c2_9592c60,R_255c4_96e8940,R_255c6_96e89e8,R_255c8_9d30278,R_255ca_96e8be0,R_255cc_9592f00,R_255ce_9d29588,R_255d0_9d296d8,R_255d2_9d30518,
        R_255d6_9d29828,R_255d8_96e9120,R_255da_96e93c0,R_255dc_96e9510,R_255de_9d307b8,R_255e0_9d29cc0,R_255e2_9592fa8,R_255e4_9593050,R_255e6_96e9858,R_255e8_96e9a50,
        R_255ec_95930f8,R_255ee_9d29eb8,R_255f0_96ea038,R_255f2_95931a0,R_253bc_96eacb0,R_253be_9593248,R_253c0_9d29f60,R_253c2_95932f0,R_253c4_96eae00,R_253c6_9536b58,
        R_253c8_9593398,R_253ca_9d2a350,R_253cc_b7dc210,R_253ce_b7dcd38,R_253d0_b7dcde0,R_253d2_9593590,R_253d4_96376b8,R_253d6_9d2a4a0,R_253d8_9596038,R_253da_b7dc2b8,
        R_253dc_96eb0a0,R_253de_9596578,R_253e0_9536f48,R_253e2_96eb298,R_253e4_9537098,R_253e6_96eb340,R_253e8_95373e0,R_253ea_9596a10,R_253ec_9d30860,R_253ee_9ef0090,
        R_253f0_9d30f98,R_253f2_9ef05d0,R_253f4_9d31040,R_253f6_9d31238,R_253f8_9d314d8,R_253fa_9d316d0,R_25666_96346d0,R_1a4_b821b50,R_1a3_b821aa8,R_23ca4_96329f0,
        R_23cba_9f596e0,R_23cd0_962b7c0,R_23ce6_955f268,R_23cfc_9f5c4d0,R_23d12_9d225e8,R_23d1c_962b910,R_23d1e_95a3470,R_23d20_9632c90,R_23d22_95a3710,R_23ca6_9ee76c0,
        R_23ca8_9ee7810,R_23caa_9ee78b8,R_23cac_9ee8140,R_23cae_962bbb0,R_23cb0_9ee8920,R_23cb2_9d22d20,R_23cb4_9ee8bc0,R_23cb6_9632d38,R_23cb8_9d23110,R_23cbc_962bc58,
        R_23cbe_9ee9ad8,R_23cc0_9d23260,R_23cc2_9632f30,R_23cc4_9eec430,R_23cc6_9d23308,R_23cc8_9eef4c0,R_23cca_9eefca0,R_23ccc_9d23650,R_23cce_9ef0678,R_23cd2_95a3908,
        R_23cd4_962bd00,R_23cd6_9632fd8,R_23cd8_962be50,R_23cda_96331d0,R_23cdc_962bef8,R_23cde_9d30ef0,R_23ce0_9d238f0,R_23ce2_9d23b90,R_23ce4_962bfa0,R_23ce8_962c048,
        R_23cea_95a3a58,R_23cec_9d23ed8,R_23cee_9ef09c0,R_23cf0_9ef4380,R_23cf2_95a3ba8,R_23cf4_9ef4a10,R_23cf6_962c0f0,R_23cf8_96c3060,R_23cfa_96c6d68,R_23cfe_9d310e8,
        R_23d00_96c72a8,R_23d02_962c390,R_23d04_96c74a0,R_23d06_962da88,R_23d08_9d24178,R_23d0a_962df20,R_23d0c_9633278,R_23d0e_9633320,R_23d10_95a3e48,R_23d14_95a4040,
        R_23d16_9d24370,R_23d18_96c7e78,R_23d1a_96333c8,R_23d24_9633470,R_23d3a_9633518,R_23d50_962dfc8,R_23d66_9629b88,R_23d7c_95547c8,R_23d92_96335c0,R_23d9c_96337b8,
        R_23d9e_9633908,R_23da0_9633a58,R_23da2_962e7a8,R_23d26_9554870,R_23d28_962a560,R_23d2a_962ee38,R_23d2c_962a8a8,R_23d2e_962f2d0,R_23d30_95549c0,R_23d32_9633cf8,
        R_23d34_962f4c8,R_23d36_9633da0,R_23d38_9633e48,R_23d3c_9633ef0,R_23d3e_962c4e0,R_23d40_9554bb8,R_23d42_9554d08,R_23d44_9634040,R_23d46_962f6c0,R_23d48_9554f00,
        R_23d4a_962c8d0,R_23d4c_9635000,R_23d4e_962fab0,R_23d52_95552f0,R_23d54_96350a8,R_23d56_96351f8,R_23d58_962fc00,R_23d5a_95554e8,R_23d5c_9555638,R_23d5e_9635540,
        R_23d60_96355e8,R_23d62_9635738,R_23d64_96359d8,R_23d68_962ca20,R_23d6a_9635f18,R_23d6c_962ff48,R_23d6e_9636068,R_23d70_96363b0,R_23d72_9636ae8,R_23d74_9637220,
        R_23d76_9637e98,R_23d78_9638b10,R_23d7a_962d4a0,R_23d7e_96305d8,R_23d80_9638bb8,R_23d82_9638fa8,R_23d84_962d548,R_23d86_9639398,R_23d88_95556e0,R_23d8a_9639440,
        R_23d8c_9d18d00,R_23d8e_9d19d68,R_23d90_9630a70,R_23d94_9d1a008,R_23d96_9d1a350,R_23d98_9d1a9e0,R_23d9a_96314f0,R_23da4_9634430,R_23dba_95558d8,R_23dd0_9555a28,
        R_23de6_9d1ac80,R_23dfc_962d9e0,R_23e12_9555b78,R_23e1c_96344d8,R_23e1e_9555e18,R_23e20_9d1b070,R_23e22_9d1b8f8,R_23da6_9634a18,R_23da8_9555f68,R_23daa_9635150,
        R_23dac_96352a0,R_23dae_9556010,R_23db0_9557078,R_23db2_96353f0,R_23db4_9d1ba48,R_23db6_962db30,R_23db8_96357e0,R_23dbc_9559730,R_23dbe_955bde8,R_23dc0_955dd68,
        R_23dc2_9d1baf0,R_23dc4_955e158,R_23dc6_9638db0,R_23dc8_9d1bb98,R_23dca_9639248,R_23dcc_9d1bce8,R_23dce_96c81c0,R_23dd2_955e4a0,R_23dd4_955ea88,R_23dd6_96392f0,
        R_23dd8_9d15d18,R_23dda_955ee78,R_23ddc_9d168e8,R_23dde_9d16ae0,R_23de0_962e310,R_23de2_9d16c30,R_23de4_9d16e28,R_23de8_9d170c8,R_23dea_955f1c0,R_23dec_96c87a8,
        R_23dee_955f310,R_23df0_9d1bee0,R_23df2_955f3b8,R_23df4_95a39b0,R_23df6_96c8af0,R_23df8_95a3b00,R_23dfa_95a40e8,R_23dfe_95a44d8,R_23e00_9d1bf88,R_23e02_95a4580,
        R_23e04_95a4c10,R_23e06_9d17218,R_23e08_95a5348,R_23e0a_962ec40,R_23e0c_9d17608,R_23e0e_95a57e0,R_23e10_95a5930,R_23e14_9d18910,R_23e16_9d19630,R_23e18_95a5c78,
        R_23e1a_95a6260,R_23e24_9d1c030,R_23e3a_95a4628,R_23e50_95a48c8,R_23e66_95a4b68,R_23e7c_95b1438,R_23e92_9d19780,R_23e9c_95a6d88,R_23e9e_95b1780,R_23ea0_95a7028,
        R_23ea2_95a70d0,R_23e26_95b1828,R_23e28_95a7220,R_23e2a_95b2bd8,R_23e2c_95b3310,R_23e2e_95818b0,R_23e30_9582138,R_23e32_9582288,R_23e34_95a7760,R_23e36_9582870,
        R_23e38_95a78b0,R_23e3c_9d1c0d8,R_23e3e_9582a68,R_23e40_9d1b118,R_23e42_9582e58,R_23e44_9582f00,R_23e46_95830f8,R_23e48_958cbd8,R_23e4a_958cc80,R_23e4c_95a7aa8,
        R_23e4e_958f5d8,R_23e52_958f920,R_23e54_9590058,R_23e56_95a7bf8,R_23e58_95a7ca0,R_23e5a_95901a8,R_23e5c_959fdb8,R_23e5e_95a0b80,R_23e60_9d1c4c8,R_23e62_9625b28,
        R_23e64_96261b8,R_23e68_9d1b268,R_23e6a_9d1c570,R_23e6c_95a7d48,R_23e6e_9626458,R_23e70_95a8090,R_23e72_9628330,R_23e74_9628480,R_23e76_9628528,R_23e78_95a8138,
        R_23e7a_96285d0,R_23e7e_9628720,R_23e80_9628bb8,R_23e82_962c198,R_23e84_9d1c618,R_23e86_95a8288,R_23e88_9634238,R_23e8a_9d1c6c0,R_23e8c_96342e0,R_23e8e_9634970,
        R_23e90_9d1c8b8,R_23e94_9639830,R_23e96_9d159d0,R_23e98_9d15e68,R_23e9a_95a83d8,R_23c64_96c9a08,R_23c66_9d1b658,R_23c68_96ca920,R_23c6a_9d244c0,R_23c6c_96cb4f0,
        R_23c6e_9d1b700,R_23c70_9d1ca08,R_23c72_96cb640,R_23c74_962f030,R_23c76_9d1cc00,R_23c78_9d1cd50,R_23c7a_9d1cdf8,R_23c7c_9d1b7a8,R_23c7e_9d1cf48,R_23c80_9d1d098,
        R_23c82_9d1d1e8,R_23c84_95a8528,R_23c86_9d1b9a0,R_23c88_95a8720,R_23c8a_9d1be38,R_23c8c_9d246b8,R_23c8e_96cb838,R_23c90_9d24760,R_23c92_9d1c2d0,R_23c94_9d1d3e0,
        R_23c96_95a87c8,R_23c98_9d19438,R_23c9a_9d1c378,R_23c9c_9d1c768,R_23c9e_9d1d488,R_23ca0_9d1c960,R_23ca2_9d1e8e0,R_23ebc_9667ae0,R_23ebe_965f6f8,R_23ec0_9667b88,
        R_23ec2_96688a8,R_23ec4_95ac230,R_23ec6_95ac428,R_23ec8_966a780,R_23eca_966a8d0,R_23eba_965f8f0,R_23ecc_95ac620,R_23ece_95ac770,R_23ed0_966a978,R_23ed2_966aa20,
        R_23eb8_966aac8,R_23eea_95b1588,R_23eec_9d1e448,R_23eee_9d1e790,R_23a0c_95b1630,R_23a22_95b1c18,R_23a38_966acc0,R_23a4e_95b1d68,R_23a64_966ad68,R_23a7a_95b2c80,
        R_23a84_9661a68,R_23a86_9d1d7d0,R_23a88_966ae10,R_23a8a_966b0b0,R_23a0e_962f420,R_23a10_966ba88,R_23a12_95b2fc8,R_23a14_9d1f6a8,R_23a16_952daf8,R_23a18_95b3268,
        R_23a1a_9581220,R_23a1c_9d1d878,R_23a1e_9663160,R_23a20_9d1e250,R_23a24_9d1fb40,R_23a26_95305a0,R_23a28_95812c8,R_23a2a_9530798,R_23a2c_95816b8,R_23a2e_9663550,
        R_23a30_9531e90,R_23a32_9531f38,R_23a34_9532130,R_23a36_9532280,R_23a3a_9532328,R_23a3c_9581760,R_23a3e_9581f40,R_23a40_95323d0,R_23a42_9532868,R_23a44_9582720,
        R_23a46_9532b08,R_23a48_9532c58,R_23a4a_9582918,R_23a4c_966a4e0,R_23a50_9532e50,R_23a52_9d24808,R_23a54_9533390,R_23a56_9d20668,R_23a58_9582db0,R_23a5a_9583050,
        R_23a5c_9533978,R_23a5e_9534158,R_23a60_9d20710,R_23a62_95349e0,R_23a66_9537290,R_23a68_9d1f750,R_23a6a_966a6d8,R_23a6c_966aeb8,R_23a6e_966b158,R_23a70_9537a70,
        R_23a72_9539f30,R_23a74_95831a0,R_23a76_9537c68,R_23a78_9d20a58,R_23a7c_9537d10,R_23a7e_9537e60,R_23a80_9538250,R_23a82_95382f8,R_23a8c_9d21e08,R_23aa2_9583440,
        R_23ab8_9d1f8a0,R_23ace_9d1ff30,R_23ae4_9d23ce0,R_23afa_95834e8,R_23b04_9583590,R_23b06_9d20860,R_23b08_9d24958,R_23b0a_9d24ca0,R_23a8e_95836e0,R_23a90_9583e18,
        R_23a92_9d25288,R_23a94_9d20908,R_23a96_9d25330,R_23a98_9d22348,R_23a9a_9d253d8,R_23a9c_9d233b0,R_23a9e_9d25528,R_23aa0_9d255d0,R_23aa4_9d23500,R_23aa6_9d25678,
        R_23aa8_9d23a40,R_23aaa_9d24610,R_23aac_9d25880,R_23aae_9d248b0,R_23ab0_9d26258,R_23ab2_9584898,R_23ab4_9d24a00,R_23ab6_9d26450,R_23aba_9d26648,R_23abc_9d26e28,
        R_23abe_9d270c8,R_23ac0_9584c88,R_23ac2_9d24aa8,R_23ac4_9d24d48,R_23ac6_9585270,R_23ac8_9585708,R_23aca_9d27bf0,R_23acc_9d28910,R_23ad0_9d29198,R_23ad2_9d29630,
        R_23ad4_9d24fe8,R_23ad6_95857b0,R_23ad8_9d2a0b0,R_23ada_9585900,R_23adc_9d2a200,R_23ade_9d2a3f8,R_23ae0_9d2a7e8,R_23ae2_9d25138,R_23ae6_9d2ad28,R_23ae8_95860e0,
        R_23aea_9d25480,R_23aec_9d25928,R_23aee_9d25bc8,R_23af0_95864d0,R_23af2_9d25e68,R_23af4_95866c8,R_23af6_9586770,R_23af8_9587688,R_23afc_9d26ed0,R_23afe_9587730,
        R_23b00_9d27aa0,R_23b02_9d2add0,R_23b0c_95877d8,R_23b22_95386e8,R_23b38_95388e0,R_23b4e_9588108,R_23b64_9538ad8,R_23b7a_9d2b118,R_23b84_95881b0,R_23b86_95899f8,
        R_23b88_9589aa0,R_23b8a_9d2b460,R_23b0e_958d268,R_23b10_95390c0,R_23b12_9539168,R_23b14_95394b0,R_23b16_95399f0,R_23b18_9539c90,R_23b1a_953ba18,R_23b1c_953bac0,
        R_23b1e_958d460,R_23b20_9d2b508,R_23b24_953bf58,R_23b26_953c0a8,R_23b28_953c1f8,R_23b2a_953c540,R_23b2c_9d2b5b0,R_23b2e_953c888,R_23b30_953cdc8,R_23b32_958da48,
        R_23b34_9d2b700,R_23b36_953cf18,R_23b3a_958de38,R_23b3c_958e180,R_23b3e_96ddca8,R_23b40_96dddf8,R_23b42_958e570,R_23b44_958e810,R_23b46_96de098,R_23b48_9d285c8,
        R_23b4a_96de3e0,R_23b4c_9d28b08,R_23b50_96de530,R_23b52_958ef48,R_23b54_9d24b50,R_23b56_9d25d18,R_23b58_958ff08,R_23b5a_96e6c60,R_23b5c_96e8160,R_23b5e_96ebc70,
        R_23b60_95903a0,R_23b62_95906e8,R_23b66_96ebdc0,R_23b68_95efb90,R_23b6a_9596d58,R_23b6c_9d2b7a8,R_23b6e_9598c30,R_23b70_95f0220,R_23b72_9598cd8,R_23b74_95f1918,
        R_23b76_9599170,R_23b78_9d28bb0,R_23b7c_95f37f0,R_23b7e_95f41c8,R_23b80_95f4318,R_23b82_95992c0,R_23b8c_9599608,R_23ba2_9599758,R_23bb8_9599800,R_23bce_9599950,
        R_23be4_962f570,R_23bfa_9599b48,R_23c04_959a088,R_23c06_959a130,R_23c08_959a1d8,R_23c0a_962f618,R_23b8e_959a5c8,R_23b90_959a9b8,R_23b92_959ac58,R_23b94_959aef8,
        R_23b96_962f8b8,R_23b98_959afa0,R_23b9a_959b048,R_23b9c_959b0f0,R_23b9e_959b198,R_23ba0_959b240,R_23ba4_959b6d8,R_23ba6_959b828,R_23ba8_959b8d0,R_23baa_959ba20,
        R_23bac_9d28da8,R_23bae_959bac8,R_23bb0_959d268,R_23bb2_959d508,R_23bb4_959dce8,R_23bb6_959e420,R_23bba_9d28fa0,R_23bbc_962f960,R_23bbe_9d298d0,R_23bc0_959e618,
        R_23bc2_959eea0,R_23bc4_959f098,R_23bc6_9d29978,R_23bc8_9d25dc0,R_23bca_959f9c8,R_23bcc_9d29a20,R_23bd0_95a0e20,R_23bd2_9d29b70,R_23bd4_962fb58,R_23bd6_95a0f70,
        R_23bd8_9d29c18,R_23bda_9619ae0,R_23bdc_9619b88,R_23bde_9619d80,R_23be0_9619e28,R_23be2_961a020,R_23be6_961a0c8,R_23be8_961a218,R_23bea_961a4b8,R_23bec_961a800,
        R_23bee_961a8a8,R_23bf0_961a950,R_23bf2_961ad40,R_23bf4_961ade8,R_23bf6_961ae90,R_23bf8_961af38,R_23bfc_9d26060,R_23bfe_961b088,R_23c00_9d29d68,R_23c02_961b1d8,
        R_239cc_95f4af8,R_239ce_962fd50,R_239d0_9558e00,R_239d2_9d261b0,R_239d4_95f52d8,R_239d6_9558ea8,R_239d8_961b670,R_239da_95f5620,R_239dc_961b910,R_239de_9d2b850,
        R_239e0_9d2b9a0,R_239e2_9d29e10,R_239e4_9d2a158,R_239e6_961bb08,R_239e8_961c978,R_239ea_961cd68,R_239ec_9d2baf0,R_239ee_95f5968,R_239f0_95f5ab8,R_239f2_9d2a2a8,
        R_239f4_961ce10,R_239f6_9634e08,R_239f8_9d2bb98,R_239fa_9d2bd90,R_239fc_962fdf8,R_239fe_962fea0,R_23a00_961d200,R_23a02_961d5f0,R_23a04_961d698,R_23a06_962fff0,
        R_23a08_961d740,R_23a0a_961d938,R_23c24_9d2a698,R_23c26_9d2c420,R_23c28_962ac98,R_23c2a_9d2c4c8,R_23c2c_9d2c570,R_23c2e_95f63e8,R_23c30_9d2a890,R_23c32_962ad40,
        R_23c22_9d2aa88,R_23c34_9d2c810,R_23c36_9d2ab30,R_23c38_9d2c8b8,R_23c3a_9d2cab0,R_23c20_9635e70,R_23c52_962b868,R_23c54_9d2af20,R_23c56_9d2b310,R_23774_9630098,
        R_2378a_962b9b8,R_237a0_9d2cd50,R_237b6_962bb08,R_237cc_9d2cff0,R_237e2_9d2d098,R_237ec_9d2d140,R_237ee_9d2d290,R_237f0_962c240,R_237f2_9559688,R_23776_96301e8,
        R_23778_9d2d7d0,R_2377a_962c2e8,R_2377c_9d2d878,R_2377e_962ce10,R_23780_9d2d920,R_23782_962d938,R_23784_962e5b0,R_23786_9d2d9c8,R_23788_9d2dc68,R_2378c_9d2dd10,
        R_2378e_9d2ddb8,R_23790_9d2e100,R_23792_9d2e1a8,R_23794_9d2f0c0,R_23796_9630290,R_23798_96303e0,R_2379a_9d2f210,R_2379c_9d2f7f8,R_2379e_9630728,R_237a2_96307d0,
        R_237a4_9d2fb40,R_237a6_9d301d0,R_237a8_9559bc8,R_237aa_9630140,R_237ac_96312f8,R_237ae_9d30710,R_237b0_9630b18,R_237b2_9630c68,R_237b4_9d309b0,R_237b8_9630d10,
        R_237ba_9630fb0,R_237bc_9631100,R_237be_9d30a58,R_237c0_9d30da0,R_237c2_96311a8,R_237c4_96313a0,R_237c6_96318e0,R_237c8_9631a30,R_237ca_9d30e48,R_237ce_9d31190,
        R_237d0_9631b80,R_237d2_9d31f58,R_237d4_9631448,R_237d6_9631790,R_237d8_9d323f0,R_237da_9631ad8,R_237dc_9d32540,R_237de_9632018,R_237e0_9631cd0,R_237e4_9632210,
        R_237e6_9d32690,R_237e8_96322b8,R_237ea_9d32888,R_237f4_9631e20,R_2380a_9d329d8,R_23820_9d32a80,R_23836_9d32f18,R_2384c_9d2b3b8,R_23862_9631ec8,R_2386c_9632360,
        R_2386e_9632a98,R_23870_9d32fc0,R_23872_9632408,R_237f6_9632600,R_237f8_9d33500,R_237fa_96326a8,R_237fc_9d33650,R_237fe_9d336f8,R_23800_9d33a40,R_23802_9632750,
        R_23804_96328a0,R_23806_9d340d0,R_23808_9632948,R_2380c_9d2b658,R_2380e_9d34418,R_23810_9d34760,R_23812_9d34fe8,R_23814_9632de0,R_23816_9632e88,R_23818_9d35720,
        R_2381a_9d2bc40,R_2381c_b805670,R_2381e_b805868,R_23822_9633080,R_23824_b8060f0,R_23826_9633128,R_23828_9633b00,R_2382a_9632b40,R_2382c_9634190,R_2382e_9638720,
        R_23830_9d2c180,R_23832_96389c0,R_23834_9638a68,R_23838_9d15880,R_2383a_b806198,R_2383c_9d2c768,R_2383e_9d16a38,R_23840_9d2ca08,R_23842_b806240,R_23844_9d17170,
        R_23846_9d17c98,R_23848_b8062e8,R_2384a_b806390,R_2384e_9d2cca8,R_23850_9d17fe0,R_23852_9d18328,R_23854_9d2d1e8,R_23856_9d1fd38,R_23858_b8064e0,R_2385a_9d2d3e0,
        R_2385c_9d220a8,R_2385e_9535d90,R_23860_b806588,R_23864_9d25720,R_23866_b8066d8,R_23868_b806780,R_2386a_9d2d530,R_23874_95f7840,R_2388a_95f7e28,R_238a0_9d28e50,
        R_238b6_95f8170,R_238cc_95fcd90,R_238e2_95fda08,R_238ec_95fdb58,R_238ee_95fdca8,R_238f0_95fdd50,R_238f2_9d2d728,R_23876_95ff6e8,R_23878_9535e38,R_2387a_9633668,
        R_2387c_9f4ddd0,R_2387e_9f51b80,R_23880_9f51e20,R_23882_9d29ac8,R_23884_9f53278,R_23886_9f53320,R_23888_9f54580,R_2388c_9f54778,R_2388e_9d2dbc0,R_23890_9d2e250,
        R_23892_9f548c8,R_23894_9f54970,R_23896_9f54c10,R_23898_9f55348,R_2389a_9f55498,R_2389c_9d2a740,R_2389e_9d2e3a0,R_238a2_9d2b070,R_238a4_9633710,R_238a6_9f55b28,
        R_238a8_9f56260,R_238aa_9f56500,R_238ac_9f5baf8,R_238ae_9ee9d78,R_238b0_9d2ba48,R_238b2_9d2bce8,R_238b4_9eea0c0,R_238b8_9eeb518,R_238ba_9eedf18,R_238bc_9eee6f8,
        R_238be_9ef2010,R_238c0_9537530,R_238c2_9ef2208,R_238c4_9ef3660,R_238c6_9ef3858,R_238c8_9633860,R_238ca_9ef3a50,R_238ce_9ef3af8,R_238d0_9ef3ba0,R_238d2_9ef3c48,
        R_238d4_9ef4620,R_238d6_9d2c2d0,R_238d8_9ef4770,R_238da_9d2cb58,R_238dc_9ef4ab8,R_238de_9ef4c08,R_238e0_9ef4ff8,R_238e4_9ef5148,R_238e6_9ef51f0,R_238e8_9d2cf48,
        R_238ea_9ef53e8,R_238f4_9d2e4f0,R_2390a_96339b0,R_23920_9633c50,R_23936_9d266f0,R_2394c_9d2e838,R_23962_9d2ecd0,R_2396c_9d2ed78,R_2396e_9d2f018,R_23970_9d2f168,
        R_23972_b8068d0,R_238f6_9d2f2b8,R_238f8_9d2f9f0,R_238fa_9d2fde0,R_238fc_9633f98,R_238fe_b806a20,R_23900_96340e8,R_23902_9d30320,R_23904_9634580,R_23906_9d305c0,
        R_23908_9634b68,R_2390c_9d30ba8,R_2390e_9d30c50,R_23910_b806ac8,R_23912_9d32000,R_23914_b806b70,R_23916_9d320a8,R_23918_9634c10,R_2391a_9d32150,R_2391c_9634cb8,
        R_2391e_9d32498,R_23922_9d32738,R_23924_9d327e0,R_23926_9d32b28,R_23928_9d32bd0,R_2392a_9635348,R_2392c_9635690,R_2392e_9d32c78,R_23930_9d32d20,R_23932_9635a80,
        R_23934_9d32dc8,R_23938_9d331b8,R_2393a_9d2d488,R_2393c_9d333b0,R_2393e_9d335a8,R_23940_9d337a0,R_23942_9635b28,R_23944_9d2d5d8,R_23946_9d338f0,R_23948_9635bd0,
        R_2394a_9d33998,R_2394e_9d33ae8,R_23950_9d33b90,R_23952_9636110,R_23954_9d33ce0,R_23956_b806c18,R_23958_9d33ed8,R_2395a_9d33f80,R_2395c_9636308,R_2395e_b806cc0,
        R_23960_9d34028,R_23964_9d34178,R_23966_9d2db18,R_23968_96365a8,R_2396a_9636848,R_23734_96368f0,R_23736_9636998,R_23738_9636a40,R_2373a_b7dc0c0,R_2373c_9636b90,
        R_2373e_9636c38,R_23740_b7dc168,R_23742_b806d68,R_23744_b806e10,R_23746_9636ed8,R_23748_b806eb8,R_2374a_9637028,R_2374c_b806f60,R_2374e_b8070b0,R_23750_9d33308,
        R_23752_b807158,R_23754_9ef5880,R_23756_9d26798,R_23758_9d342c8,R_2375a_9ef5928,R_2375c_96c2b20,R_2375e_9d31820,R_23760_9d31970,R_23762_9637178,R_23764_9d26840,
        R_23766_96372c8,R_23768_9d268e8,R_2376a_9d26a38,R_2376c_9d26ae0,R_2376e_9637370,R_23770_9d26b88,R_23772_9637418,R_2398c_96c2fb8,R_2398e_9559c70,R_23990_96c35a0,
        R_23992_96e8010,R_23994_955a300,R_23996_955a450,R_23998_9d34ca0,R_2399a_96c3840,R_2398a_9d34d48,R_2399c_96c3a38,R_2399e_96c3d80,R_239a0_955a840,R_239a2_96c59b8,
        R_23988_96eaf50,R_239ba_96ca728,R_239bc_955b8a8,R_239be_b7db6e8,R_234dc_b8085b0,R_234f2_b80b988,R_23508_b808658,R_2351e_b808700,R_23534_b8087a8,R_2354a_b8088f8,
        R_23554_b80ba30,R_23556_b80bb80,R_23558_b80bec8,R_2355a_b80bf70,R_234de_b8089a0,R_234e0_b808a48,R_234e2_b809768,R_234e4_b809df8,R_234e6_b80c2b8,R_234e8_b80e040,
        R_234ea_b80e580,R_234ec_b80c600,R_234ee_b80f0a8,R_234f0_b80fd20,R_234f4_b80c750,R_234f6_b80ffc0,R_234f8_b7ddf98,R_234fa_b80c7f8,R_234fc_b7de0e8,R_234fe_b7de388,
        R_23500_b7de430,R_23502_b80c9f0,R_23504_b7de580,R_23506_b80ca98,R_2350a_b7de820,R_2350c_b7dea18,R_2350e_b7dee08,R_23510_b80cc90,R_23512_b80cd38,R_23514_b7df1f8,
        R_23516_b80ce88,R_23518_b7df348,R_2351a_b7df540,R_2351c_b80cf30,R_23520_b7dfc78,R_23522_b80d080,R_23524_b80d278,R_23526_b7dff18,R_23528_b80d320,R_2352a_b7e0068,
        R_2352c_b80d5c0,R_2352e_b7e01b8,R_23530_b80d668,R_23532_b7e0458,R_23536_b7e05a8,R_23538_b80d7b8,R_2353a_b80de48,R_2353c_b7e0998,R_2353e_b7e0b90,R_23540_b7e1178,
        R_23542_b80e430,R_23544_b80e628,R_23546_b80e778,R_23548_b7e1568,R_2354c_b80e970,R_2354e_b7e16b8,R_23550_b80eb68,R_23552_b7e1808,R_2355c_b7e18b0,R_23572_b805c58,
        R_23588_b7e1958,R_2359e_b80ed60,R_235b4_95ad7d8,R_235ca_b806438,R_235d4_b7e1a00,R_235d6_b80f000,R_235d8_b7e1bf8,R_235da_b7e1ca0,R_2355e_b7e1e98,R_23560_95ad9d0,
        R_23562_b7e1f40,R_23564_95adb20,R_23566_b7e1fe8,R_23568_b80f3f0,R_2356a_b80f5e8,R_2356c_b806630,R_2356e_b7e2090,R_23570_b80f690,R_23574_b7e2138,R_23576_b7e21e0,
        R_23578_b7e23d8,R_2357a_b7e2720,R_2357c_b7e2870,R_2357e_b7e29c0,R_23580_b806828,R_23582_b7e2a68,R_23584_b7e2c60,R_23586_b7e2f00,R_2358a_b80f7e0,R_2358c_96cb8e0,
        R_2358e_b7e2fa8,R_23590_b7e30f8,R_23592_b806978,R_23594_b807008,R_23596_b7e32f0,R_23598_b80fb28,R_2359a_b7e3398,R_2359c_b807698,R_235a0_b7e34e8,R_235a2_96cbb80,
        R_235a4_b80fbd0,R_235a6_96cc018,R_235a8_95adf10,R_235aa_b7e36e0,R_235ac_b807890,R_235ae_b7e3788,R_235b0_b7e38d8,R_235b2_b7e3ad0,R_235b6_b7e3cc8,R_235b8_b7e3f68,
        R_235ba_b807f20,R_235bc_b807fc8,R_235be_b8101b8,R_235c0_b7e40b8,R_235c2_b7e4208,R_235c4_b8105a8,R_235c6_b810650,R_235c8_96cc210,R_235cc_b7e42b0,R_235ce_b7e4400,
        R_235d0_b7e4550,R_235d2_b7e45f8,R_235dc_b8106f8,R_235f2_b7e46a0,R_23608_b808118,R_2361e_b7e47f0,R_23634_b7e49e8,R_2364a_b7dd860,R_23654_95ae060,R_23656_b7dd908,
        R_23658_b7ddda0,R_2365a_b7dde48,R_235de_9637b50,R_235e0_95ae1b0,R_235e2_b7ddef0,R_235e4_b7de238,R_235e6_b7e4b38,R_235e8_9637fe8,R_235ea_b7de2e0,R_235ec_b808310,
        R_235ee_9638138,R_235f0_96381e0,R_235f4_b7e4d30,R_235f6_96383d8,R_235f8_b7de6d0,R_235fa_9638480,R_235fc_b7de8c8,R_235fe_9638528,R_23600_96385d0,R_23602_b7de970,
        R_23604_b7deac0,R_23606_9638678,R_2360a_96387c8;

wire \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 ,
         \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 ,
         \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 ,
         \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 ,
         \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 ,
         \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 ,
         \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 ,
         \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 ,
         \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 ,
         \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 ,
         \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 ,
         \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 ,
         \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 ,
         \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 ,
         \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 ,
         \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 ,
         \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 ,
         \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 ,
         \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 ,
         \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 ,
         \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 ,
         \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 ,
         \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 ,
         \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 ,
         \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 ,
         \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 ,
         \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 ,
         \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 ,
         \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 ,
         \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 ,
         \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 ,
         \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 ,
         \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 ,
         \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 ,
         \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 ,
         \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 ,
         \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 ,
         \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 ,
         \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 ,
         \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 ,
         \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 ,
         \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 ,
         \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 ,
         \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 ,
         \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 ,
         \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 ,
         \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 ,
         \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 ,
         \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 ,
         \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 ,
         \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 ,
         \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 ,
         \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 ,
         \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 ,
         \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 ,
         \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 ,
         \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 ,
         \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 ,
         \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 ,
         \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 ,
         \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 ,
         \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 ,
         \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 ,
         \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 ,
         \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 ,
         \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 ,
         \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 ,
         \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 ,
         \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 ,
         \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 ,
         \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 ,
         \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 ,
         \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 ,
         \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 ,
         \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 ,
         \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 ,
         \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 ,
         \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 ,
         \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 ,
         \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 ,
         \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 ,
         \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 ,
         \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 ,
         \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 ,
         \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 ,
         \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 ,
         \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 ,
         \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 ,
         \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 ,
         \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 ,
         \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 ,
         \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 ,
         \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 ,
         \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 ,
         \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 ,
         \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 ,
         \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 ,
         \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 ,
         \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 ,
         \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 ,
         \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 ,
         \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 ,
         \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 ,
         \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 ,
         \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 ,
         \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 ,
         \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 ,
         \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 ,
         \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 ,
         \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 ,
         \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 ,
         \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 ,
         \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 ,
         \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 ,
         \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 ,
         \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 ,
         \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 ,
         \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 ,
         \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 , \4473 , \4474 ,
         \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 ,
         \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 ,
         \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 ,
         \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514 ,
         \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 ,
         \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 ,
         \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 ,
         \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 , \4553 , \4554 ,
         \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 ,
         \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 ,
         \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 ,
         \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 , \4593 , \4594 ,
         \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 ,
         \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 ,
         \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 ,
         \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 , \4633 , \4634 ,
         \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 ,
         \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 ,
         \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 ,
         \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 , \4673 , \4674 ,
         \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 , \4683 , \4684 ,
         \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 , \4693 , \4694 ,
         \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 , \4703 , \4704 ,
         \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 , \4713 , \4714 ,
         \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 ,
         \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 ,
         \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 ,
         \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 ,
         \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 , \4763 , \4764 ,
         \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 , \4773 , \4774 ,
         \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 , \4783 , \4784 ,
         \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 , \4793 , \4794 ,
         \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 , \4803 , \4804 ,
         \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 , \4813 , \4814 ,
         \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 , \4823 , \4824 ,
         \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 , \4833 , \4834 ,
         \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 , \4843 , \4844 ,
         \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 , \4853 , \4854 ,
         \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 , \4863 , \4864 ,
         \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 , \4873 , \4874 ,
         \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 , \4883 , \4884 ,
         \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 , \4893 , \4894 ,
         \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 , \4903 , \4904 ,
         \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 , \4913 , \4914 ,
         \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 , \4923 , \4924 ,
         \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 , \4933 , \4934 ,
         \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 ,
         \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 , \4953 , \4954 ,
         \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 , \4963 , \4964 ,
         \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 , \4973 , \4974 ,
         \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 , \4983 , \4984 ,
         \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 ,
         \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 ,
         \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 , \5013 , \5014 ,
         \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 ,
         \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 , \5033 , \5034 ,
         \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 ,
         \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 ,
         \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 , \5063 , \5064 ,
         \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 ,
         \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 ,
         \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 ,
         \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 ,
         \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 , \5113 , \5114 ,
         \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 ,
         \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 ,
         \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 ,
         \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 ,
         \5155 , \5156 , \5157_N$2 , \5158_N$5 , \5159_N$7 , \5160_N$8 , \5161_N$9 , \5162_N$10 , \5163_N$11 , \5164_N$12 ,
         \5165_N$13 , \5166_N$14 , \5167_N$15 , \5168_N$16 , \5169_N$17 , \5170_N$19 , \5171_N$22 , \5172_N$24 , \5173_N$25 , \5174_N$26 ,
         \5175_N$27 , \5176_N$28 , \5177_N$29 , \5178_N$30 , \5179_N$31 , \5180_N$32 , \5181_N$33 , \5182_N$35 , \5183_N$38 , \5184_N$40 ,
         \5185_N$41 , \5186_N$42 , \5187_N$43 , \5188_N$44 , \5189_N$45 , \5190_N$46 , \5191_N$47 , \5192_N$48 , \5193_N$49 , \5194_N$50 ,
         \5195_N$53 , \5196_N$56 , \5197_N$58 , \5198_N$59 , \5199_N$60 , \5200_N$61 , \5201_N$62 , \5202_N$63 , \5203_N$64 , \5204_N$65 ,
         \5205_N$66 , \5206_N$67 , \5207_N$68 , \5208_N$69 , \5209_N$70 , \5210_N$71 , \5211_N$72 , \5212_N$73 , \5213_N$74 , \5214_N$75 ,
         \5215_N$76 , \5216_N$77 , \5217_N$78 , \5218_N$79 , \5219_N$80 , \5220_N$81 , \5221_N$82 , \5222_N$83 , \5223_N$84 , \5224_N$85 ,
         \5225_N$86 , \5226_N$87 , \5227_N$88 , \5228_N$89 , \5229_N$90 , \5230_N$91 , \5231_N$92 , \5232_N$93 , \5233_N$94 , \5234_N$95 ,
         \5235_N$96 , \5236_N$97 , \5237_N$98 , \5238_N$99 , \5239_N$100 , \5240_N$101 , \5241_N$102 , \5242_N$103 , \5243_N$104 , \5244_N$105 ,
         \5245_N$106 , \5246_N$107 , \5247_N$108 , \5248_N$109 , \5249_N$110 , \5250_N$111 , \5251_N$112 , \5252_N$113 , \5253_N$114 , \5254_N$115 ,
         \5255_N$116 , \5256_N$117 , \5257_N$118 , \5258_N$119 , \5259_N$120 , \5260_N$121 , \5261_N$122 , \5262_N$123 , \5263_N$124 , \5264_N$125 ,
         \5265_N$126 , \5266_N$127 , \5267_N$128 , \5268_N$129 , \5269_N$130 , \5270_N$131 , \5271_N$132 , \5272_N$133 , \5273_N$134 , \5274_N$135 ,
         \5275_N$136 , \5276_N$137 , \5277_N$138 , \5278_N$139 , \5279_N$140 , \5280_N$141 , \5281_N$142 , \5282_N$143 , \5283_N$144 , \5284_N$145 ,
         \5285_N$146 , \5286_N$147 , \5287_N$148 , \5288_N$149 , \5289_N$150 , \5290_N$151 , \5291_N$152 , \5292_N$153 , \5293_N$154 , \5294_N$155 ,
         \5295_N$156 , \5296_N$157 , \5297_N$158 , \5298_N$159 , \5299_N$160 , \5300_N$161 , \5301_N$162 , \5302_N$163 , \5303_N$164 , \5304_N$165 ,
         \5305_N$166 , \5306_N$167 , \5307_N$168 , \5308_N$169 , \5309_N$170 , \5310_N$171 , \5311_N$172 , \5312_N$173 , \5313_N$174 , \5314_N$175 ,
         \5315_N$176 , \5316_N$177 , \5317_N$178 , \5318_N$179 , \5319_N$180 , \5320_N$181 , \5321_N$182 , \5322_N$183 , \5323_N$184 , \5324_N$185 ,
         \5325_N$186 , \5326_N$187 , \5327_N$188 , \5328_N$189 , \5329_N$190 , \5330_N$191 , \5331_N$192 , \5332_N$193 , \5333_N$194 , \5334_N$195 ,
         \5335_N$196 , \5336_N$197 , \5337_N$198 , \5338_N$199 , \5339_N$200 , \5340_N$201 , \5341_N$202 , \5342_N$203 , \5343_N$204 , \5344_N$205 ,
         \5345_N$206 , \5346_N$207 , \5347_N$208 , \5348_N$209 , \5349_N$210 , \5350_N$211 , \5351_N$212 , \5352_N$213 , \5353_N$214 , \5354_N$215 ,
         \5355_N$216 , \5356_N$217 , \5357_N$218 , \5358_N$219 , \5359_N$220 , \5360_N$221 , \5361_N$222 , \5362_N$223 , \5363_N$224 , \5364_N$225 ,
         \5365_N$226 , \5366_N$227 , \5367_N$228 , \5368_N$229 , \5369_N$230 , \5370_N$231 , \5371_N$232 , \5372_N$233 , \5373_N$234 , \5374_N$235 ,
         \5375_N$236 , \5376_N$237 , \5377_N$238 , \5378_N$239 , \5379_N$240 , \5380_N$241 , \5381_N$242 , \5382_N$243 , \5383_N$244 , \5384_N$245 ,
         \5385_N$246 , \5386_N$247 , \5387_N$248 , \5388_N$249 , \5389_N$250 , \5390_N$251 , \5391_N$252 , \5392_N$253 , \5393_N$254 , \5394_N$255 ,
         \5395_N$256 , \5396_N$257 , \5397_N$258 , \5398_N$259 , \5399_N$260 , \5400_N$261 , \5401_N$262 , \5402_N$263 , \5403_N$264 , \5404_N$265 ,
         \5405_N$266 , \5406_N$267 , \5407_N$268 , \5408_N$269 , \5409_N$270 , \5410_N$271 , \5411_N$272 , \5412_N$273 , \5413_N$274 , \5414_N$275 ,
         \5415_N$276 , \5416_N$277 , \5417_N$278 , \5418_N$279 , \5419_N$280 , \5420_N$281 , \5421_N$282 , \5422_N$283 , \5423_N$284 , \5424_N$285 ,
         \5425_N$286 , \5426_N$287 , \5427_N$288 , \5428_N$289 , \5429_N$290 , \5430_N$291 , \5431_N$292 , \5432_N$293 , \5433_N$294 , \5434_N$295 ,
         \5435_N$296 , \5436_N$297 , \5437_N$298 , \5438_N$299 , \5439_N$300 , \5440_N$301 , \5441_N$302 , \5442_N$303 , \5443_N$304 , \5444_N$305 ,
         \5445_N$306 , \5446_N$307 , \5447_N$308 , \5448_N$309 , \5449_N$310 , \5450_N$311 , \5451_N$312 , \5452_N$313 , \5453_N$314 , \5454_N$315 ,
         \5455_N$316 , \5456_N$317 , \5457_N$318 , \5458_N$319 , \5459_N$320 , \5460_N$321 , \5461_N$322 , \5462_N$323 , \5463_N$324 , \5464_N$325 ,
         \5465_N$326 , \5466_N$327 , \5467_N$328 , \5468_N$329 , \5469_N$330 , \5470_N$331 , \5471_N$332 , \5472_N$333 , \5473_N$334 , \5474_N$335 ,
         \5475_N$336 , \5476_N$337 , \5477_N$338 , \5478_N$339 , \5479_N$340 , \5480_N$341 , \5481_N$342 , \5482_N$343 , \5483_N$344 , \5484_N$345 ,
         \5485_N$346 , \5486_N$347 , \5487_N$348 , \5488_N$349 , \5489_N$350 , \5490_N$351 , \5491_N$352 , \5492_N$353 , \5493_N$354 , \5494_N$355 ,
         \5495_N$356 , \5496_N$357 , \5497_N$358 , \5498_N$359 , \5499_N$360 , \5500_N$361 , \5501_N$362 , \5502_N$363 , \5503_N$364 , \5504_N$365 ,
         \5505_N$366 , \5506_N$367 , \5507_N$368 , \5508_N$369 , \5509_N$370 , \5510_N$371 , \5511_N$372 , \5512_N$373 , \5513_N$374 , \5514_N$375 ,
         \5515_N$376 , \5516_N$377 , \5517_N$378 , \5518_N$379 , \5519_N$380 , \5520_N$381 , \5521_N$382 , \5522_N$383 , \5523_N$384 , \5524_N$385 ,
         \5525_N$386 , \5526_N$387 , \5527_N$388 , \5528_N$389 , \5529_N$390 , \5530_N$391 , \5531_N$392 , \5532_N$393 , \5533_N$394 , \5534_N$395 ,
         \5535_N$396 , \5536_N$397 , \5537_N$398 , \5538_N$399 , \5539_N$400 , \5540_N$401 , \5541_N$402 , \5542_N$403 , \5543_N$404 , \5544_N$405 ,
         \5545_N$406 , \5546_N$407 , \5547_N$408 , \5548_N$409 , \5549_N$410 , \5550_N$411 , \5551_N$412 , \5552_N$413 , \5553_N$414 , \5554_N$415 ,
         \5555_N$416 , \5556_N$417 , \5557_N$418 , \5558_N$419 , \5559_N$420 , \5560_N$421 , \5561_N$422 , \5562_N$423 , \5563_N$424 , \5564_N$425 ,
         \5565_N$426 , \5566_N$427 , \5567_N$428 , \5568_N$429 , \5569_N$430 , \5570_N$431 , \5571_N$432 , \5572_N$433 , \5573_N$434 , \5574_N$435 ,
         \5575_N$436 , \5576_N$437 , \5577_N$438 , \5578_N$439 , \5579_N$440 , \5580_N$441 , \5581_N$442 , \5582_N$443 , \5583_N$444 , \5584_N$445 ,
         \5585_N$446 , \5586_N$447 , \5587_N$448 , \5588_N$449 , \5589_N$450 , \5590_N$451 , \5591_N$452 , \5592_N$453 , \5593_N$454 , \5594_N$455 ,
         \5595_N$456 , \5596_N$457 , \5597_N$458 , \5598_N$459 , \5599_N$460 , \5600_N$461 , \5601_N$462 , \5602_N$463 , \5603_N$464 , \5604_N$465 ,
         \5605_N$466 , \5606_N$467 , \5607_N$468 , \5608_N$469 , \5609_N$470 , \5610_N$471 , \5611_N$472 , \5612_N$473 , \5613_N$474 , \5614_N$475 ,
         \5615_N$476 , \5616_N$477 , \5617_N$478 , \5618_N$479 , \5619_N$480 , \5620_N$481 , \5621_N$482 , \5622_N$483 , \5623_N$484 , \5624_N$485 ,
         \5625_N$486 , \5626_N$487 , \5627_N$488 , \5628_N$489 , \5629_N$490 , \5630_N$491 , \5631_N$492 , \5632_N$493 , \5633_N$494 , \5634_N$495 ,
         \5635_N$496 , \5636_N$497 , \5637_N$498 , \5638_N$499 , \5639_N$500 , \5640_N$501 , \5641_N$502 , \5642_N$503 , \5643_N$504 , \5644_N$505 ,
         \5645_N$506 , \5646_N$507 , \5647_N$508 , \5648_N$509 , \5649_N$510 , \5650_N$511 , \5651_N$512 , \5652_N$513 , \5653_N$514 , \5654_N$515 ,
         \5655_N$516 , \5656_N$517 , \5657_N$518 , \5658_N$519 , \5659_N$520 , \5660_N$521 , \5661_N$522 , \5662_N$523 , \5663_N$524 , \5664_N$525 ,
         \5665_N$526 , \5666_N$527 , \5667_N$528 , \5668_N$529 , \5669_N$530 , \5670_N$531 , \5671_N$532 , \5672_N$533 , \5673_N$534 , \5674_N$535 ,
         \5675_N$536 , \5676_N$537 , \5677_N$538 , \5678_N$539 , \5679_N$540 , \5680_N$541 , \5681_N$542 , \5682_N$543 , \5683_N$544 , \5684_N$545 ,
         \5685_N$546 , \5686_N$547 , \5687_N$548 , \5688_N$549 , \5689_N$550 , \5690_N$551 , \5691_N$552 , \5692_N$553 , \5693_N$554 , \5694_N$555 ,
         \5695_N$556 , \5696_N$557 , \5697_N$558 , \5698_N$559 , \5699_N$560 , \5700_N$561 , \5701_N$562 , \5702_N$563 , \5703_N$564 , \5704_N$565 ,
         \5705_N$566 , \5706_N$567 , \5707_N$568 , \5708_N$569 , \5709_N$570 , \5710_N$571 , \5711_N$572 , \5712_N$573 , \5713_N$574 , \5714_N$575 ,
         \5715_N$576 , \5716_N$577 , \5717_N$578 , \5718_N$579 , \5719_N$580 , \5720_N$581 , \5721_N$582 , \5722_N$583 , \5723_N$584 , \5724_N$585 ,
         \5725_N$586 , \5726_N$587 , \5727_N$588 , \5728_N$589 , \5729_N$590 , \5730_N$591 , \5731_N$592 , \5732_N$593 , \5733_N$594 , \5734_N$595 ,
         \5735_N$596 , \5736_N$597 , \5737_N$598 , \5738_N$599 , \5739_N$600 , \5740_N$601 , \5741_N$602 , \5742_N$603 , \5743_N$604 , \5744_N$605 ,
         \5745_N$606 , \5746_N$607 , \5747_N$608 , \5748_N$609 , \5749_N$610 , \5750_N$611 , \5751_N$612 , \5752_N$613 , \5753_N$614 , \5754_N$615 ,
         \5755_N$616 , \5756_N$617 , \5757_N$618 , \5758_N$619 , \5759_N$620 , \5760_N$621 , \5761_N$622 , \5762_N$623 , \5763_N$624 , \5764_N$625 ,
         \5765_N$626 , \5766_N$627 , \5767_N$628 , \5768_N$629 , \5769_N$630 , \5770_N$631 , \5771_N$632 , \5772_N$633 , \5773_N$634 , \5774_N$635 ,
         \5775_N$636 , \5776_N$637 , \5777_N$638 , \5778_N$639 , \5779_N$640 , \5780_N$641 , \5781_N$642 , \5782_N$643 , \5783_N$644 , \5784_N$645 ,
         \5785_N$646 , \5786_N$647 , \5787_N$648 , \5788_N$649 , \5789_N$650 , \5790_N$651 , \5791_N$652 , \5792_N$653 , \5793_N$654 , \5794_N$655 ,
         \5795_N$656 , \5796_N$657 , \5797_N$658 , \5798_N$659 , \5799_N$660 , \5800_N$661 , \5801_N$662 , \5802_N$663 , \5803_N$664 , \5804_N$665 ,
         \5805_N$666 , \5806_N$667 , \5807_N$668 , \5808_N$669 , \5809_N$670 , \5810_N$671 , \5811_N$672 , \5812_N$673 , \5813_N$674 , \5814_N$675 ,
         \5815_N$676 , \5816_N$677 , \5817_N$678 , \5818_N$679 , \5819_N$680 , \5820_N$681 , \5821_N$682 , \5822_N$683 , \5823_N$684 , \5824_N$685 ,
         \5825_N$686 , \5826_N$687 , \5827_N$688 , \5828_N$689 , \5829_N$690 , \5830_N$691 , \5831_N$692 , \5832_N$693 , \5833_N$694 , \5834_N$695 ,
         \5835_N$696 , \5836_N$697 , \5837_N$698 , \5838_N$699 , \5839_N$700 , \5840_N$701 , \5841_N$702 , \5842_N$703 , \5843_N$704 , \5844_N$705 ,
         \5845_N$706 , \5846_N$707 , \5847_N$708 , \5848_N$709 , \5849_N$710 , \5850_N$711 , \5851_N$712 , \5852_N$713 , \5853_N$714 , \5854_N$715 ,
         \5855_N$716 , \5856_N$717 , \5857_N$718 , \5858_N$719 , \5859_N$720 , \5860_N$721 , \5861_N$722 , \5862_N$723 , \5863_N$724 , \5864_N$725 ,
         \5865_N$726 , \5866_N$727 , \5867_N$728 , \5868_N$729 , \5869_N$730 , \5870_N$731 , \5871_N$732 , \5872_N$733 , \5873_N$734 , \5874_N$735 ,
         \5875_N$736 , \5876_N$737 , \5877_N$738 , \5878_N$739 , \5879_N$740 , \5880_N$741 , \5881_N$742 , \5882_N$743 , \5883_N$744 , \5884_N$745 ,
         \5885_N$746 , \5886_N$747 , \5887_N$748 , \5888_N$749 , \5889_N$750 , \5890_N$751 , \5891_N$752 , \5892_N$753 , \5893_N$754 , \5894_N$755 ,
         \5895_N$756 , \5896_N$757 , \5897_N$758 , \5898_N$759 , \5899_N$760 , \5900_N$761 , \5901_N$762 , \5902_N$763 , \5903_N$764 , \5904_N$765 ,
         \5905_N$766 , \5906_N$767 , \5907_N$768 , \5908_N$769 , \5909_N$770 , \5910_N$771 , \5911_N$772 , \5912_N$773 , \5913_N$774 , \5914_N$775 ,
         \5915_N$776 , \5916_N$777 , \5917_N$778 , \5918_N$779 , \5919_N$780 , \5920_N$781 , \5921_N$782 , \5922_N$783 , \5923_N$784 , \5924_N$785 ,
         \5925_N$786 , \5926_N$787 , \5927_N$788 , \5928_N$789 , \5929_N$790 , \5930_N$791 , \5931_N$792 , \5932_N$793 , \5933_N$794 , \5934_N$795 ,
         \5935_N$796 , \5936_N$797 , \5937_N$798 , \5938_N$799 , \5939_N$800 , \5940_N$801 , \5941_N$802 , \5942_N$803 , \5943_N$804 , \5944_N$805 ,
         \5945_N$806 , \5946_N$807 , \5947_N$808 , \5948_N$809 , \5949_N$810 , \5950_N$811 , \5951_N$812 , \5952_N$813 , \5953_N$814 , \5954_N$815 ,
         \5955_N$816 , \5956_N$817 , \5957_N$818 , \5958_N$819 , \5959_N$820 , \5960_N$821 , \5961_N$822 , \5962_N$823 , \5963_N$824 , \5964_N$825 ,
         \5965_N$826 , \5966_N$827 , \5967_N$828 , \5968_N$829 , \5969_N$830 , \5970_N$831 , \5971_N$832 , \5972_N$833 , \5973_N$834 , \5974_N$835 ,
         \5975_N$836 , \5976_N$837 , \5977_N$838 , \5978_N$839 , \5979_N$840 , \5980_N$841 , \5981_N$842 , \5982_N$843 , \5983_N$844 , \5984_N$845 ,
         \5985_N$846 , \5986_N$847 , \5987_N$848 , \5988_N$849 , \5989_N$850 , \5990_N$851 , \5991_N$852 , \5992_N$853 , \5993_N$854 , \5994_N$855 ,
         \5995_N$856 , \5996_N$857 , \5997_N$858 , \5998_N$859 , \5999_N$860 , \6000_N$861 , \6001_N$862 , \6002_N$863 , \6003_N$864 , \6004_N$865 ,
         \6005_N$866 , \6006_N$867 , \6007_N$868 , \6008_N$869 , \6009_N$870 , \6010_N$871 , \6011_N$872 , \6012_N$873 , \6013_N$874 , \6014_N$875 ,
         \6015_N$876 , \6016_N$877 , \6017_N$878 , \6018_N$879 , \6019_N$880 , \6020_N$881 , \6021_N$882 , \6022_N$883 , \6023_N$884 , \6024_N$885 ,
         \6025_N$886 , \6026_N$887 , \6027_N$888 , \6028_N$889 , \6029_N$890 , \6030_N$891 , \6031_N$892 , \6032_N$893 , \6033_N$894 , \6034_N$895 ,
         \6035_N$896 , \6036_N$897 , \6037_N$898 , \6038_N$899 , \6039_N$900 , \6040_N$901 , \6041_N$902 , \6042_N$903 , \6043_N$904 , \6044_N$905 ,
         \6045_N$906 , \6046_N$907 , \6047_N$908 , \6048_N$909 , \6049_N$910 , \6050_N$911 , \6051_N$912 , \6052_N$913 , \6053_N$914 , \6054_N$915 ,
         \6055_N$916 , \6056_N$917 , \6057_N$918 , \6058_N$919 , \6059_N$920 , \6060_N$921 , \6061_N$922 , \6062_N$923 , \6063_N$924 , \6064_N$925 ,
         \6065_N$926 , \6066_N$927 , \6067_N$928 , \6068_N$929 , \6069_N$930 , \6070_N$931 , \6071_N$932 , \6072_N$933 , \6073_N$934 , \6074_N$935 ,
         \6075_N$936 , \6076_N$937 , \6077_N$938 , \6078_N$939 , \6079_N$940 , \6080_N$941 , \6081_N$942 , \6082_N$943 , \6083_N$944 , \6084_N$945 ,
         \6085_N$946 , \6086_N$947 , \6087_N$948 , \6088_N$949 , \6089_N$950 , \6090_N$951 , \6091_N$952 , \6092_N$953 , \6093_N$954 , \6094_N$955 ,
         \6095_N$956 , \6096_N$957 , \6097_N$958 , \6098_N$959 , \6099_N$960 , \6100_N$961 , \6101_N$962 , \6102_N$963 , \6103_N$964 , \6104_N$965 ,
         \6105_N$966 , \6106_N$967 , \6107_N$968 , \6108_N$969 , \6109_N$970 , \6110_N$971 , \6111_N$972 , \6112_N$973 , \6113_N$974 , \6114_N$975 ,
         \6115_N$976 , \6116_N$977 , \6117_N$978 , \6118_N$979 , \6119_N$980 , \6120_N$981 , \6121_N$982 , \6122_N$983 , \6123_N$984 , \6124_N$985 ,
         \6125_N$986 , \6126_N$987 , \6127_N$988 , \6128_N$989 , \6129_N$990 , \6130_N$991 , \6131_N$992 , \6132_N$993 , \6133_N$994 , \6134_N$995 ,
         \6135_N$996 , \6136_N$997 , \6137_N$998 , \6138_N$999 , \6139_N$1000 , \6140_N$1001 , \6141_N$1002 , \6142_N$1003 , \6143_N$1004 , \6144_N$1005 ,
         \6145_N$1006 , \6146_N$1007 , \6147_N$1008 , \6148_N$1009 , \6149_N$1010 , \6150_N$1011 , \6151_N$1012 , \6152_N$1013 , \6153_N$1014 , \6154_N$1015 ,
         \6155_N$1016 , \6156_N$1017 , \6157_N$1018 , \6158_N$1019 , \6159_N$1020 , \6160_N$1021 , \6161_N$1022 , \6162_N$1023 , \6163_N$1024 , \6164_N$1025 ,
         \6165_N$1026 , \6166_N$1027 , \6167_N$1028 , \6168_N$1029 , \6169_N$1030 , \6170_N$1031 , \6171_N$1032 , \6172_N$1033 , \6173_N$1034 , \6174_N$1035 ,
         \6175_N$1036 , \6176_N$1037 , \6177_N$1038 , \6178_N$1039 , \6179_N$1040 , \6180_N$1041 , \6181_N$1042 , \6182_N$1043 , \6183_N$1044 , \6184_N$1045 ,
         \6185_N$1046 , \6186_N$1047 , \6187_N$1048 , \6188_N$1049 , \6189_N$1050 , \6190_N$1051 , \6191_N$1052 , \6192_N$1053 , \6193_N$1054 , \6194_N$1055 ,
         \6195_N$1056 , \6196_N$1057 , \6197_N$1058 , \6198_N$1059 , \6199_N$1060 , \6200_N$1061 , \6201_N$1062 , \6202_N$1063 , \6203_N$1064 , \6204_N$1065 ,
         \6205_N$1066 , \6206_N$1067 , \6207_N$1068 , \6208_N$1069 , \6209_N$1070 , \6210_N$1071 , \6211_N$1072 , \6212_N$1073 , \6213_N$1074 , \6214_N$1075 ,
         \6215_N$1076 , \6216_N$1077 , \6217_N$1078 , \6218_N$1079 , \6219_N$1080 , \6220_N$1081 , \6221_N$1082 , \6222_N$1083 , \6223_N$1084 , \6224_N$1085 ,
         \6225_N$1086 , \6226_N$1087 , \6227_N$1088 , \6228_N$1089 , \6229_N$1090 , \6230_N$1091 , \6231_N$1092 , \6232_N$1093 , \6233_N$1094 , \6234_N$1095 ,
         \6235_N$1096 , \6236_N$1097 , \6237_N$1098 , \6238_N$1099 , \6239_N$1100 , \6240_N$1101 , \6241_N$1102 , \6242_N$1103 , \6243_N$1104 , \6244_N$1105 ,
         \6245_N$1106 , \6246_N$1107 , \6247_N$1108 , \6248_N$1109 , \6249_N$1110 , \6250_N$1111 , \6251_N$1112 , \6252_N$1113 , \6253_N$1114 , \6254_N$1115 ,
         \6255_N$1116 , \6256_N$1117 , \6257_N$1118 , \6258_N$1119 , \6259_N$1120 , \6260_N$1121 , \6261_N$1122 , \6262_N$1123 , \6263_N$1124 , \6264_N$1125 ,
         \6265_N$1126 , \6266_N$1127 , \6267_N$1128 , \6268_N$1129 , \6269_N$1130 , \6270_N$1131 , \6271_N$1132 , \6272_N$1133 , \6273_N$1134 , \6274_N$1135 ,
         \6275_N$1136 , \6276_N$1137 , \6277_N$1138 , \6278_N$1139 , \6279_N$1140 , \6280_N$1141 , \6281_N$1142 , \6282_N$1143 , \6283_N$1144 , \6284_N$1145 ,
         \6285_N$1146 , \6286_N$1147 , \6287_N$1148 , \6288_N$1149 , \6289_N$1150 , \6290_N$1151 , \6291_N$1152 , \6292_N$1153 , \6293_N$1154 , \6294_N$1155 ,
         \6295_N$1156 , \6296_N$1157 , \6297_N$1158 , \6298_N$1159 , \6299_N$1160 , \6300_N$1161 , \6301_N$1162 , \6302_N$1163 , \6303_N$1164 , \6304_N$1165 ,
         \6305_N$1166 , \6306_N$1167 , \6307_N$1168 , \6308_N$1169 , \6309_N$1170 , \6310_N$1171 , \6311_N$1172 , \6312_N$1173 , \6313_N$1174 , \6314_N$1175 ,
         \6315_N$1176 , \6316_N$1177 , \6317_N$1178 , \6318_N$1179 , \6319_N$1180 , \6320_N$1181 , \6321_N$1182 , \6322_N$1183 , \6323_N$1184 , \6324_N$1185 ,
         \6325_N$1186 , \6326_N$1187 , \6327_N$1188 , \6328_N$1189 , \6329_N$1190 , \6330_N$1191 , \6331_N$1192 , \6332_N$1193 , \6333_N$1194 , \6334_N$1195 ,
         \6335_N$1196 , \6336_N$1197 , \6337_N$1198 , \6338_N$1199 , \6339_N$1200 , \6340_N$1201 , \6341_N$1202 , \6342_N$1203 , \6343_N$1204 , \6344_N$1205 ,
         \6345_N$1206 , \6346_N$1207 , \6347_N$1208 , \6348_N$1209 , \6349_N$1210 , \6350_N$1211 , \6351_N$1212 , \6352_N$1213 , \6353_N$1214 , \6354_N$1215 ,
         \6355_N$1216 , \6356_N$1217 , \6357_N$1218 , \6358_N$1219 , \6359_N$1220 , \6360_N$1221 , \6361_N$1222 , \6362_N$1223 , \6363_N$1224 , \6364_N$1225 ,
         \6365_N$1226 , \6366_N$1227 , \6367_N$1228 , \6368_N$1229 , \6369_N$1230 , \6370_N$1231 , \6371_N$1232 , \6372_N$1233 , \6373_N$1234 , \6374_N$1235 ,
         \6375_N$1236 , \6376_N$1237 , \6377_N$1238 , \6378_N$1239 , \6379_N$1240 , \6380_N$1241 , \6381_N$1242 , \6382_N$1243 , \6383_N$1244 , \6384_N$1245 ,
         \6385_N$1246 , \6386_N$1247 , \6387_N$1248 , \6388_N$1249 , \6389_N$1250 , \6390_N$1251 , \6391_N$1252 , \6392_N$1253 , \6393_N$1254 , \6394_N$1255 ,
         \6395_N$1256 , \6396_N$1257 , \6397_N$1258 , \6398_N$1259 , \6399_N$1260 , \6400_N$1261 , \6401_N$1262 , \6402_N$1263 , \6403_N$1264 , \6404_N$1265 ,
         \6405_N$1266 , \6406_N$1267 , \6407_N$1268 , \6408_N$1269 , \6409_N$1270 , \6410_N$1271 , \6411_N$1272 , \6412_N$1273 , \6413_N$1274 , \6414_N$1275 ,
         \6415_N$1276 , \6416_N$1277 , \6417_N$1278 , \6418_N$1279 , \6419_N$1280 , \6420_N$1281 , \6421_N$1282 , \6422_N$1283 , \6423_N$1284 , \6424_N$1285 ,
         \6425_N$1286 , \6426_N$1287 , \6427_N$1288 , \6428_N$1289 , \6429_N$1290 , \6430_N$1291 , \6431_N$1292 , \6432_N$1293 , \6433_N$1294 , \6434_N$1295 ,
         \6435_N$1296 , \6436_N$1297 , \6437_N$1298 , \6438_N$1299 , \6439_N$1300 , \6440_N$1301 , \6441_N$1302 , \6442_N$1303 , \6443_N$1304 , \6444_N$1305 ,
         \6445_N$1306 , \6446_N$1307 , \6447_N$1308 , \6448_N$1309 , \6449_N$1310 , \6450_N$1311 , \6451_N$1312 , \6452_N$1313 , \6453_N$1314 , \6454_N$1315 ,
         \6455_N$1316 , \6456_N$1317 , \6457_N$1318 , \6458_N$1319 , \6459_N$1320 , \6460_N$1321 , \6461_N$1322 , \6462_N$1323 , \6463_N$1324 , \6464_N$1325 ,
         \6465_N$1326 , \6466_N$1327 , \6467_N$1328 , \6468_N$1329 , \6469_N$1330 , \6470_N$1331 , \6471_N$1332 , \6472_N$1333 , \6473_N$1334 , \6474_N$1335 ,
         \6475_N$1336 , \6476_N$1337 , \6477_N$1338 , \6478_N$1339 , \6479_N$1340 , \6480_N$1341 , \6481_N$1342 , \6482_N$1343 , \6483_N$1344 , \6484_N$1345 ,
         \6485_N$1346 , \6486_N$1347 , \6487_N$1348 , \6488_N$1349 , \6489_N$1350 , \6490_N$1351 , \6491_N$1352 , \6492_N$1353 , \6493_N$1354 , \6494_N$1355 ,
         \6495_N$1356 , \6496_N$1357 , \6497_N$1358 , \6498_N$1359 , \6499_N$1360 , \6500_N$1361 , \6501_N$1362 , \6502_N$1363 , \6503_N$1364 , \6504_N$1365 ,
         \6505_N$1366 , \6506_N$1367 , \6507_N$1368 , \6508_N$1369 , \6509_N$1370 , \6510_N$1371 , \6511_N$1372 , \6512_N$1373 , \6513_N$1374 , \6514_N$1375 ,
         \6515_N$1376 , \6516_N$1377 , \6517_N$1378 , \6518_N$1379 , \6519_N$1380 , \6520_N$1381 , \6521_N$1382 , \6522_N$1383 , \6523_N$1384 , \6524_N$1385 ,
         \6525_N$1386 , \6526_N$1387 , \6527_N$1388 , \6528_N$1389 , \6529_N$1390 , \6530_N$1391 , \6531_N$1392 , \6532_N$1393 , \6533_N$1394 , \6534_N$1395 ,
         \6535_N$1396 , \6536_N$1397 , \6537_N$1398 , \6538_N$1399 , \6539_N$1400 , \6540_N$1401 , \6541_N$1402 , \6542_N$1403 , \6543_N$1404 , \6544_N$1405 ,
         \6545_N$1406 , \6546_N$1407 , \6547_N$1408 , \6548_N$1409 , \6549_N$1410 , \6550_N$1411 , \6551_N$1412 , \6552_N$1413 , \6553_N$1414 , \6554_N$1415 ,
         \6555_N$1416 , \6556_N$1417 , \6557_N$1418 , \6558_N$1419 , \6559_N$1420 , \6560_N$1421 , \6561_N$1422 , \6562_N$1423 , \6563_N$1424 , \6564_N$1425 ,
         \6565_N$1426 , \6566_N$1427 , \6567_N$1428 , \6568_N$1429 , \6569_N$1430 , \6570_N$1431 , \6571_N$1432 , \6572_N$1433 , \6573_N$1434 , \6574_N$1435 ,
         \6575_N$1436 , \6576_N$1437 , \6577_N$1438 , \6578_N$1439 , \6579_N$1440 , \6580_N$1441 , \6581_N$1442 , \6582_N$1443 , \6583_N$1444 , \6584_N$1445 ,
         \6585_N$1446 , \6586_N$1447 , \6587_N$1448 , \6588_N$1449 , \6589_N$1450 , \6590_N$1451 , \6591_N$1452 , \6592_N$1453 , \6593_N$1454 , \6594_N$1455 ,
         \6595_N$1456 , \6596_N$1457 , \6597_N$1458 , \6598_N$1459 , \6599_N$1460 , \6600_N$1461 , \6601_N$1462 , \6602_N$1463 , \6603_N$1464 , \6604_N$1465 ,
         \6605_N$1466 , \6606_N$1467 , \6607_N$1468 , \6608_N$1469 , \6609_N$1470 , \6610_N$1471 , \6611_N$1472 , \6612_N$1473 , \6613_N$1474 , \6614_N$1475 ,
         \6615_N$1476 , \6616_N$1477 , \6617_N$1478 , \6618_N$1479 , \6619_N$1480 , \6620_N$1481 , \6621_N$1482 , \6622_N$1483 , \6623_N$1484 , \6624_N$1485 ,
         \6625_N$1486 , \6626_N$1487 , \6627_N$1488 , \6628_N$1489 , \6629_N$1490 , \6630_N$1491 , \6631_N$1492 , \6632_N$1493 , \6633_N$1494 , \6634_N$1495 ,
         \6635_N$1496 , \6636_N$1497 , \6637_N$1498 , \6638_N$1499 , \6639_N$1500 , \6640_N$1501 , \6641_N$1502 , \6642_N$1503 , \6643_N$1504 , \6644_N$1505 ,
         \6645_N$1506 , \6646_N$1507 , \6647_N$1508 , \6648_N$1509 , \6649_N$1510 , \6650_N$1511 , \6651_N$1512 , \6652_N$1513 , \6653_N$1514 , \6654_N$1515 ,
         \6655_N$1516 , \6656_N$1517 , \6657_N$1518 , \6658_N$1519 , \6659_N$1520 , \6660_N$1521 , \6661_N$1522 , \6662_N$1523 , \6663_N$1524 , \6664_N$1525 ,
         \6665_N$1526 , \6666_N$1527 , \6667_N$1528 , \6668_N$1529 , \6669_N$1530 , \6670_N$1531 , \6671_N$1532 , \6672_N$1533 , \6673_N$1534 , \6674_N$1535 ,
         \6675_N$1536 , \6676_N$1537 , \6677_N$1538 , \6678_N$1539 , \6679_N$1540 , \6680_N$1541 , \6681_N$1542 , \6682_N$1543 , \6683_N$1544 , \6684_N$1545 ,
         \6685_N$1546 , \6686_N$1547 , \6687_N$1548 , \6688_N$1549 , \6689_N$1550 , \6690_N$1551 , \6691_N$1552 , \6692_N$1553 , \6693_N$1554 , \6694_N$1555 ,
         \6695_N$1556 , \6696_N$1557 , \6697_N$1558 , \6698_N$1559 , \6699_N$1560 , \6700_N$1561 , \6701_N$1562 , \6702_N$1563 , \6703_N$1564 , \6704_N$1565 ,
         \6705_N$1566 , \6706_N$1567 , \6707_N$1568 , \6708_N$1569 , \6709_N$1570 , \6710_N$1571 , \6711_N$1572 , \6712_N$1573 , \6713_N$1574 , \6714_N$1575 ,
         \6715_N$1576 , \6716_N$1577 , \6717_N$1578 , \6718_N$1579 , \6719_N$1580 , \6720_N$1581 , \6721_N$1582 , \6722_N$1583 , \6723_N$1584 , \6724_N$1585 ,
         \6725_N$1586 , \6726_N$1587 , \6727_N$1588 , \6728_N$1589 , \6729_N$1590 , \6730_N$1591 , \6731_N$1592 , \6732_N$1593 , \6733_N$1594 , \6734_N$1595 ,
         \6735_N$1596 , \6736_N$1597 , \6737_N$1598 , \6738_N$1599 , \6739_N$1600 , \6740_N$1601 , \6741_N$1602 , \6742_N$1603 , \6743_N$1604 , \6744_N$1605 ,
         \6745_N$1606 , \6746_N$1607 , \6747_N$1608 , \6748_N$1609 , \6749_N$1610 , \6750_N$1611 , \6751_N$1612 , \6752_N$1613 , \6753_N$1614 , \6754_N$1615 ,
         \6755_N$1616 , \6756_N$1617 , \6757_N$1618 , \6758_N$1619 , \6759_N$1620 , \6760_N$1621 , \6761_N$1622 , \6762_N$1623 , \6763_N$1624 , \6764_N$1625 ,
         \6765_N$1626 , \6766_N$1627 , \6767_N$1628 , \6768_N$1629 , \6769_N$1630 , \6770_N$1631 , \6771_N$1632 , \6772_N$1633 , \6773_N$1634 , \6774_N$1635 ,
         \6775_N$1636 , \6776_N$1637 , \6777_N$1638 , \6778_N$1639 , \6779_N$1640 , \6780_N$1641 , \6781_N$1642 , \6782_N$1643 , \6783_N$1644 , \6784_N$1645 ,
         \6785_N$1646 , \6786_N$1647 , \6787_N$1648 , \6788_N$1649 , \6789_N$1650 , \6790_N$1651 , \6791_N$1652 , \6792_N$1653 , \6793_N$1654 , \6794_N$1655 ,
         \6795_N$1656 , \6796_N$1657 , \6797_N$1658 , \6798_N$1659 , \6799_N$1660 , \6800_N$1661 , \6801_N$1662 , \6802_N$1663 , \6803_N$1664 , \6804_N$1665 ,
         \6805_N$1666 , \6806_N$1667 , \6807_N$1668 , \6808_N$1669 , \6809_N$1670 , \6810_N$1671 , \6811_N$1672 , \6812_N$1673 , \6813_N$1674 , \6814_N$1675 ,
         \6815_N$1676 , \6816_N$1677 , \6817_N$1678 , \6818_N$1679 , \6819_N$1680 , \6820_N$1681 , \6821_N$1682 , \6822_N$1683 , \6823_N$1684 , \6824_N$1685 ,
         \6825_N$1686 , \6826_N$1687 , \6827_N$1688 , \6828_N$1689 , \6829_N$1690 , \6830_N$1691 , \6831_N$1692 , \6832_N$1693 , \6833_N$1694 , \6834_N$1695 ,
         \6835_N$1696 , \6836_N$1697 , \6837_N$1698 , \6838_N$1699 , \6839_N$1700 , \6840_N$1701 , \6841_N$1702 , \6842_N$1703 , \6843_N$1704 , \6844_N$1705 ,
         \6845_N$1706 , \6846_N$1707 , \6847_N$1708 , \6848_N$1709 , \6849_N$1710 , \6850_N$1711 , \6851_N$1712 , \6852_N$1713 , \6853_N$1714 , \6854_N$1715 ,
         \6855_N$1716 , \6856_N$1717 , \6857_N$1718 , \6858_N$1719 , \6859_N$1720 , \6860_N$1721 , \6861_N$1722 , \6862_N$1723 , \6863_N$1724 , \6864_N$1725 ,
         \6865_N$1726 , \6866_N$1727 , \6867_N$1728 , \6868_N$1729 , \6869_N$1730 , \6870_N$1731 , \6871_N$1732 , \6872_N$1733 , \6873_N$1734 , \6874_N$1735 ,
         \6875_N$1736 , \6876_N$1737 , \6877_N$1738 , \6878_N$1739 , \6879_N$1740 , \6880_N$1741 , \6881_N$1742 , \6882_N$1743 , \6883_N$1744 , \6884_N$1745 ,
         \6885_N$1746 , \6886_N$1747 , \6887_N$1748 , \6888_N$1749 , \6889_N$1750 , \6890_N$1751 , \6891_N$1752 , \6892_N$1753 , \6893_N$1754 , \6894_N$1755 ,
         \6895_N$1756 , \6896_N$1757 , \6897_N$1758 , \6898_N$1759 , \6899_N$1760 , \6900_N$1761 , \6901_N$1762 , \6902_N$1763 , \6903_N$1764 , \6904_N$1765 ,
         \6905_N$1766 , \6906_N$1767 , \6907_N$1768 , \6908_N$1769 , \6909_N$1770 , \6910_N$1771 , \6911_N$1772 , \6912_N$1773 , \6913_N$1774 , \6914_N$1775 ,
         \6915_N$1776 , \6916_N$1777 , \6917_N$1778 , \6918_N$1779 , \6919_N$1780 , \6920_N$1781 , \6921_N$1782 , \6922_N$1783 , \6923_N$1784 , \6924_N$1785 ,
         \6925_N$1786 , \6926_N$1787 , \6927_N$1788 , \6928_N$1789 , \6929_N$1790 , \6930_N$1791 , \6931_N$1792 , \6932_N$1793 , \6933_N$1794 , \6934_N$1795 ,
         \6935_N$1796 , \6936_N$1797 , \6937_N$1798 , \6938_N$1799 , \6939_N$1800 , \6940_N$1801 , \6941_N$1802 , \6942_N$1803 , \6943_N$1804 , \6944_N$1805 ,
         \6945_N$1806 , \6946_N$1807 , \6947_N$1808 , \6948_N$1809 , \6949_N$1810 , \6950_N$1811 , \6951_N$1812 , \6952_N$1813 , \6953_N$1814 , \6954_N$1815 ,
         \6955_N$1816 , \6956_N$1817 , \6957_N$1818 , \6958_N$1819 , \6959_N$1820 , \6960_N$1821 , \6961_N$1822 , \6962_N$1823 , \6963_N$1824 , \6964_N$1825 ,
         \6965_N$1826 , \6966_N$1827 , \6967_N$1828 , \6968_N$1829 , \6969_N$1830 , \6970_N$1831 , \6971_N$1832 , \6972_N$1833 , \6973_N$1834 , \6974_N$1835 ,
         \6975_N$1836 , \6976_N$1837 , \6977_N$1838 , \6978_N$1839 , \6979_N$1840 , \6980_N$1841 , \6981_N$1842 , \6982_N$1843 , \6983_N$1844 , \6984_N$1845 ,
         \6985_N$1846 , \6986_N$1847 , \6987_N$1848 , \6988_N$1849 , \6989_N$1850 , \6990_N$1851 , \6991_N$1852 , \6992_N$1853 , \6993_N$1854 , \6994_N$1855 ,
         \6995_N$1856 , \6996_N$1857 , \6997_N$1858 , \6998_N$1859 , \6999_N$1860 , \7000_N$1861 , \7001_N$1862 , \7002_N$1863 , \7003_N$1864 , \7004_N$1865 ,
         \7005_N$1866 , \7006_N$1867 , \7007_N$1868 , \7008_N$1869 , \7009_N$1870 , \7010_N$1871 , \7011_N$1872 , \7012_N$1873 , \7013_N$1874 , \7014_N$1875 ,
         \7015_N$1876 , \7016_N$1877 , \7017_N$1878 , \7018_N$1879 , \7019_N$1880 , \7020_N$1881 , \7021_N$1882 , \7022_N$1883 , \7023_N$1884 , \7024_N$1885 ,
         \7025_N$1886 , \7026_N$1887 , \7027_N$1888 , \7028_ZERO , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 ,
         \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042_N$1 , \7043_N$3 , \7044_N$6 ,
         \7045_N$18 , \7046_N$20 , \7047_N$23 , \7048_N$34 , \7049_N$36 , \7050_N$39 , \7051_N$51 , \7052_N$52 , \7053_N$54 , \7054_N$57 ,
         \7055_ONE , \7056 , \7057 , \7058 , \7059 , \7060_nG14890 , \7061 , \7062 , \7063 , \7064 ,
         \7065 , \7066 , \7067 , \7068_nG14891 , \7069 , \7070 , \7071 , \7072 , \7073 , \7074_nG14897 ,
         \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 , \7083 , \7084 ,
         \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 , \7093 , \7094 ,
         \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 ,
         \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114_nG32b3 ,
         \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122_nG32bb , \7123 , \7124 ,
         \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131_nG32c4 , \7132 , \7133 , \7134 ,
         \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141_nG32ce , \7142 , \7143 , \7144 ,
         \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151_nG32d8 , \7152 , \7153 , \7154 ,
         \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161_nG32e2 , \7162 , \7163 , \7164 ,
         \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171_nG32ec , \7172 , \7173 , \7174 ,
         \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181_nG32f6 , \7182 , \7183 , \7184 ,
         \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191_nG3300 , \7192 , \7193 , \7194 ,
         \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 , \7203_nG330c , \7204 ,
         \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212_nG3315 , \7213 , \7214 ,
         \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222_nG331f , \7223 , \7224 ,
         \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232_nG3329 , \7233 , \7234 ,
         \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242_nG3331 , \7243 , \7244 ,
         \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252_nG3339 , \7253 , \7254 ,
         \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262_nG3341 , \7263 , \7264 ,
         \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272_nG3349 , \7273 , \7274 ,
         \7275 , \7276 , \7277 , \7278 , \7279 , \7280_nG3351 , \7281 , \7282 , \7283 , \7284 ,
         \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 , \7293 , \7294 ,
         \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 , \7303 , \7304 ,
         \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 , \7313 , \7314 ,
         \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 , \7322 , \7323 , \7324 ,
         \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 , \7333 , \7334 ,
         \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 , \7343 , \7344 ,
         \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 , \7352 , \7353 , \7354 ,
         \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 , \7363 , \7364 ,
         \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 , \7373 , \7374 ,
         \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 , \7382 , \7383 , \7384 ,
         \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 , \7393 , \7394 ,
         \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 , \7403 , \7404 ,
         \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 , \7413 , \7414 ,
         \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 , \7423 , \7424 ,
         \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 , \7432 , \7433 , \7434 ,
         \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 , \7442 , \7443 , \7444 ,
         \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 , \7452 , \7453 , \7454 ,
         \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 , \7462 , \7463 , \7464 ,
         \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 , \7472 , \7473 , \7474 ,
         \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 , \7482 , \7483 , \7484 ,
         \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 , \7492 , \7493 , \7494 ,
         \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 , \7502 , \7503 , \7504 ,
         \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 , \7512 , \7513 , \7514 ,
         \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 , \7522 , \7523 , \7524 ,
         \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 , \7532 , \7533 , \7534 ,
         \7535 , \7536 , \7537 , \7538 , \7539 , \7540 , \7541 , \7542 , \7543 , \7544 ,
         \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 , \7552 , \7553 , \7554 ,
         \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 , \7562 , \7563 , \7564 ,
         \7565 , \7566 , \7567 , \7568 , \7569 , \7570 , \7571 , \7572 , \7573 , \7574 ,
         \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 , \7582 , \7583 , \7584 ,
         \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 , \7592 , \7593 , \7594 ,
         \7595 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 , \7602 , \7603 , \7604 ,
         \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 , \7612 , \7613 , \7614 ,
         \7615 , \7616 , \7617 , \7618 , \7619 , \7620 , \7621 , \7622 , \7623 , \7624 ,
         \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 , \7632 , \7633 , \7634 ,
         \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 , \7642 , \7643 , \7644 ,
         \7645 , \7646 , \7647 , \7648 , \7649 , \7650 , \7651 , \7652 , \7653 , \7654 ,
         \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 , \7662 , \7663 , \7664 ,
         \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 , \7672 , \7673 , \7674 ,
         \7675 , \7676 , \7677 , \7678 , \7679 , \7680 , \7681 , \7682 , \7683 , \7684 ,
         \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 , \7692 , \7693 , \7694 ,
         \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 , \7702 , \7703 , \7704 ,
         \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 , \7712 , \7713 , \7714 ,
         \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 , \7722 , \7723 , \7724 ,
         \7725 , \7726 , \7727 , \7728 , \7729 , \7730 , \7731 , \7732 , \7733 , \7734 ,
         \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 , \7742 , \7743 , \7744 ,
         \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 , \7752 , \7753 , \7754 ,
         \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 , \7762 , \7763 , \7764 ,
         \7765 , \7766 , \7767 , \7768 , \7769 , \7770 , \7771 , \7772 , \7773 , \7774 ,
         \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 , \7782 , \7783 , \7784 ,
         \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791 , \7792 , \7793 , \7794 ,
         \7795 , \7796 , \7797 , \7798 , \7799 , \7800 , \7801 , \7802 , \7803 , \7804 ,
         \7805 , \7806 , \7807_nG3568 , \7808 , \7809 , \7810 , \7811 , \7812 , \7813 , \7814 ,
         \7815 , \7816 , \7817 , \7818 , \7819 , \7820 , \7821 , \7822 , \7823 , \7824 ,
         \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 , \7832 , \7833 , \7834 ,
         \7835 , \7836 , \7837 , \7838 , \7839 , \7840 , \7841 , \7842 , \7843 , \7844 ,
         \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 , \7852 , \7853 , \7854 ,
         \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 , \7862 , \7863 , \7864 ,
         \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 , \7872 , \7873 , \7874 ,
         \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 , \7883 , \7884 ,
         \7885 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891 , \7892 , \7893 , \7894 ,
         \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 , \7903 , \7904 ,
         \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 , \7913 , \7914 ,
         \7915 , \7916 , \7917 , \7918 , \7919 , \7920 , \7921 , \7922 , \7923 , \7924 ,
         \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 , \7933 , \7934 ,
         \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 , \7942 , \7943 , \7944 ,
         \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 , \7952 , \7953 , \7954 ,
         \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 , \7963 , \7964 ,
         \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 , \7972 , \7973 , \7974 ,
         \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 , \7983 , \7984 ,
         \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 , \7992 , \7993 , \7994 ,
         \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 , \8002 , \8003 , \8004 ,
         \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 , \8013 , \8014 ,
         \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 , \8022 , \8023 , \8024 ,
         \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 , \8032 , \8033 , \8034 ,
         \8035 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 , \8042 , \8043 , \8044 ,
         \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 , \8053 , \8054 ,
         \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 , \8062 , \8063 , \8064 ,
         \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 , \8072 , \8073 , \8074 ,
         \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 , \8082 , \8083 , \8084 ,
         \8085 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 , \8092 , \8093 , \8094 ,
         \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 , \8103 , \8104 ,
         \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 , \8112 , \8113 , \8114 ,
         \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 , \8122 , \8123 , \8124 ,
         \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 , \8132 , \8133 , \8134 ,
         \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 , \8142 , \8143 , \8144 ,
         \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 , \8152 , \8153 , \8154 ,
         \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 , \8162 , \8163 , \8164 ,
         \8165 , \8166 , \8167 , \8168 , \8169 , \8170 , \8171 , \8172 , \8173 , \8174 ,
         \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 , \8182 , \8183 , \8184 ,
         \8185 , \8186 , \8187 , \8188 , \8189 , \8190 , \8191 , \8192 , \8193 , \8194 ,
         \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 , \8202 , \8203 , \8204 ,
         \8205 , \8206 , \8207 , \8208 , \8209 , \8210 , \8211 , \8212 , \8213 , \8214 ,
         \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 , \8222 , \8223 , \8224 ,
         \8225 , \8226 , \8227 , \8228 , \8229 , \8230 , \8231 , \8232 , \8233 , \8234 ,
         \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 , \8242 , \8243 , \8244 ,
         \8245 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 , \8252 , \8253 , \8254 ,
         \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 , \8262 , \8263 , \8264 ,
         \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271 , \8272 , \8273 , \8274 ,
         \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 , \8282 , \8283 , \8284 ,
         \8285 , \8286 , \8287 , \8288 , \8289 , \8290 , \8291 , \8292 , \8293 , \8294 ,
         \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 , \8302 , \8303 , \8304 ,
         \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 , \8312 , \8313 , \8314 ,
         \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 , \8322 , \8323 , \8324 ,
         \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 , \8332_nG3775 , \8333 , \8334 ,
         \8335 , \8336 , \8337 , \8338 , \8339 , \8340 , \8341 , \8342 , \8343 , \8344 ,
         \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 , \8352 , \8353 , \8354 ,
         \8355 , \8356 , \8357 , \8358 , \8359 , \8360 , \8361 , \8362 , \8363 , \8364 ,
         \8365 , \8366 , \8367_nG3798 , \8368 , \8369 , \8370 , \8371 , \8372 , \8373 , \8374 ,
         \8375 , \8376 , \8377 , \8378 , \8379 , \8380 , \8381 , \8382 , \8383 , \8384 ,
         \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 , \8392 , \8393 , \8394 ,
         \8395 , \8396 , \8397 , \8398 , \8399 , \8400 , \8401 , \8402 , \8403_nG37bc , \8404 ,
         \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 , \8412 , \8413 , \8414 ,
         \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 , \8422 , \8423 , \8424 ,
         \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 , \8432 , \8433 , \8434 ,
         \8435 , \8436 , \8437 , \8438 , \8439_nG37e0 , \8440 , \8441 , \8442 , \8443 , \8444 ,
         \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 , \8452 , \8453 , \8454 ,
         \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 , \8462 , \8463 , \8464 ,
         \8465 , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 , \8472 , \8473 , \8474 ,
         \8475_nG3804 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 , \8482 , \8483 , \8484 ,
         \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 , \8492 , \8493 , \8494 ,
         \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 , \8502 , \8503 , \8504 ,
         \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511_nG3828 , \8512 , \8513 , \8514 ,
         \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 , \8522 , \8523 , \8524 ,
         \8525 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 , \8532 , \8533 , \8534 ,
         \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 , \8542 , \8543 , \8544 ,
         \8545 , \8546 , \8547_nG384c , \8548 , \8549 , \8550 , \8551 , \8552 , \8553 , \8554 ,
         \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 , \8562 , \8563 , \8564 ,
         \8565 , \8566 , \8567 , \8568 , \8569 , \8570 , \8571 , \8572 , \8573 , \8574 ,
         \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 , \8582 , \8583_nG3870 , \8584 ,
         \8585 , \8586 , \8587 , \8588 , \8589 , \8590 , \8591 , \8592 , \8593 , \8594 ,
         \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 ,
         \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 , \8612 , \8613 , \8614 ,
         \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 , \8622 , \8623 , \8624 ,
         \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 , \8632 , \8633 , \8634 ,
         \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 , \8643 , \8644 ,
         \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 , \8653 , \8654 ,
         \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 , \8663 , \8664 ,
         \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 , \8672 , \8673 , \8674 ,
         \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 , \8682 , \8683 , \8684 ,
         \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 ,
         \8695 , \8696 , \8697 , \8698 , \8699 , \8700 , \8701 , \8702 , \8703 , \8704 ,
         \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 ,
         \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 , \8722 , \8723 , \8724 ,
         \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 , \8732 , \8733 , \8734 ,
         \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 , \8742 , \8743 , \8744 ,
         \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 ,
         \8755 , \8756 , \8757 , \8758 , \8759 , \8760 , \8761 , \8762 , \8763 , \8764 ,
         \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 , \8772 , \8773 , \8774 ,
         \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 , \8782 , \8783 , \8784 ,
         \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 , \8792 , \8793 , \8794 ,
         \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 , \8802 , \8803 , \8804 ,
         \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 , \8812 , \8813 , \8814 ,
         \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 , \8822 , \8823 , \8824 ,
         \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 , \8832 , \8833 , \8834 ,
         \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 , \8842 , \8843 , \8844 ,
         \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 , \8852 , \8853 , \8854 ,
         \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 , \8862 , \8863 , \8864 ,
         \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 , \8872 , \8873 , \8874 ,
         \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 , \8882 , \8883 , \8884 ,
         \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 , \8892 , \8893 , \8894 ,
         \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 , \8902 , \8903 , \8904 ,
         \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 , \8912 , \8913 , \8914 ,
         \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 , \8922 , \8923 , \8924 ,
         \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 , \8932 , \8933 , \8934 ,
         \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 , \8942 , \8943 , \8944 ,
         \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 , \8952 , \8953 , \8954 ,
         \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 , \8962 , \8963 , \8964 ,
         \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 , \8972 , \8973 , \8974 ,
         \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 , \8982 , \8983 , \8984 ,
         \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 , \8992 , \8993 , \8994 ,
         \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 , \9002 , \9003 , \9004 ,
         \9005 , \9006 , \9007 , \9008 , \9009 , \9010 , \9011 , \9012 , \9013 , \9014 ,
         \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 , \9022 , \9023 , \9024 ,
         \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 , \9032 , \9033 , \9034 ,
         \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 , \9042 , \9043 , \9044 ,
         \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 , \9052 , \9053 , \9054 ,
         \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 , \9062 , \9063 , \9064 ,
         \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 , \9072 , \9073 , \9074 ,
         \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 , \9082 , \9083 , \9084 ,
         \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 , \9092 , \9093 , \9094 ,
         \9095 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 , \9102 , \9103 , \9104 ,
         \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 , \9112 , \9113_nG3a82 , \9114 ,
         \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 , \9122 , \9123 , \9124 ,
         \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 , \9132 , \9133 , \9134 ,
         \9135 , \9136 , \9137 , \9138 , \9139 , \9140 , \9141 , \9142 , \9143 , \9144 ,
         \9145 , \9146 , \9147 , \9148_nG3aa5 , \9149 , \9150 , \9151 , \9152 , \9153 , \9154 ,
         \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 , \9162 , \9163 , \9164 ,
         \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 , \9172 , \9173 , \9174 ,
         \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 , \9182 , \9183 , \9184_nG3ac9 ,
         \9185 , \9186 , \9187 , \9188 , \9189 , \9190 , \9191 , \9192 , \9193 , \9194 ,
         \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 , \9202 , \9203 , \9204 ,
         \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 , \9212 , \9213 , \9214 ,
         \9215 , \9216 , \9217 , \9218 , \9219 , \9220_nG3aed , \9221 , \9222 , \9223 , \9224 ,
         \9225 , \9226 , \9227 , \9228 , \9229 , \9230 , \9231 , \9232 , \9233 , \9234 ,
         \9235 , \9236 , \9237 , \9238 , \9239 , \9240 , \9241 , \9242 , \9243 , \9244 ,
         \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 , \9252 , \9253 , \9254 ,
         \9255 , \9256_nG3b03 , \9257 , \9258 , \9259 , \9260 , \9261 , \9262 , \9263 , \9264 ,
         \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 , \9272 , \9273 , \9274 ,
         \9275 , \9276 , \9277 , \9278 , \9279 , \9280 , \9281 , \9282 , \9283 , \9284 ,
         \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 , \9292_nG3b19 , \9293 , \9294 ,
         \9295 , \9296 , \9297 , \9298 , \9299 , \9300 , \9301 , \9302 , \9303 , \9304 ,
         \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 , \9312 , \9313 , \9314 ,
         \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 , \9322 , \9323 , \9324 ,
         \9325 , \9326 , \9327 , \9328_nG3b2f , \9329 , \9330 , \9331 , \9332 , \9333 , \9334 ,
         \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 , \9342 , \9343 , \9344 ,
         \9345 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 , \9352 , \9353 , \9354 ,
         \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 , \9362 , \9363 , \9364_nG3b45 ,
         \9365 , \9366 , \9367 , \9368 , \9369 , \9370 , \9371_nG3b4c , \9372 , \9373 , \9374 ,
         \9375 , \9376 , \9377 , \9378 , \9379 , \9380 , \9381 , \9382_nG3b57 , \9383 , \9384 ,
         \9385 , \9386 , \9387 , \9388 , \9389 , \9390 , \9391 , \9392 , \9393 , \9394 ,
         \9395 , \9396 , \9397 , \9398 , \9399 , \9400 , \9401 , \9402 , \9403 , \9404 ,
         \9405 , \9406 , \9407 , \9408 , \9409 , \9410 , \9411 , \9412 , \9413 , \9414 ,
         \9415 , \9416 , \9417 , \9418 , \9419 , \9420 , \9421 , \9422_nG3b80 , \9423 , \9424 ,
         \9425 , \9426 , \9427 , \9428 , \9429_nG3b87 , \9430 , \9431 , \9432 , \9433 , \9434 ,
         \9435 , \9436 , \9437_nG3b8f , \9438 , \9439 , \9440 , \9441 , \9442 , \9443 , \9444 ,
         \9445 , \9446_nG3b98 , \9447 , \9448 , \9449 , \9450 , \9451 , \9452 , \9453 , \9454 ,
         \9455_nG3ba1 , \9456 , \9457 , \9458 , \9459 , \9460 , \9461 , \9462 , \9463 , \9464_nG3baa ,
         \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471 , \9472 , \9473_nG3bb3 , \9474 ,
         \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 , \9482_nG3bbc , \9483 , \9484 ,
         \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491_nG3bc5 , \9492 , \9493 , \9494 ,
         \9495 , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 , \9502_nG3bd0 , \9503 , \9504 ,
         \9505 , \9506 , \9507 , \9508 , \9509 , \9510_nG3bd8 , \9511 , \9512 , \9513 , \9514 ,
         \9515 , \9516 , \9517 , \9518 , \9519_nG3be1 , \9520 , \9521 , \9522 , \9523 , \9524 ,
         \9525 , \9526 , \9527 , \9528_nG3bea , \9529 , \9530 , \9531 , \9532 , \9533 , \9534 ,
         \9535 , \9536 , \9537_nG3bf3 , \9538 , \9539 , \9540 , \9541 , \9542 , \9543 , \9544 ,
         \9545 , \9546_nG3bfc , \9547 , \9548 , \9549 , \9550 , \9551 , \9552 , \9553 , \9554 ,
         \9555_nG3c05 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 , \9562 , \9563 , \9564_nG3c0e ,
         \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 , \9572_nG3c16 , \9573 , \9574 ,
         \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 , \9582 , \9583 , \9584 ,
         \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 , \9592 , \9593 , \9594 ,
         \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 , \9602 , \9603 , \9604 ,
         \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 , \9612 , \9613 , \9614 ,
         \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 , \9622 , \9623 , \9624 ,
         \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 , \9633 , \9634 ,
         \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 , \9643 , \9644 ,
         \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 , \9653 , \9654 ,
         \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 , \9663 , \9664 ,
         \9665 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 , \9672 , \9673 , \9674 ,
         \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 , \9683 , \9684 ,
         \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 , \9693 , \9694 ,
         \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 ,
         \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 ,
         \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 , \9723 , \9724 ,
         \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 , \9733 , \9734 ,
         \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 ,
         \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 ,
         \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 ,
         \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 , \9773 , \9774 ,
         \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 ,
         \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 ,
         \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 ,
         \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 ,
         \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 , \9823 , \9824 ,
         \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 ,
         \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 ,
         \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 ,
         \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 , \9863 , \9864 ,
         \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 ,
         \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 ,
         \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 ,
         \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 ,
         \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 ,
         \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 ,
         \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 ,
         \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 ,
         \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 ,
         \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 ,
         \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974 ,
         \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 ,
         \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 ,
         \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 , \10003 , \10004 ,
         \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 ,
         \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 , \10023 , \10024 ,
         \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 ,
         \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 ,
         \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 ,
         \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 , \10062 , \10063 , \10064 ,
         \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 ,
         \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 , \10083 , \10084 ,
         \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 , \10093 , \10094 ,
         \10095 , \10096 , \10097 , \10098 , \10099_nG3e2d , \10100 , \10101 , \10102 , \10103 , \10104 ,
         \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 ,
         \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 ,
         \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 , \10132 , \10133 , \10134 ,
         \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 ,
         \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 , \10153 , \10154 ,
         \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 ,
         \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 ,
         \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 ,
         \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 ,
         \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 ,
         \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 , \10212 , \10213 , \10214 ,
         \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 ,
         \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 ,
         \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 , \10243 , \10244 ,
         \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 ,
         \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 , \10262 , \10263 , \10264 ,
         \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 ,
         \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 ,
         \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 , \10292 , \10293 , \10294 ,
         \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 ,
         \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 ,
         \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 ,
         \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 ,
         \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 , \10343 , \10344 ,
         \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 ,
         \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 ,
         \10365 , \10366 , \10367 , \10368 , \10369 , \10370 , \10371 , \10372 , \10373 , \10374 ,
         \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 ,
         \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 ,
         \10395 , \10396 , \10397 , \10398 , \10399 , \10400 , \10401 , \10402 , \10403 , \10404 ,
         \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 , \10413 , \10414 ,
         \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 , \10422 , \10423 , \10424 ,
         \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 ,
         \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444 ,
         \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 ,
         \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 ,
         \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 ,
         \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 ,
         \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 ,
         \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504 ,
         \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 ,
         \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 ,
         \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 , \10532 , \10533 , \10534 ,
         \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 ,
         \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 , \10553 , \10554 ,
         \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 , \10563 , \10564 ,
         \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 ,
         \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 ,
         \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 , \10593 , \10594 ,
         \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 ,
         \10605 , \10606 , \10607 , \10608 , \10609 , \10610_nG402c , \10611 , \10612 , \10613 , \10614 ,
         \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 ,
         \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631_nG4041 , \10632 , \10633 , \10634 ,
         \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 ,
         \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 , \10653_nG4057 , \10654 ,
         \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 ,
         \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 ,
         \10675_nG406d , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 , \10682 , \10683 , \10684 ,
         \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 ,
         \10695 , \10696 , \10697_nG4083 , \10698 , \10699 , \10700 , \10701 , \10702 , \10703 , \10704 ,
         \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 , \10712 , \10713 , \10714 ,
         \10715 , \10716 , \10717 , \10718 , \10719_nG4099 , \10720 , \10721 , \10722 , \10723 , \10724 ,
         \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 ,
         \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741_nG40af , \10742 , \10743 , \10744 ,
         \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 ,
         \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 , \10763_nG40c5 , \10764 ,
         \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 ,
         \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 , \10783 , \10784 ,
         \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 ,
         \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 , \10802 , \10803 , \10804 ,
         \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 ,
         \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 ,
         \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 ,
         \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 ,
         \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 , \10853 , \10854 ,
         \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 ,
         \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 ,
         \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 ,
         \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 ,
         \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 ,
         \10905 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 , \10912 , \10913 , \10914 ,
         \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 ,
         \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 , \10932 , \10933 , \10934 ,
         \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 ,
         \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 ,
         \10955 , \10956 , \10957 , \10958 , \10959 , \10960 , \10961 , \10962 , \10963 , \10964 ,
         \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 ,
         \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 , \10982 , \10983 , \10984 ,
         \10985 , \10986 , \10987 , \10988 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 ,
         \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 ,
         \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 , \11012 , \11013 , \11014 ,
         \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 ,
         \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 ,
         \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 , \11042 , \11043 , \11044 ,
         \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 ,
         \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 ,
         \11065 , \11066 , \11067 , \11068 , \11069 , \11070 , \11071 , \11072 , \11073 , \11074 ,
         \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 ,
         \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 , \11092 , \11093 , \11094 ,
         \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 ,
         \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 ,
         \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 , \11122 , \11123 , \11124 ,
         \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 , \11132 , \11133 , \11134 ,
         \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 ,
         \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 ,
         \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 ,
         \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 , \11172 , \11173 , \11174 ,
         \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 ,
         \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 ,
         \11195 , \11196 , \11197 , \11198 , \11199 , \11200 , \11201 , \11202 , \11203 , \11204 ,
         \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 ,
         \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 ,
         \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 ,
         \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 , \11242 , \11243 , \11244 ,
         \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 ,
         \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 ,
         \11265 , \11266 , \11267 , \11268 , \11269 , \11270 , \11271 , \11272 , \11273 , \11274 ,
         \11275 , \11276 , \11277 , \11278 , \11279_nG42c9 , \11280 , \11281 , \11282 , \11283 , \11284 ,
         \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 , \11292 , \11293 , \11294 ,
         \11295 , \11296 , \11297 , \11298 , \11299 , \11300_nG42de , \11301 , \11302 , \11303 , \11304 ,
         \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 ,
         \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 , \11322_nG42f4 , \11323 , \11324 ,
         \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 ,
         \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 , \11342 , \11343 , \11344_nG430a ,
         \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 ,
         \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 ,
         \11365 , \11366_nG4320 , \11367 , \11368 , \11369 , \11370 , \11371 , \11372 , \11373 , \11374 ,
         \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 ,
         \11385 , \11386 , \11387 , \11388_nG4336 , \11389 , \11390 , \11391 , \11392 , \11393 , \11394 ,
         \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 , \11402 , \11403 , \11404 ,
         \11405 , \11406 , \11407 , \11408 , \11409 , \11410_nG434c , \11411 , \11412 , \11413 , \11414 ,
         \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 ,
         \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 , \11432_nG4362 , \11433 , \11434 ,
         \11435 , \11436 , \11437 , \11438 , \11439_nG4369 , \11440 , \11441 , \11442 , \11443 , \11444 ,
         \11445 , \11446 , \11447 , \11448 , \11449 , \11450_nG4374 , \11451 , \11452 , \11453 , \11454 ,
         \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 , \11462 , \11463 , \11464 ,
         \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 , \11472 , \11473 , \11474 ,
         \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 , \11482 , \11483 , \11484 ,
         \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 , \11492 , \11493 , \11494 ,
         \11495_nG43a1 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 , \11502 , \11503_nG43a9 , \11504 ,
         \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 , \11512_nG43b2 , \11513 , \11514 ,
         \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 , \11522_nG43bc , \11523 , \11524 ,
         \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 , \11532_nG43c6 , \11533 , \11534 ,
         \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 , \11542_nG43d0 , \11543 , \11544 ,
         \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 , \11552_nG43da , \11553 , \11554 ,
         \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 , \11562_nG43e4 , \11563 , \11564 ,
         \11565 , \11566 , \11567 , \11568 , \11569 , \11570 , \11571 , \11572_nG43ee , \11573 , \11574 ,
         \11575 , \11576 , \11577 , \11578 , \11579 , \11580 , \11581 , \11582 , \11583 , \11584_nG43fa ,
         \11585 , \11586 , \11587 , \11588 , \11589 , \11590 , \11591 , \11592 , \11593_nG4403 , \11594 ,
         \11595 , \11596 , \11597 , \11598 , \11599 , \11600 , \11601 , \11602 , \11603_nG440d , \11604 ,
         \11605 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 , \11612 , \11613_nG4417 , \11614 ,
         \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 , \11622 , \11623_nG4421 , \11624 ,
         \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 , \11632 , \11633_nG442b , \11634 ,
         \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 , \11642 , \11643_nG4435 , \11644 ,
         \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 , \11652 , \11653_nG443f , \11654 ,
         \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661_nG4447 , \11662 , \11663 , \11664 ,
         \11665 , \11666 , \11667 , \11668 , \11669 , \11670 , \11671 , \11672 , \11673 , \11674 ,
         \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 ,
         \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 , \11692 , \11693 , \11694 ,
         \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 , \11702 , \11703 , \11704 ,
         \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 ,
         \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 ,
         \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 , \11732 , \11733 , \11734 ,
         \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 ,
         \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 ,
         \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 , \11762 , \11763 , \11764 ,
         \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 ,
         \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 , \11782 , \11783 , \11784 ,
         \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 ,
         \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 , \11802 , \11803 , \11804 ,
         \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 , \11812 , \11813 , \11814 ,
         \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 , \11822 , \11823 , \11824 ,
         \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 , \11832 , \11833 , \11834 ,
         \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 , \11842 , \11843 , \11844 ,
         \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 ,
         \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 ,
         \11865 , \11866 , \11867 , \11868 , \11869 , \11870 , \11871 , \11872 , \11873 , \11874 ,
         \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 , \11882 , \11883 , \11884 ,
         \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 , \11892 , \11893 , \11894 ,
         \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 ,
         \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 ,
         \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 , \11922 , \11923 , \11924 ,
         \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 ,
         \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 ,
         \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 , \11952 , \11953 , \11954 ,
         \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 ,
         \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 , \11972 , \11973 , \11974 ,
         \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 , \11982 , \11983 , \11984 ,
         \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 ,
         \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 , \12002 , \12003 , \12004 ,
         \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 , \12012 , \12013 , \12014 ,
         \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 ,
         \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 , \12032 , \12033 , \12034 ,
         \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 , \12042 , \12043 , \12044 ,
         \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 ,
         \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 ,
         \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 , \12072 , \12073 , \12074 ,
         \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 , \12082 , \12083 , \12084 ,
         \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 , \12092 , \12093 , \12094 ,
         \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 , \12102 , \12103 , \12104 ,
         \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 , \12112 , \12113 , \12114 ,
         \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 ,
         \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 , \12132 , \12133 , \12134 ,
         \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 , \12142 , \12143 , \12144 ,
         \12145 , \12146 , \12147 , \12148 , \12149 , \12150 , \12151 , \12152 , \12153 , \12154 ,
         \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 , \12162 , \12163 , \12164 ,
         \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 , \12172 , \12173 , \12174 ,
         \12175 , \12176 , \12177 , \12178 , \12179 , \12180 , \12181 , \12182 , \12183 , \12184 ,
         \12185 , \12186 , \12187 , \12188_nG465e , \12189 , \12190 , \12191 , \12192 , \12193 , \12194 ,
         \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 ,
         \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 , \12212 , \12213 , \12214 ,
         \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 , \12222 , \12223 , \12224 ,
         \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 ,
         \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 , \12242 , \12243 , \12244 ,
         \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 , \12252 , \12253 , \12254 ,
         \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 ,
         \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 , \12272 , \12273 , \12274 ,
         \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 ,
         \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 ,
         \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 ,
         \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 , \12312 , \12313 , \12314 ,
         \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 , \12322 , \12323 , \12324 ,
         \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 ,
         \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 ,
         \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 , \12352 , \12353 , \12354 ,
         \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 ,
         \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 , \12372 , \12373 , \12374 ,
         \12375 , \12376 , \12377 , \12378 , \12379 , \12380 , \12381 , \12382 , \12383 , \12384 ,
         \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 ,
         \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 ,
         \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 ,
         \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 ,
         \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 , \12432 , \12433 , \12434 ,
         \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 , \12442 , \12443 , \12444 ,
         \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 , \12452 , \12453 , \12454 ,
         \12455 , \12456 , \12457 , \12458 , \12459 , \12460 , \12461 , \12462 , \12463 , \12464 ,
         \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 , \12472 , \12473 , \12474 ,
         \12475 , \12476 , \12477 , \12478 , \12479 , \12480 , \12481 , \12482 , \12483 , \12484 ,
         \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 ,
         \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12504 ,
         \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 ,
         \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 ,
         \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 ,
         \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 , \12542 , \12543 , \12544 ,
         \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 , \12552 , \12553 , \12554 ,
         \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 ,
         \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 ,
         \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 ,
         \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 ,
         \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 ,
         \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 ,
         \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 , \12622 , \12623 , \12624 ,
         \12625 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 , \12633 , \12634 ,
         \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 ,
         \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 ,
         \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 ,
         \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 ,
         \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 ,
         \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 , \12693 , \12694 ,
         \12695 , \12696 , \12697 , \12698 , \12699_nG485d , \12700 , \12701 , \12702 , \12703 , \12704 ,
         \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 ,
         \12715 , \12716 , \12717 , \12718 , \12719 , \12720_nG4872 , \12721 , \12722 , \12723 , \12724 ,
         \12725 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 ,
         \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742_nG4888 , \12743 , \12744 ,
         \12745 , \12746 , \12747 , \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 ,
         \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764_nG489e ,
         \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 , \12772 , \12773 , \12774 ,
         \12775 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 ,
         \12785 , \12786_nG48b4 , \12787 , \12788 , \12789 , \12790 , \12791 , \12792 , \12793 , \12794 ,
         \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801 , \12802 , \12803 , \12804 ,
         \12805 , \12806 , \12807 , \12808_nG48ca , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 ,
         \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 ,
         \12825 , \12826 , \12827 , \12828 , \12829 , \12830_nG48e0 , \12831 , \12832 , \12833 , \12834 ,
         \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844 ,
         \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851 , \12852_nG48f6 , \12853 , \12854 ,
         \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 ,
         \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 ,
         \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 , \12883 , \12884 ,
         \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 ,
         \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 ,
         \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 ,
         \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 ,
         \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 ,
         \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 ,
         \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 , \12952 , \12953 , \12954 ,
         \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 ,
         \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 ,
         \12975 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 ,
         \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 ,
         \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 ,
         \13005 , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 ,
         \13015 , \13016 , \13017 , \13018 , \13019 , \13020 , \13021 , \13022 , \13023 , \13024 ,
         \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 ,
         \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 ,
         \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 ,
         \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 , \13062 , \13063 , \13064 ,
         \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 , \13072 , \13073 , \13074 ,
         \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 , \13082 , \13083 , \13084 ,
         \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 , \13092 , \13093 , \13094 ,
         \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 , \13102 , \13103 , \13104 ,
         \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 ,
         \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 ,
         \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 ,
         \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 , \13142 , \13143 , \13144 ,
         \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 ,
         \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 , \13163 , \13164 ,
         \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 ,
         \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 , \13182 , \13183 , \13184 ,
         \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 ,
         \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 ,
         \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 , \13212 , \13213 , \13214 ,
         \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 ,
         \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 ,
         \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 ,
         \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 ,
         \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 ,
         \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 ,
         \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 ,
         \13285 , \13286 , \13287 , \13288 , \13289 , \13290 , \13291 , \13292 , \13293 , \13294 ,
         \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 ,
         \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 , \13312 , \13313 , \13314 ,
         \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 , \13322 , \13323 , \13324 ,
         \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 ,
         \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 ,
         \13345 , \13346 , \13347 , \13348 , \13349 , \13350 , \13351 , \13352 , \13353 , \13354 ,
         \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 , \13362 , \13363 , \13364 ,
         \13365 , \13366 , \13367 , \13368_nG4afa , \13369 , \13370 , \13371 , \13372 , \13373 , \13374 ,
         \13375 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 , \13382 , \13383 , \13384 ,
         \13385 , \13386 , \13387 , \13388 , \13389_nG4b0f , \13390 , \13391 , \13392 , \13393 , \13394 ,
         \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 , \13403 , \13404 ,
         \13405 , \13406 , \13407 , \13408 , \13409 , \13410 , \13411_nG4b25 , \13412 , \13413 , \13414 ,
         \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 ,
         \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 , \13432 , \13433_nG4b3b , \13434 ,
         \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 ,
         \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 ,
         \13455_nG4b51 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 ,
         \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 , \13473 , \13474 ,
         \13475 , \13476 , \13477_nG4b67 , \13478 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 ,
         \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 ,
         \13495 , \13496 , \13497 , \13498 , \13499_nG4b7d , \13500 , \13501 , \13502 , \13503 , \13504 ,
         \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 ,
         \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521_nG4b93 , \13522 , \13523 , \13524 ,
         \13525 , \13526 , \13527 , \13528_nG4b9a , \13529 , \13530 , \13531 , \13532 , \13533 , \13534 ,
         \13535 , \13536 , \13537 , \13538 , \13539_nG4ba5 , \13540 , \13541 , \13542 , \13543 , \13544 ,
         \13545 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 ,
         \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 ,
         \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 ,
         \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 , \13582_nG4bd2 , \13583 , \13584 ,
         \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591_nG4bdb , \13592 , \13593 , \13594 ,
         \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601_nG4be5 , \13602 , \13603 , \13604 ,
         \13605 , \13606 , \13607 , \13608 , \13609 , \13610 , \13611 , \13612_nG4bf0 , \13613 , \13614 ,
         \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 , \13622 , \13623_nG4bfb , \13624 ,
         \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634_nG4c06 ,
         \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 ,
         \13645_nG4c11 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 , \13652 , \13653 , \13654 ,
         \13655 , \13656_nG4c1c , \13657 , \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 ,
         \13665 , \13666 , \13667_nG4c27 , \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 ,
         \13675 , \13676 , \13677 , \13678 , \13679 , \13680_nG4c34 , \13681 , \13682 , \13683 , \13684 ,
         \13685 , \13686 , \13687 , \13688 , \13689 , \13690_nG4c3e , \13691 , \13692 , \13693 , \13694 ,
         \13695 , \13696 , \13697 , \13698 , \13699 , \13700 , \13701_nG4c49 , \13702 , \13703 , \13704 ,
         \13705 , \13706 , \13707 , \13708 , \13709 , \13710 , \13711 , \13712_nG4c54 , \13713 , \13714 ,
         \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 , \13722 , \13723_nG4c5f , \13724 ,
         \13725 , \13726 , \13727 , \13728 , \13729 , \13730 , \13731 , \13732 , \13733 , \13734_nG4c6a ,
         \13735 , \13736 , \13737 , \13738 , \13739 , \13740 , \13741 , \13742 , \13743 , \13744 ,
         \13745_nG4c75 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 , \13752 , \13753 , \13754 ,
         \13755 , \13756_nG4c80 , \13757 , \13758 , \13759 , \13760 , \13761 , \13762 , \13763 , \13764_nG4c88 ,
         \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 ,
         \13775 , \13776 , \13777 , \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 ,
         \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 ,
         \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 , \13802 , \13803 , \13804 ,
         \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 , \13812 , \13813 , \13814 ,
         \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 , \13822 , \13823 , \13824 ,
         \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 ,
         \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 ,
         \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 , \13852 , \13853 , \13854 ,
         \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 , \13862 , \13863 , \13864 ,
         \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 ,
         \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 ,
         \13885 , \13886 , \13887 , \13888 , \13889 , \13890 , \13891 , \13892 , \13893 , \13894 ,
         \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 ,
         \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 ,
         \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 ,
         \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 ,
         \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 , \13942 , \13943 , \13944 ,
         \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 ,
         \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 ,
         \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 , \13972 , \13973 , \13974 ,
         \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 ,
         \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 ,
         \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 ,
         \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 ,
         \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 , \14022 , \14023 , \14024 ,
         \14025 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 , \14032 , \14033 , \14034 ,
         \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 , \14042 , \14043 , \14044 ,
         \14045 , \14046 , \14047 , \14048 , \14049 , \14050 , \14051 , \14052 , \14053 , \14054 ,
         \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 , \14062 , \14063 , \14064 ,
         \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 , \14072 , \14073 , \14074 ,
         \14075 , \14076 , \14077 , \14078 , \14079 , \14080 , \14081 , \14082 , \14083 , \14084 ,
         \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 ,
         \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 ,
         \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 ,
         \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 ,
         \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 , \14132 , \14133 , \14134 ,
         \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 , \14142 , \14143 , \14144 ,
         \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 ,
         \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 , \14162 , \14163 , \14164 ,
         \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 , \14172 , \14173 , \14174 ,
         \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 ,
         \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 ,
         \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 ,
         \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 , \14212 , \14213 , \14214 ,
         \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 ,
         \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 ,
         \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 ,
         \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 , \14252 , \14253 , \14254 ,
         \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 ,
         \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 ,
         \14275 , \14276 , \14277 , \14278 , \14279 , \14280 , \14281 , \14282 , \14283 , \14284 ,
         \14285 , \14286 , \14287 , \14288 , \14289 , \14290 , \14291_nG4e9f , \14292 , \14293 , \14294 ,
         \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 ,
         \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 ,
         \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 , \14322 , \14323 , \14324 ,
         \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 ,
         \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 , \14342 , \14343 , \14344 ,
         \14345 , \14346 , \14347 , \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 ,
         \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 ,
         \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 , \14372 , \14373 , \14374 ,
         \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 ,
         \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 ,
         \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 , \14402 , \14403 , \14404 ,
         \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 , \14412 , \14413 , \14414 ,
         \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 ,
         \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 ,
         \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 ,
         \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 , \14452 , \14453 , \14454 ,
         \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 ,
         \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 ,
         \14475 , \14476 , \14477 , \14478 , \14479 , \14480 , \14481 , \14482 , \14483 , \14484 ,
         \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 ,
         \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 ,
         \14505 , \14506 , \14507 , \14508 , \14509 , \14510 , \14511 , \14512 , \14513 , \14514 ,
         \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 ,
         \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 ,
         \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 , \14542 , \14543 , \14544 ,
         \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 ,
         \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 , \14562 , \14563 , \14564 ,
         \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 , \14572 , \14573 , \14574 ,
         \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 , \14582 , \14583 , \14584 ,
         \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 , \14592 , \14593 , \14594 ,
         \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 , \14602 , \14603 , \14604 ,
         \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 , \14612 , \14613 , \14614 ,
         \14615 , \14616 , \14617 , \14618 , \14619 , \14620 , \14621 , \14622 , \14623 , \14624 ,
         \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 , \14632 , \14633 , \14634 ,
         \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 , \14642 , \14643 , \14644 ,
         \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 , \14652 , \14653 , \14654 ,
         \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 , \14662 , \14663 , \14664 ,
         \14665 , \14666 , \14667 , \14668 , \14669 , \14670 , \14671 , \14672 , \14673 , \14674 ,
         \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 , \14682 , \14683 , \14684 ,
         \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 , \14692 , \14693 , \14694 ,
         \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 , \14702 , \14703 , \14704 ,
         \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 , \14712 , \14713 , \14714 ,
         \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 , \14722 , \14723 , \14724 ,
         \14725 , \14726 , \14727 , \14728 , \14729 , \14730 , \14731 , \14732 , \14733 , \14734 ,
         \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 , \14742 , \14743 , \14744 ,
         \14745 , \14746 , \14747 , \14748 , \14749 , \14750 , \14751 , \14752 , \14753 , \14754 ,
         \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 , \14762 , \14763 , \14764 ,
         \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 , \14772 , \14773 , \14774 ,
         \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 , \14782 , \14783 , \14784 ,
         \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14791 , \14792 , \14793 , \14794 ,
         \14795 , \14796 , \14797 , \14798 , \14799 , \14800 , \14801 , \14802_nG509e , \14803 , \14804 ,
         \14805 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 , \14812 , \14813 , \14814 ,
         \14815 , \14816 , \14817 , \14818 , \14819 , \14820 , \14821 , \14822 , \14823_nG50b3 , \14824 ,
         \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831 , \14832 , \14833 , \14834 ,
         \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 , \14842 , \14843 , \14844 ,
         \14845_nG50c9 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 , \14852 , \14853 , \14854 ,
         \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 , \14862 , \14863 , \14864 ,
         \14865 , \14866 , \14867_nG50df , \14868 , \14869 , \14870 , \14871 , \14872 , \14873 , \14874 ,
         \14875 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 , \14882 , \14883 , \14884 ,
         \14885 , \14886 , \14887 , \14888 , \14889_nG50f5 , \14890 , \14891 , \14892 , \14893 , \14894 ,
         \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 , \14902 , \14903 , \14904 ,
         \14905 , \14906 , \14907 , \14908 , \14909 , \14910 , \14911_nG510b , \14912 , \14913 , \14914 ,
         \14915 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 , \14922 , \14923 , \14924 ,
         \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 , \14932 , \14933_nG5121 , \14934 ,
         \14935 , \14936 , \14937 , \14938 , \14939 , \14940 , \14941 , \14942 , \14943 , \14944 ,
         \14945 , \14946 , \14947 , \14948 , \14949 , \14950 , \14951 , \14952 , \14953 , \14954 ,
         \14955_nG5137 , \14956 , \14957 , \14958 , \14959 , \14960 , \14961 , \14962 , \14963 , \14964 ,
         \14965 , \14966 , \14967 , \14968 , \14969 , \14970 , \14971 , \14972 , \14973 , \14974 ,
         \14975 , \14976 , \14977 , \14978 , \14979 , \14980 , \14981 , \14982 , \14983 , \14984 ,
         \14985 , \14986 , \14987 , \14988 , \14989 , \14990 , \14991 , \14992 , \14993 , \14994 ,
         \14995 , \14996 , \14997 , \14998 , \14999 , \15000 , \15001 , \15002 , \15003 , \15004 ,
         \15005 , \15006 , \15007 , \15008 , \15009 , \15010 , \15011 , \15012 , \15013 , \15014 ,
         \15015 , \15016 , \15017 , \15018 , \15019 , \15020 , \15021 , \15022 , \15023 , \15024 ,
         \15025 , \15026 , \15027 , \15028 , \15029 , \15030 , \15031 , \15032 , \15033 , \15034 ,
         \15035 , \15036 , \15037 , \15038 , \15039 , \15040 , \15041 , \15042 , \15043 , \15044 ,
         \15045 , \15046 , \15047 , \15048 , \15049 , \15050 , \15051 , \15052 , \15053 , \15054 ,
         \15055 , \15056 , \15057 , \15058 , \15059 , \15060 , \15061 , \15062 , \15063 , \15064 ,
         \15065 , \15066 , \15067 , \15068 , \15069 , \15070 , \15071 , \15072 , \15073 , \15074 ,
         \15075 , \15076 , \15077 , \15078 , \15079 , \15080 , \15081 , \15082 , \15083 , \15084 ,
         \15085 , \15086 , \15087 , \15088 , \15089 , \15090 , \15091 , \15092 , \15093 , \15094 ,
         \15095 , \15096 , \15097 , \15098 , \15099 , \15100 , \15101 , \15102 , \15103 , \15104 ,
         \15105 , \15106 , \15107 , \15108 , \15109 , \15110 , \15111 , \15112 , \15113 , \15114 ,
         \15115 , \15116 , \15117 , \15118 , \15119 , \15120 , \15121 , \15122 , \15123 , \15124 ,
         \15125 , \15126 , \15127 , \15128 , \15129 , \15130 , \15131 , \15132 , \15133 , \15134 ,
         \15135 , \15136 , \15137 , \15138 , \15139 , \15140 , \15141 , \15142 , \15143 , \15144 ,
         \15145 , \15146 , \15147 , \15148 , \15149 , \15150 , \15151 , \15152 , \15153 , \15154 ,
         \15155 , \15156 , \15157 , \15158 , \15159 , \15160 , \15161 , \15162 , \15163 , \15164 ,
         \15165 , \15166 , \15167 , \15168 , \15169 , \15170 , \15171 , \15172 , \15173 , \15174 ,
         \15175 , \15176 , \15177 , \15178 , \15179 , \15180 , \15181 , \15182 , \15183 , \15184 ,
         \15185 , \15186 , \15187 , \15188 , \15189 , \15190 , \15191 , \15192 , \15193 , \15194 ,
         \15195 , \15196 , \15197 , \15198 , \15199 , \15200 , \15201 , \15202 , \15203 , \15204 ,
         \15205 , \15206 , \15207 , \15208 , \15209 , \15210 , \15211 , \15212 , \15213 , \15214 ,
         \15215 , \15216 , \15217 , \15218 , \15219 , \15220 , \15221 , \15222 , \15223 , \15224 ,
         \15225 , \15226 , \15227 , \15228 , \15229 , \15230 , \15231 , \15232 , \15233 , \15234 ,
         \15235 , \15236 , \15237 , \15238 , \15239 , \15240 , \15241 , \15242 , \15243 , \15244 ,
         \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 , \15252 , \15253 , \15254 ,
         \15255 , \15256 , \15257 , \15258 , \15259 , \15260 , \15261 , \15262 , \15263 , \15264 ,
         \15265 , \15266 , \15267 , \15268 , \15269 , \15270 , \15271 , \15272 , \15273 , \15274 ,
         \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 , \15282 , \15283 , \15284 ,
         \15285 , \15286 , \15287 , \15288 , \15289 , \15290 , \15291 , \15292 , \15293 , \15294 ,
         \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 , \15302 , \15303 , \15304 ,
         \15305 , \15306 , \15307 , \15308 , \15309 , \15310 , \15311 , \15312 , \15313 , \15314 ,
         \15315 , \15316 , \15317 , \15318 , \15319 , \15320 , \15321 , \15322 , \15323 , \15324 ,
         \15325 , \15326 , \15327 , \15328 , \15329 , \15330 , \15331 , \15332 , \15333 , \15334 ,
         \15335 , \15336 , \15337 , \15338 , \15339 , \15340 , \15341 , \15342 , \15343 , \15344 ,
         \15345 , \15346 , \15347 , \15348 , \15349 , \15350 , \15351 , \15352 , \15353 , \15354 ,
         \15355 , \15356 , \15357 , \15358 , \15359 , \15360 , \15361 , \15362 , \15363 , \15364 ,
         \15365 , \15366 , \15367 , \15368 , \15369 , \15370 , \15371 , \15372 , \15373 , \15374 ,
         \15375 , \15376 , \15377 , \15378 , \15379 , \15380 , \15381 , \15382 , \15383 , \15384 ,
         \15385 , \15386 , \15387 , \15388 , \15389 , \15390 , \15391 , \15392 , \15393 , \15394 ,
         \15395 , \15396 , \15397 , \15398 , \15399 , \15400 , \15401 , \15402 , \15403 , \15404 ,
         \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411 , \15412 , \15413 , \15414 ,
         \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 , \15422 , \15423 , \15424 ,
         \15425 , \15426 , \15427 , \15428 , \15429 , \15430 , \15431 , \15432 , \15433 , \15434 ,
         \15435 , \15436 , \15437 , \15438 , \15439 , \15440 , \15441 , \15442 , \15443 , \15444 ,
         \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 , \15452 , \15453 , \15454 ,
         \15455 , \15456 , \15457 , \15458 , \15459 , \15460 , \15461 , \15462 , \15463 , \15464 ,
         \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15471_nG533b , \15472 , \15473 , \15474 ,
         \15475 , \15476 , \15477 , \15478 , \15479 , \15480 , \15481 , \15482 , \15483 , \15484 ,
         \15485 , \15486 , \15487 , \15488 , \15489 , \15490 , \15491 , \15492_nG5350 , \15493 , \15494 ,
         \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 , \15502 , \15503 , \15504 ,
         \15505 , \15506 , \15507 , \15508 , \15509 , \15510 , \15511 , \15512 , \15513 , \15514_nG5366 ,
         \15515 , \15516 , \15517 , \15518 , \15519 , \15520 , \15521 , \15522 , \15523 , \15524 ,
         \15525 , \15526 , \15527 , \15528 , \15529 , \15530 , \15531 , \15532 , \15533 , \15534 ,
         \15535 , \15536_nG537c , \15537 , \15538 , \15539 , \15540 , \15541 , \15542 , \15543 , \15544 ,
         \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 , \15552 , \15553 , \15554 ,
         \15555 , \15556 , \15557 , \15558_nG5392 , \15559 , \15560 , \15561 , \15562 , \15563 , \15564 ,
         \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 , \15572 , \15573 , \15574 ,
         \15575 , \15576 , \15577 , \15578 , \15579 , \15580_nG53a8 , \15581 , \15582 , \15583 , \15584 ,
         \15585 , \15586 , \15587 , \15588 , \15589 , \15590 , \15591 , \15592 , \15593 , \15594 ,
         \15595 , \15596 , \15597 , \15598 , \15599 , \15600 , \15601 , \15602_nG53be , \15603 , \15604 ,
         \15605 , \15606 , \15607 , \15608 , \15609 , \15610 , \15611 , \15612 , \15613 , \15614 ,
         \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 , \15622 , \15623 , \15624_nG53d4 ,
         \15625 , \15626 , \15627 , \15628 , \15629 , \15630 , \15631_nG53db , \15632 , \15633 , \15634 ,
         \15635 , \15636 , \15637 , \15638 , \15639 , \15640 , \15641 , \15642_nG53e6 , \15643 , \15644 ,
         \15645 , \15646 , \15647 , \15648 , \15649 , \15650 , \15651 , \15652 , \15653 , \15654 ,
         \15655 , \15656 , \15657 , \15658 , \15659 , \15660 , \15661 , \15662 , \15663 , \15664 ,
         \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 , \15672 , \15673 , \15674 ,
         \15675 , \15676 , \15677 , \15678 , \15679 , \15680 , \15681 , \15682 , \15683 , \15684 ,
         \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 , \15692_nG5418 , \15693 , \15694 ,
         \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 , \15702_nG5422 , \15703 , \15704 ,
         \15705 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 , \15712 , \15713_nG542d , \15714 ,
         \15715 , \15716 , \15717 , \15718 , \15719 , \15720 , \15721 , \15722 , \15723 , \15724 ,
         \15725_nG5439 , \15726 , \15727 , \15728 , \15729 , \15730 , \15731 , \15732 , \15733 , \15734 ,
         \15735 , \15736 , \15737_nG5445 , \15738 , \15739 , \15740 , \15741 , \15742 , \15743 , \15744 ,
         \15745 , \15746 , \15747 , \15748 , \15749_nG5451 , \15750 , \15751 , \15752 , \15753 , \15754 ,
         \15755 , \15756 , \15757 , \15758 , \15759 , \15760 , \15761_nG545d , \15762 , \15763 , \15764 ,
         \15765 , \15766 , \15767 , \15768 , \15769 , \15770 , \15771 , \15772 , \15773_nG5469 , \15774 ,
         \15775 , \15776 , \15777 , \15778 , \15779 , \15780 , \15781 , \15782 , \15783 , \15784 ,
         \15785_nG5475 , \15786 , \15787 , \15788 , \15789 , \15790 , \15791 , \15792 , \15793 , \15794 ,
         \15795 , \15796 , \15797 , \15798 , \15799_nG5483 , \15800 , \15801 , \15802 , \15803 , \15804 ,
         \15805 , \15806 , \15807 , \15808 , \15809 , \15810_nG548e , \15811 , \15812 , \15813 , \15814 ,
         \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , \15821 , \15822_nG549a , \15823 , \15824 ,
         \15825 , \15826 , \15827 , \15828 , \15829 , \15830 , \15831 , \15832 , \15833 , \15834_nG54a6 ,
         \15835 , \15836 , \15837 , \15838 , \15839 , \15840 , \15841 , \15842 , \15843 , \15844 ,
         \15845 , \15846_nG54b2 , \15847 , \15848 , \15849 , \15850 , \15851 , \15852 , \15853 , \15854 ,
         \15855 , \15856 , \15857 , \15858_nG54be , \15859 , \15860 , \15861 , \15862 , \15863 , \15864 ,
         \15865 , \15866 , \15867 , \15868 , \15869 , \15870_nG54ca , \15871 , \15872 , \15873 , \15874 ,
         \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 , \15882_nG54d6 , \15883 , \15884 ,
         \15885 , \15886 , \15887 , \15888 , \15889 , \15890_nG54de , \15891 , \15892 , \15893 , \15894 ,
         \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 , \15902 , \15903 , \15904 ,
         \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 , \15912 , \15913 , \15914 ,
         \15915 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 , \15922 , \15923 , \15924 ,
         \15925 , \15926 , \15927 , \15928 , \15929 , \15930 , \15931 , \15932 , \15933 , \15934 ,
         \15935 , \15936 , \15937 , \15938 , \15939 , \15940 , \15941 , \15942 , \15943 , \15944 ,
         \15945 , \15946 , \15947 , \15948 , \15949 , \15950 , \15951 , \15952 , \15953 , \15954 ,
         \15955 , \15956 , \15957 , \15958 , \15959 , \15960 , \15961 , \15962 , \15963 , \15964 ,
         \15965 , \15966 , \15967 , \15968 , \15969 , \15970 , \15971 , \15972 , \15973 , \15974 ,
         \15975 , \15976 , \15977 , \15978 , \15979 , \15980 , \15981 , \15982 , \15983 , \15984 ,
         \15985 , \15986 , \15987 , \15988 , \15989 , \15990 , \15991 , \15992 , \15993 , \15994 ,
         \15995 , \15996 , \15997 , \15998 , \15999 , \16000 , \16001 , \16002 , \16003 , \16004 ,
         \16005 , \16006 , \16007 , \16008 , \16009 , \16010 , \16011 , \16012 , \16013 , \16014 ,
         \16015 , \16016 , \16017 , \16018 , \16019 , \16020 , \16021 , \16022 , \16023 , \16024 ,
         \16025 , \16026 , \16027 , \16028 , \16029 , \16030 , \16031 , \16032 , \16033 , \16034 ,
         \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 , \16042 , \16043 , \16044 ,
         \16045 , \16046 , \16047 , \16048 , \16049 , \16050 , \16051 , \16052 , \16053 , \16054 ,
         \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 , \16062 , \16063 , \16064 ,
         \16065 , \16066 , \16067 , \16068 , \16069 , \16070 , \16071 , \16072 , \16073 , \16074 ,
         \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 , \16082 , \16083 , \16084 ,
         \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 , \16092 , \16093 , \16094 ,
         \16095 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 , \16102 , \16103 , \16104 ,
         \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 , \16112 , \16113 , \16114 ,
         \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 , \16122 , \16123 , \16124 ,
         \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 , \16132 , \16133 , \16134 ,
         \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 , \16142 , \16143 , \16144 ,
         \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 , \16152 , \16153 , \16154 ,
         \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 , \16162 , \16163 , \16164 ,
         \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 , \16172 , \16173 , \16174 ,
         \16175 , \16176 , \16177 , \16178 , \16179 , \16180 , \16181 , \16182 , \16183 , \16184 ,
         \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 , \16192 , \16193 , \16194 ,
         \16195 , \16196 , \16197 , \16198 , \16199 , \16200 , \16201 , \16202 , \16203 , \16204 ,
         \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 , \16212 , \16213 , \16214 ,
         \16215 , \16216 , \16217 , \16218 , \16219 , \16220 , \16221 , \16222 , \16223 , \16224 ,
         \16225 , \16226 , \16227 , \16228 , \16229 , \16230 , \16231 , \16232 , \16233 , \16234 ,
         \16235 , \16236 , \16237 , \16238 , \16239 , \16240 , \16241 , \16242 , \16243 , \16244 ,
         \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 , \16252 , \16253 , \16254 ,
         \16255 , \16256 , \16257 , \16258 , \16259 , \16260 , \16261 , \16262 , \16263 , \16264 ,
         \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 , \16272 , \16273 , \16274 ,
         \16275 , \16276 , \16277 , \16278 , \16279 , \16280 , \16281 , \16282 , \16283 , \16284 ,
         \16285 , \16286 , \16287 , \16288 , \16289 , \16290 , \16291 , \16292 , \16293 , \16294 ,
         \16295 , \16296 , \16297 , \16298 , \16299 , \16300 , \16301 , \16302 , \16303 , \16304 ,
         \16305 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 , \16312 , \16313 , \16314 ,
         \16315 , \16316 , \16317 , \16318 , \16319 , \16320 , \16321 , \16322 , \16323 , \16324 ,
         \16325 , \16326 , \16327 , \16328 , \16329 , \16330 , \16331 , \16332 , \16333 , \16334 ,
         \16335 , \16336 , \16337 , \16338 , \16339 , \16340 , \16341 , \16342 , \16343 , \16344 ,
         \16345 , \16346 , \16347 , \16348 , \16349 , \16350 , \16351 , \16352 , \16353 , \16354 ,
         \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 , \16362 , \16363 , \16364 ,
         \16365 , \16366 , \16367 , \16368 , \16369 , \16370 , \16371 , \16372 , \16373 , \16374 ,
         \16375 , \16376 , \16377 , \16378 , \16379 , \16380 , \16381 , \16382 , \16383 , \16384 ,
         \16385 , \16386 , \16387 , \16388 , \16389 , \16390 , \16391 , \16392 , \16393 , \16394 ,
         \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 , \16402 , \16403 , \16404 ,
         \16405 , \16406 , \16407 , \16408 , \16409 , \16410 , \16411 , \16412 , \16413 , \16414 ,
         \16415 , \16416 , \16417_nG56f5 , \16418 , \16419 , \16420 , \16421 , \16422 , \16423 , \16424 ,
         \16425 , \16426 , \16427 , \16428 , \16429 , \16430 , \16431 , \16432 , \16433 , \16434 ,
         \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 , \16442 , \16443 , \16444 ,
         \16445 , \16446 , \16447 , \16448 , \16449 , \16450 , \16451 , \16452 , \16453 , \16454 ,
         \16455 , \16456 , \16457 , \16458 , \16459 , \16460 , \16461 , \16462 , \16463 , \16464 ,
         \16465 , \16466 , \16467 , \16468 , \16469 , \16470 , \16471 , \16472 , \16473 , \16474 ,
         \16475 , \16476 , \16477 , \16478 , \16479 , \16480 , \16481 , \16482 , \16483 , \16484 ,
         \16485 , \16486 , \16487 , \16488 , \16489 , \16490 , \16491 , \16492 , \16493 , \16494 ,
         \16495 , \16496 , \16497 , \16498 , \16499 , \16500 , \16501 , \16502 , \16503 , \16504 ,
         \16505 , \16506 , \16507 , \16508 , \16509 , \16510 , \16511 , \16512 , \16513 , \16514 ,
         \16515 , \16516 , \16517 , \16518 , \16519 , \16520 , \16521 , \16522 , \16523 , \16524 ,
         \16525 , \16526 , \16527 , \16528 , \16529 , \16530 , \16531 , \16532 , \16533 , \16534 ,
         \16535 , \16536 , \16537 , \16538 , \16539 , \16540 , \16541 , \16542 , \16543 , \16544 ,
         \16545 , \16546 , \16547 , \16548 , \16549 , \16550 , \16551 , \16552 , \16553 , \16554 ,
         \16555 , \16556 , \16557 , \16558 , \16559 , \16560 , \16561 , \16562 , \16563 , \16564 ,
         \16565 , \16566 , \16567 , \16568 , \16569 , \16570 , \16571 , \16572 , \16573 , \16574 ,
         \16575 , \16576 , \16577 , \16578 , \16579 , \16580 , \16581 , \16582 , \16583 , \16584 ,
         \16585 , \16586 , \16587 , \16588 , \16589 , \16590 , \16591 , \16592 , \16593 , \16594 ,
         \16595 , \16596 , \16597 , \16598 , \16599 , \16600 , \16601 , \16602 , \16603 , \16604 ,
         \16605 , \16606 , \16607 , \16608 , \16609 , \16610 , \16611 , \16612 , \16613 , \16614 ,
         \16615 , \16616 , \16617 , \16618 , \16619 , \16620 , \16621 , \16622 , \16623 , \16624 ,
         \16625 , \16626 , \16627 , \16628 , \16629 , \16630 , \16631 , \16632 , \16633 , \16634 ,
         \16635 , \16636 , \16637 , \16638 , \16639 , \16640 , \16641 , \16642 , \16643 , \16644 ,
         \16645 , \16646 , \16647 , \16648 , \16649 , \16650 , \16651 , \16652 , \16653 , \16654 ,
         \16655 , \16656 , \16657 , \16658 , \16659 , \16660 , \16661 , \16662 , \16663 , \16664 ,
         \16665 , \16666 , \16667 , \16668 , \16669 , \16670 , \16671 , \16672 , \16673 , \16674 ,
         \16675 , \16676 , \16677 , \16678 , \16679 , \16680 , \16681 , \16682 , \16683 , \16684 ,
         \16685 , \16686 , \16687 , \16688 , \16689 , \16690 , \16691 , \16692 , \16693 , \16694 ,
         \16695 , \16696 , \16697 , \16698 , \16699 , \16700 , \16701 , \16702 , \16703 , \16704 ,
         \16705 , \16706 , \16707 , \16708 , \16709 , \16710 , \16711 , \16712 , \16713 , \16714 ,
         \16715 , \16716 , \16717 , \16718 , \16719 , \16720 , \16721 , \16722 , \16723 , \16724 ,
         \16725 , \16726 , \16727 , \16728 , \16729 , \16730 , \16731 , \16732 , \16733 , \16734 ,
         \16735 , \16736 , \16737 , \16738 , \16739 , \16740 , \16741 , \16742 , \16743 , \16744 ,
         \16745 , \16746 , \16747 , \16748 , \16749 , \16750 , \16751 , \16752 , \16753 , \16754 ,
         \16755 , \16756 , \16757 , \16758 , \16759 , \16760 , \16761 , \16762 , \16763 , \16764 ,
         \16765 , \16766 , \16767 , \16768 , \16769 , \16770 , \16771 , \16772 , \16773 , \16774 ,
         \16775 , \16776 , \16777 , \16778 , \16779 , \16780 , \16781 , \16782 , \16783 , \16784 ,
         \16785 , \16786 , \16787 , \16788 , \16789 , \16790 , \16791 , \16792 , \16793 , \16794 ,
         \16795 , \16796 , \16797 , \16798 , \16799 , \16800 , \16801 , \16802 , \16803 , \16804 ,
         \16805 , \16806 , \16807 , \16808 , \16809 , \16810 , \16811 , \16812 , \16813 , \16814 ,
         \16815 , \16816 , \16817 , \16818 , \16819 , \16820 , \16821 , \16822 , \16823 , \16824 ,
         \16825 , \16826 , \16827 , \16828 , \16829 , \16830 , \16831 , \16832 , \16833 , \16834 ,
         \16835 , \16836 , \16837 , \16838 , \16839 , \16840 , \16841 , \16842 , \16843 , \16844 ,
         \16845 , \16846 , \16847 , \16848 , \16849 , \16850 , \16851 , \16852 , \16853 , \16854 ,
         \16855 , \16856 , \16857 , \16858 , \16859 , \16860 , \16861 , \16862 , \16863 , \16864 ,
         \16865 , \16866 , \16867 , \16868 , \16869 , \16870 , \16871 , \16872 , \16873 , \16874 ,
         \16875 , \16876 , \16877 , \16878 , \16879 , \16880 , \16881 , \16882 , \16883 , \16884 ,
         \16885 , \16886 , \16887 , \16888 , \16889 , \16890 , \16891 , \16892 , \16893 , \16894 ,
         \16895 , \16896 , \16897 , \16898 , \16899 , \16900 , \16901 , \16902 , \16903 , \16904 ,
         \16905 , \16906 , \16907 , \16908 , \16909 , \16910 , \16911 , \16912 , \16913 , \16914 ,
         \16915 , \16916 , \16917 , \16918 , \16919 , \16920 , \16921 , \16922 , \16923 , \16924 ,
         \16925 , \16926 , \16927 , \16928_nG58f4 , \16929 , \16930 , \16931 , \16932 , \16933 , \16934 ,
         \16935 , \16936 , \16937 , \16938 , \16939 , \16940 , \16941 , \16942 , \16943 , \16944 ,
         \16945 , \16946 , \16947 , \16948 , \16949_nG5909 , \16950 , \16951 , \16952 , \16953 , \16954 ,
         \16955 , \16956 , \16957 , \16958 , \16959 , \16960 , \16961 , \16962 , \16963 , \16964 ,
         \16965 , \16966 , \16967 , \16968 , \16969 , \16970 , \16971_nG591f , \16972 , \16973 , \16974 ,
         \16975 , \16976 , \16977 , \16978 , \16979 , \16980 , \16981 , \16982 , \16983 , \16984 ,
         \16985 , \16986 , \16987 , \16988 , \16989 , \16990 , \16991 , \16992 , \16993_nG5935 , \16994 ,
         \16995 , \16996 , \16997 , \16998 , \16999 , \17000 , \17001 , \17002 , \17003 , \17004 ,
         \17005 , \17006 , \17007 , \17008 , \17009 , \17010 , \17011 , \17012 , \17013 , \17014 ,
         \17015_nG594b , \17016 , \17017 , \17018 , \17019 , \17020 , \17021 , \17022 , \17023 , \17024 ,
         \17025 , \17026 , \17027 , \17028 , \17029 , \17030 , \17031 , \17032 , \17033 , \17034 ,
         \17035 , \17036 , \17037_nG5961 , \17038 , \17039 , \17040 , \17041 , \17042 , \17043 , \17044 ,
         \17045 , \17046 , \17047 , \17048 , \17049 , \17050 , \17051 , \17052 , \17053 , \17054 ,
         \17055 , \17056 , \17057 , \17058 , \17059_nG5977 , \17060 , \17061 , \17062 , \17063 , \17064 ,
         \17065 , \17066 , \17067 , \17068 , \17069 , \17070 , \17071 , \17072 , \17073 , \17074 ,
         \17075 , \17076 , \17077 , \17078 , \17079 , \17080 , \17081_nG598d , \17082 , \17083 , \17084 ,
         \17085 , \17086 , \17087 , \17088 , \17089 , \17090 , \17091 , \17092 , \17093 , \17094 ,
         \17095 , \17096 , \17097 , \17098 , \17099 , \17100 , \17101 , \17102 , \17103 , \17104 ,
         \17105 , \17106 , \17107 , \17108 , \17109 , \17110 , \17111 , \17112 , \17113 , \17114 ,
         \17115 , \17116 , \17117 , \17118 , \17119 , \17120 , \17121 , \17122 , \17123 , \17124 ,
         \17125 , \17126 , \17127 , \17128 , \17129 , \17130 , \17131 , \17132 , \17133 , \17134 ,
         \17135 , \17136 , \17137 , \17138 , \17139 , \17140 , \17141 , \17142 , \17143 , \17144 ,
         \17145 , \17146 , \17147 , \17148 , \17149 , \17150 , \17151 , \17152 , \17153 , \17154 ,
         \17155 , \17156 , \17157 , \17158 , \17159 , \17160 , \17161 , \17162 , \17163 , \17164 ,
         \17165 , \17166 , \17167 , \17168 , \17169 , \17170 , \17171 , \17172 , \17173 , \17174 ,
         \17175 , \17176 , \17177 , \17178 , \17179 , \17180 , \17181 , \17182 , \17183 , \17184 ,
         \17185 , \17186 , \17187 , \17188 , \17189 , \17190 , \17191 , \17192 , \17193 , \17194 ,
         \17195 , \17196 , \17197 , \17198 , \17199 , \17200 , \17201 , \17202 , \17203 , \17204 ,
         \17205 , \17206 , \17207 , \17208 , \17209 , \17210 , \17211 , \17212 , \17213 , \17214 ,
         \17215 , \17216 , \17217 , \17218 , \17219 , \17220 , \17221 , \17222 , \17223 , \17224 ,
         \17225 , \17226 , \17227 , \17228 , \17229 , \17230 , \17231 , \17232 , \17233 , \17234 ,
         \17235 , \17236 , \17237 , \17238 , \17239 , \17240 , \17241 , \17242 , \17243 , \17244 ,
         \17245 , \17246 , \17247 , \17248 , \17249 , \17250 , \17251 , \17252 , \17253 , \17254 ,
         \17255 , \17256 , \17257 , \17258 , \17259 , \17260 , \17261 , \17262 , \17263 , \17264 ,
         \17265 , \17266 , \17267 , \17268 , \17269 , \17270 , \17271 , \17272 , \17273 , \17274 ,
         \17275 , \17276 , \17277 , \17278 , \17279 , \17280 , \17281 , \17282 , \17283 , \17284 ,
         \17285 , \17286 , \17287 , \17288 , \17289 , \17290 , \17291 , \17292 , \17293 , \17294 ,
         \17295 , \17296 , \17297 , \17298 , \17299 , \17300 , \17301 , \17302 , \17303 , \17304 ,
         \17305 , \17306 , \17307 , \17308 , \17309 , \17310 , \17311 , \17312 , \17313 , \17314 ,
         \17315 , \17316 , \17317 , \17318 , \17319 , \17320 , \17321 , \17322 , \17323 , \17324 ,
         \17325 , \17326 , \17327 , \17328 , \17329 , \17330 , \17331 , \17332 , \17333 , \17334 ,
         \17335 , \17336 , \17337 , \17338 , \17339 , \17340 , \17341 , \17342 , \17343 , \17344 ,
         \17345 , \17346 , \17347 , \17348 , \17349 , \17350 , \17351 , \17352 , \17353 , \17354 ,
         \17355 , \17356 , \17357 , \17358 , \17359 , \17360 , \17361 , \17362 , \17363 , \17364 ,
         \17365 , \17366 , \17367 , \17368 , \17369 , \17370 , \17371 , \17372 , \17373 , \17374 ,
         \17375 , \17376 , \17377 , \17378 , \17379 , \17380 , \17381 , \17382 , \17383 , \17384 ,
         \17385 , \17386 , \17387 , \17388 , \17389 , \17390 , \17391 , \17392 , \17393 , \17394 ,
         \17395 , \17396 , \17397 , \17398 , \17399 , \17400 , \17401 , \17402 , \17403 , \17404 ,
         \17405 , \17406 , \17407 , \17408 , \17409 , \17410 , \17411 , \17412 , \17413 , \17414 ,
         \17415 , \17416 , \17417 , \17418 , \17419 , \17420 , \17421 , \17422 , \17423 , \17424 ,
         \17425 , \17426 , \17427 , \17428 , \17429 , \17430 , \17431 , \17432 , \17433 , \17434 ,
         \17435 , \17436 , \17437 , \17438 , \17439 , \17440 , \17441 , \17442 , \17443 , \17444 ,
         \17445 , \17446 , \17447 , \17448 , \17449 , \17450 , \17451 , \17452 , \17453 , \17454 ,
         \17455 , \17456 , \17457 , \17458 , \17459 , \17460 , \17461 , \17462 , \17463 , \17464 ,
         \17465 , \17466 , \17467 , \17468 , \17469 , \17470 , \17471 , \17472 , \17473 , \17474 ,
         \17475 , \17476 , \17477 , \17478 , \17479 , \17480 , \17481 , \17482 , \17483 , \17484 ,
         \17485 , \17486 , \17487 , \17488 , \17489 , \17490 , \17491 , \17492 , \17493 , \17494 ,
         \17495 , \17496 , \17497 , \17498 , \17499 , \17500 , \17501 , \17502 , \17503 , \17504 ,
         \17505 , \17506 , \17507 , \17508 , \17509 , \17510 , \17511 , \17512 , \17513 , \17514 ,
         \17515 , \17516 , \17517 , \17518 , \17519 , \17520 , \17521 , \17522 , \17523 , \17524 ,
         \17525 , \17526 , \17527 , \17528 , \17529 , \17530 , \17531 , \17532 , \17533 , \17534 ,
         \17535 , \17536 , \17537 , \17538 , \17539 , \17540 , \17541 , \17542 , \17543 , \17544 ,
         \17545 , \17546 , \17547 , \17548 , \17549 , \17550 , \17551 , \17552 , \17553 , \17554 ,
         \17555 , \17556 , \17557 , \17558 , \17559 , \17560 , \17561 , \17562 , \17563 , \17564 ,
         \17565 , \17566 , \17567 , \17568 , \17569 , \17570 , \17571 , \17572 , \17573 , \17574 ,
         \17575 , \17576 , \17577 , \17578 , \17579 , \17580 , \17581 , \17582 , \17583 , \17584 ,
         \17585 , \17586 , \17587 , \17588 , \17589 , \17590 , \17591 , \17592 , \17593 , \17594 ,
         \17595 , \17596 , \17597_nG5b91 , \17598 , \17599 , \17600 , \17601 , \17602 , \17603 , \17604 ,
         \17605 , \17606 , \17607 , \17608 , \17609 , \17610 , \17611 , \17612 , \17613 , \17614 ,
         \17615 , \17616 , \17617 , \17618_nG5ba6 , \17619 , \17620 , \17621 , \17622 , \17623 , \17624 ,
         \17625 , \17626 , \17627 , \17628 , \17629 , \17630 , \17631 , \17632 , \17633 , \17634 ,
         \17635 , \17636 , \17637 , \17638 , \17639 , \17640_nG5bbc , \17641 , \17642 , \17643 , \17644 ,
         \17645 , \17646 , \17647 , \17648 , \17649 , \17650 , \17651 , \17652 , \17653 , \17654 ,
         \17655 , \17656 , \17657 , \17658 , \17659 , \17660 , \17661 , \17662_nG5bd2 , \17663 , \17664 ,
         \17665 , \17666 , \17667 , \17668 , \17669 , \17670 , \17671 , \17672 , \17673 , \17674 ,
         \17675 , \17676 , \17677 , \17678 , \17679 , \17680 , \17681 , \17682 , \17683 , \17684_nG5be8 ,
         \17685 , \17686 , \17687 , \17688 , \17689 , \17690 , \17691 , \17692 , \17693 , \17694 ,
         \17695 , \17696 , \17697 , \17698 , \17699 , \17700 , \17701 , \17702 , \17703 , \17704 ,
         \17705 , \17706_nG5bfe , \17707 , \17708 , \17709 , \17710 , \17711 , \17712 , \17713 , \17714 ,
         \17715 , \17716 , \17717 , \17718 , \17719 , \17720 , \17721 , \17722 , \17723 , \17724 ,
         \17725 , \17726 , \17727 , \17728_nG5c14 , \17729 , \17730 , \17731 , \17732 , \17733 , \17734 ,
         \17735 , \17736 , \17737 , \17738 , \17739 , \17740 , \17741 , \17742 , \17743 , \17744 ,
         \17745 , \17746 , \17747 , \17748 , \17749 , \17750_nG5c2a , \17751 , \17752 , \17753 , \17754 ,
         \17755 , \17756 , \17757_nG5c31 , \17758 , \17759 , \17760 , \17761 , \17762 , \17763 , \17764 ,
         \17765 , \17766 , \17767 , \17768_nG5c3c , \17769 , \17770 , \17771 , \17772 , \17773 , \17774 ,
         \17775 , \17776 , \17777 , \17778 , \17779 , \17780 , \17781 , \17782 , \17783 , \17784 ,
         \17785 , \17786 , \17787 , \17788 , \17789 , \17790 , \17791 , \17792 , \17793 , \17794 ,
         \17795 , \17796 , \17797 , \17798 , \17799 , \17800 , \17801 , \17802 , \17803 , \17804 ,
         \17805 , \17806 , \17807 , \17808 , \17809 , \17810 , \17811 , \17812 , \17813 , \17814 ,
         \17815 , \17816 , \17817 , \17818_nG5c6f , \17819 , \17820 , \17821 , \17822 , \17823 , \17824 ,
         \17825 , \17826 , \17827 , \17828 , \17829_nG5c7a , \17830 , \17831 , \17832 , \17833 , \17834 ,
         \17835 , \17836 , \17837 , \17838 , \17839 , \17840 , \17841_nG5c86 , \17842 , \17843 , \17844 ,
         \17845 , \17846 , \17847 , \17848 , \17849 , \17850 , \17851 , \17852 , \17853 , \17854_nG5c93 ,
         \17855 , \17856 , \17857 , \17858 , \17859 , \17860 , \17861 , \17862 , \17863 , \17864 ,
         \17865 , \17866 , \17867_nG5ca0 , \17868 , \17869 , \17870 , \17871 , \17872 , \17873 , \17874 ,
         \17875 , \17876 , \17877 , \17878 , \17879 , \17880_nG5cad , \17881 , \17882 , \17883 , \17884 ,
         \17885 , \17886 , \17887 , \17888 , \17889 , \17890 , \17891 , \17892 , \17893_nG5cba , \17894 ,
         \17895 , \17896 , \17897 , \17898 , \17899 , \17900 , \17901 , \17902 , \17903 , \17904 ,
         \17905 , \17906_nG5cc7 , \17907 , \17908 , \17909 , \17910 , \17911 , \17912 , \17913 , \17914 ,
         \17915 , \17916 , \17917 , \17918 , \17919_nG5cd4 , \17920 , \17921 , \17922 , \17923 , \17924 ,
         \17925 , \17926 , \17927 , \17928 , \17929 , \17930 , \17931 , \17932 , \17933 , \17934_nG5ce3 ,
         \17935 , \17936 , \17937 , \17938 , \17939 , \17940 , \17941 , \17942 , \17943 , \17944 ,
         \17945 , \17946_nG5cef , \17947 , \17948 , \17949 , \17950 , \17951 , \17952 , \17953 , \17954 ,
         \17955 , \17956 , \17957 , \17958 , \17959_nG5cfc , \17960 , \17961 , \17962 , \17963 , \17964 ,
         \17965 , \17966 , \17967 , \17968 , \17969 , \17970 , \17971 , \17972_nG5d09 , \17973 , \17974 ,
         \17975 , \17976 , \17977 , \17978 , \17979 , \17980 , \17981 , \17982 , \17983 , \17984 ,
         \17985_nG5d16 , \17986 , \17987 , \17988 , \17989 , \17990 , \17991 , \17992 , \17993 , \17994 ,
         \17995 , \17996 , \17997 , \17998_nG5d23 , \17999 , \18000 , \18001 , \18002 , \18003 , \18004 ,
         \18005 , \18006 , \18007 , \18008 , \18009 , \18010 , \18011_nG5d30 , \18012 , \18013 , \18014 ,
         \18015 , \18016 , \18017 , \18018 , \18019 , \18020 , \18021 , \18022 , \18023 , \18024_nG5d3d ,
         \18025 , \18026 , \18027 , \18028 , \18029 , \18030 , \18031 , \18032_nG5d45 , \18033 , \18034 ,
         \18035 , \18036 , \18037 , \18038 , \18039 , \18040 , \18041 , \18042 , \18043 , \18044 ,
         \18045 , \18046 , \18047 , \18048 , \18049 , \18050 , \18051 , \18052 , \18053 , \18054 ,
         \18055 , \18056 , \18057 , \18058 , \18059 , \18060 , \18061 , \18062 , \18063 , \18064 ,
         \18065 , \18066 , \18067 , \18068 , \18069 , \18070 , \18071 , \18072 , \18073 , \18074 ,
         \18075 , \18076 , \18077 , \18078 , \18079 , \18080 , \18081 , \18082 , \18083 , \18084 ,
         \18085 , \18086 , \18087 , \18088 , \18089 , \18090 , \18091 , \18092 , \18093 , \18094 ,
         \18095 , \18096 , \18097 , \18098 , \18099 , \18100 , \18101 , \18102 , \18103 , \18104 ,
         \18105 , \18106 , \18107 , \18108 , \18109 , \18110 , \18111 , \18112 , \18113 , \18114 ,
         \18115 , \18116 , \18117 , \18118 , \18119 , \18120 , \18121 , \18122 , \18123 , \18124 ,
         \18125 , \18126 , \18127 , \18128 , \18129 , \18130 , \18131 , \18132 , \18133 , \18134 ,
         \18135 , \18136 , \18137 , \18138 , \18139 , \18140 , \18141 , \18142 , \18143 , \18144 ,
         \18145 , \18146 , \18147 , \18148 , \18149 , \18150 , \18151 , \18152 , \18153 , \18154 ,
         \18155 , \18156 , \18157 , \18158 , \18159 , \18160 , \18161 , \18162 , \18163 , \18164 ,
         \18165 , \18166 , \18167 , \18168 , \18169 , \18170 , \18171 , \18172 , \18173 , \18174 ,
         \18175 , \18176 , \18177 , \18178 , \18179 , \18180 , \18181 , \18182 , \18183 , \18184 ,
         \18185 , \18186 , \18187 , \18188 , \18189 , \18190 , \18191 , \18192 , \18193 , \18194 ,
         \18195 , \18196 , \18197 , \18198 , \18199 , \18200 , \18201 , \18202 , \18203 , \18204 ,
         \18205 , \18206 , \18207 , \18208 , \18209 , \18210 , \18211 , \18212 , \18213 , \18214 ,
         \18215 , \18216 , \18217 , \18218 , \18219 , \18220 , \18221 , \18222 , \18223 , \18224 ,
         \18225 , \18226 , \18227 , \18228 , \18229 , \18230 , \18231 , \18232 , \18233 , \18234 ,
         \18235 , \18236 , \18237 , \18238 , \18239 , \18240 , \18241 , \18242 , \18243 , \18244 ,
         \18245 , \18246 , \18247 , \18248 , \18249 , \18250 , \18251 , \18252 , \18253 , \18254 ,
         \18255 , \18256 , \18257 , \18258 , \18259 , \18260 , \18261 , \18262 , \18263 , \18264 ,
         \18265 , \18266 , \18267 , \18268 , \18269 , \18270 , \18271 , \18272 , \18273 , \18274 ,
         \18275 , \18276 , \18277 , \18278 , \18279 , \18280 , \18281 , \18282 , \18283 , \18284 ,
         \18285 , \18286 , \18287 , \18288 , \18289 , \18290 , \18291 , \18292 , \18293 , \18294 ,
         \18295 , \18296 , \18297 , \18298 , \18299 , \18300 , \18301 , \18302 , \18303 , \18304 ,
         \18305 , \18306 , \18307 , \18308 , \18309 , \18310 , \18311 , \18312 , \18313 , \18314 ,
         \18315 , \18316 , \18317 , \18318 , \18319 , \18320 , \18321 , \18322 , \18323 , \18324 ,
         \18325 , \18326 , \18327 , \18328 , \18329 , \18330 , \18331 , \18332 , \18333 , \18334 ,
         \18335 , \18336 , \18337 , \18338 , \18339 , \18340 , \18341 , \18342 , \18343 , \18344 ,
         \18345 , \18346 , \18347 , \18348 , \18349 , \18350 , \18351 , \18352 , \18353 , \18354 ,
         \18355 , \18356 , \18357 , \18358 , \18359 , \18360 , \18361 , \18362 , \18363 , \18364 ,
         \18365 , \18366 , \18367 , \18368 , \18369 , \18370 , \18371 , \18372 , \18373 , \18374 ,
         \18375 , \18376 , \18377 , \18378 , \18379 , \18380 , \18381 , \18382 , \18383 , \18384 ,
         \18385 , \18386 , \18387 , \18388 , \18389 , \18390 , \18391 , \18392 , \18393 , \18394 ,
         \18395 , \18396 , \18397 , \18398 , \18399 , \18400 , \18401 , \18402 , \18403 , \18404 ,
         \18405 , \18406 , \18407 , \18408 , \18409 , \18410 , \18411 , \18412 , \18413 , \18414 ,
         \18415 , \18416 , \18417 , \18418 , \18419 , \18420 , \18421 , \18422 , \18423 , \18424 ,
         \18425 , \18426 , \18427 , \18428 , \18429 , \18430 , \18431 , \18432 , \18433 , \18434 ,
         \18435 , \18436 , \18437 , \18438 , \18439 , \18440 , \18441 , \18442 , \18443 , \18444 ,
         \18445 , \18446 , \18447 , \18448 , \18449 , \18450 , \18451 , \18452 , \18453 , \18454 ,
         \18455 , \18456 , \18457 , \18458 , \18459 , \18460 , \18461 , \18462 , \18463 , \18464 ,
         \18465 , \18466 , \18467 , \18468 , \18469 , \18470 , \18471 , \18472 , \18473 , \18474 ,
         \18475 , \18476 , \18477 , \18478 , \18479 , \18480 , \18481 , \18482 , \18483 , \18484 ,
         \18485 , \18486 , \18487 , \18488 , \18489 , \18490 , \18491 , \18492 , \18493 , \18494 ,
         \18495 , \18496 , \18497 , \18498 , \18499 , \18500 , \18501 , \18502 , \18503 , \18504 ,
         \18505 , \18506 , \18507 , \18508 , \18509 , \18510 , \18511 , \18512 , \18513 , \18514 ,
         \18515 , \18516 , \18517 , \18518 , \18519 , \18520 , \18521 , \18522 , \18523 , \18524 ,
         \18525 , \18526 , \18527 , \18528 , \18529 , \18530 , \18531 , \18532 , \18533 , \18534 ,
         \18535 , \18536 , \18537 , \18538 , \18539 , \18540 , \18541 , \18542 , \18543 , \18544 ,
         \18545 , \18546 , \18547 , \18548 , \18549 , \18550 , \18551 , \18552 , \18553 , \18554 ,
         \18555 , \18556 , \18557 , \18558 , \18559_nG5f5c , \18560 , \18561 , \18562 , \18563 , \18564 ,
         \18565 , \18566 , \18567 , \18568 , \18569 , \18570 , \18571 , \18572 , \18573 , \18574 ,
         \18575 , \18576 , \18577 , \18578 , \18579 , \18580 , \18581 , \18582 , \18583 , \18584 ,
         \18585 , \18586 , \18587 , \18588 , \18589 , \18590 , \18591 , \18592 , \18593 , \18594 ,
         \18595 , \18596 , \18597 , \18598 , \18599 , \18600 , \18601 , \18602 , \18603 , \18604 ,
         \18605 , \18606 , \18607 , \18608 , \18609 , \18610 , \18611 , \18612 , \18613 , \18614 ,
         \18615 , \18616 , \18617 , \18618 , \18619 , \18620 , \18621 , \18622 , \18623 , \18624 ,
         \18625 , \18626 , \18627 , \18628 , \18629 , \18630 , \18631 , \18632 , \18633 , \18634 ,
         \18635 , \18636 , \18637 , \18638 , \18639 , \18640 , \18641 , \18642 , \18643 , \18644 ,
         \18645 , \18646 , \18647 , \18648 , \18649 , \18650 , \18651 , \18652 , \18653 , \18654 ,
         \18655 , \18656 , \18657 , \18658 , \18659 , \18660 , \18661 , \18662 , \18663 , \18664 ,
         \18665 , \18666 , \18667 , \18668 , \18669 , \18670 , \18671 , \18672 , \18673 , \18674 ,
         \18675 , \18676 , \18677 , \18678 , \18679 , \18680 , \18681 , \18682 , \18683 , \18684 ,
         \18685 , \18686 , \18687 , \18688 , \18689 , \18690 , \18691 , \18692 , \18693 , \18694 ,
         \18695 , \18696 , \18697 , \18698 , \18699 , \18700 , \18701 , \18702 , \18703 , \18704 ,
         \18705 , \18706 , \18707 , \18708 , \18709 , \18710 , \18711 , \18712 , \18713 , \18714 ,
         \18715 , \18716 , \18717 , \18718 , \18719 , \18720 , \18721 , \18722 , \18723 , \18724 ,
         \18725 , \18726 , \18727 , \18728 , \18729 , \18730 , \18731 , \18732 , \18733 , \18734 ,
         \18735 , \18736 , \18737 , \18738 , \18739 , \18740 , \18741 , \18742 , \18743 , \18744 ,
         \18745 , \18746 , \18747 , \18748 , \18749 , \18750 , \18751 , \18752 , \18753 , \18754 ,
         \18755 , \18756 , \18757 , \18758 , \18759 , \18760 , \18761 , \18762 , \18763 , \18764 ,
         \18765 , \18766 , \18767 , \18768 , \18769 , \18770 , \18771 , \18772 , \18773 , \18774 ,
         \18775 , \18776 , \18777 , \18778 , \18779 , \18780 , \18781 , \18782 , \18783 , \18784 ,
         \18785 , \18786 , \18787 , \18788 , \18789 , \18790 , \18791 , \18792 , \18793 , \18794 ,
         \18795 , \18796 , \18797 , \18798 , \18799 , \18800 , \18801 , \18802 , \18803 , \18804 ,
         \18805 , \18806 , \18807 , \18808 , \18809 , \18810 , \18811 , \18812 , \18813 , \18814 ,
         \18815 , \18816 , \18817 , \18818 , \18819 , \18820 , \18821 , \18822 , \18823 , \18824 ,
         \18825 , \18826 , \18827 , \18828 , \18829 , \18830 , \18831 , \18832 , \18833 , \18834 ,
         \18835 , \18836 , \18837 , \18838 , \18839 , \18840 , \18841 , \18842 , \18843 , \18844 ,
         \18845 , \18846 , \18847 , \18848 , \18849 , \18850 , \18851 , \18852 , \18853 , \18854 ,
         \18855 , \18856 , \18857 , \18858 , \18859 , \18860 , \18861 , \18862 , \18863 , \18864 ,
         \18865 , \18866 , \18867 , \18868 , \18869 , \18870 , \18871 , \18872 , \18873 , \18874 ,
         \18875 , \18876 , \18877 , \18878 , \18879 , \18880 , \18881 , \18882 , \18883 , \18884 ,
         \18885 , \18886 , \18887 , \18888 , \18889 , \18890 , \18891 , \18892 , \18893 , \18894 ,
         \18895 , \18896 , \18897 , \18898 , \18899 , \18900 , \18901 , \18902 , \18903 , \18904 ,
         \18905 , \18906 , \18907 , \18908 , \18909 , \18910 , \18911 , \18912 , \18913 , \18914 ,
         \18915 , \18916 , \18917 , \18918 , \18919 , \18920 , \18921 , \18922 , \18923 , \18924 ,
         \18925 , \18926 , \18927 , \18928 , \18929 , \18930 , \18931 , \18932 , \18933 , \18934 ,
         \18935 , \18936 , \18937 , \18938 , \18939 , \18940 , \18941 , \18942 , \18943 , \18944 ,
         \18945 , \18946 , \18947 , \18948 , \18949 , \18950 , \18951 , \18952 , \18953 , \18954 ,
         \18955 , \18956 , \18957 , \18958 , \18959 , \18960 , \18961 , \18962 , \18963 , \18964 ,
         \18965 , \18966 , \18967 , \18968 , \18969 , \18970 , \18971 , \18972 , \18973 , \18974 ,
         \18975 , \18976 , \18977 , \18978 , \18979 , \18980 , \18981 , \18982 , \18983 , \18984 ,
         \18985 , \18986 , \18987 , \18988 , \18989 , \18990 , \18991 , \18992 , \18993 , \18994 ,
         \18995 , \18996 , \18997 , \18998 , \18999 , \19000 , \19001 , \19002 , \19003 , \19004 ,
         \19005 , \19006 , \19007 , \19008 , \19009 , \19010 , \19011 , \19012 , \19013 , \19014 ,
         \19015 , \19016 , \19017 , \19018 , \19019 , \19020 , \19021 , \19022 , \19023 , \19024 ,
         \19025 , \19026 , \19027 , \19028 , \19029 , \19030 , \19031 , \19032 , \19033 , \19034 ,
         \19035 , \19036 , \19037 , \19038 , \19039 , \19040 , \19041 , \19042 , \19043 , \19044 ,
         \19045 , \19046 , \19047 , \19048 , \19049 , \19050 , \19051 , \19052 , \19053 , \19054 ,
         \19055 , \19056 , \19057 , \19058 , \19059 , \19060 , \19061 , \19062 , \19063 , \19064 ,
         \19065 , \19066 , \19067 , \19068 , \19069 , \19070_nG615b , \19071 , \19072 , \19073 , \19074 ,
         \19075 , \19076 , \19077 , \19078 , \19079 , \19080 , \19081 , \19082 , \19083 , \19084 ,
         \19085 , \19086 , \19087 , \19088 , \19089 , \19090 , \19091_nG6170 , \19092 , \19093 , \19094 ,
         \19095 , \19096 , \19097 , \19098 , \19099 , \19100 , \19101 , \19102 , \19103 , \19104 ,
         \19105 , \19106 , \19107 , \19108 , \19109 , \19110 , \19111 , \19112 , \19113_nG6186 , \19114 ,
         \19115 , \19116 , \19117 , \19118 , \19119 , \19120 , \19121 , \19122 , \19123 , \19124 ,
         \19125 , \19126 , \19127 , \19128 , \19129 , \19130 , \19131 , \19132 , \19133 , \19134 ,
         \19135_nG619c , \19136 , \19137 , \19138 , \19139 , \19140 , \19141 , \19142 , \19143 , \19144 ,
         \19145 , \19146 , \19147 , \19148 , \19149 , \19150 , \19151 , \19152 , \19153 , \19154 ,
         \19155 , \19156 , \19157_nG61b2 , \19158 , \19159 , \19160 , \19161 , \19162 , \19163 , \19164 ,
         \19165 , \19166 , \19167 , \19168 , \19169 , \19170 , \19171 , \19172 , \19173 , \19174 ,
         \19175 , \19176 , \19177 , \19178 , \19179_nG61c8 , \19180 , \19181 , \19182 , \19183 , \19184 ,
         \19185 , \19186 , \19187 , \19188 , \19189 , \19190 , \19191 , \19192 , \19193 , \19194 ,
         \19195 , \19196 , \19197 , \19198 , \19199 , \19200 , \19201_nG61de , \19202 , \19203 , \19204 ,
         \19205 , \19206 , \19207 , \19208 , \19209 , \19210 , \19211 , \19212 , \19213 , \19214 ,
         \19215 , \19216 , \19217 , \19218 , \19219 , \19220 , \19221 , \19222 , \19223_nG61f4 , \19224 ,
         \19225 , \19226 , \19227 , \19228 , \19229 , \19230 , \19231 , \19232 , \19233 , \19234 ,
         \19235 , \19236 , \19237 , \19238 , \19239 , \19240 , \19241 , \19242 , \19243 , \19244 ,
         \19245 , \19246 , \19247 , \19248 , \19249 , \19250 , \19251 , \19252 , \19253 , \19254 ,
         \19255 , \19256 , \19257 , \19258 , \19259 , \19260 , \19261 , \19262 , \19263 , \19264 ,
         \19265 , \19266 , \19267 , \19268 , \19269 , \19270 , \19271 , \19272 , \19273 , \19274 ,
         \19275 , \19276 , \19277 , \19278 , \19279 , \19280 , \19281 , \19282 , \19283 , \19284 ,
         \19285 , \19286 , \19287 , \19288 , \19289 , \19290 , \19291 , \19292 , \19293 , \19294 ,
         \19295 , \19296 , \19297 , \19298 , \19299 , \19300 , \19301 , \19302 , \19303 , \19304 ,
         \19305 , \19306 , \19307 , \19308 , \19309 , \19310 , \19311 , \19312 , \19313 , \19314 ,
         \19315 , \19316 , \19317 , \19318 , \19319 , \19320 , \19321 , \19322 , \19323 , \19324 ,
         \19325 , \19326 , \19327 , \19328 , \19329 , \19330 , \19331 , \19332 , \19333 , \19334 ,
         \19335 , \19336 , \19337 , \19338 , \19339 , \19340 , \19341 , \19342 , \19343 , \19344 ,
         \19345 , \19346 , \19347 , \19348 , \19349 , \19350 , \19351 , \19352 , \19353 , \19354 ,
         \19355 , \19356 , \19357 , \19358 , \19359 , \19360 , \19361 , \19362 , \19363 , \19364 ,
         \19365 , \19366 , \19367 , \19368 , \19369 , \19370 , \19371 , \19372 , \19373 , \19374 ,
         \19375 , \19376 , \19377 , \19378 , \19379 , \19380 , \19381 , \19382 , \19383 , \19384 ,
         \19385 , \19386 , \19387 , \19388 , \19389 , \19390 , \19391 , \19392 , \19393 , \19394 ,
         \19395 , \19396 , \19397 , \19398 , \19399 , \19400 , \19401 , \19402 , \19403 , \19404 ,
         \19405 , \19406 , \19407 , \19408 , \19409 , \19410 , \19411 , \19412 , \19413 , \19414 ,
         \19415 , \19416 , \19417 , \19418 , \19419 , \19420 , \19421 , \19422 , \19423 , \19424 ,
         \19425 , \19426 , \19427 , \19428 , \19429 , \19430 , \19431 , \19432 , \19433 , \19434 ,
         \19435 , \19436 , \19437 , \19438 , \19439 , \19440 , \19441 , \19442 , \19443 , \19444 ,
         \19445 , \19446 , \19447 , \19448 , \19449 , \19450 , \19451 , \19452 , \19453 , \19454 ,
         \19455 , \19456 , \19457 , \19458 , \19459 , \19460 , \19461 , \19462 , \19463 , \19464 ,
         \19465 , \19466 , \19467 , \19468 , \19469 , \19470 , \19471 , \19472 , \19473 , \19474 ,
         \19475 , \19476 , \19477 , \19478 , \19479 , \19480 , \19481 , \19482 , \19483 , \19484 ,
         \19485 , \19486 , \19487 , \19488 , \19489 , \19490 , \19491 , \19492 , \19493 , \19494 ,
         \19495 , \19496 , \19497 , \19498 , \19499 , \19500 , \19501 , \19502 , \19503 , \19504 ,
         \19505 , \19506 , \19507 , \19508 , \19509 , \19510 , \19511 , \19512 , \19513 , \19514 ,
         \19515 , \19516 , \19517 , \19518 , \19519 , \19520 , \19521 , \19522 , \19523 , \19524 ,
         \19525 , \19526 , \19527 , \19528 , \19529 , \19530 , \19531 , \19532 , \19533 , \19534 ,
         \19535 , \19536 , \19537 , \19538 , \19539 , \19540 , \19541 , \19542 , \19543 , \19544 ,
         \19545 , \19546 , \19547 , \19548 , \19549 , \19550 , \19551 , \19552 , \19553 , \19554 ,
         \19555 , \19556 , \19557 , \19558 , \19559 , \19560 , \19561 , \19562 , \19563 , \19564 ,
         \19565 , \19566 , \19567 , \19568 , \19569 , \19570 , \19571 , \19572 , \19573 , \19574 ,
         \19575 , \19576 , \19577 , \19578 , \19579 , \19580 , \19581 , \19582 , \19583 , \19584 ,
         \19585 , \19586 , \19587 , \19588 , \19589 , \19590 , \19591 , \19592 , \19593 , \19594 ,
         \19595 , \19596 , \19597 , \19598 , \19599 , \19600 , \19601 , \19602 , \19603 , \19604 ,
         \19605 , \19606 , \19607 , \19608 , \19609 , \19610 , \19611 , \19612 , \19613 , \19614 ,
         \19615 , \19616 , \19617 , \19618 , \19619 , \19620 , \19621 , \19622 , \19623 , \19624 ,
         \19625 , \19626 , \19627 , \19628 , \19629 , \19630 , \19631 , \19632 , \19633 , \19634 ,
         \19635 , \19636 , \19637 , \19638 , \19639 , \19640 , \19641 , \19642 , \19643 , \19644 ,
         \19645 , \19646 , \19647 , \19648 , \19649 , \19650 , \19651 , \19652 , \19653 , \19654 ,
         \19655 , \19656 , \19657 , \19658 , \19659 , \19660 , \19661 , \19662 , \19663 , \19664 ,
         \19665 , \19666 , \19667 , \19668 , \19669 , \19670 , \19671 , \19672 , \19673 , \19674 ,
         \19675 , \19676 , \19677 , \19678 , \19679 , \19680 , \19681 , \19682 , \19683 , \19684 ,
         \19685 , \19686 , \19687 , \19688 , \19689 , \19690 , \19691 , \19692 , \19693 , \19694 ,
         \19695 , \19696 , \19697 , \19698 , \19699 , \19700 , \19701 , \19702 , \19703 , \19704 ,
         \19705 , \19706 , \19707 , \19708 , \19709 , \19710 , \19711 , \19712 , \19713 , \19714 ,
         \19715 , \19716 , \19717 , \19718 , \19719 , \19720 , \19721 , \19722 , \19723 , \19724 ,
         \19725 , \19726 , \19727 , \19728 , \19729 , \19730 , \19731 , \19732 , \19733 , \19734 ,
         \19735 , \19736 , \19737 , \19738 , \19739_nG63f8 , \19740 , \19741 , \19742 , \19743 , \19744 ,
         \19745 , \19746 , \19747 , \19748 , \19749 , \19750 , \19751 , \19752 , \19753 , \19754 ,
         \19755 , \19756 , \19757 , \19758 , \19759 , \19760_nG640d , \19761 , \19762 , \19763 , \19764 ,
         \19765 , \19766 , \19767 , \19768 , \19769 , \19770 , \19771 , \19772 , \19773 , \19774 ,
         \19775 , \19776 , \19777 , \19778 , \19779 , \19780 , \19781 , \19782_nG6423 , \19783 , \19784 ,
         \19785 , \19786 , \19787 , \19788 , \19789 , \19790 , \19791 , \19792 , \19793 , \19794 ,
         \19795 , \19796 , \19797 , \19798 , \19799 , \19800 , \19801 , \19802 , \19803 , \19804_nG6439 ,
         \19805 , \19806 , \19807 , \19808 , \19809 , \19810 , \19811 , \19812 , \19813 , \19814 ,
         \19815 , \19816 , \19817 , \19818 , \19819 , \19820 , \19821 , \19822 , \19823 , \19824 ,
         \19825 , \19826_nG644f , \19827 , \19828 , \19829 , \19830 , \19831 , \19832 , \19833 , \19834 ,
         \19835 , \19836 , \19837 , \19838 , \19839 , \19840 , \19841 , \19842 , \19843 , \19844 ,
         \19845 , \19846 , \19847 , \19848_nG6465 , \19849 , \19850 , \19851 , \19852 , \19853 , \19854 ,
         \19855 , \19856 , \19857 , \19858 , \19859 , \19860 , \19861 , \19862 , \19863 , \19864 ,
         \19865 , \19866 , \19867 , \19868 , \19869 , \19870_nG647b , \19871 , \19872 , \19873 , \19874 ,
         \19875 , \19876 , \19877 , \19878 , \19879 , \19880 , \19881 , \19882 , \19883 , \19884 ,
         \19885 , \19886 , \19887 , \19888 , \19889 , \19890 , \19891 , \19892_nG6491 , \19893 , \19894 ,
         \19895 , \19896 , \19897 , \19898 , \19899_nG6498 , \19900 , \19901 , \19902 , \19903 , \19904 ,
         \19905 , \19906 , \19907 , \19908 , \19909 , \19910_nG64a3 , \19911 , \19912 , \19913 , \19914 ,
         \19915 , \19916 , \19917 , \19918 , \19919 , \19920 , \19921 , \19922 , \19923 , \19924 ,
         \19925 , \19926 , \19927 , \19928 , \19929 , \19930 , \19931 , \19932 , \19933 , \19934 ,
         \19935 , \19936 , \19937 , \19938 , \19939 , \19940 , \19941 , \19942 , \19943 , \19944 ,
         \19945 , \19946 , \19947 , \19948 , \19949 , \19950 , \19951 , \19952 , \19953 , \19954 ,
         \19955 , \19956 , \19957 , \19958 , \19959 , \19960 , \19961 , \19962 , \19963 , \19964_nG64d9 ,
         \19965 , \19966 , \19967 , \19968 , \19969 , \19970 , \19971 , \19972 , \19973 , \19974 ,
         \19975 , \19976_nG64e5 , \19977 , \19978 , \19979 , \19980 , \19981 , \19982 , \19983 , \19984 ,
         \19985 , \19986 , \19987 , \19988 , \19989_nG64f2 , \19990 , \19991 , \19992 , \19993 , \19994 ,
         \19995 , \19996 , \19997 , \19998 , \19999 , \20000 , \20001 , \20002 , \20003_nG6500 , \20004 ,
         \20005 , \20006 , \20007 , \20008 , \20009 , \20010 , \20011 , \20012 , \20013 , \20014 ,
         \20015 , \20016 , \20017_nG650e , \20018 , \20019 , \20020 , \20021 , \20022 , \20023 , \20024 ,
         \20025 , \20026 , \20027 , \20028 , \20029 , \20030 , \20031_nG651c , \20032 , \20033 , \20034 ,
         \20035 , \20036 , \20037 , \20038 , \20039 , \20040 , \20041 , \20042 , \20043 , \20044 ,
         \20045_nG652a , \20046 , \20047 , \20048 , \20049 , \20050 , \20051 , \20052 , \20053 , \20054 ,
         \20055 , \20056 , \20057 , \20058 , \20059_nG6538 , \20060 , \20061 , \20062 , \20063 , \20064 ,
         \20065 , \20066 , \20067 , \20068 , \20069 , \20070 , \20071 , \20072 , \20073_nG6546 , \20074 ,
         \20075 , \20076 , \20077 , \20078 , \20079 , \20080 , \20081 , \20082 , \20083 , \20084 ,
         \20085 , \20086 , \20087 , \20088 , \20089_nG6556 , \20090 , \20091 , \20092 , \20093 , \20094 ,
         \20095 , \20096 , \20097 , \20098 , \20099 , \20100 , \20101 , \20102_nG6563 , \20103 , \20104 ,
         \20105 , \20106 , \20107 , \20108 , \20109 , \20110 , \20111 , \20112 , \20113 , \20114 ,
         \20115 , \20116_nG6571 , \20117 , \20118 , \20119 , \20120 , \20121 , \20122 , \20123 , \20124 ,
         \20125 , \20126 , \20127 , \20128 , \20129 , \20130_nG657f , \20131 , \20132 , \20133 , \20134 ,
         \20135 , \20136 , \20137 , \20138 , \20139 , \20140 , \20141 , \20142 , \20143 , \20144_nG658d ,
         \20145 , \20146 , \20147 , \20148 , \20149 , \20150 , \20151 , \20152 , \20153 , \20154 ,
         \20155 , \20156 , \20157 , \20158_nG659b , \20159 , \20160 , \20161 , \20162 , \20163 , \20164 ,
         \20165 , \20166 , \20167 , \20168 , \20169 , \20170 , \20171 , \20172_nG65a9 , \20173 , \20174 ,
         \20175 , \20176 , \20177 , \20178 , \20179 , \20180 , \20181 , \20182 , \20183 , \20184 ,
         \20185 , \20186_nG65b7 , \20187 , \20188 , \20189 , \20190 , \20191 , \20192 , \20193 , \20194_nG65bf ,
         \20195 , \20196 , \20197 , \20198 , \20199 , \20200 , \20201 , \20202 , \20203 , \20204 ,
         \20205 , \20206 , \20207 , \20208 , \20209 , \20210 , \20211 , \20212 , \20213 , \20214 ,
         \20215 , \20216 , \20217 , \20218 , \20219 , \20220 , \20221 , \20222 , \20223 , \20224 ,
         \20225 , \20226 , \20227 , \20228 , \20229 , \20230 , \20231 , \20232 , \20233 , \20234 ,
         \20235 , \20236 , \20237 , \20238 , \20239 , \20240 , \20241 , \20242 , \20243 , \20244 ,
         \20245 , \20246 , \20247 , \20248 , \20249 , \20250 , \20251 , \20252 , \20253 , \20254 ,
         \20255 , \20256 , \20257 , \20258 , \20259 , \20260 , \20261 , \20262 , \20263 , \20264 ,
         \20265 , \20266 , \20267 , \20268 , \20269 , \20270 , \20271 , \20272 , \20273 , \20274 ,
         \20275 , \20276 , \20277 , \20278 , \20279 , \20280 , \20281 , \20282 , \20283 , \20284 ,
         \20285 , \20286 , \20287 , \20288 , \20289 , \20290 , \20291 , \20292 , \20293 , \20294 ,
         \20295 , \20296 , \20297 , \20298 , \20299 , \20300 , \20301 , \20302 , \20303 , \20304 ,
         \20305 , \20306 , \20307 , \20308 , \20309 , \20310 , \20311 , \20312 , \20313 , \20314 ,
         \20315 , \20316 , \20317 , \20318 , \20319 , \20320 , \20321 , \20322 , \20323 , \20324 ,
         \20325 , \20326 , \20327 , \20328 , \20329 , \20330 , \20331 , \20332 , \20333 , \20334 ,
         \20335 , \20336 , \20337 , \20338 , \20339 , \20340 , \20341 , \20342 , \20343 , \20344 ,
         \20345 , \20346 , \20347 , \20348 , \20349 , \20350 , \20351 , \20352 , \20353 , \20354 ,
         \20355 , \20356 , \20357 , \20358 , \20359 , \20360 , \20361 , \20362 , \20363 , \20364 ,
         \20365 , \20366 , \20367 , \20368 , \20369 , \20370 , \20371 , \20372 , \20373 , \20374 ,
         \20375 , \20376 , \20377 , \20378 , \20379 , \20380 , \20381 , \20382 , \20383 , \20384 ,
         \20385 , \20386 , \20387 , \20388 , \20389 , \20390 , \20391 , \20392 , \20393 , \20394 ,
         \20395 , \20396 , \20397 , \20398 , \20399 , \20400 , \20401 , \20402 , \20403 , \20404 ,
         \20405 , \20406 , \20407 , \20408 , \20409 , \20410 , \20411 , \20412 , \20413 , \20414 ,
         \20415 , \20416 , \20417 , \20418 , \20419 , \20420 , \20421 , \20422 , \20423 , \20424 ,
         \20425 , \20426 , \20427 , \20428 , \20429 , \20430 , \20431 , \20432 , \20433 , \20434 ,
         \20435 , \20436 , \20437 , \20438 , \20439 , \20440 , \20441 , \20442 , \20443 , \20444 ,
         \20445 , \20446 , \20447 , \20448 , \20449 , \20450 , \20451 , \20452 , \20453 , \20454 ,
         \20455 , \20456 , \20457 , \20458 , \20459 , \20460 , \20461 , \20462 , \20463 , \20464 ,
         \20465 , \20466 , \20467 , \20468 , \20469 , \20470 , \20471 , \20472 , \20473 , \20474 ,
         \20475 , \20476 , \20477 , \20478 , \20479 , \20480 , \20481 , \20482 , \20483 , \20484 ,
         \20485 , \20486 , \20487 , \20488 , \20489 , \20490 , \20491 , \20492 , \20493 , \20494 ,
         \20495 , \20496 , \20497 , \20498 , \20499 , \20500 , \20501 , \20502 , \20503 , \20504 ,
         \20505 , \20506 , \20507 , \20508 , \20509 , \20510 , \20511 , \20512 , \20513 , \20514 ,
         \20515 , \20516 , \20517 , \20518 , \20519 , \20520 , \20521 , \20522 , \20523 , \20524 ,
         \20525 , \20526 , \20527 , \20528 , \20529 , \20530 , \20531 , \20532 , \20533 , \20534 ,
         \20535 , \20536 , \20537 , \20538 , \20539 , \20540 , \20541 , \20542 , \20543 , \20544 ,
         \20545 , \20546 , \20547 , \20548 , \20549 , \20550 , \20551 , \20552 , \20553 , \20554 ,
         \20555 , \20556 , \20557 , \20558 , \20559 , \20560 , \20561 , \20562 , \20563 , \20564 ,
         \20565 , \20566 , \20567 , \20568 , \20569 , \20570 , \20571 , \20572 , \20573 , \20574 ,
         \20575 , \20576 , \20577 , \20578 , \20579 , \20580 , \20581 , \20582 , \20583 , \20584 ,
         \20585 , \20586 , \20587 , \20588 , \20589 , \20590 , \20591 , \20592 , \20593 , \20594 ,
         \20595 , \20596 , \20597 , \20598 , \20599 , \20600 , \20601 , \20602 , \20603 , \20604 ,
         \20605 , \20606 , \20607 , \20608 , \20609 , \20610 , \20611 , \20612 , \20613 , \20614 ,
         \20615 , \20616 , \20617 , \20618 , \20619 , \20620 , \20621 , \20622 , \20623 , \20624 ,
         \20625 , \20626 , \20627 , \20628 , \20629 , \20630 , \20631 , \20632 , \20633 , \20634 ,
         \20635 , \20636 , \20637 , \20638 , \20639 , \20640 , \20641 , \20642 , \20643 , \20644 ,
         \20645 , \20646 , \20647 , \20648 , \20649 , \20650 , \20651 , \20652 , \20653 , \20654 ,
         \20655 , \20656 , \20657 , \20658 , \20659 , \20660 , \20661 , \20662 , \20663 , \20664 ,
         \20665 , \20666 , \20667 , \20668 , \20669 , \20670 , \20671 , \20672 , \20673 , \20674 ,
         \20675 , \20676 , \20677 , \20678 , \20679 , \20680 , \20681 , \20682 , \20683 , \20684 ,
         \20685 , \20686 , \20687 , \20688 , \20689 , \20690 , \20691 , \20692 , \20693 , \20694 ,
         \20695 , \20696 , \20697 , \20698 , \20699 , \20700 , \20701 , \20702 , \20703 , \20704 ,
         \20705 , \20706 , \20707 , \20708 , \20709 , \20710 , \20711 , \20712 , \20713 , \20714 ,
         \20715 , \20716 , \20717 , \20718 , \20719 , \20720 , \20721_nG67d6 , \20722 , \20723 , \20724 ,
         \20725 , \20726 , \20727 , \20728 , \20729 , \20730 , \20731 , \20732 , \20733 , \20734 ,
         \20735 , \20736 , \20737 , \20738 , \20739 , \20740 , \20741 , \20742 , \20743 , \20744 ,
         \20745 , \20746 , \20747 , \20748 , \20749 , \20750 , \20751 , \20752 , \20753 , \20754 ,
         \20755 , \20756 , \20757 , \20758 , \20759 , \20760 , \20761 , \20762 , \20763 , \20764 ,
         \20765 , \20766 , \20767 , \20768 , \20769 , \20770 , \20771 , \20772 , \20773 , \20774 ,
         \20775 , \20776 , \20777 , \20778 , \20779 , \20780 , \20781 , \20782 , \20783 , \20784 ,
         \20785 , \20786 , \20787 , \20788 , \20789 , \20790 , \20791 , \20792 , \20793 , \20794 ,
         \20795 , \20796 , \20797 , \20798 , \20799 , \20800 , \20801 , \20802 , \20803 , \20804 ,
         \20805 , \20806 , \20807 , \20808 , \20809 , \20810 , \20811 , \20812 , \20813 , \20814 ,
         \20815 , \20816 , \20817 , \20818 , \20819 , \20820 , \20821 , \20822 , \20823 , \20824 ,
         \20825 , \20826 , \20827 , \20828 , \20829 , \20830 , \20831 , \20832 , \20833 , \20834 ,
         \20835 , \20836 , \20837 , \20838 , \20839 , \20840 , \20841 , \20842 , \20843 , \20844 ,
         \20845 , \20846 , \20847 , \20848 , \20849 , \20850 , \20851 , \20852 , \20853 , \20854 ,
         \20855 , \20856 , \20857 , \20858 , \20859 , \20860 , \20861 , \20862 , \20863 , \20864 ,
         \20865 , \20866 , \20867 , \20868 , \20869 , \20870 , \20871 , \20872 , \20873 , \20874 ,
         \20875 , \20876 , \20877 , \20878 , \20879 , \20880 , \20881 , \20882 , \20883 , \20884 ,
         \20885 , \20886 , \20887 , \20888 , \20889 , \20890 , \20891 , \20892 , \20893 , \20894 ,
         \20895 , \20896 , \20897 , \20898 , \20899 , \20900 , \20901 , \20902 , \20903 , \20904 ,
         \20905 , \20906 , \20907 , \20908 , \20909 , \20910 , \20911 , \20912 , \20913 , \20914 ,
         \20915 , \20916 , \20917 , \20918 , \20919 , \20920 , \20921 , \20922 , \20923 , \20924 ,
         \20925 , \20926 , \20927 , \20928 , \20929 , \20930 , \20931 , \20932 , \20933 , \20934 ,
         \20935 , \20936 , \20937 , \20938 , \20939 , \20940 , \20941 , \20942 , \20943 , \20944 ,
         \20945 , \20946 , \20947 , \20948 , \20949 , \20950 , \20951 , \20952 , \20953 , \20954 ,
         \20955 , \20956 , \20957 , \20958 , \20959 , \20960 , \20961 , \20962 , \20963 , \20964 ,
         \20965 , \20966 , \20967 , \20968 , \20969 , \20970 , \20971 , \20972 , \20973 , \20974 ,
         \20975 , \20976 , \20977 , \20978 , \20979 , \20980 , \20981 , \20982 , \20983 , \20984 ,
         \20985 , \20986 , \20987 , \20988 , \20989 , \20990 , \20991 , \20992 , \20993 , \20994 ,
         \20995 , \20996 , \20997 , \20998 , \20999 , \21000 , \21001 , \21002 , \21003 , \21004 ,
         \21005 , \21006 , \21007 , \21008 , \21009 , \21010 , \21011 , \21012 , \21013 , \21014 ,
         \21015 , \21016 , \21017 , \21018 , \21019 , \21020 , \21021 , \21022 , \21023 , \21024 ,
         \21025 , \21026 , \21027 , \21028 , \21029 , \21030 , \21031 , \21032 , \21033 , \21034 ,
         \21035 , \21036 , \21037 , \21038 , \21039 , \21040 , \21041 , \21042 , \21043 , \21044 ,
         \21045 , \21046 , \21047 , \21048 , \21049 , \21050 , \21051 , \21052 , \21053 , \21054 ,
         \21055 , \21056 , \21057 , \21058 , \21059 , \21060 , \21061 , \21062 , \21063 , \21064 ,
         \21065 , \21066 , \21067 , \21068 , \21069 , \21070 , \21071 , \21072 , \21073 , \21074 ,
         \21075 , \21076 , \21077 , \21078 , \21079 , \21080 , \21081 , \21082 , \21083 , \21084 ,
         \21085 , \21086 , \21087 , \21088 , \21089 , \21090 , \21091 , \21092 , \21093 , \21094 ,
         \21095 , \21096 , \21097 , \21098 , \21099 , \21100 , \21101 , \21102 , \21103 , \21104 ,
         \21105 , \21106 , \21107 , \21108 , \21109 , \21110 , \21111 , \21112 , \21113 , \21114 ,
         \21115 , \21116 , \21117 , \21118 , \21119 , \21120 , \21121 , \21122 , \21123 , \21124 ,
         \21125 , \21126 , \21127 , \21128 , \21129 , \21130 , \21131 , \21132 , \21133 , \21134 ,
         \21135 , \21136 , \21137 , \21138 , \21139 , \21140 , \21141 , \21142 , \21143 , \21144 ,
         \21145 , \21146 , \21147 , \21148 , \21149 , \21150 , \21151 , \21152 , \21153 , \21154 ,
         \21155 , \21156 , \21157 , \21158 , \21159 , \21160 , \21161 , \21162 , \21163 , \21164 ,
         \21165 , \21166 , \21167 , \21168 , \21169 , \21170 , \21171 , \21172 , \21173 , \21174 ,
         \21175 , \21176 , \21177 , \21178 , \21179 , \21180 , \21181 , \21182 , \21183 , \21184 ,
         \21185 , \21186 , \21187 , \21188 , \21189 , \21190 , \21191 , \21192 , \21193 , \21194 ,
         \21195 , \21196 , \21197 , \21198 , \21199 , \21200 , \21201 , \21202 , \21203 , \21204 ,
         \21205 , \21206 , \21207 , \21208 , \21209 , \21210 , \21211 , \21212 , \21213 , \21214 ,
         \21215 , \21216 , \21217 , \21218 , \21219 , \21220 , \21221 , \21222 , \21223 , \21224 ,
         \21225 , \21226 , \21227 , \21228 , \21229 , \21230 , \21231 , \21232_nG69d5 , \21233 , \21234 ,
         \21235 , \21236 , \21237 , \21238 , \21239 , \21240 , \21241 , \21242 , \21243 , \21244 ,
         \21245 , \21246 , \21247 , \21248 , \21249 , \21250 , \21251 , \21252 , \21253_nG69ea , \21254 ,
         \21255 , \21256 , \21257 , \21258 , \21259 , \21260 , \21261 , \21262 , \21263 , \21264 ,
         \21265 , \21266 , \21267 , \21268 , \21269 , \21270 , \21271 , \21272 , \21273 , \21274 ,
         \21275_nG6a00 , \21276 , \21277 , \21278 , \21279 , \21280 , \21281 , \21282 , \21283 , \21284 ,
         \21285 , \21286 , \21287 , \21288 , \21289 , \21290 , \21291 , \21292 , \21293 , \21294 ,
         \21295 , \21296 , \21297_nG6a16 , \21298 , \21299 , \21300 , \21301 , \21302 , \21303 , \21304 ,
         \21305 , \21306 , \21307 , \21308 , \21309 , \21310 , \21311 , \21312 , \21313 , \21314 ,
         \21315 , \21316 , \21317 , \21318 , \21319_nG6a2c , \21320 , \21321 , \21322 , \21323 , \21324 ,
         \21325 , \21326 , \21327 , \21328 , \21329 , \21330 , \21331 , \21332 , \21333 , \21334 ,
         \21335 , \21336 , \21337 , \21338 , \21339 , \21340 , \21341_nG6a42 , \21342 , \21343 , \21344 ,
         \21345 , \21346 , \21347 , \21348 , \21349 , \21350 , \21351 , \21352 , \21353 , \21354 ,
         \21355 , \21356 , \21357 , \21358 , \21359 , \21360 , \21361 , \21362 , \21363_nG6a58 , \21364 ,
         \21365 , \21366 , \21367 , \21368 , \21369 , \21370 , \21371 , \21372 , \21373 , \21374 ,
         \21375 , \21376 , \21377 , \21378 , \21379 , \21380 , \21381 , \21382 , \21383 , \21384 ,
         \21385_nG6a6e , \21386 , \21387 , \21388 , \21389 , \21390 , \21391 , \21392 , \21393 , \21394 ,
         \21395 , \21396 , \21397 , \21398 , \21399 , \21400 , \21401 , \21402 , \21403 , \21404 ,
         \21405 , \21406 , \21407 , \21408 , \21409 , \21410 , \21411 , \21412 , \21413 , \21414 ,
         \21415 , \21416 , \21417 , \21418 , \21419 , \21420 , \21421 , \21422 , \21423 , \21424 ,
         \21425 , \21426 , \21427 , \21428 , \21429 , \21430 , \21431 , \21432 , \21433 , \21434 ,
         \21435 , \21436 , \21437 , \21438 , \21439 , \21440 , \21441 , \21442 , \21443 , \21444 ,
         \21445 , \21446 , \21447 , \21448 , \21449 , \21450 , \21451 , \21452 , \21453 , \21454 ,
         \21455 , \21456 , \21457 , \21458 , \21459 , \21460 , \21461 , \21462 , \21463 , \21464 ,
         \21465 , \21466 , \21467 , \21468 , \21469 , \21470 , \21471 , \21472 , \21473 , \21474 ,
         \21475 , \21476 , \21477 , \21478 , \21479 , \21480 , \21481 , \21482 , \21483 , \21484 ,
         \21485 , \21486 , \21487 , \21488 , \21489 , \21490 , \21491 , \21492 , \21493 , \21494 ,
         \21495 , \21496 , \21497 , \21498 , \21499 , \21500 , \21501 , \21502 , \21503 , \21504 ,
         \21505 , \21506 , \21507 , \21508 , \21509 , \21510 , \21511 , \21512 , \21513 , \21514 ,
         \21515 , \21516 , \21517 , \21518 , \21519 , \21520 , \21521 , \21522 , \21523 , \21524 ,
         \21525 , \21526 , \21527 , \21528 , \21529 , \21530 , \21531 , \21532 , \21533 , \21534 ,
         \21535 , \21536 , \21537 , \21538 , \21539 , \21540 , \21541 , \21542 , \21543 , \21544 ,
         \21545 , \21546 , \21547 , \21548 , \21549 , \21550 , \21551 , \21552 , \21553 , \21554 ,
         \21555 , \21556 , \21557 , \21558 , \21559 , \21560 , \21561 , \21562 , \21563 , \21564 ,
         \21565 , \21566 , \21567 , \21568 , \21569 , \21570 , \21571 , \21572 , \21573 , \21574 ,
         \21575 , \21576 , \21577 , \21578 , \21579 , \21580 , \21581 , \21582 , \21583 , \21584 ,
         \21585 , \21586 , \21587 , \21588 , \21589 , \21590 , \21591 , \21592 , \21593 , \21594 ,
         \21595 , \21596 , \21597 , \21598 , \21599 , \21600 , \21601 , \21602 , \21603 , \21604 ,
         \21605 , \21606 , \21607 , \21608 , \21609 , \21610 , \21611 , \21612 , \21613 , \21614 ,
         \21615 , \21616 , \21617 , \21618 , \21619 , \21620 , \21621 , \21622 , \21623 , \21624 ,
         \21625 , \21626 , \21627 , \21628 , \21629 , \21630 , \21631 , \21632 , \21633 , \21634 ,
         \21635 , \21636 , \21637 , \21638 , \21639 , \21640 , \21641 , \21642 , \21643 , \21644 ,
         \21645 , \21646 , \21647 , \21648 , \21649 , \21650 , \21651 , \21652 , \21653 , \21654 ,
         \21655 , \21656 , \21657 , \21658 , \21659 , \21660 , \21661 , \21662 , \21663 , \21664 ,
         \21665 , \21666 , \21667 , \21668 , \21669 , \21670 , \21671 , \21672 , \21673 , \21674 ,
         \21675 , \21676 , \21677 , \21678 , \21679 , \21680 , \21681 , \21682 , \21683 , \21684 ,
         \21685 , \21686 , \21687 , \21688 , \21689 , \21690 , \21691 , \21692 , \21693 , \21694 ,
         \21695 , \21696 , \21697 , \21698 , \21699 , \21700 , \21701 , \21702 , \21703 , \21704 ,
         \21705 , \21706 , \21707 , \21708 , \21709 , \21710 , \21711 , \21712 , \21713 , \21714 ,
         \21715 , \21716 , \21717 , \21718 , \21719 , \21720 , \21721 , \21722 , \21723 , \21724 ,
         \21725 , \21726 , \21727 , \21728 , \21729 , \21730 , \21731 , \21732 , \21733 , \21734 ,
         \21735 , \21736 , \21737 , \21738 , \21739 , \21740 , \21741 , \21742 , \21743 , \21744 ,
         \21745 , \21746 , \21747 , \21748 , \21749 , \21750 , \21751 , \21752 , \21753 , \21754 ,
         \21755 , \21756 , \21757 , \21758 , \21759 , \21760 , \21761 , \21762 , \21763 , \21764 ,
         \21765 , \21766 , \21767 , \21768 , \21769 , \21770 , \21771 , \21772 , \21773 , \21774 ,
         \21775 , \21776 , \21777 , \21778 , \21779 , \21780 , \21781 , \21782 , \21783 , \21784 ,
         \21785 , \21786 , \21787 , \21788 , \21789 , \21790 , \21791 , \21792 , \21793 , \21794 ,
         \21795 , \21796 , \21797 , \21798 , \21799 , \21800 , \21801 , \21802 , \21803 , \21804 ,
         \21805 , \21806 , \21807 , \21808 , \21809 , \21810 , \21811 , \21812 , \21813 , \21814 ,
         \21815 , \21816 , \21817 , \21818 , \21819 , \21820 , \21821 , \21822 , \21823 , \21824 ,
         \21825 , \21826 , \21827 , \21828 , \21829 , \21830 , \21831 , \21832 , \21833 , \21834 ,
         \21835 , \21836 , \21837 , \21838 , \21839 , \21840 , \21841 , \21842 , \21843 , \21844 ,
         \21845 , \21846 , \21847 , \21848 , \21849 , \21850 , \21851 , \21852 , \21853 , \21854 ,
         \21855 , \21856 , \21857 , \21858 , \21859 , \21860 , \21861 , \21862 , \21863 , \21864 ,
         \21865 , \21866 , \21867 , \21868 , \21869 , \21870 , \21871 , \21872 , \21873 , \21874 ,
         \21875 , \21876 , \21877 , \21878 , \21879 , \21880 , \21881 , \21882 , \21883 , \21884 ,
         \21885 , \21886 , \21887 , \21888 , \21889 , \21890 , \21891 , \21892 , \21893 , \21894 ,
         \21895 , \21896 , \21897 , \21898 , \21899 , \21900 , \21901_nG6c72 , \21902 , \21903 , \21904 ,
         \21905 , \21906 , \21907 , \21908 , \21909 , \21910 , \21911 , \21912 , \21913 , \21914 ,
         \21915 , \21916 , \21917 , \21918 , \21919 , \21920 , \21921 , \21922_nG6c87 , \21923 , \21924 ,
         \21925 , \21926 , \21927 , \21928 , \21929 , \21930 , \21931 , \21932 , \21933 , \21934 ,
         \21935 , \21936 , \21937 , \21938 , \21939 , \21940 , \21941 , \21942 , \21943 , \21944_nG6c9d ,
         \21945 , \21946 , \21947 , \21948 , \21949 , \21950 , \21951 , \21952 , \21953 , \21954 ,
         \21955 , \21956 , \21957 , \21958 , \21959 , \21960 , \21961 , \21962 , \21963 , \21964 ,
         \21965 , \21966_nG6cb3 , \21967 , \21968 , \21969 , \21970 , \21971 , \21972 , \21973 , \21974 ,
         \21975 , \21976 , \21977 , \21978 , \21979 , \21980 , \21981 , \21982 , \21983 , \21984 ,
         \21985 , \21986 , \21987 , \21988_nG6cc9 , \21989 , \21990 , \21991 , \21992 , \21993 , \21994 ,
         \21995 , \21996 , \21997 , \21998 , \21999 , \22000 , \22001 , \22002 , \22003 , \22004 ,
         \22005 , \22006 , \22007 , \22008 , \22009 , \22010_nG6cdf , \22011 , \22012 , \22013 , \22014 ,
         \22015 , \22016 , \22017 , \22018 , \22019 , \22020 , \22021 , \22022 , \22023 , \22024 ,
         \22025 , \22026 , \22027 , \22028 , \22029 , \22030 , \22031 , \22032_nG6cf5 , \22033 , \22034 ,
         \22035 , \22036 , \22037 , \22038 , \22039 , \22040 , \22041 , \22042 , \22043 , \22044 ,
         \22045 , \22046 , \22047 , \22048 , \22049 , \22050 , \22051 , \22052 , \22053 , \22054_nG6d0b ,
         \22055 , \22056 , \22057 , \22058 , \22059 , \22060 , \22061_nG6d12 , \22062 , \22063 , \22064 ,
         \22065 , \22066 , \22067 , \22068 , \22069 , \22070 , \22071 , \22072_nG6d1d , \22073 , \22074 ,
         \22075 , \22076 , \22077 , \22078 , \22079 , \22080 , \22081 , \22082 , \22083 , \22084 ,
         \22085 , \22086 , \22087 , \22088 , \22089 , \22090 , \22091 , \22092 , \22093 , \22094 ,
         \22095 , \22096 , \22097 , \22098 , \22099 , \22100 , \22101 , \22102 , \22103 , \22104 ,
         \22105 , \22106 , \22107 , \22108 , \22109 , \22110 , \22111 , \22112 , \22113 , \22114 ,
         \22115 , \22116 , \22117 , \22118 , \22119 , \22120 , \22121 , \22122_nG6d52 , \22123 , \22124 ,
         \22125 , \22126 , \22127 , \22128 , \22129 , \22130 , \22131 , \22132 , \22133 , \22134 ,
         \22135_nG6d5f , \22136 , \22137 , \22138 , \22139 , \22140 , \22141 , \22142 , \22143 , \22144 ,
         \22145 , \22146 , \22147 , \22148 , \22149_nG6d6d , \22150 , \22151 , \22152 , \22153 , \22154 ,
         \22155 , \22156 , \22157 , \22158 , \22159 , \22160 , \22161 , \22162 , \22163 , \22164_nG6d7c ,
         \22165 , \22166 , \22167 , \22168 , \22169 , \22170 , \22171 , \22172 , \22173 , \22174 ,
         \22175 , \22176 , \22177 , \22178 , \22179_nG6d8b , \22180 , \22181 , \22182 , \22183 , \22184 ,
         \22185 , \22186 , \22187 , \22188 , \22189 , \22190 , \22191 , \22192 , \22193 , \22194_nG6d9a ,
         \22195 , \22196 , \22197 , \22198 , \22199 , \22200 , \22201 , \22202 , \22203 , \22204 ,
         \22205 , \22206 , \22207 , \22208 , \22209_nG6da9 , \22210 , \22211 , \22212 , \22213 , \22214 ,
         \22215 , \22216 , \22217 , \22218 , \22219 , \22220 , \22221 , \22222 , \22223 , \22224_nG6db8 ,
         \22225 , \22226 , \22227 , \22228 , \22229 , \22230 , \22231 , \22232 , \22233 , \22234 ,
         \22235 , \22236 , \22237 , \22238 , \22239_nG6dc7 , \22240 , \22241 , \22242 , \22243 , \22244 ,
         \22245 , \22246 , \22247 , \22248 , \22249 , \22250 , \22251 , \22252 , \22253 , \22254 ,
         \22255 , \22256_nG6dd8 , \22257 , \22258 , \22259 , \22260 , \22261 , \22262 , \22263 , \22264 ,
         \22265 , \22266 , \22267 , \22268 , \22269 , \22270_nG6de6 , \22271 , \22272 , \22273 , \22274 ,
         \22275 , \22276 , \22277 , \22278 , \22279 , \22280 , \22281 , \22282 , \22283 , \22284 ,
         \22285_nG6df5 , \22286 , \22287 , \22288 , \22289 , \22290 , \22291 , \22292 , \22293 , \22294 ,
         \22295 , \22296 , \22297 , \22298 , \22299 , \22300_nG6e04 , \22301 , \22302 , \22303 , \22304 ,
         \22305 , \22306 , \22307 , \22308 , \22309 , \22310 , \22311 , \22312 , \22313 , \22314 ,
         \22315_nG6e13 , \22316 , \22317 , \22318 , \22319 , \22320 , \22321 , \22322 , \22323 , \22324 ,
         \22325 , \22326 , \22327 , \22328 , \22329 , \22330_nG6e22 , \22331 , \22332 , \22333 , \22334 ,
         \22335 , \22336 , \22337 , \22338 , \22339 , \22340 , \22341 , \22342 , \22343 , \22344 ,
         \22345_nG6e31 , \22346 , \22347 , \22348 , \22349 , \22350 , \22351 , \22352 , \22353 , \22354 ,
         \22355 , \22356 , \22357 , \22358 , \22359 , \22360_nG6e40 , \22361 , \22362 , \22363 , \22364 ,
         \22365 , \22366 , \22367 , \22368_nG6e48 , \22369 , \22370 , \22371 , \22372 , \22373 , \22374 ,
         \22375 , \22376 , \22377 , \22378 , \22379 , \22380 , \22381 , \22382 , \22383 , \22384 ,
         \22385 , \22386 , \22387 , \22388 , \22389 , \22390 , \22391 , \22392 , \22393 , \22394 ,
         \22395 , \22396 , \22397 , \22398 , \22399 , \22400 , \22401 , \22402 , \22403 , \22404 ,
         \22405 , \22406 , \22407 , \22408 , \22409 , \22410 , \22411 , \22412 , \22413 , \22414 ,
         \22415 , \22416 , \22417 , \22418 , \22419 , \22420 , \22421 , \22422 , \22423 , \22424 ,
         \22425 , \22426 , \22427 , \22428 , \22429 , \22430 , \22431 , \22432 , \22433 , \22434 ,
         \22435 , \22436 , \22437 , \22438 , \22439 , \22440 , \22441 , \22442 , \22443 , \22444 ,
         \22445 , \22446 , \22447 , \22448 , \22449 , \22450 , \22451 , \22452 , \22453 , \22454 ,
         \22455 , \22456 , \22457 , \22458 , \22459 , \22460 , \22461 , \22462 , \22463 , \22464 ,
         \22465 , \22466 , \22467 , \22468 , \22469 , \22470 , \22471 , \22472 , \22473 , \22474 ,
         \22475 , \22476 , \22477 , \22478 , \22479 , \22480 , \22481 , \22482 , \22483 , \22484 ,
         \22485 , \22486 , \22487 , \22488 , \22489 , \22490 , \22491 , \22492 , \22493 , \22494 ,
         \22495 , \22496 , \22497 , \22498 , \22499 , \22500 , \22501 , \22502 , \22503 , \22504 ,
         \22505 , \22506 , \22507 , \22508 , \22509 , \22510 , \22511 , \22512 , \22513 , \22514 ,
         \22515 , \22516 , \22517 , \22518 , \22519 , \22520 , \22521 , \22522 , \22523 , \22524 ,
         \22525 , \22526 , \22527 , \22528 , \22529 , \22530 , \22531 , \22532 , \22533 , \22534 ,
         \22535 , \22536 , \22537 , \22538 , \22539 , \22540 , \22541 , \22542 , \22543 , \22544 ,
         \22545 , \22546 , \22547 , \22548 , \22549 , \22550 , \22551 , \22552 , \22553 , \22554 ,
         \22555 , \22556 , \22557 , \22558 , \22559 , \22560 , \22561 , \22562 , \22563 , \22564 ,
         \22565 , \22566 , \22567 , \22568 , \22569 , \22570 , \22571 , \22572 , \22573 , \22574 ,
         \22575 , \22576 , \22577 , \22578 , \22579 , \22580 , \22581 , \22582 , \22583 , \22584 ,
         \22585 , \22586 , \22587 , \22588 , \22589 , \22590 , \22591 , \22592 , \22593 , \22594 ,
         \22595 , \22596 , \22597 , \22598 , \22599 , \22600 , \22601 , \22602 , \22603 , \22604 ,
         \22605 , \22606 , \22607 , \22608 , \22609 , \22610 , \22611 , \22612 , \22613 , \22614 ,
         \22615 , \22616 , \22617 , \22618 , \22619 , \22620 , \22621 , \22622 , \22623 , \22624 ,
         \22625 , \22626 , \22627 , \22628 , \22629 , \22630 , \22631 , \22632 , \22633 , \22634 ,
         \22635 , \22636 , \22637 , \22638 , \22639 , \22640 , \22641 , \22642 , \22643 , \22644 ,
         \22645 , \22646 , \22647 , \22648 , \22649 , \22650 , \22651 , \22652 , \22653 , \22654 ,
         \22655 , \22656 , \22657 , \22658 , \22659 , \22660 , \22661 , \22662 , \22663 , \22664 ,
         \22665 , \22666 , \22667 , \22668 , \22669 , \22670 , \22671 , \22672 , \22673 , \22674 ,
         \22675 , \22676 , \22677 , \22678 , \22679 , \22680 , \22681 , \22682 , \22683 , \22684 ,
         \22685 , \22686 , \22687 , \22688 , \22689 , \22690 , \22691 , \22692 , \22693 , \22694 ,
         \22695 , \22696 , \22697 , \22698 , \22699 , \22700 , \22701 , \22702 , \22703 , \22704 ,
         \22705 , \22706 , \22707 , \22708 , \22709 , \22710 , \22711 , \22712 , \22713 , \22714 ,
         \22715 , \22716 , \22717 , \22718 , \22719 , \22720 , \22721 , \22722 , \22723 , \22724 ,
         \22725 , \22726 , \22727 , \22728 , \22729 , \22730 , \22731 , \22732 , \22733 , \22734 ,
         \22735 , \22736 , \22737 , \22738 , \22739 , \22740 , \22741 , \22742 , \22743 , \22744 ,
         \22745 , \22746 , \22747 , \22748 , \22749 , \22750 , \22751 , \22752 , \22753 , \22754 ,
         \22755 , \22756 , \22757 , \22758 , \22759 , \22760 , \22761 , \22762 , \22763 , \22764 ,
         \22765 , \22766 , \22767 , \22768 , \22769 , \22770 , \22771 , \22772 , \22773 , \22774 ,
         \22775 , \22776 , \22777 , \22778 , \22779 , \22780 , \22781 , \22782 , \22783 , \22784 ,
         \22785 , \22786 , \22787 , \22788 , \22789 , \22790 , \22791 , \22792 , \22793 , \22794 ,
         \22795 , \22796 , \22797 , \22798 , \22799 , \22800 , \22801 , \22802 , \22803 , \22804 ,
         \22805 , \22806 , \22807 , \22808 , \22809 , \22810 , \22811 , \22812 , \22813 , \22814 ,
         \22815 , \22816 , \22817 , \22818 , \22819 , \22820 , \22821 , \22822 , \22823 , \22824 ,
         \22825 , \22826 , \22827 , \22828 , \22829 , \22830 , \22831 , \22832 , \22833 , \22834 ,
         \22835 , \22836 , \22837 , \22838 , \22839 , \22840 , \22841 , \22842 , \22843 , \22844 ,
         \22845 , \22846 , \22847 , \22848 , \22849 , \22850 , \22851 , \22852 , \22853 , \22854 ,
         \22855 , \22856 , \22857 , \22858 , \22859 , \22860 , \22861 , \22862 , \22863 , \22864 ,
         \22865 , \22866 , \22867 , \22868 , \22869 , \22870 , \22871 , \22872 , \22873 , \22874 ,
         \22875 , \22876 , \22877 , \22878 , \22879 , \22880 , \22881 , \22882 , \22883 , \22884 ,
         \22885 , \22886 , \22887 , \22888 , \22889 , \22890 , \22891 , \22892 , \22893 , \22894 ,
         \22895_nG705f , \22896 , \22897 , \22898 , \22899 , \22900 , \22901 , \22902 , \22903 , \22904 ,
         \22905 , \22906 , \22907 , \22908 , \22909 , \22910 , \22911 , \22912 , \22913 , \22914 ,
         \22915 , \22916 , \22917 , \22918 , \22919 , \22920 , \22921 , \22922 , \22923 , \22924 ,
         \22925 , \22926 , \22927 , \22928 , \22929 , \22930 , \22931 , \22932 , \22933 , \22934 ,
         \22935 , \22936 , \22937 , \22938 , \22939 , \22940 , \22941 , \22942 , \22943 , \22944 ,
         \22945 , \22946 , \22947 , \22948 , \22949 , \22950 , \22951 , \22952 , \22953 , \22954 ,
         \22955 , \22956 , \22957 , \22958 , \22959 , \22960 , \22961 , \22962 , \22963 , \22964 ,
         \22965 , \22966 , \22967 , \22968 , \22969 , \22970 , \22971 , \22972 , \22973 , \22974 ,
         \22975 , \22976 , \22977 , \22978 , \22979 , \22980 , \22981 , \22982 , \22983 , \22984 ,
         \22985 , \22986 , \22987 , \22988 , \22989 , \22990 , \22991 , \22992 , \22993 , \22994 ,
         \22995 , \22996 , \22997 , \22998 , \22999 , \23000 , \23001 , \23002 , \23003 , \23004 ,
         \23005 , \23006 , \23007 , \23008 , \23009 , \23010 , \23011 , \23012 , \23013 , \23014 ,
         \23015 , \23016 , \23017 , \23018 , \23019 , \23020 , \23021 , \23022 , \23023 , \23024 ,
         \23025 , \23026 , \23027 , \23028 , \23029 , \23030 , \23031 , \23032 , \23033 , \23034 ,
         \23035 , \23036 , \23037 , \23038 , \23039 , \23040 , \23041 , \23042 , \23043 , \23044 ,
         \23045 , \23046 , \23047 , \23048 , \23049 , \23050 , \23051 , \23052 , \23053 , \23054 ,
         \23055 , \23056 , \23057 , \23058 , \23059 , \23060 , \23061 , \23062 , \23063 , \23064 ,
         \23065 , \23066 , \23067 , \23068 , \23069 , \23070 , \23071 , \23072 , \23073 , \23074 ,
         \23075 , \23076 , \23077 , \23078 , \23079 , \23080 , \23081 , \23082 , \23083 , \23084 ,
         \23085 , \23086 , \23087 , \23088 , \23089 , \23090 , \23091 , \23092 , \23093 , \23094 ,
         \23095 , \23096 , \23097 , \23098 , \23099 , \23100 , \23101 , \23102 , \23103 , \23104 ,
         \23105 , \23106 , \23107 , \23108 , \23109 , \23110 , \23111 , \23112 , \23113 , \23114 ,
         \23115 , \23116 , \23117 , \23118 , \23119 , \23120 , \23121 , \23122 , \23123 , \23124 ,
         \23125 , \23126 , \23127 , \23128 , \23129 , \23130 , \23131 , \23132 , \23133 , \23134 ,
         \23135 , \23136 , \23137 , \23138 , \23139 , \23140 , \23141 , \23142 , \23143 , \23144 ,
         \23145 , \23146 , \23147 , \23148 , \23149 , \23150 , \23151 , \23152 , \23153 , \23154 ,
         \23155 , \23156 , \23157 , \23158 , \23159 , \23160 , \23161 , \23162 , \23163 , \23164 ,
         \23165 , \23166 , \23167 , \23168 , \23169 , \23170 , \23171 , \23172 , \23173 , \23174 ,
         \23175 , \23176 , \23177 , \23178 , \23179 , \23180 , \23181 , \23182 , \23183 , \23184 ,
         \23185 , \23186 , \23187 , \23188 , \23189 , \23190 , \23191 , \23192 , \23193 , \23194 ,
         \23195 , \23196 , \23197 , \23198 , \23199 , \23200 , \23201 , \23202 , \23203 , \23204 ,
         \23205 , \23206 , \23207 , \23208 , \23209 , \23210 , \23211 , \23212 , \23213 , \23214 ,
         \23215 , \23216 , \23217 , \23218 , \23219 , \23220 , \23221 , \23222 , \23223 , \23224 ,
         \23225 , \23226 , \23227 , \23228 , \23229 , \23230 , \23231 , \23232 , \23233 , \23234 ,
         \23235 , \23236 , \23237 , \23238 , \23239 , \23240 , \23241 , \23242 , \23243 , \23244 ,
         \23245 , \23246 , \23247 , \23248 , \23249 , \23250 , \23251 , \23252 , \23253 , \23254 ,
         \23255 , \23256 , \23257 , \23258 , \23259 , \23260 , \23261 , \23262 , \23263 , \23264 ,
         \23265 , \23266 , \23267 , \23268 , \23269 , \23270 , \23271 , \23272 , \23273 , \23274 ,
         \23275 , \23276 , \23277 , \23278 , \23279 , \23280 , \23281 , \23282 , \23283 , \23284 ,
         \23285 , \23286 , \23287 , \23288 , \23289 , \23290 , \23291 , \23292 , \23293 , \23294 ,
         \23295 , \23296 , \23297 , \23298 , \23299 , \23300 , \23301 , \23302 , \23303 , \23304 ,
         \23305 , \23306 , \23307 , \23308 , \23309 , \23310 , \23311 , \23312 , \23313 , \23314 ,
         \23315 , \23316 , \23317 , \23318 , \23319 , \23320 , \23321 , \23322 , \23323 , \23324 ,
         \23325 , \23326 , \23327 , \23328 , \23329 , \23330 , \23331 , \23332 , \23333 , \23334 ,
         \23335 , \23336 , \23337 , \23338 , \23339 , \23340 , \23341 , \23342 , \23343 , \23344 ,
         \23345 , \23346 , \23347 , \23348 , \23349 , \23350 , \23351 , \23352 , \23353 , \23354 ,
         \23355 , \23356 , \23357 , \23358 , \23359 , \23360 , \23361 , \23362 , \23363 , \23364 ,
         \23365 , \23366 , \23367 , \23368 , \23369 , \23370 , \23371 , \23372 , \23373 , \23374 ,
         \23375 , \23376 , \23377 , \23378 , \23379 , \23380 , \23381 , \23382 , \23383 , \23384 ,
         \23385 , \23386 , \23387 , \23388 , \23389 , \23390 , \23391 , \23392 , \23393 , \23394 ,
         \23395 , \23396 , \23397 , \23398 , \23399 , \23400 , \23401 , \23402 , \23403 , \23404 ,
         \23405 , \23406_nG725e , \23407 , \23408 , \23409 , \23410 , \23411 , \23412 , \23413 , \23414 ,
         \23415 , \23416 , \23417 , \23418 , \23419 , \23420 , \23421 , \23422 , \23423 , \23424 ,
         \23425 , \23426 , \23427_nG7273 , \23428 , \23429 , \23430 , \23431 , \23432 , \23433 , \23434 ,
         \23435 , \23436 , \23437 , \23438 , \23439 , \23440 , \23441 , \23442 , \23443 , \23444 ,
         \23445 , \23446 , \23447 , \23448 , \23449_nG7289 , \23450 , \23451 , \23452 , \23453 , \23454 ,
         \23455 , \23456 , \23457 , \23458 , \23459 , \23460 , \23461 , \23462 , \23463 , \23464 ,
         \23465 , \23466 , \23467 , \23468 , \23469 , \23470 , \23471_nG729f , \23472 , \23473 , \23474 ,
         \23475 , \23476 , \23477 , \23478 , \23479 , \23480 , \23481 , \23482 , \23483 , \23484 ,
         \23485 , \23486 , \23487 , \23488 , \23489 , \23490 , \23491 , \23492 , \23493_nG72b5 , \23494 ,
         \23495 , \23496 , \23497 , \23498 , \23499 , \23500 , \23501 , \23502 , \23503 , \23504 ,
         \23505 , \23506 , \23507 , \23508 , \23509 , \23510 , \23511 , \23512 , \23513 , \23514 ,
         \23515_nG72cb , \23516 , \23517 , \23518 , \23519 , \23520 , \23521 , \23522 , \23523 , \23524 ,
         \23525 , \23526 , \23527 , \23528 , \23529 , \23530 , \23531 , \23532 , \23533 , \23534 ,
         \23535 , \23536 , \23537_nG72e1 , \23538 , \23539 , \23540 , \23541 , \23542 , \23543 , \23544 ,
         \23545 , \23546 , \23547 , \23548 , \23549 , \23550 , \23551 , \23552 , \23553 , \23554 ,
         \23555 , \23556 , \23557 , \23558 , \23559_nG72f7 , \23560 , \23561 , \23562 , \23563 , \23564 ,
         \23565 , \23566 , \23567 , \23568 , \23569 , \23570 , \23571 , \23572 , \23573 , \23574 ,
         \23575 , \23576 , \23577 , \23578 , \23579 , \23580 , \23581 , \23582 , \23583 , \23584 ,
         \23585 , \23586 , \23587 , \23588 , \23589 , \23590 , \23591 , \23592 , \23593 , \23594 ,
         \23595 , \23596 , \23597 , \23598 , \23599 , \23600 , \23601 , \23602 , \23603 , \23604 ,
         \23605 , \23606 , \23607 , \23608 , \23609 , \23610 , \23611 , \23612 , \23613 , \23614 ,
         \23615 , \23616 , \23617 , \23618 , \23619 , \23620 , \23621 , \23622 , \23623 , \23624 ,
         \23625 , \23626 , \23627 , \23628 , \23629 , \23630 , \23631 , \23632 , \23633 , \23634 ,
         \23635 , \23636 , \23637 , \23638 , \23639 , \23640 , \23641 , \23642 , \23643 , \23644 ,
         \23645 , \23646 , \23647 , \23648 , \23649 , \23650 , \23651 , \23652 , \23653 , \23654 ,
         \23655 , \23656 , \23657 , \23658 , \23659 , \23660 , \23661 , \23662 , \23663 , \23664 ,
         \23665 , \23666 , \23667 , \23668 , \23669 , \23670 , \23671 , \23672 , \23673 , \23674 ,
         \23675 , \23676 , \23677 , \23678 , \23679 , \23680 , \23681 , \23682 , \23683 , \23684 ,
         \23685 , \23686 , \23687 , \23688 , \23689 , \23690 , \23691 , \23692 , \23693 , \23694 ,
         \23695 , \23696 , \23697 , \23698 , \23699 , \23700 , \23701 , \23702 , \23703 , \23704 ,
         \23705 , \23706 , \23707 , \23708 , \23709 , \23710 , \23711 , \23712 , \23713 , \23714 ,
         \23715 , \23716 , \23717 , \23718 , \23719 , \23720 , \23721 , \23722 , \23723 , \23724 ,
         \23725 , \23726 , \23727 , \23728 , \23729 , \23730 , \23731 , \23732 , \23733 , \23734 ,
         \23735 , \23736 , \23737 , \23738 , \23739 , \23740 , \23741 , \23742 , \23743 , \23744 ,
         \23745 , \23746 , \23747 , \23748 , \23749 , \23750 , \23751 , \23752 , \23753 , \23754 ,
         \23755 , \23756 , \23757 , \23758 , \23759 , \23760 , \23761 , \23762 , \23763 , \23764 ,
         \23765 , \23766 , \23767 , \23768 , \23769 , \23770 , \23771 , \23772 , \23773 , \23774 ,
         \23775 , \23776 , \23777 , \23778 , \23779 , \23780 , \23781 , \23782 , \23783 , \23784 ,
         \23785 , \23786 , \23787 , \23788 , \23789 , \23790 , \23791 , \23792 , \23793 , \23794 ,
         \23795 , \23796 , \23797 , \23798 , \23799 , \23800 , \23801 , \23802 , \23803 , \23804 ,
         \23805 , \23806 , \23807 , \23808 , \23809 , \23810 , \23811 , \23812 , \23813 , \23814 ,
         \23815 , \23816 , \23817 , \23818 , \23819 , \23820 , \23821 , \23822 , \23823 , \23824 ,
         \23825 , \23826 , \23827 , \23828 , \23829 , \23830 , \23831 , \23832 , \23833 , \23834 ,
         \23835 , \23836 , \23837 , \23838 , \23839 , \23840 , \23841 , \23842 , \23843 , \23844 ,
         \23845 , \23846 , \23847 , \23848 , \23849 , \23850 , \23851 , \23852 , \23853 , \23854 ,
         \23855 , \23856 , \23857 , \23858 , \23859 , \23860 , \23861 , \23862 , \23863 , \23864 ,
         \23865 , \23866 , \23867 , \23868 , \23869 , \23870 , \23871 , \23872 , \23873 , \23874 ,
         \23875 , \23876 , \23877 , \23878 , \23879 , \23880 , \23881 , \23882 , \23883 , \23884 ,
         \23885 , \23886 , \23887 , \23888 , \23889 , \23890 , \23891 , \23892 , \23893 , \23894 ,
         \23895 , \23896 , \23897 , \23898 , \23899 , \23900 , \23901 , \23902 , \23903 , \23904 ,
         \23905 , \23906 , \23907 , \23908 , \23909 , \23910 , \23911 , \23912 , \23913 , \23914 ,
         \23915 , \23916 , \23917 , \23918 , \23919 , \23920 , \23921 , \23922 , \23923 , \23924 ,
         \23925 , \23926 , \23927 , \23928 , \23929 , \23930 , \23931 , \23932 , \23933 , \23934 ,
         \23935 , \23936 , \23937 , \23938 , \23939 , \23940 , \23941 , \23942 , \23943 , \23944 ,
         \23945 , \23946 , \23947 , \23948 , \23949 , \23950 , \23951 , \23952 , \23953 , \23954 ,
         \23955 , \23956 , \23957 , \23958 , \23959 , \23960 , \23961 , \23962 , \23963 , \23964 ,
         \23965 , \23966 , \23967 , \23968 , \23969 , \23970 , \23971 , \23972 , \23973 , \23974 ,
         \23975 , \23976 , \23977 , \23978 , \23979 , \23980 , \23981 , \23982 , \23983 , \23984 ,
         \23985 , \23986 , \23987 , \23988 , \23989 , \23990 , \23991 , \23992 , \23993 , \23994 ,
         \23995 , \23996 , \23997 , \23998 , \23999 , \24000 , \24001 , \24002 , \24003 , \24004 ,
         \24005 , \24006 , \24007 , \24008 , \24009 , \24010 , \24011 , \24012 , \24013 , \24014 ,
         \24015 , \24016 , \24017 , \24018 , \24019 , \24020 , \24021 , \24022 , \24023 , \24024 ,
         \24025 , \24026 , \24027 , \24028 , \24029 , \24030 , \24031 , \24032 , \24033 , \24034 ,
         \24035 , \24036 , \24037 , \24038 , \24039 , \24040 , \24041 , \24042 , \24043 , \24044 ,
         \24045 , \24046 , \24047 , \24048 , \24049 , \24050 , \24051 , \24052 , \24053 , \24054 ,
         \24055 , \24056 , \24057 , \24058 , \24059 , \24060 , \24061 , \24062 , \24063 , \24064 ,
         \24065 , \24066 , \24067 , \24068 , \24069 , \24070 , \24071 , \24072 , \24073 , \24074 ,
         \24075_nG74fb , \24076 , \24077 , \24078 , \24079 , \24080 , \24081 , \24082 , \24083 , \24084 ,
         \24085 , \24086 , \24087 , \24088 , \24089 , \24090 , \24091 , \24092 , \24093 , \24094 ,
         \24095 , \24096_nG7510 , \24097 , \24098 , \24099 , \24100 , \24101 , \24102 , \24103 , \24104 ,
         \24105 , \24106 , \24107 , \24108 , \24109 , \24110 , \24111 , \24112 , \24113 , \24114 ,
         \24115 , \24116 , \24117 , \24118_nG7526 , \24119 , \24120 , \24121 , \24122 , \24123 , \24124 ,
         \24125 , \24126 , \24127 , \24128 , \24129 , \24130 , \24131 , \24132 , \24133 , \24134 ,
         \24135 , \24136 , \24137 , \24138 , \24139 , \24140_nG753c , \24141 , \24142 , \24143 , \24144 ,
         \24145 , \24146 , \24147 , \24148 , \24149 , \24150 , \24151 , \24152 , \24153 , \24154 ,
         \24155 , \24156 , \24157 , \24158 , \24159 , \24160 , \24161 , \24162_nG7552 , \24163 , \24164 ,
         \24165 , \24166 , \24167 , \24168 , \24169 , \24170 , \24171 , \24172 , \24173 , \24174 ,
         \24175 , \24176 , \24177 , \24178 , \24179 , \24180 , \24181 , \24182 , \24183 , \24184_nG7568 ,
         \24185 , \24186 , \24187 , \24188 , \24189 , \24190 , \24191 , \24192 , \24193 , \24194 ,
         \24195 , \24196 , \24197 , \24198 , \24199 , \24200 , \24201 , \24202 , \24203 , \24204 ,
         \24205 , \24206_nG757e , \24207 , \24208 , \24209 , \24210 , \24211 , \24212 , \24213 , \24214 ,
         \24215 , \24216 , \24217 , \24218 , \24219 , \24220 , \24221 , \24222 , \24223 , \24224 ,
         \24225 , \24226 , \24227 , \24228_nG7594 , \24229 , \24230 , \24231 , \24232 , \24233 , \24234 ,
         \24235_nG759b , \24236 , \24237 , \24238 , \24239 , \24240 , \24241 , \24242 , \24243 , \24244 ,
         \24245 , \24246_nG75a6 , \24247 , \24248 , \24249 , \24250 , \24251 , \24252 , \24253 , \24254 ,
         \24255 , \24256 , \24257 , \24258 , \24259 , \24260 , \24261 , \24262 , \24263 , \24264 ,
         \24265 , \24266 , \24267 , \24268 , \24269 , \24270 , \24271 , \24272 , \24273 , \24274 ,
         \24275 , \24276 , \24277 , \24278 , \24279 , \24280 , \24281 , \24282 , \24283 , \24284 ,
         \24285 , \24286 , \24287 , \24288 , \24289 , \24290 , \24291 , \24292 , \24293 , \24294 ,
         \24295 , \24296 , \24297 , \24298 , \24299 , \24300 , \24301 , \24302 , \24303 , \24304_nG75e0 ,
         \24305 , \24306 , \24307 , \24308 , \24309 , \24310 , \24311 , \24312 , \24313 , \24314 ,
         \24315 , \24316 , \24317 , \24318_nG75ee , \24319 , \24320 , \24321 , \24322 , \24323 , \24324 ,
         \24325 , \24326 , \24327 , \24328 , \24329 , \24330 , \24331 , \24332 , \24333_nG75fd , \24334 ,
         \24335 , \24336 , \24337 , \24338 , \24339 , \24340 , \24341 , \24342 , \24343 , \24344 ,
         \24345 , \24346 , \24347 , \24348 , \24349_nG760d , \24350 , \24351 , \24352 , \24353 , \24354 ,
         \24355 , \24356 , \24357 , \24358 , \24359 , \24360 , \24361 , \24362 , \24363 , \24364 ,
         \24365_nG761d , \24366 , \24367 , \24368 , \24369 , \24370 , \24371 , \24372 , \24373 , \24374 ,
         \24375 , \24376 , \24377 , \24378 , \24379 , \24380 , \24381_nG762d , \24382 , \24383 , \24384 ,
         \24385 , \24386 , \24387 , \24388 , \24389 , \24390 , \24391 , \24392 , \24393 , \24394 ,
         \24395 , \24396 , \24397_nG763d , \24398 , \24399 , \24400 , \24401 , \24402 , \24403 , \24404 ,
         \24405 , \24406 , \24407 , \24408 , \24409 , \24410 , \24411 , \24412 , \24413_nG764d , \24414 ,
         \24415 , \24416 , \24417 , \24418 , \24419 , \24420 , \24421 , \24422 , \24423 , \24424 ,
         \24425 , \24426 , \24427 , \24428 , \24429_nG765d , \24430 , \24431 , \24432 , \24433 , \24434 ,
         \24435 , \24436 , \24437 , \24438 , \24439 , \24440 , \24441 , \24442 , \24443 , \24444 ,
         \24445 , \24446 , \24447_nG766f , \24448 , \24449 , \24450 , \24451 , \24452 , \24453 , \24454 ,
         \24455 , \24456 , \24457 , \24458 , \24459 , \24460 , \24461 , \24462_nG767e , \24463 , \24464 ,
         \24465 , \24466 , \24467 , \24468 , \24469 , \24470 , \24471 , \24472 , \24473 , \24474 ,
         \24475 , \24476 , \24477 , \24478_nG768e , \24479 , \24480 , \24481 , \24482 , \24483 , \24484 ,
         \24485 , \24486 , \24487 , \24488 , \24489 , \24490 , \24491 , \24492 , \24493 , \24494_nG769e ,
         \24495 , \24496 , \24497 , \24498 , \24499 , \24500 , \24501 , \24502 , \24503 , \24504 ,
         \24505 , \24506 , \24507 , \24508 , \24509 , \24510_nG76ae , \24511 , \24512 , \24513 , \24514 ,
         \24515 , \24516 , \24517 , \24518 , \24519 , \24520 , \24521 , \24522 , \24523 , \24524 ,
         \24525 , \24526_nG76be , \24527 , \24528 , \24529 , \24530 , \24531 , \24532 , \24533 , \24534 ,
         \24535 , \24536 , \24537 , \24538 , \24539 , \24540 , \24541 , \24542_nG76ce , \24543 , \24544 ,
         \24545 , \24546 , \24547 , \24548 , \24549 , \24550 , \24551 , \24552 , \24553 , \24554 ,
         \24555 , \24556 , \24557 , \24558_nG76de , \24559 , \24560 , \24561 , \24562 , \24563 , \24564 ,
         \24565 , \24566_nG76e6 , \24567 , \24568 , \24569 , \24570 , \24571 , \24572 , \24573 , \24574 ,
         \24575 , \24576 , \24577 , \24578 , \24579 , \24580 , \24581 , \24582 , \24583 , \24584 ,
         \24585 , \24586 , \24587 , \24588 , \24589 , \24590 , \24591 , \24592 , \24593 , \24594 ,
         \24595 , \24596 , \24597 , \24598 , \24599 , \24600 , \24601 , \24602 , \24603 , \24604 ,
         \24605 , \24606 , \24607 , \24608 , \24609 , \24610 , \24611 , \24612 , \24613 , \24614 ,
         \24615 , \24616 , \24617 , \24618 , \24619 , \24620 , \24621 , \24622 , \24623 , \24624 ,
         \24625 , \24626 , \24627 , \24628 , \24629 , \24630 , \24631 , \24632 , \24633 , \24634 ,
         \24635 , \24636 , \24637 , \24638 , \24639 , \24640 , \24641 , \24642 , \24643 , \24644 ,
         \24645 , \24646 , \24647 , \24648 , \24649 , \24650 , \24651 , \24652 , \24653 , \24654 ,
         \24655 , \24656 , \24657 , \24658 , \24659 , \24660 , \24661 , \24662 , \24663 , \24664 ,
         \24665 , \24666 , \24667 , \24668 , \24669 , \24670 , \24671 , \24672 , \24673 , \24674 ,
         \24675 , \24676 , \24677 , \24678 , \24679 , \24680 , \24681 , \24682 , \24683 , \24684 ,
         \24685 , \24686 , \24687 , \24688 , \24689 , \24690 , \24691 , \24692 , \24693 , \24694 ,
         \24695 , \24696 , \24697 , \24698 , \24699 , \24700 , \24701 , \24702 , \24703 , \24704 ,
         \24705 , \24706 , \24707 , \24708 , \24709 , \24710 , \24711 , \24712 , \24713 , \24714 ,
         \24715 , \24716 , \24717 , \24718 , \24719 , \24720 , \24721 , \24722 , \24723 , \24724 ,
         \24725 , \24726 , \24727 , \24728 , \24729 , \24730 , \24731 , \24732 , \24733 , \24734 ,
         \24735 , \24736 , \24737 , \24738 , \24739 , \24740 , \24741 , \24742 , \24743 , \24744 ,
         \24745 , \24746 , \24747 , \24748 , \24749 , \24750 , \24751 , \24752 , \24753 , \24754 ,
         \24755 , \24756 , \24757 , \24758 , \24759 , \24760 , \24761 , \24762 , \24763 , \24764 ,
         \24765 , \24766 , \24767 , \24768 , \24769 , \24770 , \24771 , \24772 , \24773 , \24774 ,
         \24775 , \24776 , \24777 , \24778 , \24779 , \24780 , \24781 , \24782 , \24783 , \24784 ,
         \24785 , \24786 , \24787 , \24788 , \24789 , \24790 , \24791 , \24792 , \24793 , \24794 ,
         \24795 , \24796 , \24797 , \24798 , \24799 , \24800 , \24801 , \24802 , \24803 , \24804 ,
         \24805 , \24806 , \24807 , \24808 , \24809 , \24810 , \24811 , \24812 , \24813 , \24814 ,
         \24815 , \24816 , \24817 , \24818 , \24819 , \24820 , \24821 , \24822 , \24823 , \24824 ,
         \24825 , \24826 , \24827 , \24828 , \24829 , \24830 , \24831 , \24832 , \24833 , \24834 ,
         \24835 , \24836 , \24837 , \24838 , \24839 , \24840 , \24841 , \24842 , \24843 , \24844 ,
         \24845 , \24846 , \24847 , \24848 , \24849 , \24850 , \24851 , \24852 , \24853 , \24854 ,
         \24855 , \24856 , \24857 , \24858 , \24859 , \24860 , \24861 , \24862 , \24863 , \24864 ,
         \24865 , \24866 , \24867 , \24868 , \24869 , \24870 , \24871 , \24872 , \24873 , \24874 ,
         \24875 , \24876 , \24877 , \24878 , \24879 , \24880 , \24881 , \24882 , \24883 , \24884 ,
         \24885 , \24886 , \24887 , \24888 , \24889 , \24890 , \24891 , \24892 , \24893 , \24894 ,
         \24895 , \24896 , \24897 , \24898 , \24899 , \24900 , \24901 , \24902 , \24903 , \24904 ,
         \24905 , \24906 , \24907 , \24908 , \24909 , \24910 , \24911 , \24912 , \24913 , \24914 ,
         \24915 , \24916 , \24917 , \24918 , \24919 , \24920 , \24921 , \24922 , \24923 , \24924 ,
         \24925 , \24926 , \24927 , \24928 , \24929 , \24930 , \24931 , \24932 , \24933 , \24934 ,
         \24935 , \24936 , \24937 , \24938 , \24939 , \24940 , \24941 , \24942 , \24943 , \24944 ,
         \24945 , \24946 , \24947 , \24948 , \24949 , \24950 , \24951 , \24952 , \24953 , \24954 ,
         \24955 , \24956 , \24957 , \24958 , \24959 , \24960 , \24961 , \24962 , \24963 , \24964 ,
         \24965 , \24966 , \24967 , \24968 , \24969 , \24970 , \24971 , \24972 , \24973 , \24974 ,
         \24975 , \24976 , \24977 , \24978 , \24979 , \24980 , \24981 , \24982 , \24983 , \24984 ,
         \24985 , \24986 , \24987 , \24988 , \24989 , \24990 , \24991 , \24992 , \24993 , \24994 ,
         \24995 , \24996 , \24997 , \24998 , \24999 , \25000 , \25001 , \25002 , \25003 , \25004 ,
         \25005 , \25006 , \25007 , \25008 , \25009 , \25010 , \25011 , \25012 , \25013 , \25014 ,
         \25015 , \25016 , \25017 , \25018 , \25019 , \25020 , \25021 , \25022 , \25023 , \25024 ,
         \25025 , \25026 , \25027 , \25028 , \25029 , \25030 , \25031 , \25032 , \25033 , \25034 ,
         \25035 , \25036 , \25037 , \25038 , \25039 , \25040 , \25041 , \25042 , \25043 , \25044 ,
         \25045 , \25046 , \25047 , \25048 , \25049 , \25050 , \25051 , \25052 , \25053 , \25054 ,
         \25055 , \25056 , \25057 , \25058 , \25059 , \25060 , \25061 , \25062 , \25063 , \25064 ,
         \25065 , \25066 , \25067 , \25068 , \25069 , \25070 , \25071 , \25072 , \25073 , \25074 ,
         \25075 , \25076 , \25077 , \25078 , \25079 , \25080 , \25081 , \25082 , \25083 , \25084 ,
         \25085 , \25086 , \25087 , \25088 , \25089 , \25090 , \25091 , \25092 , \25093_nG78fd , \25094 ,
         \25095 , \25096 , \25097 , \25098 , \25099 , \25100 , \25101 , \25102 , \25103 , \25104 ,
         \25105 , \25106 , \25107 , \25108 , \25109 , \25110 , \25111 , \25112 , \25113 , \25114 ,
         \25115 , \25116 , \25117 , \25118 , \25119 , \25120 , \25121 , \25122 , \25123 , \25124 ,
         \25125 , \25126 , \25127 , \25128 , \25129 , \25130 , \25131 , \25132 , \25133 , \25134 ,
         \25135 , \25136 , \25137 , \25138 , \25139 , \25140 , \25141 , \25142 , \25143 , \25144 ,
         \25145 , \25146 , \25147 , \25148 , \25149 , \25150 , \25151 , \25152 , \25153 , \25154 ,
         \25155 , \25156 , \25157 , \25158 , \25159 , \25160 , \25161 , \25162 , \25163 , \25164 ,
         \25165 , \25166 , \25167 , \25168 , \25169 , \25170 , \25171 , \25172 , \25173 , \25174 ,
         \25175 , \25176 , \25177 , \25178 , \25179 , \25180 , \25181 , \25182 , \25183 , \25184 ,
         \25185 , \25186 , \25187 , \25188 , \25189 , \25190 , \25191 , \25192 , \25193 , \25194 ,
         \25195 , \25196 , \25197 , \25198 , \25199 , \25200 , \25201 , \25202 , \25203 , \25204 ,
         \25205 , \25206 , \25207 , \25208 , \25209 , \25210 , \25211 , \25212 , \25213 , \25214 ,
         \25215 , \25216 , \25217 , \25218 , \25219 , \25220 , \25221 , \25222 , \25223 , \25224 ,
         \25225 , \25226 , \25227 , \25228 , \25229 , \25230 , \25231 , \25232 , \25233 , \25234 ,
         \25235 , \25236 , \25237 , \25238 , \25239 , \25240 , \25241 , \25242 , \25243 , \25244 ,
         \25245 , \25246 , \25247 , \25248 , \25249 , \25250 , \25251 , \25252 , \25253 , \25254 ,
         \25255 , \25256 , \25257 , \25258 , \25259 , \25260 , \25261 , \25262 , \25263 , \25264 ,
         \25265 , \25266 , \25267 , \25268 , \25269 , \25270 , \25271 , \25272 , \25273 , \25274 ,
         \25275 , \25276 , \25277 , \25278 , \25279 , \25280 , \25281 , \25282 , \25283 , \25284 ,
         \25285 , \25286 , \25287 , \25288 , \25289 , \25290 , \25291 , \25292 , \25293 , \25294 ,
         \25295 , \25296 , \25297 , \25298 , \25299 , \25300 , \25301 , \25302 , \25303 , \25304 ,
         \25305 , \25306 , \25307 , \25308 , \25309 , \25310 , \25311 , \25312 , \25313 , \25314 ,
         \25315 , \25316 , \25317 , \25318 , \25319 , \25320 , \25321 , \25322 , \25323 , \25324 ,
         \25325 , \25326 , \25327 , \25328 , \25329 , \25330 , \25331 , \25332 , \25333 , \25334 ,
         \25335 , \25336 , \25337 , \25338 , \25339 , \25340 , \25341 , \25342 , \25343 , \25344 ,
         \25345 , \25346 , \25347 , \25348 , \25349 , \25350 , \25351 , \25352 , \25353 , \25354 ,
         \25355 , \25356 , \25357 , \25358 , \25359 , \25360 , \25361 , \25362 , \25363 , \25364 ,
         \25365 , \25366 , \25367 , \25368 , \25369 , \25370 , \25371 , \25372 , \25373 , \25374 ,
         \25375 , \25376 , \25377 , \25378 , \25379 , \25380 , \25381 , \25382 , \25383 , \25384 ,
         \25385 , \25386 , \25387 , \25388 , \25389 , \25390 , \25391 , \25392 , \25393 , \25394 ,
         \25395 , \25396 , \25397 , \25398 , \25399 , \25400 , \25401 , \25402 , \25403 , \25404 ,
         \25405 , \25406 , \25407 , \25408 , \25409 , \25410 , \25411 , \25412 , \25413 , \25414 ,
         \25415 , \25416 , \25417 , \25418 , \25419 , \25420 , \25421 , \25422 , \25423 , \25424 ,
         \25425 , \25426 , \25427 , \25428 , \25429 , \25430 , \25431 , \25432 , \25433 , \25434 ,
         \25435 , \25436 , \25437 , \25438 , \25439 , \25440 , \25441 , \25442 , \25443 , \25444 ,
         \25445 , \25446 , \25447 , \25448 , \25449 , \25450 , \25451 , \25452 , \25453 , \25454 ,
         \25455 , \25456 , \25457 , \25458 , \25459 , \25460 , \25461 , \25462 , \25463 , \25464 ,
         \25465 , \25466 , \25467 , \25468 , \25469 , \25470 , \25471 , \25472 , \25473 , \25474 ,
         \25475 , \25476 , \25477 , \25478 , \25479 , \25480 , \25481 , \25482 , \25483 , \25484 ,
         \25485 , \25486 , \25487 , \25488 , \25489 , \25490 , \25491 , \25492 , \25493 , \25494 ,
         \25495 , \25496 , \25497 , \25498 , \25499 , \25500 , \25501 , \25502 , \25503 , \25504 ,
         \25505 , \25506 , \25507 , \25508 , \25509 , \25510 , \25511 , \25512 , \25513 , \25514 ,
         \25515 , \25516 , \25517 , \25518 , \25519 , \25520 , \25521 , \25522 , \25523 , \25524 ,
         \25525 , \25526 , \25527 , \25528 , \25529 , \25530 , \25531 , \25532 , \25533 , \25534 ,
         \25535 , \25536 , \25537 , \25538 , \25539 , \25540 , \25541 , \25542 , \25543 , \25544 ,
         \25545 , \25546 , \25547 , \25548 , \25549 , \25550 , \25551 , \25552 , \25553 , \25554 ,
         \25555 , \25556 , \25557 , \25558 , \25559 , \25560 , \25561 , \25562 , \25563 , \25564 ,
         \25565 , \25566 , \25567 , \25568 , \25569 , \25570 , \25571 , \25572 , \25573 , \25574 ,
         \25575 , \25576 , \25577 , \25578 , \25579 , \25580 , \25581 , \25582 , \25583 , \25584 ,
         \25585 , \25586 , \25587 , \25588 , \25589 , \25590 , \25591 , \25592 , \25593 , \25594 ,
         \25595 , \25596 , \25597 , \25598 , \25599 , \25600 , \25601 , \25602 , \25603 , \25604_nG7afc ,
         \25605 , \25606 , \25607 , \25608 , \25609 , \25610 , \25611 , \25612 , \25613 , \25614 ,
         \25615 , \25616 , \25617 , \25618 , \25619 , \25620 , \25621 , \25622 , \25623 , \25624 ,
         \25625_nG7b11 , \25626 , \25627 , \25628 , \25629 , \25630 , \25631 , \25632 , \25633 , \25634 ,
         \25635 , \25636 , \25637 , \25638 , \25639 , \25640 , \25641 , \25642 , \25643 , \25644 ,
         \25645 , \25646 , \25647_nG7b27 , \25648 , \25649 , \25650 , \25651 , \25652 , \25653 , \25654 ,
         \25655 , \25656 , \25657 , \25658 , \25659 , \25660 , \25661 , \25662 , \25663 , \25664 ,
         \25665 , \25666 , \25667 , \25668 , \25669_nG7b3d , \25670 , \25671 , \25672 , \25673 , \25674 ,
         \25675 , \25676 , \25677 , \25678 , \25679 , \25680 , \25681 , \25682 , \25683 , \25684 ,
         \25685 , \25686 , \25687 , \25688 , \25689 , \25690 , \25691_nG7b53 , \25692 , \25693 , \25694 ,
         \25695 , \25696 , \25697 , \25698 , \25699 , \25700 , \25701 , \25702 , \25703 , \25704 ,
         \25705 , \25706 , \25707 , \25708 , \25709 , \25710 , \25711 , \25712 , \25713_nG7b69 , \25714 ,
         \25715 , \25716 , \25717 , \25718 , \25719 , \25720 , \25721 , \25722 , \25723 , \25724 ,
         \25725 , \25726 , \25727 , \25728 , \25729 , \25730 , \25731 , \25732 , \25733 , \25734 ,
         \25735_nG7b7f , \25736 , \25737 , \25738 , \25739 , \25740 , \25741 , \25742 , \25743 , \25744 ,
         \25745 , \25746 , \25747 , \25748 , \25749 , \25750 , \25751 , \25752 , \25753 , \25754 ,
         \25755 , \25756 , \25757_nG7b95 , \25758 , \25759 , \25760 , \25761 , \25762 , \25763 , \25764 ,
         \25765 , \25766 , \25767 , \25768 , \25769 , \25770 , \25771 , \25772 , \25773 , \25774 ,
         \25775 , \25776 , \25777 , \25778 , \25779 , \25780 , \25781 , \25782 , \25783 , \25784 ,
         \25785 , \25786 , \25787 , \25788 , \25789 , \25790 , \25791 , \25792 , \25793 , \25794 ,
         \25795 , \25796 , \25797 , \25798 , \25799 , \25800 , \25801 , \25802 , \25803 , \25804 ,
         \25805 , \25806 , \25807 , \25808 , \25809 , \25810 , \25811 , \25812 , \25813 , \25814 ,
         \25815 , \25816 , \25817 , \25818 , \25819 , \25820 , \25821 , \25822 , \25823 , \25824 ,
         \25825 , \25826 , \25827 , \25828 , \25829 , \25830 , \25831 , \25832 , \25833 , \25834 ,
         \25835 , \25836 , \25837 , \25838 , \25839 , \25840 , \25841 , \25842 , \25843 , \25844 ,
         \25845 , \25846 , \25847 , \25848 , \25849 , \25850 , \25851 , \25852 , \25853 , \25854 ,
         \25855 , \25856 , \25857 , \25858 , \25859 , \25860 , \25861 , \25862 , \25863 , \25864 ,
         \25865 , \25866 , \25867 , \25868 , \25869 , \25870 , \25871 , \25872 , \25873 , \25874 ,
         \25875 , \25876 , \25877 , \25878 , \25879 , \25880 , \25881 , \25882 , \25883 , \25884 ,
         \25885 , \25886 , \25887 , \25888 , \25889 , \25890 , \25891 , \25892 , \25893 , \25894 ,
         \25895 , \25896 , \25897 , \25898 , \25899 , \25900 , \25901 , \25902 , \25903 , \25904 ,
         \25905 , \25906 , \25907 , \25908 , \25909 , \25910 , \25911 , \25912 , \25913 , \25914 ,
         \25915 , \25916 , \25917 , \25918 , \25919 , \25920 , \25921 , \25922 , \25923 , \25924 ,
         \25925 , \25926 , \25927 , \25928 , \25929 , \25930 , \25931 , \25932 , \25933 , \25934 ,
         \25935 , \25936 , \25937 , \25938 , \25939 , \25940 , \25941 , \25942 , \25943 , \25944 ,
         \25945 , \25946 , \25947 , \25948 , \25949 , \25950 , \25951 , \25952 , \25953 , \25954 ,
         \25955 , \25956 , \25957 , \25958 , \25959 , \25960 , \25961 , \25962 , \25963 , \25964 ,
         \25965 , \25966 , \25967 , \25968 , \25969 , \25970 , \25971 , \25972 , \25973 , \25974 ,
         \25975 , \25976 , \25977 , \25978 , \25979 , \25980 , \25981 , \25982 , \25983 , \25984 ,
         \25985 , \25986 , \25987 , \25988 , \25989 , \25990 , \25991 , \25992 , \25993 , \25994 ,
         \25995 , \25996 , \25997 , \25998 , \25999 , \26000 , \26001 , \26002 , \26003 , \26004 ,
         \26005 , \26006 , \26007 , \26008 , \26009 , \26010 , \26011 , \26012 , \26013 , \26014 ,
         \26015 , \26016 , \26017 , \26018 , \26019 , \26020 , \26021 , \26022 , \26023 , \26024 ,
         \26025 , \26026 , \26027 , \26028 , \26029 , \26030 , \26031 , \26032 , \26033 , \26034 ,
         \26035 , \26036 , \26037 , \26038 , \26039 , \26040 , \26041 , \26042 , \26043 , \26044 ,
         \26045 , \26046 , \26047 , \26048 , \26049 , \26050 , \26051 , \26052 , \26053 , \26054 ,
         \26055 , \26056 , \26057 , \26058 , \26059 , \26060 , \26061 , \26062 , \26063 , \26064 ,
         \26065 , \26066 , \26067 , \26068 , \26069 , \26070 , \26071 , \26072 , \26073 , \26074 ,
         \26075 , \26076 , \26077 , \26078 , \26079 , \26080 , \26081 , \26082 , \26083 , \26084 ,
         \26085 , \26086 , \26087 , \26088 , \26089 , \26090 , \26091 , \26092 , \26093 , \26094 ,
         \26095 , \26096 , \26097 , \26098 , \26099 , \26100 , \26101 , \26102 , \26103 , \26104 ,
         \26105 , \26106 , \26107 , \26108 , \26109 , \26110 , \26111 , \26112 , \26113 , \26114 ,
         \26115 , \26116 , \26117 , \26118 , \26119 , \26120 , \26121 , \26122 , \26123 , \26124 ,
         \26125 , \26126 , \26127 , \26128 , \26129 , \26130 , \26131 , \26132 , \26133 , \26134 ,
         \26135 , \26136 , \26137 , \26138 , \26139 , \26140 , \26141 , \26142 , \26143 , \26144 ,
         \26145 , \26146 , \26147 , \26148 , \26149 , \26150 , \26151 , \26152 , \26153 , \26154 ,
         \26155 , \26156 , \26157 , \26158 , \26159 , \26160 , \26161 , \26162 , \26163 , \26164 ,
         \26165 , \26166 , \26167 , \26168 , \26169 , \26170 , \26171 , \26172 , \26173 , \26174 ,
         \26175 , \26176 , \26177 , \26178 , \26179 , \26180 , \26181 , \26182 , \26183 , \26184 ,
         \26185 , \26186 , \26187 , \26188 , \26189 , \26190 , \26191 , \26192 , \26193 , \26194 ,
         \26195 , \26196 , \26197 , \26198 , \26199 , \26200 , \26201 , \26202 , \26203 , \26204 ,
         \26205 , \26206 , \26207 , \26208 , \26209 , \26210 , \26211 , \26212 , \26213 , \26214 ,
         \26215 , \26216 , \26217 , \26218 , \26219 , \26220 , \26221 , \26222 , \26223 , \26224 ,
         \26225 , \26226 , \26227 , \26228 , \26229 , \26230 , \26231 , \26232 , \26233 , \26234 ,
         \26235 , \26236 , \26237 , \26238 , \26239 , \26240 , \26241 , \26242 , \26243 , \26244 ,
         \26245 , \26246 , \26247 , \26248 , \26249 , \26250 , \26251 , \26252 , \26253 , \26254 ,
         \26255 , \26256 , \26257 , \26258 , \26259 , \26260 , \26261 , \26262 , \26263 , \26264 ,
         \26265 , \26266 , \26267 , \26268 , \26269 , \26270 , \26271 , \26272 , \26273_nG7d99 , \26274 ,
         \26275 , \26276 , \26277 , \26278 , \26279 , \26280 , \26281 , \26282 , \26283 , \26284 ,
         \26285 , \26286 , \26287 , \26288 , \26289 , \26290 , \26291 , \26292 , \26293 , \26294_nG7dae ,
         \26295 , \26296 , \26297 , \26298 , \26299 , \26300 , \26301 , \26302 , \26303 , \26304 ,
         \26305 , \26306 , \26307 , \26308 , \26309 , \26310 , \26311 , \26312 , \26313 , \26314 ,
         \26315 , \26316_nG7dc4 , \26317 , \26318 , \26319 , \26320 , \26321 , \26322 , \26323 , \26324 ,
         \26325 , \26326 , \26327 , \26328 , \26329 , \26330 , \26331 , \26332 , \26333 , \26334 ,
         \26335 , \26336 , \26337 , \26338_nG7dda , \26339 , \26340 , \26341 , \26342 , \26343 , \26344 ,
         \26345 , \26346 , \26347 , \26348 , \26349 , \26350 , \26351 , \26352 , \26353 , \26354 ,
         \26355 , \26356 , \26357 , \26358 , \26359 , \26360_nG7df0 , \26361 , \26362 , \26363 , \26364 ,
         \26365 , \26366 , \26367 , \26368 , \26369 , \26370 , \26371 , \26372 , \26373 , \26374 ,
         \26375 , \26376 , \26377 , \26378 , \26379 , \26380 , \26381 , \26382_nG7e06 , \26383 , \26384 ,
         \26385 , \26386 , \26387 , \26388 , \26389 , \26390 , \26391 , \26392 , \26393 , \26394 ,
         \26395 , \26396 , \26397 , \26398 , \26399 , \26400 , \26401 , \26402 , \26403 , \26404_nG7e1c ,
         \26405 , \26406 , \26407 , \26408 , \26409 , \26410 , \26411 , \26412 , \26413 , \26414 ,
         \26415 , \26416 , \26417 , \26418 , \26419 , \26420 , \26421 , \26422 , \26423 , \26424 ,
         \26425 , \26426_nG7e32 , \26427 , \26428 , \26429 , \26430 , \26431 , \26432 , \26433_nG7e39 , \26434 ,
         \26435 , \26436 , \26437 , \26438 , \26439 , \26440 , \26441 , \26442 , \26443 , \26444_nG7e44 ,
         \26445 , \26446 , \26447 , \26448 , \26449 , \26450 , \26451 , \26452 , \26453 , \26454 ,
         \26455 , \26456 , \26457 , \26458 , \26459 , \26460 , \26461 , \26462 , \26463 , \26464 ,
         \26465 , \26466 , \26467 , \26468 , \26469 , \26470 , \26471 , \26472 , \26473 , \26474 ,
         \26475 , \26476 , \26477 , \26478 , \26479 , \26480 , \26481 , \26482 , \26483 , \26484 ,
         \26485 , \26486 , \26487 , \26488 , \26489 , \26490 , \26491 , \26492 , \26493 , \26494 ,
         \26495 , \26496 , \26497 , \26498 , \26499 , \26500 , \26501 , \26502_nG7e7f , \26503 , \26504 ,
         \26505 , \26506 , \26507 , \26508 , \26509 , \26510 , \26511 , \26512 , \26513 , \26514 ,
         \26515 , \26516 , \26517_nG7e8e , \26518 , \26519 , \26520 , \26521 , \26522 , \26523 , \26524 ,
         \26525 , \26526 , \26527 , \26528 , \26529 , \26530 , \26531 , \26532 , \26533_nG7e9e , \26534 ,
         \26535 , \26536 , \26537 , \26538 , \26539 , \26540 , \26541 , \26542 , \26543 , \26544 ,
         \26545 , \26546 , \26547 , \26548 , \26549 , \26550_nG7eaf , \26551 , \26552 , \26553 , \26554 ,
         \26555 , \26556 , \26557 , \26558 , \26559 , \26560 , \26561 , \26562 , \26563 , \26564 ,
         \26565 , \26566 , \26567_nG7ec0 , \26568 , \26569 , \26570 , \26571 , \26572 , \26573 , \26574 ,
         \26575 , \26576 , \26577 , \26578 , \26579 , \26580 , \26581 , \26582 , \26583 , \26584_nG7ed1 ,
         \26585 , \26586 , \26587 , \26588 , \26589 , \26590 , \26591 , \26592 , \26593 , \26594 ,
         \26595 , \26596 , \26597 , \26598 , \26599 , \26600 , \26601_nG7ee2 , \26602 , \26603 , \26604 ,
         \26605 , \26606 , \26607 , \26608 , \26609 , \26610 , \26611 , \26612 , \26613 , \26614 ,
         \26615 , \26616 , \26617 , \26618_nG7ef3 , \26619 , \26620 , \26621 , \26622 , \26623 , \26624 ,
         \26625 , \26626 , \26627 , \26628 , \26629 , \26630 , \26631 , \26632 , \26633 , \26634 ,
         \26635_nG7f04 , \26636 , \26637 , \26638 , \26639 , \26640 , \26641 , \26642 , \26643 , \26644 ,
         \26645 , \26646 , \26647 , \26648 , \26649 , \26650 , \26651 , \26652 , \26653 , \26654_nG7f17 ,
         \26655 , \26656 , \26657 , \26658 , \26659 , \26660 , \26661 , \26662 , \26663 , \26664 ,
         \26665 , \26666 , \26667 , \26668 , \26669 , \26670_nG7f27 , \26671 , \26672 , \26673 , \26674 ,
         \26675 , \26676 , \26677 , \26678 , \26679 , \26680 , \26681 , \26682 , \26683 , \26684 ,
         \26685 , \26686 , \26687_nG7f38 , \26688 , \26689 , \26690 , \26691 , \26692 , \26693 , \26694 ,
         \26695 , \26696 , \26697 , \26698 , \26699 , \26700 , \26701 , \26702 , \26703 , \26704_nG7f49 ,
         \26705 , \26706 , \26707 , \26708 , \26709 , \26710 , \26711 , \26712 , \26713 , \26714 ,
         \26715 , \26716 , \26717 , \26718 , \26719 , \26720 , \26721_nG7f5a , \26722 , \26723 , \26724 ,
         \26725 , \26726 , \26727 , \26728 , \26729 , \26730 , \26731 , \26732 , \26733 , \26734 ,
         \26735 , \26736 , \26737 , \26738_nG7f6b , \26739 , \26740 , \26741 , \26742 , \26743 , \26744 ,
         \26745 , \26746 , \26747 , \26748 , \26749 , \26750 , \26751 , \26752 , \26753 , \26754 ,
         \26755_nG7f7c , \26756 , \26757 , \26758 , \26759 , \26760 , \26761 , \26762 , \26763 , \26764 ,
         \26765 , \26766 , \26767 , \26768 , \26769 , \26770 , \26771 , \26772_nG7f8d , \26773 , \26774 ,
         \26775 , \26776 , \26777 , \26778 , \26779 , \26780_nG7f95 , \26781 , \26782 , \26783 , \26784 ,
         \26785 , \26786 , \26787 , \26788 , \26789 , \26790 , \26791 , \26792 , \26793 , \26794 ,
         \26795 , \26796 , \26797 , \26798 , \26799 , \26800 , \26801 , \26802 , \26803 , \26804 ,
         \26805 , \26806 , \26807 , \26808 , \26809 , \26810 , \26811 , \26812 , \26813 , \26814 ,
         \26815 , \26816 , \26817 , \26818 , \26819 , \26820 , \26821 , \26822 , \26823 , \26824 ,
         \26825 , \26826 , \26827 , \26828 , \26829 , \26830 , \26831 , \26832 , \26833 , \26834 ,
         \26835 , \26836 , \26837 , \26838 , \26839 , \26840 , \26841 , \26842 , \26843 , \26844 ,
         \26845 , \26846 , \26847 , \26848 , \26849 , \26850 , \26851 , \26852 , \26853 , \26854 ,
         \26855 , \26856 , \26857 , \26858 , \26859 , \26860 , \26861 , \26862 , \26863 , \26864 ,
         \26865 , \26866 , \26867 , \26868 , \26869 , \26870 , \26871 , \26872 , \26873 , \26874 ,
         \26875 , \26876 , \26877 , \26878 , \26879 , \26880 , \26881 , \26882 , \26883 , \26884 ,
         \26885 , \26886 , \26887 , \26888 , \26889 , \26890 , \26891 , \26892 , \26893 , \26894 ,
         \26895 , \26896 , \26897 , \26898 , \26899 , \26900 , \26901 , \26902 , \26903 , \26904 ,
         \26905 , \26906 , \26907 , \26908 , \26909 , \26910 , \26911 , \26912 , \26913 , \26914 ,
         \26915 , \26916 , \26917 , \26918 , \26919 , \26920 , \26921 , \26922 , \26923 , \26924 ,
         \26925 , \26926 , \26927 , \26928 , \26929 , \26930 , \26931 , \26932 , \26933 , \26934 ,
         \26935 , \26936 , \26937 , \26938 , \26939 , \26940 , \26941 , \26942 , \26943 , \26944 ,
         \26945 , \26946 , \26947 , \26948 , \26949 , \26950 , \26951 , \26952 , \26953 , \26954 ,
         \26955 , \26956 , \26957 , \26958 , \26959 , \26960 , \26961 , \26962 , \26963 , \26964 ,
         \26965 , \26966 , \26967 , \26968 , \26969 , \26970 , \26971 , \26972 , \26973 , \26974 ,
         \26975 , \26976 , \26977 , \26978 , \26979 , \26980 , \26981 , \26982 , \26983 , \26984 ,
         \26985 , \26986 , \26987 , \26988 , \26989 , \26990 , \26991 , \26992 , \26993 , \26994 ,
         \26995 , \26996 , \26997 , \26998 , \26999 , \27000 , \27001 , \27002 , \27003 , \27004 ,
         \27005 , \27006 , \27007 , \27008 , \27009 , \27010 , \27011 , \27012 , \27013 , \27014 ,
         \27015 , \27016 , \27017 , \27018 , \27019 , \27020 , \27021 , \27022 , \27023 , \27024 ,
         \27025 , \27026 , \27027 , \27028 , \27029 , \27030 , \27031 , \27032 , \27033 , \27034 ,
         \27035 , \27036 , \27037 , \27038 , \27039 , \27040 , \27041 , \27042 , \27043 , \27044 ,
         \27045 , \27046 , \27047 , \27048 , \27049 , \27050 , \27051 , \27052 , \27053 , \27054 ,
         \27055 , \27056 , \27057 , \27058 , \27059 , \27060 , \27061 , \27062 , \27063 , \27064 ,
         \27065 , \27066 , \27067 , \27068 , \27069 , \27070 , \27071 , \27072 , \27073 , \27074 ,
         \27075 , \27076 , \27077 , \27078 , \27079 , \27080 , \27081 , \27082 , \27083 , \27084 ,
         \27085 , \27086 , \27087 , \27088 , \27089 , \27090 , \27091 , \27092 , \27093 , \27094 ,
         \27095 , \27096 , \27097 , \27098 , \27099 , \27100 , \27101 , \27102 , \27103 , \27104 ,
         \27105 , \27106 , \27107 , \27108 , \27109 , \27110 , \27111 , \27112 , \27113 , \27114 ,
         \27115 , \27116 , \27117 , \27118 , \27119 , \27120 , \27121 , \27122 , \27123 , \27124 ,
         \27125 , \27126 , \27127 , \27128 , \27129 , \27130 , \27131 , \27132 , \27133 , \27134 ,
         \27135 , \27136 , \27137 , \27138 , \27139 , \27140 , \27141 , \27142 , \27143 , \27144 ,
         \27145 , \27146 , \27147 , \27148 , \27149 , \27150 , \27151 , \27152 , \27153 , \27154 ,
         \27155 , \27156 , \27157 , \27158 , \27159 , \27160 , \27161 , \27162 , \27163 , \27164 ,
         \27165 , \27166 , \27167 , \27168 , \27169 , \27170 , \27171 , \27172 , \27173 , \27174 ,
         \27175 , \27176 , \27177 , \27178 , \27179 , \27180 , \27181 , \27182 , \27183 , \27184 ,
         \27185 , \27186 , \27187 , \27188 , \27189 , \27190 , \27191 , \27192 , \27193 , \27194 ,
         \27195 , \27196 , \27197 , \27198 , \27199 , \27200 , \27201 , \27202 , \27203 , \27204 ,
         \27205 , \27206 , \27207 , \27208 , \27209 , \27210 , \27211 , \27212 , \27213 , \27214 ,
         \27215 , \27216 , \27217 , \27218 , \27219 , \27220 , \27221 , \27222 , \27223 , \27224 ,
         \27225 , \27226 , \27227 , \27228 , \27229 , \27230 , \27231 , \27232 , \27233 , \27234 ,
         \27235 , \27236 , \27237 , \27238 , \27239 , \27240 , \27241 , \27242 , \27243 , \27244 ,
         \27245 , \27246 , \27247 , \27248 , \27249 , \27250 , \27251 , \27252 , \27253 , \27254 ,
         \27255 , \27256 , \27257 , \27258 , \27259 , \27260 , \27261 , \27262 , \27263 , \27264 ,
         \27265 , \27266 , \27267 , \27268 , \27269 , \27270 , \27271 , \27272 , \27273 , \27274 ,
         \27275 , \27276 , \27277 , \27278 , \27279 , \27280 , \27281 , \27282 , \27283 , \27284 ,
         \27285 , \27286 , \27287 , \27288 , \27289 , \27290 , \27291 , \27292 , \27293 , \27294 ,
         \27295 , \27296 , \27297 , \27298 , \27299 , \27300 , \27301 , \27302 , \27303 , \27304 ,
         \27305 , \27306 , \27307_nG81ac , \27308 , \27309 , \27310 , \27311 , \27312 , \27313 , \27314 ,
         \27315 , \27316 , \27317 , \27318 , \27319 , \27320 , \27321 , \27322 , \27323 , \27324 ,
         \27325 , \27326 , \27327 , \27328 , \27329 , \27330 , \27331 , \27332 , \27333 , \27334 ,
         \27335 , \27336 , \27337 , \27338 , \27339 , \27340 , \27341 , \27342 , \27343 , \27344 ,
         \27345 , \27346 , \27347 , \27348 , \27349 , \27350 , \27351 , \27352 , \27353 , \27354 ,
         \27355 , \27356 , \27357 , \27358 , \27359 , \27360 , \27361 , \27362 , \27363 , \27364 ,
         \27365 , \27366 , \27367 , \27368 , \27369 , \27370 , \27371 , \27372 , \27373 , \27374 ,
         \27375 , \27376 , \27377 , \27378 , \27379 , \27380 , \27381 , \27382 , \27383 , \27384 ,
         \27385 , \27386 , \27387 , \27388 , \27389 , \27390 , \27391 , \27392 , \27393 , \27394 ,
         \27395 , \27396 , \27397 , \27398 , \27399 , \27400 , \27401 , \27402 , \27403 , \27404 ,
         \27405 , \27406 , \27407 , \27408 , \27409 , \27410 , \27411 , \27412 , \27413 , \27414 ,
         \27415 , \27416 , \27417 , \27418 , \27419 , \27420 , \27421 , \27422 , \27423 , \27424 ,
         \27425 , \27426 , \27427 , \27428 , \27429 , \27430 , \27431 , \27432 , \27433 , \27434 ,
         \27435 , \27436 , \27437 , \27438 , \27439 , \27440 , \27441 , \27442 , \27443 , \27444 ,
         \27445 , \27446 , \27447 , \27448 , \27449 , \27450 , \27451 , \27452 , \27453 , \27454 ,
         \27455 , \27456 , \27457 , \27458 , \27459 , \27460 , \27461 , \27462 , \27463 , \27464 ,
         \27465 , \27466 , \27467 , \27468 , \27469 , \27470 , \27471 , \27472 , \27473 , \27474 ,
         \27475 , \27476 , \27477 , \27478 , \27479 , \27480 , \27481 , \27482 , \27483 , \27484 ,
         \27485 , \27486 , \27487 , \27488 , \27489 , \27490 , \27491 , \27492 , \27493 , \27494 ,
         \27495 , \27496 , \27497 , \27498 , \27499 , \27500 , \27501 , \27502 , \27503 , \27504 ,
         \27505 , \27506 , \27507 , \27508 , \27509 , \27510 , \27511 , \27512 , \27513 , \27514 ,
         \27515 , \27516 , \27517 , \27518 , \27519 , \27520 , \27521 , \27522 , \27523 , \27524 ,
         \27525 , \27526 , \27527 , \27528 , \27529 , \27530 , \27531 , \27532 , \27533 , \27534 ,
         \27535 , \27536 , \27537 , \27538 , \27539 , \27540 , \27541 , \27542 , \27543 , \27544 ,
         \27545 , \27546 , \27547 , \27548 , \27549 , \27550 , \27551 , \27552 , \27553 , \27554 ,
         \27555 , \27556 , \27557 , \27558 , \27559 , \27560 , \27561 , \27562 , \27563 , \27564 ,
         \27565 , \27566 , \27567 , \27568 , \27569 , \27570 , \27571 , \27572 , \27573 , \27574 ,
         \27575 , \27576 , \27577 , \27578 , \27579 , \27580 , \27581 , \27582 , \27583 , \27584 ,
         \27585 , \27586 , \27587 , \27588 , \27589 , \27590 , \27591 , \27592 , \27593 , \27594 ,
         \27595 , \27596 , \27597 , \27598 , \27599 , \27600 , \27601 , \27602 , \27603 , \27604 ,
         \27605 , \27606 , \27607 , \27608 , \27609 , \27610 , \27611 , \27612 , \27613 , \27614 ,
         \27615 , \27616 , \27617 , \27618 , \27619 , \27620 , \27621 , \27622 , \27623 , \27624 ,
         \27625 , \27626 , \27627 , \27628 , \27629 , \27630 , \27631 , \27632 , \27633 , \27634 ,
         \27635 , \27636 , \27637 , \27638 , \27639 , \27640 , \27641 , \27642 , \27643 , \27644 ,
         \27645 , \27646 , \27647 , \27648 , \27649 , \27650 , \27651 , \27652 , \27653 , \27654 ,
         \27655 , \27656 , \27657 , \27658 , \27659 , \27660 , \27661 , \27662 , \27663 , \27664 ,
         \27665 , \27666 , \27667 , \27668 , \27669 , \27670 , \27671 , \27672 , \27673 , \27674 ,
         \27675 , \27676 , \27677 , \27678 , \27679 , \27680 , \27681 , \27682 , \27683 , \27684 ,
         \27685 , \27686 , \27687 , \27688 , \27689 , \27690 , \27691 , \27692 , \27693 , \27694 ,
         \27695 , \27696 , \27697 , \27698 , \27699 , \27700 , \27701 , \27702 , \27703 , \27704 ,
         \27705 , \27706 , \27707 , \27708 , \27709 , \27710 , \27711 , \27712 , \27713 , \27714 ,
         \27715 , \27716 , \27717 , \27718 , \27719 , \27720 , \27721 , \27722 , \27723 , \27724 ,
         \27725 , \27726 , \27727 , \27728 , \27729 , \27730 , \27731 , \27732 , \27733 , \27734 ,
         \27735 , \27736 , \27737 , \27738 , \27739 , \27740 , \27741 , \27742 , \27743 , \27744 ,
         \27745 , \27746 , \27747 , \27748 , \27749 , \27750 , \27751 , \27752 , \27753 , \27754 ,
         \27755 , \27756 , \27757 , \27758 , \27759 , \27760 , \27761 , \27762 , \27763 , \27764 ,
         \27765 , \27766 , \27767 , \27768 , \27769 , \27770 , \27771 , \27772 , \27773 , \27774 ,
         \27775 , \27776 , \27777 , \27778 , \27779 , \27780 , \27781 , \27782 , \27783 , \27784 ,
         \27785 , \27786 , \27787 , \27788 , \27789 , \27790 , \27791 , \27792 , \27793 , \27794 ,
         \27795 , \27796 , \27797 , \27798 , \27799 , \27800 , \27801 , \27802 , \27803 , \27804 ,
         \27805 , \27806 , \27807 , \27808 , \27809 , \27810 , \27811 , \27812 , \27813 , \27814 ,
         \27815 , \27816 , \27817 , \27818_nG83ab , \27819 , \27820 , \27821 , \27822 , \27823 , \27824 ,
         \27825 , \27826 , \27827 , \27828 , \27829 , \27830 , \27831 , \27832 , \27833 , \27834 ,
         \27835 , \27836 , \27837 , \27838 , \27839_nG83c0 , \27840 , \27841 , \27842 , \27843 , \27844 ,
         \27845 , \27846 , \27847 , \27848 , \27849 , \27850 , \27851 , \27852 , \27853 , \27854 ,
         \27855 , \27856 , \27857 , \27858 , \27859 , \27860 , \27861_nG83d6 , \27862 , \27863 , \27864 ,
         \27865 , \27866 , \27867 , \27868 , \27869 , \27870 , \27871 , \27872 , \27873 , \27874 ,
         \27875 , \27876 , \27877 , \27878 , \27879 , \27880 , \27881 , \27882 , \27883_nG83ec , \27884 ,
         \27885 , \27886 , \27887 , \27888 , \27889 , \27890 , \27891 , \27892 , \27893 , \27894 ,
         \27895 , \27896 , \27897 , \27898 , \27899 , \27900 , \27901 , \27902 , \27903 , \27904 ,
         \27905_nG8402 , \27906 , \27907 , \27908 , \27909 , \27910 , \27911 , \27912 , \27913 , \27914 ,
         \27915 , \27916 , \27917 , \27918 , \27919 , \27920 , \27921 , \27922 , \27923 , \27924 ,
         \27925 , \27926 , \27927_nG8418 , \27928 , \27929 , \27930 , \27931 , \27932 , \27933 , \27934 ,
         \27935 , \27936 , \27937 , \27938 , \27939 , \27940 , \27941 , \27942 , \27943 , \27944 ,
         \27945 , \27946 , \27947 , \27948 , \27949_nG842e , \27950 , \27951 , \27952 , \27953 , \27954 ,
         \27955 , \27956 , \27957 , \27958 , \27959 , \27960 , \27961 , \27962 , \27963 , \27964 ,
         \27965 , \27966 , \27967 , \27968 , \27969 , \27970 , \27971_nG8444 , \27972 , \27973 , \27974 ,
         \27975 , \27976 , \27977 , \27978 , \27979 , \27980 , \27981 , \27982 , \27983 , \27984 ,
         \27985 , \27986 , \27987 , \27988 , \27989 , \27990 , \27991 , \27992 , \27993 , \27994 ,
         \27995 , \27996 , \27997 , \27998 , \27999 , \28000 , \28001 , \28002 , \28003 , \28004 ,
         \28005 , \28006 , \28007 , \28008 , \28009 , \28010 , \28011 , \28012 , \28013 , \28014 ,
         \28015 , \28016 , \28017 , \28018 , \28019 , \28020 , \28021 , \28022 , \28023 , \28024 ,
         \28025 , \28026 , \28027 , \28028 , \28029 , \28030 , \28031 , \28032 , \28033 , \28034 ,
         \28035 , \28036 , \28037 , \28038 , \28039 , \28040 , \28041 , \28042 , \28043 , \28044 ,
         \28045 , \28046 , \28047 , \28048 , \28049 , \28050 , \28051 , \28052 , \28053 , \28054 ,
         \28055 , \28056 , \28057 , \28058 , \28059 , \28060 , \28061 , \28062 , \28063 , \28064 ,
         \28065 , \28066 , \28067 , \28068 , \28069 , \28070 , \28071 , \28072 , \28073 , \28074 ,
         \28075 , \28076 , \28077 , \28078 , \28079 , \28080 , \28081 , \28082 , \28083 , \28084 ,
         \28085 , \28086 , \28087 , \28088 , \28089 , \28090 , \28091 , \28092 , \28093 , \28094 ,
         \28095 , \28096 , \28097 , \28098 , \28099 , \28100 , \28101 , \28102 , \28103 , \28104 ,
         \28105 , \28106 , \28107 , \28108 , \28109 , \28110 , \28111 , \28112 , \28113 , \28114 ,
         \28115 , \28116 , \28117 , \28118 , \28119 , \28120 , \28121 , \28122 , \28123 , \28124 ,
         \28125 , \28126 , \28127 , \28128 , \28129 , \28130 , \28131 , \28132 , \28133 , \28134 ,
         \28135 , \28136 , \28137 , \28138 , \28139 , \28140 , \28141 , \28142 , \28143 , \28144 ,
         \28145 , \28146 , \28147 , \28148 , \28149 , \28150 , \28151 , \28152 , \28153 , \28154 ,
         \28155 , \28156 , \28157 , \28158 , \28159 , \28160 , \28161 , \28162 , \28163 , \28164 ,
         \28165 , \28166 , \28167 , \28168 , \28169 , \28170 , \28171 , \28172 , \28173 , \28174 ,
         \28175 , \28176 , \28177 , \28178 , \28179 , \28180 , \28181 , \28182 , \28183 , \28184 ,
         \28185 , \28186 , \28187 , \28188 , \28189 , \28190 , \28191 , \28192 , \28193 , \28194 ,
         \28195 , \28196 , \28197 , \28198 , \28199 , \28200 , \28201 , \28202 , \28203 , \28204 ,
         \28205 , \28206 , \28207 , \28208 , \28209 , \28210 , \28211 , \28212 , \28213 , \28214 ,
         \28215 , \28216 , \28217 , \28218 , \28219 , \28220 , \28221 , \28222 , \28223 , \28224 ,
         \28225 , \28226 , \28227 , \28228 , \28229 , \28230 , \28231 , \28232 , \28233 , \28234 ,
         \28235 , \28236 , \28237 , \28238 , \28239 , \28240 , \28241 , \28242 , \28243 , \28244 ,
         \28245 , \28246 , \28247 , \28248 , \28249 , \28250 , \28251 , \28252 , \28253 , \28254 ,
         \28255 , \28256 , \28257 , \28258 , \28259 , \28260 , \28261 , \28262 , \28263 , \28264 ,
         \28265 , \28266 , \28267 , \28268 , \28269 , \28270 , \28271 , \28272 , \28273 , \28274 ,
         \28275 , \28276 , \28277 , \28278 , \28279 , \28280 , \28281 , \28282 , \28283 , \28284 ,
         \28285 , \28286 , \28287 , \28288 , \28289 , \28290 , \28291 , \28292 , \28293 , \28294 ,
         \28295 , \28296 , \28297 , \28298 , \28299 , \28300 , \28301 , \28302 , \28303 , \28304 ,
         \28305 , \28306 , \28307 , \28308 , \28309 , \28310 , \28311 , \28312 , \28313 , \28314 ,
         \28315 , \28316 , \28317 , \28318 , \28319 , \28320 , \28321 , \28322 , \28323 , \28324 ,
         \28325 , \28326 , \28327 , \28328 , \28329 , \28330 , \28331 , \28332 , \28333 , \28334 ,
         \28335 , \28336 , \28337 , \28338 , \28339 , \28340 , \28341 , \28342 , \28343 , \28344 ,
         \28345 , \28346 , \28347 , \28348 , \28349 , \28350 , \28351 , \28352 , \28353 , \28354 ,
         \28355 , \28356 , \28357 , \28358 , \28359 , \28360 , \28361 , \28362 , \28363 , \28364 ,
         \28365 , \28366 , \28367 , \28368 , \28369 , \28370 , \28371 , \28372 , \28373 , \28374 ,
         \28375 , \28376 , \28377 , \28378 , \28379 , \28380 , \28381 , \28382 , \28383 , \28384 ,
         \28385 , \28386 , \28387 , \28388 , \28389 , \28390 , \28391 , \28392 , \28393 , \28394 ,
         \28395 , \28396 , \28397 , \28398 , \28399 , \28400 , \28401 , \28402 , \28403 , \28404 ,
         \28405 , \28406 , \28407 , \28408 , \28409 , \28410 , \28411 , \28412 , \28413 , \28414 ,
         \28415 , \28416 , \28417 , \28418 , \28419 , \28420 , \28421 , \28422 , \28423 , \28424 ,
         \28425 , \28426 , \28427 , \28428 , \28429 , \28430 , \28431 , \28432 , \28433 , \28434 ,
         \28435 , \28436 , \28437 , \28438 , \28439 , \28440 , \28441 , \28442 , \28443 , \28444 ,
         \28445 , \28446 , \28447 , \28448 , \28449 , \28450 , \28451 , \28452 , \28453 , \28454 ,
         \28455 , \28456 , \28457 , \28458 , \28459 , \28460 , \28461 , \28462 , \28463 , \28464 ,
         \28465 , \28466 , \28467 , \28468 , \28469 , \28470 , \28471 , \28472 , \28473 , \28474 ,
         \28475 , \28476 , \28477 , \28478 , \28479 , \28480 , \28481 , \28482 , \28483 , \28484 ,
         \28485 , \28486 , \28487_nG8648 , \28488 , \28489 , \28490 , \28491 , \28492 , \28493 , \28494 ,
         \28495 , \28496 , \28497 , \28498 , \28499 , \28500 , \28501 , \28502 , \28503 , \28504 ,
         \28505 , \28506 , \28507 , \28508_nG865d , \28509 , \28510 , \28511 , \28512 , \28513 , \28514 ,
         \28515 , \28516 , \28517 , \28518 , \28519 , \28520 , \28521 , \28522 , \28523 , \28524 ,
         \28525 , \28526 , \28527 , \28528 , \28529 , \28530_nG8673 , \28531 , \28532 , \28533 , \28534 ,
         \28535 , \28536 , \28537 , \28538 , \28539 , \28540 , \28541 , \28542 , \28543 , \28544 ,
         \28545 , \28546 , \28547 , \28548 , \28549 , \28550 , \28551 , \28552_nG8689 , \28553 , \28554 ,
         \28555 , \28556 , \28557 , \28558 , \28559 , \28560 , \28561 , \28562 , \28563 , \28564 ,
         \28565 , \28566 , \28567 , \28568 , \28569 , \28570 , \28571 , \28572 , \28573 , \28574_nG869f ,
         \28575 , \28576 , \28577 , \28578 , \28579 , \28580 , \28581 , \28582 , \28583 , \28584 ,
         \28585 , \28586 , \28587 , \28588 , \28589 , \28590 , \28591 , \28592 , \28593 , \28594 ,
         \28595 , \28596_nG86b5 , \28597 , \28598 , \28599 , \28600 , \28601 , \28602 , \28603 , \28604 ,
         \28605 , \28606 , \28607 , \28608 , \28609 , \28610 , \28611 , \28612 , \28613 , \28614 ,
         \28615 , \28616 , \28617 , \28618_nG86cb , \28619 , \28620 , \28621 , \28622 , \28623 , \28624 ,
         \28625 , \28626 , \28627 , \28628 , \28629 , \28630 , \28631 , \28632 , \28633 , \28634 ,
         \28635 , \28636 , \28637 , \28638 , \28639 , \28640_nG86e1 , \28641 , \28642 , \28643 , \28644 ,
         \28645 , \28646 , \28647_nG86e8 , \28648 , \28649 , \28650 , \28651 , \28652 , \28653 , \28654 ,
         \28655 , \28656 , \28657 , \28658_nG86f3 , \28659 , \28660 , \28661 , \28662 , \28663 , \28664 ,
         \28665 , \28666 , \28667 , \28668 , \28669 , \28670 , \28671 , \28672 , \28673 , \28674 ,
         \28675 , \28676 , \28677 , \28678 , \28679 , \28680 , \28681 , \28682 , \28683 , \28684 ,
         \28685 , \28686 , \28687 , \28688 , \28689 , \28690 , \28691 , \28692 , \28693 , \28694 ,
         \28695 , \28696 , \28697 , \28698 , \28699 , \28700 , \28701 , \28702 , \28703 , \28704 ,
         \28705 , \28706 , \28707 , \28708 , \28709 , \28710 , \28711 , \28712 , \28713 , \28714 ,
         \28715 , \28716 , \28717 , \28718 , \28719 , \28720_nG8731 , \28721 , \28722 , \28723 , \28724 ,
         \28725 , \28726 , \28727 , \28728 , \28729 , \28730 , \28731 , \28732 , \28733 , \28734 ,
         \28735 , \28736_nG8741 , \28737 , \28738 , \28739 , \28740 , \28741 , \28742 , \28743 , \28744 ,
         \28745 , \28746 , \28747 , \28748 , \28749 , \28750 , \28751 , \28752 , \28753_nG8752 , \28754 ,
         \28755 , \28756 , \28757 , \28758 , \28759 , \28760 , \28761 , \28762 , \28763 , \28764 ,
         \28765 , \28766 , \28767 , \28768 , \28769 , \28770 , \28771_nG8764 , \28772 , \28773 , \28774 ,
         \28775 , \28776 , \28777 , \28778 , \28779 , \28780 , \28781 , \28782 , \28783 , \28784 ,
         \28785 , \28786 , \28787 , \28788 , \28789_nG8776 , \28790 , \28791 , \28792 , \28793 , \28794 ,
         \28795 , \28796 , \28797 , \28798 , \28799 , \28800 , \28801 , \28802 , \28803 , \28804 ,
         \28805 , \28806 , \28807_nG8788 , \28808 , \28809 , \28810 , \28811 , \28812 , \28813 , \28814 ,
         \28815 , \28816 , \28817 , \28818 , \28819 , \28820 , \28821 , \28822 , \28823 , \28824 ,
         \28825_nG879a , \28826 , \28827 , \28828 , \28829 , \28830 , \28831 , \28832 , \28833 , \28834 ,
         \28835 , \28836 , \28837 , \28838 , \28839 , \28840 , \28841 , \28842 , \28843_nG87ac , \28844 ,
         \28845 , \28846 , \28847 , \28848 , \28849 , \28850 , \28851 , \28852 , \28853 , \28854 ,
         \28855 , \28856 , \28857 , \28858 , \28859 , \28860 , \28861_nG87be , \28862 , \28863 , \28864 ,
         \28865 , \28866 , \28867 , \28868 , \28869 , \28870 , \28871 , \28872 , \28873 , \28874 ,
         \28875 , \28876 , \28877 , \28878 , \28879 , \28880 , \28881_nG87d2 , \28882 , \28883 , \28884 ,
         \28885 , \28886 , \28887 , \28888 , \28889 , \28890 , \28891 , \28892 , \28893 , \28894 ,
         \28895 , \28896 , \28897 , \28898_nG87e3 , \28899 , \28900 , \28901 , \28902 , \28903 , \28904 ,
         \28905 , \28906 , \28907 , \28908 , \28909 , \28910 , \28911 , \28912 , \28913 , \28914 ,
         \28915 , \28916_nG87f5 , \28917 , \28918 , \28919 , \28920 , \28921 , \28922 , \28923 , \28924 ,
         \28925 , \28926 , \28927 , \28928 , \28929 , \28930 , \28931 , \28932 , \28933 , \28934_nG8807 ,
         \28935 , \28936 , \28937 , \28938 , \28939 , \28940 , \28941 , \28942 , \28943 , \28944 ,
         \28945 , \28946 , \28947 , \28948 , \28949 , \28950 , \28951 , \28952_nG8819 , \28953 , \28954 ,
         \28955 , \28956 , \28957 , \28958 , \28959 , \28960 , \28961 , \28962 , \28963 , \28964 ,
         \28965 , \28966 , \28967 , \28968 , \28969 , \28970_nG882b , \28971 , \28972 , \28973 , \28974 ,
         \28975 , \28976 , \28977 , \28978 , \28979 , \28980 , \28981 , \28982 , \28983 , \28984 ,
         \28985 , \28986 , \28987 , \28988_nG883d , \28989 , \28990 , \28991 , \28992 , \28993 , \28994 ,
         \28995 , \28996 , \28997 , \28998 , \28999 , \29000 , \29001 , \29002 , \29003 , \29004 ,
         \29005 , \29006_nG884f , \29007 , \29008 , \29009 , \29010 , \29011 , \29012 , \29013 , \29014_nG8857 ,
         \29015 , \29016 , \29017 , \29018 , \29019 , \29020 , \29021 , \29022 , \29023 , \29024 ,
         \29025 , \29026 , \29027 , \29028 , \29029 , \29030 , \29031 , \29032 , \29033 , \29034 ,
         \29035 , \29036 , \29037 , \29038 , \29039 , \29040 , \29041 , \29042 , \29043 , \29044 ,
         \29045 , \29046 , \29047 , \29048 , \29049 , \29050 , \29051 , \29052 , \29053 , \29054 ,
         \29055 , \29056 , \29057 , \29058 , \29059 , \29060 , \29061 , \29062 , \29063 , \29064 ,
         \29065 , \29066 , \29067 , \29068 , \29069 , \29070 , \29071 , \29072 , \29073 , \29074 ,
         \29075 , \29076 , \29077 , \29078 , \29079 , \29080 , \29081 , \29082 , \29083 , \29084 ,
         \29085 , \29086 , \29087 , \29088 , \29089 , \29090 , \29091 , \29092 , \29093 , \29094 ,
         \29095 , \29096 , \29097 , \29098 , \29099 , \29100 , \29101 , \29102 , \29103 , \29104 ,
         \29105 , \29106 , \29107 , \29108 , \29109 , \29110 , \29111 , \29112 , \29113 , \29114 ,
         \29115 , \29116 , \29117 , \29118 , \29119 , \29120 , \29121 , \29122 , \29123 , \29124 ,
         \29125 , \29126 , \29127 , \29128 , \29129 , \29130 , \29131 , \29132 , \29133 , \29134 ,
         \29135 , \29136 , \29137 , \29138 , \29139 , \29140 , \29141 , \29142 , \29143 , \29144 ,
         \29145 , \29146 , \29147 , \29148 , \29149 , \29150 , \29151 , \29152 , \29153 , \29154 ,
         \29155 , \29156 , \29157 , \29158 , \29159 , \29160 , \29161 , \29162 , \29163 , \29164 ,
         \29165 , \29166 , \29167 , \29168 , \29169 , \29170 , \29171 , \29172 , \29173 , \29174 ,
         \29175 , \29176 , \29177 , \29178 , \29179 , \29180 , \29181 , \29182 , \29183 , \29184 ,
         \29185 , \29186 , \29187 , \29188 , \29189 , \29190 , \29191 , \29192 , \29193 , \29194 ,
         \29195 , \29196 , \29197 , \29198 , \29199 , \29200 , \29201 , \29202 , \29203 , \29204 ,
         \29205 , \29206 , \29207 , \29208 , \29209 , \29210 , \29211 , \29212 , \29213 , \29214 ,
         \29215 , \29216 , \29217 , \29218 , \29219 , \29220 , \29221 , \29222 , \29223 , \29224 ,
         \29225 , \29226 , \29227 , \29228 , \29229 , \29230 , \29231 , \29232 , \29233 , \29234 ,
         \29235 , \29236 , \29237 , \29238 , \29239 , \29240 , \29241 , \29242 , \29243 , \29244 ,
         \29245 , \29246 , \29247 , \29248 , \29249 , \29250 , \29251 , \29252 , \29253 , \29254 ,
         \29255 , \29256 , \29257 , \29258 , \29259 , \29260 , \29261 , \29262 , \29263 , \29264 ,
         \29265 , \29266 , \29267 , \29268 , \29269 , \29270 , \29271 , \29272 , \29273 , \29274 ,
         \29275 , \29276 , \29277 , \29278 , \29279 , \29280 , \29281 , \29282 , \29283 , \29284 ,
         \29285 , \29286 , \29287 , \29288 , \29289 , \29290 , \29291 , \29292 , \29293 , \29294 ,
         \29295 , \29296 , \29297 , \29298 , \29299 , \29300 , \29301 , \29302 , \29303 , \29304 ,
         \29305 , \29306 , \29307 , \29308 , \29309 , \29310 , \29311 , \29312 , \29313 , \29314 ,
         \29315 , \29316 , \29317 , \29318 , \29319 , \29320 , \29321 , \29322 , \29323 , \29324 ,
         \29325 , \29326 , \29327 , \29328 , \29329 , \29330 , \29331 , \29332 , \29333 , \29334 ,
         \29335 , \29336 , \29337 , \29338 , \29339 , \29340 , \29341 , \29342 , \29343 , \29344 ,
         \29345 , \29346 , \29347 , \29348 , \29349 , \29350 , \29351 , \29352 , \29353 , \29354 ,
         \29355 , \29356 , \29357 , \29358 , \29359 , \29360 , \29361 , \29362 , \29363 , \29364 ,
         \29365 , \29366 , \29367 , \29368 , \29369 , \29370 , \29371 , \29372 , \29373 , \29374 ,
         \29375 , \29376 , \29377 , \29378 , \29379 , \29380 , \29381 , \29382 , \29383 , \29384 ,
         \29385 , \29386 , \29387 , \29388 , \29389 , \29390 , \29391 , \29392 , \29393 , \29394 ,
         \29395 , \29396 , \29397 , \29398 , \29399 , \29400 , \29401 , \29402 , \29403 , \29404 ,
         \29405 , \29406 , \29407 , \29408 , \29409 , \29410 , \29411 , \29412 , \29413 , \29414 ,
         \29415 , \29416 , \29417 , \29418 , \29419 , \29420 , \29421 , \29422 , \29423 , \29424 ,
         \29425 , \29426 , \29427 , \29428 , \29429 , \29430 , \29431 , \29432 , \29433 , \29434 ,
         \29435 , \29436 , \29437 , \29438 , \29439 , \29440 , \29441 , \29442 , \29443 , \29444 ,
         \29445 , \29446 , \29447 , \29448 , \29449 , \29450 , \29451 , \29452 , \29453 , \29454 ,
         \29455 , \29456 , \29457 , \29458 , \29459 , \29460 , \29461 , \29462 , \29463 , \29464 ,
         \29465 , \29466 , \29467 , \29468 , \29469 , \29470 , \29471 , \29472 , \29473 , \29474 ,
         \29475 , \29476 , \29477 , \29478 , \29479 , \29480 , \29481 , \29482 , \29483 , \29484 ,
         \29485 , \29486 , \29487 , \29488 , \29489 , \29490 , \29491 , \29492 , \29493 , \29494 ,
         \29495 , \29496 , \29497 , \29498 , \29499 , \29500 , \29501 , \29502 , \29503 , \29504 ,
         \29505 , \29506 , \29507 , \29508 , \29509 , \29510 , \29511 , \29512 , \29513 , \29514 ,
         \29515 , \29516 , \29517 , \29518 , \29519 , \29520 , \29521 , \29522 , \29523 , \29524 ,
         \29525 , \29526 , \29527 , \29528 , \29529 , \29530 , \29531 , \29532 , \29533 , \29534 ,
         \29535 , \29536 , \29537 , \29538 , \29539 , \29540 , \29541_nG8a6e , \29542 , \29543 , \29544 ,
         \29545 , \29546 , \29547 , \29548 , \29549 , \29550 , \29551 , \29552 , \29553 , \29554 ,
         \29555 , \29556 , \29557 , \29558 , \29559 , \29560 , \29561 , \29562 , \29563 , \29564 ,
         \29565 , \29566 , \29567 , \29568 , \29569 , \29570 , \29571 , \29572 , \29573 , \29574 ,
         \29575 , \29576 , \29577 , \29578 , \29579 , \29580 , \29581 , \29582 , \29583 , \29584 ,
         \29585 , \29586 , \29587 , \29588 , \29589 , \29590 , \29591 , \29592 , \29593 , \29594 ,
         \29595 , \29596 , \29597 , \29598 , \29599 , \29600 , \29601 , \29602 , \29603 , \29604 ,
         \29605 , \29606 , \29607 , \29608 , \29609 , \29610 , \29611 , \29612 , \29613 , \29614 ,
         \29615 , \29616 , \29617 , \29618 , \29619 , \29620 , \29621 , \29622 , \29623 , \29624 ,
         \29625 , \29626 , \29627 , \29628 , \29629 , \29630 , \29631 , \29632 , \29633 , \29634 ,
         \29635 , \29636 , \29637 , \29638 , \29639 , \29640 , \29641 , \29642 , \29643 , \29644 ,
         \29645 , \29646 , \29647 , \29648 , \29649 , \29650 , \29651 , \29652 , \29653 , \29654 ,
         \29655 , \29656 , \29657 , \29658 , \29659 , \29660 , \29661 , \29662 , \29663 , \29664 ,
         \29665 , \29666 , \29667 , \29668 , \29669 , \29670 , \29671 , \29672 , \29673 , \29674 ,
         \29675 , \29676 , \29677 , \29678 , \29679 , \29680 , \29681 , \29682 , \29683 , \29684 ,
         \29685 , \29686 , \29687 , \29688 , \29689 , \29690 , \29691 , \29692 , \29693 , \29694 ,
         \29695 , \29696 , \29697 , \29698 , \29699 , \29700 , \29701 , \29702 , \29703 , \29704 ,
         \29705 , \29706 , \29707 , \29708 , \29709 , \29710 , \29711 , \29712 , \29713 , \29714 ,
         \29715 , \29716 , \29717 , \29718 , \29719 , \29720 , \29721 , \29722 , \29723 , \29724 ,
         \29725 , \29726 , \29727 , \29728 , \29729 , \29730 , \29731 , \29732 , \29733 , \29734 ,
         \29735 , \29736 , \29737 , \29738 , \29739 , \29740 , \29741 , \29742 , \29743 , \29744 ,
         \29745 , \29746 , \29747 , \29748 , \29749 , \29750 , \29751 , \29752 , \29753 , \29754 ,
         \29755 , \29756 , \29757 , \29758 , \29759 , \29760 , \29761 , \29762 , \29763 , \29764 ,
         \29765 , \29766 , \29767 , \29768 , \29769 , \29770 , \29771 , \29772 , \29773 , \29774 ,
         \29775 , \29776 , \29777 , \29778 , \29779 , \29780 , \29781 , \29782 , \29783 , \29784 ,
         \29785 , \29786 , \29787 , \29788 , \29789 , \29790 , \29791 , \29792 , \29793 , \29794 ,
         \29795 , \29796 , \29797 , \29798 , \29799 , \29800 , \29801 , \29802 , \29803 , \29804 ,
         \29805 , \29806 , \29807 , \29808 , \29809 , \29810 , \29811 , \29812 , \29813 , \29814 ,
         \29815 , \29816 , \29817 , \29818 , \29819 , \29820 , \29821 , \29822 , \29823 , \29824 ,
         \29825 , \29826 , \29827 , \29828 , \29829 , \29830 , \29831 , \29832 , \29833 , \29834 ,
         \29835 , \29836 , \29837 , \29838 , \29839 , \29840 , \29841 , \29842 , \29843 , \29844 ,
         \29845 , \29846 , \29847 , \29848 , \29849 , \29850 , \29851 , \29852 , \29853 , \29854 ,
         \29855 , \29856 , \29857 , \29858 , \29859 , \29860 , \29861 , \29862 , \29863 , \29864 ,
         \29865 , \29866 , \29867 , \29868 , \29869 , \29870 , \29871 , \29872 , \29873 , \29874 ,
         \29875 , \29876 , \29877 , \29878 , \29879 , \29880 , \29881 , \29882 , \29883 , \29884 ,
         \29885 , \29886 , \29887 , \29888 , \29889 , \29890 , \29891 , \29892 , \29893 , \29894 ,
         \29895 , \29896 , \29897 , \29898 , \29899 , \29900 , \29901 , \29902 , \29903 , \29904 ,
         \29905 , \29906 , \29907 , \29908 , \29909 , \29910 , \29911 , \29912 , \29913 , \29914 ,
         \29915 , \29916 , \29917 , \29918 , \29919 , \29920 , \29921 , \29922 , \29923 , \29924 ,
         \29925 , \29926 , \29927 , \29928 , \29929 , \29930 , \29931 , \29932 , \29933 , \29934 ,
         \29935 , \29936 , \29937 , \29938 , \29939 , \29940 , \29941 , \29942 , \29943 , \29944 ,
         \29945 , \29946 , \29947 , \29948 , \29949 , \29950 , \29951 , \29952 , \29953 , \29954 ,
         \29955 , \29956 , \29957 , \29958 , \29959 , \29960 , \29961 , \29962 , \29963 , \29964 ,
         \29965 , \29966 , \29967 , \29968 , \29969 , \29970 , \29971 , \29972 , \29973 , \29974 ,
         \29975 , \29976 , \29977 , \29978 , \29979 , \29980 , \29981 , \29982 , \29983 , \29984 ,
         \29985 , \29986 , \29987 , \29988 , \29989 , \29990 , \29991 , \29992 , \29993 , \29994 ,
         \29995 , \29996 , \29997 , \29998 , \29999 , \30000 , \30001 , \30002 , \30003 , \30004 ,
         \30005 , \30006 , \30007 , \30008 , \30009 , \30010 , \30011 , \30012 , \30013 , \30014 ,
         \30015 , \30016 , \30017 , \30018 , \30019 , \30020 , \30021 , \30022 , \30023 , \30024 ,
         \30025 , \30026 , \30027 , \30028 , \30029 , \30030 , \30031 , \30032 , \30033 , \30034 ,
         \30035 , \30036 , \30037 , \30038 , \30039 , \30040 , \30041 , \30042 , \30043 , \30044 ,
         \30045 , \30046 , \30047 , \30048 , \30049 , \30050 , \30051 , \30052_nG8c6d , \30053 , \30054 ,
         \30055 , \30056 , \30057 , \30058 , \30059 , \30060 , \30061 , \30062 , \30063 , \30064 ,
         \30065 , \30066 , \30067 , \30068 , \30069 , \30070 , \30071 , \30072 , \30073_nG8c82 , \30074 ,
         \30075 , \30076 , \30077 , \30078 , \30079 , \30080 , \30081 , \30082 , \30083 , \30084 ,
         \30085 , \30086 , \30087 , \30088 , \30089 , \30090 , \30091 , \30092 , \30093 , \30094 ,
         \30095_nG8c98 , \30096 , \30097 , \30098 , \30099 , \30100 , \30101 , \30102 , \30103 , \30104 ,
         \30105 , \30106 , \30107 , \30108 , \30109 , \30110 , \30111 , \30112 , \30113 , \30114 ,
         \30115 , \30116 , \30117_nG8cae , \30118 , \30119 , \30120 , \30121 , \30122 , \30123 , \30124 ,
         \30125 , \30126 , \30127 , \30128 , \30129 , \30130 , \30131 , \30132 , \30133 , \30134 ,
         \30135 , \30136 , \30137 , \30138 , \30139_nG8cc4 , \30140 , \30141 , \30142 , \30143 , \30144 ,
         \30145 , \30146 , \30147 , \30148 , \30149 , \30150 , \30151 , \30152 , \30153 , \30154 ,
         \30155 , \30156 , \30157 , \30158 , \30159 , \30160 , \30161_nG8cda , \30162 , \30163 , \30164 ,
         \30165 , \30166 , \30167 , \30168 , \30169 , \30170 , \30171 , \30172 , \30173 , \30174 ,
         \30175 , \30176 , \30177 , \30178 , \30179 , \30180 , \30181 , \30182 , \30183_nG8cf0 , \30184 ,
         \30185 , \30186 , \30187 , \30188 , \30189 , \30190 , \30191 , \30192 , \30193 , \30194 ,
         \30195 , \30196 , \30197 , \30198 , \30199 , \30200 , \30201 , \30202 , \30203 , \30204 ,
         \30205_nG8d06 , \30206 , \30207 , \30208 , \30209 , \30210 , \30211 , \30212 , \30213 , \30214 ,
         \30215 , \30216 , \30217 , \30218 , \30219 , \30220 , \30221 , \30222 , \30223 , \30224 ,
         \30225 , \30226 , \30227 , \30228 , \30229 , \30230 , \30231 , \30232 , \30233 , \30234 ,
         \30235 , \30236 , \30237 , \30238 , \30239 , \30240 , \30241 , \30242 , \30243 , \30244 ,
         \30245 , \30246 , \30247 , \30248 , \30249 , \30250 , \30251 , \30252 , \30253 , \30254 ,
         \30255 , \30256 , \30257 , \30258 , \30259 , \30260 , \30261 , \30262 , \30263 , \30264 ,
         \30265 , \30266 , \30267 , \30268 , \30269 , \30270 , \30271 , \30272 , \30273 , \30274 ,
         \30275 , \30276 , \30277 , \30278 , \30279 , \30280 , \30281 , \30282 , \30283 , \30284 ,
         \30285 , \30286 , \30287 , \30288 , \30289 , \30290 , \30291 , \30292 , \30293 , \30294 ,
         \30295 , \30296 , \30297 , \30298 , \30299 , \30300 , \30301 , \30302 , \30303 , \30304 ,
         \30305 , \30306 , \30307 , \30308 , \30309 , \30310 , \30311 , \30312 , \30313 , \30314 ,
         \30315 , \30316 , \30317 , \30318 , \30319 , \30320 , \30321 , \30322 , \30323 , \30324 ,
         \30325 , \30326 , \30327 , \30328 , \30329 , \30330 , \30331 , \30332 , \30333 , \30334 ,
         \30335 , \30336 , \30337 , \30338 , \30339 , \30340 , \30341 , \30342 , \30343 , \30344 ,
         \30345 , \30346 , \30347 , \30348 , \30349 , \30350 , \30351 , \30352 , \30353 , \30354 ,
         \30355 , \30356 , \30357 , \30358 , \30359 , \30360 , \30361 , \30362 , \30363 , \30364 ,
         \30365 , \30366 , \30367 , \30368 , \30369 , \30370 , \30371 , \30372 , \30373 , \30374 ,
         \30375 , \30376 , \30377 , \30378 , \30379 , \30380 , \30381 , \30382 , \30383 , \30384 ,
         \30385 , \30386 , \30387 , \30388 , \30389 , \30390 , \30391 , \30392 , \30393 , \30394 ,
         \30395 , \30396 , \30397 , \30398 , \30399 , \30400 , \30401 , \30402 , \30403 , \30404 ,
         \30405 , \30406 , \30407 , \30408 , \30409 , \30410 , \30411 , \30412 , \30413 , \30414 ,
         \30415 , \30416 , \30417 , \30418 , \30419 , \30420 , \30421 , \30422 , \30423 , \30424 ,
         \30425 , \30426 , \30427 , \30428 , \30429 , \30430 , \30431 , \30432 , \30433 , \30434 ,
         \30435 , \30436 , \30437 , \30438 , \30439 , \30440 , \30441 , \30442 , \30443 , \30444 ,
         \30445 , \30446 , \30447 , \30448 , \30449 , \30450 , \30451 , \30452 , \30453 , \30454 ,
         \30455 , \30456 , \30457 , \30458 , \30459 , \30460 , \30461 , \30462 , \30463 , \30464 ,
         \30465 , \30466 , \30467 , \30468 , \30469 , \30470 , \30471 , \30472 , \30473 , \30474 ,
         \30475 , \30476 , \30477 , \30478 , \30479 , \30480 , \30481 , \30482 , \30483 , \30484 ,
         \30485 , \30486 , \30487 , \30488 , \30489 , \30490 , \30491 , \30492 , \30493 , \30494 ,
         \30495 , \30496 , \30497 , \30498 , \30499 , \30500 , \30501 , \30502 , \30503 , \30504 ,
         \30505 , \30506 , \30507 , \30508 , \30509 , \30510 , \30511 , \30512 , \30513 , \30514 ,
         \30515 , \30516 , \30517 , \30518 , \30519 , \30520 , \30521 , \30522 , \30523 , \30524 ,
         \30525 , \30526 , \30527 , \30528 , \30529 , \30530 , \30531 , \30532 , \30533 , \30534 ,
         \30535 , \30536 , \30537 , \30538 , \30539 , \30540 , \30541 , \30542 , \30543 , \30544 ,
         \30545 , \30546 , \30547 , \30548 , \30549 , \30550 , \30551 , \30552 , \30553 , \30554 ,
         \30555 , \30556 , \30557 , \30558 , \30559 , \30560 , \30561 , \30562 , \30563 , \30564 ,
         \30565 , \30566 , \30567 , \30568 , \30569 , \30570 , \30571 , \30572 , \30573 , \30574 ,
         \30575 , \30576 , \30577 , \30578 , \30579 , \30580 , \30581 , \30582 , \30583 , \30584 ,
         \30585 , \30586 , \30587 , \30588 , \30589 , \30590 , \30591 , \30592 , \30593 , \30594 ,
         \30595 , \30596 , \30597 , \30598 , \30599 , \30600 , \30601 , \30602 , \30603 , \30604 ,
         \30605 , \30606 , \30607 , \30608 , \30609 , \30610 , \30611 , \30612 , \30613 , \30614 ,
         \30615 , \30616 , \30617 , \30618 , \30619 , \30620 , \30621 , \30622 , \30623 , \30624 ,
         \30625 , \30626 , \30627 , \30628 , \30629 , \30630 , \30631 , \30632 , \30633 , \30634 ,
         \30635 , \30636 , \30637 , \30638 , \30639 , \30640 , \30641 , \30642 , \30643 , \30644 ,
         \30645 , \30646 , \30647 , \30648 , \30649 , \30650 , \30651 , \30652 , \30653 , \30654 ,
         \30655 , \30656 , \30657 , \30658 , \30659 , \30660 , \30661 , \30662 , \30663 , \30664 ,
         \30665 , \30666 , \30667 , \30668 , \30669 , \30670 , \30671 , \30672 , \30673 , \30674 ,
         \30675 , \30676 , \30677 , \30678 , \30679 , \30680 , \30681 , \30682 , \30683 , \30684 ,
         \30685 , \30686 , \30687 , \30688 , \30689 , \30690 , \30691 , \30692 , \30693 , \30694 ,
         \30695 , \30696 , \30697 , \30698 , \30699 , \30700 , \30701 , \30702 , \30703 , \30704 ,
         \30705 , \30706 , \30707 , \30708 , \30709 , \30710 , \30711 , \30712 , \30713 , \30714 ,
         \30715 , \30716 , \30717 , \30718 , \30719 , \30720 , \30721_nG8f0a , \30722 , \30723 , \30724 ,
         \30725 , \30726 , \30727 , \30728 , \30729 , \30730 , \30731 , \30732 , \30733 , \30734 ,
         \30735 , \30736 , \30737 , \30738 , \30739 , \30740 , \30741 , \30742_nG8f1f , \30743 , \30744 ,
         \30745 , \30746 , \30747 , \30748 , \30749 , \30750 , \30751 , \30752 , \30753 , \30754 ,
         \30755 , \30756 , \30757 , \30758 , \30759 , \30760 , \30761 , \30762 , \30763 , \30764_nG8f35 ,
         \30765 , \30766 , \30767 , \30768 , \30769 , \30770 , \30771 , \30772 , \30773 , \30774 ,
         \30775 , \30776 , \30777 , \30778 , \30779 , \30780 , \30781 , \30782 , \30783 , \30784 ,
         \30785 , \30786_nG8f4b , \30787 , \30788 , \30789 , \30790 , \30791 , \30792 , \30793 , \30794 ,
         \30795 , \30796 , \30797 , \30798 , \30799 , \30800 , \30801 , \30802 , \30803 , \30804 ,
         \30805 , \30806 , \30807 , \30808_nG8f61 , \30809 , \30810 , \30811 , \30812 , \30813 , \30814 ,
         \30815 , \30816 , \30817 , \30818 , \30819 , \30820 , \30821 , \30822 , \30823 , \30824 ,
         \30825 , \30826 , \30827 , \30828 , \30829 , \30830_nG8f77 , \30831 , \30832 , \30833 , \30834 ,
         \30835 , \30836 , \30837 , \30838 , \30839 , \30840 , \30841 , \30842 , \30843 , \30844 ,
         \30845 , \30846 , \30847 , \30848 , \30849 , \30850 , \30851 , \30852_nG8f8d , \30853 , \30854 ,
         \30855 , \30856 , \30857 , \30858 , \30859 , \30860 , \30861 , \30862 , \30863 , \30864 ,
         \30865 , \30866 , \30867 , \30868 , \30869 , \30870 , \30871 , \30872 , \30873 , \30874_nG8fa3 ,
         \30875 , \30876 , \30877 , \30878 , \30879 , \30880 , \30881_nG8faa , \30882 , \30883 , \30884 ,
         \30885 , \30886 , \30887 , \30888 , \30889 , \30890 , \30891 , \30892_nG8fb5 , \30893 , \30894 ,
         \30895 , \30896 , \30897 , \30898 , \30899 , \30900 , \30901 , \30902 , \30903 , \30904 ,
         \30905 , \30906 , \30907 , \30908 , \30909 , \30910 , \30911 , \30912 , \30913 , \30914 ,
         \30915 , \30916 , \30917 , \30918 , \30919 , \30920 , \30921 , \30922 , \30923 , \30924 ,
         \30925 , \30926 , \30927 , \30928 , \30929 , \30930 , \30931 , \30932 , \30933 , \30934 ,
         \30935 , \30936 , \30937 , \30938 , \30939 , \30940 , \30941 , \30942 , \30943 , \30944 ,
         \30945 , \30946 , \30947 , \30948 , \30949 , \30950 , \30951 , \30952_nG8ff3 , \30953 , \30954 ,
         \30955 , \30956 , \30957 , \30958 , \30959 , \30960 , \30961 , \30962 , \30963 , \30964 ,
         \30965 , \30966 , \30967 , \30968 , \30969_nG9004 , \30970 , \30971 , \30972 , \30973 , \30974 ,
         \30975 , \30976 , \30977 , \30978 , \30979 , \30980 , \30981 , \30982 , \30983 , \30984 ,
         \30985 , \30986 , \30987_nG9016 , \30988 , \30989 , \30990 , \30991 , \30992 , \30993 , \30994 ,
         \30995 , \30996 , \30997 , \30998 , \30999 , \31000 , \31001 , \31002 , \31003 , \31004 ,
         \31005 , \31006_nG9029 , \31007 , \31008 , \31009 , \31010 , \31011 , \31012 , \31013 , \31014 ,
         \31015 , \31016 , \31017 , \31018 , \31019 , \31020 , \31021 , \31022 , \31023 , \31024 ,
         \31025_nG903c , \31026 , \31027 , \31028 , \31029 , \31030 , \31031 , \31032 , \31033 , \31034 ,
         \31035 , \31036 , \31037 , \31038 , \31039 , \31040 , \31041 , \31042 , \31043 , \31044_nG904f ,
         \31045 , \31046 , \31047 , \31048 , \31049 , \31050 , \31051 , \31052 , \31053 , \31054 ,
         \31055 , \31056 , \31057 , \31058 , \31059 , \31060 , \31061 , \31062 , \31063_nG9062 , \31064 ,
         \31065 , \31066 , \31067 , \31068 , \31069 , \31070 , \31071 , \31072 , \31073 , \31074 ,
         \31075 , \31076 , \31077 , \31078 , \31079 , \31080 , \31081 , \31082_nG9075 , \31083 , \31084 ,
         \31085 , \31086 , \31087 , \31088 , \31089 , \31090 , \31091 , \31092 , \31093 , \31094 ,
         \31095 , \31096 , \31097 , \31098 , \31099 , \31100 , \31101_nG9088 , \31102 , \31103 , \31104 ,
         \31105 , \31106 , \31107 , \31108 , \31109 , \31110 , \31111 , \31112 , \31113 , \31114 ,
         \31115 , \31116 , \31117 , \31118 , \31119 , \31120 , \31121 , \31122_nG909d , \31123 , \31124 ,
         \31125 , \31126 , \31127 , \31128 , \31129 , \31130 , \31131 , \31132 , \31133 , \31134 ,
         \31135 , \31136 , \31137 , \31138 , \31139 , \31140_nG90af , \31141 , \31142 , \31143 , \31144 ,
         \31145 , \31146 , \31147 , \31148 , \31149 , \31150 , \31151 , \31152 , \31153 , \31154 ,
         \31155 , \31156 , \31157 , \31158 , \31159_nG90c2 , \31160 , \31161 , \31162 , \31163 , \31164 ,
         \31165 , \31166 , \31167 , \31168 , \31169 , \31170 , \31171 , \31172 , \31173 , \31174 ,
         \31175 , \31176 , \31177 , \31178_nG90d5 , \31179 , \31180 , \31181 , \31182 , \31183 , \31184 ,
         \31185 , \31186 , \31187 , \31188 , \31189 , \31190 , \31191 , \31192 , \31193 , \31194 ,
         \31195 , \31196 , \31197_nG90e8 , \31198 , \31199 , \31200 , \31201 , \31202 , \31203 , \31204 ,
         \31205 , \31206 , \31207 , \31208 , \31209 , \31210 , \31211 , \31212 , \31213 , \31214 ,
         \31215 , \31216_nG90fb , \31217 , \31218 , \31219 , \31220 , \31221 , \31222 , \31223 , \31224 ,
         \31225 , \31226 , \31227 , \31228 , \31229 , \31230 , \31231 , \31232 , \31233 , \31234 ,
         \31235_nG910e , \31236 , \31237 , \31238 , \31239 , \31240 , \31241 , \31242 , \31243 , \31244 ,
         \31245 , \31246 , \31247 , \31248 , \31249 , \31250 , \31251 , \31252 , \31253 , \31254_nG9121 ,
         \31255 , \31256 , \31257 , \31258 , \31259 , \31260 , \31261 , \31262_nG9129 , \31263 , \31264 ,
         \31265 , \31266 , \31267 , \31268 , \31269 , \31270 , \31271 , \31272 , \31273 , \31274 ,
         \31275 , \31276 , \31277 , \31278 , \31279 , \31280 , \31281 , \31282 , \31283 , \31284 ,
         \31285 , \31286 , \31287 , \31288 , \31289 , \31290 , \31291 , \31292 , \31293 , \31294 ,
         \31295 , \31296 , \31297 , \31298 , \31299 , \31300 , \31301 , \31302 , \31303 , \31304 ,
         \31305 , \31306 , \31307 , \31308 , \31309 , \31310 , \31311 , \31312 , \31313 , \31314 ,
         \31315 , \31316 , \31317 , \31318 , \31319 , \31320 , \31321 , \31322 , \31323 , \31324 ,
         \31325 , \31326 , \31327 , \31328 , \31329 , \31330 , \31331 , \31332 , \31333 , \31334 ,
         \31335 , \31336 , \31337 , \31338 , \31339 , \31340 , \31341 , \31342 , \31343 , \31344 ,
         \31345 , \31346 , \31347 , \31348 , \31349 , \31350 , \31351 , \31352 , \31353 , \31354 ,
         \31355 , \31356 , \31357 , \31358 , \31359 , \31360 , \31361 , \31362 , \31363 , \31364 ,
         \31365 , \31366 , \31367 , \31368 , \31369 , \31370 , \31371 , \31372 , \31373 , \31374 ,
         \31375 , \31376 , \31377 , \31378 , \31379 , \31380 , \31381 , \31382 , \31383 , \31384 ,
         \31385 , \31386 , \31387 , \31388 , \31389 , \31390 , \31391 , \31392 , \31393 , \31394 ,
         \31395 , \31396 , \31397 , \31398 , \31399 , \31400 , \31401 , \31402 , \31403 , \31404 ,
         \31405 , \31406 , \31407 , \31408 , \31409 , \31410 , \31411 , \31412 , \31413 , \31414 ,
         \31415 , \31416 , \31417 , \31418 , \31419 , \31420 , \31421 , \31422 , \31423 , \31424 ,
         \31425 , \31426 , \31427 , \31428 , \31429 , \31430 , \31431 , \31432 , \31433 , \31434 ,
         \31435 , \31436 , \31437 , \31438 , \31439 , \31440 , \31441 , \31442 , \31443 , \31444 ,
         \31445 , \31446 , \31447 , \31448 , \31449 , \31450 , \31451 , \31452 , \31453 , \31454 ,
         \31455 , \31456 , \31457 , \31458 , \31459 , \31460 , \31461 , \31462 , \31463 , \31464 ,
         \31465 , \31466 , \31467 , \31468 , \31469 , \31470 , \31471 , \31472 , \31473 , \31474 ,
         \31475 , \31476 , \31477 , \31478 , \31479 , \31480 , \31481 , \31482 , \31483 , \31484 ,
         \31485 , \31486 , \31487 , \31488 , \31489 , \31490 , \31491 , \31492 , \31493 , \31494 ,
         \31495 , \31496 , \31497 , \31498 , \31499 , \31500 , \31501 , \31502 , \31503 , \31504 ,
         \31505 , \31506 , \31507 , \31508 , \31509 , \31510 , \31511 , \31512 , \31513 , \31514 ,
         \31515 , \31516 , \31517 , \31518 , \31519 , \31520 , \31521 , \31522 , \31523 , \31524 ,
         \31525 , \31526 , \31527 , \31528 , \31529 , \31530 , \31531 , \31532 , \31533 , \31534 ,
         \31535 , \31536 , \31537 , \31538 , \31539 , \31540 , \31541 , \31542 , \31543 , \31544 ,
         \31545 , \31546 , \31547 , \31548 , \31549 , \31550 , \31551 , \31552 , \31553 , \31554 ,
         \31555 , \31556 , \31557 , \31558 , \31559 , \31560 , \31561 , \31562 , \31563 , \31564 ,
         \31565 , \31566 , \31567 , \31568 , \31569 , \31570 , \31571 , \31572 , \31573 , \31574 ,
         \31575 , \31576 , \31577 , \31578 , \31579 , \31580 , \31581 , \31582 , \31583 , \31584 ,
         \31585 , \31586 , \31587 , \31588 , \31589 , \31590 , \31591 , \31592 , \31593 , \31594 ,
         \31595 , \31596 , \31597 , \31598 , \31599 , \31600 , \31601 , \31602 , \31603 , \31604 ,
         \31605 , \31606 , \31607 , \31608 , \31609 , \31610 , \31611 , \31612 , \31613 , \31614 ,
         \31615 , \31616 , \31617 , \31618 , \31619 , \31620 , \31621 , \31622 , \31623 , \31624 ,
         \31625 , \31626 , \31627 , \31628 , \31629 , \31630 , \31631 , \31632 , \31633 , \31634 ,
         \31635 , \31636 , \31637 , \31638 , \31639 , \31640 , \31641 , \31642 , \31643 , \31644 ,
         \31645 , \31646 , \31647 , \31648 , \31649 , \31650 , \31651 , \31652 , \31653 , \31654 ,
         \31655 , \31656 , \31657 , \31658 , \31659 , \31660 , \31661 , \31662 , \31663 , \31664 ,
         \31665 , \31666 , \31667 , \31668 , \31669 , \31670 , \31671 , \31672 , \31673 , \31674 ,
         \31675 , \31676 , \31677 , \31678 , \31679 , \31680 , \31681 , \31682 , \31683 , \31684 ,
         \31685 , \31686 , \31687 , \31688 , \31689 , \31690 , \31691 , \31692 , \31693 , \31694 ,
         \31695 , \31696 , \31697 , \31698 , \31699 , \31700 , \31701 , \31702 , \31703 , \31704 ,
         \31705 , \31706 , \31707 , \31708 , \31709 , \31710 , \31711 , \31712 , \31713 , \31714 ,
         \31715 , \31716 , \31717 , \31718 , \31719 , \31720 , \31721 , \31722 , \31723 , \31724 ,
         \31725 , \31726 , \31727 , \31728 , \31729 , \31730 , \31731 , \31732 , \31733 , \31734 ,
         \31735 , \31736 , \31737 , \31738 , \31739 , \31740 , \31741 , \31742 , \31743 , \31744 ,
         \31745 , \31746 , \31747 , \31748 , \31749 , \31750 , \31751 , \31752 , \31753 , \31754 ,
         \31755 , \31756 , \31757 , \31758 , \31759 , \31760 , \31761 , \31762 , \31763 , \31764 ,
         \31765 , \31766 , \31767 , \31768 , \31769 , \31770 , \31771 , \31772 , \31773 , \31774 ,
         \31775 , \31776 , \31777 , \31778 , \31779 , \31780 , \31781 , \31782 , \31783 , \31784 ,
         \31785 , \31786 , \31787 , \31788 , \31789_nG9340 , \31790 , \31791 , \31792 , \31793 , \31794 ,
         \31795 , \31796 , \31797 , \31798 , \31799 , \31800 , \31801 , \31802 , \31803 , \31804 ,
         \31805 , \31806 , \31807 , \31808 , \31809 , \31810 , \31811 , \31812 , \31813 , \31814 ,
         \31815 , \31816 , \31817 , \31818 , \31819 , \31820 , \31821 , \31822 , \31823 , \31824 ,
         \31825 , \31826 , \31827 , \31828 , \31829 , \31830 , \31831 , \31832 , \31833 , \31834 ,
         \31835 , \31836 , \31837 , \31838 , \31839 , \31840 , \31841 , \31842 , \31843 , \31844 ,
         \31845 , \31846 , \31847 , \31848 , \31849 , \31850 , \31851 , \31852 , \31853 , \31854 ,
         \31855 , \31856 , \31857 , \31858 , \31859 , \31860 , \31861 , \31862 , \31863 , \31864 ,
         \31865 , \31866 , \31867 , \31868 , \31869 , \31870 , \31871 , \31872 , \31873 , \31874 ,
         \31875 , \31876 , \31877 , \31878 , \31879 , \31880 , \31881 , \31882 , \31883 , \31884 ,
         \31885 , \31886 , \31887 , \31888 , \31889 , \31890 , \31891 , \31892 , \31893 , \31894 ,
         \31895 , \31896 , \31897 , \31898 , \31899 , \31900 , \31901 , \31902 , \31903 , \31904 ,
         \31905 , \31906 , \31907 , \31908 , \31909 , \31910 , \31911 , \31912 , \31913 , \31914 ,
         \31915 , \31916 , \31917 , \31918 , \31919 , \31920 , \31921 , \31922 , \31923 , \31924 ,
         \31925 , \31926 , \31927 , \31928 , \31929 , \31930 , \31931 , \31932 , \31933 , \31934 ,
         \31935 , \31936 , \31937 , \31938 , \31939 , \31940 , \31941 , \31942 , \31943 , \31944 ,
         \31945 , \31946 , \31947 , \31948 , \31949 , \31950 , \31951 , \31952 , \31953 , \31954 ,
         \31955 , \31956 , \31957 , \31958 , \31959 , \31960 , \31961 , \31962 , \31963 , \31964 ,
         \31965 , \31966 , \31967 , \31968 , \31969 , \31970 , \31971 , \31972 , \31973 , \31974 ,
         \31975 , \31976 , \31977 , \31978 , \31979 , \31980 , \31981 , \31982 , \31983 , \31984 ,
         \31985 , \31986 , \31987 , \31988 , \31989 , \31990 , \31991 , \31992 , \31993 , \31994 ,
         \31995 , \31996 , \31997 , \31998 , \31999 , \32000 , \32001 , \32002 , \32003 , \32004 ,
         \32005 , \32006 , \32007 , \32008 , \32009 , \32010 , \32011 , \32012 , \32013 , \32014 ,
         \32015 , \32016 , \32017 , \32018 , \32019 , \32020 , \32021 , \32022 , \32023 , \32024 ,
         \32025 , \32026 , \32027 , \32028 , \32029 , \32030 , \32031 , \32032 , \32033 , \32034 ,
         \32035 , \32036 , \32037 , \32038 , \32039 , \32040 , \32041 , \32042 , \32043 , \32044 ,
         \32045 , \32046 , \32047 , \32048 , \32049 , \32050 , \32051 , \32052 , \32053 , \32054 ,
         \32055 , \32056 , \32057 , \32058 , \32059 , \32060 , \32061 , \32062 , \32063 , \32064 ,
         \32065 , \32066 , \32067 , \32068 , \32069 , \32070 , \32071 , \32072 , \32073 , \32074 ,
         \32075 , \32076 , \32077 , \32078 , \32079 , \32080 , \32081 , \32082 , \32083 , \32084 ,
         \32085 , \32086 , \32087 , \32088 , \32089 , \32090 , \32091 , \32092 , \32093 , \32094 ,
         \32095 , \32096 , \32097 , \32098 , \32099 , \32100 , \32101 , \32102 , \32103 , \32104 ,
         \32105 , \32106 , \32107 , \32108 , \32109 , \32110 , \32111 , \32112 , \32113 , \32114 ,
         \32115 , \32116 , \32117 , \32118 , \32119 , \32120 , \32121 , \32122 , \32123 , \32124 ,
         \32125 , \32126 , \32127 , \32128 , \32129 , \32130 , \32131 , \32132 , \32133 , \32134 ,
         \32135 , \32136 , \32137 , \32138 , \32139 , \32140 , \32141 , \32142 , \32143 , \32144 ,
         \32145 , \32146 , \32147 , \32148 , \32149 , \32150 , \32151 , \32152 , \32153 , \32154 ,
         \32155 , \32156 , \32157 , \32158 , \32159 , \32160 , \32161 , \32162 , \32163 , \32164 ,
         \32165 , \32166 , \32167 , \32168 , \32169 , \32170 , \32171 , \32172 , \32173 , \32174 ,
         \32175 , \32176 , \32177 , \32178 , \32179 , \32180 , \32181 , \32182 , \32183 , \32184 ,
         \32185 , \32186 , \32187 , \32188 , \32189 , \32190 , \32191 , \32192 , \32193 , \32194 ,
         \32195 , \32196 , \32197 , \32198 , \32199 , \32200 , \32201 , \32202 , \32203 , \32204 ,
         \32205 , \32206 , \32207 , \32208 , \32209 , \32210 , \32211 , \32212 , \32213 , \32214 ,
         \32215 , \32216 , \32217 , \32218 , \32219 , \32220 , \32221 , \32222 , \32223 , \32224 ,
         \32225 , \32226 , \32227 , \32228 , \32229 , \32230 , \32231 , \32232 , \32233 , \32234 ,
         \32235 , \32236 , \32237 , \32238 , \32239 , \32240 , \32241 , \32242 , \32243 , \32244 ,
         \32245 , \32246 , \32247 , \32248 , \32249 , \32250 , \32251 , \32252 , \32253 , \32254 ,
         \32255 , \32256 , \32257 , \32258 , \32259 , \32260 , \32261 , \32262 , \32263 , \32264 ,
         \32265 , \32266 , \32267 , \32268 , \32269 , \32270 , \32271 , \32272 , \32273 , \32274 ,
         \32275 , \32276 , \32277 , \32278 , \32279 , \32280 , \32281 , \32282 , \32283 , \32284 ,
         \32285 , \32286 , \32287 , \32288 , \32289 , \32290 , \32291 , \32292 , \32293 , \32294 ,
         \32295 , \32296 , \32297 , \32298 , \32299 , \32300_nG953f , \32301 , \32302 , \32303 , \32304 ,
         \32305 , \32306 , \32307 , \32308 , \32309 , \32310 , \32311 , \32312 , \32313 , \32314 ,
         \32315 , \32316 , \32317 , \32318 , \32319 , \32320 , \32321_nG9554 , \32322 , \32323 , \32324 ,
         \32325 , \32326 , \32327 , \32328 , \32329 , \32330 , \32331 , \32332 , \32333 , \32334 ,
         \32335 , \32336 , \32337 , \32338 , \32339 , \32340 , \32341 , \32342 , \32343_nG956a , \32344 ,
         \32345 , \32346 , \32347 , \32348 , \32349 , \32350 , \32351 , \32352 , \32353 , \32354 ,
         \32355 , \32356 , \32357 , \32358 , \32359 , \32360 , \32361 , \32362 , \32363 , \32364 ,
         \32365_nG9580 , \32366 , \32367 , \32368 , \32369 , \32370 , \32371 , \32372 , \32373 , \32374 ,
         \32375 , \32376 , \32377 , \32378 , \32379 , \32380 , \32381 , \32382 , \32383 , \32384 ,
         \32385 , \32386 , \32387_nG9596 , \32388 , \32389 , \32390 , \32391 , \32392 , \32393 , \32394 ,
         \32395 , \32396 , \32397 , \32398 , \32399 , \32400 , \32401 , \32402 , \32403 , \32404 ,
         \32405 , \32406 , \32407 , \32408 , \32409_nG95ac , \32410 , \32411 , \32412 , \32413 , \32414 ,
         \32415 , \32416 , \32417 , \32418 , \32419 , \32420 , \32421 , \32422 , \32423 , \32424 ,
         \32425 , \32426 , \32427 , \32428 , \32429 , \32430 , \32431_nG95c2 , \32432 , \32433 , \32434 ,
         \32435 , \32436 , \32437 , \32438 , \32439 , \32440 , \32441 , \32442 , \32443 , \32444 ,
         \32445 , \32446 , \32447 , \32448 , \32449 , \32450 , \32451 , \32452 , \32453_nG95d8 , \32454 ,
         \32455 , \32456 , \32457 , \32458 , \32459 , \32460 , \32461 , \32462 , \32463 , \32464 ,
         \32465 , \32466 , \32467 , \32468 , \32469 , \32470 , \32471 , \32472 , \32473 , \32474 ,
         \32475 , \32476 , \32477 , \32478 , \32479 , \32480 , \32481 , \32482 , \32483 , \32484 ,
         \32485 , \32486 , \32487 , \32488 , \32489 , \32490 , \32491 , \32492 , \32493 , \32494 ,
         \32495 , \32496 , \32497 , \32498 , \32499 , \32500 , \32501 , \32502 , \32503 , \32504 ,
         \32505 , \32506 , \32507 , \32508 , \32509 , \32510 , \32511 , \32512 , \32513 , \32514 ,
         \32515 , \32516 , \32517 , \32518 , \32519 , \32520 , \32521 , \32522 , \32523 , \32524 ,
         \32525 , \32526 , \32527 , \32528 , \32529 , \32530 , \32531 , \32532 , \32533 , \32534 ,
         \32535 , \32536 , \32537 , \32538 , \32539 , \32540 , \32541 , \32542 , \32543 , \32544 ,
         \32545 , \32546 , \32547 , \32548 , \32549 , \32550 , \32551 , \32552 , \32553 , \32554 ,
         \32555 , \32556 , \32557 , \32558 , \32559 , \32560 , \32561 , \32562 , \32563 , \32564 ,
         \32565 , \32566 , \32567 , \32568 , \32569 , \32570 , \32571 , \32572 , \32573 , \32574 ,
         \32575 , \32576 , \32577 , \32578 , \32579 , \32580 , \32581 , \32582 , \32583 , \32584 ,
         \32585 , \32586 , \32587 , \32588 , \32589 , \32590 , \32591 , \32592 , \32593 , \32594 ,
         \32595 , \32596 , \32597 , \32598 , \32599 , \32600 , \32601 , \32602 , \32603 , \32604 ,
         \32605 , \32606 , \32607 , \32608 , \32609 , \32610 , \32611 , \32612 , \32613 , \32614 ,
         \32615 , \32616 , \32617 , \32618 , \32619 , \32620 , \32621 , \32622 , \32623 , \32624 ,
         \32625 , \32626 , \32627 , \32628 , \32629 , \32630 , \32631 , \32632 , \32633 , \32634 ,
         \32635 , \32636 , \32637 , \32638 , \32639 , \32640 , \32641 , \32642 , \32643 , \32644 ,
         \32645 , \32646 , \32647 , \32648 , \32649 , \32650 , \32651 , \32652 , \32653 , \32654 ,
         \32655 , \32656 , \32657 , \32658 , \32659 , \32660 , \32661 , \32662 , \32663 , \32664 ,
         \32665 , \32666 , \32667 , \32668 , \32669 , \32670 , \32671 , \32672 , \32673 , \32674 ,
         \32675 , \32676 , \32677 , \32678 , \32679 , \32680 , \32681 , \32682 , \32683 , \32684 ,
         \32685 , \32686 , \32687 , \32688 , \32689 , \32690 , \32691 , \32692 , \32693 , \32694 ,
         \32695 , \32696 , \32697 , \32698 , \32699 , \32700 , \32701 , \32702 , \32703 , \32704 ,
         \32705 , \32706 , \32707 , \32708 , \32709 , \32710 , \32711 , \32712 , \32713 , \32714 ,
         \32715 , \32716 , \32717 , \32718 , \32719 , \32720 , \32721 , \32722 , \32723 , \32724 ,
         \32725 , \32726 , \32727 , \32728 , \32729 , \32730 , \32731 , \32732 , \32733 , \32734 ,
         \32735 , \32736 , \32737 , \32738 , \32739 , \32740 , \32741 , \32742 , \32743 , \32744 ,
         \32745 , \32746 , \32747 , \32748 , \32749 , \32750 , \32751 , \32752 , \32753 , \32754 ,
         \32755 , \32756 , \32757 , \32758 , \32759 , \32760 , \32761 , \32762 , \32763 , \32764 ,
         \32765 , \32766 , \32767 , \32768 , \32769 , \32770 , \32771 , \32772 , \32773 , \32774 ,
         \32775 , \32776 , \32777 , \32778 , \32779 , \32780 , \32781 , \32782 , \32783 , \32784 ,
         \32785 , \32786 , \32787 , \32788 , \32789 , \32790 , \32791 , \32792 , \32793 , \32794 ,
         \32795 , \32796 , \32797 , \32798 , \32799 , \32800 , \32801 , \32802 , \32803 , \32804 ,
         \32805 , \32806 , \32807 , \32808 , \32809 , \32810 , \32811 , \32812 , \32813 , \32814 ,
         \32815 , \32816 , \32817 , \32818 , \32819 , \32820 , \32821 , \32822 , \32823 , \32824 ,
         \32825 , \32826 , \32827 , \32828 , \32829 , \32830 , \32831 , \32832 , \32833 , \32834 ,
         \32835 , \32836 , \32837 , \32838 , \32839 , \32840 , \32841 , \32842 , \32843 , \32844 ,
         \32845 , \32846 , \32847 , \32848 , \32849 , \32850 , \32851 , \32852 , \32853 , \32854 ,
         \32855 , \32856 , \32857 , \32858 , \32859 , \32860 , \32861 , \32862 , \32863 , \32864 ,
         \32865 , \32866 , \32867 , \32868 , \32869 , \32870 , \32871 , \32872 , \32873 , \32874 ,
         \32875 , \32876 , \32877 , \32878 , \32879 , \32880 , \32881 , \32882 , \32883 , \32884 ,
         \32885 , \32886 , \32887 , \32888 , \32889 , \32890 , \32891 , \32892 , \32893 , \32894 ,
         \32895 , \32896 , \32897 , \32898 , \32899 , \32900 , \32901 , \32902 , \32903 , \32904 ,
         \32905 , \32906 , \32907 , \32908 , \32909 , \32910 , \32911 , \32912 , \32913 , \32914 ,
         \32915 , \32916 , \32917 , \32918 , \32919 , \32920 , \32921 , \32922 , \32923 , \32924 ,
         \32925 , \32926 , \32927 , \32928 , \32929 , \32930 , \32931 , \32932 , \32933 , \32934 ,
         \32935 , \32936 , \32937 , \32938 , \32939 , \32940 , \32941 , \32942 , \32943 , \32944 ,
         \32945 , \32946 , \32947 , \32948 , \32949 , \32950 , \32951 , \32952 , \32953 , \32954 ,
         \32955 , \32956 , \32957 , \32958 , \32959 , \32960 , \32961 , \32962 , \32963 , \32964 ,
         \32965 , \32966 , \32967 , \32968 , \32969_nG97dc , \32970 , \32971 , \32972 , \32973 , \32974 ,
         \32975 , \32976 , \32977 , \32978 , \32979 , \32980 , \32981 , \32982 , \32983 , \32984 ,
         \32985 , \32986 , \32987 , \32988 , \32989 , \32990_nG97f1 , \32991 , \32992 , \32993 , \32994 ,
         \32995 , \32996 , \32997 , \32998 , \32999 , \33000 , \33001 , \33002 , \33003 , \33004 ,
         \33005 , \33006 , \33007 , \33008 , \33009 , \33010 , \33011 , \33012_nG9807 , \33013 , \33014 ,
         \33015 , \33016 , \33017 , \33018 , \33019 , \33020 , \33021 , \33022 , \33023 , \33024 ,
         \33025 , \33026 , \33027 , \33028 , \33029 , \33030 , \33031 , \33032 , \33033 , \33034_nG981d ,
         \33035 , \33036 , \33037 , \33038 , \33039 , \33040 , \33041 , \33042 , \33043 , \33044 ,
         \33045 , \33046 , \33047 , \33048 , \33049 , \33050 , \33051 , \33052 , \33053 , \33054 ,
         \33055 , \33056_nG9833 , \33057 , \33058 , \33059 , \33060 , \33061 , \33062 , \33063 , \33064 ,
         \33065 , \33066 , \33067 , \33068 , \33069 , \33070 , \33071 , \33072 , \33073 , \33074 ,
         \33075 , \33076 , \33077 , \33078_nG9849 , \33079 , \33080 , \33081 , \33082 , \33083 , \33084 ,
         \33085 , \33086 , \33087 , \33088 , \33089 , \33090 , \33091 , \33092 , \33093 , \33094 ,
         \33095 , \33096 , \33097 , \33098 , \33099 , \33100_nG985f , \33101 , \33102 , \33103 , \33104 ,
         \33105 , \33106 , \33107 , \33108 , \33109 , \33110 , \33111 , \33112 , \33113 , \33114 ,
         \33115 , \33116 , \33117 , \33118 , \33119 , \33120 , \33121 , \33122_nG9875 , \33123 , \33124 ,
         \33125 , \33126 , \33127 , \33128 , \33129_nG987c , \33130 , \33131 , \33132 , \33133 , \33134 ,
         \33135 , \33136 , \33137 , \33138 , \33139 , \33140_nG9887 , \33141 , \33142 , \33143 , \33144 ,
         \33145 , \33146 , \33147 , \33148 , \33149 , \33150 , \33151 , \33152 , \33153 , \33154 ,
         \33155 , \33156 , \33157 , \33158 , \33159 , \33160 , \33161 , \33162 , \33163 , \33164 ,
         \33165 , \33166 , \33167 , \33168 , \33169 , \33170 , \33171 , \33172 , \33173 , \33174 ,
         \33175 , \33176 , \33177 , \33178 , \33179 , \33180 , \33181 , \33182 , \33183 , \33184 ,
         \33185 , \33186 , \33187 , \33188 , \33189 , \33190 , \33191 , \33192 , \33193 , \33194 ,
         \33195 , \33196 , \33197 , \33198 , \33199 , \33200 , \33201 , \33202 , \33203 , \33204 ,
         \33205 , \33206_nG98c9 , \33207 , \33208 , \33209 , \33210 , \33211 , \33212 , \33213 , \33214 ,
         \33215 , \33216 , \33217 , \33218 , \33219 , \33220 , \33221 , \33222 , \33223 , \33224_nG98db ,
         \33225 , \33226 , \33227 , \33228 , \33229 , \33230 , \33231 , \33232 , \33233 , \33234 ,
         \33235 , \33236 , \33237 , \33238 , \33239 , \33240 , \33241 , \33242 , \33243_nG98ee , \33244 ,
         \33245 , \33246 , \33247 , \33248 , \33249 , \33250 , \33251 , \33252 , \33253 , \33254 ,
         \33255 , \33256 , \33257 , \33258 , \33259 , \33260 , \33261 , \33262 , \33263_nG9902 , \33264 ,
         \33265 , \33266 , \33267 , \33268 , \33269 , \33270 , \33271 , \33272 , \33273 , \33274 ,
         \33275 , \33276 , \33277 , \33278 , \33279 , \33280 , \33281 , \33282 , \33283_nG9916 , \33284 ,
         \33285 , \33286 , \33287 , \33288 , \33289 , \33290 , \33291 , \33292 , \33293 , \33294 ,
         \33295 , \33296 , \33297 , \33298 , \33299 , \33300 , \33301 , \33302 , \33303_nG992a , \33304 ,
         \33305 , \33306 , \33307 , \33308 , \33309 , \33310 , \33311 , \33312 , \33313 , \33314 ,
         \33315 , \33316 , \33317 , \33318 , \33319 , \33320 , \33321 , \33322 , \33323_nG993e , \33324 ,
         \33325 , \33326 , \33327 , \33328 , \33329 , \33330 , \33331 , \33332 , \33333 , \33334 ,
         \33335 , \33336 , \33337 , \33338 , \33339 , \33340 , \33341 , \33342 , \33343_nG9952 , \33344 ,
         \33345 , \33346 , \33347 , \33348 , \33349 , \33350 , \33351 , \33352 , \33353 , \33354 ,
         \33355 , \33356 , \33357 , \33358 , \33359 , \33360 , \33361 , \33362 , \33363_nG9966 , \33364 ,
         \33365 , \33366 , \33367 , \33368 , \33369 , \33370 , \33371 , \33372 , \33373 , \33374 ,
         \33375 , \33376 , \33377 , \33378 , \33379 , \33380 , \33381 , \33382 , \33383 , \33384 ,
         \33385_nG997c , \33386 , \33387 , \33388 , \33389 , \33390 , \33391 , \33392 , \33393 , \33394 ,
         \33395 , \33396 , \33397 , \33398 , \33399 , \33400 , \33401 , \33402 , \33403 , \33404_nG998f ,
         \33405 , \33406 , \33407 , \33408 , \33409 , \33410 , \33411 , \33412 , \33413 , \33414 ,
         \33415 , \33416 , \33417 , \33418 , \33419 , \33420 , \33421 , \33422 , \33423 , \33424_nG99a3 ,
         \33425 , \33426 , \33427 , \33428 , \33429 , \33430 , \33431 , \33432 , \33433 , \33434 ,
         \33435 , \33436 , \33437 , \33438 , \33439 , \33440 , \33441 , \33442 , \33443 , \33444_nG99b7 ,
         \33445 , \33446 , \33447 , \33448 , \33449 , \33450 , \33451 , \33452 , \33453 , \33454 ,
         \33455 , \33456 , \33457 , \33458 , \33459 , \33460 , \33461 , \33462 , \33463 , \33464_nG99cb ,
         \33465 , \33466 , \33467 , \33468 , \33469 , \33470 , \33471 , \33472 , \33473 , \33474 ,
         \33475 , \33476 , \33477 , \33478 , \33479 , \33480 , \33481 , \33482 , \33483 , \33484_nG99df ,
         \33485 , \33486 , \33487 , \33488 , \33489 , \33490 , \33491 , \33492 , \33493 , \33494 ,
         \33495 , \33496 , \33497 , \33498 , \33499 , \33500 , \33501 , \33502 , \33503 , \33504_nG99f3 ,
         \33505 , \33506 , \33507 , \33508 , \33509 , \33510 , \33511 , \33512 , \33513 , \33514 ,
         \33515 , \33516 , \33517 , \33518 , \33519 , \33520 , \33521 , \33522 , \33523 , \33524_nG9a07 ,
         \33525 , \33526 , \33527 , \33528 , \33529 , \33530 , \33531 , \33532_nG9a0f , \33533 , \33534 ,
         \33535 , \33536 , \33537 , \33538 , \33539 , \33540 , \33541 , \33542 , \33543 , \33544 ,
         \33545 , \33546 , \33547 , \33548 , \33549 , \33550 , \33551 , \33552 , \33553 , \33554 ,
         \33555 , \33556 , \33557 , \33558 , \33559 , \33560 , \33561 , \33562 , \33563 , \33564 ,
         \33565 , \33566 , \33567 , \33568 , \33569 , \33570 , \33571 , \33572 , \33573 , \33574 ,
         \33575 , \33576 , \33577 , \33578 , \33579 , \33580 , \33581 , \33582 , \33583 , \33584 ,
         \33585 , \33586 , \33587 , \33588 , \33589 , \33590 , \33591 , \33592 , \33593 , \33594 ,
         \33595 , \33596 , \33597 , \33598 , \33599 , \33600 , \33601 , \33602 , \33603 , \33604 ,
         \33605 , \33606 , \33607 , \33608 , \33609 , \33610 , \33611 , \33612 , \33613 , \33614 ,
         \33615 , \33616 , \33617 , \33618 , \33619 , \33620 , \33621 , \33622 , \33623 , \33624 ,
         \33625 , \33626 , \33627 , \33628 , \33629 , \33630 , \33631 , \33632 , \33633 , \33634 ,
         \33635 , \33636 , \33637 , \33638 , \33639 , \33640 , \33641 , \33642 , \33643 , \33644 ,
         \33645 , \33646 , \33647 , \33648 , \33649 , \33650 , \33651 , \33652 , \33653 , \33654 ,
         \33655 , \33656 , \33657 , \33658 , \33659 , \33660 , \33661 , \33662 , \33663 , \33664 ,
         \33665 , \33666 , \33667 , \33668 , \33669 , \33670 , \33671 , \33672 , \33673 , \33674 ,
         \33675 , \33676 , \33677 , \33678 , \33679 , \33680 , \33681 , \33682 , \33683 , \33684 ,
         \33685 , \33686 , \33687 , \33688 , \33689 , \33690 , \33691 , \33692 , \33693 , \33694 ,
         \33695 , \33696 , \33697 , \33698 , \33699 , \33700 , \33701 , \33702 , \33703 , \33704 ,
         \33705 , \33706 , \33707 , \33708 , \33709 , \33710 , \33711 , \33712 , \33713 , \33714 ,
         \33715 , \33716 , \33717 , \33718 , \33719 , \33720 , \33721 , \33722 , \33723 , \33724 ,
         \33725 , \33726 , \33727 , \33728 , \33729 , \33730 , \33731 , \33732 , \33733 , \33734 ,
         \33735 , \33736 , \33737 , \33738 , \33739 , \33740 , \33741 , \33742 , \33743 , \33744 ,
         \33745 , \33746 , \33747 , \33748 , \33749 , \33750 , \33751 , \33752 , \33753 , \33754 ,
         \33755 , \33756 , \33757 , \33758 , \33759 , \33760 , \33761 , \33762 , \33763 , \33764 ,
         \33765 , \33766 , \33767 , \33768 , \33769 , \33770 , \33771 , \33772 , \33773 , \33774 ,
         \33775 , \33776 , \33777 , \33778 , \33779 , \33780 , \33781 , \33782 , \33783 , \33784 ,
         \33785 , \33786 , \33787 , \33788 , \33789 , \33790 , \33791 , \33792 , \33793 , \33794 ,
         \33795 , \33796 , \33797 , \33798 , \33799 , \33800 , \33801 , \33802 , \33803 , \33804 ,
         \33805 , \33806 , \33807 , \33808 , \33809 , \33810 , \33811 , \33812 , \33813 , \33814 ,
         \33815 , \33816 , \33817 , \33818 , \33819 , \33820 , \33821 , \33822 , \33823 , \33824 ,
         \33825 , \33826 , \33827 , \33828 , \33829 , \33830 , \33831 , \33832 , \33833 , \33834 ,
         \33835 , \33836 , \33837 , \33838 , \33839 , \33840 , \33841 , \33842 , \33843 , \33844 ,
         \33845 , \33846 , \33847 , \33848 , \33849 , \33850 , \33851 , \33852 , \33853 , \33854 ,
         \33855 , \33856 , \33857 , \33858 , \33859 , \33860 , \33861 , \33862 , \33863 , \33864 ,
         \33865 , \33866 , \33867 , \33868 , \33869 , \33870 , \33871 , \33872 , \33873 , \33874 ,
         \33875 , \33876 , \33877 , \33878 , \33879 , \33880 , \33881 , \33882 , \33883 , \33884 ,
         \33885 , \33886 , \33887 , \33888 , \33889 , \33890 , \33891 , \33892 , \33893 , \33894 ,
         \33895 , \33896 , \33897 , \33898 , \33899 , \33900 , \33901 , \33902 , \33903 , \33904 ,
         \33905 , \33906 , \33907 , \33908 , \33909 , \33910 , \33911 , \33912 , \33913 , \33914 ,
         \33915 , \33916 , \33917 , \33918 , \33919 , \33920 , \33921 , \33922 , \33923 , \33924 ,
         \33925 , \33926 , \33927 , \33928 , \33929 , \33930 , \33931 , \33932 , \33933 , \33934 ,
         \33935 , \33936 , \33937 , \33938 , \33939 , \33940 , \33941 , \33942 , \33943 , \33944 ,
         \33945 , \33946 , \33947 , \33948 , \33949 , \33950 , \33951 , \33952 , \33953 , \33954 ,
         \33955 , \33956 , \33957 , \33958 , \33959 , \33960 , \33961 , \33962 , \33963 , \33964 ,
         \33965 , \33966 , \33967 , \33968 , \33969 , \33970 , \33971 , \33972 , \33973 , \33974 ,
         \33975 , \33976 , \33977 , \33978 , \33979 , \33980 , \33981 , \33982 , \33983 , \33984 ,
         \33985 , \33986 , \33987 , \33988 , \33989 , \33990 , \33991 , \33992 , \33993 , \33994 ,
         \33995 , \33996 , \33997 , \33998 , \33999 , \34000 , \34001 , \34002 , \34003 , \34004 ,
         \34005 , \34006 , \34007 , \34008 , \34009 , \34010 , \34011 , \34012 , \34013 , \34014 ,
         \34015 , \34016 , \34017 , \34018 , \34019 , \34020 , \34021 , \34022 , \34023 , \34024 ,
         \34025 , \34026 , \34027 , \34028 , \34029 , \34030 , \34031 , \34032 , \34033 , \34034 ,
         \34035 , \34036 , \34037 , \34038 , \34039 , \34040 , \34041 , \34042 , \34043 , \34044 ,
         \34045 , \34046 , \34047 , \34048 , \34049 , \34050 , \34051 , \34052 , \34053 , \34054 ,
         \34055 , \34056 , \34057 , \34058 , \34059_nG9c26 , \34060 , \34061 , \34062 , \34063 , \34064 ,
         \34065 , \34066 , \34067 , \34068 , \34069 , \34070 , \34071 , \34072 , \34073 , \34074 ,
         \34075 , \34076 , \34077 , \34078 , \34079 , \34080 , \34081 , \34082 , \34083 , \34084 ,
         \34085 , \34086 , \34087 , \34088 , \34089 , \34090 , \34091 , \34092 , \34093 , \34094 ,
         \34095 , \34096 , \34097 , \34098 , \34099 , \34100 , \34101 , \34102 , \34103 , \34104 ,
         \34105 , \34106 , \34107 , \34108 , \34109 , \34110 , \34111 , \34112 , \34113 , \34114 ,
         \34115 , \34116 , \34117 , \34118 , \34119 , \34120 , \34121 , \34122 , \34123 , \34124 ,
         \34125 , \34126 , \34127 , \34128 , \34129 , \34130 , \34131 , \34132 , \34133 , \34134 ,
         \34135 , \34136 , \34137 , \34138 , \34139 , \34140 , \34141 , \34142 , \34143 , \34144 ,
         \34145 , \34146 , \34147 , \34148 , \34149 , \34150 , \34151 , \34152 , \34153 , \34154 ,
         \34155 , \34156 , \34157 , \34158 , \34159 , \34160 , \34161 , \34162 , \34163 , \34164 ,
         \34165 , \34166 , \34167 , \34168 , \34169 , \34170 , \34171 , \34172 , \34173 , \34174 ,
         \34175 , \34176 , \34177 , \34178 , \34179 , \34180 , \34181 , \34182 , \34183 , \34184 ,
         \34185 , \34186 , \34187 , \34188 , \34189 , \34190 , \34191 , \34192 , \34193 , \34194 ,
         \34195 , \34196 , \34197 , \34198 , \34199 , \34200 , \34201 , \34202 , \34203 , \34204 ,
         \34205 , \34206 , \34207 , \34208 , \34209 , \34210 , \34211 , \34212 , \34213 , \34214 ,
         \34215 , \34216 , \34217 , \34218 , \34219 , \34220 , \34221 , \34222 , \34223 , \34224 ,
         \34225 , \34226 , \34227 , \34228 , \34229 , \34230 , \34231 , \34232 , \34233 , \34234 ,
         \34235 , \34236 , \34237 , \34238 , \34239 , \34240 , \34241 , \34242 , \34243 , \34244 ,
         \34245 , \34246 , \34247 , \34248 , \34249 , \34250 , \34251 , \34252 , \34253 , \34254 ,
         \34255 , \34256 , \34257 , \34258 , \34259 , \34260 , \34261 , \34262 , \34263 , \34264 ,
         \34265 , \34266 , \34267 , \34268 , \34269 , \34270 , \34271 , \34272 , \34273 , \34274 ,
         \34275 , \34276 , \34277 , \34278 , \34279 , \34280 , \34281 , \34282 , \34283 , \34284 ,
         \34285 , \34286 , \34287 , \34288 , \34289 , \34290 , \34291 , \34292 , \34293 , \34294 ,
         \34295 , \34296 , \34297 , \34298 , \34299 , \34300 , \34301 , \34302 , \34303 , \34304 ,
         \34305 , \34306 , \34307 , \34308 , \34309 , \34310 , \34311 , \34312 , \34313 , \34314 ,
         \34315 , \34316 , \34317 , \34318 , \34319 , \34320 , \34321 , \34322 , \34323 , \34324 ,
         \34325 , \34326 , \34327 , \34328 , \34329 , \34330 , \34331 , \34332 , \34333 , \34334 ,
         \34335 , \34336 , \34337 , \34338 , \34339 , \34340 , \34341 , \34342 , \34343 , \34344 ,
         \34345 , \34346 , \34347 , \34348 , \34349 , \34350 , \34351 , \34352 , \34353 , \34354 ,
         \34355 , \34356 , \34357 , \34358 , \34359 , \34360 , \34361 , \34362 , \34363 , \34364 ,
         \34365 , \34366 , \34367 , \34368 , \34369 , \34370 , \34371 , \34372 , \34373 , \34374 ,
         \34375 , \34376 , \34377 , \34378 , \34379 , \34380 , \34381 , \34382 , \34383 , \34384 ,
         \34385 , \34386 , \34387 , \34388 , \34389 , \34390 , \34391 , \34392 , \34393 , \34394 ,
         \34395 , \34396 , \34397 , \34398 , \34399 , \34400 , \34401 , \34402 , \34403 , \34404 ,
         \34405 , \34406 , \34407 , \34408 , \34409 , \34410 , \34411 , \34412 , \34413 , \34414 ,
         \34415 , \34416 , \34417 , \34418 , \34419 , \34420 , \34421 , \34422 , \34423 , \34424 ,
         \34425 , \34426 , \34427 , \34428 , \34429 , \34430 , \34431 , \34432 , \34433 , \34434 ,
         \34435 , \34436 , \34437 , \34438 , \34439 , \34440 , \34441 , \34442 , \34443 , \34444 ,
         \34445 , \34446 , \34447 , \34448 , \34449 , \34450 , \34451 , \34452 , \34453 , \34454 ,
         \34455 , \34456 , \34457 , \34458 , \34459 , \34460 , \34461 , \34462 , \34463 , \34464 ,
         \34465 , \34466 , \34467 , \34468 , \34469 , \34470 , \34471 , \34472 , \34473 , \34474 ,
         \34475 , \34476 , \34477 , \34478 , \34479 , \34480 , \34481 , \34482 , \34483 , \34484 ,
         \34485 , \34486 , \34487 , \34488 , \34489 , \34490 , \34491 , \34492 , \34493 , \34494 ,
         \34495 , \34496 , \34497 , \34498 , \34499 , \34500 , \34501 , \34502 , \34503 , \34504 ,
         \34505 , \34506 , \34507 , \34508 , \34509 , \34510 , \34511 , \34512 , \34513 , \34514 ,
         \34515 , \34516 , \34517 , \34518 , \34519 , \34520 , \34521 , \34522 , \34523 , \34524 ,
         \34525 , \34526 , \34527 , \34528 , \34529 , \34530 , \34531 , \34532 , \34533 , \34534 ,
         \34535 , \34536 , \34537 , \34538 , \34539 , \34540 , \34541 , \34542 , \34543 , \34544 ,
         \34545 , \34546 , \34547 , \34548 , \34549 , \34550 , \34551 , \34552 , \34553 , \34554 ,
         \34555 , \34556 , \34557 , \34558 , \34559 , \34560 , \34561 , \34562 , \34563 , \34564 ,
         \34565 , \34566 , \34567 , \34568 , \34569 , \34570_nG9e25 , \34571 , \34572 , \34573 , \34574 ,
         \34575 , \34576 , \34577 , \34578 , \34579 , \34580 , \34581 , \34582 , \34583 , \34584 ,
         \34585 , \34586 , \34587 , \34588 , \34589 , \34590 , \34591_nG9e3a , \34592 , \34593 , \34594 ,
         \34595 , \34596 , \34597 , \34598 , \34599 , \34600 , \34601 , \34602 , \34603 , \34604 ,
         \34605 , \34606 , \34607 , \34608 , \34609 , \34610 , \34611 , \34612 , \34613_nG9e50 , \34614 ,
         \34615 , \34616 , \34617 , \34618 , \34619 , \34620 , \34621 , \34622 , \34623 , \34624 ,
         \34625 , \34626 , \34627 , \34628 , \34629 , \34630 , \34631 , \34632 , \34633 , \34634 ,
         \34635_nG9e66 , \34636 , \34637 , \34638 , \34639 , \34640 , \34641 , \34642 , \34643 , \34644 ,
         \34645 , \34646 , \34647 , \34648 , \34649 , \34650 , \34651 , \34652 , \34653 , \34654 ,
         \34655 , \34656 , \34657_nG9e7c , \34658 , \34659 , \34660 , \34661 , \34662 , \34663 , \34664 ,
         \34665 , \34666 , \34667 , \34668 , \34669 , \34670 , \34671 , \34672 , \34673 , \34674 ,
         \34675 , \34676 , \34677 , \34678 , \34679_nG9e92 , \34680 , \34681 , \34682 , \34683 , \34684 ,
         \34685 , \34686 , \34687 , \34688 , \34689 , \34690 , \34691 , \34692 , \34693 , \34694 ,
         \34695 , \34696 , \34697 , \34698 , \34699 , \34700 , \34701_nG9ea8 , \34702 , \34703 , \34704 ,
         \34705 , \34706 , \34707 , \34708 , \34709 , \34710 , \34711 , \34712 , \34713 , \34714 ,
         \34715 , \34716 , \34717 , \34718 , \34719 , \34720 , \34721 , \34722 , \34723_nG9ebe , \34724 ,
         \34725 , \34726 , \34727 , \34728 , \34729 , \34730 , \34731 , \34732 , \34733 , \34734 ,
         \34735 , \34736 , \34737 , \34738 , \34739 , \34740 , \34741 , \34742 , \34743 , \34744 ,
         \34745 , \34746 , \34747 , \34748 , \34749 , \34750 , \34751 , \34752 , \34753 , \34754 ,
         \34755 , \34756 , \34757 , \34758 , \34759 , \34760 , \34761 , \34762 , \34763 , \34764 ,
         \34765 , \34766 , \34767 , \34768 , \34769 , \34770 , \34771 , \34772 , \34773 , \34774 ,
         \34775 , \34776 , \34777 , \34778 , \34779 , \34780 , \34781 , \34782 , \34783 , \34784 ,
         \34785 , \34786 , \34787 , \34788 , \34789 , \34790 , \34791 , \34792 , \34793 , \34794 ,
         \34795 , \34796 , \34797 , \34798 , \34799 , \34800 , \34801 , \34802 , \34803 , \34804 ,
         \34805 , \34806 , \34807 , \34808 , \34809 , \34810 , \34811 , \34812 , \34813 , \34814 ,
         \34815 , \34816 , \34817 , \34818 , \34819 , \34820 , \34821 , \34822 , \34823 , \34824 ,
         \34825 , \34826 , \34827 , \34828 , \34829 , \34830 , \34831 , \34832 , \34833 , \34834 ,
         \34835 , \34836 , \34837 , \34838 , \34839 , \34840 , \34841 , \34842 , \34843 , \34844 ,
         \34845 , \34846 , \34847 , \34848 , \34849 , \34850 , \34851 , \34852 , \34853 , \34854 ,
         \34855 , \34856 , \34857 , \34858 , \34859 , \34860 , \34861 , \34862 , \34863 , \34864 ,
         \34865 , \34866 , \34867 , \34868 , \34869 , \34870 , \34871 , \34872 , \34873 , \34874 ,
         \34875 , \34876 , \34877 , \34878 , \34879 , \34880 , \34881 , \34882 , \34883 , \34884 ,
         \34885 , \34886 , \34887 , \34888 , \34889 , \34890 , \34891 , \34892 , \34893 , \34894 ,
         \34895 , \34896 , \34897 , \34898 , \34899 , \34900 , \34901 , \34902 , \34903 , \34904 ,
         \34905 , \34906 , \34907 , \34908 , \34909 , \34910 , \34911 , \34912 , \34913 , \34914 ,
         \34915 , \34916 , \34917 , \34918 , \34919 , \34920 , \34921 , \34922 , \34923 , \34924 ,
         \34925 , \34926 , \34927 , \34928 , \34929 , \34930 , \34931 , \34932 , \34933 , \34934 ,
         \34935 , \34936 , \34937 , \34938 , \34939 , \34940 , \34941 , \34942 , \34943 , \34944 ,
         \34945 , \34946 , \34947 , \34948 , \34949 , \34950 , \34951 , \34952 , \34953 , \34954 ,
         \34955 , \34956 , \34957 , \34958 , \34959 , \34960 , \34961 , \34962 , \34963 , \34964 ,
         \34965 , \34966 , \34967 , \34968 , \34969 , \34970 , \34971 , \34972 , \34973 , \34974 ,
         \34975 , \34976 , \34977 , \34978 , \34979 , \34980 , \34981 , \34982 , \34983 , \34984 ,
         \34985 , \34986 , \34987 , \34988 , \34989 , \34990 , \34991 , \34992 , \34993 , \34994 ,
         \34995 , \34996 , \34997 , \34998 , \34999 , \35000 , \35001 , \35002 , \35003 , \35004 ,
         \35005 , \35006 , \35007 , \35008 , \35009 , \35010 , \35011 , \35012 , \35013 , \35014 ,
         \35015 , \35016 , \35017 , \35018 , \35019 , \35020 , \35021 , \35022 , \35023 , \35024 ,
         \35025 , \35026 , \35027 , \35028 , \35029 , \35030 , \35031 , \35032 , \35033 , \35034 ,
         \35035 , \35036 , \35037 , \35038 , \35039 , \35040 , \35041 , \35042 , \35043 , \35044 ,
         \35045 , \35046 , \35047 , \35048 , \35049 , \35050 , \35051 , \35052 , \35053 , \35054 ,
         \35055 , \35056 , \35057 , \35058 , \35059 , \35060 , \35061 , \35062 , \35063 , \35064 ,
         \35065 , \35066 , \35067 , \35068 , \35069 , \35070 , \35071 , \35072 , \35073 , \35074 ,
         \35075 , \35076 , \35077 , \35078 , \35079 , \35080 , \35081 , \35082 , \35083 , \35084 ,
         \35085 , \35086 , \35087 , \35088 , \35089 , \35090 , \35091 , \35092 , \35093 , \35094 ,
         \35095 , \35096 , \35097 , \35098 , \35099 , \35100 , \35101 , \35102 , \35103 , \35104 ,
         \35105 , \35106 , \35107 , \35108 , \35109 , \35110 , \35111 , \35112 , \35113 , \35114 ,
         \35115 , \35116 , \35117 , \35118 , \35119 , \35120 , \35121 , \35122 , \35123 , \35124 ,
         \35125 , \35126 , \35127 , \35128 , \35129 , \35130 , \35131 , \35132 , \35133 , \35134 ,
         \35135 , \35136 , \35137 , \35138 , \35139 , \35140 , \35141 , \35142 , \35143 , \35144 ,
         \35145 , \35146 , \35147 , \35148 , \35149 , \35150 , \35151 , \35152 , \35153 , \35154 ,
         \35155 , \35156 , \35157 , \35158 , \35159 , \35160 , \35161 , \35162 , \35163 , \35164 ,
         \35165 , \35166 , \35167 , \35168 , \35169 , \35170 , \35171 , \35172 , \35173 , \35174 ,
         \35175 , \35176 , \35177 , \35178 , \35179 , \35180 , \35181 , \35182 , \35183 , \35184 ,
         \35185 , \35186 , \35187 , \35188 , \35189 , \35190 , \35191 , \35192 , \35193 , \35194 ,
         \35195 , \35196 , \35197 , \35198 , \35199 , \35200 , \35201 , \35202 , \35203 , \35204 ,
         \35205 , \35206 , \35207 , \35208 , \35209 , \35210 , \35211 , \35212 , \35213 , \35214 ,
         \35215 , \35216 , \35217 , \35218 , \35219 , \35220 , \35221 , \35222 , \35223 , \35224 ,
         \35225 , \35226 , \35227 , \35228 , \35229 , \35230 , \35231 , \35232 , \35233 , \35234 ,
         \35235 , \35236 , \35237 , \35238 , \35239_nGa0c2 , \35240 , \35241 , \35242 , \35243 , \35244 ,
         \35245 , \35246 , \35247 , \35248 , \35249 , \35250 , \35251 , \35252 , \35253 , \35254 ,
         \35255 , \35256 , \35257 , \35258 , \35259 , \35260_nGa0d7 , \35261 , \35262 , \35263 , \35264 ,
         \35265 , \35266 , \35267 , \35268 , \35269 , \35270 , \35271 , \35272 , \35273 , \35274 ,
         \35275 , \35276 , \35277 , \35278 , \35279 , \35280 , \35281 , \35282_nGa0ed , \35283 , \35284 ,
         \35285 , \35286 , \35287 , \35288 , \35289 , \35290 , \35291 , \35292 , \35293 , \35294 ,
         \35295 , \35296 , \35297 , \35298 , \35299 , \35300 , \35301 , \35302 , \35303 , \35304_nGa103 ,
         \35305 , \35306 , \35307 , \35308 , \35309 , \35310 , \35311 , \35312 , \35313 , \35314 ,
         \35315 , \35316 , \35317 , \35318 , \35319 , \35320 , \35321 , \35322 , \35323 , \35324 ,
         \35325 , \35326_nGa119 , \35327 , \35328 , \35329 , \35330 , \35331 , \35332 , \35333 , \35334 ,
         \35335 , \35336 , \35337 , \35338 , \35339 , \35340 , \35341 , \35342 , \35343 , \35344 ,
         \35345 , \35346 , \35347 , \35348_nGa12f , \35349 , \35350 , \35351 , \35352 , \35353 , \35354 ,
         \35355 , \35356 , \35357 , \35358 , \35359 , \35360 , \35361 , \35362 , \35363 , \35364 ,
         \35365 , \35366 , \35367 , \35368 , \35369 , \35370_nGa145 , \35371 , \35372 , \35373 , \35374 ,
         \35375 , \35376 , \35377 , \35378 , \35379 , \35380 , \35381 , \35382 , \35383 , \35384 ,
         \35385 , \35386 , \35387 , \35388 , \35389 , \35390 , \35391 , \35392_nGa15b , \35393 , \35394 ,
         \35395 , \35396 , \35397 , \35398 , \35399_nGa162 , \35400 , \35401 , \35402 , \35403 , \35404 ,
         \35405 , \35406 , \35407 , \35408 , \35409 , \35410_nGa16d , \35411 , \35412 , \35413 , \35414 ,
         \35415 , \35416 , \35417 , \35418 , \35419 , \35420 , \35421 , \35422 , \35423 , \35424 ,
         \35425 , \35426 , \35427 , \35428 , \35429 , \35430 , \35431 , \35432 , \35433 , \35434 ,
         \35435 , \35436 , \35437 , \35438 , \35439 , \35440 , \35441 , \35442 , \35443 , \35444 ,
         \35445 , \35446 , \35447 , \35448 , \35449 , \35450 , \35451 , \35452 , \35453 , \35454 ,
         \35455 , \35456 , \35457 , \35458 , \35459 , \35460 , \35461 , \35462 , \35463 , \35464 ,
         \35465 , \35466 , \35467 , \35468 , \35469 , \35470 , \35471 , \35472 , \35473 , \35474 ,
         \35475 , \35476_nGa1b0 , \35477 , \35478 , \35479 , \35480 , \35481 , \35482 , \35483 , \35484 ,
         \35485 , \35486 , \35487 , \35488 , \35489 , \35490 , \35491 , \35492 , \35493 , \35494 ,
         \35495_nGa1c3 , \35496 , \35497 , \35498 , \35499 , \35500 , \35501 , \35502 , \35503 , \35504 ,
         \35505 , \35506 , \35507 , \35508 , \35509 , \35510 , \35511 , \35512 , \35513 , \35514 ,
         \35515_nGa1d7 , \35516 , \35517 , \35518 , \35519 , \35520 , \35521 , \35522 , \35523 , \35524 ,
         \35525 , \35526 , \35527 , \35528 , \35529 , \35530 , \35531 , \35532 , \35533 , \35534 ,
         \35535 , \35536_nGa1ec , \35537 , \35538 , \35539 , \35540 , \35541 , \35542 , \35543 , \35544 ,
         \35545 , \35546 , \35547 , \35548 , \35549 , \35550 , \35551 , \35552 , \35553 , \35554 ,
         \35555 , \35556 , \35557_nGa201 , \35558 , \35559 , \35560 , \35561 , \35562 , \35563 , \35564 ,
         \35565 , \35566 , \35567 , \35568 , \35569 , \35570 , \35571 , \35572 , \35573 , \35574 ,
         \35575 , \35576 , \35577 , \35578_nGa216 , \35579 , \35580 , \35581 , \35582 , \35583 , \35584 ,
         \35585 , \35586 , \35587 , \35588 , \35589 , \35590 , \35591 , \35592 , \35593 , \35594 ,
         \35595 , \35596 , \35597 , \35598 , \35599_nGa22b , \35600 , \35601 , \35602 , \35603 , \35604 ,
         \35605 , \35606 , \35607 , \35608 , \35609 , \35610 , \35611 , \35612 , \35613 , \35614 ,
         \35615 , \35616 , \35617 , \35618 , \35619 , \35620_nGa240 , \35621 , \35622 , \35623 , \35624 ,
         \35625 , \35626 , \35627 , \35628 , \35629 , \35630 , \35631 , \35632 , \35633 , \35634 ,
         \35635 , \35636 , \35637 , \35638 , \35639 , \35640 , \35641_nGa255 , \35642 , \35643 , \35644 ,
         \35645 , \35646 , \35647 , \35648 , \35649 , \35650 , \35651 , \35652 , \35653 , \35654 ,
         \35655 , \35656 , \35657 , \35658 , \35659 , \35660 , \35661 , \35662 , \35663 , \35664_nGa26c ,
         \35665 , \35666 , \35667 , \35668 , \35669 , \35670 , \35671 , \35672 , \35673 , \35674 ,
         \35675 , \35676 , \35677 , \35678 , \35679 , \35680 , \35681 , \35682 , \35683 , \35684_nGa280 ,
         \35685 , \35686 , \35687 , \35688 , \35689 , \35690 , \35691 , \35692 , \35693 , \35694 ,
         \35695 , \35696 , \35697 , \35698 , \35699 , \35700 , \35701 , \35702 , \35703 , \35704 ,
         \35705_nGa295 , \35706 , \35707 , \35708 , \35709 , \35710 , \35711 , \35712 , \35713 , \35714 ,
         \35715 , \35716 , \35717 , \35718 , \35719 , \35720 , \35721 , \35722 , \35723 , \35724 ,
         \35725 , \35726_nGa2aa , \35727 , \35728 , \35729 , \35730 , \35731 , \35732 , \35733 , \35734 ,
         \35735 , \35736 , \35737 , \35738 , \35739 , \35740 , \35741 , \35742 , \35743 , \35744 ,
         \35745 , \35746 , \35747_nGa2bf , \35748 , \35749 , \35750 , \35751 , \35752 , \35753 , \35754 ,
         \35755 , \35756 , \35757 , \35758 , \35759 , \35760 , \35761 , \35762 , \35763 , \35764 ,
         \35765 , \35766 , \35767 , \35768_nGa2d4 , \35769 , \35770 , \35771 , \35772 , \35773 , \35774 ,
         \35775 , \35776 , \35777 , \35778 , \35779 , \35780 , \35781 , \35782 , \35783 , \35784 ,
         \35785 , \35786 , \35787 , \35788 , \35789_nGa2e9 , \35790 , \35791 , \35792 , \35793 , \35794 ,
         \35795 , \35796 , \35797 , \35798 , \35799 , \35800 , \35801 , \35802 , \35803 , \35804 ,
         \35805 , \35806 , \35807 , \35808 , \35809 , \35810_nGa2fe , \35811 , \35812 , \35813 , \35814 ,
         \35815 , \35816 , \35817 , \35818_nGa306 , \35819 , \35820 , \35821 , \35822 , \35823 , \35824 ,
         \35825 , \35826 , \35827 , \35828 , \35829 , \35830 , \35831 , \35832 , \35833 , \35834 ,
         \35835 , \35836 , \35837 , \35838 , \35839 , \35840 , \35841 , \35842 , \35843 , \35844 ,
         \35845 , \35846 , \35847 , \35848 , \35849 , \35850 , \35851 , \35852 , \35853 , \35854 ,
         \35855 , \35856 , \35857 , \35858 , \35859 , \35860 , \35861 , \35862 , \35863 , \35864 ,
         \35865 , \35866 , \35867 , \35868 , \35869 , \35870 , \35871 , \35872 , \35873 , \35874 ,
         \35875 , \35876 , \35877 , \35878 , \35879 , \35880 , \35881 , \35882 , \35883 , \35884 ,
         \35885 , \35886 , \35887 , \35888 , \35889 , \35890 , \35891 , \35892 , \35893 , \35894 ,
         \35895 , \35896 , \35897 , \35898 , \35899 , \35900 , \35901 , \35902 , \35903 , \35904 ,
         \35905 , \35906 , \35907 , \35908 , \35909 , \35910 , \35911 , \35912 , \35913 , \35914 ,
         \35915 , \35916 , \35917 , \35918 , \35919 , \35920 , \35921 , \35922 , \35923 , \35924 ,
         \35925 , \35926 , \35927 , \35928 , \35929 , \35930 , \35931 , \35932 , \35933 , \35934 ,
         \35935 , \35936 , \35937 , \35938 , \35939 , \35940 , \35941 , \35942 , \35943 , \35944 ,
         \35945 , \35946 , \35947 , \35948 , \35949 , \35950 , \35951 , \35952 , \35953 , \35954 ,
         \35955 , \35956 , \35957 , \35958 , \35959 , \35960 , \35961 , \35962 , \35963 , \35964 ,
         \35965 , \35966 , \35967 , \35968 , \35969 , \35970 , \35971 , \35972 , \35973 , \35974 ,
         \35975 , \35976 , \35977 , \35978 , \35979 , \35980 , \35981 , \35982 , \35983 , \35984 ,
         \35985 , \35986 , \35987 , \35988 , \35989 , \35990 , \35991 , \35992 , \35993 , \35994 ,
         \35995 , \35996 , \35997 , \35998 , \35999 , \36000 , \36001 , \36002 , \36003 , \36004 ,
         \36005 , \36006 , \36007 , \36008 , \36009 , \36010 , \36011 , \36012 , \36013 , \36014 ,
         \36015 , \36016 , \36017 , \36018 , \36019 , \36020 , \36021 , \36022 , \36023 , \36024 ,
         \36025 , \36026 , \36027 , \36028 , \36029 , \36030 , \36031 , \36032 , \36033 , \36034 ,
         \36035 , \36036 , \36037 , \36038 , \36039 , \36040 , \36041 , \36042 , \36043 , \36044 ,
         \36045 , \36046 , \36047 , \36048 , \36049 , \36050 , \36051 , \36052 , \36053 , \36054 ,
         \36055 , \36056 , \36057 , \36058 , \36059 , \36060 , \36061 , \36062 , \36063 , \36064 ,
         \36065 , \36066 , \36067 , \36068 , \36069 , \36070 , \36071 , \36072 , \36073 , \36074 ,
         \36075 , \36076 , \36077 , \36078 , \36079 , \36080 , \36081 , \36082 , \36083 , \36084 ,
         \36085 , \36086 , \36087 , \36088 , \36089 , \36090 , \36091 , \36092 , \36093 , \36094 ,
         \36095 , \36096 , \36097 , \36098 , \36099 , \36100 , \36101 , \36102 , \36103 , \36104 ,
         \36105 , \36106 , \36107 , \36108 , \36109 , \36110 , \36111 , \36112 , \36113 , \36114 ,
         \36115 , \36116 , \36117 , \36118 , \36119 , \36120 , \36121 , \36122 , \36123 , \36124 ,
         \36125 , \36126 , \36127 , \36128 , \36129 , \36130 , \36131 , \36132 , \36133 , \36134 ,
         \36135 , \36136 , \36137 , \36138 , \36139 , \36140 , \36141 , \36142 , \36143 , \36144 ,
         \36145 , \36146 , \36147 , \36148 , \36149 , \36150 , \36151 , \36152 , \36153 , \36154 ,
         \36155 , \36156 , \36157 , \36158 , \36159 , \36160 , \36161 , \36162 , \36163 , \36164 ,
         \36165 , \36166 , \36167 , \36168 , \36169 , \36170 , \36171 , \36172 , \36173 , \36174 ,
         \36175 , \36176 , \36177 , \36178 , \36179 , \36180 , \36181 , \36182 , \36183 , \36184 ,
         \36185 , \36186 , \36187 , \36188 , \36189 , \36190 , \36191 , \36192 , \36193 , \36194 ,
         \36195 , \36196 , \36197 , \36198 , \36199 , \36200 , \36201 , \36202 , \36203 , \36204 ,
         \36205 , \36206 , \36207 , \36208 , \36209 , \36210 , \36211 , \36212 , \36213 , \36214 ,
         \36215 , \36216 , \36217 , \36218 , \36219 , \36220 , \36221 , \36222 , \36223 , \36224 ,
         \36225 , \36226 , \36227 , \36228 , \36229 , \36230 , \36231 , \36232 , \36233 , \36234 ,
         \36235 , \36236 , \36237 , \36238 , \36239 , \36240 , \36241 , \36242 , \36243 , \36244 ,
         \36245 , \36246 , \36247 , \36248 , \36249 , \36250 , \36251 , \36252 , \36253 , \36254 ,
         \36255 , \36256 , \36257 , \36258 , \36259 , \36260 , \36261 , \36262 , \36263 , \36264 ,
         \36265 , \36266 , \36267 , \36268 , \36269 , \36270 , \36271 , \36272 , \36273 , \36274 ,
         \36275 , \36276 , \36277 , \36278 , \36279 , \36280 , \36281 , \36282 , \36283 , \36284 ,
         \36285 , \36286 , \36287 , \36288 , \36289 , \36290 , \36291 , \36292 , \36293 , \36294 ,
         \36295 , \36296 , \36297 , \36298 , \36299 , \36300 , \36301 , \36302 , \36303 , \36304 ,
         \36305 , \36306 , \36307 , \36308 , \36309 , \36310 , \36311 , \36312 , \36313 , \36314 ,
         \36315 , \36316 , \36317 , \36318 , \36319 , \36320 , \36321 , \36322 , \36323 , \36324 ,
         \36325 , \36326 , \36327 , \36328 , \36329 , \36330 , \36331 , \36332 , \36333 , \36334 ,
         \36335 , \36336 , \36337 , \36338 , \36339 , \36340 , \36341 , \36342 , \36343 , \36344 ,
         \36345_nGa51d , \36346 , \36347 , \36348 , \36349 , \36350 , \36351 , \36352 , \36353 , \36354 ,
         \36355 , \36356 , \36357 , \36358 , \36359 , \36360 , \36361 , \36362 , \36363 , \36364 ,
         \36365 , \36366 , \36367 , \36368 , \36369 , \36370 , \36371 , \36372 , \36373 , \36374 ,
         \36375 , \36376 , \36377 , \36378 , \36379 , \36380 , \36381 , \36382 , \36383 , \36384 ,
         \36385 , \36386 , \36387 , \36388 , \36389 , \36390 , \36391 , \36392 , \36393 , \36394 ,
         \36395 , \36396 , \36397 , \36398 , \36399 , \36400 , \36401 , \36402 , \36403 , \36404 ,
         \36405 , \36406 , \36407 , \36408 , \36409 , \36410 , \36411 , \36412 , \36413 , \36414 ,
         \36415 , \36416 , \36417 , \36418 , \36419 , \36420 , \36421 , \36422 , \36423 , \36424 ,
         \36425 , \36426 , \36427 , \36428 , \36429 , \36430 , \36431 , \36432 , \36433 , \36434 ,
         \36435 , \36436 , \36437 , \36438 , \36439 , \36440 , \36441 , \36442 , \36443 , \36444 ,
         \36445 , \36446 , \36447 , \36448 , \36449 , \36450 , \36451 , \36452 , \36453 , \36454 ,
         \36455 , \36456 , \36457 , \36458 , \36459 , \36460 , \36461 , \36462 , \36463 , \36464 ,
         \36465 , \36466 , \36467 , \36468 , \36469 , \36470 , \36471 , \36472 , \36473 , \36474 ,
         \36475 , \36476 , \36477 , \36478 , \36479 , \36480 , \36481 , \36482 , \36483 , \36484 ,
         \36485 , \36486 , \36487 , \36488 , \36489 , \36490 , \36491 , \36492 , \36493 , \36494 ,
         \36495 , \36496 , \36497 , \36498 , \36499 , \36500 , \36501 , \36502 , \36503 , \36504 ,
         \36505 , \36506 , \36507 , \36508 , \36509 , \36510 , \36511 , \36512 , \36513 , \36514 ,
         \36515 , \36516 , \36517 , \36518 , \36519 , \36520 , \36521 , \36522 , \36523 , \36524 ,
         \36525 , \36526 , \36527 , \36528 , \36529 , \36530 , \36531 , \36532 , \36533 , \36534 ,
         \36535 , \36536 , \36537 , \36538 , \36539 , \36540 , \36541 , \36542 , \36543 , \36544 ,
         \36545 , \36546 , \36547 , \36548 , \36549 , \36550 , \36551 , \36552 , \36553 , \36554 ,
         \36555 , \36556 , \36557 , \36558 , \36559 , \36560 , \36561 , \36562 , \36563 , \36564 ,
         \36565 , \36566 , \36567 , \36568 , \36569 , \36570 , \36571 , \36572 , \36573 , \36574 ,
         \36575 , \36576 , \36577 , \36578 , \36579 , \36580 , \36581 , \36582 , \36583 , \36584 ,
         \36585 , \36586 , \36587 , \36588 , \36589 , \36590 , \36591 , \36592 , \36593 , \36594 ,
         \36595 , \36596 , \36597 , \36598 , \36599 , \36600 , \36601 , \36602 , \36603 , \36604 ,
         \36605 , \36606 , \36607 , \36608 , \36609 , \36610 , \36611 , \36612 , \36613 , \36614 ,
         \36615 , \36616 , \36617 , \36618 , \36619 , \36620 , \36621 , \36622 , \36623 , \36624 ,
         \36625 , \36626 , \36627 , \36628 , \36629 , \36630 , \36631 , \36632 , \36633 , \36634 ,
         \36635 , \36636 , \36637 , \36638 , \36639 , \36640 , \36641 , \36642 , \36643 , \36644 ,
         \36645 , \36646 , \36647 , \36648 , \36649 , \36650 , \36651 , \36652 , \36653 , \36654 ,
         \36655 , \36656 , \36657 , \36658 , \36659 , \36660 , \36661 , \36662 , \36663 , \36664 ,
         \36665 , \36666 , \36667 , \36668 , \36669 , \36670 , \36671 , \36672 , \36673 , \36674 ,
         \36675 , \36676 , \36677 , \36678 , \36679 , \36680 , \36681 , \36682 , \36683 , \36684 ,
         \36685 , \36686 , \36687 , \36688 , \36689 , \36690 , \36691 , \36692 , \36693 , \36694 ,
         \36695 , \36696 , \36697 , \36698 , \36699 , \36700 , \36701 , \36702 , \36703 , \36704 ,
         \36705 , \36706 , \36707 , \36708 , \36709 , \36710 , \36711 , \36712 , \36713 , \36714 ,
         \36715 , \36716 , \36717 , \36718 , \36719 , \36720 , \36721 , \36722 , \36723 , \36724 ,
         \36725 , \36726 , \36727 , \36728 , \36729 , \36730 , \36731 , \36732 , \36733 , \36734 ,
         \36735 , \36736 , \36737 , \36738 , \36739 , \36740 , \36741 , \36742 , \36743 , \36744 ,
         \36745 , \36746 , \36747 , \36748 , \36749 , \36750 , \36751 , \36752 , \36753 , \36754 ,
         \36755 , \36756 , \36757 , \36758 , \36759 , \36760 , \36761 , \36762 , \36763 , \36764 ,
         \36765 , \36766 , \36767 , \36768 , \36769 , \36770 , \36771 , \36772 , \36773 , \36774 ,
         \36775 , \36776 , \36777 , \36778 , \36779 , \36780 , \36781 , \36782 , \36783 , \36784 ,
         \36785 , \36786 , \36787 , \36788 , \36789 , \36790 , \36791 , \36792 , \36793 , \36794 ,
         \36795 , \36796 , \36797 , \36798 , \36799 , \36800 , \36801 , \36802 , \36803 , \36804 ,
         \36805 , \36806 , \36807 , \36808 , \36809 , \36810 , \36811 , \36812 , \36813 , \36814 ,
         \36815 , \36816 , \36817 , \36818 , \36819 , \36820 , \36821 , \36822 , \36823 , \36824 ,
         \36825 , \36826 , \36827 , \36828 , \36829 , \36830 , \36831 , \36832 , \36833 , \36834 ,
         \36835 , \36836 , \36837 , \36838 , \36839 , \36840 , \36841 , \36842 , \36843 , \36844 ,
         \36845 , \36846 , \36847 , \36848 , \36849 , \36850 , \36851 , \36852 , \36853 , \36854 ,
         \36855 , \36856_nGa71c , \36857 , \36858 , \36859 , \36860 , \36861 , \36862 , \36863 , \36864 ,
         \36865 , \36866 , \36867 , \36868 , \36869 , \36870 , \36871 , \36872 , \36873 , \36874 ,
         \36875 , \36876 , \36877_nGa731 , \36878 , \36879 , \36880 , \36881 , \36882 , \36883 , \36884 ,
         \36885 , \36886 , \36887 , \36888 , \36889 , \36890 , \36891 , \36892 , \36893 , \36894 ,
         \36895 , \36896 , \36897 , \36898 , \36899_nGa747 , \36900 , \36901 , \36902 , \36903 , \36904 ,
         \36905 , \36906 , \36907 , \36908 , \36909 , \36910 , \36911 , \36912 , \36913 , \36914 ,
         \36915 , \36916 , \36917 , \36918 , \36919 , \36920 , \36921_nGa75d , \36922 , \36923 , \36924 ,
         \36925 , \36926 , \36927 , \36928 , \36929 , \36930 , \36931 , \36932 , \36933 , \36934 ,
         \36935 , \36936 , \36937 , \36938 , \36939 , \36940 , \36941 , \36942 , \36943_nGa773 , \36944 ,
         \36945 , \36946 , \36947 , \36948 , \36949 , \36950 , \36951 , \36952 , \36953 , \36954 ,
         \36955 , \36956 , \36957 , \36958 , \36959 , \36960 , \36961 , \36962 , \36963 , \36964 ,
         \36965_nGa789 , \36966 , \36967 , \36968 , \36969 , \36970 , \36971 , \36972 , \36973 , \36974 ,
         \36975 , \36976 , \36977 , \36978 , \36979 , \36980 , \36981 , \36982 , \36983 , \36984 ,
         \36985 , \36986 , \36987_nGa79f , \36988 , \36989 , \36990 , \36991 , \36992 , \36993 , \36994 ,
         \36995 , \36996 , \36997 , \36998 , \36999 , \37000 , \37001 , \37002 , \37003 , \37004 ,
         \37005 , \37006 , \37007 , \37008 , \37009_nGa7b5 , \37010 , \37011 , \37012 , \37013 , \37014 ,
         \37015 , \37016 , \37017 , \37018 , \37019 , \37020 , \37021 , \37022 , \37023 , \37024 ,
         \37025 , \37026 , \37027 , \37028 , \37029 , \37030 , \37031 , \37032 , \37033 , \37034 ,
         \37035 , \37036 , \37037 , \37038 , \37039 , \37040 , \37041 , \37042 , \37043 , \37044 ,
         \37045 , \37046 , \37047 , \37048 , \37049 , \37050 , \37051 , \37052 , \37053 , \37054 ,
         \37055 , \37056 , \37057 , \37058 , \37059 , \37060 , \37061 , \37062 , \37063 , \37064 ,
         \37065 , \37066 , \37067 , \37068 , \37069 , \37070 , \37071 , \37072 , \37073 , \37074 ,
         \37075 , \37076 , \37077 , \37078 , \37079 , \37080 , \37081 , \37082 , \37083 , \37084 ,
         \37085 , \37086 , \37087 , \37088 , \37089 , \37090 , \37091 , \37092 , \37093 , \37094 ,
         \37095 , \37096 , \37097 , \37098 , \37099 , \37100 , \37101 , \37102 , \37103 , \37104 ,
         \37105 , \37106 , \37107 , \37108 , \37109 , \37110 , \37111 , \37112 , \37113 , \37114 ,
         \37115 , \37116 , \37117 , \37118 , \37119 , \37120 , \37121 , \37122 , \37123 , \37124 ,
         \37125 , \37126 , \37127 , \37128 , \37129 , \37130 , \37131 , \37132 , \37133 , \37134 ,
         \37135 , \37136 , \37137 , \37138 , \37139 , \37140 , \37141 , \37142 , \37143 , \37144 ,
         \37145 , \37146 , \37147 , \37148 , \37149 , \37150 , \37151 , \37152 , \37153 , \37154 ,
         \37155 , \37156 , \37157 , \37158 , \37159 , \37160 , \37161 , \37162 , \37163 , \37164 ,
         \37165 , \37166 , \37167 , \37168 , \37169 , \37170 , \37171 , \37172 , \37173 , \37174 ,
         \37175 , \37176 , \37177 , \37178 , \37179 , \37180 , \37181 , \37182 , \37183 , \37184 ,
         \37185 , \37186 , \37187 , \37188 , \37189 , \37190 , \37191 , \37192 , \37193 , \37194 ,
         \37195 , \37196 , \37197 , \37198 , \37199 , \37200 , \37201 , \37202 , \37203 , \37204 ,
         \37205 , \37206 , \37207 , \37208 , \37209 , \37210 , \37211 , \37212 , \37213 , \37214 ,
         \37215 , \37216 , \37217 , \37218 , \37219 , \37220 , \37221 , \37222 , \37223 , \37224 ,
         \37225 , \37226 , \37227 , \37228 , \37229 , \37230 , \37231 , \37232 , \37233 , \37234 ,
         \37235 , \37236 , \37237 , \37238 , \37239 , \37240 , \37241 , \37242 , \37243 , \37244 ,
         \37245 , \37246 , \37247 , \37248 , \37249 , \37250 , \37251 , \37252 , \37253 , \37254 ,
         \37255 , \37256 , \37257 , \37258 , \37259 , \37260 , \37261 , \37262 , \37263 , \37264 ,
         \37265 , \37266 , \37267 , \37268 , \37269 , \37270 , \37271 , \37272 , \37273 , \37274 ,
         \37275 , \37276 , \37277 , \37278 , \37279 , \37280 , \37281 , \37282 , \37283 , \37284 ,
         \37285 , \37286 , \37287 , \37288 , \37289 , \37290 , \37291 , \37292 , \37293 , \37294 ,
         \37295 , \37296 , \37297 , \37298 , \37299 , \37300 , \37301 , \37302 , \37303 , \37304 ,
         \37305 , \37306 , \37307 , \37308 , \37309 , \37310 , \37311 , \37312 , \37313 , \37314 ,
         \37315 , \37316 , \37317 , \37318 , \37319 , \37320 , \37321 , \37322 , \37323 , \37324 ,
         \37325 , \37326 , \37327 , \37328 , \37329 , \37330 , \37331 , \37332 , \37333 , \37334 ,
         \37335 , \37336 , \37337 , \37338 , \37339 , \37340 , \37341 , \37342 , \37343 , \37344 ,
         \37345 , \37346 , \37347 , \37348 , \37349 , \37350 , \37351 , \37352 , \37353 , \37354 ,
         \37355 , \37356 , \37357 , \37358 , \37359 , \37360 , \37361 , \37362 , \37363 , \37364 ,
         \37365 , \37366 , \37367 , \37368 , \37369 , \37370 , \37371 , \37372 , \37373 , \37374 ,
         \37375 , \37376 , \37377 , \37378 , \37379 , \37380 , \37381 , \37382 , \37383 , \37384 ,
         \37385 , \37386 , \37387 , \37388 , \37389 , \37390 , \37391 , \37392 , \37393 , \37394 ,
         \37395 , \37396 , \37397 , \37398 , \37399 , \37400 , \37401 , \37402 , \37403 , \37404 ,
         \37405 , \37406 , \37407 , \37408 , \37409 , \37410 , \37411 , \37412 , \37413 , \37414 ,
         \37415 , \37416 , \37417 , \37418 , \37419 , \37420 , \37421 , \37422 , \37423 , \37424 ,
         \37425 , \37426 , \37427 , \37428 , \37429 , \37430 , \37431 , \37432 , \37433 , \37434 ,
         \37435 , \37436 , \37437 , \37438 , \37439 , \37440 , \37441 , \37442 , \37443 , \37444 ,
         \37445 , \37446 , \37447 , \37448 , \37449 , \37450 , \37451 , \37452 , \37453 , \37454 ,
         \37455 , \37456 , \37457 , \37458 , \37459 , \37460 , \37461 , \37462 , \37463 , \37464 ,
         \37465 , \37466 , \37467 , \37468 , \37469 , \37470 , \37471 , \37472 , \37473 , \37474 ,
         \37475 , \37476 , \37477 , \37478 , \37479 , \37480 , \37481 , \37482 , \37483 , \37484 ,
         \37485 , \37486 , \37487 , \37488 , \37489 , \37490 , \37491 , \37492 , \37493 , \37494 ,
         \37495 , \37496 , \37497 , \37498 , \37499 , \37500 , \37501 , \37502 , \37503 , \37504 ,
         \37505 , \37506 , \37507 , \37508 , \37509 , \37510 , \37511 , \37512 , \37513 , \37514 ,
         \37515 , \37516 , \37517 , \37518 , \37519 , \37520 , \37521 , \37522 , \37523 , \37524 ,
         \37525_nGa9b9 , \37526 , \37527 , \37528 , \37529 , \37530 , \37531 , \37532 , \37533 , \37534 ,
         \37535 , \37536 , \37537 , \37538 , \37539 , \37540 , \37541 , \37542 , \37543 , \37544 ,
         \37545 , \37546_nGa9ce , \37547 , \37548 , \37549 , \37550 , \37551 , \37552 , \37553 , \37554 ,
         \37555 , \37556 , \37557 , \37558 , \37559 , \37560 , \37561 , \37562 , \37563 , \37564 ,
         \37565 , \37566 , \37567 , \37568_nGa9e4 , \37569 , \37570 , \37571 , \37572 , \37573 , \37574 ,
         \37575 , \37576 , \37577 , \37578 , \37579 , \37580 , \37581 , \37582 , \37583 , \37584 ,
         \37585 , \37586 , \37587 , \37588 , \37589 , \37590_nGa9fa , \37591 , \37592 , \37593 , \37594 ,
         \37595 , \37596 , \37597 , \37598 , \37599 , \37600 , \37601 , \37602 , \37603 , \37604 ,
         \37605 , \37606 , \37607 , \37608 , \37609 , \37610 , \37611 , \37612_nGaa10 , \37613 , \37614 ,
         \37615 , \37616 , \37617 , \37618 , \37619 , \37620 , \37621 , \37622 , \37623 , \37624 ,
         \37625 , \37626 , \37627 , \37628 , \37629 , \37630 , \37631 , \37632 , \37633 , \37634_nGaa26 ,
         \37635 , \37636 , \37637 , \37638 , \37639 , \37640 , \37641 , \37642 , \37643 , \37644 ,
         \37645 , \37646 , \37647 , \37648 , \37649 , \37650 , \37651 , \37652 , \37653 , \37654 ,
         \37655 , \37656_nGaa3c , \37657 , \37658 , \37659 , \37660 , \37661 , \37662 , \37663 , \37664 ,
         \37665 , \37666 , \37667 , \37668 , \37669 , \37670 , \37671 , \37672 , \37673 , \37674 ,
         \37675 , \37676 , \37677 , \37678_nGaa52 , \37679 , \37680 , \37681 , \37682 , \37683 , \37684 ,
         \37685_nGaa59 , \37686 , \37687 , \37688 , \37689 , \37690 , \37691 , \37692 , \37693 , \37694 ,
         \37695 , \37696_nGaa64 , \37697 , \37698 , \37699 , \37700 , \37701 , \37702 , \37703 , \37704 ,
         \37705 , \37706 , \37707 , \37708 , \37709 , \37710 , \37711 , \37712 , \37713 , \37714 ,
         \37715 , \37716 , \37717 , \37718 , \37719 , \37720 , \37721 , \37722 , \37723 , \37724 ,
         \37725 , \37726 , \37727 , \37728 , \37729 , \37730 , \37731 , \37732 , \37733 , \37734 ,
         \37735 , \37736 , \37737 , \37738 , \37739 , \37740 , \37741 , \37742 , \37743 , \37744 ,
         \37745 , \37746 , \37747 , \37748 , \37749 , \37750 , \37751 , \37752 , \37753 , \37754 ,
         \37755 , \37756 , \37757 , \37758 , \37759 , \37760 , \37761 , \37762 , \37763 , \37764 ,
         \37765 , \37766_nGaaaa , \37767 , \37768 , \37769 , \37770 , \37771 , \37772 , \37773 , \37774 ,
         \37775 , \37776 , \37777 , \37778 , \37779 , \37780 , \37781 , \37782 , \37783 , \37784 ,
         \37785 , \37786_nGaabe , \37787 , \37788 , \37789 , \37790 , \37791 , \37792 , \37793 , \37794 ,
         \37795 , \37796 , \37797 , \37798 , \37799 , \37800 , \37801 , \37802 , \37803 , \37804 ,
         \37805 , \37806 , \37807_nGaad3 , \37808 , \37809 , \37810 , \37811 , \37812 , \37813 , \37814 ,
         \37815 , \37816 , \37817 , \37818 , \37819 , \37820 , \37821 , \37822 , \37823 , \37824 ,
         \37825 , \37826 , \37827 , \37828 , \37829_nGaae9 , \37830 , \37831 , \37832 , \37833 , \37834 ,
         \37835 , \37836 , \37837 , \37838 , \37839 , \37840 , \37841 , \37842 , \37843 , \37844 ,
         \37845 , \37846 , \37847 , \37848 , \37849 , \37850 , \37851_nGaaff , \37852 , \37853 , \37854 ,
         \37855 , \37856 , \37857 , \37858 , \37859 , \37860 , \37861 , \37862 , \37863 , \37864 ,
         \37865 , \37866 , \37867 , \37868 , \37869 , \37870 , \37871 , \37872 , \37873_nGab15 , \37874 ,
         \37875 , \37876 , \37877 , \37878 , \37879 , \37880 , \37881 , \37882 , \37883 , \37884 ,
         \37885 , \37886 , \37887 , \37888 , \37889 , \37890 , \37891 , \37892 , \37893 , \37894 ,
         \37895_nGab2b , \37896 , \37897 , \37898 , \37899 , \37900 , \37901 , \37902 , \37903 , \37904 ,
         \37905 , \37906 , \37907 , \37908 , \37909 , \37910 , \37911 , \37912 , \37913 , \37914 ,
         \37915 , \37916 , \37917_nGab41 , \37918 , \37919 , \37920 , \37921 , \37922 , \37923 , \37924 ,
         \37925 , \37926 , \37927 , \37928 , \37929 , \37930 , \37931 , \37932 , \37933 , \37934 ,
         \37935 , \37936 , \37937 , \37938 , \37939_nGab57 , \37940 , \37941 , \37942 , \37943 , \37944 ,
         \37945 , \37946 , \37947 , \37948 , \37949 , \37950 , \37951 , \37952 , \37953 , \37954 ,
         \37955 , \37956 , \37957 , \37958 , \37959 , \37960 , \37961 , \37962 , \37963_nGab6f , \37964 ,
         \37965 , \37966 , \37967 , \37968 , \37969 , \37970 , \37971 , \37972 , \37973 , \37974 ,
         \37975 , \37976 , \37977 , \37978 , \37979 , \37980 , \37981 , \37982 , \37983 , \37984_nGab84 ,
         \37985 , \37986 , \37987 , \37988 , \37989 , \37990 , \37991 , \37992 , \37993 , \37994 ,
         \37995 , \37996 , \37997 , \37998 , \37999 , \38000 , \38001 , \38002 , \38003 , \38004 ,
         \38005 , \38006_nGab9a , \38007 , \38008 , \38009 , \38010 , \38011 , \38012 , \38013 , \38014 ,
         \38015 , \38016 , \38017 , \38018 , \38019 , \38020 , \38021 , \38022 , \38023 , \38024 ,
         \38025 , \38026 , \38027 , \38028_nGabb0 , \38029 , \38030 , \38031 , \38032 , \38033 , \38034 ,
         \38035 , \38036 , \38037 , \38038 , \38039 , \38040 , \38041 , \38042 , \38043 , \38044 ,
         \38045 , \38046 , \38047 , \38048 , \38049 , \38050_nGabc6 , \38051 , \38052 , \38053 , \38054 ,
         \38055 , \38056 , \38057 , \38058 , \38059 , \38060 , \38061 , \38062 , \38063 , \38064 ,
         \38065 , \38066 , \38067 , \38068 , \38069 , \38070 , \38071 , \38072_nGabdc , \38073 , \38074 ,
         \38075 , \38076 , \38077 , \38078 , \38079 , \38080 , \38081 , \38082 , \38083 , \38084 ,
         \38085 , \38086 , \38087 , \38088 , \38089 , \38090 , \38091 , \38092 , \38093 , \38094_nGabf2 ,
         \38095 , \38096 , \38097 , \38098 , \38099 , \38100 , \38101 , \38102 , \38103 , \38104 ,
         \38105 , \38106 , \38107 , \38108 , \38109 , \38110 , \38111 , \38112 , \38113 , \38114 ,
         \38115 , \38116_nGac08 , \38117 , \38118 , \38119 , \38120 , \38121 , \38122 , \38123 , \38124_nGac10 ,
         \38125 , \38126 , \38127 , \38128 , \38129 , \38130 , \38131 , \38132 , \38133 , \38134 ,
         \38135 , \38136 , \38137 , \38138 , \38139 , \38140 , \38141 , \38142 , \38143 , \38144 ,
         \38145 , \38146 , \38147 , \38148 , \38149 , \38150 , \38151 , \38152 , \38153 , \38154 ,
         \38155 , \38156 , \38157 , \38158 , \38159 , \38160 , \38161 , \38162 , \38163 , \38164 ,
         \38165 , \38166 , \38167 , \38168 , \38169 , \38170 , \38171 , \38172 , \38173 , \38174 ,
         \38175 , \38176 , \38177 , \38178 , \38179 , \38180 , \38181 , \38182 , \38183 , \38184 ,
         \38185 , \38186 , \38187 , \38188 , \38189 , \38190 , \38191 , \38192 , \38193 , \38194 ,
         \38195 , \38196 , \38197 , \38198 , \38199 , \38200 , \38201 , \38202 , \38203 , \38204 ,
         \38205 , \38206 , \38207 , \38208 , \38209 , \38210 , \38211 , \38212 , \38213 , \38214 ,
         \38215 , \38216 , \38217 , \38218 , \38219 , \38220 , \38221 , \38222 , \38223 , \38224 ,
         \38225 , \38226 , \38227 , \38228 , \38229 , \38230 , \38231 , \38232 , \38233 , \38234 ,
         \38235 , \38236 , \38237 , \38238 , \38239 , \38240 , \38241 , \38242 , \38243 , \38244 ,
         \38245 , \38246 , \38247 , \38248 , \38249 , \38250 , \38251 , \38252 , \38253 , \38254 ,
         \38255 , \38256 , \38257 , \38258 , \38259 , \38260 , \38261 , \38262 , \38263 , \38264 ,
         \38265 , \38266 , \38267 , \38268 , \38269 , \38270 , \38271 , \38272 , \38273 , \38274 ,
         \38275 , \38276 , \38277 , \38278 , \38279 , \38280 , \38281 , \38282 , \38283 , \38284 ,
         \38285 , \38286 , \38287 , \38288 , \38289 , \38290 , \38291 , \38292 , \38293 , \38294 ,
         \38295 , \38296 , \38297 , \38298 , \38299 , \38300 , \38301 , \38302 , \38303 , \38304 ,
         \38305 , \38306 , \38307 , \38308 , \38309 , \38310 , \38311 , \38312 , \38313 , \38314 ,
         \38315 , \38316 , \38317 , \38318 , \38319 , \38320 , \38321 , \38322 , \38323 , \38324 ,
         \38325 , \38326 , \38327 , \38328 , \38329 , \38330 , \38331 , \38332 , \38333 , \38334 ,
         \38335 , \38336 , \38337 , \38338 , \38339 , \38340 , \38341 , \38342 , \38343 , \38344 ,
         \38345 , \38346 , \38347 , \38348 , \38349 , \38350 , \38351 , \38352 , \38353 , \38354 ,
         \38355 , \38356 , \38357 , \38358 , \38359 , \38360 , \38361 , \38362 , \38363 , \38364 ,
         \38365 , \38366 , \38367 , \38368 , \38369 , \38370 , \38371 , \38372 , \38373 , \38374 ,
         \38375 , \38376 , \38377 , \38378 , \38379 , \38380 , \38381 , \38382 , \38383 , \38384 ,
         \38385 , \38386 , \38387 , \38388 , \38389 , \38390 , \38391 , \38392 , \38393 , \38394 ,
         \38395 , \38396 , \38397 , \38398 , \38399 , \38400 , \38401 , \38402 , \38403 , \38404 ,
         \38405 , \38406 , \38407 , \38408 , \38409 , \38410 , \38411 , \38412 , \38413 , \38414 ,
         \38415 , \38416 , \38417 , \38418 , \38419 , \38420 , \38421 , \38422 , \38423 , \38424 ,
         \38425 , \38426 , \38427 , \38428 , \38429 , \38430 , \38431 , \38432 , \38433 , \38434 ,
         \38435 , \38436 , \38437 , \38438 , \38439 , \38440 , \38441 , \38442 , \38443 , \38444 ,
         \38445 , \38446 , \38447 , \38448 , \38449 , \38450 , \38451 , \38452 , \38453 , \38454 ,
         \38455 , \38456 , \38457 , \38458 , \38459 , \38460 , \38461 , \38462 , \38463 , \38464 ,
         \38465 , \38466 , \38467 , \38468 , \38469 , \38470 , \38471 , \38472 , \38473 , \38474 ,
         \38475 , \38476 , \38477 , \38478 , \38479 , \38480 , \38481 , \38482 , \38483 , \38484 ,
         \38485 , \38486 , \38487 , \38488 , \38489 , \38490 , \38491 , \38492 , \38493 , \38494 ,
         \38495 , \38496 , \38497 , \38498 , \38499 , \38500 , \38501 , \38502 , \38503 , \38504 ,
         \38505 , \38506 , \38507 , \38508 , \38509 , \38510 , \38511 , \38512 , \38513 , \38514 ,
         \38515 , \38516 , \38517 , \38518 , \38519 , \38520 , \38521 , \38522 , \38523 , \38524 ,
         \38525 , \38526 , \38527 , \38528 , \38529 , \38530 , \38531 , \38532 , \38533 , \38534 ,
         \38535 , \38536 , \38537 , \38538 , \38539 , \38540 , \38541 , \38542 , \38543 , \38544 ,
         \38545 , \38546 , \38547 , \38548 , \38549 , \38550 , \38551 , \38552 , \38553 , \38554 ,
         \38555 , \38556 , \38557 , \38558 , \38559 , \38560 , \38561 , \38562 , \38563 , \38564 ,
         \38565 , \38566 , \38567 , \38568 , \38569 , \38570 , \38571 , \38572 , \38573 , \38574 ,
         \38575 , \38576 , \38577 , \38578 , \38579 , \38580 , \38581 , \38582 , \38583 , \38584 ,
         \38585 , \38586 , \38587 , \38588 , \38589 , \38590 , \38591 , \38592 , \38593 , \38594 ,
         \38595 , \38596 , \38597 , \38598 , \38599 , \38600 , \38601 , \38602 , \38603 , \38604 ,
         \38605 , \38606 , \38607 , \38608 , \38609 , \38610 , \38611 , \38612 , \38613 , \38614 ,
         \38615 , \38616 , \38617 , \38618 , \38619 , \38620 , \38621 , \38622 , \38623 , \38624 ,
         \38625 , \38626 , \38627 , \38628 , \38629 , \38630 , \38631 , \38632 , \38633 , \38634 ,
         \38635 , \38636 , \38637 , \38638 , \38639 , \38640 , \38641 , \38642 , \38643 , \38644 ,
         \38645 , \38646 , \38647 , \38648 , \38649 , \38650 , \38651_nGae27 , \38652 , \38653 , \38654 ,
         \38655 , \38656 , \38657 , \38658 , \38659 , \38660 , \38661 , \38662 , \38663 , \38664 ,
         \38665 , \38666 , \38667 , \38668 , \38669 , \38670 , \38671 , \38672 , \38673 , \38674 ,
         \38675 , \38676 , \38677 , \38678 , \38679 , \38680 , \38681 , \38682 , \38683 , \38684 ,
         \38685 , \38686 , \38687 , \38688 , \38689 , \38690 , \38691 , \38692 , \38693 , \38694 ,
         \38695 , \38696 , \38697 , \38698 , \38699 , \38700 , \38701 , \38702 , \38703 , \38704 ,
         \38705 , \38706 , \38707 , \38708 , \38709 , \38710 , \38711 , \38712 , \38713 , \38714 ,
         \38715 , \38716 , \38717 , \38718 , \38719 , \38720 , \38721 , \38722 , \38723 , \38724 ,
         \38725 , \38726 , \38727 , \38728 , \38729 , \38730 , \38731 , \38732 , \38733 , \38734 ,
         \38735 , \38736 , \38737 , \38738 , \38739 , \38740 , \38741 , \38742 , \38743 , \38744 ,
         \38745 , \38746 , \38747 , \38748 , \38749 , \38750 , \38751 , \38752 , \38753 , \38754 ,
         \38755 , \38756 , \38757 , \38758 , \38759 , \38760 , \38761 , \38762 , \38763 , \38764 ,
         \38765 , \38766 , \38767 , \38768 , \38769 , \38770 , \38771 , \38772 , \38773 , \38774 ,
         \38775 , \38776 , \38777 , \38778 , \38779 , \38780 , \38781 , \38782 , \38783 , \38784 ,
         \38785 , \38786 , \38787 , \38788 , \38789 , \38790 , \38791 , \38792 , \38793 , \38794 ,
         \38795 , \38796 , \38797 , \38798 , \38799 , \38800 , \38801 , \38802 , \38803 , \38804 ,
         \38805 , \38806 , \38807 , \38808 , \38809 , \38810 , \38811 , \38812 , \38813 , \38814 ,
         \38815 , \38816 , \38817 , \38818 , \38819 , \38820 , \38821 , \38822 , \38823 , \38824 ,
         \38825 , \38826 , \38827 , \38828 , \38829 , \38830 , \38831 , \38832 , \38833 , \38834 ,
         \38835 , \38836 , \38837 , \38838 , \38839 , \38840 , \38841 , \38842 , \38843 , \38844 ,
         \38845 , \38846 , \38847 , \38848 , \38849 , \38850 , \38851 , \38852 , \38853 , \38854 ,
         \38855 , \38856 , \38857 , \38858 , \38859 , \38860 , \38861 , \38862 , \38863 , \38864 ,
         \38865 , \38866 , \38867 , \38868 , \38869 , \38870 , \38871 , \38872 , \38873 , \38874 ,
         \38875 , \38876 , \38877 , \38878 , \38879 , \38880 , \38881 , \38882 , \38883 , \38884 ,
         \38885 , \38886 , \38887 , \38888 , \38889 , \38890 , \38891 , \38892 , \38893 , \38894 ,
         \38895 , \38896 , \38897 , \38898 , \38899 , \38900 , \38901 , \38902 , \38903 , \38904 ,
         \38905 , \38906 , \38907 , \38908 , \38909 , \38910 , \38911 , \38912 , \38913 , \38914 ,
         \38915 , \38916 , \38917 , \38918 , \38919 , \38920 , \38921 , \38922 , \38923 , \38924 ,
         \38925 , \38926 , \38927 , \38928 , \38929 , \38930 , \38931 , \38932 , \38933 , \38934 ,
         \38935 , \38936 , \38937 , \38938 , \38939 , \38940 , \38941 , \38942 , \38943 , \38944 ,
         \38945 , \38946 , \38947 , \38948 , \38949 , \38950 , \38951 , \38952 , \38953 , \38954 ,
         \38955 , \38956 , \38957 , \38958 , \38959 , \38960 , \38961 , \38962 , \38963 , \38964 ,
         \38965 , \38966 , \38967 , \38968 , \38969 , \38970 , \38971 , \38972 , \38973 , \38974 ,
         \38975 , \38976 , \38977 , \38978 , \38979 , \38980 , \38981 , \38982 , \38983 , \38984 ,
         \38985 , \38986 , \38987 , \38988 , \38989 , \38990 , \38991 , \38992 , \38993 , \38994 ,
         \38995 , \38996 , \38997 , \38998 , \38999 , \39000 , \39001 , \39002 , \39003 , \39004 ,
         \39005 , \39006 , \39007 , \39008 , \39009 , \39010 , \39011 , \39012 , \39013 , \39014 ,
         \39015 , \39016 , \39017 , \39018 , \39019 , \39020 , \39021 , \39022 , \39023 , \39024 ,
         \39025 , \39026 , \39027 , \39028 , \39029 , \39030 , \39031 , \39032 , \39033 , \39034 ,
         \39035 , \39036 , \39037 , \39038 , \39039 , \39040 , \39041 , \39042 , \39043 , \39044 ,
         \39045 , \39046 , \39047 , \39048 , \39049 , \39050 , \39051 , \39052 , \39053 , \39054 ,
         \39055 , \39056 , \39057 , \39058 , \39059 , \39060 , \39061 , \39062 , \39063 , \39064 ,
         \39065 , \39066 , \39067 , \39068 , \39069 , \39070 , \39071 , \39072 , \39073 , \39074 ,
         \39075 , \39076 , \39077 , \39078 , \39079 , \39080 , \39081 , \39082 , \39083 , \39084 ,
         \39085 , \39086 , \39087 , \39088 , \39089 , \39090 , \39091 , \39092 , \39093 , \39094 ,
         \39095 , \39096 , \39097 , \39098 , \39099 , \39100 , \39101 , \39102 , \39103 , \39104 ,
         \39105 , \39106 , \39107 , \39108 , \39109 , \39110 , \39111 , \39112 , \39113 , \39114 ,
         \39115 , \39116 , \39117 , \39118 , \39119 , \39120 , \39121 , \39122 , \39123 , \39124 ,
         \39125 , \39126 , \39127 , \39128 , \39129 , \39130 , \39131 , \39132 , \39133 , \39134 ,
         \39135 , \39136 , \39137 , \39138 , \39139 , \39140 , \39141 , \39142 , \39143 , \39144 ,
         \39145 , \39146 , \39147 , \39148 , \39149 , \39150 , \39151 , \39152 , \39153 , \39154 ,
         \39155 , \39156 , \39157 , \39158 , \39159 , \39160 , \39161 , \39162_nGb026 , \39163 , \39164 ,
         \39165 , \39166 , \39167 , \39168 , \39169 , \39170 , \39171 , \39172 , \39173 , \39174 ,
         \39175 , \39176 , \39177 , \39178 , \39179 , \39180 , \39181 , \39182 , \39183_nGb03b , \39184 ,
         \39185 , \39186 , \39187 , \39188 , \39189 , \39190 , \39191 , \39192 , \39193 , \39194 ,
         \39195 , \39196 , \39197 , \39198 , \39199 , \39200 , \39201 , \39202 , \39203 , \39204 ,
         \39205_nGb051 , \39206 , \39207 , \39208 , \39209 , \39210 , \39211 , \39212 , \39213 , \39214 ,
         \39215 , \39216 , \39217 , \39218 , \39219 , \39220 , \39221 , \39222 , \39223 , \39224 ,
         \39225 , \39226 , \39227_nGb067 , \39228 , \39229 , \39230 , \39231 , \39232 , \39233 , \39234 ,
         \39235 , \39236 , \39237 , \39238 , \39239 , \39240 , \39241 , \39242 , \39243 , \39244 ,
         \39245 , \39246 , \39247 , \39248 , \39249_nGb07d , \39250 , \39251 , \39252 , \39253 , \39254 ,
         \39255 , \39256 , \39257 , \39258 , \39259 , \39260 , \39261 , \39262 , \39263 , \39264 ,
         \39265 , \39266 , \39267 , \39268 , \39269 , \39270 , \39271_nGb093 , \39272 , \39273 , \39274 ,
         \39275 , \39276 , \39277 , \39278 , \39279 , \39280 , \39281 , \39282 , \39283 , \39284 ,
         \39285 , \39286 , \39287 , \39288 , \39289 , \39290 , \39291 , \39292 , \39293_nGb0a9 , \39294 ,
         \39295 , \39296 , \39297 , \39298 , \39299 , \39300 , \39301 , \39302 , \39303 , \39304 ,
         \39305 , \39306 , \39307 , \39308 , \39309 , \39310 , \39311 , \39312 , \39313 , \39314 ,
         \39315_nGb0bf , \39316 , \39317 , \39318 , \39319 , \39320 , \39321 , \39322 , \39323 , \39324 ,
         \39325 , \39326 , \39327 , \39328 , \39329 , \39330 , \39331 , \39332 , \39333 , \39334 ,
         \39335 , \39336 , \39337 , \39338 , \39339 , \39340 , \39341 , \39342 , \39343 , \39344 ,
         \39345 , \39346 , \39347 , \39348 , \39349 , \39350 , \39351 , \39352 , \39353 , \39354 ,
         \39355 , \39356 , \39357 , \39358 , \39359 , \39360 , \39361 , \39362 , \39363 , \39364 ,
         \39365 , \39366 , \39367 , \39368 , \39369 , \39370 , \39371 , \39372 , \39373 , \39374 ,
         \39375 , \39376 , \39377 , \39378 , \39379 , \39380 , \39381 , \39382 , \39383 , \39384 ,
         \39385 , \39386 , \39387 , \39388 , \39389 , \39390 , \39391 , \39392 , \39393 , \39394 ,
         \39395 , \39396 , \39397 , \39398 , \39399 , \39400 , \39401 , \39402 , \39403 , \39404 ,
         \39405 , \39406 , \39407 , \39408 , \39409 , \39410 , \39411 , \39412 , \39413 , \39414 ,
         \39415 , \39416 , \39417 , \39418 , \39419 , \39420 , \39421 , \39422 , \39423 , \39424 ,
         \39425 , \39426 , \39427 , \39428 , \39429 , \39430 , \39431 , \39432 , \39433 , \39434 ,
         \39435 , \39436 , \39437 , \39438 , \39439 , \39440 , \39441 , \39442 , \39443 , \39444 ,
         \39445 , \39446 , \39447 , \39448 , \39449 , \39450 , \39451 , \39452 , \39453 , \39454 ,
         \39455 , \39456 , \39457 , \39458 , \39459 , \39460 , \39461 , \39462 , \39463 , \39464 ,
         \39465 , \39466 , \39467 , \39468 , \39469 , \39470 , \39471 , \39472 , \39473 , \39474 ,
         \39475 , \39476 , \39477 , \39478 , \39479 , \39480 , \39481 , \39482 , \39483 , \39484 ,
         \39485 , \39486 , \39487 , \39488 , \39489 , \39490 , \39491 , \39492 , \39493 , \39494 ,
         \39495 , \39496 , \39497 , \39498 , \39499 , \39500 , \39501 , \39502 , \39503 , \39504 ,
         \39505 , \39506 , \39507 , \39508 , \39509 , \39510 , \39511 , \39512 , \39513 , \39514 ,
         \39515 , \39516 , \39517 , \39518 , \39519 , \39520 , \39521 , \39522 , \39523 , \39524 ,
         \39525 , \39526 , \39527 , \39528 , \39529 , \39530 , \39531 , \39532 , \39533 , \39534 ,
         \39535 , \39536 , \39537 , \39538 , \39539 , \39540 , \39541 , \39542 , \39543 , \39544 ,
         \39545 , \39546 , \39547 , \39548 , \39549 , \39550 , \39551 , \39552 , \39553 , \39554 ,
         \39555 , \39556 , \39557 , \39558 , \39559 , \39560 , \39561 , \39562 , \39563 , \39564 ,
         \39565 , \39566 , \39567 , \39568 , \39569 , \39570 , \39571 , \39572 , \39573 , \39574 ,
         \39575 , \39576 , \39577 , \39578 , \39579 , \39580 , \39581 , \39582 , \39583 , \39584 ,
         \39585 , \39586 , \39587 , \39588 , \39589 , \39590 , \39591 , \39592 , \39593 , \39594 ,
         \39595 , \39596 , \39597 , \39598 , \39599 , \39600 , \39601 , \39602 , \39603 , \39604 ,
         \39605 , \39606 , \39607 , \39608 , \39609 , \39610 , \39611 , \39612 , \39613 , \39614 ,
         \39615 , \39616 , \39617 , \39618 , \39619 , \39620 , \39621 , \39622 , \39623 , \39624 ,
         \39625 , \39626 , \39627 , \39628 , \39629 , \39630 , \39631 , \39632 , \39633 , \39634 ,
         \39635 , \39636 , \39637 , \39638 , \39639 , \39640 , \39641 , \39642 , \39643 , \39644 ,
         \39645 , \39646 , \39647 , \39648 , \39649 , \39650 , \39651 , \39652 , \39653 , \39654 ,
         \39655 , \39656 , \39657 , \39658 , \39659 , \39660 , \39661 , \39662 , \39663 , \39664 ,
         \39665 , \39666 , \39667 , \39668 , \39669 , \39670 , \39671 , \39672 , \39673 , \39674 ,
         \39675 , \39676 , \39677 , \39678 , \39679 , \39680 , \39681 , \39682 , \39683 , \39684 ,
         \39685 , \39686 , \39687 , \39688 , \39689 , \39690 , \39691 , \39692 , \39693 , \39694 ,
         \39695 , \39696 , \39697 , \39698 , \39699 , \39700 , \39701 , \39702 , \39703 , \39704 ,
         \39705 , \39706 , \39707 , \39708 , \39709 , \39710 , \39711 , \39712 , \39713 , \39714 ,
         \39715 , \39716 , \39717 , \39718 , \39719 , \39720 , \39721 , \39722 , \39723 , \39724 ,
         \39725 , \39726 , \39727 , \39728 , \39729 , \39730 , \39731 , \39732 , \39733 , \39734 ,
         \39735 , \39736 , \39737 , \39738 , \39739 , \39740 , \39741 , \39742 , \39743 , \39744 ,
         \39745 , \39746 , \39747 , \39748 , \39749 , \39750 , \39751 , \39752 , \39753 , \39754 ,
         \39755 , \39756 , \39757 , \39758 , \39759 , \39760 , \39761 , \39762 , \39763 , \39764 ,
         \39765 , \39766 , \39767 , \39768 , \39769 , \39770 , \39771 , \39772 , \39773 , \39774 ,
         \39775 , \39776 , \39777 , \39778 , \39779 , \39780 , \39781 , \39782 , \39783 , \39784 ,
         \39785 , \39786 , \39787 , \39788 , \39789 , \39790 , \39791 , \39792 , \39793 , \39794 ,
         \39795 , \39796 , \39797 , \39798 , \39799 , \39800 , \39801 , \39802 , \39803 , \39804 ,
         \39805 , \39806 , \39807 , \39808 , \39809 , \39810 , \39811 , \39812 , \39813 , \39814 ,
         \39815 , \39816 , \39817 , \39818 , \39819 , \39820 , \39821 , \39822 , \39823 , \39824 ,
         \39825 , \39826 , \39827 , \39828 , \39829 , \39830 , \39831_nGb2c3 , \39832 , \39833 , \39834 ,
         \39835 , \39836 , \39837 , \39838 , \39839 , \39840 , \39841 , \39842 , \39843 , \39844 ,
         \39845 , \39846 , \39847 , \39848 , \39849 , \39850 , \39851 , \39852_nGb2d8 , \39853 , \39854 ,
         \39855 , \39856 , \39857 , \39858 , \39859 , \39860 , \39861 , \39862 , \39863 , \39864 ,
         \39865 , \39866 , \39867 , \39868 , \39869 , \39870 , \39871 , \39872 , \39873 , \39874_nGb2ee ,
         \39875 , \39876 , \39877 , \39878 , \39879 , \39880 , \39881 , \39882 , \39883 , \39884 ,
         \39885 , \39886 , \39887 , \39888 , \39889 , \39890 , \39891 , \39892 , \39893 , \39894 ,
         \39895 , \39896_nGb304 , \39897 , \39898 , \39899 , \39900 , \39901 , \39902 , \39903 , \39904 ,
         \39905 , \39906 , \39907 , \39908 , \39909 , \39910 , \39911 , \39912 , \39913 , \39914 ,
         \39915 , \39916 , \39917 , \39918_nGb31a , \39919 , \39920 , \39921 , \39922 , \39923 , \39924 ,
         \39925 , \39926 , \39927 , \39928 , \39929 , \39930 , \39931 , \39932 , \39933 , \39934 ,
         \39935 , \39936 , \39937 , \39938 , \39939 , \39940_nGb330 , \39941 , \39942 , \39943 , \39944 ,
         \39945 , \39946 , \39947 , \39948 , \39949 , \39950 , \39951 , \39952 , \39953 , \39954 ,
         \39955 , \39956 , \39957 , \39958 , \39959 , \39960 , \39961 , \39962_nGb346 , \39963 , \39964 ,
         \39965 , \39966 , \39967 , \39968 , \39969 , \39970 , \39971 , \39972 , \39973 , \39974 ,
         \39975 , \39976 , \39977 , \39978 , \39979 , \39980 , \39981 , \39982 , \39983 , \39984_nGb35c ,
         \39985 , \39986 , \39987 , \39988 , \39989 , \39990 , \39991_nGb363 , \39992 , \39993 , \39994 ,
         \39995 , \39996 , \39997 , \39998 , \39999 , \40000 , \40001 , \40002_nGb36e , \40003 , \40004 ,
         \40005 , \40006 , \40007 , \40008 , \40009 , \40010 , \40011 , \40012 , \40013 , \40014 ,
         \40015 , \40016 , \40017 , \40018 , \40019 , \40020 , \40021 , \40022 , \40023 , \40024 ,
         \40025 , \40026 , \40027 , \40028 , \40029 , \40030 , \40031 , \40032 , \40033 , \40034 ,
         \40035 , \40036 , \40037 , \40038 , \40039 , \40040 , \40041 , \40042 , \40043 , \40044 ,
         \40045 , \40046 , \40047 , \40048 , \40049 , \40050 , \40051 , \40052 , \40053_nGb3a4 , \40054 ,
         \40055 , \40056 , \40057 , \40058 , \40059 , \40060 , \40061 , \40062 , \40063 , \40064 ,
         \40065 , \40066 , \40067 , \40068 , \40069 , \40070 , \40071 , \40072 , \40073_nGb3b8 , \40074 ,
         \40075 , \40076 , \40077 , \40078 , \40079 , \40080 , \40081 , \40082 , \40083 , \40084 ,
         \40085 , \40086 , \40087 , \40088 , \40089 , \40090 , \40091 , \40092 , \40093 , \40094_nGb3cd ,
         \40095 , \40096 , \40097 , \40098 , \40099 , \40100 , \40101 , \40102 , \40103 , \40104 ,
         \40105 , \40106 , \40107 , \40108 , \40109 , \40110 , \40111 , \40112 , \40113 , \40114 ,
         \40115 , \40116_nGb3e3 , \40117 , \40118 , \40119 , \40120 , \40121 , \40122 , \40123 , \40124 ,
         \40125 , \40126 , \40127 , \40128 , \40129 , \40130 , \40131 , \40132 , \40133 , \40134 ,
         \40135 , \40136 , \40137 , \40138_nGb3f9 , \40139 , \40140 , \40141 , \40142 , \40143 , \40144 ,
         \40145 , \40146 , \40147 , \40148 , \40149 , \40150 , \40151 , \40152 , \40153 , \40154 ,
         \40155 , \40156 , \40157 , \40158 , \40159 , \40160_nGb40f , \40161 , \40162 , \40163 , \40164 ,
         \40165 , \40166 , \40167 , \40168 , \40169 , \40170 , \40171 , \40172 , \40173 , \40174 ,
         \40175 , \40176 , \40177 , \40178 , \40179 , \40180 , \40181 , \40182_nGb425 , \40183 , \40184 ,
         \40185 , \40186 , \40187 , \40188 , \40189 , \40190 , \40191 , \40192 , \40193 , \40194 ,
         \40195 , \40196 , \40197 , \40198 , \40199 , \40200 , \40201 , \40202 , \40203 , \40204_nGb43b ,
         \40205 , \40206 , \40207 , \40208 , \40209 , \40210 , \40211 , \40212 , \40213 , \40214 ,
         \40215 , \40216 , \40217 , \40218 , \40219 , \40220 , \40221 , \40222 , \40223 , \40224 ,
         \40225 , \40226_nGb451 , \40227 , \40228 , \40229 , \40230 , \40231 , \40232 , \40233 , \40234 ,
         \40235 , \40236 , \40237 , \40238 , \40239 , \40240 , \40241 , \40242 , \40243 , \40244 ,
         \40245 , \40246 , \40247 , \40248 , \40249 , \40250_nGb469 , \40251 , \40252 , \40253 , \40254 ,
         \40255 , \40256 , \40257 , \40258 , \40259 , \40260 , \40261 , \40262 , \40263 , \40264 ,
         \40265 , \40266 , \40267 , \40268 , \40269 , \40270 , \40271_nGb47e , \40272 , \40273 , \40274 ,
         \40275 , \40276 , \40277 , \40278 , \40279 , \40280 , \40281 , \40282 , \40283 , \40284 ,
         \40285 , \40286 , \40287 , \40288 , \40289 , \40290 , \40291 , \40292 , \40293_nGb494 , \40294 ,
         \40295 , \40296 , \40297 , \40298 , \40299 , \40300 , \40301 , \40302 , \40303 , \40304 ,
         \40305 , \40306 , \40307 , \40308 , \40309 , \40310 , \40311 , \40312 , \40313 , \40314 ,
         \40315_nGb4aa , \40316 , \40317 , \40318 , \40319 , \40320 , \40321 , \40322 , \40323 , \40324 ,
         \40325 , \40326 , \40327 , \40328 , \40329 , \40330 , \40331 , \40332 , \40333 , \40334 ,
         \40335 , \40336 , \40337_nGb4c0 , \40338 , \40339 , \40340 , \40341 , \40342 , \40343 , \40344 ,
         \40345 , \40346 , \40347 , \40348 , \40349 , \40350 , \40351 , \40352 , \40353 , \40354 ,
         \40355 , \40356 , \40357 , \40358 , \40359_nGb4d6 , \40360 , \40361 , \40362 , \40363 , \40364 ,
         \40365 , \40366 , \40367 , \40368 , \40369 , \40370 , \40371 , \40372 , \40373 , \40374 ,
         \40375 , \40376 , \40377 , \40378 , \40379 , \40380 , \40381_nGb4ec , \40382 , \40383 , \40384 ,
         \40385 , \40386 , \40387 , \40388 , \40389 , \40390 , \40391 , \40392 , \40393 , \40394 ,
         \40395 , \40396 , \40397 , \40398 , \40399 , \40400 , \40401 , \40402 , \40403_nGb502 , \40404 ,
         \40405 , \40406 , \40407 , \40408 , \40409 , \40410 , \40411_nGb50a , \40412 , \40413 , \40414 ,
         \40415 , \40416 , \40417 , \40418 , \40419 , \40420 , \40421 , \40422 , \40423 , \40424 ,
         \40425 , \40426 , \40427 , \40428 , \40429 , \40430 , \40431 , \40432 , \40433 , \40434 ,
         \40435 , \40436 , \40437 , \40438 , \40439 , \40440 , \40441 , \40442 , \40443 , \40444 ,
         \40445 , \40446 , \40447 , \40448 , \40449 , \40450 , \40451 , \40452 , \40453 , \40454 ,
         \40455 , \40456 , \40457 , \40458 , \40459 , \40460 , \40461 , \40462 , \40463 , \40464 ,
         \40465 , \40466 , \40467 , \40468 , \40469 , \40470 , \40471 , \40472 , \40473 , \40474 ,
         \40475 , \40476 , \40477 , \40478 , \40479 , \40480 , \40481 , \40482 , \40483 , \40484 ,
         \40485 , \40486 , \40487 , \40488 , \40489 , \40490 , \40491 , \40492 , \40493 , \40494 ,
         \40495 , \40496 , \40497 , \40498 , \40499 , \40500 , \40501 , \40502 , \40503 , \40504 ,
         \40505 , \40506 , \40507 , \40508 , \40509 , \40510 , \40511 , \40512 , \40513 , \40514 ,
         \40515 , \40516 , \40517 , \40518 , \40519 , \40520 , \40521 , \40522 , \40523 , \40524 ,
         \40525 , \40526 , \40527 , \40528 , \40529 , \40530 , \40531 , \40532 , \40533 , \40534 ,
         \40535 , \40536 , \40537 , \40538 , \40539 , \40540 , \40541 , \40542 , \40543 , \40544 ,
         \40545 , \40546 , \40547 , \40548 , \40549 , \40550 , \40551 , \40552 , \40553 , \40554 ,
         \40555 , \40556 , \40557 , \40558 , \40559 , \40560 , \40561 , \40562 , \40563 , \40564 ,
         \40565 , \40566 , \40567 , \40568 , \40569 , \40570 , \40571 , \40572 , \40573 , \40574 ,
         \40575 , \40576 , \40577 , \40578 , \40579 , \40580 , \40581 , \40582 , \40583 , \40584 ,
         \40585 , \40586 , \40587 , \40588 , \40589 , \40590 , \40591 , \40592 , \40593 , \40594 ,
         \40595 , \40596 , \40597 , \40598 , \40599 , \40600 , \40601 , \40602 , \40603 , \40604 ,
         \40605 , \40606 , \40607 , \40608 , \40609 , \40610 , \40611 , \40612 , \40613 , \40614 ,
         \40615 , \40616 , \40617 , \40618 , \40619 , \40620 , \40621 , \40622 , \40623 , \40624 ,
         \40625 , \40626 , \40627 , \40628 , \40629 , \40630 , \40631 , \40632 , \40633 , \40634 ,
         \40635 , \40636 , \40637 , \40638 , \40639 , \40640 , \40641 , \40642 , \40643 , \40644 ,
         \40645 , \40646 , \40647 , \40648 , \40649 , \40650 , \40651 , \40652 , \40653 , \40654 ,
         \40655 , \40656 , \40657 , \40658 , \40659 , \40660 , \40661 , \40662 , \40663 , \40664 ,
         \40665 , \40666 , \40667 , \40668 , \40669 , \40670 , \40671 , \40672 , \40673 , \40674 ,
         \40675 , \40676 , \40677 , \40678 , \40679 , \40680 , \40681 , \40682 , \40683 , \40684 ,
         \40685 , \40686 , \40687 , \40688 , \40689 , \40690 , \40691 , \40692 , \40693 , \40694 ,
         \40695 , \40696 , \40697 , \40698 , \40699 , \40700 , \40701 , \40702 , \40703 , \40704 ,
         \40705 , \40706 , \40707 , \40708 , \40709 , \40710 , \40711 , \40712 , \40713 , \40714 ,
         \40715 , \40716 , \40717 , \40718 , \40719 , \40720 , \40721 , \40722 , \40723 , \40724 ,
         \40725 , \40726 , \40727 , \40728 , \40729 , \40730 , \40731 , \40732 , \40733 , \40734 ,
         \40735 , \40736 , \40737 , \40738 , \40739 , \40740 , \40741 , \40742 , \40743 , \40744 ,
         \40745 , \40746 , \40747 , \40748 , \40749 , \40750 , \40751 , \40752 , \40753 , \40754 ,
         \40755 , \40756 , \40757 , \40758 , \40759 , \40760 , \40761 , \40762 , \40763 , \40764 ,
         \40765 , \40766 , \40767 , \40768 , \40769 , \40770 , \40771 , \40772 , \40773 , \40774 ,
         \40775 , \40776 , \40777 , \40778 , \40779 , \40780 , \40781 , \40782 , \40783 , \40784 ,
         \40785 , \40786 , \40787 , \40788 , \40789 , \40790 , \40791 , \40792 , \40793 , \40794 ,
         \40795 , \40796 , \40797 , \40798 , \40799 , \40800 , \40801 , \40802 , \40803 , \40804 ,
         \40805 , \40806 , \40807 , \40808 , \40809 , \40810 , \40811 , \40812 , \40813 , \40814 ,
         \40815 , \40816 , \40817 , \40818 , \40819 , \40820 , \40821 , \40822 , \40823 , \40824 ,
         \40825 , \40826 , \40827 , \40828 , \40829 , \40830 , \40831 , \40832 , \40833 , \40834 ,
         \40835 , \40836 , \40837 , \40838 , \40839 , \40840 , \40841 , \40842 , \40843 , \40844 ,
         \40845 , \40846 , \40847 , \40848 , \40849 , \40850 , \40851 , \40852 , \40853 , \40854 ,
         \40855 , \40856 , \40857 , \40858 , \40859 , \40860 , \40861 , \40862 , \40863 , \40864 ,
         \40865 , \40866 , \40867 , \40868 , \40869 , \40870 , \40871 , \40872 , \40873 , \40874 ,
         \40875 , \40876 , \40877 , \40878 , \40879 , \40880 , \40881 , \40882 , \40883 , \40884 ,
         \40885 , \40886_nGb6e9 , \40887 , \40888 , \40889 , \40890 , \40891 , \40892 , \40893 , \40894 ,
         \40895 , \40896 , \40897 , \40898 , \40899 , \40900 , \40901 , \40902 , \40903 , \40904 ,
         \40905 , \40906 , \40907 , \40908 , \40909 , \40910 , \40911 , \40912 , \40913 , \40914 ,
         \40915 , \40916 , \40917 , \40918 , \40919 , \40920 , \40921 , \40922 , \40923 , \40924 ,
         \40925 , \40926 , \40927 , \40928 , \40929 , \40930 , \40931 , \40932 , \40933 , \40934 ,
         \40935 , \40936 , \40937 , \40938 , \40939 , \40940 , \40941 , \40942 , \40943 , \40944 ,
         \40945 , \40946 , \40947 , \40948 , \40949 , \40950 , \40951 , \40952 , \40953 , \40954 ,
         \40955 , \40956 , \40957 , \40958 , \40959 , \40960 , \40961 , \40962 , \40963 , \40964 ,
         \40965 , \40966 , \40967 , \40968 , \40969 , \40970 , \40971 , \40972 , \40973 , \40974 ,
         \40975 , \40976 , \40977 , \40978 , \40979 , \40980 , \40981 , \40982 , \40983 , \40984 ,
         \40985 , \40986 , \40987 , \40988 , \40989 , \40990 , \40991 , \40992 , \40993 , \40994 ,
         \40995 , \40996 , \40997 , \40998 , \40999 , \41000 , \41001 , \41002 , \41003 , \41004 ,
         \41005 , \41006 , \41007 , \41008 , \41009 , \41010 , \41011 , \41012 , \41013 , \41014 ,
         \41015 , \41016 , \41017 , \41018 , \41019 , \41020 , \41021 , \41022 , \41023 , \41024 ,
         \41025 , \41026 , \41027 , \41028 , \41029 , \41030 , \41031 , \41032 , \41033 , \41034 ,
         \41035 , \41036 , \41037 , \41038 , \41039 , \41040 , \41041 , \41042 , \41043 , \41044 ,
         \41045 , \41046 , \41047 , \41048 , \41049 , \41050 , \41051 , \41052 , \41053 , \41054 ,
         \41055 , \41056 , \41057 , \41058 , \41059 , \41060 , \41061 , \41062 , \41063 , \41064 ,
         \41065 , \41066 , \41067 , \41068 , \41069 , \41070 , \41071 , \41072 , \41073 , \41074 ,
         \41075 , \41076 , \41077 , \41078 , \41079 , \41080 , \41081 , \41082 , \41083 , \41084 ,
         \41085 , \41086 , \41087 , \41088 , \41089 , \41090 , \41091 , \41092 , \41093 , \41094 ,
         \41095 , \41096 , \41097 , \41098 , \41099 , \41100 , \41101 , \41102 , \41103 , \41104 ,
         \41105 , \41106 , \41107 , \41108 , \41109 , \41110 , \41111 , \41112 , \41113 , \41114 ,
         \41115 , \41116 , \41117 , \41118 , \41119 , \41120 , \41121 , \41122 , \41123 , \41124 ,
         \41125 , \41126 , \41127 , \41128 , \41129 , \41130 , \41131 , \41132 , \41133 , \41134 ,
         \41135 , \41136 , \41137 , \41138 , \41139 , \41140 , \41141 , \41142 , \41143 , \41144 ,
         \41145 , \41146 , \41147 , \41148 , \41149 , \41150 , \41151 , \41152 , \41153 , \41154 ,
         \41155 , \41156 , \41157 , \41158 , \41159 , \41160 , \41161 , \41162 , \41163 , \41164 ,
         \41165 , \41166 , \41167 , \41168 , \41169 , \41170 , \41171 , \41172 , \41173 , \41174 ,
         \41175 , \41176 , \41177 , \41178 , \41179 , \41180 , \41181 , \41182 , \41183 , \41184 ,
         \41185 , \41186 , \41187 , \41188 , \41189 , \41190 , \41191 , \41192 , \41193 , \41194 ,
         \41195 , \41196 , \41197 , \41198 , \41199 , \41200 , \41201 , \41202 , \41203 , \41204 ,
         \41205 , \41206 , \41207 , \41208 , \41209 , \41210 , \41211 , \41212 , \41213 , \41214 ,
         \41215 , \41216 , \41217 , \41218 , \41219 , \41220 , \41221 , \41222 , \41223 , \41224 ,
         \41225 , \41226 , \41227 , \41228 , \41229 , \41230 , \41231 , \41232 , \41233 , \41234 ,
         \41235 , \41236 , \41237 , \41238 , \41239 , \41240 , \41241 , \41242 , \41243 , \41244 ,
         \41245 , \41246 , \41247 , \41248 , \41249 , \41250 , \41251 , \41252 , \41253 , \41254 ,
         \41255 , \41256 , \41257 , \41258 , \41259 , \41260 , \41261 , \41262 , \41263 , \41264 ,
         \41265 , \41266 , \41267 , \41268 , \41269 , \41270 , \41271 , \41272 , \41273 , \41274 ,
         \41275 , \41276 , \41277 , \41278 , \41279 , \41280 , \41281 , \41282 , \41283 , \41284 ,
         \41285 , \41286 , \41287 , \41288 , \41289 , \41290 , \41291 , \41292 , \41293 , \41294 ,
         \41295 , \41296 , \41297 , \41298 , \41299 , \41300 , \41301 , \41302 , \41303 , \41304 ,
         \41305 , \41306 , \41307 , \41308 , \41309 , \41310 , \41311 , \41312 , \41313 , \41314 ,
         \41315 , \41316 , \41317 , \41318 , \41319 , \41320 , \41321 , \41322 , \41323 , \41324 ,
         \41325 , \41326 , \41327 , \41328 , \41329 , \41330 , \41331 , \41332 , \41333 , \41334 ,
         \41335 , \41336 , \41337 , \41338 , \41339 , \41340 , \41341 , \41342 , \41343 , \41344 ,
         \41345 , \41346 , \41347_nGb8b6 , \41348 , \41349 , \41350 , \41351 , \41352 , \41353 , \41354 ,
         \41355 , \41356 , \41357 , \41358 , \41359 , \41360 , \41361 , \41362 , \41363 , \41364 ,
         \41365 , \41366 , \41367_nGb8ca , \41368 , \41369 , \41370 , \41371 , \41372 , \41373 , \41374 ,
         \41375 , \41376 , \41377 , \41378 , \41379 , \41380 , \41381 , \41382 , \41383 , \41384 ,
         \41385 , \41386 , \41387 , \41388_nGb8df , \41389 , \41390 , \41391 , \41392 , \41393 , \41394 ,
         \41395 , \41396 , \41397 , \41398 , \41399 , \41400 , \41401 , \41402 , \41403 , \41404 ,
         \41405 , \41406 , \41407 , \41408 , \41409_nGb8f4 , \41410 , \41411 , \41412 , \41413 , \41414 ,
         \41415 , \41416 , \41417 , \41418 , \41419 , \41420 , \41421 , \41422 , \41423 , \41424 ,
         \41425 , \41426 , \41427 , \41428 , \41429 , \41430_nGb909 , \41431 , \41432 , \41433 , \41434 ,
         \41435 , \41436 , \41437 , \41438 , \41439 , \41440 , \41441 , \41442 , \41443 , \41444 ,
         \41445 , \41446 , \41447 , \41448 , \41449 , \41450 , \41451_nGb91e , \41452 , \41453 , \41454 ,
         \41455 , \41456 , \41457 , \41458 , \41459 , \41460 , \41461 , \41462 , \41463 , \41464 ,
         \41465 , \41466 , \41467 , \41468 , \41469 , \41470 , \41471 , \41472_nGb933 , \41473 , \41474 ,
         \41475 , \41476 , \41477 , \41478 , \41479 , \41480 , \41481 , \41482 , \41483 , \41484 ,
         \41485 , \41486 , \41487 , \41488 , \41489 , \41490 , \41491 , \41492 , \41493_nGb948 , \41494 ,
         \41495 , \41496 , \41497 , \41498 , \41499 , \41500 , \41501 , \41502 , \41503 , \41504 ,
         \41505 , \41506 , \41507 , \41508 , \41509 , \41510 , \41511 , \41512 , \41513 , \41514 ,
         \41515 , \41516 , \41517 , \41518 , \41519 , \41520 , \41521 , \41522 , \41523 , \41524 ,
         \41525 , \41526 , \41527 , \41528 , \41529 , \41530 , \41531 , \41532 , \41533 , \41534 ,
         \41535 , \41536 , \41537 , \41538 , \41539 , \41540 , \41541 , \41542 , \41543 , \41544 ,
         \41545 , \41546 , \41547 , \41548 , \41549 , \41550 , \41551 , \41552 , \41553 , \41554 ,
         \41555 , \41556 , \41557 , \41558 , \41559 , \41560 , \41561 , \41562 , \41563 , \41564 ,
         \41565 , \41566 , \41567 , \41568 , \41569 , \41570 , \41571 , \41572 , \41573 , \41574 ,
         \41575 , \41576 , \41577 , \41578 , \41579 , \41580 , \41581 , \41582 , \41583 , \41584 ,
         \41585 , \41586 , \41587 , \41588 , \41589 , \41590 , \41591 , \41592 , \41593 , \41594 ,
         \41595 , \41596 , \41597 , \41598 , \41599 , \41600 , \41601 , \41602 , \41603 , \41604 ,
         \41605 , \41606 , \41607 , \41608 , \41609 , \41610 , \41611 , \41612 , \41613 , \41614 ,
         \41615 , \41616 , \41617 , \41618 , \41619 , \41620 , \41621 , \41622 , \41623 , \41624 ,
         \41625 , \41626 , \41627 , \41628 , \41629 , \41630 , \41631 , \41632 , \41633 , \41634 ,
         \41635 , \41636 , \41637 , \41638 , \41639 , \41640 , \41641 , \41642 , \41643 , \41644 ,
         \41645 , \41646 , \41647 , \41648 , \41649 , \41650 , \41651 , \41652 , \41653 , \41654 ,
         \41655 , \41656 , \41657 , \41658 , \41659 , \41660 , \41661 , \41662 , \41663 , \41664 ,
         \41665 , \41666 , \41667 , \41668 , \41669 , \41670 , \41671 , \41672 , \41673 , \41674 ,
         \41675 , \41676 , \41677 , \41678 , \41679 , \41680 , \41681 , \41682 , \41683 , \41684 ,
         \41685 , \41686 , \41687 , \41688 , \41689 , \41690 , \41691 , \41692 , \41693 , \41694 ,
         \41695 , \41696 , \41697 , \41698 , \41699 , \41700 , \41701 , \41702 , \41703 , \41704 ,
         \41705 , \41706 , \41707 , \41708 , \41709 , \41710 , \41711 , \41712 , \41713 , \41714 ,
         \41715 , \41716 , \41717 , \41718 , \41719 , \41720 , \41721 , \41722 , \41723 , \41724 ,
         \41725 , \41726 , \41727 , \41728 , \41729 , \41730 , \41731 , \41732 , \41733 , \41734 ,
         \41735 , \41736 , \41737 , \41738 , \41739 , \41740 , \41741 , \41742 , \41743 , \41744 ,
         \41745 , \41746 , \41747 , \41748 , \41749 , \41750 , \41751 , \41752 , \41753 , \41754 ,
         \41755 , \41756 , \41757 , \41758 , \41759 , \41760 , \41761 , \41762 , \41763 , \41764 ,
         \41765 , \41766 , \41767 , \41768 , \41769 , \41770 , \41771 , \41772 , \41773 , \41774 ,
         \41775 , \41776 , \41777 , \41778 , \41779 , \41780 , \41781 , \41782 , \41783 , \41784 ,
         \41785 , \41786 , \41787 , \41788 , \41789 , \41790 , \41791 , \41792 , \41793 , \41794 ,
         \41795 , \41796 , \41797 , \41798 , \41799 , \41800 , \41801 , \41802 , \41803 , \41804 ,
         \41805 , \41806 , \41807 , \41808 , \41809 , \41810 , \41811 , \41812 , \41813 , \41814 ,
         \41815 , \41816 , \41817 , \41818 , \41819 , \41820 , \41821 , \41822 , \41823 , \41824 ,
         \41825 , \41826 , \41827 , \41828 , \41829 , \41830 , \41831 , \41832 , \41833 , \41834 ,
         \41835 , \41836 , \41837 , \41838 , \41839 , \41840 , \41841 , \41842 , \41843 , \41844 ,
         \41845 , \41846 , \41847 , \41848 , \41849 , \41850 , \41851 , \41852 , \41853 , \41854 ,
         \41855 , \41856 , \41857 , \41858 , \41859 , \41860 , \41861 , \41862 , \41863 , \41864 ,
         \41865 , \41866 , \41867 , \41868 , \41869 , \41870 , \41871 , \41872 , \41873 , \41874 ,
         \41875 , \41876 , \41877 , \41878 , \41879 , \41880 , \41881 , \41882 , \41883 , \41884 ,
         \41885 , \41886 , \41887 , \41888 , \41889 , \41890 , \41891 , \41892 , \41893 , \41894 ,
         \41895 , \41896 , \41897 , \41898 , \41899 , \41900 , \41901 , \41902 , \41903 , \41904 ,
         \41905 , \41906 , \41907 , \41908 , \41909 , \41910 , \41911 , \41912 , \41913 , \41914 ,
         \41915 , \41916 , \41917 , \41918 , \41919 , \41920 , \41921 , \41922 , \41923 , \41924 ,
         \41925 , \41926 , \41927 , \41928 , \41929 , \41930 , \41931 , \41932 , \41933 , \41934 ,
         \41935 , \41936 , \41937 , \41938 , \41939 , \41940 , \41941 , \41942 , \41943 , \41944 ,
         \41945 , \41946 , \41947 , \41948 , \41949 , \41950 , \41951 , \41952 , \41953 , \41954 ,
         \41955 , \41956 , \41957 , \41958 , \41959_nGbb1a , \41960 , \41961 , \41962 , \41963 , \41964 ,
         \41965 , \41966 , \41967 , \41968 , \41969 , \41970 , \41971 , \41972 , \41973 , \41974 ,
         \41975 , \41976 , \41977 , \41978 , \41979_nGbb2e , \41980 , \41981 , \41982 , \41983 , \41984 ,
         \41985 , \41986 , \41987 , \41988 , \41989 , \41990 , \41991 , \41992 , \41993 , \41994 ,
         \41995 , \41996 , \41997 , \41998 , \41999 , \42000_nGbb43 , \42001 , \42002 , \42003 , \42004 ,
         \42005 , \42006 , \42007 , \42008 , \42009 , \42010 , \42011 , \42012 , \42013 , \42014 ,
         \42015 , \42016 , \42017 , \42018 , \42019 , \42020 , \42021_nGbb58 , \42022 , \42023 , \42024 ,
         \42025 , \42026 , \42027 , \42028 , \42029 , \42030 , \42031 , \42032 , \42033 , \42034 ,
         \42035 , \42036 , \42037 , \42038 , \42039 , \42040 , \42041 , \42042_nGbb6d , \42043 , \42044 ,
         \42045 , \42046 , \42047 , \42048 , \42049 , \42050 , \42051 , \42052 , \42053 , \42054 ,
         \42055 , \42056 , \42057 , \42058 , \42059 , \42060 , \42061 , \42062 , \42063_nGbb82 , \42064 ,
         \42065 , \42066 , \42067 , \42068 , \42069 , \42070 , \42071 , \42072 , \42073 , \42074 ,
         \42075 , \42076 , \42077 , \42078 , \42079 , \42080 , \42081 , \42082 , \42083 , \42084_nGbb97 ,
         \42085 , \42086 , \42087 , \42088 , \42089 , \42090 , \42091 , \42092 , \42093 , \42094 ,
         \42095 , \42096 , \42097 , \42098 , \42099 , \42100 , \42101 , \42102 , \42103 , \42104 ,
         \42105_nGbbac , \42106 , \42107 , \42108 , \42109 , \42110 , \42111 , \42112_nGbbb3 , \42113 , \42114 ,
         \42115 , \42116 , \42117 , \42118 , \42119 , \42120 , \42121_nGbbbc , \42122_nGbbbd , \42123_nGbbbe , \42124_nGbbbf ,
         \42125_nGbbc0 , \42126_nGbbc1 , \42127_nGbbc2 , \42128_nGbbc3 , \42129_nGbbc4 , \42130_nGbbc5 , \42131_nGbbc6 , \42132_nGbbc7 , \42133_nGbbc8 , \42134_nGbbc9 ,
         \42135_nGbbca , \42136_nGbbcb , \42137_nGbbcc , \42138_nGbbcd , \42139_nGbbce , \42140_nGbbcf , \42141_nGbbd0 , \42142_nGbbd1 , \42143_nGbbd2 , \42144_nGbbd3 ,
         \42145_nGbbd4 , \42146_nGbbd5 , \42147_nGbbd6 , \42148_nGbbd7 , \42149_nGbbd8 , \42150_nGbbd9 , \42151_nGbbda , \42152_nGbbdb , \42153_nGbbdc , \42154_nGbbdd ,
         \42155_nGbbde , \42156_nGbbdf , \42157_nGbbe0 , \42158_nGbbe1 , \42159_nGbbe2 , \42160_nGbbe3 , \42161_nGbbe4 , \42162_nGbbe5 , \42163_nGbbe6 , \42164_nGbbe7 ,
         \42165_nGbbe8 , \42166_nGbbe9 , \42167_nGbbea , \42168_nGbbeb , \42169_nGbbec , \42170 , \42171_nGbbed , \42172_nGbbee , \42173_nGbbef , \42174_nGbbf0 ,
         \42175_nGbbf1 , \42176_nGbbf2 , \42177_nGbbf3 , \42178_nGbbf4 , \42179_nGbbf5 , \42180_nGbbf6 , \42181_nGbbf7 , \42182_nGbbf8 , \42183_nGbbf9 , \42184_nGbbfa ,
         \42185_nGbbfb , \42186_nGbbfc , \42187_nGbbfd , \42188_nGbbfe , \42189_nGbbff , \42190_nGbc00 , \42191_nGbc01 , \42192_nGbc02 , \42193_nGbc03 , \42194_nGbc04 ,
         \42195_nGbc05 , \42196_nGbc06 , \42197_nGbc07 , \42198_nGbc08 , \42199_nGbc09 , \42200_nGbc0a , \42201_nGbc0b , \42202_nGbc0c , \42203_nGbc0d , \42204_nGbc0e ,
         \42205_nGbc0f , \42206_nGbc10 , \42207_nGbc11 , \42208_nGbc12 , \42209_nGbc13 , \42210_nGbc14 , \42211_nGbc15 , \42212_nGbc16 , \42213_nGbc17 , \42214_nGbc18 ,
         \42215_nGbc19 , \42216_nGbc1a , \42217_nGbc1b , \42218_nGbc1c , \42219 , \42220_nGbc1d , \42221_nGbc1e , \42222_nGbc1f , \42223_nGbc20 , \42224_nGbc21 ,
         \42225_nGbc22 , \42226_nGbc23 , \42227_nGbc24 , \42228_nGbc25 , \42229_nGbc26 , \42230_nGbc27 , \42231_nGbc28 , \42232_nGbc29 , \42233_nGbc2a , \42234_nGbc2b ,
         \42235_nGbc2c , \42236_nGbc2d , \42237_nGbc2e , \42238_nGbc2f , \42239_nGbc30 , \42240_nGbc31 , \42241_nGbc32 , \42242_nGbc33 , \42243_nGbc34 , \42244_nGbc35 ,
         \42245_nGbc36 , \42246_nGbc37 , \42247_nGbc38 , \42248_nGbc39 , \42249_nGbc3a , \42250_nGbc3b , \42251_nGbc3c , \42252_nGbc3d , \42253_nGbc3e , \42254_nGbc3f ,
         \42255_nGbc40 , \42256_nGbc41 , \42257_nGbc42 , \42258_nGbc43 , \42259_nGbc44 , \42260_nGbc45 , \42261_nGbc46 , \42262_nGbc47 , \42263_nGbc48 , \42264_nGbc49 ,
         \42265_nGbc4a , \42266_nGbc4b , \42267_nGbc4c , \42268_nGbc4d , \42269_nGbc4e , \42270_nGbc4f , \42271_nGbc50 , \42272_nGbc51 , \42273_nGbc52 , \42274_nGbc53 ,
         \42275_nGbc54 , \42276_nGbc55 , \42277_nGbc56 , \42278_nGbc57 , \42279_nGbc58 , \42280_nGbc59 , \42281_nGbc5a , \42282_nGbc5b , \42283_nGbc5c , \42284_nGbc5d ,
         \42285_nGbc5e , \42286_nGbc5f , \42287_nGbc60 , \42288_nGbc61 , \42289_nGbc62 , \42290_nGbc63 , \42291_nGbc64 , \42292_nGbc65 , \42293_nGbc66 , \42294_nGbc67 ,
         \42295_nGbc68 , \42296_nGbc69 , \42297_nGbc6a , \42298_nGbc6b , \42299_nGbc6c , \42300_nGbc6d , \42301_nGbc6e , \42302_nGbc6f , \42303_nGbc70 , \42304_nGbc71 ,
         \42305_nGbc72 , \42306_nGbc73 , \42307_nGbc74 , \42308_nGbc75 , \42309_nGbc76 , \42310_nGbc77 , \42311_nGbc78 , \42312_nGbc79 , \42313_nGbc7a , \42314_nGbc7b ,
         \42315_nGbc7c , \42316 , \42317 , \42318 , \42319 , \42320_nG1489b , \42321 , \42322 , \42323_nG1489e , \42324 ,
         \42325 , \42326 , \42327 , \42328 , \42329 , \42330_nG148a5 , \42331 , \42332 , \42333_nG148a6 , \42334 ,
         \42335 , \42336 , \42337 , \42338_nG148aa , \42339_nG148ab , \42340 , \42341 , \42342 , \42343_nG148af , \42344_nG148b0 ,
         \42345_nG148b1 , \42346_nG148b2 , \42347_nG148b3 , \42348 , \42349 , \42350 , \42351 , \42352 , \42353_nG148b8 , \42354_nG148b9 ,
         \42355 , \42356 , \42357 , \42358 , \42359_nG148be , \42360_nG148bf , \42361_nG148c0 , \42362_nG148c1 , \42363_nG148c2 , \42364 ,
         \42365 , \42366 , \42367 , \42368 , \42369 , \42370 , \42371 , \42372 , \42373 , \42374 ,
         \42375 , \42376 , \42377_nG14887 , \42378_nG14888 , \42379 , \42380 , \42381 , \42382 , \42383 , \42384 ,
         \42385 , \42386 , \42387 , \42388 , \42389 , \42390 , \42391 , \42392 , \42393 , \42394 ,
         \42395 , \42396 , \42397 , \42398_nG14945 , \42399 , \42400 , \42401 , \42402 , \42403 , \42404 ,
         \42405 , \42406_nG14949 , \42407 , \42408 , \42409_nG1494a , \42410 , \42411 , \42412_nG1494b , \42413 , \42414_nG1494c ,
         \42415 , \42416 , \42417 , \42418 , \42419_nG14881 , \42420_nG14882 , \42421 , \42422 , \42423 , \42424 ,
         \42425_nG14936 , \42426 , \42427 , \42428_nG1493d , \42429_nG1493e , \42430_nG1493f , \42431_nG14940 , \42432 , \42433 , \42434 ,
         \42435 , \42436_nG1487a , \42437_nG1487d , \42438 , \42439 , \42440 , \42441 , \42442_nG14926 , \42443 , \42444_nG1492a ,
         \42445_nG1492d , \42446_nG14930 , \42447_nG14932 , \42448 , \42449 , \42450 , \42451 , \42452 , \42453 , \42454 ,
         \42455 , \42456 , \42457 , \42458 , \42459 , \42460_nG149bd , \42461 , \42462 , \42463 , \42464_nG149c1 ,
         \42465 , \42466 , \42467 , \42468 , \42469 , \42470 , \42471 , \42472 , \42473 , \42474 ,
         \42475 , \42476 , \42477 , \42478 , \42479 , \42480 , \42481 , \42482 , \42483 , \42484 ,
         \42485 , \42486 , \42487 , \42488 , \42489 , \42490 , \42491 , \42492 , \42493 , \42494 ,
         \42495 , \42496 , \42497 , \42498 , \42499 , \42500 , \42501 , \42502 , \42503 , \42504_nG1a9a6 ,
         \42505 , \42506 , \42507_nG1abf3 , \42508 , \42509 , \42510_nG1abf4 , \42511 , \42512 , \42513_nG1abf5 , \42514 ,
         \42515 , \42516_nG1abef , \42517 , \42518 , \42519_nG14a2a , \42520 , \42521_nG1a98c , \42522 , \42523 , \42524_nG14a2c ,
         \42525 , \42526_nG1a98e , \42527 , \42528 , \42529_nG14a2e , \42530 , \42531_nG1a990 , \42532 , \42533 , \42534_nG14a30 ,
         \42535 , \42536_nG1a992 , \42537 , \42538 , \42539_nG14a32 , \42540 , \42541_nG1a994 , \42542 , \42543 , \42544_nG14a34 ,
         \42545 , \42546_nG1a996 , \42547 , \42548 , \42549_nG14a36 , \42550 , \42551_nG1a998 , \42552 , \42553 , \42554_nG14a28 ,
         \42555 , \42556_nG1a98a , \42557 , \42558 , \42559_nG14a20 , \42560 , \42561_nG1a982 , \42562 , \42563 , \42564_nG14a22 ,
         \42565 , \42566_nG1a984 , \42567 , \42568 , \42569_nG14a24 , \42570 , \42571_nG1a986 , \42572 , \42573 , \42574_nG14a26 ,
         \42575 , \42576_nG1a988 , \42577 , \42578 , \42579 , \42580 , \42581 , \42582_nG14ebe , \42583 , \42584 ,
         \42585 , \42586 , \42587 , \42588 , \42589 , \42590 , \42591_nG14ebf , \42592 , \42593 , \42594 ,
         \42595 , \42596_nG14ec1 , \42597 , \42598 , \42599 , \42600_nG14ec2 , \42601 , \42602_nG1ab60 , \42603 , \42604 ,
         \42605_nG14ec3 , \42606_nG14ec4 , \42607 , \42608_nG14ec5 , \42609_nG14ec6 , \42610 , \42611_nG1ab76 , \42612 , \42613 , \42614_nG14ec7 ,
         \42615_nG14ec8 , \42616 , \42617_nG14ec9 , \42618_nG14eca , \42619 , \42620_nG1ab8c , \42621 , \42622 , \42623_nG14ecb , \42624_nG14ecc ,
         \42625 , \42626_nG14ecd , \42627_nG14ece , \42628 , \42629_nG1aba2 , \42630 , \42631 , \42632_nG14ecf , \42633_nG14ed0 , \42634 ,
         \42635_nG14ed1 , \42636_nG14ed2 , \42637 , \42638_nG1abb8 , \42639 , \42640 , \42641_nG14ed3 , \42642_nG14ed4 , \42643 , \42644_nG14ed5 ,
         \42645_nG14ed6 , \42646 , \42647_nG1abce , \42648 , \42649 , \42650_nG14ed7 , \42651_nG14ed8 , \42652 , \42653_nG14ed9 , \42654_nG14eda ,
         \42655 , \42656_nG1abda , \42657 , \42658 , \42659_nG14edb , \42660_nG14edc , \42661 , \42662_nG14edd , \42663_nG14ede , \42664 ,
         \42665_nG1abdc , \42666 , \42667 , \42668_nG14edf , \42669_nG14ee0 , \42670 , \42671_nG14ee1 , \42672_nG14ee2 , \42673 , \42674_nG1abde ,
         \42675 , \42676 , \42677_nG14ee3 , \42678_nG14ee4 , \42679 , \42680_nG14ee5 , \42681_nG14ee6 , \42682 , \42683_nG1ab62 , \42684 ,
         \42685 , \42686_nG14ee7 , \42687_nG14ee8 , \42688 , \42689_nG14ee9 , \42690_nG14eea , \42691 , \42692_nG1ab64 , \42693 , \42694 ,
         \42695_nG14eeb , \42696_nG14eec , \42697 , \42698_nG14eed , \42699_nG14eee , \42700 , \42701_nG1ab66 , \42702 , \42703 , \42704_nG14eef ,
         \42705_nG14ef0 , \42706 , \42707_nG14ef1 , \42708_nG14ef2 , \42709 , \42710_nG1ab68 , \42711 , \42712 , \42713_nG14ef3 , \42714_nG14ef4 ,
         \42715 , \42716_nG14ef5 , \42717_nG14ef6 , \42718 , \42719_nG1ab6a , \42720 , \42721 , \42722_nG14ef7 , \42723_nG14ef8 , \42724 ,
         \42725_nG14ef9 , \42726_nG14efa , \42727 , \42728_nG1ab6c , \42729 , \42730 , \42731_nG14efb , \42732_nG14efc , \42733 , \42734_nG14efd ,
         \42735_nG14efe , \42736 , \42737_nG1ab6e , \42738 , \42739 , \42740_nG14eff , \42741_nG14f00 , \42742 , \42743_nG14f01 , \42744_nG14f02 ,
         \42745 , \42746_nG1ab70 , \42747 , \42748 , \42749_nG14f03 , \42750_nG14f04 , \42751 , \42752_nG14f05 , \42753_nG14f06 , \42754 ,
         \42755_nG1ab72 , \42756 , \42757 , \42758_nG14f07 , \42759_nG14f08 , \42760 , \42761_nG14f09 , \42762_nG14f0a , \42763 , \42764_nG1ab74 ,
         \42765 , \42766 , \42767_nG14f0b , \42768_nG14f0c , \42769 , \42770_nG14f0d , \42771_nG14f0e , \42772 , \42773_nG1ab78 , \42774 ,
         \42775 , \42776_nG14f0f , \42777_nG14f10 , \42778 , \42779_nG14f11 , \42780_nG14f12 , \42781 , \42782_nG1ab7a , \42783 , \42784 ,
         \42785_nG14f13 , \42786_nG14f14 , \42787 , \42788_nG14f15 , \42789_nG14f16 , \42790 , \42791_nG1ab7c , \42792 , \42793 , \42794_nG14f17 ,
         \42795_nG14f18 , \42796 , \42797_nG14f19 , \42798_nG14f1a , \42799 , \42800_nG1ab7e , \42801 , \42802 , \42803_nG14f1b , \42804_nG14f1c ,
         \42805 , \42806_nG14f1d , \42807_nG14f1e , \42808 , \42809_nG1ab80 , \42810 , \42811 , \42812_nG14f1f , \42813_nG14f20 , \42814 ,
         \42815_nG14f21 , \42816_nG14f22 , \42817 , \42818_nG1ab82 , \42819 , \42820 , \42821_nG14f23 , \42822_nG14f24 , \42823 , \42824_nG14f25 ,
         \42825_nG14f26 , \42826 , \42827_nG1ab84 , \42828 , \42829 , \42830_nG14f27 , \42831_nG14f28 , \42832 , \42833_nG14f29 , \42834_nG14f2a ,
         \42835 , \42836_nG1ab86 , \42837 , \42838 , \42839_nG14f2b , \42840_nG14f2c , \42841 , \42842_nG14f2d , \42843_nG14f2e , \42844 ,
         \42845_nG1ab88 , \42846 , \42847 , \42848_nG14f2f , \42849_nG14f30 , \42850 , \42851_nG14f31 , \42852_nG14f32 , \42853 , \42854_nG1ab8a ,
         \42855 , \42856 , \42857_nG14f33 , \42858_nG14f34 , \42859 , \42860_nG14f35 , \42861_nG14f36 , \42862 , \42863_nG1ab8e , \42864 ,
         \42865 , \42866_nG14f37 , \42867_nG14f38 , \42868 , \42869_nG14f39 , \42870_nG14f3a , \42871 , \42872_nG1ab90 , \42873 , \42874 ,
         \42875_nG14f3b , \42876_nG14f3c , \42877 , \42878_nG14f3d , \42879_nG14f3e , \42880 , \42881_nG1ab92 , \42882 , \42883 , \42884_nG14f3f ,
         \42885_nG14f40 , \42886 , \42887_nG14f41 , \42888_nG14f42 , \42889 , \42890_nG1ab94 , \42891 , \42892 , \42893_nG14f43 , \42894_nG14f44 ,
         \42895 , \42896_nG14f45 , \42897_nG14f46 , \42898 , \42899_nG1ab96 , \42900 , \42901 , \42902_nG14f47 , \42903_nG14f48 , \42904 ,
         \42905_nG14f49 , \42906_nG14f4a , \42907 , \42908_nG1ab98 , \42909 , \42910 , \42911_nG14f4b , \42912_nG14f4c , \42913 , \42914_nG14f4d ,
         \42915_nG14f4e , \42916 , \42917_nG1ab9a , \42918 , \42919 , \42920_nG14f4f , \42921_nG14f50 , \42922 , \42923_nG14f51 , \42924_nG14f52 ,
         \42925 , \42926_nG1ab9c , \42927 , \42928 , \42929_nG14f53 , \42930_nG14f54 , \42931 , \42932_nG14f55 , \42933_nG14f56 , \42934 ,
         \42935_nG1ab9e , \42936 , \42937 , \42938_nG14f57 , \42939_nG14f58 , \42940 , \42941_nG14f59 , \42942_nG14f5a , \42943 , \42944_nG1aba0 ,
         \42945 , \42946 , \42947_nG14f5b , \42948_nG14f5c , \42949 , \42950_nG14f5d , \42951_nG14f5e , \42952 , \42953_nG1aba4 , \42954 ,
         \42955 , \42956_nG14f5f , \42957_nG14f60 , \42958 , \42959_nG14f61 , \42960_nG14f62 , \42961 , \42962_nG1aba6 , \42963 , \42964 ,
         \42965_nG14f63 , \42966_nG14f64 , \42967 , \42968_nG14f65 , \42969_nG14f66 , \42970 , \42971_nG1aba8 , \42972 , \42973 , \42974_nG14f67 ,
         \42975_nG14f68 , \42976 , \42977_nG14f69 , \42978_nG14f6a , \42979 , \42980_nG1abaa , \42981 , \42982 , \42983_nG14f6b , \42984_nG14f6c ,
         \42985 , \42986_nG14f6d , \42987_nG14f6e , \42988 , \42989_nG1abac , \42990 , \42991 , \42992_nG14f6f , \42993_nG14f70 , \42994 ,
         \42995_nG14f71 , \42996_nG14f72 , \42997 , \42998_nG1abae , \42999 , \43000 , \43001_nG14f73 , \43002_nG14f74 , \43003 , \43004_nG14f75 ,
         \43005_nG14f76 , \43006 , \43007_nG1abb0 , \43008 , \43009 , \43010_nG14f77 , \43011_nG14f78 , \43012 , \43013_nG14f79 , \43014_nG14f7a ,
         \43015 , \43016_nG1abb2 , \43017 , \43018 , \43019_nG14f7b , \43020_nG14f7c , \43021 , \43022_nG14f7d , \43023_nG14f7e , \43024 ,
         \43025_nG1abb4 , \43026 , \43027 , \43028_nG14f7f , \43029_nG14f80 , \43030 , \43031_nG14f81 , \43032_nG14f82 , \43033 , \43034_nG1abb6 ,
         \43035 , \43036 , \43037_nG14f83 , \43038_nG14f84 , \43039 , \43040_nG14f85 , \43041_nG14f86 , \43042 , \43043_nG1abba , \43044 ,
         \43045 , \43046_nG14f87 , \43047_nG14f88 , \43048 , \43049_nG14f89 , \43050_nG14f8a , \43051 , \43052_nG1abbc , \43053 , \43054 ,
         \43055_nG14f8b , \43056_nG14f8c , \43057 , \43058_nG14f8d , \43059_nG14f8e , \43060 , \43061_nG1abbe , \43062 , \43063 , \43064_nG14f8f ,
         \43065_nG14f90 , \43066 , \43067_nG14f91 , \43068_nG14f92 , \43069 , \43070_nG1abc0 , \43071 , \43072 , \43073_nG14f93 , \43074_nG14f94 ,
         \43075 , \43076_nG14f95 , \43077_nG14f96 , \43078 , \43079_nG1abc2 , \43080 , \43081 , \43082_nG14f97 , \43083_nG14f98 , \43084 ,
         \43085_nG14f99 , \43086_nG14f9a , \43087 , \43088_nG1abc4 , \43089 , \43090 , \43091_nG14f9b , \43092_nG14f9c , \43093 , \43094_nG14f9d ,
         \43095_nG14f9e , \43096 , \43097_nG1abc6 , \43098 , \43099 , \43100_nG14f9f , \43101_nG14fa0 , \43102 , \43103_nG14fa1 , \43104_nG14fa2 ,
         \43105 , \43106_nG1abc8 , \43107 , \43108 , \43109_nG14fa3 , \43110_nG14fa4 , \43111 , \43112_nG14fa5 , \43113_nG14fa6 , \43114 ,
         \43115_nG1abca , \43116 , \43117 , \43118_nG14fa7 , \43119_nG14fa8 , \43120 , \43121_nG14fa9 , \43122_nG14faa , \43123 , \43124_nG1abcc ,
         \43125 , \43126 , \43127_nG14fab , \43128_nG14fac , \43129 , \43130_nG14fad , \43131_nG14fae , \43132 , \43133_nG1abd0 , \43134 ,
         \43135 , \43136_nG14faf , \43137_nG14fb0 , \43138 , \43139_nG14fb1 , \43140_nG14fb2 , \43141 , \43142_nG1abd2 , \43143 , \43144 ,
         \43145_nG14fb3 , \43146_nG14fb4 , \43147 , \43148_nG14fb5 , \43149_nG14fb6 , \43150 , \43151_nG1abd4 , \43152 , \43153 , \43154_nG14fb7 ,
         \43155_nG14fb8 , \43156 , \43157_nG14fb9 , \43158_nG14fba , \43159 , \43160_nG1abd6 , \43161 , \43162 , \43163_nG14fbb , \43164_nG14fbc ,
         \43165 , \43166_nG14fbd , \43167_nG14fbe , \43168 , \43169_nG1abd8 , \43170 , \43171 , \43172 , \43173_nG14dbd , \43174_nG14dbe ,
         \43175 , \43176 , \43177_nG14dc0 , \43178_nG14dc1 , \43179 , \43180_nG1aae0 , \43181 , \43182_nG14dc2 , \43183_nG14dc3 , \43184_nG14dc4 ,
         \43185_nG14dc5 , \43186 , \43187_nG1aaf6 , \43188 , \43189_nG14dc6 , \43190_nG14dc7 , \43191_nG14dc8 , \43192_nG14dc9 , \43193 , \43194_nG1ab0c ,
         \43195 , \43196_nG14dca , \43197_nG14dcb , \43198_nG14dcc , \43199_nG14dcd , \43200 , \43201_nG1ab22 , \43202 , \43203_nG14dce , \43204_nG14dcf ,
         \43205_nG14dd0 , \43206_nG14dd1 , \43207 , \43208_nG1ab38 , \43209 , \43210_nG14dd2 , \43211_nG14dd3 , \43212_nG14dd4 , \43213_nG14dd5 , \43214 ,
         \43215_nG1ab4e , \43216 , \43217_nG14dd6 , \43218_nG14dd7 , \43219_nG14dd8 , \43220_nG14dd9 , \43221 , \43222_nG1ab5a , \43223 , \43224_nG14dda ,
         \43225_nG14ddb , \43226_nG14ddc , \43227_nG14ddd , \43228 , \43229_nG1ab5c , \43230 , \43231_nG14dde , \43232_nG14ddf , \43233_nG14de0 , \43234_nG14de1 ,
         \43235 , \43236_nG1ab5e , \43237 , \43238_nG14de2 , \43239_nG14de3 , \43240_nG14de4 , \43241_nG14de5 , \43242 , \43243_nG1aae2 , \43244 ,
         \43245_nG14de6 , \43246_nG14de7 , \43247_nG14de8 , \43248_nG14de9 , \43249 , \43250_nG1aae4 , \43251 , \43252_nG14dea , \43253_nG14deb , \43254_nG14dec ,
         \43255_nG14ded , \43256 , \43257_nG1aae6 , \43258 , \43259_nG14dee , \43260_nG14def , \43261_nG14df0 , \43262_nG14df1 , \43263 , \43264_nG1aae8 ,
         \43265 , \43266_nG14df2 , \43267_nG14df3 , \43268_nG14df4 , \43269_nG14df5 , \43270 , \43271_nG1aaea , \43272 , \43273_nG14df6 , \43274_nG14df7 ,
         \43275_nG14df8 , \43276_nG14df9 , \43277 , \43278_nG1aaec , \43279 , \43280_nG14dfa , \43281_nG14dfb , \43282_nG14dfc , \43283_nG14dfd , \43284 ,
         \43285_nG1aaee , \43286 , \43287_nG14dfe , \43288_nG14dff , \43289_nG14e00 , \43290_nG14e01 , \43291 , \43292_nG1aaf0 , \43293 , \43294_nG14e02 ,
         \43295_nG14e03 , \43296_nG14e04 , \43297_nG14e05 , \43298 , \43299_nG1aaf2 , \43300 , \43301_nG14e06 , \43302_nG14e07 , \43303_nG14e08 , \43304_nG14e09 ,
         \43305 , \43306_nG1aaf4 , \43307 , \43308_nG14e0a , \43309_nG14e0b , \43310_nG14e0c , \43311_nG14e0d , \43312 , \43313_nG1aaf8 , \43314 ,
         \43315_nG14e0e , \43316_nG14e0f , \43317_nG14e10 , \43318_nG14e11 , \43319 , \43320_nG1aafa , \43321 , \43322_nG14e12 , \43323_nG14e13 , \43324_nG14e14 ,
         \43325_nG14e15 , \43326 , \43327_nG1aafc , \43328 , \43329_nG14e16 , \43330_nG14e17 , \43331_nG14e18 , \43332_nG14e19 , \43333 , \43334_nG1aafe ,
         \43335 , \43336_nG14e1a , \43337_nG14e1b , \43338_nG14e1c , \43339_nG14e1d , \43340 , \43341_nG1ab00 , \43342 , \43343_nG14e1e , \43344_nG14e1f ,
         \43345_nG14e20 , \43346_nG14e21 , \43347 , \43348_nG1ab02 , \43349 , \43350_nG14e22 , \43351_nG14e23 , \43352_nG14e24 , \43353_nG14e25 , \43354 ,
         \43355_nG1ab04 , \43356 , \43357_nG14e26 , \43358_nG14e27 , \43359_nG14e28 , \43360_nG14e29 , \43361 , \43362_nG1ab06 , \43363 , \43364_nG14e2a ,
         \43365_nG14e2b , \43366_nG14e2c , \43367_nG14e2d , \43368 , \43369_nG1ab08 , \43370 , \43371_nG14e2e , \43372_nG14e2f , \43373_nG14e30 , \43374_nG14e31 ,
         \43375 , \43376_nG1ab0a , \43377 , \43378_nG14e32 , \43379_nG14e33 , \43380_nG14e34 , \43381_nG14e35 , \43382 , \43383_nG1ab0e , \43384 ,
         \43385_nG14e36 , \43386_nG14e37 , \43387_nG14e38 , \43388_nG14e39 , \43389 , \43390_nG1ab10 , \43391 , \43392_nG14e3a , \43393_nG14e3b , \43394_nG14e3c ,
         \43395_nG14e3d , \43396 , \43397_nG1ab12 , \43398 , \43399_nG14e3e , \43400_nG14e3f , \43401_nG14e40 , \43402_nG14e41 , \43403 , \43404_nG1ab14 ,
         \43405 , \43406_nG14e42 , \43407_nG14e43 , \43408_nG14e44 , \43409_nG14e45 , \43410 , \43411_nG1ab16 , \43412 , \43413_nG14e46 , \43414_nG14e47 ,
         \43415_nG14e48 , \43416_nG14e49 , \43417 , \43418_nG1ab18 , \43419 , \43420_nG14e4a , \43421_nG14e4b , \43422_nG14e4c , \43423_nG14e4d , \43424 ,
         \43425_nG1ab1a , \43426 , \43427_nG14e4e , \43428_nG14e4f , \43429_nG14e50 , \43430_nG14e51 , \43431 , \43432_nG1ab1c , \43433 , \43434_nG14e52 ,
         \43435_nG14e53 , \43436_nG14e54 , \43437_nG14e55 , \43438 , \43439_nG1ab1e , \43440 , \43441_nG14e56 , \43442_nG14e57 , \43443_nG14e58 , \43444_nG14e59 ,
         \43445 , \43446_nG1ab20 , \43447 , \43448_nG14e5a , \43449_nG14e5b , \43450_nG14e5c , \43451_nG14e5d , \43452 , \43453_nG1ab24 , \43454 ,
         \43455_nG14e5e , \43456_nG14e5f , \43457_nG14e60 , \43458_nG14e61 , \43459 , \43460_nG1ab26 , \43461 , \43462_nG14e62 , \43463_nG14e63 , \43464_nG14e64 ,
         \43465_nG14e65 , \43466 , \43467_nG1ab28 , \43468 , \43469_nG14e66 , \43470_nG14e67 , \43471_nG14e68 , \43472_nG14e69 , \43473 , \43474_nG1ab2a ,
         \43475 , \43476_nG14e6a , \43477_nG14e6b , \43478_nG14e6c , \43479_nG14e6d , \43480 , \43481_nG1ab2c , \43482 , \43483_nG14e6e , \43484_nG14e6f ,
         \43485_nG14e70 , \43486_nG14e71 , \43487 , \43488_nG1ab2e , \43489 , \43490_nG14e72 , \43491_nG14e73 , \43492_nG14e74 , \43493_nG14e75 , \43494 ,
         \43495_nG1ab30 , \43496 , \43497_nG14e76 , \43498_nG14e77 , \43499_nG14e78 , \43500_nG14e79 , \43501 , \43502_nG1ab32 , \43503 , \43504_nG14e7a ,
         \43505_nG14e7b , \43506_nG14e7c , \43507_nG14e7d , \43508 , \43509_nG1ab34 , \43510 , \43511_nG14e7e , \43512_nG14e7f , \43513_nG14e80 , \43514_nG14e81 ,
         \43515 , \43516_nG1ab36 , \43517 , \43518_nG14e82 , \43519_nG14e83 , \43520_nG14e84 , \43521_nG14e85 , \43522 , \43523_nG1ab3a , \43524 ,
         \43525_nG14e86 , \43526_nG14e87 , \43527_nG14e88 , \43528_nG14e89 , \43529 , \43530_nG1ab3c , \43531 , \43532_nG14e8a , \43533_nG14e8b , \43534_nG14e8c ,
         \43535_nG14e8d , \43536 , \43537_nG1ab3e , \43538 , \43539_nG14e8e , \43540_nG14e8f , \43541_nG14e90 , \43542_nG14e91 , \43543 , \43544_nG1ab40 ,
         \43545 , \43546_nG14e92 , \43547_nG14e93 , \43548_nG14e94 , \43549_nG14e95 , \43550 , \43551_nG1ab42 , \43552 , \43553_nG14e96 , \43554_nG14e97 ,
         \43555_nG14e98 , \43556_nG14e99 , \43557 , \43558_nG1ab44 , \43559 , \43560_nG14e9a , \43561_nG14e9b , \43562_nG14e9c , \43563_nG14e9d , \43564 ,
         \43565_nG1ab46 , \43566 , \43567_nG14e9e , \43568_nG14e9f , \43569_nG14ea0 , \43570_nG14ea1 , \43571 , \43572_nG1ab48 , \43573 , \43574_nG14ea2 ,
         \43575_nG14ea3 , \43576_nG14ea4 , \43577_nG14ea5 , \43578 , \43579_nG1ab4a , \43580 , \43581_nG14ea6 , \43582_nG14ea7 , \43583_nG14ea8 , \43584_nG14ea9 ,
         \43585 , \43586_nG1ab4c , \43587 , \43588_nG14eaa , \43589_nG14eab , \43590_nG14eac , \43591_nG14ead , \43592 , \43593_nG1ab50 , \43594 ,
         \43595_nG14eae , \43596_nG14eaf , \43597_nG14eb0 , \43598_nG14eb1 , \43599 , \43600_nG1ab52 , \43601 , \43602_nG14eb2 , \43603_nG14eb3 , \43604_nG14eb4 ,
         \43605_nG14eb5 , \43606 , \43607_nG1ab54 , \43608 , \43609_nG14eb6 , \43610_nG14eb7 , \43611_nG14eb8 , \43612_nG14eb9 , \43613 , \43614_nG1ab56 ,
         \43615 , \43616_nG14eba , \43617_nG14ebb , \43618_nG14ebc , \43619_nG14ebd , \43620 , \43621_nG1ab58 , \43622 , \43623 , \43624_nG14cbb ,
         \43625_nG14cbc , \43626 , \43627_nG14cbf , \43628_nG14cc0 , \43629 , \43630_nG1aa60 , \43631 , \43632_nG14cc1 , \43633_nG14cc2 , \43634_nG14cc3 ,
         \43635_nG14cc4 , \43636 , \43637_nG1aa76 , \43638 , \43639_nG14cc5 , \43640_nG14cc6 , \43641_nG14cc7 , \43642_nG14cc8 , \43643 , \43644_nG1aa8c ,
         \43645 , \43646_nG14cc9 , \43647_nG14cca , \43648_nG14ccb , \43649_nG14ccc , \43650 , \43651_nG1aaa2 , \43652 , \43653_nG14ccd , \43654_nG14cce ,
         \43655_nG14ccf , \43656_nG14cd0 , \43657 , \43658_nG1aab8 , \43659 , \43660_nG14cd1 , \43661_nG14cd2 , \43662_nG14cd3 , \43663_nG14cd4 , \43664 ,
         \43665_nG1aace , \43666 , \43667_nG14cd5 , \43668_nG14cd6 , \43669_nG14cd7 , \43670_nG14cd8 , \43671 , \43672_nG1aada , \43673 , \43674_nG14cd9 ,
         \43675_nG14cda , \43676_nG14cdb , \43677_nG14cdc , \43678 , \43679_nG1aadc , \43680 , \43681_nG14cdd , \43682_nG14cde , \43683_nG14cdf , \43684_nG14ce0 ,
         \43685 , \43686_nG1aade , \43687 , \43688_nG14ce1 , \43689_nG14ce2 , \43690_nG14ce3 , \43691_nG14ce4 , \43692 , \43693_nG1aa62 , \43694 ,
         \43695_nG14ce5 , \43696_nG14ce6 , \43697_nG14ce7 , \43698_nG14ce8 , \43699 , \43700_nG1aa64 , \43701 , \43702_nG14ce9 , \43703_nG14cea , \43704_nG14ceb ,
         \43705_nG14cec , \43706 , \43707_nG1aa66 , \43708 , \43709_nG14ced , \43710_nG14cee , \43711_nG14cef , \43712_nG14cf0 , \43713 , \43714_nG1aa68 ,
         \43715 , \43716_nG14cf1 , \43717_nG14cf2 , \43718_nG14cf3 , \43719_nG14cf4 , \43720 , \43721_nG1aa6a , \43722 , \43723_nG14cf5 , \43724_nG14cf6 ,
         \43725_nG14cf7 , \43726_nG14cf8 , \43727 , \43728_nG1aa6c , \43729 , \43730_nG14cf9 , \43731_nG14cfa , \43732_nG14cfb , \43733_nG14cfc , \43734 ,
         \43735_nG1aa6e , \43736 , \43737_nG14cfd , \43738_nG14cfe , \43739_nG14cff , \43740_nG14d00 , \43741 , \43742_nG1aa70 , \43743 , \43744_nG14d01 ,
         \43745_nG14d02 , \43746_nG14d03 , \43747_nG14d04 , \43748 , \43749_nG1aa72 , \43750 , \43751_nG14d05 , \43752_nG14d06 , \43753_nG14d07 , \43754_nG14d08 ,
         \43755 , \43756_nG1aa74 , \43757 , \43758_nG14d09 , \43759_nG14d0a , \43760_nG14d0b , \43761_nG14d0c , \43762 , \43763_nG1aa78 , \43764 ,
         \43765_nG14d0d , \43766_nG14d0e , \43767_nG14d0f , \43768_nG14d10 , \43769 , \43770_nG1aa7a , \43771 , \43772_nG14d11 , \43773_nG14d12 , \43774_nG14d13 ,
         \43775_nG14d14 , \43776 , \43777_nG1aa7c , \43778 , \43779_nG14d15 , \43780_nG14d16 , \43781_nG14d17 , \43782_nG14d18 , \43783 , \43784_nG1aa7e ,
         \43785 , \43786_nG14d19 , \43787_nG14d1a , \43788_nG14d1b , \43789_nG14d1c , \43790 , \43791_nG1aa80 , \43792 , \43793_nG14d1d , \43794_nG14d1e ,
         \43795_nG14d1f , \43796_nG14d20 , \43797 , \43798_nG1aa82 , \43799 , \43800_nG14d21 , \43801_nG14d22 , \43802_nG14d23 , \43803_nG14d24 , \43804 ,
         \43805_nG1aa84 , \43806 , \43807_nG14d25 , \43808_nG14d26 , \43809_nG14d27 , \43810_nG14d28 , \43811 , \43812_nG1aa86 , \43813 , \43814_nG14d29 ,
         \43815_nG14d2a , \43816_nG14d2b , \43817_nG14d2c , \43818 , \43819_nG1aa88 , \43820 , \43821_nG14d2d , \43822_nG14d2e , \43823_nG14d2f , \43824_nG14d30 ,
         \43825 , \43826_nG1aa8a , \43827 , \43828_nG14d31 , \43829_nG14d32 , \43830_nG14d33 , \43831_nG14d34 , \43832 , \43833_nG1aa8e , \43834 ,
         \43835_nG14d35 , \43836_nG14d36 , \43837_nG14d37 , \43838_nG14d38 , \43839 , \43840_nG1aa90 , \43841 , \43842_nG14d39 , \43843_nG14d3a , \43844_nG14d3b ,
         \43845_nG14d3c , \43846 , \43847_nG1aa92 , \43848 , \43849_nG14d3d , \43850_nG14d3e , \43851_nG14d3f , \43852_nG14d40 , \43853 , \43854_nG1aa94 ,
         \43855 , \43856_nG14d41 , \43857_nG14d42 , \43858_nG14d43 , \43859_nG14d44 , \43860 , \43861_nG1aa96 , \43862 , \43863_nG14d45 , \43864_nG14d46 ,
         \43865_nG14d47 , \43866_nG14d48 , \43867 , \43868_nG1aa98 , \43869 , \43870_nG14d49 , \43871_nG14d4a , \43872_nG14d4b , \43873_nG14d4c , \43874 ,
         \43875_nG1aa9a , \43876 , \43877_nG14d4d , \43878_nG14d4e , \43879_nG14d4f , \43880_nG14d50 , \43881 , \43882_nG1aa9c , \43883 , \43884_nG14d51 ,
         \43885_nG14d52 , \43886_nG14d53 , \43887_nG14d54 , \43888 , \43889_nG1aa9e , \43890 , \43891_nG14d55 , \43892_nG14d56 , \43893_nG14d57 , \43894_nG14d58 ,
         \43895 , \43896_nG1aaa0 , \43897 , \43898_nG14d59 , \43899_nG14d5a , \43900_nG14d5b , \43901_nG14d5c , \43902 , \43903_nG1aaa4 , \43904 ,
         \43905_nG14d5d , \43906_nG14d5e , \43907_nG14d5f , \43908_nG14d60 , \43909 , \43910_nG1aaa6 , \43911 , \43912_nG14d61 , \43913_nG14d62 , \43914_nG14d63 ,
         \43915_nG14d64 , \43916 , \43917_nG1aaa8 , \43918 , \43919_nG14d65 , \43920_nG14d66 , \43921_nG14d67 , \43922_nG14d68 , \43923 , \43924_nG1aaaa ,
         \43925 , \43926_nG14d69 , \43927_nG14d6a , \43928_nG14d6b , \43929_nG14d6c , \43930 , \43931_nG1aaac , \43932 , \43933_nG14d6d , \43934_nG14d6e ,
         \43935_nG14d6f , \43936_nG14d70 , \43937 , \43938_nG1aaae , \43939 , \43940_nG14d71 , \43941_nG14d72 , \43942_nG14d73 , \43943_nG14d74 , \43944 ,
         \43945_nG1aab0 , \43946 , \43947_nG14d75 , \43948_nG14d76 , \43949_nG14d77 , \43950_nG14d78 , \43951 , \43952_nG1aab2 , \43953 , \43954_nG14d79 ,
         \43955_nG14d7a , \43956_nG14d7b , \43957_nG14d7c , \43958 , \43959_nG1aab4 , \43960 , \43961_nG14d7d , \43962_nG14d7e , \43963_nG14d7f , \43964_nG14d80 ,
         \43965 , \43966_nG1aab6 , \43967 , \43968_nG14d81 , \43969_nG14d82 , \43970_nG14d83 , \43971_nG14d84 , \43972 , \43973_nG1aaba , \43974 ,
         \43975_nG14d85 , \43976_nG14d86 , \43977_nG14d87 , \43978_nG14d88 , \43979 , \43980_nG1aabc , \43981 , \43982_nG14d89 , \43983_nG14d8a , \43984_nG14d8b ,
         \43985_nG14d8c , \43986 , \43987_nG1aabe , \43988 , \43989_nG14d8d , \43990_nG14d8e , \43991_nG14d8f , \43992_nG14d90 , \43993 , \43994_nG1aac0 ,
         \43995 , \43996_nG14d91 , \43997_nG14d92 , \43998_nG14d93 , \43999_nG14d94 , \44000 , \44001_nG1aac2 , \44002 , \44003_nG14d95 , \44004_nG14d96 ,
         \44005_nG14d97 , \44006_nG14d98 , \44007 , \44008_nG1aac4 , \44009 , \44010_nG14d99 , \44011_nG14d9a , \44012_nG14d9b , \44013_nG14d9c , \44014 ,
         \44015_nG1aac6 , \44016 , \44017_nG14d9d , \44018_nG14d9e , \44019_nG14d9f , \44020_nG14da0 , \44021 , \44022_nG1aac8 , \44023 , \44024_nG14da1 ,
         \44025_nG14da2 , \44026_nG14da3 , \44027_nG14da4 , \44028 , \44029_nG1aaca , \44030 , \44031_nG14da5 , \44032_nG14da6 , \44033_nG14da7 , \44034_nG14da8 ,
         \44035 , \44036_nG1aacc , \44037 , \44038_nG14da9 , \44039_nG14daa , \44040_nG14dab , \44041_nG14dac , \44042 , \44043_nG1aad0 , \44044 ,
         \44045_nG14dad , \44046_nG14dae , \44047_nG14daf , \44048_nG14db0 , \44049 , \44050_nG1aad2 , \44051 , \44052_nG14db1 , \44053_nG14db2 , \44054_nG14db3 ,
         \44055_nG14db4 , \44056 , \44057_nG1aad4 , \44058 , \44059_nG14db5 , \44060_nG14db6 , \44061_nG14db7 , \44062_nG14db8 , \44063 , \44064_nG1aad6 ,
         \44065 , \44066_nG14db9 , \44067_nG14dba , \44068_nG14dbb , \44069_nG14dbc , \44070 , \44071_nG1aad8 , \44072 , \44073 , \44074_nG14b39 ,
         \44075_nG14b3a , \44076 , \44077_nG14b3f , \44078_nG14b40 , \44079 , \44080_nG1a9e0 , \44081 , \44082_nG14b42 , \44083_nG14b43 , \44084_nG14b45 ,
         \44085_nG14b46 , \44086 , \44087_nG1a9f6 , \44088 , \44089_nG14b48 , \44090_nG14b49 , \44091_nG14b4b , \44092_nG14b4c , \44093 , \44094_nG1aa0c ,
         \44095 , \44096_nG14b4e , \44097_nG14b4f , \44098_nG14b51 , \44099_nG14b52 , \44100 , \44101_nG1aa22 , \44102 , \44103_nG14b54 , \44104_nG14b55 ,
         \44105_nG14b57 , \44106_nG14b58 , \44107 , \44108_nG1aa38 , \44109 , \44110_nG14b5a , \44111_nG14b5b , \44112_nG14b5d , \44113_nG14b5e , \44114 ,
         \44115_nG1aa4e , \44116 , \44117_nG14b60 , \44118_nG14b61 , \44119_nG14b63 , \44120_nG14b64 , \44121 , \44122_nG1aa5a , \44123 , \44124_nG14b66 ,
         \44125_nG14b67 , \44126_nG14b69 , \44127_nG14b6a , \44128 , \44129_nG1aa5c , \44130 , \44131_nG14b6c , \44132_nG14b6d , \44133_nG14b6f , \44134_nG14b70 ,
         \44135 , \44136_nG1aa5e , \44137 , \44138_nG14b72 , \44139_nG14b73 , \44140_nG14b75 , \44141_nG14b76 , \44142 , \44143_nG1a9e2 , \44144 ,
         \44145_nG14b78 , \44146_nG14b79 , \44147_nG14b7b , \44148_nG14b7c , \44149 , \44150_nG1a9e4 , \44151 , \44152_nG14b7e , \44153_nG14b7f , \44154_nG14b81 ,
         \44155_nG14b82 , \44156 , \44157_nG1a9e6 , \44158 , \44159_nG14b84 , \44160_nG14b85 , \44161_nG14b87 , \44162_nG14b88 , \44163 , \44164_nG1a9e8 ,
         \44165 , \44166_nG14b8a , \44167_nG14b8b , \44168_nG14b8d , \44169_nG14b8e , \44170 , \44171_nG1a9ea , \44172 , \44173_nG14b90 , \44174_nG14b91 ,
         \44175_nG14b93 , \44176_nG14b94 , \44177 , \44178_nG1a9ec , \44179 , \44180_nG14b96 , \44181_nG14b97 , \44182_nG14b99 , \44183_nG14b9a , \44184 ,
         \44185_nG1a9ee , \44186 , \44187_nG14b9c , \44188_nG14b9d , \44189_nG14b9f , \44190_nG14ba0 , \44191 , \44192_nG1a9f0 , \44193 , \44194_nG14ba2 ,
         \44195_nG14ba3 , \44196_nG14ba5 , \44197_nG14ba6 , \44198 , \44199_nG1a9f2 , \44200 , \44201_nG14ba8 , \44202_nG14ba9 , \44203_nG14bab , \44204_nG14bac ,
         \44205 , \44206_nG1a9f4 , \44207 , \44208_nG14bae , \44209_nG14baf , \44210_nG14bb1 , \44211_nG14bb2 , \44212 , \44213_nG1a9f8 , \44214 ,
         \44215_nG14bb4 , \44216_nG14bb5 , \44217_nG14bb7 , \44218_nG14bb8 , \44219 , \44220_nG1a9fa , \44221 , \44222_nG14bba , \44223_nG14bbb , \44224_nG14bbd ,
         \44225_nG14bbe , \44226 , \44227_nG1a9fc , \44228 , \44229_nG14bc0 , \44230_nG14bc1 , \44231_nG14bc3 , \44232_nG14bc4 , \44233 , \44234_nG1a9fe ,
         \44235 , \44236_nG14bc6 , \44237_nG14bc7 , \44238_nG14bc9 , \44239_nG14bca , \44240 , \44241_nG1aa00 , \44242 , \44243_nG14bcc , \44244_nG14bcd ,
         \44245_nG14bcf , \44246_nG14bd0 , \44247 , \44248_nG1aa02 , \44249 , \44250_nG14bd2 , \44251_nG14bd3 , \44252_nG14bd5 , \44253_nG14bd6 , \44254 ,
         \44255_nG1aa04 , \44256 , \44257_nG14bd8 , \44258_nG14bd9 , \44259_nG14bdb , \44260_nG14bdc , \44261 , \44262_nG1aa06 , \44263 , \44264_nG14bde ,
         \44265_nG14bdf , \44266_nG14be1 , \44267_nG14be2 , \44268 , \44269_nG1aa08 , \44270 , \44271_nG14be4 , \44272_nG14be5 , \44273_nG14be7 , \44274_nG14be8 ,
         \44275 , \44276_nG1aa0a , \44277 , \44278_nG14bea , \44279_nG14beb , \44280_nG14bed , \44281_nG14bee , \44282 , \44283_nG1aa0e , \44284 ,
         \44285_nG14bf0 , \44286_nG14bf1 , \44287_nG14bf3 , \44288_nG14bf4 , \44289 , \44290_nG1aa10 , \44291 , \44292_nG14bf6 , \44293_nG14bf7 , \44294_nG14bf9 ,
         \44295_nG14bfa , \44296 , \44297_nG1aa12 , \44298 , \44299_nG14bfc , \44300_nG14bfd , \44301_nG14bff , \44302_nG14c00 , \44303 , \44304_nG1aa14 ,
         \44305 , \44306_nG14c02 , \44307_nG14c03 , \44308_nG14c05 , \44309_nG14c06 , \44310 , \44311_nG1aa16 , \44312 , \44313_nG14c08 , \44314_nG14c09 ,
         \44315_nG14c0b , \44316_nG14c0c , \44317 , \44318_nG1aa18 , \44319 , \44320_nG14c0e , \44321_nG14c0f , \44322_nG14c11 , \44323_nG14c12 , \44324 ,
         \44325_nG1aa1a , \44326 , \44327_nG14c14 , \44328_nG14c15 , \44329_nG14c17 , \44330_nG14c18 , \44331 , \44332_nG1aa1c , \44333 , \44334_nG14c1a ,
         \44335_nG14c1b , \44336_nG14c1d , \44337_nG14c1e , \44338 , \44339_nG1aa1e , \44340 , \44341_nG14c20 , \44342_nG14c21 , \44343_nG14c23 , \44344_nG14c24 ,
         \44345 , \44346_nG1aa20 , \44347 , \44348_nG14c26 , \44349_nG14c27 , \44350_nG14c29 , \44351_nG14c2a , \44352 , \44353_nG1aa24 , \44354 ,
         \44355_nG14c2c , \44356_nG14c2d , \44357_nG14c2f , \44358_nG14c30 , \44359 , \44360_nG1aa26 , \44361 , \44362_nG14c32 , \44363_nG14c33 , \44364_nG14c35 ,
         \44365_nG14c36 , \44366 , \44367_nG1aa28 , \44368 , \44369_nG14c38 , \44370_nG14c39 , \44371_nG14c3b , \44372_nG14c3c , \44373 , \44374_nG1aa2a ,
         \44375 , \44376_nG14c3e , \44377_nG14c3f , \44378_nG14c41 , \44379_nG14c42 , \44380 , \44381_nG1aa2c , \44382 , \44383_nG14c44 , \44384_nG14c45 ,
         \44385_nG14c47 , \44386_nG14c48 , \44387 , \44388_nG1aa2e , \44389 , \44390_nG14c4a , \44391_nG14c4b , \44392_nG14c4d , \44393_nG14c4e , \44394 ,
         \44395_nG1aa30 , \44396 , \44397_nG14c50 , \44398_nG14c51 , \44399_nG14c53 , \44400_nG14c54 , \44401 , \44402_nG1aa32 , \44403 , \44404_nG14c56 ,
         \44405_nG14c57 , \44406_nG14c59 , \44407_nG14c5a , \44408 , \44409_nG1aa34 , \44410 , \44411_nG14c5c , \44412_nG14c5d , \44413_nG14c5f , \44414_nG14c60 ,
         \44415 , \44416_nG1aa36 , \44417 , \44418_nG14c62 , \44419_nG14c63 , \44420_nG14c65 , \44421_nG14c66 , \44422 , \44423_nG1aa3a , \44424 ,
         \44425_nG14c68 , \44426_nG14c69 , \44427_nG14c6b , \44428_nG14c6c , \44429 , \44430_nG1aa3c , \44431 , \44432_nG14c6e , \44433_nG14c6f , \44434_nG14c71 ,
         \44435_nG14c72 , \44436 , \44437_nG1aa3e , \44438 , \44439_nG14c74 , \44440_nG14c75 , \44441_nG14c77 , \44442_nG14c78 , \44443 , \44444_nG1aa40 ,
         \44445 , \44446_nG14c7a , \44447_nG14c7b , \44448_nG14c7d , \44449_nG14c7e , \44450 , \44451_nG1aa42 , \44452 , \44453_nG14c80 , \44454_nG14c81 ,
         \44455_nG14c83 , \44456_nG14c84 , \44457 , \44458_nG1aa44 , \44459 , \44460_nG14c86 , \44461_nG14c87 , \44462_nG14c89 , \44463_nG14c8a , \44464 ,
         \44465_nG1aa46 , \44466 , \44467_nG14c8c , \44468_nG14c8d , \44469_nG14c8f , \44470_nG14c90 , \44471 , \44472_nG1aa48 , \44473 , \44474_nG14c92 ,
         \44475_nG14c93 , \44476_nG14c95 , \44477_nG14c96 , \44478 , \44479_nG1aa4a , \44480 , \44481_nG14c98 , \44482_nG14c99 , \44483_nG14c9b , \44484_nG14c9c ,
         \44485 , \44486_nG1aa4c , \44487 , \44488_nG14c9e , \44489_nG14c9f , \44490_nG14ca1 , \44491_nG14ca2 , \44492 , \44493_nG1aa50 , \44494 ,
         \44495_nG14ca4 , \44496_nG14ca5 , \44497_nG14ca7 , \44498_nG14ca8 , \44499 , \44500_nG1aa52 , \44501 , \44502_nG14caa , \44503_nG14cab , \44504_nG14cad ,
         \44505_nG14cae , \44506 , \44507_nG1aa54 , \44508 , \44509_nG14cb0 , \44510_nG14cb1 , \44511_nG14cb3 , \44512_nG14cb4 , \44513 , \44514_nG1aa56 ,
         \44515 , \44516_nG14cb6 , \44517_nG14cb7 , \44518_nG14cb9 , \44519_nG14cba , \44520 , \44521_nG1aa58 , \44522 , \44523 , \44524_nG14b0b ,
         \44525 , \44526 , \44527_nG14b0c , \44528 , \44529_nG1a9c8 , \44530 , \44531 , \44532_nG14b0d , \44533_nG14b0e , \44534 ,
         \44535_nG1a9ca , \44536 , \44537 , \44538_nG14b0f , \44539_nG14b10 , \44540 , \44541_nG1a9cc , \44542 , \44543 , \44544_nG14b11 ,
         \44545_nG14b12 , \44546 , \44547_nG1a9ce , \44548 , \44549 , \44550_nG14b13 , \44551_nG14b14 , \44552 , \44553_nG1a9d0 , \44554 ,
         \44555 , \44556_nG14b15 , \44557_nG14b16 , \44558 , \44559_nG1a9d2 , \44560 , \44561 , \44562_nG14b17 , \44563_nG14b18 , \44564 ,
         \44565_nG1a9d4 , \44566 , \44567 , \44568_nG14b19 , \44569_nG14b1a , \44570 , \44571_nG1a9d6 , \44572 , \44573_nG14afa , \44574_nG14afb ,
         \44575 , \44576_nG1a9b8 , \44577 , \44578_nG14afc , \44579_nG14afd , \44580 , \44581_nG1a9ba , \44582 , \44583_nG14afe , \44584_nG14aff ,
         \44585 , \44586_nG1a9bc , \44587 , \44588_nG14b00 , \44589_nG14b01 , \44590 , \44591_nG1a9be , \44592 , \44593_nG14b02 , \44594_nG14b03 ,
         \44595 , \44596_nG1a9c0 , \44597 , \44598_nG14b04 , \44599_nG14b05 , \44600 , \44601_nG1a9c2 , \44602 , \44603_nG14b06 , \44604_nG14b07 ,
         \44605 , \44606_nG1a9c4 , \44607 , \44608_nG14b08 , \44609_nG14b09 , \44610 , \44611_nG1a9c6 , \44612 , \44613_nG14ae9 , \44614_nG14aea ,
         \44615 , \44616_nG1a9a8 , \44617 , \44618_nG14aeb , \44619_nG14aec , \44620 , \44621_nG1a9aa , \44622 , \44623_nG14aed , \44624_nG14aee ,
         \44625 , \44626_nG1a9ac , \44627 , \44628_nG14aef , \44629_nG14af0 , \44630 , \44631_nG1a9ae , \44632 , \44633_nG14af1 , \44634_nG14af2 ,
         \44635 , \44636_nG1a9b0 , \44637 , \44638_nG14af3 , \44639_nG14af4 , \44640 , \44641_nG1a9b2 , \44642 , \44643_nG14af5 , \44644_nG14af6 ,
         \44645 , \44646_nG1a9b4 , \44647 , \44648_nG14af7 , \44649_nG14af8 , \44650 , \44651_nG1a9b6 , \44652 , \44653_nG14ac8 , \44654_nG14ad1 ,
         \44655 , \44656_nG1abe0 , \44657 , \44658_nG14ad3 , \44659_nG14ad4 , \44660 , \44661_nG1abe2 , \44662 , \44663_nG14ad6 , \44664_nG14ad7 ,
         \44665 , \44666_nG1abe4 , \44667 , \44668_nG14ad9 , \44669_nG14ada , \44670 , \44671_nG1abe6 , \44672 , \44673_nG14adc , \44674_nG14add ,
         \44675 , \44676_nG1abe8 , \44677 , \44678_nG14adf , \44679_nG14ae0 , \44680 , \44681_nG1abea , \44682 , \44683_nG14ae2 , \44684_nG14ae3 ,
         \44685 , \44686_nG1abec , \44687 , \44688_nG14ae5 , \44689_nG14ae6 , \44690 , \44691_nG1abee , \44692 , \44693 , \44694_nGbcb6 ,
         \44695 , \44696 , \44697 , \44698_nG1ac03 , \44699 , \44700 , \44701 , \44702 , \44703 , \44704 ,
         \44705 , \44706 , \44707 , \44708 , \44709 , \44710 , \44711 , \44712 , \44713 , \44714 ,
         \44715 , \44716 , \44717 , \44718 , \44719 , \44720 , \44721 , \44722 , \44723 , \44724 ,
         \44725 , \44726 , \44727 , \44728 , \44729 , \44730 , \44731 , \44732 , \44733 , \44734 ,
         \44735 , \44736 , \44737 , \44738 , \44739 , \44740 , \44741 , \44742 , \44743 , \44744 ,
         \44745 , \44746 , \44747 , \44748 , \44749 , \44750 , \44751 , \44752 , \44753 , \44754 ,
         \44755 , \44756 , \44757 , \44758 , \44759 , \44760 , \44761 , \44762 , \44763 , \44764 ,
         \44765 , \44766_nGe706 , \44767 , \44768_nG1ade5 , \44769 , \44770 , \44771 , \44772 , \44773 , \44774 ,
         \44775 , \44776 , \44777 , \44778 , \44779 , \44780 , \44781 , \44782 , \44783 , \44784 ,
         \44785 , \44786 , \44787 , \44788 , \44789 , \44790 , \44791 , \44792 , \44793 , \44794 ,
         \44795 , \44796 , \44797 , \44798 , \44799 , \44800 , \44801 , \44802 , \44803_nGe728 , \44804 ,
         \44805_nG1ac11 , \44806 , \44807 , \44808 , \44809 , \44810 , \44811_nG17ab0 , \44812 , \44813 , \44814 ,
         \44815 , \44816 , \44817 , \44818_nG17ab1 , \44819 , \44820 , \44821 , \44822 , \44823_nG17ab3 , \44824 ,
         \44825 , \44826 , \44827 , \44828 , \44829 , \44830_nG17ab4 , \44831 , \44832_nG1927e , \44833 , \44834 ,
         \44835_nG17ab5 , \44836_nG17ab6 , \44837 , \44838_nG17ab7 , \44839_nG17ab8 , \44840 , \44841_nG19294 , \44842 , \44843 , \44844_nG17ab9 ,
         \44845_nG17aba , \44846 , \44847_nG17abb , \44848_nG17abc , \44849 , \44850_nG192aa , \44851 , \44852 , \44853_nG17abd , \44854_nG17abe ,
         \44855 , \44856_nG17abf , \44857_nG17ac0 , \44858 , \44859_nG192c0 , \44860 , \44861 , \44862_nG17ac1 , \44863_nG17ac2 , \44864 ,
         \44865_nG17ac3 , \44866_nG17ac4 , \44867 , \44868_nG192d6 , \44869 , \44870 , \44871_nG17ac5 , \44872_nG17ac6 , \44873 , \44874_nG17ac7 ,
         \44875_nG17ac8 , \44876 , \44877_nG192ec , \44878 , \44879 , \44880_nG17ac9 , \44881_nG17aca , \44882 , \44883_nG17acb , \44884_nG17acc ,
         \44885 , \44886_nG192f8 , \44887 , \44888 , \44889_nG17acd , \44890_nG17ace , \44891 , \44892_nG17acf , \44893_nG17ad0 , \44894 ,
         \44895_nG192fa , \44896 , \44897 , \44898_nG17ad1 , \44899_nG17ad2 , \44900 , \44901_nG17ad3 , \44902_nG17ad4 , \44903 , \44904_nG192fc ,
         \44905 , \44906 , \44907_nG17ad5 , \44908_nG17ad6 , \44909 , \44910_nG17ad7 , \44911_nG17ad8 , \44912 , \44913_nG19280 , \44914 ,
         \44915 , \44916_nG17ad9 , \44917_nG17ada , \44918 , \44919_nG17adb , \44920_nG17adc , \44921 , \44922_nG19282 , \44923 , \44924 ,
         \44925_nG17add , \44926_nG17ade , \44927 , \44928_nG17adf , \44929_nG17ae0 , \44930 , \44931_nG19284 , \44932 , \44933 , \44934_nG17ae1 ,
         \44935_nG17ae2 , \44936 , \44937_nG17ae3 , \44938_nG17ae4 , \44939 , \44940_nG19286 , \44941 , \44942 , \44943_nG17ae5 , \44944_nG17ae6 ,
         \44945 , \44946_nG17ae7 , \44947_nG17ae8 , \44948 , \44949_nG19288 , \44950 , \44951 , \44952_nG17ae9 , \44953_nG17aea , \44954 ,
         \44955_nG17aeb , \44956_nG17aec , \44957 , \44958_nG1928a , \44959 , \44960 , \44961_nG17aed , \44962_nG17aee , \44963 , \44964_nG17aef ,
         \44965_nG17af0 , \44966 , \44967_nG1928c , \44968 , \44969 , \44970_nG17af1 , \44971_nG17af2 , \44972 , \44973_nG17af3 , \44974_nG17af4 ,
         \44975 , \44976_nG1928e , \44977 , \44978 , \44979_nG17af5 , \44980_nG17af6 , \44981 , \44982_nG17af7 , \44983_nG17af8 , \44984 ,
         \44985_nG19290 , \44986 , \44987 , \44988_nG17af9 , \44989_nG17afa , \44990 , \44991_nG17afb , \44992_nG17afc , \44993 , \44994_nG19292 ,
         \44995 , \44996 , \44997_nG17afd , \44998_nG17afe , \44999 , \45000_nG17aff , \45001_nG17b00 , \45002 , \45003_nG19296 , \45004 ,
         \45005 , \45006_nG17b01 , \45007_nG17b02 , \45008 , \45009_nG17b03 , \45010_nG17b04 , \45011 , \45012_nG19298 , \45013 , \45014 ,
         \45015_nG17b05 , \45016_nG17b06 , \45017 , \45018_nG17b07 , \45019_nG17b08 , \45020 , \45021_nG1929a , \45022 , \45023 , \45024_nG17b09 ,
         \45025_nG17b0a , \45026 , \45027_nG17b0b , \45028_nG17b0c , \45029 , \45030_nG1929c , \45031 , \45032 , \45033_nG17b0d , \45034_nG17b0e ,
         \45035 , \45036_nG17b0f , \45037_nG17b10 , \45038 , \45039_nG1929e , \45040 , \45041 , \45042_nG17b11 , \45043_nG17b12 , \45044 ,
         \45045_nG17b13 , \45046_nG17b14 , \45047 , \45048_nG192a0 , \45049 , \45050 , \45051_nG17b15 , \45052_nG17b16 , \45053 , \45054_nG17b17 ,
         \45055_nG17b18 , \45056 , \45057_nG192a2 , \45058 , \45059 , \45060_nG17b19 , \45061_nG17b1a , \45062 , \45063_nG17b1b , \45064_nG17b1c ,
         \45065 , \45066_nG192a4 , \45067 , \45068 , \45069_nG17b1d , \45070_nG17b1e , \45071 , \45072_nG17b1f , \45073_nG17b20 , \45074 ,
         \45075_nG192a6 , \45076 , \45077 , \45078_nG17b21 , \45079_nG17b22 , \45080 , \45081_nG17b23 , \45082_nG17b24 , \45083 , \45084_nG192a8 ,
         \45085 , \45086 , \45087_nG17b25 , \45088_nG17b26 , \45089 , \45090_nG17b27 , \45091_nG17b28 , \45092 , \45093_nG192ac , \45094 ,
         \45095 , \45096_nG17b29 , \45097_nG17b2a , \45098 , \45099_nG17b2b , \45100_nG17b2c , \45101 , \45102_nG192ae , \45103 , \45104 ,
         \45105_nG17b2d , \45106_nG17b2e , \45107 , \45108_nG17b2f , \45109_nG17b30 , \45110 , \45111_nG192b0 , \45112 , \45113 , \45114_nG17b31 ,
         \45115_nG17b32 , \45116 , \45117_nG17b33 , \45118_nG17b34 , \45119 , \45120_nG192b2 , \45121 , \45122 , \45123_nG17b35 , \45124_nG17b36 ,
         \45125 , \45126_nG17b37 , \45127_nG17b38 , \45128 , \45129_nG192b4 , \45130 , \45131 , \45132_nG17b39 , \45133_nG17b3a , \45134 ,
         \45135_nG17b3b , \45136_nG17b3c , \45137 , \45138_nG192b6 , \45139 , \45140 , \45141_nG17b3d , \45142_nG17b3e , \45143 , \45144_nG17b3f ,
         \45145_nG17b40 , \45146 , \45147_nG192b8 , \45148 , \45149 , \45150_nG17b41 , \45151_nG17b42 , \45152 , \45153_nG17b43 , \45154_nG17b44 ,
         \45155 , \45156_nG192ba , \45157 , \45158 , \45159_nG17b45 , \45160_nG17b46 , \45161 , \45162_nG17b47 , \45163_nG17b48 , \45164 ,
         \45165_nG192bc , \45166 , \45167 , \45168_nG17b49 , \45169_nG17b4a , \45170 , \45171_nG17b4b , \45172_nG17b4c , \45173 , \45174_nG192be ,
         \45175 , \45176 , \45177_nG17b4d , \45178_nG17b4e , \45179 , \45180_nG17b4f , \45181_nG17b50 , \45182 , \45183_nG192c2 , \45184 ,
         \45185 , \45186_nG17b51 , \45187_nG17b52 , \45188 , \45189_nG17b53 , \45190_nG17b54 , \45191 , \45192_nG192c4 , \45193 , \45194 ,
         \45195_nG17b55 , \45196_nG17b56 , \45197 , \45198_nG17b57 , \45199_nG17b58 , \45200 , \45201_nG192c6 , \45202 , \45203 , \45204_nG17b59 ,
         \45205_nG17b5a , \45206 , \45207_nG17b5b , \45208_nG17b5c , \45209 , \45210_nG192c8 , \45211 , \45212 , \45213_nG17b5d , \45214_nG17b5e ,
         \45215 , \45216_nG17b5f , \45217_nG17b60 , \45218 , \45219_nG192ca , \45220 , \45221 , \45222_nG17b61 , \45223_nG17b62 , \45224 ,
         \45225_nG17b63 , \45226_nG17b64 , \45227 , \45228_nG192cc , \45229 , \45230 , \45231_nG17b65 , \45232_nG17b66 , \45233 , \45234_nG17b67 ,
         \45235_nG17b68 , \45236 , \45237_nG192ce , \45238 , \45239 , \45240_nG17b69 , \45241_nG17b6a , \45242 , \45243_nG17b6b , \45244_nG17b6c ,
         \45245 , \45246_nG192d0 , \45247 , \45248 , \45249_nG17b6d , \45250_nG17b6e , \45251 , \45252_nG17b6f , \45253_nG17b70 , \45254 ,
         \45255_nG192d2 , \45256 , \45257 , \45258_nG17b71 , \45259_nG17b72 , \45260 , \45261_nG17b73 , \45262_nG17b74 , \45263 , \45264_nG192d4 ,
         \45265 , \45266 , \45267_nG17b75 , \45268_nG17b76 , \45269 , \45270_nG17b77 , \45271_nG17b78 , \45272 , \45273_nG192d8 , \45274 ,
         \45275 , \45276_nG17b79 , \45277_nG17b7a , \45278 , \45279_nG17b7b , \45280_nG17b7c , \45281 , \45282_nG192da , \45283 , \45284 ,
         \45285_nG17b7d , \45286_nG17b7e , \45287 , \45288_nG17b7f , \45289_nG17b80 , \45290 , \45291_nG192dc , \45292 , \45293 , \45294_nG17b81 ,
         \45295_nG17b82 , \45296 , \45297_nG17b83 , \45298_nG17b84 , \45299 , \45300_nG192de , \45301 , \45302 , \45303_nG17b85 , \45304_nG17b86 ,
         \45305 , \45306_nG17b87 , \45307_nG17b88 , \45308 , \45309_nG192e0 , \45310 , \45311 , \45312_nG17b89 , \45313_nG17b8a , \45314 ,
         \45315_nG17b8b , \45316_nG17b8c , \45317 , \45318_nG192e2 , \45319 , \45320 , \45321_nG17b8d , \45322_nG17b8e , \45323 , \45324_nG17b8f ,
         \45325_nG17b90 , \45326 , \45327_nG192e4 , \45328 , \45329 , \45330_nG17b91 , \45331_nG17b92 , \45332 , \45333_nG17b93 , \45334_nG17b94 ,
         \45335 , \45336_nG192e6 , \45337 , \45338 , \45339_nG17b95 , \45340_nG17b96 , \45341 , \45342_nG17b97 , \45343_nG17b98 , \45344 ,
         \45345_nG192e8 , \45346 , \45347 , \45348_nG17b99 , \45349_nG17b9a , \45350 , \45351_nG17b9b , \45352_nG17b9c , \45353 , \45354_nG192ea ,
         \45355 , \45356 , \45357_nG17b9d , \45358_nG17b9e , \45359 , \45360_nG17b9f , \45361_nG17ba0 , \45362 , \45363_nG192ee , \45364 ,
         \45365 , \45366_nG17ba1 , \45367_nG17ba2 , \45368 , \45369_nG17ba3 , \45370_nG17ba4 , \45371 , \45372_nG192f0 , \45373 , \45374 ,
         \45375_nG17ba5 , \45376_nG17ba6 , \45377 , \45378_nG17ba7 , \45379_nG17ba8 , \45380 , \45381_nG192f2 , \45382 , \45383 , \45384_nG17ba9 ,
         \45385_nG17baa , \45386 , \45387_nG17bab , \45388_nG17bac , \45389 , \45390_nG192f4 , \45391 , \45392 , \45393_nG17bad , \45394_nG17bae ,
         \45395 , \45396_nG17baf , \45397_nG17bb0 , \45398 , \45399_nG192f6 , \45400 , \45401 , \45402 , \45403_nG179af , \45404_nG179b0 ,
         \45405 , \45406 , \45407_nG179b2 , \45408_nG179b3 , \45409 , \45410_nG191fe , \45411 , \45412_nG179b4 , \45413_nG179b5 , \45414_nG179b6 ,
         \45415_nG179b7 , \45416 , \45417_nG19214 , \45418 , \45419_nG179b8 , \45420_nG179b9 , \45421_nG179ba , \45422_nG179bb , \45423 , \45424_nG1922a ,
         \45425 , \45426_nG179bc , \45427_nG179bd , \45428_nG179be , \45429_nG179bf , \45430 , \45431_nG19240 , \45432 , \45433_nG179c0 , \45434_nG179c1 ,
         \45435_nG179c2 , \45436_nG179c3 , \45437 , \45438_nG19256 , \45439 , \45440_nG179c4 , \45441_nG179c5 , \45442_nG179c6 , \45443_nG179c7 , \45444 ,
         \45445_nG1926c , \45446 , \45447_nG179c8 , \45448_nG179c9 , \45449_nG179ca , \45450_nG179cb , \45451 , \45452_nG19278 , \45453 , \45454_nG179cc ,
         \45455_nG179cd , \45456_nG179ce , \45457_nG179cf , \45458 , \45459_nG1927a , \45460 , \45461_nG179d0 , \45462_nG179d1 , \45463_nG179d2 , \45464_nG179d3 ,
         \45465 , \45466_nG1927c , \45467 , \45468_nG179d4 , \45469_nG179d5 , \45470_nG179d6 , \45471_nG179d7 , \45472 , \45473_nG19200 , \45474 ,
         \45475_nG179d8 , \45476_nG179d9 , \45477_nG179da , \45478_nG179db , \45479 , \45480_nG19202 , \45481 , \45482_nG179dc , \45483_nG179dd , \45484_nG179de ,
         \45485_nG179df , \45486 , \45487_nG19204 , \45488 , \45489_nG179e0 , \45490_nG179e1 , \45491_nG179e2 , \45492_nG179e3 , \45493 , \45494_nG19206 ,
         \45495 , \45496_nG179e4 , \45497_nG179e5 , \45498_nG179e6 , \45499_nG179e7 , \45500 , \45501_nG19208 , \45502 , \45503_nG179e8 , \45504_nG179e9 ,
         \45505_nG179ea , \45506_nG179eb , \45507 , \45508_nG1920a , \45509 , \45510_nG179ec , \45511_nG179ed , \45512_nG179ee , \45513_nG179ef , \45514 ,
         \45515_nG1920c , \45516 , \45517_nG179f0 , \45518_nG179f1 , \45519_nG179f2 , \45520_nG179f3 , \45521 , \45522_nG1920e , \45523 , \45524_nG179f4 ,
         \45525_nG179f5 , \45526_nG179f6 , \45527_nG179f7 , \45528 , \45529_nG19210 , \45530 , \45531_nG179f8 , \45532_nG179f9 , \45533_nG179fa , \45534_nG179fb ,
         \45535 , \45536_nG19212 , \45537 , \45538_nG179fc , \45539_nG179fd , \45540_nG179fe , \45541_nG179ff , \45542 , \45543_nG19216 , \45544 ,
         \45545_nG17a00 , \45546_nG17a01 , \45547_nG17a02 , \45548_nG17a03 , \45549 , \45550_nG19218 , \45551 , \45552_nG17a04 , \45553_nG17a05 , \45554_nG17a06 ,
         \45555_nG17a07 , \45556 , \45557_nG1921a , \45558 , \45559_nG17a08 , \45560_nG17a09 , \45561_nG17a0a , \45562_nG17a0b , \45563 , \45564_nG1921c ,
         \45565 , \45566_nG17a0c , \45567_nG17a0d , \45568_nG17a0e , \45569_nG17a0f , \45570 , \45571_nG1921e , \45572 , \45573_nG17a10 , \45574_nG17a11 ,
         \45575_nG17a12 , \45576_nG17a13 , \45577 , \45578_nG19220 , \45579 , \45580_nG17a14 , \45581_nG17a15 , \45582_nG17a16 , \45583_nG17a17 , \45584 ,
         \45585_nG19222 , \45586 , \45587_nG17a18 , \45588_nG17a19 , \45589_nG17a1a , \45590_nG17a1b , \45591 , \45592_nG19224 , \45593 , \45594_nG17a1c ,
         \45595_nG17a1d , \45596_nG17a1e , \45597_nG17a1f , \45598 , \45599_nG19226 , \45600 , \45601_nG17a20 , \45602_nG17a21 , \45603_nG17a22 , \45604_nG17a23 ,
         \45605 , \45606_nG19228 , \45607 , \45608_nG17a24 , \45609_nG17a25 , \45610_nG17a26 , \45611_nG17a27 , \45612 , \45613_nG1922c , \45614 ,
         \45615_nG17a28 , \45616_nG17a29 , \45617_nG17a2a , \45618_nG17a2b , \45619 , \45620_nG1922e , \45621 , \45622_nG17a2c , \45623_nG17a2d , \45624_nG17a2e ,
         \45625_nG17a2f , \45626 , \45627_nG19230 , \45628 , \45629_nG17a30 , \45630_nG17a31 , \45631_nG17a32 , \45632_nG17a33 , \45633 , \45634_nG19232 ,
         \45635 , \45636_nG17a34 , \45637_nG17a35 , \45638_nG17a36 , \45639_nG17a37 , \45640 , \45641_nG19234 , \45642 , \45643_nG17a38 , \45644_nG17a39 ,
         \45645_nG17a3a , \45646_nG17a3b , \45647 , \45648_nG19236 , \45649 , \45650_nG17a3c , \45651_nG17a3d , \45652_nG17a3e , \45653_nG17a3f , \45654 ,
         \45655_nG19238 , \45656 , \45657_nG17a40 , \45658_nG17a41 , \45659_nG17a42 , \45660_nG17a43 , \45661 , \45662_nG1923a , \45663 , \45664_nG17a44 ,
         \45665_nG17a45 , \45666_nG17a46 , \45667_nG17a47 , \45668 , \45669_nG1923c , \45670 , \45671_nG17a48 , \45672_nG17a49 , \45673_nG17a4a , \45674_nG17a4b ,
         \45675 , \45676_nG1923e , \45677 , \45678_nG17a4c , \45679_nG17a4d , \45680_nG17a4e , \45681_nG17a4f , \45682 , \45683_nG19242 , \45684 ,
         \45685_nG17a50 , \45686_nG17a51 , \45687_nG17a52 , \45688_nG17a53 , \45689 , \45690_nG19244 , \45691 , \45692_nG17a54 , \45693_nG17a55 , \45694_nG17a56 ,
         \45695_nG17a57 , \45696 , \45697_nG19246 , \45698 , \45699_nG17a58 , \45700_nG17a59 , \45701_nG17a5a , \45702_nG17a5b , \45703 , \45704_nG19248 ,
         \45705 , \45706_nG17a5c , \45707_nG17a5d , \45708_nG17a5e , \45709_nG17a5f , \45710 , \45711_nG1924a , \45712 , \45713_nG17a60 , \45714_nG17a61 ,
         \45715_nG17a62 , \45716_nG17a63 , \45717 , \45718_nG1924c , \45719 , \45720_nG17a64 , \45721_nG17a65 , \45722_nG17a66 , \45723_nG17a67 , \45724 ,
         \45725_nG1924e , \45726 , \45727_nG17a68 , \45728_nG17a69 , \45729_nG17a6a , \45730_nG17a6b , \45731 , \45732_nG19250 , \45733 , \45734_nG17a6c ,
         \45735_nG17a6d , \45736_nG17a6e , \45737_nG17a6f , \45738 , \45739_nG19252 , \45740 , \45741_nG17a70 , \45742_nG17a71 , \45743_nG17a72 , \45744_nG17a73 ,
         \45745 , \45746_nG19254 , \45747 , \45748_nG17a74 , \45749_nG17a75 , \45750_nG17a76 , \45751_nG17a77 , \45752 , \45753_nG19258 , \45754 ,
         \45755_nG17a78 , \45756_nG17a79 , \45757_nG17a7a , \45758_nG17a7b , \45759 , \45760_nG1925a , \45761 , \45762_nG17a7c , \45763_nG17a7d , \45764_nG17a7e ,
         \45765_nG17a7f , \45766 , \45767_nG1925c , \45768 , \45769_nG17a80 , \45770_nG17a81 , \45771_nG17a82 , \45772_nG17a83 , \45773 , \45774_nG1925e ,
         \45775 , \45776_nG17a84 , \45777_nG17a85 , \45778_nG17a86 , \45779_nG17a87 , \45780 , \45781_nG19260 , \45782 , \45783_nG17a88 , \45784_nG17a89 ,
         \45785_nG17a8a , \45786_nG17a8b , \45787 , \45788_nG19262 , \45789 , \45790_nG17a8c , \45791_nG17a8d , \45792_nG17a8e , \45793_nG17a8f , \45794 ,
         \45795_nG19264 , \45796 , \45797_nG17a90 , \45798_nG17a91 , \45799_nG17a92 , \45800_nG17a93 , \45801 , \45802_nG19266 , \45803 , \45804_nG17a94 ,
         \45805_nG17a95 , \45806_nG17a96 , \45807_nG17a97 , \45808 , \45809_nG19268 , \45810 , \45811_nG17a98 , \45812_nG17a99 , \45813_nG17a9a , \45814_nG17a9b ,
         \45815 , \45816_nG1926a , \45817 , \45818_nG17a9c , \45819_nG17a9d , \45820_nG17a9e , \45821_nG17a9f , \45822 , \45823_nG1926e , \45824 ,
         \45825_nG17aa0 , \45826_nG17aa1 , \45827_nG17aa2 , \45828_nG17aa3 , \45829 , \45830_nG19270 , \45831 , \45832_nG17aa4 , \45833_nG17aa5 , \45834_nG17aa6 ,
         \45835_nG17aa7 , \45836 , \45837_nG19272 , \45838 , \45839_nG17aa8 , \45840_nG17aa9 , \45841_nG17aaa , \45842_nG17aab , \45843 , \45844_nG19274 ,
         \45845 , \45846_nG17aac , \45847_nG17aad , \45848_nG17aae , \45849_nG17aaf , \45850 , \45851_nG19276 , \45852 , \45853 , \45854_nG178ad ,
         \45855_nG178ae , \45856 , \45857_nG178b1 , \45858_nG178b2 , \45859 , \45860_nG1917e , \45861 , \45862_nG178b3 , \45863_nG178b4 , \45864_nG178b5 ,
         \45865_nG178b6 , \45866 , \45867_nG19194 , \45868 , \45869_nG178b7 , \45870_nG178b8 , \45871_nG178b9 , \45872_nG178ba , \45873 , \45874_nG191aa ,
         \45875 , \45876_nG178bb , \45877_nG178bc , \45878_nG178bd , \45879_nG178be , \45880 , \45881_nG191c0 , \45882 , \45883_nG178bf , \45884_nG178c0 ,
         \45885_nG178c1 , \45886_nG178c2 , \45887 , \45888_nG191d6 , \45889 , \45890_nG178c3 , \45891_nG178c4 , \45892_nG178c5 , \45893_nG178c6 , \45894 ,
         \45895_nG191ec , \45896 , \45897_nG178c7 , \45898_nG178c8 , \45899_nG178c9 , \45900_nG178ca , \45901 , \45902_nG191f8 , \45903 , \45904_nG178cb ,
         \45905_nG178cc , \45906_nG178cd , \45907_nG178ce , \45908 , \45909_nG191fa , \45910 , \45911_nG178cf , \45912_nG178d0 , \45913_nG178d1 , \45914_nG178d2 ,
         \45915 , \45916_nG191fc , \45917 , \45918_nG178d3 , \45919_nG178d4 , \45920_nG178d5 , \45921_nG178d6 , \45922 , \45923_nG19180 , \45924 ,
         \45925_nG178d7 , \45926_nG178d8 , \45927_nG178d9 , \45928_nG178da , \45929 , \45930_nG19182 , \45931 , \45932_nG178db , \45933_nG178dc , \45934_nG178dd ,
         \45935_nG178de , \45936 , \45937_nG19184 , \45938 , \45939_nG178df , \45940_nG178e0 , \45941_nG178e1 , \45942_nG178e2 , \45943 , \45944_nG19186 ,
         \45945 , \45946_nG178e3 , \45947_nG178e4 , \45948_nG178e5 , \45949_nG178e6 , \45950 , \45951_nG19188 , \45952 , \45953_nG178e7 , \45954_nG178e8 ,
         \45955_nG178e9 , \45956_nG178ea , \45957 , \45958_nG1918a , \45959 , \45960_nG178eb , \45961_nG178ec , \45962_nG178ed , \45963_nG178ee , \45964 ,
         \45965_nG1918c , \45966 , \45967_nG178ef , \45968_nG178f0 , \45969_nG178f1 , \45970_nG178f2 , \45971 , \45972_nG1918e , \45973 , \45974_nG178f3 ,
         \45975_nG178f4 , \45976_nG178f5 , \45977_nG178f6 , \45978 , \45979_nG19190 , \45980 , \45981_nG178f7 , \45982_nG178f8 , \45983_nG178f9 , \45984_nG178fa ,
         \45985 , \45986_nG19192 , \45987 , \45988_nG178fb , \45989_nG178fc , \45990_nG178fd , \45991_nG178fe , \45992 , \45993_nG19196 , \45994 ,
         \45995_nG178ff , \45996_nG17900 , \45997_nG17901 , \45998_nG17902 , \45999 , \46000_nG19198 , \46001 , \46002_nG17903 , \46003_nG17904 , \46004_nG17905 ,
         \46005_nG17906 , \46006 , \46007_nG1919a , \46008 , \46009_nG17907 , \46010_nG17908 , \46011_nG17909 , \46012_nG1790a , \46013 , \46014_nG1919c ,
         \46015 , \46016_nG1790b , \46017_nG1790c , \46018_nG1790d , \46019_nG1790e , \46020 , \46021_nG1919e , \46022 , \46023_nG1790f , \46024_nG17910 ,
         \46025_nG17911 , \46026_nG17912 , \46027 , \46028_nG191a0 , \46029 , \46030_nG17913 , \46031_nG17914 , \46032_nG17915 , \46033_nG17916 , \46034 ,
         \46035_nG191a2 , \46036 , \46037_nG17917 , \46038_nG17918 , \46039_nG17919 , \46040_nG1791a , \46041 , \46042_nG191a4 , \46043 , \46044_nG1791b ,
         \46045_nG1791c , \46046_nG1791d , \46047_nG1791e , \46048 , \46049_nG191a6 , \46050 , \46051_nG1791f , \46052_nG17920 , \46053_nG17921 , \46054_nG17922 ,
         \46055 , \46056_nG191a8 , \46057 , \46058_nG17923 , \46059_nG17924 , \46060_nG17925 , \46061_nG17926 , \46062 , \46063_nG191ac , \46064 ,
         \46065_nG17927 , \46066_nG17928 , \46067_nG17929 , \46068_nG1792a , \46069 , \46070_nG191ae , \46071 , \46072_nG1792b , \46073_nG1792c , \46074_nG1792d ,
         \46075_nG1792e , \46076 , \46077_nG191b0 , \46078 , \46079_nG1792f , \46080_nG17930 , \46081_nG17931 , \46082_nG17932 , \46083 , \46084_nG191b2 ,
         \46085 , \46086_nG17933 , \46087_nG17934 , \46088_nG17935 , \46089_nG17936 , \46090 , \46091_nG191b4 , \46092 , \46093_nG17937 , \46094_nG17938 ,
         \46095_nG17939 , \46096_nG1793a , \46097 , \46098_nG191b6 , \46099 , \46100_nG1793b , \46101_nG1793c , \46102_nG1793d , \46103_nG1793e , \46104 ,
         \46105_nG191b8 , \46106 , \46107_nG1793f , \46108_nG17940 , \46109_nG17941 , \46110_nG17942 , \46111 , \46112_nG191ba , \46113 , \46114_nG17943 ,
         \46115_nG17944 , \46116_nG17945 , \46117_nG17946 , \46118 , \46119_nG191bc , \46120 , \46121_nG17947 , \46122_nG17948 , \46123_nG17949 , \46124_nG1794a ,
         \46125 , \46126_nG191be , \46127 , \46128_nG1794b , \46129_nG1794c , \46130_nG1794d , \46131_nG1794e , \46132 , \46133_nG191c2 , \46134 ,
         \46135_nG1794f , \46136_nG17950 , \46137_nG17951 , \46138_nG17952 , \46139 , \46140_nG191c4 , \46141 , \46142_nG17953 , \46143_nG17954 , \46144_nG17955 ,
         \46145_nG17956 , \46146 , \46147_nG191c6 , \46148 , \46149_nG17957 , \46150_nG17958 , \46151_nG17959 , \46152_nG1795a , \46153 , \46154_nG191c8 ,
         \46155 , \46156_nG1795b , \46157_nG1795c , \46158_nG1795d , \46159_nG1795e , \46160 , \46161_nG191ca , \46162 , \46163_nG1795f , \46164_nG17960 ,
         \46165_nG17961 , \46166_nG17962 , \46167 , \46168_nG191cc , \46169 , \46170_nG17963 , \46171_nG17964 , \46172_nG17965 , \46173_nG17966 , \46174 ,
         \46175_nG191ce , \46176 , \46177_nG17967 , \46178_nG17968 , \46179_nG17969 , \46180_nG1796a , \46181 , \46182_nG191d0 , \46183 , \46184_nG1796b ,
         \46185_nG1796c , \46186_nG1796d , \46187_nG1796e , \46188 , \46189_nG191d2 , \46190 , \46191_nG1796f , \46192_nG17970 , \46193_nG17971 , \46194_nG17972 ,
         \46195 , \46196_nG191d4 , \46197 , \46198_nG17973 , \46199_nG17974 , \46200_nG17975 , \46201_nG17976 , \46202 , \46203_nG191d8 , \46204 ,
         \46205_nG17977 , \46206_nG17978 , \46207_nG17979 , \46208_nG1797a , \46209 , \46210_nG191da , \46211 , \46212_nG1797b , \46213_nG1797c , \46214_nG1797d ,
         \46215_nG1797e , \46216 , \46217_nG191dc , \46218 , \46219_nG1797f , \46220_nG17980 , \46221_nG17981 , \46222_nG17982 , \46223 , \46224_nG191de ,
         \46225 , \46226_nG17983 , \46227_nG17984 , \46228_nG17985 , \46229_nG17986 , \46230 , \46231_nG191e0 , \46232 , \46233_nG17987 , \46234_nG17988 ,
         \46235_nG17989 , \46236_nG1798a , \46237 , \46238_nG191e2 , \46239 , \46240_nG1798b , \46241_nG1798c , \46242_nG1798d , \46243_nG1798e , \46244 ,
         \46245_nG191e4 , \46246 , \46247_nG1798f , \46248_nG17990 , \46249_nG17991 , \46250_nG17992 , \46251 , \46252_nG191e6 , \46253 , \46254_nG17993 ,
         \46255_nG17994 , \46256_nG17995 , \46257_nG17996 , \46258 , \46259_nG191e8 , \46260 , \46261_nG17997 , \46262_nG17998 , \46263_nG17999 , \46264_nG1799a ,
         \46265 , \46266_nG191ea , \46267 , \46268_nG1799b , \46269_nG1799c , \46270_nG1799d , \46271_nG1799e , \46272 , \46273_nG191ee , \46274 ,
         \46275_nG1799f , \46276_nG179a0 , \46277_nG179a1 , \46278_nG179a2 , \46279 , \46280_nG191f0 , \46281 , \46282_nG179a3 , \46283_nG179a4 , \46284_nG179a5 ,
         \46285_nG179a6 , \46286 , \46287_nG191f2 , \46288 , \46289_nG179a7 , \46290_nG179a8 , \46291_nG179a9 , \46292_nG179aa , \46293 , \46294_nG191f4 ,
         \46295 , \46296_nG179ab , \46297_nG179ac , \46298_nG179ad , \46299_nG179ae , \46300 , \46301_nG191f6 , \46302 , \46303 , \46304_nG1772b ,
         \46305_nG1772c , \46306 , \46307_nG17731 , \46308_nG17732 , \46309 , \46310_nG190fe , \46311 , \46312_nG17734 , \46313_nG17735 , \46314_nG17737 ,
         \46315_nG17738 , \46316 , \46317_nG19114 , \46318 , \46319_nG1773a , \46320_nG1773b , \46321_nG1773d , \46322_nG1773e , \46323 , \46324_nG1912a ,
         \46325 , \46326_nG17740 , \46327_nG17741 , \46328_nG17743 , \46329_nG17744 , \46330 , \46331_nG19140 , \46332 , \46333_nG17746 , \46334_nG17747 ,
         \46335_nG17749 , \46336_nG1774a , \46337 , \46338_nG19156 , \46339 , \46340_nG1774c , \46341_nG1774d , \46342_nG1774f , \46343_nG17750 , \46344 ,
         \46345_nG1916c , \46346 , \46347_nG17752 , \46348_nG17753 , \46349_nG17755 , \46350_nG17756 , \46351 , \46352_nG19178 , \46353 , \46354_nG17758 ,
         \46355_nG17759 , \46356_nG1775b , \46357_nG1775c , \46358 , \46359_nG1917a , \46360 , \46361_nG1775e , \46362_nG1775f , \46363_nG17761 , \46364_nG17762 ,
         \46365 , \46366_nG1917c , \46367 , \46368_nG17764 , \46369_nG17765 , \46370_nG17767 , \46371_nG17768 , \46372 , \46373_nG19100 , \46374 ,
         \46375_nG1776a , \46376_nG1776b , \46377_nG1776d , \46378_nG1776e , \46379 , \46380_nG19102 , \46381 , \46382_nG17770 , \46383_nG17771 , \46384_nG17773 ,
         \46385_nG17774 , \46386 , \46387_nG19104 , \46388 , \46389_nG17776 , \46390_nG17777 , \46391_nG17779 , \46392_nG1777a , \46393 , \46394_nG19106 ,
         \46395 , \46396_nG1777c , \46397_nG1777d , \46398_nG1777f , \46399_nG17780 , \46400 , \46401_nG19108 , \46402 , \46403_nG17782 , \46404_nG17783 ,
         \46405_nG17785 , \46406_nG17786 , \46407 , \46408_nG1910a , \46409 , \46410_nG17788 , \46411_nG17789 , \46412_nG1778b , \46413_nG1778c , \46414 ,
         \46415_nG1910c , \46416 , \46417_nG1778e , \46418_nG1778f , \46419_nG17791 , \46420_nG17792 , \46421 , \46422_nG1910e , \46423 , \46424_nG17794 ,
         \46425_nG17795 , \46426_nG17797 , \46427_nG17798 , \46428 , \46429_nG19110 , \46430 , \46431_nG1779a , \46432_nG1779b , \46433_nG1779d , \46434_nG1779e ,
         \46435 , \46436_nG19112 , \46437 , \46438_nG177a0 , \46439_nG177a1 , \46440_nG177a3 , \46441_nG177a4 , \46442 , \46443_nG19116 , \46444 ,
         \46445_nG177a6 , \46446_nG177a7 , \46447_nG177a9 , \46448_nG177aa , \46449 , \46450_nG19118 , \46451 , \46452_nG177ac , \46453_nG177ad , \46454_nG177af ,
         \46455_nG177b0 , \46456 , \46457_nG1911a , \46458 , \46459_nG177b2 , \46460_nG177b3 , \46461_nG177b5 , \46462_nG177b6 , \46463 , \46464_nG1911c ,
         \46465 , \46466_nG177b8 , \46467_nG177b9 , \46468_nG177bb , \46469_nG177bc , \46470 , \46471_nG1911e , \46472 , \46473_nG177be , \46474_nG177bf ,
         \46475_nG177c1 , \46476_nG177c2 , \46477 , \46478_nG19120 , \46479 , \46480_nG177c4 , \46481_nG177c5 , \46482_nG177c7 , \46483_nG177c8 , \46484 ,
         \46485_nG19122 , \46486 , \46487_nG177ca , \46488_nG177cb , \46489_nG177cd , \46490_nG177ce , \46491 , \46492_nG19124 , \46493 , \46494_nG177d0 ,
         \46495_nG177d1 , \46496_nG177d3 , \46497_nG177d4 , \46498 , \46499_nG19126 , \46500 , \46501_nG177d6 , \46502_nG177d7 , \46503_nG177d9 , \46504_nG177da ,
         \46505 , \46506_nG19128 , \46507 , \46508_nG177dc , \46509_nG177dd , \46510_nG177df , \46511_nG177e0 , \46512 , \46513_nG1912c , \46514 ,
         \46515_nG177e2 , \46516_nG177e3 , \46517_nG177e5 , \46518_nG177e6 , \46519 , \46520_nG1912e , \46521 , \46522_nG177e8 , \46523_nG177e9 , \46524_nG177eb ,
         \46525_nG177ec , \46526 , \46527_nG19130 , \46528 , \46529_nG177ee , \46530_nG177ef , \46531_nG177f1 , \46532_nG177f2 , \46533 , \46534_nG19132 ,
         \46535 , \46536_nG177f4 , \46537_nG177f5 , \46538_nG177f7 , \46539_nG177f8 , \46540 , \46541_nG19134 , \46542 , \46543_nG177fa , \46544_nG177fb ,
         \46545_nG177fd , \46546_nG177fe , \46547 , \46548_nG19136 , \46549 , \46550_nG17800 , \46551_nG17801 , \46552_nG17803 , \46553_nG17804 , \46554 ,
         \46555_nG19138 , \46556 , \46557_nG17806 , \46558_nG17807 , \46559_nG17809 , \46560_nG1780a , \46561 , \46562_nG1913a , \46563 , \46564_nG1780c ,
         \46565_nG1780d , \46566_nG1780f , \46567_nG17810 , \46568 , \46569_nG1913c , \46570 , \46571_nG17812 , \46572_nG17813 , \46573_nG17815 , \46574_nG17816 ,
         \46575 , \46576_nG1913e , \46577 , \46578_nG17818 , \46579_nG17819 , \46580_nG1781b , \46581_nG1781c , \46582 , \46583_nG19142 , \46584 ,
         \46585_nG1781e , \46586_nG1781f , \46587_nG17821 , \46588_nG17822 , \46589 , \46590_nG19144 , \46591 , \46592_nG17824 , \46593_nG17825 , \46594_nG17827 ,
         \46595_nG17828 , \46596 , \46597_nG19146 , \46598 , \46599_nG1782a , \46600_nG1782b , \46601_nG1782d , \46602_nG1782e , \46603 , \46604_nG19148 ,
         \46605 , \46606_nG17830 , \46607_nG17831 , \46608_nG17833 , \46609_nG17834 , \46610 , \46611_nG1914a , \46612 , \46613_nG17836 , \46614_nG17837 ,
         \46615_nG17839 , \46616_nG1783a , \46617 , \46618_nG1914c , \46619 , \46620_nG1783c , \46621_nG1783d , \46622_nG1783f , \46623_nG17840 , \46624 ,
         \46625_nG1914e , \46626 , \46627_nG17842 , \46628_nG17843 , \46629_nG17845 , \46630_nG17846 , \46631 , \46632_nG19150 , \46633 , \46634_nG17848 ,
         \46635_nG17849 , \46636_nG1784b , \46637_nG1784c , \46638 , \46639_nG19152 , \46640 , \46641_nG1784e , \46642_nG1784f , \46643_nG17851 , \46644_nG17852 ,
         \46645 , \46646_nG19154 , \46647 , \46648_nG17854 , \46649_nG17855 , \46650_nG17857 , \46651_nG17858 , \46652 , \46653_nG19158 , \46654 ,
         \46655_nG1785a , \46656_nG1785b , \46657_nG1785d , \46658_nG1785e , \46659 , \46660_nG1915a , \46661 , \46662_nG17860 , \46663_nG17861 , \46664_nG17863 ,
         \46665_nG17864 , \46666 , \46667_nG1915c , \46668 , \46669_nG17866 , \46670_nG17867 , \46671_nG17869 , \46672_nG1786a , \46673 , \46674_nG1915e ,
         \46675 , \46676_nG1786c , \46677_nG1786d , \46678_nG1786f , \46679_nG17870 , \46680 , \46681_nG19160 , \46682 , \46683_nG17872 , \46684_nG17873 ,
         \46685_nG17875 , \46686_nG17876 , \46687 , \46688_nG19162 , \46689 , \46690_nG17878 , \46691_nG17879 , \46692_nG1787b , \46693_nG1787c , \46694 ,
         \46695_nG19164 , \46696 , \46697_nG1787e , \46698_nG1787f , \46699_nG17881 , \46700_nG17882 , \46701 , \46702_nG19166 , \46703 , \46704_nG17884 ,
         \46705_nG17885 , \46706_nG17887 , \46707_nG17888 , \46708 , \46709_nG19168 , \46710 , \46711_nG1788a , \46712_nG1788b , \46713_nG1788d , \46714_nG1788e ,
         \46715 , \46716_nG1916a , \46717 , \46718_nG17890 , \46719_nG17891 , \46720_nG17893 , \46721_nG17894 , \46722 , \46723_nG1916e , \46724 ,
         \46725_nG17896 , \46726_nG17897 , \46727_nG17899 , \46728_nG1789a , \46729 , \46730_nG19170 , \46731 , \46732_nG1789c , \46733_nG1789d , \46734_nG1789f ,
         \46735_nG178a0 , \46736 , \46737_nG19172 , \46738 , \46739_nG178a2 , \46740_nG178a3 , \46741_nG178a5 , \46742_nG178a6 , \46743 , \46744_nG19174 ,
         \46745 , \46746_nG178a8 , \46747_nG178a9 , \46748_nG178ab , \46749_nG178ac , \46750 , \46751_nG19176 , \46752 , \46753 , \46754_nG176fd ,
         \46755 , \46756 , \46757_nG176fe , \46758 , \46759_nG190e6 , \46760 , \46761 , \46762_nG176ff , \46763_nG17700 , \46764 ,
         \46765_nG190e8 , \46766 , \46767 , \46768_nG17701 , \46769_nG17702 , \46770 , \46771_nG190ea , \46772 , \46773 , \46774_nG17703 ,
         \46775_nG17704 , \46776 , \46777_nG190ec , \46778 , \46779 , \46780_nG17705 , \46781_nG17706 , \46782 , \46783_nG190ee , \46784 ,
         \46785 , \46786_nG17707 , \46787_nG17708 , \46788 , \46789_nG190f0 , \46790 , \46791 , \46792_nG17709 , \46793_nG1770a , \46794 ,
         \46795_nG190f2 , \46796 , \46797 , \46798_nG1770b , \46799_nG1770c , \46800 , \46801_nG190f4 , \46802 , \46803_nG176ec , \46804_nG176ed ,
         \46805 , \46806_nG190d6 , \46807 , \46808_nG176ee , \46809_nG176ef , \46810 , \46811_nG190d8 , \46812 , \46813_nG176f0 , \46814_nG176f1 ,
         \46815 , \46816_nG190da , \46817 , \46818_nG176f2 , \46819_nG176f3 , \46820 , \46821_nG190dc , \46822 , \46823_nG176f4 , \46824_nG176f5 ,
         \46825 , \46826_nG190de , \46827 , \46828_nG176f6 , \46829_nG176f7 , \46830 , \46831_nG190e0 , \46832 , \46833_nG176f8 , \46834_nG176f9 ,
         \46835 , \46836_nG190e2 , \46837 , \46838_nG176fa , \46839_nG176fb , \46840 , \46841_nG190e4 , \46842 , \46843_nG176db , \46844_nG176dc ,
         \46845 , \46846_nG190c6 , \46847 , \46848_nG176dd , \46849_nG176de , \46850 , \46851_nG190c8 , \46852 , \46853_nG176df , \46854_nG176e0 ,
         \46855 , \46856_nG190ca , \46857 , \46858_nG176e1 , \46859_nG176e2 , \46860 , \46861_nG190cc , \46862 , \46863_nG176e3 , \46864_nG176e4 ,
         \46865 , \46866_nG190ce , \46867 , \46868_nG176e5 , \46869_nG176e6 , \46870 , \46871_nG190d0 , \46872 , \46873_nG176e7 , \46874_nG176e8 ,
         \46875 , \46876_nG190d2 , \46877 , \46878_nG176e9 , \46879_nG176ea , \46880 , \46881_nG190d4 , \46882 , \46883_nG176ba , \46884_nG176c3 ,
         \46885 , \46886_nG192fe , \46887 , \46888_nG176c5 , \46889_nG176c6 , \46890 , \46891_nG19300 , \46892 , \46893_nG176c8 , \46894_nG176c9 ,
         \46895 , \46896_nG19302 , \46897 , \46898_nG176cb , \46899_nG176cc , \46900 , \46901_nG19304 , \46902 , \46903_nG176ce , \46904_nG176cf ,
         \46905 , \46906_nG19306 , \46907 , \46908_nG176d1 , \46909_nG176d2 , \46910 , \46911_nG19308 , \46912 , \46913_nG176d4 , \46914_nG176d5 ,
         \46915 , \46916_nG1930a , \46917 , \46918_nG176d7 , \46919_nG176d8 , \46920 , \46921_nG1930c , \46922 , \46923 , \46924 ,
         \46925 , \46926_nG175af , \46927 , \46928_nG1930d , \46929 , \46930 , \46931_nG1761c , \46932 , \46933_nG190aa , \46934 ,
         \46935 , \46936_nG1761e , \46937 , \46938_nG190ac , \46939 , \46940 , \46941_nG17620 , \46942 , \46943_nG190ae , \46944 ,
         \46945 , \46946_nG17622 , \46947 , \46948_nG190b0 , \46949 , \46950 , \46951_nG17624 , \46952 , \46953_nG190b2 , \46954 ,
         \46955 , \46956_nG17626 , \46957 , \46958_nG190b4 , \46959 , \46960 , \46961_nG17628 , \46962 , \46963_nG190b6 , \46964 ,
         \46965 , \46966_nG1761a , \46967 , \46968_nG190a8 , \46969 , \46970 , \46971_nG17612 , \46972 , \46973_nG190a0 , \46974 ,
         \46975 , \46976_nG17614 , \46977 , \46978_nG190a2 , \46979 , \46980 , \46981_nG17616 , \46982 , \46983_nG190a4 , \46984 ,
         \46985 , \46986_nG17618 , \46987 , \46988_nG190a6 , \46989 , \46990 , \46991 , \46992 , \46993 , \46994_nG17482 ,
         \46995 , \46996 , \46997 , \46998 , \46999_nG17483 , \47000 , \47001 , \47002 , \47003 , \47004 ,
         \47005_nG17489 , \47006 , \47007_nG1748d , \47008 , \47009 , \47010_nG17490 , \47011 , \47012 , \47013 , \47014 ,
         \47015 , \47016_nG17497 , \47017 , \47018 , \47019_nG17498 , \47020 , \47021 , \47022 , \47023 , \47024_nG1749c ,
         \47025_nG1749d , \47026 , \47027 , \47028 , \47029_nG174a1 , \47030_nG174a2 , \47031_nG174a3 , \47032_nG174a4 , \47033_nG174a5 , \47034 ,
         \47035 , \47036 , \47037 , \47038 , \47039_nG174aa , \47040_nG174ab , \47041 , \47042 , \47043 , \47044 ,
         \47045_nG174b0 , \47046_nG174b1 , \47047_nG174b2 , \47048_nG174b3 , \47049_nG174b4 , \47050 , \47051 , \47052 , \47053 , \47054 ,
         \47055 , \47056 , \47057 , \47058 , \47059 , \47060 , \47061 , \47062 , \47063_nG17479 , \47064_nG1747a ,
         \47065 , \47066 , \47067 , \47068 , \47069 , \47070 , \47071 , \47072 , \47073 , \47074 ,
         \47075 , \47076 , \47077 , \47078 , \47079_nG17537 , \47080 , \47081 , \47082 , \47083 , \47084 ,
         \47085 , \47086 , \47087_nG1753b , \47088 , \47089 , \47090_nG1753c , \47091 , \47092 , \47093_nG1753d , \47094 ,
         \47095_nG1753e , \47096 , \47097 , \47098 , \47099 , \47100_nG17473 , \47101_nG17474 , \47102 , \47103 , \47104 ,
         \47105 , \47106_nG17528 , \47107 , \47108 , \47109_nG1752f , \47110_nG17530 , \47111_nG17531 , \47112_nG17532 , \47113 , \47114 ,
         \47115 , \47116 , \47117_nG1746c , \47118_nG1746f , \47119 , \47120 , \47121 , \47122 , \47123_nG17518 , \47124 ,
         \47125_nG1751c , \47126_nG1751f , \47127_nG17522 , \47128_nG17524 , \47129 , \47130 , \47131 , \47132 , \47133 , \47134 ,
         \47135 , \47136 , \47137 , \47138 , \47139 , \47140 , \47141 , \47142_nG175b3 , \47143 , \47144_nG190c4 ,
         \47145 , \47146 , \47147_nG19311 , \47148 , \47149 , \47150_nG19312 , \47151 , \47152 , \47153_nG19313 , \47154 ,
         \47155 , \47156 , \47157 , \47158 , \47159_nG1735d , \47160 , \47161 , \47162 , \47163 , \47164 ,
         \47165 , \47166 , \47167_nG1735e , \47168 , \47169 , \47170 , \47171 , \47172_nG17360 , \47173 , \47174 ,
         \47175 , \47176 , \47177 , \47178 , \47179_nG17361 , \47180 , \47181_nG19001 , \47182 , \47183 , \47184_nG17362 ,
         \47185_nG17363 , \47186 , \47187_nG17364 , \47188_nG17365 , \47189 , \47190_nG19017 , \47191 , \47192 , \47193_nG17366 , \47194_nG17367 ,
         \47195 , \47196_nG17368 , \47197_nG17369 , \47198 , \47199_nG1902d , \47200 , \47201 , \47202_nG1736a , \47203_nG1736b , \47204 ,
         \47205_nG1736c , \47206_nG1736d , \47207 , \47208_nG19043 , \47209 , \47210 , \47211_nG1736e , \47212_nG1736f , \47213 , \47214_nG17370 ,
         \47215_nG17371 , \47216 , \47217_nG19059 , \47218 , \47219 , \47220_nG17372 , \47221_nG17373 , \47222 , \47223_nG17374 , \47224_nG17375 ,
         \47225 , \47226_nG1906f , \47227 , \47228 , \47229_nG17376 , \47230_nG17377 , \47231 , \47232_nG17378 , \47233_nG17379 , \47234 ,
         \47235_nG1907b , \47236 , \47237 , \47238_nG1737a , \47239_nG1737b , \47240 , \47241_nG1737c , \47242_nG1737d , \47243 , \47244_nG1907d ,
         \47245 , \47246 , \47247_nG1737e , \47248_nG1737f , \47249 , \47250_nG17380 , \47251_nG17381 , \47252 , \47253_nG1907f , \47254 ,
         \47255 , \47256_nG17382 , \47257_nG17383 , \47258 , \47259_nG17384 , \47260_nG17385 , \47261 , \47262_nG19003 , \47263 , \47264 ,
         \47265_nG17386 , \47266_nG17387 , \47267 , \47268_nG17388 , \47269_nG17389 , \47270 , \47271_nG19005 , \47272 , \47273 , \47274_nG1738a ,
         \47275_nG1738b , \47276 , \47277_nG1738c , \47278_nG1738d , \47279 , \47280_nG19007 , \47281 , \47282 , \47283_nG1738e , \47284_nG1738f ,
         \47285 , \47286_nG17390 , \47287_nG17391 , \47288 , \47289_nG19009 , \47290 , \47291 , \47292_nG17392 , \47293_nG17393 , \47294 ,
         \47295_nG17394 , \47296_nG17395 , \47297 , \47298_nG1900b , \47299 , \47300 , \47301_nG17396 , \47302_nG17397 , \47303 , \47304_nG17398 ,
         \47305_nG17399 , \47306 , \47307_nG1900d , \47308 , \47309 , \47310_nG1739a , \47311_nG1739b , \47312 , \47313_nG1739c , \47314_nG1739d ,
         \47315 , \47316_nG1900f , \47317 , \47318 , \47319_nG1739e , \47320_nG1739f , \47321 , \47322_nG173a0 , \47323_nG173a1 , \47324 ,
         \47325_nG19011 , \47326 , \47327 , \47328_nG173a2 , \47329_nG173a3 , \47330 , \47331_nG173a4 , \47332_nG173a5 , \47333 , \47334_nG19013 ,
         \47335 , \47336 , \47337_nG173a6 , \47338_nG173a7 , \47339 , \47340_nG173a8 , \47341_nG173a9 , \47342 , \47343_nG19015 , \47344 ,
         \47345 , \47346_nG173aa , \47347_nG173ab , \47348 , \47349_nG173ac , \47350_nG173ad , \47351 , \47352_nG19019 , \47353 , \47354 ,
         \47355_nG173ae , \47356_nG173af , \47357 , \47358_nG173b0 , \47359_nG173b1 , \47360 , \47361_nG1901b , \47362 , \47363 , \47364_nG173b2 ,
         \47365_nG173b3 , \47366 , \47367_nG173b4 , \47368_nG173b5 , \47369 , \47370_nG1901d , \47371 , \47372 , \47373_nG173b6 , \47374_nG173b7 ,
         \47375 , \47376_nG173b8 , \47377_nG173b9 , \47378 , \47379_nG1901f , \47380 , \47381 , \47382_nG173ba , \47383_nG173bb , \47384 ,
         \47385_nG173bc , \47386_nG173bd , \47387 , \47388_nG19021 , \47389 , \47390 , \47391_nG173be , \47392_nG173bf , \47393 , \47394_nG173c0 ,
         \47395_nG173c1 , \47396 , \47397_nG19023 , \47398 , \47399 , \47400_nG173c2 , \47401_nG173c3 , \47402 , \47403_nG173c4 , \47404_nG173c5 ,
         \47405 , \47406_nG19025 , \47407 , \47408 , \47409_nG173c6 , \47410_nG173c7 , \47411 , \47412_nG173c8 , \47413_nG173c9 , \47414 ,
         \47415_nG19027 , \47416 , \47417 , \47418_nG173ca , \47419_nG173cb , \47420 , \47421_nG173cc , \47422_nG173cd , \47423 , \47424_nG19029 ,
         \47425 , \47426 , \47427_nG173ce , \47428_nG173cf , \47429 , \47430_nG173d0 , \47431_nG173d1 , \47432 , \47433_nG1902b , \47434 ,
         \47435 , \47436_nG173d2 , \47437_nG173d3 , \47438 , \47439_nG173d4 , \47440_nG173d5 , \47441 , \47442_nG1902f , \47443 , \47444 ,
         \47445_nG173d6 , \47446_nG173d7 , \47447 , \47448_nG173d8 , \47449_nG173d9 , \47450 , \47451_nG19031 , \47452 , \47453 , \47454_nG173da ,
         \47455_nG173db , \47456 , \47457_nG173dc , \47458_nG173dd , \47459 , \47460_nG19033 , \47461 , \47462 , \47463_nG173de , \47464_nG173df ,
         \47465 , \47466_nG173e0 , \47467_nG173e1 , \47468 , \47469_nG19035 , \47470 , \47471 , \47472_nG173e2 , \47473_nG173e3 , \47474 ,
         \47475_nG173e4 , \47476_nG173e5 , \47477 , \47478_nG19037 , \47479 , \47480 , \47481_nG173e6 , \47482_nG173e7 , \47483 , \47484_nG173e8 ,
         \47485_nG173e9 , \47486 , \47487_nG19039 , \47488 , \47489 , \47490_nG173ea , \47491_nG173eb , \47492 , \47493_nG173ec , \47494_nG173ed ,
         \47495 , \47496_nG1903b , \47497 , \47498 , \47499_nG173ee , \47500_nG173ef , \47501 , \47502_nG173f0 , \47503_nG173f1 , \47504 ,
         \47505_nG1903d , \47506 , \47507 , \47508_nG173f2 , \47509_nG173f3 , \47510 , \47511_nG173f4 , \47512_nG173f5 , \47513 , \47514_nG1903f ,
         \47515 , \47516 , \47517_nG173f6 , \47518_nG173f7 , \47519 , \47520_nG173f8 , \47521_nG173f9 , \47522 , \47523_nG19041 , \47524 ,
         \47525 , \47526_nG173fa , \47527_nG173fb , \47528 , \47529_nG173fc , \47530_nG173fd , \47531 , \47532_nG19045 , \47533 , \47534 ,
         \47535_nG173fe , \47536_nG173ff , \47537 , \47538_nG17400 , \47539_nG17401 , \47540 , \47541_nG19047 , \47542 , \47543 , \47544_nG17402 ,
         \47545_nG17403 , \47546 , \47547_nG17404 , \47548_nG17405 , \47549 , \47550_nG19049 , \47551 , \47552 , \47553_nG17406 , \47554_nG17407 ,
         \47555 , \47556_nG17408 , \47557_nG17409 , \47558 , \47559_nG1904b , \47560 , \47561 , \47562_nG1740a , \47563_nG1740b , \47564 ,
         \47565_nG1740c , \47566_nG1740d , \47567 , \47568_nG1904d , \47569 , \47570 , \47571_nG1740e , \47572_nG1740f , \47573 , \47574_nG17410 ,
         \47575_nG17411 , \47576 , \47577_nG1904f , \47578 , \47579 , \47580_nG17412 , \47581_nG17413 , \47582 , \47583_nG17414 , \47584_nG17415 ,
         \47585 , \47586_nG19051 , \47587 , \47588 , \47589_nG17416 , \47590_nG17417 , \47591 , \47592_nG17418 , \47593_nG17419 , \47594 ,
         \47595_nG19053 , \47596 , \47597 , \47598_nG1741a , \47599_nG1741b , \47600 , \47601_nG1741c , \47602_nG1741d , \47603 , \47604_nG19055 ,
         \47605 , \47606 , \47607_nG1741e , \47608_nG1741f , \47609 , \47610_nG17420 , \47611_nG17421 , \47612 , \47613_nG19057 , \47614 ,
         \47615 , \47616_nG17422 , \47617_nG17423 , \47618 , \47619_nG17424 , \47620_nG17425 , \47621 , \47622_nG1905b , \47623 , \47624 ,
         \47625_nG17426 , \47626_nG17427 , \47627 , \47628_nG17428 , \47629_nG17429 , \47630 , \47631_nG1905d , \47632 , \47633 , \47634_nG1742a ,
         \47635_nG1742b , \47636 , \47637_nG1742c , \47638_nG1742d , \47639 , \47640_nG1905f , \47641 , \47642 , \47643_nG1742e , \47644_nG1742f ,
         \47645 , \47646_nG17430 , \47647_nG17431 , \47648 , \47649_nG19061 , \47650 , \47651 , \47652_nG17432 , \47653_nG17433 , \47654 ,
         \47655_nG17434 , \47656_nG17435 , \47657 , \47658_nG19063 , \47659 , \47660 , \47661_nG17436 , \47662_nG17437 , \47663 , \47664_nG17438 ,
         \47665_nG17439 , \47666 , \47667_nG19065 , \47668 , \47669 , \47670_nG1743a , \47671_nG1743b , \47672 , \47673_nG1743c , \47674_nG1743d ,
         \47675 , \47676_nG19067 , \47677 , \47678 , \47679_nG1743e , \47680_nG1743f , \47681 , \47682_nG17440 , \47683_nG17441 , \47684 ,
         \47685_nG19069 , \47686 , \47687 , \47688_nG17442 , \47689_nG17443 , \47690 , \47691_nG17444 , \47692_nG17445 , \47693 , \47694_nG1906b ,
         \47695 , \47696 , \47697_nG17446 , \47698_nG17447 , \47699 , \47700_nG17448 , \47701_nG17449 , \47702 , \47703_nG1906d , \47704 ,
         \47705 , \47706_nG1744a , \47707_nG1744b , \47708 , \47709_nG1744c , \47710_nG1744d , \47711 , \47712_nG19071 , \47713 , \47714 ,
         \47715_nG1744e , \47716_nG1744f , \47717 , \47718_nG17450 , \47719_nG17451 , \47720 , \47721_nG19073 , \47722 , \47723 , \47724_nG17452 ,
         \47725_nG17453 , \47726 , \47727_nG17454 , \47728_nG17455 , \47729 , \47730_nG19075 , \47731 , \47732 , \47733_nG17456 , \47734_nG17457 ,
         \47735 , \47736_nG17458 , \47737_nG17459 , \47738 , \47739_nG19077 , \47740 , \47741 , \47742_nG1745a , \47743_nG1745b , \47744 ,
         \47745_nG1745c , \47746_nG1745d , \47747 , \47748_nG19079 , \47749 , \47750 , \47751 , \47752_nG1725c , \47753_nG1725d , \47754 ,
         \47755 , \47756_nG1725f , \47757_nG17260 , \47758 , \47759_nG18f81 , \47760 , \47761_nG17261 , \47762_nG17262 , \47763_nG17263 , \47764_nG17264 ,
         \47765 , \47766_nG18f97 , \47767 , \47768_nG17265 , \47769_nG17266 , \47770_nG17267 , \47771_nG17268 , \47772 , \47773_nG18fad , \47774 ,
         \47775_nG17269 , \47776_nG1726a , \47777_nG1726b , \47778_nG1726c , \47779 , \47780_nG18fc3 , \47781 , \47782_nG1726d , \47783_nG1726e , \47784_nG1726f ,
         \47785_nG17270 , \47786 , \47787_nG18fd9 , \47788 , \47789_nG17271 , \47790_nG17272 , \47791_nG17273 , \47792_nG17274 , \47793 , \47794_nG18fef ,
         \47795 , \47796_nG17275 , \47797_nG17276 , \47798_nG17277 , \47799_nG17278 , \47800 , \47801_nG18ffb , \47802 , \47803_nG17279 , \47804_nG1727a ,
         \47805_nG1727b , \47806_nG1727c , \47807 , \47808_nG18ffd , \47809 , \47810_nG1727d , \47811_nG1727e , \47812_nG1727f , \47813_nG17280 , \47814 ,
         \47815_nG18fff , \47816 , \47817_nG17281 , \47818_nG17282 , \47819_nG17283 , \47820_nG17284 , \47821 , \47822_nG18f83 , \47823 , \47824_nG17285 ,
         \47825_nG17286 , \47826_nG17287 , \47827_nG17288 , \47828 , \47829_nG18f85 , \47830 , \47831_nG17289 , \47832_nG1728a , \47833_nG1728b , \47834_nG1728c ,
         \47835 , \47836_nG18f87 , \47837 , \47838_nG1728d , \47839_nG1728e , \47840_nG1728f , \47841_nG17290 , \47842 , \47843_nG18f89 , \47844 ,
         \47845_nG17291 , \47846_nG17292 , \47847_nG17293 , \47848_nG17294 , \47849 , \47850_nG18f8b , \47851 , \47852_nG17295 , \47853_nG17296 , \47854_nG17297 ,
         \47855_nG17298 , \47856 , \47857_nG18f8d , \47858 , \47859_nG17299 , \47860_nG1729a , \47861_nG1729b , \47862_nG1729c , \47863 , \47864_nG18f8f ,
         \47865 , \47866_nG1729d , \47867_nG1729e , \47868_nG1729f , \47869_nG172a0 , \47870 , \47871_nG18f91 , \47872 , \47873_nG172a1 , \47874_nG172a2 ,
         \47875_nG172a3 , \47876_nG172a4 , \47877 , \47878_nG18f93 , \47879 , \47880_nG172a5 , \47881_nG172a6 , \47882_nG172a7 , \47883_nG172a8 , \47884 ,
         \47885_nG18f95 , \47886 , \47887_nG172a9 , \47888_nG172aa , \47889_nG172ab , \47890_nG172ac , \47891 , \47892_nG18f99 , \47893 , \47894_nG172ad ,
         \47895_nG172ae , \47896_nG172af , \47897_nG172b0 , \47898 , \47899_nG18f9b , \47900 , \47901_nG172b1 , \47902_nG172b2 , \47903_nG172b3 , \47904_nG172b4 ,
         \47905 , \47906_nG18f9d , \47907 , \47908_nG172b5 , \47909_nG172b6 , \47910_nG172b7 , \47911_nG172b8 , \47912 , \47913_nG18f9f , \47914 ,
         \47915_nG172b9 , \47916_nG172ba , \47917_nG172bb , \47918_nG172bc , \47919 , \47920_nG18fa1 , \47921 , \47922_nG172bd , \47923_nG172be , \47924_nG172bf ,
         \47925_nG172c0 , \47926 , \47927_nG18fa3 , \47928 , \47929_nG172c1 , \47930_nG172c2 , \47931_nG172c3 , \47932_nG172c4 , \47933 , \47934_nG18fa5 ,
         \47935 , \47936_nG172c5 , \47937_nG172c6 , \47938_nG172c7 , \47939_nG172c8 , \47940 , \47941_nG18fa7 , \47942 , \47943_nG172c9 , \47944_nG172ca ,
         \47945_nG172cb , \47946_nG172cc , \47947 , \47948_nG18fa9 , \47949 , \47950_nG172cd , \47951_nG172ce , \47952_nG172cf , \47953_nG172d0 , \47954 ,
         \47955_nG18fab , \47956 , \47957_nG172d1 , \47958_nG172d2 , \47959_nG172d3 , \47960_nG172d4 , \47961 , \47962_nG18faf , \47963 , \47964_nG172d5 ,
         \47965_nG172d6 , \47966_nG172d7 , \47967_nG172d8 , \47968 , \47969_nG18fb1 , \47970 , \47971_nG172d9 , \47972_nG172da , \47973_nG172db , \47974_nG172dc ,
         \47975 , \47976_nG18fb3 , \47977 , \47978_nG172dd , \47979_nG172de , \47980_nG172df , \47981_nG172e0 , \47982 , \47983_nG18fb5 , \47984 ,
         \47985_nG172e1 , \47986_nG172e2 , \47987_nG172e3 , \47988_nG172e4 , \47989 , \47990_nG18fb7 , \47991 , \47992_nG172e5 , \47993_nG172e6 , \47994_nG172e7 ,
         \47995_nG172e8 , \47996 , \47997_nG18fb9 , \47998 , \47999_nG172e9 , \48000_nG172ea , \48001_nG172eb , \48002_nG172ec , \48003 , \48004_nG18fbb ,
         \48005 , \48006_nG172ed , \48007_nG172ee , \48008_nG172ef , \48009_nG172f0 , \48010 , \48011_nG18fbd , \48012 , \48013_nG172f1 , \48014_nG172f2 ,
         \48015_nG172f3 , \48016_nG172f4 , \48017 , \48018_nG18fbf , \48019 , \48020_nG172f5 , \48021_nG172f6 , \48022_nG172f7 , \48023_nG172f8 , \48024 ,
         \48025_nG18fc1 , \48026 , \48027_nG172f9 , \48028_nG172fa , \48029_nG172fb , \48030_nG172fc , \48031 , \48032_nG18fc5 , \48033 , \48034_nG172fd ,
         \48035_nG172fe , \48036_nG172ff , \48037_nG17300 , \48038 , \48039_nG18fc7 , \48040 , \48041_nG17301 , \48042_nG17302 , \48043_nG17303 , \48044_nG17304 ,
         \48045 , \48046_nG18fc9 , \48047 , \48048_nG17305 , \48049_nG17306 , \48050_nG17307 , \48051_nG17308 , \48052 , \48053_nG18fcb , \48054 ,
         \48055_nG17309 , \48056_nG1730a , \48057_nG1730b , \48058_nG1730c , \48059 , \48060_nG18fcd , \48061 , \48062_nG1730d , \48063_nG1730e , \48064_nG1730f ,
         \48065_nG17310 , \48066 , \48067_nG18fcf , \48068 , \48069_nG17311 , \48070_nG17312 , \48071_nG17313 , \48072_nG17314 , \48073 , \48074_nG18fd1 ,
         \48075 , \48076_nG17315 , \48077_nG17316 , \48078_nG17317 , \48079_nG17318 , \48080 , \48081_nG18fd3 , \48082 , \48083_nG17319 , \48084_nG1731a ,
         \48085_nG1731b , \48086_nG1731c , \48087 , \48088_nG18fd5 , \48089 , \48090_nG1731d , \48091_nG1731e , \48092_nG1731f , \48093_nG17320 , \48094 ,
         \48095_nG18fd7 , \48096 , \48097_nG17321 , \48098_nG17322 , \48099_nG17323 , \48100_nG17324 , \48101 , \48102_nG18fdb , \48103 , \48104_nG17325 ,
         \48105_nG17326 , \48106_nG17327 , \48107_nG17328 , \48108 , \48109_nG18fdd , \48110 , \48111_nG17329 , \48112_nG1732a , \48113_nG1732b , \48114_nG1732c ,
         \48115 , \48116_nG18fdf , \48117 , \48118_nG1732d , \48119_nG1732e , \48120_nG1732f , \48121_nG17330 , \48122 , \48123_nG18fe1 , \48124 ,
         \48125_nG17331 , \48126_nG17332 , \48127_nG17333 , \48128_nG17334 , \48129 , \48130_nG18fe3 , \48131 , \48132_nG17335 , \48133_nG17336 , \48134_nG17337 ,
         \48135_nG17338 , \48136 , \48137_nG18fe5 , \48138 , \48139_nG17339 , \48140_nG1733a , \48141_nG1733b , \48142_nG1733c , \48143 , \48144_nG18fe7 ,
         \48145 , \48146_nG1733d , \48147_nG1733e , \48148_nG1733f , \48149_nG17340 , \48150 , \48151_nG18fe9 , \48152 , \48153_nG17341 , \48154_nG17342 ,
         \48155_nG17343 , \48156_nG17344 , \48157 , \48158_nG18feb , \48159 , \48160_nG17345 , \48161_nG17346 , \48162_nG17347 , \48163_nG17348 , \48164 ,
         \48165_nG18fed , \48166 , \48167_nG17349 , \48168_nG1734a , \48169_nG1734b , \48170_nG1734c , \48171 , \48172_nG18ff1 , \48173 , \48174_nG1734d ,
         \48175_nG1734e , \48176_nG1734f , \48177_nG17350 , \48178 , \48179_nG18ff3 , \48180 , \48181_nG17351 , \48182_nG17352 , \48183_nG17353 , \48184_nG17354 ,
         \48185 , \48186_nG18ff5 , \48187 , \48188_nG17355 , \48189_nG17356 , \48190_nG17357 , \48191_nG17358 , \48192 , \48193_nG18ff7 , \48194 ,
         \48195_nG17359 , \48196_nG1735a , \48197_nG1735b , \48198_nG1735c , \48199 , \48200_nG18ff9 , \48201 , \48202 , \48203_nG1715a , \48204_nG1715b ,
         \48205 , \48206_nG1715e , \48207_nG1715f , \48208 , \48209_nG18f01 , \48210 , \48211_nG17160 , \48212_nG17161 , \48213_nG17162 , \48214_nG17163 ,
         \48215 , \48216_nG18f17 , \48217 , \48218_nG17164 , \48219_nG17165 , \48220_nG17166 , \48221_nG17167 , \48222 , \48223_nG18f2d , \48224 ,
         \48225_nG17168 , \48226_nG17169 , \48227_nG1716a , \48228_nG1716b , \48229 , \48230_nG18f43 , \48231 , \48232_nG1716c , \48233_nG1716d , \48234_nG1716e ,
         \48235_nG1716f , \48236 , \48237_nG18f59 , \48238 , \48239_nG17170 , \48240_nG17171 , \48241_nG17172 , \48242_nG17173 , \48243 , \48244_nG18f6f ,
         \48245 , \48246_nG17174 , \48247_nG17175 , \48248_nG17176 , \48249_nG17177 , \48250 , \48251_nG18f7b , \48252 , \48253_nG17178 , \48254_nG17179 ,
         \48255_nG1717a , \48256_nG1717b , \48257 , \48258_nG18f7d , \48259 , \48260_nG1717c , \48261_nG1717d , \48262_nG1717e , \48263_nG1717f , \48264 ,
         \48265_nG18f7f , \48266 , \48267_nG17180 , \48268_nG17181 , \48269_nG17182 , \48270_nG17183 , \48271 , \48272_nG18f03 , \48273 , \48274_nG17184 ,
         \48275_nG17185 , \48276_nG17186 , \48277_nG17187 , \48278 , \48279_nG18f05 , \48280 , \48281_nG17188 , \48282_nG17189 , \48283_nG1718a , \48284_nG1718b ,
         \48285 , \48286_nG18f07 , \48287 , \48288_nG1718c , \48289_nG1718d , \48290_nG1718e , \48291_nG1718f , \48292 , \48293_nG18f09 , \48294 ,
         \48295_nG17190 , \48296_nG17191 , \48297_nG17192 , \48298_nG17193 , \48299 , \48300_nG18f0b , \48301 , \48302_nG17194 , \48303_nG17195 , \48304_nG17196 ,
         \48305_nG17197 , \48306 , \48307_nG18f0d , \48308 , \48309_nG17198 , \48310_nG17199 , \48311_nG1719a , \48312_nG1719b , \48313 , \48314_nG18f0f ,
         \48315 , \48316_nG1719c , \48317_nG1719d , \48318_nG1719e , \48319_nG1719f , \48320 , \48321_nG18f11 , \48322 , \48323_nG171a0 , \48324_nG171a1 ,
         \48325_nG171a2 , \48326_nG171a3 , \48327 , \48328_nG18f13 , \48329 , \48330_nG171a4 , \48331_nG171a5 , \48332_nG171a6 , \48333_nG171a7 , \48334 ,
         \48335_nG18f15 , \48336 , \48337_nG171a8 , \48338_nG171a9 , \48339_nG171aa , \48340_nG171ab , \48341 , \48342_nG18f19 , \48343 , \48344_nG171ac ,
         \48345_nG171ad , \48346_nG171ae , \48347_nG171af , \48348 , \48349_nG18f1b , \48350 , \48351_nG171b0 , \48352_nG171b1 , \48353_nG171b2 , \48354_nG171b3 ,
         \48355 , \48356_nG18f1d , \48357 , \48358_nG171b4 , \48359_nG171b5 , \48360_nG171b6 , \48361_nG171b7 , \48362 , \48363_nG18f1f , \48364 ,
         \48365_nG171b8 , \48366_nG171b9 , \48367_nG171ba , \48368_nG171bb , \48369 , \48370_nG18f21 , \48371 , \48372_nG171bc , \48373_nG171bd , \48374_nG171be ,
         \48375_nG171bf , \48376 , \48377_nG18f23 , \48378 , \48379_nG171c0 , \48380_nG171c1 , \48381_nG171c2 , \48382_nG171c3 , \48383 , \48384_nG18f25 ,
         \48385 , \48386_nG171c4 , \48387_nG171c5 , \48388_nG171c6 , \48389_nG171c7 , \48390 , \48391_nG18f27 , \48392 , \48393_nG171c8 , \48394_nG171c9 ,
         \48395_nG171ca , \48396_nG171cb , \48397 , \48398_nG18f29 , \48399 , \48400_nG171cc , \48401_nG171cd , \48402_nG171ce , \48403_nG171cf , \48404 ,
         \48405_nG18f2b , \48406 , \48407_nG171d0 , \48408_nG171d1 , \48409_nG171d2 , \48410_nG171d3 , \48411 , \48412_nG18f2f , \48413 , \48414_nG171d4 ,
         \48415_nG171d5 , \48416_nG171d6 , \48417_nG171d7 , \48418 , \48419_nG18f31 , \48420 , \48421_nG171d8 , \48422_nG171d9 , \48423_nG171da , \48424_nG171db ,
         \48425 , \48426_nG18f33 , \48427 , \48428_nG171dc , \48429_nG171dd , \48430_nG171de , \48431_nG171df , \48432 , \48433_nG18f35 , \48434 ,
         \48435_nG171e0 , \48436_nG171e1 , \48437_nG171e2 , \48438_nG171e3 , \48439 , \48440_nG18f37 , \48441 , \48442_nG171e4 , \48443_nG171e5 , \48444_nG171e6 ,
         \48445_nG171e7 , \48446 , \48447_nG18f39 , \48448 , \48449_nG171e8 , \48450_nG171e9 , \48451_nG171ea , \48452_nG171eb , \48453 , \48454_nG18f3b ,
         \48455 , \48456_nG171ec , \48457_nG171ed , \48458_nG171ee , \48459_nG171ef , \48460 , \48461_nG18f3d , \48462 , \48463_nG171f0 , \48464_nG171f1 ,
         \48465_nG171f2 , \48466_nG171f3 , \48467 , \48468_nG18f3f , \48469 , \48470_nG171f4 , \48471_nG171f5 , \48472_nG171f6 , \48473_nG171f7 , \48474 ,
         \48475_nG18f41 , \48476 , \48477_nG171f8 , \48478_nG171f9 , \48479_nG171fa , \48480_nG171fb , \48481 , \48482_nG18f45 , \48483 , \48484_nG171fc ,
         \48485_nG171fd , \48486_nG171fe , \48487_nG171ff , \48488 , \48489_nG18f47 , \48490 , \48491_nG17200 , \48492_nG17201 , \48493_nG17202 , \48494_nG17203 ,
         \48495 , \48496_nG18f49 , \48497 , \48498_nG17204 , \48499_nG17205 , \48500_nG17206 , \48501_nG17207 , \48502 , \48503_nG18f4b , \48504 ,
         \48505_nG17208 , \48506_nG17209 , \48507_nG1720a , \48508_nG1720b , \48509 , \48510_nG18f4d , \48511 , \48512_nG1720c , \48513_nG1720d , \48514_nG1720e ,
         \48515_nG1720f , \48516 , \48517_nG18f4f , \48518 , \48519_nG17210 , \48520_nG17211 , \48521_nG17212 , \48522_nG17213 , \48523 , \48524_nG18f51 ,
         \48525 , \48526_nG17214 , \48527_nG17215 , \48528_nG17216 , \48529_nG17217 , \48530 , \48531_nG18f53 , \48532 , \48533_nG17218 , \48534_nG17219 ,
         \48535_nG1721a , \48536_nG1721b , \48537 , \48538_nG18f55 , \48539 , \48540_nG1721c , \48541_nG1721d , \48542_nG1721e , \48543_nG1721f , \48544 ,
         \48545_nG18f57 , \48546 , \48547_nG17220 , \48548_nG17221 , \48549_nG17222 , \48550_nG17223 , \48551 , \48552_nG18f5b , \48553 , \48554_nG17224 ,
         \48555_nG17225 , \48556_nG17226 , \48557_nG17227 , \48558 , \48559_nG18f5d , \48560 , \48561_nG17228 , \48562_nG17229 , \48563_nG1722a , \48564_nG1722b ,
         \48565 , \48566_nG18f5f , \48567 , \48568_nG1722c , \48569_nG1722d , \48570_nG1722e , \48571_nG1722f , \48572 , \48573_nG18f61 , \48574 ,
         \48575_nG17230 , \48576_nG17231 , \48577_nG17232 , \48578_nG17233 , \48579 , \48580_nG18f63 , \48581 , \48582_nG17234 , \48583_nG17235 , \48584_nG17236 ,
         \48585_nG17237 , \48586 , \48587_nG18f65 , \48588 , \48589_nG17238 , \48590_nG17239 , \48591_nG1723a , \48592_nG1723b , \48593 , \48594_nG18f67 ,
         \48595 , \48596_nG1723c , \48597_nG1723d , \48598_nG1723e , \48599_nG1723f , \48600 , \48601_nG18f69 , \48602 , \48603_nG17240 , \48604_nG17241 ,
         \48605_nG17242 , \48606_nG17243 , \48607 , \48608_nG18f6b , \48609 , \48610_nG17244 , \48611_nG17245 , \48612_nG17246 , \48613_nG17247 , \48614 ,
         \48615_nG18f6d , \48616 , \48617_nG17248 , \48618_nG17249 , \48619_nG1724a , \48620_nG1724b , \48621 , \48622_nG18f71 , \48623 , \48624_nG1724c ,
         \48625_nG1724d , \48626_nG1724e , \48627_nG1724f , \48628 , \48629_nG18f73 , \48630 , \48631_nG17250 , \48632_nG17251 , \48633_nG17252 , \48634_nG17253 ,
         \48635 , \48636_nG18f75 , \48637 , \48638_nG17254 , \48639_nG17255 , \48640_nG17256 , \48641_nG17257 , \48642 , \48643_nG18f77 , \48644 ,
         \48645_nG17258 , \48646_nG17259 , \48647_nG1725a , \48648_nG1725b , \48649 , \48650_nG18f79 , \48651 , \48652 , \48653_nG16fd8 , \48654_nG16fd9 ,
         \48655 , \48656_nG16fde , \48657_nG16fdf , \48658 , \48659_nG18e81 , \48660 , \48661_nG16fe1 , \48662_nG16fe2 , \48663_nG16fe4 , \48664_nG16fe5 ,
         \48665 , \48666_nG18e97 , \48667 , \48668_nG16fe7 , \48669_nG16fe8 , \48670_nG16fea , \48671_nG16feb , \48672 , \48673_nG18ead , \48674 ,
         \48675_nG16fed , \48676_nG16fee , \48677_nG16ff0 , \48678_nG16ff1 , \48679 , \48680_nG18ec3 , \48681 , \48682_nG16ff3 , \48683_nG16ff4 , \48684_nG16ff6 ,
         \48685_nG16ff7 , \48686 , \48687_nG18ed9 , \48688 , \48689_nG16ff9 , \48690_nG16ffa , \48691_nG16ffc , \48692_nG16ffd , \48693 , \48694_nG18eef ,
         \48695 , \48696_nG16fff , \48697_nG17000 , \48698_nG17002 , \48699_nG17003 , \48700 , \48701_nG18efb , \48702 , \48703_nG17005 , \48704_nG17006 ,
         \48705_nG17008 , \48706_nG17009 , \48707 , \48708_nG18efd , \48709 , \48710_nG1700b , \48711_nG1700c , \48712_nG1700e , \48713_nG1700f , \48714 ,
         \48715_nG18eff , \48716 , \48717_nG17011 , \48718_nG17012 , \48719_nG17014 , \48720_nG17015 , \48721 , \48722_nG18e83 , \48723 , \48724_nG17017 ,
         \48725_nG17018 , \48726_nG1701a , \48727_nG1701b , \48728 , \48729_nG18e85 , \48730 , \48731_nG1701d , \48732_nG1701e , \48733_nG17020 , \48734_nG17021 ,
         \48735 , \48736_nG18e87 , \48737 , \48738_nG17023 , \48739_nG17024 , \48740_nG17026 , \48741_nG17027 , \48742 , \48743_nG18e89 , \48744 ,
         \48745_nG17029 , \48746_nG1702a , \48747_nG1702c , \48748_nG1702d , \48749 , \48750_nG18e8b , \48751 , \48752_nG1702f , \48753_nG17030 , \48754_nG17032 ,
         \48755_nG17033 , \48756 , \48757_nG18e8d , \48758 , \48759_nG17035 , \48760_nG17036 , \48761_nG17038 , \48762_nG17039 , \48763 , \48764_nG18e8f ,
         \48765 , \48766_nG1703b , \48767_nG1703c , \48768_nG1703e , \48769_nG1703f , \48770 , \48771_nG18e91 , \48772 , \48773_nG17041 , \48774_nG17042 ,
         \48775_nG17044 , \48776_nG17045 , \48777 , \48778_nG18e93 , \48779 , \48780_nG17047 , \48781_nG17048 , \48782_nG1704a , \48783_nG1704b , \48784 ,
         \48785_nG18e95 , \48786 , \48787_nG1704d , \48788_nG1704e , \48789_nG17050 , \48790_nG17051 , \48791 , \48792_nG18e99 , \48793 , \48794_nG17053 ,
         \48795_nG17054 , \48796_nG17056 , \48797_nG17057 , \48798 , \48799_nG18e9b , \48800 , \48801_nG17059 , \48802_nG1705a , \48803_nG1705c , \48804_nG1705d ,
         \48805 , \48806_nG18e9d , \48807 , \48808_nG1705f , \48809_nG17060 , \48810_nG17062 , \48811_nG17063 , \48812 , \48813_nG18e9f , \48814 ,
         \48815_nG17065 , \48816_nG17066 , \48817_nG17068 , \48818_nG17069 , \48819 , \48820_nG18ea1 , \48821 , \48822_nG1706b , \48823_nG1706c , \48824_nG1706e ,
         \48825_nG1706f , \48826 , \48827_nG18ea3 , \48828 , \48829_nG17071 , \48830_nG17072 , \48831_nG17074 , \48832_nG17075 , \48833 , \48834_nG18ea5 ,
         \48835 , \48836_nG17077 , \48837_nG17078 , \48838_nG1707a , \48839_nG1707b , \48840 , \48841_nG18ea7 , \48842 , \48843_nG1707d , \48844_nG1707e ,
         \48845_nG17080 , \48846_nG17081 , \48847 , \48848_nG18ea9 , \48849 , \48850_nG17083 , \48851_nG17084 , \48852_nG17086 , \48853_nG17087 , \48854 ,
         \48855_nG18eab , \48856 , \48857_nG17089 , \48858_nG1708a , \48859_nG1708c , \48860_nG1708d , \48861 , \48862_nG18eaf , \48863 , \48864_nG1708f ,
         \48865_nG17090 , \48866_nG17092 , \48867_nG17093 , \48868 , \48869_nG18eb1 , \48870 , \48871_nG17095 , \48872_nG17096 , \48873_nG17098 , \48874_nG17099 ,
         \48875 , \48876_nG18eb3 , \48877 , \48878_nG1709b , \48879_nG1709c , \48880_nG1709e , \48881_nG1709f , \48882 , \48883_nG18eb5 , \48884 ,
         \48885_nG170a1 , \48886_nG170a2 , \48887_nG170a4 , \48888_nG170a5 , \48889 , \48890_nG18eb7 , \48891 , \48892_nG170a7 , \48893_nG170a8 , \48894_nG170aa ,
         \48895_nG170ab , \48896 , \48897_nG18eb9 , \48898 , \48899_nG170ad , \48900_nG170ae , \48901_nG170b0 , \48902_nG170b1 , \48903 , \48904_nG18ebb ,
         \48905 , \48906_nG170b3 , \48907_nG170b4 , \48908_nG170b6 , \48909_nG170b7 , \48910 , \48911_nG18ebd , \48912 , \48913_nG170b9 , \48914_nG170ba ,
         \48915_nG170bc , \48916_nG170bd , \48917 , \48918_nG18ebf , \48919 , \48920_nG170bf , \48921_nG170c0 , \48922_nG170c2 , \48923_nG170c3 , \48924 ,
         \48925_nG18ec1 , \48926 , \48927_nG170c5 , \48928_nG170c6 , \48929_nG170c8 , \48930_nG170c9 , \48931 , \48932_nG18ec5 , \48933 , \48934_nG170cb ,
         \48935_nG170cc , \48936_nG170ce , \48937_nG170cf , \48938 , \48939_nG18ec7 , \48940 , \48941_nG170d1 , \48942_nG170d2 , \48943_nG170d4 , \48944_nG170d5 ,
         \48945 , \48946_nG18ec9 , \48947 , \48948_nG170d7 , \48949_nG170d8 , \48950_nG170da , \48951_nG170db , \48952 , \48953_nG18ecb , \48954 ,
         \48955_nG170dd , \48956_nG170de , \48957_nG170e0 , \48958_nG170e1 , \48959 , \48960_nG18ecd , \48961 , \48962_nG170e3 , \48963_nG170e4 , \48964_nG170e6 ,
         \48965_nG170e7 , \48966 , \48967_nG18ecf , \48968 , \48969_nG170e9 , \48970_nG170ea , \48971_nG170ec , \48972_nG170ed , \48973 , \48974_nG18ed1 ,
         \48975 , \48976_nG170ef , \48977_nG170f0 , \48978_nG170f2 , \48979_nG170f3 , \48980 , \48981_nG18ed3 , \48982 , \48983_nG170f5 , \48984_nG170f6 ,
         \48985_nG170f8 , \48986_nG170f9 , \48987 , \48988_nG18ed5 , \48989 , \48990_nG170fb , \48991_nG170fc , \48992_nG170fe , \48993_nG170ff , \48994 ,
         \48995_nG18ed7 , \48996 , \48997_nG17101 , \48998_nG17102 , \48999_nG17104 , \49000_nG17105 , \49001 , \49002_nG18edb , \49003 , \49004_nG17107 ,
         \49005_nG17108 , \49006_nG1710a , \49007_nG1710b , \49008 , \49009_nG18edd , \49010 , \49011_nG1710d , \49012_nG1710e , \49013_nG17110 , \49014_nG17111 ,
         \49015 , \49016_nG18edf , \49017 , \49018_nG17113 , \49019_nG17114 , \49020_nG17116 , \49021_nG17117 , \49022 , \49023_nG18ee1 , \49024 ,
         \49025_nG17119 , \49026_nG1711a , \49027_nG1711c , \49028_nG1711d , \49029 , \49030_nG18ee3 , \49031 , \49032_nG1711f , \49033_nG17120 , \49034_nG17122 ,
         \49035_nG17123 , \49036 , \49037_nG18ee5 , \49038 , \49039_nG17125 , \49040_nG17126 , \49041_nG17128 , \49042_nG17129 , \49043 , \49044_nG18ee7 ,
         \49045 , \49046_nG1712b , \49047_nG1712c , \49048_nG1712e , \49049_nG1712f , \49050 , \49051_nG18ee9 , \49052 , \49053_nG17131 , \49054_nG17132 ,
         \49055_nG17134 , \49056_nG17135 , \49057 , \49058_nG18eeb , \49059 , \49060_nG17137 , \49061_nG17138 , \49062_nG1713a , \49063_nG1713b , \49064 ,
         \49065_nG18eed , \49066 , \49067_nG1713d , \49068_nG1713e , \49069_nG17140 , \49070_nG17141 , \49071 , \49072_nG18ef1 , \49073 , \49074_nG17143 ,
         \49075_nG17144 , \49076_nG17146 , \49077_nG17147 , \49078 , \49079_nG18ef3 , \49080 , \49081_nG17149 , \49082_nG1714a , \49083_nG1714c , \49084_nG1714d ,
         \49085 , \49086_nG18ef5 , \49087 , \49088_nG1714f , \49089_nG17150 , \49090_nG17152 , \49091_nG17153 , \49092 , \49093_nG18ef7 , \49094 ,
         \49095_nG17155 , \49096_nG17156 , \49097_nG17158 , \49098_nG17159 , \49099 , \49100_nG18ef9 , \49101 , \49102 , \49103_nG16faa , \49104 ,
         \49105 , \49106_nG16fab , \49107 , \49108_nG18e69 , \49109 , \49110 , \49111_nG16fac , \49112_nG16fad , \49113 , \49114_nG18e6b ,
         \49115 , \49116 , \49117_nG16fae , \49118_nG16faf , \49119 , \49120_nG18e6d , \49121 , \49122 , \49123_nG16fb0 , \49124_nG16fb1 ,
         \49125 , \49126_nG18e6f , \49127 , \49128 , \49129_nG16fb2 , \49130_nG16fb3 , \49131 , \49132_nG18e71 , \49133 , \49134 ,
         \49135_nG16fb4 , \49136_nG16fb5 , \49137 , \49138_nG18e73 , \49139 , \49140 , \49141_nG16fb6 , \49142_nG16fb7 , \49143 , \49144_nG18e75 ,
         \49145 , \49146 , \49147_nG16fb8 , \49148_nG16fb9 , \49149 , \49150_nG18e77 , \49151 , \49152_nG16f99 , \49153_nG16f9a , \49154 ,
         \49155_nG18e59 , \49156 , \49157_nG16f9b , \49158_nG16f9c , \49159 , \49160_nG18e5b , \49161 , \49162_nG16f9d , \49163_nG16f9e , \49164 ,
         \49165_nG18e5d , \49166 , \49167_nG16f9f , \49168_nG16fa0 , \49169 , \49170_nG18e5f , \49171 , \49172_nG16fa1 , \49173_nG16fa2 , \49174 ,
         \49175_nG18e61 , \49176 , \49177_nG16fa3 , \49178_nG16fa4 , \49179 , \49180_nG18e63 , \49181 , \49182_nG16fa5 , \49183_nG16fa6 , \49184 ,
         \49185_nG18e65 , \49186 , \49187_nG16fa7 , \49188_nG16fa8 , \49189 , \49190_nG18e67 , \49191 , \49192_nG16f88 , \49193_nG16f89 , \49194 ,
         \49195_nG18e49 , \49196 , \49197_nG16f8a , \49198_nG16f8b , \49199 , \49200_nG18e4b , \49201 , \49202_nG16f8c , \49203_nG16f8d , \49204 ,
         \49205_nG18e4d , \49206 , \49207_nG16f8e , \49208_nG16f8f , \49209 , \49210_nG18e4f , \49211 , \49212_nG16f90 , \49213_nG16f91 , \49214 ,
         \49215_nG18e51 , \49216 , \49217_nG16f92 , \49218_nG16f93 , \49219 , \49220_nG18e53 , \49221 , \49222_nG16f94 , \49223_nG16f95 , \49224 ,
         \49225_nG18e55 , \49226 , \49227_nG16f96 , \49228_nG16f97 , \49229 , \49230_nG18e57 , \49231 , \49232_nG16f67 , \49233_nG16f70 , \49234 ,
         \49235_nG19081 , \49236 , \49237_nG16f72 , \49238_nG16f73 , \49239 , \49240_nG19083 , \49241 , \49242_nG16f75 , \49243_nG16f76 , \49244 ,
         \49245_nG19085 , \49246 , \49247_nG16f78 , \49248_nG16f79 , \49249 , \49250_nG19087 , \49251 , \49252_nG16f7b , \49253_nG16f7c , \49254 ,
         \49255_nG19089 , \49256 , \49257_nG16f7e , \49258_nG16f7f , \49259 , \49260_nG1908b , \49261 , \49262_nG16f81 , \49263_nG16f82 , \49264 ,
         \49265_nG1908d , \49266 , \49267_nG16f84 , \49268_nG16f85 , \49269 , \49270_nG1908f , \49271 , \49272 , \49273 , \49274 ,
         \49275_nG16e5c , \49276 , \49277_nG19090 , \49278 , \49279 , \49280_nG16ec9 , \49281 , \49282_nG18e2d , \49283 , \49284 ,
         \49285_nG16ecb , \49286 , \49287_nG18e2f , \49288 , \49289 , \49290_nG16ecd , \49291 , \49292_nG18e31 , \49293 , \49294 ,
         \49295_nG16ecf , \49296 , \49297_nG18e33 , \49298 , \49299 , \49300_nG16ed1 , \49301 , \49302_nG18e35 , \49303 , \49304 ,
         \49305_nG16ed3 , \49306 , \49307_nG18e37 , \49308 , \49309 , \49310_nG16ed5 , \49311 , \49312_nG18e39 , \49313 , \49314 ,
         \49315_nG16ec7 , \49316 , \49317_nG18e2b , \49318 , \49319 , \49320_nG16ebf , \49321 , \49322_nG18e23 , \49323 , \49324 ,
         \49325_nG16ec1 , \49326 , \49327_nG18e25 , \49328 , \49329 , \49330_nG16ec3 , \49331 , \49332_nG18e27 , \49333 , \49334 ,
         \49335_nG16ec5 , \49336 , \49337_nG18e29 , \49338 , \49339 , \49340 , \49341 , \49342 , \49343_nG16d2f , \49344 ,
         \49345 , \49346 , \49347 , \49348_nG16d30 , \49349 , \49350 , \49351 , \49352 , \49353 , \49354_nG16d36 ,
         \49355 , \49356_nG16d3a , \49357 , \49358 , \49359_nG16d3d , \49360 , \49361 , \49362 , \49363 , \49364 ,
         \49365_nG16d44 , \49366 , \49367 , \49368_nG16d45 , \49369 , \49370 , \49371 , \49372 , \49373_nG16d49 , \49374_nG16d4a ,
         \49375 , \49376 , \49377 , \49378_nG16d4e , \49379_nG16d4f , \49380_nG16d50 , \49381_nG16d51 , \49382_nG16d52 , \49383 , \49384 ,
         \49385 , \49386 , \49387 , \49388_nG16d57 , \49389_nG16d58 , \49390 , \49391 , \49392 , \49393 , \49394_nG16d5d ,
         \49395_nG16d5e , \49396_nG16d5f , \49397_nG16d60 , \49398_nG16d61 , \49399 , \49400 , \49401 , \49402 , \49403 , \49404 ,
         \49405 , \49406 , \49407 , \49408 , \49409 , \49410 , \49411 , \49412_nG16d26 , \49413_nG16d27 , \49414 ,
         \49415 , \49416 , \49417 , \49418 , \49419 , \49420 , \49421 , \49422 , \49423 , \49424 ,
         \49425 , \49426 , \49427 , \49428_nG16de4 , \49429 , \49430 , \49431 , \49432 , \49433 , \49434 ,
         \49435 , \49436_nG16de8 , \49437 , \49438 , \49439_nG16de9 , \49440 , \49441 , \49442_nG16dea , \49443 , \49444_nG16deb ,
         \49445 , \49446 , \49447 , \49448 , \49449_nG16d20 , \49450_nG16d21 , \49451 , \49452 , \49453 , \49454 ,
         \49455_nG16dd5 , \49456 , \49457 , \49458_nG16ddc , \49459_nG16ddd , \49460_nG16dde , \49461_nG16ddf , \49462 , \49463 , \49464 ,
         \49465 , \49466_nG16d19 , \49467_nG16d1c , \49468 , \49469 , \49470 , \49471 , \49472_nG16dc5 , \49473 , \49474_nG16dc9 ,
         \49475_nG16dcc , \49476_nG16dcf , \49477_nG16dd1 , \49478 , \49479 , \49480 , \49481 , \49482 , \49483 , \49484 ,
         \49485 , \49486 , \49487 , \49488 , \49489 , \49490 , \49491_nG16e60 , \49492 , \49493_nG18e47 , \49494 ,
         \49495 , \49496_nG19094 , \49497 , \49498 , \49499_nG19095 , \49500 , \49501 , \49502_nG19096 , \49503 , \49504 ,
         \49505 , \49506 , \49507 , \49508_nG16c0a , \49509 , \49510 , \49511 , \49512 , \49513 , \49514 ,
         \49515_nG16c0b , \49516 , \49517 , \49518 , \49519 , \49520_nG16c0d , \49521 , \49522 , \49523 , \49524 ,
         \49525 , \49526 , \49527_nG16c0e , \49528 , \49529_nG18d84 , \49530 , \49531 , \49532_nG16c0f , \49533_nG16c10 , \49534 ,
         \49535_nG16c11 , \49536_nG16c12 , \49537 , \49538_nG18d9a , \49539 , \49540 , \49541_nG16c13 , \49542_nG16c14 , \49543 , \49544_nG16c15 ,
         \49545_nG16c16 , \49546 , \49547_nG18db0 , \49548 , \49549 , \49550_nG16c17 , \49551_nG16c18 , \49552 , \49553_nG16c19 , \49554_nG16c1a ,
         \49555 , \49556_nG18dc6 , \49557 , \49558 , \49559_nG16c1b , \49560_nG16c1c , \49561 , \49562_nG16c1d , \49563_nG16c1e , \49564 ,
         \49565_nG18ddc , \49566 , \49567 , \49568_nG16c1f , \49569_nG16c20 , \49570 , \49571_nG16c21 , \49572_nG16c22 , \49573 , \49574_nG18df2 ,
         \49575 , \49576 , \49577_nG16c23 , \49578_nG16c24 , \49579 , \49580_nG16c25 , \49581_nG16c26 , \49582 , \49583_nG18dfe , \49584 ,
         \49585 , \49586_nG16c27 , \49587_nG16c28 , \49588 , \49589_nG16c29 , \49590_nG16c2a , \49591 , \49592_nG18e00 , \49593 , \49594 ,
         \49595_nG16c2b , \49596_nG16c2c , \49597 , \49598_nG16c2d , \49599_nG16c2e , \49600 , \49601_nG18e02 , \49602 , \49603 , \49604_nG16c2f ,
         \49605_nG16c30 , \49606 , \49607_nG16c31 , \49608_nG16c32 , \49609 , \49610_nG18d86 , \49611 , \49612 , \49613_nG16c33 , \49614_nG16c34 ,
         \49615 , \49616_nG16c35 , \49617_nG16c36 , \49618 , \49619_nG18d88 , \49620 , \49621 , \49622_nG16c37 , \49623_nG16c38 , \49624 ,
         \49625_nG16c39 , \49626_nG16c3a , \49627 , \49628_nG18d8a , \49629 , \49630 , \49631_nG16c3b , \49632_nG16c3c , \49633 , \49634_nG16c3d ,
         \49635_nG16c3e , \49636 , \49637_nG18d8c , \49638 , \49639 , \49640_nG16c3f , \49641_nG16c40 , \49642 , \49643_nG16c41 , \49644_nG16c42 ,
         \49645 , \49646_nG18d8e , \49647 , \49648 , \49649_nG16c43 , \49650_nG16c44 , \49651 , \49652_nG16c45 , \49653_nG16c46 , \49654 ,
         \49655_nG18d90 , \49656 , \49657 , \49658_nG16c47 , \49659_nG16c48 , \49660 , \49661_nG16c49 , \49662_nG16c4a , \49663 , \49664_nG18d92 ,
         \49665 , \49666 , \49667_nG16c4b , \49668_nG16c4c , \49669 , \49670_nG16c4d , \49671_nG16c4e , \49672 , \49673_nG18d94 , \49674 ,
         \49675 , \49676_nG16c4f , \49677_nG16c50 , \49678 , \49679_nG16c51 , \49680_nG16c52 , \49681 , \49682_nG18d96 , \49683 , \49684 ,
         \49685_nG16c53 , \49686_nG16c54 , \49687 , \49688_nG16c55 , \49689_nG16c56 , \49690 , \49691_nG18d98 , \49692 , \49693 , \49694_nG16c57 ,
         \49695_nG16c58 , \49696 , \49697_nG16c59 , \49698_nG16c5a , \49699 , \49700_nG18d9c , \49701 , \49702 , \49703_nG16c5b , \49704_nG16c5c ,
         \49705 , \49706_nG16c5d , \49707_nG16c5e , \49708 , \49709_nG18d9e , \49710 , \49711 , \49712_nG16c5f , \49713_nG16c60 , \49714 ,
         \49715_nG16c61 , \49716_nG16c62 , \49717 , \49718_nG18da0 , \49719 , \49720 , \49721_nG16c63 , \49722_nG16c64 , \49723 , \49724_nG16c65 ,
         \49725_nG16c66 , \49726 , \49727_nG18da2 , \49728 , \49729 , \49730_nG16c67 , \49731_nG16c68 , \49732 , \49733_nG16c69 , \49734_nG16c6a ,
         \49735 , \49736_nG18da4 , \49737 , \49738 , \49739_nG16c6b , \49740_nG16c6c , \49741 , \49742_nG16c6d , \49743_nG16c6e , \49744 ,
         \49745_nG18da6 , \49746 , \49747 , \49748_nG16c6f , \49749_nG16c70 , \49750 , \49751_nG16c71 , \49752_nG16c72 , \49753 , \49754_nG18da8 ,
         \49755 , \49756 , \49757_nG16c73 , \49758_nG16c74 , \49759 , \49760_nG16c75 , \49761_nG16c76 , \49762 , \49763_nG18daa , \49764 ,
         \49765 , \49766_nG16c77 , \49767_nG16c78 , \49768 , \49769_nG16c79 , \49770_nG16c7a , \49771 , \49772_nG18dac , \49773 , \49774 ,
         \49775_nG16c7b , \49776_nG16c7c , \49777 , \49778_nG16c7d , \49779_nG16c7e , \49780 , \49781_nG18dae , \49782 , \49783 , \49784_nG16c7f ,
         \49785_nG16c80 , \49786 , \49787_nG16c81 , \49788_nG16c82 , \49789 , \49790_nG18db2 , \49791 , \49792 , \49793_nG16c83 , \49794_nG16c84 ,
         \49795 , \49796_nG16c85 , \49797_nG16c86 , \49798 , \49799_nG18db4 , \49800 , \49801 , \49802_nG16c87 , \49803_nG16c88 , \49804 ,
         \49805_nG16c89 , \49806_nG16c8a , \49807 , \49808_nG18db6 , \49809 , \49810 , \49811_nG16c8b , \49812_nG16c8c , \49813 , \49814_nG16c8d ,
         \49815_nG16c8e , \49816 , \49817_nG18db8 , \49818 , \49819 , \49820_nG16c8f , \49821_nG16c90 , \49822 , \49823_nG16c91 , \49824_nG16c92 ,
         \49825 , \49826_nG18dba , \49827 , \49828 , \49829_nG16c93 , \49830_nG16c94 , \49831 , \49832_nG16c95 , \49833_nG16c96 , \49834 ,
         \49835_nG18dbc , \49836 , \49837 , \49838_nG16c97 , \49839_nG16c98 , \49840 , \49841_nG16c99 , \49842_nG16c9a , \49843 , \49844_nG18dbe ,
         \49845 , \49846 , \49847_nG16c9b , \49848_nG16c9c , \49849 , \49850_nG16c9d , \49851_nG16c9e , \49852 , \49853_nG18dc0 , \49854 ,
         \49855 , \49856_nG16c9f , \49857_nG16ca0 , \49858 , \49859_nG16ca1 , \49860_nG16ca2 , \49861 , \49862_nG18dc2 , \49863 , \49864 ,
         \49865_nG16ca3 , \49866_nG16ca4 , \49867 , \49868_nG16ca5 , \49869_nG16ca6 , \49870 , \49871_nG18dc4 , \49872 , \49873 , \49874_nG16ca7 ,
         \49875_nG16ca8 , \49876 , \49877_nG16ca9 , \49878_nG16caa , \49879 , \49880_nG18dc8 , \49881 , \49882 , \49883_nG16cab , \49884_nG16cac ,
         \49885 , \49886_nG16cad , \49887_nG16cae , \49888 , \49889_nG18dca , \49890 , \49891 , \49892_nG16caf , \49893_nG16cb0 , \49894 ,
         \49895_nG16cb1 , \49896_nG16cb2 , \49897 , \49898_nG18dcc , \49899 , \49900 , \49901_nG16cb3 , \49902_nG16cb4 , \49903 , \49904_nG16cb5 ,
         \49905_nG16cb6 , \49906 , \49907_nG18dce , \49908 , \49909 , \49910_nG16cb7 , \49911_nG16cb8 , \49912 , \49913_nG16cb9 , \49914_nG16cba ,
         \49915 , \49916_nG18dd0 , \49917 , \49918 , \49919_nG16cbb , \49920_nG16cbc , \49921 , \49922_nG16cbd , \49923_nG16cbe , \49924 ,
         \49925_nG18dd2 , \49926 , \49927 , \49928_nG16cbf , \49929_nG16cc0 , \49930 , \49931_nG16cc1 , \49932_nG16cc2 , \49933 , \49934_nG18dd4 ,
         \49935 , \49936 , \49937_nG16cc3 , \49938_nG16cc4 , \49939 , \49940_nG16cc5 , \49941_nG16cc6 , \49942 , \49943_nG18dd6 , \49944 ,
         \49945 , \49946_nG16cc7 , \49947_nG16cc8 , \49948 , \49949_nG16cc9 , \49950_nG16cca , \49951 , \49952_nG18dd8 , \49953 , \49954 ,
         \49955_nG16ccb , \49956_nG16ccc , \49957 , \49958_nG16ccd , \49959_nG16cce , \49960 , \49961_nG18dda , \49962 , \49963 , \49964_nG16ccf ,
         \49965_nG16cd0 , \49966 , \49967_nG16cd1 , \49968_nG16cd2 , \49969 , \49970_nG18dde , \49971 , \49972 , \49973_nG16cd3 , \49974_nG16cd4 ,
         \49975 , \49976_nG16cd5 , \49977_nG16cd6 , \49978 , \49979_nG18de0 , \49980 , \49981 , \49982_nG16cd7 , \49983_nG16cd8 , \49984 ,
         \49985_nG16cd9 , \49986_nG16cda , \49987 , \49988_nG18de2 , \49989 , \49990 , \49991_nG16cdb , \49992_nG16cdc , \49993 , \49994_nG16cdd ,
         \49995_nG16cde , \49996 , \49997_nG18de4 , \49998 , \49999 , \50000_nG16cdf , \50001_nG16ce0 , \50002 , \50003_nG16ce1 , \50004_nG16ce2 ,
         \50005 , \50006_nG18de6 , \50007 , \50008 , \50009_nG16ce3 , \50010_nG16ce4 , \50011 , \50012_nG16ce5 , \50013_nG16ce6 , \50014 ,
         \50015_nG18de8 , \50016 , \50017 , \50018_nG16ce7 , \50019_nG16ce8 , \50020 , \50021_nG16ce9 , \50022_nG16cea , \50023 , \50024_nG18dea ,
         \50025 , \50026 , \50027_nG16ceb , \50028_nG16cec , \50029 , \50030_nG16ced , \50031_nG16cee , \50032 , \50033_nG18dec , \50034 ,
         \50035 , \50036_nG16cef , \50037_nG16cf0 , \50038 , \50039_nG16cf1 , \50040_nG16cf2 , \50041 , \50042_nG18dee , \50043 , \50044 ,
         \50045_nG16cf3 , \50046_nG16cf4 , \50047 , \50048_nG16cf5 , \50049_nG16cf6 , \50050 , \50051_nG18df0 , \50052 , \50053 , \50054_nG16cf7 ,
         \50055_nG16cf8 , \50056 , \50057_nG16cf9 , \50058_nG16cfa , \50059 , \50060_nG18df4 , \50061 , \50062 , \50063_nG16cfb , \50064_nG16cfc ,
         \50065 , \50066_nG16cfd , \50067_nG16cfe , \50068 , \50069_nG18df6 , \50070 , \50071 , \50072_nG16cff , \50073_nG16d00 , \50074 ,
         \50075_nG16d01 , \50076_nG16d02 , \50077 , \50078_nG18df8 , \50079 , \50080 , \50081_nG16d03 , \50082_nG16d04 , \50083 , \50084_nG16d05 ,
         \50085_nG16d06 , \50086 , \50087_nG18dfa , \50088 , \50089 , \50090_nG16d07 , \50091_nG16d08 , \50092 , \50093_nG16d09 , \50094_nG16d0a ,
         \50095 , \50096_nG18dfc , \50097 , \50098 , \50099 , \50100_nG16b09 , \50101_nG16b0a , \50102 , \50103 , \50104_nG16b0c ,
         \50105_nG16b0d , \50106 , \50107_nG18d04 , \50108 , \50109_nG16b0e , \50110_nG16b0f , \50111_nG16b10 , \50112_nG16b11 , \50113 , \50114_nG18d1a ,
         \50115 , \50116_nG16b12 , \50117_nG16b13 , \50118_nG16b14 , \50119_nG16b15 , \50120 , \50121_nG18d30 , \50122 , \50123_nG16b16 , \50124_nG16b17 ,
         \50125_nG16b18 , \50126_nG16b19 , \50127 , \50128_nG18d46 , \50129 , \50130_nG16b1a , \50131_nG16b1b , \50132_nG16b1c , \50133_nG16b1d , \50134 ,
         \50135_nG18d5c , \50136 , \50137_nG16b1e , \50138_nG16b1f , \50139_nG16b20 , \50140_nG16b21 , \50141 , \50142_nG18d72 , \50143 , \50144_nG16b22 ,
         \50145_nG16b23 , \50146_nG16b24 , \50147_nG16b25 , \50148 , \50149_nG18d7e , \50150 , \50151_nG16b26 , \50152_nG16b27 , \50153_nG16b28 , \50154_nG16b29 ,
         \50155 , \50156_nG18d80 , \50157 , \50158_nG16b2a , \50159_nG16b2b , \50160_nG16b2c , \50161_nG16b2d , \50162 , \50163_nG18d82 , \50164 ,
         \50165_nG16b2e , \50166_nG16b2f , \50167_nG16b30 , \50168_nG16b31 , \50169 , \50170_nG18d06 , \50171 , \50172_nG16b32 , \50173_nG16b33 , \50174_nG16b34 ,
         \50175_nG16b35 , \50176 , \50177_nG18d08 , \50178 , \50179_nG16b36 , \50180_nG16b37 , \50181_nG16b38 , \50182_nG16b39 , \50183 , \50184_nG18d0a ,
         \50185 , \50186_nG16b3a , \50187_nG16b3b , \50188_nG16b3c , \50189_nG16b3d , \50190 , \50191_nG18d0c , \50192 , \50193_nG16b3e , \50194_nG16b3f ,
         \50195_nG16b40 , \50196_nG16b41 , \50197 , \50198_nG18d0e , \50199 , \50200_nG16b42 , \50201_nG16b43 , \50202_nG16b44 , \50203_nG16b45 , \50204 ,
         \50205_nG18d10 , \50206 , \50207_nG16b46 , \50208_nG16b47 , \50209_nG16b48 , \50210_nG16b49 , \50211 , \50212_nG18d12 , \50213 , \50214_nG16b4a ,
         \50215_nG16b4b , \50216_nG16b4c , \50217_nG16b4d , \50218 , \50219_nG18d14 , \50220 , \50221_nG16b4e , \50222_nG16b4f , \50223_nG16b50 , \50224_nG16b51 ,
         \50225 , \50226_nG18d16 , \50227 , \50228_nG16b52 , \50229_nG16b53 , \50230_nG16b54 , \50231_nG16b55 , \50232 , \50233_nG18d18 , \50234 ,
         \50235_nG16b56 , \50236_nG16b57 , \50237_nG16b58 , \50238_nG16b59 , \50239 , \50240_nG18d1c , \50241 , \50242_nG16b5a , \50243_nG16b5b , \50244_nG16b5c ,
         \50245_nG16b5d , \50246 , \50247_nG18d1e , \50248 , \50249_nG16b5e , \50250_nG16b5f , \50251_nG16b60 , \50252_nG16b61 , \50253 , \50254_nG18d20 ,
         \50255 , \50256_nG16b62 , \50257_nG16b63 , \50258_nG16b64 , \50259_nG16b65 , \50260 , \50261_nG18d22 , \50262 , \50263_nG16b66 , \50264_nG16b67 ,
         \50265_nG16b68 , \50266_nG16b69 , \50267 , \50268_nG18d24 , \50269 , \50270_nG16b6a , \50271_nG16b6b , \50272_nG16b6c , \50273_nG16b6d , \50274 ,
         \50275_nG18d26 , \50276 , \50277_nG16b6e , \50278_nG16b6f , \50279_nG16b70 , \50280_nG16b71 , \50281 , \50282_nG18d28 , \50283 , \50284_nG16b72 ,
         \50285_nG16b73 , \50286_nG16b74 , \50287_nG16b75 , \50288 , \50289_nG18d2a , \50290 , \50291_nG16b76 , \50292_nG16b77 , \50293_nG16b78 , \50294_nG16b79 ,
         \50295 , \50296_nG18d2c , \50297 , \50298_nG16b7a , \50299_nG16b7b , \50300_nG16b7c , \50301_nG16b7d , \50302 , \50303_nG18d2e , \50304 ,
         \50305_nG16b7e , \50306_nG16b7f , \50307_nG16b80 , \50308_nG16b81 , \50309 , \50310_nG18d32 , \50311 , \50312_nG16b82 , \50313_nG16b83 , \50314_nG16b84 ,
         \50315_nG16b85 , \50316 , \50317_nG18d34 , \50318 , \50319_nG16b86 , \50320_nG16b87 , \50321_nG16b88 , \50322_nG16b89 , \50323 , \50324_nG18d36 ,
         \50325 , \50326_nG16b8a , \50327_nG16b8b , \50328_nG16b8c , \50329_nG16b8d , \50330 , \50331_nG18d38 , \50332 , \50333_nG16b8e , \50334_nG16b8f ,
         \50335_nG16b90 , \50336_nG16b91 , \50337 , \50338_nG18d3a , \50339 , \50340_nG16b92 , \50341_nG16b93 , \50342_nG16b94 , \50343_nG16b95 , \50344 ,
         \50345_nG18d3c , \50346 , \50347_nG16b96 , \50348_nG16b97 , \50349_nG16b98 , \50350_nG16b99 , \50351 , \50352_nG18d3e , \50353 , \50354_nG16b9a ,
         \50355_nG16b9b , \50356_nG16b9c , \50357_nG16b9d , \50358 , \50359_nG18d40 , \50360 , \50361_nG16b9e , \50362_nG16b9f , \50363_nG16ba0 , \50364_nG16ba1 ,
         \50365 , \50366_nG18d42 , \50367 , \50368_nG16ba2 , \50369_nG16ba3 , \50370_nG16ba4 , \50371_nG16ba5 , \50372 , \50373_nG18d44 , \50374 ,
         \50375_nG16ba6 , \50376_nG16ba7 , \50377_nG16ba8 , \50378_nG16ba9 , \50379 , \50380_nG18d48 , \50381 , \50382_nG16baa , \50383_nG16bab , \50384_nG16bac ,
         \50385_nG16bad , \50386 , \50387_nG18d4a , \50388 , \50389_nG16bae , \50390_nG16baf , \50391_nG16bb0 , \50392_nG16bb1 , \50393 , \50394_nG18d4c ,
         \50395 , \50396_nG16bb2 , \50397_nG16bb3 , \50398_nG16bb4 , \50399_nG16bb5 , \50400 , \50401_nG18d4e , \50402 , \50403_nG16bb6 , \50404_nG16bb7 ,
         \50405_nG16bb8 , \50406_nG16bb9 , \50407 , \50408_nG18d50 , \50409 , \50410_nG16bba , \50411_nG16bbb , \50412_nG16bbc , \50413_nG16bbd , \50414 ,
         \50415_nG18d52 , \50416 , \50417_nG16bbe , \50418_nG16bbf , \50419_nG16bc0 , \50420_nG16bc1 , \50421 , \50422_nG18d54 , \50423 , \50424_nG16bc2 ,
         \50425_nG16bc3 , \50426_nG16bc4 , \50427_nG16bc5 , \50428 , \50429_nG18d56 , \50430 , \50431_nG16bc6 , \50432_nG16bc7 , \50433_nG16bc8 , \50434_nG16bc9 ,
         \50435 , \50436_nG18d58 , \50437 , \50438_nG16bca , \50439_nG16bcb , \50440_nG16bcc , \50441_nG16bcd , \50442 , \50443_nG18d5a , \50444 ,
         \50445_nG16bce , \50446_nG16bcf , \50447_nG16bd0 , \50448_nG16bd1 , \50449 , \50450_nG18d5e , \50451 , \50452_nG16bd2 , \50453_nG16bd3 , \50454_nG16bd4 ,
         \50455_nG16bd5 , \50456 , \50457_nG18d60 , \50458 , \50459_nG16bd6 , \50460_nG16bd7 , \50461_nG16bd8 , \50462_nG16bd9 , \50463 , \50464_nG18d62 ,
         \50465 , \50466_nG16bda , \50467_nG16bdb , \50468_nG16bdc , \50469_nG16bdd , \50470 , \50471_nG18d64 , \50472 , \50473_nG16bde , \50474_nG16bdf ,
         \50475_nG16be0 , \50476_nG16be1 , \50477 , \50478_nG18d66 , \50479 , \50480_nG16be2 , \50481_nG16be3 , \50482_nG16be4 , \50483_nG16be5 , \50484 ,
         \50485_nG18d68 , \50486 , \50487_nG16be6 , \50488_nG16be7 , \50489_nG16be8 , \50490_nG16be9 , \50491 , \50492_nG18d6a , \50493 , \50494_nG16bea ,
         \50495_nG16beb , \50496_nG16bec , \50497_nG16bed , \50498 , \50499_nG18d6c , \50500 , \50501_nG16bee , \50502_nG16bef , \50503_nG16bf0 , \50504_nG16bf1 ,
         \50505 , \50506_nG18d6e , \50507 , \50508_nG16bf2 , \50509_nG16bf3 , \50510_nG16bf4 , \50511_nG16bf5 , \50512 , \50513_nG18d70 , \50514 ,
         \50515_nG16bf6 , \50516_nG16bf7 , \50517_nG16bf8 , \50518_nG16bf9 , \50519 , \50520_nG18d74 , \50521 , \50522_nG16bfa , \50523_nG16bfb , \50524_nG16bfc ,
         \50525_nG16bfd , \50526 , \50527_nG18d76 , \50528 , \50529_nG16bfe , \50530_nG16bff , \50531_nG16c00 , \50532_nG16c01 , \50533 , \50534_nG18d78 ,
         \50535 , \50536_nG16c02 , \50537_nG16c03 , \50538_nG16c04 , \50539_nG16c05 , \50540 , \50541_nG18d7a , \50542 , \50543_nG16c06 , \50544_nG16c07 ,
         \50545_nG16c08 , \50546_nG16c09 , \50547 , \50548_nG18d7c , \50549 , \50550 , \50551_nG16a07 , \50552_nG16a08 , \50553 , \50554_nG16a0b ,
         \50555_nG16a0c , \50556 , \50557_nG18c84 , \50558 , \50559_nG16a0d , \50560_nG16a0e , \50561_nG16a0f , \50562_nG16a10 , \50563 , \50564_nG18c9a ,
         \50565 , \50566_nG16a11 , \50567_nG16a12 , \50568_nG16a13 , \50569_nG16a14 , \50570 , \50571_nG18cb0 , \50572 , \50573_nG16a15 , \50574_nG16a16 ,
         \50575_nG16a17 , \50576_nG16a18 , \50577 , \50578_nG18cc6 , \50579 , \50580_nG16a19 , \50581_nG16a1a , \50582_nG16a1b , \50583_nG16a1c , \50584 ,
         \50585_nG18cdc , \50586 , \50587_nG16a1d , \50588_nG16a1e , \50589_nG16a1f , \50590_nG16a20 , \50591 , \50592_nG18cf2 , \50593 , \50594_nG16a21 ,
         \50595_nG16a22 , \50596_nG16a23 , \50597_nG16a24 , \50598 , \50599_nG18cfe , \50600 , \50601_nG16a25 , \50602_nG16a26 , \50603_nG16a27 , \50604_nG16a28 ,
         \50605 , \50606_nG18d00 , \50607 , \50608_nG16a29 , \50609_nG16a2a , \50610_nG16a2b , \50611_nG16a2c , \50612 , \50613_nG18d02 , \50614 ,
         \50615_nG16a2d , \50616_nG16a2e , \50617_nG16a2f , \50618_nG16a30 , \50619 , \50620_nG18c86 , \50621 , \50622_nG16a31 , \50623_nG16a32 , \50624_nG16a33 ,
         \50625_nG16a34 , \50626 , \50627_nG18c88 , \50628 , \50629_nG16a35 , \50630_nG16a36 , \50631_nG16a37 , \50632_nG16a38 , \50633 , \50634_nG18c8a ,
         \50635 , \50636_nG16a39 , \50637_nG16a3a , \50638_nG16a3b , \50639_nG16a3c , \50640 , \50641_nG18c8c , \50642 , \50643_nG16a3d , \50644_nG16a3e ,
         \50645_nG16a3f , \50646_nG16a40 , \50647 , \50648_nG18c8e , \50649 , \50650_nG16a41 , \50651_nG16a42 , \50652_nG16a43 , \50653_nG16a44 , \50654 ,
         \50655_nG18c90 , \50656 , \50657_nG16a45 , \50658_nG16a46 , \50659_nG16a47 , \50660_nG16a48 , \50661 , \50662_nG18c92 , \50663 , \50664_nG16a49 ,
         \50665_nG16a4a , \50666_nG16a4b , \50667_nG16a4c , \50668 , \50669_nG18c94 , \50670 , \50671_nG16a4d , \50672_nG16a4e , \50673_nG16a4f , \50674_nG16a50 ,
         \50675 , \50676_nG18c96 , \50677 , \50678_nG16a51 , \50679_nG16a52 , \50680_nG16a53 , \50681_nG16a54 , \50682 , \50683_nG18c98 , \50684 ,
         \50685_nG16a55 , \50686_nG16a56 , \50687_nG16a57 , \50688_nG16a58 , \50689 , \50690_nG18c9c , \50691 , \50692_nG16a59 , \50693_nG16a5a , \50694_nG16a5b ,
         \50695_nG16a5c , \50696 , \50697_nG18c9e , \50698 , \50699_nG16a5d , \50700_nG16a5e , \50701_nG16a5f , \50702_nG16a60 , \50703 , \50704_nG18ca0 ,
         \50705 , \50706_nG16a61 , \50707_nG16a62 , \50708_nG16a63 , \50709_nG16a64 , \50710 , \50711_nG18ca2 , \50712 , \50713_nG16a65 , \50714_nG16a66 ,
         \50715_nG16a67 , \50716_nG16a68 , \50717 , \50718_nG18ca4 , \50719 , \50720_nG16a69 , \50721_nG16a6a , \50722_nG16a6b , \50723_nG16a6c , \50724 ,
         \50725_nG18ca6 , \50726 , \50727_nG16a6d , \50728_nG16a6e , \50729_nG16a6f , \50730_nG16a70 , \50731 , \50732_nG18ca8 , \50733 , \50734_nG16a71 ,
         \50735_nG16a72 , \50736_nG16a73 , \50737_nG16a74 , \50738 , \50739_nG18caa , \50740 , \50741_nG16a75 , \50742_nG16a76 , \50743_nG16a77 , \50744_nG16a78 ,
         \50745 , \50746_nG18cac , \50747 , \50748_nG16a79 , \50749_nG16a7a , \50750_nG16a7b , \50751_nG16a7c , \50752 , \50753_nG18cae , \50754 ,
         \50755_nG16a7d , \50756_nG16a7e , \50757_nG16a7f , \50758_nG16a80 , \50759 , \50760_nG18cb2 , \50761 , \50762_nG16a81 , \50763_nG16a82 , \50764_nG16a83 ,
         \50765_nG16a84 , \50766 , \50767_nG18cb4 , \50768 , \50769_nG16a85 , \50770_nG16a86 , \50771_nG16a87 , \50772_nG16a88 , \50773 , \50774_nG18cb6 ,
         \50775 , \50776_nG16a89 , \50777_nG16a8a , \50778_nG16a8b , \50779_nG16a8c , \50780 , \50781_nG18cb8 , \50782 , \50783_nG16a8d , \50784_nG16a8e ,
         \50785_nG16a8f , \50786_nG16a90 , \50787 , \50788_nG18cba , \50789 , \50790_nG16a91 , \50791_nG16a92 , \50792_nG16a93 , \50793_nG16a94 , \50794 ,
         \50795_nG18cbc , \50796 , \50797_nG16a95 , \50798_nG16a96 , \50799_nG16a97 , \50800_nG16a98 , \50801 , \50802_nG18cbe , \50803 , \50804_nG16a99 ,
         \50805_nG16a9a , \50806_nG16a9b , \50807_nG16a9c , \50808 , \50809_nG18cc0 , \50810 , \50811_nG16a9d , \50812_nG16a9e , \50813_nG16a9f , \50814_nG16aa0 ,
         \50815 , \50816_nG18cc2 , \50817 , \50818_nG16aa1 , \50819_nG16aa2 , \50820_nG16aa3 , \50821_nG16aa4 , \50822 , \50823_nG18cc4 , \50824 ,
         \50825_nG16aa5 , \50826_nG16aa6 , \50827_nG16aa7 , \50828_nG16aa8 , \50829 , \50830_nG18cc8 , \50831 , \50832_nG16aa9 , \50833_nG16aaa , \50834_nG16aab ,
         \50835_nG16aac , \50836 , \50837_nG18cca , \50838 , \50839_nG16aad , \50840_nG16aae , \50841_nG16aaf , \50842_nG16ab0 , \50843 , \50844_nG18ccc ,
         \50845 , \50846_nG16ab1 , \50847_nG16ab2 , \50848_nG16ab3 , \50849_nG16ab4 , \50850 , \50851_nG18cce , \50852 , \50853_nG16ab5 , \50854_nG16ab6 ,
         \50855_nG16ab7 , \50856_nG16ab8 , \50857 , \50858_nG18cd0 , \50859 , \50860_nG16ab9 , \50861_nG16aba , \50862_nG16abb , \50863_nG16abc , \50864 ,
         \50865_nG18cd2 , \50866 , \50867_nG16abd , \50868_nG16abe , \50869_nG16abf , \50870_nG16ac0 , \50871 , \50872_nG18cd4 , \50873 , \50874_nG16ac1 ,
         \50875_nG16ac2 , \50876_nG16ac3 , \50877_nG16ac4 , \50878 , \50879_nG18cd6 , \50880 , \50881_nG16ac5 , \50882_nG16ac6 , \50883_nG16ac7 , \50884_nG16ac8 ,
         \50885 , \50886_nG18cd8 , \50887 , \50888_nG16ac9 , \50889_nG16aca , \50890_nG16acb , \50891_nG16acc , \50892 , \50893_nG18cda , \50894 ,
         \50895_nG16acd , \50896_nG16ace , \50897_nG16acf , \50898_nG16ad0 , \50899 , \50900_nG18cde , \50901 , \50902_nG16ad1 , \50903_nG16ad2 , \50904_nG16ad3 ,
         \50905_nG16ad4 , \50906 , \50907_nG18ce0 , \50908 , \50909_nG16ad5 , \50910_nG16ad6 , \50911_nG16ad7 , \50912_nG16ad8 , \50913 , \50914_nG18ce2 ,
         \50915 , \50916_nG16ad9 , \50917_nG16ada , \50918_nG16adb , \50919_nG16adc , \50920 , \50921_nG18ce4 , \50922 , \50923_nG16add , \50924_nG16ade ,
         \50925_nG16adf , \50926_nG16ae0 , \50927 , \50928_nG18ce6 , \50929 , \50930_nG16ae1 , \50931_nG16ae2 , \50932_nG16ae3 , \50933_nG16ae4 , \50934 ,
         \50935_nG18ce8 , \50936 , \50937_nG16ae5 , \50938_nG16ae6 , \50939_nG16ae7 , \50940_nG16ae8 , \50941 , \50942_nG18cea , \50943 , \50944_nG16ae9 ,
         \50945_nG16aea , \50946_nG16aeb , \50947_nG16aec , \50948 , \50949_nG18cec , \50950 , \50951_nG16aed , \50952_nG16aee , \50953_nG16aef , \50954_nG16af0 ,
         \50955 , \50956_nG18cee , \50957 , \50958_nG16af1 , \50959_nG16af2 , \50960_nG16af3 , \50961_nG16af4 , \50962 , \50963_nG18cf0 , \50964 ,
         \50965_nG16af5 , \50966_nG16af6 , \50967_nG16af7 , \50968_nG16af8 , \50969 , \50970_nG18cf4 , \50971 , \50972_nG16af9 , \50973_nG16afa , \50974_nG16afb ,
         \50975_nG16afc , \50976 , \50977_nG18cf6 , \50978 , \50979_nG16afd , \50980_nG16afe , \50981_nG16aff , \50982_nG16b00 , \50983 , \50984_nG18cf8 ,
         \50985 , \50986_nG16b01 , \50987_nG16b02 , \50988_nG16b03 , \50989_nG16b04 , \50990 , \50991_nG18cfa , \50992 , \50993_nG16b05 , \50994_nG16b06 ,
         \50995_nG16b07 , \50996_nG16b08 , \50997 , \50998_nG18cfc , \50999 , \51000 , \51001_nG16885 , \51002_nG16886 , \51003 , \51004_nG1688b ,
         \51005_nG1688c , \51006 , \51007_nG18c04 , \51008 , \51009_nG1688e , \51010_nG1688f , \51011_nG16891 , \51012_nG16892 , \51013 , \51014_nG18c1a ,
         \51015 , \51016_nG16894 , \51017_nG16895 , \51018_nG16897 , \51019_nG16898 , \51020 , \51021_nG18c30 , \51022 , \51023_nG1689a , \51024_nG1689b ,
         \51025_nG1689d , \51026_nG1689e , \51027 , \51028_nG18c46 , \51029 , \51030_nG168a0 , \51031_nG168a1 , \51032_nG168a3 , \51033_nG168a4 , \51034 ,
         \51035_nG18c5c , \51036 , \51037_nG168a6 , \51038_nG168a7 , \51039_nG168a9 , \51040_nG168aa , \51041 , \51042_nG18c72 , \51043 , \51044_nG168ac ,
         \51045_nG168ad , \51046_nG168af , \51047_nG168b0 , \51048 , \51049_nG18c7e , \51050 , \51051_nG168b2 , \51052_nG168b3 , \51053_nG168b5 , \51054_nG168b6 ,
         \51055 , \51056_nG18c80 , \51057 , \51058_nG168b8 , \51059_nG168b9 , \51060_nG168bb , \51061_nG168bc , \51062 , \51063_nG18c82 , \51064 ,
         \51065_nG168be , \51066_nG168bf , \51067_nG168c1 , \51068_nG168c2 , \51069 , \51070_nG18c06 , \51071 , \51072_nG168c4 , \51073_nG168c5 , \51074_nG168c7 ,
         \51075_nG168c8 , \51076 , \51077_nG18c08 , \51078 , \51079_nG168ca , \51080_nG168cb , \51081_nG168cd , \51082_nG168ce , \51083 , \51084_nG18c0a ,
         \51085 , \51086_nG168d0 , \51087_nG168d1 , \51088_nG168d3 , \51089_nG168d4 , \51090 , \51091_nG18c0c , \51092 , \51093_nG168d6 , \51094_nG168d7 ,
         \51095_nG168d9 , \51096_nG168da , \51097 , \51098_nG18c0e , \51099 , \51100_nG168dc , \51101_nG168dd , \51102_nG168df , \51103_nG168e0 , \51104 ,
         \51105_nG18c10 , \51106 , \51107_nG168e2 , \51108_nG168e3 , \51109_nG168e5 , \51110_nG168e6 , \51111 , \51112_nG18c12 , \51113 , \51114_nG168e8 ,
         \51115_nG168e9 , \51116_nG168eb , \51117_nG168ec , \51118 , \51119_nG18c14 , \51120 , \51121_nG168ee , \51122_nG168ef , \51123_nG168f1 , \51124_nG168f2 ,
         \51125 , \51126_nG18c16 , \51127 , \51128_nG168f4 , \51129_nG168f5 , \51130_nG168f7 , \51131_nG168f8 , \51132 , \51133_nG18c18 , \51134 ,
         \51135_nG168fa , \51136_nG168fb , \51137_nG168fd , \51138_nG168fe , \51139 , \51140_nG18c1c , \51141 , \51142_nG16900 , \51143_nG16901 , \51144_nG16903 ,
         \51145_nG16904 , \51146 , \51147_nG18c1e , \51148 , \51149_nG16906 , \51150_nG16907 , \51151_nG16909 , \51152_nG1690a , \51153 , \51154_nG18c20 ,
         \51155 , \51156_nG1690c , \51157_nG1690d , \51158_nG1690f , \51159_nG16910 , \51160 , \51161_nG18c22 , \51162 , \51163_nG16912 , \51164_nG16913 ,
         \51165_nG16915 , \51166_nG16916 , \51167 , \51168_nG18c24 , \51169 , \51170_nG16918 , \51171_nG16919 , \51172_nG1691b , \51173_nG1691c , \51174 ,
         \51175_nG18c26 , \51176 , \51177_nG1691e , \51178_nG1691f , \51179_nG16921 , \51180_nG16922 , \51181 , \51182_nG18c28 , \51183 , \51184_nG16924 ,
         \51185_nG16925 , \51186_nG16927 , \51187_nG16928 , \51188 , \51189_nG18c2a , \51190 , \51191_nG1692a , \51192_nG1692b , \51193_nG1692d , \51194_nG1692e ,
         \51195 , \51196_nG18c2c , \51197 , \51198_nG16930 , \51199_nG16931 , \51200_nG16933 , \51201_nG16934 , \51202 , \51203_nG18c2e , \51204 ,
         \51205_nG16936 , \51206_nG16937 , \51207_nG16939 , \51208_nG1693a , \51209 , \51210_nG18c32 , \51211 , \51212_nG1693c , \51213_nG1693d , \51214_nG1693f ,
         \51215_nG16940 , \51216 , \51217_nG18c34 , \51218 , \51219_nG16942 , \51220_nG16943 , \51221_nG16945 , \51222_nG16946 , \51223 , \51224_nG18c36 ,
         \51225 , \51226_nG16948 , \51227_nG16949 , \51228_nG1694b , \51229_nG1694c , \51230 , \51231_nG18c38 , \51232 , \51233_nG1694e , \51234_nG1694f ,
         \51235_nG16951 , \51236_nG16952 , \51237 , \51238_nG18c3a , \51239 , \51240_nG16954 , \51241_nG16955 , \51242_nG16957 , \51243_nG16958 , \51244 ,
         \51245_nG18c3c , \51246 , \51247_nG1695a , \51248_nG1695b , \51249_nG1695d , \51250_nG1695e , \51251 , \51252_nG18c3e , \51253 , \51254_nG16960 ,
         \51255_nG16961 , \51256_nG16963 , \51257_nG16964 , \51258 , \51259_nG18c40 , \51260 , \51261_nG16966 , \51262_nG16967 , \51263_nG16969 , \51264_nG1696a ,
         \51265 , \51266_nG18c42 , \51267 , \51268_nG1696c , \51269_nG1696d , \51270_nG1696f , \51271_nG16970 , \51272 , \51273_nG18c44 , \51274 ,
         \51275_nG16972 , \51276_nG16973 , \51277_nG16975 , \51278_nG16976 , \51279 , \51280_nG18c48 , \51281 , \51282_nG16978 , \51283_nG16979 , \51284_nG1697b ,
         \51285_nG1697c , \51286 , \51287_nG18c4a , \51288 , \51289_nG1697e , \51290_nG1697f , \51291_nG16981 , \51292_nG16982 , \51293 , \51294_nG18c4c ,
         \51295 , \51296_nG16984 , \51297_nG16985 , \51298_nG16987 , \51299_nG16988 , \51300 , \51301_nG18c4e , \51302 , \51303_nG1698a , \51304_nG1698b ,
         \51305_nG1698d , \51306_nG1698e , \51307 , \51308_nG18c50 , \51309 , \51310_nG16990 , \51311_nG16991 , \51312_nG16993 , \51313_nG16994 , \51314 ,
         \51315_nG18c52 , \51316 , \51317_nG16996 , \51318_nG16997 , \51319_nG16999 , \51320_nG1699a , \51321 , \51322_nG18c54 , \51323 , \51324_nG1699c ,
         \51325_nG1699d , \51326_nG1699f , \51327_nG169a0 , \51328 , \51329_nG18c56 , \51330 , \51331_nG169a2 , \51332_nG169a3 , \51333_nG169a5 , \51334_nG169a6 ,
         \51335 , \51336_nG18c58 , \51337 , \51338_nG169a8 , \51339_nG169a9 , \51340_nG169ab , \51341_nG169ac , \51342 , \51343_nG18c5a , \51344 ,
         \51345_nG169ae , \51346_nG169af , \51347_nG169b1 , \51348_nG169b2 , \51349 , \51350_nG18c5e , \51351 , \51352_nG169b4 , \51353_nG169b5 , \51354_nG169b7 ,
         \51355_nG169b8 , \51356 , \51357_nG18c60 , \51358 , \51359_nG169ba , \51360_nG169bb , \51361_nG169bd , \51362_nG169be , \51363 , \51364_nG18c62 ,
         \51365 , \51366_nG169c0 , \51367_nG169c1 , \51368_nG169c3 , \51369_nG169c4 , \51370 , \51371_nG18c64 , \51372 , \51373_nG169c6 , \51374_nG169c7 ,
         \51375_nG169c9 , \51376_nG169ca , \51377 , \51378_nG18c66 , \51379 , \51380_nG169cc , \51381_nG169cd , \51382_nG169cf , \51383_nG169d0 , \51384 ,
         \51385_nG18c68 , \51386 , \51387_nG169d2 , \51388_nG169d3 , \51389_nG169d5 , \51390_nG169d6 , \51391 , \51392_nG18c6a , \51393 , \51394_nG169d8 ,
         \51395_nG169d9 , \51396_nG169db , \51397_nG169dc , \51398 , \51399_nG18c6c , \51400 , \51401_nG169de , \51402_nG169df , \51403_nG169e1 , \51404_nG169e2 ,
         \51405 , \51406_nG18c6e , \51407 , \51408_nG169e4 , \51409_nG169e5 , \51410_nG169e7 , \51411_nG169e8 , \51412 , \51413_nG18c70 , \51414 ,
         \51415_nG169ea , \51416_nG169eb , \51417_nG169ed , \51418_nG169ee , \51419 , \51420_nG18c74 , \51421 , \51422_nG169f0 , \51423_nG169f1 , \51424_nG169f3 ,
         \51425_nG169f4 , \51426 , \51427_nG18c76 , \51428 , \51429_nG169f6 , \51430_nG169f7 , \51431_nG169f9 , \51432_nG169fa , \51433 , \51434_nG18c78 ,
         \51435 , \51436_nG169fc , \51437_nG169fd , \51438_nG169ff , \51439_nG16a00 , \51440 , \51441_nG18c7a , \51442 , \51443_nG16a02 , \51444_nG16a03 ,
         \51445_nG16a05 , \51446_nG16a06 , \51447 , \51448_nG18c7c , \51449 , \51450 , \51451_nG16857 , \51452 , \51453 , \51454_nG16858 ,
         \51455 , \51456_nG18bec , \51457 , \51458 , \51459_nG16859 , \51460_nG1685a , \51461 , \51462_nG18bee , \51463 , \51464 ,
         \51465_nG1685b , \51466_nG1685c , \51467 , \51468_nG18bf0 , \51469 , \51470 , \51471_nG1685d , \51472_nG1685e , \51473 , \51474_nG18bf2 ,
         \51475 , \51476 , \51477_nG1685f , \51478_nG16860 , \51479 , \51480_nG18bf4 , \51481 , \51482 , \51483_nG16861 , \51484_nG16862 ,
         \51485 , \51486_nG18bf6 , \51487 , \51488 , \51489_nG16863 , \51490_nG16864 , \51491 , \51492_nG18bf8 , \51493 , \51494 ,
         \51495_nG16865 , \51496_nG16866 , \51497 , \51498_nG18bfa , \51499 , \51500_nG16846 , \51501_nG16847 , \51502 , \51503_nG18bdc , \51504 ,
         \51505_nG16848 , \51506_nG16849 , \51507 , \51508_nG18bde , \51509 , \51510_nG1684a , \51511_nG1684b , \51512 , \51513_nG18be0 , \51514 ,
         \51515_nG1684c , \51516_nG1684d , \51517 , \51518_nG18be2 , \51519 , \51520_nG1684e , \51521_nG1684f , \51522 , \51523_nG18be4 , \51524 ,
         \51525_nG16850 , \51526_nG16851 , \51527 , \51528_nG18be6 , \51529 , \51530_nG16852 , \51531_nG16853 , \51532 , \51533_nG18be8 , \51534 ,
         \51535_nG16854 , \51536_nG16855 , \51537 , \51538_nG18bea , \51539 , \51540_nG16835 , \51541_nG16836 , \51542 , \51543_nG18bcc , \51544 ,
         \51545_nG16837 , \51546_nG16838 , \51547 , \51548_nG18bce , \51549 , \51550_nG16839 , \51551_nG1683a , \51552 , \51553_nG18bd0 , \51554 ,
         \51555_nG1683b , \51556_nG1683c , \51557 , \51558_nG18bd2 , \51559 , \51560_nG1683d , \51561_nG1683e , \51562 , \51563_nG18bd4 , \51564 ,
         \51565_nG1683f , \51566_nG16840 , \51567 , \51568_nG18bd6 , \51569 , \51570_nG16841 , \51571_nG16842 , \51572 , \51573_nG18bd8 , \51574 ,
         \51575_nG16843 , \51576_nG16844 , \51577 , \51578_nG18bda , \51579 , \51580_nG16814 , \51581_nG1681d , \51582 , \51583_nG18e04 , \51584 ,
         \51585_nG1681f , \51586_nG16820 , \51587 , \51588_nG18e06 , \51589 , \51590_nG16822 , \51591_nG16823 , \51592 , \51593_nG18e08 , \51594 ,
         \51595_nG16825 , \51596_nG16826 , \51597 , \51598_nG18e0a , \51599 , \51600_nG16828 , \51601_nG16829 , \51602 , \51603_nG18e0c , \51604 ,
         \51605_nG1682b , \51606_nG1682c , \51607 , \51608_nG18e0e , \51609 , \51610_nG1682e , \51611_nG1682f , \51612 , \51613_nG18e10 , \51614 ,
         \51615_nG16831 , \51616_nG16832 , \51617 , \51618_nG18e12 , \51619 , \51620 , \51621 , \51622 , \51623_nG16709 , \51624 ,
         \51625_nG18e13 , \51626 , \51627 , \51628_nG16776 , \51629 , \51630_nG18bb0 , \51631 , \51632 , \51633_nG16778 , \51634 ,
         \51635_nG18bb2 , \51636 , \51637 , \51638_nG1677a , \51639 , \51640_nG18bb4 , \51641 , \51642 , \51643_nG1677c , \51644 ,
         \51645_nG18bb6 , \51646 , \51647 , \51648_nG1677e , \51649 , \51650_nG18bb8 , \51651 , \51652 , \51653_nG16780 , \51654 ,
         \51655_nG18bba , \51656 , \51657 , \51658_nG16782 , \51659 , \51660_nG18bbc , \51661 , \51662 , \51663_nG16774 , \51664 ,
         \51665_nG18bae , \51666 , \51667 , \51668_nG1676c , \51669 , \51670_nG18ba6 , \51671 , \51672 , \51673_nG1676e , \51674 ,
         \51675_nG18ba8 , \51676 , \51677 , \51678_nG16770 , \51679 , \51680_nG18baa , \51681 , \51682 , \51683_nG16772 , \51684 ,
         \51685_nG18bac , \51686 , \51687 , \51688 , \51689 , \51690 , \51691_nG165dc , \51692 , \51693 , \51694 ,
         \51695 , \51696_nG165dd , \51697 , \51698 , \51699 , \51700 , \51701 , \51702_nG165e3 , \51703 , \51704_nG165e7 ,
         \51705 , \51706 , \51707_nG165ea , \51708 , \51709 , \51710 , \51711 , \51712 , \51713_nG165f1 , \51714 ,
         \51715 , \51716_nG165f2 , \51717 , \51718 , \51719 , \51720 , \51721_nG165f6 , \51722_nG165f7 , \51723 , \51724 ,
         \51725 , \51726_nG165fb , \51727_nG165fc , \51728_nG165fd , \51729_nG165fe , \51730_nG165ff , \51731 , \51732 , \51733 , \51734 ,
         \51735 , \51736_nG16604 , \51737_nG16605 , \51738 , \51739 , \51740 , \51741 , \51742_nG1660a , \51743_nG1660b , \51744_nG1660c ,
         \51745_nG1660d , \51746_nG1660e , \51747 , \51748 , \51749 , \51750 , \51751 , \51752 , \51753 , \51754 ,
         \51755 , \51756 , \51757 , \51758 , \51759 , \51760_nG165d3 , \51761_nG165d4 , \51762 , \51763 , \51764 ,
         \51765 , \51766 , \51767 , \51768 , \51769 , \51770 , \51771 , \51772 , \51773 , \51774 ,
         \51775 , \51776_nG16691 , \51777 , \51778 , \51779 , \51780 , \51781 , \51782 , \51783 , \51784_nG16695 ,
         \51785 , \51786 , \51787_nG16696 , \51788 , \51789 , \51790_nG16697 , \51791 , \51792_nG16698 , \51793 , \51794 ,
         \51795 , \51796 , \51797_nG165cd , \51798_nG165ce , \51799 , \51800 , \51801 , \51802 , \51803_nG16682 , \51804 ,
         \51805 , \51806_nG16689 , \51807_nG1668a , \51808_nG1668b , \51809_nG1668c , \51810 , \51811 , \51812 , \51813 , \51814_nG165c6 ,
         \51815_nG165c9 , \51816 , \51817 , \51818 , \51819 , \51820_nG16672 , \51821 , \51822_nG16676 , \51823_nG16679 , \51824_nG1667c ,
         \51825_nG1667e , \51826 , \51827 , \51828 , \51829 , \51830 , \51831 , \51832 , \51833 , \51834 ,
         \51835 , \51836 , \51837 , \51838 , \51839_nG1670d , \51840 , \51841_nG18bca , \51842 , \51843 , \51844_nG18e17 ,
         \51845 , \51846 , \51847_nG18e18 , \51848 , \51849 , \51850_nG18e19 , \51851 , \51852 , \51853 , \51854 ,
         \51855 , \51856_nG164b7 , \51857 , \51858 , \51859 , \51860 , \51861 , \51862 , \51863_nG164b8 , \51864 ,
         \51865 , \51866 , \51867 , \51868_nG164ba , \51869 , \51870 , \51871 , \51872 , \51873 , \51874 ,
         \51875_nG164bb , \51876 , \51877_nG18b07 , \51878 , \51879 , \51880_nG164bc , \51881_nG164bd , \51882 , \51883_nG164be , \51884_nG164bf ,
         \51885 , \51886_nG18b1d , \51887 , \51888 , \51889_nG164c0 , \51890_nG164c1 , \51891 , \51892_nG164c2 , \51893_nG164c3 , \51894 ,
         \51895_nG18b33 , \51896 , \51897 , \51898_nG164c4 , \51899_nG164c5 , \51900 , \51901_nG164c6 , \51902_nG164c7 , \51903 , \51904_nG18b49 ,
         \51905 , \51906 , \51907_nG164c8 , \51908_nG164c9 , \51909 , \51910_nG164ca , \51911_nG164cb , \51912 , \51913_nG18b5f , \51914 ,
         \51915 , \51916_nG164cc , \51917_nG164cd , \51918 , \51919_nG164ce , \51920_nG164cf , \51921 , \51922_nG18b75 , \51923 , \51924 ,
         \51925_nG164d0 , \51926_nG164d1 , \51927 , \51928_nG164d2 , \51929_nG164d3 , \51930 , \51931_nG18b81 , \51932 , \51933 , \51934_nG164d4 ,
         \51935_nG164d5 , \51936 , \51937_nG164d6 , \51938_nG164d7 , \51939 , \51940_nG18b83 , \51941 , \51942 , \51943_nG164d8 , \51944_nG164d9 ,
         \51945 , \51946_nG164da , \51947_nG164db , \51948 , \51949_nG18b85 , \51950 , \51951 , \51952_nG164dc , \51953_nG164dd , \51954 ,
         \51955_nG164de , \51956_nG164df , \51957 , \51958_nG18b09 , \51959 , \51960 , \51961_nG164e0 , \51962_nG164e1 , \51963 , \51964_nG164e2 ,
         \51965_nG164e3 , \51966 , \51967_nG18b0b , \51968 , \51969 , \51970_nG164e4 , \51971_nG164e5 , \51972 , \51973_nG164e6 , \51974_nG164e7 ,
         \51975 , \51976_nG18b0d , \51977 , \51978 , \51979_nG164e8 , \51980_nG164e9 , \51981 , \51982_nG164ea , \51983_nG164eb , \51984 ,
         \51985_nG18b0f , \51986 , \51987 , \51988_nG164ec , \51989_nG164ed , \51990 , \51991_nG164ee , \51992_nG164ef , \51993 , \51994_nG18b11 ,
         \51995 , \51996 , \51997_nG164f0 , \51998_nG164f1 , \51999 , \52000_nG164f2 , \52001_nG164f3 , \52002 , \52003_nG18b13 , \52004 ,
         \52005 , \52006_nG164f4 , \52007_nG164f5 , \52008 , \52009_nG164f6 , \52010_nG164f7 , \52011 , \52012_nG18b15 , \52013 , \52014 ,
         \52015_nG164f8 , \52016_nG164f9 , \52017 , \52018_nG164fa , \52019_nG164fb , \52020 , \52021_nG18b17 , \52022 , \52023 , \52024_nG164fc ,
         \52025_nG164fd , \52026 , \52027_nG164fe , \52028_nG164ff , \52029 , \52030_nG18b19 , \52031 , \52032 , \52033_nG16500 , \52034_nG16501 ,
         \52035 , \52036_nG16502 , \52037_nG16503 , \52038 , \52039_nG18b1b , \52040 , \52041 , \52042_nG16504 , \52043_nG16505 , \52044 ,
         \52045_nG16506 , \52046_nG16507 , \52047 , \52048_nG18b1f , \52049 , \52050 , \52051_nG16508 , \52052_nG16509 , \52053 , \52054_nG1650a ,
         \52055_nG1650b , \52056 , \52057_nG18b21 , \52058 , \52059 , \52060_nG1650c , \52061_nG1650d , \52062 , \52063_nG1650e , \52064_nG1650f ,
         \52065 , \52066_nG18b23 , \52067 , \52068 , \52069_nG16510 , \52070_nG16511 , \52071 , \52072_nG16512 , \52073_nG16513 , \52074 ,
         \52075_nG18b25 , \52076 , \52077 , \52078_nG16514 , \52079_nG16515 , \52080 , \52081_nG16516 , \52082_nG16517 , \52083 , \52084_nG18b27 ,
         \52085 , \52086 , \52087_nG16518 , \52088_nG16519 , \52089 , \52090_nG1651a , \52091_nG1651b , \52092 , \52093_nG18b29 , \52094 ,
         \52095 , \52096_nG1651c , \52097_nG1651d , \52098 , \52099_nG1651e , \52100_nG1651f , \52101 , \52102_nG18b2b , \52103 , \52104 ,
         \52105_nG16520 , \52106_nG16521 , \52107 , \52108_nG16522 , \52109_nG16523 , \52110 , \52111_nG18b2d , \52112 , \52113 , \52114_nG16524 ,
         \52115_nG16525 , \52116 , \52117_nG16526 , \52118_nG16527 , \52119 , \52120_nG18b2f , \52121 , \52122 , \52123_nG16528 , \52124_nG16529 ,
         \52125 , \52126_nG1652a , \52127_nG1652b , \52128 , \52129_nG18b31 , \52130 , \52131 , \52132_nG1652c , \52133_nG1652d , \52134 ,
         \52135_nG1652e , \52136_nG1652f , \52137 , \52138_nG18b35 , \52139 , \52140 , \52141_nG16530 , \52142_nG16531 , \52143 , \52144_nG16532 ,
         \52145_nG16533 , \52146 , \52147_nG18b37 , \52148 , \52149 , \52150_nG16534 , \52151_nG16535 , \52152 , \52153_nG16536 , \52154_nG16537 ,
         \52155 , \52156_nG18b39 , \52157 , \52158 , \52159_nG16538 , \52160_nG16539 , \52161 , \52162_nG1653a , \52163_nG1653b , \52164 ,
         \52165_nG18b3b , \52166 , \52167 , \52168_nG1653c , \52169_nG1653d , \52170 , \52171_nG1653e , \52172_nG1653f , \52173 , \52174_nG18b3d ,
         \52175 , \52176 , \52177_nG16540 , \52178_nG16541 , \52179 , \52180_nG16542 , \52181_nG16543 , \52182 , \52183_nG18b3f , \52184 ,
         \52185 , \52186_nG16544 , \52187_nG16545 , \52188 , \52189_nG16546 , \52190_nG16547 , \52191 , \52192_nG18b41 , \52193 , \52194 ,
         \52195_nG16548 , \52196_nG16549 , \52197 , \52198_nG1654a , \52199_nG1654b , \52200 , \52201_nG18b43 , \52202 , \52203 , \52204_nG1654c ,
         \52205_nG1654d , \52206 , \52207_nG1654e , \52208_nG1654f , \52209 , \52210_nG18b45 , \52211 , \52212 , \52213_nG16550 , \52214_nG16551 ,
         \52215 , \52216_nG16552 , \52217_nG16553 , \52218 , \52219_nG18b47 , \52220 , \52221 , \52222_nG16554 , \52223_nG16555 , \52224 ,
         \52225_nG16556 , \52226_nG16557 , \52227 , \52228_nG18b4b , \52229 , \52230 , \52231_nG16558 , \52232_nG16559 , \52233 , \52234_nG1655a ,
         \52235_nG1655b , \52236 , \52237_nG18b4d , \52238 , \52239 , \52240_nG1655c , \52241_nG1655d , \52242 , \52243_nG1655e , \52244_nG1655f ,
         \52245 , \52246_nG18b4f , \52247 , \52248 , \52249_nG16560 , \52250_nG16561 , \52251 , \52252_nG16562 , \52253_nG16563 , \52254 ,
         \52255_nG18b51 , \52256 , \52257 , \52258_nG16564 , \52259_nG16565 , \52260 , \52261_nG16566 , \52262_nG16567 , \52263 , \52264_nG18b53 ,
         \52265 , \52266 , \52267_nG16568 , \52268_nG16569 , \52269 , \52270_nG1656a , \52271_nG1656b , \52272 , \52273_nG18b55 , \52274 ,
         \52275 , \52276_nG1656c , \52277_nG1656d , \52278 , \52279_nG1656e , \52280_nG1656f , \52281 , \52282_nG18b57 , \52283 , \52284 ,
         \52285_nG16570 , \52286_nG16571 , \52287 , \52288_nG16572 , \52289_nG16573 , \52290 , \52291_nG18b59 , \52292 , \52293 , \52294_nG16574 ,
         \52295_nG16575 , \52296 , \52297_nG16576 , \52298_nG16577 , \52299 , \52300_nG18b5b , \52301 , \52302 , \52303_nG16578 , \52304_nG16579 ,
         \52305 , \52306_nG1657a , \52307_nG1657b , \52308 , \52309_nG18b5d , \52310 , \52311 , \52312_nG1657c , \52313_nG1657d , \52314 ,
         \52315_nG1657e , \52316_nG1657f , \52317 , \52318_nG18b61 , \52319 , \52320 , \52321_nG16580 , \52322_nG16581 , \52323 , \52324_nG16582 ,
         \52325_nG16583 , \52326 , \52327_nG18b63 , \52328 , \52329 , \52330_nG16584 , \52331_nG16585 , \52332 , \52333_nG16586 , \52334_nG16587 ,
         \52335 , \52336_nG18b65 , \52337 , \52338 , \52339_nG16588 , \52340_nG16589 , \52341 , \52342_nG1658a , \52343_nG1658b , \52344 ,
         \52345_nG18b67 , \52346 , \52347 , \52348_nG1658c , \52349_nG1658d , \52350 , \52351_nG1658e , \52352_nG1658f , \52353 , \52354_nG18b69 ,
         \52355 , \52356 , \52357_nG16590 , \52358_nG16591 , \52359 , \52360_nG16592 , \52361_nG16593 , \52362 , \52363_nG18b6b , \52364 ,
         \52365 , \52366_nG16594 , \52367_nG16595 , \52368 , \52369_nG16596 , \52370_nG16597 , \52371 , \52372_nG18b6d , \52373 , \52374 ,
         \52375_nG16598 , \52376_nG16599 , \52377 , \52378_nG1659a , \52379_nG1659b , \52380 , \52381_nG18b6f , \52382 , \52383 , \52384_nG1659c ,
         \52385_nG1659d , \52386 , \52387_nG1659e , \52388_nG1659f , \52389 , \52390_nG18b71 , \52391 , \52392 , \52393_nG165a0 , \52394_nG165a1 ,
         \52395 , \52396_nG165a2 , \52397_nG165a3 , \52398 , \52399_nG18b73 , \52400 , \52401 , \52402_nG165a4 , \52403_nG165a5 , \52404 ,
         \52405_nG165a6 , \52406_nG165a7 , \52407 , \52408_nG18b77 , \52409 , \52410 , \52411_nG165a8 , \52412_nG165a9 , \52413 , \52414_nG165aa ,
         \52415_nG165ab , \52416 , \52417_nG18b79 , \52418 , \52419 , \52420_nG165ac , \52421_nG165ad , \52422 , \52423_nG165ae , \52424_nG165af ,
         \52425 , \52426_nG18b7b , \52427 , \52428 , \52429_nG165b0 , \52430_nG165b1 , \52431 , \52432_nG165b2 , \52433_nG165b3 , \52434 ,
         \52435_nG18b7d , \52436 , \52437 , \52438_nG165b4 , \52439_nG165b5 , \52440 , \52441_nG165b6 , \52442_nG165b7 , \52443 , \52444_nG18b7f ,
         \52445 , \52446 , \52447 , \52448_nG163b6 , \52449_nG163b7 , \52450 , \52451 , \52452_nG163b9 , \52453_nG163ba , \52454 ,
         \52455_nG18a87 , \52456 , \52457_nG163bb , \52458_nG163bc , \52459_nG163bd , \52460_nG163be , \52461 , \52462_nG18a9d , \52463 , \52464_nG163bf ,
         \52465_nG163c0 , \52466_nG163c1 , \52467_nG163c2 , \52468 , \52469_nG18ab3 , \52470 , \52471_nG163c3 , \52472_nG163c4 , \52473_nG163c5 , \52474_nG163c6 ,
         \52475 , \52476_nG18ac9 , \52477 , \52478_nG163c7 , \52479_nG163c8 , \52480_nG163c9 , \52481_nG163ca , \52482 , \52483_nG18adf , \52484 ,
         \52485_nG163cb , \52486_nG163cc , \52487_nG163cd , \52488_nG163ce , \52489 , \52490_nG18af5 , \52491 , \52492_nG163cf , \52493_nG163d0 , \52494_nG163d1 ,
         \52495_nG163d2 , \52496 , \52497_nG18b01 , \52498 , \52499_nG163d3 , \52500_nG163d4 , \52501_nG163d5 , \52502_nG163d6 , \52503 , \52504_nG18b03 ,
         \52505 , \52506_nG163d7 , \52507_nG163d8 , \52508_nG163d9 , \52509_nG163da , \52510 , \52511_nG18b05 , \52512 , \52513_nG163db , \52514_nG163dc ,
         \52515_nG163dd , \52516_nG163de , \52517 , \52518_nG18a89 , \52519 , \52520_nG163df , \52521_nG163e0 , \52522_nG163e1 , \52523_nG163e2 , \52524 ,
         \52525_nG18a8b , \52526 , \52527_nG163e3 , \52528_nG163e4 , \52529_nG163e5 , \52530_nG163e6 , \52531 , \52532_nG18a8d , \52533 , \52534_nG163e7 ,
         \52535_nG163e8 , \52536_nG163e9 , \52537_nG163ea , \52538 , \52539_nG18a8f , \52540 , \52541_nG163eb , \52542_nG163ec , \52543_nG163ed , \52544_nG163ee ,
         \52545 , \52546_nG18a91 , \52547 , \52548_nG163ef , \52549_nG163f0 , \52550_nG163f1 , \52551_nG163f2 , \52552 , \52553_nG18a93 , \52554 ,
         \52555_nG163f3 , \52556_nG163f4 , \52557_nG163f5 , \52558_nG163f6 , \52559 , \52560_nG18a95 , \52561 , \52562_nG163f7 , \52563_nG163f8 , \52564_nG163f9 ,
         \52565_nG163fa , \52566 , \52567_nG18a97 , \52568 , \52569_nG163fb , \52570_nG163fc , \52571_nG163fd , \52572_nG163fe , \52573 , \52574_nG18a99 ,
         \52575 , \52576_nG163ff , \52577_nG16400 , \52578_nG16401 , \52579_nG16402 , \52580 , \52581_nG18a9b , \52582 , \52583_nG16403 , \52584_nG16404 ,
         \52585_nG16405 , \52586_nG16406 , \52587 , \52588_nG18a9f , \52589 , \52590_nG16407 , \52591_nG16408 , \52592_nG16409 , \52593_nG1640a , \52594 ,
         \52595_nG18aa1 , \52596 , \52597_nG1640b , \52598_nG1640c , \52599_nG1640d , \52600_nG1640e , \52601 , \52602_nG18aa3 , \52603 , \52604_nG1640f ,
         \52605_nG16410 , \52606_nG16411 , \52607_nG16412 , \52608 , \52609_nG18aa5 , \52610 , \52611_nG16413 , \52612_nG16414 , \52613_nG16415 , \52614_nG16416 ,
         \52615 , \52616_nG18aa7 , \52617 , \52618_nG16417 , \52619_nG16418 , \52620_nG16419 , \52621_nG1641a , \52622 , \52623_nG18aa9 , \52624 ,
         \52625_nG1641b , \52626_nG1641c , \52627_nG1641d , \52628_nG1641e , \52629 , \52630_nG18aab , \52631 , \52632_nG1641f , \52633_nG16420 , \52634_nG16421 ,
         \52635_nG16422 , \52636 , \52637_nG18aad , \52638 , \52639_nG16423 , \52640_nG16424 , \52641_nG16425 , \52642_nG16426 , \52643 , \52644_nG18aaf ,
         \52645 , \52646_nG16427 , \52647_nG16428 , \52648_nG16429 , \52649_nG1642a , \52650 , \52651_nG18ab1 , \52652 , \52653_nG1642b , \52654_nG1642c ,
         \52655_nG1642d , \52656_nG1642e , \52657 , \52658_nG18ab5 , \52659 , \52660_nG1642f , \52661_nG16430 , \52662_nG16431 , \52663_nG16432 , \52664 ,
         \52665_nG18ab7 , \52666 , \52667_nG16433 , \52668_nG16434 , \52669_nG16435 , \52670_nG16436 , \52671 , \52672_nG18ab9 , \52673 , \52674_nG16437 ,
         \52675_nG16438 , \52676_nG16439 , \52677_nG1643a , \52678 , \52679_nG18abb , \52680 , \52681_nG1643b , \52682_nG1643c , \52683_nG1643d , \52684_nG1643e ,
         \52685 , \52686_nG18abd , \52687 , \52688_nG1643f , \52689_nG16440 , \52690_nG16441 , \52691_nG16442 , \52692 , \52693_nG18abf , \52694 ,
         \52695_nG16443 , \52696_nG16444 , \52697_nG16445 , \52698_nG16446 , \52699 , \52700_nG18ac1 , \52701 , \52702_nG16447 , \52703_nG16448 , \52704_nG16449 ,
         \52705_nG1644a , \52706 , \52707_nG18ac3 , \52708 , \52709_nG1644b , \52710_nG1644c , \52711_nG1644d , \52712_nG1644e , \52713 , \52714_nG18ac5 ,
         \52715 , \52716_nG1644f , \52717_nG16450 , \52718_nG16451 , \52719_nG16452 , \52720 , \52721_nG18ac7 , \52722 , \52723_nG16453 , \52724_nG16454 ,
         \52725_nG16455 , \52726_nG16456 , \52727 , \52728_nG18acb , \52729 , \52730_nG16457 , \52731_nG16458 , \52732_nG16459 , \52733_nG1645a , \52734 ,
         \52735_nG18acd , \52736 , \52737_nG1645b , \52738_nG1645c , \52739_nG1645d , \52740_nG1645e , \52741 , \52742_nG18acf , \52743 , \52744_nG1645f ,
         \52745_nG16460 , \52746_nG16461 , \52747_nG16462 , \52748 , \52749_nG18ad1 , \52750 , \52751_nG16463 , \52752_nG16464 , \52753_nG16465 , \52754_nG16466 ,
         \52755 , \52756_nG18ad3 , \52757 , \52758_nG16467 , \52759_nG16468 , \52760_nG16469 , \52761_nG1646a , \52762 , \52763_nG18ad5 , \52764 ,
         \52765_nG1646b , \52766_nG1646c , \52767_nG1646d , \52768_nG1646e , \52769 , \52770_nG18ad7 , \52771 , \52772_nG1646f , \52773_nG16470 , \52774_nG16471 ,
         \52775_nG16472 , \52776 , \52777_nG18ad9 , \52778 , \52779_nG16473 , \52780_nG16474 , \52781_nG16475 , \52782_nG16476 , \52783 , \52784_nG18adb ,
         \52785 , \52786_nG16477 , \52787_nG16478 , \52788_nG16479 , \52789_nG1647a , \52790 , \52791_nG18add , \52792 , \52793_nG1647b , \52794_nG1647c ,
         \52795_nG1647d , \52796_nG1647e , \52797 , \52798_nG18ae1 , \52799 , \52800_nG1647f , \52801_nG16480 , \52802_nG16481 , \52803_nG16482 , \52804 ,
         \52805_nG18ae3 , \52806 , \52807_nG16483 , \52808_nG16484 , \52809_nG16485 , \52810_nG16486 , \52811 , \52812_nG18ae5 , \52813 , \52814_nG16487 ,
         \52815_nG16488 , \52816_nG16489 , \52817_nG1648a , \52818 , \52819_nG18ae7 , \52820 , \52821_nG1648b , \52822_nG1648c , \52823_nG1648d , \52824_nG1648e ,
         \52825 , \52826_nG18ae9 , \52827 , \52828_nG1648f , \52829_nG16490 , \52830_nG16491 , \52831_nG16492 , \52832 , \52833_nG18aeb , \52834 ,
         \52835_nG16493 , \52836_nG16494 , \52837_nG16495 , \52838_nG16496 , \52839 , \52840_nG18aed , \52841 , \52842_nG16497 , \52843_nG16498 , \52844_nG16499 ,
         \52845_nG1649a , \52846 , \52847_nG18aef , \52848 , \52849_nG1649b , \52850_nG1649c , \52851_nG1649d , \52852_nG1649e , \52853 , \52854_nG18af1 ,
         \52855 , \52856_nG1649f , \52857_nG164a0 , \52858_nG164a1 , \52859_nG164a2 , \52860 , \52861_nG18af3 , \52862 , \52863_nG164a3 , \52864_nG164a4 ,
         \52865_nG164a5 , \52866_nG164a6 , \52867 , \52868_nG18af7 , \52869 , \52870_nG164a7 , \52871_nG164a8 , \52872_nG164a9 , \52873_nG164aa , \52874 ,
         \52875_nG18af9 , \52876 , \52877_nG164ab , \52878_nG164ac , \52879_nG164ad , \52880_nG164ae , \52881 , \52882_nG18afb , \52883 , \52884_nG164af ,
         \52885_nG164b0 , \52886_nG164b1 , \52887_nG164b2 , \52888 , \52889_nG18afd , \52890 , \52891_nG164b3 , \52892_nG164b4 , \52893_nG164b5 , \52894_nG164b6 ,
         \52895 , \52896_nG18aff , \52897 , \52898 , \52899_nG162b4 , \52900_nG162b5 , \52901 , \52902_nG162b8 , \52903_nG162b9 , \52904 ,
         \52905_nG18a07 , \52906 , \52907_nG162ba , \52908_nG162bb , \52909_nG162bc , \52910_nG162bd , \52911 , \52912_nG18a1d , \52913 , \52914_nG162be ,
         \52915_nG162bf , \52916_nG162c0 , \52917_nG162c1 , \52918 , \52919_nG18a33 , \52920 , \52921_nG162c2 , \52922_nG162c3 , \52923_nG162c4 , \52924_nG162c5 ,
         \52925 , \52926_nG18a49 , \52927 , \52928_nG162c6 , \52929_nG162c7 , \52930_nG162c8 , \52931_nG162c9 , \52932 , \52933_nG18a5f , \52934 ,
         \52935_nG162ca , \52936_nG162cb , \52937_nG162cc , \52938_nG162cd , \52939 , \52940_nG18a75 , \52941 , \52942_nG162ce , \52943_nG162cf , \52944_nG162d0 ,
         \52945_nG162d1 , \52946 , \52947_nG18a81 , \52948 , \52949_nG162d2 , \52950_nG162d3 , \52951_nG162d4 , \52952_nG162d5 , \52953 , \52954_nG18a83 ,
         \52955 , \52956_nG162d6 , \52957_nG162d7 , \52958_nG162d8 , \52959_nG162d9 , \52960 , \52961_nG18a85 , \52962 , \52963_nG162da , \52964_nG162db ,
         \52965_nG162dc , \52966_nG162dd , \52967 , \52968_nG18a09 , \52969 , \52970_nG162de , \52971_nG162df , \52972_nG162e0 , \52973_nG162e1 , \52974 ,
         \52975_nG18a0b , \52976 , \52977_nG162e2 , \52978_nG162e3 , \52979_nG162e4 , \52980_nG162e5 , \52981 , \52982_nG18a0d , \52983 , \52984_nG162e6 ,
         \52985_nG162e7 , \52986_nG162e8 , \52987_nG162e9 , \52988 , \52989_nG18a0f , \52990 , \52991_nG162ea , \52992_nG162eb , \52993_nG162ec , \52994_nG162ed ,
         \52995 , \52996_nG18a11 , \52997 , \52998_nG162ee , \52999_nG162ef , \53000_nG162f0 , \53001_nG162f1 , \53002 , \53003_nG18a13 , \53004 ,
         \53005_nG162f2 , \53006_nG162f3 , \53007_nG162f4 , \53008_nG162f5 , \53009 , \53010_nG18a15 , \53011 , \53012_nG162f6 , \53013_nG162f7 , \53014_nG162f8 ,
         \53015_nG162f9 , \53016 , \53017_nG18a17 , \53018 , \53019_nG162fa , \53020_nG162fb , \53021_nG162fc , \53022_nG162fd , \53023 , \53024_nG18a19 ,
         \53025 , \53026_nG162fe , \53027_nG162ff , \53028_nG16300 , \53029_nG16301 , \53030 , \53031_nG18a1b , \53032 , \53033_nG16302 , \53034_nG16303 ,
         \53035_nG16304 , \53036_nG16305 , \53037 , \53038_nG18a1f , \53039 , \53040_nG16306 , \53041_nG16307 , \53042_nG16308 , \53043_nG16309 , \53044 ,
         \53045_nG18a21 , \53046 , \53047_nG1630a , \53048_nG1630b , \53049_nG1630c , \53050_nG1630d , \53051 , \53052_nG18a23 , \53053 , \53054_nG1630e ,
         \53055_nG1630f , \53056_nG16310 , \53057_nG16311 , \53058 , \53059_nG18a25 , \53060 , \53061_nG16312 , \53062_nG16313 , \53063_nG16314 , \53064_nG16315 ,
         \53065 , \53066_nG18a27 , \53067 , \53068_nG16316 , \53069_nG16317 , \53070_nG16318 , \53071_nG16319 , \53072 , \53073_nG18a29 , \53074 ,
         \53075_nG1631a , \53076_nG1631b , \53077_nG1631c , \53078_nG1631d , \53079 , \53080_nG18a2b , \53081 , \53082_nG1631e , \53083_nG1631f , \53084_nG16320 ,
         \53085_nG16321 , \53086 , \53087_nG18a2d , \53088 , \53089_nG16322 , \53090_nG16323 , \53091_nG16324 , \53092_nG16325 , \53093 , \53094_nG18a2f ,
         \53095 , \53096_nG16326 , \53097_nG16327 , \53098_nG16328 , \53099_nG16329 , \53100 , \53101_nG18a31 , \53102 , \53103_nG1632a , \53104_nG1632b ,
         \53105_nG1632c , \53106_nG1632d , \53107 , \53108_nG18a35 , \53109 , \53110_nG1632e , \53111_nG1632f , \53112_nG16330 , \53113_nG16331 , \53114 ,
         \53115_nG18a37 , \53116 ;
buf \U$labaj5648 ( R_25610_96cc360, \42505 );
buf \U$labaj5649 ( R_25642_95f0d48, \42508 );
buf \U$labaj5650 ( R_25644_9598060, \42511 );
buf \U$labaj5651 ( R_25646_95984f8, \42514 );
buf \U$labaj5652 ( R_25614_953c348, \42517 );
buf \U$labaj5653 ( R_25616_96251f8, \42522 );
buf \U$labaj5654 ( R_25618_96ed6b0, \42527 );
buf \U$labaj5655 ( R_2561a_95f00d0, \42532 );
buf \U$labaj5656 ( R_2561c_95f0418, \42537 );
buf \U$labaj5657 ( R_2561e_95f0760, \42542 );
buf \U$labaj5658 ( R_25620_953c3f0, \42547 );
buf \U$labaj5659 ( R_25622_953c690, \42552 );
buf \U$labaj5660 ( R_25612_953c9d8, \42557 );
buf \U$labaj5661 ( R_25624_95f08b0, \42562 );
buf \U$labaj5662 ( R_25626_953ca80, \42567 );
buf \U$labaj5663 ( R_25628_96253f0, \42572 );
buf \U$labaj5664 ( R_2562a_9632be8, \42577 );
buf \U$labaj5665 ( R_253fc_9d20ef0, \42603 );
buf \U$labaj5666 ( R_25412_9530108, \42612 );
buf \U$labaj5667 ( R_25428_95f75a0, \42621 );
buf \U$labaj5668 ( R_2543e_95301b0, \42630 );
buf \U$labaj5669 ( R_25454_95304f8, \42639 );
buf \U$labaj5670 ( R_2546a_9533198, \42648 );
buf \U$labaj5671 ( R_25474_95332e8, \42657 );
buf \U$labaj5672 ( R_25476_96dee60, \42666 );
buf \U$labaj5673 ( R_25478_95f7798, \42675 );
buf \U$labaj5674 ( R_2547a_96def08, \42684 );
buf \U$labaj5675 ( R_253fe_95f7990, \42693 );
buf \U$labaj5676 ( R_25400_9d21190, \42702 );
buf \U$labaj5677 ( R_25402_9d21388, \42711 );
buf \U$labaj5678 ( R_25404_9589e90, \42720 );
buf \U$labaj5679 ( R_25406_9d21430, \42729 );
buf \U$labaj5680 ( R_25408_9533780, \42738 );
buf \U$labaj5681 ( R_2540a_9533b70, \42747 );
buf \U$labaj5682 ( R_2540c_9d216d0, \42756 );
buf \U$labaj5683 ( R_2540e_958a5c8, \42765 );
buf \U$labaj5684 ( R_25410_96defb0, \42774 );
buf \U$labaj5685 ( R_25414_9d21778, \42783 );
buf \U$labaj5686 ( R_25416_9d21cb8, \42792 );
buf \U$labaj5687 ( R_25418_95f7ae0, \42801 );
buf \U$labaj5688 ( R_2541a_9d21d60, \42810 );
buf \U$labaj5689 ( R_2541c_96df100, \42819 );
buf \U$labaj5690 ( R_2541e_9d221f8, \42828 );
buf \U$labaj5691 ( R_25420_958ac58, \42837 );
buf \U$labaj5692 ( R_25422_95f7b88, \42846 );
buf \U$labaj5693 ( R_25424_9533c18, \42855 );
buf \U$labaj5694 ( R_25426_958b630, \42864 );
buf \U$labaj5695 ( R_2542a_9d222a0, \42873 );
buf \U$labaj5696 ( R_2542c_9533d68, \42882 );
buf \U$labaj5697 ( R_2542e_95f7c30, \42891 );
buf \U$labaj5698 ( R_25430_9d22498, \42900 );
buf \U$labaj5699 ( R_25432_9d22540, \42909 );
buf \U$labaj5700 ( R_25434_9533f60, \42918 );
buf \U$labaj5701 ( R_25436_96df1a8, \42927 );
buf \U$labaj5702 ( R_25438_95f7f78, \42936 );
buf \U$labaj5703 ( R_2543a_9534008, \42945 );
buf \U$labaj5704 ( R_2543c_9534200, \42954 );
buf \U$labaj5705 ( R_25440_95f80c8, \42963 );
buf \U$labaj5706 ( R_25442_96df250, \42972 );
buf \U$labaj5707 ( R_25444_9d22690, \42981 );
buf \U$labaj5708 ( R_25446_95fa438, \42990 );
buf \U$labaj5709 ( R_25448_95fa4e0, \42999 );
buf \U$labaj5710 ( R_2544a_958bcc0, \43008 );
buf \U$labaj5711 ( R_2544c_9d22738, \43017 );
buf \U$labaj5712 ( R_2544e_9d227e0, \43026 );
buf \U$labaj5713 ( R_25450_9d22888, \43035 );
buf \U$labaj5714 ( R_25452_9d22930, \43044 );
buf \U$labaj5715 ( R_25456_9d229d8, \43053 );
buf \U$labaj5716 ( R_25458_95fa588, \43062 );
buf \U$labaj5717 ( R_2545a_9534350, \43071 );
buf \U$labaj5718 ( R_2545c_95fa828, \43080 );
buf \U$labaj5719 ( R_2545e_9d22a80, \43089 );
buf \U$labaj5720 ( R_25460_96df2f8, \43098 );
buf \U$labaj5721 ( R_25462_96df3a0, \43107 );
buf \U$labaj5722 ( R_25464_95343f8, \43116 );
buf \U$labaj5723 ( R_25466_95fa8d0, \43125 );
buf \U$labaj5724 ( R_25468_95faac8, \43134 );
buf \U$labaj5725 ( R_2546c_958bd68, \43143 );
buf \U$labaj5726 ( R_2546e_958be10, \43152 );
buf \U$labaj5727 ( R_25470_95fab70, \43161 );
buf \U$labaj5728 ( R_25472_9d22b28, \43170 );
buf \U$labaj5729 ( R_2547c_958beb8, \43181 );
buf \U$labaj5730 ( R_25492_9d22bd0, \43188 );
buf \U$labaj5731 ( R_254a8_958bf60, \43195 );
buf \U$labaj5732 ( R_254be_9d22c78, \43202 );
buf \U$labaj5733 ( R_254d4_9d22dc8, \43209 );
buf \U$labaj5734 ( R_254ea_9d22e70, \43216 );
buf \U$labaj5735 ( R_254f4_958c0b0, \43223 );
buf \U$labaj5736 ( R_254f6_9d22f18, \43230 );
buf \U$labaj5737 ( R_254f8_958c158, \43237 );
buf \U$labaj5738 ( R_254fa_9d22fc0, \43244 );
buf \U$labaj5739 ( R_2547e_958c200, \43251 );
buf \U$labaj5740 ( R_25480_9d23068, \43258 );
buf \U$labaj5741 ( R_25482_9d231b8, \43265 );
buf \U$labaj5742 ( R_25484_958c2a8, \43272 );
buf \U$labaj5743 ( R_25486_958c350, \43279 );
buf \U$labaj5744 ( R_25488_9d23458, \43286 );
buf \U$labaj5745 ( R_2548a_958c4a0, \43293 );
buf \U$labaj5746 ( R_2548c_9d235a8, \43300 );
buf \U$labaj5747 ( R_2548e_9d236f8, \43307 );
buf \U$labaj5748 ( R_25490_958c548, \43314 );
buf \U$labaj5749 ( R_25494_958c5f0, \43321 );
buf \U$labaj5750 ( R_25496_9d237a0, \43328 );
buf \U$labaj5751 ( R_25498_958c698, \43335 );
buf \U$labaj5752 ( R_2549a_958f728, \43342 );
buf \U$labaj5753 ( R_2549c_9d23848, \43349 );
buf \U$labaj5754 ( R_2549e_958f7d0, \43356 );
buf \U$labaj5755 ( R_254a0_958f878, \43363 );
buf \U$labaj5756 ( R_254a2_9d23998, \43370 );
buf \U$labaj5757 ( R_254a4_9d23ae8, \43377 );
buf \U$labaj5758 ( R_254a6_9d23c38, \43384 );
buf \U$labaj5759 ( R_254aa_9d23d88, \43391 );
buf \U$labaj5760 ( R_254ac_9d23e30, \43398 );
buf \U$labaj5761 ( R_254ae_9d23f80, \43405 );
buf \U$labaj5762 ( R_254b0_9d24028, \43412 );
buf \U$labaj5763 ( R_254b2_9d240d0, \43419 );
buf \U$labaj5764 ( R_254b4_9d24220, \43426 );
buf \U$labaj5765 ( R_254b6_9d242c8, \43433 );
buf \U$labaj5766 ( R_254b8_9590988, \43440 );
buf \U$labaj5767 ( R_254ba_9590a30, \43447 );
buf \U$labaj5768 ( R_254bc_9590cd0, \43454 );
buf \U$labaj5769 ( R_254c0_9d24418, \43461 );
buf \U$labaj5770 ( R_254c2_9590d78, \43468 );
buf \U$labaj5771 ( R_254c4_9590f70, \43475 );
buf \U$labaj5772 ( R_254c6_9591178, \43482 );
buf \U$labaj5773 ( R_254c8_9d24568, \43489 );
buf \U$labaj5774 ( R_254ca_9d24bf8, \43496 );
buf \U$labaj5775 ( R_254cc_9d25090, \43503 );
buf \U$labaj5776 ( R_254ce_95916b8, \43510 );
buf \U$labaj5777 ( R_254d0_9591808, \43517 );
buf \U$labaj5778 ( R_254d2_9d251e0, \43524 );
buf \U$labaj5779 ( R_254d6_9d25f10, \43531 );
buf \U$labaj5780 ( R_254d8_9d25fb8, \43538 );
buf \U$labaj5781 ( R_254da_95918b0, \43545 );
buf \U$labaj5782 ( R_254dc_9d265a0, \43552 );
buf \U$labaj5783 ( R_254de_9591958, \43559 );
buf \U$labaj5784 ( R_254e0_9d26990, \43566 );
buf \U$labaj5785 ( R_254e2_9d26c30, \43573 );
buf \U$labaj5786 ( R_254e4_9591a00, \43580 );
buf \U$labaj5787 ( R_254e6_95347e8, \43587 );
buf \U$labaj5788 ( R_254e8_9591b50, \43594 );
buf \U$labaj5789 ( R_254ec_9591bf8, \43601 );
buf \U$labaj5790 ( R_254ee_9d26d80, \43608 );
buf \U$labaj5791 ( R_254f0_9d27368, \43615 );
buf \U$labaj5792 ( R_254f2_9d27410, \43622 );
buf \U$labaj5793 ( R_254fc_96df4f0, \43631 );
buf \U$labaj5794 ( R_25512_9d276b0, \43638 );
buf \U$labaj5795 ( R_25528_96df598, \43645 );
buf \U$labaj5796 ( R_2553e_9534890, \43652 );
buf \U$labaj5797 ( R_25554_9d27c98, \43659 );
buf \U$labaj5798 ( R_2556a_96df640, \43666 );
buf \U$labaj5799 ( R_25574_9d27de8, \43673 );
buf \U$labaj5800 ( R_25576_96df6e8, \43680 );
buf \U$labaj5801 ( R_25578_9534bd8, \43687 );
buf \U$labaj5802 ( R_2557a_96df838, \43694 );
buf \U$labaj5803 ( R_254fe_96dfad8, \43701 );
buf \U$labaj5804 ( R_25500_9534d28, \43708 );
buf \U$labaj5805 ( R_25502_9534dd0, \43715 );
buf \U$labaj5806 ( R_25504_9534f20, \43722 );
buf \U$labaj5807 ( R_25506_9d281d8, \43729 );
buf \U$labaj5808 ( R_25508_96dfb80, \43736 );
buf \U$labaj5809 ( R_2550a_9d28328, \43743 );
buf \U$labaj5810 ( R_2550c_9d283d0, \43750 );
buf \U$labaj5811 ( R_2550e_96dfc28, \43757 );
buf \U$labaj5812 ( R_25510_9534fc8, \43764 );
buf \U$labaj5813 ( R_25514_96dfcd0, \43771 );
buf \U$labaj5814 ( R_25516_9d28520, \43778 );
buf \U$labaj5815 ( R_25518_96dfe20, \43785 );
buf \U$labaj5816 ( R_2551a_96dfec8, \43792 );
buf \U$labaj5817 ( R_2551c_9535070, \43799 );
buf \U$labaj5818 ( R_2551e_95351c0, \43806 );
buf \U$labaj5819 ( R_25520_9535268, \43813 );
buf \U$labaj5820 ( R_25522_96dff70, \43820 );
buf \U$labaj5821 ( R_25524_96e0018, \43827 );
buf \U$labaj5822 ( R_25526_96e00c0, \43834 );
buf \U$labaj5823 ( R_2552a_9535310, \43841 );
buf \U$labaj5824 ( R_2552c_96e0168, \43848 );
buf \U$labaj5825 ( R_2552e_96e0210, \43855 );
buf \U$labaj5826 ( R_25530_96e02b8, \43862 );
buf \U$labaj5827 ( R_25532_96e0408, \43869 );
buf \U$labaj5828 ( R_25534_96e0558, \43876 );
buf \U$labaj5829 ( R_25536_96e0600, \43883 );
buf \U$labaj5830 ( R_25538_9535658, \43890 );
buf \U$labaj5831 ( R_2553a_9d289b8, \43897 );
buf \U$labaj5832 ( R_2553c_96e06a8, \43904 );
buf \U$labaj5833 ( R_25540_95358f8, \43911 );
buf \U$labaj5834 ( R_25542_96e0750, \43918 );
buf \U$labaj5835 ( R_25544_96e0b40, \43925 );
buf \U$labaj5836 ( R_25546_96e0be8, \43932 );
buf \U$labaj5837 ( R_25548_96e0c90, \43939 );
buf \U$labaj5838 ( R_2554a_96e0d38, \43946 );
buf \U$labaj5839 ( R_2554c_95359a0, \43953 );
buf \U$labaj5840 ( R_2554e_9d28a60, \43960 );
buf \U$labaj5841 ( R_25550_96e0e88, \43967 );
buf \U$labaj5842 ( R_25552_9535a48, \43974 );
buf \U$labaj5843 ( R_25556_96e0f30, \43981 );
buf \U$labaj5844 ( R_25558_9535b98, \43988 );
buf \U$labaj5845 ( R_2555a_9d28c58, \43995 );
buf \U$labaj5846 ( R_2555c_96e0fd8, \44002 );
buf \U$labaj5847 ( R_2555e_9d28d00, \44009 );
buf \U$labaj5848 ( R_25560_9535c40, \44016 );
buf \U$labaj5849 ( R_25562_95362d0, \44023 );
buf \U$labaj5850 ( R_25564_9536810, \44030 );
buf \U$labaj5851 ( R_25566_9536a08, \44037 );
buf \U$labaj5852 ( R_25568_96e1080, \44044 );
buf \U$labaj5853 ( R_2556c_96e1128, \44051 );
buf \U$labaj5854 ( R_2556e_9d28ef8, \44058 );
buf \U$labaj5855 ( R_25570_96e11d0, \44065 );
buf \U$labaj5856 ( R_25572_96e1c50, \44072 );
buf \U$labaj5857 ( R_2557c_9591d48, \44081 );
buf \U$labaj5858 ( R_25592_9591df0, \44088 );
buf \U$labaj5859 ( R_255a8_96e2e08, \44095 );
buf \U$labaj5860 ( R_255be_9591e98, \44102 );
buf \U$labaj5861 ( R_255d4_9591f40, \44109 );
buf \U$labaj5862 ( R_255ea_96e3690, \44116 );
buf \U$labaj5863 ( R_255f4_96e6918, \44123 );
buf \U$labaj5864 ( R_255f6_96e69c0, \44130 );
buf \U$labaj5865 ( R_255f8_9d29048, \44137 );
buf \U$labaj5866 ( R_255fa_9d28718, \44144 );
buf \U$labaj5867 ( R_2557e_9591fe8, \44151 );
buf \U$labaj5868 ( R_25580_96e6fa8, \44158 );
buf \U$labaj5869 ( R_25582_96e72f0, \44165 );
buf \U$labaj5870 ( R_25584_9d287c0, \44172 );
buf \U$labaj5871 ( R_25586_9592090, \44179 );
buf \U$labaj5872 ( R_25588_9592138, \44186 );
buf \U$labaj5873 ( R_2558a_96e7398, \44193 );
buf \U$labaj5874 ( R_2558c_9d28868, \44200 );
buf \U$labaj5875 ( R_2558e_9d290f0, \44207 );
buf \U$labaj5876 ( R_25590_9d29240, \44214 );
buf \U$labaj5877 ( R_25594_96e7cc8, \44221 );
buf \U$labaj5878 ( R_25596_95921e0, \44228 );
buf \U$labaj5879 ( R_25598_9592288, \44235 );
buf \U$labaj5880 ( R_2559a_9592330, \44242 );
buf \U$labaj5881 ( R_2559c_96e82b0, \44249 );
buf \U$labaj5882 ( R_2559e_9d292e8, \44256 );
buf \U$labaj5883 ( R_255a0_9d2dfb0, \44263 );
buf \U$labaj5884 ( R_255a2_9592528, \44270 );
buf \U$labaj5885 ( R_255a4_9592678, \44277 );
buf \U$labaj5886 ( R_255a6_9d2e058, \44284 );
buf \U$labaj5887 ( R_255aa_96e8358, \44291 );
buf \U$labaj5888 ( R_255ac_9592918, \44298 );
buf \U$labaj5889 ( R_255ae_96e86a0, \44305 );
buf \U$labaj5890 ( R_255b0_9d2e988, \44312 );
buf \U$labaj5891 ( R_255b2_9d29390, \44319 );
buf \U$labaj5892 ( R_255b4_9d2ec28, \44326 );
buf \U$labaj5893 ( R_255b6_9d294e0, \44333 );
buf \U$labaj5894 ( R_255b8_9d2f360, \44340 );
buf \U$labaj5895 ( R_255ba_9592a68, \44347 );
buf \U$labaj5896 ( R_255bc_9592b10, \44354 );
buf \U$labaj5897 ( R_255c0_9d30128, \44361 );
buf \U$labaj5898 ( R_255c2_9592c60, \44368 );
buf \U$labaj5899 ( R_255c4_96e8940, \44375 );
buf \U$labaj5900 ( R_255c6_96e89e8, \44382 );
buf \U$labaj5901 ( R_255c8_9d30278, \44389 );
buf \U$labaj5902 ( R_255ca_96e8be0, \44396 );
buf \U$labaj5903 ( R_255cc_9592f00, \44403 );
buf \U$labaj5904 ( R_255ce_9d29588, \44410 );
buf \U$labaj5905 ( R_255d0_9d296d8, \44417 );
buf \U$labaj5906 ( R_255d2_9d30518, \44424 );
buf \U$labaj5907 ( R_255d6_9d29828, \44431 );
buf \U$labaj5908 ( R_255d8_96e9120, \44438 );
buf \U$labaj5909 ( R_255da_96e93c0, \44445 );
buf \U$labaj5910 ( R_255dc_96e9510, \44452 );
buf \U$labaj5911 ( R_255de_9d307b8, \44459 );
buf \U$labaj5912 ( R_255e0_9d29cc0, \44466 );
buf \U$labaj5913 ( R_255e2_9592fa8, \44473 );
buf \U$labaj5914 ( R_255e4_9593050, \44480 );
buf \U$labaj5915 ( R_255e6_96e9858, \44487 );
buf \U$labaj5916 ( R_255e8_96e9a50, \44494 );
buf \U$labaj5917 ( R_255ec_95930f8, \44501 );
buf \U$labaj5918 ( R_255ee_9d29eb8, \44508 );
buf \U$labaj5919 ( R_255f0_96ea038, \44515 );
buf \U$labaj5920 ( R_255f2_95931a0, \44522 );
buf \U$labaj5921 ( R_253bc_96eacb0, \44530 );
buf \U$labaj5922 ( R_253be_9593248, \44536 );
buf \U$labaj5923 ( R_253c0_9d29f60, \44542 );
buf \U$labaj5924 ( R_253c2_95932f0, \44548 );
buf \U$labaj5925 ( R_253c4_96eae00, \44554 );
buf \U$labaj5926 ( R_253c6_9536b58, \44560 );
buf \U$labaj5927 ( R_253c8_9593398, \44566 );
buf \U$labaj5928 ( R_253ca_9d2a350, \44572 );
buf \U$labaj5929 ( R_253cc_b7dc210, \44577 );
buf \U$labaj5930 ( R_253ce_b7dcd38, \44582 );
buf \U$labaj5931 ( R_253d0_b7dcde0, \44587 );
buf \U$labaj5932 ( R_253d2_9593590, \44592 );
buf \U$labaj5933 ( R_253d4_96376b8, \44597 );
buf \U$labaj5934 ( R_253d6_9d2a4a0, \44602 );
buf \U$labaj5935 ( R_253d8_9596038, \44607 );
buf \U$labaj5936 ( R_253da_b7dc2b8, \44612 );
buf \U$labaj5937 ( R_253dc_96eb0a0, \44617 );
buf \U$labaj5938 ( R_253de_9596578, \44622 );
buf \U$labaj5939 ( R_253e0_9536f48, \44627 );
buf \U$labaj5940 ( R_253e2_96eb298, \44632 );
buf \U$labaj5941 ( R_253e4_9537098, \44637 );
buf \U$labaj5942 ( R_253e6_96eb340, \44642 );
buf \U$labaj5943 ( R_253e8_95373e0, \44647 );
buf \U$labaj5944 ( R_253ea_9596a10, \44652 );
buf \U$labaj5945 ( R_253ec_9d30860, \44657 );
buf \U$labaj5946 ( R_253ee_9ef0090, \44662 );
buf \U$labaj5947 ( R_253f0_9d30f98, \44667 );
buf \U$labaj5948 ( R_253f2_9ef05d0, \44672 );
buf \U$labaj5949 ( R_253f4_9d31040, \44677 );
buf \U$labaj5950 ( R_253f6_9d31238, \44682 );
buf \U$labaj5951 ( R_253f8_9d314d8, \44687 );
buf \U$labaj5952 ( R_253fa_9d316d0, \44692 );
buf \U$labaj5953 ( R_25666_96346d0, \44699 );
buf \U$labaj5954 ( R_1a4_b821b50, \44769 );
buf \U$labaj5955 ( R_1a3_b821aa8, \44806 );
buf \U$labaj5956 ( R_23ca4_96329f0, \44833 );
buf \U$labaj5957 ( R_23cba_9f596e0, \44842 );
buf \U$labaj5958 ( R_23cd0_962b7c0, \44851 );
buf \U$labaj5959 ( R_23ce6_955f268, \44860 );
buf \U$labaj5960 ( R_23cfc_9f5c4d0, \44869 );
buf \U$labaj5961 ( R_23d12_9d225e8, \44878 );
buf \U$labaj5962 ( R_23d1c_962b910, \44887 );
buf \U$labaj5963 ( R_23d1e_95a3470, \44896 );
buf \U$labaj5964 ( R_23d20_9632c90, \44905 );
buf \U$labaj5965 ( R_23d22_95a3710, \44914 );
buf \U$labaj5966 ( R_23ca6_9ee76c0, \44923 );
buf \U$labaj5967 ( R_23ca8_9ee7810, \44932 );
buf \U$labaj5968 ( R_23caa_9ee78b8, \44941 );
buf \U$labaj5969 ( R_23cac_9ee8140, \44950 );
buf \U$labaj5970 ( R_23cae_962bbb0, \44959 );
buf \U$labaj5971 ( R_23cb0_9ee8920, \44968 );
buf \U$labaj5972 ( R_23cb2_9d22d20, \44977 );
buf \U$labaj5973 ( R_23cb4_9ee8bc0, \44986 );
buf \U$labaj5974 ( R_23cb6_9632d38, \44995 );
buf \U$labaj5975 ( R_23cb8_9d23110, \45004 );
buf \U$labaj5976 ( R_23cbc_962bc58, \45013 );
buf \U$labaj5977 ( R_23cbe_9ee9ad8, \45022 );
buf \U$labaj5978 ( R_23cc0_9d23260, \45031 );
buf \U$labaj5979 ( R_23cc2_9632f30, \45040 );
buf \U$labaj5980 ( R_23cc4_9eec430, \45049 );
buf \U$labaj5981 ( R_23cc6_9d23308, \45058 );
buf \U$labaj5982 ( R_23cc8_9eef4c0, \45067 );
buf \U$labaj5983 ( R_23cca_9eefca0, \45076 );
buf \U$labaj5984 ( R_23ccc_9d23650, \45085 );
buf \U$labaj5985 ( R_23cce_9ef0678, \45094 );
buf \U$labaj5986 ( R_23cd2_95a3908, \45103 );
buf \U$labaj5987 ( R_23cd4_962bd00, \45112 );
buf \U$labaj5988 ( R_23cd6_9632fd8, \45121 );
buf \U$labaj5989 ( R_23cd8_962be50, \45130 );
buf \U$labaj5990 ( R_23cda_96331d0, \45139 );
buf \U$labaj5991 ( R_23cdc_962bef8, \45148 );
buf \U$labaj5992 ( R_23cde_9d30ef0, \45157 );
buf \U$labaj5993 ( R_23ce0_9d238f0, \45166 );
buf \U$labaj5994 ( R_23ce2_9d23b90, \45175 );
buf \U$labaj5995 ( R_23ce4_962bfa0, \45184 );
buf \U$labaj5996 ( R_23ce8_962c048, \45193 );
buf \U$labaj5997 ( R_23cea_95a3a58, \45202 );
buf \U$labaj5998 ( R_23cec_9d23ed8, \45211 );
buf \U$labaj5999 ( R_23cee_9ef09c0, \45220 );
buf \U$labaj6000 ( R_23cf0_9ef4380, \45229 );
buf \U$labaj6001 ( R_23cf2_95a3ba8, \45238 );
buf \U$labaj6002 ( R_23cf4_9ef4a10, \45247 );
buf \U$labaj6003 ( R_23cf6_962c0f0, \45256 );
buf \U$labaj6004 ( R_23cf8_96c3060, \45265 );
buf \U$labaj6005 ( R_23cfa_96c6d68, \45274 );
buf \U$labaj6006 ( R_23cfe_9d310e8, \45283 );
buf \U$labaj6007 ( R_23d00_96c72a8, \45292 );
buf \U$labaj6008 ( R_23d02_962c390, \45301 );
buf \U$labaj6009 ( R_23d04_96c74a0, \45310 );
buf \U$labaj6010 ( R_23d06_962da88, \45319 );
buf \U$labaj6011 ( R_23d08_9d24178, \45328 );
buf \U$labaj6012 ( R_23d0a_962df20, \45337 );
buf \U$labaj6013 ( R_23d0c_9633278, \45346 );
buf \U$labaj6014 ( R_23d0e_9633320, \45355 );
buf \U$labaj6015 ( R_23d10_95a3e48, \45364 );
buf \U$labaj6016 ( R_23d14_95a4040, \45373 );
buf \U$labaj6017 ( R_23d16_9d24370, \45382 );
buf \U$labaj6018 ( R_23d18_96c7e78, \45391 );
buf \U$labaj6019 ( R_23d1a_96333c8, \45400 );
buf \U$labaj6020 ( R_23d24_9633470, \45411 );
buf \U$labaj6021 ( R_23d3a_9633518, \45418 );
buf \U$labaj6022 ( R_23d50_962dfc8, \45425 );
buf \U$labaj6023 ( R_23d66_9629b88, \45432 );
buf \U$labaj6024 ( R_23d7c_95547c8, \45439 );
buf \U$labaj6025 ( R_23d92_96335c0, \45446 );
buf \U$labaj6026 ( R_23d9c_96337b8, \45453 );
buf \U$labaj6027 ( R_23d9e_9633908, \45460 );
buf \U$labaj6028 ( R_23da0_9633a58, \45467 );
buf \U$labaj6029 ( R_23da2_962e7a8, \45474 );
buf \U$labaj6030 ( R_23d26_9554870, \45481 );
buf \U$labaj6031 ( R_23d28_962a560, \45488 );
buf \U$labaj6032 ( R_23d2a_962ee38, \45495 );
buf \U$labaj6033 ( R_23d2c_962a8a8, \45502 );
buf \U$labaj6034 ( R_23d2e_962f2d0, \45509 );
buf \U$labaj6035 ( R_23d30_95549c0, \45516 );
buf \U$labaj6036 ( R_23d32_9633cf8, \45523 );
buf \U$labaj6037 ( R_23d34_962f4c8, \45530 );
buf \U$labaj6038 ( R_23d36_9633da0, \45537 );
buf \U$labaj6039 ( R_23d38_9633e48, \45544 );
buf \U$labaj6040 ( R_23d3c_9633ef0, \45551 );
buf \U$labaj6041 ( R_23d3e_962c4e0, \45558 );
buf \U$labaj6042 ( R_23d40_9554bb8, \45565 );
buf \U$labaj6043 ( R_23d42_9554d08, \45572 );
buf \U$labaj6044 ( R_23d44_9634040, \45579 );
buf \U$labaj6045 ( R_23d46_962f6c0, \45586 );
buf \U$labaj6046 ( R_23d48_9554f00, \45593 );
buf \U$labaj6047 ( R_23d4a_962c8d0, \45600 );
buf \U$labaj6048 ( R_23d4c_9635000, \45607 );
buf \U$labaj6049 ( R_23d4e_962fab0, \45614 );
buf \U$labaj6050 ( R_23d52_95552f0, \45621 );
buf \U$labaj6051 ( R_23d54_96350a8, \45628 );
buf \U$labaj6052 ( R_23d56_96351f8, \45635 );
buf \U$labaj6053 ( R_23d58_962fc00, \45642 );
buf \U$labaj6054 ( R_23d5a_95554e8, \45649 );
buf \U$labaj6055 ( R_23d5c_9555638, \45656 );
buf \U$labaj6056 ( R_23d5e_9635540, \45663 );
buf \U$labaj6057 ( R_23d60_96355e8, \45670 );
buf \U$labaj6058 ( R_23d62_9635738, \45677 );
buf \U$labaj6059 ( R_23d64_96359d8, \45684 );
buf \U$labaj6060 ( R_23d68_962ca20, \45691 );
buf \U$labaj6061 ( R_23d6a_9635f18, \45698 );
buf \U$labaj6062 ( R_23d6c_962ff48, \45705 );
buf \U$labaj6063 ( R_23d6e_9636068, \45712 );
buf \U$labaj6064 ( R_23d70_96363b0, \45719 );
buf \U$labaj6065 ( R_23d72_9636ae8, \45726 );
buf \U$labaj6066 ( R_23d74_9637220, \45733 );
buf \U$labaj6067 ( R_23d76_9637e98, \45740 );
buf \U$labaj6068 ( R_23d78_9638b10, \45747 );
buf \U$labaj6069 ( R_23d7a_962d4a0, \45754 );
buf \U$labaj6070 ( R_23d7e_96305d8, \45761 );
buf \U$labaj6071 ( R_23d80_9638bb8, \45768 );
buf \U$labaj6072 ( R_23d82_9638fa8, \45775 );
buf \U$labaj6073 ( R_23d84_962d548, \45782 );
buf \U$labaj6074 ( R_23d86_9639398, \45789 );
buf \U$labaj6075 ( R_23d88_95556e0, \45796 );
buf \U$labaj6076 ( R_23d8a_9639440, \45803 );
buf \U$labaj6077 ( R_23d8c_9d18d00, \45810 );
buf \U$labaj6078 ( R_23d8e_9d19d68, \45817 );
buf \U$labaj6079 ( R_23d90_9630a70, \45824 );
buf \U$labaj6080 ( R_23d94_9d1a008, \45831 );
buf \U$labaj6081 ( R_23d96_9d1a350, \45838 );
buf \U$labaj6082 ( R_23d98_9d1a9e0, \45845 );
buf \U$labaj6083 ( R_23d9a_96314f0, \45852 );
buf \U$labaj6084 ( R_23da4_9634430, \45861 );
buf \U$labaj6085 ( R_23dba_95558d8, \45868 );
buf \U$labaj6086 ( R_23dd0_9555a28, \45875 );
buf \U$labaj6087 ( R_23de6_9d1ac80, \45882 );
buf \U$labaj6088 ( R_23dfc_962d9e0, \45889 );
buf \U$labaj6089 ( R_23e12_9555b78, \45896 );
buf \U$labaj6090 ( R_23e1c_96344d8, \45903 );
buf \U$labaj6091 ( R_23e1e_9555e18, \45910 );
buf \U$labaj6092 ( R_23e20_9d1b070, \45917 );
buf \U$labaj6093 ( R_23e22_9d1b8f8, \45924 );
buf \U$labaj6094 ( R_23da6_9634a18, \45931 );
buf \U$labaj6095 ( R_23da8_9555f68, \45938 );
buf \U$labaj6096 ( R_23daa_9635150, \45945 );
buf \U$labaj6097 ( R_23dac_96352a0, \45952 );
buf \U$labaj6098 ( R_23dae_9556010, \45959 );
buf \U$labaj6099 ( R_23db0_9557078, \45966 );
buf \U$labaj6100 ( R_23db2_96353f0, \45973 );
buf \U$labaj6101 ( R_23db4_9d1ba48, \45980 );
buf \U$labaj6102 ( R_23db6_962db30, \45987 );
buf \U$labaj6103 ( R_23db8_96357e0, \45994 );
buf \U$labaj6104 ( R_23dbc_9559730, \46001 );
buf \U$labaj6105 ( R_23dbe_955bde8, \46008 );
buf \U$labaj6106 ( R_23dc0_955dd68, \46015 );
buf \U$labaj6107 ( R_23dc2_9d1baf0, \46022 );
buf \U$labaj6108 ( R_23dc4_955e158, \46029 );
buf \U$labaj6109 ( R_23dc6_9638db0, \46036 );
buf \U$labaj6110 ( R_23dc8_9d1bb98, \46043 );
buf \U$labaj6111 ( R_23dca_9639248, \46050 );
buf \U$labaj6112 ( R_23dcc_9d1bce8, \46057 );
buf \U$labaj6113 ( R_23dce_96c81c0, \46064 );
buf \U$labaj6114 ( R_23dd2_955e4a0, \46071 );
buf \U$labaj6115 ( R_23dd4_955ea88, \46078 );
buf \U$labaj6116 ( R_23dd6_96392f0, \46085 );
buf \U$labaj6117 ( R_23dd8_9d15d18, \46092 );
buf \U$labaj6118 ( R_23dda_955ee78, \46099 );
buf \U$labaj6119 ( R_23ddc_9d168e8, \46106 );
buf \U$labaj6120 ( R_23dde_9d16ae0, \46113 );
buf \U$labaj6121 ( R_23de0_962e310, \46120 );
buf \U$labaj6122 ( R_23de2_9d16c30, \46127 );
buf \U$labaj6123 ( R_23de4_9d16e28, \46134 );
buf \U$labaj6124 ( R_23de8_9d170c8, \46141 );
buf \U$labaj6125 ( R_23dea_955f1c0, \46148 );
buf \U$labaj6126 ( R_23dec_96c87a8, \46155 );
buf \U$labaj6127 ( R_23dee_955f310, \46162 );
buf \U$labaj6128 ( R_23df0_9d1bee0, \46169 );
buf \U$labaj6129 ( R_23df2_955f3b8, \46176 );
buf \U$labaj6130 ( R_23df4_95a39b0, \46183 );
buf \U$labaj6131 ( R_23df6_96c8af0, \46190 );
buf \U$labaj6132 ( R_23df8_95a3b00, \46197 );
buf \U$labaj6133 ( R_23dfa_95a40e8, \46204 );
buf \U$labaj6134 ( R_23dfe_95a44d8, \46211 );
buf \U$labaj6135 ( R_23e00_9d1bf88, \46218 );
buf \U$labaj6136 ( R_23e02_95a4580, \46225 );
buf \U$labaj6137 ( R_23e04_95a4c10, \46232 );
buf \U$labaj6138 ( R_23e06_9d17218, \46239 );
buf \U$labaj6139 ( R_23e08_95a5348, \46246 );
buf \U$labaj6140 ( R_23e0a_962ec40, \46253 );
buf \U$labaj6141 ( R_23e0c_9d17608, \46260 );
buf \U$labaj6142 ( R_23e0e_95a57e0, \46267 );
buf \U$labaj6143 ( R_23e10_95a5930, \46274 );
buf \U$labaj6144 ( R_23e14_9d18910, \46281 );
buf \U$labaj6145 ( R_23e16_9d19630, \46288 );
buf \U$labaj6146 ( R_23e18_95a5c78, \46295 );
buf \U$labaj6147 ( R_23e1a_95a6260, \46302 );
buf \U$labaj6148 ( R_23e24_9d1c030, \46311 );
buf \U$labaj6149 ( R_23e3a_95a4628, \46318 );
buf \U$labaj6150 ( R_23e50_95a48c8, \46325 );
buf \U$labaj6151 ( R_23e66_95a4b68, \46332 );
buf \U$labaj6152 ( R_23e7c_95b1438, \46339 );
buf \U$labaj6153 ( R_23e92_9d19780, \46346 );
buf \U$labaj6154 ( R_23e9c_95a6d88, \46353 );
buf \U$labaj6155 ( R_23e9e_95b1780, \46360 );
buf \U$labaj6156 ( R_23ea0_95a7028, \46367 );
buf \U$labaj6157 ( R_23ea2_95a70d0, \46374 );
buf \U$labaj6158 ( R_23e26_95b1828, \46381 );
buf \U$labaj6159 ( R_23e28_95a7220, \46388 );
buf \U$labaj6160 ( R_23e2a_95b2bd8, \46395 );
buf \U$labaj6161 ( R_23e2c_95b3310, \46402 );
buf \U$labaj6162 ( R_23e2e_95818b0, \46409 );
buf \U$labaj6163 ( R_23e30_9582138, \46416 );
buf \U$labaj6164 ( R_23e32_9582288, \46423 );
buf \U$labaj6165 ( R_23e34_95a7760, \46430 );
buf \U$labaj6166 ( R_23e36_9582870, \46437 );
buf \U$labaj6167 ( R_23e38_95a78b0, \46444 );
buf \U$labaj6168 ( R_23e3c_9d1c0d8, \46451 );
buf \U$labaj6169 ( R_23e3e_9582a68, \46458 );
buf \U$labaj6170 ( R_23e40_9d1b118, \46465 );
buf \U$labaj6171 ( R_23e42_9582e58, \46472 );
buf \U$labaj6172 ( R_23e44_9582f00, \46479 );
buf \U$labaj6173 ( R_23e46_95830f8, \46486 );
buf \U$labaj6174 ( R_23e48_958cbd8, \46493 );
buf \U$labaj6175 ( R_23e4a_958cc80, \46500 );
buf \U$labaj6176 ( R_23e4c_95a7aa8, \46507 );
buf \U$labaj6177 ( R_23e4e_958f5d8, \46514 );
buf \U$labaj6178 ( R_23e52_958f920, \46521 );
buf \U$labaj6179 ( R_23e54_9590058, \46528 );
buf \U$labaj6180 ( R_23e56_95a7bf8, \46535 );
buf \U$labaj6181 ( R_23e58_95a7ca0, \46542 );
buf \U$labaj6182 ( R_23e5a_95901a8, \46549 );
buf \U$labaj6183 ( R_23e5c_959fdb8, \46556 );
buf \U$labaj6184 ( R_23e5e_95a0b80, \46563 );
buf \U$labaj6185 ( R_23e60_9d1c4c8, \46570 );
buf \U$labaj6186 ( R_23e62_9625b28, \46577 );
buf \U$labaj6187 ( R_23e64_96261b8, \46584 );
buf \U$labaj6188 ( R_23e68_9d1b268, \46591 );
buf \U$labaj6189 ( R_23e6a_9d1c570, \46598 );
buf \U$labaj6190 ( R_23e6c_95a7d48, \46605 );
buf \U$labaj6191 ( R_23e6e_9626458, \46612 );
buf \U$labaj6192 ( R_23e70_95a8090, \46619 );
buf \U$labaj6193 ( R_23e72_9628330, \46626 );
buf \U$labaj6194 ( R_23e74_9628480, \46633 );
buf \U$labaj6195 ( R_23e76_9628528, \46640 );
buf \U$labaj6196 ( R_23e78_95a8138, \46647 );
buf \U$labaj6197 ( R_23e7a_96285d0, \46654 );
buf \U$labaj6198 ( R_23e7e_9628720, \46661 );
buf \U$labaj6199 ( R_23e80_9628bb8, \46668 );
buf \U$labaj6200 ( R_23e82_962c198, \46675 );
buf \U$labaj6201 ( R_23e84_9d1c618, \46682 );
buf \U$labaj6202 ( R_23e86_95a8288, \46689 );
buf \U$labaj6203 ( R_23e88_9634238, \46696 );
buf \U$labaj6204 ( R_23e8a_9d1c6c0, \46703 );
buf \U$labaj6205 ( R_23e8c_96342e0, \46710 );
buf \U$labaj6206 ( R_23e8e_9634970, \46717 );
buf \U$labaj6207 ( R_23e90_9d1c8b8, \46724 );
buf \U$labaj6208 ( R_23e94_9639830, \46731 );
buf \U$labaj6209 ( R_23e96_9d159d0, \46738 );
buf \U$labaj6210 ( R_23e98_9d15e68, \46745 );
buf \U$labaj6211 ( R_23e9a_95a83d8, \46752 );
buf \U$labaj6212 ( R_23c64_96c9a08, \46760 );
buf \U$labaj6213 ( R_23c66_9d1b658, \46766 );
buf \U$labaj6214 ( R_23c68_96ca920, \46772 );
buf \U$labaj6215 ( R_23c6a_9d244c0, \46778 );
buf \U$labaj6216 ( R_23c6c_96cb4f0, \46784 );
buf \U$labaj6217 ( R_23c6e_9d1b700, \46790 );
buf \U$labaj6218 ( R_23c70_9d1ca08, \46796 );
buf \U$labaj6219 ( R_23c72_96cb640, \46802 );
buf \U$labaj6220 ( R_23c74_962f030, \46807 );
buf \U$labaj6221 ( R_23c76_9d1cc00, \46812 );
buf \U$labaj6222 ( R_23c78_9d1cd50, \46817 );
buf \U$labaj6223 ( R_23c7a_9d1cdf8, \46822 );
buf \U$labaj6224 ( R_23c7c_9d1b7a8, \46827 );
buf \U$labaj6225 ( R_23c7e_9d1cf48, \46832 );
buf \U$labaj6226 ( R_23c80_9d1d098, \46837 );
buf \U$labaj6227 ( R_23c82_9d1d1e8, \46842 );
buf \U$labaj6228 ( R_23c84_95a8528, \46847 );
buf \U$labaj6229 ( R_23c86_9d1b9a0, \46852 );
buf \U$labaj6230 ( R_23c88_95a8720, \46857 );
buf \U$labaj6231 ( R_23c8a_9d1be38, \46862 );
buf \U$labaj6232 ( R_23c8c_9d246b8, \46867 );
buf \U$labaj6233 ( R_23c8e_96cb838, \46872 );
buf \U$labaj6234 ( R_23c90_9d24760, \46877 );
buf \U$labaj6235 ( R_23c92_9d1c2d0, \46882 );
buf \U$labaj6236 ( R_23c94_9d1d3e0, \46887 );
buf \U$labaj6237 ( R_23c96_95a87c8, \46892 );
buf \U$labaj6238 ( R_23c98_9d19438, \46897 );
buf \U$labaj6239 ( R_23c9a_9d1c378, \46902 );
buf \U$labaj6240 ( R_23c9c_9d1c768, \46907 );
buf \U$labaj6241 ( R_23c9e_9d1d488, \46912 );
buf \U$labaj6242 ( R_23ca0_9d1c960, \46917 );
buf \U$labaj6243 ( R_23ca2_9d1e8e0, \46922 );
buf \U$labaj6244 ( R_23ebc_9667ae0, \46929 );
buf \U$labaj6245 ( R_23ebe_965f6f8, \46934 );
buf \U$labaj6246 ( R_23ec0_9667b88, \46939 );
buf \U$labaj6247 ( R_23ec2_96688a8, \46944 );
buf \U$labaj6248 ( R_23ec4_95ac230, \46949 );
buf \U$labaj6249 ( R_23ec6_95ac428, \46954 );
buf \U$labaj6250 ( R_23ec8_966a780, \46959 );
buf \U$labaj6251 ( R_23eca_966a8d0, \46964 );
buf \U$labaj6252 ( R_23eba_965f8f0, \46969 );
buf \U$labaj6253 ( R_23ecc_95ac620, \46974 );
buf \U$labaj6254 ( R_23ece_95ac770, \46979 );
buf \U$labaj6255 ( R_23ed0_966a978, \46984 );
buf \U$labaj6256 ( R_23ed2_966aa20, \46989 );
buf \U$labaj6257 ( R_23eb8_966aac8, \47145 );
buf \U$labaj6258 ( R_23eea_95b1588, \47148 );
buf \U$labaj6259 ( R_23eec_9d1e448, \47151 );
buf \U$labaj6260 ( R_23eee_9d1e790, \47154 );
buf \U$labaj6261 ( R_23a0c_95b1630, \47182 );
buf \U$labaj6262 ( R_23a22_95b1c18, \47191 );
buf \U$labaj6263 ( R_23a38_966acc0, \47200 );
buf \U$labaj6264 ( R_23a4e_95b1d68, \47209 );
buf \U$labaj6265 ( R_23a64_966ad68, \47218 );
buf \U$labaj6266 ( R_23a7a_95b2c80, \47227 );
buf \U$labaj6267 ( R_23a84_9661a68, \47236 );
buf \U$labaj6268 ( R_23a86_9d1d7d0, \47245 );
buf \U$labaj6269 ( R_23a88_966ae10, \47254 );
buf \U$labaj6270 ( R_23a8a_966b0b0, \47263 );
buf \U$labaj6271 ( R_23a0e_962f420, \47272 );
buf \U$labaj6272 ( R_23a10_966ba88, \47281 );
buf \U$labaj6273 ( R_23a12_95b2fc8, \47290 );
buf \U$labaj6274 ( R_23a14_9d1f6a8, \47299 );
buf \U$labaj6275 ( R_23a16_952daf8, \47308 );
buf \U$labaj6276 ( R_23a18_95b3268, \47317 );
buf \U$labaj6277 ( R_23a1a_9581220, \47326 );
buf \U$labaj6278 ( R_23a1c_9d1d878, \47335 );
buf \U$labaj6279 ( R_23a1e_9663160, \47344 );
buf \U$labaj6280 ( R_23a20_9d1e250, \47353 );
buf \U$labaj6281 ( R_23a24_9d1fb40, \47362 );
buf \U$labaj6282 ( R_23a26_95305a0, \47371 );
buf \U$labaj6283 ( R_23a28_95812c8, \47380 );
buf \U$labaj6284 ( R_23a2a_9530798, \47389 );
buf \U$labaj6285 ( R_23a2c_95816b8, \47398 );
buf \U$labaj6286 ( R_23a2e_9663550, \47407 );
buf \U$labaj6287 ( R_23a30_9531e90, \47416 );
buf \U$labaj6288 ( R_23a32_9531f38, \47425 );
buf \U$labaj6289 ( R_23a34_9532130, \47434 );
buf \U$labaj6290 ( R_23a36_9532280, \47443 );
buf \U$labaj6291 ( R_23a3a_9532328, \47452 );
buf \U$labaj6292 ( R_23a3c_9581760, \47461 );
buf \U$labaj6293 ( R_23a3e_9581f40, \47470 );
buf \U$labaj6294 ( R_23a40_95323d0, \47479 );
buf \U$labaj6295 ( R_23a42_9532868, \47488 );
buf \U$labaj6296 ( R_23a44_9582720, \47497 );
buf \U$labaj6297 ( R_23a46_9532b08, \47506 );
buf \U$labaj6298 ( R_23a48_9532c58, \47515 );
buf \U$labaj6299 ( R_23a4a_9582918, \47524 );
buf \U$labaj6300 ( R_23a4c_966a4e0, \47533 );
buf \U$labaj6301 ( R_23a50_9532e50, \47542 );
buf \U$labaj6302 ( R_23a52_9d24808, \47551 );
buf \U$labaj6303 ( R_23a54_9533390, \47560 );
buf \U$labaj6304 ( R_23a56_9d20668, \47569 );
buf \U$labaj6305 ( R_23a58_9582db0, \47578 );
buf \U$labaj6306 ( R_23a5a_9583050, \47587 );
buf \U$labaj6307 ( R_23a5c_9533978, \47596 );
buf \U$labaj6308 ( R_23a5e_9534158, \47605 );
buf \U$labaj6309 ( R_23a60_9d20710, \47614 );
buf \U$labaj6310 ( R_23a62_95349e0, \47623 );
buf \U$labaj6311 ( R_23a66_9537290, \47632 );
buf \U$labaj6312 ( R_23a68_9d1f750, \47641 );
buf \U$labaj6313 ( R_23a6a_966a6d8, \47650 );
buf \U$labaj6314 ( R_23a6c_966aeb8, \47659 );
buf \U$labaj6315 ( R_23a6e_966b158, \47668 );
buf \U$labaj6316 ( R_23a70_9537a70, \47677 );
buf \U$labaj6317 ( R_23a72_9539f30, \47686 );
buf \U$labaj6318 ( R_23a74_95831a0, \47695 );
buf \U$labaj6319 ( R_23a76_9537c68, \47704 );
buf \U$labaj6320 ( R_23a78_9d20a58, \47713 );
buf \U$labaj6321 ( R_23a7c_9537d10, \47722 );
buf \U$labaj6322 ( R_23a7e_9537e60, \47731 );
buf \U$labaj6323 ( R_23a80_9538250, \47740 );
buf \U$labaj6324 ( R_23a82_95382f8, \47749 );
buf \U$labaj6325 ( R_23a8c_9d21e08, \47760 );
buf \U$labaj6326 ( R_23aa2_9583440, \47767 );
buf \U$labaj6327 ( R_23ab8_9d1f8a0, \47774 );
buf \U$labaj6328 ( R_23ace_9d1ff30, \47781 );
buf \U$labaj6329 ( R_23ae4_9d23ce0, \47788 );
buf \U$labaj6330 ( R_23afa_95834e8, \47795 );
buf \U$labaj6331 ( R_23b04_9583590, \47802 );
buf \U$labaj6332 ( R_23b06_9d20860, \47809 );
buf \U$labaj6333 ( R_23b08_9d24958, \47816 );
buf \U$labaj6334 ( R_23b0a_9d24ca0, \47823 );
buf \U$labaj6335 ( R_23a8e_95836e0, \47830 );
buf \U$labaj6336 ( R_23a90_9583e18, \47837 );
buf \U$labaj6337 ( R_23a92_9d25288, \47844 );
buf \U$labaj6338 ( R_23a94_9d20908, \47851 );
buf \U$labaj6339 ( R_23a96_9d25330, \47858 );
buf \U$labaj6340 ( R_23a98_9d22348, \47865 );
buf \U$labaj6341 ( R_23a9a_9d253d8, \47872 );
buf \U$labaj6342 ( R_23a9c_9d233b0, \47879 );
buf \U$labaj6343 ( R_23a9e_9d25528, \47886 );
buf \U$labaj6344 ( R_23aa0_9d255d0, \47893 );
buf \U$labaj6345 ( R_23aa4_9d23500, \47900 );
buf \U$labaj6346 ( R_23aa6_9d25678, \47907 );
buf \U$labaj6347 ( R_23aa8_9d23a40, \47914 );
buf \U$labaj6348 ( R_23aaa_9d24610, \47921 );
buf \U$labaj6349 ( R_23aac_9d25880, \47928 );
buf \U$labaj6350 ( R_23aae_9d248b0, \47935 );
buf \U$labaj6351 ( R_23ab0_9d26258, \47942 );
buf \U$labaj6352 ( R_23ab2_9584898, \47949 );
buf \U$labaj6353 ( R_23ab4_9d24a00, \47956 );
buf \U$labaj6354 ( R_23ab6_9d26450, \47963 );
buf \U$labaj6355 ( R_23aba_9d26648, \47970 );
buf \U$labaj6356 ( R_23abc_9d26e28, \47977 );
buf \U$labaj6357 ( R_23abe_9d270c8, \47984 );
buf \U$labaj6358 ( R_23ac0_9584c88, \47991 );
buf \U$labaj6359 ( R_23ac2_9d24aa8, \47998 );
buf \U$labaj6360 ( R_23ac4_9d24d48, \48005 );
buf \U$labaj6361 ( R_23ac6_9585270, \48012 );
buf \U$labaj6362 ( R_23ac8_9585708, \48019 );
buf \U$labaj6363 ( R_23aca_9d27bf0, \48026 );
buf \U$labaj6364 ( R_23acc_9d28910, \48033 );
buf \U$labaj6365 ( R_23ad0_9d29198, \48040 );
buf \U$labaj6366 ( R_23ad2_9d29630, \48047 );
buf \U$labaj6367 ( R_23ad4_9d24fe8, \48054 );
buf \U$labaj6368 ( R_23ad6_95857b0, \48061 );
buf \U$labaj6369 ( R_23ad8_9d2a0b0, \48068 );
buf \U$labaj6370 ( R_23ada_9585900, \48075 );
buf \U$labaj6371 ( R_23adc_9d2a200, \48082 );
buf \U$labaj6372 ( R_23ade_9d2a3f8, \48089 );
buf \U$labaj6373 ( R_23ae0_9d2a7e8, \48096 );
buf \U$labaj6374 ( R_23ae2_9d25138, \48103 );
buf \U$labaj6375 ( R_23ae6_9d2ad28, \48110 );
buf \U$labaj6376 ( R_23ae8_95860e0, \48117 );
buf \U$labaj6377 ( R_23aea_9d25480, \48124 );
buf \U$labaj6378 ( R_23aec_9d25928, \48131 );
buf \U$labaj6379 ( R_23aee_9d25bc8, \48138 );
buf \U$labaj6380 ( R_23af0_95864d0, \48145 );
buf \U$labaj6381 ( R_23af2_9d25e68, \48152 );
buf \U$labaj6382 ( R_23af4_95866c8, \48159 );
buf \U$labaj6383 ( R_23af6_9586770, \48166 );
buf \U$labaj6384 ( R_23af8_9587688, \48173 );
buf \U$labaj6385 ( R_23afc_9d26ed0, \48180 );
buf \U$labaj6386 ( R_23afe_9587730, \48187 );
buf \U$labaj6387 ( R_23b00_9d27aa0, \48194 );
buf \U$labaj6388 ( R_23b02_9d2add0, \48201 );
buf \U$labaj6389 ( R_23b0c_95877d8, \48210 );
buf \U$labaj6390 ( R_23b22_95386e8, \48217 );
buf \U$labaj6391 ( R_23b38_95388e0, \48224 );
buf \U$labaj6392 ( R_23b4e_9588108, \48231 );
buf \U$labaj6393 ( R_23b64_9538ad8, \48238 );
buf \U$labaj6394 ( R_23b7a_9d2b118, \48245 );
buf \U$labaj6395 ( R_23b84_95881b0, \48252 );
buf \U$labaj6396 ( R_23b86_95899f8, \48259 );
buf \U$labaj6397 ( R_23b88_9589aa0, \48266 );
buf \U$labaj6398 ( R_23b8a_9d2b460, \48273 );
buf \U$labaj6399 ( R_23b0e_958d268, \48280 );
buf \U$labaj6400 ( R_23b10_95390c0, \48287 );
buf \U$labaj6401 ( R_23b12_9539168, \48294 );
buf \U$labaj6402 ( R_23b14_95394b0, \48301 );
buf \U$labaj6403 ( R_23b16_95399f0, \48308 );
buf \U$labaj6404 ( R_23b18_9539c90, \48315 );
buf \U$labaj6405 ( R_23b1a_953ba18, \48322 );
buf \U$labaj6406 ( R_23b1c_953bac0, \48329 );
buf \U$labaj6407 ( R_23b1e_958d460, \48336 );
buf \U$labaj6408 ( R_23b20_9d2b508, \48343 );
buf \U$labaj6409 ( R_23b24_953bf58, \48350 );
buf \U$labaj6410 ( R_23b26_953c0a8, \48357 );
buf \U$labaj6411 ( R_23b28_953c1f8, \48364 );
buf \U$labaj6412 ( R_23b2a_953c540, \48371 );
buf \U$labaj6413 ( R_23b2c_9d2b5b0, \48378 );
buf \U$labaj6414 ( R_23b2e_953c888, \48385 );
buf \U$labaj6415 ( R_23b30_953cdc8, \48392 );
buf \U$labaj6416 ( R_23b32_958da48, \48399 );
buf \U$labaj6417 ( R_23b34_9d2b700, \48406 );
buf \U$labaj6418 ( R_23b36_953cf18, \48413 );
buf \U$labaj6419 ( R_23b3a_958de38, \48420 );
buf \U$labaj6420 ( R_23b3c_958e180, \48427 );
buf \U$labaj6421 ( R_23b3e_96ddca8, \48434 );
buf \U$labaj6422 ( R_23b40_96dddf8, \48441 );
buf \U$labaj6423 ( R_23b42_958e570, \48448 );
buf \U$labaj6424 ( R_23b44_958e810, \48455 );
buf \U$labaj6425 ( R_23b46_96de098, \48462 );
buf \U$labaj6426 ( R_23b48_9d285c8, \48469 );
buf \U$labaj6427 ( R_23b4a_96de3e0, \48476 );
buf \U$labaj6428 ( R_23b4c_9d28b08, \48483 );
buf \U$labaj6429 ( R_23b50_96de530, \48490 );
buf \U$labaj6430 ( R_23b52_958ef48, \48497 );
buf \U$labaj6431 ( R_23b54_9d24b50, \48504 );
buf \U$labaj6432 ( R_23b56_9d25d18, \48511 );
buf \U$labaj6433 ( R_23b58_958ff08, \48518 );
buf \U$labaj6434 ( R_23b5a_96e6c60, \48525 );
buf \U$labaj6435 ( R_23b5c_96e8160, \48532 );
buf \U$labaj6436 ( R_23b5e_96ebc70, \48539 );
buf \U$labaj6437 ( R_23b60_95903a0, \48546 );
buf \U$labaj6438 ( R_23b62_95906e8, \48553 );
buf \U$labaj6439 ( R_23b66_96ebdc0, \48560 );
buf \U$labaj6440 ( R_23b68_95efb90, \48567 );
buf \U$labaj6441 ( R_23b6a_9596d58, \48574 );
buf \U$labaj6442 ( R_23b6c_9d2b7a8, \48581 );
buf \U$labaj6443 ( R_23b6e_9598c30, \48588 );
buf \U$labaj6444 ( R_23b70_95f0220, \48595 );
buf \U$labaj6445 ( R_23b72_9598cd8, \48602 );
buf \U$labaj6446 ( R_23b74_95f1918, \48609 );
buf \U$labaj6447 ( R_23b76_9599170, \48616 );
buf \U$labaj6448 ( R_23b78_9d28bb0, \48623 );
buf \U$labaj6449 ( R_23b7c_95f37f0, \48630 );
buf \U$labaj6450 ( R_23b7e_95f41c8, \48637 );
buf \U$labaj6451 ( R_23b80_95f4318, \48644 );
buf \U$labaj6452 ( R_23b82_95992c0, \48651 );
buf \U$labaj6453 ( R_23b8c_9599608, \48660 );
buf \U$labaj6454 ( R_23ba2_9599758, \48667 );
buf \U$labaj6455 ( R_23bb8_9599800, \48674 );
buf \U$labaj6456 ( R_23bce_9599950, \48681 );
buf \U$labaj6457 ( R_23be4_962f570, \48688 );
buf \U$labaj6458 ( R_23bfa_9599b48, \48695 );
buf \U$labaj6459 ( R_23c04_959a088, \48702 );
buf \U$labaj6460 ( R_23c06_959a130, \48709 );
buf \U$labaj6461 ( R_23c08_959a1d8, \48716 );
buf \U$labaj6462 ( R_23c0a_962f618, \48723 );
buf \U$labaj6463 ( R_23b8e_959a5c8, \48730 );
buf \U$labaj6464 ( R_23b90_959a9b8, \48737 );
buf \U$labaj6465 ( R_23b92_959ac58, \48744 );
buf \U$labaj6466 ( R_23b94_959aef8, \48751 );
buf \U$labaj6467 ( R_23b96_962f8b8, \48758 );
buf \U$labaj6468 ( R_23b98_959afa0, \48765 );
buf \U$labaj6469 ( R_23b9a_959b048, \48772 );
buf \U$labaj6470 ( R_23b9c_959b0f0, \48779 );
buf \U$labaj6471 ( R_23b9e_959b198, \48786 );
buf \U$labaj6472 ( R_23ba0_959b240, \48793 );
buf \U$labaj6473 ( R_23ba4_959b6d8, \48800 );
buf \U$labaj6474 ( R_23ba6_959b828, \48807 );
buf \U$labaj6475 ( R_23ba8_959b8d0, \48814 );
buf \U$labaj6476 ( R_23baa_959ba20, \48821 );
buf \U$labaj6477 ( R_23bac_9d28da8, \48828 );
buf \U$labaj6478 ( R_23bae_959bac8, \48835 );
buf \U$labaj6479 ( R_23bb0_959d268, \48842 );
buf \U$labaj6480 ( R_23bb2_959d508, \48849 );
buf \U$labaj6481 ( R_23bb4_959dce8, \48856 );
buf \U$labaj6482 ( R_23bb6_959e420, \48863 );
buf \U$labaj6483 ( R_23bba_9d28fa0, \48870 );
buf \U$labaj6484 ( R_23bbc_962f960, \48877 );
buf \U$labaj6485 ( R_23bbe_9d298d0, \48884 );
buf \U$labaj6486 ( R_23bc0_959e618, \48891 );
buf \U$labaj6487 ( R_23bc2_959eea0, \48898 );
buf \U$labaj6488 ( R_23bc4_959f098, \48905 );
buf \U$labaj6489 ( R_23bc6_9d29978, \48912 );
buf \U$labaj6490 ( R_23bc8_9d25dc0, \48919 );
buf \U$labaj6491 ( R_23bca_959f9c8, \48926 );
buf \U$labaj6492 ( R_23bcc_9d29a20, \48933 );
buf \U$labaj6493 ( R_23bd0_95a0e20, \48940 );
buf \U$labaj6494 ( R_23bd2_9d29b70, \48947 );
buf \U$labaj6495 ( R_23bd4_962fb58, \48954 );
buf \U$labaj6496 ( R_23bd6_95a0f70, \48961 );
buf \U$labaj6497 ( R_23bd8_9d29c18, \48968 );
buf \U$labaj6498 ( R_23bda_9619ae0, \48975 );
buf \U$labaj6499 ( R_23bdc_9619b88, \48982 );
buf \U$labaj6500 ( R_23bde_9619d80, \48989 );
buf \U$labaj6501 ( R_23be0_9619e28, \48996 );
buf \U$labaj6502 ( R_23be2_961a020, \49003 );
buf \U$labaj6503 ( R_23be6_961a0c8, \49010 );
buf \U$labaj6504 ( R_23be8_961a218, \49017 );
buf \U$labaj6505 ( R_23bea_961a4b8, \49024 );
buf \U$labaj6506 ( R_23bec_961a800, \49031 );
buf \U$labaj6507 ( R_23bee_961a8a8, \49038 );
buf \U$labaj6508 ( R_23bf0_961a950, \49045 );
buf \U$labaj6509 ( R_23bf2_961ad40, \49052 );
buf \U$labaj6510 ( R_23bf4_961ade8, \49059 );
buf \U$labaj6511 ( R_23bf6_961ae90, \49066 );
buf \U$labaj6512 ( R_23bf8_961af38, \49073 );
buf \U$labaj6513 ( R_23bfc_9d26060, \49080 );
buf \U$labaj6514 ( R_23bfe_961b088, \49087 );
buf \U$labaj6515 ( R_23c00_9d29d68, \49094 );
buf \U$labaj6516 ( R_23c02_961b1d8, \49101 );
buf \U$labaj6517 ( R_239cc_95f4af8, \49109 );
buf \U$labaj6518 ( R_239ce_962fd50, \49115 );
buf \U$labaj6519 ( R_239d0_9558e00, \49121 );
buf \U$labaj6520 ( R_239d2_9d261b0, \49127 );
buf \U$labaj6521 ( R_239d4_95f52d8, \49133 );
buf \U$labaj6522 ( R_239d6_9558ea8, \49139 );
buf \U$labaj6523 ( R_239d8_961b670, \49145 );
buf \U$labaj6524 ( R_239da_95f5620, \49151 );
buf \U$labaj6525 ( R_239dc_961b910, \49156 );
buf \U$labaj6526 ( R_239de_9d2b850, \49161 );
buf \U$labaj6527 ( R_239e0_9d2b9a0, \49166 );
buf \U$labaj6528 ( R_239e2_9d29e10, \49171 );
buf \U$labaj6529 ( R_239e4_9d2a158, \49176 );
buf \U$labaj6530 ( R_239e6_961bb08, \49181 );
buf \U$labaj6531 ( R_239e8_961c978, \49186 );
buf \U$labaj6532 ( R_239ea_961cd68, \49191 );
buf \U$labaj6533 ( R_239ec_9d2baf0, \49196 );
buf \U$labaj6534 ( R_239ee_95f5968, \49201 );
buf \U$labaj6535 ( R_239f0_95f5ab8, \49206 );
buf \U$labaj6536 ( R_239f2_9d2a2a8, \49211 );
buf \U$labaj6537 ( R_239f4_961ce10, \49216 );
buf \U$labaj6538 ( R_239f6_9634e08, \49221 );
buf \U$labaj6539 ( R_239f8_9d2bb98, \49226 );
buf \U$labaj6540 ( R_239fa_9d2bd90, \49231 );
buf \U$labaj6541 ( R_239fc_962fdf8, \49236 );
buf \U$labaj6542 ( R_239fe_962fea0, \49241 );
buf \U$labaj6543 ( R_23a00_961d200, \49246 );
buf \U$labaj6544 ( R_23a02_961d5f0, \49251 );
buf \U$labaj6545 ( R_23a04_961d698, \49256 );
buf \U$labaj6546 ( R_23a06_962fff0, \49261 );
buf \U$labaj6547 ( R_23a08_961d740, \49266 );
buf \U$labaj6548 ( R_23a0a_961d938, \49271 );
buf \U$labaj6549 ( R_23c24_9d2a698, \49278 );
buf \U$labaj6550 ( R_23c26_9d2c420, \49283 );
buf \U$labaj6551 ( R_23c28_962ac98, \49288 );
buf \U$labaj6552 ( R_23c2a_9d2c4c8, \49293 );
buf \U$labaj6553 ( R_23c2c_9d2c570, \49298 );
buf \U$labaj6554 ( R_23c2e_95f63e8, \49303 );
buf \U$labaj6555 ( R_23c30_9d2a890, \49308 );
buf \U$labaj6556 ( R_23c32_962ad40, \49313 );
buf \U$labaj6557 ( R_23c22_9d2aa88, \49318 );
buf \U$labaj6558 ( R_23c34_9d2c810, \49323 );
buf \U$labaj6559 ( R_23c36_9d2ab30, \49328 );
buf \U$labaj6560 ( R_23c38_9d2c8b8, \49333 );
buf \U$labaj6561 ( R_23c3a_9d2cab0, \49338 );
buf \U$labaj6562 ( R_23c20_9635e70, \49494 );
buf \U$labaj6563 ( R_23c52_962b868, \49497 );
buf \U$labaj6564 ( R_23c54_9d2af20, \49500 );
buf \U$labaj6565 ( R_23c56_9d2b310, \49503 );
buf \U$labaj6566 ( R_23774_9630098, \49530 );
buf \U$labaj6567 ( R_2378a_962b9b8, \49539 );
buf \U$labaj6568 ( R_237a0_9d2cd50, \49548 );
buf \U$labaj6569 ( R_237b6_962bb08, \49557 );
buf \U$labaj6570 ( R_237cc_9d2cff0, \49566 );
buf \U$labaj6571 ( R_237e2_9d2d098, \49575 );
buf \U$labaj6572 ( R_237ec_9d2d140, \49584 );
buf \U$labaj6573 ( R_237ee_9d2d290, \49593 );
buf \U$labaj6574 ( R_237f0_962c240, \49602 );
buf \U$labaj6575 ( R_237f2_9559688, \49611 );
buf \U$labaj6576 ( R_23776_96301e8, \49620 );
buf \U$labaj6577 ( R_23778_9d2d7d0, \49629 );
buf \U$labaj6578 ( R_2377a_962c2e8, \49638 );
buf \U$labaj6579 ( R_2377c_9d2d878, \49647 );
buf \U$labaj6580 ( R_2377e_962ce10, \49656 );
buf \U$labaj6581 ( R_23780_9d2d920, \49665 );
buf \U$labaj6582 ( R_23782_962d938, \49674 );
buf \U$labaj6583 ( R_23784_962e5b0, \49683 );
buf \U$labaj6584 ( R_23786_9d2d9c8, \49692 );
buf \U$labaj6585 ( R_23788_9d2dc68, \49701 );
buf \U$labaj6586 ( R_2378c_9d2dd10, \49710 );
buf \U$labaj6587 ( R_2378e_9d2ddb8, \49719 );
buf \U$labaj6588 ( R_23790_9d2e100, \49728 );
buf \U$labaj6589 ( R_23792_9d2e1a8, \49737 );
buf \U$labaj6590 ( R_23794_9d2f0c0, \49746 );
buf \U$labaj6591 ( R_23796_9630290, \49755 );
buf \U$labaj6592 ( R_23798_96303e0, \49764 );
buf \U$labaj6593 ( R_2379a_9d2f210, \49773 );
buf \U$labaj6594 ( R_2379c_9d2f7f8, \49782 );
buf \U$labaj6595 ( R_2379e_9630728, \49791 );
buf \U$labaj6596 ( R_237a2_96307d0, \49800 );
buf \U$labaj6597 ( R_237a4_9d2fb40, \49809 );
buf \U$labaj6598 ( R_237a6_9d301d0, \49818 );
buf \U$labaj6599 ( R_237a8_9559bc8, \49827 );
buf \U$labaj6600 ( R_237aa_9630140, \49836 );
buf \U$labaj6601 ( R_237ac_96312f8, \49845 );
buf \U$labaj6602 ( R_237ae_9d30710, \49854 );
buf \U$labaj6603 ( R_237b0_9630b18, \49863 );
buf \U$labaj6604 ( R_237b2_9630c68, \49872 );
buf \U$labaj6605 ( R_237b4_9d309b0, \49881 );
buf \U$labaj6606 ( R_237b8_9630d10, \49890 );
buf \U$labaj6607 ( R_237ba_9630fb0, \49899 );
buf \U$labaj6608 ( R_237bc_9631100, \49908 );
buf \U$labaj6609 ( R_237be_9d30a58, \49917 );
buf \U$labaj6610 ( R_237c0_9d30da0, \49926 );
buf \U$labaj6611 ( R_237c2_96311a8, \49935 );
buf \U$labaj6612 ( R_237c4_96313a0, \49944 );
buf \U$labaj6613 ( R_237c6_96318e0, \49953 );
buf \U$labaj6614 ( R_237c8_9631a30, \49962 );
buf \U$labaj6615 ( R_237ca_9d30e48, \49971 );
buf \U$labaj6616 ( R_237ce_9d31190, \49980 );
buf \U$labaj6617 ( R_237d0_9631b80, \49989 );
buf \U$labaj6618 ( R_237d2_9d31f58, \49998 );
buf \U$labaj6619 ( R_237d4_9631448, \50007 );
buf \U$labaj6620 ( R_237d6_9631790, \50016 );
buf \U$labaj6621 ( R_237d8_9d323f0, \50025 );
buf \U$labaj6622 ( R_237da_9631ad8, \50034 );
buf \U$labaj6623 ( R_237dc_9d32540, \50043 );
buf \U$labaj6624 ( R_237de_9632018, \50052 );
buf \U$labaj6625 ( R_237e0_9631cd0, \50061 );
buf \U$labaj6626 ( R_237e4_9632210, \50070 );
buf \U$labaj6627 ( R_237e6_9d32690, \50079 );
buf \U$labaj6628 ( R_237e8_96322b8, \50088 );
buf \U$labaj6629 ( R_237ea_9d32888, \50097 );
buf \U$labaj6630 ( R_237f4_9631e20, \50108 );
buf \U$labaj6631 ( R_2380a_9d329d8, \50115 );
buf \U$labaj6632 ( R_23820_9d32a80, \50122 );
buf \U$labaj6633 ( R_23836_9d32f18, \50129 );
buf \U$labaj6634 ( R_2384c_9d2b3b8, \50136 );
buf \U$labaj6635 ( R_23862_9631ec8, \50143 );
buf \U$labaj6636 ( R_2386c_9632360, \50150 );
buf \U$labaj6637 ( R_2386e_9632a98, \50157 );
buf \U$labaj6638 ( R_23870_9d32fc0, \50164 );
buf \U$labaj6639 ( R_23872_9632408, \50171 );
buf \U$labaj6640 ( R_237f6_9632600, \50178 );
buf \U$labaj6641 ( R_237f8_9d33500, \50185 );
buf \U$labaj6642 ( R_237fa_96326a8, \50192 );
buf \U$labaj6643 ( R_237fc_9d33650, \50199 );
buf \U$labaj6644 ( R_237fe_9d336f8, \50206 );
buf \U$labaj6645 ( R_23800_9d33a40, \50213 );
buf \U$labaj6646 ( R_23802_9632750, \50220 );
buf \U$labaj6647 ( R_23804_96328a0, \50227 );
buf \U$labaj6648 ( R_23806_9d340d0, \50234 );
buf \U$labaj6649 ( R_23808_9632948, \50241 );
buf \U$labaj6650 ( R_2380c_9d2b658, \50248 );
buf \U$labaj6651 ( R_2380e_9d34418, \50255 );
buf \U$labaj6652 ( R_23810_9d34760, \50262 );
buf \U$labaj6653 ( R_23812_9d34fe8, \50269 );
buf \U$labaj6654 ( R_23814_9632de0, \50276 );
buf \U$labaj6655 ( R_23816_9632e88, \50283 );
buf \U$labaj6656 ( R_23818_9d35720, \50290 );
buf \U$labaj6657 ( R_2381a_9d2bc40, \50297 );
buf \U$labaj6658 ( R_2381c_b805670, \50304 );
buf \U$labaj6659 ( R_2381e_b805868, \50311 );
buf \U$labaj6660 ( R_23822_9633080, \50318 );
buf \U$labaj6661 ( R_23824_b8060f0, \50325 );
buf \U$labaj6662 ( R_23826_9633128, \50332 );
buf \U$labaj6663 ( R_23828_9633b00, \50339 );
buf \U$labaj6664 ( R_2382a_9632b40, \50346 );
buf \U$labaj6665 ( R_2382c_9634190, \50353 );
buf \U$labaj6666 ( R_2382e_9638720, \50360 );
buf \U$labaj6667 ( R_23830_9d2c180, \50367 );
buf \U$labaj6668 ( R_23832_96389c0, \50374 );
buf \U$labaj6669 ( R_23834_9638a68, \50381 );
buf \U$labaj6670 ( R_23838_9d15880, \50388 );
buf \U$labaj6671 ( R_2383a_b806198, \50395 );
buf \U$labaj6672 ( R_2383c_9d2c768, \50402 );
buf \U$labaj6673 ( R_2383e_9d16a38, \50409 );
buf \U$labaj6674 ( R_23840_9d2ca08, \50416 );
buf \U$labaj6675 ( R_23842_b806240, \50423 );
buf \U$labaj6676 ( R_23844_9d17170, \50430 );
buf \U$labaj6677 ( R_23846_9d17c98, \50437 );
buf \U$labaj6678 ( R_23848_b8062e8, \50444 );
buf \U$labaj6679 ( R_2384a_b806390, \50451 );
buf \U$labaj6680 ( R_2384e_9d2cca8, \50458 );
buf \U$labaj6681 ( R_23850_9d17fe0, \50465 );
buf \U$labaj6682 ( R_23852_9d18328, \50472 );
buf \U$labaj6683 ( R_23854_9d2d1e8, \50479 );
buf \U$labaj6684 ( R_23856_9d1fd38, \50486 );
buf \U$labaj6685 ( R_23858_b8064e0, \50493 );
buf \U$labaj6686 ( R_2385a_9d2d3e0, \50500 );
buf \U$labaj6687 ( R_2385c_9d220a8, \50507 );
buf \U$labaj6688 ( R_2385e_9535d90, \50514 );
buf \U$labaj6689 ( R_23860_b806588, \50521 );
buf \U$labaj6690 ( R_23864_9d25720, \50528 );
buf \U$labaj6691 ( R_23866_b8066d8, \50535 );
buf \U$labaj6692 ( R_23868_b806780, \50542 );
buf \U$labaj6693 ( R_2386a_9d2d530, \50549 );
buf \U$labaj6694 ( R_23874_95f7840, \50558 );
buf \U$labaj6695 ( R_2388a_95f7e28, \50565 );
buf \U$labaj6696 ( R_238a0_9d28e50, \50572 );
buf \U$labaj6697 ( R_238b6_95f8170, \50579 );
buf \U$labaj6698 ( R_238cc_95fcd90, \50586 );
buf \U$labaj6699 ( R_238e2_95fda08, \50593 );
buf \U$labaj6700 ( R_238ec_95fdb58, \50600 );
buf \U$labaj6701 ( R_238ee_95fdca8, \50607 );
buf \U$labaj6702 ( R_238f0_95fdd50, \50614 );
buf \U$labaj6703 ( R_238f2_9d2d728, \50621 );
buf \U$labaj6704 ( R_23876_95ff6e8, \50628 );
buf \U$labaj6705 ( R_23878_9535e38, \50635 );
buf \U$labaj6706 ( R_2387a_9633668, \50642 );
buf \U$labaj6707 ( R_2387c_9f4ddd0, \50649 );
buf \U$labaj6708 ( R_2387e_9f51b80, \50656 );
buf \U$labaj6709 ( R_23880_9f51e20, \50663 );
buf \U$labaj6710 ( R_23882_9d29ac8, \50670 );
buf \U$labaj6711 ( R_23884_9f53278, \50677 );
buf \U$labaj6712 ( R_23886_9f53320, \50684 );
buf \U$labaj6713 ( R_23888_9f54580, \50691 );
buf \U$labaj6714 ( R_2388c_9f54778, \50698 );
buf \U$labaj6715 ( R_2388e_9d2dbc0, \50705 );
buf \U$labaj6716 ( R_23890_9d2e250, \50712 );
buf \U$labaj6717 ( R_23892_9f548c8, \50719 );
buf \U$labaj6718 ( R_23894_9f54970, \50726 );
buf \U$labaj6719 ( R_23896_9f54c10, \50733 );
buf \U$labaj6720 ( R_23898_9f55348, \50740 );
buf \U$labaj6721 ( R_2389a_9f55498, \50747 );
buf \U$labaj6722 ( R_2389c_9d2a740, \50754 );
buf \U$labaj6723 ( R_2389e_9d2e3a0, \50761 );
buf \U$labaj6724 ( R_238a2_9d2b070, \50768 );
buf \U$labaj6725 ( R_238a4_9633710, \50775 );
buf \U$labaj6726 ( R_238a6_9f55b28, \50782 );
buf \U$labaj6727 ( R_238a8_9f56260, \50789 );
buf \U$labaj6728 ( R_238aa_9f56500, \50796 );
buf \U$labaj6729 ( R_238ac_9f5baf8, \50803 );
buf \U$labaj6730 ( R_238ae_9ee9d78, \50810 );
buf \U$labaj6731 ( R_238b0_9d2ba48, \50817 );
buf \U$labaj6732 ( R_238b2_9d2bce8, \50824 );
buf \U$labaj6733 ( R_238b4_9eea0c0, \50831 );
buf \U$labaj6734 ( R_238b8_9eeb518, \50838 );
buf \U$labaj6735 ( R_238ba_9eedf18, \50845 );
buf \U$labaj6736 ( R_238bc_9eee6f8, \50852 );
buf \U$labaj6737 ( R_238be_9ef2010, \50859 );
buf \U$labaj6738 ( R_238c0_9537530, \50866 );
buf \U$labaj6739 ( R_238c2_9ef2208, \50873 );
buf \U$labaj6740 ( R_238c4_9ef3660, \50880 );
buf \U$labaj6741 ( R_238c6_9ef3858, \50887 );
buf \U$labaj6742 ( R_238c8_9633860, \50894 );
buf \U$labaj6743 ( R_238ca_9ef3a50, \50901 );
buf \U$labaj6744 ( R_238ce_9ef3af8, \50908 );
buf \U$labaj6745 ( R_238d0_9ef3ba0, \50915 );
buf \U$labaj6746 ( R_238d2_9ef3c48, \50922 );
buf \U$labaj6747 ( R_238d4_9ef4620, \50929 );
buf \U$labaj6748 ( R_238d6_9d2c2d0, \50936 );
buf \U$labaj6749 ( R_238d8_9ef4770, \50943 );
buf \U$labaj6750 ( R_238da_9d2cb58, \50950 );
buf \U$labaj6751 ( R_238dc_9ef4ab8, \50957 );
buf \U$labaj6752 ( R_238de_9ef4c08, \50964 );
buf \U$labaj6753 ( R_238e0_9ef4ff8, \50971 );
buf \U$labaj6754 ( R_238e4_9ef5148, \50978 );
buf \U$labaj6755 ( R_238e6_9ef51f0, \50985 );
buf \U$labaj6756 ( R_238e8_9d2cf48, \50992 );
buf \U$labaj6757 ( R_238ea_9ef53e8, \50999 );
buf \U$labaj6758 ( R_238f4_9d2e4f0, \51008 );
buf \U$labaj6759 ( R_2390a_96339b0, \51015 );
buf \U$labaj6760 ( R_23920_9633c50, \51022 );
buf \U$labaj6761 ( R_23936_9d266f0, \51029 );
buf \U$labaj6762 ( R_2394c_9d2e838, \51036 );
buf \U$labaj6763 ( R_23962_9d2ecd0, \51043 );
buf \U$labaj6764 ( R_2396c_9d2ed78, \51050 );
buf \U$labaj6765 ( R_2396e_9d2f018, \51057 );
buf \U$labaj6766 ( R_23970_9d2f168, \51064 );
buf \U$labaj6767 ( R_23972_b8068d0, \51071 );
buf \U$labaj6768 ( R_238f6_9d2f2b8, \51078 );
buf \U$labaj6769 ( R_238f8_9d2f9f0, \51085 );
buf \U$labaj6770 ( R_238fa_9d2fde0, \51092 );
buf \U$labaj6771 ( R_238fc_9633f98, \51099 );
buf \U$labaj6772 ( R_238fe_b806a20, \51106 );
buf \U$labaj6773 ( R_23900_96340e8, \51113 );
buf \U$labaj6774 ( R_23902_9d30320, \51120 );
buf \U$labaj6775 ( R_23904_9634580, \51127 );
buf \U$labaj6776 ( R_23906_9d305c0, \51134 );
buf \U$labaj6777 ( R_23908_9634b68, \51141 );
buf \U$labaj6778 ( R_2390c_9d30ba8, \51148 );
buf \U$labaj6779 ( R_2390e_9d30c50, \51155 );
buf \U$labaj6780 ( R_23910_b806ac8, \51162 );
buf \U$labaj6781 ( R_23912_9d32000, \51169 );
buf \U$labaj6782 ( R_23914_b806b70, \51176 );
buf \U$labaj6783 ( R_23916_9d320a8, \51183 );
buf \U$labaj6784 ( R_23918_9634c10, \51190 );
buf \U$labaj6785 ( R_2391a_9d32150, \51197 );
buf \U$labaj6786 ( R_2391c_9634cb8, \51204 );
buf \U$labaj6787 ( R_2391e_9d32498, \51211 );
buf \U$labaj6788 ( R_23922_9d32738, \51218 );
buf \U$labaj6789 ( R_23924_9d327e0, \51225 );
buf \U$labaj6790 ( R_23926_9d32b28, \51232 );
buf \U$labaj6791 ( R_23928_9d32bd0, \51239 );
buf \U$labaj6792 ( R_2392a_9635348, \51246 );
buf \U$labaj6793 ( R_2392c_9635690, \51253 );
buf \U$labaj6794 ( R_2392e_9d32c78, \51260 );
buf \U$labaj6795 ( R_23930_9d32d20, \51267 );
buf \U$labaj6796 ( R_23932_9635a80, \51274 );
buf \U$labaj6797 ( R_23934_9d32dc8, \51281 );
buf \U$labaj6798 ( R_23938_9d331b8, \51288 );
buf \U$labaj6799 ( R_2393a_9d2d488, \51295 );
buf \U$labaj6800 ( R_2393c_9d333b0, \51302 );
buf \U$labaj6801 ( R_2393e_9d335a8, \51309 );
buf \U$labaj6802 ( R_23940_9d337a0, \51316 );
buf \U$labaj6803 ( R_23942_9635b28, \51323 );
buf \U$labaj6804 ( R_23944_9d2d5d8, \51330 );
buf \U$labaj6805 ( R_23946_9d338f0, \51337 );
buf \U$labaj6806 ( R_23948_9635bd0, \51344 );
buf \U$labaj6807 ( R_2394a_9d33998, \51351 );
buf \U$labaj6808 ( R_2394e_9d33ae8, \51358 );
buf \U$labaj6809 ( R_23950_9d33b90, \51365 );
buf \U$labaj6810 ( R_23952_9636110, \51372 );
buf \U$labaj6811 ( R_23954_9d33ce0, \51379 );
buf \U$labaj6812 ( R_23956_b806c18, \51386 );
buf \U$labaj6813 ( R_23958_9d33ed8, \51393 );
buf \U$labaj6814 ( R_2395a_9d33f80, \51400 );
buf \U$labaj6815 ( R_2395c_9636308, \51407 );
buf \U$labaj6816 ( R_2395e_b806cc0, \51414 );
buf \U$labaj6817 ( R_23960_9d34028, \51421 );
buf \U$labaj6818 ( R_23964_9d34178, \51428 );
buf \U$labaj6819 ( R_23966_9d2db18, \51435 );
buf \U$labaj6820 ( R_23968_96365a8, \51442 );
buf \U$labaj6821 ( R_2396a_9636848, \51449 );
buf \U$labaj6822 ( R_23734_96368f0, \51457 );
buf \U$labaj6823 ( R_23736_9636998, \51463 );
buf \U$labaj6824 ( R_23738_9636a40, \51469 );
buf \U$labaj6825 ( R_2373a_b7dc0c0, \51475 );
buf \U$labaj6826 ( R_2373c_9636b90, \51481 );
buf \U$labaj6827 ( R_2373e_9636c38, \51487 );
buf \U$labaj6828 ( R_23740_b7dc168, \51493 );
buf \U$labaj6829 ( R_23742_b806d68, \51499 );
buf \U$labaj6830 ( R_23744_b806e10, \51504 );
buf \U$labaj6831 ( R_23746_9636ed8, \51509 );
buf \U$labaj6832 ( R_23748_b806eb8, \51514 );
buf \U$labaj6833 ( R_2374a_9637028, \51519 );
buf \U$labaj6834 ( R_2374c_b806f60, \51524 );
buf \U$labaj6835 ( R_2374e_b8070b0, \51529 );
buf \U$labaj6836 ( R_23750_9d33308, \51534 );
buf \U$labaj6837 ( R_23752_b807158, \51539 );
buf \U$labaj6838 ( R_23754_9ef5880, \51544 );
buf \U$labaj6839 ( R_23756_9d26798, \51549 );
buf \U$labaj6840 ( R_23758_9d342c8, \51554 );
buf \U$labaj6841 ( R_2375a_9ef5928, \51559 );
buf \U$labaj6842 ( R_2375c_96c2b20, \51564 );
buf \U$labaj6843 ( R_2375e_9d31820, \51569 );
buf \U$labaj6844 ( R_23760_9d31970, \51574 );
buf \U$labaj6845 ( R_23762_9637178, \51579 );
buf \U$labaj6846 ( R_23764_9d26840, \51584 );
buf \U$labaj6847 ( R_23766_96372c8, \51589 );
buf \U$labaj6848 ( R_23768_9d268e8, \51594 );
buf \U$labaj6849 ( R_2376a_9d26a38, \51599 );
buf \U$labaj6850 ( R_2376c_9d26ae0, \51604 );
buf \U$labaj6851 ( R_2376e_9637370, \51609 );
buf \U$labaj6852 ( R_23770_9d26b88, \51614 );
buf \U$labaj6853 ( R_23772_9637418, \51619 );
buf \U$labaj6854 ( R_2398c_96c2fb8, \51626 );
buf \U$labaj6855 ( R_2398e_9559c70, \51631 );
buf \U$labaj6856 ( R_23990_96c35a0, \51636 );
buf \U$labaj6857 ( R_23992_96e8010, \51641 );
buf \U$labaj6858 ( R_23994_955a300, \51646 );
buf \U$labaj6859 ( R_23996_955a450, \51651 );
buf \U$labaj6860 ( R_23998_9d34ca0, \51656 );
buf \U$labaj6861 ( R_2399a_96c3840, \51661 );
buf \U$labaj6862 ( R_2398a_9d34d48, \51666 );
buf \U$labaj6863 ( R_2399c_96c3a38, \51671 );
buf \U$labaj6864 ( R_2399e_96c3d80, \51676 );
buf \U$labaj6865 ( R_239a0_955a840, \51681 );
buf \U$labaj6866 ( R_239a2_96c59b8, \51686 );
buf \U$labaj6867 ( R_23988_96eaf50, \51842 );
buf \U$labaj6868 ( R_239ba_96ca728, \51845 );
buf \U$labaj6869 ( R_239bc_955b8a8, \51848 );
buf \U$labaj6870 ( R_239be_b7db6e8, \51851 );
buf \U$labaj6871 ( R_234dc_b8085b0, \51878 );
buf \U$labaj6872 ( R_234f2_b80b988, \51887 );
buf \U$labaj6873 ( R_23508_b808658, \51896 );
buf \U$labaj6874 ( R_2351e_b808700, \51905 );
buf \U$labaj6875 ( R_23534_b8087a8, \51914 );
buf \U$labaj6876 ( R_2354a_b8088f8, \51923 );
buf \U$labaj6877 ( R_23554_b80ba30, \51932 );
buf \U$labaj6878 ( R_23556_b80bb80, \51941 );
buf \U$labaj6879 ( R_23558_b80bec8, \51950 );
buf \U$labaj6880 ( R_2355a_b80bf70, \51959 );
buf \U$labaj6881 ( R_234de_b8089a0, \51968 );
buf \U$labaj6882 ( R_234e0_b808a48, \51977 );
buf \U$labaj6883 ( R_234e2_b809768, \51986 );
buf \U$labaj6884 ( R_234e4_b809df8, \51995 );
buf \U$labaj6885 ( R_234e6_b80c2b8, \52004 );
buf \U$labaj6886 ( R_234e8_b80e040, \52013 );
buf \U$labaj6887 ( R_234ea_b80e580, \52022 );
buf \U$labaj6888 ( R_234ec_b80c600, \52031 );
buf \U$labaj6889 ( R_234ee_b80f0a8, \52040 );
buf \U$labaj6890 ( R_234f0_b80fd20, \52049 );
buf \U$labaj6891 ( R_234f4_b80c750, \52058 );
buf \U$labaj6892 ( R_234f6_b80ffc0, \52067 );
buf \U$labaj6893 ( R_234f8_b7ddf98, \52076 );
buf \U$labaj6894 ( R_234fa_b80c7f8, \52085 );
buf \U$labaj6895 ( R_234fc_b7de0e8, \52094 );
buf \U$labaj6896 ( R_234fe_b7de388, \52103 );
buf \U$labaj6897 ( R_23500_b7de430, \52112 );
buf \U$labaj6898 ( R_23502_b80c9f0, \52121 );
buf \U$labaj6899 ( R_23504_b7de580, \52130 );
buf \U$labaj6900 ( R_23506_b80ca98, \52139 );
buf \U$labaj6901 ( R_2350a_b7de820, \52148 );
buf \U$labaj6902 ( R_2350c_b7dea18, \52157 );
buf \U$labaj6903 ( R_2350e_b7dee08, \52166 );
buf \U$labaj6904 ( R_23510_b80cc90, \52175 );
buf \U$labaj6905 ( R_23512_b80cd38, \52184 );
buf \U$labaj6906 ( R_23514_b7df1f8, \52193 );
buf \U$labaj6907 ( R_23516_b80ce88, \52202 );
buf \U$labaj6908 ( R_23518_b7df348, \52211 );
buf \U$labaj6909 ( R_2351a_b7df540, \52220 );
buf \U$labaj6910 ( R_2351c_b80cf30, \52229 );
buf \U$labaj6911 ( R_23520_b7dfc78, \52238 );
buf \U$labaj6912 ( R_23522_b80d080, \52247 );
buf \U$labaj6913 ( R_23524_b80d278, \52256 );
buf \U$labaj6914 ( R_23526_b7dff18, \52265 );
buf \U$labaj6915 ( R_23528_b80d320, \52274 );
buf \U$labaj6916 ( R_2352a_b7e0068, \52283 );
buf \U$labaj6917 ( R_2352c_b80d5c0, \52292 );
buf \U$labaj6918 ( R_2352e_b7e01b8, \52301 );
buf \U$labaj6919 ( R_23530_b80d668, \52310 );
buf \U$labaj6920 ( R_23532_b7e0458, \52319 );
buf \U$labaj6921 ( R_23536_b7e05a8, \52328 );
buf \U$labaj6922 ( R_23538_b80d7b8, \52337 );
buf \U$labaj6923 ( R_2353a_b80de48, \52346 );
buf \U$labaj6924 ( R_2353c_b7e0998, \52355 );
buf \U$labaj6925 ( R_2353e_b7e0b90, \52364 );
buf \U$labaj6926 ( R_23540_b7e1178, \52373 );
buf \U$labaj6927 ( R_23542_b80e430, \52382 );
buf \U$labaj6928 ( R_23544_b80e628, \52391 );
buf \U$labaj6929 ( R_23546_b80e778, \52400 );
buf \U$labaj6930 ( R_23548_b7e1568, \52409 );
buf \U$labaj6931 ( R_2354c_b80e970, \52418 );
buf \U$labaj6932 ( R_2354e_b7e16b8, \52427 );
buf \U$labaj6933 ( R_23550_b80eb68, \52436 );
buf \U$labaj6934 ( R_23552_b7e1808, \52445 );
buf \U$labaj6935 ( R_2355c_b7e18b0, \52456 );
buf \U$labaj6936 ( R_23572_b805c58, \52463 );
buf \U$labaj6937 ( R_23588_b7e1958, \52470 );
buf \U$labaj6938 ( R_2359e_b80ed60, \52477 );
buf \U$labaj6939 ( R_235b4_95ad7d8, \52484 );
buf \U$labaj6940 ( R_235ca_b806438, \52491 );
buf \U$labaj6941 ( R_235d4_b7e1a00, \52498 );
buf \U$labaj6942 ( R_235d6_b80f000, \52505 );
buf \U$labaj6943 ( R_235d8_b7e1bf8, \52512 );
buf \U$labaj6944 ( R_235da_b7e1ca0, \52519 );
buf \U$labaj6945 ( R_2355e_b7e1e98, \52526 );
buf \U$labaj6946 ( R_23560_95ad9d0, \52533 );
buf \U$labaj6947 ( R_23562_b7e1f40, \52540 );
buf \U$labaj6948 ( R_23564_95adb20, \52547 );
buf \U$labaj6949 ( R_23566_b7e1fe8, \52554 );
buf \U$labaj6950 ( R_23568_b80f3f0, \52561 );
buf \U$labaj6951 ( R_2356a_b80f5e8, \52568 );
buf \U$labaj6952 ( R_2356c_b806630, \52575 );
buf \U$labaj6953 ( R_2356e_b7e2090, \52582 );
buf \U$labaj6954 ( R_23570_b80f690, \52589 );
buf \U$labaj6955 ( R_23574_b7e2138, \52596 );
buf \U$labaj6956 ( R_23576_b7e21e0, \52603 );
buf \U$labaj6957 ( R_23578_b7e23d8, \52610 );
buf \U$labaj6958 ( R_2357a_b7e2720, \52617 );
buf \U$labaj6959 ( R_2357c_b7e2870, \52624 );
buf \U$labaj6960 ( R_2357e_b7e29c0, \52631 );
buf \U$labaj6961 ( R_23580_b806828, \52638 );
buf \U$labaj6962 ( R_23582_b7e2a68, \52645 );
buf \U$labaj6963 ( R_23584_b7e2c60, \52652 );
buf \U$labaj6964 ( R_23586_b7e2f00, \52659 );
buf \U$labaj6965 ( R_2358a_b80f7e0, \52666 );
buf \U$labaj6966 ( R_2358c_96cb8e0, \52673 );
buf \U$labaj6967 ( R_2358e_b7e2fa8, \52680 );
buf \U$labaj6968 ( R_23590_b7e30f8, \52687 );
buf \U$labaj6969 ( R_23592_b806978, \52694 );
buf \U$labaj6970 ( R_23594_b807008, \52701 );
buf \U$labaj6971 ( R_23596_b7e32f0, \52708 );
buf \U$labaj6972 ( R_23598_b80fb28, \52715 );
buf \U$labaj6973 ( R_2359a_b7e3398, \52722 );
buf \U$labaj6974 ( R_2359c_b807698, \52729 );
buf \U$labaj6975 ( R_235a0_b7e34e8, \52736 );
buf \U$labaj6976 ( R_235a2_96cbb80, \52743 );
buf \U$labaj6977 ( R_235a4_b80fbd0, \52750 );
buf \U$labaj6978 ( R_235a6_96cc018, \52757 );
buf \U$labaj6979 ( R_235a8_95adf10, \52764 );
buf \U$labaj6980 ( R_235aa_b7e36e0, \52771 );
buf \U$labaj6981 ( R_235ac_b807890, \52778 );
buf \U$labaj6982 ( R_235ae_b7e3788, \52785 );
buf \U$labaj6983 ( R_235b0_b7e38d8, \52792 );
buf \U$labaj6984 ( R_235b2_b7e3ad0, \52799 );
buf \U$labaj6985 ( R_235b6_b7e3cc8, \52806 );
buf \U$labaj6986 ( R_235b8_b7e3f68, \52813 );
buf \U$labaj6987 ( R_235ba_b807f20, \52820 );
buf \U$labaj6988 ( R_235bc_b807fc8, \52827 );
buf \U$labaj6989 ( R_235be_b8101b8, \52834 );
buf \U$labaj6990 ( R_235c0_b7e40b8, \52841 );
buf \U$labaj6991 ( R_235c2_b7e4208, \52848 );
buf \U$labaj6992 ( R_235c4_b8105a8, \52855 );
buf \U$labaj6993 ( R_235c6_b810650, \52862 );
buf \U$labaj6994 ( R_235c8_96cc210, \52869 );
buf \U$labaj6995 ( R_235cc_b7e42b0, \52876 );
buf \U$labaj6996 ( R_235ce_b7e4400, \52883 );
buf \U$labaj6997 ( R_235d0_b7e4550, \52890 );
buf \U$labaj6998 ( R_235d2_b7e45f8, \52897 );
buf \U$labaj6999 ( R_235dc_b8106f8, \52906 );
buf \U$labaj7000 ( R_235f2_b7e46a0, \52913 );
buf \U$labaj7001 ( R_23608_b808118, \52920 );
buf \U$labaj7002 ( R_2361e_b7e47f0, \52927 );
buf \U$labaj7003 ( R_23634_b7e49e8, \52934 );
buf \U$labaj7004 ( R_2364a_b7dd860, \52941 );
buf \U$labaj7005 ( R_23654_95ae060, \52948 );
buf \U$labaj7006 ( R_23656_b7dd908, \52955 );
buf \U$labaj7007 ( R_23658_b7ddda0, \52962 );
buf \U$labaj7008 ( R_2365a_b7dde48, \52969 );
buf \U$labaj7009 ( R_235de_9637b50, \52976 );
buf \U$labaj7010 ( R_235e0_95ae1b0, \52983 );
buf \U$labaj7011 ( R_235e2_b7ddef0, \52990 );
buf \U$labaj7012 ( R_235e4_b7de238, \52997 );
buf \U$labaj7013 ( R_235e6_b7e4b38, \53004 );
buf \U$labaj7014 ( R_235e8_9637fe8, \53011 );
buf \U$labaj7015 ( R_235ea_b7de2e0, \53018 );
buf \U$labaj7016 ( R_235ec_b808310, \53025 );
buf \U$labaj7017 ( R_235ee_9638138, \53032 );
buf \U$labaj7018 ( R_235f0_96381e0, \53039 );
buf \U$labaj7019 ( R_235f4_b7e4d30, \53046 );
buf \U$labaj7020 ( R_235f6_96383d8, \53053 );
buf \U$labaj7021 ( R_235f8_b7de6d0, \53060 );
buf \U$labaj7022 ( R_235fa_9638480, \53067 );
buf \U$labaj7023 ( R_235fc_b7de8c8, \53074 );
buf \U$labaj7024 ( R_235fe_9638528, \53081 );
buf \U$labaj7025 ( R_23600_96385d0, \53088 );
buf \U$labaj7026 ( R_23602_b7de970, \53095 );
buf \U$labaj7027 ( R_23604_b7deac0, \53102 );
buf \U$labaj7028 ( R_23606_9638678, \53109 );
buf \U$labaj7029 ( R_2360a_96387c8, \53116 );
buf \U$1 ( \7056 , RIde67cd8_3982);
not \U$2 ( \7057 , \7056 );
buf \U$3 ( \7058 , \7057 );
nor \U$5 ( \7059 , RIde67cd8_3982, RIde68638_3981, RIde68f20_3980);
_HMUX g14890 ( \7060_nG14890 , \7058 , 1'b0 , \7059 );
not \U$6 ( \7061 , RIe549ef0_6842);
not \U$7 ( \7062 , RIe549770_6843);
not \U$8 ( \7063 , RIea91330_6888);
and \U$9 ( \7064 , RIe5319e0_6884, \7061 , \7062 , RIe548ff0_6844, \7063 );
buf \U$10 ( \7065 , \7064 );
buf \U$11 ( \7066 , RIb79b4a0_271);
and \U$12 ( \7067 , \7065 , \7066 );
_HMUX g14891 ( \7068_nG14891 , RIde67cd8_3982 , \7060_nG14890 , \7067 );
buf \U$13 ( \7069 , RIde67cd8_3982);
not \U$14 ( \7070 , \7069 );
buf \U$15 ( \7071 , \7070 );
not \U$16 ( \7072 , RIde68f20_3980);
nor \U$17 ( \7073 , RIde67cd8_3982, RIde68638_3981, \7072 );
_HMUX g14897 ( \7074_nG14897 , \7071 , RIde67cd8_3982 , \7073 );
buf \U$18 ( \7075 , RIb79b518_270);
buf \U$19 ( \7076 , RIe5319e0_6884);
not \U$20 ( \7077 , \7076 );
buf \U$21 ( \7078 , \7077 );
buf \U$22 ( \7079 , RIe549ef0_6842);
xnor \U$23 ( \7080 , \7079 , \7076 );
buf \U$24 ( \7081 , \7080 );
buf \U$25 ( \7082 , RIe549770_6843);
or \U$26 ( \7083 , \7079 , \7076 );
xnor \U$27 ( \7084 , \7082 , \7083 );
buf \U$28 ( \7085 , \7084 );
buf \U$29 ( \7086 , RIe548ff0_6844);
or \U$30 ( \7087 , \7082 , \7083 );
xnor \U$31 ( \7088 , \7086 , \7087 );
buf \U$32 ( \7089 , \7088 );
buf \U$33 ( \7090 , RIea91330_6888);
or \U$34 ( \7091 , \7086 , \7087 );
xor \U$35 ( \7092 , \7090 , \7091 );
buf \U$36 ( \7093 , \7092 );
not \U$37 ( \7094 , \7093 );
and \U$38 ( \7095 , \7090 , \7091 );
buf \U$39 ( \7096 , \7095 );
nor \U$40 ( \7097 , \7078 , \7081 , \7085 , \7089 , \7094 , \7096 );
and \U$41 ( \7098 , RIe5329d0_6883, \7097 );
not \U$42 ( \7099 , \7096 );
and \U$43 ( \7100 , \7078 , \7081 , \7085 , \7089 , \7094 , \7099 );
and \U$44 ( \7101 , RIeb72150_6905, \7100 );
or \U$59 ( \7102 , \7098 , \7101 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
buf \U$61 ( \7103 , \7096 );
buf \U$62 ( \7104 , \7093 );
buf \U$63 ( \7105 , \7078 );
buf \U$64 ( \7106 , \7081 );
buf \U$65 ( \7107 , \7085 );
buf \U$66 ( \7108 , \7089 );
or \U$67 ( \7109 , \7105 , \7106 , \7107 , \7108 );
and \U$68 ( \7110 , \7104 , \7109 );
or \U$69 ( \7111 , \7103 , \7110 );
buf \U$70 ( \7112 , \7111 );
or \U$71 ( \7113 , 1'b0 , \7112 );
_DC g32b3 ( \7114_nG32b3 , \7102 , \7113 );
not \U$72 ( \7115 , \7114_nG32b3 );
buf \U$73 ( \7116 , RIb7b9608_246);
buf \U$74 ( \7117 , RIe5c6738_6786);
and \U$75 ( \7118 , \7117 , \7097 );
buf \U$76 ( \7119 , RIe4fc9e8_6393);
and \U$77 ( \7120 , \7119 , \7100 );
or \U$92 ( \7121 , \7118 , \7120 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g32bb ( \7122_nG32bb , \7121 , \7113 );
buf \U$93 ( \7123 , \7122_nG32bb );
xor \U$94 ( \7124 , \7116 , \7123 );
buf \U$95 ( \7125 , RIb7b9590_247);
buf \U$96 ( \7126 , RIe5c5bf8_6787);
and \U$97 ( \7127 , \7126 , \7097 );
buf \U$98 ( \7128 , RIe4fbcc8_6394);
and \U$99 ( \7129 , \7128 , \7100 );
or \U$114 ( \7130 , \7127 , \7129 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g32c4 ( \7131_nG32c4 , \7130 , \7113 );
buf \U$115 ( \7132 , \7131_nG32c4 );
xor \U$116 ( \7133 , \7125 , \7132 );
or \U$117 ( \7134 , \7124 , \7133 );
buf \U$118 ( \7135 , RIb7b9518_248);
buf \U$119 ( \7136 , RIe5c4fc8_6788);
and \U$120 ( \7137 , \7136 , \7097 );
buf \U$121 ( \7138 , RIe4faf30_6395);
and \U$122 ( \7139 , \7138 , \7100 );
or \U$137 ( \7140 , \7137 , \7139 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g32ce ( \7141_nG32ce , \7140 , \7113 );
buf \U$138 ( \7142 , \7141_nG32ce );
xor \U$139 ( \7143 , \7135 , \7142 );
or \U$140 ( \7144 , \7134 , \7143 );
buf \U$141 ( \7145 , RIb7b94a0_249);
buf \U$142 ( \7146 , RIe5c4500_6789);
and \U$143 ( \7147 , \7146 , \7097 );
buf \U$144 ( \7148 , RIe4fa198_6396);
and \U$145 ( \7149 , \7148 , \7100 );
or \U$160 ( \7150 , \7147 , \7149 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g32d8 ( \7151_nG32d8 , \7150 , \7113 );
buf \U$161 ( \7152 , \7151_nG32d8 );
xor \U$162 ( \7153 , \7145 , \7152 );
or \U$163 ( \7154 , \7144 , \7153 );
buf \U$164 ( \7155 , RIb7b9428_250);
buf \U$165 ( \7156 , RIe5c3948_6790);
and \U$166 ( \7157 , \7156 , \7097 );
buf \U$167 ( \7158 , RIe4f9388_6397);
and \U$168 ( \7159 , \7158 , \7100 );
or \U$183 ( \7160 , \7157 , \7159 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g32e2 ( \7161_nG32e2 , \7160 , \7113 );
buf \U$184 ( \7162 , \7161_nG32e2 );
xor \U$185 ( \7163 , \7155 , \7162 );
or \U$186 ( \7164 , \7154 , \7163 );
buf \U$187 ( \7165 , RIb7b93b0_251);
buf \U$188 ( \7166 , RIe5c2e08_6791);
and \U$189 ( \7167 , \7166 , \7097 );
buf \U$190 ( \7168 , RIe4f85f0_6398);
and \U$191 ( \7169 , \7168 , \7100 );
or \U$206 ( \7170 , \7167 , \7169 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g32ec ( \7171_nG32ec , \7170 , \7113 );
buf \U$207 ( \7172 , \7171_nG32ec );
xor \U$208 ( \7173 , \7165 , \7172 );
or \U$209 ( \7174 , \7164 , \7173 );
buf \U$210 ( \7175 , RIb7af720_252);
buf \U$211 ( \7176 , RIe5c22c8_6792);
and \U$212 ( \7177 , \7176 , \7097 );
buf \U$213 ( \7178 , RIe4f7a38_6399);
and \U$214 ( \7179 , \7178 , \7100 );
or \U$229 ( \7180 , \7177 , \7179 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g32f6 ( \7181_nG32f6 , \7180 , \7113 );
buf \U$230 ( \7182 , \7181_nG32f6 );
xor \U$231 ( \7183 , \7175 , \7182 );
or \U$232 ( \7184 , \7174 , \7183 );
buf \U$233 ( \7185 , RIb7af6a8_253);
buf \U$234 ( \7186 , RIe5c1710_6793);
and \U$235 ( \7187 , \7186 , \7097 );
buf \U$236 ( \7188 , RIe4f6ef8_6400);
and \U$237 ( \7189 , \7188 , \7100 );
or \U$252 ( \7190 , \7187 , \7189 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3300 ( \7191_nG3300 , \7190 , \7113 );
buf \U$253 ( \7192 , \7191_nG3300 );
xor \U$254 ( \7193 , \7185 , \7192 );
or \U$255 ( \7194 , \7184 , \7193 );
not \U$256 ( \7195 , \7194 );
buf \U$257 ( \7196 , \7195 );
buf \U$258 ( \7197 , RIb7af630_254);
buf \U$259 ( \7198 , RIe5e09d0_6767);
and \U$260 ( \7199 , \7198 , \7097 );
buf \U$261 ( \7200 , RIe4af828_6445);
and \U$262 ( \7201 , \7200 , \7100 );
or \U$277 ( \7202 , \7199 , \7201 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g330c ( \7203_nG330c , \7202 , \7113 );
buf \U$278 ( \7204 , \7203_nG330c );
xor \U$279 ( \7205 , \7197 , \7204 );
buf \U$280 ( \7206 , RIb7af5b8_255);
buf \U$281 ( \7207 , RIe5e1330_6766);
and \U$282 ( \7208 , \7207 , \7097 );
buf \U$283 ( \7209 , RIe519818_6368);
and \U$284 ( \7210 , \7209 , \7100 );
or \U$299 ( \7211 , \7208 , \7210 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3315 ( \7212_nG3315 , \7211 , \7113 );
buf \U$300 ( \7213 , \7212_nG3315 );
xor \U$301 ( \7214 , \7206 , \7213 );
or \U$302 ( \7215 , \7205 , \7214 );
buf \U$303 ( \7216 , RIb7af540_256);
buf \U$304 ( \7217 , RIe5e1ba0_6765);
and \U$305 ( \7218 , \7217 , \7097 );
buf \U$306 ( \7219 , RIe4b0200_6444);
and \U$307 ( \7220 , \7219 , \7100 );
or \U$322 ( \7221 , \7218 , \7220 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g331f ( \7222_nG331f , \7221 , \7113 );
buf \U$323 ( \7223 , \7222_nG331f );
xor \U$324 ( \7224 , \7216 , \7223 );
or \U$325 ( \7225 , \7215 , \7224 );
buf \U$326 ( \7226 , RIb7af4c8_257);
buf \U$327 ( \7227 , RIe5e2488_6764);
and \U$328 ( \7228 , \7227 , \7097 );
buf \U$329 ( \7229 , RIe51a2e0_6367);
and \U$330 ( \7230 , \7229 , \7100 );
or \U$345 ( \7231 , \7228 , \7230 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3329 ( \7232_nG3329 , \7231 , \7113 );
buf \U$346 ( \7233 , \7232_nG3329 );
xor \U$347 ( \7234 , \7226 , \7233 );
or \U$348 ( \7235 , \7225 , \7234 );
buf \U$349 ( \7236 , RIb7af450_258);
buf \U$350 ( \7237 , RIe5e2d70_6763);
and \U$351 ( \7238 , \7237 , \7097 );
buf \U$352 ( \7239 , RIe4bdce8_6441);
and \U$353 ( \7240 , \7239 , \7100 );
or \U$368 ( \7241 , \7238 , \7240 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3331 ( \7242_nG3331 , \7241 , \7113 );
buf \U$369 ( \7243 , \7242_nG3331 );
xor \U$370 ( \7244 , \7236 , \7243 );
or \U$371 ( \7245 , \7235 , \7244 );
buf \U$372 ( \7246 , RIb7af3d8_259);
buf \U$373 ( \7247 , RIe5e3568_6762);
and \U$374 ( \7248 , \7247 , \7097 );
buf \U$375 ( \7249 , RIe51acb8_6366);
and \U$376 ( \7250 , \7249 , \7100 );
or \U$391 ( \7251 , \7248 , \7250 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3339 ( \7252_nG3339 , \7251 , \7113 );
buf \U$392 ( \7253 , \7252_nG3339 );
xor \U$393 ( \7254 , \7246 , \7253 );
or \U$394 ( \7255 , \7245 , \7254 );
buf \U$395 ( \7256 , RIb7a5bf8_260);
buf \U$396 ( \7257 , RIe588848_6840);
and \U$397 ( \7258 , \7257 , \7097 );
buf \U$398 ( \7259 , RIe4bd310_6442);
and \U$399 ( \7260 , \7259 , \7100 );
or \U$414 ( \7261 , \7258 , \7260 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3341 ( \7262_nG3341 , \7261 , \7113 );
buf \U$415 ( \7263 , \7262_nG3341 );
xor \U$416 ( \7264 , \7256 , \7263 );
or \U$417 ( \7265 , \7255 , \7264 );
buf \U$418 ( \7266 , RIb7a0c48_261);
buf \U$419 ( \7267 , RIe5e3e50_6761);
and \U$420 ( \7268 , \7267 , \7097 );
buf \U$421 ( \7269 , RIe4b0a70_6443);
and \U$422 ( \7270 , \7269 , \7100 );
or \U$437 ( \7271 , \7268 , \7270 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3349 ( \7272_nG3349 , \7271 , \7113 );
buf \U$438 ( \7273 , \7272_nG3349 );
xor \U$439 ( \7274 , \7266 , \7273 );
or \U$440 ( \7275 , \7265 , \7274 );
not \U$441 ( \7276 , \7275 );
buf \U$442 ( \7277 , \7276 );
and \U$443 ( \7278 , \7196 , \7277 );
and \U$444 ( \7279 , \7115 , \7278 );
_HMUX g3351 ( \7280_nG3351 , RIe5319e0_6884 , \7078 , \7279 );
buf \U$447 ( \7281 , \7078 );
buf \U$450 ( \7282 , \7081 );
buf \U$453 ( \7283 , \7085 );
buf \U$456 ( \7284 , \7089 );
buf \U$457 ( \7285 , \7093 );
not \U$458 ( \7286 , \7285 );
buf \U$459 ( \7287 , \7286 );
not \U$460 ( \7288 , \7287 );
buf \U$461 ( \7289 , \7096 );
xnor \U$462 ( \7290 , \7289 , \7285 );
buf \U$463 ( \7291 , \7290 );
or \U$464 ( \7292 , \7289 , \7285 );
not \U$465 ( \7293 , \7292 );
buf \U$466 ( \7294 , \7293 );
buf \U$467 ( \7295 , \7294 );
buf \U$468 ( \7296 , \7294 );
buf \U$469 ( \7297 , \7294 );
buf \U$470 ( \7298 , \7294 );
buf \U$471 ( \7299 , \7294 );
buf \U$472 ( \7300 , \7294 );
buf \U$473 ( \7301 , \7294 );
buf \U$474 ( \7302 , \7294 );
buf \U$475 ( \7303 , \7294 );
buf \U$476 ( \7304 , \7294 );
buf \U$477 ( \7305 , \7294 );
buf \U$478 ( \7306 , \7294 );
buf \U$479 ( \7307 , \7294 );
buf \U$480 ( \7308 , \7294 );
buf \U$481 ( \7309 , \7294 );
buf \U$482 ( \7310 , \7294 );
buf \U$483 ( \7311 , \7294 );
buf \U$484 ( \7312 , \7294 );
buf \U$485 ( \7313 , \7294 );
buf \U$486 ( \7314 , \7294 );
buf \U$487 ( \7315 , \7294 );
buf \U$488 ( \7316 , \7294 );
buf \U$489 ( \7317 , \7294 );
buf \U$490 ( \7318 , \7294 );
buf \U$491 ( \7319 , \7294 );
nor \U$492 ( \7320 , \7281 , \7282 , \7283 , \7284 , \7288 , \7291 , \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 , \7303 , \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 , \7313 , \7314 , \7315 , \7316 , \7317 , \7318 , \7319 );
and \U$493 ( \7321 , RIe5329d0_6883, \7320 );
not \U$494 ( \7322 , \7281 );
not \U$495 ( \7323 , \7282 );
not \U$496 ( \7324 , \7283 );
not \U$497 ( \7325 , \7284 );
buf \U$498 ( \7326 , \7294 );
buf \U$499 ( \7327 , \7294 );
buf \U$500 ( \7328 , \7294 );
buf \U$501 ( \7329 , \7294 );
buf \U$502 ( \7330 , \7294 );
buf \U$503 ( \7331 , \7294 );
buf \U$504 ( \7332 , \7294 );
buf \U$505 ( \7333 , \7294 );
buf \U$506 ( \7334 , \7294 );
buf \U$507 ( \7335 , \7294 );
buf \U$508 ( \7336 , \7294 );
buf \U$509 ( \7337 , \7294 );
buf \U$510 ( \7338 , \7294 );
buf \U$511 ( \7339 , \7294 );
buf \U$512 ( \7340 , \7294 );
buf \U$513 ( \7341 , \7294 );
buf \U$514 ( \7342 , \7294 );
buf \U$515 ( \7343 , \7294 );
buf \U$516 ( \7344 , \7294 );
buf \U$517 ( \7345 , \7294 );
buf \U$518 ( \7346 , \7294 );
buf \U$519 ( \7347 , \7294 );
buf \U$520 ( \7348 , \7294 );
buf \U$521 ( \7349 , \7294 );
buf \U$522 ( \7350 , \7294 );
nor \U$523 ( \7351 , \7322 , \7323 , \7324 , \7325 , \7287 , \7291 , \7294 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 , \7333 , \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 , \7343 , \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 );
and \U$524 ( \7352 , RIeb72150_6905, \7351 );
buf \U$525 ( \7353 , \7294 );
buf \U$526 ( \7354 , \7294 );
buf \U$527 ( \7355 , \7294 );
buf \U$528 ( \7356 , \7294 );
buf \U$529 ( \7357 , \7294 );
buf \U$530 ( \7358 , \7294 );
buf \U$531 ( \7359 , \7294 );
buf \U$532 ( \7360 , \7294 );
buf \U$533 ( \7361 , \7294 );
buf \U$534 ( \7362 , \7294 );
buf \U$535 ( \7363 , \7294 );
buf \U$536 ( \7364 , \7294 );
buf \U$537 ( \7365 , \7294 );
buf \U$538 ( \7366 , \7294 );
buf \U$539 ( \7367 , \7294 );
buf \U$540 ( \7368 , \7294 );
buf \U$541 ( \7369 , \7294 );
buf \U$542 ( \7370 , \7294 );
buf \U$543 ( \7371 , \7294 );
buf \U$544 ( \7372 , \7294 );
buf \U$545 ( \7373 , \7294 );
buf \U$546 ( \7374 , \7294 );
buf \U$547 ( \7375 , \7294 );
buf \U$548 ( \7376 , \7294 );
buf \U$549 ( \7377 , \7294 );
nor \U$550 ( \7378 , \7281 , \7323 , \7324 , \7325 , \7287 , \7291 , \7294 , \7353 , \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 , \7363 , \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 , \7373 , \7374 , \7375 , \7376 , \7377 );
and \U$551 ( \7379 , RIeab80c0_6897, \7378 );
buf \U$552 ( \7380 , \7294 );
buf \U$553 ( \7381 , \7294 );
buf \U$554 ( \7382 , \7294 );
buf \U$555 ( \7383 , \7294 );
buf \U$556 ( \7384 , \7294 );
buf \U$557 ( \7385 , \7294 );
buf \U$558 ( \7386 , \7294 );
buf \U$559 ( \7387 , \7294 );
buf \U$560 ( \7388 , \7294 );
buf \U$561 ( \7389 , \7294 );
buf \U$562 ( \7390 , \7294 );
buf \U$563 ( \7391 , \7294 );
buf \U$564 ( \7392 , \7294 );
buf \U$565 ( \7393 , \7294 );
buf \U$566 ( \7394 , \7294 );
buf \U$567 ( \7395 , \7294 );
buf \U$568 ( \7396 , \7294 );
buf \U$569 ( \7397 , \7294 );
buf \U$570 ( \7398 , \7294 );
buf \U$571 ( \7399 , \7294 );
buf \U$572 ( \7400 , \7294 );
buf \U$573 ( \7401 , \7294 );
buf \U$574 ( \7402 , \7294 );
buf \U$575 ( \7403 , \7294 );
buf \U$576 ( \7404 , \7294 );
nor \U$577 ( \7405 , \7322 , \7282 , \7324 , \7325 , \7287 , \7291 , \7294 , \7380 , \7381 , \7382 , \7383 , \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 , \7393 , \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 , \7403 , \7404 );
and \U$578 ( \7406 , RIe5331c8_6882, \7405 );
buf \U$579 ( \7407 , \7294 );
buf \U$580 ( \7408 , \7294 );
buf \U$581 ( \7409 , \7294 );
buf \U$582 ( \7410 , \7294 );
buf \U$583 ( \7411 , \7294 );
buf \U$584 ( \7412 , \7294 );
buf \U$585 ( \7413 , \7294 );
buf \U$586 ( \7414 , \7294 );
buf \U$587 ( \7415 , \7294 );
buf \U$588 ( \7416 , \7294 );
buf \U$589 ( \7417 , \7294 );
buf \U$590 ( \7418 , \7294 );
buf \U$591 ( \7419 , \7294 );
buf \U$592 ( \7420 , \7294 );
buf \U$593 ( \7421 , \7294 );
buf \U$594 ( \7422 , \7294 );
buf \U$595 ( \7423 , \7294 );
buf \U$596 ( \7424 , \7294 );
buf \U$597 ( \7425 , \7294 );
buf \U$598 ( \7426 , \7294 );
buf \U$599 ( \7427 , \7294 );
buf \U$600 ( \7428 , \7294 );
buf \U$601 ( \7429 , \7294 );
buf \U$602 ( \7430 , \7294 );
buf \U$603 ( \7431 , \7294 );
nor \U$604 ( \7432 , \7281 , \7282 , \7324 , \7325 , \7287 , \7291 , \7294 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 , \7413 , \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 , \7423 , \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 );
and \U$605 ( \7433 , RIe5339c0_6881, \7432 );
buf \U$606 ( \7434 , \7294 );
buf \U$607 ( \7435 , \7294 );
buf \U$608 ( \7436 , \7294 );
buf \U$609 ( \7437 , \7294 );
buf \U$610 ( \7438 , \7294 );
buf \U$611 ( \7439 , \7294 );
buf \U$612 ( \7440 , \7294 );
buf \U$613 ( \7441 , \7294 );
buf \U$614 ( \7442 , \7294 );
buf \U$615 ( \7443 , \7294 );
buf \U$616 ( \7444 , \7294 );
buf \U$617 ( \7445 , \7294 );
buf \U$618 ( \7446 , \7294 );
buf \U$619 ( \7447 , \7294 );
buf \U$620 ( \7448 , \7294 );
buf \U$621 ( \7449 , \7294 );
buf \U$622 ( \7450 , \7294 );
buf \U$623 ( \7451 , \7294 );
buf \U$624 ( \7452 , \7294 );
buf \U$625 ( \7453 , \7294 );
buf \U$626 ( \7454 , \7294 );
buf \U$627 ( \7455 , \7294 );
buf \U$628 ( \7456 , \7294 );
buf \U$629 ( \7457 , \7294 );
buf \U$630 ( \7458 , \7294 );
nor \U$631 ( \7459 , \7322 , \7323 , \7283 , \7325 , \7287 , \7291 , \7294 , \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 , \7442 , \7443 , \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 , \7452 , \7453 , \7454 , \7455 , \7456 , \7457 , \7458 );
and \U$632 ( \7460 , RIeab87c8_6898, \7459 );
buf \U$633 ( \7461 , \7294 );
buf \U$634 ( \7462 , \7294 );
buf \U$635 ( \7463 , \7294 );
buf \U$636 ( \7464 , \7294 );
buf \U$637 ( \7465 , \7294 );
buf \U$638 ( \7466 , \7294 );
buf \U$639 ( \7467 , \7294 );
buf \U$640 ( \7468 , \7294 );
buf \U$641 ( \7469 , \7294 );
buf \U$642 ( \7470 , \7294 );
buf \U$643 ( \7471 , \7294 );
buf \U$644 ( \7472 , \7294 );
buf \U$645 ( \7473 , \7294 );
buf \U$646 ( \7474 , \7294 );
buf \U$647 ( \7475 , \7294 );
buf \U$648 ( \7476 , \7294 );
buf \U$649 ( \7477 , \7294 );
buf \U$650 ( \7478 , \7294 );
buf \U$651 ( \7479 , \7294 );
buf \U$652 ( \7480 , \7294 );
buf \U$653 ( \7481 , \7294 );
buf \U$654 ( \7482 , \7294 );
buf \U$655 ( \7483 , \7294 );
buf \U$656 ( \7484 , \7294 );
buf \U$657 ( \7485 , \7294 );
nor \U$658 ( \7486 , \7281 , \7323 , \7283 , \7325 , \7287 , \7291 , \7294 , \7461 , \7462 , \7463 , \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 , \7472 , \7473 , \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 , \7482 , \7483 , \7484 , \7485 );
and \U$659 ( \7487 , RIe5341b8_6880, \7486 );
buf \U$660 ( \7488 , \7294 );
buf \U$661 ( \7489 , \7294 );
buf \U$662 ( \7490 , \7294 );
buf \U$663 ( \7491 , \7294 );
buf \U$664 ( \7492 , \7294 );
buf \U$665 ( \7493 , \7294 );
buf \U$666 ( \7494 , \7294 );
buf \U$667 ( \7495 , \7294 );
buf \U$668 ( \7496 , \7294 );
buf \U$669 ( \7497 , \7294 );
buf \U$670 ( \7498 , \7294 );
buf \U$671 ( \7499 , \7294 );
buf \U$672 ( \7500 , \7294 );
buf \U$673 ( \7501 , \7294 );
buf \U$674 ( \7502 , \7294 );
buf \U$675 ( \7503 , \7294 );
buf \U$676 ( \7504 , \7294 );
buf \U$677 ( \7505 , \7294 );
buf \U$678 ( \7506 , \7294 );
buf \U$679 ( \7507 , \7294 );
buf \U$680 ( \7508 , \7294 );
buf \U$681 ( \7509 , \7294 );
buf \U$682 ( \7510 , \7294 );
buf \U$683 ( \7511 , \7294 );
buf \U$684 ( \7512 , \7294 );
nor \U$685 ( \7513 , \7322 , \7282 , \7283 , \7325 , \7287 , \7291 , \7294 , \7488 , \7489 , \7490 , \7491 , \7492 , \7493 , \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 , \7502 , \7503 , \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 , \7512 );
and \U$686 ( \7514 , RIe5349b0_6879, \7513 );
buf \U$687 ( \7515 , \7294 );
buf \U$688 ( \7516 , \7294 );
buf \U$689 ( \7517 , \7294 );
buf \U$690 ( \7518 , \7294 );
buf \U$691 ( \7519 , \7294 );
buf \U$692 ( \7520 , \7294 );
buf \U$693 ( \7521 , \7294 );
buf \U$694 ( \7522 , \7294 );
buf \U$695 ( \7523 , \7294 );
buf \U$696 ( \7524 , \7294 );
buf \U$697 ( \7525 , \7294 );
buf \U$698 ( \7526 , \7294 );
buf \U$699 ( \7527 , \7294 );
buf \U$700 ( \7528 , \7294 );
buf \U$701 ( \7529 , \7294 );
buf \U$702 ( \7530 , \7294 );
buf \U$703 ( \7531 , \7294 );
buf \U$704 ( \7532 , \7294 );
buf \U$705 ( \7533 , \7294 );
buf \U$706 ( \7534 , \7294 );
buf \U$707 ( \7535 , \7294 );
buf \U$708 ( \7536 , \7294 );
buf \U$709 ( \7537 , \7294 );
buf \U$710 ( \7538 , \7294 );
buf \U$711 ( \7539 , \7294 );
nor \U$712 ( \7540 , \7281 , \7282 , \7283 , \7325 , \7287 , \7291 , \7294 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 , \7522 , \7523 , \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 , \7532 , \7533 , \7534 , \7535 , \7536 , \7537 , \7538 , \7539 );
and \U$713 ( \7541 , RIea94af8_6890, \7540 );
buf \U$714 ( \7542 , \7294 );
buf \U$715 ( \7543 , \7294 );
buf \U$716 ( \7544 , \7294 );
buf \U$717 ( \7545 , \7294 );
buf \U$718 ( \7546 , \7294 );
buf \U$719 ( \7547 , \7294 );
buf \U$720 ( \7548 , \7294 );
buf \U$721 ( \7549 , \7294 );
buf \U$722 ( \7550 , \7294 );
buf \U$723 ( \7551 , \7294 );
buf \U$724 ( \7552 , \7294 );
buf \U$725 ( \7553 , \7294 );
buf \U$726 ( \7554 , \7294 );
buf \U$727 ( \7555 , \7294 );
buf \U$728 ( \7556 , \7294 );
buf \U$729 ( \7557 , \7294 );
buf \U$730 ( \7558 , \7294 );
buf \U$731 ( \7559 , \7294 );
buf \U$732 ( \7560 , \7294 );
buf \U$733 ( \7561 , \7294 );
buf \U$734 ( \7562 , \7294 );
buf \U$735 ( \7563 , \7294 );
buf \U$736 ( \7564 , \7294 );
buf \U$737 ( \7565 , \7294 );
buf \U$738 ( \7566 , \7294 );
nor \U$739 ( \7567 , \7322 , \7323 , \7324 , \7284 , \7287 , \7291 , \7294 , \7542 , \7543 , \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 , \7552 , \7553 , \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 , \7562 , \7563 , \7564 , \7565 , \7566 );
and \U$740 ( \7568 , RIe5351a8_6878, \7567 );
buf \U$741 ( \7569 , \7294 );
buf \U$742 ( \7570 , \7294 );
buf \U$743 ( \7571 , \7294 );
buf \U$744 ( \7572 , \7294 );
buf \U$745 ( \7573 , \7294 );
buf \U$746 ( \7574 , \7294 );
buf \U$747 ( \7575 , \7294 );
buf \U$748 ( \7576 , \7294 );
buf \U$749 ( \7577 , \7294 );
buf \U$750 ( \7578 , \7294 );
buf \U$751 ( \7579 , \7294 );
buf \U$752 ( \7580 , \7294 );
buf \U$753 ( \7581 , \7294 );
buf \U$754 ( \7582 , \7294 );
buf \U$755 ( \7583 , \7294 );
buf \U$756 ( \7584 , \7294 );
buf \U$757 ( \7585 , \7294 );
buf \U$758 ( \7586 , \7294 );
buf \U$759 ( \7587 , \7294 );
buf \U$760 ( \7588 , \7294 );
buf \U$761 ( \7589 , \7294 );
buf \U$762 ( \7590 , \7294 );
buf \U$763 ( \7591 , \7294 );
buf \U$764 ( \7592 , \7294 );
buf \U$765 ( \7593 , \7294 );
nor \U$766 ( \7594 , \7281 , \7323 , \7324 , \7284 , \7287 , \7291 , \7294 , \7569 , \7570 , \7571 , \7572 , \7573 , \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 , \7582 , \7583 , \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 , \7592 , \7593 );
and \U$767 ( \7595 , RIe5359a0_6877, \7594 );
buf \U$768 ( \7596 , \7294 );
buf \U$769 ( \7597 , \7294 );
buf \U$770 ( \7598 , \7294 );
buf \U$771 ( \7599 , \7294 );
buf \U$772 ( \7600 , \7294 );
buf \U$773 ( \7601 , \7294 );
buf \U$774 ( \7602 , \7294 );
buf \U$775 ( \7603 , \7294 );
buf \U$776 ( \7604 , \7294 );
buf \U$777 ( \7605 , \7294 );
buf \U$778 ( \7606 , \7294 );
buf \U$779 ( \7607 , \7294 );
buf \U$780 ( \7608 , \7294 );
buf \U$781 ( \7609 , \7294 );
buf \U$782 ( \7610 , \7294 );
buf \U$783 ( \7611 , \7294 );
buf \U$784 ( \7612 , \7294 );
buf \U$785 ( \7613 , \7294 );
buf \U$786 ( \7614 , \7294 );
buf \U$787 ( \7615 , \7294 );
buf \U$788 ( \7616 , \7294 );
buf \U$789 ( \7617 , \7294 );
buf \U$790 ( \7618 , \7294 );
buf \U$791 ( \7619 , \7294 );
buf \U$792 ( \7620 , \7294 );
nor \U$793 ( \7621 , \7322 , \7282 , \7324 , \7284 , \7287 , \7291 , \7294 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 , \7612 , \7613 , \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 );
and \U$794 ( \7622 , RIeab78c8_6895, \7621 );
buf \U$795 ( \7623 , \7294 );
buf \U$796 ( \7624 , \7294 );
buf \U$797 ( \7625 , \7294 );
buf \U$798 ( \7626 , \7294 );
buf \U$799 ( \7627 , \7294 );
buf \U$800 ( \7628 , \7294 );
buf \U$801 ( \7629 , \7294 );
buf \U$802 ( \7630 , \7294 );
buf \U$803 ( \7631 , \7294 );
buf \U$804 ( \7632 , \7294 );
buf \U$805 ( \7633 , \7294 );
buf \U$806 ( \7634 , \7294 );
buf \U$807 ( \7635 , \7294 );
buf \U$808 ( \7636 , \7294 );
buf \U$809 ( \7637 , \7294 );
buf \U$810 ( \7638 , \7294 );
buf \U$811 ( \7639 , \7294 );
buf \U$812 ( \7640 , \7294 );
buf \U$813 ( \7641 , \7294 );
buf \U$814 ( \7642 , \7294 );
buf \U$815 ( \7643 , \7294 );
buf \U$816 ( \7644 , \7294 );
buf \U$817 ( \7645 , \7294 );
buf \U$818 ( \7646 , \7294 );
buf \U$819 ( \7647 , \7294 );
nor \U$820 ( \7648 , \7281 , \7282 , \7324 , \7284 , \7287 , \7291 , \7294 , \7623 , \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 , \7632 , \7633 , \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 , \7642 , \7643 , \7644 , \7645 , \7646 , \7647 );
and \U$821 ( \7649 , RIeab7d00_6896, \7648 );
buf \U$822 ( \7650 , \7294 );
buf \U$823 ( \7651 , \7294 );
buf \U$824 ( \7652 , \7294 );
buf \U$825 ( \7653 , \7294 );
buf \U$826 ( \7654 , \7294 );
buf \U$827 ( \7655 , \7294 );
buf \U$828 ( \7656 , \7294 );
buf \U$829 ( \7657 , \7294 );
buf \U$830 ( \7658 , \7294 );
buf \U$831 ( \7659 , \7294 );
buf \U$832 ( \7660 , \7294 );
buf \U$833 ( \7661 , \7294 );
buf \U$834 ( \7662 , \7294 );
buf \U$835 ( \7663 , \7294 );
buf \U$836 ( \7664 , \7294 );
buf \U$837 ( \7665 , \7294 );
buf \U$838 ( \7666 , \7294 );
buf \U$839 ( \7667 , \7294 );
buf \U$840 ( \7668 , \7294 );
buf \U$841 ( \7669 , \7294 );
buf \U$842 ( \7670 , \7294 );
buf \U$843 ( \7671 , \7294 );
buf \U$844 ( \7672 , \7294 );
buf \U$845 ( \7673 , \7294 );
buf \U$846 ( \7674 , \7294 );
nor \U$847 ( \7675 , \7322 , \7323 , \7283 , \7284 , \7287 , \7291 , \7294 , \7650 , \7651 , \7652 , \7653 , \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 , \7662 , \7663 , \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 , \7672 , \7673 , \7674 );
and \U$848 ( \7676 , RIeacfa18_6902, \7675 );
buf \U$849 ( \7677 , \7294 );
buf \U$850 ( \7678 , \7294 );
buf \U$851 ( \7679 , \7294 );
buf \U$852 ( \7680 , \7294 );
buf \U$853 ( \7681 , \7294 );
buf \U$854 ( \7682 , \7294 );
buf \U$855 ( \7683 , \7294 );
buf \U$856 ( \7684 , \7294 );
buf \U$857 ( \7685 , \7294 );
buf \U$858 ( \7686 , \7294 );
buf \U$859 ( \7687 , \7294 );
buf \U$860 ( \7688 , \7294 );
buf \U$861 ( \7689 , \7294 );
buf \U$862 ( \7690 , \7294 );
buf \U$863 ( \7691 , \7294 );
buf \U$864 ( \7692 , \7294 );
buf \U$865 ( \7693 , \7294 );
buf \U$866 ( \7694 , \7294 );
buf \U$867 ( \7695 , \7294 );
buf \U$868 ( \7696 , \7294 );
buf \U$869 ( \7697 , \7294 );
buf \U$870 ( \7698 , \7294 );
buf \U$871 ( \7699 , \7294 );
buf \U$872 ( \7700 , \7294 );
buf \U$873 ( \7701 , \7294 );
nor \U$874 ( \7702 , \7281 , \7323 , \7283 , \7284 , \7287 , \7291 , \7294 , \7677 , \7678 , \7679 , \7680 , \7681 , \7682 , \7683 , \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 , \7692 , \7693 , \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 );
and \U$875 ( \7703 , RIeab6518_6891, \7702 );
buf \U$876 ( \7704 , \7294 );
buf \U$877 ( \7705 , \7294 );
buf \U$878 ( \7706 , \7294 );
buf \U$879 ( \7707 , \7294 );
buf \U$880 ( \7708 , \7294 );
buf \U$881 ( \7709 , \7294 );
buf \U$882 ( \7710 , \7294 );
buf \U$883 ( \7711 , \7294 );
buf \U$884 ( \7712 , \7294 );
buf \U$885 ( \7713 , \7294 );
buf \U$886 ( \7714 , \7294 );
buf \U$887 ( \7715 , \7294 );
buf \U$888 ( \7716 , \7294 );
buf \U$889 ( \7717 , \7294 );
buf \U$890 ( \7718 , \7294 );
buf \U$891 ( \7719 , \7294 );
buf \U$892 ( \7720 , \7294 );
buf \U$893 ( \7721 , \7294 );
buf \U$894 ( \7722 , \7294 );
buf \U$895 ( \7723 , \7294 );
buf \U$896 ( \7724 , \7294 );
buf \U$897 ( \7725 , \7294 );
buf \U$898 ( \7726 , \7294 );
buf \U$899 ( \7727 , \7294 );
buf \U$900 ( \7728 , \7294 );
nor \U$901 ( \7729 , \7322 , \7282 , \7283 , \7284 , \7287 , \7291 , \7294 , \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 , \7712 , \7713 , \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 , \7722 , \7723 , \7724 , \7725 , \7726 , \7727 , \7728 );
and \U$902 ( \7730 , RIeb352c8_6904, \7729 );
or \U$903 ( \7731 , \7321 , \7352 , \7379 , \7406 , \7433 , \7460 , \7487 , \7514 , \7541 , \7568 , \7595 , \7622 , \7649 , \7676 , \7703 , \7730 );
buf \U$904 ( \7732 , \7294 );
not \U$905 ( \7733 , \7732 );
buf \U$906 ( \7734 , \7282 );
buf \U$907 ( \7735 , \7283 );
buf \U$908 ( \7736 , \7284 );
buf \U$909 ( \7737 , \7287 );
buf \U$910 ( \7738 , \7291 );
buf \U$911 ( \7739 , \7294 );
buf \U$912 ( \7740 , \7294 );
buf \U$913 ( \7741 , \7294 );
buf \U$914 ( \7742 , \7294 );
buf \U$915 ( \7743 , \7294 );
buf \U$916 ( \7744 , \7294 );
buf \U$917 ( \7745 , \7294 );
buf \U$918 ( \7746 , \7294 );
buf \U$919 ( \7747 , \7294 );
buf \U$920 ( \7748 , \7294 );
buf \U$921 ( \7749 , \7294 );
buf \U$922 ( \7750 , \7294 );
buf \U$923 ( \7751 , \7294 );
buf \U$924 ( \7752 , \7294 );
buf \U$925 ( \7753 , \7294 );
buf \U$926 ( \7754 , \7294 );
buf \U$927 ( \7755 , \7294 );
buf \U$928 ( \7756 , \7294 );
buf \U$929 ( \7757 , \7294 );
buf \U$930 ( \7758 , \7294 );
buf \U$931 ( \7759 , \7294 );
buf \U$932 ( \7760 , \7294 );
buf \U$933 ( \7761 , \7294 );
buf \U$934 ( \7762 , \7294 );
buf \U$935 ( \7763 , \7294 );
buf \U$936 ( \7764 , \7281 );
or \U$937 ( \7765 , \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 , \7742 , \7743 , \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 , \7752 , \7753 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 , \7762 , \7763 , \7764 );
nand \U$938 ( \7766 , \7733 , \7765 );
buf \U$939 ( \7767 , \7766 );
buf \U$940 ( \7768 , \7294 );
not \U$941 ( \7769 , \7768 );
buf \U$942 ( \7770 , \7291 );
buf \U$943 ( \7771 , \7294 );
buf \U$944 ( \7772 , \7294 );
buf \U$945 ( \7773 , \7294 );
buf \U$946 ( \7774 , \7294 );
buf \U$947 ( \7775 , \7294 );
buf \U$948 ( \7776 , \7294 );
buf \U$949 ( \7777 , \7294 );
buf \U$950 ( \7778 , \7294 );
buf \U$951 ( \7779 , \7294 );
buf \U$952 ( \7780 , \7294 );
buf \U$953 ( \7781 , \7294 );
buf \U$954 ( \7782 , \7294 );
buf \U$955 ( \7783 , \7294 );
buf \U$956 ( \7784 , \7294 );
buf \U$957 ( \7785 , \7294 );
buf \U$958 ( \7786 , \7294 );
buf \U$959 ( \7787 , \7294 );
buf \U$960 ( \7788 , \7294 );
buf \U$961 ( \7789 , \7294 );
buf \U$962 ( \7790 , \7294 );
buf \U$963 ( \7791 , \7294 );
buf \U$964 ( \7792 , \7294 );
buf \U$965 ( \7793 , \7294 );
buf \U$966 ( \7794 , \7294 );
buf \U$967 ( \7795 , \7294 );
buf \U$968 ( \7796 , \7287 );
buf \U$969 ( \7797 , \7281 );
buf \U$970 ( \7798 , \7282 );
buf \U$971 ( \7799 , \7283 );
buf \U$972 ( \7800 , \7284 );
or \U$973 ( \7801 , \7797 , \7798 , \7799 , \7800 );
and \U$974 ( \7802 , \7796 , \7801 );
or \U$975 ( \7803 , \7770 , \7771 , \7772 , \7773 , \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 , \7782 , \7783 , \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791 , \7792 , \7793 , \7794 , \7795 , \7802 );
and \U$976 ( \7804 , \7769 , \7803 );
buf \U$977 ( \7805 , \7804 );
or \U$978 ( \7806 , \7767 , \7805 );
_DC g3568 ( \7807_nG3568 , \7731 , \7806 );
not \U$979 ( \7808 , \7807_nG3568 );
buf \U$980 ( \7809 , RIb7b9608_246);
buf \U$981 ( \7810 , \7294 );
buf \U$982 ( \7811 , \7294 );
buf \U$983 ( \7812 , \7294 );
buf \U$984 ( \7813 , \7294 );
buf \U$985 ( \7814 , \7294 );
buf \U$986 ( \7815 , \7294 );
buf \U$987 ( \7816 , \7294 );
buf \U$988 ( \7817 , \7294 );
buf \U$989 ( \7818 , \7294 );
buf \U$990 ( \7819 , \7294 );
buf \U$991 ( \7820 , \7294 );
buf \U$992 ( \7821 , \7294 );
buf \U$993 ( \7822 , \7294 );
buf \U$994 ( \7823 , \7294 );
buf \U$995 ( \7824 , \7294 );
buf \U$996 ( \7825 , \7294 );
buf \U$997 ( \7826 , \7294 );
buf \U$998 ( \7827 , \7294 );
buf \U$999 ( \7828 , \7294 );
buf \U$1000 ( \7829 , \7294 );
buf \U$1001 ( \7830 , \7294 );
buf \U$1002 ( \7831 , \7294 );
buf \U$1003 ( \7832 , \7294 );
buf \U$1004 ( \7833 , \7294 );
buf \U$1005 ( \7834 , \7294 );
nor \U$1006 ( \7835 , \7281 , \7282 , \7283 , \7284 , \7288 , \7291 , \7294 , \7810 , \7811 , \7812 , \7813 , \7814 , \7815 , \7816 , \7817 , \7818 , \7819 , \7820 , \7821 , \7822 , \7823 , \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 , \7832 , \7833 , \7834 );
and \U$1007 ( \7836 , \7117 , \7835 );
buf \U$1008 ( \7837 , \7294 );
buf \U$1009 ( \7838 , \7294 );
buf \U$1010 ( \7839 , \7294 );
buf \U$1011 ( \7840 , \7294 );
buf \U$1012 ( \7841 , \7294 );
buf \U$1013 ( \7842 , \7294 );
buf \U$1014 ( \7843 , \7294 );
buf \U$1015 ( \7844 , \7294 );
buf \U$1016 ( \7845 , \7294 );
buf \U$1017 ( \7846 , \7294 );
buf \U$1018 ( \7847 , \7294 );
buf \U$1019 ( \7848 , \7294 );
buf \U$1020 ( \7849 , \7294 );
buf \U$1021 ( \7850 , \7294 );
buf \U$1022 ( \7851 , \7294 );
buf \U$1023 ( \7852 , \7294 );
buf \U$1024 ( \7853 , \7294 );
buf \U$1025 ( \7854 , \7294 );
buf \U$1026 ( \7855 , \7294 );
buf \U$1027 ( \7856 , \7294 );
buf \U$1028 ( \7857 , \7294 );
buf \U$1029 ( \7858 , \7294 );
buf \U$1030 ( \7859 , \7294 );
buf \U$1031 ( \7860 , \7294 );
buf \U$1032 ( \7861 , \7294 );
nor \U$1033 ( \7862 , \7322 , \7323 , \7324 , \7325 , \7287 , \7291 , \7294 , \7837 , \7838 , \7839 , \7840 , \7841 , \7842 , \7843 , \7844 , \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 , \7852 , \7853 , \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 );
and \U$1034 ( \7863 , \7119 , \7862 );
buf \U$1035 ( \7864 , RIe4340c0_5995);
buf \U$1036 ( \7865 , \7294 );
buf \U$1037 ( \7866 , \7294 );
buf \U$1038 ( \7867 , \7294 );
buf \U$1039 ( \7868 , \7294 );
buf \U$1040 ( \7869 , \7294 );
buf \U$1041 ( \7870 , \7294 );
buf \U$1042 ( \7871 , \7294 );
buf \U$1043 ( \7872 , \7294 );
buf \U$1044 ( \7873 , \7294 );
buf \U$1045 ( \7874 , \7294 );
buf \U$1046 ( \7875 , \7294 );
buf \U$1047 ( \7876 , \7294 );
buf \U$1048 ( \7877 , \7294 );
buf \U$1049 ( \7878 , \7294 );
buf \U$1050 ( \7879 , \7294 );
buf \U$1051 ( \7880 , \7294 );
buf \U$1052 ( \7881 , \7294 );
buf \U$1053 ( \7882 , \7294 );
buf \U$1054 ( \7883 , \7294 );
buf \U$1055 ( \7884 , \7294 );
buf \U$1056 ( \7885 , \7294 );
buf \U$1057 ( \7886 , \7294 );
buf \U$1058 ( \7887 , \7294 );
buf \U$1059 ( \7888 , \7294 );
buf \U$1060 ( \7889 , \7294 );
nor \U$1061 ( \7890 , \7281 , \7323 , \7324 , \7325 , \7287 , \7291 , \7294 , \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 , \7872 , \7873 , \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 , \7883 , \7884 , \7885 , \7886 , \7887 , \7888 , \7889 );
and \U$1062 ( \7891 , \7864 , \7890 );
buf \U$1063 ( \7892 , RIe26ce10_5604);
buf \U$1064 ( \7893 , \7294 );
buf \U$1065 ( \7894 , \7294 );
buf \U$1066 ( \7895 , \7294 );
buf \U$1067 ( \7896 , \7294 );
buf \U$1068 ( \7897 , \7294 );
buf \U$1069 ( \7898 , \7294 );
buf \U$1070 ( \7899 , \7294 );
buf \U$1071 ( \7900 , \7294 );
buf \U$1072 ( \7901 , \7294 );
buf \U$1073 ( \7902 , \7294 );
buf \U$1074 ( \7903 , \7294 );
buf \U$1075 ( \7904 , \7294 );
buf \U$1076 ( \7905 , \7294 );
buf \U$1077 ( \7906 , \7294 );
buf \U$1078 ( \7907 , \7294 );
buf \U$1079 ( \7908 , \7294 );
buf \U$1080 ( \7909 , \7294 );
buf \U$1081 ( \7910 , \7294 );
buf \U$1082 ( \7911 , \7294 );
buf \U$1083 ( \7912 , \7294 );
buf \U$1084 ( \7913 , \7294 );
buf \U$1085 ( \7914 , \7294 );
buf \U$1086 ( \7915 , \7294 );
buf \U$1087 ( \7916 , \7294 );
buf \U$1088 ( \7917 , \7294 );
nor \U$1089 ( \7918 , \7322 , \7282 , \7324 , \7325 , \7287 , \7291 , \7294 , \7893 , \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 , \7903 , \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 , \7913 , \7914 , \7915 , \7916 , \7917 );
and \U$1090 ( \7919 , \7892 , \7918 );
buf \U$1091 ( \7920 , RIe162368_5252);
buf \U$1092 ( \7921 , \7294 );
buf \U$1093 ( \7922 , \7294 );
buf \U$1094 ( \7923 , \7294 );
buf \U$1095 ( \7924 , \7294 );
buf \U$1096 ( \7925 , \7294 );
buf \U$1097 ( \7926 , \7294 );
buf \U$1098 ( \7927 , \7294 );
buf \U$1099 ( \7928 , \7294 );
buf \U$1100 ( \7929 , \7294 );
buf \U$1101 ( \7930 , \7294 );
buf \U$1102 ( \7931 , \7294 );
buf \U$1103 ( \7932 , \7294 );
buf \U$1104 ( \7933 , \7294 );
buf \U$1105 ( \7934 , \7294 );
buf \U$1106 ( \7935 , \7294 );
buf \U$1107 ( \7936 , \7294 );
buf \U$1108 ( \7937 , \7294 );
buf \U$1109 ( \7938 , \7294 );
buf \U$1110 ( \7939 , \7294 );
buf \U$1111 ( \7940 , \7294 );
buf \U$1112 ( \7941 , \7294 );
buf \U$1113 ( \7942 , \7294 );
buf \U$1114 ( \7943 , \7294 );
buf \U$1115 ( \7944 , \7294 );
buf \U$1116 ( \7945 , \7294 );
nor \U$1117 ( \7946 , \7281 , \7282 , \7324 , \7325 , \7287 , \7291 , \7294 , \7921 , \7922 , \7923 , \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 , \7933 , \7934 , \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 , \7942 , \7943 , \7944 , \7945 );
and \U$1118 ( \7947 , \7920 , \7946 );
buf \U$1119 ( \7948 , RIe0d89b0_4811);
buf \U$1120 ( \7949 , \7294 );
buf \U$1121 ( \7950 , \7294 );
buf \U$1122 ( \7951 , \7294 );
buf \U$1123 ( \7952 , \7294 );
buf \U$1124 ( \7953 , \7294 );
buf \U$1125 ( \7954 , \7294 );
buf \U$1126 ( \7955 , \7294 );
buf \U$1127 ( \7956 , \7294 );
buf \U$1128 ( \7957 , \7294 );
buf \U$1129 ( \7958 , \7294 );
buf \U$1130 ( \7959 , \7294 );
buf \U$1131 ( \7960 , \7294 );
buf \U$1132 ( \7961 , \7294 );
buf \U$1133 ( \7962 , \7294 );
buf \U$1134 ( \7963 , \7294 );
buf \U$1135 ( \7964 , \7294 );
buf \U$1136 ( \7965 , \7294 );
buf \U$1137 ( \7966 , \7294 );
buf \U$1138 ( \7967 , \7294 );
buf \U$1139 ( \7968 , \7294 );
buf \U$1140 ( \7969 , \7294 );
buf \U$1141 ( \7970 , \7294 );
buf \U$1142 ( \7971 , \7294 );
buf \U$1143 ( \7972 , \7294 );
buf \U$1144 ( \7973 , \7294 );
nor \U$1145 ( \7974 , \7322 , \7323 , \7283 , \7325 , \7287 , \7291 , \7294 , \7949 , \7950 , \7951 , \7952 , \7953 , \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 , \7963 , \7964 , \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 , \7972 , \7973 );
and \U$1146 ( \7975 , \7948 , \7974 );
buf \U$1147 ( \7976 , RIe00f6b0_4415);
buf \U$1148 ( \7977 , \7294 );
buf \U$1149 ( \7978 , \7294 );
buf \U$1150 ( \7979 , \7294 );
buf \U$1151 ( \7980 , \7294 );
buf \U$1152 ( \7981 , \7294 );
buf \U$1153 ( \7982 , \7294 );
buf \U$1154 ( \7983 , \7294 );
buf \U$1155 ( \7984 , \7294 );
buf \U$1156 ( \7985 , \7294 );
buf \U$1157 ( \7986 , \7294 );
buf \U$1158 ( \7987 , \7294 );
buf \U$1159 ( \7988 , \7294 );
buf \U$1160 ( \7989 , \7294 );
buf \U$1161 ( \7990 , \7294 );
buf \U$1162 ( \7991 , \7294 );
buf \U$1163 ( \7992 , \7294 );
buf \U$1164 ( \7993 , \7294 );
buf \U$1165 ( \7994 , \7294 );
buf \U$1166 ( \7995 , \7294 );
buf \U$1167 ( \7996 , \7294 );
buf \U$1168 ( \7997 , \7294 );
buf \U$1169 ( \7998 , \7294 );
buf \U$1170 ( \7999 , \7294 );
buf \U$1171 ( \8000 , \7294 );
buf \U$1172 ( \8001 , \7294 );
nor \U$1173 ( \8002 , \7281 , \7323 , \7283 , \7325 , \7287 , \7291 , \7294 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 , \7983 , \7984 , \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 , \7992 , \7993 , \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 );
and \U$1174 ( \8003 , \7976 , \8002 );
buf \U$1175 ( \8004 , RIde415d8_4022);
buf \U$1176 ( \8005 , \7294 );
buf \U$1177 ( \8006 , \7294 );
buf \U$1178 ( \8007 , \7294 );
buf \U$1179 ( \8008 , \7294 );
buf \U$1180 ( \8009 , \7294 );
buf \U$1181 ( \8010 , \7294 );
buf \U$1182 ( \8011 , \7294 );
buf \U$1183 ( \8012 , \7294 );
buf \U$1184 ( \8013 , \7294 );
buf \U$1185 ( \8014 , \7294 );
buf \U$1186 ( \8015 , \7294 );
buf \U$1187 ( \8016 , \7294 );
buf \U$1188 ( \8017 , \7294 );
buf \U$1189 ( \8018 , \7294 );
buf \U$1190 ( \8019 , \7294 );
buf \U$1191 ( \8020 , \7294 );
buf \U$1192 ( \8021 , \7294 );
buf \U$1193 ( \8022 , \7294 );
buf \U$1194 ( \8023 , \7294 );
buf \U$1195 ( \8024 , \7294 );
buf \U$1196 ( \8025 , \7294 );
buf \U$1197 ( \8026 , \7294 );
buf \U$1198 ( \8027 , \7294 );
buf \U$1199 ( \8028 , \7294 );
buf \U$1200 ( \8029 , \7294 );
nor \U$1201 ( \8030 , \7322 , \7282 , \7283 , \7325 , \7287 , \7291 , \7294 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 , \8013 , \8014 , \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 , \8022 , \8023 , \8024 , \8025 , \8026 , \8027 , \8028 , \8029 );
and \U$1202 ( \8031 , \8004 , \8030 );
buf \U$1203 ( \8032 , RIdd731d8_3637);
buf \U$1204 ( \8033 , \7294 );
buf \U$1205 ( \8034 , \7294 );
buf \U$1206 ( \8035 , \7294 );
buf \U$1207 ( \8036 , \7294 );
buf \U$1208 ( \8037 , \7294 );
buf \U$1209 ( \8038 , \7294 );
buf \U$1210 ( \8039 , \7294 );
buf \U$1211 ( \8040 , \7294 );
buf \U$1212 ( \8041 , \7294 );
buf \U$1213 ( \8042 , \7294 );
buf \U$1214 ( \8043 , \7294 );
buf \U$1215 ( \8044 , \7294 );
buf \U$1216 ( \8045 , \7294 );
buf \U$1217 ( \8046 , \7294 );
buf \U$1218 ( \8047 , \7294 );
buf \U$1219 ( \8048 , \7294 );
buf \U$1220 ( \8049 , \7294 );
buf \U$1221 ( \8050 , \7294 );
buf \U$1222 ( \8051 , \7294 );
buf \U$1223 ( \8052 , \7294 );
buf \U$1224 ( \8053 , \7294 );
buf \U$1225 ( \8054 , \7294 );
buf \U$1226 ( \8055 , \7294 );
buf \U$1227 ( \8056 , \7294 );
buf \U$1228 ( \8057 , \7294 );
nor \U$1229 ( \8058 , \7281 , \7282 , \7283 , \7325 , \7287 , \7291 , \7294 , \8033 , \8034 , \8035 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 , \8042 , \8043 , \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 , \8053 , \8054 , \8055 , \8056 , \8057 );
and \U$1230 ( \8059 , \8032 , \8058 );
buf \U$1231 ( \8060 , RIdba6bb8_3248);
buf \U$1232 ( \8061 , \7294 );
buf \U$1233 ( \8062 , \7294 );
buf \U$1234 ( \8063 , \7294 );
buf \U$1235 ( \8064 , \7294 );
buf \U$1236 ( \8065 , \7294 );
buf \U$1237 ( \8066 , \7294 );
buf \U$1238 ( \8067 , \7294 );
buf \U$1239 ( \8068 , \7294 );
buf \U$1240 ( \8069 , \7294 );
buf \U$1241 ( \8070 , \7294 );
buf \U$1242 ( \8071 , \7294 );
buf \U$1243 ( \8072 , \7294 );
buf \U$1244 ( \8073 , \7294 );
buf \U$1245 ( \8074 , \7294 );
buf \U$1246 ( \8075 , \7294 );
buf \U$1247 ( \8076 , \7294 );
buf \U$1248 ( \8077 , \7294 );
buf \U$1249 ( \8078 , \7294 );
buf \U$1250 ( \8079 , \7294 );
buf \U$1251 ( \8080 , \7294 );
buf \U$1252 ( \8081 , \7294 );
buf \U$1253 ( \8082 , \7294 );
buf \U$1254 ( \8083 , \7294 );
buf \U$1255 ( \8084 , \7294 );
buf \U$1256 ( \8085 , \7294 );
nor \U$1257 ( \8086 , \7322 , \7323 , \7324 , \7284 , \7287 , \7291 , \7294 , \8061 , \8062 , \8063 , \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 , \8072 , \8073 , \8074 , \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 , \8082 , \8083 , \8084 , \8085 );
and \U$1258 ( \8087 , \8060 , \8086 );
buf \U$1259 ( \8088 , RIdad7918_2858);
buf \U$1260 ( \8089 , \7294 );
buf \U$1261 ( \8090 , \7294 );
buf \U$1262 ( \8091 , \7294 );
buf \U$1263 ( \8092 , \7294 );
buf \U$1264 ( \8093 , \7294 );
buf \U$1265 ( \8094 , \7294 );
buf \U$1266 ( \8095 , \7294 );
buf \U$1267 ( \8096 , \7294 );
buf \U$1268 ( \8097 , \7294 );
buf \U$1269 ( \8098 , \7294 );
buf \U$1270 ( \8099 , \7294 );
buf \U$1271 ( \8100 , \7294 );
buf \U$1272 ( \8101 , \7294 );
buf \U$1273 ( \8102 , \7294 );
buf \U$1274 ( \8103 , \7294 );
buf \U$1275 ( \8104 , \7294 );
buf \U$1276 ( \8105 , \7294 );
buf \U$1277 ( \8106 , \7294 );
buf \U$1278 ( \8107 , \7294 );
buf \U$1279 ( \8108 , \7294 );
buf \U$1280 ( \8109 , \7294 );
buf \U$1281 ( \8110 , \7294 );
buf \U$1282 ( \8111 , \7294 );
buf \U$1283 ( \8112 , \7294 );
buf \U$1284 ( \8113 , \7294 );
nor \U$1285 ( \8114 , \7281 , \7323 , \7324 , \7284 , \7287 , \7291 , \7294 , \8089 , \8090 , \8091 , \8092 , \8093 , \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 , \8103 , \8104 , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 , \8112 , \8113 );
and \U$1286 ( \8115 , \8088 , \8114 );
buf \U$1287 ( \8116 , RIda15da0_2441);
buf \U$1288 ( \8117 , \7294 );
buf \U$1289 ( \8118 , \7294 );
buf \U$1290 ( \8119 , \7294 );
buf \U$1291 ( \8120 , \7294 );
buf \U$1292 ( \8121 , \7294 );
buf \U$1293 ( \8122 , \7294 );
buf \U$1294 ( \8123 , \7294 );
buf \U$1295 ( \8124 , \7294 );
buf \U$1296 ( \8125 , \7294 );
buf \U$1297 ( \8126 , \7294 );
buf \U$1298 ( \8127 , \7294 );
buf \U$1299 ( \8128 , \7294 );
buf \U$1300 ( \8129 , \7294 );
buf \U$1301 ( \8130 , \7294 );
buf \U$1302 ( \8131 , \7294 );
buf \U$1303 ( \8132 , \7294 );
buf \U$1304 ( \8133 , \7294 );
buf \U$1305 ( \8134 , \7294 );
buf \U$1306 ( \8135 , \7294 );
buf \U$1307 ( \8136 , \7294 );
buf \U$1308 ( \8137 , \7294 );
buf \U$1309 ( \8138 , \7294 );
buf \U$1310 ( \8139 , \7294 );
buf \U$1311 ( \8140 , \7294 );
buf \U$1312 ( \8141 , \7294 );
nor \U$1313 ( \8142 , \7322 , \7282 , \7324 , \7284 , \7287 , \7291 , \7294 , \8117 , \8118 , \8119 , \8120 , \8121 , \8122 , \8123 , \8124 , \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 , \8132 , \8133 , \8134 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 );
and \U$1314 ( \8143 , \8116 , \8142 );
buf \U$1315 ( \8144 , RId95c8b0_2053);
buf \U$1316 ( \8145 , \7294 );
buf \U$1317 ( \8146 , \7294 );
buf \U$1318 ( \8147 , \7294 );
buf \U$1319 ( \8148 , \7294 );
buf \U$1320 ( \8149 , \7294 );
buf \U$1321 ( \8150 , \7294 );
buf \U$1322 ( \8151 , \7294 );
buf \U$1323 ( \8152 , \7294 );
buf \U$1324 ( \8153 , \7294 );
buf \U$1325 ( \8154 , \7294 );
buf \U$1326 ( \8155 , \7294 );
buf \U$1327 ( \8156 , \7294 );
buf \U$1328 ( \8157 , \7294 );
buf \U$1329 ( \8158 , \7294 );
buf \U$1330 ( \8159 , \7294 );
buf \U$1331 ( \8160 , \7294 );
buf \U$1332 ( \8161 , \7294 );
buf \U$1333 ( \8162 , \7294 );
buf \U$1334 ( \8163 , \7294 );
buf \U$1335 ( \8164 , \7294 );
buf \U$1336 ( \8165 , \7294 );
buf \U$1337 ( \8166 , \7294 );
buf \U$1338 ( \8167 , \7294 );
buf \U$1339 ( \8168 , \7294 );
buf \U$1340 ( \8169 , \7294 );
nor \U$1341 ( \8170 , \7281 , \7282 , \7324 , \7284 , \7287 , \7291 , \7294 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 , \8152 , \8153 , \8154 , \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 , \8162 , \8163 , \8164 , \8165 , \8166 , \8167 , \8168 , \8169 );
and \U$1342 ( \8171 , \8144 , \8170 );
buf \U$1343 ( \8172 , RId88c728_1664);
buf \U$1344 ( \8173 , \7294 );
buf \U$1345 ( \8174 , \7294 );
buf \U$1346 ( \8175 , \7294 );
buf \U$1347 ( \8176 , \7294 );
buf \U$1348 ( \8177 , \7294 );
buf \U$1349 ( \8178 , \7294 );
buf \U$1350 ( \8179 , \7294 );
buf \U$1351 ( \8180 , \7294 );
buf \U$1352 ( \8181 , \7294 );
buf \U$1353 ( \8182 , \7294 );
buf \U$1354 ( \8183 , \7294 );
buf \U$1355 ( \8184 , \7294 );
buf \U$1356 ( \8185 , \7294 );
buf \U$1357 ( \8186 , \7294 );
buf \U$1358 ( \8187 , \7294 );
buf \U$1359 ( \8188 , \7294 );
buf \U$1360 ( \8189 , \7294 );
buf \U$1361 ( \8190 , \7294 );
buf \U$1362 ( \8191 , \7294 );
buf \U$1363 ( \8192 , \7294 );
buf \U$1364 ( \8193 , \7294 );
buf \U$1365 ( \8194 , \7294 );
buf \U$1366 ( \8195 , \7294 );
buf \U$1367 ( \8196 , \7294 );
buf \U$1368 ( \8197 , \7294 );
nor \U$1369 ( \8198 , \7322 , \7323 , \7283 , \7284 , \7287 , \7291 , \7294 , \8173 , \8174 , \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 , \8182 , \8183 , \8184 , \8185 , \8186 , \8187 , \8188 , \8189 , \8190 , \8191 , \8192 , \8193 , \8194 , \8195 , \8196 , \8197 );
and \U$1370 ( \8199 , \8172 , \8198 );
buf \U$1371 ( \8200 , RId7c3590_1267);
buf \U$1372 ( \8201 , \7294 );
buf \U$1373 ( \8202 , \7294 );
buf \U$1374 ( \8203 , \7294 );
buf \U$1375 ( \8204 , \7294 );
buf \U$1376 ( \8205 , \7294 );
buf \U$1377 ( \8206 , \7294 );
buf \U$1378 ( \8207 , \7294 );
buf \U$1379 ( \8208 , \7294 );
buf \U$1380 ( \8209 , \7294 );
buf \U$1381 ( \8210 , \7294 );
buf \U$1382 ( \8211 , \7294 );
buf \U$1383 ( \8212 , \7294 );
buf \U$1384 ( \8213 , \7294 );
buf \U$1385 ( \8214 , \7294 );
buf \U$1386 ( \8215 , \7294 );
buf \U$1387 ( \8216 , \7294 );
buf \U$1388 ( \8217 , \7294 );
buf \U$1389 ( \8218 , \7294 );
buf \U$1390 ( \8219 , \7294 );
buf \U$1391 ( \8220 , \7294 );
buf \U$1392 ( \8221 , \7294 );
buf \U$1393 ( \8222 , \7294 );
buf \U$1394 ( \8223 , \7294 );
buf \U$1395 ( \8224 , \7294 );
buf \U$1396 ( \8225 , \7294 );
nor \U$1397 ( \8226 , \7281 , \7323 , \7283 , \7284 , \7287 , \7291 , \7294 , \8201 , \8202 , \8203 , \8204 , \8205 , \8206 , \8207 , \8208 , \8209 , \8210 , \8211 , \8212 , \8213 , \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 , \8222 , \8223 , \8224 , \8225 );
and \U$1398 ( \8227 , \8200 , \8226 );
buf \U$1399 ( \8228 , RId6f73b0_878);
buf \U$1400 ( \8229 , \7294 );
buf \U$1401 ( \8230 , \7294 );
buf \U$1402 ( \8231 , \7294 );
buf \U$1403 ( \8232 , \7294 );
buf \U$1404 ( \8233 , \7294 );
buf \U$1405 ( \8234 , \7294 );
buf \U$1406 ( \8235 , \7294 );
buf \U$1407 ( \8236 , \7294 );
buf \U$1408 ( \8237 , \7294 );
buf \U$1409 ( \8238 , \7294 );
buf \U$1410 ( \8239 , \7294 );
buf \U$1411 ( \8240 , \7294 );
buf \U$1412 ( \8241 , \7294 );
buf \U$1413 ( \8242 , \7294 );
buf \U$1414 ( \8243 , \7294 );
buf \U$1415 ( \8244 , \7294 );
buf \U$1416 ( \8245 , \7294 );
buf \U$1417 ( \8246 , \7294 );
buf \U$1418 ( \8247 , \7294 );
buf \U$1419 ( \8248 , \7294 );
buf \U$1420 ( \8249 , \7294 );
buf \U$1421 ( \8250 , \7294 );
buf \U$1422 ( \8251 , \7294 );
buf \U$1423 ( \8252 , \7294 );
buf \U$1424 ( \8253 , \7294 );
nor \U$1425 ( \8254 , \7322 , \7282 , \7283 , \7284 , \7287 , \7291 , \7294 , \8229 , \8230 , \8231 , \8232 , \8233 , \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 , \8242 , \8243 , \8244 , \8245 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 , \8252 , \8253 );
and \U$1426 ( \8255 , \8228 , \8254 );
or \U$1427 ( \8256 , \7836 , \7863 , \7891 , \7919 , \7947 , \7975 , \8003 , \8031 , \8059 , \8087 , \8115 , \8143 , \8171 , \8199 , \8227 , \8255 );
buf \U$1428 ( \8257 , \7294 );
not \U$1429 ( \8258 , \8257 );
buf \U$1430 ( \8259 , \7282 );
buf \U$1431 ( \8260 , \7283 );
buf \U$1432 ( \8261 , \7284 );
buf \U$1433 ( \8262 , \7287 );
buf \U$1434 ( \8263 , \7291 );
buf \U$1435 ( \8264 , \7294 );
buf \U$1436 ( \8265 , \7294 );
buf \U$1437 ( \8266 , \7294 );
buf \U$1438 ( \8267 , \7294 );
buf \U$1439 ( \8268 , \7294 );
buf \U$1440 ( \8269 , \7294 );
buf \U$1441 ( \8270 , \7294 );
buf \U$1442 ( \8271 , \7294 );
buf \U$1443 ( \8272 , \7294 );
buf \U$1444 ( \8273 , \7294 );
buf \U$1445 ( \8274 , \7294 );
buf \U$1446 ( \8275 , \7294 );
buf \U$1447 ( \8276 , \7294 );
buf \U$1448 ( \8277 , \7294 );
buf \U$1449 ( \8278 , \7294 );
buf \U$1450 ( \8279 , \7294 );
buf \U$1451 ( \8280 , \7294 );
buf \U$1452 ( \8281 , \7294 );
buf \U$1453 ( \8282 , \7294 );
buf \U$1454 ( \8283 , \7294 );
buf \U$1455 ( \8284 , \7294 );
buf \U$1456 ( \8285 , \7294 );
buf \U$1457 ( \8286 , \7294 );
buf \U$1458 ( \8287 , \7294 );
buf \U$1459 ( \8288 , \7294 );
buf \U$1460 ( \8289 , \7281 );
or \U$1461 ( \8290 , \8259 , \8260 , \8261 , \8262 , \8263 , \8264 , \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271 , \8272 , \8273 , \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 , \8282 , \8283 , \8284 , \8285 , \8286 , \8287 , \8288 , \8289 );
nand \U$1462 ( \8291 , \8258 , \8290 );
buf \U$1463 ( \8292 , \8291 );
buf \U$1464 ( \8293 , \7294 );
not \U$1465 ( \8294 , \8293 );
buf \U$1466 ( \8295 , \7291 );
buf \U$1467 ( \8296 , \7294 );
buf \U$1468 ( \8297 , \7294 );
buf \U$1469 ( \8298 , \7294 );
buf \U$1470 ( \8299 , \7294 );
buf \U$1471 ( \8300 , \7294 );
buf \U$1472 ( \8301 , \7294 );
buf \U$1473 ( \8302 , \7294 );
buf \U$1474 ( \8303 , \7294 );
buf \U$1475 ( \8304 , \7294 );
buf \U$1476 ( \8305 , \7294 );
buf \U$1477 ( \8306 , \7294 );
buf \U$1478 ( \8307 , \7294 );
buf \U$1479 ( \8308 , \7294 );
buf \U$1480 ( \8309 , \7294 );
buf \U$1481 ( \8310 , \7294 );
buf \U$1482 ( \8311 , \7294 );
buf \U$1483 ( \8312 , \7294 );
buf \U$1484 ( \8313 , \7294 );
buf \U$1485 ( \8314 , \7294 );
buf \U$1486 ( \8315 , \7294 );
buf \U$1487 ( \8316 , \7294 );
buf \U$1488 ( \8317 , \7294 );
buf \U$1489 ( \8318 , \7294 );
buf \U$1490 ( \8319 , \7294 );
buf \U$1491 ( \8320 , \7294 );
buf \U$1492 ( \8321 , \7287 );
buf \U$1493 ( \8322 , \7281 );
buf \U$1494 ( \8323 , \7282 );
buf \U$1495 ( \8324 , \7283 );
buf \U$1496 ( \8325 , \7284 );
or \U$1497 ( \8326 , \8322 , \8323 , \8324 , \8325 );
and \U$1498 ( \8327 , \8321 , \8326 );
or \U$1499 ( \8328 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 , \8302 , \8303 , \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 , \8312 , \8313 , \8314 , \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8327 );
and \U$1500 ( \8329 , \8294 , \8328 );
buf \U$1501 ( \8330 , \8329 );
or \U$1502 ( \8331 , \8292 , \8330 );
_DC g3775 ( \8332_nG3775 , \8256 , \8331 );
buf \U$1503 ( \8333 , \8332_nG3775 );
xor \U$1504 ( \8334 , \7809 , \8333 );
buf \U$1505 ( \8335 , RIb7b9590_247);
and \U$1506 ( \8336 , \7126 , \7835 );
and \U$1507 ( \8337 , \7128 , \7862 );
buf \U$1508 ( \8338 , RIe4333a0_5996);
and \U$1509 ( \8339 , \8338 , \7890 );
buf \U$1510 ( \8340 , RIe26c000_5605);
and \U$1511 ( \8341 , \8340 , \7918 );
buf \U$1512 ( \8342 , RIe1658d8_5248);
and \U$1513 ( \8343 , \8342 , \7946 );
buf \U$1514 ( \8344 , RIe0d7d08_4812);
and \U$1515 ( \8345 , \8344 , \7974 );
buf \U$1516 ( \8346 , RIe00e918_4416);
and \U$1517 ( \8347 , \8346 , \8002 );
buf \U$1518 ( \8348 , RIde408b8_4023);
and \U$1519 ( \8349 , \8348 , \8030 );
buf \U$1520 ( \8350 , RIdc72420_3638);
and \U$1521 ( \8351 , \8350 , \8058 );
buf \U$1522 ( \8352 , RIdba5e98_3249);
and \U$1523 ( \8353 , \8352 , \8086 );
buf \U$1524 ( \8354 , RIdad6b80_2859);
and \U$1525 ( \8355 , \8354 , \8114 );
buf \U$1526 ( \8356 , RIda150f8_2442);
and \U$1527 ( \8357 , \8356 , \8142 );
buf \U$1528 ( \8358 , RId95bcf8_2054);
and \U$1529 ( \8359 , \8358 , \8170 );
buf \U$1530 ( \8360 , RId88bbe8_1665);
and \U$1531 ( \8361 , \8360 , \8198 );
buf \U$1532 ( \8362 , RId7c2870_1268);
and \U$1533 ( \8363 , \8362 , \8226 );
buf \U$1534 ( \8364 , RId6f68e8_879);
and \U$1535 ( \8365 , \8364 , \8254 );
or \U$1536 ( \8366 , \8336 , \8337 , \8339 , \8341 , \8343 , \8345 , \8347 , \8349 , \8351 , \8353 , \8355 , \8357 , \8359 , \8361 , \8363 , \8365 );
_DC g3798 ( \8367_nG3798 , \8366 , \8331 );
buf \U$1537 ( \8368 , \8367_nG3798 );
xor \U$1538 ( \8369 , \8335 , \8368 );
or \U$1539 ( \8370 , \8334 , \8369 );
buf \U$1540 ( \8371 , RIb7b9518_248);
and \U$1541 ( \8372 , \7136 , \7835 );
and \U$1542 ( \8373 , \7138 , \7862 );
buf \U$1543 ( \8374 , RIe4326f8_5997);
and \U$1544 ( \8375 , \8374 , \7890 );
buf \U$1545 ( \8376 , RIe26b2e0_5606);
and \U$1546 ( \8377 , \8376 , \7918 );
buf \U$1547 ( \8378 , RIe164b40_5249);
and \U$1548 ( \8379 , \8378 , \7946 );
buf \U$1549 ( \8380 , RIe0d6fe8_4813);
and \U$1550 ( \8381 , \8380 , \7974 );
buf \U$1551 ( \8382 , RIe00db80_4417);
and \U$1552 ( \8383 , \8382 , \8002 );
buf \U$1553 ( \8384 , RIde3fb20_4024);
and \U$1554 ( \8385 , \8384 , \8030 );
buf \U$1555 ( \8386 , RIdc71610_3639);
and \U$1556 ( \8387 , \8386 , \8058 );
buf \U$1557 ( \8388 , RIdba51f0_3250);
and \U$1558 ( \8389 , \8388 , \8086 );
buf \U$1559 ( \8390 , RIdad5d70_2860);
and \U$1560 ( \8391 , \8390 , \8114 );
buf \U$1561 ( \8392 , RIda143d8_2443);
and \U$1562 ( \8393 , \8392 , \8142 );
buf \U$1563 ( \8394 , RId95b1b8_2055);
and \U$1564 ( \8395 , \8394 , \8170 );
buf \U$1565 ( \8396 , RId88b030_1666);
and \U$1566 ( \8397 , \8396 , \8198 );
buf \U$1567 ( \8398 , RId7c1b50_1269);
and \U$1568 ( \8399 , \8398 , \8226 );
buf \U$1569 ( \8400 , RId6f5cb8_880);
and \U$1570 ( \8401 , \8400 , \8254 );
or \U$1571 ( \8402 , \8372 , \8373 , \8375 , \8377 , \8379 , \8381 , \8383 , \8385 , \8387 , \8389 , \8391 , \8393 , \8395 , \8397 , \8399 , \8401 );
_DC g37bc ( \8403_nG37bc , \8402 , \8331 );
buf \U$1572 ( \8404 , \8403_nG37bc );
xor \U$1573 ( \8405 , \8371 , \8404 );
or \U$1574 ( \8406 , \8370 , \8405 );
buf \U$1575 ( \8407 , RIb7b94a0_249);
and \U$1576 ( \8408 , \7146 , \7835 );
and \U$1577 ( \8409 , \7148 , \7862 );
buf \U$1578 ( \8410 , RIe431ac8_5998);
and \U$1579 ( \8411 , \8410 , \7890 );
buf \U$1580 ( \8412 , RIe26a7a0_5607);
and \U$1581 ( \8413 , \8412 , \7918 );
buf \U$1582 ( \8414 , RIe1615d0_5253);
and \U$1583 ( \8415 , \8414 , \7946 );
buf \U$1584 ( \8416 , RIe0d62c8_4814);
and \U$1585 ( \8417 , \8416 , \7974 );
buf \U$1586 ( \8418 , RIe00ce60_4418);
and \U$1587 ( \8419 , \8418 , \8002 );
buf \U$1588 ( \8420 , RIde3ed88_4025);
and \U$1589 ( \8421 , \8420 , \8030 );
buf \U$1590 ( \8422 , RIdc70800_3640);
and \U$1591 ( \8423 , \8422 , \8058 );
buf \U$1592 ( \8424 , RIdba4548_3251);
and \U$1593 ( \8425 , \8424 , \8086 );
buf \U$1594 ( \8426 , RIdaebc88_2833);
and \U$1595 ( \8427 , \8426 , \8114 );
buf \U$1596 ( \8428 , RIda13640_2444);
and \U$1597 ( \8429 , \8428 , \8142 );
buf \U$1598 ( \8430 , RId95a600_2056);
and \U$1599 ( \8431 , \8430 , \8170 );
buf \U$1600 ( \8432 , RId88a478_1667);
and \U$1601 ( \8433 , \8432 , \8198 );
buf \U$1602 ( \8434 , RId7c0e30_1270);
and \U$1603 ( \8435 , \8434 , \8226 );
buf \U$1604 ( \8436 , RId6f5100_881);
and \U$1605 ( \8437 , \8436 , \8254 );
or \U$1606 ( \8438 , \8408 , \8409 , \8411 , \8413 , \8415 , \8417 , \8419 , \8421 , \8423 , \8425 , \8427 , \8429 , \8431 , \8433 , \8435 , \8437 );
_DC g37e0 ( \8439_nG37e0 , \8438 , \8331 );
buf \U$1607 ( \8440 , \8439_nG37e0 );
xor \U$1608 ( \8441 , \8407 , \8440 );
or \U$1609 ( \8442 , \8406 , \8441 );
buf \U$1610 ( \8443 , RIb7b9428_250);
and \U$1611 ( \8444 , \7156 , \7835 );
and \U$1612 ( \8445 , \7158 , \7862 );
buf \U$1613 ( \8446 , RIe430e20_5999);
and \U$1614 ( \8447 , \8446 , \7890 );
buf \U$1615 ( \8448 , RIe269c60_5608);
and \U$1616 ( \8449 , \8448 , \7918 );
buf \U$1617 ( \8450 , RIe163088_5251);
and \U$1618 ( \8451 , \8450 , \7946 );
buf \U$1619 ( \8452 , RIe0d55a8_4815);
and \U$1620 ( \8453 , \8452 , \7974 );
buf \U$1621 ( \8454 , RIe00c0c8_4419);
and \U$1622 ( \8455 , \8454 , \8002 );
buf \U$1623 ( \8456 , RIde3df00_4026);
and \U$1624 ( \8457 , \8456 , \8030 );
buf \U$1625 ( \8458 , RIdc6f9f0_3641);
and \U$1626 ( \8459 , \8458 , \8058 );
buf \U$1627 ( \8460 , RIdba3828_3252);
and \U$1628 ( \8461 , \8460 , \8086 );
buf \U$1629 ( \8462 , RIdaeb0d0_2834);
and \U$1630 ( \8463 , \8462 , \8114 );
buf \U$1631 ( \8464 , RIda12920_2445);
and \U$1632 ( \8465 , \8464 , \8142 );
buf \U$1633 ( \8466 , RId959a48_2057);
and \U$1634 ( \8467 , \8466 , \8170 );
buf \U$1635 ( \8468 , RId889938_1668);
and \U$1636 ( \8469 , \8468 , \8198 );
buf \U$1637 ( \8470 , RId7c0110_1271);
and \U$1638 ( \8471 , \8470 , \8226 );
buf \U$1639 ( \8472 , RId6f4638_882);
and \U$1640 ( \8473 , \8472 , \8254 );
or \U$1641 ( \8474 , \8444 , \8445 , \8447 , \8449 , \8451 , \8453 , \8455 , \8457 , \8459 , \8461 , \8463 , \8465 , \8467 , \8469 , \8471 , \8473 );
_DC g3804 ( \8475_nG3804 , \8474 , \8331 );
buf \U$1642 ( \8476 , \8475_nG3804 );
xor \U$1643 ( \8477 , \8443 , \8476 );
or \U$1644 ( \8478 , \8442 , \8477 );
buf \U$1645 ( \8479 , RIb7b93b0_251);
and \U$1646 ( \8480 , \7166 , \7835 );
and \U$1647 ( \8481 , \7168 , \7862 );
buf \U$1648 ( \8482 , RIe4301f0_6000);
and \U$1649 ( \8483 , \8482 , \7890 );
buf \U$1650 ( \8484 , RIe269120_5609);
and \U$1651 ( \8485 , \8484 , \7918 );
buf \U$1652 ( \8486 , RIe160838_5254);
and \U$1653 ( \8487 , \8486 , \7946 );
buf \U$1654 ( \8488 , RIe0d49f0_4816);
and \U$1655 ( \8489 , \8488 , \7974 );
buf \U$1656 ( \8490 , RIe00b330_4420);
and \U$1657 ( \8491 , \8490 , \8002 );
buf \U$1658 ( \8492 , RIde3d1e0_4027);
and \U$1659 ( \8493 , \8492 , \8030 );
buf \U$1660 ( \8494 , RIdc6ed48_3642);
and \U$1661 ( \8495 , \8494 , \8058 );
buf \U$1662 ( \8496 , RIdbb8138_3227);
and \U$1663 ( \8497 , \8496 , \8086 );
buf \U$1664 ( \8498 , RIdaea590_2835);
and \U$1665 ( \8499 , \8498 , \8114 );
buf \U$1666 ( \8500 , RIda11c00_2446);
and \U$1667 ( \8501 , \8500 , \8142 );
buf \U$1668 ( \8502 , RId958f08_2058);
and \U$1669 ( \8503 , \8502 , \8170 );
buf \U$1670 ( \8504 , RId888d80_1669);
and \U$1671 ( \8505 , \8504 , \8198 );
buf \U$1672 ( \8506 , RId7bf4e0_1272);
and \U$1673 ( \8507 , \8506 , \8226 );
buf \U$1674 ( \8508 , RId6f3a80_883);
and \U$1675 ( \8509 , \8508 , \8254 );
or \U$1676 ( \8510 , \8480 , \8481 , \8483 , \8485 , \8487 , \8489 , \8491 , \8493 , \8495 , \8497 , \8499 , \8501 , \8503 , \8505 , \8507 , \8509 );
_DC g3828 ( \8511_nG3828 , \8510 , \8331 );
buf \U$1677 ( \8512 , \8511_nG3828 );
xor \U$1678 ( \8513 , \8479 , \8512 );
or \U$1679 ( \8514 , \8478 , \8513 );
buf \U$1680 ( \8515 , RIb7af720_252);
and \U$1681 ( \8516 , \7176 , \7835 );
and \U$1682 ( \8517 , \7178 , \7862 );
buf \U$1683 ( \8518 , RIe42f4d0_6001);
and \U$1684 ( \8519 , \8518 , \7890 );
buf \U$1685 ( \8520 , RIe268568_5610);
and \U$1686 ( \8521 , \8520 , \7918 );
buf \U$1687 ( \8522 , RIe172718_5244);
and \U$1688 ( \8523 , \8522 , \7946 );
buf \U$1689 ( \8524 , RIe0d3dc0_4817);
and \U$1690 ( \8525 , \8524 , \7974 );
buf \U$1691 ( \8526 , RIe00a598_4421);
and \U$1692 ( \8527 , \8526 , \8002 );
buf \U$1693 ( \8528 , RIde3c448_4028);
and \U$1694 ( \8529 , \8528 , \8030 );
buf \U$1695 ( \8530 , RIdc6e280_3643);
and \U$1696 ( \8531 , \8530 , \8058 );
buf \U$1697 ( \8532 , RIdbb7328_3228);
and \U$1698 ( \8533 , \8532 , \8086 );
buf \U$1699 ( \8534 , RIdae97f8_2836);
and \U$1700 ( \8535 , \8534 , \8114 );
buf \U$1701 ( \8536 , RIda10df0_2447);
and \U$1702 ( \8537 , \8536 , \8142 );
buf \U$1703 ( \8538 , RId9582d8_2059);
and \U$1704 ( \8539 , \8538 , \8170 );
buf \U$1705 ( \8540 , RId888240_1670);
and \U$1706 ( \8541 , \8540 , \8198 );
buf \U$1707 ( \8542 , RId7be838_1273);
and \U$1708 ( \8543 , \8542 , \8226 );
buf \U$1709 ( \8544 , RId7064a0_859);
and \U$1710 ( \8545 , \8544 , \8254 );
or \U$1711 ( \8546 , \8516 , \8517 , \8519 , \8521 , \8523 , \8525 , \8527 , \8529 , \8531 , \8533 , \8535 , \8537 , \8539 , \8541 , \8543 , \8545 );
_DC g384c ( \8547_nG384c , \8546 , \8331 );
buf \U$1712 ( \8548 , \8547_nG384c );
xor \U$1713 ( \8549 , \8515 , \8548 );
or \U$1714 ( \8550 , \8514 , \8549 );
buf \U$1715 ( \8551 , RIb7af6a8_253);
and \U$1716 ( \8552 , \7186 , \7835 );
and \U$1717 ( \8553 , \7188 , \7862 );
buf \U$1718 ( \8554 , RIe42e8a0_6002);
and \U$1719 ( \8555 , \8554 , \7890 );
buf \U$1720 ( \8556 , RIe2679b0_5611);
and \U$1721 ( \8557 , \8556 , \7918 );
buf \U$1722 ( \8558 , RIe163e20_5250);
and \U$1723 ( \8559 , \8558 , \7946 );
buf \U$1724 ( \8560 , RIe0d2e48_4818);
and \U$1725 ( \8561 , \8560 , \7974 );
buf \U$1726 ( \8562 , RIe009710_4422);
and \U$1727 ( \8563 , \8562 , \8002 );
buf \U$1728 ( \8564 , RIde3b728_4029);
and \U$1729 ( \8565 , \8564 , \8030 );
buf \U$1730 ( \8566 , RIdc6d740_3644);
and \U$1731 ( \8567 , \8566 , \8058 );
buf \U$1732 ( \8568 , RIdbb6518_3229);
and \U$1733 ( \8569 , \8568 , \8086 );
buf \U$1734 ( \8570 , RIdae8a60_2837);
and \U$1735 ( \8571 , \8570 , \8114 );
buf \U$1736 ( \8572 , RIda101c0_2448);
and \U$1737 ( \8573 , \8572 , \8142 );
buf \U$1738 ( \8574 , RId957720_2060);
and \U$1739 ( \8575 , \8574 , \8170 );
buf \U$1740 ( \8576 , RId89b638_1645);
and \U$1741 ( \8577 , \8576 , \8198 );
buf \U$1742 ( \8578 , RId7d2338_1248);
and \U$1743 ( \8579 , \8578 , \8226 );
buf \U$1744 ( \8580 , RId705780_860);
and \U$1745 ( \8581 , \8580 , \8254 );
or \U$1746 ( \8582 , \8552 , \8553 , \8555 , \8557 , \8559 , \8561 , \8563 , \8565 , \8567 , \8569 , \8571 , \8573 , \8575 , \8577 , \8579 , \8581 );
_DC g3870 ( \8583_nG3870 , \8582 , \8331 );
buf \U$1747 ( \8584 , \8583_nG3870 );
xor \U$1748 ( \8585 , \8551 , \8584 );
or \U$1749 ( \8586 , \8550 , \8585 );
not \U$1750 ( \8587 , \8586 );
buf \U$1751 ( \8588 , \8587 );
and \U$1752 ( \8589 , \7808 , \8588 );
buf \U$1753 ( \8590 , RIb7af630_254);
buf \U$1754 ( \8591 , \7294 );
buf \U$1755 ( \8592 , \7294 );
buf \U$1756 ( \8593 , \7294 );
buf \U$1757 ( \8594 , \7294 );
buf \U$1758 ( \8595 , \7294 );
buf \U$1759 ( \8596 , \7294 );
buf \U$1760 ( \8597 , \7294 );
buf \U$1761 ( \8598 , \7294 );
buf \U$1762 ( \8599 , \7294 );
buf \U$1763 ( \8600 , \7294 );
buf \U$1764 ( \8601 , \7294 );
buf \U$1765 ( \8602 , \7294 );
buf \U$1766 ( \8603 , \7294 );
buf \U$1767 ( \8604 , \7294 );
buf \U$1768 ( \8605 , \7294 );
buf \U$1769 ( \8606 , \7294 );
buf \U$1770 ( \8607 , \7294 );
buf \U$1771 ( \8608 , \7294 );
buf \U$1772 ( \8609 , \7294 );
buf \U$1773 ( \8610 , \7294 );
buf \U$1774 ( \8611 , \7294 );
buf \U$1775 ( \8612 , \7294 );
buf \U$1776 ( \8613 , \7294 );
buf \U$1777 ( \8614 , \7294 );
buf \U$1778 ( \8615 , \7294 );
nor \U$1779 ( \8616 , \7281 , \7282 , \7283 , \7284 , \7288 , \7291 , \7294 , \8591 , \8592 , \8593 , \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 , \8612 , \8613 , \8614 , \8615 );
and \U$1780 ( \8617 , \7198 , \8616 );
buf \U$1781 ( \8618 , \7294 );
buf \U$1782 ( \8619 , \7294 );
buf \U$1783 ( \8620 , \7294 );
buf \U$1784 ( \8621 , \7294 );
buf \U$1785 ( \8622 , \7294 );
buf \U$1786 ( \8623 , \7294 );
buf \U$1787 ( \8624 , \7294 );
buf \U$1788 ( \8625 , \7294 );
buf \U$1789 ( \8626 , \7294 );
buf \U$1790 ( \8627 , \7294 );
buf \U$1791 ( \8628 , \7294 );
buf \U$1792 ( \8629 , \7294 );
buf \U$1793 ( \8630 , \7294 );
buf \U$1794 ( \8631 , \7294 );
buf \U$1795 ( \8632 , \7294 );
buf \U$1796 ( \8633 , \7294 );
buf \U$1797 ( \8634 , \7294 );
buf \U$1798 ( \8635 , \7294 );
buf \U$1799 ( \8636 , \7294 );
buf \U$1800 ( \8637 , \7294 );
buf \U$1801 ( \8638 , \7294 );
buf \U$1802 ( \8639 , \7294 );
buf \U$1803 ( \8640 , \7294 );
buf \U$1804 ( \8641 , \7294 );
buf \U$1805 ( \8642 , \7294 );
nor \U$1806 ( \8643 , \7322 , \7323 , \7324 , \7325 , \7287 , \7291 , \7294 , \8618 , \8619 , \8620 , \8621 , \8622 , \8623 , \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 , \8632 , \8633 , \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 );
and \U$1807 ( \8644 , \7200 , \8643 );
buf \U$1808 ( \8645 , RIe3f8a98_6047);
buf \U$1809 ( \8646 , \7294 );
buf \U$1810 ( \8647 , \7294 );
buf \U$1811 ( \8648 , \7294 );
buf \U$1812 ( \8649 , \7294 );
buf \U$1813 ( \8650 , \7294 );
buf \U$1814 ( \8651 , \7294 );
buf \U$1815 ( \8652 , \7294 );
buf \U$1816 ( \8653 , \7294 );
buf \U$1817 ( \8654 , \7294 );
buf \U$1818 ( \8655 , \7294 );
buf \U$1819 ( \8656 , \7294 );
buf \U$1820 ( \8657 , \7294 );
buf \U$1821 ( \8658 , \7294 );
buf \U$1822 ( \8659 , \7294 );
buf \U$1823 ( \8660 , \7294 );
buf \U$1824 ( \8661 , \7294 );
buf \U$1825 ( \8662 , \7294 );
buf \U$1826 ( \8663 , \7294 );
buf \U$1827 ( \8664 , \7294 );
buf \U$1828 ( \8665 , \7294 );
buf \U$1829 ( \8666 , \7294 );
buf \U$1830 ( \8667 , \7294 );
buf \U$1831 ( \8668 , \7294 );
buf \U$1832 ( \8669 , \7294 );
buf \U$1833 ( \8670 , \7294 );
nor \U$1834 ( \8671 , \7281 , \7323 , \7324 , \7325 , \7287 , \7291 , \7294 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 , \8653 , \8654 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 , \8663 , \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 );
and \U$1835 ( \8672 , \8645 , \8671 );
buf \U$1836 ( \8673 , RIe385d90_5583);
buf \U$1837 ( \8674 , \7294 );
buf \U$1838 ( \8675 , \7294 );
buf \U$1839 ( \8676 , \7294 );
buf \U$1840 ( \8677 , \7294 );
buf \U$1841 ( \8678 , \7294 );
buf \U$1842 ( \8679 , \7294 );
buf \U$1843 ( \8680 , \7294 );
buf \U$1844 ( \8681 , \7294 );
buf \U$1845 ( \8682 , \7294 );
buf \U$1846 ( \8683 , \7294 );
buf \U$1847 ( \8684 , \7294 );
buf \U$1848 ( \8685 , \7294 );
buf \U$1849 ( \8686 , \7294 );
buf \U$1850 ( \8687 , \7294 );
buf \U$1851 ( \8688 , \7294 );
buf \U$1852 ( \8689 , \7294 );
buf \U$1853 ( \8690 , \7294 );
buf \U$1854 ( \8691 , \7294 );
buf \U$1855 ( \8692 , \7294 );
buf \U$1856 ( \8693 , \7294 );
buf \U$1857 ( \8694 , \7294 );
buf \U$1858 ( \8695 , \7294 );
buf \U$1859 ( \8696 , \7294 );
buf \U$1860 ( \8697 , \7294 );
buf \U$1861 ( \8698 , \7294 );
nor \U$1862 ( \8699 , \7322 , \7282 , \7324 , \7325 , \7287 , \7291 , \7294 , \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 , \8682 , \8683 , \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 , \8695 , \8696 , \8697 , \8698 );
and \U$1863 ( \8700 , \8673 , \8699 );
buf \U$1864 ( \8701 , RIe182a68_5243);
buf \U$1865 ( \8702 , \7294 );
buf \U$1866 ( \8703 , \7294 );
buf \U$1867 ( \8704 , \7294 );
buf \U$1868 ( \8705 , \7294 );
buf \U$1869 ( \8706 , \7294 );
buf \U$1870 ( \8707 , \7294 );
buf \U$1871 ( \8708 , \7294 );
buf \U$1872 ( \8709 , \7294 );
buf \U$1873 ( \8710 , \7294 );
buf \U$1874 ( \8711 , \7294 );
buf \U$1875 ( \8712 , \7294 );
buf \U$1876 ( \8713 , \7294 );
buf \U$1877 ( \8714 , \7294 );
buf \U$1878 ( \8715 , \7294 );
buf \U$1879 ( \8716 , \7294 );
buf \U$1880 ( \8717 , \7294 );
buf \U$1881 ( \8718 , \7294 );
buf \U$1882 ( \8719 , \7294 );
buf \U$1883 ( \8720 , \7294 );
buf \U$1884 ( \8721 , \7294 );
buf \U$1885 ( \8722 , \7294 );
buf \U$1886 ( \8723 , \7294 );
buf \U$1887 ( \8724 , \7294 );
buf \U$1888 ( \8725 , \7294 );
buf \U$1889 ( \8726 , \7294 );
nor \U$1890 ( \8727 , \7281 , \7282 , \7324 , \7325 , \7287 , \7291 , \7294 , \8702 , \8703 , \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 , \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 , \8722 , \8723 , \8724 , \8725 , \8726 );
and \U$1891 ( \8728 , \8701 , \8727 );
buf \U$1892 ( \8729 , RIe0f3008_4788);
buf \U$1893 ( \8730 , \7294 );
buf \U$1894 ( \8731 , \7294 );
buf \U$1895 ( \8732 , \7294 );
buf \U$1896 ( \8733 , \7294 );
buf \U$1897 ( \8734 , \7294 );
buf \U$1898 ( \8735 , \7294 );
buf \U$1899 ( \8736 , \7294 );
buf \U$1900 ( \8737 , \7294 );
buf \U$1901 ( \8738 , \7294 );
buf \U$1902 ( \8739 , \7294 );
buf \U$1903 ( \8740 , \7294 );
buf \U$1904 ( \8741 , \7294 );
buf \U$1905 ( \8742 , \7294 );
buf \U$1906 ( \8743 , \7294 );
buf \U$1907 ( \8744 , \7294 );
buf \U$1908 ( \8745 , \7294 );
buf \U$1909 ( \8746 , \7294 );
buf \U$1910 ( \8747 , \7294 );
buf \U$1911 ( \8748 , \7294 );
buf \U$1912 ( \8749 , \7294 );
buf \U$1913 ( \8750 , \7294 );
buf \U$1914 ( \8751 , \7294 );
buf \U$1915 ( \8752 , \7294 );
buf \U$1916 ( \8753 , \7294 );
buf \U$1917 ( \8754 , \7294 );
nor \U$1918 ( \8755 , \7322 , \7323 , \7283 , \7325 , \7287 , \7291 , \7294 , \8730 , \8731 , \8732 , \8733 , \8734 , \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 , \8742 , \8743 , \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 );
and \U$1919 ( \8756 , \8729 , \8755 );
buf \U$1920 ( \8757 , RIdfc11b8_4469);
buf \U$1921 ( \8758 , \7294 );
buf \U$1922 ( \8759 , \7294 );
buf \U$1923 ( \8760 , \7294 );
buf \U$1924 ( \8761 , \7294 );
buf \U$1925 ( \8762 , \7294 );
buf \U$1926 ( \8763 , \7294 );
buf \U$1927 ( \8764 , \7294 );
buf \U$1928 ( \8765 , \7294 );
buf \U$1929 ( \8766 , \7294 );
buf \U$1930 ( \8767 , \7294 );
buf \U$1931 ( \8768 , \7294 );
buf \U$1932 ( \8769 , \7294 );
buf \U$1933 ( \8770 , \7294 );
buf \U$1934 ( \8771 , \7294 );
buf \U$1935 ( \8772 , \7294 );
buf \U$1936 ( \8773 , \7294 );
buf \U$1937 ( \8774 , \7294 );
buf \U$1938 ( \8775 , \7294 );
buf \U$1939 ( \8776 , \7294 );
buf \U$1940 ( \8777 , \7294 );
buf \U$1941 ( \8778 , \7294 );
buf \U$1942 ( \8779 , \7294 );
buf \U$1943 ( \8780 , \7294 );
buf \U$1944 ( \8781 , \7294 );
buf \U$1945 ( \8782 , \7294 );
nor \U$1946 ( \8783 , \7281 , \7323 , \7283 , \7325 , \7287 , \7291 , \7294 , \8758 , \8759 , \8760 , \8761 , \8762 , \8763 , \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 , \8772 , \8773 , \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 , \8782 );
and \U$1947 ( \8784 , \8757 , \8783 );
buf \U$1948 ( \8785 , RIde5ad30_4003);
buf \U$1949 ( \8786 , \7294 );
buf \U$1950 ( \8787 , \7294 );
buf \U$1951 ( \8788 , \7294 );
buf \U$1952 ( \8789 , \7294 );
buf \U$1953 ( \8790 , \7294 );
buf \U$1954 ( \8791 , \7294 );
buf \U$1955 ( \8792 , \7294 );
buf \U$1956 ( \8793 , \7294 );
buf \U$1957 ( \8794 , \7294 );
buf \U$1958 ( \8795 , \7294 );
buf \U$1959 ( \8796 , \7294 );
buf \U$1960 ( \8797 , \7294 );
buf \U$1961 ( \8798 , \7294 );
buf \U$1962 ( \8799 , \7294 );
buf \U$1963 ( \8800 , \7294 );
buf \U$1964 ( \8801 , \7294 );
buf \U$1965 ( \8802 , \7294 );
buf \U$1966 ( \8803 , \7294 );
buf \U$1967 ( \8804 , \7294 );
buf \U$1968 ( \8805 , \7294 );
buf \U$1969 ( \8806 , \7294 );
buf \U$1970 ( \8807 , \7294 );
buf \U$1971 ( \8808 , \7294 );
buf \U$1972 ( \8809 , \7294 );
buf \U$1973 ( \8810 , \7294 );
nor \U$1974 ( \8811 , \7322 , \7282 , \7283 , \7325 , \7287 , \7291 , \7294 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 , \8792 , \8793 , \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 , \8802 , \8803 , \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 );
and \U$1975 ( \8812 , \8785 , \8811 );
buf \U$1976 ( \8813 , RIdd93500_3608);
buf \U$1977 ( \8814 , \7294 );
buf \U$1978 ( \8815 , \7294 );
buf \U$1979 ( \8816 , \7294 );
buf \U$1980 ( \8817 , \7294 );
buf \U$1981 ( \8818 , \7294 );
buf \U$1982 ( \8819 , \7294 );
buf \U$1983 ( \8820 , \7294 );
buf \U$1984 ( \8821 , \7294 );
buf \U$1985 ( \8822 , \7294 );
buf \U$1986 ( \8823 , \7294 );
buf \U$1987 ( \8824 , \7294 );
buf \U$1988 ( \8825 , \7294 );
buf \U$1989 ( \8826 , \7294 );
buf \U$1990 ( \8827 , \7294 );
buf \U$1991 ( \8828 , \7294 );
buf \U$1992 ( \8829 , \7294 );
buf \U$1993 ( \8830 , \7294 );
buf \U$1994 ( \8831 , \7294 );
buf \U$1995 ( \8832 , \7294 );
buf \U$1996 ( \8833 , \7294 );
buf \U$1997 ( \8834 , \7294 );
buf \U$1998 ( \8835 , \7294 );
buf \U$1999 ( \8836 , \7294 );
buf \U$2000 ( \8837 , \7294 );
buf \U$2001 ( \8838 , \7294 );
nor \U$2002 ( \8839 , \7281 , \7282 , \7283 , \7325 , \7287 , \7291 , \7294 , \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 , \8822 , \8823 , \8824 , \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 , \8832 , \8833 , \8834 , \8835 , \8836 , \8837 , \8838 );
and \U$2003 ( \8840 , \8813 , \8839 );
buf \U$2004 ( \8841 , RIdbcac48_3211);
buf \U$2005 ( \8842 , \7294 );
buf \U$2006 ( \8843 , \7294 );
buf \U$2007 ( \8844 , \7294 );
buf \U$2008 ( \8845 , \7294 );
buf \U$2009 ( \8846 , \7294 );
buf \U$2010 ( \8847 , \7294 );
buf \U$2011 ( \8848 , \7294 );
buf \U$2012 ( \8849 , \7294 );
buf \U$2013 ( \8850 , \7294 );
buf \U$2014 ( \8851 , \7294 );
buf \U$2015 ( \8852 , \7294 );
buf \U$2016 ( \8853 , \7294 );
buf \U$2017 ( \8854 , \7294 );
buf \U$2018 ( \8855 , \7294 );
buf \U$2019 ( \8856 , \7294 );
buf \U$2020 ( \8857 , \7294 );
buf \U$2021 ( \8858 , \7294 );
buf \U$2022 ( \8859 , \7294 );
buf \U$2023 ( \8860 , \7294 );
buf \U$2024 ( \8861 , \7294 );
buf \U$2025 ( \8862 , \7294 );
buf \U$2026 ( \8863 , \7294 );
buf \U$2027 ( \8864 , \7294 );
buf \U$2028 ( \8865 , \7294 );
buf \U$2029 ( \8866 , \7294 );
nor \U$2030 ( \8867 , \7322 , \7323 , \7324 , \7284 , \7287 , \7291 , \7294 , \8842 , \8843 , \8844 , \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 , \8852 , \8853 , \8854 , \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 , \8862 , \8863 , \8864 , \8865 , \8866 );
and \U$2031 ( \8868 , \8841 , \8867 );
buf \U$2032 ( \8869 , RIdaff2d8_2817);
buf \U$2033 ( \8870 , \7294 );
buf \U$2034 ( \8871 , \7294 );
buf \U$2035 ( \8872 , \7294 );
buf \U$2036 ( \8873 , \7294 );
buf \U$2037 ( \8874 , \7294 );
buf \U$2038 ( \8875 , \7294 );
buf \U$2039 ( \8876 , \7294 );
buf \U$2040 ( \8877 , \7294 );
buf \U$2041 ( \8878 , \7294 );
buf \U$2042 ( \8879 , \7294 );
buf \U$2043 ( \8880 , \7294 );
buf \U$2044 ( \8881 , \7294 );
buf \U$2045 ( \8882 , \7294 );
buf \U$2046 ( \8883 , \7294 );
buf \U$2047 ( \8884 , \7294 );
buf \U$2048 ( \8885 , \7294 );
buf \U$2049 ( \8886 , \7294 );
buf \U$2050 ( \8887 , \7294 );
buf \U$2051 ( \8888 , \7294 );
buf \U$2052 ( \8889 , \7294 );
buf \U$2053 ( \8890 , \7294 );
buf \U$2054 ( \8891 , \7294 );
buf \U$2055 ( \8892 , \7294 );
buf \U$2056 ( \8893 , \7294 );
buf \U$2057 ( \8894 , \7294 );
nor \U$2058 ( \8895 , \7281 , \7323 , \7324 , \7284 , \7287 , \7291 , \7294 , \8870 , \8871 , \8872 , \8873 , \8874 , \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 , \8882 , \8883 , \8884 , \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 , \8892 , \8893 , \8894 );
and \U$2059 ( \8896 , \8869 , \8895 );
buf \U$2060 ( \8897 , RIda2b970_2422);
buf \U$2061 ( \8898 , \7294 );
buf \U$2062 ( \8899 , \7294 );
buf \U$2063 ( \8900 , \7294 );
buf \U$2064 ( \8901 , \7294 );
buf \U$2065 ( \8902 , \7294 );
buf \U$2066 ( \8903 , \7294 );
buf \U$2067 ( \8904 , \7294 );
buf \U$2068 ( \8905 , \7294 );
buf \U$2069 ( \8906 , \7294 );
buf \U$2070 ( \8907 , \7294 );
buf \U$2071 ( \8908 , \7294 );
buf \U$2072 ( \8909 , \7294 );
buf \U$2073 ( \8910 , \7294 );
buf \U$2074 ( \8911 , \7294 );
buf \U$2075 ( \8912 , \7294 );
buf \U$2076 ( \8913 , \7294 );
buf \U$2077 ( \8914 , \7294 );
buf \U$2078 ( \8915 , \7294 );
buf \U$2079 ( \8916 , \7294 );
buf \U$2080 ( \8917 , \7294 );
buf \U$2081 ( \8918 , \7294 );
buf \U$2082 ( \8919 , \7294 );
buf \U$2083 ( \8920 , \7294 );
buf \U$2084 ( \8921 , \7294 );
buf \U$2085 ( \8922 , \7294 );
nor \U$2086 ( \8923 , \7322 , \7282 , \7324 , \7284 , \7287 , \7291 , \7294 , \8898 , \8899 , \8900 , \8901 , \8902 , \8903 , \8904 , \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 , \8912 , \8913 , \8914 , \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 , \8922 );
and \U$2087 ( \8924 , \8897 , \8923 );
buf \U$2088 ( \8925 , RId977f88_2027);
buf \U$2089 ( \8926 , \7294 );
buf \U$2090 ( \8927 , \7294 );
buf \U$2091 ( \8928 , \7294 );
buf \U$2092 ( \8929 , \7294 );
buf \U$2093 ( \8930 , \7294 );
buf \U$2094 ( \8931 , \7294 );
buf \U$2095 ( \8932 , \7294 );
buf \U$2096 ( \8933 , \7294 );
buf \U$2097 ( \8934 , \7294 );
buf \U$2098 ( \8935 , \7294 );
buf \U$2099 ( \8936 , \7294 );
buf \U$2100 ( \8937 , \7294 );
buf \U$2101 ( \8938 , \7294 );
buf \U$2102 ( \8939 , \7294 );
buf \U$2103 ( \8940 , \7294 );
buf \U$2104 ( \8941 , \7294 );
buf \U$2105 ( \8942 , \7294 );
buf \U$2106 ( \8943 , \7294 );
buf \U$2107 ( \8944 , \7294 );
buf \U$2108 ( \8945 , \7294 );
buf \U$2109 ( \8946 , \7294 );
buf \U$2110 ( \8947 , \7294 );
buf \U$2111 ( \8948 , \7294 );
buf \U$2112 ( \8949 , \7294 );
buf \U$2113 ( \8950 , \7294 );
nor \U$2114 ( \8951 , \7281 , \7282 , \7324 , \7284 , \7287 , \7291 , \7294 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 , \8932 , \8933 , \8934 , \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 , \8942 , \8943 , \8944 , \8945 , \8946 , \8947 , \8948 , \8949 , \8950 );
and \U$2115 ( \8952 , \8925 , \8951 );
buf \U$2116 ( \8953 , RId8ab538_1631);
buf \U$2117 ( \8954 , \7294 );
buf \U$2118 ( \8955 , \7294 );
buf \U$2119 ( \8956 , \7294 );
buf \U$2120 ( \8957 , \7294 );
buf \U$2121 ( \8958 , \7294 );
buf \U$2122 ( \8959 , \7294 );
buf \U$2123 ( \8960 , \7294 );
buf \U$2124 ( \8961 , \7294 );
buf \U$2125 ( \8962 , \7294 );
buf \U$2126 ( \8963 , \7294 );
buf \U$2127 ( \8964 , \7294 );
buf \U$2128 ( \8965 , \7294 );
buf \U$2129 ( \8966 , \7294 );
buf \U$2130 ( \8967 , \7294 );
buf \U$2131 ( \8968 , \7294 );
buf \U$2132 ( \8969 , \7294 );
buf \U$2133 ( \8970 , \7294 );
buf \U$2134 ( \8971 , \7294 );
buf \U$2135 ( \8972 , \7294 );
buf \U$2136 ( \8973 , \7294 );
buf \U$2137 ( \8974 , \7294 );
buf \U$2138 ( \8975 , \7294 );
buf \U$2139 ( \8976 , \7294 );
buf \U$2140 ( \8977 , \7294 );
buf \U$2141 ( \8978 , \7294 );
nor \U$2142 ( \8979 , \7322 , \7323 , \7283 , \7284 , \7287 , \7291 , \7294 , \8954 , \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 , \8962 , \8963 , \8964 , \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 , \8972 , \8973 , \8974 , \8975 , \8976 , \8977 , \8978 );
and \U$2143 ( \8980 , \8953 , \8979 );
buf \U$2144 ( \8981 , RId7e5f28_1234);
buf \U$2145 ( \8982 , \7294 );
buf \U$2146 ( \8983 , \7294 );
buf \U$2147 ( \8984 , \7294 );
buf \U$2148 ( \8985 , \7294 );
buf \U$2149 ( \8986 , \7294 );
buf \U$2150 ( \8987 , \7294 );
buf \U$2151 ( \8988 , \7294 );
buf \U$2152 ( \8989 , \7294 );
buf \U$2153 ( \8990 , \7294 );
buf \U$2154 ( \8991 , \7294 );
buf \U$2155 ( \8992 , \7294 );
buf \U$2156 ( \8993 , \7294 );
buf \U$2157 ( \8994 , \7294 );
buf \U$2158 ( \8995 , \7294 );
buf \U$2159 ( \8996 , \7294 );
buf \U$2160 ( \8997 , \7294 );
buf \U$2161 ( \8998 , \7294 );
buf \U$2162 ( \8999 , \7294 );
buf \U$2163 ( \9000 , \7294 );
buf \U$2164 ( \9001 , \7294 );
buf \U$2165 ( \9002 , \7294 );
buf \U$2166 ( \9003 , \7294 );
buf \U$2167 ( \9004 , \7294 );
buf \U$2168 ( \9005 , \7294 );
buf \U$2169 ( \9006 , \7294 );
nor \U$2170 ( \9007 , \7281 , \7323 , \7283 , \7284 , \7287 , \7291 , \7294 , \8982 , \8983 , \8984 , \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 , \8992 , \8993 , \8994 , \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 , \9002 , \9003 , \9004 , \9005 , \9006 );
and \U$2171 ( \9008 , \8981 , \9007 );
buf \U$2172 ( \9009 , RId71bad0_843);
buf \U$2173 ( \9010 , \7294 );
buf \U$2174 ( \9011 , \7294 );
buf \U$2175 ( \9012 , \7294 );
buf \U$2176 ( \9013 , \7294 );
buf \U$2177 ( \9014 , \7294 );
buf \U$2178 ( \9015 , \7294 );
buf \U$2179 ( \9016 , \7294 );
buf \U$2180 ( \9017 , \7294 );
buf \U$2181 ( \9018 , \7294 );
buf \U$2182 ( \9019 , \7294 );
buf \U$2183 ( \9020 , \7294 );
buf \U$2184 ( \9021 , \7294 );
buf \U$2185 ( \9022 , \7294 );
buf \U$2186 ( \9023 , \7294 );
buf \U$2187 ( \9024 , \7294 );
buf \U$2188 ( \9025 , \7294 );
buf \U$2189 ( \9026 , \7294 );
buf \U$2190 ( \9027 , \7294 );
buf \U$2191 ( \9028 , \7294 );
buf \U$2192 ( \9029 , \7294 );
buf \U$2193 ( \9030 , \7294 );
buf \U$2194 ( \9031 , \7294 );
buf \U$2195 ( \9032 , \7294 );
buf \U$2196 ( \9033 , \7294 );
buf \U$2197 ( \9034 , \7294 );
nor \U$2198 ( \9035 , \7322 , \7282 , \7283 , \7284 , \7287 , \7291 , \7294 , \9010 , \9011 , \9012 , \9013 , \9014 , \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 , \9022 , \9023 , \9024 , \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 , \9032 , \9033 , \9034 );
and \U$2199 ( \9036 , \9009 , \9035 );
or \U$2200 ( \9037 , \8617 , \8644 , \8672 , \8700 , \8728 , \8756 , \8784 , \8812 , \8840 , \8868 , \8896 , \8924 , \8952 , \8980 , \9008 , \9036 );
buf \U$2201 ( \9038 , \7294 );
not \U$2202 ( \9039 , \9038 );
buf \U$2203 ( \9040 , \7282 );
buf \U$2204 ( \9041 , \7283 );
buf \U$2205 ( \9042 , \7284 );
buf \U$2206 ( \9043 , \7287 );
buf \U$2207 ( \9044 , \7291 );
buf \U$2208 ( \9045 , \7294 );
buf \U$2209 ( \9046 , \7294 );
buf \U$2210 ( \9047 , \7294 );
buf \U$2211 ( \9048 , \7294 );
buf \U$2212 ( \9049 , \7294 );
buf \U$2213 ( \9050 , \7294 );
buf \U$2214 ( \9051 , \7294 );
buf \U$2215 ( \9052 , \7294 );
buf \U$2216 ( \9053 , \7294 );
buf \U$2217 ( \9054 , \7294 );
buf \U$2218 ( \9055 , \7294 );
buf \U$2219 ( \9056 , \7294 );
buf \U$2220 ( \9057 , \7294 );
buf \U$2221 ( \9058 , \7294 );
buf \U$2222 ( \9059 , \7294 );
buf \U$2223 ( \9060 , \7294 );
buf \U$2224 ( \9061 , \7294 );
buf \U$2225 ( \9062 , \7294 );
buf \U$2226 ( \9063 , \7294 );
buf \U$2227 ( \9064 , \7294 );
buf \U$2228 ( \9065 , \7294 );
buf \U$2229 ( \9066 , \7294 );
buf \U$2230 ( \9067 , \7294 );
buf \U$2231 ( \9068 , \7294 );
buf \U$2232 ( \9069 , \7294 );
buf \U$2233 ( \9070 , \7281 );
or \U$2234 ( \9071 , \9040 , \9041 , \9042 , \9043 , \9044 , \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 , \9052 , \9053 , \9054 , \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 , \9062 , \9063 , \9064 , \9065 , \9066 , \9067 , \9068 , \9069 , \9070 );
nand \U$2235 ( \9072 , \9039 , \9071 );
buf \U$2236 ( \9073 , \9072 );
buf \U$2237 ( \9074 , \7294 );
not \U$2238 ( \9075 , \9074 );
buf \U$2239 ( \9076 , \7291 );
buf \U$2240 ( \9077 , \7294 );
buf \U$2241 ( \9078 , \7294 );
buf \U$2242 ( \9079 , \7294 );
buf \U$2243 ( \9080 , \7294 );
buf \U$2244 ( \9081 , \7294 );
buf \U$2245 ( \9082 , \7294 );
buf \U$2246 ( \9083 , \7294 );
buf \U$2247 ( \9084 , \7294 );
buf \U$2248 ( \9085 , \7294 );
buf \U$2249 ( \9086 , \7294 );
buf \U$2250 ( \9087 , \7294 );
buf \U$2251 ( \9088 , \7294 );
buf \U$2252 ( \9089 , \7294 );
buf \U$2253 ( \9090 , \7294 );
buf \U$2254 ( \9091 , \7294 );
buf \U$2255 ( \9092 , \7294 );
buf \U$2256 ( \9093 , \7294 );
buf \U$2257 ( \9094 , \7294 );
buf \U$2258 ( \9095 , \7294 );
buf \U$2259 ( \9096 , \7294 );
buf \U$2260 ( \9097 , \7294 );
buf \U$2261 ( \9098 , \7294 );
buf \U$2262 ( \9099 , \7294 );
buf \U$2263 ( \9100 , \7294 );
buf \U$2264 ( \9101 , \7294 );
buf \U$2265 ( \9102 , \7287 );
buf \U$2266 ( \9103 , \7281 );
buf \U$2267 ( \9104 , \7282 );
buf \U$2268 ( \9105 , \7283 );
buf \U$2269 ( \9106 , \7284 );
or \U$2270 ( \9107 , \9103 , \9104 , \9105 , \9106 );
and \U$2271 ( \9108 , \9102 , \9107 );
or \U$2272 ( \9109 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 , \9082 , \9083 , \9084 , \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 , \9092 , \9093 , \9094 , \9095 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 , \9108 );
and \U$2273 ( \9110 , \9075 , \9109 );
buf \U$2274 ( \9111 , \9110 );
or \U$2275 ( \9112 , \9073 , \9111 );
_DC g3a82 ( \9113_nG3a82 , \9037 , \9112 );
buf \U$2276 ( \9114 , \9113_nG3a82 );
xor \U$2277 ( \9115 , \8590 , \9114 );
buf \U$2278 ( \9116 , RIb7af5b8_255);
and \U$2279 ( \9117 , \7207 , \8616 );
and \U$2280 ( \9118 , \7209 , \8643 );
buf \U$2281 ( \9119 , RIe450d88_5972);
and \U$2282 ( \9120 , \9119 , \8671 );
buf \U$2283 ( \9121 , RIe386678_5582);
and \U$2284 ( \9122 , \9121 , \8699 );
buf \U$2285 ( \9123 , RIe1bcc68_5184);
and \U$2286 ( \9124 , \9123 , \8727 );
buf \U$2287 ( \9125 , RIe088e38_4865);
and \U$2288 ( \9126 , \9125 , \8755 );
buf \U$2289 ( \9127 , RIdfc07e0_4470);
and \U$2290 ( \9128 , \9127 , \8783 );
buf \U$2291 ( \9129 , RIde5b618_4002);
and \U$2292 ( \9130 , \9129 , \8811 );
buf \U$2293 ( \9131 , RIdd93ed8_3607);
and \U$2294 ( \9132 , \9131 , \8839 );
buf \U$2295 ( \9133 , RIdb62338_3285);
and \U$2296 ( \9134 , \9133 , \8867 );
buf \U$2297 ( \9135 , RIdaffda0_2816);
and \U$2298 ( \9136 , \9135 , \8895 );
buf \U$2299 ( \9137 , RIda2c258_2421);
and \U$2300 ( \9138 , \9137 , \8923 );
buf \U$2301 ( \9139 , RId978960_2026);
and \U$2302 ( \9140 , \9139 , \8951 );
buf \U$2303 ( \9141 , RId8ae508_1629);
and \U$2304 ( \9142 , \9141 , \8979 );
buf \U$2305 ( \9143 , RId7827c0_1310);
and \U$2306 ( \9144 , \9143 , \9007 );
buf \U$2307 ( \9145 , RId71c2c8_842);
and \U$2308 ( \9146 , \9145 , \9035 );
or \U$2309 ( \9147 , \9117 , \9118 , \9120 , \9122 , \9124 , \9126 , \9128 , \9130 , \9132 , \9134 , \9136 , \9138 , \9140 , \9142 , \9144 , \9146 );
_DC g3aa5 ( \9148_nG3aa5 , \9147 , \9112 );
buf \U$2310 ( \9149 , \9148_nG3aa5 );
xor \U$2311 ( \9150 , \9116 , \9149 );
or \U$2312 ( \9151 , \9115 , \9150 );
buf \U$2313 ( \9152 , RIb7af540_256);
and \U$2314 ( \9153 , \7217 , \8616 );
and \U$2315 ( \9154 , \7219 , \8643 );
buf \U$2316 ( \9155 , RIe3f8048_6048);
and \U$2317 ( \9156 , \9155 , \8671 );
buf \U$2318 ( \9157 , RIe386e70_5581);
and \U$2319 ( \9158 , \9157 , \8699 );
buf \U$2320 ( \9159 , RIe1bd4d8_5183);
and \U$2321 ( \9160 , \9159 , \8727 );
buf \U$2322 ( \9161 , RIe0af538_4863);
and \U$2323 ( \9162 , \9161 , \8755 );
buf \U$2324 ( \9163 , RIe02a050_4392);
and \U$2325 ( \9164 , \9163 , \8783 );
buf \U$2326 ( \9165 , RIde5be10_4001);
and \U$2327 ( \9166 , \9165 , \8811 );
buf \U$2328 ( \9167 , RIdd94928_3606);
and \U$2329 ( \9168 , \9167 , \8839 );
buf \U$2330 ( \9169 , RIdbcb530_3210);
and \U$2331 ( \9170 , \9169 , \8867 );
buf \U$2332 ( \9171 , RIdb00bb0_2815);
and \U$2333 ( \9172 , \9171 , \8895 );
buf \U$2334 ( \9173 , RId9cdfc8_2495);
and \U$2335 ( \9174 , \9173 , \8923 );
buf \U$2336 ( \9175 , RId9791d0_2025);
and \U$2337 ( \9176 , \9175 , \8951 );
buf \U$2338 ( \9177 , RId86cf28_1704);
and \U$2339 ( \9178 , \9177 , \8979 );
buf \U$2340 ( \9179 , RId7e6798_1233);
and \U$2341 ( \9180 , \9179 , \9007 );
buf \U$2342 ( \9181 , RId71cb38_841);
and \U$2343 ( \9182 , \9181 , \9035 );
or \U$2344 ( \9183 , \9153 , \9154 , \9156 , \9158 , \9160 , \9162 , \9164 , \9166 , \9168 , \9170 , \9172 , \9174 , \9176 , \9178 , \9180 , \9182 );
_DC g3ac9 ( \9184_nG3ac9 , \9183 , \9112 );
buf \U$2345 ( \9185 , \9184_nG3ac9 );
xor \U$2346 ( \9186 , \9152 , \9185 );
or \U$2347 ( \9187 , \9151 , \9186 );
buf \U$2348 ( \9188 , RIb7af4c8_257);
and \U$2349 ( \9189 , \7227 , \8616 );
and \U$2350 ( \9190 , \7229 , \8643 );
buf \U$2351 ( \9191 , RIe3e5628_6050);
and \U$2352 ( \9192 , \9191 , \8671 );
buf \U$2353 ( \9193 , RIe3876e0_5580);
and \U$2354 ( \9194 , \9193 , \8699 );
buf \U$2355 ( \9195 , RIe1bdd48_5182);
and \U$2356 ( \9196 , \9195 , \8727 );
buf \U$2357 ( \9197 , RIe0aeb60_4864);
and \U$2358 ( \9198 , \9197 , \8755 );
buf \U$2359 ( \9199 , RIe02a8c0_4391);
and \U$2360 ( \9200 , \9199 , \8783 );
buf \U$2361 ( \9201 , RIde5c6f8_4000);
and \U$2362 ( \9202 , \9201 , \8811 );
buf \U$2363 ( \9203 , RIdd95288_3605);
and \U$2364 ( \9204 , \9203 , \8839 );
buf \U$2365 ( \9205 , RIdb8a760_3284);
and \U$2366 ( \9206 , \9205 , \8867 );
buf \U$2367 ( \9207 , RIdabee68_2890);
and \U$2368 ( \9208 , \9207 , \8895 );
buf \U$2369 ( \9209 , RIda2cbb8_2420);
and \U$2370 ( \9210 , \9209 , \8923 );
buf \U$2371 ( \9211 , RId9799c8_2024);
and \U$2372 ( \9212 , \9211 , \8951 );
buf \U$2373 ( \9213 , RId8aed00_1628);
and \U$2374 ( \9214 , \9213 , \8979 );
buf \U$2375 ( \9215 , RId790848_1309);
and \U$2376 ( \9216 , \9215 , \9007 );
buf \U$2377 ( \9217 , RId71d330_840);
and \U$2378 ( \9218 , \9217 , \9035 );
or \U$2379 ( \9219 , \9189 , \9190 , \9192 , \9194 , \9196 , \9198 , \9200 , \9202 , \9204 , \9206 , \9208 , \9210 , \9212 , \9214 , \9216 , \9218 );
_DC g3aed ( \9220_nG3aed , \9219 , \9112 );
buf \U$2380 ( \9221 , \9220_nG3aed );
xor \U$2381 ( \9222 , \9188 , \9221 );
or \U$2382 ( \9223 , \9187 , \9222 );
buf \U$2383 ( \9224 , RIb7af450_258);
and \U$2384 ( \9225 , \7237 , \8616 );
and \U$2385 ( \9226 , \7239 , \8643 );
buf \U$2386 ( \9227 , RIe3f9e48_6045);
and \U$2387 ( \9228 , \9227 , \8671 );
buf \U$2388 ( \9229 , RIe387ed8_5579);
and \U$2389 ( \9230 , \9229 , \8699 );
buf \U$2390 ( \9231 , RIe183440_5242);
and \U$2391 ( \9232 , \9231 , \8727 );
buf \U$2392 ( \9233 , RIe0aff10_4862);
and \U$2393 ( \9234 , \9233 , \8755 );
buf \U$2394 ( \9235 , RIdfcdc38_4468);
and \U$2395 ( \9236 , \9235 , \8783 );
buf \U$2396 ( \9237 , RIde5cf68_3999);
and \U$2397 ( \9238 , \9237 , \8811 );
buf \U$2398 ( \9239 , RIdd95b70_3604);
and \U$2399 ( \9240 , \9239 , \8839 );
buf \U$2400 ( \9241 , RIdbcbe18_3209);
and \U$2401 ( \9242 , \9241 , \8867 );
buf \U$2402 ( \9243 , RIdb01498_2814);
and \U$2403 ( \9244 , \9243 , \8895 );
buf \U$2404 ( \9245 , RIda2d4a0_2419);
and \U$2405 ( \9246 , \9245 , \8923 );
buf \U$2406 ( \9247 , RId97a238_2023);
and \U$2407 ( \9248 , \9247 , \8951 );
buf \U$2408 ( \9249 , RId8af7c8_1627);
and \U$2409 ( \9250 , \9249 , \8979 );
buf \U$2410 ( \9251 , RId7a41e0_1308);
and \U$2411 ( \9252 , \9251 , \9007 );
buf \U$2412 ( \9253 , RId71dba0_839);
and \U$2413 ( \9254 , \9253 , \9035 );
or \U$2414 ( \9255 , \9225 , \9226 , \9228 , \9230 , \9232 , \9234 , \9236 , \9238 , \9240 , \9242 , \9244 , \9246 , \9248 , \9250 , \9252 , \9254 );
_DC g3b03 ( \9256_nG3b03 , \9255 , \9112 );
buf \U$2415 ( \9257 , \9256_nG3b03 );
xor \U$2416 ( \9258 , \9224 , \9257 );
or \U$2417 ( \9259 , \9223 , \9258 );
buf \U$2418 ( \9260 , RIb7af3d8_259);
and \U$2419 ( \9261 , \7247 , \8616 );
and \U$2420 ( \9262 , \7249 , \8643 );
buf \U$2421 ( \9263 , RIe3f7760_6049);
and \U$2422 ( \9264 , \9263 , \8671 );
buf \U$2423 ( \9265 , RIe3887c0_5578);
and \U$2424 ( \9266 , \9265 , \8699 );
buf \U$2425 ( \9267 , RIe15c260_5259);
and \U$2426 ( \9268 , \9267 , \8727 );
buf \U$2427 ( \9269 , RIe0f3878_4787);
and \U$2428 ( \9270 , \9269 , \8755 );
buf \U$2429 ( \9271 , RIdfce700_4467);
and \U$2430 ( \9272 , \9271 , \8783 );
buf \U$2431 ( \9273 , RIde5d760_3998);
and \U$2432 ( \9274 , \9273 , \8811 );
buf \U$2433 ( \9275 , RIdd963e0_3603);
and \U$2434 ( \9276 , \9275 , \8839 );
buf \U$2435 ( \9277 , RIdbcc7f0_3208);
and \U$2436 ( \9278 , \9277 , \8867 );
buf \U$2437 ( \9279 , RIdb01d80_2813);
and \U$2438 ( \9280 , \9279 , \8895 );
buf \U$2439 ( \9281 , RIda2def0_2418);
and \U$2440 ( \9282 , \9281 , \8923 );
buf \U$2441 ( \9283 , RId97ab20_2022);
and \U$2442 ( \9284 , \9283 , \8951 );
buf \U$2443 ( \9285 , RId8ac078_1630);
and \U$2444 ( \9286 , \9285 , \8979 );
buf \U$2445 ( \9287 , RId7e6f90_1232);
and \U$2446 ( \9288 , \9287 , \9007 );
buf \U$2447 ( \9289 , RId71e398_838);
and \U$2448 ( \9290 , \9289 , \9035 );
or \U$2449 ( \9291 , \9261 , \9262 , \9264 , \9266 , \9268 , \9270 , \9272 , \9274 , \9276 , \9278 , \9280 , \9282 , \9284 , \9286 , \9288 , \9290 );
_DC g3b19 ( \9292_nG3b19 , \9291 , \9112 );
buf \U$2450 ( \9293 , \9292_nG3b19 );
xor \U$2451 ( \9294 , \9260 , \9293 );
or \U$2452 ( \9295 , \9259 , \9294 );
buf \U$2453 ( \9296 , RIb7a5bf8_260);
and \U$2454 ( \9297 , \7257 , \8616 );
and \U$2455 ( \9298 , \7259 , \8643 );
buf \U$2456 ( \9299 , RIe451670_5971);
and \U$2457 ( \9300 , \9299 , \8671 );
buf \U$2458 ( \9301 , RIe388fb8_5577);
and \U$2459 ( \9302 , \9301 , \8699 );
buf \U$2460 ( \9303 , RIe1be5b8_5181);
and \U$2461 ( \9304 , \9303 , \8727 );
buf \U$2462 ( \9305 , RIe0b0870_4861);
and \U$2463 ( \9306 , \9305 , \8755 );
buf \U$2464 ( \9307 , RIdfcf2b8_4466);
and \U$2465 ( \9308 , \9307 , \8783 );
buf \U$2466 ( \9309 , RIde5dfd0_3997);
and \U$2467 ( \9310 , \9309 , \8811 );
buf \U$2468 ( \9311 , RIdd96cc8_3602);
and \U$2469 ( \9312 , \9311 , \8839 );
buf \U$2470 ( \9313 , RIdbcd0d8_3207);
and \U$2471 ( \9314 , \9313 , \8867 );
buf \U$2472 ( \9315 , RIdb02668_2812);
and \U$2473 ( \9316 , \9315 , \8895 );
buf \U$2474 ( \9317 , RIda2e760_2417);
and \U$2475 ( \9318 , \9317 , \8923 );
buf \U$2476 ( \9319 , RId97b318_2021);
and \U$2477 ( \9320 , \9319 , \8951 );
buf \U$2478 ( \9321 , RId86c4d8_1705);
and \U$2479 ( \9322 , \9321 , \8979 );
buf \U$2480 ( \9323 , RId7a4bb8_1307);
and \U$2481 ( \9324 , \9323 , \9007 );
buf \U$2482 ( \9325 , RId71ec08_837);
and \U$2483 ( \9326 , \9325 , \9035 );
or \U$2484 ( \9327 , \9297 , \9298 , \9300 , \9302 , \9304 , \9306 , \9308 , \9310 , \9312 , \9314 , \9316 , \9318 , \9320 , \9322 , \9324 , \9326 );
_DC g3b2f ( \9328_nG3b2f , \9327 , \9112 );
buf \U$2485 ( \9329 , \9328_nG3b2f );
xor \U$2486 ( \9330 , \9296 , \9329 );
or \U$2487 ( \9331 , \9295 , \9330 );
buf \U$2488 ( \9332 , RIb7a0c48_261);
and \U$2489 ( \9333 , \7267 , \8616 );
and \U$2490 ( \9334 , \7269 , \8643 );
buf \U$2491 ( \9335 , RIe3f9470_6046);
and \U$2492 ( \9336 , \9335 , \8671 );
buf \U$2493 ( \9337 , RIe3898a0_5576);
and \U$2494 ( \9338 , \9337 , \8699 );
buf \U$2495 ( \9339 , RIe15b900_5260);
and \U$2496 ( \9340 , \9339 , \8727 );
buf \U$2497 ( \9341 , RIe0f4070_4786);
and \U$2498 ( \9342 , \9341 , \8755 );
buf \U$2499 ( \9343 , RIdfcfc90_4465);
and \U$2500 ( \9344 , \9343 , \8783 );
buf \U$2501 ( \9345 , RIde5e840_3996);
and \U$2502 ( \9346 , \9345 , \8811 );
buf \U$2503 ( \9347 , RIdd97538_3601);
and \U$2504 ( \9348 , \9347 , \8839 );
buf \U$2505 ( \9349 , RIdbcd9c0_3206);
and \U$2506 ( \9350 , \9349 , \8867 );
buf \U$2507 ( \9351 , RIdb02f50_2811);
and \U$2508 ( \9352 , \9351 , \8895 );
buf \U$2509 ( \9353 , RIda2f0c0_2416);
and \U$2510 ( \9354 , \9353 , \8923 );
buf \U$2511 ( \9355 , RId97bc00_2020);
and \U$2512 ( \9356 , \9355 , \8951 );
buf \U$2513 ( \9357 , RId8b0290_1626);
and \U$2514 ( \9358 , \9357 , \8979 );
buf \U$2515 ( \9359 , RId7e7800_1231);
and \U$2516 ( \9360 , \9359 , \9007 );
buf \U$2517 ( \9361 , RId71f400_836);
and \U$2518 ( \9362 , \9361 , \9035 );
or \U$2519 ( \9363 , \9333 , \9334 , \9336 , \9338 , \9340 , \9342 , \9344 , \9346 , \9348 , \9350 , \9352 , \9354 , \9356 , \9358 , \9360 , \9362 );
_DC g3b45 ( \9364_nG3b45 , \9363 , \9112 );
buf \U$2520 ( \9365 , \9364_nG3b45 );
xor \U$2521 ( \9366 , \9332 , \9365 );
or \U$2522 ( \9367 , \9331 , \9366 );
not \U$2523 ( \9368 , \9367 );
buf \U$2524 ( \9369 , \9368 );
and \U$2525 ( \9370 , \8589 , \9369 );
_HMUX g3b4c ( \9371_nG3b4c , RIe5319e0_6884 , \7281 , \9370 );
buf \U$2526 ( \9372 , \7096 );
buf \U$2527 ( \9373 , \7093 );
buf \U$2528 ( \9374 , \7078 );
buf \U$2529 ( \9375 , \7081 );
buf \U$2530 ( \9376 , \7085 );
buf \U$2531 ( \9377 , \7089 );
or \U$2532 ( \9378 , \9374 , \9375 , \9376 , \9377 );
and \U$2533 ( \9379 , \9373 , \9378 );
or \U$2534 ( \9380 , \9372 , \9379 );
buf \U$2535 ( \9381 , \9380 );
_HMUX g3b57 ( \9382_nG3b57 , \7280_nG3351 , \9371_nG3b4c , \9381 );
buf \U$2536 ( \9383 , RIe5319e0_6884);
buf \U$2538 ( \9384 , \9383 );
buf \U$2539 ( \9385 , RIe549ef0_6842);
not \U$2540 ( \9386 , \9385 );
buf \U$2541 ( \9387 , \9386 );
buf \U$2542 ( \9388 , RIe549770_6843);
xnor \U$2543 ( \9389 , \9388 , \9385 );
buf \U$2544 ( \9390 , \9389 );
buf \U$2545 ( \9391 , RIe548ff0_6844);
or \U$2546 ( \9392 , \9388 , \9385 );
xnor \U$2547 ( \9393 , \9391 , \9392 );
buf \U$2548 ( \9394 , \9393 );
buf \U$2549 ( \9395 , RIea91330_6888);
or \U$2550 ( \9396 , \9391 , \9392 );
xor \U$2551 ( \9397 , \9395 , \9396 );
buf \U$2552 ( \9398 , \9397 );
not \U$2553 ( \9399 , \9398 );
and \U$2554 ( \9400 , \9395 , \9396 );
buf \U$2555 ( \9401 , \9400 );
nor \U$2556 ( \9402 , \9384 , \9387 , \9390 , \9394 , \9399 , \9401 );
and \U$2557 ( \9403 , RIe5329d0_6883, \9402 );
not \U$2558 ( \9404 , \9401 );
and \U$2559 ( \9405 , \9384 , \9387 , \9390 , \9394 , \9399 , \9404 );
and \U$2560 ( \9406 , RIeb72150_6905, \9405 );
not \U$2561 ( \9407 , \9384 );
and \U$2562 ( \9408 , \9407 , \9387 , \9390 , \9394 , \9399 , \9404 );
and \U$2563 ( \9409 , RIeab80c0_6897, \9408 );
or \U$2577 ( \9410 , \9403 , \9406 , \9409 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
buf \U$2579 ( \9411 , \9401 );
buf \U$2580 ( \9412 , \9398 );
buf \U$2581 ( \9413 , \9384 );
buf \U$2582 ( \9414 , \9387 );
buf \U$2583 ( \9415 , \9390 );
buf \U$2584 ( \9416 , \9394 );
or \U$2585 ( \9417 , \9413 , \9414 , \9415 , \9416 );
and \U$2586 ( \9418 , \9412 , \9417 );
or \U$2587 ( \9419 , \9411 , \9418 );
buf \U$2588 ( \9420 , \9419 );
or \U$2589 ( \9421 , 1'b0 , \9420 );
_DC g3b80 ( \9422_nG3b80 , \9410 , \9421 );
not \U$2590 ( \9423 , \9422_nG3b80 );
buf \U$2591 ( \9424 , RIb7b9608_246);
and \U$2592 ( \9425 , \7117 , \9402 );
and \U$2593 ( \9426 , \7119 , \9405 );
and \U$2594 ( \9427 , \7864 , \9408 );
or \U$2608 ( \9428 , \9425 , \9426 , \9427 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3b87 ( \9429_nG3b87 , \9428 , \9421 );
buf \U$2609 ( \9430 , \9429_nG3b87 );
xor \U$2610 ( \9431 , \9424 , \9430 );
buf \U$2611 ( \9432 , RIb7b9590_247);
and \U$2612 ( \9433 , \7126 , \9402 );
and \U$2613 ( \9434 , \7128 , \9405 );
and \U$2614 ( \9435 , \8338 , \9408 );
or \U$2628 ( \9436 , \9433 , \9434 , \9435 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3b8f ( \9437_nG3b8f , \9436 , \9421 );
buf \U$2629 ( \9438 , \9437_nG3b8f );
xor \U$2630 ( \9439 , \9432 , \9438 );
or \U$2631 ( \9440 , \9431 , \9439 );
buf \U$2632 ( \9441 , RIb7b9518_248);
and \U$2633 ( \9442 , \7136 , \9402 );
and \U$2634 ( \9443 , \7138 , \9405 );
and \U$2635 ( \9444 , \8374 , \9408 );
or \U$2649 ( \9445 , \9442 , \9443 , \9444 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3b98 ( \9446_nG3b98 , \9445 , \9421 );
buf \U$2650 ( \9447 , \9446_nG3b98 );
xor \U$2651 ( \9448 , \9441 , \9447 );
or \U$2652 ( \9449 , \9440 , \9448 );
buf \U$2653 ( \9450 , RIb7b94a0_249);
and \U$2654 ( \9451 , \7146 , \9402 );
and \U$2655 ( \9452 , \7148 , \9405 );
and \U$2656 ( \9453 , \8410 , \9408 );
or \U$2670 ( \9454 , \9451 , \9452 , \9453 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3ba1 ( \9455_nG3ba1 , \9454 , \9421 );
buf \U$2671 ( \9456 , \9455_nG3ba1 );
xor \U$2672 ( \9457 , \9450 , \9456 );
or \U$2673 ( \9458 , \9449 , \9457 );
buf \U$2674 ( \9459 , RIb7b9428_250);
and \U$2675 ( \9460 , \7156 , \9402 );
and \U$2676 ( \9461 , \7158 , \9405 );
and \U$2677 ( \9462 , \8446 , \9408 );
or \U$2691 ( \9463 , \9460 , \9461 , \9462 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3baa ( \9464_nG3baa , \9463 , \9421 );
buf \U$2692 ( \9465 , \9464_nG3baa );
xor \U$2693 ( \9466 , \9459 , \9465 );
or \U$2694 ( \9467 , \9458 , \9466 );
buf \U$2695 ( \9468 , RIb7b93b0_251);
and \U$2696 ( \9469 , \7166 , \9402 );
and \U$2697 ( \9470 , \7168 , \9405 );
and \U$2698 ( \9471 , \8482 , \9408 );
or \U$2712 ( \9472 , \9469 , \9470 , \9471 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3bb3 ( \9473_nG3bb3 , \9472 , \9421 );
buf \U$2713 ( \9474 , \9473_nG3bb3 );
xor \U$2714 ( \9475 , \9468 , \9474 );
or \U$2715 ( \9476 , \9467 , \9475 );
buf \U$2716 ( \9477 , RIb7af720_252);
and \U$2717 ( \9478 , \7176 , \9402 );
and \U$2718 ( \9479 , \7178 , \9405 );
and \U$2719 ( \9480 , \8518 , \9408 );
or \U$2733 ( \9481 , \9478 , \9479 , \9480 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3bbc ( \9482_nG3bbc , \9481 , \9421 );
buf \U$2734 ( \9483 , \9482_nG3bbc );
xor \U$2735 ( \9484 , \9477 , \9483 );
or \U$2736 ( \9485 , \9476 , \9484 );
buf \U$2737 ( \9486 , RIb7af6a8_253);
and \U$2738 ( \9487 , \7186 , \9402 );
and \U$2739 ( \9488 , \7188 , \9405 );
and \U$2740 ( \9489 , \8554 , \9408 );
or \U$2754 ( \9490 , \9487 , \9488 , \9489 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3bc5 ( \9491_nG3bc5 , \9490 , \9421 );
buf \U$2755 ( \9492 , \9491_nG3bc5 );
xor \U$2756 ( \9493 , \9486 , \9492 );
or \U$2757 ( \9494 , \9485 , \9493 );
not \U$2758 ( \9495 , \9494 );
buf \U$2759 ( \9496 , \9495 );
buf \U$2760 ( \9497 , RIb7af630_254);
and \U$2761 ( \9498 , \7198 , \9402 );
and \U$2762 ( \9499 , \7200 , \9405 );
and \U$2763 ( \9500 , \8645 , \9408 );
or \U$2777 ( \9501 , \9498 , \9499 , \9500 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3bd0 ( \9502_nG3bd0 , \9501 , \9421 );
buf \U$2778 ( \9503 , \9502_nG3bd0 );
xor \U$2779 ( \9504 , \9497 , \9503 );
buf \U$2780 ( \9505 , RIb7af5b8_255);
and \U$2781 ( \9506 , \7207 , \9402 );
and \U$2782 ( \9507 , \7209 , \9405 );
and \U$2783 ( \9508 , \9119 , \9408 );
or \U$2797 ( \9509 , \9506 , \9507 , \9508 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3bd8 ( \9510_nG3bd8 , \9509 , \9421 );
buf \U$2798 ( \9511 , \9510_nG3bd8 );
xor \U$2799 ( \9512 , \9505 , \9511 );
or \U$2800 ( \9513 , \9504 , \9512 );
buf \U$2801 ( \9514 , RIb7af540_256);
and \U$2802 ( \9515 , \7217 , \9402 );
and \U$2803 ( \9516 , \7219 , \9405 );
and \U$2804 ( \9517 , \9155 , \9408 );
or \U$2818 ( \9518 , \9515 , \9516 , \9517 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3be1 ( \9519_nG3be1 , \9518 , \9421 );
buf \U$2819 ( \9520 , \9519_nG3be1 );
xor \U$2820 ( \9521 , \9514 , \9520 );
or \U$2821 ( \9522 , \9513 , \9521 );
buf \U$2822 ( \9523 , RIb7af4c8_257);
and \U$2823 ( \9524 , \7227 , \9402 );
and \U$2824 ( \9525 , \7229 , \9405 );
and \U$2825 ( \9526 , \9191 , \9408 );
or \U$2839 ( \9527 , \9524 , \9525 , \9526 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3bea ( \9528_nG3bea , \9527 , \9421 );
buf \U$2840 ( \9529 , \9528_nG3bea );
xor \U$2841 ( \9530 , \9523 , \9529 );
or \U$2842 ( \9531 , \9522 , \9530 );
buf \U$2843 ( \9532 , RIb7af450_258);
and \U$2844 ( \9533 , \7237 , \9402 );
and \U$2845 ( \9534 , \7239 , \9405 );
and \U$2846 ( \9535 , \9227 , \9408 );
or \U$2860 ( \9536 , \9533 , \9534 , \9535 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3bf3 ( \9537_nG3bf3 , \9536 , \9421 );
buf \U$2861 ( \9538 , \9537_nG3bf3 );
xor \U$2862 ( \9539 , \9532 , \9538 );
or \U$2863 ( \9540 , \9531 , \9539 );
buf \U$2864 ( \9541 , RIb7af3d8_259);
and \U$2865 ( \9542 , \7247 , \9402 );
and \U$2866 ( \9543 , \7249 , \9405 );
and \U$2867 ( \9544 , \9263 , \9408 );
or \U$2881 ( \9545 , \9542 , \9543 , \9544 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3bfc ( \9546_nG3bfc , \9545 , \9421 );
buf \U$2882 ( \9547 , \9546_nG3bfc );
xor \U$2883 ( \9548 , \9541 , \9547 );
or \U$2884 ( \9549 , \9540 , \9548 );
buf \U$2885 ( \9550 , RIb7a5bf8_260);
and \U$2886 ( \9551 , \7257 , \9402 );
and \U$2887 ( \9552 , \7259 , \9405 );
and \U$2888 ( \9553 , \9299 , \9408 );
or \U$2902 ( \9554 , \9551 , \9552 , \9553 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3c05 ( \9555_nG3c05 , \9554 , \9421 );
buf \U$2903 ( \9556 , \9555_nG3c05 );
xor \U$2904 ( \9557 , \9550 , \9556 );
or \U$2905 ( \9558 , \9549 , \9557 );
buf \U$2906 ( \9559 , RIb7a0c48_261);
and \U$2907 ( \9560 , \7267 , \9402 );
and \U$2908 ( \9561 , \7269 , \9405 );
and \U$2909 ( \9562 , \9335 , \9408 );
or \U$2923 ( \9563 , \9560 , \9561 , \9562 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g3c0e ( \9564_nG3c0e , \9563 , \9421 );
buf \U$2924 ( \9565 , \9564_nG3c0e );
xor \U$2925 ( \9566 , \9559 , \9565 );
or \U$2926 ( \9567 , \9558 , \9566 );
not \U$2927 ( \9568 , \9567 );
buf \U$2928 ( \9569 , \9568 );
and \U$2929 ( \9570 , \9496 , \9569 );
and \U$2930 ( \9571 , \9423 , \9570 );
_HMUX g3c16 ( \9572_nG3c16 , \9382_nG3b57 , \9384 , \9571 );
buf \U$2933 ( \9573 , \9384 );
buf \U$2936 ( \9574 , \9387 );
buf \U$2939 ( \9575 , \9390 );
buf \U$2942 ( \9576 , \9394 );
buf \U$2943 ( \9577 , \9398 );
not \U$2944 ( \9578 , \9577 );
buf \U$2945 ( \9579 , \9578 );
not \U$2946 ( \9580 , \9579 );
buf \U$2947 ( \9581 , \9401 );
xnor \U$2948 ( \9582 , \9581 , \9577 );
buf \U$2949 ( \9583 , \9582 );
or \U$2950 ( \9584 , \9581 , \9577 );
not \U$2951 ( \9585 , \9584 );
buf \U$2952 ( \9586 , \9585 );
buf \U$2953 ( \9587 , \9586 );
buf \U$2954 ( \9588 , \9586 );
buf \U$2955 ( \9589 , \9586 );
buf \U$2956 ( \9590 , \9586 );
buf \U$2957 ( \9591 , \9586 );
buf \U$2958 ( \9592 , \9586 );
buf \U$2959 ( \9593 , \9586 );
buf \U$2960 ( \9594 , \9586 );
buf \U$2961 ( \9595 , \9586 );
buf \U$2962 ( \9596 , \9586 );
buf \U$2963 ( \9597 , \9586 );
buf \U$2964 ( \9598 , \9586 );
buf \U$2965 ( \9599 , \9586 );
buf \U$2966 ( \9600 , \9586 );
buf \U$2967 ( \9601 , \9586 );
buf \U$2968 ( \9602 , \9586 );
buf \U$2969 ( \9603 , \9586 );
buf \U$2970 ( \9604 , \9586 );
buf \U$2971 ( \9605 , \9586 );
buf \U$2972 ( \9606 , \9586 );
buf \U$2973 ( \9607 , \9586 );
buf \U$2974 ( \9608 , \9586 );
buf \U$2975 ( \9609 , \9586 );
buf \U$2976 ( \9610 , \9586 );
buf \U$2977 ( \9611 , \9586 );
nor \U$2978 ( \9612 , \9573 , \9574 , \9575 , \9576 , \9580 , \9583 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 , \9592 , \9593 , \9594 , \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 , \9602 , \9603 , \9604 , \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 );
and \U$2979 ( \9613 , RIe5329d0_6883, \9612 );
not \U$2980 ( \9614 , \9573 );
not \U$2981 ( \9615 , \9574 );
not \U$2982 ( \9616 , \9575 );
not \U$2983 ( \9617 , \9576 );
buf \U$2984 ( \9618 , \9586 );
buf \U$2985 ( \9619 , \9586 );
buf \U$2986 ( \9620 , \9586 );
buf \U$2987 ( \9621 , \9586 );
buf \U$2988 ( \9622 , \9586 );
buf \U$2989 ( \9623 , \9586 );
buf \U$2990 ( \9624 , \9586 );
buf \U$2991 ( \9625 , \9586 );
buf \U$2992 ( \9626 , \9586 );
buf \U$2993 ( \9627 , \9586 );
buf \U$2994 ( \9628 , \9586 );
buf \U$2995 ( \9629 , \9586 );
buf \U$2996 ( \9630 , \9586 );
buf \U$2997 ( \9631 , \9586 );
buf \U$2998 ( \9632 , \9586 );
buf \U$2999 ( \9633 , \9586 );
buf \U$3000 ( \9634 , \9586 );
buf \U$3001 ( \9635 , \9586 );
buf \U$3002 ( \9636 , \9586 );
buf \U$3003 ( \9637 , \9586 );
buf \U$3004 ( \9638 , \9586 );
buf \U$3005 ( \9639 , \9586 );
buf \U$3006 ( \9640 , \9586 );
buf \U$3007 ( \9641 , \9586 );
buf \U$3008 ( \9642 , \9586 );
nor \U$3009 ( \9643 , \9614 , \9615 , \9616 , \9617 , \9579 , \9583 , \9586 , \9618 , \9619 , \9620 , \9621 , \9622 , \9623 , \9624 , \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 , \9633 , \9634 , \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 );
and \U$3010 ( \9644 , RIeb72150_6905, \9643 );
buf \U$3011 ( \9645 , \9586 );
buf \U$3012 ( \9646 , \9586 );
buf \U$3013 ( \9647 , \9586 );
buf \U$3014 ( \9648 , \9586 );
buf \U$3015 ( \9649 , \9586 );
buf \U$3016 ( \9650 , \9586 );
buf \U$3017 ( \9651 , \9586 );
buf \U$3018 ( \9652 , \9586 );
buf \U$3019 ( \9653 , \9586 );
buf \U$3020 ( \9654 , \9586 );
buf \U$3021 ( \9655 , \9586 );
buf \U$3022 ( \9656 , \9586 );
buf \U$3023 ( \9657 , \9586 );
buf \U$3024 ( \9658 , \9586 );
buf \U$3025 ( \9659 , \9586 );
buf \U$3026 ( \9660 , \9586 );
buf \U$3027 ( \9661 , \9586 );
buf \U$3028 ( \9662 , \9586 );
buf \U$3029 ( \9663 , \9586 );
buf \U$3030 ( \9664 , \9586 );
buf \U$3031 ( \9665 , \9586 );
buf \U$3032 ( \9666 , \9586 );
buf \U$3033 ( \9667 , \9586 );
buf \U$3034 ( \9668 , \9586 );
buf \U$3035 ( \9669 , \9586 );
nor \U$3036 ( \9670 , \9573 , \9615 , \9616 , \9617 , \9579 , \9583 , \9586 , \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 , \9653 , \9654 , \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 , \9663 , \9664 , \9665 , \9666 , \9667 , \9668 , \9669 );
and \U$3037 ( \9671 , RIeab80c0_6897, \9670 );
buf \U$3038 ( \9672 , \9586 );
buf \U$3039 ( \9673 , \9586 );
buf \U$3040 ( \9674 , \9586 );
buf \U$3041 ( \9675 , \9586 );
buf \U$3042 ( \9676 , \9586 );
buf \U$3043 ( \9677 , \9586 );
buf \U$3044 ( \9678 , \9586 );
buf \U$3045 ( \9679 , \9586 );
buf \U$3046 ( \9680 , \9586 );
buf \U$3047 ( \9681 , \9586 );
buf \U$3048 ( \9682 , \9586 );
buf \U$3049 ( \9683 , \9586 );
buf \U$3050 ( \9684 , \9586 );
buf \U$3051 ( \9685 , \9586 );
buf \U$3052 ( \9686 , \9586 );
buf \U$3053 ( \9687 , \9586 );
buf \U$3054 ( \9688 , \9586 );
buf \U$3055 ( \9689 , \9586 );
buf \U$3056 ( \9690 , \9586 );
buf \U$3057 ( \9691 , \9586 );
buf \U$3058 ( \9692 , \9586 );
buf \U$3059 ( \9693 , \9586 );
buf \U$3060 ( \9694 , \9586 );
buf \U$3061 ( \9695 , \9586 );
buf \U$3062 ( \9696 , \9586 );
nor \U$3063 ( \9697 , \9614 , \9574 , \9616 , \9617 , \9579 , \9583 , \9586 , \9672 , \9673 , \9674 , \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 , \9683 , \9684 , \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 , \9693 , \9694 , \9695 , \9696 );
and \U$3064 ( \9698 , RIe5331c8_6882, \9697 );
buf \U$3065 ( \9699 , \9586 );
buf \U$3066 ( \9700 , \9586 );
buf \U$3067 ( \9701 , \9586 );
buf \U$3068 ( \9702 , \9586 );
buf \U$3069 ( \9703 , \9586 );
buf \U$3070 ( \9704 , \9586 );
buf \U$3071 ( \9705 , \9586 );
buf \U$3072 ( \9706 , \9586 );
buf \U$3073 ( \9707 , \9586 );
buf \U$3074 ( \9708 , \9586 );
buf \U$3075 ( \9709 , \9586 );
buf \U$3076 ( \9710 , \9586 );
buf \U$3077 ( \9711 , \9586 );
buf \U$3078 ( \9712 , \9586 );
buf \U$3079 ( \9713 , \9586 );
buf \U$3080 ( \9714 , \9586 );
buf \U$3081 ( \9715 , \9586 );
buf \U$3082 ( \9716 , \9586 );
buf \U$3083 ( \9717 , \9586 );
buf \U$3084 ( \9718 , \9586 );
buf \U$3085 ( \9719 , \9586 );
buf \U$3086 ( \9720 , \9586 );
buf \U$3087 ( \9721 , \9586 );
buf \U$3088 ( \9722 , \9586 );
buf \U$3089 ( \9723 , \9586 );
nor \U$3090 ( \9724 , \9573 , \9574 , \9616 , \9617 , \9579 , \9583 , \9586 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 , \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 , \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 , \9723 );
and \U$3091 ( \9725 , RIe5339c0_6881, \9724 );
buf \U$3092 ( \9726 , \9586 );
buf \U$3093 ( \9727 , \9586 );
buf \U$3094 ( \9728 , \9586 );
buf \U$3095 ( \9729 , \9586 );
buf \U$3096 ( \9730 , \9586 );
buf \U$3097 ( \9731 , \9586 );
buf \U$3098 ( \9732 , \9586 );
buf \U$3099 ( \9733 , \9586 );
buf \U$3100 ( \9734 , \9586 );
buf \U$3101 ( \9735 , \9586 );
buf \U$3102 ( \9736 , \9586 );
buf \U$3103 ( \9737 , \9586 );
buf \U$3104 ( \9738 , \9586 );
buf \U$3105 ( \9739 , \9586 );
buf \U$3106 ( \9740 , \9586 );
buf \U$3107 ( \9741 , \9586 );
buf \U$3108 ( \9742 , \9586 );
buf \U$3109 ( \9743 , \9586 );
buf \U$3110 ( \9744 , \9586 );
buf \U$3111 ( \9745 , \9586 );
buf \U$3112 ( \9746 , \9586 );
buf \U$3113 ( \9747 , \9586 );
buf \U$3114 ( \9748 , \9586 );
buf \U$3115 ( \9749 , \9586 );
buf \U$3116 ( \9750 , \9586 );
nor \U$3117 ( \9751 , \9614 , \9615 , \9575 , \9617 , \9579 , \9583 , \9586 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 , \9733 , \9734 , \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 , \9745 , \9746 , \9747 , \9748 , \9749 , \9750 );
and \U$3118 ( \9752 , RIeab87c8_6898, \9751 );
buf \U$3119 ( \9753 , \9586 );
buf \U$3120 ( \9754 , \9586 );
buf \U$3121 ( \9755 , \9586 );
buf \U$3122 ( \9756 , \9586 );
buf \U$3123 ( \9757 , \9586 );
buf \U$3124 ( \9758 , \9586 );
buf \U$3125 ( \9759 , \9586 );
buf \U$3126 ( \9760 , \9586 );
buf \U$3127 ( \9761 , \9586 );
buf \U$3128 ( \9762 , \9586 );
buf \U$3129 ( \9763 , \9586 );
buf \U$3130 ( \9764 , \9586 );
buf \U$3131 ( \9765 , \9586 );
buf \U$3132 ( \9766 , \9586 );
buf \U$3133 ( \9767 , \9586 );
buf \U$3134 ( \9768 , \9586 );
buf \U$3135 ( \9769 , \9586 );
buf \U$3136 ( \9770 , \9586 );
buf \U$3137 ( \9771 , \9586 );
buf \U$3138 ( \9772 , \9586 );
buf \U$3139 ( \9773 , \9586 );
buf \U$3140 ( \9774 , \9586 );
buf \U$3141 ( \9775 , \9586 );
buf \U$3142 ( \9776 , \9586 );
buf \U$3143 ( \9777 , \9586 );
nor \U$3144 ( \9778 , \9573 , \9615 , \9575 , \9617 , \9579 , \9583 , \9586 , \9753 , \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 , \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 , \9773 , \9774 , \9775 , \9776 , \9777 );
and \U$3145 ( \9779 , RIe5341b8_6880, \9778 );
buf \U$3146 ( \9780 , \9586 );
buf \U$3147 ( \9781 , \9586 );
buf \U$3148 ( \9782 , \9586 );
buf \U$3149 ( \9783 , \9586 );
buf \U$3150 ( \9784 , \9586 );
buf \U$3151 ( \9785 , \9586 );
buf \U$3152 ( \9786 , \9586 );
buf \U$3153 ( \9787 , \9586 );
buf \U$3154 ( \9788 , \9586 );
buf \U$3155 ( \9789 , \9586 );
buf \U$3156 ( \9790 , \9586 );
buf \U$3157 ( \9791 , \9586 );
buf \U$3158 ( \9792 , \9586 );
buf \U$3159 ( \9793 , \9586 );
buf \U$3160 ( \9794 , \9586 );
buf \U$3161 ( \9795 , \9586 );
buf \U$3162 ( \9796 , \9586 );
buf \U$3163 ( \9797 , \9586 );
buf \U$3164 ( \9798 , \9586 );
buf \U$3165 ( \9799 , \9586 );
buf \U$3166 ( \9800 , \9586 );
buf \U$3167 ( \9801 , \9586 );
buf \U$3168 ( \9802 , \9586 );
buf \U$3169 ( \9803 , \9586 );
buf \U$3170 ( \9804 , \9586 );
nor \U$3171 ( \9805 , \9614 , \9574 , \9575 , \9617 , \9579 , \9583 , \9586 , \9780 , \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 , \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 );
and \U$3172 ( \9806 , RIe5349b0_6879, \9805 );
buf \U$3173 ( \9807 , \9586 );
buf \U$3174 ( \9808 , \9586 );
buf \U$3175 ( \9809 , \9586 );
buf \U$3176 ( \9810 , \9586 );
buf \U$3177 ( \9811 , \9586 );
buf \U$3178 ( \9812 , \9586 );
buf \U$3179 ( \9813 , \9586 );
buf \U$3180 ( \9814 , \9586 );
buf \U$3181 ( \9815 , \9586 );
buf \U$3182 ( \9816 , \9586 );
buf \U$3183 ( \9817 , \9586 );
buf \U$3184 ( \9818 , \9586 );
buf \U$3185 ( \9819 , \9586 );
buf \U$3186 ( \9820 , \9586 );
buf \U$3187 ( \9821 , \9586 );
buf \U$3188 ( \9822 , \9586 );
buf \U$3189 ( \9823 , \9586 );
buf \U$3190 ( \9824 , \9586 );
buf \U$3191 ( \9825 , \9586 );
buf \U$3192 ( \9826 , \9586 );
buf \U$3193 ( \9827 , \9586 );
buf \U$3194 ( \9828 , \9586 );
buf \U$3195 ( \9829 , \9586 );
buf \U$3196 ( \9830 , \9586 );
buf \U$3197 ( \9831 , \9586 );
nor \U$3198 ( \9832 , \9573 , \9574 , \9575 , \9617 , \9579 , \9583 , \9586 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 , \9823 , \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 );
and \U$3199 ( \9833 , RIea94af8_6890, \9832 );
buf \U$3200 ( \9834 , \9586 );
buf \U$3201 ( \9835 , \9586 );
buf \U$3202 ( \9836 , \9586 );
buf \U$3203 ( \9837 , \9586 );
buf \U$3204 ( \9838 , \9586 );
buf \U$3205 ( \9839 , \9586 );
buf \U$3206 ( \9840 , \9586 );
buf \U$3207 ( \9841 , \9586 );
buf \U$3208 ( \9842 , \9586 );
buf \U$3209 ( \9843 , \9586 );
buf \U$3210 ( \9844 , \9586 );
buf \U$3211 ( \9845 , \9586 );
buf \U$3212 ( \9846 , \9586 );
buf \U$3213 ( \9847 , \9586 );
buf \U$3214 ( \9848 , \9586 );
buf \U$3215 ( \9849 , \9586 );
buf \U$3216 ( \9850 , \9586 );
buf \U$3217 ( \9851 , \9586 );
buf \U$3218 ( \9852 , \9586 );
buf \U$3219 ( \9853 , \9586 );
buf \U$3220 ( \9854 , \9586 );
buf \U$3221 ( \9855 , \9586 );
buf \U$3222 ( \9856 , \9586 );
buf \U$3223 ( \9857 , \9586 );
buf \U$3224 ( \9858 , \9586 );
nor \U$3225 ( \9859 , \9614 , \9615 , \9616 , \9576 , \9579 , \9583 , \9586 , \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 , \9855 , \9856 , \9857 , \9858 );
and \U$3226 ( \9860 , RIe5351a8_6878, \9859 );
buf \U$3227 ( \9861 , \9586 );
buf \U$3228 ( \9862 , \9586 );
buf \U$3229 ( \9863 , \9586 );
buf \U$3230 ( \9864 , \9586 );
buf \U$3231 ( \9865 , \9586 );
buf \U$3232 ( \9866 , \9586 );
buf \U$3233 ( \9867 , \9586 );
buf \U$3234 ( \9868 , \9586 );
buf \U$3235 ( \9869 , \9586 );
buf \U$3236 ( \9870 , \9586 );
buf \U$3237 ( \9871 , \9586 );
buf \U$3238 ( \9872 , \9586 );
buf \U$3239 ( \9873 , \9586 );
buf \U$3240 ( \9874 , \9586 );
buf \U$3241 ( \9875 , \9586 );
buf \U$3242 ( \9876 , \9586 );
buf \U$3243 ( \9877 , \9586 );
buf \U$3244 ( \9878 , \9586 );
buf \U$3245 ( \9879 , \9586 );
buf \U$3246 ( \9880 , \9586 );
buf \U$3247 ( \9881 , \9586 );
buf \U$3248 ( \9882 , \9586 );
buf \U$3249 ( \9883 , \9586 );
buf \U$3250 ( \9884 , \9586 );
buf \U$3251 ( \9885 , \9586 );
nor \U$3252 ( \9886 , \9573 , \9615 , \9616 , \9576 , \9579 , \9583 , \9586 , \9861 , \9862 , \9863 , \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 , \9885 );
and \U$3253 ( \9887 , RIe5359a0_6877, \9886 );
buf \U$3254 ( \9888 , \9586 );
buf \U$3255 ( \9889 , \9586 );
buf \U$3256 ( \9890 , \9586 );
buf \U$3257 ( \9891 , \9586 );
buf \U$3258 ( \9892 , \9586 );
buf \U$3259 ( \9893 , \9586 );
buf \U$3260 ( \9894 , \9586 );
buf \U$3261 ( \9895 , \9586 );
buf \U$3262 ( \9896 , \9586 );
buf \U$3263 ( \9897 , \9586 );
buf \U$3264 ( \9898 , \9586 );
buf \U$3265 ( \9899 , \9586 );
buf \U$3266 ( \9900 , \9586 );
buf \U$3267 ( \9901 , \9586 );
buf \U$3268 ( \9902 , \9586 );
buf \U$3269 ( \9903 , \9586 );
buf \U$3270 ( \9904 , \9586 );
buf \U$3271 ( \9905 , \9586 );
buf \U$3272 ( \9906 , \9586 );
buf \U$3273 ( \9907 , \9586 );
buf \U$3274 ( \9908 , \9586 );
buf \U$3275 ( \9909 , \9586 );
buf \U$3276 ( \9910 , \9586 );
buf \U$3277 ( \9911 , \9586 );
buf \U$3278 ( \9912 , \9586 );
nor \U$3279 ( \9913 , \9614 , \9574 , \9616 , \9576 , \9579 , \9583 , \9586 , \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 );
and \U$3280 ( \9914 , RIeab78c8_6895, \9913 );
buf \U$3281 ( \9915 , \9586 );
buf \U$3282 ( \9916 , \9586 );
buf \U$3283 ( \9917 , \9586 );
buf \U$3284 ( \9918 , \9586 );
buf \U$3285 ( \9919 , \9586 );
buf \U$3286 ( \9920 , \9586 );
buf \U$3287 ( \9921 , \9586 );
buf \U$3288 ( \9922 , \9586 );
buf \U$3289 ( \9923 , \9586 );
buf \U$3290 ( \9924 , \9586 );
buf \U$3291 ( \9925 , \9586 );
buf \U$3292 ( \9926 , \9586 );
buf \U$3293 ( \9927 , \9586 );
buf \U$3294 ( \9928 , \9586 );
buf \U$3295 ( \9929 , \9586 );
buf \U$3296 ( \9930 , \9586 );
buf \U$3297 ( \9931 , \9586 );
buf \U$3298 ( \9932 , \9586 );
buf \U$3299 ( \9933 , \9586 );
buf \U$3300 ( \9934 , \9586 );
buf \U$3301 ( \9935 , \9586 );
buf \U$3302 ( \9936 , \9586 );
buf \U$3303 ( \9937 , \9586 );
buf \U$3304 ( \9938 , \9586 );
buf \U$3305 ( \9939 , \9586 );
nor \U$3306 ( \9940 , \9573 , \9574 , \9616 , \9576 , \9579 , \9583 , \9586 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 , \9935 , \9936 , \9937 , \9938 , \9939 );
and \U$3307 ( \9941 , RIeab7d00_6896, \9940 );
buf \U$3308 ( \9942 , \9586 );
buf \U$3309 ( \9943 , \9586 );
buf \U$3310 ( \9944 , \9586 );
buf \U$3311 ( \9945 , \9586 );
buf \U$3312 ( \9946 , \9586 );
buf \U$3313 ( \9947 , \9586 );
buf \U$3314 ( \9948 , \9586 );
buf \U$3315 ( \9949 , \9586 );
buf \U$3316 ( \9950 , \9586 );
buf \U$3317 ( \9951 , \9586 );
buf \U$3318 ( \9952 , \9586 );
buf \U$3319 ( \9953 , \9586 );
buf \U$3320 ( \9954 , \9586 );
buf \U$3321 ( \9955 , \9586 );
buf \U$3322 ( \9956 , \9586 );
buf \U$3323 ( \9957 , \9586 );
buf \U$3324 ( \9958 , \9586 );
buf \U$3325 ( \9959 , \9586 );
buf \U$3326 ( \9960 , \9586 );
buf \U$3327 ( \9961 , \9586 );
buf \U$3328 ( \9962 , \9586 );
buf \U$3329 ( \9963 , \9586 );
buf \U$3330 ( \9964 , \9586 );
buf \U$3331 ( \9965 , \9586 );
buf \U$3332 ( \9966 , \9586 );
nor \U$3333 ( \9967 , \9614 , \9615 , \9575 , \9576 , \9579 , \9583 , \9586 , \9942 , \9943 , \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 , \9965 , \9966 );
and \U$3334 ( \9968 , RIeacfa18_6902, \9967 );
buf \U$3335 ( \9969 , \9586 );
buf \U$3336 ( \9970 , \9586 );
buf \U$3337 ( \9971 , \9586 );
buf \U$3338 ( \9972 , \9586 );
buf \U$3339 ( \9973 , \9586 );
buf \U$3340 ( \9974 , \9586 );
buf \U$3341 ( \9975 , \9586 );
buf \U$3342 ( \9976 , \9586 );
buf \U$3343 ( \9977 , \9586 );
buf \U$3344 ( \9978 , \9586 );
buf \U$3345 ( \9979 , \9586 );
buf \U$3346 ( \9980 , \9586 );
buf \U$3347 ( \9981 , \9586 );
buf \U$3348 ( \9982 , \9586 );
buf \U$3349 ( \9983 , \9586 );
buf \U$3350 ( \9984 , \9586 );
buf \U$3351 ( \9985 , \9586 );
buf \U$3352 ( \9986 , \9586 );
buf \U$3353 ( \9987 , \9586 );
buf \U$3354 ( \9988 , \9586 );
buf \U$3355 ( \9989 , \9586 );
buf \U$3356 ( \9990 , \9586 );
buf \U$3357 ( \9991 , \9586 );
buf \U$3358 ( \9992 , \9586 );
buf \U$3359 ( \9993 , \9586 );
nor \U$3360 ( \9994 , \9573 , \9615 , \9575 , \9576 , \9579 , \9583 , \9586 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 , \9993 );
and \U$3361 ( \9995 , RIeab6518_6891, \9994 );
buf \U$3362 ( \9996 , \9586 );
buf \U$3363 ( \9997 , \9586 );
buf \U$3364 ( \9998 , \9586 );
buf \U$3365 ( \9999 , \9586 );
buf \U$3366 ( \10000 , \9586 );
buf \U$3367 ( \10001 , \9586 );
buf \U$3368 ( \10002 , \9586 );
buf \U$3369 ( \10003 , \9586 );
buf \U$3370 ( \10004 , \9586 );
buf \U$3371 ( \10005 , \9586 );
buf \U$3372 ( \10006 , \9586 );
buf \U$3373 ( \10007 , \9586 );
buf \U$3374 ( \10008 , \9586 );
buf \U$3375 ( \10009 , \9586 );
buf \U$3376 ( \10010 , \9586 );
buf \U$3377 ( \10011 , \9586 );
buf \U$3378 ( \10012 , \9586 );
buf \U$3379 ( \10013 , \9586 );
buf \U$3380 ( \10014 , \9586 );
buf \U$3381 ( \10015 , \9586 );
buf \U$3382 ( \10016 , \9586 );
buf \U$3383 ( \10017 , \9586 );
buf \U$3384 ( \10018 , \9586 );
buf \U$3385 ( \10019 , \9586 );
buf \U$3386 ( \10020 , \9586 );
nor \U$3387 ( \10021 , \9614 , \9574 , \9575 , \9576 , \9579 , \9583 , \9586 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 , \10003 , \10004 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 );
and \U$3388 ( \10022 , RIeb352c8_6904, \10021 );
or \U$3389 ( \10023 , \9613 , \9644 , \9671 , \9698 , \9725 , \9752 , \9779 , \9806 , \9833 , \9860 , \9887 , \9914 , \9941 , \9968 , \9995 , \10022 );
buf \U$3390 ( \10024 , \9586 );
not \U$3391 ( \10025 , \10024 );
buf \U$3392 ( \10026 , \9574 );
buf \U$3393 ( \10027 , \9575 );
buf \U$3394 ( \10028 , \9576 );
buf \U$3395 ( \10029 , \9579 );
buf \U$3396 ( \10030 , \9583 );
buf \U$3397 ( \10031 , \9586 );
buf \U$3398 ( \10032 , \9586 );
buf \U$3399 ( \10033 , \9586 );
buf \U$3400 ( \10034 , \9586 );
buf \U$3401 ( \10035 , \9586 );
buf \U$3402 ( \10036 , \9586 );
buf \U$3403 ( \10037 , \9586 );
buf \U$3404 ( \10038 , \9586 );
buf \U$3405 ( \10039 , \9586 );
buf \U$3406 ( \10040 , \9586 );
buf \U$3407 ( \10041 , \9586 );
buf \U$3408 ( \10042 , \9586 );
buf \U$3409 ( \10043 , \9586 );
buf \U$3410 ( \10044 , \9586 );
buf \U$3411 ( \10045 , \9586 );
buf \U$3412 ( \10046 , \9586 );
buf \U$3413 ( \10047 , \9586 );
buf \U$3414 ( \10048 , \9586 );
buf \U$3415 ( \10049 , \9586 );
buf \U$3416 ( \10050 , \9586 );
buf \U$3417 ( \10051 , \9586 );
buf \U$3418 ( \10052 , \9586 );
buf \U$3419 ( \10053 , \9586 );
buf \U$3420 ( \10054 , \9586 );
buf \U$3421 ( \10055 , \9586 );
buf \U$3422 ( \10056 , \9573 );
or \U$3423 ( \10057 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 , \10055 , \10056 );
nand \U$3424 ( \10058 , \10025 , \10057 );
buf \U$3425 ( \10059 , \10058 );
buf \U$3426 ( \10060 , \9586 );
not \U$3427 ( \10061 , \10060 );
buf \U$3428 ( \10062 , \9583 );
buf \U$3429 ( \10063 , \9586 );
buf \U$3430 ( \10064 , \9586 );
buf \U$3431 ( \10065 , \9586 );
buf \U$3432 ( \10066 , \9586 );
buf \U$3433 ( \10067 , \9586 );
buf \U$3434 ( \10068 , \9586 );
buf \U$3435 ( \10069 , \9586 );
buf \U$3436 ( \10070 , \9586 );
buf \U$3437 ( \10071 , \9586 );
buf \U$3438 ( \10072 , \9586 );
buf \U$3439 ( \10073 , \9586 );
buf \U$3440 ( \10074 , \9586 );
buf \U$3441 ( \10075 , \9586 );
buf \U$3442 ( \10076 , \9586 );
buf \U$3443 ( \10077 , \9586 );
buf \U$3444 ( \10078 , \9586 );
buf \U$3445 ( \10079 , \9586 );
buf \U$3446 ( \10080 , \9586 );
buf \U$3447 ( \10081 , \9586 );
buf \U$3448 ( \10082 , \9586 );
buf \U$3449 ( \10083 , \9586 );
buf \U$3450 ( \10084 , \9586 );
buf \U$3451 ( \10085 , \9586 );
buf \U$3452 ( \10086 , \9586 );
buf \U$3453 ( \10087 , \9586 );
buf \U$3454 ( \10088 , \9579 );
buf \U$3455 ( \10089 , \9573 );
buf \U$3456 ( \10090 , \9574 );
buf \U$3457 ( \10091 , \9575 );
buf \U$3458 ( \10092 , \9576 );
or \U$3459 ( \10093 , \10089 , \10090 , \10091 , \10092 );
and \U$3460 ( \10094 , \10088 , \10093 );
or \U$3461 ( \10095 , \10062 , \10063 , \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 , \10083 , \10084 , \10085 , \10086 , \10087 , \10094 );
and \U$3462 ( \10096 , \10061 , \10095 );
buf \U$3463 ( \10097 , \10096 );
or \U$3464 ( \10098 , \10059 , \10097 );
_DC g3e2d ( \10099_nG3e2d , \10023 , \10098 );
not \U$3465 ( \10100 , \10099_nG3e2d );
buf \U$3466 ( \10101 , RIb7b9608_246);
buf \U$3467 ( \10102 , \9586 );
buf \U$3468 ( \10103 , \9586 );
buf \U$3469 ( \10104 , \9586 );
buf \U$3470 ( \10105 , \9586 );
buf \U$3471 ( \10106 , \9586 );
buf \U$3472 ( \10107 , \9586 );
buf \U$3473 ( \10108 , \9586 );
buf \U$3474 ( \10109 , \9586 );
buf \U$3475 ( \10110 , \9586 );
buf \U$3476 ( \10111 , \9586 );
buf \U$3477 ( \10112 , \9586 );
buf \U$3478 ( \10113 , \9586 );
buf \U$3479 ( \10114 , \9586 );
buf \U$3480 ( \10115 , \9586 );
buf \U$3481 ( \10116 , \9586 );
buf \U$3482 ( \10117 , \9586 );
buf \U$3483 ( \10118 , \9586 );
buf \U$3484 ( \10119 , \9586 );
buf \U$3485 ( \10120 , \9586 );
buf \U$3486 ( \10121 , \9586 );
buf \U$3487 ( \10122 , \9586 );
buf \U$3488 ( \10123 , \9586 );
buf \U$3489 ( \10124 , \9586 );
buf \U$3490 ( \10125 , \9586 );
buf \U$3491 ( \10126 , \9586 );
nor \U$3492 ( \10127 , \9573 , \9574 , \9575 , \9576 , \9580 , \9583 , \9586 , \10102 , \10103 , \10104 , \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 , \10125 , \10126 );
and \U$3493 ( \10128 , \7117 , \10127 );
buf \U$3494 ( \10129 , \9586 );
buf \U$3495 ( \10130 , \9586 );
buf \U$3496 ( \10131 , \9586 );
buf \U$3497 ( \10132 , \9586 );
buf \U$3498 ( \10133 , \9586 );
buf \U$3499 ( \10134 , \9586 );
buf \U$3500 ( \10135 , \9586 );
buf \U$3501 ( \10136 , \9586 );
buf \U$3502 ( \10137 , \9586 );
buf \U$3503 ( \10138 , \9586 );
buf \U$3504 ( \10139 , \9586 );
buf \U$3505 ( \10140 , \9586 );
buf \U$3506 ( \10141 , \9586 );
buf \U$3507 ( \10142 , \9586 );
buf \U$3508 ( \10143 , \9586 );
buf \U$3509 ( \10144 , \9586 );
buf \U$3510 ( \10145 , \9586 );
buf \U$3511 ( \10146 , \9586 );
buf \U$3512 ( \10147 , \9586 );
buf \U$3513 ( \10148 , \9586 );
buf \U$3514 ( \10149 , \9586 );
buf \U$3515 ( \10150 , \9586 );
buf \U$3516 ( \10151 , \9586 );
buf \U$3517 ( \10152 , \9586 );
buf \U$3518 ( \10153 , \9586 );
nor \U$3519 ( \10154 , \9614 , \9615 , \9616 , \9617 , \9579 , \9583 , \9586 , \10129 , \10130 , \10131 , \10132 , \10133 , \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 , \10153 );
and \U$3520 ( \10155 , \7119 , \10154 );
buf \U$3521 ( \10156 , \9586 );
buf \U$3522 ( \10157 , \9586 );
buf \U$3523 ( \10158 , \9586 );
buf \U$3524 ( \10159 , \9586 );
buf \U$3525 ( \10160 , \9586 );
buf \U$3526 ( \10161 , \9586 );
buf \U$3527 ( \10162 , \9586 );
buf \U$3528 ( \10163 , \9586 );
buf \U$3529 ( \10164 , \9586 );
buf \U$3530 ( \10165 , \9586 );
buf \U$3531 ( \10166 , \9586 );
buf \U$3532 ( \10167 , \9586 );
buf \U$3533 ( \10168 , \9586 );
buf \U$3534 ( \10169 , \9586 );
buf \U$3535 ( \10170 , \9586 );
buf \U$3536 ( \10171 , \9586 );
buf \U$3537 ( \10172 , \9586 );
buf \U$3538 ( \10173 , \9586 );
buf \U$3539 ( \10174 , \9586 );
buf \U$3540 ( \10175 , \9586 );
buf \U$3541 ( \10176 , \9586 );
buf \U$3542 ( \10177 , \9586 );
buf \U$3543 ( \10178 , \9586 );
buf \U$3544 ( \10179 , \9586 );
buf \U$3545 ( \10180 , \9586 );
nor \U$3546 ( \10181 , \9573 , \9615 , \9616 , \9617 , \9579 , \9583 , \9586 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 , \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 );
and \U$3547 ( \10182 , \7864 , \10181 );
buf \U$3548 ( \10183 , \9586 );
buf \U$3549 ( \10184 , \9586 );
buf \U$3550 ( \10185 , \9586 );
buf \U$3551 ( \10186 , \9586 );
buf \U$3552 ( \10187 , \9586 );
buf \U$3553 ( \10188 , \9586 );
buf \U$3554 ( \10189 , \9586 );
buf \U$3555 ( \10190 , \9586 );
buf \U$3556 ( \10191 , \9586 );
buf \U$3557 ( \10192 , \9586 );
buf \U$3558 ( \10193 , \9586 );
buf \U$3559 ( \10194 , \9586 );
buf \U$3560 ( \10195 , \9586 );
buf \U$3561 ( \10196 , \9586 );
buf \U$3562 ( \10197 , \9586 );
buf \U$3563 ( \10198 , \9586 );
buf \U$3564 ( \10199 , \9586 );
buf \U$3565 ( \10200 , \9586 );
buf \U$3566 ( \10201 , \9586 );
buf \U$3567 ( \10202 , \9586 );
buf \U$3568 ( \10203 , \9586 );
buf \U$3569 ( \10204 , \9586 );
buf \U$3570 ( \10205 , \9586 );
buf \U$3571 ( \10206 , \9586 );
buf \U$3572 ( \10207 , \9586 );
nor \U$3573 ( \10208 , \9614 , \9574 , \9616 , \9617 , \9579 , \9583 , \9586 , \10183 , \10184 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10207 );
and \U$3574 ( \10209 , \7892 , \10208 );
buf \U$3575 ( \10210 , \9586 );
buf \U$3576 ( \10211 , \9586 );
buf \U$3577 ( \10212 , \9586 );
buf \U$3578 ( \10213 , \9586 );
buf \U$3579 ( \10214 , \9586 );
buf \U$3580 ( \10215 , \9586 );
buf \U$3581 ( \10216 , \9586 );
buf \U$3582 ( \10217 , \9586 );
buf \U$3583 ( \10218 , \9586 );
buf \U$3584 ( \10219 , \9586 );
buf \U$3585 ( \10220 , \9586 );
buf \U$3586 ( \10221 , \9586 );
buf \U$3587 ( \10222 , \9586 );
buf \U$3588 ( \10223 , \9586 );
buf \U$3589 ( \10224 , \9586 );
buf \U$3590 ( \10225 , \9586 );
buf \U$3591 ( \10226 , \9586 );
buf \U$3592 ( \10227 , \9586 );
buf \U$3593 ( \10228 , \9586 );
buf \U$3594 ( \10229 , \9586 );
buf \U$3595 ( \10230 , \9586 );
buf \U$3596 ( \10231 , \9586 );
buf \U$3597 ( \10232 , \9586 );
buf \U$3598 ( \10233 , \9586 );
buf \U$3599 ( \10234 , \9586 );
nor \U$3600 ( \10235 , \9573 , \9574 , \9616 , \9617 , \9579 , \9583 , \9586 , \10210 , \10211 , \10212 , \10213 , \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 );
and \U$3601 ( \10236 , \7920 , \10235 );
buf \U$3602 ( \10237 , \9586 );
buf \U$3603 ( \10238 , \9586 );
buf \U$3604 ( \10239 , \9586 );
buf \U$3605 ( \10240 , \9586 );
buf \U$3606 ( \10241 , \9586 );
buf \U$3607 ( \10242 , \9586 );
buf \U$3608 ( \10243 , \9586 );
buf \U$3609 ( \10244 , \9586 );
buf \U$3610 ( \10245 , \9586 );
buf \U$3611 ( \10246 , \9586 );
buf \U$3612 ( \10247 , \9586 );
buf \U$3613 ( \10248 , \9586 );
buf \U$3614 ( \10249 , \9586 );
buf \U$3615 ( \10250 , \9586 );
buf \U$3616 ( \10251 , \9586 );
buf \U$3617 ( \10252 , \9586 );
buf \U$3618 ( \10253 , \9586 );
buf \U$3619 ( \10254 , \9586 );
buf \U$3620 ( \10255 , \9586 );
buf \U$3621 ( \10256 , \9586 );
buf \U$3622 ( \10257 , \9586 );
buf \U$3623 ( \10258 , \9586 );
buf \U$3624 ( \10259 , \9586 );
buf \U$3625 ( \10260 , \9586 );
buf \U$3626 ( \10261 , \9586 );
nor \U$3627 ( \10262 , \9614 , \9615 , \9575 , \9617 , \9579 , \9583 , \9586 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 , \10243 , \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 );
and \U$3628 ( \10263 , \7948 , \10262 );
buf \U$3629 ( \10264 , \9586 );
buf \U$3630 ( \10265 , \9586 );
buf \U$3631 ( \10266 , \9586 );
buf \U$3632 ( \10267 , \9586 );
buf \U$3633 ( \10268 , \9586 );
buf \U$3634 ( \10269 , \9586 );
buf \U$3635 ( \10270 , \9586 );
buf \U$3636 ( \10271 , \9586 );
buf \U$3637 ( \10272 , \9586 );
buf \U$3638 ( \10273 , \9586 );
buf \U$3639 ( \10274 , \9586 );
buf \U$3640 ( \10275 , \9586 );
buf \U$3641 ( \10276 , \9586 );
buf \U$3642 ( \10277 , \9586 );
buf \U$3643 ( \10278 , \9586 );
buf \U$3644 ( \10279 , \9586 );
buf \U$3645 ( \10280 , \9586 );
buf \U$3646 ( \10281 , \9586 );
buf \U$3647 ( \10282 , \9586 );
buf \U$3648 ( \10283 , \9586 );
buf \U$3649 ( \10284 , \9586 );
buf \U$3650 ( \10285 , \9586 );
buf \U$3651 ( \10286 , \9586 );
buf \U$3652 ( \10287 , \9586 );
buf \U$3653 ( \10288 , \9586 );
nor \U$3654 ( \10289 , \9573 , \9615 , \9575 , \9617 , \9579 , \9583 , \9586 , \10264 , \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 , \10285 , \10286 , \10287 , \10288 );
and \U$3655 ( \10290 , \7976 , \10289 );
buf \U$3656 ( \10291 , \9586 );
buf \U$3657 ( \10292 , \9586 );
buf \U$3658 ( \10293 , \9586 );
buf \U$3659 ( \10294 , \9586 );
buf \U$3660 ( \10295 , \9586 );
buf \U$3661 ( \10296 , \9586 );
buf \U$3662 ( \10297 , \9586 );
buf \U$3663 ( \10298 , \9586 );
buf \U$3664 ( \10299 , \9586 );
buf \U$3665 ( \10300 , \9586 );
buf \U$3666 ( \10301 , \9586 );
buf \U$3667 ( \10302 , \9586 );
buf \U$3668 ( \10303 , \9586 );
buf \U$3669 ( \10304 , \9586 );
buf \U$3670 ( \10305 , \9586 );
buf \U$3671 ( \10306 , \9586 );
buf \U$3672 ( \10307 , \9586 );
buf \U$3673 ( \10308 , \9586 );
buf \U$3674 ( \10309 , \9586 );
buf \U$3675 ( \10310 , \9586 );
buf \U$3676 ( \10311 , \9586 );
buf \U$3677 ( \10312 , \9586 );
buf \U$3678 ( \10313 , \9586 );
buf \U$3679 ( \10314 , \9586 );
buf \U$3680 ( \10315 , \9586 );
nor \U$3681 ( \10316 , \9614 , \9574 , \9575 , \9617 , \9579 , \9583 , \9586 , \10291 , \10292 , \10293 , \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 , \10315 );
and \U$3682 ( \10317 , \8004 , \10316 );
buf \U$3683 ( \10318 , \9586 );
buf \U$3684 ( \10319 , \9586 );
buf \U$3685 ( \10320 , \9586 );
buf \U$3686 ( \10321 , \9586 );
buf \U$3687 ( \10322 , \9586 );
buf \U$3688 ( \10323 , \9586 );
buf \U$3689 ( \10324 , \9586 );
buf \U$3690 ( \10325 , \9586 );
buf \U$3691 ( \10326 , \9586 );
buf \U$3692 ( \10327 , \9586 );
buf \U$3693 ( \10328 , \9586 );
buf \U$3694 ( \10329 , \9586 );
buf \U$3695 ( \10330 , \9586 );
buf \U$3696 ( \10331 , \9586 );
buf \U$3697 ( \10332 , \9586 );
buf \U$3698 ( \10333 , \9586 );
buf \U$3699 ( \10334 , \9586 );
buf \U$3700 ( \10335 , \9586 );
buf \U$3701 ( \10336 , \9586 );
buf \U$3702 ( \10337 , \9586 );
buf \U$3703 ( \10338 , \9586 );
buf \U$3704 ( \10339 , \9586 );
buf \U$3705 ( \10340 , \9586 );
buf \U$3706 ( \10341 , \9586 );
buf \U$3707 ( \10342 , \9586 );
nor \U$3708 ( \10343 , \9573 , \9574 , \9575 , \9617 , \9579 , \9583 , \9586 , \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 );
and \U$3709 ( \10344 , \8032 , \10343 );
buf \U$3710 ( \10345 , \9586 );
buf \U$3711 ( \10346 , \9586 );
buf \U$3712 ( \10347 , \9586 );
buf \U$3713 ( \10348 , \9586 );
buf \U$3714 ( \10349 , \9586 );
buf \U$3715 ( \10350 , \9586 );
buf \U$3716 ( \10351 , \9586 );
buf \U$3717 ( \10352 , \9586 );
buf \U$3718 ( \10353 , \9586 );
buf \U$3719 ( \10354 , \9586 );
buf \U$3720 ( \10355 , \9586 );
buf \U$3721 ( \10356 , \9586 );
buf \U$3722 ( \10357 , \9586 );
buf \U$3723 ( \10358 , \9586 );
buf \U$3724 ( \10359 , \9586 );
buf \U$3725 ( \10360 , \9586 );
buf \U$3726 ( \10361 , \9586 );
buf \U$3727 ( \10362 , \9586 );
buf \U$3728 ( \10363 , \9586 );
buf \U$3729 ( \10364 , \9586 );
buf \U$3730 ( \10365 , \9586 );
buf \U$3731 ( \10366 , \9586 );
buf \U$3732 ( \10367 , \9586 );
buf \U$3733 ( \10368 , \9586 );
buf \U$3734 ( \10369 , \9586 );
nor \U$3735 ( \10370 , \9614 , \9615 , \9616 , \9576 , \9579 , \9583 , \9586 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 , \10365 , \10366 , \10367 , \10368 , \10369 );
and \U$3736 ( \10371 , \8060 , \10370 );
buf \U$3737 ( \10372 , \9586 );
buf \U$3738 ( \10373 , \9586 );
buf \U$3739 ( \10374 , \9586 );
buf \U$3740 ( \10375 , \9586 );
buf \U$3741 ( \10376 , \9586 );
buf \U$3742 ( \10377 , \9586 );
buf \U$3743 ( \10378 , \9586 );
buf \U$3744 ( \10379 , \9586 );
buf \U$3745 ( \10380 , \9586 );
buf \U$3746 ( \10381 , \9586 );
buf \U$3747 ( \10382 , \9586 );
buf \U$3748 ( \10383 , \9586 );
buf \U$3749 ( \10384 , \9586 );
buf \U$3750 ( \10385 , \9586 );
buf \U$3751 ( \10386 , \9586 );
buf \U$3752 ( \10387 , \9586 );
buf \U$3753 ( \10388 , \9586 );
buf \U$3754 ( \10389 , \9586 );
buf \U$3755 ( \10390 , \9586 );
buf \U$3756 ( \10391 , \9586 );
buf \U$3757 ( \10392 , \9586 );
buf \U$3758 ( \10393 , \9586 );
buf \U$3759 ( \10394 , \9586 );
buf \U$3760 ( \10395 , \9586 );
buf \U$3761 ( \10396 , \9586 );
nor \U$3762 ( \10397 , \9573 , \9615 , \9616 , \9576 , \9579 , \9583 , \9586 , \10372 , \10373 , \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 , \10395 , \10396 );
and \U$3763 ( \10398 , \8088 , \10397 );
buf \U$3764 ( \10399 , \9586 );
buf \U$3765 ( \10400 , \9586 );
buf \U$3766 ( \10401 , \9586 );
buf \U$3767 ( \10402 , \9586 );
buf \U$3768 ( \10403 , \9586 );
buf \U$3769 ( \10404 , \9586 );
buf \U$3770 ( \10405 , \9586 );
buf \U$3771 ( \10406 , \9586 );
buf \U$3772 ( \10407 , \9586 );
buf \U$3773 ( \10408 , \9586 );
buf \U$3774 ( \10409 , \9586 );
buf \U$3775 ( \10410 , \9586 );
buf \U$3776 ( \10411 , \9586 );
buf \U$3777 ( \10412 , \9586 );
buf \U$3778 ( \10413 , \9586 );
buf \U$3779 ( \10414 , \9586 );
buf \U$3780 ( \10415 , \9586 );
buf \U$3781 ( \10416 , \9586 );
buf \U$3782 ( \10417 , \9586 );
buf \U$3783 ( \10418 , \9586 );
buf \U$3784 ( \10419 , \9586 );
buf \U$3785 ( \10420 , \9586 );
buf \U$3786 ( \10421 , \9586 );
buf \U$3787 ( \10422 , \9586 );
buf \U$3788 ( \10423 , \9586 );
nor \U$3789 ( \10424 , \9614 , \9574 , \9616 , \9576 , \9579 , \9583 , \9586 , \10399 , \10400 , \10401 , \10402 , \10403 , \10404 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 , \10413 , \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 , \10422 , \10423 );
and \U$3790 ( \10425 , \8116 , \10424 );
buf \U$3791 ( \10426 , \9586 );
buf \U$3792 ( \10427 , \9586 );
buf \U$3793 ( \10428 , \9586 );
buf \U$3794 ( \10429 , \9586 );
buf \U$3795 ( \10430 , \9586 );
buf \U$3796 ( \10431 , \9586 );
buf \U$3797 ( \10432 , \9586 );
buf \U$3798 ( \10433 , \9586 );
buf \U$3799 ( \10434 , \9586 );
buf \U$3800 ( \10435 , \9586 );
buf \U$3801 ( \10436 , \9586 );
buf \U$3802 ( \10437 , \9586 );
buf \U$3803 ( \10438 , \9586 );
buf \U$3804 ( \10439 , \9586 );
buf \U$3805 ( \10440 , \9586 );
buf \U$3806 ( \10441 , \9586 );
buf \U$3807 ( \10442 , \9586 );
buf \U$3808 ( \10443 , \9586 );
buf \U$3809 ( \10444 , \9586 );
buf \U$3810 ( \10445 , \9586 );
buf \U$3811 ( \10446 , \9586 );
buf \U$3812 ( \10447 , \9586 );
buf \U$3813 ( \10448 , \9586 );
buf \U$3814 ( \10449 , \9586 );
buf \U$3815 ( \10450 , \9586 );
nor \U$3816 ( \10451 , \9573 , \9574 , \9616 , \9576 , \9579 , \9583 , \9586 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 );
and \U$3817 ( \10452 , \8144 , \10451 );
buf \U$3818 ( \10453 , \9586 );
buf \U$3819 ( \10454 , \9586 );
buf \U$3820 ( \10455 , \9586 );
buf \U$3821 ( \10456 , \9586 );
buf \U$3822 ( \10457 , \9586 );
buf \U$3823 ( \10458 , \9586 );
buf \U$3824 ( \10459 , \9586 );
buf \U$3825 ( \10460 , \9586 );
buf \U$3826 ( \10461 , \9586 );
buf \U$3827 ( \10462 , \9586 );
buf \U$3828 ( \10463 , \9586 );
buf \U$3829 ( \10464 , \9586 );
buf \U$3830 ( \10465 , \9586 );
buf \U$3831 ( \10466 , \9586 );
buf \U$3832 ( \10467 , \9586 );
buf \U$3833 ( \10468 , \9586 );
buf \U$3834 ( \10469 , \9586 );
buf \U$3835 ( \10470 , \9586 );
buf \U$3836 ( \10471 , \9586 );
buf \U$3837 ( \10472 , \9586 );
buf \U$3838 ( \10473 , \9586 );
buf \U$3839 ( \10474 , \9586 );
buf \U$3840 ( \10475 , \9586 );
buf \U$3841 ( \10476 , \9586 );
buf \U$3842 ( \10477 , \9586 );
nor \U$3843 ( \10478 , \9614 , \9615 , \9575 , \9576 , \9579 , \9583 , \9586 , \10453 , \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 , \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 , \10475 , \10476 , \10477 );
and \U$3844 ( \10479 , \8172 , \10478 );
buf \U$3845 ( \10480 , \9586 );
buf \U$3846 ( \10481 , \9586 );
buf \U$3847 ( \10482 , \9586 );
buf \U$3848 ( \10483 , \9586 );
buf \U$3849 ( \10484 , \9586 );
buf \U$3850 ( \10485 , \9586 );
buf \U$3851 ( \10486 , \9586 );
buf \U$3852 ( \10487 , \9586 );
buf \U$3853 ( \10488 , \9586 );
buf \U$3854 ( \10489 , \9586 );
buf \U$3855 ( \10490 , \9586 );
buf \U$3856 ( \10491 , \9586 );
buf \U$3857 ( \10492 , \9586 );
buf \U$3858 ( \10493 , \9586 );
buf \U$3859 ( \10494 , \9586 );
buf \U$3860 ( \10495 , \9586 );
buf \U$3861 ( \10496 , \9586 );
buf \U$3862 ( \10497 , \9586 );
buf \U$3863 ( \10498 , \9586 );
buf \U$3864 ( \10499 , \9586 );
buf \U$3865 ( \10500 , \9586 );
buf \U$3866 ( \10501 , \9586 );
buf \U$3867 ( \10502 , \9586 );
buf \U$3868 ( \10503 , \9586 );
buf \U$3869 ( \10504 , \9586 );
nor \U$3870 ( \10505 , \9573 , \9615 , \9575 , \9576 , \9579 , \9583 , \9586 , \10480 , \10481 , \10482 , \10483 , \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504 );
and \U$3871 ( \10506 , \8200 , \10505 );
buf \U$3872 ( \10507 , \9586 );
buf \U$3873 ( \10508 , \9586 );
buf \U$3874 ( \10509 , \9586 );
buf \U$3875 ( \10510 , \9586 );
buf \U$3876 ( \10511 , \9586 );
buf \U$3877 ( \10512 , \9586 );
buf \U$3878 ( \10513 , \9586 );
buf \U$3879 ( \10514 , \9586 );
buf \U$3880 ( \10515 , \9586 );
buf \U$3881 ( \10516 , \9586 );
buf \U$3882 ( \10517 , \9586 );
buf \U$3883 ( \10518 , \9586 );
buf \U$3884 ( \10519 , \9586 );
buf \U$3885 ( \10520 , \9586 );
buf \U$3886 ( \10521 , \9586 );
buf \U$3887 ( \10522 , \9586 );
buf \U$3888 ( \10523 , \9586 );
buf \U$3889 ( \10524 , \9586 );
buf \U$3890 ( \10525 , \9586 );
buf \U$3891 ( \10526 , \9586 );
buf \U$3892 ( \10527 , \9586 );
buf \U$3893 ( \10528 , \9586 );
buf \U$3894 ( \10529 , \9586 );
buf \U$3895 ( \10530 , \9586 );
buf \U$3896 ( \10531 , \9586 );
nor \U$3897 ( \10532 , \9614 , \9574 , \9575 , \9576 , \9579 , \9583 , \9586 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 , \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 );
and \U$3898 ( \10533 , \8228 , \10532 );
or \U$3899 ( \10534 , \10128 , \10155 , \10182 , \10209 , \10236 , \10263 , \10290 , \10317 , \10344 , \10371 , \10398 , \10425 , \10452 , \10479 , \10506 , \10533 );
buf \U$3900 ( \10535 , \9586 );
not \U$3901 ( \10536 , \10535 );
buf \U$3902 ( \10537 , \9574 );
buf \U$3903 ( \10538 , \9575 );
buf \U$3904 ( \10539 , \9576 );
buf \U$3905 ( \10540 , \9579 );
buf \U$3906 ( \10541 , \9583 );
buf \U$3907 ( \10542 , \9586 );
buf \U$3908 ( \10543 , \9586 );
buf \U$3909 ( \10544 , \9586 );
buf \U$3910 ( \10545 , \9586 );
buf \U$3911 ( \10546 , \9586 );
buf \U$3912 ( \10547 , \9586 );
buf \U$3913 ( \10548 , \9586 );
buf \U$3914 ( \10549 , \9586 );
buf \U$3915 ( \10550 , \9586 );
buf \U$3916 ( \10551 , \9586 );
buf \U$3917 ( \10552 , \9586 );
buf \U$3918 ( \10553 , \9586 );
buf \U$3919 ( \10554 , \9586 );
buf \U$3920 ( \10555 , \9586 );
buf \U$3921 ( \10556 , \9586 );
buf \U$3922 ( \10557 , \9586 );
buf \U$3923 ( \10558 , \9586 );
buf \U$3924 ( \10559 , \9586 );
buf \U$3925 ( \10560 , \9586 );
buf \U$3926 ( \10561 , \9586 );
buf \U$3927 ( \10562 , \9586 );
buf \U$3928 ( \10563 , \9586 );
buf \U$3929 ( \10564 , \9586 );
buf \U$3930 ( \10565 , \9586 );
buf \U$3931 ( \10566 , \9586 );
buf \U$3932 ( \10567 , \9573 );
or \U$3933 ( \10568 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 , \10553 , \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 , \10563 , \10564 , \10565 , \10566 , \10567 );
nand \U$3934 ( \10569 , \10536 , \10568 );
buf \U$3935 ( \10570 , \10569 );
buf \U$3936 ( \10571 , \9586 );
not \U$3937 ( \10572 , \10571 );
buf \U$3938 ( \10573 , \9583 );
buf \U$3939 ( \10574 , \9586 );
buf \U$3940 ( \10575 , \9586 );
buf \U$3941 ( \10576 , \9586 );
buf \U$3942 ( \10577 , \9586 );
buf \U$3943 ( \10578 , \9586 );
buf \U$3944 ( \10579 , \9586 );
buf \U$3945 ( \10580 , \9586 );
buf \U$3946 ( \10581 , \9586 );
buf \U$3947 ( \10582 , \9586 );
buf \U$3948 ( \10583 , \9586 );
buf \U$3949 ( \10584 , \9586 );
buf \U$3950 ( \10585 , \9586 );
buf \U$3951 ( \10586 , \9586 );
buf \U$3952 ( \10587 , \9586 );
buf \U$3953 ( \10588 , \9586 );
buf \U$3954 ( \10589 , \9586 );
buf \U$3955 ( \10590 , \9586 );
buf \U$3956 ( \10591 , \9586 );
buf \U$3957 ( \10592 , \9586 );
buf \U$3958 ( \10593 , \9586 );
buf \U$3959 ( \10594 , \9586 );
buf \U$3960 ( \10595 , \9586 );
buf \U$3961 ( \10596 , \9586 );
buf \U$3962 ( \10597 , \9586 );
buf \U$3963 ( \10598 , \9586 );
buf \U$3964 ( \10599 , \9579 );
buf \U$3965 ( \10600 , \9573 );
buf \U$3966 ( \10601 , \9574 );
buf \U$3967 ( \10602 , \9575 );
buf \U$3968 ( \10603 , \9576 );
or \U$3969 ( \10604 , \10600 , \10601 , \10602 , \10603 );
and \U$3970 ( \10605 , \10599 , \10604 );
or \U$3971 ( \10606 , \10573 , \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 , \10593 , \10594 , \10595 , \10596 , \10597 , \10598 , \10605 );
and \U$3972 ( \10607 , \10572 , \10606 );
buf \U$3973 ( \10608 , \10607 );
or \U$3974 ( \10609 , \10570 , \10608 );
_DC g402c ( \10610_nG402c , \10534 , \10609 );
buf \U$3975 ( \10611 , \10610_nG402c );
xor \U$3976 ( \10612 , \10101 , \10611 );
buf \U$3977 ( \10613 , RIb7b9590_247);
and \U$3978 ( \10614 , \7126 , \10127 );
and \U$3979 ( \10615 , \7128 , \10154 );
and \U$3980 ( \10616 , \8338 , \10181 );
and \U$3981 ( \10617 , \8340 , \10208 );
and \U$3982 ( \10618 , \8342 , \10235 );
and \U$3983 ( \10619 , \8344 , \10262 );
and \U$3984 ( \10620 , \8346 , \10289 );
and \U$3985 ( \10621 , \8348 , \10316 );
and \U$3986 ( \10622 , \8350 , \10343 );
and \U$3987 ( \10623 , \8352 , \10370 );
and \U$3988 ( \10624 , \8354 , \10397 );
and \U$3989 ( \10625 , \8356 , \10424 );
and \U$3990 ( \10626 , \8358 , \10451 );
and \U$3991 ( \10627 , \8360 , \10478 );
and \U$3992 ( \10628 , \8362 , \10505 );
and \U$3993 ( \10629 , \8364 , \10532 );
or \U$3994 ( \10630 , \10614 , \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 );
_DC g4041 ( \10631_nG4041 , \10630 , \10609 );
buf \U$3995 ( \10632 , \10631_nG4041 );
xor \U$3996 ( \10633 , \10613 , \10632 );
or \U$3997 ( \10634 , \10612 , \10633 );
buf \U$3998 ( \10635 , RIb7b9518_248);
and \U$3999 ( \10636 , \7136 , \10127 );
and \U$4000 ( \10637 , \7138 , \10154 );
and \U$4001 ( \10638 , \8374 , \10181 );
and \U$4002 ( \10639 , \8376 , \10208 );
and \U$4003 ( \10640 , \8378 , \10235 );
and \U$4004 ( \10641 , \8380 , \10262 );
and \U$4005 ( \10642 , \8382 , \10289 );
and \U$4006 ( \10643 , \8384 , \10316 );
and \U$4007 ( \10644 , \8386 , \10343 );
and \U$4008 ( \10645 , \8388 , \10370 );
and \U$4009 ( \10646 , \8390 , \10397 );
and \U$4010 ( \10647 , \8392 , \10424 );
and \U$4011 ( \10648 , \8394 , \10451 );
and \U$4012 ( \10649 , \8396 , \10478 );
and \U$4013 ( \10650 , \8398 , \10505 );
and \U$4014 ( \10651 , \8400 , \10532 );
or \U$4015 ( \10652 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 );
_DC g4057 ( \10653_nG4057 , \10652 , \10609 );
buf \U$4016 ( \10654 , \10653_nG4057 );
xor \U$4017 ( \10655 , \10635 , \10654 );
or \U$4018 ( \10656 , \10634 , \10655 );
buf \U$4019 ( \10657 , RIb7b94a0_249);
and \U$4020 ( \10658 , \7146 , \10127 );
and \U$4021 ( \10659 , \7148 , \10154 );
and \U$4022 ( \10660 , \8410 , \10181 );
and \U$4023 ( \10661 , \8412 , \10208 );
and \U$4024 ( \10662 , \8414 , \10235 );
and \U$4025 ( \10663 , \8416 , \10262 );
and \U$4026 ( \10664 , \8418 , \10289 );
and \U$4027 ( \10665 , \8420 , \10316 );
and \U$4028 ( \10666 , \8422 , \10343 );
and \U$4029 ( \10667 , \8424 , \10370 );
and \U$4030 ( \10668 , \8426 , \10397 );
and \U$4031 ( \10669 , \8428 , \10424 );
and \U$4032 ( \10670 , \8430 , \10451 );
and \U$4033 ( \10671 , \8432 , \10478 );
and \U$4034 ( \10672 , \8434 , \10505 );
and \U$4035 ( \10673 , \8436 , \10532 );
or \U$4036 ( \10674 , \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 , \10673 );
_DC g406d ( \10675_nG406d , \10674 , \10609 );
buf \U$4037 ( \10676 , \10675_nG406d );
xor \U$4038 ( \10677 , \10657 , \10676 );
or \U$4039 ( \10678 , \10656 , \10677 );
buf \U$4040 ( \10679 , RIb7b9428_250);
and \U$4041 ( \10680 , \7156 , \10127 );
and \U$4042 ( \10681 , \7158 , \10154 );
and \U$4043 ( \10682 , \8446 , \10181 );
and \U$4044 ( \10683 , \8448 , \10208 );
and \U$4045 ( \10684 , \8450 , \10235 );
and \U$4046 ( \10685 , \8452 , \10262 );
and \U$4047 ( \10686 , \8454 , \10289 );
and \U$4048 ( \10687 , \8456 , \10316 );
and \U$4049 ( \10688 , \8458 , \10343 );
and \U$4050 ( \10689 , \8460 , \10370 );
and \U$4051 ( \10690 , \8462 , \10397 );
and \U$4052 ( \10691 , \8464 , \10424 );
and \U$4053 ( \10692 , \8466 , \10451 );
and \U$4054 ( \10693 , \8468 , \10478 );
and \U$4055 ( \10694 , \8470 , \10505 );
and \U$4056 ( \10695 , \8472 , \10532 );
or \U$4057 ( \10696 , \10680 , \10681 , \10682 , \10683 , \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 , \10695 );
_DC g4083 ( \10697_nG4083 , \10696 , \10609 );
buf \U$4058 ( \10698 , \10697_nG4083 );
xor \U$4059 ( \10699 , \10679 , \10698 );
or \U$4060 ( \10700 , \10678 , \10699 );
buf \U$4061 ( \10701 , RIb7b93b0_251);
and \U$4062 ( \10702 , \7166 , \10127 );
and \U$4063 ( \10703 , \7168 , \10154 );
and \U$4064 ( \10704 , \8482 , \10181 );
and \U$4065 ( \10705 , \8484 , \10208 );
and \U$4066 ( \10706 , \8486 , \10235 );
and \U$4067 ( \10707 , \8488 , \10262 );
and \U$4068 ( \10708 , \8490 , \10289 );
and \U$4069 ( \10709 , \8492 , \10316 );
and \U$4070 ( \10710 , \8494 , \10343 );
and \U$4071 ( \10711 , \8496 , \10370 );
and \U$4072 ( \10712 , \8498 , \10397 );
and \U$4073 ( \10713 , \8500 , \10424 );
and \U$4074 ( \10714 , \8502 , \10451 );
and \U$4075 ( \10715 , \8504 , \10478 );
and \U$4076 ( \10716 , \8506 , \10505 );
and \U$4077 ( \10717 , \8508 , \10532 );
or \U$4078 ( \10718 , \10702 , \10703 , \10704 , \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 , \10712 , \10713 , \10714 , \10715 , \10716 , \10717 );
_DC g4099 ( \10719_nG4099 , \10718 , \10609 );
buf \U$4079 ( \10720 , \10719_nG4099 );
xor \U$4080 ( \10721 , \10701 , \10720 );
or \U$4081 ( \10722 , \10700 , \10721 );
buf \U$4082 ( \10723 , RIb7af720_252);
and \U$4083 ( \10724 , \7176 , \10127 );
and \U$4084 ( \10725 , \7178 , \10154 );
and \U$4085 ( \10726 , \8518 , \10181 );
and \U$4086 ( \10727 , \8520 , \10208 );
and \U$4087 ( \10728 , \8522 , \10235 );
and \U$4088 ( \10729 , \8524 , \10262 );
and \U$4089 ( \10730 , \8526 , \10289 );
and \U$4090 ( \10731 , \8528 , \10316 );
and \U$4091 ( \10732 , \8530 , \10343 );
and \U$4092 ( \10733 , \8532 , \10370 );
and \U$4093 ( \10734 , \8534 , \10397 );
and \U$4094 ( \10735 , \8536 , \10424 );
and \U$4095 ( \10736 , \8538 , \10451 );
and \U$4096 ( \10737 , \8540 , \10478 );
and \U$4097 ( \10738 , \8542 , \10505 );
and \U$4098 ( \10739 , \8544 , \10532 );
or \U$4099 ( \10740 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 , \10735 , \10736 , \10737 , \10738 , \10739 );
_DC g40af ( \10741_nG40af , \10740 , \10609 );
buf \U$4100 ( \10742 , \10741_nG40af );
xor \U$4101 ( \10743 , \10723 , \10742 );
or \U$4102 ( \10744 , \10722 , \10743 );
buf \U$4103 ( \10745 , RIb7af6a8_253);
and \U$4104 ( \10746 , \7186 , \10127 );
and \U$4105 ( \10747 , \7188 , \10154 );
and \U$4106 ( \10748 , \8554 , \10181 );
and \U$4107 ( \10749 , \8556 , \10208 );
and \U$4108 ( \10750 , \8558 , \10235 );
and \U$4109 ( \10751 , \8560 , \10262 );
and \U$4110 ( \10752 , \8562 , \10289 );
and \U$4111 ( \10753 , \8564 , \10316 );
and \U$4112 ( \10754 , \8566 , \10343 );
and \U$4113 ( \10755 , \8568 , \10370 );
and \U$4114 ( \10756 , \8570 , \10397 );
and \U$4115 ( \10757 , \8572 , \10424 );
and \U$4116 ( \10758 , \8574 , \10451 );
and \U$4117 ( \10759 , \8576 , \10478 );
and \U$4118 ( \10760 , \8578 , \10505 );
and \U$4119 ( \10761 , \8580 , \10532 );
or \U$4120 ( \10762 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 );
_DC g40c5 ( \10763_nG40c5 , \10762 , \10609 );
buf \U$4121 ( \10764 , \10763_nG40c5 );
xor \U$4122 ( \10765 , \10745 , \10764 );
or \U$4123 ( \10766 , \10744 , \10765 );
not \U$4124 ( \10767 , \10766 );
buf \U$4125 ( \10768 , \10767 );
and \U$4126 ( \10769 , \10100 , \10768 );
buf \U$4127 ( \10770 , RIb7af630_254);
buf \U$4128 ( \10771 , \9586 );
buf \U$4129 ( \10772 , \9586 );
buf \U$4130 ( \10773 , \9586 );
buf \U$4131 ( \10774 , \9586 );
buf \U$4132 ( \10775 , \9586 );
buf \U$4133 ( \10776 , \9586 );
buf \U$4134 ( \10777 , \9586 );
buf \U$4135 ( \10778 , \9586 );
buf \U$4136 ( \10779 , \9586 );
buf \U$4137 ( \10780 , \9586 );
buf \U$4138 ( \10781 , \9586 );
buf \U$4139 ( \10782 , \9586 );
buf \U$4140 ( \10783 , \9586 );
buf \U$4141 ( \10784 , \9586 );
buf \U$4142 ( \10785 , \9586 );
buf \U$4143 ( \10786 , \9586 );
buf \U$4144 ( \10787 , \9586 );
buf \U$4145 ( \10788 , \9586 );
buf \U$4146 ( \10789 , \9586 );
buf \U$4147 ( \10790 , \9586 );
buf \U$4148 ( \10791 , \9586 );
buf \U$4149 ( \10792 , \9586 );
buf \U$4150 ( \10793 , \9586 );
buf \U$4151 ( \10794 , \9586 );
buf \U$4152 ( \10795 , \9586 );
nor \U$4153 ( \10796 , \9573 , \9574 , \9575 , \9576 , \9580 , \9583 , \9586 , \10771 , \10772 , \10773 , \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 , \10783 , \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 , \10795 );
and \U$4154 ( \10797 , \7198 , \10796 );
buf \U$4155 ( \10798 , \9586 );
buf \U$4156 ( \10799 , \9586 );
buf \U$4157 ( \10800 , \9586 );
buf \U$4158 ( \10801 , \9586 );
buf \U$4159 ( \10802 , \9586 );
buf \U$4160 ( \10803 , \9586 );
buf \U$4161 ( \10804 , \9586 );
buf \U$4162 ( \10805 , \9586 );
buf \U$4163 ( \10806 , \9586 );
buf \U$4164 ( \10807 , \9586 );
buf \U$4165 ( \10808 , \9586 );
buf \U$4166 ( \10809 , \9586 );
buf \U$4167 ( \10810 , \9586 );
buf \U$4168 ( \10811 , \9586 );
buf \U$4169 ( \10812 , \9586 );
buf \U$4170 ( \10813 , \9586 );
buf \U$4171 ( \10814 , \9586 );
buf \U$4172 ( \10815 , \9586 );
buf \U$4173 ( \10816 , \9586 );
buf \U$4174 ( \10817 , \9586 );
buf \U$4175 ( \10818 , \9586 );
buf \U$4176 ( \10819 , \9586 );
buf \U$4177 ( \10820 , \9586 );
buf \U$4178 ( \10821 , \9586 );
buf \U$4179 ( \10822 , \9586 );
nor \U$4180 ( \10823 , \9614 , \9615 , \9616 , \9617 , \9579 , \9583 , \9586 , \10798 , \10799 , \10800 , \10801 , \10802 , \10803 , \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 );
and \U$4181 ( \10824 , \7200 , \10823 );
buf \U$4182 ( \10825 , \9586 );
buf \U$4183 ( \10826 , \9586 );
buf \U$4184 ( \10827 , \9586 );
buf \U$4185 ( \10828 , \9586 );
buf \U$4186 ( \10829 , \9586 );
buf \U$4187 ( \10830 , \9586 );
buf \U$4188 ( \10831 , \9586 );
buf \U$4189 ( \10832 , \9586 );
buf \U$4190 ( \10833 , \9586 );
buf \U$4191 ( \10834 , \9586 );
buf \U$4192 ( \10835 , \9586 );
buf \U$4193 ( \10836 , \9586 );
buf \U$4194 ( \10837 , \9586 );
buf \U$4195 ( \10838 , \9586 );
buf \U$4196 ( \10839 , \9586 );
buf \U$4197 ( \10840 , \9586 );
buf \U$4198 ( \10841 , \9586 );
buf \U$4199 ( \10842 , \9586 );
buf \U$4200 ( \10843 , \9586 );
buf \U$4201 ( \10844 , \9586 );
buf \U$4202 ( \10845 , \9586 );
buf \U$4203 ( \10846 , \9586 );
buf \U$4204 ( \10847 , \9586 );
buf \U$4205 ( \10848 , \9586 );
buf \U$4206 ( \10849 , \9586 );
nor \U$4207 ( \10850 , \9573 , \9615 , \9616 , \9617 , \9579 , \9583 , \9586 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 , \10845 , \10846 , \10847 , \10848 , \10849 );
and \U$4208 ( \10851 , \8645 , \10850 );
buf \U$4209 ( \10852 , \9586 );
buf \U$4210 ( \10853 , \9586 );
buf \U$4211 ( \10854 , \9586 );
buf \U$4212 ( \10855 , \9586 );
buf \U$4213 ( \10856 , \9586 );
buf \U$4214 ( \10857 , \9586 );
buf \U$4215 ( \10858 , \9586 );
buf \U$4216 ( \10859 , \9586 );
buf \U$4217 ( \10860 , \9586 );
buf \U$4218 ( \10861 , \9586 );
buf \U$4219 ( \10862 , \9586 );
buf \U$4220 ( \10863 , \9586 );
buf \U$4221 ( \10864 , \9586 );
buf \U$4222 ( \10865 , \9586 );
buf \U$4223 ( \10866 , \9586 );
buf \U$4224 ( \10867 , \9586 );
buf \U$4225 ( \10868 , \9586 );
buf \U$4226 ( \10869 , \9586 );
buf \U$4227 ( \10870 , \9586 );
buf \U$4228 ( \10871 , \9586 );
buf \U$4229 ( \10872 , \9586 );
buf \U$4230 ( \10873 , \9586 );
buf \U$4231 ( \10874 , \9586 );
buf \U$4232 ( \10875 , \9586 );
buf \U$4233 ( \10876 , \9586 );
nor \U$4234 ( \10877 , \9614 , \9574 , \9616 , \9617 , \9579 , \9583 , \9586 , \10852 , \10853 , \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 , \10875 , \10876 );
and \U$4235 ( \10878 , \8673 , \10877 );
buf \U$4236 ( \10879 , \9586 );
buf \U$4237 ( \10880 , \9586 );
buf \U$4238 ( \10881 , \9586 );
buf \U$4239 ( \10882 , \9586 );
buf \U$4240 ( \10883 , \9586 );
buf \U$4241 ( \10884 , \9586 );
buf \U$4242 ( \10885 , \9586 );
buf \U$4243 ( \10886 , \9586 );
buf \U$4244 ( \10887 , \9586 );
buf \U$4245 ( \10888 , \9586 );
buf \U$4246 ( \10889 , \9586 );
buf \U$4247 ( \10890 , \9586 );
buf \U$4248 ( \10891 , \9586 );
buf \U$4249 ( \10892 , \9586 );
buf \U$4250 ( \10893 , \9586 );
buf \U$4251 ( \10894 , \9586 );
buf \U$4252 ( \10895 , \9586 );
buf \U$4253 ( \10896 , \9586 );
buf \U$4254 ( \10897 , \9586 );
buf \U$4255 ( \10898 , \9586 );
buf \U$4256 ( \10899 , \9586 );
buf \U$4257 ( \10900 , \9586 );
buf \U$4258 ( \10901 , \9586 );
buf \U$4259 ( \10902 , \9586 );
buf \U$4260 ( \10903 , \9586 );
nor \U$4261 ( \10904 , \9573 , \9574 , \9616 , \9617 , \9579 , \9583 , \9586 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 , \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 , \10903 );
and \U$4262 ( \10905 , \8701 , \10904 );
buf \U$4263 ( \10906 , \9586 );
buf \U$4264 ( \10907 , \9586 );
buf \U$4265 ( \10908 , \9586 );
buf \U$4266 ( \10909 , \9586 );
buf \U$4267 ( \10910 , \9586 );
buf \U$4268 ( \10911 , \9586 );
buf \U$4269 ( \10912 , \9586 );
buf \U$4270 ( \10913 , \9586 );
buf \U$4271 ( \10914 , \9586 );
buf \U$4272 ( \10915 , \9586 );
buf \U$4273 ( \10916 , \9586 );
buf \U$4274 ( \10917 , \9586 );
buf \U$4275 ( \10918 , \9586 );
buf \U$4276 ( \10919 , \9586 );
buf \U$4277 ( \10920 , \9586 );
buf \U$4278 ( \10921 , \9586 );
buf \U$4279 ( \10922 , \9586 );
buf \U$4280 ( \10923 , \9586 );
buf \U$4281 ( \10924 , \9586 );
buf \U$4282 ( \10925 , \9586 );
buf \U$4283 ( \10926 , \9586 );
buf \U$4284 ( \10927 , \9586 );
buf \U$4285 ( \10928 , \9586 );
buf \U$4286 ( \10929 , \9586 );
buf \U$4287 ( \10930 , \9586 );
nor \U$4288 ( \10931 , \9614 , \9615 , \9575 , \9617 , \9579 , \9583 , \9586 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 , \10912 , \10913 , \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 );
and \U$4289 ( \10932 , \8729 , \10931 );
buf \U$4290 ( \10933 , \9586 );
buf \U$4291 ( \10934 , \9586 );
buf \U$4292 ( \10935 , \9586 );
buf \U$4293 ( \10936 , \9586 );
buf \U$4294 ( \10937 , \9586 );
buf \U$4295 ( \10938 , \9586 );
buf \U$4296 ( \10939 , \9586 );
buf \U$4297 ( \10940 , \9586 );
buf \U$4298 ( \10941 , \9586 );
buf \U$4299 ( \10942 , \9586 );
buf \U$4300 ( \10943 , \9586 );
buf \U$4301 ( \10944 , \9586 );
buf \U$4302 ( \10945 , \9586 );
buf \U$4303 ( \10946 , \9586 );
buf \U$4304 ( \10947 , \9586 );
buf \U$4305 ( \10948 , \9586 );
buf \U$4306 ( \10949 , \9586 );
buf \U$4307 ( \10950 , \9586 );
buf \U$4308 ( \10951 , \9586 );
buf \U$4309 ( \10952 , \9586 );
buf \U$4310 ( \10953 , \9586 );
buf \U$4311 ( \10954 , \9586 );
buf \U$4312 ( \10955 , \9586 );
buf \U$4313 ( \10956 , \9586 );
buf \U$4314 ( \10957 , \9586 );
nor \U$4315 ( \10958 , \9573 , \9615 , \9575 , \9617 , \9579 , \9583 , \9586 , \10933 , \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 , \10955 , \10956 , \10957 );
and \U$4316 ( \10959 , \8757 , \10958 );
buf \U$4317 ( \10960 , \9586 );
buf \U$4318 ( \10961 , \9586 );
buf \U$4319 ( \10962 , \9586 );
buf \U$4320 ( \10963 , \9586 );
buf \U$4321 ( \10964 , \9586 );
buf \U$4322 ( \10965 , \9586 );
buf \U$4323 ( \10966 , \9586 );
buf \U$4324 ( \10967 , \9586 );
buf \U$4325 ( \10968 , \9586 );
buf \U$4326 ( \10969 , \9586 );
buf \U$4327 ( \10970 , \9586 );
buf \U$4328 ( \10971 , \9586 );
buf \U$4329 ( \10972 , \9586 );
buf \U$4330 ( \10973 , \9586 );
buf \U$4331 ( \10974 , \9586 );
buf \U$4332 ( \10975 , \9586 );
buf \U$4333 ( \10976 , \9586 );
buf \U$4334 ( \10977 , \9586 );
buf \U$4335 ( \10978 , \9586 );
buf \U$4336 ( \10979 , \9586 );
buf \U$4337 ( \10980 , \9586 );
buf \U$4338 ( \10981 , \9586 );
buf \U$4339 ( \10982 , \9586 );
buf \U$4340 ( \10983 , \9586 );
buf \U$4341 ( \10984 , \9586 );
nor \U$4342 ( \10985 , \9614 , \9574 , \9575 , \9617 , \9579 , \9583 , \9586 , \10960 , \10961 , \10962 , \10963 , \10964 , \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 , \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 , \10982 , \10983 , \10984 );
and \U$4343 ( \10986 , \8785 , \10985 );
buf \U$4344 ( \10987 , \9586 );
buf \U$4345 ( \10988 , \9586 );
buf \U$4346 ( \10989 , \9586 );
buf \U$4347 ( \10990 , \9586 );
buf \U$4348 ( \10991 , \9586 );
buf \U$4349 ( \10992 , \9586 );
buf \U$4350 ( \10993 , \9586 );
buf \U$4351 ( \10994 , \9586 );
buf \U$4352 ( \10995 , \9586 );
buf \U$4353 ( \10996 , \9586 );
buf \U$4354 ( \10997 , \9586 );
buf \U$4355 ( \10998 , \9586 );
buf \U$4356 ( \10999 , \9586 );
buf \U$4357 ( \11000 , \9586 );
buf \U$4358 ( \11001 , \9586 );
buf \U$4359 ( \11002 , \9586 );
buf \U$4360 ( \11003 , \9586 );
buf \U$4361 ( \11004 , \9586 );
buf \U$4362 ( \11005 , \9586 );
buf \U$4363 ( \11006 , \9586 );
buf \U$4364 ( \11007 , \9586 );
buf \U$4365 ( \11008 , \9586 );
buf \U$4366 ( \11009 , \9586 );
buf \U$4367 ( \11010 , \9586 );
buf \U$4368 ( \11011 , \9586 );
nor \U$4369 ( \11012 , \9573 , \9574 , \9575 , \9617 , \9579 , \9583 , \9586 , \10987 , \10988 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 , \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 , \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 );
and \U$4370 ( \11013 , \8813 , \11012 );
buf \U$4371 ( \11014 , \9586 );
buf \U$4372 ( \11015 , \9586 );
buf \U$4373 ( \11016 , \9586 );
buf \U$4374 ( \11017 , \9586 );
buf \U$4375 ( \11018 , \9586 );
buf \U$4376 ( \11019 , \9586 );
buf \U$4377 ( \11020 , \9586 );
buf \U$4378 ( \11021 , \9586 );
buf \U$4379 ( \11022 , \9586 );
buf \U$4380 ( \11023 , \9586 );
buf \U$4381 ( \11024 , \9586 );
buf \U$4382 ( \11025 , \9586 );
buf \U$4383 ( \11026 , \9586 );
buf \U$4384 ( \11027 , \9586 );
buf \U$4385 ( \11028 , \9586 );
buf \U$4386 ( \11029 , \9586 );
buf \U$4387 ( \11030 , \9586 );
buf \U$4388 ( \11031 , \9586 );
buf \U$4389 ( \11032 , \9586 );
buf \U$4390 ( \11033 , \9586 );
buf \U$4391 ( \11034 , \9586 );
buf \U$4392 ( \11035 , \9586 );
buf \U$4393 ( \11036 , \9586 );
buf \U$4394 ( \11037 , \9586 );
buf \U$4395 ( \11038 , \9586 );
nor \U$4396 ( \11039 , \9614 , \9615 , \9616 , \9576 , \9579 , \9583 , \9586 , \11014 , \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 , \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 , \11035 , \11036 , \11037 , \11038 );
and \U$4397 ( \11040 , \8841 , \11039 );
buf \U$4398 ( \11041 , \9586 );
buf \U$4399 ( \11042 , \9586 );
buf \U$4400 ( \11043 , \9586 );
buf \U$4401 ( \11044 , \9586 );
buf \U$4402 ( \11045 , \9586 );
buf \U$4403 ( \11046 , \9586 );
buf \U$4404 ( \11047 , \9586 );
buf \U$4405 ( \11048 , \9586 );
buf \U$4406 ( \11049 , \9586 );
buf \U$4407 ( \11050 , \9586 );
buf \U$4408 ( \11051 , \9586 );
buf \U$4409 ( \11052 , \9586 );
buf \U$4410 ( \11053 , \9586 );
buf \U$4411 ( \11054 , \9586 );
buf \U$4412 ( \11055 , \9586 );
buf \U$4413 ( \11056 , \9586 );
buf \U$4414 ( \11057 , \9586 );
buf \U$4415 ( \11058 , \9586 );
buf \U$4416 ( \11059 , \9586 );
buf \U$4417 ( \11060 , \9586 );
buf \U$4418 ( \11061 , \9586 );
buf \U$4419 ( \11062 , \9586 );
buf \U$4420 ( \11063 , \9586 );
buf \U$4421 ( \11064 , \9586 );
buf \U$4422 ( \11065 , \9586 );
nor \U$4423 ( \11066 , \9573 , \9615 , \9616 , \9576 , \9579 , \9583 , \9586 , \11041 , \11042 , \11043 , \11044 , \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 , \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 , \11065 );
and \U$4424 ( \11067 , \8869 , \11066 );
buf \U$4425 ( \11068 , \9586 );
buf \U$4426 ( \11069 , \9586 );
buf \U$4427 ( \11070 , \9586 );
buf \U$4428 ( \11071 , \9586 );
buf \U$4429 ( \11072 , \9586 );
buf \U$4430 ( \11073 , \9586 );
buf \U$4431 ( \11074 , \9586 );
buf \U$4432 ( \11075 , \9586 );
buf \U$4433 ( \11076 , \9586 );
buf \U$4434 ( \11077 , \9586 );
buf \U$4435 ( \11078 , \9586 );
buf \U$4436 ( \11079 , \9586 );
buf \U$4437 ( \11080 , \9586 );
buf \U$4438 ( \11081 , \9586 );
buf \U$4439 ( \11082 , \9586 );
buf \U$4440 ( \11083 , \9586 );
buf \U$4441 ( \11084 , \9586 );
buf \U$4442 ( \11085 , \9586 );
buf \U$4443 ( \11086 , \9586 );
buf \U$4444 ( \11087 , \9586 );
buf \U$4445 ( \11088 , \9586 );
buf \U$4446 ( \11089 , \9586 );
buf \U$4447 ( \11090 , \9586 );
buf \U$4448 ( \11091 , \9586 );
buf \U$4449 ( \11092 , \9586 );
nor \U$4450 ( \11093 , \9614 , \9574 , \9616 , \9576 , \9579 , \9583 , \9586 , \11068 , \11069 , \11070 , \11071 , \11072 , \11073 , \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 , \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 , \11092 );
and \U$4451 ( \11094 , \8897 , \11093 );
buf \U$4452 ( \11095 , \9586 );
buf \U$4453 ( \11096 , \9586 );
buf \U$4454 ( \11097 , \9586 );
buf \U$4455 ( \11098 , \9586 );
buf \U$4456 ( \11099 , \9586 );
buf \U$4457 ( \11100 , \9586 );
buf \U$4458 ( \11101 , \9586 );
buf \U$4459 ( \11102 , \9586 );
buf \U$4460 ( \11103 , \9586 );
buf \U$4461 ( \11104 , \9586 );
buf \U$4462 ( \11105 , \9586 );
buf \U$4463 ( \11106 , \9586 );
buf \U$4464 ( \11107 , \9586 );
buf \U$4465 ( \11108 , \9586 );
buf \U$4466 ( \11109 , \9586 );
buf \U$4467 ( \11110 , \9586 );
buf \U$4468 ( \11111 , \9586 );
buf \U$4469 ( \11112 , \9586 );
buf \U$4470 ( \11113 , \9586 );
buf \U$4471 ( \11114 , \9586 );
buf \U$4472 ( \11115 , \9586 );
buf \U$4473 ( \11116 , \9586 );
buf \U$4474 ( \11117 , \9586 );
buf \U$4475 ( \11118 , \9586 );
buf \U$4476 ( \11119 , \9586 );
nor \U$4477 ( \11120 , \9573 , \9574 , \9616 , \9576 , \9579 , \9583 , \9586 , \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 , \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 , \11115 , \11116 , \11117 , \11118 , \11119 );
and \U$4478 ( \11121 , \8925 , \11120 );
buf \U$4479 ( \11122 , \9586 );
buf \U$4480 ( \11123 , \9586 );
buf \U$4481 ( \11124 , \9586 );
buf \U$4482 ( \11125 , \9586 );
buf \U$4483 ( \11126 , \9586 );
buf \U$4484 ( \11127 , \9586 );
buf \U$4485 ( \11128 , \9586 );
buf \U$4486 ( \11129 , \9586 );
buf \U$4487 ( \11130 , \9586 );
buf \U$4488 ( \11131 , \9586 );
buf \U$4489 ( \11132 , \9586 );
buf \U$4490 ( \11133 , \9586 );
buf \U$4491 ( \11134 , \9586 );
buf \U$4492 ( \11135 , \9586 );
buf \U$4493 ( \11136 , \9586 );
buf \U$4494 ( \11137 , \9586 );
buf \U$4495 ( \11138 , \9586 );
buf \U$4496 ( \11139 , \9586 );
buf \U$4497 ( \11140 , \9586 );
buf \U$4498 ( \11141 , \9586 );
buf \U$4499 ( \11142 , \9586 );
buf \U$4500 ( \11143 , \9586 );
buf \U$4501 ( \11144 , \9586 );
buf \U$4502 ( \11145 , \9586 );
buf \U$4503 ( \11146 , \9586 );
nor \U$4504 ( \11147 , \9614 , \9615 , \9575 , \9576 , \9579 , \9583 , \9586 , \11122 , \11123 , \11124 , \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 , \11132 , \11133 , \11134 , \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 , \11145 , \11146 );
and \U$4505 ( \11148 , \8953 , \11147 );
buf \U$4506 ( \11149 , \9586 );
buf \U$4507 ( \11150 , \9586 );
buf \U$4508 ( \11151 , \9586 );
buf \U$4509 ( \11152 , \9586 );
buf \U$4510 ( \11153 , \9586 );
buf \U$4511 ( \11154 , \9586 );
buf \U$4512 ( \11155 , \9586 );
buf \U$4513 ( \11156 , \9586 );
buf \U$4514 ( \11157 , \9586 );
buf \U$4515 ( \11158 , \9586 );
buf \U$4516 ( \11159 , \9586 );
buf \U$4517 ( \11160 , \9586 );
buf \U$4518 ( \11161 , \9586 );
buf \U$4519 ( \11162 , \9586 );
buf \U$4520 ( \11163 , \9586 );
buf \U$4521 ( \11164 , \9586 );
buf \U$4522 ( \11165 , \9586 );
buf \U$4523 ( \11166 , \9586 );
buf \U$4524 ( \11167 , \9586 );
buf \U$4525 ( \11168 , \9586 );
buf \U$4526 ( \11169 , \9586 );
buf \U$4527 ( \11170 , \9586 );
buf \U$4528 ( \11171 , \9586 );
buf \U$4529 ( \11172 , \9586 );
buf \U$4530 ( \11173 , \9586 );
nor \U$4531 ( \11174 , \9573 , \9615 , \9575 , \9576 , \9579 , \9583 , \9586 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 , \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 , \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 , \11172 , \11173 );
and \U$4532 ( \11175 , \8981 , \11174 );
buf \U$4533 ( \11176 , \9586 );
buf \U$4534 ( \11177 , \9586 );
buf \U$4535 ( \11178 , \9586 );
buf \U$4536 ( \11179 , \9586 );
buf \U$4537 ( \11180 , \9586 );
buf \U$4538 ( \11181 , \9586 );
buf \U$4539 ( \11182 , \9586 );
buf \U$4540 ( \11183 , \9586 );
buf \U$4541 ( \11184 , \9586 );
buf \U$4542 ( \11185 , \9586 );
buf \U$4543 ( \11186 , \9586 );
buf \U$4544 ( \11187 , \9586 );
buf \U$4545 ( \11188 , \9586 );
buf \U$4546 ( \11189 , \9586 );
buf \U$4547 ( \11190 , \9586 );
buf \U$4548 ( \11191 , \9586 );
buf \U$4549 ( \11192 , \9586 );
buf \U$4550 ( \11193 , \9586 );
buf \U$4551 ( \11194 , \9586 );
buf \U$4552 ( \11195 , \9586 );
buf \U$4553 ( \11196 , \9586 );
buf \U$4554 ( \11197 , \9586 );
buf \U$4555 ( \11198 , \9586 );
buf \U$4556 ( \11199 , \9586 );
buf \U$4557 ( \11200 , \9586 );
nor \U$4558 ( \11201 , \9614 , \9574 , \9575 , \9576 , \9579 , \9583 , \9586 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 , \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 , \11195 , \11196 , \11197 , \11198 , \11199 , \11200 );
and \U$4559 ( \11202 , \9009 , \11201 );
or \U$4560 ( \11203 , \10797 , \10824 , \10851 , \10878 , \10905 , \10932 , \10959 , \10986 , \11013 , \11040 , \11067 , \11094 , \11121 , \11148 , \11175 , \11202 );
buf \U$4561 ( \11204 , \9586 );
not \U$4562 ( \11205 , \11204 );
buf \U$4563 ( \11206 , \9574 );
buf \U$4564 ( \11207 , \9575 );
buf \U$4565 ( \11208 , \9576 );
buf \U$4566 ( \11209 , \9579 );
buf \U$4567 ( \11210 , \9583 );
buf \U$4568 ( \11211 , \9586 );
buf \U$4569 ( \11212 , \9586 );
buf \U$4570 ( \11213 , \9586 );
buf \U$4571 ( \11214 , \9586 );
buf \U$4572 ( \11215 , \9586 );
buf \U$4573 ( \11216 , \9586 );
buf \U$4574 ( \11217 , \9586 );
buf \U$4575 ( \11218 , \9586 );
buf \U$4576 ( \11219 , \9586 );
buf \U$4577 ( \11220 , \9586 );
buf \U$4578 ( \11221 , \9586 );
buf \U$4579 ( \11222 , \9586 );
buf \U$4580 ( \11223 , \9586 );
buf \U$4581 ( \11224 , \9586 );
buf \U$4582 ( \11225 , \9586 );
buf \U$4583 ( \11226 , \9586 );
buf \U$4584 ( \11227 , \9586 );
buf \U$4585 ( \11228 , \9586 );
buf \U$4586 ( \11229 , \9586 );
buf \U$4587 ( \11230 , \9586 );
buf \U$4588 ( \11231 , \9586 );
buf \U$4589 ( \11232 , \9586 );
buf \U$4590 ( \11233 , \9586 );
buf \U$4591 ( \11234 , \9586 );
buf \U$4592 ( \11235 , \9586 );
buf \U$4593 ( \11236 , \9573 );
or \U$4594 ( \11237 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 , \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 , \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 , \11235 , \11236 );
nand \U$4595 ( \11238 , \11205 , \11237 );
buf \U$4596 ( \11239 , \11238 );
buf \U$4597 ( \11240 , \9586 );
not \U$4598 ( \11241 , \11240 );
buf \U$4599 ( \11242 , \9583 );
buf \U$4600 ( \11243 , \9586 );
buf \U$4601 ( \11244 , \9586 );
buf \U$4602 ( \11245 , \9586 );
buf \U$4603 ( \11246 , \9586 );
buf \U$4604 ( \11247 , \9586 );
buf \U$4605 ( \11248 , \9586 );
buf \U$4606 ( \11249 , \9586 );
buf \U$4607 ( \11250 , \9586 );
buf \U$4608 ( \11251 , \9586 );
buf \U$4609 ( \11252 , \9586 );
buf \U$4610 ( \11253 , \9586 );
buf \U$4611 ( \11254 , \9586 );
buf \U$4612 ( \11255 , \9586 );
buf \U$4613 ( \11256 , \9586 );
buf \U$4614 ( \11257 , \9586 );
buf \U$4615 ( \11258 , \9586 );
buf \U$4616 ( \11259 , \9586 );
buf \U$4617 ( \11260 , \9586 );
buf \U$4618 ( \11261 , \9586 );
buf \U$4619 ( \11262 , \9586 );
buf \U$4620 ( \11263 , \9586 );
buf \U$4621 ( \11264 , \9586 );
buf \U$4622 ( \11265 , \9586 );
buf \U$4623 ( \11266 , \9586 );
buf \U$4624 ( \11267 , \9586 );
buf \U$4625 ( \11268 , \9579 );
buf \U$4626 ( \11269 , \9573 );
buf \U$4627 ( \11270 , \9574 );
buf \U$4628 ( \11271 , \9575 );
buf \U$4629 ( \11272 , \9576 );
or \U$4630 ( \11273 , \11269 , \11270 , \11271 , \11272 );
and \U$4631 ( \11274 , \11268 , \11273 );
or \U$4632 ( \11275 , \11242 , \11243 , \11244 , \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 , \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 , \11265 , \11266 , \11267 , \11274 );
and \U$4633 ( \11276 , \11241 , \11275 );
buf \U$4634 ( \11277 , \11276 );
or \U$4635 ( \11278 , \11239 , \11277 );
_DC g42c9 ( \11279_nG42c9 , \11203 , \11278 );
buf \U$4636 ( \11280 , \11279_nG42c9 );
xor \U$4637 ( \11281 , \10770 , \11280 );
buf \U$4638 ( \11282 , RIb7af5b8_255);
and \U$4639 ( \11283 , \7207 , \10796 );
and \U$4640 ( \11284 , \7209 , \10823 );
and \U$4641 ( \11285 , \9119 , \10850 );
and \U$4642 ( \11286 , \9121 , \10877 );
and \U$4643 ( \11287 , \9123 , \10904 );
and \U$4644 ( \11288 , \9125 , \10931 );
and \U$4645 ( \11289 , \9127 , \10958 );
and \U$4646 ( \11290 , \9129 , \10985 );
and \U$4647 ( \11291 , \9131 , \11012 );
and \U$4648 ( \11292 , \9133 , \11039 );
and \U$4649 ( \11293 , \9135 , \11066 );
and \U$4650 ( \11294 , \9137 , \11093 );
and \U$4651 ( \11295 , \9139 , \11120 );
and \U$4652 ( \11296 , \9141 , \11147 );
and \U$4653 ( \11297 , \9143 , \11174 );
and \U$4654 ( \11298 , \9145 , \11201 );
or \U$4655 ( \11299 , \11283 , \11284 , \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 , \11292 , \11293 , \11294 , \11295 , \11296 , \11297 , \11298 );
_DC g42de ( \11300_nG42de , \11299 , \11278 );
buf \U$4656 ( \11301 , \11300_nG42de );
xor \U$4657 ( \11302 , \11282 , \11301 );
or \U$4658 ( \11303 , \11281 , \11302 );
buf \U$4659 ( \11304 , RIb7af540_256);
and \U$4660 ( \11305 , \7217 , \10796 );
and \U$4661 ( \11306 , \7219 , \10823 );
and \U$4662 ( \11307 , \9155 , \10850 );
and \U$4663 ( \11308 , \9157 , \10877 );
and \U$4664 ( \11309 , \9159 , \10904 );
and \U$4665 ( \11310 , \9161 , \10931 );
and \U$4666 ( \11311 , \9163 , \10958 );
and \U$4667 ( \11312 , \9165 , \10985 );
and \U$4668 ( \11313 , \9167 , \11012 );
and \U$4669 ( \11314 , \9169 , \11039 );
and \U$4670 ( \11315 , \9171 , \11066 );
and \U$4671 ( \11316 , \9173 , \11093 );
and \U$4672 ( \11317 , \9175 , \11120 );
and \U$4673 ( \11318 , \9177 , \11147 );
and \U$4674 ( \11319 , \9179 , \11174 );
and \U$4675 ( \11320 , \9181 , \11201 );
or \U$4676 ( \11321 , \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 , \11315 , \11316 , \11317 , \11318 , \11319 , \11320 );
_DC g42f4 ( \11322_nG42f4 , \11321 , \11278 );
buf \U$4677 ( \11323 , \11322_nG42f4 );
xor \U$4678 ( \11324 , \11304 , \11323 );
or \U$4679 ( \11325 , \11303 , \11324 );
buf \U$4680 ( \11326 , RIb7af4c8_257);
and \U$4681 ( \11327 , \7227 , \10796 );
and \U$4682 ( \11328 , \7229 , \10823 );
and \U$4683 ( \11329 , \9191 , \10850 );
and \U$4684 ( \11330 , \9193 , \10877 );
and \U$4685 ( \11331 , \9195 , \10904 );
and \U$4686 ( \11332 , \9197 , \10931 );
and \U$4687 ( \11333 , \9199 , \10958 );
and \U$4688 ( \11334 , \9201 , \10985 );
and \U$4689 ( \11335 , \9203 , \11012 );
and \U$4690 ( \11336 , \9205 , \11039 );
and \U$4691 ( \11337 , \9207 , \11066 );
and \U$4692 ( \11338 , \9209 , \11093 );
and \U$4693 ( \11339 , \9211 , \11120 );
and \U$4694 ( \11340 , \9213 , \11147 );
and \U$4695 ( \11341 , \9215 , \11174 );
and \U$4696 ( \11342 , \9217 , \11201 );
or \U$4697 ( \11343 , \11327 , \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 , \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 , \11342 );
_DC g430a ( \11344_nG430a , \11343 , \11278 );
buf \U$4698 ( \11345 , \11344_nG430a );
xor \U$4699 ( \11346 , \11326 , \11345 );
or \U$4700 ( \11347 , \11325 , \11346 );
buf \U$4701 ( \11348 , RIb7af450_258);
and \U$4702 ( \11349 , \7237 , \10796 );
and \U$4703 ( \11350 , \7239 , \10823 );
and \U$4704 ( \11351 , \9227 , \10850 );
and \U$4705 ( \11352 , \9229 , \10877 );
and \U$4706 ( \11353 , \9231 , \10904 );
and \U$4707 ( \11354 , \9233 , \10931 );
and \U$4708 ( \11355 , \9235 , \10958 );
and \U$4709 ( \11356 , \9237 , \10985 );
and \U$4710 ( \11357 , \9239 , \11012 );
and \U$4711 ( \11358 , \9241 , \11039 );
and \U$4712 ( \11359 , \9243 , \11066 );
and \U$4713 ( \11360 , \9245 , \11093 );
and \U$4714 ( \11361 , \9247 , \11120 );
and \U$4715 ( \11362 , \9249 , \11147 );
and \U$4716 ( \11363 , \9251 , \11174 );
and \U$4717 ( \11364 , \9253 , \11201 );
or \U$4718 ( \11365 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 , \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 );
_DC g4320 ( \11366_nG4320 , \11365 , \11278 );
buf \U$4719 ( \11367 , \11366_nG4320 );
xor \U$4720 ( \11368 , \11348 , \11367 );
or \U$4721 ( \11369 , \11347 , \11368 );
buf \U$4722 ( \11370 , RIb7af3d8_259);
and \U$4723 ( \11371 , \7247 , \10796 );
and \U$4724 ( \11372 , \7249 , \10823 );
and \U$4725 ( \11373 , \9263 , \10850 );
and \U$4726 ( \11374 , \9265 , \10877 );
and \U$4727 ( \11375 , \9267 , \10904 );
and \U$4728 ( \11376 , \9269 , \10931 );
and \U$4729 ( \11377 , \9271 , \10958 );
and \U$4730 ( \11378 , \9273 , \10985 );
and \U$4731 ( \11379 , \9275 , \11012 );
and \U$4732 ( \11380 , \9277 , \11039 );
and \U$4733 ( \11381 , \9279 , \11066 );
and \U$4734 ( \11382 , \9281 , \11093 );
and \U$4735 ( \11383 , \9283 , \11120 );
and \U$4736 ( \11384 , \9285 , \11147 );
and \U$4737 ( \11385 , \9287 , \11174 );
and \U$4738 ( \11386 , \9289 , \11201 );
or \U$4739 ( \11387 , \11371 , \11372 , \11373 , \11374 , \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 , \11385 , \11386 );
_DC g4336 ( \11388_nG4336 , \11387 , \11278 );
buf \U$4740 ( \11389 , \11388_nG4336 );
xor \U$4741 ( \11390 , \11370 , \11389 );
or \U$4742 ( \11391 , \11369 , \11390 );
buf \U$4743 ( \11392 , RIb7a5bf8_260);
and \U$4744 ( \11393 , \7257 , \10796 );
and \U$4745 ( \11394 , \7259 , \10823 );
and \U$4746 ( \11395 , \9299 , \10850 );
and \U$4747 ( \11396 , \9301 , \10877 );
and \U$4748 ( \11397 , \9303 , \10904 );
and \U$4749 ( \11398 , \9305 , \10931 );
and \U$4750 ( \11399 , \9307 , \10958 );
and \U$4751 ( \11400 , \9309 , \10985 );
and \U$4752 ( \11401 , \9311 , \11012 );
and \U$4753 ( \11402 , \9313 , \11039 );
and \U$4754 ( \11403 , \9315 , \11066 );
and \U$4755 ( \11404 , \9317 , \11093 );
and \U$4756 ( \11405 , \9319 , \11120 );
and \U$4757 ( \11406 , \9321 , \11147 );
and \U$4758 ( \11407 , \9323 , \11174 );
and \U$4759 ( \11408 , \9325 , \11201 );
or \U$4760 ( \11409 , \11393 , \11394 , \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 , \11402 , \11403 , \11404 , \11405 , \11406 , \11407 , \11408 );
_DC g434c ( \11410_nG434c , \11409 , \11278 );
buf \U$4761 ( \11411 , \11410_nG434c );
xor \U$4762 ( \11412 , \11392 , \11411 );
or \U$4763 ( \11413 , \11391 , \11412 );
buf \U$4764 ( \11414 , RIb7a0c48_261);
and \U$4765 ( \11415 , \7267 , \10796 );
and \U$4766 ( \11416 , \7269 , \10823 );
and \U$4767 ( \11417 , \9335 , \10850 );
and \U$4768 ( \11418 , \9337 , \10877 );
and \U$4769 ( \11419 , \9339 , \10904 );
and \U$4770 ( \11420 , \9341 , \10931 );
and \U$4771 ( \11421 , \9343 , \10958 );
and \U$4772 ( \11422 , \9345 , \10985 );
and \U$4773 ( \11423 , \9347 , \11012 );
and \U$4774 ( \11424 , \9349 , \11039 );
and \U$4775 ( \11425 , \9351 , \11066 );
and \U$4776 ( \11426 , \9353 , \11093 );
and \U$4777 ( \11427 , \9355 , \11120 );
and \U$4778 ( \11428 , \9357 , \11147 );
and \U$4779 ( \11429 , \9359 , \11174 );
and \U$4780 ( \11430 , \9361 , \11201 );
or \U$4781 ( \11431 , \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 , \11425 , \11426 , \11427 , \11428 , \11429 , \11430 );
_DC g4362 ( \11432_nG4362 , \11431 , \11278 );
buf \U$4782 ( \11433 , \11432_nG4362 );
xor \U$4783 ( \11434 , \11414 , \11433 );
or \U$4784 ( \11435 , \11413 , \11434 );
not \U$4785 ( \11436 , \11435 );
buf \U$4786 ( \11437 , \11436 );
and \U$4787 ( \11438 , \10769 , \11437 );
_HMUX g4369 ( \11439_nG4369 , \9382_nG3b57 , \9573 , \11438 );
buf \U$4788 ( \11440 , \9401 );
buf \U$4789 ( \11441 , \9398 );
buf \U$4790 ( \11442 , \9384 );
buf \U$4791 ( \11443 , \9387 );
buf \U$4792 ( \11444 , \9390 );
buf \U$4793 ( \11445 , \9394 );
or \U$4794 ( \11446 , \11442 , \11443 , \11444 , \11445 );
and \U$4795 ( \11447 , \11441 , \11446 );
or \U$4796 ( \11448 , \11440 , \11447 );
buf \U$4797 ( \11449 , \11448 );
_HMUX g4374 ( \11450_nG4374 , \9572_nG3c16 , \11439_nG4369 , \11449 );
buf \U$4798 ( \11451 , RIe5319e0_6884);
not \U$4799 ( \11452 , \11451 );
buf \U$4800 ( \11453 , \11452 );
buf \U$4801 ( \11454 , RIe549ef0_6842);
xor \U$4802 ( \11455 , \11454 , \11451 );
buf \U$4803 ( \11456 , \11455 );
buf \U$4804 ( \11457 , RIe549770_6843);
and \U$4805 ( \11458 , \11454 , \11451 );
xnor \U$4806 ( \11459 , \11457 , \11458 );
buf \U$4807 ( \11460 , \11459 );
buf \U$4808 ( \11461 , RIe548ff0_6844);
or \U$4809 ( \11462 , \11457 , \11458 );
xnor \U$4810 ( \11463 , \11461 , \11462 );
buf \U$4811 ( \11464 , \11463 );
buf \U$4812 ( \11465 , RIea91330_6888);
or \U$4813 ( \11466 , \11461 , \11462 );
xor \U$4814 ( \11467 , \11465 , \11466 );
buf \U$4815 ( \11468 , \11467 );
not \U$4816 ( \11469 , \11468 );
and \U$4817 ( \11470 , \11465 , \11466 );
buf \U$4818 ( \11471 , \11470 );
nor \U$4819 ( \11472 , \11453 , \11456 , \11460 , \11464 , \11469 , \11471 );
and \U$4820 ( \11473 , RIe5329d0_6883, \11472 );
not \U$4821 ( \11474 , \11471 );
and \U$4822 ( \11475 , \11453 , \11456 , \11460 , \11464 , \11469 , \11474 );
and \U$4823 ( \11476 , RIeb72150_6905, \11475 );
not \U$4824 ( \11477 , \11453 );
and \U$4825 ( \11478 , \11477 , \11456 , \11460 , \11464 , \11469 , \11474 );
and \U$4826 ( \11479 , RIeab80c0_6897, \11478 );
not \U$4827 ( \11480 , \11456 );
and \U$4828 ( \11481 , \11453 , \11480 , \11460 , \11464 , \11469 , \11474 );
and \U$4829 ( \11482 , RIe5331c8_6882, \11481 );
or \U$4842 ( \11483 , \11473 , \11476 , \11479 , \11482 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
buf \U$4844 ( \11484 , \11471 );
buf \U$4845 ( \11485 , \11468 );
buf \U$4846 ( \11486 , \11453 );
buf \U$4847 ( \11487 , \11456 );
buf \U$4848 ( \11488 , \11460 );
buf \U$4849 ( \11489 , \11464 );
or \U$4850 ( \11490 , \11486 , \11487 , \11488 , \11489 );
and \U$4851 ( \11491 , \11485 , \11490 );
or \U$4852 ( \11492 , \11484 , \11491 );
buf \U$4853 ( \11493 , \11492 );
or \U$4854 ( \11494 , 1'b0 , \11493 );
_DC g43a1 ( \11495_nG43a1 , \11483 , \11494 );
not \U$4855 ( \11496 , \11495_nG43a1 );
buf \U$4856 ( \11497 , RIb7b9608_246);
and \U$4857 ( \11498 , \7117 , \11472 );
and \U$4858 ( \11499 , \7119 , \11475 );
and \U$4859 ( \11500 , \7864 , \11478 );
and \U$4860 ( \11501 , \7892 , \11481 );
or \U$4873 ( \11502 , \11498 , \11499 , \11500 , \11501 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g43a9 ( \11503_nG43a9 , \11502 , \11494 );
buf \U$4874 ( \11504 , \11503_nG43a9 );
xor \U$4875 ( \11505 , \11497 , \11504 );
buf \U$4876 ( \11506 , RIb7b9590_247);
and \U$4877 ( \11507 , \7126 , \11472 );
and \U$4878 ( \11508 , \7128 , \11475 );
and \U$4879 ( \11509 , \8338 , \11478 );
and \U$4880 ( \11510 , \8340 , \11481 );
or \U$4893 ( \11511 , \11507 , \11508 , \11509 , \11510 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g43b2 ( \11512_nG43b2 , \11511 , \11494 );
buf \U$4894 ( \11513 , \11512_nG43b2 );
xor \U$4895 ( \11514 , \11506 , \11513 );
or \U$4896 ( \11515 , \11505 , \11514 );
buf \U$4897 ( \11516 , RIb7b9518_248);
and \U$4898 ( \11517 , \7136 , \11472 );
and \U$4899 ( \11518 , \7138 , \11475 );
and \U$4900 ( \11519 , \8374 , \11478 );
and \U$4901 ( \11520 , \8376 , \11481 );
or \U$4914 ( \11521 , \11517 , \11518 , \11519 , \11520 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g43bc ( \11522_nG43bc , \11521 , \11494 );
buf \U$4915 ( \11523 , \11522_nG43bc );
xor \U$4916 ( \11524 , \11516 , \11523 );
or \U$4917 ( \11525 , \11515 , \11524 );
buf \U$4918 ( \11526 , RIb7b94a0_249);
and \U$4919 ( \11527 , \7146 , \11472 );
and \U$4920 ( \11528 , \7148 , \11475 );
and \U$4921 ( \11529 , \8410 , \11478 );
and \U$4922 ( \11530 , \8412 , \11481 );
or \U$4935 ( \11531 , \11527 , \11528 , \11529 , \11530 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g43c6 ( \11532_nG43c6 , \11531 , \11494 );
buf \U$4936 ( \11533 , \11532_nG43c6 );
xor \U$4937 ( \11534 , \11526 , \11533 );
or \U$4938 ( \11535 , \11525 , \11534 );
buf \U$4939 ( \11536 , RIb7b9428_250);
and \U$4940 ( \11537 , \7156 , \11472 );
and \U$4941 ( \11538 , \7158 , \11475 );
and \U$4942 ( \11539 , \8446 , \11478 );
and \U$4943 ( \11540 , \8448 , \11481 );
or \U$4956 ( \11541 , \11537 , \11538 , \11539 , \11540 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g43d0 ( \11542_nG43d0 , \11541 , \11494 );
buf \U$4957 ( \11543 , \11542_nG43d0 );
xor \U$4958 ( \11544 , \11536 , \11543 );
or \U$4959 ( \11545 , \11535 , \11544 );
buf \U$4960 ( \11546 , RIb7b93b0_251);
and \U$4961 ( \11547 , \7166 , \11472 );
and \U$4962 ( \11548 , \7168 , \11475 );
and \U$4963 ( \11549 , \8482 , \11478 );
and \U$4964 ( \11550 , \8484 , \11481 );
or \U$4977 ( \11551 , \11547 , \11548 , \11549 , \11550 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g43da ( \11552_nG43da , \11551 , \11494 );
buf \U$4978 ( \11553 , \11552_nG43da );
xor \U$4979 ( \11554 , \11546 , \11553 );
or \U$4980 ( \11555 , \11545 , \11554 );
buf \U$4981 ( \11556 , RIb7af720_252);
and \U$4982 ( \11557 , \7176 , \11472 );
and \U$4983 ( \11558 , \7178 , \11475 );
and \U$4984 ( \11559 , \8518 , \11478 );
and \U$4985 ( \11560 , \8520 , \11481 );
or \U$4998 ( \11561 , \11557 , \11558 , \11559 , \11560 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g43e4 ( \11562_nG43e4 , \11561 , \11494 );
buf \U$4999 ( \11563 , \11562_nG43e4 );
xor \U$5000 ( \11564 , \11556 , \11563 );
or \U$5001 ( \11565 , \11555 , \11564 );
buf \U$5002 ( \11566 , RIb7af6a8_253);
and \U$5003 ( \11567 , \7186 , \11472 );
and \U$5004 ( \11568 , \7188 , \11475 );
and \U$5005 ( \11569 , \8554 , \11478 );
and \U$5006 ( \11570 , \8556 , \11481 );
or \U$5019 ( \11571 , \11567 , \11568 , \11569 , \11570 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g43ee ( \11572_nG43ee , \11571 , \11494 );
buf \U$5020 ( \11573 , \11572_nG43ee );
xor \U$5021 ( \11574 , \11566 , \11573 );
or \U$5022 ( \11575 , \11565 , \11574 );
not \U$5023 ( \11576 , \11575 );
buf \U$5024 ( \11577 , \11576 );
buf \U$5025 ( \11578 , RIb7af630_254);
and \U$5026 ( \11579 , \7198 , \11472 );
and \U$5027 ( \11580 , \7200 , \11475 );
and \U$5028 ( \11581 , \8645 , \11478 );
and \U$5029 ( \11582 , \8673 , \11481 );
or \U$5042 ( \11583 , \11579 , \11580 , \11581 , \11582 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g43fa ( \11584_nG43fa , \11583 , \11494 );
buf \U$5043 ( \11585 , \11584_nG43fa );
xor \U$5044 ( \11586 , \11578 , \11585 );
buf \U$5045 ( \11587 , RIb7af5b8_255);
and \U$5046 ( \11588 , \7207 , \11472 );
and \U$5047 ( \11589 , \7209 , \11475 );
and \U$5048 ( \11590 , \9119 , \11478 );
and \U$5049 ( \11591 , \9121 , \11481 );
or \U$5062 ( \11592 , \11588 , \11589 , \11590 , \11591 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4403 ( \11593_nG4403 , \11592 , \11494 );
buf \U$5063 ( \11594 , \11593_nG4403 );
xor \U$5064 ( \11595 , \11587 , \11594 );
or \U$5065 ( \11596 , \11586 , \11595 );
buf \U$5066 ( \11597 , RIb7af540_256);
and \U$5067 ( \11598 , \7217 , \11472 );
and \U$5068 ( \11599 , \7219 , \11475 );
and \U$5069 ( \11600 , \9155 , \11478 );
and \U$5070 ( \11601 , \9157 , \11481 );
or \U$5083 ( \11602 , \11598 , \11599 , \11600 , \11601 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g440d ( \11603_nG440d , \11602 , \11494 );
buf \U$5084 ( \11604 , \11603_nG440d );
xor \U$5085 ( \11605 , \11597 , \11604 );
or \U$5086 ( \11606 , \11596 , \11605 );
buf \U$5087 ( \11607 , RIb7af4c8_257);
and \U$5088 ( \11608 , \7227 , \11472 );
and \U$5089 ( \11609 , \7229 , \11475 );
and \U$5090 ( \11610 , \9191 , \11478 );
and \U$5091 ( \11611 , \9193 , \11481 );
or \U$5104 ( \11612 , \11608 , \11609 , \11610 , \11611 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4417 ( \11613_nG4417 , \11612 , \11494 );
buf \U$5105 ( \11614 , \11613_nG4417 );
xor \U$5106 ( \11615 , \11607 , \11614 );
or \U$5107 ( \11616 , \11606 , \11615 );
buf \U$5108 ( \11617 , RIb7af450_258);
and \U$5109 ( \11618 , \7237 , \11472 );
and \U$5110 ( \11619 , \7239 , \11475 );
and \U$5111 ( \11620 , \9227 , \11478 );
and \U$5112 ( \11621 , \9229 , \11481 );
or \U$5125 ( \11622 , \11618 , \11619 , \11620 , \11621 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4421 ( \11623_nG4421 , \11622 , \11494 );
buf \U$5126 ( \11624 , \11623_nG4421 );
xor \U$5127 ( \11625 , \11617 , \11624 );
or \U$5128 ( \11626 , \11616 , \11625 );
buf \U$5129 ( \11627 , RIb7af3d8_259);
and \U$5130 ( \11628 , \7247 , \11472 );
and \U$5131 ( \11629 , \7249 , \11475 );
and \U$5132 ( \11630 , \9263 , \11478 );
and \U$5133 ( \11631 , \9265 , \11481 );
or \U$5146 ( \11632 , \11628 , \11629 , \11630 , \11631 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g442b ( \11633_nG442b , \11632 , \11494 );
buf \U$5147 ( \11634 , \11633_nG442b );
xor \U$5148 ( \11635 , \11627 , \11634 );
or \U$5149 ( \11636 , \11626 , \11635 );
buf \U$5150 ( \11637 , RIb7a5bf8_260);
and \U$5151 ( \11638 , \7257 , \11472 );
and \U$5152 ( \11639 , \7259 , \11475 );
and \U$5153 ( \11640 , \9299 , \11478 );
and \U$5154 ( \11641 , \9301 , \11481 );
or \U$5167 ( \11642 , \11638 , \11639 , \11640 , \11641 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4435 ( \11643_nG4435 , \11642 , \11494 );
buf \U$5168 ( \11644 , \11643_nG4435 );
xor \U$5169 ( \11645 , \11637 , \11644 );
or \U$5170 ( \11646 , \11636 , \11645 );
buf \U$5171 ( \11647 , RIb7a0c48_261);
and \U$5172 ( \11648 , \7267 , \11472 );
and \U$5173 ( \11649 , \7269 , \11475 );
and \U$5174 ( \11650 , \9335 , \11478 );
and \U$5175 ( \11651 , \9337 , \11481 );
or \U$5188 ( \11652 , \11648 , \11649 , \11650 , \11651 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g443f ( \11653_nG443f , \11652 , \11494 );
buf \U$5189 ( \11654 , \11653_nG443f );
xor \U$5190 ( \11655 , \11647 , \11654 );
or \U$5191 ( \11656 , \11646 , \11655 );
not \U$5192 ( \11657 , \11656 );
buf \U$5193 ( \11658 , \11657 );
and \U$5194 ( \11659 , \11577 , \11658 );
and \U$5195 ( \11660 , \11496 , \11659 );
_HMUX g4447 ( \11661_nG4447 , \11450_nG4374 , \11453 , \11660 );
buf \U$5198 ( \11662 , \11453 );
buf \U$5201 ( \11663 , \11456 );
buf \U$5204 ( \11664 , \11460 );
buf \U$5207 ( \11665 , \11464 );
buf \U$5208 ( \11666 , \11468 );
not \U$5209 ( \11667 , \11666 );
buf \U$5210 ( \11668 , \11667 );
not \U$5211 ( \11669 , \11668 );
buf \U$5212 ( \11670 , \11471 );
xnor \U$5213 ( \11671 , \11670 , \11666 );
buf \U$5214 ( \11672 , \11671 );
or \U$5215 ( \11673 , \11670 , \11666 );
not \U$5216 ( \11674 , \11673 );
buf \U$5217 ( \11675 , \11674 );
buf \U$5218 ( \11676 , \11675 );
buf \U$5219 ( \11677 , \11675 );
buf \U$5220 ( \11678 , \11675 );
buf \U$5221 ( \11679 , \11675 );
buf \U$5222 ( \11680 , \11675 );
buf \U$5223 ( \11681 , \11675 );
buf \U$5224 ( \11682 , \11675 );
buf \U$5225 ( \11683 , \11675 );
buf \U$5226 ( \11684 , \11675 );
buf \U$5227 ( \11685 , \11675 );
buf \U$5228 ( \11686 , \11675 );
buf \U$5229 ( \11687 , \11675 );
buf \U$5230 ( \11688 , \11675 );
buf \U$5231 ( \11689 , \11675 );
buf \U$5232 ( \11690 , \11675 );
buf \U$5233 ( \11691 , \11675 );
buf \U$5234 ( \11692 , \11675 );
buf \U$5235 ( \11693 , \11675 );
buf \U$5236 ( \11694 , \11675 );
buf \U$5237 ( \11695 , \11675 );
buf \U$5238 ( \11696 , \11675 );
buf \U$5239 ( \11697 , \11675 );
buf \U$5240 ( \11698 , \11675 );
buf \U$5241 ( \11699 , \11675 );
buf \U$5242 ( \11700 , \11675 );
nor \U$5243 ( \11701 , \11662 , \11663 , \11664 , \11665 , \11669 , \11672 , \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 , \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 , \11692 , \11693 , \11694 , \11695 , \11696 , \11697 , \11698 , \11699 , \11700 );
and \U$5244 ( \11702 , RIe5329d0_6883, \11701 );
not \U$5245 ( \11703 , \11662 );
not \U$5246 ( \11704 , \11663 );
not \U$5247 ( \11705 , \11664 );
not \U$5248 ( \11706 , \11665 );
buf \U$5249 ( \11707 , \11675 );
buf \U$5250 ( \11708 , \11675 );
buf \U$5251 ( \11709 , \11675 );
buf \U$5252 ( \11710 , \11675 );
buf \U$5253 ( \11711 , \11675 );
buf \U$5254 ( \11712 , \11675 );
buf \U$5255 ( \11713 , \11675 );
buf \U$5256 ( \11714 , \11675 );
buf \U$5257 ( \11715 , \11675 );
buf \U$5258 ( \11716 , \11675 );
buf \U$5259 ( \11717 , \11675 );
buf \U$5260 ( \11718 , \11675 );
buf \U$5261 ( \11719 , \11675 );
buf \U$5262 ( \11720 , \11675 );
buf \U$5263 ( \11721 , \11675 );
buf \U$5264 ( \11722 , \11675 );
buf \U$5265 ( \11723 , \11675 );
buf \U$5266 ( \11724 , \11675 );
buf \U$5267 ( \11725 , \11675 );
buf \U$5268 ( \11726 , \11675 );
buf \U$5269 ( \11727 , \11675 );
buf \U$5270 ( \11728 , \11675 );
buf \U$5271 ( \11729 , \11675 );
buf \U$5272 ( \11730 , \11675 );
buf \U$5273 ( \11731 , \11675 );
nor \U$5274 ( \11732 , \11703 , \11704 , \11705 , \11706 , \11668 , \11672 , \11675 , \11707 , \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 , \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 , \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 );
and \U$5275 ( \11733 , RIeb72150_6905, \11732 );
buf \U$5276 ( \11734 , \11675 );
buf \U$5277 ( \11735 , \11675 );
buf \U$5278 ( \11736 , \11675 );
buf \U$5279 ( \11737 , \11675 );
buf \U$5280 ( \11738 , \11675 );
buf \U$5281 ( \11739 , \11675 );
buf \U$5282 ( \11740 , \11675 );
buf \U$5283 ( \11741 , \11675 );
buf \U$5284 ( \11742 , \11675 );
buf \U$5285 ( \11743 , \11675 );
buf \U$5286 ( \11744 , \11675 );
buf \U$5287 ( \11745 , \11675 );
buf \U$5288 ( \11746 , \11675 );
buf \U$5289 ( \11747 , \11675 );
buf \U$5290 ( \11748 , \11675 );
buf \U$5291 ( \11749 , \11675 );
buf \U$5292 ( \11750 , \11675 );
buf \U$5293 ( \11751 , \11675 );
buf \U$5294 ( \11752 , \11675 );
buf \U$5295 ( \11753 , \11675 );
buf \U$5296 ( \11754 , \11675 );
buf \U$5297 ( \11755 , \11675 );
buf \U$5298 ( \11756 , \11675 );
buf \U$5299 ( \11757 , \11675 );
buf \U$5300 ( \11758 , \11675 );
nor \U$5301 ( \11759 , \11662 , \11704 , \11705 , \11706 , \11668 , \11672 , \11675 , \11734 , \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 , \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 , \11755 , \11756 , \11757 , \11758 );
and \U$5302 ( \11760 , RIeab80c0_6897, \11759 );
buf \U$5303 ( \11761 , \11675 );
buf \U$5304 ( \11762 , \11675 );
buf \U$5305 ( \11763 , \11675 );
buf \U$5306 ( \11764 , \11675 );
buf \U$5307 ( \11765 , \11675 );
buf \U$5308 ( \11766 , \11675 );
buf \U$5309 ( \11767 , \11675 );
buf \U$5310 ( \11768 , \11675 );
buf \U$5311 ( \11769 , \11675 );
buf \U$5312 ( \11770 , \11675 );
buf \U$5313 ( \11771 , \11675 );
buf \U$5314 ( \11772 , \11675 );
buf \U$5315 ( \11773 , \11675 );
buf \U$5316 ( \11774 , \11675 );
buf \U$5317 ( \11775 , \11675 );
buf \U$5318 ( \11776 , \11675 );
buf \U$5319 ( \11777 , \11675 );
buf \U$5320 ( \11778 , \11675 );
buf \U$5321 ( \11779 , \11675 );
buf \U$5322 ( \11780 , \11675 );
buf \U$5323 ( \11781 , \11675 );
buf \U$5324 ( \11782 , \11675 );
buf \U$5325 ( \11783 , \11675 );
buf \U$5326 ( \11784 , \11675 );
buf \U$5327 ( \11785 , \11675 );
nor \U$5328 ( \11786 , \11703 , \11663 , \11705 , \11706 , \11668 , \11672 , \11675 , \11761 , \11762 , \11763 , \11764 , \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 , \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 , \11782 , \11783 , \11784 , \11785 );
and \U$5329 ( \11787 , RIe5331c8_6882, \11786 );
buf \U$5330 ( \11788 , \11675 );
buf \U$5331 ( \11789 , \11675 );
buf \U$5332 ( \11790 , \11675 );
buf \U$5333 ( \11791 , \11675 );
buf \U$5334 ( \11792 , \11675 );
buf \U$5335 ( \11793 , \11675 );
buf \U$5336 ( \11794 , \11675 );
buf \U$5337 ( \11795 , \11675 );
buf \U$5338 ( \11796 , \11675 );
buf \U$5339 ( \11797 , \11675 );
buf \U$5340 ( \11798 , \11675 );
buf \U$5341 ( \11799 , \11675 );
buf \U$5342 ( \11800 , \11675 );
buf \U$5343 ( \11801 , \11675 );
buf \U$5344 ( \11802 , \11675 );
buf \U$5345 ( \11803 , \11675 );
buf \U$5346 ( \11804 , \11675 );
buf \U$5347 ( \11805 , \11675 );
buf \U$5348 ( \11806 , \11675 );
buf \U$5349 ( \11807 , \11675 );
buf \U$5350 ( \11808 , \11675 );
buf \U$5351 ( \11809 , \11675 );
buf \U$5352 ( \11810 , \11675 );
buf \U$5353 ( \11811 , \11675 );
buf \U$5354 ( \11812 , \11675 );
nor \U$5355 ( \11813 , \11662 , \11663 , \11705 , \11706 , \11668 , \11672 , \11675 , \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 , \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 , \11802 , \11803 , \11804 , \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 , \11812 );
and \U$5356 ( \11814 , RIe5339c0_6881, \11813 );
buf \U$5357 ( \11815 , \11675 );
buf \U$5358 ( \11816 , \11675 );
buf \U$5359 ( \11817 , \11675 );
buf \U$5360 ( \11818 , \11675 );
buf \U$5361 ( \11819 , \11675 );
buf \U$5362 ( \11820 , \11675 );
buf \U$5363 ( \11821 , \11675 );
buf \U$5364 ( \11822 , \11675 );
buf \U$5365 ( \11823 , \11675 );
buf \U$5366 ( \11824 , \11675 );
buf \U$5367 ( \11825 , \11675 );
buf \U$5368 ( \11826 , \11675 );
buf \U$5369 ( \11827 , \11675 );
buf \U$5370 ( \11828 , \11675 );
buf \U$5371 ( \11829 , \11675 );
buf \U$5372 ( \11830 , \11675 );
buf \U$5373 ( \11831 , \11675 );
buf \U$5374 ( \11832 , \11675 );
buf \U$5375 ( \11833 , \11675 );
buf \U$5376 ( \11834 , \11675 );
buf \U$5377 ( \11835 , \11675 );
buf \U$5378 ( \11836 , \11675 );
buf \U$5379 ( \11837 , \11675 );
buf \U$5380 ( \11838 , \11675 );
buf \U$5381 ( \11839 , \11675 );
nor \U$5382 ( \11840 , \11703 , \11704 , \11664 , \11706 , \11668 , \11672 , \11675 , \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 , \11822 , \11823 , \11824 , \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 , \11832 , \11833 , \11834 , \11835 , \11836 , \11837 , \11838 , \11839 );
and \U$5383 ( \11841 , RIeab87c8_6898, \11840 );
buf \U$5384 ( \11842 , \11675 );
buf \U$5385 ( \11843 , \11675 );
buf \U$5386 ( \11844 , \11675 );
buf \U$5387 ( \11845 , \11675 );
buf \U$5388 ( \11846 , \11675 );
buf \U$5389 ( \11847 , \11675 );
buf \U$5390 ( \11848 , \11675 );
buf \U$5391 ( \11849 , \11675 );
buf \U$5392 ( \11850 , \11675 );
buf \U$5393 ( \11851 , \11675 );
buf \U$5394 ( \11852 , \11675 );
buf \U$5395 ( \11853 , \11675 );
buf \U$5396 ( \11854 , \11675 );
buf \U$5397 ( \11855 , \11675 );
buf \U$5398 ( \11856 , \11675 );
buf \U$5399 ( \11857 , \11675 );
buf \U$5400 ( \11858 , \11675 );
buf \U$5401 ( \11859 , \11675 );
buf \U$5402 ( \11860 , \11675 );
buf \U$5403 ( \11861 , \11675 );
buf \U$5404 ( \11862 , \11675 );
buf \U$5405 ( \11863 , \11675 );
buf \U$5406 ( \11864 , \11675 );
buf \U$5407 ( \11865 , \11675 );
buf \U$5408 ( \11866 , \11675 );
nor \U$5409 ( \11867 , \11662 , \11704 , \11664 , \11706 , \11668 , \11672 , \11675 , \11842 , \11843 , \11844 , \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 , \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 , \11865 , \11866 );
and \U$5410 ( \11868 , RIe5341b8_6880, \11867 );
buf \U$5411 ( \11869 , \11675 );
buf \U$5412 ( \11870 , \11675 );
buf \U$5413 ( \11871 , \11675 );
buf \U$5414 ( \11872 , \11675 );
buf \U$5415 ( \11873 , \11675 );
buf \U$5416 ( \11874 , \11675 );
buf \U$5417 ( \11875 , \11675 );
buf \U$5418 ( \11876 , \11675 );
buf \U$5419 ( \11877 , \11675 );
buf \U$5420 ( \11878 , \11675 );
buf \U$5421 ( \11879 , \11675 );
buf \U$5422 ( \11880 , \11675 );
buf \U$5423 ( \11881 , \11675 );
buf \U$5424 ( \11882 , \11675 );
buf \U$5425 ( \11883 , \11675 );
buf \U$5426 ( \11884 , \11675 );
buf \U$5427 ( \11885 , \11675 );
buf \U$5428 ( \11886 , \11675 );
buf \U$5429 ( \11887 , \11675 );
buf \U$5430 ( \11888 , \11675 );
buf \U$5431 ( \11889 , \11675 );
buf \U$5432 ( \11890 , \11675 );
buf \U$5433 ( \11891 , \11675 );
buf \U$5434 ( \11892 , \11675 );
buf \U$5435 ( \11893 , \11675 );
nor \U$5436 ( \11894 , \11703 , \11663 , \11664 , \11706 , \11668 , \11672 , \11675 , \11869 , \11870 , \11871 , \11872 , \11873 , \11874 , \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 , \11882 , \11883 , \11884 , \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 , \11892 , \11893 );
and \U$5437 ( \11895 , RIe5349b0_6879, \11894 );
buf \U$5438 ( \11896 , \11675 );
buf \U$5439 ( \11897 , \11675 );
buf \U$5440 ( \11898 , \11675 );
buf \U$5441 ( \11899 , \11675 );
buf \U$5442 ( \11900 , \11675 );
buf \U$5443 ( \11901 , \11675 );
buf \U$5444 ( \11902 , \11675 );
buf \U$5445 ( \11903 , \11675 );
buf \U$5446 ( \11904 , \11675 );
buf \U$5447 ( \11905 , \11675 );
buf \U$5448 ( \11906 , \11675 );
buf \U$5449 ( \11907 , \11675 );
buf \U$5450 ( \11908 , \11675 );
buf \U$5451 ( \11909 , \11675 );
buf \U$5452 ( \11910 , \11675 );
buf \U$5453 ( \11911 , \11675 );
buf \U$5454 ( \11912 , \11675 );
buf \U$5455 ( \11913 , \11675 );
buf \U$5456 ( \11914 , \11675 );
buf \U$5457 ( \11915 , \11675 );
buf \U$5458 ( \11916 , \11675 );
buf \U$5459 ( \11917 , \11675 );
buf \U$5460 ( \11918 , \11675 );
buf \U$5461 ( \11919 , \11675 );
buf \U$5462 ( \11920 , \11675 );
nor \U$5463 ( \11921 , \11662 , \11663 , \11664 , \11706 , \11668 , \11672 , \11675 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 , \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 , \11915 , \11916 , \11917 , \11918 , \11919 , \11920 );
and \U$5464 ( \11922 , RIea94af8_6890, \11921 );
buf \U$5465 ( \11923 , \11675 );
buf \U$5466 ( \11924 , \11675 );
buf \U$5467 ( \11925 , \11675 );
buf \U$5468 ( \11926 , \11675 );
buf \U$5469 ( \11927 , \11675 );
buf \U$5470 ( \11928 , \11675 );
buf \U$5471 ( \11929 , \11675 );
buf \U$5472 ( \11930 , \11675 );
buf \U$5473 ( \11931 , \11675 );
buf \U$5474 ( \11932 , \11675 );
buf \U$5475 ( \11933 , \11675 );
buf \U$5476 ( \11934 , \11675 );
buf \U$5477 ( \11935 , \11675 );
buf \U$5478 ( \11936 , \11675 );
buf \U$5479 ( \11937 , \11675 );
buf \U$5480 ( \11938 , \11675 );
buf \U$5481 ( \11939 , \11675 );
buf \U$5482 ( \11940 , \11675 );
buf \U$5483 ( \11941 , \11675 );
buf \U$5484 ( \11942 , \11675 );
buf \U$5485 ( \11943 , \11675 );
buf \U$5486 ( \11944 , \11675 );
buf \U$5487 ( \11945 , \11675 );
buf \U$5488 ( \11946 , \11675 );
buf \U$5489 ( \11947 , \11675 );
nor \U$5490 ( \11948 , \11703 , \11704 , \11705 , \11665 , \11668 , \11672 , \11675 , \11923 , \11924 , \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 , \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 , \11945 , \11946 , \11947 );
and \U$5491 ( \11949 , RIe5351a8_6878, \11948 );
buf \U$5492 ( \11950 , \11675 );
buf \U$5493 ( \11951 , \11675 );
buf \U$5494 ( \11952 , \11675 );
buf \U$5495 ( \11953 , \11675 );
buf \U$5496 ( \11954 , \11675 );
buf \U$5497 ( \11955 , \11675 );
buf \U$5498 ( \11956 , \11675 );
buf \U$5499 ( \11957 , \11675 );
buf \U$5500 ( \11958 , \11675 );
buf \U$5501 ( \11959 , \11675 );
buf \U$5502 ( \11960 , \11675 );
buf \U$5503 ( \11961 , \11675 );
buf \U$5504 ( \11962 , \11675 );
buf \U$5505 ( \11963 , \11675 );
buf \U$5506 ( \11964 , \11675 );
buf \U$5507 ( \11965 , \11675 );
buf \U$5508 ( \11966 , \11675 );
buf \U$5509 ( \11967 , \11675 );
buf \U$5510 ( \11968 , \11675 );
buf \U$5511 ( \11969 , \11675 );
buf \U$5512 ( \11970 , \11675 );
buf \U$5513 ( \11971 , \11675 );
buf \U$5514 ( \11972 , \11675 );
buf \U$5515 ( \11973 , \11675 );
buf \U$5516 ( \11974 , \11675 );
nor \U$5517 ( \11975 , \11662 , \11704 , \11705 , \11665 , \11668 , \11672 , \11675 , \11950 , \11951 , \11952 , \11953 , \11954 , \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 , \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 , \11972 , \11973 , \11974 );
and \U$5518 ( \11976 , RIe5359a0_6877, \11975 );
buf \U$5519 ( \11977 , \11675 );
buf \U$5520 ( \11978 , \11675 );
buf \U$5521 ( \11979 , \11675 );
buf \U$5522 ( \11980 , \11675 );
buf \U$5523 ( \11981 , \11675 );
buf \U$5524 ( \11982 , \11675 );
buf \U$5525 ( \11983 , \11675 );
buf \U$5526 ( \11984 , \11675 );
buf \U$5527 ( \11985 , \11675 );
buf \U$5528 ( \11986 , \11675 );
buf \U$5529 ( \11987 , \11675 );
buf \U$5530 ( \11988 , \11675 );
buf \U$5531 ( \11989 , \11675 );
buf \U$5532 ( \11990 , \11675 );
buf \U$5533 ( \11991 , \11675 );
buf \U$5534 ( \11992 , \11675 );
buf \U$5535 ( \11993 , \11675 );
buf \U$5536 ( \11994 , \11675 );
buf \U$5537 ( \11995 , \11675 );
buf \U$5538 ( \11996 , \11675 );
buf \U$5539 ( \11997 , \11675 );
buf \U$5540 ( \11998 , \11675 );
buf \U$5541 ( \11999 , \11675 );
buf \U$5542 ( \12000 , \11675 );
buf \U$5543 ( \12001 , \11675 );
nor \U$5544 ( \12002 , \11703 , \11663 , \11705 , \11665 , \11668 , \11672 , \11675 , \11977 , \11978 , \11979 , \11980 , \11981 , \11982 , \11983 , \11984 , \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 , \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 );
and \U$5545 ( \12003 , RIeab78c8_6895, \12002 );
buf \U$5546 ( \12004 , \11675 );
buf \U$5547 ( \12005 , \11675 );
buf \U$5548 ( \12006 , \11675 );
buf \U$5549 ( \12007 , \11675 );
buf \U$5550 ( \12008 , \11675 );
buf \U$5551 ( \12009 , \11675 );
buf \U$5552 ( \12010 , \11675 );
buf \U$5553 ( \12011 , \11675 );
buf \U$5554 ( \12012 , \11675 );
buf \U$5555 ( \12013 , \11675 );
buf \U$5556 ( \12014 , \11675 );
buf \U$5557 ( \12015 , \11675 );
buf \U$5558 ( \12016 , \11675 );
buf \U$5559 ( \12017 , \11675 );
buf \U$5560 ( \12018 , \11675 );
buf \U$5561 ( \12019 , \11675 );
buf \U$5562 ( \12020 , \11675 );
buf \U$5563 ( \12021 , \11675 );
buf \U$5564 ( \12022 , \11675 );
buf \U$5565 ( \12023 , \11675 );
buf \U$5566 ( \12024 , \11675 );
buf \U$5567 ( \12025 , \11675 );
buf \U$5568 ( \12026 , \11675 );
buf \U$5569 ( \12027 , \11675 );
buf \U$5570 ( \12028 , \11675 );
nor \U$5571 ( \12029 , \11662 , \11663 , \11705 , \11665 , \11668 , \11672 , \11675 , \12004 , \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 , \12012 , \12013 , \12014 , \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 , \12025 , \12026 , \12027 , \12028 );
and \U$5572 ( \12030 , RIeab7d00_6896, \12029 );
buf \U$5573 ( \12031 , \11675 );
buf \U$5574 ( \12032 , \11675 );
buf \U$5575 ( \12033 , \11675 );
buf \U$5576 ( \12034 , \11675 );
buf \U$5577 ( \12035 , \11675 );
buf \U$5578 ( \12036 , \11675 );
buf \U$5579 ( \12037 , \11675 );
buf \U$5580 ( \12038 , \11675 );
buf \U$5581 ( \12039 , \11675 );
buf \U$5582 ( \12040 , \11675 );
buf \U$5583 ( \12041 , \11675 );
buf \U$5584 ( \12042 , \11675 );
buf \U$5585 ( \12043 , \11675 );
buf \U$5586 ( \12044 , \11675 );
buf \U$5587 ( \12045 , \11675 );
buf \U$5588 ( \12046 , \11675 );
buf \U$5589 ( \12047 , \11675 );
buf \U$5590 ( \12048 , \11675 );
buf \U$5591 ( \12049 , \11675 );
buf \U$5592 ( \12050 , \11675 );
buf \U$5593 ( \12051 , \11675 );
buf \U$5594 ( \12052 , \11675 );
buf \U$5595 ( \12053 , \11675 );
buf \U$5596 ( \12054 , \11675 );
buf \U$5597 ( \12055 , \11675 );
nor \U$5598 ( \12056 , \11703 , \11704 , \11664 , \11665 , \11668 , \11672 , \11675 , \12031 , \12032 , \12033 , \12034 , \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 , \12042 , \12043 , \12044 , \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 , \12055 );
and \U$5599 ( \12057 , RIeacfa18_6902, \12056 );
buf \U$5600 ( \12058 , \11675 );
buf \U$5601 ( \12059 , \11675 );
buf \U$5602 ( \12060 , \11675 );
buf \U$5603 ( \12061 , \11675 );
buf \U$5604 ( \12062 , \11675 );
buf \U$5605 ( \12063 , \11675 );
buf \U$5606 ( \12064 , \11675 );
buf \U$5607 ( \12065 , \11675 );
buf \U$5608 ( \12066 , \11675 );
buf \U$5609 ( \12067 , \11675 );
buf \U$5610 ( \12068 , \11675 );
buf \U$5611 ( \12069 , \11675 );
buf \U$5612 ( \12070 , \11675 );
buf \U$5613 ( \12071 , \11675 );
buf \U$5614 ( \12072 , \11675 );
buf \U$5615 ( \12073 , \11675 );
buf \U$5616 ( \12074 , \11675 );
buf \U$5617 ( \12075 , \11675 );
buf \U$5618 ( \12076 , \11675 );
buf \U$5619 ( \12077 , \11675 );
buf \U$5620 ( \12078 , \11675 );
buf \U$5621 ( \12079 , \11675 );
buf \U$5622 ( \12080 , \11675 );
buf \U$5623 ( \12081 , \11675 );
buf \U$5624 ( \12082 , \11675 );
nor \U$5625 ( \12083 , \11662 , \11704 , \11664 , \11665 , \11668 , \11672 , \11675 , \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 , \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 , \12072 , \12073 , \12074 , \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 , \12082 );
and \U$5626 ( \12084 , RIeab6518_6891, \12083 );
buf \U$5627 ( \12085 , \11675 );
buf \U$5628 ( \12086 , \11675 );
buf \U$5629 ( \12087 , \11675 );
buf \U$5630 ( \12088 , \11675 );
buf \U$5631 ( \12089 , \11675 );
buf \U$5632 ( \12090 , \11675 );
buf \U$5633 ( \12091 , \11675 );
buf \U$5634 ( \12092 , \11675 );
buf \U$5635 ( \12093 , \11675 );
buf \U$5636 ( \12094 , \11675 );
buf \U$5637 ( \12095 , \11675 );
buf \U$5638 ( \12096 , \11675 );
buf \U$5639 ( \12097 , \11675 );
buf \U$5640 ( \12098 , \11675 );
buf \U$5641 ( \12099 , \11675 );
buf \U$5642 ( \12100 , \11675 );
buf \U$5643 ( \12101 , \11675 );
buf \U$5644 ( \12102 , \11675 );
buf \U$5645 ( \12103 , \11675 );
buf \U$5646 ( \12104 , \11675 );
buf \U$5647 ( \12105 , \11675 );
buf \U$5648 ( \12106 , \11675 );
buf \U$5649 ( \12107 , \11675 );
buf \U$5650 ( \12108 , \11675 );
buf \U$5651 ( \12109 , \11675 );
nor \U$5652 ( \12110 , \11703 , \11663 , \11664 , \11665 , \11668 , \11672 , \11675 , \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 , \12092 , \12093 , \12094 , \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 , \12102 , \12103 , \12104 , \12105 , \12106 , \12107 , \12108 , \12109 );
and \U$5653 ( \12111 , RIeb352c8_6904, \12110 );
or \U$5654 ( \12112 , \11702 , \11733 , \11760 , \11787 , \11814 , \11841 , \11868 , \11895 , \11922 , \11949 , \11976 , \12003 , \12030 , \12057 , \12084 , \12111 );
buf \U$5655 ( \12113 , \11675 );
not \U$5656 ( \12114 , \12113 );
buf \U$5657 ( \12115 , \11663 );
buf \U$5658 ( \12116 , \11664 );
buf \U$5659 ( \12117 , \11665 );
buf \U$5660 ( \12118 , \11668 );
buf \U$5661 ( \12119 , \11672 );
buf \U$5662 ( \12120 , \11675 );
buf \U$5663 ( \12121 , \11675 );
buf \U$5664 ( \12122 , \11675 );
buf \U$5665 ( \12123 , \11675 );
buf \U$5666 ( \12124 , \11675 );
buf \U$5667 ( \12125 , \11675 );
buf \U$5668 ( \12126 , \11675 );
buf \U$5669 ( \12127 , \11675 );
buf \U$5670 ( \12128 , \11675 );
buf \U$5671 ( \12129 , \11675 );
buf \U$5672 ( \12130 , \11675 );
buf \U$5673 ( \12131 , \11675 );
buf \U$5674 ( \12132 , \11675 );
buf \U$5675 ( \12133 , \11675 );
buf \U$5676 ( \12134 , \11675 );
buf \U$5677 ( \12135 , \11675 );
buf \U$5678 ( \12136 , \11675 );
buf \U$5679 ( \12137 , \11675 );
buf \U$5680 ( \12138 , \11675 );
buf \U$5681 ( \12139 , \11675 );
buf \U$5682 ( \12140 , \11675 );
buf \U$5683 ( \12141 , \11675 );
buf \U$5684 ( \12142 , \11675 );
buf \U$5685 ( \12143 , \11675 );
buf \U$5686 ( \12144 , \11675 );
buf \U$5687 ( \12145 , \11662 );
or \U$5688 ( \12146 , \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 , \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 , \12132 , \12133 , \12134 , \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 , \12142 , \12143 , \12144 , \12145 );
nand \U$5689 ( \12147 , \12114 , \12146 );
buf \U$5690 ( \12148 , \12147 );
buf \U$5691 ( \12149 , \11675 );
not \U$5692 ( \12150 , \12149 );
buf \U$5693 ( \12151 , \11672 );
buf \U$5694 ( \12152 , \11675 );
buf \U$5695 ( \12153 , \11675 );
buf \U$5696 ( \12154 , \11675 );
buf \U$5697 ( \12155 , \11675 );
buf \U$5698 ( \12156 , \11675 );
buf \U$5699 ( \12157 , \11675 );
buf \U$5700 ( \12158 , \11675 );
buf \U$5701 ( \12159 , \11675 );
buf \U$5702 ( \12160 , \11675 );
buf \U$5703 ( \12161 , \11675 );
buf \U$5704 ( \12162 , \11675 );
buf \U$5705 ( \12163 , \11675 );
buf \U$5706 ( \12164 , \11675 );
buf \U$5707 ( \12165 , \11675 );
buf \U$5708 ( \12166 , \11675 );
buf \U$5709 ( \12167 , \11675 );
buf \U$5710 ( \12168 , \11675 );
buf \U$5711 ( \12169 , \11675 );
buf \U$5712 ( \12170 , \11675 );
buf \U$5713 ( \12171 , \11675 );
buf \U$5714 ( \12172 , \11675 );
buf \U$5715 ( \12173 , \11675 );
buf \U$5716 ( \12174 , \11675 );
buf \U$5717 ( \12175 , \11675 );
buf \U$5718 ( \12176 , \11675 );
buf \U$5719 ( \12177 , \11668 );
buf \U$5720 ( \12178 , \11662 );
buf \U$5721 ( \12179 , \11663 );
buf \U$5722 ( \12180 , \11664 );
buf \U$5723 ( \12181 , \11665 );
or \U$5724 ( \12182 , \12178 , \12179 , \12180 , \12181 );
and \U$5725 ( \12183 , \12177 , \12182 );
or \U$5726 ( \12184 , \12151 , \12152 , \12153 , \12154 , \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 , \12162 , \12163 , \12164 , \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 , \12172 , \12173 , \12174 , \12175 , \12176 , \12183 );
and \U$5727 ( \12185 , \12150 , \12184 );
buf \U$5728 ( \12186 , \12185 );
or \U$5729 ( \12187 , \12148 , \12186 );
_DC g465e ( \12188_nG465e , \12112 , \12187 );
not \U$5730 ( \12189 , \12188_nG465e );
buf \U$5731 ( \12190 , RIb7b9608_246);
buf \U$5732 ( \12191 , \11675 );
buf \U$5733 ( \12192 , \11675 );
buf \U$5734 ( \12193 , \11675 );
buf \U$5735 ( \12194 , \11675 );
buf \U$5736 ( \12195 , \11675 );
buf \U$5737 ( \12196 , \11675 );
buf \U$5738 ( \12197 , \11675 );
buf \U$5739 ( \12198 , \11675 );
buf \U$5740 ( \12199 , \11675 );
buf \U$5741 ( \12200 , \11675 );
buf \U$5742 ( \12201 , \11675 );
buf \U$5743 ( \12202 , \11675 );
buf \U$5744 ( \12203 , \11675 );
buf \U$5745 ( \12204 , \11675 );
buf \U$5746 ( \12205 , \11675 );
buf \U$5747 ( \12206 , \11675 );
buf \U$5748 ( \12207 , \11675 );
buf \U$5749 ( \12208 , \11675 );
buf \U$5750 ( \12209 , \11675 );
buf \U$5751 ( \12210 , \11675 );
buf \U$5752 ( \12211 , \11675 );
buf \U$5753 ( \12212 , \11675 );
buf \U$5754 ( \12213 , \11675 );
buf \U$5755 ( \12214 , \11675 );
buf \U$5756 ( \12215 , \11675 );
nor \U$5757 ( \12216 , \11662 , \11663 , \11664 , \11665 , \11669 , \11672 , \11675 , \12191 , \12192 , \12193 , \12194 , \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 , \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 , \12212 , \12213 , \12214 , \12215 );
and \U$5758 ( \12217 , \7117 , \12216 );
buf \U$5759 ( \12218 , \11675 );
buf \U$5760 ( \12219 , \11675 );
buf \U$5761 ( \12220 , \11675 );
buf \U$5762 ( \12221 , \11675 );
buf \U$5763 ( \12222 , \11675 );
buf \U$5764 ( \12223 , \11675 );
buf \U$5765 ( \12224 , \11675 );
buf \U$5766 ( \12225 , \11675 );
buf \U$5767 ( \12226 , \11675 );
buf \U$5768 ( \12227 , \11675 );
buf \U$5769 ( \12228 , \11675 );
buf \U$5770 ( \12229 , \11675 );
buf \U$5771 ( \12230 , \11675 );
buf \U$5772 ( \12231 , \11675 );
buf \U$5773 ( \12232 , \11675 );
buf \U$5774 ( \12233 , \11675 );
buf \U$5775 ( \12234 , \11675 );
buf \U$5776 ( \12235 , \11675 );
buf \U$5777 ( \12236 , \11675 );
buf \U$5778 ( \12237 , \11675 );
buf \U$5779 ( \12238 , \11675 );
buf \U$5780 ( \12239 , \11675 );
buf \U$5781 ( \12240 , \11675 );
buf \U$5782 ( \12241 , \11675 );
buf \U$5783 ( \12242 , \11675 );
nor \U$5784 ( \12243 , \11703 , \11704 , \11705 , \11706 , \11668 , \11672 , \11675 , \12218 , \12219 , \12220 , \12221 , \12222 , \12223 , \12224 , \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 , \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 , \12242 );
and \U$5785 ( \12244 , \7119 , \12243 );
buf \U$5786 ( \12245 , \11675 );
buf \U$5787 ( \12246 , \11675 );
buf \U$5788 ( \12247 , \11675 );
buf \U$5789 ( \12248 , \11675 );
buf \U$5790 ( \12249 , \11675 );
buf \U$5791 ( \12250 , \11675 );
buf \U$5792 ( \12251 , \11675 );
buf \U$5793 ( \12252 , \11675 );
buf \U$5794 ( \12253 , \11675 );
buf \U$5795 ( \12254 , \11675 );
buf \U$5796 ( \12255 , \11675 );
buf \U$5797 ( \12256 , \11675 );
buf \U$5798 ( \12257 , \11675 );
buf \U$5799 ( \12258 , \11675 );
buf \U$5800 ( \12259 , \11675 );
buf \U$5801 ( \12260 , \11675 );
buf \U$5802 ( \12261 , \11675 );
buf \U$5803 ( \12262 , \11675 );
buf \U$5804 ( \12263 , \11675 );
buf \U$5805 ( \12264 , \11675 );
buf \U$5806 ( \12265 , \11675 );
buf \U$5807 ( \12266 , \11675 );
buf \U$5808 ( \12267 , \11675 );
buf \U$5809 ( \12268 , \11675 );
buf \U$5810 ( \12269 , \11675 );
nor \U$5811 ( \12270 , \11662 , \11704 , \11705 , \11706 , \11668 , \11672 , \11675 , \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 , \12252 , \12253 , \12254 , \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 , \12265 , \12266 , \12267 , \12268 , \12269 );
and \U$5812 ( \12271 , \7864 , \12270 );
buf \U$5813 ( \12272 , \11675 );
buf \U$5814 ( \12273 , \11675 );
buf \U$5815 ( \12274 , \11675 );
buf \U$5816 ( \12275 , \11675 );
buf \U$5817 ( \12276 , \11675 );
buf \U$5818 ( \12277 , \11675 );
buf \U$5819 ( \12278 , \11675 );
buf \U$5820 ( \12279 , \11675 );
buf \U$5821 ( \12280 , \11675 );
buf \U$5822 ( \12281 , \11675 );
buf \U$5823 ( \12282 , \11675 );
buf \U$5824 ( \12283 , \11675 );
buf \U$5825 ( \12284 , \11675 );
buf \U$5826 ( \12285 , \11675 );
buf \U$5827 ( \12286 , \11675 );
buf \U$5828 ( \12287 , \11675 );
buf \U$5829 ( \12288 , \11675 );
buf \U$5830 ( \12289 , \11675 );
buf \U$5831 ( \12290 , \11675 );
buf \U$5832 ( \12291 , \11675 );
buf \U$5833 ( \12292 , \11675 );
buf \U$5834 ( \12293 , \11675 );
buf \U$5835 ( \12294 , \11675 );
buf \U$5836 ( \12295 , \11675 );
buf \U$5837 ( \12296 , \11675 );
nor \U$5838 ( \12297 , \11703 , \11663 , \11705 , \11706 , \11668 , \11672 , \11675 , \12272 , \12273 , \12274 , \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 , \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 , \12295 , \12296 );
and \U$5839 ( \12298 , \7892 , \12297 );
buf \U$5840 ( \12299 , \11675 );
buf \U$5841 ( \12300 , \11675 );
buf \U$5842 ( \12301 , \11675 );
buf \U$5843 ( \12302 , \11675 );
buf \U$5844 ( \12303 , \11675 );
buf \U$5845 ( \12304 , \11675 );
buf \U$5846 ( \12305 , \11675 );
buf \U$5847 ( \12306 , \11675 );
buf \U$5848 ( \12307 , \11675 );
buf \U$5849 ( \12308 , \11675 );
buf \U$5850 ( \12309 , \11675 );
buf \U$5851 ( \12310 , \11675 );
buf \U$5852 ( \12311 , \11675 );
buf \U$5853 ( \12312 , \11675 );
buf \U$5854 ( \12313 , \11675 );
buf \U$5855 ( \12314 , \11675 );
buf \U$5856 ( \12315 , \11675 );
buf \U$5857 ( \12316 , \11675 );
buf \U$5858 ( \12317 , \11675 );
buf \U$5859 ( \12318 , \11675 );
buf \U$5860 ( \12319 , \11675 );
buf \U$5861 ( \12320 , \11675 );
buf \U$5862 ( \12321 , \11675 );
buf \U$5863 ( \12322 , \11675 );
buf \U$5864 ( \12323 , \11675 );
nor \U$5865 ( \12324 , \11662 , \11663 , \11705 , \11706 , \11668 , \11672 , \11675 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 , \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 , \12312 , \12313 , \12314 , \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 , \12322 , \12323 );
and \U$5866 ( \12325 , \7920 , \12324 );
buf \U$5867 ( \12326 , \11675 );
buf \U$5868 ( \12327 , \11675 );
buf \U$5869 ( \12328 , \11675 );
buf \U$5870 ( \12329 , \11675 );
buf \U$5871 ( \12330 , \11675 );
buf \U$5872 ( \12331 , \11675 );
buf \U$5873 ( \12332 , \11675 );
buf \U$5874 ( \12333 , \11675 );
buf \U$5875 ( \12334 , \11675 );
buf \U$5876 ( \12335 , \11675 );
buf \U$5877 ( \12336 , \11675 );
buf \U$5878 ( \12337 , \11675 );
buf \U$5879 ( \12338 , \11675 );
buf \U$5880 ( \12339 , \11675 );
buf \U$5881 ( \12340 , \11675 );
buf \U$5882 ( \12341 , \11675 );
buf \U$5883 ( \12342 , \11675 );
buf \U$5884 ( \12343 , \11675 );
buf \U$5885 ( \12344 , \11675 );
buf \U$5886 ( \12345 , \11675 );
buf \U$5887 ( \12346 , \11675 );
buf \U$5888 ( \12347 , \11675 );
buf \U$5889 ( \12348 , \11675 );
buf \U$5890 ( \12349 , \11675 );
buf \U$5891 ( \12350 , \11675 );
nor \U$5892 ( \12351 , \11703 , \11704 , \11664 , \11706 , \11668 , \11672 , \11675 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 , \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 , \12345 , \12346 , \12347 , \12348 , \12349 , \12350 );
and \U$5893 ( \12352 , \7948 , \12351 );
buf \U$5894 ( \12353 , \11675 );
buf \U$5895 ( \12354 , \11675 );
buf \U$5896 ( \12355 , \11675 );
buf \U$5897 ( \12356 , \11675 );
buf \U$5898 ( \12357 , \11675 );
buf \U$5899 ( \12358 , \11675 );
buf \U$5900 ( \12359 , \11675 );
buf \U$5901 ( \12360 , \11675 );
buf \U$5902 ( \12361 , \11675 );
buf \U$5903 ( \12362 , \11675 );
buf \U$5904 ( \12363 , \11675 );
buf \U$5905 ( \12364 , \11675 );
buf \U$5906 ( \12365 , \11675 );
buf \U$5907 ( \12366 , \11675 );
buf \U$5908 ( \12367 , \11675 );
buf \U$5909 ( \12368 , \11675 );
buf \U$5910 ( \12369 , \11675 );
buf \U$5911 ( \12370 , \11675 );
buf \U$5912 ( \12371 , \11675 );
buf \U$5913 ( \12372 , \11675 );
buf \U$5914 ( \12373 , \11675 );
buf \U$5915 ( \12374 , \11675 );
buf \U$5916 ( \12375 , \11675 );
buf \U$5917 ( \12376 , \11675 );
buf \U$5918 ( \12377 , \11675 );
nor \U$5919 ( \12378 , \11662 , \11704 , \11664 , \11706 , \11668 , \11672 , \11675 , \12353 , \12354 , \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 , \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 , \12372 , \12373 , \12374 , \12375 , \12376 , \12377 );
and \U$5920 ( \12379 , \7976 , \12378 );
buf \U$5921 ( \12380 , \11675 );
buf \U$5922 ( \12381 , \11675 );
buf \U$5923 ( \12382 , \11675 );
buf \U$5924 ( \12383 , \11675 );
buf \U$5925 ( \12384 , \11675 );
buf \U$5926 ( \12385 , \11675 );
buf \U$5927 ( \12386 , \11675 );
buf \U$5928 ( \12387 , \11675 );
buf \U$5929 ( \12388 , \11675 );
buf \U$5930 ( \12389 , \11675 );
buf \U$5931 ( \12390 , \11675 );
buf \U$5932 ( \12391 , \11675 );
buf \U$5933 ( \12392 , \11675 );
buf \U$5934 ( \12393 , \11675 );
buf \U$5935 ( \12394 , \11675 );
buf \U$5936 ( \12395 , \11675 );
buf \U$5937 ( \12396 , \11675 );
buf \U$5938 ( \12397 , \11675 );
buf \U$5939 ( \12398 , \11675 );
buf \U$5940 ( \12399 , \11675 );
buf \U$5941 ( \12400 , \11675 );
buf \U$5942 ( \12401 , \11675 );
buf \U$5943 ( \12402 , \11675 );
buf \U$5944 ( \12403 , \11675 );
buf \U$5945 ( \12404 , \11675 );
nor \U$5946 ( \12405 , \11703 , \11663 , \11664 , \11706 , \11668 , \11672 , \11675 , \12380 , \12381 , \12382 , \12383 , \12384 , \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 );
and \U$5947 ( \12406 , \8004 , \12405 );
buf \U$5948 ( \12407 , \11675 );
buf \U$5949 ( \12408 , \11675 );
buf \U$5950 ( \12409 , \11675 );
buf \U$5951 ( \12410 , \11675 );
buf \U$5952 ( \12411 , \11675 );
buf \U$5953 ( \12412 , \11675 );
buf \U$5954 ( \12413 , \11675 );
buf \U$5955 ( \12414 , \11675 );
buf \U$5956 ( \12415 , \11675 );
buf \U$5957 ( \12416 , \11675 );
buf \U$5958 ( \12417 , \11675 );
buf \U$5959 ( \12418 , \11675 );
buf \U$5960 ( \12419 , \11675 );
buf \U$5961 ( \12420 , \11675 );
buf \U$5962 ( \12421 , \11675 );
buf \U$5963 ( \12422 , \11675 );
buf \U$5964 ( \12423 , \11675 );
buf \U$5965 ( \12424 , \11675 );
buf \U$5966 ( \12425 , \11675 );
buf \U$5967 ( \12426 , \11675 );
buf \U$5968 ( \12427 , \11675 );
buf \U$5969 ( \12428 , \11675 );
buf \U$5970 ( \12429 , \11675 );
buf \U$5971 ( \12430 , \11675 );
buf \U$5972 ( \12431 , \11675 );
nor \U$5973 ( \12432 , \11662 , \11663 , \11664 , \11706 , \11668 , \11672 , \11675 , \12407 , \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 , \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 , \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 );
and \U$5974 ( \12433 , \8032 , \12432 );
buf \U$5975 ( \12434 , \11675 );
buf \U$5976 ( \12435 , \11675 );
buf \U$5977 ( \12436 , \11675 );
buf \U$5978 ( \12437 , \11675 );
buf \U$5979 ( \12438 , \11675 );
buf \U$5980 ( \12439 , \11675 );
buf \U$5981 ( \12440 , \11675 );
buf \U$5982 ( \12441 , \11675 );
buf \U$5983 ( \12442 , \11675 );
buf \U$5984 ( \12443 , \11675 );
buf \U$5985 ( \12444 , \11675 );
buf \U$5986 ( \12445 , \11675 );
buf \U$5987 ( \12446 , \11675 );
buf \U$5988 ( \12447 , \11675 );
buf \U$5989 ( \12448 , \11675 );
buf \U$5990 ( \12449 , \11675 );
buf \U$5991 ( \12450 , \11675 );
buf \U$5992 ( \12451 , \11675 );
buf \U$5993 ( \12452 , \11675 );
buf \U$5994 ( \12453 , \11675 );
buf \U$5995 ( \12454 , \11675 );
buf \U$5996 ( \12455 , \11675 );
buf \U$5997 ( \12456 , \11675 );
buf \U$5998 ( \12457 , \11675 );
buf \U$5999 ( \12458 , \11675 );
nor \U$6000 ( \12459 , \11703 , \11704 , \11705 , \11665 , \11668 , \11672 , \11675 , \12434 , \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 , \12442 , \12443 , \12444 , \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 , \12452 , \12453 , \12454 , \12455 , \12456 , \12457 , \12458 );
and \U$6001 ( \12460 , \8060 , \12459 );
buf \U$6002 ( \12461 , \11675 );
buf \U$6003 ( \12462 , \11675 );
buf \U$6004 ( \12463 , \11675 );
buf \U$6005 ( \12464 , \11675 );
buf \U$6006 ( \12465 , \11675 );
buf \U$6007 ( \12466 , \11675 );
buf \U$6008 ( \12467 , \11675 );
buf \U$6009 ( \12468 , \11675 );
buf \U$6010 ( \12469 , \11675 );
buf \U$6011 ( \12470 , \11675 );
buf \U$6012 ( \12471 , \11675 );
buf \U$6013 ( \12472 , \11675 );
buf \U$6014 ( \12473 , \11675 );
buf \U$6015 ( \12474 , \11675 );
buf \U$6016 ( \12475 , \11675 );
buf \U$6017 ( \12476 , \11675 );
buf \U$6018 ( \12477 , \11675 );
buf \U$6019 ( \12478 , \11675 );
buf \U$6020 ( \12479 , \11675 );
buf \U$6021 ( \12480 , \11675 );
buf \U$6022 ( \12481 , \11675 );
buf \U$6023 ( \12482 , \11675 );
buf \U$6024 ( \12483 , \11675 );
buf \U$6025 ( \12484 , \11675 );
buf \U$6026 ( \12485 , \11675 );
nor \U$6027 ( \12486 , \11662 , \11704 , \11705 , \11665 , \11668 , \11672 , \11675 , \12461 , \12462 , \12463 , \12464 , \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 , \12472 , \12473 , \12474 , \12475 , \12476 , \12477 , \12478 , \12479 , \12480 , \12481 , \12482 , \12483 , \12484 , \12485 );
and \U$6028 ( \12487 , \8088 , \12486 );
buf \U$6029 ( \12488 , \11675 );
buf \U$6030 ( \12489 , \11675 );
buf \U$6031 ( \12490 , \11675 );
buf \U$6032 ( \12491 , \11675 );
buf \U$6033 ( \12492 , \11675 );
buf \U$6034 ( \12493 , \11675 );
buf \U$6035 ( \12494 , \11675 );
buf \U$6036 ( \12495 , \11675 );
buf \U$6037 ( \12496 , \11675 );
buf \U$6038 ( \12497 , \11675 );
buf \U$6039 ( \12498 , \11675 );
buf \U$6040 ( \12499 , \11675 );
buf \U$6041 ( \12500 , \11675 );
buf \U$6042 ( \12501 , \11675 );
buf \U$6043 ( \12502 , \11675 );
buf \U$6044 ( \12503 , \11675 );
buf \U$6045 ( \12504 , \11675 );
buf \U$6046 ( \12505 , \11675 );
buf \U$6047 ( \12506 , \11675 );
buf \U$6048 ( \12507 , \11675 );
buf \U$6049 ( \12508 , \11675 );
buf \U$6050 ( \12509 , \11675 );
buf \U$6051 ( \12510 , \11675 );
buf \U$6052 ( \12511 , \11675 );
buf \U$6053 ( \12512 , \11675 );
nor \U$6054 ( \12513 , \11703 , \11663 , \11705 , \11665 , \11668 , \11672 , \11675 , \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 , \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12504 , \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 , \12512 );
and \U$6055 ( \12514 , \8116 , \12513 );
buf \U$6056 ( \12515 , \11675 );
buf \U$6057 ( \12516 , \11675 );
buf \U$6058 ( \12517 , \11675 );
buf \U$6059 ( \12518 , \11675 );
buf \U$6060 ( \12519 , \11675 );
buf \U$6061 ( \12520 , \11675 );
buf \U$6062 ( \12521 , \11675 );
buf \U$6063 ( \12522 , \11675 );
buf \U$6064 ( \12523 , \11675 );
buf \U$6065 ( \12524 , \11675 );
buf \U$6066 ( \12525 , \11675 );
buf \U$6067 ( \12526 , \11675 );
buf \U$6068 ( \12527 , \11675 );
buf \U$6069 ( \12528 , \11675 );
buf \U$6070 ( \12529 , \11675 );
buf \U$6071 ( \12530 , \11675 );
buf \U$6072 ( \12531 , \11675 );
buf \U$6073 ( \12532 , \11675 );
buf \U$6074 ( \12533 , \11675 );
buf \U$6075 ( \12534 , \11675 );
buf \U$6076 ( \12535 , \11675 );
buf \U$6077 ( \12536 , \11675 );
buf \U$6078 ( \12537 , \11675 );
buf \U$6079 ( \12538 , \11675 );
buf \U$6080 ( \12539 , \11675 );
nor \U$6081 ( \12540 , \11662 , \11663 , \11705 , \11665 , \11668 , \11672 , \11675 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 , \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 , \12535 , \12536 , \12537 , \12538 , \12539 );
and \U$6082 ( \12541 , \8144 , \12540 );
buf \U$6083 ( \12542 , \11675 );
buf \U$6084 ( \12543 , \11675 );
buf \U$6085 ( \12544 , \11675 );
buf \U$6086 ( \12545 , \11675 );
buf \U$6087 ( \12546 , \11675 );
buf \U$6088 ( \12547 , \11675 );
buf \U$6089 ( \12548 , \11675 );
buf \U$6090 ( \12549 , \11675 );
buf \U$6091 ( \12550 , \11675 );
buf \U$6092 ( \12551 , \11675 );
buf \U$6093 ( \12552 , \11675 );
buf \U$6094 ( \12553 , \11675 );
buf \U$6095 ( \12554 , \11675 );
buf \U$6096 ( \12555 , \11675 );
buf \U$6097 ( \12556 , \11675 );
buf \U$6098 ( \12557 , \11675 );
buf \U$6099 ( \12558 , \11675 );
buf \U$6100 ( \12559 , \11675 );
buf \U$6101 ( \12560 , \11675 );
buf \U$6102 ( \12561 , \11675 );
buf \U$6103 ( \12562 , \11675 );
buf \U$6104 ( \12563 , \11675 );
buf \U$6105 ( \12564 , \11675 );
buf \U$6106 ( \12565 , \11675 );
buf \U$6107 ( \12566 , \11675 );
nor \U$6108 ( \12567 , \11703 , \11704 , \11664 , \11665 , \11668 , \11672 , \11675 , \12542 , \12543 , \12544 , \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 , \12552 , \12553 , \12554 , \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 , \12565 , \12566 );
and \U$6109 ( \12568 , \8172 , \12567 );
buf \U$6110 ( \12569 , \11675 );
buf \U$6111 ( \12570 , \11675 );
buf \U$6112 ( \12571 , \11675 );
buf \U$6113 ( \12572 , \11675 );
buf \U$6114 ( \12573 , \11675 );
buf \U$6115 ( \12574 , \11675 );
buf \U$6116 ( \12575 , \11675 );
buf \U$6117 ( \12576 , \11675 );
buf \U$6118 ( \12577 , \11675 );
buf \U$6119 ( \12578 , \11675 );
buf \U$6120 ( \12579 , \11675 );
buf \U$6121 ( \12580 , \11675 );
buf \U$6122 ( \12581 , \11675 );
buf \U$6123 ( \12582 , \11675 );
buf \U$6124 ( \12583 , \11675 );
buf \U$6125 ( \12584 , \11675 );
buf \U$6126 ( \12585 , \11675 );
buf \U$6127 ( \12586 , \11675 );
buf \U$6128 ( \12587 , \11675 );
buf \U$6129 ( \12588 , \11675 );
buf \U$6130 ( \12589 , \11675 );
buf \U$6131 ( \12590 , \11675 );
buf \U$6132 ( \12591 , \11675 );
buf \U$6133 ( \12592 , \11675 );
buf \U$6134 ( \12593 , \11675 );
nor \U$6135 ( \12594 , \11662 , \11704 , \11664 , \11665 , \11668 , \11672 , \11675 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 , \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 , \12593 );
and \U$6136 ( \12595 , \8200 , \12594 );
buf \U$6137 ( \12596 , \11675 );
buf \U$6138 ( \12597 , \11675 );
buf \U$6139 ( \12598 , \11675 );
buf \U$6140 ( \12599 , \11675 );
buf \U$6141 ( \12600 , \11675 );
buf \U$6142 ( \12601 , \11675 );
buf \U$6143 ( \12602 , \11675 );
buf \U$6144 ( \12603 , \11675 );
buf \U$6145 ( \12604 , \11675 );
buf \U$6146 ( \12605 , \11675 );
buf \U$6147 ( \12606 , \11675 );
buf \U$6148 ( \12607 , \11675 );
buf \U$6149 ( \12608 , \11675 );
buf \U$6150 ( \12609 , \11675 );
buf \U$6151 ( \12610 , \11675 );
buf \U$6152 ( \12611 , \11675 );
buf \U$6153 ( \12612 , \11675 );
buf \U$6154 ( \12613 , \11675 );
buf \U$6155 ( \12614 , \11675 );
buf \U$6156 ( \12615 , \11675 );
buf \U$6157 ( \12616 , \11675 );
buf \U$6158 ( \12617 , \11675 );
buf \U$6159 ( \12618 , \11675 );
buf \U$6160 ( \12619 , \11675 );
buf \U$6161 ( \12620 , \11675 );
nor \U$6162 ( \12621 , \11703 , \11663 , \11664 , \11665 , \11668 , \11672 , \11675 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 );
and \U$6163 ( \12622 , \8228 , \12621 );
or \U$6164 ( \12623 , \12217 , \12244 , \12271 , \12298 , \12325 , \12352 , \12379 , \12406 , \12433 , \12460 , \12487 , \12514 , \12541 , \12568 , \12595 , \12622 );
buf \U$6165 ( \12624 , \11675 );
not \U$6166 ( \12625 , \12624 );
buf \U$6167 ( \12626 , \11663 );
buf \U$6168 ( \12627 , \11664 );
buf \U$6169 ( \12628 , \11665 );
buf \U$6170 ( \12629 , \11668 );
buf \U$6171 ( \12630 , \11672 );
buf \U$6172 ( \12631 , \11675 );
buf \U$6173 ( \12632 , \11675 );
buf \U$6174 ( \12633 , \11675 );
buf \U$6175 ( \12634 , \11675 );
buf \U$6176 ( \12635 , \11675 );
buf \U$6177 ( \12636 , \11675 );
buf \U$6178 ( \12637 , \11675 );
buf \U$6179 ( \12638 , \11675 );
buf \U$6180 ( \12639 , \11675 );
buf \U$6181 ( \12640 , \11675 );
buf \U$6182 ( \12641 , \11675 );
buf \U$6183 ( \12642 , \11675 );
buf \U$6184 ( \12643 , \11675 );
buf \U$6185 ( \12644 , \11675 );
buf \U$6186 ( \12645 , \11675 );
buf \U$6187 ( \12646 , \11675 );
buf \U$6188 ( \12647 , \11675 );
buf \U$6189 ( \12648 , \11675 );
buf \U$6190 ( \12649 , \11675 );
buf \U$6191 ( \12650 , \11675 );
buf \U$6192 ( \12651 , \11675 );
buf \U$6193 ( \12652 , \11675 );
buf \U$6194 ( \12653 , \11675 );
buf \U$6195 ( \12654 , \11675 );
buf \U$6196 ( \12655 , \11675 );
buf \U$6197 ( \12656 , \11662 );
or \U$6198 ( \12657 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 , \12633 , \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 , \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 , \12655 , \12656 );
nand \U$6199 ( \12658 , \12625 , \12657 );
buf \U$6200 ( \12659 , \12658 );
buf \U$6201 ( \12660 , \11675 );
not \U$6202 ( \12661 , \12660 );
buf \U$6203 ( \12662 , \11672 );
buf \U$6204 ( \12663 , \11675 );
buf \U$6205 ( \12664 , \11675 );
buf \U$6206 ( \12665 , \11675 );
buf \U$6207 ( \12666 , \11675 );
buf \U$6208 ( \12667 , \11675 );
buf \U$6209 ( \12668 , \11675 );
buf \U$6210 ( \12669 , \11675 );
buf \U$6211 ( \12670 , \11675 );
buf \U$6212 ( \12671 , \11675 );
buf \U$6213 ( \12672 , \11675 );
buf \U$6214 ( \12673 , \11675 );
buf \U$6215 ( \12674 , \11675 );
buf \U$6216 ( \12675 , \11675 );
buf \U$6217 ( \12676 , \11675 );
buf \U$6218 ( \12677 , \11675 );
buf \U$6219 ( \12678 , \11675 );
buf \U$6220 ( \12679 , \11675 );
buf \U$6221 ( \12680 , \11675 );
buf \U$6222 ( \12681 , \11675 );
buf \U$6223 ( \12682 , \11675 );
buf \U$6224 ( \12683 , \11675 );
buf \U$6225 ( \12684 , \11675 );
buf \U$6226 ( \12685 , \11675 );
buf \U$6227 ( \12686 , \11675 );
buf \U$6228 ( \12687 , \11675 );
buf \U$6229 ( \12688 , \11668 );
buf \U$6230 ( \12689 , \11662 );
buf \U$6231 ( \12690 , \11663 );
buf \U$6232 ( \12691 , \11664 );
buf \U$6233 ( \12692 , \11665 );
or \U$6234 ( \12693 , \12689 , \12690 , \12691 , \12692 );
and \U$6235 ( \12694 , \12688 , \12693 );
or \U$6236 ( \12695 , \12662 , \12663 , \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 , \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 , \12685 , \12686 , \12687 , \12694 );
and \U$6237 ( \12696 , \12661 , \12695 );
buf \U$6238 ( \12697 , \12696 );
or \U$6239 ( \12698 , \12659 , \12697 );
_DC g485d ( \12699_nG485d , \12623 , \12698 );
buf \U$6240 ( \12700 , \12699_nG485d );
xor \U$6241 ( \12701 , \12190 , \12700 );
buf \U$6242 ( \12702 , RIb7b9590_247);
and \U$6243 ( \12703 , \7126 , \12216 );
and \U$6244 ( \12704 , \7128 , \12243 );
and \U$6245 ( \12705 , \8338 , \12270 );
and \U$6246 ( \12706 , \8340 , \12297 );
and \U$6247 ( \12707 , \8342 , \12324 );
and \U$6248 ( \12708 , \8344 , \12351 );
and \U$6249 ( \12709 , \8346 , \12378 );
and \U$6250 ( \12710 , \8348 , \12405 );
and \U$6251 ( \12711 , \8350 , \12432 );
and \U$6252 ( \12712 , \8352 , \12459 );
and \U$6253 ( \12713 , \8354 , \12486 );
and \U$6254 ( \12714 , \8356 , \12513 );
and \U$6255 ( \12715 , \8358 , \12540 );
and \U$6256 ( \12716 , \8360 , \12567 );
and \U$6257 ( \12717 , \8362 , \12594 );
and \U$6258 ( \12718 , \8364 , \12621 );
or \U$6259 ( \12719 , \12703 , \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 , \12718 );
_DC g4872 ( \12720_nG4872 , \12719 , \12698 );
buf \U$6260 ( \12721 , \12720_nG4872 );
xor \U$6261 ( \12722 , \12702 , \12721 );
or \U$6262 ( \12723 , \12701 , \12722 );
buf \U$6263 ( \12724 , RIb7b9518_248);
and \U$6264 ( \12725 , \7136 , \12216 );
and \U$6265 ( \12726 , \7138 , \12243 );
and \U$6266 ( \12727 , \8374 , \12270 );
and \U$6267 ( \12728 , \8376 , \12297 );
and \U$6268 ( \12729 , \8378 , \12324 );
and \U$6269 ( \12730 , \8380 , \12351 );
and \U$6270 ( \12731 , \8382 , \12378 );
and \U$6271 ( \12732 , \8384 , \12405 );
and \U$6272 ( \12733 , \8386 , \12432 );
and \U$6273 ( \12734 , \8388 , \12459 );
and \U$6274 ( \12735 , \8390 , \12486 );
and \U$6275 ( \12736 , \8392 , \12513 );
and \U$6276 ( \12737 , \8394 , \12540 );
and \U$6277 ( \12738 , \8396 , \12567 );
and \U$6278 ( \12739 , \8398 , \12594 );
and \U$6279 ( \12740 , \8400 , \12621 );
or \U$6280 ( \12741 , \12725 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 );
_DC g4888 ( \12742_nG4888 , \12741 , \12698 );
buf \U$6281 ( \12743 , \12742_nG4888 );
xor \U$6282 ( \12744 , \12724 , \12743 );
or \U$6283 ( \12745 , \12723 , \12744 );
buf \U$6284 ( \12746 , RIb7b94a0_249);
and \U$6285 ( \12747 , \7146 , \12216 );
and \U$6286 ( \12748 , \7148 , \12243 );
and \U$6287 ( \12749 , \8410 , \12270 );
and \U$6288 ( \12750 , \8412 , \12297 );
and \U$6289 ( \12751 , \8414 , \12324 );
and \U$6290 ( \12752 , \8416 , \12351 );
and \U$6291 ( \12753 , \8418 , \12378 );
and \U$6292 ( \12754 , \8420 , \12405 );
and \U$6293 ( \12755 , \8422 , \12432 );
and \U$6294 ( \12756 , \8424 , \12459 );
and \U$6295 ( \12757 , \8426 , \12486 );
and \U$6296 ( \12758 , \8428 , \12513 );
and \U$6297 ( \12759 , \8430 , \12540 );
and \U$6298 ( \12760 , \8432 , \12567 );
and \U$6299 ( \12761 , \8434 , \12594 );
and \U$6300 ( \12762 , \8436 , \12621 );
or \U$6301 ( \12763 , \12747 , \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 );
_DC g489e ( \12764_nG489e , \12763 , \12698 );
buf \U$6302 ( \12765 , \12764_nG489e );
xor \U$6303 ( \12766 , \12746 , \12765 );
or \U$6304 ( \12767 , \12745 , \12766 );
buf \U$6305 ( \12768 , RIb7b9428_250);
and \U$6306 ( \12769 , \7156 , \12216 );
and \U$6307 ( \12770 , \7158 , \12243 );
and \U$6308 ( \12771 , \8446 , \12270 );
and \U$6309 ( \12772 , \8448 , \12297 );
and \U$6310 ( \12773 , \8450 , \12324 );
and \U$6311 ( \12774 , \8452 , \12351 );
and \U$6312 ( \12775 , \8454 , \12378 );
and \U$6313 ( \12776 , \8456 , \12405 );
and \U$6314 ( \12777 , \8458 , \12432 );
and \U$6315 ( \12778 , \8460 , \12459 );
and \U$6316 ( \12779 , \8462 , \12486 );
and \U$6317 ( \12780 , \8464 , \12513 );
and \U$6318 ( \12781 , \8466 , \12540 );
and \U$6319 ( \12782 , \8468 , \12567 );
and \U$6320 ( \12783 , \8470 , \12594 );
and \U$6321 ( \12784 , \8472 , \12621 );
or \U$6322 ( \12785 , \12769 , \12770 , \12771 , \12772 , \12773 , \12774 , \12775 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 );
_DC g48b4 ( \12786_nG48b4 , \12785 , \12698 );
buf \U$6323 ( \12787 , \12786_nG48b4 );
xor \U$6324 ( \12788 , \12768 , \12787 );
or \U$6325 ( \12789 , \12767 , \12788 );
buf \U$6326 ( \12790 , RIb7b93b0_251);
and \U$6327 ( \12791 , \7166 , \12216 );
and \U$6328 ( \12792 , \7168 , \12243 );
and \U$6329 ( \12793 , \8482 , \12270 );
and \U$6330 ( \12794 , \8484 , \12297 );
and \U$6331 ( \12795 , \8486 , \12324 );
and \U$6332 ( \12796 , \8488 , \12351 );
and \U$6333 ( \12797 , \8490 , \12378 );
and \U$6334 ( \12798 , \8492 , \12405 );
and \U$6335 ( \12799 , \8494 , \12432 );
and \U$6336 ( \12800 , \8496 , \12459 );
and \U$6337 ( \12801 , \8498 , \12486 );
and \U$6338 ( \12802 , \8500 , \12513 );
and \U$6339 ( \12803 , \8502 , \12540 );
and \U$6340 ( \12804 , \8504 , \12567 );
and \U$6341 ( \12805 , \8506 , \12594 );
and \U$6342 ( \12806 , \8508 , \12621 );
or \U$6343 ( \12807 , \12791 , \12792 , \12793 , \12794 , \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801 , \12802 , \12803 , \12804 , \12805 , \12806 );
_DC g48ca ( \12808_nG48ca , \12807 , \12698 );
buf \U$6344 ( \12809 , \12808_nG48ca );
xor \U$6345 ( \12810 , \12790 , \12809 );
or \U$6346 ( \12811 , \12789 , \12810 );
buf \U$6347 ( \12812 , RIb7af720_252);
and \U$6348 ( \12813 , \7176 , \12216 );
and \U$6349 ( \12814 , \7178 , \12243 );
and \U$6350 ( \12815 , \8518 , \12270 );
and \U$6351 ( \12816 , \8520 , \12297 );
and \U$6352 ( \12817 , \8522 , \12324 );
and \U$6353 ( \12818 , \8524 , \12351 );
and \U$6354 ( \12819 , \8526 , \12378 );
and \U$6355 ( \12820 , \8528 , \12405 );
and \U$6356 ( \12821 , \8530 , \12432 );
and \U$6357 ( \12822 , \8532 , \12459 );
and \U$6358 ( \12823 , \8534 , \12486 );
and \U$6359 ( \12824 , \8536 , \12513 );
and \U$6360 ( \12825 , \8538 , \12540 );
and \U$6361 ( \12826 , \8540 , \12567 );
and \U$6362 ( \12827 , \8542 , \12594 );
and \U$6363 ( \12828 , \8544 , \12621 );
or \U$6364 ( \12829 , \12813 , \12814 , \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 , \12825 , \12826 , \12827 , \12828 );
_DC g48e0 ( \12830_nG48e0 , \12829 , \12698 );
buf \U$6365 ( \12831 , \12830_nG48e0 );
xor \U$6366 ( \12832 , \12812 , \12831 );
or \U$6367 ( \12833 , \12811 , \12832 );
buf \U$6368 ( \12834 , RIb7af6a8_253);
and \U$6369 ( \12835 , \7186 , \12216 );
and \U$6370 ( \12836 , \7188 , \12243 );
and \U$6371 ( \12837 , \8554 , \12270 );
and \U$6372 ( \12838 , \8556 , \12297 );
and \U$6373 ( \12839 , \8558 , \12324 );
and \U$6374 ( \12840 , \8560 , \12351 );
and \U$6375 ( \12841 , \8562 , \12378 );
and \U$6376 ( \12842 , \8564 , \12405 );
and \U$6377 ( \12843 , \8566 , \12432 );
and \U$6378 ( \12844 , \8568 , \12459 );
and \U$6379 ( \12845 , \8570 , \12486 );
and \U$6380 ( \12846 , \8572 , \12513 );
and \U$6381 ( \12847 , \8574 , \12540 );
and \U$6382 ( \12848 , \8576 , \12567 );
and \U$6383 ( \12849 , \8578 , \12594 );
and \U$6384 ( \12850 , \8580 , \12621 );
or \U$6385 ( \12851 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844 , \12845 , \12846 , \12847 , \12848 , \12849 , \12850 );
_DC g48f6 ( \12852_nG48f6 , \12851 , \12698 );
buf \U$6386 ( \12853 , \12852_nG48f6 );
xor \U$6387 ( \12854 , \12834 , \12853 );
or \U$6388 ( \12855 , \12833 , \12854 );
not \U$6389 ( \12856 , \12855 );
buf \U$6390 ( \12857 , \12856 );
and \U$6391 ( \12858 , \12189 , \12857 );
buf \U$6392 ( \12859 , RIb7af630_254);
buf \U$6393 ( \12860 , \11675 );
buf \U$6394 ( \12861 , \11675 );
buf \U$6395 ( \12862 , \11675 );
buf \U$6396 ( \12863 , \11675 );
buf \U$6397 ( \12864 , \11675 );
buf \U$6398 ( \12865 , \11675 );
buf \U$6399 ( \12866 , \11675 );
buf \U$6400 ( \12867 , \11675 );
buf \U$6401 ( \12868 , \11675 );
buf \U$6402 ( \12869 , \11675 );
buf \U$6403 ( \12870 , \11675 );
buf \U$6404 ( \12871 , \11675 );
buf \U$6405 ( \12872 , \11675 );
buf \U$6406 ( \12873 , \11675 );
buf \U$6407 ( \12874 , \11675 );
buf \U$6408 ( \12875 , \11675 );
buf \U$6409 ( \12876 , \11675 );
buf \U$6410 ( \12877 , \11675 );
buf \U$6411 ( \12878 , \11675 );
buf \U$6412 ( \12879 , \11675 );
buf \U$6413 ( \12880 , \11675 );
buf \U$6414 ( \12881 , \11675 );
buf \U$6415 ( \12882 , \11675 );
buf \U$6416 ( \12883 , \11675 );
buf \U$6417 ( \12884 , \11675 );
nor \U$6418 ( \12885 , \11662 , \11663 , \11664 , \11665 , \11669 , \11672 , \11675 , \12860 , \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 , \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 , \12883 , \12884 );
and \U$6419 ( \12886 , \7198 , \12885 );
buf \U$6420 ( \12887 , \11675 );
buf \U$6421 ( \12888 , \11675 );
buf \U$6422 ( \12889 , \11675 );
buf \U$6423 ( \12890 , \11675 );
buf \U$6424 ( \12891 , \11675 );
buf \U$6425 ( \12892 , \11675 );
buf \U$6426 ( \12893 , \11675 );
buf \U$6427 ( \12894 , \11675 );
buf \U$6428 ( \12895 , \11675 );
buf \U$6429 ( \12896 , \11675 );
buf \U$6430 ( \12897 , \11675 );
buf \U$6431 ( \12898 , \11675 );
buf \U$6432 ( \12899 , \11675 );
buf \U$6433 ( \12900 , \11675 );
buf \U$6434 ( \12901 , \11675 );
buf \U$6435 ( \12902 , \11675 );
buf \U$6436 ( \12903 , \11675 );
buf \U$6437 ( \12904 , \11675 );
buf \U$6438 ( \12905 , \11675 );
buf \U$6439 ( \12906 , \11675 );
buf \U$6440 ( \12907 , \11675 );
buf \U$6441 ( \12908 , \11675 );
buf \U$6442 ( \12909 , \11675 );
buf \U$6443 ( \12910 , \11675 );
buf \U$6444 ( \12911 , \11675 );
nor \U$6445 ( \12912 , \11703 , \11704 , \11705 , \11706 , \11668 , \11672 , \11675 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 , \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 , \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 );
and \U$6446 ( \12913 , \7200 , \12912 );
buf \U$6447 ( \12914 , \11675 );
buf \U$6448 ( \12915 , \11675 );
buf \U$6449 ( \12916 , \11675 );
buf \U$6450 ( \12917 , \11675 );
buf \U$6451 ( \12918 , \11675 );
buf \U$6452 ( \12919 , \11675 );
buf \U$6453 ( \12920 , \11675 );
buf \U$6454 ( \12921 , \11675 );
buf \U$6455 ( \12922 , \11675 );
buf \U$6456 ( \12923 , \11675 );
buf \U$6457 ( \12924 , \11675 );
buf \U$6458 ( \12925 , \11675 );
buf \U$6459 ( \12926 , \11675 );
buf \U$6460 ( \12927 , \11675 );
buf \U$6461 ( \12928 , \11675 );
buf \U$6462 ( \12929 , \11675 );
buf \U$6463 ( \12930 , \11675 );
buf \U$6464 ( \12931 , \11675 );
buf \U$6465 ( \12932 , \11675 );
buf \U$6466 ( \12933 , \11675 );
buf \U$6467 ( \12934 , \11675 );
buf \U$6468 ( \12935 , \11675 );
buf \U$6469 ( \12936 , \11675 );
buf \U$6470 ( \12937 , \11675 );
buf \U$6471 ( \12938 , \11675 );
nor \U$6472 ( \12939 , \11662 , \11704 , \11705 , \11706 , \11668 , \11672 , \11675 , \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 , \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 , \12935 , \12936 , \12937 , \12938 );
and \U$6473 ( \12940 , \8645 , \12939 );
buf \U$6474 ( \12941 , \11675 );
buf \U$6475 ( \12942 , \11675 );
buf \U$6476 ( \12943 , \11675 );
buf \U$6477 ( \12944 , \11675 );
buf \U$6478 ( \12945 , \11675 );
buf \U$6479 ( \12946 , \11675 );
buf \U$6480 ( \12947 , \11675 );
buf \U$6481 ( \12948 , \11675 );
buf \U$6482 ( \12949 , \11675 );
buf \U$6483 ( \12950 , \11675 );
buf \U$6484 ( \12951 , \11675 );
buf \U$6485 ( \12952 , \11675 );
buf \U$6486 ( \12953 , \11675 );
buf \U$6487 ( \12954 , \11675 );
buf \U$6488 ( \12955 , \11675 );
buf \U$6489 ( \12956 , \11675 );
buf \U$6490 ( \12957 , \11675 );
buf \U$6491 ( \12958 , \11675 );
buf \U$6492 ( \12959 , \11675 );
buf \U$6493 ( \12960 , \11675 );
buf \U$6494 ( \12961 , \11675 );
buf \U$6495 ( \12962 , \11675 );
buf \U$6496 ( \12963 , \11675 );
buf \U$6497 ( \12964 , \11675 );
buf \U$6498 ( \12965 , \11675 );
nor \U$6499 ( \12966 , \11703 , \11663 , \11705 , \11706 , \11668 , \11672 , \11675 , \12941 , \12942 , \12943 , \12944 , \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 , \12952 , \12953 , \12954 , \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 , \12965 );
and \U$6500 ( \12967 , \8673 , \12966 );
buf \U$6501 ( \12968 , \11675 );
buf \U$6502 ( \12969 , \11675 );
buf \U$6503 ( \12970 , \11675 );
buf \U$6504 ( \12971 , \11675 );
buf \U$6505 ( \12972 , \11675 );
buf \U$6506 ( \12973 , \11675 );
buf \U$6507 ( \12974 , \11675 );
buf \U$6508 ( \12975 , \11675 );
buf \U$6509 ( \12976 , \11675 );
buf \U$6510 ( \12977 , \11675 );
buf \U$6511 ( \12978 , \11675 );
buf \U$6512 ( \12979 , \11675 );
buf \U$6513 ( \12980 , \11675 );
buf \U$6514 ( \12981 , \11675 );
buf \U$6515 ( \12982 , \11675 );
buf \U$6516 ( \12983 , \11675 );
buf \U$6517 ( \12984 , \11675 );
buf \U$6518 ( \12985 , \11675 );
buf \U$6519 ( \12986 , \11675 );
buf \U$6520 ( \12987 , \11675 );
buf \U$6521 ( \12988 , \11675 );
buf \U$6522 ( \12989 , \11675 );
buf \U$6523 ( \12990 , \11675 );
buf \U$6524 ( \12991 , \11675 );
buf \U$6525 ( \12992 , \11675 );
nor \U$6526 ( \12993 , \11662 , \11663 , \11705 , \11706 , \11668 , \11672 , \11675 , \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 , \12975 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 , \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 );
and \U$6527 ( \12994 , \8701 , \12993 );
buf \U$6528 ( \12995 , \11675 );
buf \U$6529 ( \12996 , \11675 );
buf \U$6530 ( \12997 , \11675 );
buf \U$6531 ( \12998 , \11675 );
buf \U$6532 ( \12999 , \11675 );
buf \U$6533 ( \13000 , \11675 );
buf \U$6534 ( \13001 , \11675 );
buf \U$6535 ( \13002 , \11675 );
buf \U$6536 ( \13003 , \11675 );
buf \U$6537 ( \13004 , \11675 );
buf \U$6538 ( \13005 , \11675 );
buf \U$6539 ( \13006 , \11675 );
buf \U$6540 ( \13007 , \11675 );
buf \U$6541 ( \13008 , \11675 );
buf \U$6542 ( \13009 , \11675 );
buf \U$6543 ( \13010 , \11675 );
buf \U$6544 ( \13011 , \11675 );
buf \U$6545 ( \13012 , \11675 );
buf \U$6546 ( \13013 , \11675 );
buf \U$6547 ( \13014 , \11675 );
buf \U$6548 ( \13015 , \11675 );
buf \U$6549 ( \13016 , \11675 );
buf \U$6550 ( \13017 , \11675 );
buf \U$6551 ( \13018 , \11675 );
buf \U$6552 ( \13019 , \11675 );
nor \U$6553 ( \13020 , \11703 , \11704 , \11664 , \11706 , \11668 , \11672 , \11675 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 , \13005 , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 , \13015 , \13016 , \13017 , \13018 , \13019 );
and \U$6554 ( \13021 , \8729 , \13020 );
buf \U$6555 ( \13022 , \11675 );
buf \U$6556 ( \13023 , \11675 );
buf \U$6557 ( \13024 , \11675 );
buf \U$6558 ( \13025 , \11675 );
buf \U$6559 ( \13026 , \11675 );
buf \U$6560 ( \13027 , \11675 );
buf \U$6561 ( \13028 , \11675 );
buf \U$6562 ( \13029 , \11675 );
buf \U$6563 ( \13030 , \11675 );
buf \U$6564 ( \13031 , \11675 );
buf \U$6565 ( \13032 , \11675 );
buf \U$6566 ( \13033 , \11675 );
buf \U$6567 ( \13034 , \11675 );
buf \U$6568 ( \13035 , \11675 );
buf \U$6569 ( \13036 , \11675 );
buf \U$6570 ( \13037 , \11675 );
buf \U$6571 ( \13038 , \11675 );
buf \U$6572 ( \13039 , \11675 );
buf \U$6573 ( \13040 , \11675 );
buf \U$6574 ( \13041 , \11675 );
buf \U$6575 ( \13042 , \11675 );
buf \U$6576 ( \13043 , \11675 );
buf \U$6577 ( \13044 , \11675 );
buf \U$6578 ( \13045 , \11675 );
buf \U$6579 ( \13046 , \11675 );
nor \U$6580 ( \13047 , \11662 , \11704 , \11664 , \11706 , \11668 , \11672 , \11675 , \13022 , \13023 , \13024 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 , \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 , \13045 , \13046 );
and \U$6581 ( \13048 , \8757 , \13047 );
buf \U$6582 ( \13049 , \11675 );
buf \U$6583 ( \13050 , \11675 );
buf \U$6584 ( \13051 , \11675 );
buf \U$6585 ( \13052 , \11675 );
buf \U$6586 ( \13053 , \11675 );
buf \U$6587 ( \13054 , \11675 );
buf \U$6588 ( \13055 , \11675 );
buf \U$6589 ( \13056 , \11675 );
buf \U$6590 ( \13057 , \11675 );
buf \U$6591 ( \13058 , \11675 );
buf \U$6592 ( \13059 , \11675 );
buf \U$6593 ( \13060 , \11675 );
buf \U$6594 ( \13061 , \11675 );
buf \U$6595 ( \13062 , \11675 );
buf \U$6596 ( \13063 , \11675 );
buf \U$6597 ( \13064 , \11675 );
buf \U$6598 ( \13065 , \11675 );
buf \U$6599 ( \13066 , \11675 );
buf \U$6600 ( \13067 , \11675 );
buf \U$6601 ( \13068 , \11675 );
buf \U$6602 ( \13069 , \11675 );
buf \U$6603 ( \13070 , \11675 );
buf \U$6604 ( \13071 , \11675 );
buf \U$6605 ( \13072 , \11675 );
buf \U$6606 ( \13073 , \11675 );
nor \U$6607 ( \13074 , \11703 , \11663 , \11664 , \11706 , \11668 , \11672 , \11675 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 , \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 , \13062 , \13063 , \13064 , \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 , \13072 , \13073 );
and \U$6608 ( \13075 , \8785 , \13074 );
buf \U$6609 ( \13076 , \11675 );
buf \U$6610 ( \13077 , \11675 );
buf \U$6611 ( \13078 , \11675 );
buf \U$6612 ( \13079 , \11675 );
buf \U$6613 ( \13080 , \11675 );
buf \U$6614 ( \13081 , \11675 );
buf \U$6615 ( \13082 , \11675 );
buf \U$6616 ( \13083 , \11675 );
buf \U$6617 ( \13084 , \11675 );
buf \U$6618 ( \13085 , \11675 );
buf \U$6619 ( \13086 , \11675 );
buf \U$6620 ( \13087 , \11675 );
buf \U$6621 ( \13088 , \11675 );
buf \U$6622 ( \13089 , \11675 );
buf \U$6623 ( \13090 , \11675 );
buf \U$6624 ( \13091 , \11675 );
buf \U$6625 ( \13092 , \11675 );
buf \U$6626 ( \13093 , \11675 );
buf \U$6627 ( \13094 , \11675 );
buf \U$6628 ( \13095 , \11675 );
buf \U$6629 ( \13096 , \11675 );
buf \U$6630 ( \13097 , \11675 );
buf \U$6631 ( \13098 , \11675 );
buf \U$6632 ( \13099 , \11675 );
buf \U$6633 ( \13100 , \11675 );
nor \U$6634 ( \13101 , \11662 , \11663 , \11664 , \11706 , \11668 , \11672 , \11675 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 , \13082 , \13083 , \13084 , \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 , \13092 , \13093 , \13094 , \13095 , \13096 , \13097 , \13098 , \13099 , \13100 );
and \U$6635 ( \13102 , \8813 , \13101 );
buf \U$6636 ( \13103 , \11675 );
buf \U$6637 ( \13104 , \11675 );
buf \U$6638 ( \13105 , \11675 );
buf \U$6639 ( \13106 , \11675 );
buf \U$6640 ( \13107 , \11675 );
buf \U$6641 ( \13108 , \11675 );
buf \U$6642 ( \13109 , \11675 );
buf \U$6643 ( \13110 , \11675 );
buf \U$6644 ( \13111 , \11675 );
buf \U$6645 ( \13112 , \11675 );
buf \U$6646 ( \13113 , \11675 );
buf \U$6647 ( \13114 , \11675 );
buf \U$6648 ( \13115 , \11675 );
buf \U$6649 ( \13116 , \11675 );
buf \U$6650 ( \13117 , \11675 );
buf \U$6651 ( \13118 , \11675 );
buf \U$6652 ( \13119 , \11675 );
buf \U$6653 ( \13120 , \11675 );
buf \U$6654 ( \13121 , \11675 );
buf \U$6655 ( \13122 , \11675 );
buf \U$6656 ( \13123 , \11675 );
buf \U$6657 ( \13124 , \11675 );
buf \U$6658 ( \13125 , \11675 );
buf \U$6659 ( \13126 , \11675 );
buf \U$6660 ( \13127 , \11675 );
nor \U$6661 ( \13128 , \11703 , \11704 , \11705 , \11665 , \11668 , \11672 , \11675 , \13103 , \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 , \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 , \13125 , \13126 , \13127 );
and \U$6662 ( \13129 , \8841 , \13128 );
buf \U$6663 ( \13130 , \11675 );
buf \U$6664 ( \13131 , \11675 );
buf \U$6665 ( \13132 , \11675 );
buf \U$6666 ( \13133 , \11675 );
buf \U$6667 ( \13134 , \11675 );
buf \U$6668 ( \13135 , \11675 );
buf \U$6669 ( \13136 , \11675 );
buf \U$6670 ( \13137 , \11675 );
buf \U$6671 ( \13138 , \11675 );
buf \U$6672 ( \13139 , \11675 );
buf \U$6673 ( \13140 , \11675 );
buf \U$6674 ( \13141 , \11675 );
buf \U$6675 ( \13142 , \11675 );
buf \U$6676 ( \13143 , \11675 );
buf \U$6677 ( \13144 , \11675 );
buf \U$6678 ( \13145 , \11675 );
buf \U$6679 ( \13146 , \11675 );
buf \U$6680 ( \13147 , \11675 );
buf \U$6681 ( \13148 , \11675 );
buf \U$6682 ( \13149 , \11675 );
buf \U$6683 ( \13150 , \11675 );
buf \U$6684 ( \13151 , \11675 );
buf \U$6685 ( \13152 , \11675 );
buf \U$6686 ( \13153 , \11675 );
buf \U$6687 ( \13154 , \11675 );
nor \U$6688 ( \13155 , \11662 , \11704 , \11705 , \11665 , \11668 , \11672 , \11675 , \13130 , \13131 , \13132 , \13133 , \13134 , \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 );
and \U$6689 ( \13156 , \8869 , \13155 );
buf \U$6690 ( \13157 , \11675 );
buf \U$6691 ( \13158 , \11675 );
buf \U$6692 ( \13159 , \11675 );
buf \U$6693 ( \13160 , \11675 );
buf \U$6694 ( \13161 , \11675 );
buf \U$6695 ( \13162 , \11675 );
buf \U$6696 ( \13163 , \11675 );
buf \U$6697 ( \13164 , \11675 );
buf \U$6698 ( \13165 , \11675 );
buf \U$6699 ( \13166 , \11675 );
buf \U$6700 ( \13167 , \11675 );
buf \U$6701 ( \13168 , \11675 );
buf \U$6702 ( \13169 , \11675 );
buf \U$6703 ( \13170 , \11675 );
buf \U$6704 ( \13171 , \11675 );
buf \U$6705 ( \13172 , \11675 );
buf \U$6706 ( \13173 , \11675 );
buf \U$6707 ( \13174 , \11675 );
buf \U$6708 ( \13175 , \11675 );
buf \U$6709 ( \13176 , \11675 );
buf \U$6710 ( \13177 , \11675 );
buf \U$6711 ( \13178 , \11675 );
buf \U$6712 ( \13179 , \11675 );
buf \U$6713 ( \13180 , \11675 );
buf \U$6714 ( \13181 , \11675 );
nor \U$6715 ( \13182 , \11703 , \11663 , \11705 , \11665 , \11668 , \11672 , \11675 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 , \13163 , \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 , \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 );
and \U$6716 ( \13183 , \8897 , \13182 );
buf \U$6717 ( \13184 , \11675 );
buf \U$6718 ( \13185 , \11675 );
buf \U$6719 ( \13186 , \11675 );
buf \U$6720 ( \13187 , \11675 );
buf \U$6721 ( \13188 , \11675 );
buf \U$6722 ( \13189 , \11675 );
buf \U$6723 ( \13190 , \11675 );
buf \U$6724 ( \13191 , \11675 );
buf \U$6725 ( \13192 , \11675 );
buf \U$6726 ( \13193 , \11675 );
buf \U$6727 ( \13194 , \11675 );
buf \U$6728 ( \13195 , \11675 );
buf \U$6729 ( \13196 , \11675 );
buf \U$6730 ( \13197 , \11675 );
buf \U$6731 ( \13198 , \11675 );
buf \U$6732 ( \13199 , \11675 );
buf \U$6733 ( \13200 , \11675 );
buf \U$6734 ( \13201 , \11675 );
buf \U$6735 ( \13202 , \11675 );
buf \U$6736 ( \13203 , \11675 );
buf \U$6737 ( \13204 , \11675 );
buf \U$6738 ( \13205 , \11675 );
buf \U$6739 ( \13206 , \11675 );
buf \U$6740 ( \13207 , \11675 );
buf \U$6741 ( \13208 , \11675 );
nor \U$6742 ( \13209 , \11662 , \11663 , \11705 , \11665 , \11668 , \11672 , \11675 , \13184 , \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 , \13205 , \13206 , \13207 , \13208 );
and \U$6743 ( \13210 , \8925 , \13209 );
buf \U$6744 ( \13211 , \11675 );
buf \U$6745 ( \13212 , \11675 );
buf \U$6746 ( \13213 , \11675 );
buf \U$6747 ( \13214 , \11675 );
buf \U$6748 ( \13215 , \11675 );
buf \U$6749 ( \13216 , \11675 );
buf \U$6750 ( \13217 , \11675 );
buf \U$6751 ( \13218 , \11675 );
buf \U$6752 ( \13219 , \11675 );
buf \U$6753 ( \13220 , \11675 );
buf \U$6754 ( \13221 , \11675 );
buf \U$6755 ( \13222 , \11675 );
buf \U$6756 ( \13223 , \11675 );
buf \U$6757 ( \13224 , \11675 );
buf \U$6758 ( \13225 , \11675 );
buf \U$6759 ( \13226 , \11675 );
buf \U$6760 ( \13227 , \11675 );
buf \U$6761 ( \13228 , \11675 );
buf \U$6762 ( \13229 , \11675 );
buf \U$6763 ( \13230 , \11675 );
buf \U$6764 ( \13231 , \11675 );
buf \U$6765 ( \13232 , \11675 );
buf \U$6766 ( \13233 , \11675 );
buf \U$6767 ( \13234 , \11675 );
buf \U$6768 ( \13235 , \11675 );
nor \U$6769 ( \13236 , \11703 , \11704 , \11664 , \11665 , \11668 , \11672 , \11675 , \13211 , \13212 , \13213 , \13214 , \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 , \13235 );
and \U$6770 ( \13237 , \8953 , \13236 );
buf \U$6771 ( \13238 , \11675 );
buf \U$6772 ( \13239 , \11675 );
buf \U$6773 ( \13240 , \11675 );
buf \U$6774 ( \13241 , \11675 );
buf \U$6775 ( \13242 , \11675 );
buf \U$6776 ( \13243 , \11675 );
buf \U$6777 ( \13244 , \11675 );
buf \U$6778 ( \13245 , \11675 );
buf \U$6779 ( \13246 , \11675 );
buf \U$6780 ( \13247 , \11675 );
buf \U$6781 ( \13248 , \11675 );
buf \U$6782 ( \13249 , \11675 );
buf \U$6783 ( \13250 , \11675 );
buf \U$6784 ( \13251 , \11675 );
buf \U$6785 ( \13252 , \11675 );
buf \U$6786 ( \13253 , \11675 );
buf \U$6787 ( \13254 , \11675 );
buf \U$6788 ( \13255 , \11675 );
buf \U$6789 ( \13256 , \11675 );
buf \U$6790 ( \13257 , \11675 );
buf \U$6791 ( \13258 , \11675 );
buf \U$6792 ( \13259 , \11675 );
buf \U$6793 ( \13260 , \11675 );
buf \U$6794 ( \13261 , \11675 );
buf \U$6795 ( \13262 , \11675 );
nor \U$6796 ( \13263 , \11662 , \11704 , \11664 , \11665 , \11668 , \11672 , \11675 , \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 );
and \U$6797 ( \13264 , \8981 , \13263 );
buf \U$6798 ( \13265 , \11675 );
buf \U$6799 ( \13266 , \11675 );
buf \U$6800 ( \13267 , \11675 );
buf \U$6801 ( \13268 , \11675 );
buf \U$6802 ( \13269 , \11675 );
buf \U$6803 ( \13270 , \11675 );
buf \U$6804 ( \13271 , \11675 );
buf \U$6805 ( \13272 , \11675 );
buf \U$6806 ( \13273 , \11675 );
buf \U$6807 ( \13274 , \11675 );
buf \U$6808 ( \13275 , \11675 );
buf \U$6809 ( \13276 , \11675 );
buf \U$6810 ( \13277 , \11675 );
buf \U$6811 ( \13278 , \11675 );
buf \U$6812 ( \13279 , \11675 );
buf \U$6813 ( \13280 , \11675 );
buf \U$6814 ( \13281 , \11675 );
buf \U$6815 ( \13282 , \11675 );
buf \U$6816 ( \13283 , \11675 );
buf \U$6817 ( \13284 , \11675 );
buf \U$6818 ( \13285 , \11675 );
buf \U$6819 ( \13286 , \11675 );
buf \U$6820 ( \13287 , \11675 );
buf \U$6821 ( \13288 , \11675 );
buf \U$6822 ( \13289 , \11675 );
nor \U$6823 ( \13290 , \11703 , \11663 , \11664 , \11665 , \11668 , \11672 , \11675 , \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 , \13285 , \13286 , \13287 , \13288 , \13289 );
and \U$6824 ( \13291 , \9009 , \13290 );
or \U$6825 ( \13292 , \12886 , \12913 , \12940 , \12967 , \12994 , \13021 , \13048 , \13075 , \13102 , \13129 , \13156 , \13183 , \13210 , \13237 , \13264 , \13291 );
buf \U$6826 ( \13293 , \11675 );
not \U$6827 ( \13294 , \13293 );
buf \U$6828 ( \13295 , \11663 );
buf \U$6829 ( \13296 , \11664 );
buf \U$6830 ( \13297 , \11665 );
buf \U$6831 ( \13298 , \11668 );
buf \U$6832 ( \13299 , \11672 );
buf \U$6833 ( \13300 , \11675 );
buf \U$6834 ( \13301 , \11675 );
buf \U$6835 ( \13302 , \11675 );
buf \U$6836 ( \13303 , \11675 );
buf \U$6837 ( \13304 , \11675 );
buf \U$6838 ( \13305 , \11675 );
buf \U$6839 ( \13306 , \11675 );
buf \U$6840 ( \13307 , \11675 );
buf \U$6841 ( \13308 , \11675 );
buf \U$6842 ( \13309 , \11675 );
buf \U$6843 ( \13310 , \11675 );
buf \U$6844 ( \13311 , \11675 );
buf \U$6845 ( \13312 , \11675 );
buf \U$6846 ( \13313 , \11675 );
buf \U$6847 ( \13314 , \11675 );
buf \U$6848 ( \13315 , \11675 );
buf \U$6849 ( \13316 , \11675 );
buf \U$6850 ( \13317 , \11675 );
buf \U$6851 ( \13318 , \11675 );
buf \U$6852 ( \13319 , \11675 );
buf \U$6853 ( \13320 , \11675 );
buf \U$6854 ( \13321 , \11675 );
buf \U$6855 ( \13322 , \11675 );
buf \U$6856 ( \13323 , \11675 );
buf \U$6857 ( \13324 , \11675 );
buf \U$6858 ( \13325 , \11662 );
or \U$6859 ( \13326 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 , \13312 , \13313 , \13314 , \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 , \13322 , \13323 , \13324 , \13325 );
nand \U$6860 ( \13327 , \13294 , \13326 );
buf \U$6861 ( \13328 , \13327 );
buf \U$6862 ( \13329 , \11675 );
not \U$6863 ( \13330 , \13329 );
buf \U$6864 ( \13331 , \11672 );
buf \U$6865 ( \13332 , \11675 );
buf \U$6866 ( \13333 , \11675 );
buf \U$6867 ( \13334 , \11675 );
buf \U$6868 ( \13335 , \11675 );
buf \U$6869 ( \13336 , \11675 );
buf \U$6870 ( \13337 , \11675 );
buf \U$6871 ( \13338 , \11675 );
buf \U$6872 ( \13339 , \11675 );
buf \U$6873 ( \13340 , \11675 );
buf \U$6874 ( \13341 , \11675 );
buf \U$6875 ( \13342 , \11675 );
buf \U$6876 ( \13343 , \11675 );
buf \U$6877 ( \13344 , \11675 );
buf \U$6878 ( \13345 , \11675 );
buf \U$6879 ( \13346 , \11675 );
buf \U$6880 ( \13347 , \11675 );
buf \U$6881 ( \13348 , \11675 );
buf \U$6882 ( \13349 , \11675 );
buf \U$6883 ( \13350 , \11675 );
buf \U$6884 ( \13351 , \11675 );
buf \U$6885 ( \13352 , \11675 );
buf \U$6886 ( \13353 , \11675 );
buf \U$6887 ( \13354 , \11675 );
buf \U$6888 ( \13355 , \11675 );
buf \U$6889 ( \13356 , \11675 );
buf \U$6890 ( \13357 , \11668 );
buf \U$6891 ( \13358 , \11662 );
buf \U$6892 ( \13359 , \11663 );
buf \U$6893 ( \13360 , \11664 );
buf \U$6894 ( \13361 , \11665 );
or \U$6895 ( \13362 , \13358 , \13359 , \13360 , \13361 );
and \U$6896 ( \13363 , \13357 , \13362 );
or \U$6897 ( \13364 , \13331 , \13332 , \13333 , \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 , \13345 , \13346 , \13347 , \13348 , \13349 , \13350 , \13351 , \13352 , \13353 , \13354 , \13355 , \13356 , \13363 );
and \U$6898 ( \13365 , \13330 , \13364 );
buf \U$6899 ( \13366 , \13365 );
or \U$6900 ( \13367 , \13328 , \13366 );
_DC g4afa ( \13368_nG4afa , \13292 , \13367 );
buf \U$6901 ( \13369 , \13368_nG4afa );
xor \U$6902 ( \13370 , \12859 , \13369 );
buf \U$6903 ( \13371 , RIb7af5b8_255);
and \U$6904 ( \13372 , \7207 , \12885 );
and \U$6905 ( \13373 , \7209 , \12912 );
and \U$6906 ( \13374 , \9119 , \12939 );
and \U$6907 ( \13375 , \9121 , \12966 );
and \U$6908 ( \13376 , \9123 , \12993 );
and \U$6909 ( \13377 , \9125 , \13020 );
and \U$6910 ( \13378 , \9127 , \13047 );
and \U$6911 ( \13379 , \9129 , \13074 );
and \U$6912 ( \13380 , \9131 , \13101 );
and \U$6913 ( \13381 , \9133 , \13128 );
and \U$6914 ( \13382 , \9135 , \13155 );
and \U$6915 ( \13383 , \9137 , \13182 );
and \U$6916 ( \13384 , \9139 , \13209 );
and \U$6917 ( \13385 , \9141 , \13236 );
and \U$6918 ( \13386 , \9143 , \13263 );
and \U$6919 ( \13387 , \9145 , \13290 );
or \U$6920 ( \13388 , \13372 , \13373 , \13374 , \13375 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 , \13382 , \13383 , \13384 , \13385 , \13386 , \13387 );
_DC g4b0f ( \13389_nG4b0f , \13388 , \13367 );
buf \U$6921 ( \13390 , \13389_nG4b0f );
xor \U$6922 ( \13391 , \13371 , \13390 );
or \U$6923 ( \13392 , \13370 , \13391 );
buf \U$6924 ( \13393 , RIb7af540_256);
and \U$6925 ( \13394 , \7217 , \12885 );
and \U$6926 ( \13395 , \7219 , \12912 );
and \U$6927 ( \13396 , \9155 , \12939 );
and \U$6928 ( \13397 , \9157 , \12966 );
and \U$6929 ( \13398 , \9159 , \12993 );
and \U$6930 ( \13399 , \9161 , \13020 );
and \U$6931 ( \13400 , \9163 , \13047 );
and \U$6932 ( \13401 , \9165 , \13074 );
and \U$6933 ( \13402 , \9167 , \13101 );
and \U$6934 ( \13403 , \9169 , \13128 );
and \U$6935 ( \13404 , \9171 , \13155 );
and \U$6936 ( \13405 , \9173 , \13182 );
and \U$6937 ( \13406 , \9175 , \13209 );
and \U$6938 ( \13407 , \9177 , \13236 );
and \U$6939 ( \13408 , \9179 , \13263 );
and \U$6940 ( \13409 , \9181 , \13290 );
or \U$6941 ( \13410 , \13394 , \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 , \13403 , \13404 , \13405 , \13406 , \13407 , \13408 , \13409 );
_DC g4b25 ( \13411_nG4b25 , \13410 , \13367 );
buf \U$6942 ( \13412 , \13411_nG4b25 );
xor \U$6943 ( \13413 , \13393 , \13412 );
or \U$6944 ( \13414 , \13392 , \13413 );
buf \U$6945 ( \13415 , RIb7af4c8_257);
and \U$6946 ( \13416 , \7227 , \12885 );
and \U$6947 ( \13417 , \7229 , \12912 );
and \U$6948 ( \13418 , \9191 , \12939 );
and \U$6949 ( \13419 , \9193 , \12966 );
and \U$6950 ( \13420 , \9195 , \12993 );
and \U$6951 ( \13421 , \9197 , \13020 );
and \U$6952 ( \13422 , \9199 , \13047 );
and \U$6953 ( \13423 , \9201 , \13074 );
and \U$6954 ( \13424 , \9203 , \13101 );
and \U$6955 ( \13425 , \9205 , \13128 );
and \U$6956 ( \13426 , \9207 , \13155 );
and \U$6957 ( \13427 , \9209 , \13182 );
and \U$6958 ( \13428 , \9211 , \13209 );
and \U$6959 ( \13429 , \9213 , \13236 );
and \U$6960 ( \13430 , \9215 , \13263 );
and \U$6961 ( \13431 , \9217 , \13290 );
or \U$6962 ( \13432 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 );
_DC g4b3b ( \13433_nG4b3b , \13432 , \13367 );
buf \U$6963 ( \13434 , \13433_nG4b3b );
xor \U$6964 ( \13435 , \13415 , \13434 );
or \U$6965 ( \13436 , \13414 , \13435 );
buf \U$6966 ( \13437 , RIb7af450_258);
and \U$6967 ( \13438 , \7237 , \12885 );
and \U$6968 ( \13439 , \7239 , \12912 );
and \U$6969 ( \13440 , \9227 , \12939 );
and \U$6970 ( \13441 , \9229 , \12966 );
and \U$6971 ( \13442 , \9231 , \12993 );
and \U$6972 ( \13443 , \9233 , \13020 );
and \U$6973 ( \13444 , \9235 , \13047 );
and \U$6974 ( \13445 , \9237 , \13074 );
and \U$6975 ( \13446 , \9239 , \13101 );
and \U$6976 ( \13447 , \9241 , \13128 );
and \U$6977 ( \13448 , \9243 , \13155 );
and \U$6978 ( \13449 , \9245 , \13182 );
and \U$6979 ( \13450 , \9247 , \13209 );
and \U$6980 ( \13451 , \9249 , \13236 );
and \U$6981 ( \13452 , \9251 , \13263 );
and \U$6982 ( \13453 , \9253 , \13290 );
or \U$6983 ( \13454 , \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 , \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 , \13452 , \13453 );
_DC g4b51 ( \13455_nG4b51 , \13454 , \13367 );
buf \U$6984 ( \13456 , \13455_nG4b51 );
xor \U$6985 ( \13457 , \13437 , \13456 );
or \U$6986 ( \13458 , \13436 , \13457 );
buf \U$6987 ( \13459 , RIb7af3d8_259);
and \U$6988 ( \13460 , \7247 , \12885 );
and \U$6989 ( \13461 , \7249 , \12912 );
and \U$6990 ( \13462 , \9263 , \12939 );
and \U$6991 ( \13463 , \9265 , \12966 );
and \U$6992 ( \13464 , \9267 , \12993 );
and \U$6993 ( \13465 , \9269 , \13020 );
and \U$6994 ( \13466 , \9271 , \13047 );
and \U$6995 ( \13467 , \9273 , \13074 );
and \U$6996 ( \13468 , \9275 , \13101 );
and \U$6997 ( \13469 , \9277 , \13128 );
and \U$6998 ( \13470 , \9279 , \13155 );
and \U$6999 ( \13471 , \9281 , \13182 );
and \U$7000 ( \13472 , \9283 , \13209 );
and \U$7001 ( \13473 , \9285 , \13236 );
and \U$7002 ( \13474 , \9287 , \13263 );
and \U$7003 ( \13475 , \9289 , \13290 );
or \U$7004 ( \13476 , \13460 , \13461 , \13462 , \13463 , \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 , \13473 , \13474 , \13475 );
_DC g4b67 ( \13477_nG4b67 , \13476 , \13367 );
buf \U$7005 ( \13478 , \13477_nG4b67 );
xor \U$7006 ( \13479 , \13459 , \13478 );
or \U$7007 ( \13480 , \13458 , \13479 );
buf \U$7008 ( \13481 , RIb7a5bf8_260);
and \U$7009 ( \13482 , \7257 , \12885 );
and \U$7010 ( \13483 , \7259 , \12912 );
and \U$7011 ( \13484 , \9299 , \12939 );
and \U$7012 ( \13485 , \9301 , \12966 );
and \U$7013 ( \13486 , \9303 , \12993 );
and \U$7014 ( \13487 , \9305 , \13020 );
and \U$7015 ( \13488 , \9307 , \13047 );
and \U$7016 ( \13489 , \9309 , \13074 );
and \U$7017 ( \13490 , \9311 , \13101 );
and \U$7018 ( \13491 , \9313 , \13128 );
and \U$7019 ( \13492 , \9315 , \13155 );
and \U$7020 ( \13493 , \9317 , \13182 );
and \U$7021 ( \13494 , \9319 , \13209 );
and \U$7022 ( \13495 , \9321 , \13236 );
and \U$7023 ( \13496 , \9323 , \13263 );
and \U$7024 ( \13497 , \9325 , \13290 );
or \U$7025 ( \13498 , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 , \13495 , \13496 , \13497 );
_DC g4b7d ( \13499_nG4b7d , \13498 , \13367 );
buf \U$7026 ( \13500 , \13499_nG4b7d );
xor \U$7027 ( \13501 , \13481 , \13500 );
or \U$7028 ( \13502 , \13480 , \13501 );
buf \U$7029 ( \13503 , RIb7a0c48_261);
and \U$7030 ( \13504 , \7267 , \12885 );
and \U$7031 ( \13505 , \7269 , \12912 );
and \U$7032 ( \13506 , \9335 , \12939 );
and \U$7033 ( \13507 , \9337 , \12966 );
and \U$7034 ( \13508 , \9339 , \12993 );
and \U$7035 ( \13509 , \9341 , \13020 );
and \U$7036 ( \13510 , \9343 , \13047 );
and \U$7037 ( \13511 , \9345 , \13074 );
and \U$7038 ( \13512 , \9347 , \13101 );
and \U$7039 ( \13513 , \9349 , \13128 );
and \U$7040 ( \13514 , \9351 , \13155 );
and \U$7041 ( \13515 , \9353 , \13182 );
and \U$7042 ( \13516 , \9355 , \13209 );
and \U$7043 ( \13517 , \9357 , \13236 );
and \U$7044 ( \13518 , \9359 , \13263 );
and \U$7045 ( \13519 , \9361 , \13290 );
or \U$7046 ( \13520 , \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 );
_DC g4b93 ( \13521_nG4b93 , \13520 , \13367 );
buf \U$7047 ( \13522 , \13521_nG4b93 );
xor \U$7048 ( \13523 , \13503 , \13522 );
or \U$7049 ( \13524 , \13502 , \13523 );
not \U$7050 ( \13525 , \13524 );
buf \U$7051 ( \13526 , \13525 );
and \U$7052 ( \13527 , \12858 , \13526 );
_HMUX g4b9a ( \13528_nG4b9a , \11450_nG4374 , \11662 , \13527 );
buf \U$7053 ( \13529 , \11471 );
buf \U$7054 ( \13530 , \11468 );
buf \U$7055 ( \13531 , \11453 );
buf \U$7056 ( \13532 , \11456 );
buf \U$7057 ( \13533 , \11460 );
buf \U$7058 ( \13534 , \11464 );
or \U$7059 ( \13535 , \13531 , \13532 , \13533 , \13534 );
and \U$7060 ( \13536 , \13530 , \13535 );
or \U$7061 ( \13537 , \13529 , \13536 );
buf \U$7062 ( \13538 , \13537 );
_HMUX g4ba5 ( \13539_nG4ba5 , \11661_nG4447 , \13528_nG4b9a , \13538 );
buf \U$7063 ( \13540 , RIe5319e0_6884);
buf \U$7065 ( \13541 , \13540 );
buf \U$7066 ( \13542 , RIe549ef0_6842);
buf \U$7068 ( \13543 , \13542 );
buf \U$7069 ( \13544 , RIe549770_6843);
not \U$7070 ( \13545 , \13544 );
buf \U$7071 ( \13546 , \13545 );
buf \U$7072 ( \13547 , RIe548ff0_6844);
xnor \U$7073 ( \13548 , \13547 , \13544 );
buf \U$7074 ( \13549 , \13548 );
buf \U$7075 ( \13550 , RIea91330_6888);
or \U$7076 ( \13551 , \13547 , \13544 );
xor \U$7077 ( \13552 , \13550 , \13551 );
buf \U$7078 ( \13553 , \13552 );
not \U$7079 ( \13554 , \13553 );
and \U$7080 ( \13555 , \13550 , \13551 );
buf \U$7081 ( \13556 , \13555 );
nor \U$7082 ( \13557 , \13541 , \13543 , \13546 , \13549 , \13554 , \13556 );
and \U$7083 ( \13558 , RIe5329d0_6883, \13557 );
not \U$7084 ( \13559 , \13556 );
and \U$7085 ( \13560 , \13541 , \13543 , \13546 , \13549 , \13554 , \13559 );
and \U$7086 ( \13561 , RIeb72150_6905, \13560 );
not \U$7087 ( \13562 , \13541 );
and \U$7088 ( \13563 , \13562 , \13543 , \13546 , \13549 , \13554 , \13559 );
and \U$7089 ( \13564 , RIeab80c0_6897, \13563 );
not \U$7090 ( \13565 , \13543 );
and \U$7091 ( \13566 , \13541 , \13565 , \13546 , \13549 , \13554 , \13559 );
and \U$7092 ( \13567 , RIe5331c8_6882, \13566 );
and \U$7093 ( \13568 , \13562 , \13565 , \13546 , \13549 , \13554 , \13559 );
and \U$7094 ( \13569 , RIe5339c0_6881, \13568 );
or \U$7106 ( \13570 , \13558 , \13561 , \13564 , \13567 , \13569 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
buf \U$7108 ( \13571 , \13556 );
buf \U$7109 ( \13572 , \13553 );
buf \U$7110 ( \13573 , \13541 );
buf \U$7111 ( \13574 , \13543 );
buf \U$7112 ( \13575 , \13546 );
buf \U$7113 ( \13576 , \13549 );
or \U$7114 ( \13577 , \13573 , \13574 , \13575 , \13576 );
and \U$7115 ( \13578 , \13572 , \13577 );
or \U$7116 ( \13579 , \13571 , \13578 );
buf \U$7117 ( \13580 , \13579 );
or \U$7118 ( \13581 , 1'b0 , \13580 );
_DC g4bd2 ( \13582_nG4bd2 , \13570 , \13581 );
not \U$7119 ( \13583 , \13582_nG4bd2 );
buf \U$7120 ( \13584 , RIb7b9608_246);
and \U$7121 ( \13585 , \7117 , \13557 );
and \U$7122 ( \13586 , \7119 , \13560 );
and \U$7123 ( \13587 , \7864 , \13563 );
and \U$7124 ( \13588 , \7892 , \13566 );
and \U$7125 ( \13589 , \7920 , \13568 );
or \U$7137 ( \13590 , \13585 , \13586 , \13587 , \13588 , \13589 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4bdb ( \13591_nG4bdb , \13590 , \13581 );
buf \U$7138 ( \13592 , \13591_nG4bdb );
xor \U$7139 ( \13593 , \13584 , \13592 );
buf \U$7140 ( \13594 , RIb7b9590_247);
and \U$7141 ( \13595 , \7126 , \13557 );
and \U$7142 ( \13596 , \7128 , \13560 );
and \U$7143 ( \13597 , \8338 , \13563 );
and \U$7144 ( \13598 , \8340 , \13566 );
and \U$7145 ( \13599 , \8342 , \13568 );
or \U$7157 ( \13600 , \13595 , \13596 , \13597 , \13598 , \13599 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4be5 ( \13601_nG4be5 , \13600 , \13581 );
buf \U$7158 ( \13602 , \13601_nG4be5 );
xor \U$7159 ( \13603 , \13594 , \13602 );
or \U$7160 ( \13604 , \13593 , \13603 );
buf \U$7161 ( \13605 , RIb7b9518_248);
and \U$7162 ( \13606 , \7136 , \13557 );
and \U$7163 ( \13607 , \7138 , \13560 );
and \U$7164 ( \13608 , \8374 , \13563 );
and \U$7165 ( \13609 , \8376 , \13566 );
and \U$7166 ( \13610 , \8378 , \13568 );
or \U$7178 ( \13611 , \13606 , \13607 , \13608 , \13609 , \13610 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4bf0 ( \13612_nG4bf0 , \13611 , \13581 );
buf \U$7179 ( \13613 , \13612_nG4bf0 );
xor \U$7180 ( \13614 , \13605 , \13613 );
or \U$7181 ( \13615 , \13604 , \13614 );
buf \U$7182 ( \13616 , RIb7b94a0_249);
and \U$7183 ( \13617 , \7146 , \13557 );
and \U$7184 ( \13618 , \7148 , \13560 );
and \U$7185 ( \13619 , \8410 , \13563 );
and \U$7186 ( \13620 , \8412 , \13566 );
and \U$7187 ( \13621 , \8414 , \13568 );
or \U$7199 ( \13622 , \13617 , \13618 , \13619 , \13620 , \13621 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4bfb ( \13623_nG4bfb , \13622 , \13581 );
buf \U$7200 ( \13624 , \13623_nG4bfb );
xor \U$7201 ( \13625 , \13616 , \13624 );
or \U$7202 ( \13626 , \13615 , \13625 );
buf \U$7203 ( \13627 , RIb7b9428_250);
and \U$7204 ( \13628 , \7156 , \13557 );
and \U$7205 ( \13629 , \7158 , \13560 );
and \U$7206 ( \13630 , \8446 , \13563 );
and \U$7207 ( \13631 , \8448 , \13566 );
and \U$7208 ( \13632 , \8450 , \13568 );
or \U$7220 ( \13633 , \13628 , \13629 , \13630 , \13631 , \13632 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4c06 ( \13634_nG4c06 , \13633 , \13581 );
buf \U$7221 ( \13635 , \13634_nG4c06 );
xor \U$7222 ( \13636 , \13627 , \13635 );
or \U$7223 ( \13637 , \13626 , \13636 );
buf \U$7224 ( \13638 , RIb7b93b0_251);
and \U$7225 ( \13639 , \7166 , \13557 );
and \U$7226 ( \13640 , \7168 , \13560 );
and \U$7227 ( \13641 , \8482 , \13563 );
and \U$7228 ( \13642 , \8484 , \13566 );
and \U$7229 ( \13643 , \8486 , \13568 );
or \U$7241 ( \13644 , \13639 , \13640 , \13641 , \13642 , \13643 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4c11 ( \13645_nG4c11 , \13644 , \13581 );
buf \U$7242 ( \13646 , \13645_nG4c11 );
xor \U$7243 ( \13647 , \13638 , \13646 );
or \U$7244 ( \13648 , \13637 , \13647 );
buf \U$7245 ( \13649 , RIb7af720_252);
and \U$7246 ( \13650 , \7176 , \13557 );
and \U$7247 ( \13651 , \7178 , \13560 );
and \U$7248 ( \13652 , \8518 , \13563 );
and \U$7249 ( \13653 , \8520 , \13566 );
and \U$7250 ( \13654 , \8522 , \13568 );
or \U$7262 ( \13655 , \13650 , \13651 , \13652 , \13653 , \13654 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4c1c ( \13656_nG4c1c , \13655 , \13581 );
buf \U$7263 ( \13657 , \13656_nG4c1c );
xor \U$7264 ( \13658 , \13649 , \13657 );
or \U$7265 ( \13659 , \13648 , \13658 );
buf \U$7266 ( \13660 , RIb7af6a8_253);
and \U$7267 ( \13661 , \7186 , \13557 );
and \U$7268 ( \13662 , \7188 , \13560 );
and \U$7269 ( \13663 , \8554 , \13563 );
and \U$7270 ( \13664 , \8556 , \13566 );
and \U$7271 ( \13665 , \8558 , \13568 );
or \U$7283 ( \13666 , \13661 , \13662 , \13663 , \13664 , \13665 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4c27 ( \13667_nG4c27 , \13666 , \13581 );
buf \U$7284 ( \13668 , \13667_nG4c27 );
xor \U$7285 ( \13669 , \13660 , \13668 );
or \U$7286 ( \13670 , \13659 , \13669 );
not \U$7287 ( \13671 , \13670 );
buf \U$7288 ( \13672 , \13671 );
buf \U$7289 ( \13673 , RIb7af630_254);
and \U$7290 ( \13674 , \7198 , \13557 );
and \U$7291 ( \13675 , \7200 , \13560 );
and \U$7292 ( \13676 , \8645 , \13563 );
and \U$7293 ( \13677 , \8673 , \13566 );
and \U$7294 ( \13678 , \8701 , \13568 );
or \U$7306 ( \13679 , \13674 , \13675 , \13676 , \13677 , \13678 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4c34 ( \13680_nG4c34 , \13679 , \13581 );
buf \U$7307 ( \13681 , \13680_nG4c34 );
xor \U$7308 ( \13682 , \13673 , \13681 );
buf \U$7309 ( \13683 , RIb7af5b8_255);
and \U$7310 ( \13684 , \7207 , \13557 );
and \U$7311 ( \13685 , \7209 , \13560 );
and \U$7312 ( \13686 , \9119 , \13563 );
and \U$7313 ( \13687 , \9121 , \13566 );
and \U$7314 ( \13688 , \9123 , \13568 );
or \U$7326 ( \13689 , \13684 , \13685 , \13686 , \13687 , \13688 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4c3e ( \13690_nG4c3e , \13689 , \13581 );
buf \U$7327 ( \13691 , \13690_nG4c3e );
xor \U$7328 ( \13692 , \13683 , \13691 );
or \U$7329 ( \13693 , \13682 , \13692 );
buf \U$7330 ( \13694 , RIb7af540_256);
and \U$7331 ( \13695 , \7217 , \13557 );
and \U$7332 ( \13696 , \7219 , \13560 );
and \U$7333 ( \13697 , \9155 , \13563 );
and \U$7334 ( \13698 , \9157 , \13566 );
and \U$7335 ( \13699 , \9159 , \13568 );
or \U$7347 ( \13700 , \13695 , \13696 , \13697 , \13698 , \13699 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4c49 ( \13701_nG4c49 , \13700 , \13581 );
buf \U$7348 ( \13702 , \13701_nG4c49 );
xor \U$7349 ( \13703 , \13694 , \13702 );
or \U$7350 ( \13704 , \13693 , \13703 );
buf \U$7351 ( \13705 , RIb7af4c8_257);
and \U$7352 ( \13706 , \7227 , \13557 );
and \U$7353 ( \13707 , \7229 , \13560 );
and \U$7354 ( \13708 , \9191 , \13563 );
and \U$7355 ( \13709 , \9193 , \13566 );
and \U$7356 ( \13710 , \9195 , \13568 );
or \U$7368 ( \13711 , \13706 , \13707 , \13708 , \13709 , \13710 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4c54 ( \13712_nG4c54 , \13711 , \13581 );
buf \U$7369 ( \13713 , \13712_nG4c54 );
xor \U$7370 ( \13714 , \13705 , \13713 );
or \U$7371 ( \13715 , \13704 , \13714 );
buf \U$7372 ( \13716 , RIb7af450_258);
and \U$7373 ( \13717 , \7237 , \13557 );
and \U$7374 ( \13718 , \7239 , \13560 );
and \U$7375 ( \13719 , \9227 , \13563 );
and \U$7376 ( \13720 , \9229 , \13566 );
and \U$7377 ( \13721 , \9231 , \13568 );
or \U$7389 ( \13722 , \13717 , \13718 , \13719 , \13720 , \13721 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4c5f ( \13723_nG4c5f , \13722 , \13581 );
buf \U$7390 ( \13724 , \13723_nG4c5f );
xor \U$7391 ( \13725 , \13716 , \13724 );
or \U$7392 ( \13726 , \13715 , \13725 );
buf \U$7393 ( \13727 , RIb7af3d8_259);
and \U$7394 ( \13728 , \7247 , \13557 );
and \U$7395 ( \13729 , \7249 , \13560 );
and \U$7396 ( \13730 , \9263 , \13563 );
and \U$7397 ( \13731 , \9265 , \13566 );
and \U$7398 ( \13732 , \9267 , \13568 );
or \U$7410 ( \13733 , \13728 , \13729 , \13730 , \13731 , \13732 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4c6a ( \13734_nG4c6a , \13733 , \13581 );
buf \U$7411 ( \13735 , \13734_nG4c6a );
xor \U$7412 ( \13736 , \13727 , \13735 );
or \U$7413 ( \13737 , \13726 , \13736 );
buf \U$7414 ( \13738 , RIb7a5bf8_260);
and \U$7415 ( \13739 , \7257 , \13557 );
and \U$7416 ( \13740 , \7259 , \13560 );
and \U$7417 ( \13741 , \9299 , \13563 );
and \U$7418 ( \13742 , \9301 , \13566 );
and \U$7419 ( \13743 , \9303 , \13568 );
or \U$7431 ( \13744 , \13739 , \13740 , \13741 , \13742 , \13743 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4c75 ( \13745_nG4c75 , \13744 , \13581 );
buf \U$7432 ( \13746 , \13745_nG4c75 );
xor \U$7433 ( \13747 , \13738 , \13746 );
or \U$7434 ( \13748 , \13737 , \13747 );
buf \U$7435 ( \13749 , RIb7a0c48_261);
and \U$7436 ( \13750 , \7267 , \13557 );
and \U$7437 ( \13751 , \7269 , \13560 );
and \U$7438 ( \13752 , \9335 , \13563 );
and \U$7439 ( \13753 , \9337 , \13566 );
and \U$7440 ( \13754 , \9339 , \13568 );
or \U$7452 ( \13755 , \13750 , \13751 , \13752 , \13753 , \13754 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g4c80 ( \13756_nG4c80 , \13755 , \13581 );
buf \U$7453 ( \13757 , \13756_nG4c80 );
xor \U$7454 ( \13758 , \13749 , \13757 );
or \U$7455 ( \13759 , \13748 , \13758 );
not \U$7456 ( \13760 , \13759 );
buf \U$7457 ( \13761 , \13760 );
and \U$7458 ( \13762 , \13672 , \13761 );
and \U$7459 ( \13763 , \13583 , \13762 );
_HMUX g4c88 ( \13764_nG4c88 , \13539_nG4ba5 , \13541 , \13763 );
buf \U$7462 ( \13765 , \13541 );
buf \U$7465 ( \13766 , \13543 );
buf \U$7468 ( \13767 , \13546 );
buf \U$7471 ( \13768 , \13549 );
buf \U$7472 ( \13769 , \13553 );
not \U$7473 ( \13770 , \13769 );
buf \U$7474 ( \13771 , \13770 );
not \U$7475 ( \13772 , \13771 );
buf \U$7476 ( \13773 , \13556 );
xnor \U$7477 ( \13774 , \13773 , \13769 );
buf \U$7478 ( \13775 , \13774 );
or \U$7479 ( \13776 , \13773 , \13769 );
not \U$7480 ( \13777 , \13776 );
buf \U$7481 ( \13778 , \13777 );
buf \U$7482 ( \13779 , \13778 );
buf \U$7483 ( \13780 , \13778 );
buf \U$7484 ( \13781 , \13778 );
buf \U$7485 ( \13782 , \13778 );
buf \U$7486 ( \13783 , \13778 );
buf \U$7487 ( \13784 , \13778 );
buf \U$7488 ( \13785 , \13778 );
buf \U$7489 ( \13786 , \13778 );
buf \U$7490 ( \13787 , \13778 );
buf \U$7491 ( \13788 , \13778 );
buf \U$7492 ( \13789 , \13778 );
buf \U$7493 ( \13790 , \13778 );
buf \U$7494 ( \13791 , \13778 );
buf \U$7495 ( \13792 , \13778 );
buf \U$7496 ( \13793 , \13778 );
buf \U$7497 ( \13794 , \13778 );
buf \U$7498 ( \13795 , \13778 );
buf \U$7499 ( \13796 , \13778 );
buf \U$7500 ( \13797 , \13778 );
buf \U$7501 ( \13798 , \13778 );
buf \U$7502 ( \13799 , \13778 );
buf \U$7503 ( \13800 , \13778 );
buf \U$7504 ( \13801 , \13778 );
buf \U$7505 ( \13802 , \13778 );
buf \U$7506 ( \13803 , \13778 );
nor \U$7507 ( \13804 , \13765 , \13766 , \13767 , \13768 , \13772 , \13775 , \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 , \13802 , \13803 );
and \U$7508 ( \13805 , RIe5329d0_6883, \13804 );
not \U$7509 ( \13806 , \13765 );
not \U$7510 ( \13807 , \13766 );
not \U$7511 ( \13808 , \13767 );
not \U$7512 ( \13809 , \13768 );
buf \U$7513 ( \13810 , \13778 );
buf \U$7514 ( \13811 , \13778 );
buf \U$7515 ( \13812 , \13778 );
buf \U$7516 ( \13813 , \13778 );
buf \U$7517 ( \13814 , \13778 );
buf \U$7518 ( \13815 , \13778 );
buf \U$7519 ( \13816 , \13778 );
buf \U$7520 ( \13817 , \13778 );
buf \U$7521 ( \13818 , \13778 );
buf \U$7522 ( \13819 , \13778 );
buf \U$7523 ( \13820 , \13778 );
buf \U$7524 ( \13821 , \13778 );
buf \U$7525 ( \13822 , \13778 );
buf \U$7526 ( \13823 , \13778 );
buf \U$7527 ( \13824 , \13778 );
buf \U$7528 ( \13825 , \13778 );
buf \U$7529 ( \13826 , \13778 );
buf \U$7530 ( \13827 , \13778 );
buf \U$7531 ( \13828 , \13778 );
buf \U$7532 ( \13829 , \13778 );
buf \U$7533 ( \13830 , \13778 );
buf \U$7534 ( \13831 , \13778 );
buf \U$7535 ( \13832 , \13778 );
buf \U$7536 ( \13833 , \13778 );
buf \U$7537 ( \13834 , \13778 );
nor \U$7538 ( \13835 , \13806 , \13807 , \13808 , \13809 , \13771 , \13775 , \13778 , \13810 , \13811 , \13812 , \13813 , \13814 , \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 , \13822 , \13823 , \13824 , \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 );
and \U$7539 ( \13836 , RIeb72150_6905, \13835 );
buf \U$7540 ( \13837 , \13778 );
buf \U$7541 ( \13838 , \13778 );
buf \U$7542 ( \13839 , \13778 );
buf \U$7543 ( \13840 , \13778 );
buf \U$7544 ( \13841 , \13778 );
buf \U$7545 ( \13842 , \13778 );
buf \U$7546 ( \13843 , \13778 );
buf \U$7547 ( \13844 , \13778 );
buf \U$7548 ( \13845 , \13778 );
buf \U$7549 ( \13846 , \13778 );
buf \U$7550 ( \13847 , \13778 );
buf \U$7551 ( \13848 , \13778 );
buf \U$7552 ( \13849 , \13778 );
buf \U$7553 ( \13850 , \13778 );
buf \U$7554 ( \13851 , \13778 );
buf \U$7555 ( \13852 , \13778 );
buf \U$7556 ( \13853 , \13778 );
buf \U$7557 ( \13854 , \13778 );
buf \U$7558 ( \13855 , \13778 );
buf \U$7559 ( \13856 , \13778 );
buf \U$7560 ( \13857 , \13778 );
buf \U$7561 ( \13858 , \13778 );
buf \U$7562 ( \13859 , \13778 );
buf \U$7563 ( \13860 , \13778 );
buf \U$7564 ( \13861 , \13778 );
nor \U$7565 ( \13862 , \13765 , \13807 , \13808 , \13809 , \13771 , \13775 , \13778 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 , \13852 , \13853 , \13854 , \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 );
and \U$7566 ( \13863 , RIeab80c0_6897, \13862 );
buf \U$7567 ( \13864 , \13778 );
buf \U$7568 ( \13865 , \13778 );
buf \U$7569 ( \13866 , \13778 );
buf \U$7570 ( \13867 , \13778 );
buf \U$7571 ( \13868 , \13778 );
buf \U$7572 ( \13869 , \13778 );
buf \U$7573 ( \13870 , \13778 );
buf \U$7574 ( \13871 , \13778 );
buf \U$7575 ( \13872 , \13778 );
buf \U$7576 ( \13873 , \13778 );
buf \U$7577 ( \13874 , \13778 );
buf \U$7578 ( \13875 , \13778 );
buf \U$7579 ( \13876 , \13778 );
buf \U$7580 ( \13877 , \13778 );
buf \U$7581 ( \13878 , \13778 );
buf \U$7582 ( \13879 , \13778 );
buf \U$7583 ( \13880 , \13778 );
buf \U$7584 ( \13881 , \13778 );
buf \U$7585 ( \13882 , \13778 );
buf \U$7586 ( \13883 , \13778 );
buf \U$7587 ( \13884 , \13778 );
buf \U$7588 ( \13885 , \13778 );
buf \U$7589 ( \13886 , \13778 );
buf \U$7590 ( \13887 , \13778 );
buf \U$7591 ( \13888 , \13778 );
nor \U$7592 ( \13889 , \13806 , \13766 , \13808 , \13809 , \13771 , \13775 , \13778 , \13864 , \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 , \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 , \13885 , \13886 , \13887 , \13888 );
and \U$7593 ( \13890 , RIe5331c8_6882, \13889 );
buf \U$7594 ( \13891 , \13778 );
buf \U$7595 ( \13892 , \13778 );
buf \U$7596 ( \13893 , \13778 );
buf \U$7597 ( \13894 , \13778 );
buf \U$7598 ( \13895 , \13778 );
buf \U$7599 ( \13896 , \13778 );
buf \U$7600 ( \13897 , \13778 );
buf \U$7601 ( \13898 , \13778 );
buf \U$7602 ( \13899 , \13778 );
buf \U$7603 ( \13900 , \13778 );
buf \U$7604 ( \13901 , \13778 );
buf \U$7605 ( \13902 , \13778 );
buf \U$7606 ( \13903 , \13778 );
buf \U$7607 ( \13904 , \13778 );
buf \U$7608 ( \13905 , \13778 );
buf \U$7609 ( \13906 , \13778 );
buf \U$7610 ( \13907 , \13778 );
buf \U$7611 ( \13908 , \13778 );
buf \U$7612 ( \13909 , \13778 );
buf \U$7613 ( \13910 , \13778 );
buf \U$7614 ( \13911 , \13778 );
buf \U$7615 ( \13912 , \13778 );
buf \U$7616 ( \13913 , \13778 );
buf \U$7617 ( \13914 , \13778 );
buf \U$7618 ( \13915 , \13778 );
nor \U$7619 ( \13916 , \13765 , \13766 , \13808 , \13809 , \13771 , \13775 , \13778 , \13891 , \13892 , \13893 , \13894 , \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 , \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 , \13915 );
and \U$7620 ( \13917 , RIe5339c0_6881, \13916 );
buf \U$7621 ( \13918 , \13778 );
buf \U$7622 ( \13919 , \13778 );
buf \U$7623 ( \13920 , \13778 );
buf \U$7624 ( \13921 , \13778 );
buf \U$7625 ( \13922 , \13778 );
buf \U$7626 ( \13923 , \13778 );
buf \U$7627 ( \13924 , \13778 );
buf \U$7628 ( \13925 , \13778 );
buf \U$7629 ( \13926 , \13778 );
buf \U$7630 ( \13927 , \13778 );
buf \U$7631 ( \13928 , \13778 );
buf \U$7632 ( \13929 , \13778 );
buf \U$7633 ( \13930 , \13778 );
buf \U$7634 ( \13931 , \13778 );
buf \U$7635 ( \13932 , \13778 );
buf \U$7636 ( \13933 , \13778 );
buf \U$7637 ( \13934 , \13778 );
buf \U$7638 ( \13935 , \13778 );
buf \U$7639 ( \13936 , \13778 );
buf \U$7640 ( \13937 , \13778 );
buf \U$7641 ( \13938 , \13778 );
buf \U$7642 ( \13939 , \13778 );
buf \U$7643 ( \13940 , \13778 );
buf \U$7644 ( \13941 , \13778 );
buf \U$7645 ( \13942 , \13778 );
nor \U$7646 ( \13943 , \13806 , \13807 , \13767 , \13809 , \13771 , \13775 , \13778 , \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 , \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 , \13942 );
and \U$7647 ( \13944 , RIeab87c8_6898, \13943 );
buf \U$7648 ( \13945 , \13778 );
buf \U$7649 ( \13946 , \13778 );
buf \U$7650 ( \13947 , \13778 );
buf \U$7651 ( \13948 , \13778 );
buf \U$7652 ( \13949 , \13778 );
buf \U$7653 ( \13950 , \13778 );
buf \U$7654 ( \13951 , \13778 );
buf \U$7655 ( \13952 , \13778 );
buf \U$7656 ( \13953 , \13778 );
buf \U$7657 ( \13954 , \13778 );
buf \U$7658 ( \13955 , \13778 );
buf \U$7659 ( \13956 , \13778 );
buf \U$7660 ( \13957 , \13778 );
buf \U$7661 ( \13958 , \13778 );
buf \U$7662 ( \13959 , \13778 );
buf \U$7663 ( \13960 , \13778 );
buf \U$7664 ( \13961 , \13778 );
buf \U$7665 ( \13962 , \13778 );
buf \U$7666 ( \13963 , \13778 );
buf \U$7667 ( \13964 , \13778 );
buf \U$7668 ( \13965 , \13778 );
buf \U$7669 ( \13966 , \13778 );
buf \U$7670 ( \13967 , \13778 );
buf \U$7671 ( \13968 , \13778 );
buf \U$7672 ( \13969 , \13778 );
nor \U$7673 ( \13970 , \13765 , \13807 , \13767 , \13809 , \13771 , \13775 , \13778 , \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 , \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 , \13965 , \13966 , \13967 , \13968 , \13969 );
and \U$7674 ( \13971 , RIe5341b8_6880, \13970 );
buf \U$7675 ( \13972 , \13778 );
buf \U$7676 ( \13973 , \13778 );
buf \U$7677 ( \13974 , \13778 );
buf \U$7678 ( \13975 , \13778 );
buf \U$7679 ( \13976 , \13778 );
buf \U$7680 ( \13977 , \13778 );
buf \U$7681 ( \13978 , \13778 );
buf \U$7682 ( \13979 , \13778 );
buf \U$7683 ( \13980 , \13778 );
buf \U$7684 ( \13981 , \13778 );
buf \U$7685 ( \13982 , \13778 );
buf \U$7686 ( \13983 , \13778 );
buf \U$7687 ( \13984 , \13778 );
buf \U$7688 ( \13985 , \13778 );
buf \U$7689 ( \13986 , \13778 );
buf \U$7690 ( \13987 , \13778 );
buf \U$7691 ( \13988 , \13778 );
buf \U$7692 ( \13989 , \13778 );
buf \U$7693 ( \13990 , \13778 );
buf \U$7694 ( \13991 , \13778 );
buf \U$7695 ( \13992 , \13778 );
buf \U$7696 ( \13993 , \13778 );
buf \U$7697 ( \13994 , \13778 );
buf \U$7698 ( \13995 , \13778 );
buf \U$7699 ( \13996 , \13778 );
nor \U$7700 ( \13997 , \13806 , \13766 , \13767 , \13809 , \13771 , \13775 , \13778 , \13972 , \13973 , \13974 , \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 , \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 , \13995 , \13996 );
and \U$7701 ( \13998 , RIe5349b0_6879, \13997 );
buf \U$7702 ( \13999 , \13778 );
buf \U$7703 ( \14000 , \13778 );
buf \U$7704 ( \14001 , \13778 );
buf \U$7705 ( \14002 , \13778 );
buf \U$7706 ( \14003 , \13778 );
buf \U$7707 ( \14004 , \13778 );
buf \U$7708 ( \14005 , \13778 );
buf \U$7709 ( \14006 , \13778 );
buf \U$7710 ( \14007 , \13778 );
buf \U$7711 ( \14008 , \13778 );
buf \U$7712 ( \14009 , \13778 );
buf \U$7713 ( \14010 , \13778 );
buf \U$7714 ( \14011 , \13778 );
buf \U$7715 ( \14012 , \13778 );
buf \U$7716 ( \14013 , \13778 );
buf \U$7717 ( \14014 , \13778 );
buf \U$7718 ( \14015 , \13778 );
buf \U$7719 ( \14016 , \13778 );
buf \U$7720 ( \14017 , \13778 );
buf \U$7721 ( \14018 , \13778 );
buf \U$7722 ( \14019 , \13778 );
buf \U$7723 ( \14020 , \13778 );
buf \U$7724 ( \14021 , \13778 );
buf \U$7725 ( \14022 , \13778 );
buf \U$7726 ( \14023 , \13778 );
nor \U$7727 ( \14024 , \13765 , \13766 , \13767 , \13809 , \13771 , \13775 , \13778 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 , \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 , \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 , \14022 , \14023 );
and \U$7728 ( \14025 , RIea94af8_6890, \14024 );
buf \U$7729 ( \14026 , \13778 );
buf \U$7730 ( \14027 , \13778 );
buf \U$7731 ( \14028 , \13778 );
buf \U$7732 ( \14029 , \13778 );
buf \U$7733 ( \14030 , \13778 );
buf \U$7734 ( \14031 , \13778 );
buf \U$7735 ( \14032 , \13778 );
buf \U$7736 ( \14033 , \13778 );
buf \U$7737 ( \14034 , \13778 );
buf \U$7738 ( \14035 , \13778 );
buf \U$7739 ( \14036 , \13778 );
buf \U$7740 ( \14037 , \13778 );
buf \U$7741 ( \14038 , \13778 );
buf \U$7742 ( \14039 , \13778 );
buf \U$7743 ( \14040 , \13778 );
buf \U$7744 ( \14041 , \13778 );
buf \U$7745 ( \14042 , \13778 );
buf \U$7746 ( \14043 , \13778 );
buf \U$7747 ( \14044 , \13778 );
buf \U$7748 ( \14045 , \13778 );
buf \U$7749 ( \14046 , \13778 );
buf \U$7750 ( \14047 , \13778 );
buf \U$7751 ( \14048 , \13778 );
buf \U$7752 ( \14049 , \13778 );
buf \U$7753 ( \14050 , \13778 );
nor \U$7754 ( \14051 , \13806 , \13807 , \13808 , \13768 , \13771 , \13775 , \13778 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 , \14032 , \14033 , \14034 , \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 , \14042 , \14043 , \14044 , \14045 , \14046 , \14047 , \14048 , \14049 , \14050 );
and \U$7755 ( \14052 , RIe5351a8_6878, \14051 );
buf \U$7756 ( \14053 , \13778 );
buf \U$7757 ( \14054 , \13778 );
buf \U$7758 ( \14055 , \13778 );
buf \U$7759 ( \14056 , \13778 );
buf \U$7760 ( \14057 , \13778 );
buf \U$7761 ( \14058 , \13778 );
buf \U$7762 ( \14059 , \13778 );
buf \U$7763 ( \14060 , \13778 );
buf \U$7764 ( \14061 , \13778 );
buf \U$7765 ( \14062 , \13778 );
buf \U$7766 ( \14063 , \13778 );
buf \U$7767 ( \14064 , \13778 );
buf \U$7768 ( \14065 , \13778 );
buf \U$7769 ( \14066 , \13778 );
buf \U$7770 ( \14067 , \13778 );
buf \U$7771 ( \14068 , \13778 );
buf \U$7772 ( \14069 , \13778 );
buf \U$7773 ( \14070 , \13778 );
buf \U$7774 ( \14071 , \13778 );
buf \U$7775 ( \14072 , \13778 );
buf \U$7776 ( \14073 , \13778 );
buf \U$7777 ( \14074 , \13778 );
buf \U$7778 ( \14075 , \13778 );
buf \U$7779 ( \14076 , \13778 );
buf \U$7780 ( \14077 , \13778 );
nor \U$7781 ( \14078 , \13765 , \13807 , \13808 , \13768 , \13771 , \13775 , \13778 , \14053 , \14054 , \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 , \14062 , \14063 , \14064 , \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 , \14072 , \14073 , \14074 , \14075 , \14076 , \14077 );
and \U$7782 ( \14079 , RIe5359a0_6877, \14078 );
buf \U$7783 ( \14080 , \13778 );
buf \U$7784 ( \14081 , \13778 );
buf \U$7785 ( \14082 , \13778 );
buf \U$7786 ( \14083 , \13778 );
buf \U$7787 ( \14084 , \13778 );
buf \U$7788 ( \14085 , \13778 );
buf \U$7789 ( \14086 , \13778 );
buf \U$7790 ( \14087 , \13778 );
buf \U$7791 ( \14088 , \13778 );
buf \U$7792 ( \14089 , \13778 );
buf \U$7793 ( \14090 , \13778 );
buf \U$7794 ( \14091 , \13778 );
buf \U$7795 ( \14092 , \13778 );
buf \U$7796 ( \14093 , \13778 );
buf \U$7797 ( \14094 , \13778 );
buf \U$7798 ( \14095 , \13778 );
buf \U$7799 ( \14096 , \13778 );
buf \U$7800 ( \14097 , \13778 );
buf \U$7801 ( \14098 , \13778 );
buf \U$7802 ( \14099 , \13778 );
buf \U$7803 ( \14100 , \13778 );
buf \U$7804 ( \14101 , \13778 );
buf \U$7805 ( \14102 , \13778 );
buf \U$7806 ( \14103 , \13778 );
buf \U$7807 ( \14104 , \13778 );
nor \U$7808 ( \14105 , \13806 , \13766 , \13808 , \13768 , \13771 , \13775 , \13778 , \14080 , \14081 , \14082 , \14083 , \14084 , \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 , \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 );
and \U$7809 ( \14106 , RIeab78c8_6895, \14105 );
buf \U$7810 ( \14107 , \13778 );
buf \U$7811 ( \14108 , \13778 );
buf \U$7812 ( \14109 , \13778 );
buf \U$7813 ( \14110 , \13778 );
buf \U$7814 ( \14111 , \13778 );
buf \U$7815 ( \14112 , \13778 );
buf \U$7816 ( \14113 , \13778 );
buf \U$7817 ( \14114 , \13778 );
buf \U$7818 ( \14115 , \13778 );
buf \U$7819 ( \14116 , \13778 );
buf \U$7820 ( \14117 , \13778 );
buf \U$7821 ( \14118 , \13778 );
buf \U$7822 ( \14119 , \13778 );
buf \U$7823 ( \14120 , \13778 );
buf \U$7824 ( \14121 , \13778 );
buf \U$7825 ( \14122 , \13778 );
buf \U$7826 ( \14123 , \13778 );
buf \U$7827 ( \14124 , \13778 );
buf \U$7828 ( \14125 , \13778 );
buf \U$7829 ( \14126 , \13778 );
buf \U$7830 ( \14127 , \13778 );
buf \U$7831 ( \14128 , \13778 );
buf \U$7832 ( \14129 , \13778 );
buf \U$7833 ( \14130 , \13778 );
buf \U$7834 ( \14131 , \13778 );
nor \U$7835 ( \14132 , \13765 , \13766 , \13808 , \13768 , \13771 , \13775 , \13778 , \14107 , \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 , \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 , \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 );
and \U$7836 ( \14133 , RIeab7d00_6896, \14132 );
buf \U$7837 ( \14134 , \13778 );
buf \U$7838 ( \14135 , \13778 );
buf \U$7839 ( \14136 , \13778 );
buf \U$7840 ( \14137 , \13778 );
buf \U$7841 ( \14138 , \13778 );
buf \U$7842 ( \14139 , \13778 );
buf \U$7843 ( \14140 , \13778 );
buf \U$7844 ( \14141 , \13778 );
buf \U$7845 ( \14142 , \13778 );
buf \U$7846 ( \14143 , \13778 );
buf \U$7847 ( \14144 , \13778 );
buf \U$7848 ( \14145 , \13778 );
buf \U$7849 ( \14146 , \13778 );
buf \U$7850 ( \14147 , \13778 );
buf \U$7851 ( \14148 , \13778 );
buf \U$7852 ( \14149 , \13778 );
buf \U$7853 ( \14150 , \13778 );
buf \U$7854 ( \14151 , \13778 );
buf \U$7855 ( \14152 , \13778 );
buf \U$7856 ( \14153 , \13778 );
buf \U$7857 ( \14154 , \13778 );
buf \U$7858 ( \14155 , \13778 );
buf \U$7859 ( \14156 , \13778 );
buf \U$7860 ( \14157 , \13778 );
buf \U$7861 ( \14158 , \13778 );
nor \U$7862 ( \14159 , \13806 , \13807 , \13767 , \13768 , \13771 , \13775 , \13778 , \14134 , \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 , \14142 , \14143 , \14144 , \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 , \14155 , \14156 , \14157 , \14158 );
and \U$7863 ( \14160 , RIeacfa18_6902, \14159 );
buf \U$7864 ( \14161 , \13778 );
buf \U$7865 ( \14162 , \13778 );
buf \U$7866 ( \14163 , \13778 );
buf \U$7867 ( \14164 , \13778 );
buf \U$7868 ( \14165 , \13778 );
buf \U$7869 ( \14166 , \13778 );
buf \U$7870 ( \14167 , \13778 );
buf \U$7871 ( \14168 , \13778 );
buf \U$7872 ( \14169 , \13778 );
buf \U$7873 ( \14170 , \13778 );
buf \U$7874 ( \14171 , \13778 );
buf \U$7875 ( \14172 , \13778 );
buf \U$7876 ( \14173 , \13778 );
buf \U$7877 ( \14174 , \13778 );
buf \U$7878 ( \14175 , \13778 );
buf \U$7879 ( \14176 , \13778 );
buf \U$7880 ( \14177 , \13778 );
buf \U$7881 ( \14178 , \13778 );
buf \U$7882 ( \14179 , \13778 );
buf \U$7883 ( \14180 , \13778 );
buf \U$7884 ( \14181 , \13778 );
buf \U$7885 ( \14182 , \13778 );
buf \U$7886 ( \14183 , \13778 );
buf \U$7887 ( \14184 , \13778 );
buf \U$7888 ( \14185 , \13778 );
nor \U$7889 ( \14186 , \13765 , \13807 , \13767 , \13768 , \13771 , \13775 , \13778 , \14161 , \14162 , \14163 , \14164 , \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 , \14172 , \14173 , \14174 , \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 , \14185 );
and \U$7890 ( \14187 , RIeab6518_6891, \14186 );
buf \U$7891 ( \14188 , \13778 );
buf \U$7892 ( \14189 , \13778 );
buf \U$7893 ( \14190 , \13778 );
buf \U$7894 ( \14191 , \13778 );
buf \U$7895 ( \14192 , \13778 );
buf \U$7896 ( \14193 , \13778 );
buf \U$7897 ( \14194 , \13778 );
buf \U$7898 ( \14195 , \13778 );
buf \U$7899 ( \14196 , \13778 );
buf \U$7900 ( \14197 , \13778 );
buf \U$7901 ( \14198 , \13778 );
buf \U$7902 ( \14199 , \13778 );
buf \U$7903 ( \14200 , \13778 );
buf \U$7904 ( \14201 , \13778 );
buf \U$7905 ( \14202 , \13778 );
buf \U$7906 ( \14203 , \13778 );
buf \U$7907 ( \14204 , \13778 );
buf \U$7908 ( \14205 , \13778 );
buf \U$7909 ( \14206 , \13778 );
buf \U$7910 ( \14207 , \13778 );
buf \U$7911 ( \14208 , \13778 );
buf \U$7912 ( \14209 , \13778 );
buf \U$7913 ( \14210 , \13778 );
buf \U$7914 ( \14211 , \13778 );
buf \U$7915 ( \14212 , \13778 );
nor \U$7916 ( \14213 , \13806 , \13766 , \13767 , \13768 , \13771 , \13775 , \13778 , \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 , \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 , \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 , \14212 );
and \U$7917 ( \14214 , RIeb352c8_6904, \14213 );
or \U$7918 ( \14215 , \13805 , \13836 , \13863 , \13890 , \13917 , \13944 , \13971 , \13998 , \14025 , \14052 , \14079 , \14106 , \14133 , \14160 , \14187 , \14214 );
buf \U$7919 ( \14216 , \13778 );
not \U$7920 ( \14217 , \14216 );
buf \U$7921 ( \14218 , \13766 );
buf \U$7922 ( \14219 , \13767 );
buf \U$7923 ( \14220 , \13768 );
buf \U$7924 ( \14221 , \13771 );
buf \U$7925 ( \14222 , \13775 );
buf \U$7926 ( \14223 , \13778 );
buf \U$7927 ( \14224 , \13778 );
buf \U$7928 ( \14225 , \13778 );
buf \U$7929 ( \14226 , \13778 );
buf \U$7930 ( \14227 , \13778 );
buf \U$7931 ( \14228 , \13778 );
buf \U$7932 ( \14229 , \13778 );
buf \U$7933 ( \14230 , \13778 );
buf \U$7934 ( \14231 , \13778 );
buf \U$7935 ( \14232 , \13778 );
buf \U$7936 ( \14233 , \13778 );
buf \U$7937 ( \14234 , \13778 );
buf \U$7938 ( \14235 , \13778 );
buf \U$7939 ( \14236 , \13778 );
buf \U$7940 ( \14237 , \13778 );
buf \U$7941 ( \14238 , \13778 );
buf \U$7942 ( \14239 , \13778 );
buf \U$7943 ( \14240 , \13778 );
buf \U$7944 ( \14241 , \13778 );
buf \U$7945 ( \14242 , \13778 );
buf \U$7946 ( \14243 , \13778 );
buf \U$7947 ( \14244 , \13778 );
buf \U$7948 ( \14245 , \13778 );
buf \U$7949 ( \14246 , \13778 );
buf \U$7950 ( \14247 , \13778 );
buf \U$7951 ( \14248 , \13765 );
or \U$7952 ( \14249 , \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 , \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 , \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 , \14245 , \14246 , \14247 , \14248 );
nand \U$7953 ( \14250 , \14217 , \14249 );
buf \U$7954 ( \14251 , \14250 );
buf \U$7955 ( \14252 , \13778 );
not \U$7956 ( \14253 , \14252 );
buf \U$7957 ( \14254 , \13775 );
buf \U$7958 ( \14255 , \13778 );
buf \U$7959 ( \14256 , \13778 );
buf \U$7960 ( \14257 , \13778 );
buf \U$7961 ( \14258 , \13778 );
buf \U$7962 ( \14259 , \13778 );
buf \U$7963 ( \14260 , \13778 );
buf \U$7964 ( \14261 , \13778 );
buf \U$7965 ( \14262 , \13778 );
buf \U$7966 ( \14263 , \13778 );
buf \U$7967 ( \14264 , \13778 );
buf \U$7968 ( \14265 , \13778 );
buf \U$7969 ( \14266 , \13778 );
buf \U$7970 ( \14267 , \13778 );
buf \U$7971 ( \14268 , \13778 );
buf \U$7972 ( \14269 , \13778 );
buf \U$7973 ( \14270 , \13778 );
buf \U$7974 ( \14271 , \13778 );
buf \U$7975 ( \14272 , \13778 );
buf \U$7976 ( \14273 , \13778 );
buf \U$7977 ( \14274 , \13778 );
buf \U$7978 ( \14275 , \13778 );
buf \U$7979 ( \14276 , \13778 );
buf \U$7980 ( \14277 , \13778 );
buf \U$7981 ( \14278 , \13778 );
buf \U$7982 ( \14279 , \13778 );
buf \U$7983 ( \14280 , \13771 );
buf \U$7984 ( \14281 , \13765 );
buf \U$7985 ( \14282 , \13766 );
buf \U$7986 ( \14283 , \13767 );
buf \U$7987 ( \14284 , \13768 );
or \U$7988 ( \14285 , \14281 , \14282 , \14283 , \14284 );
and \U$7989 ( \14286 , \14280 , \14285 );
or \U$7990 ( \14287 , \14254 , \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 , \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 , \14275 , \14276 , \14277 , \14278 , \14279 , \14286 );
and \U$7991 ( \14288 , \14253 , \14287 );
buf \U$7992 ( \14289 , \14288 );
or \U$7993 ( \14290 , \14251 , \14289 );
_DC g4e9f ( \14291_nG4e9f , \14215 , \14290 );
not \U$7994 ( \14292 , \14291_nG4e9f );
buf \U$7995 ( \14293 , RIb7b9608_246);
buf \U$7996 ( \14294 , \13778 );
buf \U$7997 ( \14295 , \13778 );
buf \U$7998 ( \14296 , \13778 );
buf \U$7999 ( \14297 , \13778 );
buf \U$8000 ( \14298 , \13778 );
buf \U$8001 ( \14299 , \13778 );
buf \U$8002 ( \14300 , \13778 );
buf \U$8003 ( \14301 , \13778 );
buf \U$8004 ( \14302 , \13778 );
buf \U$8005 ( \14303 , \13778 );
buf \U$8006 ( \14304 , \13778 );
buf \U$8007 ( \14305 , \13778 );
buf \U$8008 ( \14306 , \13778 );
buf \U$8009 ( \14307 , \13778 );
buf \U$8010 ( \14308 , \13778 );
buf \U$8011 ( \14309 , \13778 );
buf \U$8012 ( \14310 , \13778 );
buf \U$8013 ( \14311 , \13778 );
buf \U$8014 ( \14312 , \13778 );
buf \U$8015 ( \14313 , \13778 );
buf \U$8016 ( \14314 , \13778 );
buf \U$8017 ( \14315 , \13778 );
buf \U$8018 ( \14316 , \13778 );
buf \U$8019 ( \14317 , \13778 );
buf \U$8020 ( \14318 , \13778 );
nor \U$8021 ( \14319 , \13765 , \13766 , \13767 , \13768 , \13772 , \13775 , \13778 , \14294 , \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 , \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 , \14315 , \14316 , \14317 , \14318 );
and \U$8022 ( \14320 , \7117 , \14319 );
buf \U$8023 ( \14321 , \13778 );
buf \U$8024 ( \14322 , \13778 );
buf \U$8025 ( \14323 , \13778 );
buf \U$8026 ( \14324 , \13778 );
buf \U$8027 ( \14325 , \13778 );
buf \U$8028 ( \14326 , \13778 );
buf \U$8029 ( \14327 , \13778 );
buf \U$8030 ( \14328 , \13778 );
buf \U$8031 ( \14329 , \13778 );
buf \U$8032 ( \14330 , \13778 );
buf \U$8033 ( \14331 , \13778 );
buf \U$8034 ( \14332 , \13778 );
buf \U$8035 ( \14333 , \13778 );
buf \U$8036 ( \14334 , \13778 );
buf \U$8037 ( \14335 , \13778 );
buf \U$8038 ( \14336 , \13778 );
buf \U$8039 ( \14337 , \13778 );
buf \U$8040 ( \14338 , \13778 );
buf \U$8041 ( \14339 , \13778 );
buf \U$8042 ( \14340 , \13778 );
buf \U$8043 ( \14341 , \13778 );
buf \U$8044 ( \14342 , \13778 );
buf \U$8045 ( \14343 , \13778 );
buf \U$8046 ( \14344 , \13778 );
buf \U$8047 ( \14345 , \13778 );
nor \U$8048 ( \14346 , \13806 , \13807 , \13808 , \13809 , \13771 , \13775 , \13778 , \14321 , \14322 , \14323 , \14324 , \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 , \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 , \14342 , \14343 , \14344 , \14345 );
and \U$8049 ( \14347 , \7119 , \14346 );
buf \U$8050 ( \14348 , \13778 );
buf \U$8051 ( \14349 , \13778 );
buf \U$8052 ( \14350 , \13778 );
buf \U$8053 ( \14351 , \13778 );
buf \U$8054 ( \14352 , \13778 );
buf \U$8055 ( \14353 , \13778 );
buf \U$8056 ( \14354 , \13778 );
buf \U$8057 ( \14355 , \13778 );
buf \U$8058 ( \14356 , \13778 );
buf \U$8059 ( \14357 , \13778 );
buf \U$8060 ( \14358 , \13778 );
buf \U$8061 ( \14359 , \13778 );
buf \U$8062 ( \14360 , \13778 );
buf \U$8063 ( \14361 , \13778 );
buf \U$8064 ( \14362 , \13778 );
buf \U$8065 ( \14363 , \13778 );
buf \U$8066 ( \14364 , \13778 );
buf \U$8067 ( \14365 , \13778 );
buf \U$8068 ( \14366 , \13778 );
buf \U$8069 ( \14367 , \13778 );
buf \U$8070 ( \14368 , \13778 );
buf \U$8071 ( \14369 , \13778 );
buf \U$8072 ( \14370 , \13778 );
buf \U$8073 ( \14371 , \13778 );
buf \U$8074 ( \14372 , \13778 );
nor \U$8075 ( \14373 , \13765 , \13807 , \13808 , \13809 , \13771 , \13775 , \13778 , \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 , \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 , \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 , \14372 );
and \U$8076 ( \14374 , \7864 , \14373 );
buf \U$8077 ( \14375 , \13778 );
buf \U$8078 ( \14376 , \13778 );
buf \U$8079 ( \14377 , \13778 );
buf \U$8080 ( \14378 , \13778 );
buf \U$8081 ( \14379 , \13778 );
buf \U$8082 ( \14380 , \13778 );
buf \U$8083 ( \14381 , \13778 );
buf \U$8084 ( \14382 , \13778 );
buf \U$8085 ( \14383 , \13778 );
buf \U$8086 ( \14384 , \13778 );
buf \U$8087 ( \14385 , \13778 );
buf \U$8088 ( \14386 , \13778 );
buf \U$8089 ( \14387 , \13778 );
buf \U$8090 ( \14388 , \13778 );
buf \U$8091 ( \14389 , \13778 );
buf \U$8092 ( \14390 , \13778 );
buf \U$8093 ( \14391 , \13778 );
buf \U$8094 ( \14392 , \13778 );
buf \U$8095 ( \14393 , \13778 );
buf \U$8096 ( \14394 , \13778 );
buf \U$8097 ( \14395 , \13778 );
buf \U$8098 ( \14396 , \13778 );
buf \U$8099 ( \14397 , \13778 );
buf \U$8100 ( \14398 , \13778 );
buf \U$8101 ( \14399 , \13778 );
nor \U$8102 ( \14400 , \13806 , \13766 , \13808 , \13809 , \13771 , \13775 , \13778 , \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 , \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 , \14395 , \14396 , \14397 , \14398 , \14399 );
and \U$8103 ( \14401 , \7892 , \14400 );
buf \U$8104 ( \14402 , \13778 );
buf \U$8105 ( \14403 , \13778 );
buf \U$8106 ( \14404 , \13778 );
buf \U$8107 ( \14405 , \13778 );
buf \U$8108 ( \14406 , \13778 );
buf \U$8109 ( \14407 , \13778 );
buf \U$8110 ( \14408 , \13778 );
buf \U$8111 ( \14409 , \13778 );
buf \U$8112 ( \14410 , \13778 );
buf \U$8113 ( \14411 , \13778 );
buf \U$8114 ( \14412 , \13778 );
buf \U$8115 ( \14413 , \13778 );
buf \U$8116 ( \14414 , \13778 );
buf \U$8117 ( \14415 , \13778 );
buf \U$8118 ( \14416 , \13778 );
buf \U$8119 ( \14417 , \13778 );
buf \U$8120 ( \14418 , \13778 );
buf \U$8121 ( \14419 , \13778 );
buf \U$8122 ( \14420 , \13778 );
buf \U$8123 ( \14421 , \13778 );
buf \U$8124 ( \14422 , \13778 );
buf \U$8125 ( \14423 , \13778 );
buf \U$8126 ( \14424 , \13778 );
buf \U$8127 ( \14425 , \13778 );
buf \U$8128 ( \14426 , \13778 );
nor \U$8129 ( \14427 , \13765 , \13766 , \13808 , \13809 , \13771 , \13775 , \13778 , \14402 , \14403 , \14404 , \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 , \14412 , \14413 , \14414 , \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 , \14425 , \14426 );
and \U$8130 ( \14428 , \7920 , \14427 );
buf \U$8131 ( \14429 , \13778 );
buf \U$8132 ( \14430 , \13778 );
buf \U$8133 ( \14431 , \13778 );
buf \U$8134 ( \14432 , \13778 );
buf \U$8135 ( \14433 , \13778 );
buf \U$8136 ( \14434 , \13778 );
buf \U$8137 ( \14435 , \13778 );
buf \U$8138 ( \14436 , \13778 );
buf \U$8139 ( \14437 , \13778 );
buf \U$8140 ( \14438 , \13778 );
buf \U$8141 ( \14439 , \13778 );
buf \U$8142 ( \14440 , \13778 );
buf \U$8143 ( \14441 , \13778 );
buf \U$8144 ( \14442 , \13778 );
buf \U$8145 ( \14443 , \13778 );
buf \U$8146 ( \14444 , \13778 );
buf \U$8147 ( \14445 , \13778 );
buf \U$8148 ( \14446 , \13778 );
buf \U$8149 ( \14447 , \13778 );
buf \U$8150 ( \14448 , \13778 );
buf \U$8151 ( \14449 , \13778 );
buf \U$8152 ( \14450 , \13778 );
buf \U$8153 ( \14451 , \13778 );
buf \U$8154 ( \14452 , \13778 );
buf \U$8155 ( \14453 , \13778 );
nor \U$8156 ( \14454 , \13806 , \13807 , \13767 , \13809 , \13771 , \13775 , \13778 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 , \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 , \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 , \14452 , \14453 );
and \U$8157 ( \14455 , \7948 , \14454 );
buf \U$8158 ( \14456 , \13778 );
buf \U$8159 ( \14457 , \13778 );
buf \U$8160 ( \14458 , \13778 );
buf \U$8161 ( \14459 , \13778 );
buf \U$8162 ( \14460 , \13778 );
buf \U$8163 ( \14461 , \13778 );
buf \U$8164 ( \14462 , \13778 );
buf \U$8165 ( \14463 , \13778 );
buf \U$8166 ( \14464 , \13778 );
buf \U$8167 ( \14465 , \13778 );
buf \U$8168 ( \14466 , \13778 );
buf \U$8169 ( \14467 , \13778 );
buf \U$8170 ( \14468 , \13778 );
buf \U$8171 ( \14469 , \13778 );
buf \U$8172 ( \14470 , \13778 );
buf \U$8173 ( \14471 , \13778 );
buf \U$8174 ( \14472 , \13778 );
buf \U$8175 ( \14473 , \13778 );
buf \U$8176 ( \14474 , \13778 );
buf \U$8177 ( \14475 , \13778 );
buf \U$8178 ( \14476 , \13778 );
buf \U$8179 ( \14477 , \13778 );
buf \U$8180 ( \14478 , \13778 );
buf \U$8181 ( \14479 , \13778 );
buf \U$8182 ( \14480 , \13778 );
nor \U$8183 ( \14481 , \13765 , \13807 , \13767 , \13809 , \13771 , \13775 , \13778 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 , \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 , \14475 , \14476 , \14477 , \14478 , \14479 , \14480 );
and \U$8184 ( \14482 , \7976 , \14481 );
buf \U$8185 ( \14483 , \13778 );
buf \U$8186 ( \14484 , \13778 );
buf \U$8187 ( \14485 , \13778 );
buf \U$8188 ( \14486 , \13778 );
buf \U$8189 ( \14487 , \13778 );
buf \U$8190 ( \14488 , \13778 );
buf \U$8191 ( \14489 , \13778 );
buf \U$8192 ( \14490 , \13778 );
buf \U$8193 ( \14491 , \13778 );
buf \U$8194 ( \14492 , \13778 );
buf \U$8195 ( \14493 , \13778 );
buf \U$8196 ( \14494 , \13778 );
buf \U$8197 ( \14495 , \13778 );
buf \U$8198 ( \14496 , \13778 );
buf \U$8199 ( \14497 , \13778 );
buf \U$8200 ( \14498 , \13778 );
buf \U$8201 ( \14499 , \13778 );
buf \U$8202 ( \14500 , \13778 );
buf \U$8203 ( \14501 , \13778 );
buf \U$8204 ( \14502 , \13778 );
buf \U$8205 ( \14503 , \13778 );
buf \U$8206 ( \14504 , \13778 );
buf \U$8207 ( \14505 , \13778 );
buf \U$8208 ( \14506 , \13778 );
buf \U$8209 ( \14507 , \13778 );
nor \U$8210 ( \14508 , \13806 , \13766 , \13767 , \13809 , \13771 , \13775 , \13778 , \14483 , \14484 , \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 , \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 , \14505 , \14506 , \14507 );
and \U$8211 ( \14509 , \8004 , \14508 );
buf \U$8212 ( \14510 , \13778 );
buf \U$8213 ( \14511 , \13778 );
buf \U$8214 ( \14512 , \13778 );
buf \U$8215 ( \14513 , \13778 );
buf \U$8216 ( \14514 , \13778 );
buf \U$8217 ( \14515 , \13778 );
buf \U$8218 ( \14516 , \13778 );
buf \U$8219 ( \14517 , \13778 );
buf \U$8220 ( \14518 , \13778 );
buf \U$8221 ( \14519 , \13778 );
buf \U$8222 ( \14520 , \13778 );
buf \U$8223 ( \14521 , \13778 );
buf \U$8224 ( \14522 , \13778 );
buf \U$8225 ( \14523 , \13778 );
buf \U$8226 ( \14524 , \13778 );
buf \U$8227 ( \14525 , \13778 );
buf \U$8228 ( \14526 , \13778 );
buf \U$8229 ( \14527 , \13778 );
buf \U$8230 ( \14528 , \13778 );
buf \U$8231 ( \14529 , \13778 );
buf \U$8232 ( \14530 , \13778 );
buf \U$8233 ( \14531 , \13778 );
buf \U$8234 ( \14532 , \13778 );
buf \U$8235 ( \14533 , \13778 );
buf \U$8236 ( \14534 , \13778 );
nor \U$8237 ( \14535 , \13765 , \13766 , \13767 , \13809 , \13771 , \13775 , \13778 , \14510 , \14511 , \14512 , \14513 , \14514 , \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 , \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 );
and \U$8238 ( \14536 , \8032 , \14535 );
buf \U$8239 ( \14537 , \13778 );
buf \U$8240 ( \14538 , \13778 );
buf \U$8241 ( \14539 , \13778 );
buf \U$8242 ( \14540 , \13778 );
buf \U$8243 ( \14541 , \13778 );
buf \U$8244 ( \14542 , \13778 );
buf \U$8245 ( \14543 , \13778 );
buf \U$8246 ( \14544 , \13778 );
buf \U$8247 ( \14545 , \13778 );
buf \U$8248 ( \14546 , \13778 );
buf \U$8249 ( \14547 , \13778 );
buf \U$8250 ( \14548 , \13778 );
buf \U$8251 ( \14549 , \13778 );
buf \U$8252 ( \14550 , \13778 );
buf \U$8253 ( \14551 , \13778 );
buf \U$8254 ( \14552 , \13778 );
buf \U$8255 ( \14553 , \13778 );
buf \U$8256 ( \14554 , \13778 );
buf \U$8257 ( \14555 , \13778 );
buf \U$8258 ( \14556 , \13778 );
buf \U$8259 ( \14557 , \13778 );
buf \U$8260 ( \14558 , \13778 );
buf \U$8261 ( \14559 , \13778 );
buf \U$8262 ( \14560 , \13778 );
buf \U$8263 ( \14561 , \13778 );
nor \U$8264 ( \14562 , \13806 , \13807 , \13808 , \13768 , \13771 , \13775 , \13778 , \14537 , \14538 , \14539 , \14540 , \14541 , \14542 , \14543 , \14544 , \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 , \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 );
and \U$8265 ( \14563 , \8060 , \14562 );
buf \U$8266 ( \14564 , \13778 );
buf \U$8267 ( \14565 , \13778 );
buf \U$8268 ( \14566 , \13778 );
buf \U$8269 ( \14567 , \13778 );
buf \U$8270 ( \14568 , \13778 );
buf \U$8271 ( \14569 , \13778 );
buf \U$8272 ( \14570 , \13778 );
buf \U$8273 ( \14571 , \13778 );
buf \U$8274 ( \14572 , \13778 );
buf \U$8275 ( \14573 , \13778 );
buf \U$8276 ( \14574 , \13778 );
buf \U$8277 ( \14575 , \13778 );
buf \U$8278 ( \14576 , \13778 );
buf \U$8279 ( \14577 , \13778 );
buf \U$8280 ( \14578 , \13778 );
buf \U$8281 ( \14579 , \13778 );
buf \U$8282 ( \14580 , \13778 );
buf \U$8283 ( \14581 , \13778 );
buf \U$8284 ( \14582 , \13778 );
buf \U$8285 ( \14583 , \13778 );
buf \U$8286 ( \14584 , \13778 );
buf \U$8287 ( \14585 , \13778 );
buf \U$8288 ( \14586 , \13778 );
buf \U$8289 ( \14587 , \13778 );
buf \U$8290 ( \14588 , \13778 );
nor \U$8291 ( \14589 , \13765 , \13807 , \13808 , \13768 , \13771 , \13775 , \13778 , \14564 , \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 , \14572 , \14573 , \14574 , \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 , \14582 , \14583 , \14584 , \14585 , \14586 , \14587 , \14588 );
and \U$8292 ( \14590 , \8088 , \14589 );
buf \U$8293 ( \14591 , \13778 );
buf \U$8294 ( \14592 , \13778 );
buf \U$8295 ( \14593 , \13778 );
buf \U$8296 ( \14594 , \13778 );
buf \U$8297 ( \14595 , \13778 );
buf \U$8298 ( \14596 , \13778 );
buf \U$8299 ( \14597 , \13778 );
buf \U$8300 ( \14598 , \13778 );
buf \U$8301 ( \14599 , \13778 );
buf \U$8302 ( \14600 , \13778 );
buf \U$8303 ( \14601 , \13778 );
buf \U$8304 ( \14602 , \13778 );
buf \U$8305 ( \14603 , \13778 );
buf \U$8306 ( \14604 , \13778 );
buf \U$8307 ( \14605 , \13778 );
buf \U$8308 ( \14606 , \13778 );
buf \U$8309 ( \14607 , \13778 );
buf \U$8310 ( \14608 , \13778 );
buf \U$8311 ( \14609 , \13778 );
buf \U$8312 ( \14610 , \13778 );
buf \U$8313 ( \14611 , \13778 );
buf \U$8314 ( \14612 , \13778 );
buf \U$8315 ( \14613 , \13778 );
buf \U$8316 ( \14614 , \13778 );
buf \U$8317 ( \14615 , \13778 );
nor \U$8318 ( \14616 , \13806 , \13766 , \13808 , \13768 , \13771 , \13775 , \13778 , \14591 , \14592 , \14593 , \14594 , \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 , \14602 , \14603 , \14604 , \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 , \14612 , \14613 , \14614 , \14615 );
and \U$8319 ( \14617 , \8116 , \14616 );
buf \U$8320 ( \14618 , \13778 );
buf \U$8321 ( \14619 , \13778 );
buf \U$8322 ( \14620 , \13778 );
buf \U$8323 ( \14621 , \13778 );
buf \U$8324 ( \14622 , \13778 );
buf \U$8325 ( \14623 , \13778 );
buf \U$8326 ( \14624 , \13778 );
buf \U$8327 ( \14625 , \13778 );
buf \U$8328 ( \14626 , \13778 );
buf \U$8329 ( \14627 , \13778 );
buf \U$8330 ( \14628 , \13778 );
buf \U$8331 ( \14629 , \13778 );
buf \U$8332 ( \14630 , \13778 );
buf \U$8333 ( \14631 , \13778 );
buf \U$8334 ( \14632 , \13778 );
buf \U$8335 ( \14633 , \13778 );
buf \U$8336 ( \14634 , \13778 );
buf \U$8337 ( \14635 , \13778 );
buf \U$8338 ( \14636 , \13778 );
buf \U$8339 ( \14637 , \13778 );
buf \U$8340 ( \14638 , \13778 );
buf \U$8341 ( \14639 , \13778 );
buf \U$8342 ( \14640 , \13778 );
buf \U$8343 ( \14641 , \13778 );
buf \U$8344 ( \14642 , \13778 );
nor \U$8345 ( \14643 , \13765 , \13766 , \13808 , \13768 , \13771 , \13775 , \13778 , \14618 , \14619 , \14620 , \14621 , \14622 , \14623 , \14624 , \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 , \14632 , \14633 , \14634 , \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 , \14642 );
and \U$8346 ( \14644 , \8144 , \14643 );
buf \U$8347 ( \14645 , \13778 );
buf \U$8348 ( \14646 , \13778 );
buf \U$8349 ( \14647 , \13778 );
buf \U$8350 ( \14648 , \13778 );
buf \U$8351 ( \14649 , \13778 );
buf \U$8352 ( \14650 , \13778 );
buf \U$8353 ( \14651 , \13778 );
buf \U$8354 ( \14652 , \13778 );
buf \U$8355 ( \14653 , \13778 );
buf \U$8356 ( \14654 , \13778 );
buf \U$8357 ( \14655 , \13778 );
buf \U$8358 ( \14656 , \13778 );
buf \U$8359 ( \14657 , \13778 );
buf \U$8360 ( \14658 , \13778 );
buf \U$8361 ( \14659 , \13778 );
buf \U$8362 ( \14660 , \13778 );
buf \U$8363 ( \14661 , \13778 );
buf \U$8364 ( \14662 , \13778 );
buf \U$8365 ( \14663 , \13778 );
buf \U$8366 ( \14664 , \13778 );
buf \U$8367 ( \14665 , \13778 );
buf \U$8368 ( \14666 , \13778 );
buf \U$8369 ( \14667 , \13778 );
buf \U$8370 ( \14668 , \13778 );
buf \U$8371 ( \14669 , \13778 );
nor \U$8372 ( \14670 , \13806 , \13807 , \13767 , \13768 , \13771 , \13775 , \13778 , \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 , \14652 , \14653 , \14654 , \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 , \14662 , \14663 , \14664 , \14665 , \14666 , \14667 , \14668 , \14669 );
and \U$8373 ( \14671 , \8172 , \14670 );
buf \U$8374 ( \14672 , \13778 );
buf \U$8375 ( \14673 , \13778 );
buf \U$8376 ( \14674 , \13778 );
buf \U$8377 ( \14675 , \13778 );
buf \U$8378 ( \14676 , \13778 );
buf \U$8379 ( \14677 , \13778 );
buf \U$8380 ( \14678 , \13778 );
buf \U$8381 ( \14679 , \13778 );
buf \U$8382 ( \14680 , \13778 );
buf \U$8383 ( \14681 , \13778 );
buf \U$8384 ( \14682 , \13778 );
buf \U$8385 ( \14683 , \13778 );
buf \U$8386 ( \14684 , \13778 );
buf \U$8387 ( \14685 , \13778 );
buf \U$8388 ( \14686 , \13778 );
buf \U$8389 ( \14687 , \13778 );
buf \U$8390 ( \14688 , \13778 );
buf \U$8391 ( \14689 , \13778 );
buf \U$8392 ( \14690 , \13778 );
buf \U$8393 ( \14691 , \13778 );
buf \U$8394 ( \14692 , \13778 );
buf \U$8395 ( \14693 , \13778 );
buf \U$8396 ( \14694 , \13778 );
buf \U$8397 ( \14695 , \13778 );
buf \U$8398 ( \14696 , \13778 );
nor \U$8399 ( \14697 , \13765 , \13807 , \13767 , \13768 , \13771 , \13775 , \13778 , \14672 , \14673 , \14674 , \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 , \14682 , \14683 , \14684 , \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 , \14692 , \14693 , \14694 , \14695 , \14696 );
and \U$8400 ( \14698 , \8200 , \14697 );
buf \U$8401 ( \14699 , \13778 );
buf \U$8402 ( \14700 , \13778 );
buf \U$8403 ( \14701 , \13778 );
buf \U$8404 ( \14702 , \13778 );
buf \U$8405 ( \14703 , \13778 );
buf \U$8406 ( \14704 , \13778 );
buf \U$8407 ( \14705 , \13778 );
buf \U$8408 ( \14706 , \13778 );
buf \U$8409 ( \14707 , \13778 );
buf \U$8410 ( \14708 , \13778 );
buf \U$8411 ( \14709 , \13778 );
buf \U$8412 ( \14710 , \13778 );
buf \U$8413 ( \14711 , \13778 );
buf \U$8414 ( \14712 , \13778 );
buf \U$8415 ( \14713 , \13778 );
buf \U$8416 ( \14714 , \13778 );
buf \U$8417 ( \14715 , \13778 );
buf \U$8418 ( \14716 , \13778 );
buf \U$8419 ( \14717 , \13778 );
buf \U$8420 ( \14718 , \13778 );
buf \U$8421 ( \14719 , \13778 );
buf \U$8422 ( \14720 , \13778 );
buf \U$8423 ( \14721 , \13778 );
buf \U$8424 ( \14722 , \13778 );
buf \U$8425 ( \14723 , \13778 );
nor \U$8426 ( \14724 , \13806 , \13766 , \13767 , \13768 , \13771 , \13775 , \13778 , \14699 , \14700 , \14701 , \14702 , \14703 , \14704 , \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 , \14712 , \14713 , \14714 , \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 , \14722 , \14723 );
and \U$8427 ( \14725 , \8228 , \14724 );
or \U$8428 ( \14726 , \14320 , \14347 , \14374 , \14401 , \14428 , \14455 , \14482 , \14509 , \14536 , \14563 , \14590 , \14617 , \14644 , \14671 , \14698 , \14725 );
buf \U$8429 ( \14727 , \13778 );
not \U$8430 ( \14728 , \14727 );
buf \U$8431 ( \14729 , \13766 );
buf \U$8432 ( \14730 , \13767 );
buf \U$8433 ( \14731 , \13768 );
buf \U$8434 ( \14732 , \13771 );
buf \U$8435 ( \14733 , \13775 );
buf \U$8436 ( \14734 , \13778 );
buf \U$8437 ( \14735 , \13778 );
buf \U$8438 ( \14736 , \13778 );
buf \U$8439 ( \14737 , \13778 );
buf \U$8440 ( \14738 , \13778 );
buf \U$8441 ( \14739 , \13778 );
buf \U$8442 ( \14740 , \13778 );
buf \U$8443 ( \14741 , \13778 );
buf \U$8444 ( \14742 , \13778 );
buf \U$8445 ( \14743 , \13778 );
buf \U$8446 ( \14744 , \13778 );
buf \U$8447 ( \14745 , \13778 );
buf \U$8448 ( \14746 , \13778 );
buf \U$8449 ( \14747 , \13778 );
buf \U$8450 ( \14748 , \13778 );
buf \U$8451 ( \14749 , \13778 );
buf \U$8452 ( \14750 , \13778 );
buf \U$8453 ( \14751 , \13778 );
buf \U$8454 ( \14752 , \13778 );
buf \U$8455 ( \14753 , \13778 );
buf \U$8456 ( \14754 , \13778 );
buf \U$8457 ( \14755 , \13778 );
buf \U$8458 ( \14756 , \13778 );
buf \U$8459 ( \14757 , \13778 );
buf \U$8460 ( \14758 , \13778 );
buf \U$8461 ( \14759 , \13765 );
or \U$8462 ( \14760 , \14729 , \14730 , \14731 , \14732 , \14733 , \14734 , \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 , \14742 , \14743 , \14744 , \14745 , \14746 , \14747 , \14748 , \14749 , \14750 , \14751 , \14752 , \14753 , \14754 , \14755 , \14756 , \14757 , \14758 , \14759 );
nand \U$8463 ( \14761 , \14728 , \14760 );
buf \U$8464 ( \14762 , \14761 );
buf \U$8465 ( \14763 , \13778 );
not \U$8466 ( \14764 , \14763 );
buf \U$8467 ( \14765 , \13775 );
buf \U$8468 ( \14766 , \13778 );
buf \U$8469 ( \14767 , \13778 );
buf \U$8470 ( \14768 , \13778 );
buf \U$8471 ( \14769 , \13778 );
buf \U$8472 ( \14770 , \13778 );
buf \U$8473 ( \14771 , \13778 );
buf \U$8474 ( \14772 , \13778 );
buf \U$8475 ( \14773 , \13778 );
buf \U$8476 ( \14774 , \13778 );
buf \U$8477 ( \14775 , \13778 );
buf \U$8478 ( \14776 , \13778 );
buf \U$8479 ( \14777 , \13778 );
buf \U$8480 ( \14778 , \13778 );
buf \U$8481 ( \14779 , \13778 );
buf \U$8482 ( \14780 , \13778 );
buf \U$8483 ( \14781 , \13778 );
buf \U$8484 ( \14782 , \13778 );
buf \U$8485 ( \14783 , \13778 );
buf \U$8486 ( \14784 , \13778 );
buf \U$8487 ( \14785 , \13778 );
buf \U$8488 ( \14786 , \13778 );
buf \U$8489 ( \14787 , \13778 );
buf \U$8490 ( \14788 , \13778 );
buf \U$8491 ( \14789 , \13778 );
buf \U$8492 ( \14790 , \13778 );
buf \U$8493 ( \14791 , \13771 );
buf \U$8494 ( \14792 , \13765 );
buf \U$8495 ( \14793 , \13766 );
buf \U$8496 ( \14794 , \13767 );
buf \U$8497 ( \14795 , \13768 );
or \U$8498 ( \14796 , \14792 , \14793 , \14794 , \14795 );
and \U$8499 ( \14797 , \14791 , \14796 );
or \U$8500 ( \14798 , \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 , \14772 , \14773 , \14774 , \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 , \14782 , \14783 , \14784 , \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14797 );
and \U$8501 ( \14799 , \14764 , \14798 );
buf \U$8502 ( \14800 , \14799 );
or \U$8503 ( \14801 , \14762 , \14800 );
_DC g509e ( \14802_nG509e , \14726 , \14801 );
buf \U$8504 ( \14803 , \14802_nG509e );
xor \U$8505 ( \14804 , \14293 , \14803 );
buf \U$8506 ( \14805 , RIb7b9590_247);
and \U$8507 ( \14806 , \7126 , \14319 );
and \U$8508 ( \14807 , \7128 , \14346 );
and \U$8509 ( \14808 , \8338 , \14373 );
and \U$8510 ( \14809 , \8340 , \14400 );
and \U$8511 ( \14810 , \8342 , \14427 );
and \U$8512 ( \14811 , \8344 , \14454 );
and \U$8513 ( \14812 , \8346 , \14481 );
and \U$8514 ( \14813 , \8348 , \14508 );
and \U$8515 ( \14814 , \8350 , \14535 );
and \U$8516 ( \14815 , \8352 , \14562 );
and \U$8517 ( \14816 , \8354 , \14589 );
and \U$8518 ( \14817 , \8356 , \14616 );
and \U$8519 ( \14818 , \8358 , \14643 );
and \U$8520 ( \14819 , \8360 , \14670 );
and \U$8521 ( \14820 , \8362 , \14697 );
and \U$8522 ( \14821 , \8364 , \14724 );
or \U$8523 ( \14822 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 , \14812 , \14813 , \14814 , \14815 , \14816 , \14817 , \14818 , \14819 , \14820 , \14821 );
_DC g50b3 ( \14823_nG50b3 , \14822 , \14801 );
buf \U$8524 ( \14824 , \14823_nG50b3 );
xor \U$8525 ( \14825 , \14805 , \14824 );
or \U$8526 ( \14826 , \14804 , \14825 );
buf \U$8527 ( \14827 , RIb7b9518_248);
and \U$8528 ( \14828 , \7136 , \14319 );
and \U$8529 ( \14829 , \7138 , \14346 );
and \U$8530 ( \14830 , \8374 , \14373 );
and \U$8531 ( \14831 , \8376 , \14400 );
and \U$8532 ( \14832 , \8378 , \14427 );
and \U$8533 ( \14833 , \8380 , \14454 );
and \U$8534 ( \14834 , \8382 , \14481 );
and \U$8535 ( \14835 , \8384 , \14508 );
and \U$8536 ( \14836 , \8386 , \14535 );
and \U$8537 ( \14837 , \8388 , \14562 );
and \U$8538 ( \14838 , \8390 , \14589 );
and \U$8539 ( \14839 , \8392 , \14616 );
and \U$8540 ( \14840 , \8394 , \14643 );
and \U$8541 ( \14841 , \8396 , \14670 );
and \U$8542 ( \14842 , \8398 , \14697 );
and \U$8543 ( \14843 , \8400 , \14724 );
or \U$8544 ( \14844 , \14828 , \14829 , \14830 , \14831 , \14832 , \14833 , \14834 , \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 , \14842 , \14843 );
_DC g50c9 ( \14845_nG50c9 , \14844 , \14801 );
buf \U$8545 ( \14846 , \14845_nG50c9 );
xor \U$8546 ( \14847 , \14827 , \14846 );
or \U$8547 ( \14848 , \14826 , \14847 );
buf \U$8548 ( \14849 , RIb7b94a0_249);
and \U$8549 ( \14850 , \7146 , \14319 );
and \U$8550 ( \14851 , \7148 , \14346 );
and \U$8551 ( \14852 , \8410 , \14373 );
and \U$8552 ( \14853 , \8412 , \14400 );
and \U$8553 ( \14854 , \8414 , \14427 );
and \U$8554 ( \14855 , \8416 , \14454 );
and \U$8555 ( \14856 , \8418 , \14481 );
and \U$8556 ( \14857 , \8420 , \14508 );
and \U$8557 ( \14858 , \8422 , \14535 );
and \U$8558 ( \14859 , \8424 , \14562 );
and \U$8559 ( \14860 , \8426 , \14589 );
and \U$8560 ( \14861 , \8428 , \14616 );
and \U$8561 ( \14862 , \8430 , \14643 );
and \U$8562 ( \14863 , \8432 , \14670 );
and \U$8563 ( \14864 , \8434 , \14697 );
and \U$8564 ( \14865 , \8436 , \14724 );
or \U$8565 ( \14866 , \14850 , \14851 , \14852 , \14853 , \14854 , \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 , \14862 , \14863 , \14864 , \14865 );
_DC g50df ( \14867_nG50df , \14866 , \14801 );
buf \U$8566 ( \14868 , \14867_nG50df );
xor \U$8567 ( \14869 , \14849 , \14868 );
or \U$8568 ( \14870 , \14848 , \14869 );
buf \U$8569 ( \14871 , RIb7b9428_250);
and \U$8570 ( \14872 , \7156 , \14319 );
and \U$8571 ( \14873 , \7158 , \14346 );
and \U$8572 ( \14874 , \8446 , \14373 );
and \U$8573 ( \14875 , \8448 , \14400 );
and \U$8574 ( \14876 , \8450 , \14427 );
and \U$8575 ( \14877 , \8452 , \14454 );
and \U$8576 ( \14878 , \8454 , \14481 );
and \U$8577 ( \14879 , \8456 , \14508 );
and \U$8578 ( \14880 , \8458 , \14535 );
and \U$8579 ( \14881 , \8460 , \14562 );
and \U$8580 ( \14882 , \8462 , \14589 );
and \U$8581 ( \14883 , \8464 , \14616 );
and \U$8582 ( \14884 , \8466 , \14643 );
and \U$8583 ( \14885 , \8468 , \14670 );
and \U$8584 ( \14886 , \8470 , \14697 );
and \U$8585 ( \14887 , \8472 , \14724 );
or \U$8586 ( \14888 , \14872 , \14873 , \14874 , \14875 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 , \14882 , \14883 , \14884 , \14885 , \14886 , \14887 );
_DC g50f5 ( \14889_nG50f5 , \14888 , \14801 );
buf \U$8587 ( \14890 , \14889_nG50f5 );
xor \U$8588 ( \14891 , \14871 , \14890 );
or \U$8589 ( \14892 , \14870 , \14891 );
buf \U$8590 ( \14893 , RIb7b93b0_251);
and \U$8591 ( \14894 , \7166 , \14319 );
and \U$8592 ( \14895 , \7168 , \14346 );
and \U$8593 ( \14896 , \8482 , \14373 );
and \U$8594 ( \14897 , \8484 , \14400 );
and \U$8595 ( \14898 , \8486 , \14427 );
and \U$8596 ( \14899 , \8488 , \14454 );
and \U$8597 ( \14900 , \8490 , \14481 );
and \U$8598 ( \14901 , \8492 , \14508 );
and \U$8599 ( \14902 , \8494 , \14535 );
and \U$8600 ( \14903 , \8496 , \14562 );
and \U$8601 ( \14904 , \8498 , \14589 );
and \U$8602 ( \14905 , \8500 , \14616 );
and \U$8603 ( \14906 , \8502 , \14643 );
and \U$8604 ( \14907 , \8504 , \14670 );
and \U$8605 ( \14908 , \8506 , \14697 );
and \U$8606 ( \14909 , \8508 , \14724 );
or \U$8607 ( \14910 , \14894 , \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 , \14902 , \14903 , \14904 , \14905 , \14906 , \14907 , \14908 , \14909 );
_DC g510b ( \14911_nG510b , \14910 , \14801 );
buf \U$8608 ( \14912 , \14911_nG510b );
xor \U$8609 ( \14913 , \14893 , \14912 );
or \U$8610 ( \14914 , \14892 , \14913 );
buf \U$8611 ( \14915 , RIb7af720_252);
and \U$8612 ( \14916 , \7176 , \14319 );
and \U$8613 ( \14917 , \7178 , \14346 );
and \U$8614 ( \14918 , \8518 , \14373 );
and \U$8615 ( \14919 , \8520 , \14400 );
and \U$8616 ( \14920 , \8522 , \14427 );
and \U$8617 ( \14921 , \8524 , \14454 );
and \U$8618 ( \14922 , \8526 , \14481 );
and \U$8619 ( \14923 , \8528 , \14508 );
and \U$8620 ( \14924 , \8530 , \14535 );
and \U$8621 ( \14925 , \8532 , \14562 );
and \U$8622 ( \14926 , \8534 , \14589 );
and \U$8623 ( \14927 , \8536 , \14616 );
and \U$8624 ( \14928 , \8538 , \14643 );
and \U$8625 ( \14929 , \8540 , \14670 );
and \U$8626 ( \14930 , \8542 , \14697 );
and \U$8627 ( \14931 , \8544 , \14724 );
or \U$8628 ( \14932 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 , \14922 , \14923 , \14924 , \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 );
_DC g5121 ( \14933_nG5121 , \14932 , \14801 );
buf \U$8629 ( \14934 , \14933_nG5121 );
xor \U$8630 ( \14935 , \14915 , \14934 );
or \U$8631 ( \14936 , \14914 , \14935 );
buf \U$8632 ( \14937 , RIb7af6a8_253);
and \U$8633 ( \14938 , \7186 , \14319 );
and \U$8634 ( \14939 , \7188 , \14346 );
and \U$8635 ( \14940 , \8554 , \14373 );
and \U$8636 ( \14941 , \8556 , \14400 );
and \U$8637 ( \14942 , \8558 , \14427 );
and \U$8638 ( \14943 , \8560 , \14454 );
and \U$8639 ( \14944 , \8562 , \14481 );
and \U$8640 ( \14945 , \8564 , \14508 );
and \U$8641 ( \14946 , \8566 , \14535 );
and \U$8642 ( \14947 , \8568 , \14562 );
and \U$8643 ( \14948 , \8570 , \14589 );
and \U$8644 ( \14949 , \8572 , \14616 );
and \U$8645 ( \14950 , \8574 , \14643 );
and \U$8646 ( \14951 , \8576 , \14670 );
and \U$8647 ( \14952 , \8578 , \14697 );
and \U$8648 ( \14953 , \8580 , \14724 );
or \U$8649 ( \14954 , \14938 , \14939 , \14940 , \14941 , \14942 , \14943 , \14944 , \14945 , \14946 , \14947 , \14948 , \14949 , \14950 , \14951 , \14952 , \14953 );
_DC g5137 ( \14955_nG5137 , \14954 , \14801 );
buf \U$8650 ( \14956 , \14955_nG5137 );
xor \U$8651 ( \14957 , \14937 , \14956 );
or \U$8652 ( \14958 , \14936 , \14957 );
not \U$8653 ( \14959 , \14958 );
buf \U$8654 ( \14960 , \14959 );
and \U$8655 ( \14961 , \14292 , \14960 );
buf \U$8656 ( \14962 , RIb7af630_254);
buf \U$8657 ( \14963 , \13778 );
buf \U$8658 ( \14964 , \13778 );
buf \U$8659 ( \14965 , \13778 );
buf \U$8660 ( \14966 , \13778 );
buf \U$8661 ( \14967 , \13778 );
buf \U$8662 ( \14968 , \13778 );
buf \U$8663 ( \14969 , \13778 );
buf \U$8664 ( \14970 , \13778 );
buf \U$8665 ( \14971 , \13778 );
buf \U$8666 ( \14972 , \13778 );
buf \U$8667 ( \14973 , \13778 );
buf \U$8668 ( \14974 , \13778 );
buf \U$8669 ( \14975 , \13778 );
buf \U$8670 ( \14976 , \13778 );
buf \U$8671 ( \14977 , \13778 );
buf \U$8672 ( \14978 , \13778 );
buf \U$8673 ( \14979 , \13778 );
buf \U$8674 ( \14980 , \13778 );
buf \U$8675 ( \14981 , \13778 );
buf \U$8676 ( \14982 , \13778 );
buf \U$8677 ( \14983 , \13778 );
buf \U$8678 ( \14984 , \13778 );
buf \U$8679 ( \14985 , \13778 );
buf \U$8680 ( \14986 , \13778 );
buf \U$8681 ( \14987 , \13778 );
nor \U$8682 ( \14988 , \13765 , \13766 , \13767 , \13768 , \13772 , \13775 , \13778 , \14963 , \14964 , \14965 , \14966 , \14967 , \14968 , \14969 , \14970 , \14971 , \14972 , \14973 , \14974 , \14975 , \14976 , \14977 , \14978 , \14979 , \14980 , \14981 , \14982 , \14983 , \14984 , \14985 , \14986 , \14987 );
and \U$8683 ( \14989 , \7198 , \14988 );
buf \U$8684 ( \14990 , \13778 );
buf \U$8685 ( \14991 , \13778 );
buf \U$8686 ( \14992 , \13778 );
buf \U$8687 ( \14993 , \13778 );
buf \U$8688 ( \14994 , \13778 );
buf \U$8689 ( \14995 , \13778 );
buf \U$8690 ( \14996 , \13778 );
buf \U$8691 ( \14997 , \13778 );
buf \U$8692 ( \14998 , \13778 );
buf \U$8693 ( \14999 , \13778 );
buf \U$8694 ( \15000 , \13778 );
buf \U$8695 ( \15001 , \13778 );
buf \U$8696 ( \15002 , \13778 );
buf \U$8697 ( \15003 , \13778 );
buf \U$8698 ( \15004 , \13778 );
buf \U$8699 ( \15005 , \13778 );
buf \U$8700 ( \15006 , \13778 );
buf \U$8701 ( \15007 , \13778 );
buf \U$8702 ( \15008 , \13778 );
buf \U$8703 ( \15009 , \13778 );
buf \U$8704 ( \15010 , \13778 );
buf \U$8705 ( \15011 , \13778 );
buf \U$8706 ( \15012 , \13778 );
buf \U$8707 ( \15013 , \13778 );
buf \U$8708 ( \15014 , \13778 );
nor \U$8709 ( \15015 , \13806 , \13807 , \13808 , \13809 , \13771 , \13775 , \13778 , \14990 , \14991 , \14992 , \14993 , \14994 , \14995 , \14996 , \14997 , \14998 , \14999 , \15000 , \15001 , \15002 , \15003 , \15004 , \15005 , \15006 , \15007 , \15008 , \15009 , \15010 , \15011 , \15012 , \15013 , \15014 );
and \U$8710 ( \15016 , \7200 , \15015 );
buf \U$8711 ( \15017 , \13778 );
buf \U$8712 ( \15018 , \13778 );
buf \U$8713 ( \15019 , \13778 );
buf \U$8714 ( \15020 , \13778 );
buf \U$8715 ( \15021 , \13778 );
buf \U$8716 ( \15022 , \13778 );
buf \U$8717 ( \15023 , \13778 );
buf \U$8718 ( \15024 , \13778 );
buf \U$8719 ( \15025 , \13778 );
buf \U$8720 ( \15026 , \13778 );
buf \U$8721 ( \15027 , \13778 );
buf \U$8722 ( \15028 , \13778 );
buf \U$8723 ( \15029 , \13778 );
buf \U$8724 ( \15030 , \13778 );
buf \U$8725 ( \15031 , \13778 );
buf \U$8726 ( \15032 , \13778 );
buf \U$8727 ( \15033 , \13778 );
buf \U$8728 ( \15034 , \13778 );
buf \U$8729 ( \15035 , \13778 );
buf \U$8730 ( \15036 , \13778 );
buf \U$8731 ( \15037 , \13778 );
buf \U$8732 ( \15038 , \13778 );
buf \U$8733 ( \15039 , \13778 );
buf \U$8734 ( \15040 , \13778 );
buf \U$8735 ( \15041 , \13778 );
nor \U$8736 ( \15042 , \13765 , \13807 , \13808 , \13809 , \13771 , \13775 , \13778 , \15017 , \15018 , \15019 , \15020 , \15021 , \15022 , \15023 , \15024 , \15025 , \15026 , \15027 , \15028 , \15029 , \15030 , \15031 , \15032 , \15033 , \15034 , \15035 , \15036 , \15037 , \15038 , \15039 , \15040 , \15041 );
and \U$8737 ( \15043 , \8645 , \15042 );
buf \U$8738 ( \15044 , \13778 );
buf \U$8739 ( \15045 , \13778 );
buf \U$8740 ( \15046 , \13778 );
buf \U$8741 ( \15047 , \13778 );
buf \U$8742 ( \15048 , \13778 );
buf \U$8743 ( \15049 , \13778 );
buf \U$8744 ( \15050 , \13778 );
buf \U$8745 ( \15051 , \13778 );
buf \U$8746 ( \15052 , \13778 );
buf \U$8747 ( \15053 , \13778 );
buf \U$8748 ( \15054 , \13778 );
buf \U$8749 ( \15055 , \13778 );
buf \U$8750 ( \15056 , \13778 );
buf \U$8751 ( \15057 , \13778 );
buf \U$8752 ( \15058 , \13778 );
buf \U$8753 ( \15059 , \13778 );
buf \U$8754 ( \15060 , \13778 );
buf \U$8755 ( \15061 , \13778 );
buf \U$8756 ( \15062 , \13778 );
buf \U$8757 ( \15063 , \13778 );
buf \U$8758 ( \15064 , \13778 );
buf \U$8759 ( \15065 , \13778 );
buf \U$8760 ( \15066 , \13778 );
buf \U$8761 ( \15067 , \13778 );
buf \U$8762 ( \15068 , \13778 );
nor \U$8763 ( \15069 , \13806 , \13766 , \13808 , \13809 , \13771 , \13775 , \13778 , \15044 , \15045 , \15046 , \15047 , \15048 , \15049 , \15050 , \15051 , \15052 , \15053 , \15054 , \15055 , \15056 , \15057 , \15058 , \15059 , \15060 , \15061 , \15062 , \15063 , \15064 , \15065 , \15066 , \15067 , \15068 );
and \U$8764 ( \15070 , \8673 , \15069 );
buf \U$8765 ( \15071 , \13778 );
buf \U$8766 ( \15072 , \13778 );
buf \U$8767 ( \15073 , \13778 );
buf \U$8768 ( \15074 , \13778 );
buf \U$8769 ( \15075 , \13778 );
buf \U$8770 ( \15076 , \13778 );
buf \U$8771 ( \15077 , \13778 );
buf \U$8772 ( \15078 , \13778 );
buf \U$8773 ( \15079 , \13778 );
buf \U$8774 ( \15080 , \13778 );
buf \U$8775 ( \15081 , \13778 );
buf \U$8776 ( \15082 , \13778 );
buf \U$8777 ( \15083 , \13778 );
buf \U$8778 ( \15084 , \13778 );
buf \U$8779 ( \15085 , \13778 );
buf \U$8780 ( \15086 , \13778 );
buf \U$8781 ( \15087 , \13778 );
buf \U$8782 ( \15088 , \13778 );
buf \U$8783 ( \15089 , \13778 );
buf \U$8784 ( \15090 , \13778 );
buf \U$8785 ( \15091 , \13778 );
buf \U$8786 ( \15092 , \13778 );
buf \U$8787 ( \15093 , \13778 );
buf \U$8788 ( \15094 , \13778 );
buf \U$8789 ( \15095 , \13778 );
nor \U$8790 ( \15096 , \13765 , \13766 , \13808 , \13809 , \13771 , \13775 , \13778 , \15071 , \15072 , \15073 , \15074 , \15075 , \15076 , \15077 , \15078 , \15079 , \15080 , \15081 , \15082 , \15083 , \15084 , \15085 , \15086 , \15087 , \15088 , \15089 , \15090 , \15091 , \15092 , \15093 , \15094 , \15095 );
and \U$8791 ( \15097 , \8701 , \15096 );
buf \U$8792 ( \15098 , \13778 );
buf \U$8793 ( \15099 , \13778 );
buf \U$8794 ( \15100 , \13778 );
buf \U$8795 ( \15101 , \13778 );
buf \U$8796 ( \15102 , \13778 );
buf \U$8797 ( \15103 , \13778 );
buf \U$8798 ( \15104 , \13778 );
buf \U$8799 ( \15105 , \13778 );
buf \U$8800 ( \15106 , \13778 );
buf \U$8801 ( \15107 , \13778 );
buf \U$8802 ( \15108 , \13778 );
buf \U$8803 ( \15109 , \13778 );
buf \U$8804 ( \15110 , \13778 );
buf \U$8805 ( \15111 , \13778 );
buf \U$8806 ( \15112 , \13778 );
buf \U$8807 ( \15113 , \13778 );
buf \U$8808 ( \15114 , \13778 );
buf \U$8809 ( \15115 , \13778 );
buf \U$8810 ( \15116 , \13778 );
buf \U$8811 ( \15117 , \13778 );
buf \U$8812 ( \15118 , \13778 );
buf \U$8813 ( \15119 , \13778 );
buf \U$8814 ( \15120 , \13778 );
buf \U$8815 ( \15121 , \13778 );
buf \U$8816 ( \15122 , \13778 );
nor \U$8817 ( \15123 , \13806 , \13807 , \13767 , \13809 , \13771 , \13775 , \13778 , \15098 , \15099 , \15100 , \15101 , \15102 , \15103 , \15104 , \15105 , \15106 , \15107 , \15108 , \15109 , \15110 , \15111 , \15112 , \15113 , \15114 , \15115 , \15116 , \15117 , \15118 , \15119 , \15120 , \15121 , \15122 );
and \U$8818 ( \15124 , \8729 , \15123 );
buf \U$8819 ( \15125 , \13778 );
buf \U$8820 ( \15126 , \13778 );
buf \U$8821 ( \15127 , \13778 );
buf \U$8822 ( \15128 , \13778 );
buf \U$8823 ( \15129 , \13778 );
buf \U$8824 ( \15130 , \13778 );
buf \U$8825 ( \15131 , \13778 );
buf \U$8826 ( \15132 , \13778 );
buf \U$8827 ( \15133 , \13778 );
buf \U$8828 ( \15134 , \13778 );
buf \U$8829 ( \15135 , \13778 );
buf \U$8830 ( \15136 , \13778 );
buf \U$8831 ( \15137 , \13778 );
buf \U$8832 ( \15138 , \13778 );
buf \U$8833 ( \15139 , \13778 );
buf \U$8834 ( \15140 , \13778 );
buf \U$8835 ( \15141 , \13778 );
buf \U$8836 ( \15142 , \13778 );
buf \U$8837 ( \15143 , \13778 );
buf \U$8838 ( \15144 , \13778 );
buf \U$8839 ( \15145 , \13778 );
buf \U$8840 ( \15146 , \13778 );
buf \U$8841 ( \15147 , \13778 );
buf \U$8842 ( \15148 , \13778 );
buf \U$8843 ( \15149 , \13778 );
nor \U$8844 ( \15150 , \13765 , \13807 , \13767 , \13809 , \13771 , \13775 , \13778 , \15125 , \15126 , \15127 , \15128 , \15129 , \15130 , \15131 , \15132 , \15133 , \15134 , \15135 , \15136 , \15137 , \15138 , \15139 , \15140 , \15141 , \15142 , \15143 , \15144 , \15145 , \15146 , \15147 , \15148 , \15149 );
and \U$8845 ( \15151 , \8757 , \15150 );
buf \U$8846 ( \15152 , \13778 );
buf \U$8847 ( \15153 , \13778 );
buf \U$8848 ( \15154 , \13778 );
buf \U$8849 ( \15155 , \13778 );
buf \U$8850 ( \15156 , \13778 );
buf \U$8851 ( \15157 , \13778 );
buf \U$8852 ( \15158 , \13778 );
buf \U$8853 ( \15159 , \13778 );
buf \U$8854 ( \15160 , \13778 );
buf \U$8855 ( \15161 , \13778 );
buf \U$8856 ( \15162 , \13778 );
buf \U$8857 ( \15163 , \13778 );
buf \U$8858 ( \15164 , \13778 );
buf \U$8859 ( \15165 , \13778 );
buf \U$8860 ( \15166 , \13778 );
buf \U$8861 ( \15167 , \13778 );
buf \U$8862 ( \15168 , \13778 );
buf \U$8863 ( \15169 , \13778 );
buf \U$8864 ( \15170 , \13778 );
buf \U$8865 ( \15171 , \13778 );
buf \U$8866 ( \15172 , \13778 );
buf \U$8867 ( \15173 , \13778 );
buf \U$8868 ( \15174 , \13778 );
buf \U$8869 ( \15175 , \13778 );
buf \U$8870 ( \15176 , \13778 );
nor \U$8871 ( \15177 , \13806 , \13766 , \13767 , \13809 , \13771 , \13775 , \13778 , \15152 , \15153 , \15154 , \15155 , \15156 , \15157 , \15158 , \15159 , \15160 , \15161 , \15162 , \15163 , \15164 , \15165 , \15166 , \15167 , \15168 , \15169 , \15170 , \15171 , \15172 , \15173 , \15174 , \15175 , \15176 );
and \U$8872 ( \15178 , \8785 , \15177 );
buf \U$8873 ( \15179 , \13778 );
buf \U$8874 ( \15180 , \13778 );
buf \U$8875 ( \15181 , \13778 );
buf \U$8876 ( \15182 , \13778 );
buf \U$8877 ( \15183 , \13778 );
buf \U$8878 ( \15184 , \13778 );
buf \U$8879 ( \15185 , \13778 );
buf \U$8880 ( \15186 , \13778 );
buf \U$8881 ( \15187 , \13778 );
buf \U$8882 ( \15188 , \13778 );
buf \U$8883 ( \15189 , \13778 );
buf \U$8884 ( \15190 , \13778 );
buf \U$8885 ( \15191 , \13778 );
buf \U$8886 ( \15192 , \13778 );
buf \U$8887 ( \15193 , \13778 );
buf \U$8888 ( \15194 , \13778 );
buf \U$8889 ( \15195 , \13778 );
buf \U$8890 ( \15196 , \13778 );
buf \U$8891 ( \15197 , \13778 );
buf \U$8892 ( \15198 , \13778 );
buf \U$8893 ( \15199 , \13778 );
buf \U$8894 ( \15200 , \13778 );
buf \U$8895 ( \15201 , \13778 );
buf \U$8896 ( \15202 , \13778 );
buf \U$8897 ( \15203 , \13778 );
nor \U$8898 ( \15204 , \13765 , \13766 , \13767 , \13809 , \13771 , \13775 , \13778 , \15179 , \15180 , \15181 , \15182 , \15183 , \15184 , \15185 , \15186 , \15187 , \15188 , \15189 , \15190 , \15191 , \15192 , \15193 , \15194 , \15195 , \15196 , \15197 , \15198 , \15199 , \15200 , \15201 , \15202 , \15203 );
and \U$8899 ( \15205 , \8813 , \15204 );
buf \U$8900 ( \15206 , \13778 );
buf \U$8901 ( \15207 , \13778 );
buf \U$8902 ( \15208 , \13778 );
buf \U$8903 ( \15209 , \13778 );
buf \U$8904 ( \15210 , \13778 );
buf \U$8905 ( \15211 , \13778 );
buf \U$8906 ( \15212 , \13778 );
buf \U$8907 ( \15213 , \13778 );
buf \U$8908 ( \15214 , \13778 );
buf \U$8909 ( \15215 , \13778 );
buf \U$8910 ( \15216 , \13778 );
buf \U$8911 ( \15217 , \13778 );
buf \U$8912 ( \15218 , \13778 );
buf \U$8913 ( \15219 , \13778 );
buf \U$8914 ( \15220 , \13778 );
buf \U$8915 ( \15221 , \13778 );
buf \U$8916 ( \15222 , \13778 );
buf \U$8917 ( \15223 , \13778 );
buf \U$8918 ( \15224 , \13778 );
buf \U$8919 ( \15225 , \13778 );
buf \U$8920 ( \15226 , \13778 );
buf \U$8921 ( \15227 , \13778 );
buf \U$8922 ( \15228 , \13778 );
buf \U$8923 ( \15229 , \13778 );
buf \U$8924 ( \15230 , \13778 );
nor \U$8925 ( \15231 , \13806 , \13807 , \13808 , \13768 , \13771 , \13775 , \13778 , \15206 , \15207 , \15208 , \15209 , \15210 , \15211 , \15212 , \15213 , \15214 , \15215 , \15216 , \15217 , \15218 , \15219 , \15220 , \15221 , \15222 , \15223 , \15224 , \15225 , \15226 , \15227 , \15228 , \15229 , \15230 );
and \U$8926 ( \15232 , \8841 , \15231 );
buf \U$8927 ( \15233 , \13778 );
buf \U$8928 ( \15234 , \13778 );
buf \U$8929 ( \15235 , \13778 );
buf \U$8930 ( \15236 , \13778 );
buf \U$8931 ( \15237 , \13778 );
buf \U$8932 ( \15238 , \13778 );
buf \U$8933 ( \15239 , \13778 );
buf \U$8934 ( \15240 , \13778 );
buf \U$8935 ( \15241 , \13778 );
buf \U$8936 ( \15242 , \13778 );
buf \U$8937 ( \15243 , \13778 );
buf \U$8938 ( \15244 , \13778 );
buf \U$8939 ( \15245 , \13778 );
buf \U$8940 ( \15246 , \13778 );
buf \U$8941 ( \15247 , \13778 );
buf \U$8942 ( \15248 , \13778 );
buf \U$8943 ( \15249 , \13778 );
buf \U$8944 ( \15250 , \13778 );
buf \U$8945 ( \15251 , \13778 );
buf \U$8946 ( \15252 , \13778 );
buf \U$8947 ( \15253 , \13778 );
buf \U$8948 ( \15254 , \13778 );
buf \U$8949 ( \15255 , \13778 );
buf \U$8950 ( \15256 , \13778 );
buf \U$8951 ( \15257 , \13778 );
nor \U$8952 ( \15258 , \13765 , \13807 , \13808 , \13768 , \13771 , \13775 , \13778 , \15233 , \15234 , \15235 , \15236 , \15237 , \15238 , \15239 , \15240 , \15241 , \15242 , \15243 , \15244 , \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 , \15252 , \15253 , \15254 , \15255 , \15256 , \15257 );
and \U$8953 ( \15259 , \8869 , \15258 );
buf \U$8954 ( \15260 , \13778 );
buf \U$8955 ( \15261 , \13778 );
buf \U$8956 ( \15262 , \13778 );
buf \U$8957 ( \15263 , \13778 );
buf \U$8958 ( \15264 , \13778 );
buf \U$8959 ( \15265 , \13778 );
buf \U$8960 ( \15266 , \13778 );
buf \U$8961 ( \15267 , \13778 );
buf \U$8962 ( \15268 , \13778 );
buf \U$8963 ( \15269 , \13778 );
buf \U$8964 ( \15270 , \13778 );
buf \U$8965 ( \15271 , \13778 );
buf \U$8966 ( \15272 , \13778 );
buf \U$8967 ( \15273 , \13778 );
buf \U$8968 ( \15274 , \13778 );
buf \U$8969 ( \15275 , \13778 );
buf \U$8970 ( \15276 , \13778 );
buf \U$8971 ( \15277 , \13778 );
buf \U$8972 ( \15278 , \13778 );
buf \U$8973 ( \15279 , \13778 );
buf \U$8974 ( \15280 , \13778 );
buf \U$8975 ( \15281 , \13778 );
buf \U$8976 ( \15282 , \13778 );
buf \U$8977 ( \15283 , \13778 );
buf \U$8978 ( \15284 , \13778 );
nor \U$8979 ( \15285 , \13806 , \13766 , \13808 , \13768 , \13771 , \13775 , \13778 , \15260 , \15261 , \15262 , \15263 , \15264 , \15265 , \15266 , \15267 , \15268 , \15269 , \15270 , \15271 , \15272 , \15273 , \15274 , \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 , \15282 , \15283 , \15284 );
and \U$8980 ( \15286 , \8897 , \15285 );
buf \U$8981 ( \15287 , \13778 );
buf \U$8982 ( \15288 , \13778 );
buf \U$8983 ( \15289 , \13778 );
buf \U$8984 ( \15290 , \13778 );
buf \U$8985 ( \15291 , \13778 );
buf \U$8986 ( \15292 , \13778 );
buf \U$8987 ( \15293 , \13778 );
buf \U$8988 ( \15294 , \13778 );
buf \U$8989 ( \15295 , \13778 );
buf \U$8990 ( \15296 , \13778 );
buf \U$8991 ( \15297 , \13778 );
buf \U$8992 ( \15298 , \13778 );
buf \U$8993 ( \15299 , \13778 );
buf \U$8994 ( \15300 , \13778 );
buf \U$8995 ( \15301 , \13778 );
buf \U$8996 ( \15302 , \13778 );
buf \U$8997 ( \15303 , \13778 );
buf \U$8998 ( \15304 , \13778 );
buf \U$8999 ( \15305 , \13778 );
buf \U$9000 ( \15306 , \13778 );
buf \U$9001 ( \15307 , \13778 );
buf \U$9002 ( \15308 , \13778 );
buf \U$9003 ( \15309 , \13778 );
buf \U$9004 ( \15310 , \13778 );
buf \U$9005 ( \15311 , \13778 );
nor \U$9006 ( \15312 , \13765 , \13766 , \13808 , \13768 , \13771 , \13775 , \13778 , \15287 , \15288 , \15289 , \15290 , \15291 , \15292 , \15293 , \15294 , \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 , \15302 , \15303 , \15304 , \15305 , \15306 , \15307 , \15308 , \15309 , \15310 , \15311 );
and \U$9007 ( \15313 , \8925 , \15312 );
buf \U$9008 ( \15314 , \13778 );
buf \U$9009 ( \15315 , \13778 );
buf \U$9010 ( \15316 , \13778 );
buf \U$9011 ( \15317 , \13778 );
buf \U$9012 ( \15318 , \13778 );
buf \U$9013 ( \15319 , \13778 );
buf \U$9014 ( \15320 , \13778 );
buf \U$9015 ( \15321 , \13778 );
buf \U$9016 ( \15322 , \13778 );
buf \U$9017 ( \15323 , \13778 );
buf \U$9018 ( \15324 , \13778 );
buf \U$9019 ( \15325 , \13778 );
buf \U$9020 ( \15326 , \13778 );
buf \U$9021 ( \15327 , \13778 );
buf \U$9022 ( \15328 , \13778 );
buf \U$9023 ( \15329 , \13778 );
buf \U$9024 ( \15330 , \13778 );
buf \U$9025 ( \15331 , \13778 );
buf \U$9026 ( \15332 , \13778 );
buf \U$9027 ( \15333 , \13778 );
buf \U$9028 ( \15334 , \13778 );
buf \U$9029 ( \15335 , \13778 );
buf \U$9030 ( \15336 , \13778 );
buf \U$9031 ( \15337 , \13778 );
buf \U$9032 ( \15338 , \13778 );
nor \U$9033 ( \15339 , \13806 , \13807 , \13767 , \13768 , \13771 , \13775 , \13778 , \15314 , \15315 , \15316 , \15317 , \15318 , \15319 , \15320 , \15321 , \15322 , \15323 , \15324 , \15325 , \15326 , \15327 , \15328 , \15329 , \15330 , \15331 , \15332 , \15333 , \15334 , \15335 , \15336 , \15337 , \15338 );
and \U$9034 ( \15340 , \8953 , \15339 );
buf \U$9035 ( \15341 , \13778 );
buf \U$9036 ( \15342 , \13778 );
buf \U$9037 ( \15343 , \13778 );
buf \U$9038 ( \15344 , \13778 );
buf \U$9039 ( \15345 , \13778 );
buf \U$9040 ( \15346 , \13778 );
buf \U$9041 ( \15347 , \13778 );
buf \U$9042 ( \15348 , \13778 );
buf \U$9043 ( \15349 , \13778 );
buf \U$9044 ( \15350 , \13778 );
buf \U$9045 ( \15351 , \13778 );
buf \U$9046 ( \15352 , \13778 );
buf \U$9047 ( \15353 , \13778 );
buf \U$9048 ( \15354 , \13778 );
buf \U$9049 ( \15355 , \13778 );
buf \U$9050 ( \15356 , \13778 );
buf \U$9051 ( \15357 , \13778 );
buf \U$9052 ( \15358 , \13778 );
buf \U$9053 ( \15359 , \13778 );
buf \U$9054 ( \15360 , \13778 );
buf \U$9055 ( \15361 , \13778 );
buf \U$9056 ( \15362 , \13778 );
buf \U$9057 ( \15363 , \13778 );
buf \U$9058 ( \15364 , \13778 );
buf \U$9059 ( \15365 , \13778 );
nor \U$9060 ( \15366 , \13765 , \13807 , \13767 , \13768 , \13771 , \13775 , \13778 , \15341 , \15342 , \15343 , \15344 , \15345 , \15346 , \15347 , \15348 , \15349 , \15350 , \15351 , \15352 , \15353 , \15354 , \15355 , \15356 , \15357 , \15358 , \15359 , \15360 , \15361 , \15362 , \15363 , \15364 , \15365 );
and \U$9061 ( \15367 , \8981 , \15366 );
buf \U$9062 ( \15368 , \13778 );
buf \U$9063 ( \15369 , \13778 );
buf \U$9064 ( \15370 , \13778 );
buf \U$9065 ( \15371 , \13778 );
buf \U$9066 ( \15372 , \13778 );
buf \U$9067 ( \15373 , \13778 );
buf \U$9068 ( \15374 , \13778 );
buf \U$9069 ( \15375 , \13778 );
buf \U$9070 ( \15376 , \13778 );
buf \U$9071 ( \15377 , \13778 );
buf \U$9072 ( \15378 , \13778 );
buf \U$9073 ( \15379 , \13778 );
buf \U$9074 ( \15380 , \13778 );
buf \U$9075 ( \15381 , \13778 );
buf \U$9076 ( \15382 , \13778 );
buf \U$9077 ( \15383 , \13778 );
buf \U$9078 ( \15384 , \13778 );
buf \U$9079 ( \15385 , \13778 );
buf \U$9080 ( \15386 , \13778 );
buf \U$9081 ( \15387 , \13778 );
buf \U$9082 ( \15388 , \13778 );
buf \U$9083 ( \15389 , \13778 );
buf \U$9084 ( \15390 , \13778 );
buf \U$9085 ( \15391 , \13778 );
buf \U$9086 ( \15392 , \13778 );
nor \U$9087 ( \15393 , \13806 , \13766 , \13767 , \13768 , \13771 , \13775 , \13778 , \15368 , \15369 , \15370 , \15371 , \15372 , \15373 , \15374 , \15375 , \15376 , \15377 , \15378 , \15379 , \15380 , \15381 , \15382 , \15383 , \15384 , \15385 , \15386 , \15387 , \15388 , \15389 , \15390 , \15391 , \15392 );
and \U$9088 ( \15394 , \9009 , \15393 );
or \U$9089 ( \15395 , \14989 , \15016 , \15043 , \15070 , \15097 , \15124 , \15151 , \15178 , \15205 , \15232 , \15259 , \15286 , \15313 , \15340 , \15367 , \15394 );
buf \U$9090 ( \15396 , \13778 );
not \U$9091 ( \15397 , \15396 );
buf \U$9092 ( \15398 , \13766 );
buf \U$9093 ( \15399 , \13767 );
buf \U$9094 ( \15400 , \13768 );
buf \U$9095 ( \15401 , \13771 );
buf \U$9096 ( \15402 , \13775 );
buf \U$9097 ( \15403 , \13778 );
buf \U$9098 ( \15404 , \13778 );
buf \U$9099 ( \15405 , \13778 );
buf \U$9100 ( \15406 , \13778 );
buf \U$9101 ( \15407 , \13778 );
buf \U$9102 ( \15408 , \13778 );
buf \U$9103 ( \15409 , \13778 );
buf \U$9104 ( \15410 , \13778 );
buf \U$9105 ( \15411 , \13778 );
buf \U$9106 ( \15412 , \13778 );
buf \U$9107 ( \15413 , \13778 );
buf \U$9108 ( \15414 , \13778 );
buf \U$9109 ( \15415 , \13778 );
buf \U$9110 ( \15416 , \13778 );
buf \U$9111 ( \15417 , \13778 );
buf \U$9112 ( \15418 , \13778 );
buf \U$9113 ( \15419 , \13778 );
buf \U$9114 ( \15420 , \13778 );
buf \U$9115 ( \15421 , \13778 );
buf \U$9116 ( \15422 , \13778 );
buf \U$9117 ( \15423 , \13778 );
buf \U$9118 ( \15424 , \13778 );
buf \U$9119 ( \15425 , \13778 );
buf \U$9120 ( \15426 , \13778 );
buf \U$9121 ( \15427 , \13778 );
buf \U$9122 ( \15428 , \13765 );
or \U$9123 ( \15429 , \15398 , \15399 , \15400 , \15401 , \15402 , \15403 , \15404 , \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411 , \15412 , \15413 , \15414 , \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 , \15422 , \15423 , \15424 , \15425 , \15426 , \15427 , \15428 );
nand \U$9124 ( \15430 , \15397 , \15429 );
buf \U$9125 ( \15431 , \15430 );
buf \U$9126 ( \15432 , \13778 );
not \U$9127 ( \15433 , \15432 );
buf \U$9128 ( \15434 , \13775 );
buf \U$9129 ( \15435 , \13778 );
buf \U$9130 ( \15436 , \13778 );
buf \U$9131 ( \15437 , \13778 );
buf \U$9132 ( \15438 , \13778 );
buf \U$9133 ( \15439 , \13778 );
buf \U$9134 ( \15440 , \13778 );
buf \U$9135 ( \15441 , \13778 );
buf \U$9136 ( \15442 , \13778 );
buf \U$9137 ( \15443 , \13778 );
buf \U$9138 ( \15444 , \13778 );
buf \U$9139 ( \15445 , \13778 );
buf \U$9140 ( \15446 , \13778 );
buf \U$9141 ( \15447 , \13778 );
buf \U$9142 ( \15448 , \13778 );
buf \U$9143 ( \15449 , \13778 );
buf \U$9144 ( \15450 , \13778 );
buf \U$9145 ( \15451 , \13778 );
buf \U$9146 ( \15452 , \13778 );
buf \U$9147 ( \15453 , \13778 );
buf \U$9148 ( \15454 , \13778 );
buf \U$9149 ( \15455 , \13778 );
buf \U$9150 ( \15456 , \13778 );
buf \U$9151 ( \15457 , \13778 );
buf \U$9152 ( \15458 , \13778 );
buf \U$9153 ( \15459 , \13778 );
buf \U$9154 ( \15460 , \13771 );
buf \U$9155 ( \15461 , \13765 );
buf \U$9156 ( \15462 , \13766 );
buf \U$9157 ( \15463 , \13767 );
buf \U$9158 ( \15464 , \13768 );
or \U$9159 ( \15465 , \15461 , \15462 , \15463 , \15464 );
and \U$9160 ( \15466 , \15460 , \15465 );
or \U$9161 ( \15467 , \15434 , \15435 , \15436 , \15437 , \15438 , \15439 , \15440 , \15441 , \15442 , \15443 , \15444 , \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 , \15452 , \15453 , \15454 , \15455 , \15456 , \15457 , \15458 , \15459 , \15466 );
and \U$9162 ( \15468 , \15433 , \15467 );
buf \U$9163 ( \15469 , \15468 );
or \U$9164 ( \15470 , \15431 , \15469 );
_DC g533b ( \15471_nG533b , \15395 , \15470 );
buf \U$9165 ( \15472 , \15471_nG533b );
xor \U$9166 ( \15473 , \14962 , \15472 );
buf \U$9167 ( \15474 , RIb7af5b8_255);
and \U$9168 ( \15475 , \7207 , \14988 );
and \U$9169 ( \15476 , \7209 , \15015 );
and \U$9170 ( \15477 , \9119 , \15042 );
and \U$9171 ( \15478 , \9121 , \15069 );
and \U$9172 ( \15479 , \9123 , \15096 );
and \U$9173 ( \15480 , \9125 , \15123 );
and \U$9174 ( \15481 , \9127 , \15150 );
and \U$9175 ( \15482 , \9129 , \15177 );
and \U$9176 ( \15483 , \9131 , \15204 );
and \U$9177 ( \15484 , \9133 , \15231 );
and \U$9178 ( \15485 , \9135 , \15258 );
and \U$9179 ( \15486 , \9137 , \15285 );
and \U$9180 ( \15487 , \9139 , \15312 );
and \U$9181 ( \15488 , \9141 , \15339 );
and \U$9182 ( \15489 , \9143 , \15366 );
and \U$9183 ( \15490 , \9145 , \15393 );
or \U$9184 ( \15491 , \15475 , \15476 , \15477 , \15478 , \15479 , \15480 , \15481 , \15482 , \15483 , \15484 , \15485 , \15486 , \15487 , \15488 , \15489 , \15490 );
_DC g5350 ( \15492_nG5350 , \15491 , \15470 );
buf \U$9185 ( \15493 , \15492_nG5350 );
xor \U$9186 ( \15494 , \15474 , \15493 );
or \U$9187 ( \15495 , \15473 , \15494 );
buf \U$9188 ( \15496 , RIb7af540_256);
and \U$9189 ( \15497 , \7217 , \14988 );
and \U$9190 ( \15498 , \7219 , \15015 );
and \U$9191 ( \15499 , \9155 , \15042 );
and \U$9192 ( \15500 , \9157 , \15069 );
and \U$9193 ( \15501 , \9159 , \15096 );
and \U$9194 ( \15502 , \9161 , \15123 );
and \U$9195 ( \15503 , \9163 , \15150 );
and \U$9196 ( \15504 , \9165 , \15177 );
and \U$9197 ( \15505 , \9167 , \15204 );
and \U$9198 ( \15506 , \9169 , \15231 );
and \U$9199 ( \15507 , \9171 , \15258 );
and \U$9200 ( \15508 , \9173 , \15285 );
and \U$9201 ( \15509 , \9175 , \15312 );
and \U$9202 ( \15510 , \9177 , \15339 );
and \U$9203 ( \15511 , \9179 , \15366 );
and \U$9204 ( \15512 , \9181 , \15393 );
or \U$9205 ( \15513 , \15497 , \15498 , \15499 , \15500 , \15501 , \15502 , \15503 , \15504 , \15505 , \15506 , \15507 , \15508 , \15509 , \15510 , \15511 , \15512 );
_DC g5366 ( \15514_nG5366 , \15513 , \15470 );
buf \U$9206 ( \15515 , \15514_nG5366 );
xor \U$9207 ( \15516 , \15496 , \15515 );
or \U$9208 ( \15517 , \15495 , \15516 );
buf \U$9209 ( \15518 , RIb7af4c8_257);
and \U$9210 ( \15519 , \7227 , \14988 );
and \U$9211 ( \15520 , \7229 , \15015 );
and \U$9212 ( \15521 , \9191 , \15042 );
and \U$9213 ( \15522 , \9193 , \15069 );
and \U$9214 ( \15523 , \9195 , \15096 );
and \U$9215 ( \15524 , \9197 , \15123 );
and \U$9216 ( \15525 , \9199 , \15150 );
and \U$9217 ( \15526 , \9201 , \15177 );
and \U$9218 ( \15527 , \9203 , \15204 );
and \U$9219 ( \15528 , \9205 , \15231 );
and \U$9220 ( \15529 , \9207 , \15258 );
and \U$9221 ( \15530 , \9209 , \15285 );
and \U$9222 ( \15531 , \9211 , \15312 );
and \U$9223 ( \15532 , \9213 , \15339 );
and \U$9224 ( \15533 , \9215 , \15366 );
and \U$9225 ( \15534 , \9217 , \15393 );
or \U$9226 ( \15535 , \15519 , \15520 , \15521 , \15522 , \15523 , \15524 , \15525 , \15526 , \15527 , \15528 , \15529 , \15530 , \15531 , \15532 , \15533 , \15534 );
_DC g537c ( \15536_nG537c , \15535 , \15470 );
buf \U$9227 ( \15537 , \15536_nG537c );
xor \U$9228 ( \15538 , \15518 , \15537 );
or \U$9229 ( \15539 , \15517 , \15538 );
buf \U$9230 ( \15540 , RIb7af450_258);
and \U$9231 ( \15541 , \7237 , \14988 );
and \U$9232 ( \15542 , \7239 , \15015 );
and \U$9233 ( \15543 , \9227 , \15042 );
and \U$9234 ( \15544 , \9229 , \15069 );
and \U$9235 ( \15545 , \9231 , \15096 );
and \U$9236 ( \15546 , \9233 , \15123 );
and \U$9237 ( \15547 , \9235 , \15150 );
and \U$9238 ( \15548 , \9237 , \15177 );
and \U$9239 ( \15549 , \9239 , \15204 );
and \U$9240 ( \15550 , \9241 , \15231 );
and \U$9241 ( \15551 , \9243 , \15258 );
and \U$9242 ( \15552 , \9245 , \15285 );
and \U$9243 ( \15553 , \9247 , \15312 );
and \U$9244 ( \15554 , \9249 , \15339 );
and \U$9245 ( \15555 , \9251 , \15366 );
and \U$9246 ( \15556 , \9253 , \15393 );
or \U$9247 ( \15557 , \15541 , \15542 , \15543 , \15544 , \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 , \15552 , \15553 , \15554 , \15555 , \15556 );
_DC g5392 ( \15558_nG5392 , \15557 , \15470 );
buf \U$9248 ( \15559 , \15558_nG5392 );
xor \U$9249 ( \15560 , \15540 , \15559 );
or \U$9250 ( \15561 , \15539 , \15560 );
buf \U$9251 ( \15562 , RIb7af3d8_259);
and \U$9252 ( \15563 , \7247 , \14988 );
and \U$9253 ( \15564 , \7249 , \15015 );
and \U$9254 ( \15565 , \9263 , \15042 );
and \U$9255 ( \15566 , \9265 , \15069 );
and \U$9256 ( \15567 , \9267 , \15096 );
and \U$9257 ( \15568 , \9269 , \15123 );
and \U$9258 ( \15569 , \9271 , \15150 );
and \U$9259 ( \15570 , \9273 , \15177 );
and \U$9260 ( \15571 , \9275 , \15204 );
and \U$9261 ( \15572 , \9277 , \15231 );
and \U$9262 ( \15573 , \9279 , \15258 );
and \U$9263 ( \15574 , \9281 , \15285 );
and \U$9264 ( \15575 , \9283 , \15312 );
and \U$9265 ( \15576 , \9285 , \15339 );
and \U$9266 ( \15577 , \9287 , \15366 );
and \U$9267 ( \15578 , \9289 , \15393 );
or \U$9268 ( \15579 , \15563 , \15564 , \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 , \15572 , \15573 , \15574 , \15575 , \15576 , \15577 , \15578 );
_DC g53a8 ( \15580_nG53a8 , \15579 , \15470 );
buf \U$9269 ( \15581 , \15580_nG53a8 );
xor \U$9270 ( \15582 , \15562 , \15581 );
or \U$9271 ( \15583 , \15561 , \15582 );
buf \U$9272 ( \15584 , RIb7a5bf8_260);
and \U$9273 ( \15585 , \7257 , \14988 );
and \U$9274 ( \15586 , \7259 , \15015 );
and \U$9275 ( \15587 , \9299 , \15042 );
and \U$9276 ( \15588 , \9301 , \15069 );
and \U$9277 ( \15589 , \9303 , \15096 );
and \U$9278 ( \15590 , \9305 , \15123 );
and \U$9279 ( \15591 , \9307 , \15150 );
and \U$9280 ( \15592 , \9309 , \15177 );
and \U$9281 ( \15593 , \9311 , \15204 );
and \U$9282 ( \15594 , \9313 , \15231 );
and \U$9283 ( \15595 , \9315 , \15258 );
and \U$9284 ( \15596 , \9317 , \15285 );
and \U$9285 ( \15597 , \9319 , \15312 );
and \U$9286 ( \15598 , \9321 , \15339 );
and \U$9287 ( \15599 , \9323 , \15366 );
and \U$9288 ( \15600 , \9325 , \15393 );
or \U$9289 ( \15601 , \15585 , \15586 , \15587 , \15588 , \15589 , \15590 , \15591 , \15592 , \15593 , \15594 , \15595 , \15596 , \15597 , \15598 , \15599 , \15600 );
_DC g53be ( \15602_nG53be , \15601 , \15470 );
buf \U$9290 ( \15603 , \15602_nG53be );
xor \U$9291 ( \15604 , \15584 , \15603 );
or \U$9292 ( \15605 , \15583 , \15604 );
buf \U$9293 ( \15606 , RIb7a0c48_261);
and \U$9294 ( \15607 , \7267 , \14988 );
and \U$9295 ( \15608 , \7269 , \15015 );
and \U$9296 ( \15609 , \9335 , \15042 );
and \U$9297 ( \15610 , \9337 , \15069 );
and \U$9298 ( \15611 , \9339 , \15096 );
and \U$9299 ( \15612 , \9341 , \15123 );
and \U$9300 ( \15613 , \9343 , \15150 );
and \U$9301 ( \15614 , \9345 , \15177 );
and \U$9302 ( \15615 , \9347 , \15204 );
and \U$9303 ( \15616 , \9349 , \15231 );
and \U$9304 ( \15617 , \9351 , \15258 );
and \U$9305 ( \15618 , \9353 , \15285 );
and \U$9306 ( \15619 , \9355 , \15312 );
and \U$9307 ( \15620 , \9357 , \15339 );
and \U$9308 ( \15621 , \9359 , \15366 );
and \U$9309 ( \15622 , \9361 , \15393 );
or \U$9310 ( \15623 , \15607 , \15608 , \15609 , \15610 , \15611 , \15612 , \15613 , \15614 , \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 , \15622 );
_DC g53d4 ( \15624_nG53d4 , \15623 , \15470 );
buf \U$9311 ( \15625 , \15624_nG53d4 );
xor \U$9312 ( \15626 , \15606 , \15625 );
or \U$9313 ( \15627 , \15605 , \15626 );
not \U$9314 ( \15628 , \15627 );
buf \U$9315 ( \15629 , \15628 );
and \U$9316 ( \15630 , \14961 , \15629 );
_HMUX g53db ( \15631_nG53db , \13539_nG4ba5 , \13765 , \15630 );
buf \U$9317 ( \15632 , \13556 );
buf \U$9318 ( \15633 , \13553 );
buf \U$9319 ( \15634 , \13541 );
buf \U$9320 ( \15635 , \13543 );
buf \U$9321 ( \15636 , \13546 );
buf \U$9322 ( \15637 , \13549 );
or \U$9323 ( \15638 , \15634 , \15635 , \15636 , \15637 );
and \U$9324 ( \15639 , \15633 , \15638 );
or \U$9325 ( \15640 , \15632 , \15639 );
buf \U$9326 ( \15641 , \15640 );
_HMUX g53e6 ( \15642_nG53e6 , \13764_nG4c88 , \15631_nG53db , \15641 );
buf \U$9327 ( \15643 , RIe5319e0_6884);
not \U$9328 ( \15644 , \15643 );
buf \U$9329 ( \15645 , \15644 );
buf \U$9330 ( \15646 , RIe549ef0_6842);
xnor \U$9331 ( \15647 , \15646 , \15643 );
buf \U$9332 ( \15648 , \15647 );
buf \U$9333 ( \15649 , RIe549770_6843);
or \U$9334 ( \15650 , \15646 , \15643 );
xor \U$9335 ( \15651 , \15649 , \15650 );
buf \U$9336 ( \15652 , \15651 );
buf \U$9337 ( \15653 , RIe548ff0_6844);
and \U$9338 ( \15654 , \15649 , \15650 );
xnor \U$9339 ( \15655 , \15653 , \15654 );
buf \U$9340 ( \15656 , \15655 );
buf \U$9341 ( \15657 , RIea91330_6888);
or \U$9342 ( \15658 , \15653 , \15654 );
xor \U$9343 ( \15659 , \15657 , \15658 );
buf \U$9344 ( \15660 , \15659 );
not \U$9345 ( \15661 , \15660 );
and \U$9346 ( \15662 , \15657 , \15658 );
buf \U$9347 ( \15663 , \15662 );
nor \U$9348 ( \15664 , \15645 , \15648 , \15652 , \15656 , \15661 , \15663 );
and \U$9349 ( \15665 , RIe5329d0_6883, \15664 );
not \U$9350 ( \15666 , \15663 );
and \U$9351 ( \15667 , \15645 , \15648 , \15652 , \15656 , \15661 , \15666 );
and \U$9352 ( \15668 , RIeb72150_6905, \15667 );
not \U$9353 ( \15669 , \15645 );
and \U$9354 ( \15670 , \15669 , \15648 , \15652 , \15656 , \15661 , \15666 );
and \U$9355 ( \15671 , RIeab80c0_6897, \15670 );
not \U$9356 ( \15672 , \15648 );
and \U$9357 ( \15673 , \15645 , \15672 , \15652 , \15656 , \15661 , \15666 );
and \U$9358 ( \15674 , RIe5331c8_6882, \15673 );
and \U$9359 ( \15675 , \15669 , \15672 , \15652 , \15656 , \15661 , \15666 );
and \U$9360 ( \15676 , RIe5339c0_6881, \15675 );
not \U$9361 ( \15677 , \15652 );
and \U$9362 ( \15678 , \15645 , \15648 , \15677 , \15656 , \15661 , \15666 );
and \U$9363 ( \15679 , RIeab87c8_6898, \15678 );
or \U$9374 ( \15680 , \15665 , \15668 , \15671 , \15674 , \15676 , \15679 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
buf \U$9376 ( \15681 , \15663 );
buf \U$9377 ( \15682 , \15660 );
buf \U$9378 ( \15683 , \15645 );
buf \U$9379 ( \15684 , \15648 );
buf \U$9380 ( \15685 , \15652 );
buf \U$9381 ( \15686 , \15656 );
or \U$9382 ( \15687 , \15683 , \15684 , \15685 , \15686 );
and \U$9383 ( \15688 , \15682 , \15687 );
or \U$9384 ( \15689 , \15681 , \15688 );
buf \U$9385 ( \15690 , \15689 );
or \U$9386 ( \15691 , 1'b0 , \15690 );
_DC g5418 ( \15692_nG5418 , \15680 , \15691 );
not \U$9387 ( \15693 , \15692_nG5418 );
buf \U$9388 ( \15694 , RIb7b9608_246);
and \U$9389 ( \15695 , \7117 , \15664 );
and \U$9390 ( \15696 , \7119 , \15667 );
and \U$9391 ( \15697 , \7864 , \15670 );
and \U$9392 ( \15698 , \7892 , \15673 );
and \U$9393 ( \15699 , \7920 , \15675 );
and \U$9394 ( \15700 , \7948 , \15678 );
or \U$9405 ( \15701 , \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5422 ( \15702_nG5422 , \15701 , \15691 );
buf \U$9406 ( \15703 , \15702_nG5422 );
xor \U$9407 ( \15704 , \15694 , \15703 );
buf \U$9408 ( \15705 , RIb7b9590_247);
and \U$9409 ( \15706 , \7126 , \15664 );
and \U$9410 ( \15707 , \7128 , \15667 );
and \U$9411 ( \15708 , \8338 , \15670 );
and \U$9412 ( \15709 , \8340 , \15673 );
and \U$9413 ( \15710 , \8342 , \15675 );
and \U$9414 ( \15711 , \8344 , \15678 );
or \U$9425 ( \15712 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g542d ( \15713_nG542d , \15712 , \15691 );
buf \U$9426 ( \15714 , \15713_nG542d );
xor \U$9427 ( \15715 , \15705 , \15714 );
or \U$9428 ( \15716 , \15704 , \15715 );
buf \U$9429 ( \15717 , RIb7b9518_248);
and \U$9430 ( \15718 , \7136 , \15664 );
and \U$9431 ( \15719 , \7138 , \15667 );
and \U$9432 ( \15720 , \8374 , \15670 );
and \U$9433 ( \15721 , \8376 , \15673 );
and \U$9434 ( \15722 , \8378 , \15675 );
and \U$9435 ( \15723 , \8380 , \15678 );
or \U$9446 ( \15724 , \15718 , \15719 , \15720 , \15721 , \15722 , \15723 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5439 ( \15725_nG5439 , \15724 , \15691 );
buf \U$9447 ( \15726 , \15725_nG5439 );
xor \U$9448 ( \15727 , \15717 , \15726 );
or \U$9449 ( \15728 , \15716 , \15727 );
buf \U$9450 ( \15729 , RIb7b94a0_249);
and \U$9451 ( \15730 , \7146 , \15664 );
and \U$9452 ( \15731 , \7148 , \15667 );
and \U$9453 ( \15732 , \8410 , \15670 );
and \U$9454 ( \15733 , \8412 , \15673 );
and \U$9455 ( \15734 , \8414 , \15675 );
and \U$9456 ( \15735 , \8416 , \15678 );
or \U$9467 ( \15736 , \15730 , \15731 , \15732 , \15733 , \15734 , \15735 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5445 ( \15737_nG5445 , \15736 , \15691 );
buf \U$9468 ( \15738 , \15737_nG5445 );
xor \U$9469 ( \15739 , \15729 , \15738 );
or \U$9470 ( \15740 , \15728 , \15739 );
buf \U$9471 ( \15741 , RIb7b9428_250);
and \U$9472 ( \15742 , \7156 , \15664 );
and \U$9473 ( \15743 , \7158 , \15667 );
and \U$9474 ( \15744 , \8446 , \15670 );
and \U$9475 ( \15745 , \8448 , \15673 );
and \U$9476 ( \15746 , \8450 , \15675 );
and \U$9477 ( \15747 , \8452 , \15678 );
or \U$9488 ( \15748 , \15742 , \15743 , \15744 , \15745 , \15746 , \15747 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5451 ( \15749_nG5451 , \15748 , \15691 );
buf \U$9489 ( \15750 , \15749_nG5451 );
xor \U$9490 ( \15751 , \15741 , \15750 );
or \U$9491 ( \15752 , \15740 , \15751 );
buf \U$9492 ( \15753 , RIb7b93b0_251);
and \U$9493 ( \15754 , \7166 , \15664 );
and \U$9494 ( \15755 , \7168 , \15667 );
and \U$9495 ( \15756 , \8482 , \15670 );
and \U$9496 ( \15757 , \8484 , \15673 );
and \U$9497 ( \15758 , \8486 , \15675 );
and \U$9498 ( \15759 , \8488 , \15678 );
or \U$9509 ( \15760 , \15754 , \15755 , \15756 , \15757 , \15758 , \15759 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g545d ( \15761_nG545d , \15760 , \15691 );
buf \U$9510 ( \15762 , \15761_nG545d );
xor \U$9511 ( \15763 , \15753 , \15762 );
or \U$9512 ( \15764 , \15752 , \15763 );
buf \U$9513 ( \15765 , RIb7af720_252);
and \U$9514 ( \15766 , \7176 , \15664 );
and \U$9515 ( \15767 , \7178 , \15667 );
and \U$9516 ( \15768 , \8518 , \15670 );
and \U$9517 ( \15769 , \8520 , \15673 );
and \U$9518 ( \15770 , \8522 , \15675 );
and \U$9519 ( \15771 , \8524 , \15678 );
or \U$9530 ( \15772 , \15766 , \15767 , \15768 , \15769 , \15770 , \15771 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5469 ( \15773_nG5469 , \15772 , \15691 );
buf \U$9531 ( \15774 , \15773_nG5469 );
xor \U$9532 ( \15775 , \15765 , \15774 );
or \U$9533 ( \15776 , \15764 , \15775 );
buf \U$9534 ( \15777 , RIb7af6a8_253);
and \U$9535 ( \15778 , \7186 , \15664 );
and \U$9536 ( \15779 , \7188 , \15667 );
and \U$9537 ( \15780 , \8554 , \15670 );
and \U$9538 ( \15781 , \8556 , \15673 );
and \U$9539 ( \15782 , \8558 , \15675 );
and \U$9540 ( \15783 , \8560 , \15678 );
or \U$9551 ( \15784 , \15778 , \15779 , \15780 , \15781 , \15782 , \15783 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5475 ( \15785_nG5475 , \15784 , \15691 );
buf \U$9552 ( \15786 , \15785_nG5475 );
xor \U$9553 ( \15787 , \15777 , \15786 );
or \U$9554 ( \15788 , \15776 , \15787 );
not \U$9555 ( \15789 , \15788 );
buf \U$9556 ( \15790 , \15789 );
buf \U$9557 ( \15791 , RIb7af630_254);
and \U$9558 ( \15792 , \7198 , \15664 );
and \U$9559 ( \15793 , \7200 , \15667 );
and \U$9560 ( \15794 , \8645 , \15670 );
and \U$9561 ( \15795 , \8673 , \15673 );
and \U$9562 ( \15796 , \8701 , \15675 );
and \U$9563 ( \15797 , \8729 , \15678 );
or \U$9574 ( \15798 , \15792 , \15793 , \15794 , \15795 , \15796 , \15797 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5483 ( \15799_nG5483 , \15798 , \15691 );
buf \U$9575 ( \15800 , \15799_nG5483 );
xor \U$9576 ( \15801 , \15791 , \15800 );
buf \U$9577 ( \15802 , RIb7af5b8_255);
and \U$9578 ( \15803 , \7207 , \15664 );
and \U$9579 ( \15804 , \7209 , \15667 );
and \U$9580 ( \15805 , \9119 , \15670 );
and \U$9581 ( \15806 , \9121 , \15673 );
and \U$9582 ( \15807 , \9123 , \15675 );
and \U$9583 ( \15808 , \9125 , \15678 );
or \U$9594 ( \15809 , \15803 , \15804 , \15805 , \15806 , \15807 , \15808 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g548e ( \15810_nG548e , \15809 , \15691 );
buf \U$9595 ( \15811 , \15810_nG548e );
xor \U$9596 ( \15812 , \15802 , \15811 );
or \U$9597 ( \15813 , \15801 , \15812 );
buf \U$9598 ( \15814 , RIb7af540_256);
and \U$9599 ( \15815 , \7217 , \15664 );
and \U$9600 ( \15816 , \7219 , \15667 );
and \U$9601 ( \15817 , \9155 , \15670 );
and \U$9602 ( \15818 , \9157 , \15673 );
and \U$9603 ( \15819 , \9159 , \15675 );
and \U$9604 ( \15820 , \9161 , \15678 );
or \U$9615 ( \15821 , \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g549a ( \15822_nG549a , \15821 , \15691 );
buf \U$9616 ( \15823 , \15822_nG549a );
xor \U$9617 ( \15824 , \15814 , \15823 );
or \U$9618 ( \15825 , \15813 , \15824 );
buf \U$9619 ( \15826 , RIb7af4c8_257);
and \U$9620 ( \15827 , \7227 , \15664 );
and \U$9621 ( \15828 , \7229 , \15667 );
and \U$9622 ( \15829 , \9191 , \15670 );
and \U$9623 ( \15830 , \9193 , \15673 );
and \U$9624 ( \15831 , \9195 , \15675 );
and \U$9625 ( \15832 , \9197 , \15678 );
or \U$9636 ( \15833 , \15827 , \15828 , \15829 , \15830 , \15831 , \15832 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g54a6 ( \15834_nG54a6 , \15833 , \15691 );
buf \U$9637 ( \15835 , \15834_nG54a6 );
xor \U$9638 ( \15836 , \15826 , \15835 );
or \U$9639 ( \15837 , \15825 , \15836 );
buf \U$9640 ( \15838 , RIb7af450_258);
and \U$9641 ( \15839 , \7237 , \15664 );
and \U$9642 ( \15840 , \7239 , \15667 );
and \U$9643 ( \15841 , \9227 , \15670 );
and \U$9644 ( \15842 , \9229 , \15673 );
and \U$9645 ( \15843 , \9231 , \15675 );
and \U$9646 ( \15844 , \9233 , \15678 );
or \U$9657 ( \15845 , \15839 , \15840 , \15841 , \15842 , \15843 , \15844 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g54b2 ( \15846_nG54b2 , \15845 , \15691 );
buf \U$9658 ( \15847 , \15846_nG54b2 );
xor \U$9659 ( \15848 , \15838 , \15847 );
or \U$9660 ( \15849 , \15837 , \15848 );
buf \U$9661 ( \15850 , RIb7af3d8_259);
and \U$9662 ( \15851 , \7247 , \15664 );
and \U$9663 ( \15852 , \7249 , \15667 );
and \U$9664 ( \15853 , \9263 , \15670 );
and \U$9665 ( \15854 , \9265 , \15673 );
and \U$9666 ( \15855 , \9267 , \15675 );
and \U$9667 ( \15856 , \9269 , \15678 );
or \U$9678 ( \15857 , \15851 , \15852 , \15853 , \15854 , \15855 , \15856 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g54be ( \15858_nG54be , \15857 , \15691 );
buf \U$9679 ( \15859 , \15858_nG54be );
xor \U$9680 ( \15860 , \15850 , \15859 );
or \U$9681 ( \15861 , \15849 , \15860 );
buf \U$9682 ( \15862 , RIb7a5bf8_260);
and \U$9683 ( \15863 , \7257 , \15664 );
and \U$9684 ( \15864 , \7259 , \15667 );
and \U$9685 ( \15865 , \9299 , \15670 );
and \U$9686 ( \15866 , \9301 , \15673 );
and \U$9687 ( \15867 , \9303 , \15675 );
and \U$9688 ( \15868 , \9305 , \15678 );
or \U$9699 ( \15869 , \15863 , \15864 , \15865 , \15866 , \15867 , \15868 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g54ca ( \15870_nG54ca , \15869 , \15691 );
buf \U$9700 ( \15871 , \15870_nG54ca );
xor \U$9701 ( \15872 , \15862 , \15871 );
or \U$9702 ( \15873 , \15861 , \15872 );
buf \U$9703 ( \15874 , RIb7a0c48_261);
and \U$9704 ( \15875 , \7267 , \15664 );
and \U$9705 ( \15876 , \7269 , \15667 );
and \U$9706 ( \15877 , \9335 , \15670 );
and \U$9707 ( \15878 , \9337 , \15673 );
and \U$9708 ( \15879 , \9339 , \15675 );
and \U$9709 ( \15880 , \9341 , \15678 );
or \U$9720 ( \15881 , \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g54d6 ( \15882_nG54d6 , \15881 , \15691 );
buf \U$9721 ( \15883 , \15882_nG54d6 );
xor \U$9722 ( \15884 , \15874 , \15883 );
or \U$9723 ( \15885 , \15873 , \15884 );
not \U$9724 ( \15886 , \15885 );
buf \U$9725 ( \15887 , \15886 );
and \U$9726 ( \15888 , \15790 , \15887 );
and \U$9727 ( \15889 , \15693 , \15888 );
_HMUX g54de ( \15890_nG54de , \15642_nG53e6 , \15645 , \15889 );
buf \U$9730 ( \15891 , \15645 );
buf \U$9733 ( \15892 , \15648 );
buf \U$9736 ( \15893 , \15652 );
buf \U$9739 ( \15894 , \15656 );
buf \U$9740 ( \15895 , \15660 );
not \U$9741 ( \15896 , \15895 );
buf \U$9742 ( \15897 , \15896 );
not \U$9743 ( \15898 , \15897 );
buf \U$9744 ( \15899 , \15663 );
xnor \U$9745 ( \15900 , \15899 , \15895 );
buf \U$9746 ( \15901 , \15900 );
or \U$9747 ( \15902 , \15899 , \15895 );
not \U$9748 ( \15903 , \15902 );
buf \U$9749 ( \15904 , \15903 );
buf \U$9750 ( \15905 , \15904 );
buf \U$9751 ( \15906 , \15904 );
buf \U$9752 ( \15907 , \15904 );
buf \U$9753 ( \15908 , \15904 );
buf \U$9754 ( \15909 , \15904 );
buf \U$9755 ( \15910 , \15904 );
buf \U$9756 ( \15911 , \15904 );
buf \U$9757 ( \15912 , \15904 );
buf \U$9758 ( \15913 , \15904 );
buf \U$9759 ( \15914 , \15904 );
buf \U$9760 ( \15915 , \15904 );
buf \U$9761 ( \15916 , \15904 );
buf \U$9762 ( \15917 , \15904 );
buf \U$9763 ( \15918 , \15904 );
buf \U$9764 ( \15919 , \15904 );
buf \U$9765 ( \15920 , \15904 );
buf \U$9766 ( \15921 , \15904 );
buf \U$9767 ( \15922 , \15904 );
buf \U$9768 ( \15923 , \15904 );
buf \U$9769 ( \15924 , \15904 );
buf \U$9770 ( \15925 , \15904 );
buf \U$9771 ( \15926 , \15904 );
buf \U$9772 ( \15927 , \15904 );
buf \U$9773 ( \15928 , \15904 );
buf \U$9774 ( \15929 , \15904 );
nor \U$9775 ( \15930 , \15891 , \15892 , \15893 , \15894 , \15898 , \15901 , \15904 , \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 , \15912 , \15913 , \15914 , \15915 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 , \15922 , \15923 , \15924 , \15925 , \15926 , \15927 , \15928 , \15929 );
and \U$9776 ( \15931 , RIe5329d0_6883, \15930 );
not \U$9777 ( \15932 , \15891 );
not \U$9778 ( \15933 , \15892 );
not \U$9779 ( \15934 , \15893 );
not \U$9780 ( \15935 , \15894 );
buf \U$9781 ( \15936 , \15904 );
buf \U$9782 ( \15937 , \15904 );
buf \U$9783 ( \15938 , \15904 );
buf \U$9784 ( \15939 , \15904 );
buf \U$9785 ( \15940 , \15904 );
buf \U$9786 ( \15941 , \15904 );
buf \U$9787 ( \15942 , \15904 );
buf \U$9788 ( \15943 , \15904 );
buf \U$9789 ( \15944 , \15904 );
buf \U$9790 ( \15945 , \15904 );
buf \U$9791 ( \15946 , \15904 );
buf \U$9792 ( \15947 , \15904 );
buf \U$9793 ( \15948 , \15904 );
buf \U$9794 ( \15949 , \15904 );
buf \U$9795 ( \15950 , \15904 );
buf \U$9796 ( \15951 , \15904 );
buf \U$9797 ( \15952 , \15904 );
buf \U$9798 ( \15953 , \15904 );
buf \U$9799 ( \15954 , \15904 );
buf \U$9800 ( \15955 , \15904 );
buf \U$9801 ( \15956 , \15904 );
buf \U$9802 ( \15957 , \15904 );
buf \U$9803 ( \15958 , \15904 );
buf \U$9804 ( \15959 , \15904 );
buf \U$9805 ( \15960 , \15904 );
nor \U$9806 ( \15961 , \15932 , \15933 , \15934 , \15935 , \15897 , \15901 , \15904 , \15936 , \15937 , \15938 , \15939 , \15940 , \15941 , \15942 , \15943 , \15944 , \15945 , \15946 , \15947 , \15948 , \15949 , \15950 , \15951 , \15952 , \15953 , \15954 , \15955 , \15956 , \15957 , \15958 , \15959 , \15960 );
and \U$9807 ( \15962 , RIeb72150_6905, \15961 );
buf \U$9808 ( \15963 , \15904 );
buf \U$9809 ( \15964 , \15904 );
buf \U$9810 ( \15965 , \15904 );
buf \U$9811 ( \15966 , \15904 );
buf \U$9812 ( \15967 , \15904 );
buf \U$9813 ( \15968 , \15904 );
buf \U$9814 ( \15969 , \15904 );
buf \U$9815 ( \15970 , \15904 );
buf \U$9816 ( \15971 , \15904 );
buf \U$9817 ( \15972 , \15904 );
buf \U$9818 ( \15973 , \15904 );
buf \U$9819 ( \15974 , \15904 );
buf \U$9820 ( \15975 , \15904 );
buf \U$9821 ( \15976 , \15904 );
buf \U$9822 ( \15977 , \15904 );
buf \U$9823 ( \15978 , \15904 );
buf \U$9824 ( \15979 , \15904 );
buf \U$9825 ( \15980 , \15904 );
buf \U$9826 ( \15981 , \15904 );
buf \U$9827 ( \15982 , \15904 );
buf \U$9828 ( \15983 , \15904 );
buf \U$9829 ( \15984 , \15904 );
buf \U$9830 ( \15985 , \15904 );
buf \U$9831 ( \15986 , \15904 );
buf \U$9832 ( \15987 , \15904 );
nor \U$9833 ( \15988 , \15891 , \15933 , \15934 , \15935 , \15897 , \15901 , \15904 , \15963 , \15964 , \15965 , \15966 , \15967 , \15968 , \15969 , \15970 , \15971 , \15972 , \15973 , \15974 , \15975 , \15976 , \15977 , \15978 , \15979 , \15980 , \15981 , \15982 , \15983 , \15984 , \15985 , \15986 , \15987 );
and \U$9834 ( \15989 , RIeab80c0_6897, \15988 );
buf \U$9835 ( \15990 , \15904 );
buf \U$9836 ( \15991 , \15904 );
buf \U$9837 ( \15992 , \15904 );
buf \U$9838 ( \15993 , \15904 );
buf \U$9839 ( \15994 , \15904 );
buf \U$9840 ( \15995 , \15904 );
buf \U$9841 ( \15996 , \15904 );
buf \U$9842 ( \15997 , \15904 );
buf \U$9843 ( \15998 , \15904 );
buf \U$9844 ( \15999 , \15904 );
buf \U$9845 ( \16000 , \15904 );
buf \U$9846 ( \16001 , \15904 );
buf \U$9847 ( \16002 , \15904 );
buf \U$9848 ( \16003 , \15904 );
buf \U$9849 ( \16004 , \15904 );
buf \U$9850 ( \16005 , \15904 );
buf \U$9851 ( \16006 , \15904 );
buf \U$9852 ( \16007 , \15904 );
buf \U$9853 ( \16008 , \15904 );
buf \U$9854 ( \16009 , \15904 );
buf \U$9855 ( \16010 , \15904 );
buf \U$9856 ( \16011 , \15904 );
buf \U$9857 ( \16012 , \15904 );
buf \U$9858 ( \16013 , \15904 );
buf \U$9859 ( \16014 , \15904 );
nor \U$9860 ( \16015 , \15932 , \15892 , \15934 , \15935 , \15897 , \15901 , \15904 , \15990 , \15991 , \15992 , \15993 , \15994 , \15995 , \15996 , \15997 , \15998 , \15999 , \16000 , \16001 , \16002 , \16003 , \16004 , \16005 , \16006 , \16007 , \16008 , \16009 , \16010 , \16011 , \16012 , \16013 , \16014 );
and \U$9861 ( \16016 , RIe5331c8_6882, \16015 );
buf \U$9862 ( \16017 , \15904 );
buf \U$9863 ( \16018 , \15904 );
buf \U$9864 ( \16019 , \15904 );
buf \U$9865 ( \16020 , \15904 );
buf \U$9866 ( \16021 , \15904 );
buf \U$9867 ( \16022 , \15904 );
buf \U$9868 ( \16023 , \15904 );
buf \U$9869 ( \16024 , \15904 );
buf \U$9870 ( \16025 , \15904 );
buf \U$9871 ( \16026 , \15904 );
buf \U$9872 ( \16027 , \15904 );
buf \U$9873 ( \16028 , \15904 );
buf \U$9874 ( \16029 , \15904 );
buf \U$9875 ( \16030 , \15904 );
buf \U$9876 ( \16031 , \15904 );
buf \U$9877 ( \16032 , \15904 );
buf \U$9878 ( \16033 , \15904 );
buf \U$9879 ( \16034 , \15904 );
buf \U$9880 ( \16035 , \15904 );
buf \U$9881 ( \16036 , \15904 );
buf \U$9882 ( \16037 , \15904 );
buf \U$9883 ( \16038 , \15904 );
buf \U$9884 ( \16039 , \15904 );
buf \U$9885 ( \16040 , \15904 );
buf \U$9886 ( \16041 , \15904 );
nor \U$9887 ( \16042 , \15891 , \15892 , \15934 , \15935 , \15897 , \15901 , \15904 , \16017 , \16018 , \16019 , \16020 , \16021 , \16022 , \16023 , \16024 , \16025 , \16026 , \16027 , \16028 , \16029 , \16030 , \16031 , \16032 , \16033 , \16034 , \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 );
and \U$9888 ( \16043 , RIe5339c0_6881, \16042 );
buf \U$9889 ( \16044 , \15904 );
buf \U$9890 ( \16045 , \15904 );
buf \U$9891 ( \16046 , \15904 );
buf \U$9892 ( \16047 , \15904 );
buf \U$9893 ( \16048 , \15904 );
buf \U$9894 ( \16049 , \15904 );
buf \U$9895 ( \16050 , \15904 );
buf \U$9896 ( \16051 , \15904 );
buf \U$9897 ( \16052 , \15904 );
buf \U$9898 ( \16053 , \15904 );
buf \U$9899 ( \16054 , \15904 );
buf \U$9900 ( \16055 , \15904 );
buf \U$9901 ( \16056 , \15904 );
buf \U$9902 ( \16057 , \15904 );
buf \U$9903 ( \16058 , \15904 );
buf \U$9904 ( \16059 , \15904 );
buf \U$9905 ( \16060 , \15904 );
buf \U$9906 ( \16061 , \15904 );
buf \U$9907 ( \16062 , \15904 );
buf \U$9908 ( \16063 , \15904 );
buf \U$9909 ( \16064 , \15904 );
buf \U$9910 ( \16065 , \15904 );
buf \U$9911 ( \16066 , \15904 );
buf \U$9912 ( \16067 , \15904 );
buf \U$9913 ( \16068 , \15904 );
nor \U$9914 ( \16069 , \15932 , \15933 , \15893 , \15935 , \15897 , \15901 , \15904 , \16044 , \16045 , \16046 , \16047 , \16048 , \16049 , \16050 , \16051 , \16052 , \16053 , \16054 , \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 , \16062 , \16063 , \16064 , \16065 , \16066 , \16067 , \16068 );
and \U$9915 ( \16070 , RIeab87c8_6898, \16069 );
buf \U$9916 ( \16071 , \15904 );
buf \U$9917 ( \16072 , \15904 );
buf \U$9918 ( \16073 , \15904 );
buf \U$9919 ( \16074 , \15904 );
buf \U$9920 ( \16075 , \15904 );
buf \U$9921 ( \16076 , \15904 );
buf \U$9922 ( \16077 , \15904 );
buf \U$9923 ( \16078 , \15904 );
buf \U$9924 ( \16079 , \15904 );
buf \U$9925 ( \16080 , \15904 );
buf \U$9926 ( \16081 , \15904 );
buf \U$9927 ( \16082 , \15904 );
buf \U$9928 ( \16083 , \15904 );
buf \U$9929 ( \16084 , \15904 );
buf \U$9930 ( \16085 , \15904 );
buf \U$9931 ( \16086 , \15904 );
buf \U$9932 ( \16087 , \15904 );
buf \U$9933 ( \16088 , \15904 );
buf \U$9934 ( \16089 , \15904 );
buf \U$9935 ( \16090 , \15904 );
buf \U$9936 ( \16091 , \15904 );
buf \U$9937 ( \16092 , \15904 );
buf \U$9938 ( \16093 , \15904 );
buf \U$9939 ( \16094 , \15904 );
buf \U$9940 ( \16095 , \15904 );
nor \U$9941 ( \16096 , \15891 , \15933 , \15893 , \15935 , \15897 , \15901 , \15904 , \16071 , \16072 , \16073 , \16074 , \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 , \16082 , \16083 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 , \16092 , \16093 , \16094 , \16095 );
and \U$9942 ( \16097 , RIe5341b8_6880, \16096 );
buf \U$9943 ( \16098 , \15904 );
buf \U$9944 ( \16099 , \15904 );
buf \U$9945 ( \16100 , \15904 );
buf \U$9946 ( \16101 , \15904 );
buf \U$9947 ( \16102 , \15904 );
buf \U$9948 ( \16103 , \15904 );
buf \U$9949 ( \16104 , \15904 );
buf \U$9950 ( \16105 , \15904 );
buf \U$9951 ( \16106 , \15904 );
buf \U$9952 ( \16107 , \15904 );
buf \U$9953 ( \16108 , \15904 );
buf \U$9954 ( \16109 , \15904 );
buf \U$9955 ( \16110 , \15904 );
buf \U$9956 ( \16111 , \15904 );
buf \U$9957 ( \16112 , \15904 );
buf \U$9958 ( \16113 , \15904 );
buf \U$9959 ( \16114 , \15904 );
buf \U$9960 ( \16115 , \15904 );
buf \U$9961 ( \16116 , \15904 );
buf \U$9962 ( \16117 , \15904 );
buf \U$9963 ( \16118 , \15904 );
buf \U$9964 ( \16119 , \15904 );
buf \U$9965 ( \16120 , \15904 );
buf \U$9966 ( \16121 , \15904 );
buf \U$9967 ( \16122 , \15904 );
nor \U$9968 ( \16123 , \15932 , \15892 , \15893 , \15935 , \15897 , \15901 , \15904 , \16098 , \16099 , \16100 , \16101 , \16102 , \16103 , \16104 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 , \16112 , \16113 , \16114 , \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 , \16122 );
and \U$9969 ( \16124 , RIe5349b0_6879, \16123 );
buf \U$9970 ( \16125 , \15904 );
buf \U$9971 ( \16126 , \15904 );
buf \U$9972 ( \16127 , \15904 );
buf \U$9973 ( \16128 , \15904 );
buf \U$9974 ( \16129 , \15904 );
buf \U$9975 ( \16130 , \15904 );
buf \U$9976 ( \16131 , \15904 );
buf \U$9977 ( \16132 , \15904 );
buf \U$9978 ( \16133 , \15904 );
buf \U$9979 ( \16134 , \15904 );
buf \U$9980 ( \16135 , \15904 );
buf \U$9981 ( \16136 , \15904 );
buf \U$9982 ( \16137 , \15904 );
buf \U$9983 ( \16138 , \15904 );
buf \U$9984 ( \16139 , \15904 );
buf \U$9985 ( \16140 , \15904 );
buf \U$9986 ( \16141 , \15904 );
buf \U$9987 ( \16142 , \15904 );
buf \U$9988 ( \16143 , \15904 );
buf \U$9989 ( \16144 , \15904 );
buf \U$9990 ( \16145 , \15904 );
buf \U$9991 ( \16146 , \15904 );
buf \U$9992 ( \16147 , \15904 );
buf \U$9993 ( \16148 , \15904 );
buf \U$9994 ( \16149 , \15904 );
nor \U$9995 ( \16150 , \15891 , \15892 , \15893 , \15935 , \15897 , \15901 , \15904 , \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 , \16132 , \16133 , \16134 , \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 , \16142 , \16143 , \16144 , \16145 , \16146 , \16147 , \16148 , \16149 );
and \U$9996 ( \16151 , RIea94af8_6890, \16150 );
buf \U$9997 ( \16152 , \15904 );
buf \U$9998 ( \16153 , \15904 );
buf \U$9999 ( \16154 , \15904 );
buf \U$10000 ( \16155 , \15904 );
buf \U$10001 ( \16156 , \15904 );
buf \U$10002 ( \16157 , \15904 );
buf \U$10003 ( \16158 , \15904 );
buf \U$10004 ( \16159 , \15904 );
buf \U$10005 ( \16160 , \15904 );
buf \U$10006 ( \16161 , \15904 );
buf \U$10007 ( \16162 , \15904 );
buf \U$10008 ( \16163 , \15904 );
buf \U$10009 ( \16164 , \15904 );
buf \U$10010 ( \16165 , \15904 );
buf \U$10011 ( \16166 , \15904 );
buf \U$10012 ( \16167 , \15904 );
buf \U$10013 ( \16168 , \15904 );
buf \U$10014 ( \16169 , \15904 );
buf \U$10015 ( \16170 , \15904 );
buf \U$10016 ( \16171 , \15904 );
buf \U$10017 ( \16172 , \15904 );
buf \U$10018 ( \16173 , \15904 );
buf \U$10019 ( \16174 , \15904 );
buf \U$10020 ( \16175 , \15904 );
buf \U$10021 ( \16176 , \15904 );
nor \U$10022 ( \16177 , \15932 , \15933 , \15934 , \15894 , \15897 , \15901 , \15904 , \16152 , \16153 , \16154 , \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 , \16162 , \16163 , \16164 , \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 , \16172 , \16173 , \16174 , \16175 , \16176 );
and \U$10023 ( \16178 , RIe5351a8_6878, \16177 );
buf \U$10024 ( \16179 , \15904 );
buf \U$10025 ( \16180 , \15904 );
buf \U$10026 ( \16181 , \15904 );
buf \U$10027 ( \16182 , \15904 );
buf \U$10028 ( \16183 , \15904 );
buf \U$10029 ( \16184 , \15904 );
buf \U$10030 ( \16185 , \15904 );
buf \U$10031 ( \16186 , \15904 );
buf \U$10032 ( \16187 , \15904 );
buf \U$10033 ( \16188 , \15904 );
buf \U$10034 ( \16189 , \15904 );
buf \U$10035 ( \16190 , \15904 );
buf \U$10036 ( \16191 , \15904 );
buf \U$10037 ( \16192 , \15904 );
buf \U$10038 ( \16193 , \15904 );
buf \U$10039 ( \16194 , \15904 );
buf \U$10040 ( \16195 , \15904 );
buf \U$10041 ( \16196 , \15904 );
buf \U$10042 ( \16197 , \15904 );
buf \U$10043 ( \16198 , \15904 );
buf \U$10044 ( \16199 , \15904 );
buf \U$10045 ( \16200 , \15904 );
buf \U$10046 ( \16201 , \15904 );
buf \U$10047 ( \16202 , \15904 );
buf \U$10048 ( \16203 , \15904 );
nor \U$10049 ( \16204 , \15891 , \15933 , \15934 , \15894 , \15897 , \15901 , \15904 , \16179 , \16180 , \16181 , \16182 , \16183 , \16184 , \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 , \16192 , \16193 , \16194 , \16195 , \16196 , \16197 , \16198 , \16199 , \16200 , \16201 , \16202 , \16203 );
and \U$10050 ( \16205 , RIe5359a0_6877, \16204 );
buf \U$10051 ( \16206 , \15904 );
buf \U$10052 ( \16207 , \15904 );
buf \U$10053 ( \16208 , \15904 );
buf \U$10054 ( \16209 , \15904 );
buf \U$10055 ( \16210 , \15904 );
buf \U$10056 ( \16211 , \15904 );
buf \U$10057 ( \16212 , \15904 );
buf \U$10058 ( \16213 , \15904 );
buf \U$10059 ( \16214 , \15904 );
buf \U$10060 ( \16215 , \15904 );
buf \U$10061 ( \16216 , \15904 );
buf \U$10062 ( \16217 , \15904 );
buf \U$10063 ( \16218 , \15904 );
buf \U$10064 ( \16219 , \15904 );
buf \U$10065 ( \16220 , \15904 );
buf \U$10066 ( \16221 , \15904 );
buf \U$10067 ( \16222 , \15904 );
buf \U$10068 ( \16223 , \15904 );
buf \U$10069 ( \16224 , \15904 );
buf \U$10070 ( \16225 , \15904 );
buf \U$10071 ( \16226 , \15904 );
buf \U$10072 ( \16227 , \15904 );
buf \U$10073 ( \16228 , \15904 );
buf \U$10074 ( \16229 , \15904 );
buf \U$10075 ( \16230 , \15904 );
nor \U$10076 ( \16231 , \15932 , \15892 , \15934 , \15894 , \15897 , \15901 , \15904 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 , \16212 , \16213 , \16214 , \16215 , \16216 , \16217 , \16218 , \16219 , \16220 , \16221 , \16222 , \16223 , \16224 , \16225 , \16226 , \16227 , \16228 , \16229 , \16230 );
and \U$10077 ( \16232 , RIeab78c8_6895, \16231 );
buf \U$10078 ( \16233 , \15904 );
buf \U$10079 ( \16234 , \15904 );
buf \U$10080 ( \16235 , \15904 );
buf \U$10081 ( \16236 , \15904 );
buf \U$10082 ( \16237 , \15904 );
buf \U$10083 ( \16238 , \15904 );
buf \U$10084 ( \16239 , \15904 );
buf \U$10085 ( \16240 , \15904 );
buf \U$10086 ( \16241 , \15904 );
buf \U$10087 ( \16242 , \15904 );
buf \U$10088 ( \16243 , \15904 );
buf \U$10089 ( \16244 , \15904 );
buf \U$10090 ( \16245 , \15904 );
buf \U$10091 ( \16246 , \15904 );
buf \U$10092 ( \16247 , \15904 );
buf \U$10093 ( \16248 , \15904 );
buf \U$10094 ( \16249 , \15904 );
buf \U$10095 ( \16250 , \15904 );
buf \U$10096 ( \16251 , \15904 );
buf \U$10097 ( \16252 , \15904 );
buf \U$10098 ( \16253 , \15904 );
buf \U$10099 ( \16254 , \15904 );
buf \U$10100 ( \16255 , \15904 );
buf \U$10101 ( \16256 , \15904 );
buf \U$10102 ( \16257 , \15904 );
nor \U$10103 ( \16258 , \15891 , \15892 , \15934 , \15894 , \15897 , \15901 , \15904 , \16233 , \16234 , \16235 , \16236 , \16237 , \16238 , \16239 , \16240 , \16241 , \16242 , \16243 , \16244 , \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 , \16252 , \16253 , \16254 , \16255 , \16256 , \16257 );
and \U$10104 ( \16259 , RIeab7d00_6896, \16258 );
buf \U$10105 ( \16260 , \15904 );
buf \U$10106 ( \16261 , \15904 );
buf \U$10107 ( \16262 , \15904 );
buf \U$10108 ( \16263 , \15904 );
buf \U$10109 ( \16264 , \15904 );
buf \U$10110 ( \16265 , \15904 );
buf \U$10111 ( \16266 , \15904 );
buf \U$10112 ( \16267 , \15904 );
buf \U$10113 ( \16268 , \15904 );
buf \U$10114 ( \16269 , \15904 );
buf \U$10115 ( \16270 , \15904 );
buf \U$10116 ( \16271 , \15904 );
buf \U$10117 ( \16272 , \15904 );
buf \U$10118 ( \16273 , \15904 );
buf \U$10119 ( \16274 , \15904 );
buf \U$10120 ( \16275 , \15904 );
buf \U$10121 ( \16276 , \15904 );
buf \U$10122 ( \16277 , \15904 );
buf \U$10123 ( \16278 , \15904 );
buf \U$10124 ( \16279 , \15904 );
buf \U$10125 ( \16280 , \15904 );
buf \U$10126 ( \16281 , \15904 );
buf \U$10127 ( \16282 , \15904 );
buf \U$10128 ( \16283 , \15904 );
buf \U$10129 ( \16284 , \15904 );
nor \U$10130 ( \16285 , \15932 , \15933 , \15893 , \15894 , \15897 , \15901 , \15904 , \16260 , \16261 , \16262 , \16263 , \16264 , \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 , \16272 , \16273 , \16274 , \16275 , \16276 , \16277 , \16278 , \16279 , \16280 , \16281 , \16282 , \16283 , \16284 );
and \U$10131 ( \16286 , RIeacfa18_6902, \16285 );
buf \U$10132 ( \16287 , \15904 );
buf \U$10133 ( \16288 , \15904 );
buf \U$10134 ( \16289 , \15904 );
buf \U$10135 ( \16290 , \15904 );
buf \U$10136 ( \16291 , \15904 );
buf \U$10137 ( \16292 , \15904 );
buf \U$10138 ( \16293 , \15904 );
buf \U$10139 ( \16294 , \15904 );
buf \U$10140 ( \16295 , \15904 );
buf \U$10141 ( \16296 , \15904 );
buf \U$10142 ( \16297 , \15904 );
buf \U$10143 ( \16298 , \15904 );
buf \U$10144 ( \16299 , \15904 );
buf \U$10145 ( \16300 , \15904 );
buf \U$10146 ( \16301 , \15904 );
buf \U$10147 ( \16302 , \15904 );
buf \U$10148 ( \16303 , \15904 );
buf \U$10149 ( \16304 , \15904 );
buf \U$10150 ( \16305 , \15904 );
buf \U$10151 ( \16306 , \15904 );
buf \U$10152 ( \16307 , \15904 );
buf \U$10153 ( \16308 , \15904 );
buf \U$10154 ( \16309 , \15904 );
buf \U$10155 ( \16310 , \15904 );
buf \U$10156 ( \16311 , \15904 );
nor \U$10157 ( \16312 , \15891 , \15933 , \15893 , \15894 , \15897 , \15901 , \15904 , \16287 , \16288 , \16289 , \16290 , \16291 , \16292 , \16293 , \16294 , \16295 , \16296 , \16297 , \16298 , \16299 , \16300 , \16301 , \16302 , \16303 , \16304 , \16305 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 );
and \U$10158 ( \16313 , RIeab6518_6891, \16312 );
buf \U$10159 ( \16314 , \15904 );
buf \U$10160 ( \16315 , \15904 );
buf \U$10161 ( \16316 , \15904 );
buf \U$10162 ( \16317 , \15904 );
buf \U$10163 ( \16318 , \15904 );
buf \U$10164 ( \16319 , \15904 );
buf \U$10165 ( \16320 , \15904 );
buf \U$10166 ( \16321 , \15904 );
buf \U$10167 ( \16322 , \15904 );
buf \U$10168 ( \16323 , \15904 );
buf \U$10169 ( \16324 , \15904 );
buf \U$10170 ( \16325 , \15904 );
buf \U$10171 ( \16326 , \15904 );
buf \U$10172 ( \16327 , \15904 );
buf \U$10173 ( \16328 , \15904 );
buf \U$10174 ( \16329 , \15904 );
buf \U$10175 ( \16330 , \15904 );
buf \U$10176 ( \16331 , \15904 );
buf \U$10177 ( \16332 , \15904 );
buf \U$10178 ( \16333 , \15904 );
buf \U$10179 ( \16334 , \15904 );
buf \U$10180 ( \16335 , \15904 );
buf \U$10181 ( \16336 , \15904 );
buf \U$10182 ( \16337 , \15904 );
buf \U$10183 ( \16338 , \15904 );
nor \U$10184 ( \16339 , \15932 , \15892 , \15893 , \15894 , \15897 , \15901 , \15904 , \16314 , \16315 , \16316 , \16317 , \16318 , \16319 , \16320 , \16321 , \16322 , \16323 , \16324 , \16325 , \16326 , \16327 , \16328 , \16329 , \16330 , \16331 , \16332 , \16333 , \16334 , \16335 , \16336 , \16337 , \16338 );
and \U$10185 ( \16340 , RIeb352c8_6904, \16339 );
or \U$10186 ( \16341 , \15931 , \15962 , \15989 , \16016 , \16043 , \16070 , \16097 , \16124 , \16151 , \16178 , \16205 , \16232 , \16259 , \16286 , \16313 , \16340 );
buf \U$10187 ( \16342 , \15904 );
not \U$10188 ( \16343 , \16342 );
buf \U$10189 ( \16344 , \15892 );
buf \U$10190 ( \16345 , \15893 );
buf \U$10191 ( \16346 , \15894 );
buf \U$10192 ( \16347 , \15897 );
buf \U$10193 ( \16348 , \15901 );
buf \U$10194 ( \16349 , \15904 );
buf \U$10195 ( \16350 , \15904 );
buf \U$10196 ( \16351 , \15904 );
buf \U$10197 ( \16352 , \15904 );
buf \U$10198 ( \16353 , \15904 );
buf \U$10199 ( \16354 , \15904 );
buf \U$10200 ( \16355 , \15904 );
buf \U$10201 ( \16356 , \15904 );
buf \U$10202 ( \16357 , \15904 );
buf \U$10203 ( \16358 , \15904 );
buf \U$10204 ( \16359 , \15904 );
buf \U$10205 ( \16360 , \15904 );
buf \U$10206 ( \16361 , \15904 );
buf \U$10207 ( \16362 , \15904 );
buf \U$10208 ( \16363 , \15904 );
buf \U$10209 ( \16364 , \15904 );
buf \U$10210 ( \16365 , \15904 );
buf \U$10211 ( \16366 , \15904 );
buf \U$10212 ( \16367 , \15904 );
buf \U$10213 ( \16368 , \15904 );
buf \U$10214 ( \16369 , \15904 );
buf \U$10215 ( \16370 , \15904 );
buf \U$10216 ( \16371 , \15904 );
buf \U$10217 ( \16372 , \15904 );
buf \U$10218 ( \16373 , \15904 );
buf \U$10219 ( \16374 , \15891 );
or \U$10220 ( \16375 , \16344 , \16345 , \16346 , \16347 , \16348 , \16349 , \16350 , \16351 , \16352 , \16353 , \16354 , \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 , \16362 , \16363 , \16364 , \16365 , \16366 , \16367 , \16368 , \16369 , \16370 , \16371 , \16372 , \16373 , \16374 );
nand \U$10221 ( \16376 , \16343 , \16375 );
buf \U$10222 ( \16377 , \16376 );
buf \U$10223 ( \16378 , \15904 );
not \U$10224 ( \16379 , \16378 );
buf \U$10225 ( \16380 , \15901 );
buf \U$10226 ( \16381 , \15904 );
buf \U$10227 ( \16382 , \15904 );
buf \U$10228 ( \16383 , \15904 );
buf \U$10229 ( \16384 , \15904 );
buf \U$10230 ( \16385 , \15904 );
buf \U$10231 ( \16386 , \15904 );
buf \U$10232 ( \16387 , \15904 );
buf \U$10233 ( \16388 , \15904 );
buf \U$10234 ( \16389 , \15904 );
buf \U$10235 ( \16390 , \15904 );
buf \U$10236 ( \16391 , \15904 );
buf \U$10237 ( \16392 , \15904 );
buf \U$10238 ( \16393 , \15904 );
buf \U$10239 ( \16394 , \15904 );
buf \U$10240 ( \16395 , \15904 );
buf \U$10241 ( \16396 , \15904 );
buf \U$10242 ( \16397 , \15904 );
buf \U$10243 ( \16398 , \15904 );
buf \U$10244 ( \16399 , \15904 );
buf \U$10245 ( \16400 , \15904 );
buf \U$10246 ( \16401 , \15904 );
buf \U$10247 ( \16402 , \15904 );
buf \U$10248 ( \16403 , \15904 );
buf \U$10249 ( \16404 , \15904 );
buf \U$10250 ( \16405 , \15904 );
buf \U$10251 ( \16406 , \15897 );
buf \U$10252 ( \16407 , \15891 );
buf \U$10253 ( \16408 , \15892 );
buf \U$10254 ( \16409 , \15893 );
buf \U$10255 ( \16410 , \15894 );
or \U$10256 ( \16411 , \16407 , \16408 , \16409 , \16410 );
and \U$10257 ( \16412 , \16406 , \16411 );
or \U$10258 ( \16413 , \16380 , \16381 , \16382 , \16383 , \16384 , \16385 , \16386 , \16387 , \16388 , \16389 , \16390 , \16391 , \16392 , \16393 , \16394 , \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 , \16402 , \16403 , \16404 , \16405 , \16412 );
and \U$10259 ( \16414 , \16379 , \16413 );
buf \U$10260 ( \16415 , \16414 );
or \U$10261 ( \16416 , \16377 , \16415 );
_DC g56f5 ( \16417_nG56f5 , \16341 , \16416 );
not \U$10262 ( \16418 , \16417_nG56f5 );
buf \U$10263 ( \16419 , RIb7b9608_246);
buf \U$10264 ( \16420 , \15904 );
buf \U$10265 ( \16421 , \15904 );
buf \U$10266 ( \16422 , \15904 );
buf \U$10267 ( \16423 , \15904 );
buf \U$10268 ( \16424 , \15904 );
buf \U$10269 ( \16425 , \15904 );
buf \U$10270 ( \16426 , \15904 );
buf \U$10271 ( \16427 , \15904 );
buf \U$10272 ( \16428 , \15904 );
buf \U$10273 ( \16429 , \15904 );
buf \U$10274 ( \16430 , \15904 );
buf \U$10275 ( \16431 , \15904 );
buf \U$10276 ( \16432 , \15904 );
buf \U$10277 ( \16433 , \15904 );
buf \U$10278 ( \16434 , \15904 );
buf \U$10279 ( \16435 , \15904 );
buf \U$10280 ( \16436 , \15904 );
buf \U$10281 ( \16437 , \15904 );
buf \U$10282 ( \16438 , \15904 );
buf \U$10283 ( \16439 , \15904 );
buf \U$10284 ( \16440 , \15904 );
buf \U$10285 ( \16441 , \15904 );
buf \U$10286 ( \16442 , \15904 );
buf \U$10287 ( \16443 , \15904 );
buf \U$10288 ( \16444 , \15904 );
nor \U$10289 ( \16445 , \15891 , \15892 , \15893 , \15894 , \15898 , \15901 , \15904 , \16420 , \16421 , \16422 , \16423 , \16424 , \16425 , \16426 , \16427 , \16428 , \16429 , \16430 , \16431 , \16432 , \16433 , \16434 , \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 , \16442 , \16443 , \16444 );
and \U$10290 ( \16446 , \7117 , \16445 );
buf \U$10291 ( \16447 , \15904 );
buf \U$10292 ( \16448 , \15904 );
buf \U$10293 ( \16449 , \15904 );
buf \U$10294 ( \16450 , \15904 );
buf \U$10295 ( \16451 , \15904 );
buf \U$10296 ( \16452 , \15904 );
buf \U$10297 ( \16453 , \15904 );
buf \U$10298 ( \16454 , \15904 );
buf \U$10299 ( \16455 , \15904 );
buf \U$10300 ( \16456 , \15904 );
buf \U$10301 ( \16457 , \15904 );
buf \U$10302 ( \16458 , \15904 );
buf \U$10303 ( \16459 , \15904 );
buf \U$10304 ( \16460 , \15904 );
buf \U$10305 ( \16461 , \15904 );
buf \U$10306 ( \16462 , \15904 );
buf \U$10307 ( \16463 , \15904 );
buf \U$10308 ( \16464 , \15904 );
buf \U$10309 ( \16465 , \15904 );
buf \U$10310 ( \16466 , \15904 );
buf \U$10311 ( \16467 , \15904 );
buf \U$10312 ( \16468 , \15904 );
buf \U$10313 ( \16469 , \15904 );
buf \U$10314 ( \16470 , \15904 );
buf \U$10315 ( \16471 , \15904 );
nor \U$10316 ( \16472 , \15932 , \15933 , \15934 , \15935 , \15897 , \15901 , \15904 , \16447 , \16448 , \16449 , \16450 , \16451 , \16452 , \16453 , \16454 , \16455 , \16456 , \16457 , \16458 , \16459 , \16460 , \16461 , \16462 , \16463 , \16464 , \16465 , \16466 , \16467 , \16468 , \16469 , \16470 , \16471 );
and \U$10317 ( \16473 , \7119 , \16472 );
buf \U$10318 ( \16474 , \15904 );
buf \U$10319 ( \16475 , \15904 );
buf \U$10320 ( \16476 , \15904 );
buf \U$10321 ( \16477 , \15904 );
buf \U$10322 ( \16478 , \15904 );
buf \U$10323 ( \16479 , \15904 );
buf \U$10324 ( \16480 , \15904 );
buf \U$10325 ( \16481 , \15904 );
buf \U$10326 ( \16482 , \15904 );
buf \U$10327 ( \16483 , \15904 );
buf \U$10328 ( \16484 , \15904 );
buf \U$10329 ( \16485 , \15904 );
buf \U$10330 ( \16486 , \15904 );
buf \U$10331 ( \16487 , \15904 );
buf \U$10332 ( \16488 , \15904 );
buf \U$10333 ( \16489 , \15904 );
buf \U$10334 ( \16490 , \15904 );
buf \U$10335 ( \16491 , \15904 );
buf \U$10336 ( \16492 , \15904 );
buf \U$10337 ( \16493 , \15904 );
buf \U$10338 ( \16494 , \15904 );
buf \U$10339 ( \16495 , \15904 );
buf \U$10340 ( \16496 , \15904 );
buf \U$10341 ( \16497 , \15904 );
buf \U$10342 ( \16498 , \15904 );
nor \U$10343 ( \16499 , \15891 , \15933 , \15934 , \15935 , \15897 , \15901 , \15904 , \16474 , \16475 , \16476 , \16477 , \16478 , \16479 , \16480 , \16481 , \16482 , \16483 , \16484 , \16485 , \16486 , \16487 , \16488 , \16489 , \16490 , \16491 , \16492 , \16493 , \16494 , \16495 , \16496 , \16497 , \16498 );
and \U$10344 ( \16500 , \7864 , \16499 );
buf \U$10345 ( \16501 , \15904 );
buf \U$10346 ( \16502 , \15904 );
buf \U$10347 ( \16503 , \15904 );
buf \U$10348 ( \16504 , \15904 );
buf \U$10349 ( \16505 , \15904 );
buf \U$10350 ( \16506 , \15904 );
buf \U$10351 ( \16507 , \15904 );
buf \U$10352 ( \16508 , \15904 );
buf \U$10353 ( \16509 , \15904 );
buf \U$10354 ( \16510 , \15904 );
buf \U$10355 ( \16511 , \15904 );
buf \U$10356 ( \16512 , \15904 );
buf \U$10357 ( \16513 , \15904 );
buf \U$10358 ( \16514 , \15904 );
buf \U$10359 ( \16515 , \15904 );
buf \U$10360 ( \16516 , \15904 );
buf \U$10361 ( \16517 , \15904 );
buf \U$10362 ( \16518 , \15904 );
buf \U$10363 ( \16519 , \15904 );
buf \U$10364 ( \16520 , \15904 );
buf \U$10365 ( \16521 , \15904 );
buf \U$10366 ( \16522 , \15904 );
buf \U$10367 ( \16523 , \15904 );
buf \U$10368 ( \16524 , \15904 );
buf \U$10369 ( \16525 , \15904 );
nor \U$10370 ( \16526 , \15932 , \15892 , \15934 , \15935 , \15897 , \15901 , \15904 , \16501 , \16502 , \16503 , \16504 , \16505 , \16506 , \16507 , \16508 , \16509 , \16510 , \16511 , \16512 , \16513 , \16514 , \16515 , \16516 , \16517 , \16518 , \16519 , \16520 , \16521 , \16522 , \16523 , \16524 , \16525 );
and \U$10371 ( \16527 , \7892 , \16526 );
buf \U$10372 ( \16528 , \15904 );
buf \U$10373 ( \16529 , \15904 );
buf \U$10374 ( \16530 , \15904 );
buf \U$10375 ( \16531 , \15904 );
buf \U$10376 ( \16532 , \15904 );
buf \U$10377 ( \16533 , \15904 );
buf \U$10378 ( \16534 , \15904 );
buf \U$10379 ( \16535 , \15904 );
buf \U$10380 ( \16536 , \15904 );
buf \U$10381 ( \16537 , \15904 );
buf \U$10382 ( \16538 , \15904 );
buf \U$10383 ( \16539 , \15904 );
buf \U$10384 ( \16540 , \15904 );
buf \U$10385 ( \16541 , \15904 );
buf \U$10386 ( \16542 , \15904 );
buf \U$10387 ( \16543 , \15904 );
buf \U$10388 ( \16544 , \15904 );
buf \U$10389 ( \16545 , \15904 );
buf \U$10390 ( \16546 , \15904 );
buf \U$10391 ( \16547 , \15904 );
buf \U$10392 ( \16548 , \15904 );
buf \U$10393 ( \16549 , \15904 );
buf \U$10394 ( \16550 , \15904 );
buf \U$10395 ( \16551 , \15904 );
buf \U$10396 ( \16552 , \15904 );
nor \U$10397 ( \16553 , \15891 , \15892 , \15934 , \15935 , \15897 , \15901 , \15904 , \16528 , \16529 , \16530 , \16531 , \16532 , \16533 , \16534 , \16535 , \16536 , \16537 , \16538 , \16539 , \16540 , \16541 , \16542 , \16543 , \16544 , \16545 , \16546 , \16547 , \16548 , \16549 , \16550 , \16551 , \16552 );
and \U$10398 ( \16554 , \7920 , \16553 );
buf \U$10399 ( \16555 , \15904 );
buf \U$10400 ( \16556 , \15904 );
buf \U$10401 ( \16557 , \15904 );
buf \U$10402 ( \16558 , \15904 );
buf \U$10403 ( \16559 , \15904 );
buf \U$10404 ( \16560 , \15904 );
buf \U$10405 ( \16561 , \15904 );
buf \U$10406 ( \16562 , \15904 );
buf \U$10407 ( \16563 , \15904 );
buf \U$10408 ( \16564 , \15904 );
buf \U$10409 ( \16565 , \15904 );
buf \U$10410 ( \16566 , \15904 );
buf \U$10411 ( \16567 , \15904 );
buf \U$10412 ( \16568 , \15904 );
buf \U$10413 ( \16569 , \15904 );
buf \U$10414 ( \16570 , \15904 );
buf \U$10415 ( \16571 , \15904 );
buf \U$10416 ( \16572 , \15904 );
buf \U$10417 ( \16573 , \15904 );
buf \U$10418 ( \16574 , \15904 );
buf \U$10419 ( \16575 , \15904 );
buf \U$10420 ( \16576 , \15904 );
buf \U$10421 ( \16577 , \15904 );
buf \U$10422 ( \16578 , \15904 );
buf \U$10423 ( \16579 , \15904 );
nor \U$10424 ( \16580 , \15932 , \15933 , \15893 , \15935 , \15897 , \15901 , \15904 , \16555 , \16556 , \16557 , \16558 , \16559 , \16560 , \16561 , \16562 , \16563 , \16564 , \16565 , \16566 , \16567 , \16568 , \16569 , \16570 , \16571 , \16572 , \16573 , \16574 , \16575 , \16576 , \16577 , \16578 , \16579 );
and \U$10425 ( \16581 , \7948 , \16580 );
buf \U$10426 ( \16582 , \15904 );
buf \U$10427 ( \16583 , \15904 );
buf \U$10428 ( \16584 , \15904 );
buf \U$10429 ( \16585 , \15904 );
buf \U$10430 ( \16586 , \15904 );
buf \U$10431 ( \16587 , \15904 );
buf \U$10432 ( \16588 , \15904 );
buf \U$10433 ( \16589 , \15904 );
buf \U$10434 ( \16590 , \15904 );
buf \U$10435 ( \16591 , \15904 );
buf \U$10436 ( \16592 , \15904 );
buf \U$10437 ( \16593 , \15904 );
buf \U$10438 ( \16594 , \15904 );
buf \U$10439 ( \16595 , \15904 );
buf \U$10440 ( \16596 , \15904 );
buf \U$10441 ( \16597 , \15904 );
buf \U$10442 ( \16598 , \15904 );
buf \U$10443 ( \16599 , \15904 );
buf \U$10444 ( \16600 , \15904 );
buf \U$10445 ( \16601 , \15904 );
buf \U$10446 ( \16602 , \15904 );
buf \U$10447 ( \16603 , \15904 );
buf \U$10448 ( \16604 , \15904 );
buf \U$10449 ( \16605 , \15904 );
buf \U$10450 ( \16606 , \15904 );
nor \U$10451 ( \16607 , \15891 , \15933 , \15893 , \15935 , \15897 , \15901 , \15904 , \16582 , \16583 , \16584 , \16585 , \16586 , \16587 , \16588 , \16589 , \16590 , \16591 , \16592 , \16593 , \16594 , \16595 , \16596 , \16597 , \16598 , \16599 , \16600 , \16601 , \16602 , \16603 , \16604 , \16605 , \16606 );
and \U$10452 ( \16608 , \7976 , \16607 );
buf \U$10453 ( \16609 , \15904 );
buf \U$10454 ( \16610 , \15904 );
buf \U$10455 ( \16611 , \15904 );
buf \U$10456 ( \16612 , \15904 );
buf \U$10457 ( \16613 , \15904 );
buf \U$10458 ( \16614 , \15904 );
buf \U$10459 ( \16615 , \15904 );
buf \U$10460 ( \16616 , \15904 );
buf \U$10461 ( \16617 , \15904 );
buf \U$10462 ( \16618 , \15904 );
buf \U$10463 ( \16619 , \15904 );
buf \U$10464 ( \16620 , \15904 );
buf \U$10465 ( \16621 , \15904 );
buf \U$10466 ( \16622 , \15904 );
buf \U$10467 ( \16623 , \15904 );
buf \U$10468 ( \16624 , \15904 );
buf \U$10469 ( \16625 , \15904 );
buf \U$10470 ( \16626 , \15904 );
buf \U$10471 ( \16627 , \15904 );
buf \U$10472 ( \16628 , \15904 );
buf \U$10473 ( \16629 , \15904 );
buf \U$10474 ( \16630 , \15904 );
buf \U$10475 ( \16631 , \15904 );
buf \U$10476 ( \16632 , \15904 );
buf \U$10477 ( \16633 , \15904 );
nor \U$10478 ( \16634 , \15932 , \15892 , \15893 , \15935 , \15897 , \15901 , \15904 , \16609 , \16610 , \16611 , \16612 , \16613 , \16614 , \16615 , \16616 , \16617 , \16618 , \16619 , \16620 , \16621 , \16622 , \16623 , \16624 , \16625 , \16626 , \16627 , \16628 , \16629 , \16630 , \16631 , \16632 , \16633 );
and \U$10479 ( \16635 , \8004 , \16634 );
buf \U$10480 ( \16636 , \15904 );
buf \U$10481 ( \16637 , \15904 );
buf \U$10482 ( \16638 , \15904 );
buf \U$10483 ( \16639 , \15904 );
buf \U$10484 ( \16640 , \15904 );
buf \U$10485 ( \16641 , \15904 );
buf \U$10486 ( \16642 , \15904 );
buf \U$10487 ( \16643 , \15904 );
buf \U$10488 ( \16644 , \15904 );
buf \U$10489 ( \16645 , \15904 );
buf \U$10490 ( \16646 , \15904 );
buf \U$10491 ( \16647 , \15904 );
buf \U$10492 ( \16648 , \15904 );
buf \U$10493 ( \16649 , \15904 );
buf \U$10494 ( \16650 , \15904 );
buf \U$10495 ( \16651 , \15904 );
buf \U$10496 ( \16652 , \15904 );
buf \U$10497 ( \16653 , \15904 );
buf \U$10498 ( \16654 , \15904 );
buf \U$10499 ( \16655 , \15904 );
buf \U$10500 ( \16656 , \15904 );
buf \U$10501 ( \16657 , \15904 );
buf \U$10502 ( \16658 , \15904 );
buf \U$10503 ( \16659 , \15904 );
buf \U$10504 ( \16660 , \15904 );
nor \U$10505 ( \16661 , \15891 , \15892 , \15893 , \15935 , \15897 , \15901 , \15904 , \16636 , \16637 , \16638 , \16639 , \16640 , \16641 , \16642 , \16643 , \16644 , \16645 , \16646 , \16647 , \16648 , \16649 , \16650 , \16651 , \16652 , \16653 , \16654 , \16655 , \16656 , \16657 , \16658 , \16659 , \16660 );
and \U$10506 ( \16662 , \8032 , \16661 );
buf \U$10507 ( \16663 , \15904 );
buf \U$10508 ( \16664 , \15904 );
buf \U$10509 ( \16665 , \15904 );
buf \U$10510 ( \16666 , \15904 );
buf \U$10511 ( \16667 , \15904 );
buf \U$10512 ( \16668 , \15904 );
buf \U$10513 ( \16669 , \15904 );
buf \U$10514 ( \16670 , \15904 );
buf \U$10515 ( \16671 , \15904 );
buf \U$10516 ( \16672 , \15904 );
buf \U$10517 ( \16673 , \15904 );
buf \U$10518 ( \16674 , \15904 );
buf \U$10519 ( \16675 , \15904 );
buf \U$10520 ( \16676 , \15904 );
buf \U$10521 ( \16677 , \15904 );
buf \U$10522 ( \16678 , \15904 );
buf \U$10523 ( \16679 , \15904 );
buf \U$10524 ( \16680 , \15904 );
buf \U$10525 ( \16681 , \15904 );
buf \U$10526 ( \16682 , \15904 );
buf \U$10527 ( \16683 , \15904 );
buf \U$10528 ( \16684 , \15904 );
buf \U$10529 ( \16685 , \15904 );
buf \U$10530 ( \16686 , \15904 );
buf \U$10531 ( \16687 , \15904 );
nor \U$10532 ( \16688 , \15932 , \15933 , \15934 , \15894 , \15897 , \15901 , \15904 , \16663 , \16664 , \16665 , \16666 , \16667 , \16668 , \16669 , \16670 , \16671 , \16672 , \16673 , \16674 , \16675 , \16676 , \16677 , \16678 , \16679 , \16680 , \16681 , \16682 , \16683 , \16684 , \16685 , \16686 , \16687 );
and \U$10533 ( \16689 , \8060 , \16688 );
buf \U$10534 ( \16690 , \15904 );
buf \U$10535 ( \16691 , \15904 );
buf \U$10536 ( \16692 , \15904 );
buf \U$10537 ( \16693 , \15904 );
buf \U$10538 ( \16694 , \15904 );
buf \U$10539 ( \16695 , \15904 );
buf \U$10540 ( \16696 , \15904 );
buf \U$10541 ( \16697 , \15904 );
buf \U$10542 ( \16698 , \15904 );
buf \U$10543 ( \16699 , \15904 );
buf \U$10544 ( \16700 , \15904 );
buf \U$10545 ( \16701 , \15904 );
buf \U$10546 ( \16702 , \15904 );
buf \U$10547 ( \16703 , \15904 );
buf \U$10548 ( \16704 , \15904 );
buf \U$10549 ( \16705 , \15904 );
buf \U$10550 ( \16706 , \15904 );
buf \U$10551 ( \16707 , \15904 );
buf \U$10552 ( \16708 , \15904 );
buf \U$10553 ( \16709 , \15904 );
buf \U$10554 ( \16710 , \15904 );
buf \U$10555 ( \16711 , \15904 );
buf \U$10556 ( \16712 , \15904 );
buf \U$10557 ( \16713 , \15904 );
buf \U$10558 ( \16714 , \15904 );
nor \U$10559 ( \16715 , \15891 , \15933 , \15934 , \15894 , \15897 , \15901 , \15904 , \16690 , \16691 , \16692 , \16693 , \16694 , \16695 , \16696 , \16697 , \16698 , \16699 , \16700 , \16701 , \16702 , \16703 , \16704 , \16705 , \16706 , \16707 , \16708 , \16709 , \16710 , \16711 , \16712 , \16713 , \16714 );
and \U$10560 ( \16716 , \8088 , \16715 );
buf \U$10561 ( \16717 , \15904 );
buf \U$10562 ( \16718 , \15904 );
buf \U$10563 ( \16719 , \15904 );
buf \U$10564 ( \16720 , \15904 );
buf \U$10565 ( \16721 , \15904 );
buf \U$10566 ( \16722 , \15904 );
buf \U$10567 ( \16723 , \15904 );
buf \U$10568 ( \16724 , \15904 );
buf \U$10569 ( \16725 , \15904 );
buf \U$10570 ( \16726 , \15904 );
buf \U$10571 ( \16727 , \15904 );
buf \U$10572 ( \16728 , \15904 );
buf \U$10573 ( \16729 , \15904 );
buf \U$10574 ( \16730 , \15904 );
buf \U$10575 ( \16731 , \15904 );
buf \U$10576 ( \16732 , \15904 );
buf \U$10577 ( \16733 , \15904 );
buf \U$10578 ( \16734 , \15904 );
buf \U$10579 ( \16735 , \15904 );
buf \U$10580 ( \16736 , \15904 );
buf \U$10581 ( \16737 , \15904 );
buf \U$10582 ( \16738 , \15904 );
buf \U$10583 ( \16739 , \15904 );
buf \U$10584 ( \16740 , \15904 );
buf \U$10585 ( \16741 , \15904 );
nor \U$10586 ( \16742 , \15932 , \15892 , \15934 , \15894 , \15897 , \15901 , \15904 , \16717 , \16718 , \16719 , \16720 , \16721 , \16722 , \16723 , \16724 , \16725 , \16726 , \16727 , \16728 , \16729 , \16730 , \16731 , \16732 , \16733 , \16734 , \16735 , \16736 , \16737 , \16738 , \16739 , \16740 , \16741 );
and \U$10587 ( \16743 , \8116 , \16742 );
buf \U$10588 ( \16744 , \15904 );
buf \U$10589 ( \16745 , \15904 );
buf \U$10590 ( \16746 , \15904 );
buf \U$10591 ( \16747 , \15904 );
buf \U$10592 ( \16748 , \15904 );
buf \U$10593 ( \16749 , \15904 );
buf \U$10594 ( \16750 , \15904 );
buf \U$10595 ( \16751 , \15904 );
buf \U$10596 ( \16752 , \15904 );
buf \U$10597 ( \16753 , \15904 );
buf \U$10598 ( \16754 , \15904 );
buf \U$10599 ( \16755 , \15904 );
buf \U$10600 ( \16756 , \15904 );
buf \U$10601 ( \16757 , \15904 );
buf \U$10602 ( \16758 , \15904 );
buf \U$10603 ( \16759 , \15904 );
buf \U$10604 ( \16760 , \15904 );
buf \U$10605 ( \16761 , \15904 );
buf \U$10606 ( \16762 , \15904 );
buf \U$10607 ( \16763 , \15904 );
buf \U$10608 ( \16764 , \15904 );
buf \U$10609 ( \16765 , \15904 );
buf \U$10610 ( \16766 , \15904 );
buf \U$10611 ( \16767 , \15904 );
buf \U$10612 ( \16768 , \15904 );
nor \U$10613 ( \16769 , \15891 , \15892 , \15934 , \15894 , \15897 , \15901 , \15904 , \16744 , \16745 , \16746 , \16747 , \16748 , \16749 , \16750 , \16751 , \16752 , \16753 , \16754 , \16755 , \16756 , \16757 , \16758 , \16759 , \16760 , \16761 , \16762 , \16763 , \16764 , \16765 , \16766 , \16767 , \16768 );
and \U$10614 ( \16770 , \8144 , \16769 );
buf \U$10615 ( \16771 , \15904 );
buf \U$10616 ( \16772 , \15904 );
buf \U$10617 ( \16773 , \15904 );
buf \U$10618 ( \16774 , \15904 );
buf \U$10619 ( \16775 , \15904 );
buf \U$10620 ( \16776 , \15904 );
buf \U$10621 ( \16777 , \15904 );
buf \U$10622 ( \16778 , \15904 );
buf \U$10623 ( \16779 , \15904 );
buf \U$10624 ( \16780 , \15904 );
buf \U$10625 ( \16781 , \15904 );
buf \U$10626 ( \16782 , \15904 );
buf \U$10627 ( \16783 , \15904 );
buf \U$10628 ( \16784 , \15904 );
buf \U$10629 ( \16785 , \15904 );
buf \U$10630 ( \16786 , \15904 );
buf \U$10631 ( \16787 , \15904 );
buf \U$10632 ( \16788 , \15904 );
buf \U$10633 ( \16789 , \15904 );
buf \U$10634 ( \16790 , \15904 );
buf \U$10635 ( \16791 , \15904 );
buf \U$10636 ( \16792 , \15904 );
buf \U$10637 ( \16793 , \15904 );
buf \U$10638 ( \16794 , \15904 );
buf \U$10639 ( \16795 , \15904 );
nor \U$10640 ( \16796 , \15932 , \15933 , \15893 , \15894 , \15897 , \15901 , \15904 , \16771 , \16772 , \16773 , \16774 , \16775 , \16776 , \16777 , \16778 , \16779 , \16780 , \16781 , \16782 , \16783 , \16784 , \16785 , \16786 , \16787 , \16788 , \16789 , \16790 , \16791 , \16792 , \16793 , \16794 , \16795 );
and \U$10641 ( \16797 , \8172 , \16796 );
buf \U$10642 ( \16798 , \15904 );
buf \U$10643 ( \16799 , \15904 );
buf \U$10644 ( \16800 , \15904 );
buf \U$10645 ( \16801 , \15904 );
buf \U$10646 ( \16802 , \15904 );
buf \U$10647 ( \16803 , \15904 );
buf \U$10648 ( \16804 , \15904 );
buf \U$10649 ( \16805 , \15904 );
buf \U$10650 ( \16806 , \15904 );
buf \U$10651 ( \16807 , \15904 );
buf \U$10652 ( \16808 , \15904 );
buf \U$10653 ( \16809 , \15904 );
buf \U$10654 ( \16810 , \15904 );
buf \U$10655 ( \16811 , \15904 );
buf \U$10656 ( \16812 , \15904 );
buf \U$10657 ( \16813 , \15904 );
buf \U$10658 ( \16814 , \15904 );
buf \U$10659 ( \16815 , \15904 );
buf \U$10660 ( \16816 , \15904 );
buf \U$10661 ( \16817 , \15904 );
buf \U$10662 ( \16818 , \15904 );
buf \U$10663 ( \16819 , \15904 );
buf \U$10664 ( \16820 , \15904 );
buf \U$10665 ( \16821 , \15904 );
buf \U$10666 ( \16822 , \15904 );
nor \U$10667 ( \16823 , \15891 , \15933 , \15893 , \15894 , \15897 , \15901 , \15904 , \16798 , \16799 , \16800 , \16801 , \16802 , \16803 , \16804 , \16805 , \16806 , \16807 , \16808 , \16809 , \16810 , \16811 , \16812 , \16813 , \16814 , \16815 , \16816 , \16817 , \16818 , \16819 , \16820 , \16821 , \16822 );
and \U$10668 ( \16824 , \8200 , \16823 );
buf \U$10669 ( \16825 , \15904 );
buf \U$10670 ( \16826 , \15904 );
buf \U$10671 ( \16827 , \15904 );
buf \U$10672 ( \16828 , \15904 );
buf \U$10673 ( \16829 , \15904 );
buf \U$10674 ( \16830 , \15904 );
buf \U$10675 ( \16831 , \15904 );
buf \U$10676 ( \16832 , \15904 );
buf \U$10677 ( \16833 , \15904 );
buf \U$10678 ( \16834 , \15904 );
buf \U$10679 ( \16835 , \15904 );
buf \U$10680 ( \16836 , \15904 );
buf \U$10681 ( \16837 , \15904 );
buf \U$10682 ( \16838 , \15904 );
buf \U$10683 ( \16839 , \15904 );
buf \U$10684 ( \16840 , \15904 );
buf \U$10685 ( \16841 , \15904 );
buf \U$10686 ( \16842 , \15904 );
buf \U$10687 ( \16843 , \15904 );
buf \U$10688 ( \16844 , \15904 );
buf \U$10689 ( \16845 , \15904 );
buf \U$10690 ( \16846 , \15904 );
buf \U$10691 ( \16847 , \15904 );
buf \U$10692 ( \16848 , \15904 );
buf \U$10693 ( \16849 , \15904 );
nor \U$10694 ( \16850 , \15932 , \15892 , \15893 , \15894 , \15897 , \15901 , \15904 , \16825 , \16826 , \16827 , \16828 , \16829 , \16830 , \16831 , \16832 , \16833 , \16834 , \16835 , \16836 , \16837 , \16838 , \16839 , \16840 , \16841 , \16842 , \16843 , \16844 , \16845 , \16846 , \16847 , \16848 , \16849 );
and \U$10695 ( \16851 , \8228 , \16850 );
or \U$10696 ( \16852 , \16446 , \16473 , \16500 , \16527 , \16554 , \16581 , \16608 , \16635 , \16662 , \16689 , \16716 , \16743 , \16770 , \16797 , \16824 , \16851 );
buf \U$10697 ( \16853 , \15904 );
not \U$10698 ( \16854 , \16853 );
buf \U$10699 ( \16855 , \15892 );
buf \U$10700 ( \16856 , \15893 );
buf \U$10701 ( \16857 , \15894 );
buf \U$10702 ( \16858 , \15897 );
buf \U$10703 ( \16859 , \15901 );
buf \U$10704 ( \16860 , \15904 );
buf \U$10705 ( \16861 , \15904 );
buf \U$10706 ( \16862 , \15904 );
buf \U$10707 ( \16863 , \15904 );
buf \U$10708 ( \16864 , \15904 );
buf \U$10709 ( \16865 , \15904 );
buf \U$10710 ( \16866 , \15904 );
buf \U$10711 ( \16867 , \15904 );
buf \U$10712 ( \16868 , \15904 );
buf \U$10713 ( \16869 , \15904 );
buf \U$10714 ( \16870 , \15904 );
buf \U$10715 ( \16871 , \15904 );
buf \U$10716 ( \16872 , \15904 );
buf \U$10717 ( \16873 , \15904 );
buf \U$10718 ( \16874 , \15904 );
buf \U$10719 ( \16875 , \15904 );
buf \U$10720 ( \16876 , \15904 );
buf \U$10721 ( \16877 , \15904 );
buf \U$10722 ( \16878 , \15904 );
buf \U$10723 ( \16879 , \15904 );
buf \U$10724 ( \16880 , \15904 );
buf \U$10725 ( \16881 , \15904 );
buf \U$10726 ( \16882 , \15904 );
buf \U$10727 ( \16883 , \15904 );
buf \U$10728 ( \16884 , \15904 );
buf \U$10729 ( \16885 , \15891 );
or \U$10730 ( \16886 , \16855 , \16856 , \16857 , \16858 , \16859 , \16860 , \16861 , \16862 , \16863 , \16864 , \16865 , \16866 , \16867 , \16868 , \16869 , \16870 , \16871 , \16872 , \16873 , \16874 , \16875 , \16876 , \16877 , \16878 , \16879 , \16880 , \16881 , \16882 , \16883 , \16884 , \16885 );
nand \U$10731 ( \16887 , \16854 , \16886 );
buf \U$10732 ( \16888 , \16887 );
buf \U$10733 ( \16889 , \15904 );
not \U$10734 ( \16890 , \16889 );
buf \U$10735 ( \16891 , \15901 );
buf \U$10736 ( \16892 , \15904 );
buf \U$10737 ( \16893 , \15904 );
buf \U$10738 ( \16894 , \15904 );
buf \U$10739 ( \16895 , \15904 );
buf \U$10740 ( \16896 , \15904 );
buf \U$10741 ( \16897 , \15904 );
buf \U$10742 ( \16898 , \15904 );
buf \U$10743 ( \16899 , \15904 );
buf \U$10744 ( \16900 , \15904 );
buf \U$10745 ( \16901 , \15904 );
buf \U$10746 ( \16902 , \15904 );
buf \U$10747 ( \16903 , \15904 );
buf \U$10748 ( \16904 , \15904 );
buf \U$10749 ( \16905 , \15904 );
buf \U$10750 ( \16906 , \15904 );
buf \U$10751 ( \16907 , \15904 );
buf \U$10752 ( \16908 , \15904 );
buf \U$10753 ( \16909 , \15904 );
buf \U$10754 ( \16910 , \15904 );
buf \U$10755 ( \16911 , \15904 );
buf \U$10756 ( \16912 , \15904 );
buf \U$10757 ( \16913 , \15904 );
buf \U$10758 ( \16914 , \15904 );
buf \U$10759 ( \16915 , \15904 );
buf \U$10760 ( \16916 , \15904 );
buf \U$10761 ( \16917 , \15897 );
buf \U$10762 ( \16918 , \15891 );
buf \U$10763 ( \16919 , \15892 );
buf \U$10764 ( \16920 , \15893 );
buf \U$10765 ( \16921 , \15894 );
or \U$10766 ( \16922 , \16918 , \16919 , \16920 , \16921 );
and \U$10767 ( \16923 , \16917 , \16922 );
or \U$10768 ( \16924 , \16891 , \16892 , \16893 , \16894 , \16895 , \16896 , \16897 , \16898 , \16899 , \16900 , \16901 , \16902 , \16903 , \16904 , \16905 , \16906 , \16907 , \16908 , \16909 , \16910 , \16911 , \16912 , \16913 , \16914 , \16915 , \16916 , \16923 );
and \U$10769 ( \16925 , \16890 , \16924 );
buf \U$10770 ( \16926 , \16925 );
or \U$10771 ( \16927 , \16888 , \16926 );
_DC g58f4 ( \16928_nG58f4 , \16852 , \16927 );
buf \U$10772 ( \16929 , \16928_nG58f4 );
xor \U$10773 ( \16930 , \16419 , \16929 );
buf \U$10774 ( \16931 , RIb7b9590_247);
and \U$10775 ( \16932 , \7126 , \16445 );
and \U$10776 ( \16933 , \7128 , \16472 );
and \U$10777 ( \16934 , \8338 , \16499 );
and \U$10778 ( \16935 , \8340 , \16526 );
and \U$10779 ( \16936 , \8342 , \16553 );
and \U$10780 ( \16937 , \8344 , \16580 );
and \U$10781 ( \16938 , \8346 , \16607 );
and \U$10782 ( \16939 , \8348 , \16634 );
and \U$10783 ( \16940 , \8350 , \16661 );
and \U$10784 ( \16941 , \8352 , \16688 );
and \U$10785 ( \16942 , \8354 , \16715 );
and \U$10786 ( \16943 , \8356 , \16742 );
and \U$10787 ( \16944 , \8358 , \16769 );
and \U$10788 ( \16945 , \8360 , \16796 );
and \U$10789 ( \16946 , \8362 , \16823 );
and \U$10790 ( \16947 , \8364 , \16850 );
or \U$10791 ( \16948 , \16932 , \16933 , \16934 , \16935 , \16936 , \16937 , \16938 , \16939 , \16940 , \16941 , \16942 , \16943 , \16944 , \16945 , \16946 , \16947 );
_DC g5909 ( \16949_nG5909 , \16948 , \16927 );
buf \U$10792 ( \16950 , \16949_nG5909 );
xor \U$10793 ( \16951 , \16931 , \16950 );
or \U$10794 ( \16952 , \16930 , \16951 );
buf \U$10795 ( \16953 , RIb7b9518_248);
and \U$10796 ( \16954 , \7136 , \16445 );
and \U$10797 ( \16955 , \7138 , \16472 );
and \U$10798 ( \16956 , \8374 , \16499 );
and \U$10799 ( \16957 , \8376 , \16526 );
and \U$10800 ( \16958 , \8378 , \16553 );
and \U$10801 ( \16959 , \8380 , \16580 );
and \U$10802 ( \16960 , \8382 , \16607 );
and \U$10803 ( \16961 , \8384 , \16634 );
and \U$10804 ( \16962 , \8386 , \16661 );
and \U$10805 ( \16963 , \8388 , \16688 );
and \U$10806 ( \16964 , \8390 , \16715 );
and \U$10807 ( \16965 , \8392 , \16742 );
and \U$10808 ( \16966 , \8394 , \16769 );
and \U$10809 ( \16967 , \8396 , \16796 );
and \U$10810 ( \16968 , \8398 , \16823 );
and \U$10811 ( \16969 , \8400 , \16850 );
or \U$10812 ( \16970 , \16954 , \16955 , \16956 , \16957 , \16958 , \16959 , \16960 , \16961 , \16962 , \16963 , \16964 , \16965 , \16966 , \16967 , \16968 , \16969 );
_DC g591f ( \16971_nG591f , \16970 , \16927 );
buf \U$10813 ( \16972 , \16971_nG591f );
xor \U$10814 ( \16973 , \16953 , \16972 );
or \U$10815 ( \16974 , \16952 , \16973 );
buf \U$10816 ( \16975 , RIb7b94a0_249);
and \U$10817 ( \16976 , \7146 , \16445 );
and \U$10818 ( \16977 , \7148 , \16472 );
and \U$10819 ( \16978 , \8410 , \16499 );
and \U$10820 ( \16979 , \8412 , \16526 );
and \U$10821 ( \16980 , \8414 , \16553 );
and \U$10822 ( \16981 , \8416 , \16580 );
and \U$10823 ( \16982 , \8418 , \16607 );
and \U$10824 ( \16983 , \8420 , \16634 );
and \U$10825 ( \16984 , \8422 , \16661 );
and \U$10826 ( \16985 , \8424 , \16688 );
and \U$10827 ( \16986 , \8426 , \16715 );
and \U$10828 ( \16987 , \8428 , \16742 );
and \U$10829 ( \16988 , \8430 , \16769 );
and \U$10830 ( \16989 , \8432 , \16796 );
and \U$10831 ( \16990 , \8434 , \16823 );
and \U$10832 ( \16991 , \8436 , \16850 );
or \U$10833 ( \16992 , \16976 , \16977 , \16978 , \16979 , \16980 , \16981 , \16982 , \16983 , \16984 , \16985 , \16986 , \16987 , \16988 , \16989 , \16990 , \16991 );
_DC g5935 ( \16993_nG5935 , \16992 , \16927 );
buf \U$10834 ( \16994 , \16993_nG5935 );
xor \U$10835 ( \16995 , \16975 , \16994 );
or \U$10836 ( \16996 , \16974 , \16995 );
buf \U$10837 ( \16997 , RIb7b9428_250);
and \U$10838 ( \16998 , \7156 , \16445 );
and \U$10839 ( \16999 , \7158 , \16472 );
and \U$10840 ( \17000 , \8446 , \16499 );
and \U$10841 ( \17001 , \8448 , \16526 );
and \U$10842 ( \17002 , \8450 , \16553 );
and \U$10843 ( \17003 , \8452 , \16580 );
and \U$10844 ( \17004 , \8454 , \16607 );
and \U$10845 ( \17005 , \8456 , \16634 );
and \U$10846 ( \17006 , \8458 , \16661 );
and \U$10847 ( \17007 , \8460 , \16688 );
and \U$10848 ( \17008 , \8462 , \16715 );
and \U$10849 ( \17009 , \8464 , \16742 );
and \U$10850 ( \17010 , \8466 , \16769 );
and \U$10851 ( \17011 , \8468 , \16796 );
and \U$10852 ( \17012 , \8470 , \16823 );
and \U$10853 ( \17013 , \8472 , \16850 );
or \U$10854 ( \17014 , \16998 , \16999 , \17000 , \17001 , \17002 , \17003 , \17004 , \17005 , \17006 , \17007 , \17008 , \17009 , \17010 , \17011 , \17012 , \17013 );
_DC g594b ( \17015_nG594b , \17014 , \16927 );
buf \U$10855 ( \17016 , \17015_nG594b );
xor \U$10856 ( \17017 , \16997 , \17016 );
or \U$10857 ( \17018 , \16996 , \17017 );
buf \U$10858 ( \17019 , RIb7b93b0_251);
and \U$10859 ( \17020 , \7166 , \16445 );
and \U$10860 ( \17021 , \7168 , \16472 );
and \U$10861 ( \17022 , \8482 , \16499 );
and \U$10862 ( \17023 , \8484 , \16526 );
and \U$10863 ( \17024 , \8486 , \16553 );
and \U$10864 ( \17025 , \8488 , \16580 );
and \U$10865 ( \17026 , \8490 , \16607 );
and \U$10866 ( \17027 , \8492 , \16634 );
and \U$10867 ( \17028 , \8494 , \16661 );
and \U$10868 ( \17029 , \8496 , \16688 );
and \U$10869 ( \17030 , \8498 , \16715 );
and \U$10870 ( \17031 , \8500 , \16742 );
and \U$10871 ( \17032 , \8502 , \16769 );
and \U$10872 ( \17033 , \8504 , \16796 );
and \U$10873 ( \17034 , \8506 , \16823 );
and \U$10874 ( \17035 , \8508 , \16850 );
or \U$10875 ( \17036 , \17020 , \17021 , \17022 , \17023 , \17024 , \17025 , \17026 , \17027 , \17028 , \17029 , \17030 , \17031 , \17032 , \17033 , \17034 , \17035 );
_DC g5961 ( \17037_nG5961 , \17036 , \16927 );
buf \U$10876 ( \17038 , \17037_nG5961 );
xor \U$10877 ( \17039 , \17019 , \17038 );
or \U$10878 ( \17040 , \17018 , \17039 );
buf \U$10879 ( \17041 , RIb7af720_252);
and \U$10880 ( \17042 , \7176 , \16445 );
and \U$10881 ( \17043 , \7178 , \16472 );
and \U$10882 ( \17044 , \8518 , \16499 );
and \U$10883 ( \17045 , \8520 , \16526 );
and \U$10884 ( \17046 , \8522 , \16553 );
and \U$10885 ( \17047 , \8524 , \16580 );
and \U$10886 ( \17048 , \8526 , \16607 );
and \U$10887 ( \17049 , \8528 , \16634 );
and \U$10888 ( \17050 , \8530 , \16661 );
and \U$10889 ( \17051 , \8532 , \16688 );
and \U$10890 ( \17052 , \8534 , \16715 );
and \U$10891 ( \17053 , \8536 , \16742 );
and \U$10892 ( \17054 , \8538 , \16769 );
and \U$10893 ( \17055 , \8540 , \16796 );
and \U$10894 ( \17056 , \8542 , \16823 );
and \U$10895 ( \17057 , \8544 , \16850 );
or \U$10896 ( \17058 , \17042 , \17043 , \17044 , \17045 , \17046 , \17047 , \17048 , \17049 , \17050 , \17051 , \17052 , \17053 , \17054 , \17055 , \17056 , \17057 );
_DC g5977 ( \17059_nG5977 , \17058 , \16927 );
buf \U$10897 ( \17060 , \17059_nG5977 );
xor \U$10898 ( \17061 , \17041 , \17060 );
or \U$10899 ( \17062 , \17040 , \17061 );
buf \U$10900 ( \17063 , RIb7af6a8_253);
and \U$10901 ( \17064 , \7186 , \16445 );
and \U$10902 ( \17065 , \7188 , \16472 );
and \U$10903 ( \17066 , \8554 , \16499 );
and \U$10904 ( \17067 , \8556 , \16526 );
and \U$10905 ( \17068 , \8558 , \16553 );
and \U$10906 ( \17069 , \8560 , \16580 );
and \U$10907 ( \17070 , \8562 , \16607 );
and \U$10908 ( \17071 , \8564 , \16634 );
and \U$10909 ( \17072 , \8566 , \16661 );
and \U$10910 ( \17073 , \8568 , \16688 );
and \U$10911 ( \17074 , \8570 , \16715 );
and \U$10912 ( \17075 , \8572 , \16742 );
and \U$10913 ( \17076 , \8574 , \16769 );
and \U$10914 ( \17077 , \8576 , \16796 );
and \U$10915 ( \17078 , \8578 , \16823 );
and \U$10916 ( \17079 , \8580 , \16850 );
or \U$10917 ( \17080 , \17064 , \17065 , \17066 , \17067 , \17068 , \17069 , \17070 , \17071 , \17072 , \17073 , \17074 , \17075 , \17076 , \17077 , \17078 , \17079 );
_DC g598d ( \17081_nG598d , \17080 , \16927 );
buf \U$10918 ( \17082 , \17081_nG598d );
xor \U$10919 ( \17083 , \17063 , \17082 );
or \U$10920 ( \17084 , \17062 , \17083 );
not \U$10921 ( \17085 , \17084 );
buf \U$10922 ( \17086 , \17085 );
and \U$10923 ( \17087 , \16418 , \17086 );
buf \U$10924 ( \17088 , RIb7af630_254);
buf \U$10925 ( \17089 , \15904 );
buf \U$10926 ( \17090 , \15904 );
buf \U$10927 ( \17091 , \15904 );
buf \U$10928 ( \17092 , \15904 );
buf \U$10929 ( \17093 , \15904 );
buf \U$10930 ( \17094 , \15904 );
buf \U$10931 ( \17095 , \15904 );
buf \U$10932 ( \17096 , \15904 );
buf \U$10933 ( \17097 , \15904 );
buf \U$10934 ( \17098 , \15904 );
buf \U$10935 ( \17099 , \15904 );
buf \U$10936 ( \17100 , \15904 );
buf \U$10937 ( \17101 , \15904 );
buf \U$10938 ( \17102 , \15904 );
buf \U$10939 ( \17103 , \15904 );
buf \U$10940 ( \17104 , \15904 );
buf \U$10941 ( \17105 , \15904 );
buf \U$10942 ( \17106 , \15904 );
buf \U$10943 ( \17107 , \15904 );
buf \U$10944 ( \17108 , \15904 );
buf \U$10945 ( \17109 , \15904 );
buf \U$10946 ( \17110 , \15904 );
buf \U$10947 ( \17111 , \15904 );
buf \U$10948 ( \17112 , \15904 );
buf \U$10949 ( \17113 , \15904 );
nor \U$10950 ( \17114 , \15891 , \15892 , \15893 , \15894 , \15898 , \15901 , \15904 , \17089 , \17090 , \17091 , \17092 , \17093 , \17094 , \17095 , \17096 , \17097 , \17098 , \17099 , \17100 , \17101 , \17102 , \17103 , \17104 , \17105 , \17106 , \17107 , \17108 , \17109 , \17110 , \17111 , \17112 , \17113 );
and \U$10951 ( \17115 , \7198 , \17114 );
buf \U$10952 ( \17116 , \15904 );
buf \U$10953 ( \17117 , \15904 );
buf \U$10954 ( \17118 , \15904 );
buf \U$10955 ( \17119 , \15904 );
buf \U$10956 ( \17120 , \15904 );
buf \U$10957 ( \17121 , \15904 );
buf \U$10958 ( \17122 , \15904 );
buf \U$10959 ( \17123 , \15904 );
buf \U$10960 ( \17124 , \15904 );
buf \U$10961 ( \17125 , \15904 );
buf \U$10962 ( \17126 , \15904 );
buf \U$10963 ( \17127 , \15904 );
buf \U$10964 ( \17128 , \15904 );
buf \U$10965 ( \17129 , \15904 );
buf \U$10966 ( \17130 , \15904 );
buf \U$10967 ( \17131 , \15904 );
buf \U$10968 ( \17132 , \15904 );
buf \U$10969 ( \17133 , \15904 );
buf \U$10970 ( \17134 , \15904 );
buf \U$10971 ( \17135 , \15904 );
buf \U$10972 ( \17136 , \15904 );
buf \U$10973 ( \17137 , \15904 );
buf \U$10974 ( \17138 , \15904 );
buf \U$10975 ( \17139 , \15904 );
buf \U$10976 ( \17140 , \15904 );
nor \U$10977 ( \17141 , \15932 , \15933 , \15934 , \15935 , \15897 , \15901 , \15904 , \17116 , \17117 , \17118 , \17119 , \17120 , \17121 , \17122 , \17123 , \17124 , \17125 , \17126 , \17127 , \17128 , \17129 , \17130 , \17131 , \17132 , \17133 , \17134 , \17135 , \17136 , \17137 , \17138 , \17139 , \17140 );
and \U$10978 ( \17142 , \7200 , \17141 );
buf \U$10979 ( \17143 , \15904 );
buf \U$10980 ( \17144 , \15904 );
buf \U$10981 ( \17145 , \15904 );
buf \U$10982 ( \17146 , \15904 );
buf \U$10983 ( \17147 , \15904 );
buf \U$10984 ( \17148 , \15904 );
buf \U$10985 ( \17149 , \15904 );
buf \U$10986 ( \17150 , \15904 );
buf \U$10987 ( \17151 , \15904 );
buf \U$10988 ( \17152 , \15904 );
buf \U$10989 ( \17153 , \15904 );
buf \U$10990 ( \17154 , \15904 );
buf \U$10991 ( \17155 , \15904 );
buf \U$10992 ( \17156 , \15904 );
buf \U$10993 ( \17157 , \15904 );
buf \U$10994 ( \17158 , \15904 );
buf \U$10995 ( \17159 , \15904 );
buf \U$10996 ( \17160 , \15904 );
buf \U$10997 ( \17161 , \15904 );
buf \U$10998 ( \17162 , \15904 );
buf \U$10999 ( \17163 , \15904 );
buf \U$11000 ( \17164 , \15904 );
buf \U$11001 ( \17165 , \15904 );
buf \U$11002 ( \17166 , \15904 );
buf \U$11003 ( \17167 , \15904 );
nor \U$11004 ( \17168 , \15891 , \15933 , \15934 , \15935 , \15897 , \15901 , \15904 , \17143 , \17144 , \17145 , \17146 , \17147 , \17148 , \17149 , \17150 , \17151 , \17152 , \17153 , \17154 , \17155 , \17156 , \17157 , \17158 , \17159 , \17160 , \17161 , \17162 , \17163 , \17164 , \17165 , \17166 , \17167 );
and \U$11005 ( \17169 , \8645 , \17168 );
buf \U$11006 ( \17170 , \15904 );
buf \U$11007 ( \17171 , \15904 );
buf \U$11008 ( \17172 , \15904 );
buf \U$11009 ( \17173 , \15904 );
buf \U$11010 ( \17174 , \15904 );
buf \U$11011 ( \17175 , \15904 );
buf \U$11012 ( \17176 , \15904 );
buf \U$11013 ( \17177 , \15904 );
buf \U$11014 ( \17178 , \15904 );
buf \U$11015 ( \17179 , \15904 );
buf \U$11016 ( \17180 , \15904 );
buf \U$11017 ( \17181 , \15904 );
buf \U$11018 ( \17182 , \15904 );
buf \U$11019 ( \17183 , \15904 );
buf \U$11020 ( \17184 , \15904 );
buf \U$11021 ( \17185 , \15904 );
buf \U$11022 ( \17186 , \15904 );
buf \U$11023 ( \17187 , \15904 );
buf \U$11024 ( \17188 , \15904 );
buf \U$11025 ( \17189 , \15904 );
buf \U$11026 ( \17190 , \15904 );
buf \U$11027 ( \17191 , \15904 );
buf \U$11028 ( \17192 , \15904 );
buf \U$11029 ( \17193 , \15904 );
buf \U$11030 ( \17194 , \15904 );
nor \U$11031 ( \17195 , \15932 , \15892 , \15934 , \15935 , \15897 , \15901 , \15904 , \17170 , \17171 , \17172 , \17173 , \17174 , \17175 , \17176 , \17177 , \17178 , \17179 , \17180 , \17181 , \17182 , \17183 , \17184 , \17185 , \17186 , \17187 , \17188 , \17189 , \17190 , \17191 , \17192 , \17193 , \17194 );
and \U$11032 ( \17196 , \8673 , \17195 );
buf \U$11033 ( \17197 , \15904 );
buf \U$11034 ( \17198 , \15904 );
buf \U$11035 ( \17199 , \15904 );
buf \U$11036 ( \17200 , \15904 );
buf \U$11037 ( \17201 , \15904 );
buf \U$11038 ( \17202 , \15904 );
buf \U$11039 ( \17203 , \15904 );
buf \U$11040 ( \17204 , \15904 );
buf \U$11041 ( \17205 , \15904 );
buf \U$11042 ( \17206 , \15904 );
buf \U$11043 ( \17207 , \15904 );
buf \U$11044 ( \17208 , \15904 );
buf \U$11045 ( \17209 , \15904 );
buf \U$11046 ( \17210 , \15904 );
buf \U$11047 ( \17211 , \15904 );
buf \U$11048 ( \17212 , \15904 );
buf \U$11049 ( \17213 , \15904 );
buf \U$11050 ( \17214 , \15904 );
buf \U$11051 ( \17215 , \15904 );
buf \U$11052 ( \17216 , \15904 );
buf \U$11053 ( \17217 , \15904 );
buf \U$11054 ( \17218 , \15904 );
buf \U$11055 ( \17219 , \15904 );
buf \U$11056 ( \17220 , \15904 );
buf \U$11057 ( \17221 , \15904 );
nor \U$11058 ( \17222 , \15891 , \15892 , \15934 , \15935 , \15897 , \15901 , \15904 , \17197 , \17198 , \17199 , \17200 , \17201 , \17202 , \17203 , \17204 , \17205 , \17206 , \17207 , \17208 , \17209 , \17210 , \17211 , \17212 , \17213 , \17214 , \17215 , \17216 , \17217 , \17218 , \17219 , \17220 , \17221 );
and \U$11059 ( \17223 , \8701 , \17222 );
buf \U$11060 ( \17224 , \15904 );
buf \U$11061 ( \17225 , \15904 );
buf \U$11062 ( \17226 , \15904 );
buf \U$11063 ( \17227 , \15904 );
buf \U$11064 ( \17228 , \15904 );
buf \U$11065 ( \17229 , \15904 );
buf \U$11066 ( \17230 , \15904 );
buf \U$11067 ( \17231 , \15904 );
buf \U$11068 ( \17232 , \15904 );
buf \U$11069 ( \17233 , \15904 );
buf \U$11070 ( \17234 , \15904 );
buf \U$11071 ( \17235 , \15904 );
buf \U$11072 ( \17236 , \15904 );
buf \U$11073 ( \17237 , \15904 );
buf \U$11074 ( \17238 , \15904 );
buf \U$11075 ( \17239 , \15904 );
buf \U$11076 ( \17240 , \15904 );
buf \U$11077 ( \17241 , \15904 );
buf \U$11078 ( \17242 , \15904 );
buf \U$11079 ( \17243 , \15904 );
buf \U$11080 ( \17244 , \15904 );
buf \U$11081 ( \17245 , \15904 );
buf \U$11082 ( \17246 , \15904 );
buf \U$11083 ( \17247 , \15904 );
buf \U$11084 ( \17248 , \15904 );
nor \U$11085 ( \17249 , \15932 , \15933 , \15893 , \15935 , \15897 , \15901 , \15904 , \17224 , \17225 , \17226 , \17227 , \17228 , \17229 , \17230 , \17231 , \17232 , \17233 , \17234 , \17235 , \17236 , \17237 , \17238 , \17239 , \17240 , \17241 , \17242 , \17243 , \17244 , \17245 , \17246 , \17247 , \17248 );
and \U$11086 ( \17250 , \8729 , \17249 );
buf \U$11087 ( \17251 , \15904 );
buf \U$11088 ( \17252 , \15904 );
buf \U$11089 ( \17253 , \15904 );
buf \U$11090 ( \17254 , \15904 );
buf \U$11091 ( \17255 , \15904 );
buf \U$11092 ( \17256 , \15904 );
buf \U$11093 ( \17257 , \15904 );
buf \U$11094 ( \17258 , \15904 );
buf \U$11095 ( \17259 , \15904 );
buf \U$11096 ( \17260 , \15904 );
buf \U$11097 ( \17261 , \15904 );
buf \U$11098 ( \17262 , \15904 );
buf \U$11099 ( \17263 , \15904 );
buf \U$11100 ( \17264 , \15904 );
buf \U$11101 ( \17265 , \15904 );
buf \U$11102 ( \17266 , \15904 );
buf \U$11103 ( \17267 , \15904 );
buf \U$11104 ( \17268 , \15904 );
buf \U$11105 ( \17269 , \15904 );
buf \U$11106 ( \17270 , \15904 );
buf \U$11107 ( \17271 , \15904 );
buf \U$11108 ( \17272 , \15904 );
buf \U$11109 ( \17273 , \15904 );
buf \U$11110 ( \17274 , \15904 );
buf \U$11111 ( \17275 , \15904 );
nor \U$11112 ( \17276 , \15891 , \15933 , \15893 , \15935 , \15897 , \15901 , \15904 , \17251 , \17252 , \17253 , \17254 , \17255 , \17256 , \17257 , \17258 , \17259 , \17260 , \17261 , \17262 , \17263 , \17264 , \17265 , \17266 , \17267 , \17268 , \17269 , \17270 , \17271 , \17272 , \17273 , \17274 , \17275 );
and \U$11113 ( \17277 , \8757 , \17276 );
buf \U$11114 ( \17278 , \15904 );
buf \U$11115 ( \17279 , \15904 );
buf \U$11116 ( \17280 , \15904 );
buf \U$11117 ( \17281 , \15904 );
buf \U$11118 ( \17282 , \15904 );
buf \U$11119 ( \17283 , \15904 );
buf \U$11120 ( \17284 , \15904 );
buf \U$11121 ( \17285 , \15904 );
buf \U$11122 ( \17286 , \15904 );
buf \U$11123 ( \17287 , \15904 );
buf \U$11124 ( \17288 , \15904 );
buf \U$11125 ( \17289 , \15904 );
buf \U$11126 ( \17290 , \15904 );
buf \U$11127 ( \17291 , \15904 );
buf \U$11128 ( \17292 , \15904 );
buf \U$11129 ( \17293 , \15904 );
buf \U$11130 ( \17294 , \15904 );
buf \U$11131 ( \17295 , \15904 );
buf \U$11132 ( \17296 , \15904 );
buf \U$11133 ( \17297 , \15904 );
buf \U$11134 ( \17298 , \15904 );
buf \U$11135 ( \17299 , \15904 );
buf \U$11136 ( \17300 , \15904 );
buf \U$11137 ( \17301 , \15904 );
buf \U$11138 ( \17302 , \15904 );
nor \U$11139 ( \17303 , \15932 , \15892 , \15893 , \15935 , \15897 , \15901 , \15904 , \17278 , \17279 , \17280 , \17281 , \17282 , \17283 , \17284 , \17285 , \17286 , \17287 , \17288 , \17289 , \17290 , \17291 , \17292 , \17293 , \17294 , \17295 , \17296 , \17297 , \17298 , \17299 , \17300 , \17301 , \17302 );
and \U$11140 ( \17304 , \8785 , \17303 );
buf \U$11141 ( \17305 , \15904 );
buf \U$11142 ( \17306 , \15904 );
buf \U$11143 ( \17307 , \15904 );
buf \U$11144 ( \17308 , \15904 );
buf \U$11145 ( \17309 , \15904 );
buf \U$11146 ( \17310 , \15904 );
buf \U$11147 ( \17311 , \15904 );
buf \U$11148 ( \17312 , \15904 );
buf \U$11149 ( \17313 , \15904 );
buf \U$11150 ( \17314 , \15904 );
buf \U$11151 ( \17315 , \15904 );
buf \U$11152 ( \17316 , \15904 );
buf \U$11153 ( \17317 , \15904 );
buf \U$11154 ( \17318 , \15904 );
buf \U$11155 ( \17319 , \15904 );
buf \U$11156 ( \17320 , \15904 );
buf \U$11157 ( \17321 , \15904 );
buf \U$11158 ( \17322 , \15904 );
buf \U$11159 ( \17323 , \15904 );
buf \U$11160 ( \17324 , \15904 );
buf \U$11161 ( \17325 , \15904 );
buf \U$11162 ( \17326 , \15904 );
buf \U$11163 ( \17327 , \15904 );
buf \U$11164 ( \17328 , \15904 );
buf \U$11165 ( \17329 , \15904 );
nor \U$11166 ( \17330 , \15891 , \15892 , \15893 , \15935 , \15897 , \15901 , \15904 , \17305 , \17306 , \17307 , \17308 , \17309 , \17310 , \17311 , \17312 , \17313 , \17314 , \17315 , \17316 , \17317 , \17318 , \17319 , \17320 , \17321 , \17322 , \17323 , \17324 , \17325 , \17326 , \17327 , \17328 , \17329 );
and \U$11167 ( \17331 , \8813 , \17330 );
buf \U$11168 ( \17332 , \15904 );
buf \U$11169 ( \17333 , \15904 );
buf \U$11170 ( \17334 , \15904 );
buf \U$11171 ( \17335 , \15904 );
buf \U$11172 ( \17336 , \15904 );
buf \U$11173 ( \17337 , \15904 );
buf \U$11174 ( \17338 , \15904 );
buf \U$11175 ( \17339 , \15904 );
buf \U$11176 ( \17340 , \15904 );
buf \U$11177 ( \17341 , \15904 );
buf \U$11178 ( \17342 , \15904 );
buf \U$11179 ( \17343 , \15904 );
buf \U$11180 ( \17344 , \15904 );
buf \U$11181 ( \17345 , \15904 );
buf \U$11182 ( \17346 , \15904 );
buf \U$11183 ( \17347 , \15904 );
buf \U$11184 ( \17348 , \15904 );
buf \U$11185 ( \17349 , \15904 );
buf \U$11186 ( \17350 , \15904 );
buf \U$11187 ( \17351 , \15904 );
buf \U$11188 ( \17352 , \15904 );
buf \U$11189 ( \17353 , \15904 );
buf \U$11190 ( \17354 , \15904 );
buf \U$11191 ( \17355 , \15904 );
buf \U$11192 ( \17356 , \15904 );
nor \U$11193 ( \17357 , \15932 , \15933 , \15934 , \15894 , \15897 , \15901 , \15904 , \17332 , \17333 , \17334 , \17335 , \17336 , \17337 , \17338 , \17339 , \17340 , \17341 , \17342 , \17343 , \17344 , \17345 , \17346 , \17347 , \17348 , \17349 , \17350 , \17351 , \17352 , \17353 , \17354 , \17355 , \17356 );
and \U$11194 ( \17358 , \8841 , \17357 );
buf \U$11195 ( \17359 , \15904 );
buf \U$11196 ( \17360 , \15904 );
buf \U$11197 ( \17361 , \15904 );
buf \U$11198 ( \17362 , \15904 );
buf \U$11199 ( \17363 , \15904 );
buf \U$11200 ( \17364 , \15904 );
buf \U$11201 ( \17365 , \15904 );
buf \U$11202 ( \17366 , \15904 );
buf \U$11203 ( \17367 , \15904 );
buf \U$11204 ( \17368 , \15904 );
buf \U$11205 ( \17369 , \15904 );
buf \U$11206 ( \17370 , \15904 );
buf \U$11207 ( \17371 , \15904 );
buf \U$11208 ( \17372 , \15904 );
buf \U$11209 ( \17373 , \15904 );
buf \U$11210 ( \17374 , \15904 );
buf \U$11211 ( \17375 , \15904 );
buf \U$11212 ( \17376 , \15904 );
buf \U$11213 ( \17377 , \15904 );
buf \U$11214 ( \17378 , \15904 );
buf \U$11215 ( \17379 , \15904 );
buf \U$11216 ( \17380 , \15904 );
buf \U$11217 ( \17381 , \15904 );
buf \U$11218 ( \17382 , \15904 );
buf \U$11219 ( \17383 , \15904 );
nor \U$11220 ( \17384 , \15891 , \15933 , \15934 , \15894 , \15897 , \15901 , \15904 , \17359 , \17360 , \17361 , \17362 , \17363 , \17364 , \17365 , \17366 , \17367 , \17368 , \17369 , \17370 , \17371 , \17372 , \17373 , \17374 , \17375 , \17376 , \17377 , \17378 , \17379 , \17380 , \17381 , \17382 , \17383 );
and \U$11221 ( \17385 , \8869 , \17384 );
buf \U$11222 ( \17386 , \15904 );
buf \U$11223 ( \17387 , \15904 );
buf \U$11224 ( \17388 , \15904 );
buf \U$11225 ( \17389 , \15904 );
buf \U$11226 ( \17390 , \15904 );
buf \U$11227 ( \17391 , \15904 );
buf \U$11228 ( \17392 , \15904 );
buf \U$11229 ( \17393 , \15904 );
buf \U$11230 ( \17394 , \15904 );
buf \U$11231 ( \17395 , \15904 );
buf \U$11232 ( \17396 , \15904 );
buf \U$11233 ( \17397 , \15904 );
buf \U$11234 ( \17398 , \15904 );
buf \U$11235 ( \17399 , \15904 );
buf \U$11236 ( \17400 , \15904 );
buf \U$11237 ( \17401 , \15904 );
buf \U$11238 ( \17402 , \15904 );
buf \U$11239 ( \17403 , \15904 );
buf \U$11240 ( \17404 , \15904 );
buf \U$11241 ( \17405 , \15904 );
buf \U$11242 ( \17406 , \15904 );
buf \U$11243 ( \17407 , \15904 );
buf \U$11244 ( \17408 , \15904 );
buf \U$11245 ( \17409 , \15904 );
buf \U$11246 ( \17410 , \15904 );
nor \U$11247 ( \17411 , \15932 , \15892 , \15934 , \15894 , \15897 , \15901 , \15904 , \17386 , \17387 , \17388 , \17389 , \17390 , \17391 , \17392 , \17393 , \17394 , \17395 , \17396 , \17397 , \17398 , \17399 , \17400 , \17401 , \17402 , \17403 , \17404 , \17405 , \17406 , \17407 , \17408 , \17409 , \17410 );
and \U$11248 ( \17412 , \8897 , \17411 );
buf \U$11249 ( \17413 , \15904 );
buf \U$11250 ( \17414 , \15904 );
buf \U$11251 ( \17415 , \15904 );
buf \U$11252 ( \17416 , \15904 );
buf \U$11253 ( \17417 , \15904 );
buf \U$11254 ( \17418 , \15904 );
buf \U$11255 ( \17419 , \15904 );
buf \U$11256 ( \17420 , \15904 );
buf \U$11257 ( \17421 , \15904 );
buf \U$11258 ( \17422 , \15904 );
buf \U$11259 ( \17423 , \15904 );
buf \U$11260 ( \17424 , \15904 );
buf \U$11261 ( \17425 , \15904 );
buf \U$11262 ( \17426 , \15904 );
buf \U$11263 ( \17427 , \15904 );
buf \U$11264 ( \17428 , \15904 );
buf \U$11265 ( \17429 , \15904 );
buf \U$11266 ( \17430 , \15904 );
buf \U$11267 ( \17431 , \15904 );
buf \U$11268 ( \17432 , \15904 );
buf \U$11269 ( \17433 , \15904 );
buf \U$11270 ( \17434 , \15904 );
buf \U$11271 ( \17435 , \15904 );
buf \U$11272 ( \17436 , \15904 );
buf \U$11273 ( \17437 , \15904 );
nor \U$11274 ( \17438 , \15891 , \15892 , \15934 , \15894 , \15897 , \15901 , \15904 , \17413 , \17414 , \17415 , \17416 , \17417 , \17418 , \17419 , \17420 , \17421 , \17422 , \17423 , \17424 , \17425 , \17426 , \17427 , \17428 , \17429 , \17430 , \17431 , \17432 , \17433 , \17434 , \17435 , \17436 , \17437 );
and \U$11275 ( \17439 , \8925 , \17438 );
buf \U$11276 ( \17440 , \15904 );
buf \U$11277 ( \17441 , \15904 );
buf \U$11278 ( \17442 , \15904 );
buf \U$11279 ( \17443 , \15904 );
buf \U$11280 ( \17444 , \15904 );
buf \U$11281 ( \17445 , \15904 );
buf \U$11282 ( \17446 , \15904 );
buf \U$11283 ( \17447 , \15904 );
buf \U$11284 ( \17448 , \15904 );
buf \U$11285 ( \17449 , \15904 );
buf \U$11286 ( \17450 , \15904 );
buf \U$11287 ( \17451 , \15904 );
buf \U$11288 ( \17452 , \15904 );
buf \U$11289 ( \17453 , \15904 );
buf \U$11290 ( \17454 , \15904 );
buf \U$11291 ( \17455 , \15904 );
buf \U$11292 ( \17456 , \15904 );
buf \U$11293 ( \17457 , \15904 );
buf \U$11294 ( \17458 , \15904 );
buf \U$11295 ( \17459 , \15904 );
buf \U$11296 ( \17460 , \15904 );
buf \U$11297 ( \17461 , \15904 );
buf \U$11298 ( \17462 , \15904 );
buf \U$11299 ( \17463 , \15904 );
buf \U$11300 ( \17464 , \15904 );
nor \U$11301 ( \17465 , \15932 , \15933 , \15893 , \15894 , \15897 , \15901 , \15904 , \17440 , \17441 , \17442 , \17443 , \17444 , \17445 , \17446 , \17447 , \17448 , \17449 , \17450 , \17451 , \17452 , \17453 , \17454 , \17455 , \17456 , \17457 , \17458 , \17459 , \17460 , \17461 , \17462 , \17463 , \17464 );
and \U$11302 ( \17466 , \8953 , \17465 );
buf \U$11303 ( \17467 , \15904 );
buf \U$11304 ( \17468 , \15904 );
buf \U$11305 ( \17469 , \15904 );
buf \U$11306 ( \17470 , \15904 );
buf \U$11307 ( \17471 , \15904 );
buf \U$11308 ( \17472 , \15904 );
buf \U$11309 ( \17473 , \15904 );
buf \U$11310 ( \17474 , \15904 );
buf \U$11311 ( \17475 , \15904 );
buf \U$11312 ( \17476 , \15904 );
buf \U$11313 ( \17477 , \15904 );
buf \U$11314 ( \17478 , \15904 );
buf \U$11315 ( \17479 , \15904 );
buf \U$11316 ( \17480 , \15904 );
buf \U$11317 ( \17481 , \15904 );
buf \U$11318 ( \17482 , \15904 );
buf \U$11319 ( \17483 , \15904 );
buf \U$11320 ( \17484 , \15904 );
buf \U$11321 ( \17485 , \15904 );
buf \U$11322 ( \17486 , \15904 );
buf \U$11323 ( \17487 , \15904 );
buf \U$11324 ( \17488 , \15904 );
buf \U$11325 ( \17489 , \15904 );
buf \U$11326 ( \17490 , \15904 );
buf \U$11327 ( \17491 , \15904 );
nor \U$11328 ( \17492 , \15891 , \15933 , \15893 , \15894 , \15897 , \15901 , \15904 , \17467 , \17468 , \17469 , \17470 , \17471 , \17472 , \17473 , \17474 , \17475 , \17476 , \17477 , \17478 , \17479 , \17480 , \17481 , \17482 , \17483 , \17484 , \17485 , \17486 , \17487 , \17488 , \17489 , \17490 , \17491 );
and \U$11329 ( \17493 , \8981 , \17492 );
buf \U$11330 ( \17494 , \15904 );
buf \U$11331 ( \17495 , \15904 );
buf \U$11332 ( \17496 , \15904 );
buf \U$11333 ( \17497 , \15904 );
buf \U$11334 ( \17498 , \15904 );
buf \U$11335 ( \17499 , \15904 );
buf \U$11336 ( \17500 , \15904 );
buf \U$11337 ( \17501 , \15904 );
buf \U$11338 ( \17502 , \15904 );
buf \U$11339 ( \17503 , \15904 );
buf \U$11340 ( \17504 , \15904 );
buf \U$11341 ( \17505 , \15904 );
buf \U$11342 ( \17506 , \15904 );
buf \U$11343 ( \17507 , \15904 );
buf \U$11344 ( \17508 , \15904 );
buf \U$11345 ( \17509 , \15904 );
buf \U$11346 ( \17510 , \15904 );
buf \U$11347 ( \17511 , \15904 );
buf \U$11348 ( \17512 , \15904 );
buf \U$11349 ( \17513 , \15904 );
buf \U$11350 ( \17514 , \15904 );
buf \U$11351 ( \17515 , \15904 );
buf \U$11352 ( \17516 , \15904 );
buf \U$11353 ( \17517 , \15904 );
buf \U$11354 ( \17518 , \15904 );
nor \U$11355 ( \17519 , \15932 , \15892 , \15893 , \15894 , \15897 , \15901 , \15904 , \17494 , \17495 , \17496 , \17497 , \17498 , \17499 , \17500 , \17501 , \17502 , \17503 , \17504 , \17505 , \17506 , \17507 , \17508 , \17509 , \17510 , \17511 , \17512 , \17513 , \17514 , \17515 , \17516 , \17517 , \17518 );
and \U$11356 ( \17520 , \9009 , \17519 );
or \U$11357 ( \17521 , \17115 , \17142 , \17169 , \17196 , \17223 , \17250 , \17277 , \17304 , \17331 , \17358 , \17385 , \17412 , \17439 , \17466 , \17493 , \17520 );
buf \U$11358 ( \17522 , \15904 );
not \U$11359 ( \17523 , \17522 );
buf \U$11360 ( \17524 , \15892 );
buf \U$11361 ( \17525 , \15893 );
buf \U$11362 ( \17526 , \15894 );
buf \U$11363 ( \17527 , \15897 );
buf \U$11364 ( \17528 , \15901 );
buf \U$11365 ( \17529 , \15904 );
buf \U$11366 ( \17530 , \15904 );
buf \U$11367 ( \17531 , \15904 );
buf \U$11368 ( \17532 , \15904 );
buf \U$11369 ( \17533 , \15904 );
buf \U$11370 ( \17534 , \15904 );
buf \U$11371 ( \17535 , \15904 );
buf \U$11372 ( \17536 , \15904 );
buf \U$11373 ( \17537 , \15904 );
buf \U$11374 ( \17538 , \15904 );
buf \U$11375 ( \17539 , \15904 );
buf \U$11376 ( \17540 , \15904 );
buf \U$11377 ( \17541 , \15904 );
buf \U$11378 ( \17542 , \15904 );
buf \U$11379 ( \17543 , \15904 );
buf \U$11380 ( \17544 , \15904 );
buf \U$11381 ( \17545 , \15904 );
buf \U$11382 ( \17546 , \15904 );
buf \U$11383 ( \17547 , \15904 );
buf \U$11384 ( \17548 , \15904 );
buf \U$11385 ( \17549 , \15904 );
buf \U$11386 ( \17550 , \15904 );
buf \U$11387 ( \17551 , \15904 );
buf \U$11388 ( \17552 , \15904 );
buf \U$11389 ( \17553 , \15904 );
buf \U$11390 ( \17554 , \15891 );
or \U$11391 ( \17555 , \17524 , \17525 , \17526 , \17527 , \17528 , \17529 , \17530 , \17531 , \17532 , \17533 , \17534 , \17535 , \17536 , \17537 , \17538 , \17539 , \17540 , \17541 , \17542 , \17543 , \17544 , \17545 , \17546 , \17547 , \17548 , \17549 , \17550 , \17551 , \17552 , \17553 , \17554 );
nand \U$11392 ( \17556 , \17523 , \17555 );
buf \U$11393 ( \17557 , \17556 );
buf \U$11394 ( \17558 , \15904 );
not \U$11395 ( \17559 , \17558 );
buf \U$11396 ( \17560 , \15901 );
buf \U$11397 ( \17561 , \15904 );
buf \U$11398 ( \17562 , \15904 );
buf \U$11399 ( \17563 , \15904 );
buf \U$11400 ( \17564 , \15904 );
buf \U$11401 ( \17565 , \15904 );
buf \U$11402 ( \17566 , \15904 );
buf \U$11403 ( \17567 , \15904 );
buf \U$11404 ( \17568 , \15904 );
buf \U$11405 ( \17569 , \15904 );
buf \U$11406 ( \17570 , \15904 );
buf \U$11407 ( \17571 , \15904 );
buf \U$11408 ( \17572 , \15904 );
buf \U$11409 ( \17573 , \15904 );
buf \U$11410 ( \17574 , \15904 );
buf \U$11411 ( \17575 , \15904 );
buf \U$11412 ( \17576 , \15904 );
buf \U$11413 ( \17577 , \15904 );
buf \U$11414 ( \17578 , \15904 );
buf \U$11415 ( \17579 , \15904 );
buf \U$11416 ( \17580 , \15904 );
buf \U$11417 ( \17581 , \15904 );
buf \U$11418 ( \17582 , \15904 );
buf \U$11419 ( \17583 , \15904 );
buf \U$11420 ( \17584 , \15904 );
buf \U$11421 ( \17585 , \15904 );
buf \U$11422 ( \17586 , \15897 );
buf \U$11423 ( \17587 , \15891 );
buf \U$11424 ( \17588 , \15892 );
buf \U$11425 ( \17589 , \15893 );
buf \U$11426 ( \17590 , \15894 );
or \U$11427 ( \17591 , \17587 , \17588 , \17589 , \17590 );
and \U$11428 ( \17592 , \17586 , \17591 );
or \U$11429 ( \17593 , \17560 , \17561 , \17562 , \17563 , \17564 , \17565 , \17566 , \17567 , \17568 , \17569 , \17570 , \17571 , \17572 , \17573 , \17574 , \17575 , \17576 , \17577 , \17578 , \17579 , \17580 , \17581 , \17582 , \17583 , \17584 , \17585 , \17592 );
and \U$11430 ( \17594 , \17559 , \17593 );
buf \U$11431 ( \17595 , \17594 );
or \U$11432 ( \17596 , \17557 , \17595 );
_DC g5b91 ( \17597_nG5b91 , \17521 , \17596 );
buf \U$11433 ( \17598 , \17597_nG5b91 );
xor \U$11434 ( \17599 , \17088 , \17598 );
buf \U$11435 ( \17600 , RIb7af5b8_255);
and \U$11436 ( \17601 , \7207 , \17114 );
and \U$11437 ( \17602 , \7209 , \17141 );
and \U$11438 ( \17603 , \9119 , \17168 );
and \U$11439 ( \17604 , \9121 , \17195 );
and \U$11440 ( \17605 , \9123 , \17222 );
and \U$11441 ( \17606 , \9125 , \17249 );
and \U$11442 ( \17607 , \9127 , \17276 );
and \U$11443 ( \17608 , \9129 , \17303 );
and \U$11444 ( \17609 , \9131 , \17330 );
and \U$11445 ( \17610 , \9133 , \17357 );
and \U$11446 ( \17611 , \9135 , \17384 );
and \U$11447 ( \17612 , \9137 , \17411 );
and \U$11448 ( \17613 , \9139 , \17438 );
and \U$11449 ( \17614 , \9141 , \17465 );
and \U$11450 ( \17615 , \9143 , \17492 );
and \U$11451 ( \17616 , \9145 , \17519 );
or \U$11452 ( \17617 , \17601 , \17602 , \17603 , \17604 , \17605 , \17606 , \17607 , \17608 , \17609 , \17610 , \17611 , \17612 , \17613 , \17614 , \17615 , \17616 );
_DC g5ba6 ( \17618_nG5ba6 , \17617 , \17596 );
buf \U$11453 ( \17619 , \17618_nG5ba6 );
xor \U$11454 ( \17620 , \17600 , \17619 );
or \U$11455 ( \17621 , \17599 , \17620 );
buf \U$11456 ( \17622 , RIb7af540_256);
and \U$11457 ( \17623 , \7217 , \17114 );
and \U$11458 ( \17624 , \7219 , \17141 );
and \U$11459 ( \17625 , \9155 , \17168 );
and \U$11460 ( \17626 , \9157 , \17195 );
and \U$11461 ( \17627 , \9159 , \17222 );
and \U$11462 ( \17628 , \9161 , \17249 );
and \U$11463 ( \17629 , \9163 , \17276 );
and \U$11464 ( \17630 , \9165 , \17303 );
and \U$11465 ( \17631 , \9167 , \17330 );
and \U$11466 ( \17632 , \9169 , \17357 );
and \U$11467 ( \17633 , \9171 , \17384 );
and \U$11468 ( \17634 , \9173 , \17411 );
and \U$11469 ( \17635 , \9175 , \17438 );
and \U$11470 ( \17636 , \9177 , \17465 );
and \U$11471 ( \17637 , \9179 , \17492 );
and \U$11472 ( \17638 , \9181 , \17519 );
or \U$11473 ( \17639 , \17623 , \17624 , \17625 , \17626 , \17627 , \17628 , \17629 , \17630 , \17631 , \17632 , \17633 , \17634 , \17635 , \17636 , \17637 , \17638 );
_DC g5bbc ( \17640_nG5bbc , \17639 , \17596 );
buf \U$11474 ( \17641 , \17640_nG5bbc );
xor \U$11475 ( \17642 , \17622 , \17641 );
or \U$11476 ( \17643 , \17621 , \17642 );
buf \U$11477 ( \17644 , RIb7af4c8_257);
and \U$11478 ( \17645 , \7227 , \17114 );
and \U$11479 ( \17646 , \7229 , \17141 );
and \U$11480 ( \17647 , \9191 , \17168 );
and \U$11481 ( \17648 , \9193 , \17195 );
and \U$11482 ( \17649 , \9195 , \17222 );
and \U$11483 ( \17650 , \9197 , \17249 );
and \U$11484 ( \17651 , \9199 , \17276 );
and \U$11485 ( \17652 , \9201 , \17303 );
and \U$11486 ( \17653 , \9203 , \17330 );
and \U$11487 ( \17654 , \9205 , \17357 );
and \U$11488 ( \17655 , \9207 , \17384 );
and \U$11489 ( \17656 , \9209 , \17411 );
and \U$11490 ( \17657 , \9211 , \17438 );
and \U$11491 ( \17658 , \9213 , \17465 );
and \U$11492 ( \17659 , \9215 , \17492 );
and \U$11493 ( \17660 , \9217 , \17519 );
or \U$11494 ( \17661 , \17645 , \17646 , \17647 , \17648 , \17649 , \17650 , \17651 , \17652 , \17653 , \17654 , \17655 , \17656 , \17657 , \17658 , \17659 , \17660 );
_DC g5bd2 ( \17662_nG5bd2 , \17661 , \17596 );
buf \U$11495 ( \17663 , \17662_nG5bd2 );
xor \U$11496 ( \17664 , \17644 , \17663 );
or \U$11497 ( \17665 , \17643 , \17664 );
buf \U$11498 ( \17666 , RIb7af450_258);
and \U$11499 ( \17667 , \7237 , \17114 );
and \U$11500 ( \17668 , \7239 , \17141 );
and \U$11501 ( \17669 , \9227 , \17168 );
and \U$11502 ( \17670 , \9229 , \17195 );
and \U$11503 ( \17671 , \9231 , \17222 );
and \U$11504 ( \17672 , \9233 , \17249 );
and \U$11505 ( \17673 , \9235 , \17276 );
and \U$11506 ( \17674 , \9237 , \17303 );
and \U$11507 ( \17675 , \9239 , \17330 );
and \U$11508 ( \17676 , \9241 , \17357 );
and \U$11509 ( \17677 , \9243 , \17384 );
and \U$11510 ( \17678 , \9245 , \17411 );
and \U$11511 ( \17679 , \9247 , \17438 );
and \U$11512 ( \17680 , \9249 , \17465 );
and \U$11513 ( \17681 , \9251 , \17492 );
and \U$11514 ( \17682 , \9253 , \17519 );
or \U$11515 ( \17683 , \17667 , \17668 , \17669 , \17670 , \17671 , \17672 , \17673 , \17674 , \17675 , \17676 , \17677 , \17678 , \17679 , \17680 , \17681 , \17682 );
_DC g5be8 ( \17684_nG5be8 , \17683 , \17596 );
buf \U$11516 ( \17685 , \17684_nG5be8 );
xor \U$11517 ( \17686 , \17666 , \17685 );
or \U$11518 ( \17687 , \17665 , \17686 );
buf \U$11519 ( \17688 , RIb7af3d8_259);
and \U$11520 ( \17689 , \7247 , \17114 );
and \U$11521 ( \17690 , \7249 , \17141 );
and \U$11522 ( \17691 , \9263 , \17168 );
and \U$11523 ( \17692 , \9265 , \17195 );
and \U$11524 ( \17693 , \9267 , \17222 );
and \U$11525 ( \17694 , \9269 , \17249 );
and \U$11526 ( \17695 , \9271 , \17276 );
and \U$11527 ( \17696 , \9273 , \17303 );
and \U$11528 ( \17697 , \9275 , \17330 );
and \U$11529 ( \17698 , \9277 , \17357 );
and \U$11530 ( \17699 , \9279 , \17384 );
and \U$11531 ( \17700 , \9281 , \17411 );
and \U$11532 ( \17701 , \9283 , \17438 );
and \U$11533 ( \17702 , \9285 , \17465 );
and \U$11534 ( \17703 , \9287 , \17492 );
and \U$11535 ( \17704 , \9289 , \17519 );
or \U$11536 ( \17705 , \17689 , \17690 , \17691 , \17692 , \17693 , \17694 , \17695 , \17696 , \17697 , \17698 , \17699 , \17700 , \17701 , \17702 , \17703 , \17704 );
_DC g5bfe ( \17706_nG5bfe , \17705 , \17596 );
buf \U$11537 ( \17707 , \17706_nG5bfe );
xor \U$11538 ( \17708 , \17688 , \17707 );
or \U$11539 ( \17709 , \17687 , \17708 );
buf \U$11540 ( \17710 , RIb7a5bf8_260);
and \U$11541 ( \17711 , \7257 , \17114 );
and \U$11542 ( \17712 , \7259 , \17141 );
and \U$11543 ( \17713 , \9299 , \17168 );
and \U$11544 ( \17714 , \9301 , \17195 );
and \U$11545 ( \17715 , \9303 , \17222 );
and \U$11546 ( \17716 , \9305 , \17249 );
and \U$11547 ( \17717 , \9307 , \17276 );
and \U$11548 ( \17718 , \9309 , \17303 );
and \U$11549 ( \17719 , \9311 , \17330 );
and \U$11550 ( \17720 , \9313 , \17357 );
and \U$11551 ( \17721 , \9315 , \17384 );
and \U$11552 ( \17722 , \9317 , \17411 );
and \U$11553 ( \17723 , \9319 , \17438 );
and \U$11554 ( \17724 , \9321 , \17465 );
and \U$11555 ( \17725 , \9323 , \17492 );
and \U$11556 ( \17726 , \9325 , \17519 );
or \U$11557 ( \17727 , \17711 , \17712 , \17713 , \17714 , \17715 , \17716 , \17717 , \17718 , \17719 , \17720 , \17721 , \17722 , \17723 , \17724 , \17725 , \17726 );
_DC g5c14 ( \17728_nG5c14 , \17727 , \17596 );
buf \U$11558 ( \17729 , \17728_nG5c14 );
xor \U$11559 ( \17730 , \17710 , \17729 );
or \U$11560 ( \17731 , \17709 , \17730 );
buf \U$11561 ( \17732 , RIb7a0c48_261);
and \U$11562 ( \17733 , \7267 , \17114 );
and \U$11563 ( \17734 , \7269 , \17141 );
and \U$11564 ( \17735 , \9335 , \17168 );
and \U$11565 ( \17736 , \9337 , \17195 );
and \U$11566 ( \17737 , \9339 , \17222 );
and \U$11567 ( \17738 , \9341 , \17249 );
and \U$11568 ( \17739 , \9343 , \17276 );
and \U$11569 ( \17740 , \9345 , \17303 );
and \U$11570 ( \17741 , \9347 , \17330 );
and \U$11571 ( \17742 , \9349 , \17357 );
and \U$11572 ( \17743 , \9351 , \17384 );
and \U$11573 ( \17744 , \9353 , \17411 );
and \U$11574 ( \17745 , \9355 , \17438 );
and \U$11575 ( \17746 , \9357 , \17465 );
and \U$11576 ( \17747 , \9359 , \17492 );
and \U$11577 ( \17748 , \9361 , \17519 );
or \U$11578 ( \17749 , \17733 , \17734 , \17735 , \17736 , \17737 , \17738 , \17739 , \17740 , \17741 , \17742 , \17743 , \17744 , \17745 , \17746 , \17747 , \17748 );
_DC g5c2a ( \17750_nG5c2a , \17749 , \17596 );
buf \U$11579 ( \17751 , \17750_nG5c2a );
xor \U$11580 ( \17752 , \17732 , \17751 );
or \U$11581 ( \17753 , \17731 , \17752 );
not \U$11582 ( \17754 , \17753 );
buf \U$11583 ( \17755 , \17754 );
and \U$11584 ( \17756 , \17087 , \17755 );
_HMUX g5c31 ( \17757_nG5c31 , \15642_nG53e6 , \15891 , \17756 );
buf \U$11585 ( \17758 , \15663 );
buf \U$11586 ( \17759 , \15660 );
buf \U$11587 ( \17760 , \15645 );
buf \U$11588 ( \17761 , \15648 );
buf \U$11589 ( \17762 , \15652 );
buf \U$11590 ( \17763 , \15656 );
or \U$11591 ( \17764 , \17760 , \17761 , \17762 , \17763 );
and \U$11592 ( \17765 , \17759 , \17764 );
or \U$11593 ( \17766 , \17758 , \17765 );
buf \U$11594 ( \17767 , \17766 );
_HMUX g5c3c ( \17768_nG5c3c , \15890_nG54de , \17757_nG5c31 , \17767 );
buf \U$11595 ( \17769 , RIe5319e0_6884);
buf \U$11597 ( \17770 , \17769 );
buf \U$11598 ( \17771 , RIe549ef0_6842);
not \U$11599 ( \17772 , \17771 );
buf \U$11600 ( \17773 , \17772 );
buf \U$11601 ( \17774 , RIe549770_6843);
xor \U$11602 ( \17775 , \17774 , \17771 );
buf \U$11603 ( \17776 , \17775 );
buf \U$11604 ( \17777 , RIe548ff0_6844);
and \U$11605 ( \17778 , \17774 , \17771 );
xnor \U$11606 ( \17779 , \17777 , \17778 );
buf \U$11607 ( \17780 , \17779 );
buf \U$11608 ( \17781 , RIea91330_6888);
or \U$11609 ( \17782 , \17777 , \17778 );
xor \U$11610 ( \17783 , \17781 , \17782 );
buf \U$11611 ( \17784 , \17783 );
not \U$11612 ( \17785 , \17784 );
and \U$11613 ( \17786 , \17781 , \17782 );
buf \U$11614 ( \17787 , \17786 );
nor \U$11615 ( \17788 , \17770 , \17773 , \17776 , \17780 , \17785 , \17787 );
and \U$11616 ( \17789 , RIe5329d0_6883, \17788 );
not \U$11617 ( \17790 , \17787 );
and \U$11618 ( \17791 , \17770 , \17773 , \17776 , \17780 , \17785 , \17790 );
and \U$11619 ( \17792 , RIeb72150_6905, \17791 );
not \U$11620 ( \17793 , \17770 );
and \U$11621 ( \17794 , \17793 , \17773 , \17776 , \17780 , \17785 , \17790 );
and \U$11622 ( \17795 , RIeab80c0_6897, \17794 );
not \U$11623 ( \17796 , \17773 );
and \U$11624 ( \17797 , \17770 , \17796 , \17776 , \17780 , \17785 , \17790 );
and \U$11625 ( \17798 , RIe5331c8_6882, \17797 );
and \U$11626 ( \17799 , \17793 , \17796 , \17776 , \17780 , \17785 , \17790 );
and \U$11627 ( \17800 , RIe5339c0_6881, \17799 );
not \U$11628 ( \17801 , \17776 );
and \U$11629 ( \17802 , \17770 , \17773 , \17801 , \17780 , \17785 , \17790 );
and \U$11630 ( \17803 , RIeab87c8_6898, \17802 );
and \U$11631 ( \17804 , \17793 , \17773 , \17801 , \17780 , \17785 , \17790 );
and \U$11632 ( \17805 , RIe5341b8_6880, \17804 );
or \U$11642 ( \17806 , \17789 , \17792 , \17795 , \17798 , \17800 , \17803 , \17805 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
buf \U$11644 ( \17807 , \17787 );
buf \U$11645 ( \17808 , \17784 );
buf \U$11646 ( \17809 , \17770 );
buf \U$11647 ( \17810 , \17773 );
buf \U$11648 ( \17811 , \17776 );
buf \U$11649 ( \17812 , \17780 );
or \U$11650 ( \17813 , \17809 , \17810 , \17811 , \17812 );
and \U$11651 ( \17814 , \17808 , \17813 );
or \U$11652 ( \17815 , \17807 , \17814 );
buf \U$11653 ( \17816 , \17815 );
or \U$11654 ( \17817 , 1'b0 , \17816 );
_DC g5c6f ( \17818_nG5c6f , \17806 , \17817 );
not \U$11655 ( \17819 , \17818_nG5c6f );
buf \U$11656 ( \17820 , RIb7b9608_246);
and \U$11657 ( \17821 , \7117 , \17788 );
and \U$11658 ( \17822 , \7119 , \17791 );
and \U$11659 ( \17823 , \7864 , \17794 );
and \U$11660 ( \17824 , \7892 , \17797 );
and \U$11661 ( \17825 , \7920 , \17799 );
and \U$11662 ( \17826 , \7948 , \17802 );
and \U$11663 ( \17827 , \7976 , \17804 );
or \U$11673 ( \17828 , \17821 , \17822 , \17823 , \17824 , \17825 , \17826 , \17827 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5c7a ( \17829_nG5c7a , \17828 , \17817 );
buf \U$11674 ( \17830 , \17829_nG5c7a );
xor \U$11675 ( \17831 , \17820 , \17830 );
buf \U$11676 ( \17832 , RIb7b9590_247);
and \U$11677 ( \17833 , \7126 , \17788 );
and \U$11678 ( \17834 , \7128 , \17791 );
and \U$11679 ( \17835 , \8338 , \17794 );
and \U$11680 ( \17836 , \8340 , \17797 );
and \U$11681 ( \17837 , \8342 , \17799 );
and \U$11682 ( \17838 , \8344 , \17802 );
and \U$11683 ( \17839 , \8346 , \17804 );
or \U$11693 ( \17840 , \17833 , \17834 , \17835 , \17836 , \17837 , \17838 , \17839 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5c86 ( \17841_nG5c86 , \17840 , \17817 );
buf \U$11694 ( \17842 , \17841_nG5c86 );
xor \U$11695 ( \17843 , \17832 , \17842 );
or \U$11696 ( \17844 , \17831 , \17843 );
buf \U$11697 ( \17845 , RIb7b9518_248);
and \U$11698 ( \17846 , \7136 , \17788 );
and \U$11699 ( \17847 , \7138 , \17791 );
and \U$11700 ( \17848 , \8374 , \17794 );
and \U$11701 ( \17849 , \8376 , \17797 );
and \U$11702 ( \17850 , \8378 , \17799 );
and \U$11703 ( \17851 , \8380 , \17802 );
and \U$11704 ( \17852 , \8382 , \17804 );
or \U$11714 ( \17853 , \17846 , \17847 , \17848 , \17849 , \17850 , \17851 , \17852 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5c93 ( \17854_nG5c93 , \17853 , \17817 );
buf \U$11715 ( \17855 , \17854_nG5c93 );
xor \U$11716 ( \17856 , \17845 , \17855 );
or \U$11717 ( \17857 , \17844 , \17856 );
buf \U$11718 ( \17858 , RIb7b94a0_249);
and \U$11719 ( \17859 , \7146 , \17788 );
and \U$11720 ( \17860 , \7148 , \17791 );
and \U$11721 ( \17861 , \8410 , \17794 );
and \U$11722 ( \17862 , \8412 , \17797 );
and \U$11723 ( \17863 , \8414 , \17799 );
and \U$11724 ( \17864 , \8416 , \17802 );
and \U$11725 ( \17865 , \8418 , \17804 );
or \U$11735 ( \17866 , \17859 , \17860 , \17861 , \17862 , \17863 , \17864 , \17865 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5ca0 ( \17867_nG5ca0 , \17866 , \17817 );
buf \U$11736 ( \17868 , \17867_nG5ca0 );
xor \U$11737 ( \17869 , \17858 , \17868 );
or \U$11738 ( \17870 , \17857 , \17869 );
buf \U$11739 ( \17871 , RIb7b9428_250);
and \U$11740 ( \17872 , \7156 , \17788 );
and \U$11741 ( \17873 , \7158 , \17791 );
and \U$11742 ( \17874 , \8446 , \17794 );
and \U$11743 ( \17875 , \8448 , \17797 );
and \U$11744 ( \17876 , \8450 , \17799 );
and \U$11745 ( \17877 , \8452 , \17802 );
and \U$11746 ( \17878 , \8454 , \17804 );
or \U$11756 ( \17879 , \17872 , \17873 , \17874 , \17875 , \17876 , \17877 , \17878 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5cad ( \17880_nG5cad , \17879 , \17817 );
buf \U$11757 ( \17881 , \17880_nG5cad );
xor \U$11758 ( \17882 , \17871 , \17881 );
or \U$11759 ( \17883 , \17870 , \17882 );
buf \U$11760 ( \17884 , RIb7b93b0_251);
and \U$11761 ( \17885 , \7166 , \17788 );
and \U$11762 ( \17886 , \7168 , \17791 );
and \U$11763 ( \17887 , \8482 , \17794 );
and \U$11764 ( \17888 , \8484 , \17797 );
and \U$11765 ( \17889 , \8486 , \17799 );
and \U$11766 ( \17890 , \8488 , \17802 );
and \U$11767 ( \17891 , \8490 , \17804 );
or \U$11777 ( \17892 , \17885 , \17886 , \17887 , \17888 , \17889 , \17890 , \17891 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5cba ( \17893_nG5cba , \17892 , \17817 );
buf \U$11778 ( \17894 , \17893_nG5cba );
xor \U$11779 ( \17895 , \17884 , \17894 );
or \U$11780 ( \17896 , \17883 , \17895 );
buf \U$11781 ( \17897 , RIb7af720_252);
and \U$11782 ( \17898 , \7176 , \17788 );
and \U$11783 ( \17899 , \7178 , \17791 );
and \U$11784 ( \17900 , \8518 , \17794 );
and \U$11785 ( \17901 , \8520 , \17797 );
and \U$11786 ( \17902 , \8522 , \17799 );
and \U$11787 ( \17903 , \8524 , \17802 );
and \U$11788 ( \17904 , \8526 , \17804 );
or \U$11798 ( \17905 , \17898 , \17899 , \17900 , \17901 , \17902 , \17903 , \17904 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5cc7 ( \17906_nG5cc7 , \17905 , \17817 );
buf \U$11799 ( \17907 , \17906_nG5cc7 );
xor \U$11800 ( \17908 , \17897 , \17907 );
or \U$11801 ( \17909 , \17896 , \17908 );
buf \U$11802 ( \17910 , RIb7af6a8_253);
and \U$11803 ( \17911 , \7186 , \17788 );
and \U$11804 ( \17912 , \7188 , \17791 );
and \U$11805 ( \17913 , \8554 , \17794 );
and \U$11806 ( \17914 , \8556 , \17797 );
and \U$11807 ( \17915 , \8558 , \17799 );
and \U$11808 ( \17916 , \8560 , \17802 );
and \U$11809 ( \17917 , \8562 , \17804 );
or \U$11819 ( \17918 , \17911 , \17912 , \17913 , \17914 , \17915 , \17916 , \17917 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5cd4 ( \17919_nG5cd4 , \17918 , \17817 );
buf \U$11820 ( \17920 , \17919_nG5cd4 );
xor \U$11821 ( \17921 , \17910 , \17920 );
or \U$11822 ( \17922 , \17909 , \17921 );
not \U$11823 ( \17923 , \17922 );
buf \U$11824 ( \17924 , \17923 );
buf \U$11825 ( \17925 , RIb7af630_254);
and \U$11826 ( \17926 , \7198 , \17788 );
and \U$11827 ( \17927 , \7200 , \17791 );
and \U$11828 ( \17928 , \8645 , \17794 );
and \U$11829 ( \17929 , \8673 , \17797 );
and \U$11830 ( \17930 , \8701 , \17799 );
and \U$11831 ( \17931 , \8729 , \17802 );
and \U$11832 ( \17932 , \8757 , \17804 );
or \U$11842 ( \17933 , \17926 , \17927 , \17928 , \17929 , \17930 , \17931 , \17932 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5ce3 ( \17934_nG5ce3 , \17933 , \17817 );
buf \U$11843 ( \17935 , \17934_nG5ce3 );
xor \U$11844 ( \17936 , \17925 , \17935 );
buf \U$11845 ( \17937 , RIb7af5b8_255);
and \U$11846 ( \17938 , \7207 , \17788 );
and \U$11847 ( \17939 , \7209 , \17791 );
and \U$11848 ( \17940 , \9119 , \17794 );
and \U$11849 ( \17941 , \9121 , \17797 );
and \U$11850 ( \17942 , \9123 , \17799 );
and \U$11851 ( \17943 , \9125 , \17802 );
and \U$11852 ( \17944 , \9127 , \17804 );
or \U$11862 ( \17945 , \17938 , \17939 , \17940 , \17941 , \17942 , \17943 , \17944 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5cef ( \17946_nG5cef , \17945 , \17817 );
buf \U$11863 ( \17947 , \17946_nG5cef );
xor \U$11864 ( \17948 , \17937 , \17947 );
or \U$11865 ( \17949 , \17936 , \17948 );
buf \U$11866 ( \17950 , RIb7af540_256);
and \U$11867 ( \17951 , \7217 , \17788 );
and \U$11868 ( \17952 , \7219 , \17791 );
and \U$11869 ( \17953 , \9155 , \17794 );
and \U$11870 ( \17954 , \9157 , \17797 );
and \U$11871 ( \17955 , \9159 , \17799 );
and \U$11872 ( \17956 , \9161 , \17802 );
and \U$11873 ( \17957 , \9163 , \17804 );
or \U$11883 ( \17958 , \17951 , \17952 , \17953 , \17954 , \17955 , \17956 , \17957 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5cfc ( \17959_nG5cfc , \17958 , \17817 );
buf \U$11884 ( \17960 , \17959_nG5cfc );
xor \U$11885 ( \17961 , \17950 , \17960 );
or \U$11886 ( \17962 , \17949 , \17961 );
buf \U$11887 ( \17963 , RIb7af4c8_257);
and \U$11888 ( \17964 , \7227 , \17788 );
and \U$11889 ( \17965 , \7229 , \17791 );
and \U$11890 ( \17966 , \9191 , \17794 );
and \U$11891 ( \17967 , \9193 , \17797 );
and \U$11892 ( \17968 , \9195 , \17799 );
and \U$11893 ( \17969 , \9197 , \17802 );
and \U$11894 ( \17970 , \9199 , \17804 );
or \U$11904 ( \17971 , \17964 , \17965 , \17966 , \17967 , \17968 , \17969 , \17970 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5d09 ( \17972_nG5d09 , \17971 , \17817 );
buf \U$11905 ( \17973 , \17972_nG5d09 );
xor \U$11906 ( \17974 , \17963 , \17973 );
or \U$11907 ( \17975 , \17962 , \17974 );
buf \U$11908 ( \17976 , RIb7af450_258);
and \U$11909 ( \17977 , \7237 , \17788 );
and \U$11910 ( \17978 , \7239 , \17791 );
and \U$11911 ( \17979 , \9227 , \17794 );
and \U$11912 ( \17980 , \9229 , \17797 );
and \U$11913 ( \17981 , \9231 , \17799 );
and \U$11914 ( \17982 , \9233 , \17802 );
and \U$11915 ( \17983 , \9235 , \17804 );
or \U$11925 ( \17984 , \17977 , \17978 , \17979 , \17980 , \17981 , \17982 , \17983 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5d16 ( \17985_nG5d16 , \17984 , \17817 );
buf \U$11926 ( \17986 , \17985_nG5d16 );
xor \U$11927 ( \17987 , \17976 , \17986 );
or \U$11928 ( \17988 , \17975 , \17987 );
buf \U$11929 ( \17989 , RIb7af3d8_259);
and \U$11930 ( \17990 , \7247 , \17788 );
and \U$11931 ( \17991 , \7249 , \17791 );
and \U$11932 ( \17992 , \9263 , \17794 );
and \U$11933 ( \17993 , \9265 , \17797 );
and \U$11934 ( \17994 , \9267 , \17799 );
and \U$11935 ( \17995 , \9269 , \17802 );
and \U$11936 ( \17996 , \9271 , \17804 );
or \U$11946 ( \17997 , \17990 , \17991 , \17992 , \17993 , \17994 , \17995 , \17996 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5d23 ( \17998_nG5d23 , \17997 , \17817 );
buf \U$11947 ( \17999 , \17998_nG5d23 );
xor \U$11948 ( \18000 , \17989 , \17999 );
or \U$11949 ( \18001 , \17988 , \18000 );
buf \U$11950 ( \18002 , RIb7a5bf8_260);
and \U$11951 ( \18003 , \7257 , \17788 );
and \U$11952 ( \18004 , \7259 , \17791 );
and \U$11953 ( \18005 , \9299 , \17794 );
and \U$11954 ( \18006 , \9301 , \17797 );
and \U$11955 ( \18007 , \9303 , \17799 );
and \U$11956 ( \18008 , \9305 , \17802 );
and \U$11957 ( \18009 , \9307 , \17804 );
or \U$11967 ( \18010 , \18003 , \18004 , \18005 , \18006 , \18007 , \18008 , \18009 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5d30 ( \18011_nG5d30 , \18010 , \17817 );
buf \U$11968 ( \18012 , \18011_nG5d30 );
xor \U$11969 ( \18013 , \18002 , \18012 );
or \U$11970 ( \18014 , \18001 , \18013 );
buf \U$11971 ( \18015 , RIb7a0c48_261);
and \U$11972 ( \18016 , \7267 , \17788 );
and \U$11973 ( \18017 , \7269 , \17791 );
and \U$11974 ( \18018 , \9335 , \17794 );
and \U$11975 ( \18019 , \9337 , \17797 );
and \U$11976 ( \18020 , \9339 , \17799 );
and \U$11977 ( \18021 , \9341 , \17802 );
and \U$11978 ( \18022 , \9343 , \17804 );
or \U$11988 ( \18023 , \18016 , \18017 , \18018 , \18019 , \18020 , \18021 , \18022 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g5d3d ( \18024_nG5d3d , \18023 , \17817 );
buf \U$11989 ( \18025 , \18024_nG5d3d );
xor \U$11990 ( \18026 , \18015 , \18025 );
or \U$11991 ( \18027 , \18014 , \18026 );
not \U$11992 ( \18028 , \18027 );
buf \U$11993 ( \18029 , \18028 );
and \U$11994 ( \18030 , \17924 , \18029 );
and \U$11995 ( \18031 , \17819 , \18030 );
_HMUX g5d45 ( \18032_nG5d45 , \17768_nG5c3c , \17770 , \18031 );
buf \U$11998 ( \18033 , \17770 );
buf \U$12001 ( \18034 , \17773 );
buf \U$12004 ( \18035 , \17776 );
buf \U$12007 ( \18036 , \17780 );
buf \U$12008 ( \18037 , \17784 );
not \U$12009 ( \18038 , \18037 );
buf \U$12010 ( \18039 , \18038 );
not \U$12011 ( \18040 , \18039 );
buf \U$12012 ( \18041 , \17787 );
xnor \U$12013 ( \18042 , \18041 , \18037 );
buf \U$12014 ( \18043 , \18042 );
or \U$12015 ( \18044 , \18041 , \18037 );
not \U$12016 ( \18045 , \18044 );
buf \U$12017 ( \18046 , \18045 );
buf \U$12018 ( \18047 , \18046 );
buf \U$12019 ( \18048 , \18046 );
buf \U$12020 ( \18049 , \18046 );
buf \U$12021 ( \18050 , \18046 );
buf \U$12022 ( \18051 , \18046 );
buf \U$12023 ( \18052 , \18046 );
buf \U$12024 ( \18053 , \18046 );
buf \U$12025 ( \18054 , \18046 );
buf \U$12026 ( \18055 , \18046 );
buf \U$12027 ( \18056 , \18046 );
buf \U$12028 ( \18057 , \18046 );
buf \U$12029 ( \18058 , \18046 );
buf \U$12030 ( \18059 , \18046 );
buf \U$12031 ( \18060 , \18046 );
buf \U$12032 ( \18061 , \18046 );
buf \U$12033 ( \18062 , \18046 );
buf \U$12034 ( \18063 , \18046 );
buf \U$12035 ( \18064 , \18046 );
buf \U$12036 ( \18065 , \18046 );
buf \U$12037 ( \18066 , \18046 );
buf \U$12038 ( \18067 , \18046 );
buf \U$12039 ( \18068 , \18046 );
buf \U$12040 ( \18069 , \18046 );
buf \U$12041 ( \18070 , \18046 );
buf \U$12042 ( \18071 , \18046 );
nor \U$12043 ( \18072 , \18033 , \18034 , \18035 , \18036 , \18040 , \18043 , \18046 , \18047 , \18048 , \18049 , \18050 , \18051 , \18052 , \18053 , \18054 , \18055 , \18056 , \18057 , \18058 , \18059 , \18060 , \18061 , \18062 , \18063 , \18064 , \18065 , \18066 , \18067 , \18068 , \18069 , \18070 , \18071 );
and \U$12044 ( \18073 , RIe5329d0_6883, \18072 );
not \U$12045 ( \18074 , \18033 );
not \U$12046 ( \18075 , \18034 );
not \U$12047 ( \18076 , \18035 );
not \U$12048 ( \18077 , \18036 );
buf \U$12049 ( \18078 , \18046 );
buf \U$12050 ( \18079 , \18046 );
buf \U$12051 ( \18080 , \18046 );
buf \U$12052 ( \18081 , \18046 );
buf \U$12053 ( \18082 , \18046 );
buf \U$12054 ( \18083 , \18046 );
buf \U$12055 ( \18084 , \18046 );
buf \U$12056 ( \18085 , \18046 );
buf \U$12057 ( \18086 , \18046 );
buf \U$12058 ( \18087 , \18046 );
buf \U$12059 ( \18088 , \18046 );
buf \U$12060 ( \18089 , \18046 );
buf \U$12061 ( \18090 , \18046 );
buf \U$12062 ( \18091 , \18046 );
buf \U$12063 ( \18092 , \18046 );
buf \U$12064 ( \18093 , \18046 );
buf \U$12065 ( \18094 , \18046 );
buf \U$12066 ( \18095 , \18046 );
buf \U$12067 ( \18096 , \18046 );
buf \U$12068 ( \18097 , \18046 );
buf \U$12069 ( \18098 , \18046 );
buf \U$12070 ( \18099 , \18046 );
buf \U$12071 ( \18100 , \18046 );
buf \U$12072 ( \18101 , \18046 );
buf \U$12073 ( \18102 , \18046 );
nor \U$12074 ( \18103 , \18074 , \18075 , \18076 , \18077 , \18039 , \18043 , \18046 , \18078 , \18079 , \18080 , \18081 , \18082 , \18083 , \18084 , \18085 , \18086 , \18087 , \18088 , \18089 , \18090 , \18091 , \18092 , \18093 , \18094 , \18095 , \18096 , \18097 , \18098 , \18099 , \18100 , \18101 , \18102 );
and \U$12075 ( \18104 , RIeb72150_6905, \18103 );
buf \U$12076 ( \18105 , \18046 );
buf \U$12077 ( \18106 , \18046 );
buf \U$12078 ( \18107 , \18046 );
buf \U$12079 ( \18108 , \18046 );
buf \U$12080 ( \18109 , \18046 );
buf \U$12081 ( \18110 , \18046 );
buf \U$12082 ( \18111 , \18046 );
buf \U$12083 ( \18112 , \18046 );
buf \U$12084 ( \18113 , \18046 );
buf \U$12085 ( \18114 , \18046 );
buf \U$12086 ( \18115 , \18046 );
buf \U$12087 ( \18116 , \18046 );
buf \U$12088 ( \18117 , \18046 );
buf \U$12089 ( \18118 , \18046 );
buf \U$12090 ( \18119 , \18046 );
buf \U$12091 ( \18120 , \18046 );
buf \U$12092 ( \18121 , \18046 );
buf \U$12093 ( \18122 , \18046 );
buf \U$12094 ( \18123 , \18046 );
buf \U$12095 ( \18124 , \18046 );
buf \U$12096 ( \18125 , \18046 );
buf \U$12097 ( \18126 , \18046 );
buf \U$12098 ( \18127 , \18046 );
buf \U$12099 ( \18128 , \18046 );
buf \U$12100 ( \18129 , \18046 );
nor \U$12101 ( \18130 , \18033 , \18075 , \18076 , \18077 , \18039 , \18043 , \18046 , \18105 , \18106 , \18107 , \18108 , \18109 , \18110 , \18111 , \18112 , \18113 , \18114 , \18115 , \18116 , \18117 , \18118 , \18119 , \18120 , \18121 , \18122 , \18123 , \18124 , \18125 , \18126 , \18127 , \18128 , \18129 );
and \U$12102 ( \18131 , RIeab80c0_6897, \18130 );
buf \U$12103 ( \18132 , \18046 );
buf \U$12104 ( \18133 , \18046 );
buf \U$12105 ( \18134 , \18046 );
buf \U$12106 ( \18135 , \18046 );
buf \U$12107 ( \18136 , \18046 );
buf \U$12108 ( \18137 , \18046 );
buf \U$12109 ( \18138 , \18046 );
buf \U$12110 ( \18139 , \18046 );
buf \U$12111 ( \18140 , \18046 );
buf \U$12112 ( \18141 , \18046 );
buf \U$12113 ( \18142 , \18046 );
buf \U$12114 ( \18143 , \18046 );
buf \U$12115 ( \18144 , \18046 );
buf \U$12116 ( \18145 , \18046 );
buf \U$12117 ( \18146 , \18046 );
buf \U$12118 ( \18147 , \18046 );
buf \U$12119 ( \18148 , \18046 );
buf \U$12120 ( \18149 , \18046 );
buf \U$12121 ( \18150 , \18046 );
buf \U$12122 ( \18151 , \18046 );
buf \U$12123 ( \18152 , \18046 );
buf \U$12124 ( \18153 , \18046 );
buf \U$12125 ( \18154 , \18046 );
buf \U$12126 ( \18155 , \18046 );
buf \U$12127 ( \18156 , \18046 );
nor \U$12128 ( \18157 , \18074 , \18034 , \18076 , \18077 , \18039 , \18043 , \18046 , \18132 , \18133 , \18134 , \18135 , \18136 , \18137 , \18138 , \18139 , \18140 , \18141 , \18142 , \18143 , \18144 , \18145 , \18146 , \18147 , \18148 , \18149 , \18150 , \18151 , \18152 , \18153 , \18154 , \18155 , \18156 );
and \U$12129 ( \18158 , RIe5331c8_6882, \18157 );
buf \U$12130 ( \18159 , \18046 );
buf \U$12131 ( \18160 , \18046 );
buf \U$12132 ( \18161 , \18046 );
buf \U$12133 ( \18162 , \18046 );
buf \U$12134 ( \18163 , \18046 );
buf \U$12135 ( \18164 , \18046 );
buf \U$12136 ( \18165 , \18046 );
buf \U$12137 ( \18166 , \18046 );
buf \U$12138 ( \18167 , \18046 );
buf \U$12139 ( \18168 , \18046 );
buf \U$12140 ( \18169 , \18046 );
buf \U$12141 ( \18170 , \18046 );
buf \U$12142 ( \18171 , \18046 );
buf \U$12143 ( \18172 , \18046 );
buf \U$12144 ( \18173 , \18046 );
buf \U$12145 ( \18174 , \18046 );
buf \U$12146 ( \18175 , \18046 );
buf \U$12147 ( \18176 , \18046 );
buf \U$12148 ( \18177 , \18046 );
buf \U$12149 ( \18178 , \18046 );
buf \U$12150 ( \18179 , \18046 );
buf \U$12151 ( \18180 , \18046 );
buf \U$12152 ( \18181 , \18046 );
buf \U$12153 ( \18182 , \18046 );
buf \U$12154 ( \18183 , \18046 );
nor \U$12155 ( \18184 , \18033 , \18034 , \18076 , \18077 , \18039 , \18043 , \18046 , \18159 , \18160 , \18161 , \18162 , \18163 , \18164 , \18165 , \18166 , \18167 , \18168 , \18169 , \18170 , \18171 , \18172 , \18173 , \18174 , \18175 , \18176 , \18177 , \18178 , \18179 , \18180 , \18181 , \18182 , \18183 );
and \U$12156 ( \18185 , RIe5339c0_6881, \18184 );
buf \U$12157 ( \18186 , \18046 );
buf \U$12158 ( \18187 , \18046 );
buf \U$12159 ( \18188 , \18046 );
buf \U$12160 ( \18189 , \18046 );
buf \U$12161 ( \18190 , \18046 );
buf \U$12162 ( \18191 , \18046 );
buf \U$12163 ( \18192 , \18046 );
buf \U$12164 ( \18193 , \18046 );
buf \U$12165 ( \18194 , \18046 );
buf \U$12166 ( \18195 , \18046 );
buf \U$12167 ( \18196 , \18046 );
buf \U$12168 ( \18197 , \18046 );
buf \U$12169 ( \18198 , \18046 );
buf \U$12170 ( \18199 , \18046 );
buf \U$12171 ( \18200 , \18046 );
buf \U$12172 ( \18201 , \18046 );
buf \U$12173 ( \18202 , \18046 );
buf \U$12174 ( \18203 , \18046 );
buf \U$12175 ( \18204 , \18046 );
buf \U$12176 ( \18205 , \18046 );
buf \U$12177 ( \18206 , \18046 );
buf \U$12178 ( \18207 , \18046 );
buf \U$12179 ( \18208 , \18046 );
buf \U$12180 ( \18209 , \18046 );
buf \U$12181 ( \18210 , \18046 );
nor \U$12182 ( \18211 , \18074 , \18075 , \18035 , \18077 , \18039 , \18043 , \18046 , \18186 , \18187 , \18188 , \18189 , \18190 , \18191 , \18192 , \18193 , \18194 , \18195 , \18196 , \18197 , \18198 , \18199 , \18200 , \18201 , \18202 , \18203 , \18204 , \18205 , \18206 , \18207 , \18208 , \18209 , \18210 );
and \U$12183 ( \18212 , RIeab87c8_6898, \18211 );
buf \U$12184 ( \18213 , \18046 );
buf \U$12185 ( \18214 , \18046 );
buf \U$12186 ( \18215 , \18046 );
buf \U$12187 ( \18216 , \18046 );
buf \U$12188 ( \18217 , \18046 );
buf \U$12189 ( \18218 , \18046 );
buf \U$12190 ( \18219 , \18046 );
buf \U$12191 ( \18220 , \18046 );
buf \U$12192 ( \18221 , \18046 );
buf \U$12193 ( \18222 , \18046 );
buf \U$12194 ( \18223 , \18046 );
buf \U$12195 ( \18224 , \18046 );
buf \U$12196 ( \18225 , \18046 );
buf \U$12197 ( \18226 , \18046 );
buf \U$12198 ( \18227 , \18046 );
buf \U$12199 ( \18228 , \18046 );
buf \U$12200 ( \18229 , \18046 );
buf \U$12201 ( \18230 , \18046 );
buf \U$12202 ( \18231 , \18046 );
buf \U$12203 ( \18232 , \18046 );
buf \U$12204 ( \18233 , \18046 );
buf \U$12205 ( \18234 , \18046 );
buf \U$12206 ( \18235 , \18046 );
buf \U$12207 ( \18236 , \18046 );
buf \U$12208 ( \18237 , \18046 );
nor \U$12209 ( \18238 , \18033 , \18075 , \18035 , \18077 , \18039 , \18043 , \18046 , \18213 , \18214 , \18215 , \18216 , \18217 , \18218 , \18219 , \18220 , \18221 , \18222 , \18223 , \18224 , \18225 , \18226 , \18227 , \18228 , \18229 , \18230 , \18231 , \18232 , \18233 , \18234 , \18235 , \18236 , \18237 );
and \U$12210 ( \18239 , RIe5341b8_6880, \18238 );
buf \U$12211 ( \18240 , \18046 );
buf \U$12212 ( \18241 , \18046 );
buf \U$12213 ( \18242 , \18046 );
buf \U$12214 ( \18243 , \18046 );
buf \U$12215 ( \18244 , \18046 );
buf \U$12216 ( \18245 , \18046 );
buf \U$12217 ( \18246 , \18046 );
buf \U$12218 ( \18247 , \18046 );
buf \U$12219 ( \18248 , \18046 );
buf \U$12220 ( \18249 , \18046 );
buf \U$12221 ( \18250 , \18046 );
buf \U$12222 ( \18251 , \18046 );
buf \U$12223 ( \18252 , \18046 );
buf \U$12224 ( \18253 , \18046 );
buf \U$12225 ( \18254 , \18046 );
buf \U$12226 ( \18255 , \18046 );
buf \U$12227 ( \18256 , \18046 );
buf \U$12228 ( \18257 , \18046 );
buf \U$12229 ( \18258 , \18046 );
buf \U$12230 ( \18259 , \18046 );
buf \U$12231 ( \18260 , \18046 );
buf \U$12232 ( \18261 , \18046 );
buf \U$12233 ( \18262 , \18046 );
buf \U$12234 ( \18263 , \18046 );
buf \U$12235 ( \18264 , \18046 );
nor \U$12236 ( \18265 , \18074 , \18034 , \18035 , \18077 , \18039 , \18043 , \18046 , \18240 , \18241 , \18242 , \18243 , \18244 , \18245 , \18246 , \18247 , \18248 , \18249 , \18250 , \18251 , \18252 , \18253 , \18254 , \18255 , \18256 , \18257 , \18258 , \18259 , \18260 , \18261 , \18262 , \18263 , \18264 );
and \U$12237 ( \18266 , RIe5349b0_6879, \18265 );
buf \U$12238 ( \18267 , \18046 );
buf \U$12239 ( \18268 , \18046 );
buf \U$12240 ( \18269 , \18046 );
buf \U$12241 ( \18270 , \18046 );
buf \U$12242 ( \18271 , \18046 );
buf \U$12243 ( \18272 , \18046 );
buf \U$12244 ( \18273 , \18046 );
buf \U$12245 ( \18274 , \18046 );
buf \U$12246 ( \18275 , \18046 );
buf \U$12247 ( \18276 , \18046 );
buf \U$12248 ( \18277 , \18046 );
buf \U$12249 ( \18278 , \18046 );
buf \U$12250 ( \18279 , \18046 );
buf \U$12251 ( \18280 , \18046 );
buf \U$12252 ( \18281 , \18046 );
buf \U$12253 ( \18282 , \18046 );
buf \U$12254 ( \18283 , \18046 );
buf \U$12255 ( \18284 , \18046 );
buf \U$12256 ( \18285 , \18046 );
buf \U$12257 ( \18286 , \18046 );
buf \U$12258 ( \18287 , \18046 );
buf \U$12259 ( \18288 , \18046 );
buf \U$12260 ( \18289 , \18046 );
buf \U$12261 ( \18290 , \18046 );
buf \U$12262 ( \18291 , \18046 );
nor \U$12263 ( \18292 , \18033 , \18034 , \18035 , \18077 , \18039 , \18043 , \18046 , \18267 , \18268 , \18269 , \18270 , \18271 , \18272 , \18273 , \18274 , \18275 , \18276 , \18277 , \18278 , \18279 , \18280 , \18281 , \18282 , \18283 , \18284 , \18285 , \18286 , \18287 , \18288 , \18289 , \18290 , \18291 );
and \U$12264 ( \18293 , RIea94af8_6890, \18292 );
buf \U$12265 ( \18294 , \18046 );
buf \U$12266 ( \18295 , \18046 );
buf \U$12267 ( \18296 , \18046 );
buf \U$12268 ( \18297 , \18046 );
buf \U$12269 ( \18298 , \18046 );
buf \U$12270 ( \18299 , \18046 );
buf \U$12271 ( \18300 , \18046 );
buf \U$12272 ( \18301 , \18046 );
buf \U$12273 ( \18302 , \18046 );
buf \U$12274 ( \18303 , \18046 );
buf \U$12275 ( \18304 , \18046 );
buf \U$12276 ( \18305 , \18046 );
buf \U$12277 ( \18306 , \18046 );
buf \U$12278 ( \18307 , \18046 );
buf \U$12279 ( \18308 , \18046 );
buf \U$12280 ( \18309 , \18046 );
buf \U$12281 ( \18310 , \18046 );
buf \U$12282 ( \18311 , \18046 );
buf \U$12283 ( \18312 , \18046 );
buf \U$12284 ( \18313 , \18046 );
buf \U$12285 ( \18314 , \18046 );
buf \U$12286 ( \18315 , \18046 );
buf \U$12287 ( \18316 , \18046 );
buf \U$12288 ( \18317 , \18046 );
buf \U$12289 ( \18318 , \18046 );
nor \U$12290 ( \18319 , \18074 , \18075 , \18076 , \18036 , \18039 , \18043 , \18046 , \18294 , \18295 , \18296 , \18297 , \18298 , \18299 , \18300 , \18301 , \18302 , \18303 , \18304 , \18305 , \18306 , \18307 , \18308 , \18309 , \18310 , \18311 , \18312 , \18313 , \18314 , \18315 , \18316 , \18317 , \18318 );
and \U$12291 ( \18320 , RIe5351a8_6878, \18319 );
buf \U$12292 ( \18321 , \18046 );
buf \U$12293 ( \18322 , \18046 );
buf \U$12294 ( \18323 , \18046 );
buf \U$12295 ( \18324 , \18046 );
buf \U$12296 ( \18325 , \18046 );
buf \U$12297 ( \18326 , \18046 );
buf \U$12298 ( \18327 , \18046 );
buf \U$12299 ( \18328 , \18046 );
buf \U$12300 ( \18329 , \18046 );
buf \U$12301 ( \18330 , \18046 );
buf \U$12302 ( \18331 , \18046 );
buf \U$12303 ( \18332 , \18046 );
buf \U$12304 ( \18333 , \18046 );
buf \U$12305 ( \18334 , \18046 );
buf \U$12306 ( \18335 , \18046 );
buf \U$12307 ( \18336 , \18046 );
buf \U$12308 ( \18337 , \18046 );
buf \U$12309 ( \18338 , \18046 );
buf \U$12310 ( \18339 , \18046 );
buf \U$12311 ( \18340 , \18046 );
buf \U$12312 ( \18341 , \18046 );
buf \U$12313 ( \18342 , \18046 );
buf \U$12314 ( \18343 , \18046 );
buf \U$12315 ( \18344 , \18046 );
buf \U$12316 ( \18345 , \18046 );
nor \U$12317 ( \18346 , \18033 , \18075 , \18076 , \18036 , \18039 , \18043 , \18046 , \18321 , \18322 , \18323 , \18324 , \18325 , \18326 , \18327 , \18328 , \18329 , \18330 , \18331 , \18332 , \18333 , \18334 , \18335 , \18336 , \18337 , \18338 , \18339 , \18340 , \18341 , \18342 , \18343 , \18344 , \18345 );
and \U$12318 ( \18347 , RIe5359a0_6877, \18346 );
buf \U$12319 ( \18348 , \18046 );
buf \U$12320 ( \18349 , \18046 );
buf \U$12321 ( \18350 , \18046 );
buf \U$12322 ( \18351 , \18046 );
buf \U$12323 ( \18352 , \18046 );
buf \U$12324 ( \18353 , \18046 );
buf \U$12325 ( \18354 , \18046 );
buf \U$12326 ( \18355 , \18046 );
buf \U$12327 ( \18356 , \18046 );
buf \U$12328 ( \18357 , \18046 );
buf \U$12329 ( \18358 , \18046 );
buf \U$12330 ( \18359 , \18046 );
buf \U$12331 ( \18360 , \18046 );
buf \U$12332 ( \18361 , \18046 );
buf \U$12333 ( \18362 , \18046 );
buf \U$12334 ( \18363 , \18046 );
buf \U$12335 ( \18364 , \18046 );
buf \U$12336 ( \18365 , \18046 );
buf \U$12337 ( \18366 , \18046 );
buf \U$12338 ( \18367 , \18046 );
buf \U$12339 ( \18368 , \18046 );
buf \U$12340 ( \18369 , \18046 );
buf \U$12341 ( \18370 , \18046 );
buf \U$12342 ( \18371 , \18046 );
buf \U$12343 ( \18372 , \18046 );
nor \U$12344 ( \18373 , \18074 , \18034 , \18076 , \18036 , \18039 , \18043 , \18046 , \18348 , \18349 , \18350 , \18351 , \18352 , \18353 , \18354 , \18355 , \18356 , \18357 , \18358 , \18359 , \18360 , \18361 , \18362 , \18363 , \18364 , \18365 , \18366 , \18367 , \18368 , \18369 , \18370 , \18371 , \18372 );
and \U$12345 ( \18374 , RIeab78c8_6895, \18373 );
buf \U$12346 ( \18375 , \18046 );
buf \U$12347 ( \18376 , \18046 );
buf \U$12348 ( \18377 , \18046 );
buf \U$12349 ( \18378 , \18046 );
buf \U$12350 ( \18379 , \18046 );
buf \U$12351 ( \18380 , \18046 );
buf \U$12352 ( \18381 , \18046 );
buf \U$12353 ( \18382 , \18046 );
buf \U$12354 ( \18383 , \18046 );
buf \U$12355 ( \18384 , \18046 );
buf \U$12356 ( \18385 , \18046 );
buf \U$12357 ( \18386 , \18046 );
buf \U$12358 ( \18387 , \18046 );
buf \U$12359 ( \18388 , \18046 );
buf \U$12360 ( \18389 , \18046 );
buf \U$12361 ( \18390 , \18046 );
buf \U$12362 ( \18391 , \18046 );
buf \U$12363 ( \18392 , \18046 );
buf \U$12364 ( \18393 , \18046 );
buf \U$12365 ( \18394 , \18046 );
buf \U$12366 ( \18395 , \18046 );
buf \U$12367 ( \18396 , \18046 );
buf \U$12368 ( \18397 , \18046 );
buf \U$12369 ( \18398 , \18046 );
buf \U$12370 ( \18399 , \18046 );
nor \U$12371 ( \18400 , \18033 , \18034 , \18076 , \18036 , \18039 , \18043 , \18046 , \18375 , \18376 , \18377 , \18378 , \18379 , \18380 , \18381 , \18382 , \18383 , \18384 , \18385 , \18386 , \18387 , \18388 , \18389 , \18390 , \18391 , \18392 , \18393 , \18394 , \18395 , \18396 , \18397 , \18398 , \18399 );
and \U$12372 ( \18401 , RIeab7d00_6896, \18400 );
buf \U$12373 ( \18402 , \18046 );
buf \U$12374 ( \18403 , \18046 );
buf \U$12375 ( \18404 , \18046 );
buf \U$12376 ( \18405 , \18046 );
buf \U$12377 ( \18406 , \18046 );
buf \U$12378 ( \18407 , \18046 );
buf \U$12379 ( \18408 , \18046 );
buf \U$12380 ( \18409 , \18046 );
buf \U$12381 ( \18410 , \18046 );
buf \U$12382 ( \18411 , \18046 );
buf \U$12383 ( \18412 , \18046 );
buf \U$12384 ( \18413 , \18046 );
buf \U$12385 ( \18414 , \18046 );
buf \U$12386 ( \18415 , \18046 );
buf \U$12387 ( \18416 , \18046 );
buf \U$12388 ( \18417 , \18046 );
buf \U$12389 ( \18418 , \18046 );
buf \U$12390 ( \18419 , \18046 );
buf \U$12391 ( \18420 , \18046 );
buf \U$12392 ( \18421 , \18046 );
buf \U$12393 ( \18422 , \18046 );
buf \U$12394 ( \18423 , \18046 );
buf \U$12395 ( \18424 , \18046 );
buf \U$12396 ( \18425 , \18046 );
buf \U$12397 ( \18426 , \18046 );
nor \U$12398 ( \18427 , \18074 , \18075 , \18035 , \18036 , \18039 , \18043 , \18046 , \18402 , \18403 , \18404 , \18405 , \18406 , \18407 , \18408 , \18409 , \18410 , \18411 , \18412 , \18413 , \18414 , \18415 , \18416 , \18417 , \18418 , \18419 , \18420 , \18421 , \18422 , \18423 , \18424 , \18425 , \18426 );
and \U$12399 ( \18428 , RIeacfa18_6902, \18427 );
buf \U$12400 ( \18429 , \18046 );
buf \U$12401 ( \18430 , \18046 );
buf \U$12402 ( \18431 , \18046 );
buf \U$12403 ( \18432 , \18046 );
buf \U$12404 ( \18433 , \18046 );
buf \U$12405 ( \18434 , \18046 );
buf \U$12406 ( \18435 , \18046 );
buf \U$12407 ( \18436 , \18046 );
buf \U$12408 ( \18437 , \18046 );
buf \U$12409 ( \18438 , \18046 );
buf \U$12410 ( \18439 , \18046 );
buf \U$12411 ( \18440 , \18046 );
buf \U$12412 ( \18441 , \18046 );
buf \U$12413 ( \18442 , \18046 );
buf \U$12414 ( \18443 , \18046 );
buf \U$12415 ( \18444 , \18046 );
buf \U$12416 ( \18445 , \18046 );
buf \U$12417 ( \18446 , \18046 );
buf \U$12418 ( \18447 , \18046 );
buf \U$12419 ( \18448 , \18046 );
buf \U$12420 ( \18449 , \18046 );
buf \U$12421 ( \18450 , \18046 );
buf \U$12422 ( \18451 , \18046 );
buf \U$12423 ( \18452 , \18046 );
buf \U$12424 ( \18453 , \18046 );
nor \U$12425 ( \18454 , \18033 , \18075 , \18035 , \18036 , \18039 , \18043 , \18046 , \18429 , \18430 , \18431 , \18432 , \18433 , \18434 , \18435 , \18436 , \18437 , \18438 , \18439 , \18440 , \18441 , \18442 , \18443 , \18444 , \18445 , \18446 , \18447 , \18448 , \18449 , \18450 , \18451 , \18452 , \18453 );
and \U$12426 ( \18455 , RIeab6518_6891, \18454 );
buf \U$12427 ( \18456 , \18046 );
buf \U$12428 ( \18457 , \18046 );
buf \U$12429 ( \18458 , \18046 );
buf \U$12430 ( \18459 , \18046 );
buf \U$12431 ( \18460 , \18046 );
buf \U$12432 ( \18461 , \18046 );
buf \U$12433 ( \18462 , \18046 );
buf \U$12434 ( \18463 , \18046 );
buf \U$12435 ( \18464 , \18046 );
buf \U$12436 ( \18465 , \18046 );
buf \U$12437 ( \18466 , \18046 );
buf \U$12438 ( \18467 , \18046 );
buf \U$12439 ( \18468 , \18046 );
buf \U$12440 ( \18469 , \18046 );
buf \U$12441 ( \18470 , \18046 );
buf \U$12442 ( \18471 , \18046 );
buf \U$12443 ( \18472 , \18046 );
buf \U$12444 ( \18473 , \18046 );
buf \U$12445 ( \18474 , \18046 );
buf \U$12446 ( \18475 , \18046 );
buf \U$12447 ( \18476 , \18046 );
buf \U$12448 ( \18477 , \18046 );
buf \U$12449 ( \18478 , \18046 );
buf \U$12450 ( \18479 , \18046 );
buf \U$12451 ( \18480 , \18046 );
nor \U$12452 ( \18481 , \18074 , \18034 , \18035 , \18036 , \18039 , \18043 , \18046 , \18456 , \18457 , \18458 , \18459 , \18460 , \18461 , \18462 , \18463 , \18464 , \18465 , \18466 , \18467 , \18468 , \18469 , \18470 , \18471 , \18472 , \18473 , \18474 , \18475 , \18476 , \18477 , \18478 , \18479 , \18480 );
and \U$12453 ( \18482 , RIeb352c8_6904, \18481 );
or \U$12454 ( \18483 , \18073 , \18104 , \18131 , \18158 , \18185 , \18212 , \18239 , \18266 , \18293 , \18320 , \18347 , \18374 , \18401 , \18428 , \18455 , \18482 );
buf \U$12455 ( \18484 , \18046 );
not \U$12456 ( \18485 , \18484 );
buf \U$12457 ( \18486 , \18034 );
buf \U$12458 ( \18487 , \18035 );
buf \U$12459 ( \18488 , \18036 );
buf \U$12460 ( \18489 , \18039 );
buf \U$12461 ( \18490 , \18043 );
buf \U$12462 ( \18491 , \18046 );
buf \U$12463 ( \18492 , \18046 );
buf \U$12464 ( \18493 , \18046 );
buf \U$12465 ( \18494 , \18046 );
buf \U$12466 ( \18495 , \18046 );
buf \U$12467 ( \18496 , \18046 );
buf \U$12468 ( \18497 , \18046 );
buf \U$12469 ( \18498 , \18046 );
buf \U$12470 ( \18499 , \18046 );
buf \U$12471 ( \18500 , \18046 );
buf \U$12472 ( \18501 , \18046 );
buf \U$12473 ( \18502 , \18046 );
buf \U$12474 ( \18503 , \18046 );
buf \U$12475 ( \18504 , \18046 );
buf \U$12476 ( \18505 , \18046 );
buf \U$12477 ( \18506 , \18046 );
buf \U$12478 ( \18507 , \18046 );
buf \U$12479 ( \18508 , \18046 );
buf \U$12480 ( \18509 , \18046 );
buf \U$12481 ( \18510 , \18046 );
buf \U$12482 ( \18511 , \18046 );
buf \U$12483 ( \18512 , \18046 );
buf \U$12484 ( \18513 , \18046 );
buf \U$12485 ( \18514 , \18046 );
buf \U$12486 ( \18515 , \18046 );
buf \U$12487 ( \18516 , \18033 );
or \U$12488 ( \18517 , \18486 , \18487 , \18488 , \18489 , \18490 , \18491 , \18492 , \18493 , \18494 , \18495 , \18496 , \18497 , \18498 , \18499 , \18500 , \18501 , \18502 , \18503 , \18504 , \18505 , \18506 , \18507 , \18508 , \18509 , \18510 , \18511 , \18512 , \18513 , \18514 , \18515 , \18516 );
nand \U$12489 ( \18518 , \18485 , \18517 );
buf \U$12490 ( \18519 , \18518 );
buf \U$12491 ( \18520 , \18046 );
not \U$12492 ( \18521 , \18520 );
buf \U$12493 ( \18522 , \18043 );
buf \U$12494 ( \18523 , \18046 );
buf \U$12495 ( \18524 , \18046 );
buf \U$12496 ( \18525 , \18046 );
buf \U$12497 ( \18526 , \18046 );
buf \U$12498 ( \18527 , \18046 );
buf \U$12499 ( \18528 , \18046 );
buf \U$12500 ( \18529 , \18046 );
buf \U$12501 ( \18530 , \18046 );
buf \U$12502 ( \18531 , \18046 );
buf \U$12503 ( \18532 , \18046 );
buf \U$12504 ( \18533 , \18046 );
buf \U$12505 ( \18534 , \18046 );
buf \U$12506 ( \18535 , \18046 );
buf \U$12507 ( \18536 , \18046 );
buf \U$12508 ( \18537 , \18046 );
buf \U$12509 ( \18538 , \18046 );
buf \U$12510 ( \18539 , \18046 );
buf \U$12511 ( \18540 , \18046 );
buf \U$12512 ( \18541 , \18046 );
buf \U$12513 ( \18542 , \18046 );
buf \U$12514 ( \18543 , \18046 );
buf \U$12515 ( \18544 , \18046 );
buf \U$12516 ( \18545 , \18046 );
buf \U$12517 ( \18546 , \18046 );
buf \U$12518 ( \18547 , \18046 );
buf \U$12519 ( \18548 , \18039 );
buf \U$12520 ( \18549 , \18033 );
buf \U$12521 ( \18550 , \18034 );
buf \U$12522 ( \18551 , \18035 );
buf \U$12523 ( \18552 , \18036 );
or \U$12524 ( \18553 , \18549 , \18550 , \18551 , \18552 );
and \U$12525 ( \18554 , \18548 , \18553 );
or \U$12526 ( \18555 , \18522 , \18523 , \18524 , \18525 , \18526 , \18527 , \18528 , \18529 , \18530 , \18531 , \18532 , \18533 , \18534 , \18535 , \18536 , \18537 , \18538 , \18539 , \18540 , \18541 , \18542 , \18543 , \18544 , \18545 , \18546 , \18547 , \18554 );
and \U$12527 ( \18556 , \18521 , \18555 );
buf \U$12528 ( \18557 , \18556 );
or \U$12529 ( \18558 , \18519 , \18557 );
_DC g5f5c ( \18559_nG5f5c , \18483 , \18558 );
not \U$12530 ( \18560 , \18559_nG5f5c );
buf \U$12531 ( \18561 , RIb7b9608_246);
buf \U$12532 ( \18562 , \18046 );
buf \U$12533 ( \18563 , \18046 );
buf \U$12534 ( \18564 , \18046 );
buf \U$12535 ( \18565 , \18046 );
buf \U$12536 ( \18566 , \18046 );
buf \U$12537 ( \18567 , \18046 );
buf \U$12538 ( \18568 , \18046 );
buf \U$12539 ( \18569 , \18046 );
buf \U$12540 ( \18570 , \18046 );
buf \U$12541 ( \18571 , \18046 );
buf \U$12542 ( \18572 , \18046 );
buf \U$12543 ( \18573 , \18046 );
buf \U$12544 ( \18574 , \18046 );
buf \U$12545 ( \18575 , \18046 );
buf \U$12546 ( \18576 , \18046 );
buf \U$12547 ( \18577 , \18046 );
buf \U$12548 ( \18578 , \18046 );
buf \U$12549 ( \18579 , \18046 );
buf \U$12550 ( \18580 , \18046 );
buf \U$12551 ( \18581 , \18046 );
buf \U$12552 ( \18582 , \18046 );
buf \U$12553 ( \18583 , \18046 );
buf \U$12554 ( \18584 , \18046 );
buf \U$12555 ( \18585 , \18046 );
buf \U$12556 ( \18586 , \18046 );
nor \U$12557 ( \18587 , \18033 , \18034 , \18035 , \18036 , \18040 , \18043 , \18046 , \18562 , \18563 , \18564 , \18565 , \18566 , \18567 , \18568 , \18569 , \18570 , \18571 , \18572 , \18573 , \18574 , \18575 , \18576 , \18577 , \18578 , \18579 , \18580 , \18581 , \18582 , \18583 , \18584 , \18585 , \18586 );
and \U$12558 ( \18588 , \7117 , \18587 );
buf \U$12559 ( \18589 , \18046 );
buf \U$12560 ( \18590 , \18046 );
buf \U$12561 ( \18591 , \18046 );
buf \U$12562 ( \18592 , \18046 );
buf \U$12563 ( \18593 , \18046 );
buf \U$12564 ( \18594 , \18046 );
buf \U$12565 ( \18595 , \18046 );
buf \U$12566 ( \18596 , \18046 );
buf \U$12567 ( \18597 , \18046 );
buf \U$12568 ( \18598 , \18046 );
buf \U$12569 ( \18599 , \18046 );
buf \U$12570 ( \18600 , \18046 );
buf \U$12571 ( \18601 , \18046 );
buf \U$12572 ( \18602 , \18046 );
buf \U$12573 ( \18603 , \18046 );
buf \U$12574 ( \18604 , \18046 );
buf \U$12575 ( \18605 , \18046 );
buf \U$12576 ( \18606 , \18046 );
buf \U$12577 ( \18607 , \18046 );
buf \U$12578 ( \18608 , \18046 );
buf \U$12579 ( \18609 , \18046 );
buf \U$12580 ( \18610 , \18046 );
buf \U$12581 ( \18611 , \18046 );
buf \U$12582 ( \18612 , \18046 );
buf \U$12583 ( \18613 , \18046 );
nor \U$12584 ( \18614 , \18074 , \18075 , \18076 , \18077 , \18039 , \18043 , \18046 , \18589 , \18590 , \18591 , \18592 , \18593 , \18594 , \18595 , \18596 , \18597 , \18598 , \18599 , \18600 , \18601 , \18602 , \18603 , \18604 , \18605 , \18606 , \18607 , \18608 , \18609 , \18610 , \18611 , \18612 , \18613 );
and \U$12585 ( \18615 , \7119 , \18614 );
buf \U$12586 ( \18616 , \18046 );
buf \U$12587 ( \18617 , \18046 );
buf \U$12588 ( \18618 , \18046 );
buf \U$12589 ( \18619 , \18046 );
buf \U$12590 ( \18620 , \18046 );
buf \U$12591 ( \18621 , \18046 );
buf \U$12592 ( \18622 , \18046 );
buf \U$12593 ( \18623 , \18046 );
buf \U$12594 ( \18624 , \18046 );
buf \U$12595 ( \18625 , \18046 );
buf \U$12596 ( \18626 , \18046 );
buf \U$12597 ( \18627 , \18046 );
buf \U$12598 ( \18628 , \18046 );
buf \U$12599 ( \18629 , \18046 );
buf \U$12600 ( \18630 , \18046 );
buf \U$12601 ( \18631 , \18046 );
buf \U$12602 ( \18632 , \18046 );
buf \U$12603 ( \18633 , \18046 );
buf \U$12604 ( \18634 , \18046 );
buf \U$12605 ( \18635 , \18046 );
buf \U$12606 ( \18636 , \18046 );
buf \U$12607 ( \18637 , \18046 );
buf \U$12608 ( \18638 , \18046 );
buf \U$12609 ( \18639 , \18046 );
buf \U$12610 ( \18640 , \18046 );
nor \U$12611 ( \18641 , \18033 , \18075 , \18076 , \18077 , \18039 , \18043 , \18046 , \18616 , \18617 , \18618 , \18619 , \18620 , \18621 , \18622 , \18623 , \18624 , \18625 , \18626 , \18627 , \18628 , \18629 , \18630 , \18631 , \18632 , \18633 , \18634 , \18635 , \18636 , \18637 , \18638 , \18639 , \18640 );
and \U$12612 ( \18642 , \7864 , \18641 );
buf \U$12613 ( \18643 , \18046 );
buf \U$12614 ( \18644 , \18046 );
buf \U$12615 ( \18645 , \18046 );
buf \U$12616 ( \18646 , \18046 );
buf \U$12617 ( \18647 , \18046 );
buf \U$12618 ( \18648 , \18046 );
buf \U$12619 ( \18649 , \18046 );
buf \U$12620 ( \18650 , \18046 );
buf \U$12621 ( \18651 , \18046 );
buf \U$12622 ( \18652 , \18046 );
buf \U$12623 ( \18653 , \18046 );
buf \U$12624 ( \18654 , \18046 );
buf \U$12625 ( \18655 , \18046 );
buf \U$12626 ( \18656 , \18046 );
buf \U$12627 ( \18657 , \18046 );
buf \U$12628 ( \18658 , \18046 );
buf \U$12629 ( \18659 , \18046 );
buf \U$12630 ( \18660 , \18046 );
buf \U$12631 ( \18661 , \18046 );
buf \U$12632 ( \18662 , \18046 );
buf \U$12633 ( \18663 , \18046 );
buf \U$12634 ( \18664 , \18046 );
buf \U$12635 ( \18665 , \18046 );
buf \U$12636 ( \18666 , \18046 );
buf \U$12637 ( \18667 , \18046 );
nor \U$12638 ( \18668 , \18074 , \18034 , \18076 , \18077 , \18039 , \18043 , \18046 , \18643 , \18644 , \18645 , \18646 , \18647 , \18648 , \18649 , \18650 , \18651 , \18652 , \18653 , \18654 , \18655 , \18656 , \18657 , \18658 , \18659 , \18660 , \18661 , \18662 , \18663 , \18664 , \18665 , \18666 , \18667 );
and \U$12639 ( \18669 , \7892 , \18668 );
buf \U$12640 ( \18670 , \18046 );
buf \U$12641 ( \18671 , \18046 );
buf \U$12642 ( \18672 , \18046 );
buf \U$12643 ( \18673 , \18046 );
buf \U$12644 ( \18674 , \18046 );
buf \U$12645 ( \18675 , \18046 );
buf \U$12646 ( \18676 , \18046 );
buf \U$12647 ( \18677 , \18046 );
buf \U$12648 ( \18678 , \18046 );
buf \U$12649 ( \18679 , \18046 );
buf \U$12650 ( \18680 , \18046 );
buf \U$12651 ( \18681 , \18046 );
buf \U$12652 ( \18682 , \18046 );
buf \U$12653 ( \18683 , \18046 );
buf \U$12654 ( \18684 , \18046 );
buf \U$12655 ( \18685 , \18046 );
buf \U$12656 ( \18686 , \18046 );
buf \U$12657 ( \18687 , \18046 );
buf \U$12658 ( \18688 , \18046 );
buf \U$12659 ( \18689 , \18046 );
buf \U$12660 ( \18690 , \18046 );
buf \U$12661 ( \18691 , \18046 );
buf \U$12662 ( \18692 , \18046 );
buf \U$12663 ( \18693 , \18046 );
buf \U$12664 ( \18694 , \18046 );
nor \U$12665 ( \18695 , \18033 , \18034 , \18076 , \18077 , \18039 , \18043 , \18046 , \18670 , \18671 , \18672 , \18673 , \18674 , \18675 , \18676 , \18677 , \18678 , \18679 , \18680 , \18681 , \18682 , \18683 , \18684 , \18685 , \18686 , \18687 , \18688 , \18689 , \18690 , \18691 , \18692 , \18693 , \18694 );
and \U$12666 ( \18696 , \7920 , \18695 );
buf \U$12667 ( \18697 , \18046 );
buf \U$12668 ( \18698 , \18046 );
buf \U$12669 ( \18699 , \18046 );
buf \U$12670 ( \18700 , \18046 );
buf \U$12671 ( \18701 , \18046 );
buf \U$12672 ( \18702 , \18046 );
buf \U$12673 ( \18703 , \18046 );
buf \U$12674 ( \18704 , \18046 );
buf \U$12675 ( \18705 , \18046 );
buf \U$12676 ( \18706 , \18046 );
buf \U$12677 ( \18707 , \18046 );
buf \U$12678 ( \18708 , \18046 );
buf \U$12679 ( \18709 , \18046 );
buf \U$12680 ( \18710 , \18046 );
buf \U$12681 ( \18711 , \18046 );
buf \U$12682 ( \18712 , \18046 );
buf \U$12683 ( \18713 , \18046 );
buf \U$12684 ( \18714 , \18046 );
buf \U$12685 ( \18715 , \18046 );
buf \U$12686 ( \18716 , \18046 );
buf \U$12687 ( \18717 , \18046 );
buf \U$12688 ( \18718 , \18046 );
buf \U$12689 ( \18719 , \18046 );
buf \U$12690 ( \18720 , \18046 );
buf \U$12691 ( \18721 , \18046 );
nor \U$12692 ( \18722 , \18074 , \18075 , \18035 , \18077 , \18039 , \18043 , \18046 , \18697 , \18698 , \18699 , \18700 , \18701 , \18702 , \18703 , \18704 , \18705 , \18706 , \18707 , \18708 , \18709 , \18710 , \18711 , \18712 , \18713 , \18714 , \18715 , \18716 , \18717 , \18718 , \18719 , \18720 , \18721 );
and \U$12693 ( \18723 , \7948 , \18722 );
buf \U$12694 ( \18724 , \18046 );
buf \U$12695 ( \18725 , \18046 );
buf \U$12696 ( \18726 , \18046 );
buf \U$12697 ( \18727 , \18046 );
buf \U$12698 ( \18728 , \18046 );
buf \U$12699 ( \18729 , \18046 );
buf \U$12700 ( \18730 , \18046 );
buf \U$12701 ( \18731 , \18046 );
buf \U$12702 ( \18732 , \18046 );
buf \U$12703 ( \18733 , \18046 );
buf \U$12704 ( \18734 , \18046 );
buf \U$12705 ( \18735 , \18046 );
buf \U$12706 ( \18736 , \18046 );
buf \U$12707 ( \18737 , \18046 );
buf \U$12708 ( \18738 , \18046 );
buf \U$12709 ( \18739 , \18046 );
buf \U$12710 ( \18740 , \18046 );
buf \U$12711 ( \18741 , \18046 );
buf \U$12712 ( \18742 , \18046 );
buf \U$12713 ( \18743 , \18046 );
buf \U$12714 ( \18744 , \18046 );
buf \U$12715 ( \18745 , \18046 );
buf \U$12716 ( \18746 , \18046 );
buf \U$12717 ( \18747 , \18046 );
buf \U$12718 ( \18748 , \18046 );
nor \U$12719 ( \18749 , \18033 , \18075 , \18035 , \18077 , \18039 , \18043 , \18046 , \18724 , \18725 , \18726 , \18727 , \18728 , \18729 , \18730 , \18731 , \18732 , \18733 , \18734 , \18735 , \18736 , \18737 , \18738 , \18739 , \18740 , \18741 , \18742 , \18743 , \18744 , \18745 , \18746 , \18747 , \18748 );
and \U$12720 ( \18750 , \7976 , \18749 );
buf \U$12721 ( \18751 , \18046 );
buf \U$12722 ( \18752 , \18046 );
buf \U$12723 ( \18753 , \18046 );
buf \U$12724 ( \18754 , \18046 );
buf \U$12725 ( \18755 , \18046 );
buf \U$12726 ( \18756 , \18046 );
buf \U$12727 ( \18757 , \18046 );
buf \U$12728 ( \18758 , \18046 );
buf \U$12729 ( \18759 , \18046 );
buf \U$12730 ( \18760 , \18046 );
buf \U$12731 ( \18761 , \18046 );
buf \U$12732 ( \18762 , \18046 );
buf \U$12733 ( \18763 , \18046 );
buf \U$12734 ( \18764 , \18046 );
buf \U$12735 ( \18765 , \18046 );
buf \U$12736 ( \18766 , \18046 );
buf \U$12737 ( \18767 , \18046 );
buf \U$12738 ( \18768 , \18046 );
buf \U$12739 ( \18769 , \18046 );
buf \U$12740 ( \18770 , \18046 );
buf \U$12741 ( \18771 , \18046 );
buf \U$12742 ( \18772 , \18046 );
buf \U$12743 ( \18773 , \18046 );
buf \U$12744 ( \18774 , \18046 );
buf \U$12745 ( \18775 , \18046 );
nor \U$12746 ( \18776 , \18074 , \18034 , \18035 , \18077 , \18039 , \18043 , \18046 , \18751 , \18752 , \18753 , \18754 , \18755 , \18756 , \18757 , \18758 , \18759 , \18760 , \18761 , \18762 , \18763 , \18764 , \18765 , \18766 , \18767 , \18768 , \18769 , \18770 , \18771 , \18772 , \18773 , \18774 , \18775 );
and \U$12747 ( \18777 , \8004 , \18776 );
buf \U$12748 ( \18778 , \18046 );
buf \U$12749 ( \18779 , \18046 );
buf \U$12750 ( \18780 , \18046 );
buf \U$12751 ( \18781 , \18046 );
buf \U$12752 ( \18782 , \18046 );
buf \U$12753 ( \18783 , \18046 );
buf \U$12754 ( \18784 , \18046 );
buf \U$12755 ( \18785 , \18046 );
buf \U$12756 ( \18786 , \18046 );
buf \U$12757 ( \18787 , \18046 );
buf \U$12758 ( \18788 , \18046 );
buf \U$12759 ( \18789 , \18046 );
buf \U$12760 ( \18790 , \18046 );
buf \U$12761 ( \18791 , \18046 );
buf \U$12762 ( \18792 , \18046 );
buf \U$12763 ( \18793 , \18046 );
buf \U$12764 ( \18794 , \18046 );
buf \U$12765 ( \18795 , \18046 );
buf \U$12766 ( \18796 , \18046 );
buf \U$12767 ( \18797 , \18046 );
buf \U$12768 ( \18798 , \18046 );
buf \U$12769 ( \18799 , \18046 );
buf \U$12770 ( \18800 , \18046 );
buf \U$12771 ( \18801 , \18046 );
buf \U$12772 ( \18802 , \18046 );
nor \U$12773 ( \18803 , \18033 , \18034 , \18035 , \18077 , \18039 , \18043 , \18046 , \18778 , \18779 , \18780 , \18781 , \18782 , \18783 , \18784 , \18785 , \18786 , \18787 , \18788 , \18789 , \18790 , \18791 , \18792 , \18793 , \18794 , \18795 , \18796 , \18797 , \18798 , \18799 , \18800 , \18801 , \18802 );
and \U$12774 ( \18804 , \8032 , \18803 );
buf \U$12775 ( \18805 , \18046 );
buf \U$12776 ( \18806 , \18046 );
buf \U$12777 ( \18807 , \18046 );
buf \U$12778 ( \18808 , \18046 );
buf \U$12779 ( \18809 , \18046 );
buf \U$12780 ( \18810 , \18046 );
buf \U$12781 ( \18811 , \18046 );
buf \U$12782 ( \18812 , \18046 );
buf \U$12783 ( \18813 , \18046 );
buf \U$12784 ( \18814 , \18046 );
buf \U$12785 ( \18815 , \18046 );
buf \U$12786 ( \18816 , \18046 );
buf \U$12787 ( \18817 , \18046 );
buf \U$12788 ( \18818 , \18046 );
buf \U$12789 ( \18819 , \18046 );
buf \U$12790 ( \18820 , \18046 );
buf \U$12791 ( \18821 , \18046 );
buf \U$12792 ( \18822 , \18046 );
buf \U$12793 ( \18823 , \18046 );
buf \U$12794 ( \18824 , \18046 );
buf \U$12795 ( \18825 , \18046 );
buf \U$12796 ( \18826 , \18046 );
buf \U$12797 ( \18827 , \18046 );
buf \U$12798 ( \18828 , \18046 );
buf \U$12799 ( \18829 , \18046 );
nor \U$12800 ( \18830 , \18074 , \18075 , \18076 , \18036 , \18039 , \18043 , \18046 , \18805 , \18806 , \18807 , \18808 , \18809 , \18810 , \18811 , \18812 , \18813 , \18814 , \18815 , \18816 , \18817 , \18818 , \18819 , \18820 , \18821 , \18822 , \18823 , \18824 , \18825 , \18826 , \18827 , \18828 , \18829 );
and \U$12801 ( \18831 , \8060 , \18830 );
buf \U$12802 ( \18832 , \18046 );
buf \U$12803 ( \18833 , \18046 );
buf \U$12804 ( \18834 , \18046 );
buf \U$12805 ( \18835 , \18046 );
buf \U$12806 ( \18836 , \18046 );
buf \U$12807 ( \18837 , \18046 );
buf \U$12808 ( \18838 , \18046 );
buf \U$12809 ( \18839 , \18046 );
buf \U$12810 ( \18840 , \18046 );
buf \U$12811 ( \18841 , \18046 );
buf \U$12812 ( \18842 , \18046 );
buf \U$12813 ( \18843 , \18046 );
buf \U$12814 ( \18844 , \18046 );
buf \U$12815 ( \18845 , \18046 );
buf \U$12816 ( \18846 , \18046 );
buf \U$12817 ( \18847 , \18046 );
buf \U$12818 ( \18848 , \18046 );
buf \U$12819 ( \18849 , \18046 );
buf \U$12820 ( \18850 , \18046 );
buf \U$12821 ( \18851 , \18046 );
buf \U$12822 ( \18852 , \18046 );
buf \U$12823 ( \18853 , \18046 );
buf \U$12824 ( \18854 , \18046 );
buf \U$12825 ( \18855 , \18046 );
buf \U$12826 ( \18856 , \18046 );
nor \U$12827 ( \18857 , \18033 , \18075 , \18076 , \18036 , \18039 , \18043 , \18046 , \18832 , \18833 , \18834 , \18835 , \18836 , \18837 , \18838 , \18839 , \18840 , \18841 , \18842 , \18843 , \18844 , \18845 , \18846 , \18847 , \18848 , \18849 , \18850 , \18851 , \18852 , \18853 , \18854 , \18855 , \18856 );
and \U$12828 ( \18858 , \8088 , \18857 );
buf \U$12829 ( \18859 , \18046 );
buf \U$12830 ( \18860 , \18046 );
buf \U$12831 ( \18861 , \18046 );
buf \U$12832 ( \18862 , \18046 );
buf \U$12833 ( \18863 , \18046 );
buf \U$12834 ( \18864 , \18046 );
buf \U$12835 ( \18865 , \18046 );
buf \U$12836 ( \18866 , \18046 );
buf \U$12837 ( \18867 , \18046 );
buf \U$12838 ( \18868 , \18046 );
buf \U$12839 ( \18869 , \18046 );
buf \U$12840 ( \18870 , \18046 );
buf \U$12841 ( \18871 , \18046 );
buf \U$12842 ( \18872 , \18046 );
buf \U$12843 ( \18873 , \18046 );
buf \U$12844 ( \18874 , \18046 );
buf \U$12845 ( \18875 , \18046 );
buf \U$12846 ( \18876 , \18046 );
buf \U$12847 ( \18877 , \18046 );
buf \U$12848 ( \18878 , \18046 );
buf \U$12849 ( \18879 , \18046 );
buf \U$12850 ( \18880 , \18046 );
buf \U$12851 ( \18881 , \18046 );
buf \U$12852 ( \18882 , \18046 );
buf \U$12853 ( \18883 , \18046 );
nor \U$12854 ( \18884 , \18074 , \18034 , \18076 , \18036 , \18039 , \18043 , \18046 , \18859 , \18860 , \18861 , \18862 , \18863 , \18864 , \18865 , \18866 , \18867 , \18868 , \18869 , \18870 , \18871 , \18872 , \18873 , \18874 , \18875 , \18876 , \18877 , \18878 , \18879 , \18880 , \18881 , \18882 , \18883 );
and \U$12855 ( \18885 , \8116 , \18884 );
buf \U$12856 ( \18886 , \18046 );
buf \U$12857 ( \18887 , \18046 );
buf \U$12858 ( \18888 , \18046 );
buf \U$12859 ( \18889 , \18046 );
buf \U$12860 ( \18890 , \18046 );
buf \U$12861 ( \18891 , \18046 );
buf \U$12862 ( \18892 , \18046 );
buf \U$12863 ( \18893 , \18046 );
buf \U$12864 ( \18894 , \18046 );
buf \U$12865 ( \18895 , \18046 );
buf \U$12866 ( \18896 , \18046 );
buf \U$12867 ( \18897 , \18046 );
buf \U$12868 ( \18898 , \18046 );
buf \U$12869 ( \18899 , \18046 );
buf \U$12870 ( \18900 , \18046 );
buf \U$12871 ( \18901 , \18046 );
buf \U$12872 ( \18902 , \18046 );
buf \U$12873 ( \18903 , \18046 );
buf \U$12874 ( \18904 , \18046 );
buf \U$12875 ( \18905 , \18046 );
buf \U$12876 ( \18906 , \18046 );
buf \U$12877 ( \18907 , \18046 );
buf \U$12878 ( \18908 , \18046 );
buf \U$12879 ( \18909 , \18046 );
buf \U$12880 ( \18910 , \18046 );
nor \U$12881 ( \18911 , \18033 , \18034 , \18076 , \18036 , \18039 , \18043 , \18046 , \18886 , \18887 , \18888 , \18889 , \18890 , \18891 , \18892 , \18893 , \18894 , \18895 , \18896 , \18897 , \18898 , \18899 , \18900 , \18901 , \18902 , \18903 , \18904 , \18905 , \18906 , \18907 , \18908 , \18909 , \18910 );
and \U$12882 ( \18912 , \8144 , \18911 );
buf \U$12883 ( \18913 , \18046 );
buf \U$12884 ( \18914 , \18046 );
buf \U$12885 ( \18915 , \18046 );
buf \U$12886 ( \18916 , \18046 );
buf \U$12887 ( \18917 , \18046 );
buf \U$12888 ( \18918 , \18046 );
buf \U$12889 ( \18919 , \18046 );
buf \U$12890 ( \18920 , \18046 );
buf \U$12891 ( \18921 , \18046 );
buf \U$12892 ( \18922 , \18046 );
buf \U$12893 ( \18923 , \18046 );
buf \U$12894 ( \18924 , \18046 );
buf \U$12895 ( \18925 , \18046 );
buf \U$12896 ( \18926 , \18046 );
buf \U$12897 ( \18927 , \18046 );
buf \U$12898 ( \18928 , \18046 );
buf \U$12899 ( \18929 , \18046 );
buf \U$12900 ( \18930 , \18046 );
buf \U$12901 ( \18931 , \18046 );
buf \U$12902 ( \18932 , \18046 );
buf \U$12903 ( \18933 , \18046 );
buf \U$12904 ( \18934 , \18046 );
buf \U$12905 ( \18935 , \18046 );
buf \U$12906 ( \18936 , \18046 );
buf \U$12907 ( \18937 , \18046 );
nor \U$12908 ( \18938 , \18074 , \18075 , \18035 , \18036 , \18039 , \18043 , \18046 , \18913 , \18914 , \18915 , \18916 , \18917 , \18918 , \18919 , \18920 , \18921 , \18922 , \18923 , \18924 , \18925 , \18926 , \18927 , \18928 , \18929 , \18930 , \18931 , \18932 , \18933 , \18934 , \18935 , \18936 , \18937 );
and \U$12909 ( \18939 , \8172 , \18938 );
buf \U$12910 ( \18940 , \18046 );
buf \U$12911 ( \18941 , \18046 );
buf \U$12912 ( \18942 , \18046 );
buf \U$12913 ( \18943 , \18046 );
buf \U$12914 ( \18944 , \18046 );
buf \U$12915 ( \18945 , \18046 );
buf \U$12916 ( \18946 , \18046 );
buf \U$12917 ( \18947 , \18046 );
buf \U$12918 ( \18948 , \18046 );
buf \U$12919 ( \18949 , \18046 );
buf \U$12920 ( \18950 , \18046 );
buf \U$12921 ( \18951 , \18046 );
buf \U$12922 ( \18952 , \18046 );
buf \U$12923 ( \18953 , \18046 );
buf \U$12924 ( \18954 , \18046 );
buf \U$12925 ( \18955 , \18046 );
buf \U$12926 ( \18956 , \18046 );
buf \U$12927 ( \18957 , \18046 );
buf \U$12928 ( \18958 , \18046 );
buf \U$12929 ( \18959 , \18046 );
buf \U$12930 ( \18960 , \18046 );
buf \U$12931 ( \18961 , \18046 );
buf \U$12932 ( \18962 , \18046 );
buf \U$12933 ( \18963 , \18046 );
buf \U$12934 ( \18964 , \18046 );
nor \U$12935 ( \18965 , \18033 , \18075 , \18035 , \18036 , \18039 , \18043 , \18046 , \18940 , \18941 , \18942 , \18943 , \18944 , \18945 , \18946 , \18947 , \18948 , \18949 , \18950 , \18951 , \18952 , \18953 , \18954 , \18955 , \18956 , \18957 , \18958 , \18959 , \18960 , \18961 , \18962 , \18963 , \18964 );
and \U$12936 ( \18966 , \8200 , \18965 );
buf \U$12937 ( \18967 , \18046 );
buf \U$12938 ( \18968 , \18046 );
buf \U$12939 ( \18969 , \18046 );
buf \U$12940 ( \18970 , \18046 );
buf \U$12941 ( \18971 , \18046 );
buf \U$12942 ( \18972 , \18046 );
buf \U$12943 ( \18973 , \18046 );
buf \U$12944 ( \18974 , \18046 );
buf \U$12945 ( \18975 , \18046 );
buf \U$12946 ( \18976 , \18046 );
buf \U$12947 ( \18977 , \18046 );
buf \U$12948 ( \18978 , \18046 );
buf \U$12949 ( \18979 , \18046 );
buf \U$12950 ( \18980 , \18046 );
buf \U$12951 ( \18981 , \18046 );
buf \U$12952 ( \18982 , \18046 );
buf \U$12953 ( \18983 , \18046 );
buf \U$12954 ( \18984 , \18046 );
buf \U$12955 ( \18985 , \18046 );
buf \U$12956 ( \18986 , \18046 );
buf \U$12957 ( \18987 , \18046 );
buf \U$12958 ( \18988 , \18046 );
buf \U$12959 ( \18989 , \18046 );
buf \U$12960 ( \18990 , \18046 );
buf \U$12961 ( \18991 , \18046 );
nor \U$12962 ( \18992 , \18074 , \18034 , \18035 , \18036 , \18039 , \18043 , \18046 , \18967 , \18968 , \18969 , \18970 , \18971 , \18972 , \18973 , \18974 , \18975 , \18976 , \18977 , \18978 , \18979 , \18980 , \18981 , \18982 , \18983 , \18984 , \18985 , \18986 , \18987 , \18988 , \18989 , \18990 , \18991 );
and \U$12963 ( \18993 , \8228 , \18992 );
or \U$12964 ( \18994 , \18588 , \18615 , \18642 , \18669 , \18696 , \18723 , \18750 , \18777 , \18804 , \18831 , \18858 , \18885 , \18912 , \18939 , \18966 , \18993 );
buf \U$12965 ( \18995 , \18046 );
not \U$12966 ( \18996 , \18995 );
buf \U$12967 ( \18997 , \18034 );
buf \U$12968 ( \18998 , \18035 );
buf \U$12969 ( \18999 , \18036 );
buf \U$12970 ( \19000 , \18039 );
buf \U$12971 ( \19001 , \18043 );
buf \U$12972 ( \19002 , \18046 );
buf \U$12973 ( \19003 , \18046 );
buf \U$12974 ( \19004 , \18046 );
buf \U$12975 ( \19005 , \18046 );
buf \U$12976 ( \19006 , \18046 );
buf \U$12977 ( \19007 , \18046 );
buf \U$12978 ( \19008 , \18046 );
buf \U$12979 ( \19009 , \18046 );
buf \U$12980 ( \19010 , \18046 );
buf \U$12981 ( \19011 , \18046 );
buf \U$12982 ( \19012 , \18046 );
buf \U$12983 ( \19013 , \18046 );
buf \U$12984 ( \19014 , \18046 );
buf \U$12985 ( \19015 , \18046 );
buf \U$12986 ( \19016 , \18046 );
buf \U$12987 ( \19017 , \18046 );
buf \U$12988 ( \19018 , \18046 );
buf \U$12989 ( \19019 , \18046 );
buf \U$12990 ( \19020 , \18046 );
buf \U$12991 ( \19021 , \18046 );
buf \U$12992 ( \19022 , \18046 );
buf \U$12993 ( \19023 , \18046 );
buf \U$12994 ( \19024 , \18046 );
buf \U$12995 ( \19025 , \18046 );
buf \U$12996 ( \19026 , \18046 );
buf \U$12997 ( \19027 , \18033 );
or \U$12998 ( \19028 , \18997 , \18998 , \18999 , \19000 , \19001 , \19002 , \19003 , \19004 , \19005 , \19006 , \19007 , \19008 , \19009 , \19010 , \19011 , \19012 , \19013 , \19014 , \19015 , \19016 , \19017 , \19018 , \19019 , \19020 , \19021 , \19022 , \19023 , \19024 , \19025 , \19026 , \19027 );
nand \U$12999 ( \19029 , \18996 , \19028 );
buf \U$13000 ( \19030 , \19029 );
buf \U$13001 ( \19031 , \18046 );
not \U$13002 ( \19032 , \19031 );
buf \U$13003 ( \19033 , \18043 );
buf \U$13004 ( \19034 , \18046 );
buf \U$13005 ( \19035 , \18046 );
buf \U$13006 ( \19036 , \18046 );
buf \U$13007 ( \19037 , \18046 );
buf \U$13008 ( \19038 , \18046 );
buf \U$13009 ( \19039 , \18046 );
buf \U$13010 ( \19040 , \18046 );
buf \U$13011 ( \19041 , \18046 );
buf \U$13012 ( \19042 , \18046 );
buf \U$13013 ( \19043 , \18046 );
buf \U$13014 ( \19044 , \18046 );
buf \U$13015 ( \19045 , \18046 );
buf \U$13016 ( \19046 , \18046 );
buf \U$13017 ( \19047 , \18046 );
buf \U$13018 ( \19048 , \18046 );
buf \U$13019 ( \19049 , \18046 );
buf \U$13020 ( \19050 , \18046 );
buf \U$13021 ( \19051 , \18046 );
buf \U$13022 ( \19052 , \18046 );
buf \U$13023 ( \19053 , \18046 );
buf \U$13024 ( \19054 , \18046 );
buf \U$13025 ( \19055 , \18046 );
buf \U$13026 ( \19056 , \18046 );
buf \U$13027 ( \19057 , \18046 );
buf \U$13028 ( \19058 , \18046 );
buf \U$13029 ( \19059 , \18039 );
buf \U$13030 ( \19060 , \18033 );
buf \U$13031 ( \19061 , \18034 );
buf \U$13032 ( \19062 , \18035 );
buf \U$13033 ( \19063 , \18036 );
or \U$13034 ( \19064 , \19060 , \19061 , \19062 , \19063 );
and \U$13035 ( \19065 , \19059 , \19064 );
or \U$13036 ( \19066 , \19033 , \19034 , \19035 , \19036 , \19037 , \19038 , \19039 , \19040 , \19041 , \19042 , \19043 , \19044 , \19045 , \19046 , \19047 , \19048 , \19049 , \19050 , \19051 , \19052 , \19053 , \19054 , \19055 , \19056 , \19057 , \19058 , \19065 );
and \U$13037 ( \19067 , \19032 , \19066 );
buf \U$13038 ( \19068 , \19067 );
or \U$13039 ( \19069 , \19030 , \19068 );
_DC g615b ( \19070_nG615b , \18994 , \19069 );
buf \U$13040 ( \19071 , \19070_nG615b );
xor \U$13041 ( \19072 , \18561 , \19071 );
buf \U$13042 ( \19073 , RIb7b9590_247);
and \U$13043 ( \19074 , \7126 , \18587 );
and \U$13044 ( \19075 , \7128 , \18614 );
and \U$13045 ( \19076 , \8338 , \18641 );
and \U$13046 ( \19077 , \8340 , \18668 );
and \U$13047 ( \19078 , \8342 , \18695 );
and \U$13048 ( \19079 , \8344 , \18722 );
and \U$13049 ( \19080 , \8346 , \18749 );
and \U$13050 ( \19081 , \8348 , \18776 );
and \U$13051 ( \19082 , \8350 , \18803 );
and \U$13052 ( \19083 , \8352 , \18830 );
and \U$13053 ( \19084 , \8354 , \18857 );
and \U$13054 ( \19085 , \8356 , \18884 );
and \U$13055 ( \19086 , \8358 , \18911 );
and \U$13056 ( \19087 , \8360 , \18938 );
and \U$13057 ( \19088 , \8362 , \18965 );
and \U$13058 ( \19089 , \8364 , \18992 );
or \U$13059 ( \19090 , \19074 , \19075 , \19076 , \19077 , \19078 , \19079 , \19080 , \19081 , \19082 , \19083 , \19084 , \19085 , \19086 , \19087 , \19088 , \19089 );
_DC g6170 ( \19091_nG6170 , \19090 , \19069 );
buf \U$13060 ( \19092 , \19091_nG6170 );
xor \U$13061 ( \19093 , \19073 , \19092 );
or \U$13062 ( \19094 , \19072 , \19093 );
buf \U$13063 ( \19095 , RIb7b9518_248);
and \U$13064 ( \19096 , \7136 , \18587 );
and \U$13065 ( \19097 , \7138 , \18614 );
and \U$13066 ( \19098 , \8374 , \18641 );
and \U$13067 ( \19099 , \8376 , \18668 );
and \U$13068 ( \19100 , \8378 , \18695 );
and \U$13069 ( \19101 , \8380 , \18722 );
and \U$13070 ( \19102 , \8382 , \18749 );
and \U$13071 ( \19103 , \8384 , \18776 );
and \U$13072 ( \19104 , \8386 , \18803 );
and \U$13073 ( \19105 , \8388 , \18830 );
and \U$13074 ( \19106 , \8390 , \18857 );
and \U$13075 ( \19107 , \8392 , \18884 );
and \U$13076 ( \19108 , \8394 , \18911 );
and \U$13077 ( \19109 , \8396 , \18938 );
and \U$13078 ( \19110 , \8398 , \18965 );
and \U$13079 ( \19111 , \8400 , \18992 );
or \U$13080 ( \19112 , \19096 , \19097 , \19098 , \19099 , \19100 , \19101 , \19102 , \19103 , \19104 , \19105 , \19106 , \19107 , \19108 , \19109 , \19110 , \19111 );
_DC g6186 ( \19113_nG6186 , \19112 , \19069 );
buf \U$13081 ( \19114 , \19113_nG6186 );
xor \U$13082 ( \19115 , \19095 , \19114 );
or \U$13083 ( \19116 , \19094 , \19115 );
buf \U$13084 ( \19117 , RIb7b94a0_249);
and \U$13085 ( \19118 , \7146 , \18587 );
and \U$13086 ( \19119 , \7148 , \18614 );
and \U$13087 ( \19120 , \8410 , \18641 );
and \U$13088 ( \19121 , \8412 , \18668 );
and \U$13089 ( \19122 , \8414 , \18695 );
and \U$13090 ( \19123 , \8416 , \18722 );
and \U$13091 ( \19124 , \8418 , \18749 );
and \U$13092 ( \19125 , \8420 , \18776 );
and \U$13093 ( \19126 , \8422 , \18803 );
and \U$13094 ( \19127 , \8424 , \18830 );
and \U$13095 ( \19128 , \8426 , \18857 );
and \U$13096 ( \19129 , \8428 , \18884 );
and \U$13097 ( \19130 , \8430 , \18911 );
and \U$13098 ( \19131 , \8432 , \18938 );
and \U$13099 ( \19132 , \8434 , \18965 );
and \U$13100 ( \19133 , \8436 , \18992 );
or \U$13101 ( \19134 , \19118 , \19119 , \19120 , \19121 , \19122 , \19123 , \19124 , \19125 , \19126 , \19127 , \19128 , \19129 , \19130 , \19131 , \19132 , \19133 );
_DC g619c ( \19135_nG619c , \19134 , \19069 );
buf \U$13102 ( \19136 , \19135_nG619c );
xor \U$13103 ( \19137 , \19117 , \19136 );
or \U$13104 ( \19138 , \19116 , \19137 );
buf \U$13105 ( \19139 , RIb7b9428_250);
and \U$13106 ( \19140 , \7156 , \18587 );
and \U$13107 ( \19141 , \7158 , \18614 );
and \U$13108 ( \19142 , \8446 , \18641 );
and \U$13109 ( \19143 , \8448 , \18668 );
and \U$13110 ( \19144 , \8450 , \18695 );
and \U$13111 ( \19145 , \8452 , \18722 );
and \U$13112 ( \19146 , \8454 , \18749 );
and \U$13113 ( \19147 , \8456 , \18776 );
and \U$13114 ( \19148 , \8458 , \18803 );
and \U$13115 ( \19149 , \8460 , \18830 );
and \U$13116 ( \19150 , \8462 , \18857 );
and \U$13117 ( \19151 , \8464 , \18884 );
and \U$13118 ( \19152 , \8466 , \18911 );
and \U$13119 ( \19153 , \8468 , \18938 );
and \U$13120 ( \19154 , \8470 , \18965 );
and \U$13121 ( \19155 , \8472 , \18992 );
or \U$13122 ( \19156 , \19140 , \19141 , \19142 , \19143 , \19144 , \19145 , \19146 , \19147 , \19148 , \19149 , \19150 , \19151 , \19152 , \19153 , \19154 , \19155 );
_DC g61b2 ( \19157_nG61b2 , \19156 , \19069 );
buf \U$13123 ( \19158 , \19157_nG61b2 );
xor \U$13124 ( \19159 , \19139 , \19158 );
or \U$13125 ( \19160 , \19138 , \19159 );
buf \U$13126 ( \19161 , RIb7b93b0_251);
and \U$13127 ( \19162 , \7166 , \18587 );
and \U$13128 ( \19163 , \7168 , \18614 );
and \U$13129 ( \19164 , \8482 , \18641 );
and \U$13130 ( \19165 , \8484 , \18668 );
and \U$13131 ( \19166 , \8486 , \18695 );
and \U$13132 ( \19167 , \8488 , \18722 );
and \U$13133 ( \19168 , \8490 , \18749 );
and \U$13134 ( \19169 , \8492 , \18776 );
and \U$13135 ( \19170 , \8494 , \18803 );
and \U$13136 ( \19171 , \8496 , \18830 );
and \U$13137 ( \19172 , \8498 , \18857 );
and \U$13138 ( \19173 , \8500 , \18884 );
and \U$13139 ( \19174 , \8502 , \18911 );
and \U$13140 ( \19175 , \8504 , \18938 );
and \U$13141 ( \19176 , \8506 , \18965 );
and \U$13142 ( \19177 , \8508 , \18992 );
or \U$13143 ( \19178 , \19162 , \19163 , \19164 , \19165 , \19166 , \19167 , \19168 , \19169 , \19170 , \19171 , \19172 , \19173 , \19174 , \19175 , \19176 , \19177 );
_DC g61c8 ( \19179_nG61c8 , \19178 , \19069 );
buf \U$13144 ( \19180 , \19179_nG61c8 );
xor \U$13145 ( \19181 , \19161 , \19180 );
or \U$13146 ( \19182 , \19160 , \19181 );
buf \U$13147 ( \19183 , RIb7af720_252);
and \U$13148 ( \19184 , \7176 , \18587 );
and \U$13149 ( \19185 , \7178 , \18614 );
and \U$13150 ( \19186 , \8518 , \18641 );
and \U$13151 ( \19187 , \8520 , \18668 );
and \U$13152 ( \19188 , \8522 , \18695 );
and \U$13153 ( \19189 , \8524 , \18722 );
and \U$13154 ( \19190 , \8526 , \18749 );
and \U$13155 ( \19191 , \8528 , \18776 );
and \U$13156 ( \19192 , \8530 , \18803 );
and \U$13157 ( \19193 , \8532 , \18830 );
and \U$13158 ( \19194 , \8534 , \18857 );
and \U$13159 ( \19195 , \8536 , \18884 );
and \U$13160 ( \19196 , \8538 , \18911 );
and \U$13161 ( \19197 , \8540 , \18938 );
and \U$13162 ( \19198 , \8542 , \18965 );
and \U$13163 ( \19199 , \8544 , \18992 );
or \U$13164 ( \19200 , \19184 , \19185 , \19186 , \19187 , \19188 , \19189 , \19190 , \19191 , \19192 , \19193 , \19194 , \19195 , \19196 , \19197 , \19198 , \19199 );
_DC g61de ( \19201_nG61de , \19200 , \19069 );
buf \U$13165 ( \19202 , \19201_nG61de );
xor \U$13166 ( \19203 , \19183 , \19202 );
or \U$13167 ( \19204 , \19182 , \19203 );
buf \U$13168 ( \19205 , RIb7af6a8_253);
and \U$13169 ( \19206 , \7186 , \18587 );
and \U$13170 ( \19207 , \7188 , \18614 );
and \U$13171 ( \19208 , \8554 , \18641 );
and \U$13172 ( \19209 , \8556 , \18668 );
and \U$13173 ( \19210 , \8558 , \18695 );
and \U$13174 ( \19211 , \8560 , \18722 );
and \U$13175 ( \19212 , \8562 , \18749 );
and \U$13176 ( \19213 , \8564 , \18776 );
and \U$13177 ( \19214 , \8566 , \18803 );
and \U$13178 ( \19215 , \8568 , \18830 );
and \U$13179 ( \19216 , \8570 , \18857 );
and \U$13180 ( \19217 , \8572 , \18884 );
and \U$13181 ( \19218 , \8574 , \18911 );
and \U$13182 ( \19219 , \8576 , \18938 );
and \U$13183 ( \19220 , \8578 , \18965 );
and \U$13184 ( \19221 , \8580 , \18992 );
or \U$13185 ( \19222 , \19206 , \19207 , \19208 , \19209 , \19210 , \19211 , \19212 , \19213 , \19214 , \19215 , \19216 , \19217 , \19218 , \19219 , \19220 , \19221 );
_DC g61f4 ( \19223_nG61f4 , \19222 , \19069 );
buf \U$13186 ( \19224 , \19223_nG61f4 );
xor \U$13187 ( \19225 , \19205 , \19224 );
or \U$13188 ( \19226 , \19204 , \19225 );
not \U$13189 ( \19227 , \19226 );
buf \U$13190 ( \19228 , \19227 );
and \U$13191 ( \19229 , \18560 , \19228 );
buf \U$13192 ( \19230 , RIb7af630_254);
buf \U$13193 ( \19231 , \18046 );
buf \U$13194 ( \19232 , \18046 );
buf \U$13195 ( \19233 , \18046 );
buf \U$13196 ( \19234 , \18046 );
buf \U$13197 ( \19235 , \18046 );
buf \U$13198 ( \19236 , \18046 );
buf \U$13199 ( \19237 , \18046 );
buf \U$13200 ( \19238 , \18046 );
buf \U$13201 ( \19239 , \18046 );
buf \U$13202 ( \19240 , \18046 );
buf \U$13203 ( \19241 , \18046 );
buf \U$13204 ( \19242 , \18046 );
buf \U$13205 ( \19243 , \18046 );
buf \U$13206 ( \19244 , \18046 );
buf \U$13207 ( \19245 , \18046 );
buf \U$13208 ( \19246 , \18046 );
buf \U$13209 ( \19247 , \18046 );
buf \U$13210 ( \19248 , \18046 );
buf \U$13211 ( \19249 , \18046 );
buf \U$13212 ( \19250 , \18046 );
buf \U$13213 ( \19251 , \18046 );
buf \U$13214 ( \19252 , \18046 );
buf \U$13215 ( \19253 , \18046 );
buf \U$13216 ( \19254 , \18046 );
buf \U$13217 ( \19255 , \18046 );
nor \U$13218 ( \19256 , \18033 , \18034 , \18035 , \18036 , \18040 , \18043 , \18046 , \19231 , \19232 , \19233 , \19234 , \19235 , \19236 , \19237 , \19238 , \19239 , \19240 , \19241 , \19242 , \19243 , \19244 , \19245 , \19246 , \19247 , \19248 , \19249 , \19250 , \19251 , \19252 , \19253 , \19254 , \19255 );
and \U$13219 ( \19257 , \7198 , \19256 );
buf \U$13220 ( \19258 , \18046 );
buf \U$13221 ( \19259 , \18046 );
buf \U$13222 ( \19260 , \18046 );
buf \U$13223 ( \19261 , \18046 );
buf \U$13224 ( \19262 , \18046 );
buf \U$13225 ( \19263 , \18046 );
buf \U$13226 ( \19264 , \18046 );
buf \U$13227 ( \19265 , \18046 );
buf \U$13228 ( \19266 , \18046 );
buf \U$13229 ( \19267 , \18046 );
buf \U$13230 ( \19268 , \18046 );
buf \U$13231 ( \19269 , \18046 );
buf \U$13232 ( \19270 , \18046 );
buf \U$13233 ( \19271 , \18046 );
buf \U$13234 ( \19272 , \18046 );
buf \U$13235 ( \19273 , \18046 );
buf \U$13236 ( \19274 , \18046 );
buf \U$13237 ( \19275 , \18046 );
buf \U$13238 ( \19276 , \18046 );
buf \U$13239 ( \19277 , \18046 );
buf \U$13240 ( \19278 , \18046 );
buf \U$13241 ( \19279 , \18046 );
buf \U$13242 ( \19280 , \18046 );
buf \U$13243 ( \19281 , \18046 );
buf \U$13244 ( \19282 , \18046 );
nor \U$13245 ( \19283 , \18074 , \18075 , \18076 , \18077 , \18039 , \18043 , \18046 , \19258 , \19259 , \19260 , \19261 , \19262 , \19263 , \19264 , \19265 , \19266 , \19267 , \19268 , \19269 , \19270 , \19271 , \19272 , \19273 , \19274 , \19275 , \19276 , \19277 , \19278 , \19279 , \19280 , \19281 , \19282 );
and \U$13246 ( \19284 , \7200 , \19283 );
buf \U$13247 ( \19285 , \18046 );
buf \U$13248 ( \19286 , \18046 );
buf \U$13249 ( \19287 , \18046 );
buf \U$13250 ( \19288 , \18046 );
buf \U$13251 ( \19289 , \18046 );
buf \U$13252 ( \19290 , \18046 );
buf \U$13253 ( \19291 , \18046 );
buf \U$13254 ( \19292 , \18046 );
buf \U$13255 ( \19293 , \18046 );
buf \U$13256 ( \19294 , \18046 );
buf \U$13257 ( \19295 , \18046 );
buf \U$13258 ( \19296 , \18046 );
buf \U$13259 ( \19297 , \18046 );
buf \U$13260 ( \19298 , \18046 );
buf \U$13261 ( \19299 , \18046 );
buf \U$13262 ( \19300 , \18046 );
buf \U$13263 ( \19301 , \18046 );
buf \U$13264 ( \19302 , \18046 );
buf \U$13265 ( \19303 , \18046 );
buf \U$13266 ( \19304 , \18046 );
buf \U$13267 ( \19305 , \18046 );
buf \U$13268 ( \19306 , \18046 );
buf \U$13269 ( \19307 , \18046 );
buf \U$13270 ( \19308 , \18046 );
buf \U$13271 ( \19309 , \18046 );
nor \U$13272 ( \19310 , \18033 , \18075 , \18076 , \18077 , \18039 , \18043 , \18046 , \19285 , \19286 , \19287 , \19288 , \19289 , \19290 , \19291 , \19292 , \19293 , \19294 , \19295 , \19296 , \19297 , \19298 , \19299 , \19300 , \19301 , \19302 , \19303 , \19304 , \19305 , \19306 , \19307 , \19308 , \19309 );
and \U$13273 ( \19311 , \8645 , \19310 );
buf \U$13274 ( \19312 , \18046 );
buf \U$13275 ( \19313 , \18046 );
buf \U$13276 ( \19314 , \18046 );
buf \U$13277 ( \19315 , \18046 );
buf \U$13278 ( \19316 , \18046 );
buf \U$13279 ( \19317 , \18046 );
buf \U$13280 ( \19318 , \18046 );
buf \U$13281 ( \19319 , \18046 );
buf \U$13282 ( \19320 , \18046 );
buf \U$13283 ( \19321 , \18046 );
buf \U$13284 ( \19322 , \18046 );
buf \U$13285 ( \19323 , \18046 );
buf \U$13286 ( \19324 , \18046 );
buf \U$13287 ( \19325 , \18046 );
buf \U$13288 ( \19326 , \18046 );
buf \U$13289 ( \19327 , \18046 );
buf \U$13290 ( \19328 , \18046 );
buf \U$13291 ( \19329 , \18046 );
buf \U$13292 ( \19330 , \18046 );
buf \U$13293 ( \19331 , \18046 );
buf \U$13294 ( \19332 , \18046 );
buf \U$13295 ( \19333 , \18046 );
buf \U$13296 ( \19334 , \18046 );
buf \U$13297 ( \19335 , \18046 );
buf \U$13298 ( \19336 , \18046 );
nor \U$13299 ( \19337 , \18074 , \18034 , \18076 , \18077 , \18039 , \18043 , \18046 , \19312 , \19313 , \19314 , \19315 , \19316 , \19317 , \19318 , \19319 , \19320 , \19321 , \19322 , \19323 , \19324 , \19325 , \19326 , \19327 , \19328 , \19329 , \19330 , \19331 , \19332 , \19333 , \19334 , \19335 , \19336 );
and \U$13300 ( \19338 , \8673 , \19337 );
buf \U$13301 ( \19339 , \18046 );
buf \U$13302 ( \19340 , \18046 );
buf \U$13303 ( \19341 , \18046 );
buf \U$13304 ( \19342 , \18046 );
buf \U$13305 ( \19343 , \18046 );
buf \U$13306 ( \19344 , \18046 );
buf \U$13307 ( \19345 , \18046 );
buf \U$13308 ( \19346 , \18046 );
buf \U$13309 ( \19347 , \18046 );
buf \U$13310 ( \19348 , \18046 );
buf \U$13311 ( \19349 , \18046 );
buf \U$13312 ( \19350 , \18046 );
buf \U$13313 ( \19351 , \18046 );
buf \U$13314 ( \19352 , \18046 );
buf \U$13315 ( \19353 , \18046 );
buf \U$13316 ( \19354 , \18046 );
buf \U$13317 ( \19355 , \18046 );
buf \U$13318 ( \19356 , \18046 );
buf \U$13319 ( \19357 , \18046 );
buf \U$13320 ( \19358 , \18046 );
buf \U$13321 ( \19359 , \18046 );
buf \U$13322 ( \19360 , \18046 );
buf \U$13323 ( \19361 , \18046 );
buf \U$13324 ( \19362 , \18046 );
buf \U$13325 ( \19363 , \18046 );
nor \U$13326 ( \19364 , \18033 , \18034 , \18076 , \18077 , \18039 , \18043 , \18046 , \19339 , \19340 , \19341 , \19342 , \19343 , \19344 , \19345 , \19346 , \19347 , \19348 , \19349 , \19350 , \19351 , \19352 , \19353 , \19354 , \19355 , \19356 , \19357 , \19358 , \19359 , \19360 , \19361 , \19362 , \19363 );
and \U$13327 ( \19365 , \8701 , \19364 );
buf \U$13328 ( \19366 , \18046 );
buf \U$13329 ( \19367 , \18046 );
buf \U$13330 ( \19368 , \18046 );
buf \U$13331 ( \19369 , \18046 );
buf \U$13332 ( \19370 , \18046 );
buf \U$13333 ( \19371 , \18046 );
buf \U$13334 ( \19372 , \18046 );
buf \U$13335 ( \19373 , \18046 );
buf \U$13336 ( \19374 , \18046 );
buf \U$13337 ( \19375 , \18046 );
buf \U$13338 ( \19376 , \18046 );
buf \U$13339 ( \19377 , \18046 );
buf \U$13340 ( \19378 , \18046 );
buf \U$13341 ( \19379 , \18046 );
buf \U$13342 ( \19380 , \18046 );
buf \U$13343 ( \19381 , \18046 );
buf \U$13344 ( \19382 , \18046 );
buf \U$13345 ( \19383 , \18046 );
buf \U$13346 ( \19384 , \18046 );
buf \U$13347 ( \19385 , \18046 );
buf \U$13348 ( \19386 , \18046 );
buf \U$13349 ( \19387 , \18046 );
buf \U$13350 ( \19388 , \18046 );
buf \U$13351 ( \19389 , \18046 );
buf \U$13352 ( \19390 , \18046 );
nor \U$13353 ( \19391 , \18074 , \18075 , \18035 , \18077 , \18039 , \18043 , \18046 , \19366 , \19367 , \19368 , \19369 , \19370 , \19371 , \19372 , \19373 , \19374 , \19375 , \19376 , \19377 , \19378 , \19379 , \19380 , \19381 , \19382 , \19383 , \19384 , \19385 , \19386 , \19387 , \19388 , \19389 , \19390 );
and \U$13354 ( \19392 , \8729 , \19391 );
buf \U$13355 ( \19393 , \18046 );
buf \U$13356 ( \19394 , \18046 );
buf \U$13357 ( \19395 , \18046 );
buf \U$13358 ( \19396 , \18046 );
buf \U$13359 ( \19397 , \18046 );
buf \U$13360 ( \19398 , \18046 );
buf \U$13361 ( \19399 , \18046 );
buf \U$13362 ( \19400 , \18046 );
buf \U$13363 ( \19401 , \18046 );
buf \U$13364 ( \19402 , \18046 );
buf \U$13365 ( \19403 , \18046 );
buf \U$13366 ( \19404 , \18046 );
buf \U$13367 ( \19405 , \18046 );
buf \U$13368 ( \19406 , \18046 );
buf \U$13369 ( \19407 , \18046 );
buf \U$13370 ( \19408 , \18046 );
buf \U$13371 ( \19409 , \18046 );
buf \U$13372 ( \19410 , \18046 );
buf \U$13373 ( \19411 , \18046 );
buf \U$13374 ( \19412 , \18046 );
buf \U$13375 ( \19413 , \18046 );
buf \U$13376 ( \19414 , \18046 );
buf \U$13377 ( \19415 , \18046 );
buf \U$13378 ( \19416 , \18046 );
buf \U$13379 ( \19417 , \18046 );
nor \U$13380 ( \19418 , \18033 , \18075 , \18035 , \18077 , \18039 , \18043 , \18046 , \19393 , \19394 , \19395 , \19396 , \19397 , \19398 , \19399 , \19400 , \19401 , \19402 , \19403 , \19404 , \19405 , \19406 , \19407 , \19408 , \19409 , \19410 , \19411 , \19412 , \19413 , \19414 , \19415 , \19416 , \19417 );
and \U$13381 ( \19419 , \8757 , \19418 );
buf \U$13382 ( \19420 , \18046 );
buf \U$13383 ( \19421 , \18046 );
buf \U$13384 ( \19422 , \18046 );
buf \U$13385 ( \19423 , \18046 );
buf \U$13386 ( \19424 , \18046 );
buf \U$13387 ( \19425 , \18046 );
buf \U$13388 ( \19426 , \18046 );
buf \U$13389 ( \19427 , \18046 );
buf \U$13390 ( \19428 , \18046 );
buf \U$13391 ( \19429 , \18046 );
buf \U$13392 ( \19430 , \18046 );
buf \U$13393 ( \19431 , \18046 );
buf \U$13394 ( \19432 , \18046 );
buf \U$13395 ( \19433 , \18046 );
buf \U$13396 ( \19434 , \18046 );
buf \U$13397 ( \19435 , \18046 );
buf \U$13398 ( \19436 , \18046 );
buf \U$13399 ( \19437 , \18046 );
buf \U$13400 ( \19438 , \18046 );
buf \U$13401 ( \19439 , \18046 );
buf \U$13402 ( \19440 , \18046 );
buf \U$13403 ( \19441 , \18046 );
buf \U$13404 ( \19442 , \18046 );
buf \U$13405 ( \19443 , \18046 );
buf \U$13406 ( \19444 , \18046 );
nor \U$13407 ( \19445 , \18074 , \18034 , \18035 , \18077 , \18039 , \18043 , \18046 , \19420 , \19421 , \19422 , \19423 , \19424 , \19425 , \19426 , \19427 , \19428 , \19429 , \19430 , \19431 , \19432 , \19433 , \19434 , \19435 , \19436 , \19437 , \19438 , \19439 , \19440 , \19441 , \19442 , \19443 , \19444 );
and \U$13408 ( \19446 , \8785 , \19445 );
buf \U$13409 ( \19447 , \18046 );
buf \U$13410 ( \19448 , \18046 );
buf \U$13411 ( \19449 , \18046 );
buf \U$13412 ( \19450 , \18046 );
buf \U$13413 ( \19451 , \18046 );
buf \U$13414 ( \19452 , \18046 );
buf \U$13415 ( \19453 , \18046 );
buf \U$13416 ( \19454 , \18046 );
buf \U$13417 ( \19455 , \18046 );
buf \U$13418 ( \19456 , \18046 );
buf \U$13419 ( \19457 , \18046 );
buf \U$13420 ( \19458 , \18046 );
buf \U$13421 ( \19459 , \18046 );
buf \U$13422 ( \19460 , \18046 );
buf \U$13423 ( \19461 , \18046 );
buf \U$13424 ( \19462 , \18046 );
buf \U$13425 ( \19463 , \18046 );
buf \U$13426 ( \19464 , \18046 );
buf \U$13427 ( \19465 , \18046 );
buf \U$13428 ( \19466 , \18046 );
buf \U$13429 ( \19467 , \18046 );
buf \U$13430 ( \19468 , \18046 );
buf \U$13431 ( \19469 , \18046 );
buf \U$13432 ( \19470 , \18046 );
buf \U$13433 ( \19471 , \18046 );
nor \U$13434 ( \19472 , \18033 , \18034 , \18035 , \18077 , \18039 , \18043 , \18046 , \19447 , \19448 , \19449 , \19450 , \19451 , \19452 , \19453 , \19454 , \19455 , \19456 , \19457 , \19458 , \19459 , \19460 , \19461 , \19462 , \19463 , \19464 , \19465 , \19466 , \19467 , \19468 , \19469 , \19470 , \19471 );
and \U$13435 ( \19473 , \8813 , \19472 );
buf \U$13436 ( \19474 , \18046 );
buf \U$13437 ( \19475 , \18046 );
buf \U$13438 ( \19476 , \18046 );
buf \U$13439 ( \19477 , \18046 );
buf \U$13440 ( \19478 , \18046 );
buf \U$13441 ( \19479 , \18046 );
buf \U$13442 ( \19480 , \18046 );
buf \U$13443 ( \19481 , \18046 );
buf \U$13444 ( \19482 , \18046 );
buf \U$13445 ( \19483 , \18046 );
buf \U$13446 ( \19484 , \18046 );
buf \U$13447 ( \19485 , \18046 );
buf \U$13448 ( \19486 , \18046 );
buf \U$13449 ( \19487 , \18046 );
buf \U$13450 ( \19488 , \18046 );
buf \U$13451 ( \19489 , \18046 );
buf \U$13452 ( \19490 , \18046 );
buf \U$13453 ( \19491 , \18046 );
buf \U$13454 ( \19492 , \18046 );
buf \U$13455 ( \19493 , \18046 );
buf \U$13456 ( \19494 , \18046 );
buf \U$13457 ( \19495 , \18046 );
buf \U$13458 ( \19496 , \18046 );
buf \U$13459 ( \19497 , \18046 );
buf \U$13460 ( \19498 , \18046 );
nor \U$13461 ( \19499 , \18074 , \18075 , \18076 , \18036 , \18039 , \18043 , \18046 , \19474 , \19475 , \19476 , \19477 , \19478 , \19479 , \19480 , \19481 , \19482 , \19483 , \19484 , \19485 , \19486 , \19487 , \19488 , \19489 , \19490 , \19491 , \19492 , \19493 , \19494 , \19495 , \19496 , \19497 , \19498 );
and \U$13462 ( \19500 , \8841 , \19499 );
buf \U$13463 ( \19501 , \18046 );
buf \U$13464 ( \19502 , \18046 );
buf \U$13465 ( \19503 , \18046 );
buf \U$13466 ( \19504 , \18046 );
buf \U$13467 ( \19505 , \18046 );
buf \U$13468 ( \19506 , \18046 );
buf \U$13469 ( \19507 , \18046 );
buf \U$13470 ( \19508 , \18046 );
buf \U$13471 ( \19509 , \18046 );
buf \U$13472 ( \19510 , \18046 );
buf \U$13473 ( \19511 , \18046 );
buf \U$13474 ( \19512 , \18046 );
buf \U$13475 ( \19513 , \18046 );
buf \U$13476 ( \19514 , \18046 );
buf \U$13477 ( \19515 , \18046 );
buf \U$13478 ( \19516 , \18046 );
buf \U$13479 ( \19517 , \18046 );
buf \U$13480 ( \19518 , \18046 );
buf \U$13481 ( \19519 , \18046 );
buf \U$13482 ( \19520 , \18046 );
buf \U$13483 ( \19521 , \18046 );
buf \U$13484 ( \19522 , \18046 );
buf \U$13485 ( \19523 , \18046 );
buf \U$13486 ( \19524 , \18046 );
buf \U$13487 ( \19525 , \18046 );
nor \U$13488 ( \19526 , \18033 , \18075 , \18076 , \18036 , \18039 , \18043 , \18046 , \19501 , \19502 , \19503 , \19504 , \19505 , \19506 , \19507 , \19508 , \19509 , \19510 , \19511 , \19512 , \19513 , \19514 , \19515 , \19516 , \19517 , \19518 , \19519 , \19520 , \19521 , \19522 , \19523 , \19524 , \19525 );
and \U$13489 ( \19527 , \8869 , \19526 );
buf \U$13490 ( \19528 , \18046 );
buf \U$13491 ( \19529 , \18046 );
buf \U$13492 ( \19530 , \18046 );
buf \U$13493 ( \19531 , \18046 );
buf \U$13494 ( \19532 , \18046 );
buf \U$13495 ( \19533 , \18046 );
buf \U$13496 ( \19534 , \18046 );
buf \U$13497 ( \19535 , \18046 );
buf \U$13498 ( \19536 , \18046 );
buf \U$13499 ( \19537 , \18046 );
buf \U$13500 ( \19538 , \18046 );
buf \U$13501 ( \19539 , \18046 );
buf \U$13502 ( \19540 , \18046 );
buf \U$13503 ( \19541 , \18046 );
buf \U$13504 ( \19542 , \18046 );
buf \U$13505 ( \19543 , \18046 );
buf \U$13506 ( \19544 , \18046 );
buf \U$13507 ( \19545 , \18046 );
buf \U$13508 ( \19546 , \18046 );
buf \U$13509 ( \19547 , \18046 );
buf \U$13510 ( \19548 , \18046 );
buf \U$13511 ( \19549 , \18046 );
buf \U$13512 ( \19550 , \18046 );
buf \U$13513 ( \19551 , \18046 );
buf \U$13514 ( \19552 , \18046 );
nor \U$13515 ( \19553 , \18074 , \18034 , \18076 , \18036 , \18039 , \18043 , \18046 , \19528 , \19529 , \19530 , \19531 , \19532 , \19533 , \19534 , \19535 , \19536 , \19537 , \19538 , \19539 , \19540 , \19541 , \19542 , \19543 , \19544 , \19545 , \19546 , \19547 , \19548 , \19549 , \19550 , \19551 , \19552 );
and \U$13516 ( \19554 , \8897 , \19553 );
buf \U$13517 ( \19555 , \18046 );
buf \U$13518 ( \19556 , \18046 );
buf \U$13519 ( \19557 , \18046 );
buf \U$13520 ( \19558 , \18046 );
buf \U$13521 ( \19559 , \18046 );
buf \U$13522 ( \19560 , \18046 );
buf \U$13523 ( \19561 , \18046 );
buf \U$13524 ( \19562 , \18046 );
buf \U$13525 ( \19563 , \18046 );
buf \U$13526 ( \19564 , \18046 );
buf \U$13527 ( \19565 , \18046 );
buf \U$13528 ( \19566 , \18046 );
buf \U$13529 ( \19567 , \18046 );
buf \U$13530 ( \19568 , \18046 );
buf \U$13531 ( \19569 , \18046 );
buf \U$13532 ( \19570 , \18046 );
buf \U$13533 ( \19571 , \18046 );
buf \U$13534 ( \19572 , \18046 );
buf \U$13535 ( \19573 , \18046 );
buf \U$13536 ( \19574 , \18046 );
buf \U$13537 ( \19575 , \18046 );
buf \U$13538 ( \19576 , \18046 );
buf \U$13539 ( \19577 , \18046 );
buf \U$13540 ( \19578 , \18046 );
buf \U$13541 ( \19579 , \18046 );
nor \U$13542 ( \19580 , \18033 , \18034 , \18076 , \18036 , \18039 , \18043 , \18046 , \19555 , \19556 , \19557 , \19558 , \19559 , \19560 , \19561 , \19562 , \19563 , \19564 , \19565 , \19566 , \19567 , \19568 , \19569 , \19570 , \19571 , \19572 , \19573 , \19574 , \19575 , \19576 , \19577 , \19578 , \19579 );
and \U$13543 ( \19581 , \8925 , \19580 );
buf \U$13544 ( \19582 , \18046 );
buf \U$13545 ( \19583 , \18046 );
buf \U$13546 ( \19584 , \18046 );
buf \U$13547 ( \19585 , \18046 );
buf \U$13548 ( \19586 , \18046 );
buf \U$13549 ( \19587 , \18046 );
buf \U$13550 ( \19588 , \18046 );
buf \U$13551 ( \19589 , \18046 );
buf \U$13552 ( \19590 , \18046 );
buf \U$13553 ( \19591 , \18046 );
buf \U$13554 ( \19592 , \18046 );
buf \U$13555 ( \19593 , \18046 );
buf \U$13556 ( \19594 , \18046 );
buf \U$13557 ( \19595 , \18046 );
buf \U$13558 ( \19596 , \18046 );
buf \U$13559 ( \19597 , \18046 );
buf \U$13560 ( \19598 , \18046 );
buf \U$13561 ( \19599 , \18046 );
buf \U$13562 ( \19600 , \18046 );
buf \U$13563 ( \19601 , \18046 );
buf \U$13564 ( \19602 , \18046 );
buf \U$13565 ( \19603 , \18046 );
buf \U$13566 ( \19604 , \18046 );
buf \U$13567 ( \19605 , \18046 );
buf \U$13568 ( \19606 , \18046 );
nor \U$13569 ( \19607 , \18074 , \18075 , \18035 , \18036 , \18039 , \18043 , \18046 , \19582 , \19583 , \19584 , \19585 , \19586 , \19587 , \19588 , \19589 , \19590 , \19591 , \19592 , \19593 , \19594 , \19595 , \19596 , \19597 , \19598 , \19599 , \19600 , \19601 , \19602 , \19603 , \19604 , \19605 , \19606 );
and \U$13570 ( \19608 , \8953 , \19607 );
buf \U$13571 ( \19609 , \18046 );
buf \U$13572 ( \19610 , \18046 );
buf \U$13573 ( \19611 , \18046 );
buf \U$13574 ( \19612 , \18046 );
buf \U$13575 ( \19613 , \18046 );
buf \U$13576 ( \19614 , \18046 );
buf \U$13577 ( \19615 , \18046 );
buf \U$13578 ( \19616 , \18046 );
buf \U$13579 ( \19617 , \18046 );
buf \U$13580 ( \19618 , \18046 );
buf \U$13581 ( \19619 , \18046 );
buf \U$13582 ( \19620 , \18046 );
buf \U$13583 ( \19621 , \18046 );
buf \U$13584 ( \19622 , \18046 );
buf \U$13585 ( \19623 , \18046 );
buf \U$13586 ( \19624 , \18046 );
buf \U$13587 ( \19625 , \18046 );
buf \U$13588 ( \19626 , \18046 );
buf \U$13589 ( \19627 , \18046 );
buf \U$13590 ( \19628 , \18046 );
buf \U$13591 ( \19629 , \18046 );
buf \U$13592 ( \19630 , \18046 );
buf \U$13593 ( \19631 , \18046 );
buf \U$13594 ( \19632 , \18046 );
buf \U$13595 ( \19633 , \18046 );
nor \U$13596 ( \19634 , \18033 , \18075 , \18035 , \18036 , \18039 , \18043 , \18046 , \19609 , \19610 , \19611 , \19612 , \19613 , \19614 , \19615 , \19616 , \19617 , \19618 , \19619 , \19620 , \19621 , \19622 , \19623 , \19624 , \19625 , \19626 , \19627 , \19628 , \19629 , \19630 , \19631 , \19632 , \19633 );
and \U$13597 ( \19635 , \8981 , \19634 );
buf \U$13598 ( \19636 , \18046 );
buf \U$13599 ( \19637 , \18046 );
buf \U$13600 ( \19638 , \18046 );
buf \U$13601 ( \19639 , \18046 );
buf \U$13602 ( \19640 , \18046 );
buf \U$13603 ( \19641 , \18046 );
buf \U$13604 ( \19642 , \18046 );
buf \U$13605 ( \19643 , \18046 );
buf \U$13606 ( \19644 , \18046 );
buf \U$13607 ( \19645 , \18046 );
buf \U$13608 ( \19646 , \18046 );
buf \U$13609 ( \19647 , \18046 );
buf \U$13610 ( \19648 , \18046 );
buf \U$13611 ( \19649 , \18046 );
buf \U$13612 ( \19650 , \18046 );
buf \U$13613 ( \19651 , \18046 );
buf \U$13614 ( \19652 , \18046 );
buf \U$13615 ( \19653 , \18046 );
buf \U$13616 ( \19654 , \18046 );
buf \U$13617 ( \19655 , \18046 );
buf \U$13618 ( \19656 , \18046 );
buf \U$13619 ( \19657 , \18046 );
buf \U$13620 ( \19658 , \18046 );
buf \U$13621 ( \19659 , \18046 );
buf \U$13622 ( \19660 , \18046 );
nor \U$13623 ( \19661 , \18074 , \18034 , \18035 , \18036 , \18039 , \18043 , \18046 , \19636 , \19637 , \19638 , \19639 , \19640 , \19641 , \19642 , \19643 , \19644 , \19645 , \19646 , \19647 , \19648 , \19649 , \19650 , \19651 , \19652 , \19653 , \19654 , \19655 , \19656 , \19657 , \19658 , \19659 , \19660 );
and \U$13624 ( \19662 , \9009 , \19661 );
or \U$13625 ( \19663 , \19257 , \19284 , \19311 , \19338 , \19365 , \19392 , \19419 , \19446 , \19473 , \19500 , \19527 , \19554 , \19581 , \19608 , \19635 , \19662 );
buf \U$13626 ( \19664 , \18046 );
not \U$13627 ( \19665 , \19664 );
buf \U$13628 ( \19666 , \18034 );
buf \U$13629 ( \19667 , \18035 );
buf \U$13630 ( \19668 , \18036 );
buf \U$13631 ( \19669 , \18039 );
buf \U$13632 ( \19670 , \18043 );
buf \U$13633 ( \19671 , \18046 );
buf \U$13634 ( \19672 , \18046 );
buf \U$13635 ( \19673 , \18046 );
buf \U$13636 ( \19674 , \18046 );
buf \U$13637 ( \19675 , \18046 );
buf \U$13638 ( \19676 , \18046 );
buf \U$13639 ( \19677 , \18046 );
buf \U$13640 ( \19678 , \18046 );
buf \U$13641 ( \19679 , \18046 );
buf \U$13642 ( \19680 , \18046 );
buf \U$13643 ( \19681 , \18046 );
buf \U$13644 ( \19682 , \18046 );
buf \U$13645 ( \19683 , \18046 );
buf \U$13646 ( \19684 , \18046 );
buf \U$13647 ( \19685 , \18046 );
buf \U$13648 ( \19686 , \18046 );
buf \U$13649 ( \19687 , \18046 );
buf \U$13650 ( \19688 , \18046 );
buf \U$13651 ( \19689 , \18046 );
buf \U$13652 ( \19690 , \18046 );
buf \U$13653 ( \19691 , \18046 );
buf \U$13654 ( \19692 , \18046 );
buf \U$13655 ( \19693 , \18046 );
buf \U$13656 ( \19694 , \18046 );
buf \U$13657 ( \19695 , \18046 );
buf \U$13658 ( \19696 , \18033 );
or \U$13659 ( \19697 , \19666 , \19667 , \19668 , \19669 , \19670 , \19671 , \19672 , \19673 , \19674 , \19675 , \19676 , \19677 , \19678 , \19679 , \19680 , \19681 , \19682 , \19683 , \19684 , \19685 , \19686 , \19687 , \19688 , \19689 , \19690 , \19691 , \19692 , \19693 , \19694 , \19695 , \19696 );
nand \U$13660 ( \19698 , \19665 , \19697 );
buf \U$13661 ( \19699 , \19698 );
buf \U$13662 ( \19700 , \18046 );
not \U$13663 ( \19701 , \19700 );
buf \U$13664 ( \19702 , \18043 );
buf \U$13665 ( \19703 , \18046 );
buf \U$13666 ( \19704 , \18046 );
buf \U$13667 ( \19705 , \18046 );
buf \U$13668 ( \19706 , \18046 );
buf \U$13669 ( \19707 , \18046 );
buf \U$13670 ( \19708 , \18046 );
buf \U$13671 ( \19709 , \18046 );
buf \U$13672 ( \19710 , \18046 );
buf \U$13673 ( \19711 , \18046 );
buf \U$13674 ( \19712 , \18046 );
buf \U$13675 ( \19713 , \18046 );
buf \U$13676 ( \19714 , \18046 );
buf \U$13677 ( \19715 , \18046 );
buf \U$13678 ( \19716 , \18046 );
buf \U$13679 ( \19717 , \18046 );
buf \U$13680 ( \19718 , \18046 );
buf \U$13681 ( \19719 , \18046 );
buf \U$13682 ( \19720 , \18046 );
buf \U$13683 ( \19721 , \18046 );
buf \U$13684 ( \19722 , \18046 );
buf \U$13685 ( \19723 , \18046 );
buf \U$13686 ( \19724 , \18046 );
buf \U$13687 ( \19725 , \18046 );
buf \U$13688 ( \19726 , \18046 );
buf \U$13689 ( \19727 , \18046 );
buf \U$13690 ( \19728 , \18039 );
buf \U$13691 ( \19729 , \18033 );
buf \U$13692 ( \19730 , \18034 );
buf \U$13693 ( \19731 , \18035 );
buf \U$13694 ( \19732 , \18036 );
or \U$13695 ( \19733 , \19729 , \19730 , \19731 , \19732 );
and \U$13696 ( \19734 , \19728 , \19733 );
or \U$13697 ( \19735 , \19702 , \19703 , \19704 , \19705 , \19706 , \19707 , \19708 , \19709 , \19710 , \19711 , \19712 , \19713 , \19714 , \19715 , \19716 , \19717 , \19718 , \19719 , \19720 , \19721 , \19722 , \19723 , \19724 , \19725 , \19726 , \19727 , \19734 );
and \U$13698 ( \19736 , \19701 , \19735 );
buf \U$13699 ( \19737 , \19736 );
or \U$13700 ( \19738 , \19699 , \19737 );
_DC g63f8 ( \19739_nG63f8 , \19663 , \19738 );
buf \U$13701 ( \19740 , \19739_nG63f8 );
xor \U$13702 ( \19741 , \19230 , \19740 );
buf \U$13703 ( \19742 , RIb7af5b8_255);
and \U$13704 ( \19743 , \7207 , \19256 );
and \U$13705 ( \19744 , \7209 , \19283 );
and \U$13706 ( \19745 , \9119 , \19310 );
and \U$13707 ( \19746 , \9121 , \19337 );
and \U$13708 ( \19747 , \9123 , \19364 );
and \U$13709 ( \19748 , \9125 , \19391 );
and \U$13710 ( \19749 , \9127 , \19418 );
and \U$13711 ( \19750 , \9129 , \19445 );
and \U$13712 ( \19751 , \9131 , \19472 );
and \U$13713 ( \19752 , \9133 , \19499 );
and \U$13714 ( \19753 , \9135 , \19526 );
and \U$13715 ( \19754 , \9137 , \19553 );
and \U$13716 ( \19755 , \9139 , \19580 );
and \U$13717 ( \19756 , \9141 , \19607 );
and \U$13718 ( \19757 , \9143 , \19634 );
and \U$13719 ( \19758 , \9145 , \19661 );
or \U$13720 ( \19759 , \19743 , \19744 , \19745 , \19746 , \19747 , \19748 , \19749 , \19750 , \19751 , \19752 , \19753 , \19754 , \19755 , \19756 , \19757 , \19758 );
_DC g640d ( \19760_nG640d , \19759 , \19738 );
buf \U$13721 ( \19761 , \19760_nG640d );
xor \U$13722 ( \19762 , \19742 , \19761 );
or \U$13723 ( \19763 , \19741 , \19762 );
buf \U$13724 ( \19764 , RIb7af540_256);
and \U$13725 ( \19765 , \7217 , \19256 );
and \U$13726 ( \19766 , \7219 , \19283 );
and \U$13727 ( \19767 , \9155 , \19310 );
and \U$13728 ( \19768 , \9157 , \19337 );
and \U$13729 ( \19769 , \9159 , \19364 );
and \U$13730 ( \19770 , \9161 , \19391 );
and \U$13731 ( \19771 , \9163 , \19418 );
and \U$13732 ( \19772 , \9165 , \19445 );
and \U$13733 ( \19773 , \9167 , \19472 );
and \U$13734 ( \19774 , \9169 , \19499 );
and \U$13735 ( \19775 , \9171 , \19526 );
and \U$13736 ( \19776 , \9173 , \19553 );
and \U$13737 ( \19777 , \9175 , \19580 );
and \U$13738 ( \19778 , \9177 , \19607 );
and \U$13739 ( \19779 , \9179 , \19634 );
and \U$13740 ( \19780 , \9181 , \19661 );
or \U$13741 ( \19781 , \19765 , \19766 , \19767 , \19768 , \19769 , \19770 , \19771 , \19772 , \19773 , \19774 , \19775 , \19776 , \19777 , \19778 , \19779 , \19780 );
_DC g6423 ( \19782_nG6423 , \19781 , \19738 );
buf \U$13742 ( \19783 , \19782_nG6423 );
xor \U$13743 ( \19784 , \19764 , \19783 );
or \U$13744 ( \19785 , \19763 , \19784 );
buf \U$13745 ( \19786 , RIb7af4c8_257);
and \U$13746 ( \19787 , \7227 , \19256 );
and \U$13747 ( \19788 , \7229 , \19283 );
and \U$13748 ( \19789 , \9191 , \19310 );
and \U$13749 ( \19790 , \9193 , \19337 );
and \U$13750 ( \19791 , \9195 , \19364 );
and \U$13751 ( \19792 , \9197 , \19391 );
and \U$13752 ( \19793 , \9199 , \19418 );
and \U$13753 ( \19794 , \9201 , \19445 );
and \U$13754 ( \19795 , \9203 , \19472 );
and \U$13755 ( \19796 , \9205 , \19499 );
and \U$13756 ( \19797 , \9207 , \19526 );
and \U$13757 ( \19798 , \9209 , \19553 );
and \U$13758 ( \19799 , \9211 , \19580 );
and \U$13759 ( \19800 , \9213 , \19607 );
and \U$13760 ( \19801 , \9215 , \19634 );
and \U$13761 ( \19802 , \9217 , \19661 );
or \U$13762 ( \19803 , \19787 , \19788 , \19789 , \19790 , \19791 , \19792 , \19793 , \19794 , \19795 , \19796 , \19797 , \19798 , \19799 , \19800 , \19801 , \19802 );
_DC g6439 ( \19804_nG6439 , \19803 , \19738 );
buf \U$13763 ( \19805 , \19804_nG6439 );
xor \U$13764 ( \19806 , \19786 , \19805 );
or \U$13765 ( \19807 , \19785 , \19806 );
buf \U$13766 ( \19808 , RIb7af450_258);
and \U$13767 ( \19809 , \7237 , \19256 );
and \U$13768 ( \19810 , \7239 , \19283 );
and \U$13769 ( \19811 , \9227 , \19310 );
and \U$13770 ( \19812 , \9229 , \19337 );
and \U$13771 ( \19813 , \9231 , \19364 );
and \U$13772 ( \19814 , \9233 , \19391 );
and \U$13773 ( \19815 , \9235 , \19418 );
and \U$13774 ( \19816 , \9237 , \19445 );
and \U$13775 ( \19817 , \9239 , \19472 );
and \U$13776 ( \19818 , \9241 , \19499 );
and \U$13777 ( \19819 , \9243 , \19526 );
and \U$13778 ( \19820 , \9245 , \19553 );
and \U$13779 ( \19821 , \9247 , \19580 );
and \U$13780 ( \19822 , \9249 , \19607 );
and \U$13781 ( \19823 , \9251 , \19634 );
and \U$13782 ( \19824 , \9253 , \19661 );
or \U$13783 ( \19825 , \19809 , \19810 , \19811 , \19812 , \19813 , \19814 , \19815 , \19816 , \19817 , \19818 , \19819 , \19820 , \19821 , \19822 , \19823 , \19824 );
_DC g644f ( \19826_nG644f , \19825 , \19738 );
buf \U$13784 ( \19827 , \19826_nG644f );
xor \U$13785 ( \19828 , \19808 , \19827 );
or \U$13786 ( \19829 , \19807 , \19828 );
buf \U$13787 ( \19830 , RIb7af3d8_259);
and \U$13788 ( \19831 , \7247 , \19256 );
and \U$13789 ( \19832 , \7249 , \19283 );
and \U$13790 ( \19833 , \9263 , \19310 );
and \U$13791 ( \19834 , \9265 , \19337 );
and \U$13792 ( \19835 , \9267 , \19364 );
and \U$13793 ( \19836 , \9269 , \19391 );
and \U$13794 ( \19837 , \9271 , \19418 );
and \U$13795 ( \19838 , \9273 , \19445 );
and \U$13796 ( \19839 , \9275 , \19472 );
and \U$13797 ( \19840 , \9277 , \19499 );
and \U$13798 ( \19841 , \9279 , \19526 );
and \U$13799 ( \19842 , \9281 , \19553 );
and \U$13800 ( \19843 , \9283 , \19580 );
and \U$13801 ( \19844 , \9285 , \19607 );
and \U$13802 ( \19845 , \9287 , \19634 );
and \U$13803 ( \19846 , \9289 , \19661 );
or \U$13804 ( \19847 , \19831 , \19832 , \19833 , \19834 , \19835 , \19836 , \19837 , \19838 , \19839 , \19840 , \19841 , \19842 , \19843 , \19844 , \19845 , \19846 );
_DC g6465 ( \19848_nG6465 , \19847 , \19738 );
buf \U$13805 ( \19849 , \19848_nG6465 );
xor \U$13806 ( \19850 , \19830 , \19849 );
or \U$13807 ( \19851 , \19829 , \19850 );
buf \U$13808 ( \19852 , RIb7a5bf8_260);
and \U$13809 ( \19853 , \7257 , \19256 );
and \U$13810 ( \19854 , \7259 , \19283 );
and \U$13811 ( \19855 , \9299 , \19310 );
and \U$13812 ( \19856 , \9301 , \19337 );
and \U$13813 ( \19857 , \9303 , \19364 );
and \U$13814 ( \19858 , \9305 , \19391 );
and \U$13815 ( \19859 , \9307 , \19418 );
and \U$13816 ( \19860 , \9309 , \19445 );
and \U$13817 ( \19861 , \9311 , \19472 );
and \U$13818 ( \19862 , \9313 , \19499 );
and \U$13819 ( \19863 , \9315 , \19526 );
and \U$13820 ( \19864 , \9317 , \19553 );
and \U$13821 ( \19865 , \9319 , \19580 );
and \U$13822 ( \19866 , \9321 , \19607 );
and \U$13823 ( \19867 , \9323 , \19634 );
and \U$13824 ( \19868 , \9325 , \19661 );
or \U$13825 ( \19869 , \19853 , \19854 , \19855 , \19856 , \19857 , \19858 , \19859 , \19860 , \19861 , \19862 , \19863 , \19864 , \19865 , \19866 , \19867 , \19868 );
_DC g647b ( \19870_nG647b , \19869 , \19738 );
buf \U$13826 ( \19871 , \19870_nG647b );
xor \U$13827 ( \19872 , \19852 , \19871 );
or \U$13828 ( \19873 , \19851 , \19872 );
buf \U$13829 ( \19874 , RIb7a0c48_261);
and \U$13830 ( \19875 , \7267 , \19256 );
and \U$13831 ( \19876 , \7269 , \19283 );
and \U$13832 ( \19877 , \9335 , \19310 );
and \U$13833 ( \19878 , \9337 , \19337 );
and \U$13834 ( \19879 , \9339 , \19364 );
and \U$13835 ( \19880 , \9341 , \19391 );
and \U$13836 ( \19881 , \9343 , \19418 );
and \U$13837 ( \19882 , \9345 , \19445 );
and \U$13838 ( \19883 , \9347 , \19472 );
and \U$13839 ( \19884 , \9349 , \19499 );
and \U$13840 ( \19885 , \9351 , \19526 );
and \U$13841 ( \19886 , \9353 , \19553 );
and \U$13842 ( \19887 , \9355 , \19580 );
and \U$13843 ( \19888 , \9357 , \19607 );
and \U$13844 ( \19889 , \9359 , \19634 );
and \U$13845 ( \19890 , \9361 , \19661 );
or \U$13846 ( \19891 , \19875 , \19876 , \19877 , \19878 , \19879 , \19880 , \19881 , \19882 , \19883 , \19884 , \19885 , \19886 , \19887 , \19888 , \19889 , \19890 );
_DC g6491 ( \19892_nG6491 , \19891 , \19738 );
buf \U$13847 ( \19893 , \19892_nG6491 );
xor \U$13848 ( \19894 , \19874 , \19893 );
or \U$13849 ( \19895 , \19873 , \19894 );
not \U$13850 ( \19896 , \19895 );
buf \U$13851 ( \19897 , \19896 );
and \U$13852 ( \19898 , \19229 , \19897 );
_HMUX g6498 ( \19899_nG6498 , \17768_nG5c3c , \18033 , \19898 );
buf \U$13853 ( \19900 , \17787 );
buf \U$13854 ( \19901 , \17784 );
buf \U$13855 ( \19902 , \17770 );
buf \U$13856 ( \19903 , \17773 );
buf \U$13857 ( \19904 , \17776 );
buf \U$13858 ( \19905 , \17780 );
or \U$13859 ( \19906 , \19902 , \19903 , \19904 , \19905 );
and \U$13860 ( \19907 , \19901 , \19906 );
or \U$13861 ( \19908 , \19900 , \19907 );
buf \U$13862 ( \19909 , \19908 );
_HMUX g64a3 ( \19910_nG64a3 , \18032_nG5d45 , \19899_nG6498 , \19909 );
buf \U$13863 ( \19911 , RIe5319e0_6884);
not \U$13864 ( \19912 , \19911 );
buf \U$13865 ( \19913 , \19912 );
buf \U$13866 ( \19914 , RIe549ef0_6842);
xor \U$13867 ( \19915 , \19914 , \19911 );
buf \U$13868 ( \19916 , \19915 );
buf \U$13869 ( \19917 , RIe549770_6843);
and \U$13870 ( \19918 , \19914 , \19911 );
xor \U$13871 ( \19919 , \19917 , \19918 );
buf \U$13872 ( \19920 , \19919 );
buf \U$13873 ( \19921 , RIe548ff0_6844);
and \U$13874 ( \19922 , \19917 , \19918 );
xnor \U$13875 ( \19923 , \19921 , \19922 );
buf \U$13876 ( \19924 , \19923 );
buf \U$13877 ( \19925 , RIea91330_6888);
or \U$13878 ( \19926 , \19921 , \19922 );
xor \U$13879 ( \19927 , \19925 , \19926 );
buf \U$13880 ( \19928 , \19927 );
not \U$13881 ( \19929 , \19928 );
and \U$13882 ( \19930 , \19925 , \19926 );
buf \U$13883 ( \19931 , \19930 );
nor \U$13884 ( \19932 , \19913 , \19916 , \19920 , \19924 , \19929 , \19931 );
and \U$13885 ( \19933 , RIe5329d0_6883, \19932 );
not \U$13886 ( \19934 , \19931 );
and \U$13887 ( \19935 , \19913 , \19916 , \19920 , \19924 , \19929 , \19934 );
and \U$13888 ( \19936 , RIeb72150_6905, \19935 );
not \U$13889 ( \19937 , \19913 );
and \U$13890 ( \19938 , \19937 , \19916 , \19920 , \19924 , \19929 , \19934 );
and \U$13891 ( \19939 , RIeab80c0_6897, \19938 );
not \U$13892 ( \19940 , \19916 );
and \U$13893 ( \19941 , \19913 , \19940 , \19920 , \19924 , \19929 , \19934 );
and \U$13894 ( \19942 , RIe5331c8_6882, \19941 );
and \U$13895 ( \19943 , \19937 , \19940 , \19920 , \19924 , \19929 , \19934 );
and \U$13896 ( \19944 , RIe5339c0_6881, \19943 );
not \U$13897 ( \19945 , \19920 );
and \U$13898 ( \19946 , \19913 , \19916 , \19945 , \19924 , \19929 , \19934 );
and \U$13899 ( \19947 , RIeab87c8_6898, \19946 );
and \U$13900 ( \19948 , \19937 , \19916 , \19945 , \19924 , \19929 , \19934 );
and \U$13901 ( \19949 , RIe5341b8_6880, \19948 );
and \U$13902 ( \19950 , \19913 , \19940 , \19945 , \19924 , \19929 , \19934 );
and \U$13903 ( \19951 , RIe5349b0_6879, \19950 );
or \U$13912 ( \19952 , \19933 , \19936 , \19939 , \19942 , \19944 , \19947 , \19949 , \19951 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
buf \U$13914 ( \19953 , \19931 );
buf \U$13915 ( \19954 , \19928 );
buf \U$13916 ( \19955 , \19913 );
buf \U$13917 ( \19956 , \19916 );
buf \U$13918 ( \19957 , \19920 );
buf \U$13919 ( \19958 , \19924 );
or \U$13920 ( \19959 , \19955 , \19956 , \19957 , \19958 );
and \U$13921 ( \19960 , \19954 , \19959 );
or \U$13922 ( \19961 , \19953 , \19960 );
buf \U$13923 ( \19962 , \19961 );
or \U$13924 ( \19963 , 1'b0 , \19962 );
_DC g64d9 ( \19964_nG64d9 , \19952 , \19963 );
not \U$13925 ( \19965 , \19964_nG64d9 );
buf \U$13926 ( \19966 , RIb7b9608_246);
and \U$13927 ( \19967 , \7117 , \19932 );
and \U$13928 ( \19968 , \7119 , \19935 );
and \U$13929 ( \19969 , \7864 , \19938 );
and \U$13930 ( \19970 , \7892 , \19941 );
and \U$13931 ( \19971 , \7920 , \19943 );
and \U$13932 ( \19972 , \7948 , \19946 );
and \U$13933 ( \19973 , \7976 , \19948 );
and \U$13934 ( \19974 , \8004 , \19950 );
or \U$13943 ( \19975 , \19967 , \19968 , \19969 , \19970 , \19971 , \19972 , \19973 , \19974 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g64e5 ( \19976_nG64e5 , \19975 , \19963 );
buf \U$13944 ( \19977 , \19976_nG64e5 );
xor \U$13945 ( \19978 , \19966 , \19977 );
buf \U$13946 ( \19979 , RIb7b9590_247);
and \U$13947 ( \19980 , \7126 , \19932 );
and \U$13948 ( \19981 , \7128 , \19935 );
and \U$13949 ( \19982 , \8338 , \19938 );
and \U$13950 ( \19983 , \8340 , \19941 );
and \U$13951 ( \19984 , \8342 , \19943 );
and \U$13952 ( \19985 , \8344 , \19946 );
and \U$13953 ( \19986 , \8346 , \19948 );
and \U$13954 ( \19987 , \8348 , \19950 );
or \U$13963 ( \19988 , \19980 , \19981 , \19982 , \19983 , \19984 , \19985 , \19986 , \19987 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g64f2 ( \19989_nG64f2 , \19988 , \19963 );
buf \U$13964 ( \19990 , \19989_nG64f2 );
xor \U$13965 ( \19991 , \19979 , \19990 );
or \U$13966 ( \19992 , \19978 , \19991 );
buf \U$13967 ( \19993 , RIb7b9518_248);
and \U$13968 ( \19994 , \7136 , \19932 );
and \U$13969 ( \19995 , \7138 , \19935 );
and \U$13970 ( \19996 , \8374 , \19938 );
and \U$13971 ( \19997 , \8376 , \19941 );
and \U$13972 ( \19998 , \8378 , \19943 );
and \U$13973 ( \19999 , \8380 , \19946 );
and \U$13974 ( \20000 , \8382 , \19948 );
and \U$13975 ( \20001 , \8384 , \19950 );
or \U$13984 ( \20002 , \19994 , \19995 , \19996 , \19997 , \19998 , \19999 , \20000 , \20001 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6500 ( \20003_nG6500 , \20002 , \19963 );
buf \U$13985 ( \20004 , \20003_nG6500 );
xor \U$13986 ( \20005 , \19993 , \20004 );
or \U$13987 ( \20006 , \19992 , \20005 );
buf \U$13988 ( \20007 , RIb7b94a0_249);
and \U$13989 ( \20008 , \7146 , \19932 );
and \U$13990 ( \20009 , \7148 , \19935 );
and \U$13991 ( \20010 , \8410 , \19938 );
and \U$13992 ( \20011 , \8412 , \19941 );
and \U$13993 ( \20012 , \8414 , \19943 );
and \U$13994 ( \20013 , \8416 , \19946 );
and \U$13995 ( \20014 , \8418 , \19948 );
and \U$13996 ( \20015 , \8420 , \19950 );
or \U$14005 ( \20016 , \20008 , \20009 , \20010 , \20011 , \20012 , \20013 , \20014 , \20015 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g650e ( \20017_nG650e , \20016 , \19963 );
buf \U$14006 ( \20018 , \20017_nG650e );
xor \U$14007 ( \20019 , \20007 , \20018 );
or \U$14008 ( \20020 , \20006 , \20019 );
buf \U$14009 ( \20021 , RIb7b9428_250);
and \U$14010 ( \20022 , \7156 , \19932 );
and \U$14011 ( \20023 , \7158 , \19935 );
and \U$14012 ( \20024 , \8446 , \19938 );
and \U$14013 ( \20025 , \8448 , \19941 );
and \U$14014 ( \20026 , \8450 , \19943 );
and \U$14015 ( \20027 , \8452 , \19946 );
and \U$14016 ( \20028 , \8454 , \19948 );
and \U$14017 ( \20029 , \8456 , \19950 );
or \U$14026 ( \20030 , \20022 , \20023 , \20024 , \20025 , \20026 , \20027 , \20028 , \20029 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g651c ( \20031_nG651c , \20030 , \19963 );
buf \U$14027 ( \20032 , \20031_nG651c );
xor \U$14028 ( \20033 , \20021 , \20032 );
or \U$14029 ( \20034 , \20020 , \20033 );
buf \U$14030 ( \20035 , RIb7b93b0_251);
and \U$14031 ( \20036 , \7166 , \19932 );
and \U$14032 ( \20037 , \7168 , \19935 );
and \U$14033 ( \20038 , \8482 , \19938 );
and \U$14034 ( \20039 , \8484 , \19941 );
and \U$14035 ( \20040 , \8486 , \19943 );
and \U$14036 ( \20041 , \8488 , \19946 );
and \U$14037 ( \20042 , \8490 , \19948 );
and \U$14038 ( \20043 , \8492 , \19950 );
or \U$14047 ( \20044 , \20036 , \20037 , \20038 , \20039 , \20040 , \20041 , \20042 , \20043 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g652a ( \20045_nG652a , \20044 , \19963 );
buf \U$14048 ( \20046 , \20045_nG652a );
xor \U$14049 ( \20047 , \20035 , \20046 );
or \U$14050 ( \20048 , \20034 , \20047 );
buf \U$14051 ( \20049 , RIb7af720_252);
and \U$14052 ( \20050 , \7176 , \19932 );
and \U$14053 ( \20051 , \7178 , \19935 );
and \U$14054 ( \20052 , \8518 , \19938 );
and \U$14055 ( \20053 , \8520 , \19941 );
and \U$14056 ( \20054 , \8522 , \19943 );
and \U$14057 ( \20055 , \8524 , \19946 );
and \U$14058 ( \20056 , \8526 , \19948 );
and \U$14059 ( \20057 , \8528 , \19950 );
or \U$14068 ( \20058 , \20050 , \20051 , \20052 , \20053 , \20054 , \20055 , \20056 , \20057 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6538 ( \20059_nG6538 , \20058 , \19963 );
buf \U$14069 ( \20060 , \20059_nG6538 );
xor \U$14070 ( \20061 , \20049 , \20060 );
or \U$14071 ( \20062 , \20048 , \20061 );
buf \U$14072 ( \20063 , RIb7af6a8_253);
and \U$14073 ( \20064 , \7186 , \19932 );
and \U$14074 ( \20065 , \7188 , \19935 );
and \U$14075 ( \20066 , \8554 , \19938 );
and \U$14076 ( \20067 , \8556 , \19941 );
and \U$14077 ( \20068 , \8558 , \19943 );
and \U$14078 ( \20069 , \8560 , \19946 );
and \U$14079 ( \20070 , \8562 , \19948 );
and \U$14080 ( \20071 , \8564 , \19950 );
or \U$14089 ( \20072 , \20064 , \20065 , \20066 , \20067 , \20068 , \20069 , \20070 , \20071 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6546 ( \20073_nG6546 , \20072 , \19963 );
buf \U$14090 ( \20074 , \20073_nG6546 );
xor \U$14091 ( \20075 , \20063 , \20074 );
or \U$14092 ( \20076 , \20062 , \20075 );
not \U$14093 ( \20077 , \20076 );
buf \U$14094 ( \20078 , \20077 );
buf \U$14095 ( \20079 , RIb7af630_254);
and \U$14096 ( \20080 , \7198 , \19932 );
and \U$14097 ( \20081 , \7200 , \19935 );
and \U$14098 ( \20082 , \8645 , \19938 );
and \U$14099 ( \20083 , \8673 , \19941 );
and \U$14100 ( \20084 , \8701 , \19943 );
and \U$14101 ( \20085 , \8729 , \19946 );
and \U$14102 ( \20086 , \8757 , \19948 );
and \U$14103 ( \20087 , \8785 , \19950 );
or \U$14112 ( \20088 , \20080 , \20081 , \20082 , \20083 , \20084 , \20085 , \20086 , \20087 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6556 ( \20089_nG6556 , \20088 , \19963 );
buf \U$14113 ( \20090 , \20089_nG6556 );
xor \U$14114 ( \20091 , \20079 , \20090 );
buf \U$14115 ( \20092 , RIb7af5b8_255);
and \U$14116 ( \20093 , \7207 , \19932 );
and \U$14117 ( \20094 , \7209 , \19935 );
and \U$14118 ( \20095 , \9119 , \19938 );
and \U$14119 ( \20096 , \9121 , \19941 );
and \U$14120 ( \20097 , \9123 , \19943 );
and \U$14121 ( \20098 , \9125 , \19946 );
and \U$14122 ( \20099 , \9127 , \19948 );
and \U$14123 ( \20100 , \9129 , \19950 );
or \U$14132 ( \20101 , \20093 , \20094 , \20095 , \20096 , \20097 , \20098 , \20099 , \20100 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6563 ( \20102_nG6563 , \20101 , \19963 );
buf \U$14133 ( \20103 , \20102_nG6563 );
xor \U$14134 ( \20104 , \20092 , \20103 );
or \U$14135 ( \20105 , \20091 , \20104 );
buf \U$14136 ( \20106 , RIb7af540_256);
and \U$14137 ( \20107 , \7217 , \19932 );
and \U$14138 ( \20108 , \7219 , \19935 );
and \U$14139 ( \20109 , \9155 , \19938 );
and \U$14140 ( \20110 , \9157 , \19941 );
and \U$14141 ( \20111 , \9159 , \19943 );
and \U$14142 ( \20112 , \9161 , \19946 );
and \U$14143 ( \20113 , \9163 , \19948 );
and \U$14144 ( \20114 , \9165 , \19950 );
or \U$14153 ( \20115 , \20107 , \20108 , \20109 , \20110 , \20111 , \20112 , \20113 , \20114 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6571 ( \20116_nG6571 , \20115 , \19963 );
buf \U$14154 ( \20117 , \20116_nG6571 );
xor \U$14155 ( \20118 , \20106 , \20117 );
or \U$14156 ( \20119 , \20105 , \20118 );
buf \U$14157 ( \20120 , RIb7af4c8_257);
and \U$14158 ( \20121 , \7227 , \19932 );
and \U$14159 ( \20122 , \7229 , \19935 );
and \U$14160 ( \20123 , \9191 , \19938 );
and \U$14161 ( \20124 , \9193 , \19941 );
and \U$14162 ( \20125 , \9195 , \19943 );
and \U$14163 ( \20126 , \9197 , \19946 );
and \U$14164 ( \20127 , \9199 , \19948 );
and \U$14165 ( \20128 , \9201 , \19950 );
or \U$14174 ( \20129 , \20121 , \20122 , \20123 , \20124 , \20125 , \20126 , \20127 , \20128 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g657f ( \20130_nG657f , \20129 , \19963 );
buf \U$14175 ( \20131 , \20130_nG657f );
xor \U$14176 ( \20132 , \20120 , \20131 );
or \U$14177 ( \20133 , \20119 , \20132 );
buf \U$14178 ( \20134 , RIb7af450_258);
and \U$14179 ( \20135 , \7237 , \19932 );
and \U$14180 ( \20136 , \7239 , \19935 );
and \U$14181 ( \20137 , \9227 , \19938 );
and \U$14182 ( \20138 , \9229 , \19941 );
and \U$14183 ( \20139 , \9231 , \19943 );
and \U$14184 ( \20140 , \9233 , \19946 );
and \U$14185 ( \20141 , \9235 , \19948 );
and \U$14186 ( \20142 , \9237 , \19950 );
or \U$14195 ( \20143 , \20135 , \20136 , \20137 , \20138 , \20139 , \20140 , \20141 , \20142 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g658d ( \20144_nG658d , \20143 , \19963 );
buf \U$14196 ( \20145 , \20144_nG658d );
xor \U$14197 ( \20146 , \20134 , \20145 );
or \U$14198 ( \20147 , \20133 , \20146 );
buf \U$14199 ( \20148 , RIb7af3d8_259);
and \U$14200 ( \20149 , \7247 , \19932 );
and \U$14201 ( \20150 , \7249 , \19935 );
and \U$14202 ( \20151 , \9263 , \19938 );
and \U$14203 ( \20152 , \9265 , \19941 );
and \U$14204 ( \20153 , \9267 , \19943 );
and \U$14205 ( \20154 , \9269 , \19946 );
and \U$14206 ( \20155 , \9271 , \19948 );
and \U$14207 ( \20156 , \9273 , \19950 );
or \U$14216 ( \20157 , \20149 , \20150 , \20151 , \20152 , \20153 , \20154 , \20155 , \20156 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g659b ( \20158_nG659b , \20157 , \19963 );
buf \U$14217 ( \20159 , \20158_nG659b );
xor \U$14218 ( \20160 , \20148 , \20159 );
or \U$14219 ( \20161 , \20147 , \20160 );
buf \U$14220 ( \20162 , RIb7a5bf8_260);
and \U$14221 ( \20163 , \7257 , \19932 );
and \U$14222 ( \20164 , \7259 , \19935 );
and \U$14223 ( \20165 , \9299 , \19938 );
and \U$14224 ( \20166 , \9301 , \19941 );
and \U$14225 ( \20167 , \9303 , \19943 );
and \U$14226 ( \20168 , \9305 , \19946 );
and \U$14227 ( \20169 , \9307 , \19948 );
and \U$14228 ( \20170 , \9309 , \19950 );
or \U$14237 ( \20171 , \20163 , \20164 , \20165 , \20166 , \20167 , \20168 , \20169 , \20170 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g65a9 ( \20172_nG65a9 , \20171 , \19963 );
buf \U$14238 ( \20173 , \20172_nG65a9 );
xor \U$14239 ( \20174 , \20162 , \20173 );
or \U$14240 ( \20175 , \20161 , \20174 );
buf \U$14241 ( \20176 , RIb7a0c48_261);
and \U$14242 ( \20177 , \7267 , \19932 );
and \U$14243 ( \20178 , \7269 , \19935 );
and \U$14244 ( \20179 , \9335 , \19938 );
and \U$14245 ( \20180 , \9337 , \19941 );
and \U$14246 ( \20181 , \9339 , \19943 );
and \U$14247 ( \20182 , \9341 , \19946 );
and \U$14248 ( \20183 , \9343 , \19948 );
and \U$14249 ( \20184 , \9345 , \19950 );
or \U$14258 ( \20185 , \20177 , \20178 , \20179 , \20180 , \20181 , \20182 , \20183 , \20184 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g65b7 ( \20186_nG65b7 , \20185 , \19963 );
buf \U$14259 ( \20187 , \20186_nG65b7 );
xor \U$14260 ( \20188 , \20176 , \20187 );
or \U$14261 ( \20189 , \20175 , \20188 );
not \U$14262 ( \20190 , \20189 );
buf \U$14263 ( \20191 , \20190 );
and \U$14264 ( \20192 , \20078 , \20191 );
and \U$14265 ( \20193 , \19965 , \20192 );
_HMUX g65bf ( \20194_nG65bf , \19910_nG64a3 , \19913 , \20193 );
buf \U$14268 ( \20195 , \19913 );
buf \U$14271 ( \20196 , \19916 );
buf \U$14274 ( \20197 , \19920 );
buf \U$14277 ( \20198 , \19924 );
buf \U$14278 ( \20199 , \19928 );
not \U$14279 ( \20200 , \20199 );
buf \U$14280 ( \20201 , \20200 );
not \U$14281 ( \20202 , \20201 );
buf \U$14282 ( \20203 , \19931 );
xnor \U$14283 ( \20204 , \20203 , \20199 );
buf \U$14284 ( \20205 , \20204 );
or \U$14285 ( \20206 , \20203 , \20199 );
not \U$14286 ( \20207 , \20206 );
buf \U$14287 ( \20208 , \20207 );
buf \U$14288 ( \20209 , \20208 );
buf \U$14289 ( \20210 , \20208 );
buf \U$14290 ( \20211 , \20208 );
buf \U$14291 ( \20212 , \20208 );
buf \U$14292 ( \20213 , \20208 );
buf \U$14293 ( \20214 , \20208 );
buf \U$14294 ( \20215 , \20208 );
buf \U$14295 ( \20216 , \20208 );
buf \U$14296 ( \20217 , \20208 );
buf \U$14297 ( \20218 , \20208 );
buf \U$14298 ( \20219 , \20208 );
buf \U$14299 ( \20220 , \20208 );
buf \U$14300 ( \20221 , \20208 );
buf \U$14301 ( \20222 , \20208 );
buf \U$14302 ( \20223 , \20208 );
buf \U$14303 ( \20224 , \20208 );
buf \U$14304 ( \20225 , \20208 );
buf \U$14305 ( \20226 , \20208 );
buf \U$14306 ( \20227 , \20208 );
buf \U$14307 ( \20228 , \20208 );
buf \U$14308 ( \20229 , \20208 );
buf \U$14309 ( \20230 , \20208 );
buf \U$14310 ( \20231 , \20208 );
buf \U$14311 ( \20232 , \20208 );
buf \U$14312 ( \20233 , \20208 );
nor \U$14313 ( \20234 , \20195 , \20196 , \20197 , \20198 , \20202 , \20205 , \20208 , \20209 , \20210 , \20211 , \20212 , \20213 , \20214 , \20215 , \20216 , \20217 , \20218 , \20219 , \20220 , \20221 , \20222 , \20223 , \20224 , \20225 , \20226 , \20227 , \20228 , \20229 , \20230 , \20231 , \20232 , \20233 );
and \U$14314 ( \20235 , RIe5329d0_6883, \20234 );
not \U$14315 ( \20236 , \20195 );
not \U$14316 ( \20237 , \20196 );
not \U$14317 ( \20238 , \20197 );
not \U$14318 ( \20239 , \20198 );
buf \U$14319 ( \20240 , \20208 );
buf \U$14320 ( \20241 , \20208 );
buf \U$14321 ( \20242 , \20208 );
buf \U$14322 ( \20243 , \20208 );
buf \U$14323 ( \20244 , \20208 );
buf \U$14324 ( \20245 , \20208 );
buf \U$14325 ( \20246 , \20208 );
buf \U$14326 ( \20247 , \20208 );
buf \U$14327 ( \20248 , \20208 );
buf \U$14328 ( \20249 , \20208 );
buf \U$14329 ( \20250 , \20208 );
buf \U$14330 ( \20251 , \20208 );
buf \U$14331 ( \20252 , \20208 );
buf \U$14332 ( \20253 , \20208 );
buf \U$14333 ( \20254 , \20208 );
buf \U$14334 ( \20255 , \20208 );
buf \U$14335 ( \20256 , \20208 );
buf \U$14336 ( \20257 , \20208 );
buf \U$14337 ( \20258 , \20208 );
buf \U$14338 ( \20259 , \20208 );
buf \U$14339 ( \20260 , \20208 );
buf \U$14340 ( \20261 , \20208 );
buf \U$14341 ( \20262 , \20208 );
buf \U$14342 ( \20263 , \20208 );
buf \U$14343 ( \20264 , \20208 );
nor \U$14344 ( \20265 , \20236 , \20237 , \20238 , \20239 , \20201 , \20205 , \20208 , \20240 , \20241 , \20242 , \20243 , \20244 , \20245 , \20246 , \20247 , \20248 , \20249 , \20250 , \20251 , \20252 , \20253 , \20254 , \20255 , \20256 , \20257 , \20258 , \20259 , \20260 , \20261 , \20262 , \20263 , \20264 );
and \U$14345 ( \20266 , RIeb72150_6905, \20265 );
buf \U$14346 ( \20267 , \20208 );
buf \U$14347 ( \20268 , \20208 );
buf \U$14348 ( \20269 , \20208 );
buf \U$14349 ( \20270 , \20208 );
buf \U$14350 ( \20271 , \20208 );
buf \U$14351 ( \20272 , \20208 );
buf \U$14352 ( \20273 , \20208 );
buf \U$14353 ( \20274 , \20208 );
buf \U$14354 ( \20275 , \20208 );
buf \U$14355 ( \20276 , \20208 );
buf \U$14356 ( \20277 , \20208 );
buf \U$14357 ( \20278 , \20208 );
buf \U$14358 ( \20279 , \20208 );
buf \U$14359 ( \20280 , \20208 );
buf \U$14360 ( \20281 , \20208 );
buf \U$14361 ( \20282 , \20208 );
buf \U$14362 ( \20283 , \20208 );
buf \U$14363 ( \20284 , \20208 );
buf \U$14364 ( \20285 , \20208 );
buf \U$14365 ( \20286 , \20208 );
buf \U$14366 ( \20287 , \20208 );
buf \U$14367 ( \20288 , \20208 );
buf \U$14368 ( \20289 , \20208 );
buf \U$14369 ( \20290 , \20208 );
buf \U$14370 ( \20291 , \20208 );
nor \U$14371 ( \20292 , \20195 , \20237 , \20238 , \20239 , \20201 , \20205 , \20208 , \20267 , \20268 , \20269 , \20270 , \20271 , \20272 , \20273 , \20274 , \20275 , \20276 , \20277 , \20278 , \20279 , \20280 , \20281 , \20282 , \20283 , \20284 , \20285 , \20286 , \20287 , \20288 , \20289 , \20290 , \20291 );
and \U$14372 ( \20293 , RIeab80c0_6897, \20292 );
buf \U$14373 ( \20294 , \20208 );
buf \U$14374 ( \20295 , \20208 );
buf \U$14375 ( \20296 , \20208 );
buf \U$14376 ( \20297 , \20208 );
buf \U$14377 ( \20298 , \20208 );
buf \U$14378 ( \20299 , \20208 );
buf \U$14379 ( \20300 , \20208 );
buf \U$14380 ( \20301 , \20208 );
buf \U$14381 ( \20302 , \20208 );
buf \U$14382 ( \20303 , \20208 );
buf \U$14383 ( \20304 , \20208 );
buf \U$14384 ( \20305 , \20208 );
buf \U$14385 ( \20306 , \20208 );
buf \U$14386 ( \20307 , \20208 );
buf \U$14387 ( \20308 , \20208 );
buf \U$14388 ( \20309 , \20208 );
buf \U$14389 ( \20310 , \20208 );
buf \U$14390 ( \20311 , \20208 );
buf \U$14391 ( \20312 , \20208 );
buf \U$14392 ( \20313 , \20208 );
buf \U$14393 ( \20314 , \20208 );
buf \U$14394 ( \20315 , \20208 );
buf \U$14395 ( \20316 , \20208 );
buf \U$14396 ( \20317 , \20208 );
buf \U$14397 ( \20318 , \20208 );
nor \U$14398 ( \20319 , \20236 , \20196 , \20238 , \20239 , \20201 , \20205 , \20208 , \20294 , \20295 , \20296 , \20297 , \20298 , \20299 , \20300 , \20301 , \20302 , \20303 , \20304 , \20305 , \20306 , \20307 , \20308 , \20309 , \20310 , \20311 , \20312 , \20313 , \20314 , \20315 , \20316 , \20317 , \20318 );
and \U$14399 ( \20320 , RIe5331c8_6882, \20319 );
buf \U$14400 ( \20321 , \20208 );
buf \U$14401 ( \20322 , \20208 );
buf \U$14402 ( \20323 , \20208 );
buf \U$14403 ( \20324 , \20208 );
buf \U$14404 ( \20325 , \20208 );
buf \U$14405 ( \20326 , \20208 );
buf \U$14406 ( \20327 , \20208 );
buf \U$14407 ( \20328 , \20208 );
buf \U$14408 ( \20329 , \20208 );
buf \U$14409 ( \20330 , \20208 );
buf \U$14410 ( \20331 , \20208 );
buf \U$14411 ( \20332 , \20208 );
buf \U$14412 ( \20333 , \20208 );
buf \U$14413 ( \20334 , \20208 );
buf \U$14414 ( \20335 , \20208 );
buf \U$14415 ( \20336 , \20208 );
buf \U$14416 ( \20337 , \20208 );
buf \U$14417 ( \20338 , \20208 );
buf \U$14418 ( \20339 , \20208 );
buf \U$14419 ( \20340 , \20208 );
buf \U$14420 ( \20341 , \20208 );
buf \U$14421 ( \20342 , \20208 );
buf \U$14422 ( \20343 , \20208 );
buf \U$14423 ( \20344 , \20208 );
buf \U$14424 ( \20345 , \20208 );
nor \U$14425 ( \20346 , \20195 , \20196 , \20238 , \20239 , \20201 , \20205 , \20208 , \20321 , \20322 , \20323 , \20324 , \20325 , \20326 , \20327 , \20328 , \20329 , \20330 , \20331 , \20332 , \20333 , \20334 , \20335 , \20336 , \20337 , \20338 , \20339 , \20340 , \20341 , \20342 , \20343 , \20344 , \20345 );
and \U$14426 ( \20347 , RIe5339c0_6881, \20346 );
buf \U$14427 ( \20348 , \20208 );
buf \U$14428 ( \20349 , \20208 );
buf \U$14429 ( \20350 , \20208 );
buf \U$14430 ( \20351 , \20208 );
buf \U$14431 ( \20352 , \20208 );
buf \U$14432 ( \20353 , \20208 );
buf \U$14433 ( \20354 , \20208 );
buf \U$14434 ( \20355 , \20208 );
buf \U$14435 ( \20356 , \20208 );
buf \U$14436 ( \20357 , \20208 );
buf \U$14437 ( \20358 , \20208 );
buf \U$14438 ( \20359 , \20208 );
buf \U$14439 ( \20360 , \20208 );
buf \U$14440 ( \20361 , \20208 );
buf \U$14441 ( \20362 , \20208 );
buf \U$14442 ( \20363 , \20208 );
buf \U$14443 ( \20364 , \20208 );
buf \U$14444 ( \20365 , \20208 );
buf \U$14445 ( \20366 , \20208 );
buf \U$14446 ( \20367 , \20208 );
buf \U$14447 ( \20368 , \20208 );
buf \U$14448 ( \20369 , \20208 );
buf \U$14449 ( \20370 , \20208 );
buf \U$14450 ( \20371 , \20208 );
buf \U$14451 ( \20372 , \20208 );
nor \U$14452 ( \20373 , \20236 , \20237 , \20197 , \20239 , \20201 , \20205 , \20208 , \20348 , \20349 , \20350 , \20351 , \20352 , \20353 , \20354 , \20355 , \20356 , \20357 , \20358 , \20359 , \20360 , \20361 , \20362 , \20363 , \20364 , \20365 , \20366 , \20367 , \20368 , \20369 , \20370 , \20371 , \20372 );
and \U$14453 ( \20374 , RIeab87c8_6898, \20373 );
buf \U$14454 ( \20375 , \20208 );
buf \U$14455 ( \20376 , \20208 );
buf \U$14456 ( \20377 , \20208 );
buf \U$14457 ( \20378 , \20208 );
buf \U$14458 ( \20379 , \20208 );
buf \U$14459 ( \20380 , \20208 );
buf \U$14460 ( \20381 , \20208 );
buf \U$14461 ( \20382 , \20208 );
buf \U$14462 ( \20383 , \20208 );
buf \U$14463 ( \20384 , \20208 );
buf \U$14464 ( \20385 , \20208 );
buf \U$14465 ( \20386 , \20208 );
buf \U$14466 ( \20387 , \20208 );
buf \U$14467 ( \20388 , \20208 );
buf \U$14468 ( \20389 , \20208 );
buf \U$14469 ( \20390 , \20208 );
buf \U$14470 ( \20391 , \20208 );
buf \U$14471 ( \20392 , \20208 );
buf \U$14472 ( \20393 , \20208 );
buf \U$14473 ( \20394 , \20208 );
buf \U$14474 ( \20395 , \20208 );
buf \U$14475 ( \20396 , \20208 );
buf \U$14476 ( \20397 , \20208 );
buf \U$14477 ( \20398 , \20208 );
buf \U$14478 ( \20399 , \20208 );
nor \U$14479 ( \20400 , \20195 , \20237 , \20197 , \20239 , \20201 , \20205 , \20208 , \20375 , \20376 , \20377 , \20378 , \20379 , \20380 , \20381 , \20382 , \20383 , \20384 , \20385 , \20386 , \20387 , \20388 , \20389 , \20390 , \20391 , \20392 , \20393 , \20394 , \20395 , \20396 , \20397 , \20398 , \20399 );
and \U$14480 ( \20401 , RIe5341b8_6880, \20400 );
buf \U$14481 ( \20402 , \20208 );
buf \U$14482 ( \20403 , \20208 );
buf \U$14483 ( \20404 , \20208 );
buf \U$14484 ( \20405 , \20208 );
buf \U$14485 ( \20406 , \20208 );
buf \U$14486 ( \20407 , \20208 );
buf \U$14487 ( \20408 , \20208 );
buf \U$14488 ( \20409 , \20208 );
buf \U$14489 ( \20410 , \20208 );
buf \U$14490 ( \20411 , \20208 );
buf \U$14491 ( \20412 , \20208 );
buf \U$14492 ( \20413 , \20208 );
buf \U$14493 ( \20414 , \20208 );
buf \U$14494 ( \20415 , \20208 );
buf \U$14495 ( \20416 , \20208 );
buf \U$14496 ( \20417 , \20208 );
buf \U$14497 ( \20418 , \20208 );
buf \U$14498 ( \20419 , \20208 );
buf \U$14499 ( \20420 , \20208 );
buf \U$14500 ( \20421 , \20208 );
buf \U$14501 ( \20422 , \20208 );
buf \U$14502 ( \20423 , \20208 );
buf \U$14503 ( \20424 , \20208 );
buf \U$14504 ( \20425 , \20208 );
buf \U$14505 ( \20426 , \20208 );
nor \U$14506 ( \20427 , \20236 , \20196 , \20197 , \20239 , \20201 , \20205 , \20208 , \20402 , \20403 , \20404 , \20405 , \20406 , \20407 , \20408 , \20409 , \20410 , \20411 , \20412 , \20413 , \20414 , \20415 , \20416 , \20417 , \20418 , \20419 , \20420 , \20421 , \20422 , \20423 , \20424 , \20425 , \20426 );
and \U$14507 ( \20428 , RIe5349b0_6879, \20427 );
buf \U$14508 ( \20429 , \20208 );
buf \U$14509 ( \20430 , \20208 );
buf \U$14510 ( \20431 , \20208 );
buf \U$14511 ( \20432 , \20208 );
buf \U$14512 ( \20433 , \20208 );
buf \U$14513 ( \20434 , \20208 );
buf \U$14514 ( \20435 , \20208 );
buf \U$14515 ( \20436 , \20208 );
buf \U$14516 ( \20437 , \20208 );
buf \U$14517 ( \20438 , \20208 );
buf \U$14518 ( \20439 , \20208 );
buf \U$14519 ( \20440 , \20208 );
buf \U$14520 ( \20441 , \20208 );
buf \U$14521 ( \20442 , \20208 );
buf \U$14522 ( \20443 , \20208 );
buf \U$14523 ( \20444 , \20208 );
buf \U$14524 ( \20445 , \20208 );
buf \U$14525 ( \20446 , \20208 );
buf \U$14526 ( \20447 , \20208 );
buf \U$14527 ( \20448 , \20208 );
buf \U$14528 ( \20449 , \20208 );
buf \U$14529 ( \20450 , \20208 );
buf \U$14530 ( \20451 , \20208 );
buf \U$14531 ( \20452 , \20208 );
buf \U$14532 ( \20453 , \20208 );
nor \U$14533 ( \20454 , \20195 , \20196 , \20197 , \20239 , \20201 , \20205 , \20208 , \20429 , \20430 , \20431 , \20432 , \20433 , \20434 , \20435 , \20436 , \20437 , \20438 , \20439 , \20440 , \20441 , \20442 , \20443 , \20444 , \20445 , \20446 , \20447 , \20448 , \20449 , \20450 , \20451 , \20452 , \20453 );
and \U$14534 ( \20455 , RIea94af8_6890, \20454 );
buf \U$14535 ( \20456 , \20208 );
buf \U$14536 ( \20457 , \20208 );
buf \U$14537 ( \20458 , \20208 );
buf \U$14538 ( \20459 , \20208 );
buf \U$14539 ( \20460 , \20208 );
buf \U$14540 ( \20461 , \20208 );
buf \U$14541 ( \20462 , \20208 );
buf \U$14542 ( \20463 , \20208 );
buf \U$14543 ( \20464 , \20208 );
buf \U$14544 ( \20465 , \20208 );
buf \U$14545 ( \20466 , \20208 );
buf \U$14546 ( \20467 , \20208 );
buf \U$14547 ( \20468 , \20208 );
buf \U$14548 ( \20469 , \20208 );
buf \U$14549 ( \20470 , \20208 );
buf \U$14550 ( \20471 , \20208 );
buf \U$14551 ( \20472 , \20208 );
buf \U$14552 ( \20473 , \20208 );
buf \U$14553 ( \20474 , \20208 );
buf \U$14554 ( \20475 , \20208 );
buf \U$14555 ( \20476 , \20208 );
buf \U$14556 ( \20477 , \20208 );
buf \U$14557 ( \20478 , \20208 );
buf \U$14558 ( \20479 , \20208 );
buf \U$14559 ( \20480 , \20208 );
nor \U$14560 ( \20481 , \20236 , \20237 , \20238 , \20198 , \20201 , \20205 , \20208 , \20456 , \20457 , \20458 , \20459 , \20460 , \20461 , \20462 , \20463 , \20464 , \20465 , \20466 , \20467 , \20468 , \20469 , \20470 , \20471 , \20472 , \20473 , \20474 , \20475 , \20476 , \20477 , \20478 , \20479 , \20480 );
and \U$14561 ( \20482 , RIe5351a8_6878, \20481 );
buf \U$14562 ( \20483 , \20208 );
buf \U$14563 ( \20484 , \20208 );
buf \U$14564 ( \20485 , \20208 );
buf \U$14565 ( \20486 , \20208 );
buf \U$14566 ( \20487 , \20208 );
buf \U$14567 ( \20488 , \20208 );
buf \U$14568 ( \20489 , \20208 );
buf \U$14569 ( \20490 , \20208 );
buf \U$14570 ( \20491 , \20208 );
buf \U$14571 ( \20492 , \20208 );
buf \U$14572 ( \20493 , \20208 );
buf \U$14573 ( \20494 , \20208 );
buf \U$14574 ( \20495 , \20208 );
buf \U$14575 ( \20496 , \20208 );
buf \U$14576 ( \20497 , \20208 );
buf \U$14577 ( \20498 , \20208 );
buf \U$14578 ( \20499 , \20208 );
buf \U$14579 ( \20500 , \20208 );
buf \U$14580 ( \20501 , \20208 );
buf \U$14581 ( \20502 , \20208 );
buf \U$14582 ( \20503 , \20208 );
buf \U$14583 ( \20504 , \20208 );
buf \U$14584 ( \20505 , \20208 );
buf \U$14585 ( \20506 , \20208 );
buf \U$14586 ( \20507 , \20208 );
nor \U$14587 ( \20508 , \20195 , \20237 , \20238 , \20198 , \20201 , \20205 , \20208 , \20483 , \20484 , \20485 , \20486 , \20487 , \20488 , \20489 , \20490 , \20491 , \20492 , \20493 , \20494 , \20495 , \20496 , \20497 , \20498 , \20499 , \20500 , \20501 , \20502 , \20503 , \20504 , \20505 , \20506 , \20507 );
and \U$14588 ( \20509 , RIe5359a0_6877, \20508 );
buf \U$14589 ( \20510 , \20208 );
buf \U$14590 ( \20511 , \20208 );
buf \U$14591 ( \20512 , \20208 );
buf \U$14592 ( \20513 , \20208 );
buf \U$14593 ( \20514 , \20208 );
buf \U$14594 ( \20515 , \20208 );
buf \U$14595 ( \20516 , \20208 );
buf \U$14596 ( \20517 , \20208 );
buf \U$14597 ( \20518 , \20208 );
buf \U$14598 ( \20519 , \20208 );
buf \U$14599 ( \20520 , \20208 );
buf \U$14600 ( \20521 , \20208 );
buf \U$14601 ( \20522 , \20208 );
buf \U$14602 ( \20523 , \20208 );
buf \U$14603 ( \20524 , \20208 );
buf \U$14604 ( \20525 , \20208 );
buf \U$14605 ( \20526 , \20208 );
buf \U$14606 ( \20527 , \20208 );
buf \U$14607 ( \20528 , \20208 );
buf \U$14608 ( \20529 , \20208 );
buf \U$14609 ( \20530 , \20208 );
buf \U$14610 ( \20531 , \20208 );
buf \U$14611 ( \20532 , \20208 );
buf \U$14612 ( \20533 , \20208 );
buf \U$14613 ( \20534 , \20208 );
nor \U$14614 ( \20535 , \20236 , \20196 , \20238 , \20198 , \20201 , \20205 , \20208 , \20510 , \20511 , \20512 , \20513 , \20514 , \20515 , \20516 , \20517 , \20518 , \20519 , \20520 , \20521 , \20522 , \20523 , \20524 , \20525 , \20526 , \20527 , \20528 , \20529 , \20530 , \20531 , \20532 , \20533 , \20534 );
and \U$14615 ( \20536 , RIeab78c8_6895, \20535 );
buf \U$14616 ( \20537 , \20208 );
buf \U$14617 ( \20538 , \20208 );
buf \U$14618 ( \20539 , \20208 );
buf \U$14619 ( \20540 , \20208 );
buf \U$14620 ( \20541 , \20208 );
buf \U$14621 ( \20542 , \20208 );
buf \U$14622 ( \20543 , \20208 );
buf \U$14623 ( \20544 , \20208 );
buf \U$14624 ( \20545 , \20208 );
buf \U$14625 ( \20546 , \20208 );
buf \U$14626 ( \20547 , \20208 );
buf \U$14627 ( \20548 , \20208 );
buf \U$14628 ( \20549 , \20208 );
buf \U$14629 ( \20550 , \20208 );
buf \U$14630 ( \20551 , \20208 );
buf \U$14631 ( \20552 , \20208 );
buf \U$14632 ( \20553 , \20208 );
buf \U$14633 ( \20554 , \20208 );
buf \U$14634 ( \20555 , \20208 );
buf \U$14635 ( \20556 , \20208 );
buf \U$14636 ( \20557 , \20208 );
buf \U$14637 ( \20558 , \20208 );
buf \U$14638 ( \20559 , \20208 );
buf \U$14639 ( \20560 , \20208 );
buf \U$14640 ( \20561 , \20208 );
nor \U$14641 ( \20562 , \20195 , \20196 , \20238 , \20198 , \20201 , \20205 , \20208 , \20537 , \20538 , \20539 , \20540 , \20541 , \20542 , \20543 , \20544 , \20545 , \20546 , \20547 , \20548 , \20549 , \20550 , \20551 , \20552 , \20553 , \20554 , \20555 , \20556 , \20557 , \20558 , \20559 , \20560 , \20561 );
and \U$14642 ( \20563 , RIeab7d00_6896, \20562 );
buf \U$14643 ( \20564 , \20208 );
buf \U$14644 ( \20565 , \20208 );
buf \U$14645 ( \20566 , \20208 );
buf \U$14646 ( \20567 , \20208 );
buf \U$14647 ( \20568 , \20208 );
buf \U$14648 ( \20569 , \20208 );
buf \U$14649 ( \20570 , \20208 );
buf \U$14650 ( \20571 , \20208 );
buf \U$14651 ( \20572 , \20208 );
buf \U$14652 ( \20573 , \20208 );
buf \U$14653 ( \20574 , \20208 );
buf \U$14654 ( \20575 , \20208 );
buf \U$14655 ( \20576 , \20208 );
buf \U$14656 ( \20577 , \20208 );
buf \U$14657 ( \20578 , \20208 );
buf \U$14658 ( \20579 , \20208 );
buf \U$14659 ( \20580 , \20208 );
buf \U$14660 ( \20581 , \20208 );
buf \U$14661 ( \20582 , \20208 );
buf \U$14662 ( \20583 , \20208 );
buf \U$14663 ( \20584 , \20208 );
buf \U$14664 ( \20585 , \20208 );
buf \U$14665 ( \20586 , \20208 );
buf \U$14666 ( \20587 , \20208 );
buf \U$14667 ( \20588 , \20208 );
nor \U$14668 ( \20589 , \20236 , \20237 , \20197 , \20198 , \20201 , \20205 , \20208 , \20564 , \20565 , \20566 , \20567 , \20568 , \20569 , \20570 , \20571 , \20572 , \20573 , \20574 , \20575 , \20576 , \20577 , \20578 , \20579 , \20580 , \20581 , \20582 , \20583 , \20584 , \20585 , \20586 , \20587 , \20588 );
and \U$14669 ( \20590 , RIeacfa18_6902, \20589 );
buf \U$14670 ( \20591 , \20208 );
buf \U$14671 ( \20592 , \20208 );
buf \U$14672 ( \20593 , \20208 );
buf \U$14673 ( \20594 , \20208 );
buf \U$14674 ( \20595 , \20208 );
buf \U$14675 ( \20596 , \20208 );
buf \U$14676 ( \20597 , \20208 );
buf \U$14677 ( \20598 , \20208 );
buf \U$14678 ( \20599 , \20208 );
buf \U$14679 ( \20600 , \20208 );
buf \U$14680 ( \20601 , \20208 );
buf \U$14681 ( \20602 , \20208 );
buf \U$14682 ( \20603 , \20208 );
buf \U$14683 ( \20604 , \20208 );
buf \U$14684 ( \20605 , \20208 );
buf \U$14685 ( \20606 , \20208 );
buf \U$14686 ( \20607 , \20208 );
buf \U$14687 ( \20608 , \20208 );
buf \U$14688 ( \20609 , \20208 );
buf \U$14689 ( \20610 , \20208 );
buf \U$14690 ( \20611 , \20208 );
buf \U$14691 ( \20612 , \20208 );
buf \U$14692 ( \20613 , \20208 );
buf \U$14693 ( \20614 , \20208 );
buf \U$14694 ( \20615 , \20208 );
nor \U$14695 ( \20616 , \20195 , \20237 , \20197 , \20198 , \20201 , \20205 , \20208 , \20591 , \20592 , \20593 , \20594 , \20595 , \20596 , \20597 , \20598 , \20599 , \20600 , \20601 , \20602 , \20603 , \20604 , \20605 , \20606 , \20607 , \20608 , \20609 , \20610 , \20611 , \20612 , \20613 , \20614 , \20615 );
and \U$14696 ( \20617 , RIeab6518_6891, \20616 );
buf \U$14697 ( \20618 , \20208 );
buf \U$14698 ( \20619 , \20208 );
buf \U$14699 ( \20620 , \20208 );
buf \U$14700 ( \20621 , \20208 );
buf \U$14701 ( \20622 , \20208 );
buf \U$14702 ( \20623 , \20208 );
buf \U$14703 ( \20624 , \20208 );
buf \U$14704 ( \20625 , \20208 );
buf \U$14705 ( \20626 , \20208 );
buf \U$14706 ( \20627 , \20208 );
buf \U$14707 ( \20628 , \20208 );
buf \U$14708 ( \20629 , \20208 );
buf \U$14709 ( \20630 , \20208 );
buf \U$14710 ( \20631 , \20208 );
buf \U$14711 ( \20632 , \20208 );
buf \U$14712 ( \20633 , \20208 );
buf \U$14713 ( \20634 , \20208 );
buf \U$14714 ( \20635 , \20208 );
buf \U$14715 ( \20636 , \20208 );
buf \U$14716 ( \20637 , \20208 );
buf \U$14717 ( \20638 , \20208 );
buf \U$14718 ( \20639 , \20208 );
buf \U$14719 ( \20640 , \20208 );
buf \U$14720 ( \20641 , \20208 );
buf \U$14721 ( \20642 , \20208 );
nor \U$14722 ( \20643 , \20236 , \20196 , \20197 , \20198 , \20201 , \20205 , \20208 , \20618 , \20619 , \20620 , \20621 , \20622 , \20623 , \20624 , \20625 , \20626 , \20627 , \20628 , \20629 , \20630 , \20631 , \20632 , \20633 , \20634 , \20635 , \20636 , \20637 , \20638 , \20639 , \20640 , \20641 , \20642 );
and \U$14723 ( \20644 , RIeb352c8_6904, \20643 );
or \U$14724 ( \20645 , \20235 , \20266 , \20293 , \20320 , \20347 , \20374 , \20401 , \20428 , \20455 , \20482 , \20509 , \20536 , \20563 , \20590 , \20617 , \20644 );
buf \U$14725 ( \20646 , \20208 );
not \U$14726 ( \20647 , \20646 );
buf \U$14727 ( \20648 , \20196 );
buf \U$14728 ( \20649 , \20197 );
buf \U$14729 ( \20650 , \20198 );
buf \U$14730 ( \20651 , \20201 );
buf \U$14731 ( \20652 , \20205 );
buf \U$14732 ( \20653 , \20208 );
buf \U$14733 ( \20654 , \20208 );
buf \U$14734 ( \20655 , \20208 );
buf \U$14735 ( \20656 , \20208 );
buf \U$14736 ( \20657 , \20208 );
buf \U$14737 ( \20658 , \20208 );
buf \U$14738 ( \20659 , \20208 );
buf \U$14739 ( \20660 , \20208 );
buf \U$14740 ( \20661 , \20208 );
buf \U$14741 ( \20662 , \20208 );
buf \U$14742 ( \20663 , \20208 );
buf \U$14743 ( \20664 , \20208 );
buf \U$14744 ( \20665 , \20208 );
buf \U$14745 ( \20666 , \20208 );
buf \U$14746 ( \20667 , \20208 );
buf \U$14747 ( \20668 , \20208 );
buf \U$14748 ( \20669 , \20208 );
buf \U$14749 ( \20670 , \20208 );
buf \U$14750 ( \20671 , \20208 );
buf \U$14751 ( \20672 , \20208 );
buf \U$14752 ( \20673 , \20208 );
buf \U$14753 ( \20674 , \20208 );
buf \U$14754 ( \20675 , \20208 );
buf \U$14755 ( \20676 , \20208 );
buf \U$14756 ( \20677 , \20208 );
buf \U$14757 ( \20678 , \20195 );
or \U$14758 ( \20679 , \20648 , \20649 , \20650 , \20651 , \20652 , \20653 , \20654 , \20655 , \20656 , \20657 , \20658 , \20659 , \20660 , \20661 , \20662 , \20663 , \20664 , \20665 , \20666 , \20667 , \20668 , \20669 , \20670 , \20671 , \20672 , \20673 , \20674 , \20675 , \20676 , \20677 , \20678 );
nand \U$14759 ( \20680 , \20647 , \20679 );
buf \U$14760 ( \20681 , \20680 );
buf \U$14761 ( \20682 , \20208 );
not \U$14762 ( \20683 , \20682 );
buf \U$14763 ( \20684 , \20205 );
buf \U$14764 ( \20685 , \20208 );
buf \U$14765 ( \20686 , \20208 );
buf \U$14766 ( \20687 , \20208 );
buf \U$14767 ( \20688 , \20208 );
buf \U$14768 ( \20689 , \20208 );
buf \U$14769 ( \20690 , \20208 );
buf \U$14770 ( \20691 , \20208 );
buf \U$14771 ( \20692 , \20208 );
buf \U$14772 ( \20693 , \20208 );
buf \U$14773 ( \20694 , \20208 );
buf \U$14774 ( \20695 , \20208 );
buf \U$14775 ( \20696 , \20208 );
buf \U$14776 ( \20697 , \20208 );
buf \U$14777 ( \20698 , \20208 );
buf \U$14778 ( \20699 , \20208 );
buf \U$14779 ( \20700 , \20208 );
buf \U$14780 ( \20701 , \20208 );
buf \U$14781 ( \20702 , \20208 );
buf \U$14782 ( \20703 , \20208 );
buf \U$14783 ( \20704 , \20208 );
buf \U$14784 ( \20705 , \20208 );
buf \U$14785 ( \20706 , \20208 );
buf \U$14786 ( \20707 , \20208 );
buf \U$14787 ( \20708 , \20208 );
buf \U$14788 ( \20709 , \20208 );
buf \U$14789 ( \20710 , \20201 );
buf \U$14790 ( \20711 , \20195 );
buf \U$14791 ( \20712 , \20196 );
buf \U$14792 ( \20713 , \20197 );
buf \U$14793 ( \20714 , \20198 );
or \U$14794 ( \20715 , \20711 , \20712 , \20713 , \20714 );
and \U$14795 ( \20716 , \20710 , \20715 );
or \U$14796 ( \20717 , \20684 , \20685 , \20686 , \20687 , \20688 , \20689 , \20690 , \20691 , \20692 , \20693 , \20694 , \20695 , \20696 , \20697 , \20698 , \20699 , \20700 , \20701 , \20702 , \20703 , \20704 , \20705 , \20706 , \20707 , \20708 , \20709 , \20716 );
and \U$14797 ( \20718 , \20683 , \20717 );
buf \U$14798 ( \20719 , \20718 );
or \U$14799 ( \20720 , \20681 , \20719 );
_DC g67d6 ( \20721_nG67d6 , \20645 , \20720 );
not \U$14800 ( \20722 , \20721_nG67d6 );
buf \U$14801 ( \20723 , RIb7b9608_246);
buf \U$14802 ( \20724 , \20208 );
buf \U$14803 ( \20725 , \20208 );
buf \U$14804 ( \20726 , \20208 );
buf \U$14805 ( \20727 , \20208 );
buf \U$14806 ( \20728 , \20208 );
buf \U$14807 ( \20729 , \20208 );
buf \U$14808 ( \20730 , \20208 );
buf \U$14809 ( \20731 , \20208 );
buf \U$14810 ( \20732 , \20208 );
buf \U$14811 ( \20733 , \20208 );
buf \U$14812 ( \20734 , \20208 );
buf \U$14813 ( \20735 , \20208 );
buf \U$14814 ( \20736 , \20208 );
buf \U$14815 ( \20737 , \20208 );
buf \U$14816 ( \20738 , \20208 );
buf \U$14817 ( \20739 , \20208 );
buf \U$14818 ( \20740 , \20208 );
buf \U$14819 ( \20741 , \20208 );
buf \U$14820 ( \20742 , \20208 );
buf \U$14821 ( \20743 , \20208 );
buf \U$14822 ( \20744 , \20208 );
buf \U$14823 ( \20745 , \20208 );
buf \U$14824 ( \20746 , \20208 );
buf \U$14825 ( \20747 , \20208 );
buf \U$14826 ( \20748 , \20208 );
nor \U$14827 ( \20749 , \20195 , \20196 , \20197 , \20198 , \20202 , \20205 , \20208 , \20724 , \20725 , \20726 , \20727 , \20728 , \20729 , \20730 , \20731 , \20732 , \20733 , \20734 , \20735 , \20736 , \20737 , \20738 , \20739 , \20740 , \20741 , \20742 , \20743 , \20744 , \20745 , \20746 , \20747 , \20748 );
and \U$14828 ( \20750 , \7117 , \20749 );
buf \U$14829 ( \20751 , \20208 );
buf \U$14830 ( \20752 , \20208 );
buf \U$14831 ( \20753 , \20208 );
buf \U$14832 ( \20754 , \20208 );
buf \U$14833 ( \20755 , \20208 );
buf \U$14834 ( \20756 , \20208 );
buf \U$14835 ( \20757 , \20208 );
buf \U$14836 ( \20758 , \20208 );
buf \U$14837 ( \20759 , \20208 );
buf \U$14838 ( \20760 , \20208 );
buf \U$14839 ( \20761 , \20208 );
buf \U$14840 ( \20762 , \20208 );
buf \U$14841 ( \20763 , \20208 );
buf \U$14842 ( \20764 , \20208 );
buf \U$14843 ( \20765 , \20208 );
buf \U$14844 ( \20766 , \20208 );
buf \U$14845 ( \20767 , \20208 );
buf \U$14846 ( \20768 , \20208 );
buf \U$14847 ( \20769 , \20208 );
buf \U$14848 ( \20770 , \20208 );
buf \U$14849 ( \20771 , \20208 );
buf \U$14850 ( \20772 , \20208 );
buf \U$14851 ( \20773 , \20208 );
buf \U$14852 ( \20774 , \20208 );
buf \U$14853 ( \20775 , \20208 );
nor \U$14854 ( \20776 , \20236 , \20237 , \20238 , \20239 , \20201 , \20205 , \20208 , \20751 , \20752 , \20753 , \20754 , \20755 , \20756 , \20757 , \20758 , \20759 , \20760 , \20761 , \20762 , \20763 , \20764 , \20765 , \20766 , \20767 , \20768 , \20769 , \20770 , \20771 , \20772 , \20773 , \20774 , \20775 );
and \U$14855 ( \20777 , \7119 , \20776 );
buf \U$14856 ( \20778 , \20208 );
buf \U$14857 ( \20779 , \20208 );
buf \U$14858 ( \20780 , \20208 );
buf \U$14859 ( \20781 , \20208 );
buf \U$14860 ( \20782 , \20208 );
buf \U$14861 ( \20783 , \20208 );
buf \U$14862 ( \20784 , \20208 );
buf \U$14863 ( \20785 , \20208 );
buf \U$14864 ( \20786 , \20208 );
buf \U$14865 ( \20787 , \20208 );
buf \U$14866 ( \20788 , \20208 );
buf \U$14867 ( \20789 , \20208 );
buf \U$14868 ( \20790 , \20208 );
buf \U$14869 ( \20791 , \20208 );
buf \U$14870 ( \20792 , \20208 );
buf \U$14871 ( \20793 , \20208 );
buf \U$14872 ( \20794 , \20208 );
buf \U$14873 ( \20795 , \20208 );
buf \U$14874 ( \20796 , \20208 );
buf \U$14875 ( \20797 , \20208 );
buf \U$14876 ( \20798 , \20208 );
buf \U$14877 ( \20799 , \20208 );
buf \U$14878 ( \20800 , \20208 );
buf \U$14879 ( \20801 , \20208 );
buf \U$14880 ( \20802 , \20208 );
nor \U$14881 ( \20803 , \20195 , \20237 , \20238 , \20239 , \20201 , \20205 , \20208 , \20778 , \20779 , \20780 , \20781 , \20782 , \20783 , \20784 , \20785 , \20786 , \20787 , \20788 , \20789 , \20790 , \20791 , \20792 , \20793 , \20794 , \20795 , \20796 , \20797 , \20798 , \20799 , \20800 , \20801 , \20802 );
and \U$14882 ( \20804 , \7864 , \20803 );
buf \U$14883 ( \20805 , \20208 );
buf \U$14884 ( \20806 , \20208 );
buf \U$14885 ( \20807 , \20208 );
buf \U$14886 ( \20808 , \20208 );
buf \U$14887 ( \20809 , \20208 );
buf \U$14888 ( \20810 , \20208 );
buf \U$14889 ( \20811 , \20208 );
buf \U$14890 ( \20812 , \20208 );
buf \U$14891 ( \20813 , \20208 );
buf \U$14892 ( \20814 , \20208 );
buf \U$14893 ( \20815 , \20208 );
buf \U$14894 ( \20816 , \20208 );
buf \U$14895 ( \20817 , \20208 );
buf \U$14896 ( \20818 , \20208 );
buf \U$14897 ( \20819 , \20208 );
buf \U$14898 ( \20820 , \20208 );
buf \U$14899 ( \20821 , \20208 );
buf \U$14900 ( \20822 , \20208 );
buf \U$14901 ( \20823 , \20208 );
buf \U$14902 ( \20824 , \20208 );
buf \U$14903 ( \20825 , \20208 );
buf \U$14904 ( \20826 , \20208 );
buf \U$14905 ( \20827 , \20208 );
buf \U$14906 ( \20828 , \20208 );
buf \U$14907 ( \20829 , \20208 );
nor \U$14908 ( \20830 , \20236 , \20196 , \20238 , \20239 , \20201 , \20205 , \20208 , \20805 , \20806 , \20807 , \20808 , \20809 , \20810 , \20811 , \20812 , \20813 , \20814 , \20815 , \20816 , \20817 , \20818 , \20819 , \20820 , \20821 , \20822 , \20823 , \20824 , \20825 , \20826 , \20827 , \20828 , \20829 );
and \U$14909 ( \20831 , \7892 , \20830 );
buf \U$14910 ( \20832 , \20208 );
buf \U$14911 ( \20833 , \20208 );
buf \U$14912 ( \20834 , \20208 );
buf \U$14913 ( \20835 , \20208 );
buf \U$14914 ( \20836 , \20208 );
buf \U$14915 ( \20837 , \20208 );
buf \U$14916 ( \20838 , \20208 );
buf \U$14917 ( \20839 , \20208 );
buf \U$14918 ( \20840 , \20208 );
buf \U$14919 ( \20841 , \20208 );
buf \U$14920 ( \20842 , \20208 );
buf \U$14921 ( \20843 , \20208 );
buf \U$14922 ( \20844 , \20208 );
buf \U$14923 ( \20845 , \20208 );
buf \U$14924 ( \20846 , \20208 );
buf \U$14925 ( \20847 , \20208 );
buf \U$14926 ( \20848 , \20208 );
buf \U$14927 ( \20849 , \20208 );
buf \U$14928 ( \20850 , \20208 );
buf \U$14929 ( \20851 , \20208 );
buf \U$14930 ( \20852 , \20208 );
buf \U$14931 ( \20853 , \20208 );
buf \U$14932 ( \20854 , \20208 );
buf \U$14933 ( \20855 , \20208 );
buf \U$14934 ( \20856 , \20208 );
nor \U$14935 ( \20857 , \20195 , \20196 , \20238 , \20239 , \20201 , \20205 , \20208 , \20832 , \20833 , \20834 , \20835 , \20836 , \20837 , \20838 , \20839 , \20840 , \20841 , \20842 , \20843 , \20844 , \20845 , \20846 , \20847 , \20848 , \20849 , \20850 , \20851 , \20852 , \20853 , \20854 , \20855 , \20856 );
and \U$14936 ( \20858 , \7920 , \20857 );
buf \U$14937 ( \20859 , \20208 );
buf \U$14938 ( \20860 , \20208 );
buf \U$14939 ( \20861 , \20208 );
buf \U$14940 ( \20862 , \20208 );
buf \U$14941 ( \20863 , \20208 );
buf \U$14942 ( \20864 , \20208 );
buf \U$14943 ( \20865 , \20208 );
buf \U$14944 ( \20866 , \20208 );
buf \U$14945 ( \20867 , \20208 );
buf \U$14946 ( \20868 , \20208 );
buf \U$14947 ( \20869 , \20208 );
buf \U$14948 ( \20870 , \20208 );
buf \U$14949 ( \20871 , \20208 );
buf \U$14950 ( \20872 , \20208 );
buf \U$14951 ( \20873 , \20208 );
buf \U$14952 ( \20874 , \20208 );
buf \U$14953 ( \20875 , \20208 );
buf \U$14954 ( \20876 , \20208 );
buf \U$14955 ( \20877 , \20208 );
buf \U$14956 ( \20878 , \20208 );
buf \U$14957 ( \20879 , \20208 );
buf \U$14958 ( \20880 , \20208 );
buf \U$14959 ( \20881 , \20208 );
buf \U$14960 ( \20882 , \20208 );
buf \U$14961 ( \20883 , \20208 );
nor \U$14962 ( \20884 , \20236 , \20237 , \20197 , \20239 , \20201 , \20205 , \20208 , \20859 , \20860 , \20861 , \20862 , \20863 , \20864 , \20865 , \20866 , \20867 , \20868 , \20869 , \20870 , \20871 , \20872 , \20873 , \20874 , \20875 , \20876 , \20877 , \20878 , \20879 , \20880 , \20881 , \20882 , \20883 );
and \U$14963 ( \20885 , \7948 , \20884 );
buf \U$14964 ( \20886 , \20208 );
buf \U$14965 ( \20887 , \20208 );
buf \U$14966 ( \20888 , \20208 );
buf \U$14967 ( \20889 , \20208 );
buf \U$14968 ( \20890 , \20208 );
buf \U$14969 ( \20891 , \20208 );
buf \U$14970 ( \20892 , \20208 );
buf \U$14971 ( \20893 , \20208 );
buf \U$14972 ( \20894 , \20208 );
buf \U$14973 ( \20895 , \20208 );
buf \U$14974 ( \20896 , \20208 );
buf \U$14975 ( \20897 , \20208 );
buf \U$14976 ( \20898 , \20208 );
buf \U$14977 ( \20899 , \20208 );
buf \U$14978 ( \20900 , \20208 );
buf \U$14979 ( \20901 , \20208 );
buf \U$14980 ( \20902 , \20208 );
buf \U$14981 ( \20903 , \20208 );
buf \U$14982 ( \20904 , \20208 );
buf \U$14983 ( \20905 , \20208 );
buf \U$14984 ( \20906 , \20208 );
buf \U$14985 ( \20907 , \20208 );
buf \U$14986 ( \20908 , \20208 );
buf \U$14987 ( \20909 , \20208 );
buf \U$14988 ( \20910 , \20208 );
nor \U$14989 ( \20911 , \20195 , \20237 , \20197 , \20239 , \20201 , \20205 , \20208 , \20886 , \20887 , \20888 , \20889 , \20890 , \20891 , \20892 , \20893 , \20894 , \20895 , \20896 , \20897 , \20898 , \20899 , \20900 , \20901 , \20902 , \20903 , \20904 , \20905 , \20906 , \20907 , \20908 , \20909 , \20910 );
and \U$14990 ( \20912 , \7976 , \20911 );
buf \U$14991 ( \20913 , \20208 );
buf \U$14992 ( \20914 , \20208 );
buf \U$14993 ( \20915 , \20208 );
buf \U$14994 ( \20916 , \20208 );
buf \U$14995 ( \20917 , \20208 );
buf \U$14996 ( \20918 , \20208 );
buf \U$14997 ( \20919 , \20208 );
buf \U$14998 ( \20920 , \20208 );
buf \U$14999 ( \20921 , \20208 );
buf \U$15000 ( \20922 , \20208 );
buf \U$15001 ( \20923 , \20208 );
buf \U$15002 ( \20924 , \20208 );
buf \U$15003 ( \20925 , \20208 );
buf \U$15004 ( \20926 , \20208 );
buf \U$15005 ( \20927 , \20208 );
buf \U$15006 ( \20928 , \20208 );
buf \U$15007 ( \20929 , \20208 );
buf \U$15008 ( \20930 , \20208 );
buf \U$15009 ( \20931 , \20208 );
buf \U$15010 ( \20932 , \20208 );
buf \U$15011 ( \20933 , \20208 );
buf \U$15012 ( \20934 , \20208 );
buf \U$15013 ( \20935 , \20208 );
buf \U$15014 ( \20936 , \20208 );
buf \U$15015 ( \20937 , \20208 );
nor \U$15016 ( \20938 , \20236 , \20196 , \20197 , \20239 , \20201 , \20205 , \20208 , \20913 , \20914 , \20915 , \20916 , \20917 , \20918 , \20919 , \20920 , \20921 , \20922 , \20923 , \20924 , \20925 , \20926 , \20927 , \20928 , \20929 , \20930 , \20931 , \20932 , \20933 , \20934 , \20935 , \20936 , \20937 );
and \U$15017 ( \20939 , \8004 , \20938 );
buf \U$15018 ( \20940 , \20208 );
buf \U$15019 ( \20941 , \20208 );
buf \U$15020 ( \20942 , \20208 );
buf \U$15021 ( \20943 , \20208 );
buf \U$15022 ( \20944 , \20208 );
buf \U$15023 ( \20945 , \20208 );
buf \U$15024 ( \20946 , \20208 );
buf \U$15025 ( \20947 , \20208 );
buf \U$15026 ( \20948 , \20208 );
buf \U$15027 ( \20949 , \20208 );
buf \U$15028 ( \20950 , \20208 );
buf \U$15029 ( \20951 , \20208 );
buf \U$15030 ( \20952 , \20208 );
buf \U$15031 ( \20953 , \20208 );
buf \U$15032 ( \20954 , \20208 );
buf \U$15033 ( \20955 , \20208 );
buf \U$15034 ( \20956 , \20208 );
buf \U$15035 ( \20957 , \20208 );
buf \U$15036 ( \20958 , \20208 );
buf \U$15037 ( \20959 , \20208 );
buf \U$15038 ( \20960 , \20208 );
buf \U$15039 ( \20961 , \20208 );
buf \U$15040 ( \20962 , \20208 );
buf \U$15041 ( \20963 , \20208 );
buf \U$15042 ( \20964 , \20208 );
nor \U$15043 ( \20965 , \20195 , \20196 , \20197 , \20239 , \20201 , \20205 , \20208 , \20940 , \20941 , \20942 , \20943 , \20944 , \20945 , \20946 , \20947 , \20948 , \20949 , \20950 , \20951 , \20952 , \20953 , \20954 , \20955 , \20956 , \20957 , \20958 , \20959 , \20960 , \20961 , \20962 , \20963 , \20964 );
and \U$15044 ( \20966 , \8032 , \20965 );
buf \U$15045 ( \20967 , \20208 );
buf \U$15046 ( \20968 , \20208 );
buf \U$15047 ( \20969 , \20208 );
buf \U$15048 ( \20970 , \20208 );
buf \U$15049 ( \20971 , \20208 );
buf \U$15050 ( \20972 , \20208 );
buf \U$15051 ( \20973 , \20208 );
buf \U$15052 ( \20974 , \20208 );
buf \U$15053 ( \20975 , \20208 );
buf \U$15054 ( \20976 , \20208 );
buf \U$15055 ( \20977 , \20208 );
buf \U$15056 ( \20978 , \20208 );
buf \U$15057 ( \20979 , \20208 );
buf \U$15058 ( \20980 , \20208 );
buf \U$15059 ( \20981 , \20208 );
buf \U$15060 ( \20982 , \20208 );
buf \U$15061 ( \20983 , \20208 );
buf \U$15062 ( \20984 , \20208 );
buf \U$15063 ( \20985 , \20208 );
buf \U$15064 ( \20986 , \20208 );
buf \U$15065 ( \20987 , \20208 );
buf \U$15066 ( \20988 , \20208 );
buf \U$15067 ( \20989 , \20208 );
buf \U$15068 ( \20990 , \20208 );
buf \U$15069 ( \20991 , \20208 );
nor \U$15070 ( \20992 , \20236 , \20237 , \20238 , \20198 , \20201 , \20205 , \20208 , \20967 , \20968 , \20969 , \20970 , \20971 , \20972 , \20973 , \20974 , \20975 , \20976 , \20977 , \20978 , \20979 , \20980 , \20981 , \20982 , \20983 , \20984 , \20985 , \20986 , \20987 , \20988 , \20989 , \20990 , \20991 );
and \U$15071 ( \20993 , \8060 , \20992 );
buf \U$15072 ( \20994 , \20208 );
buf \U$15073 ( \20995 , \20208 );
buf \U$15074 ( \20996 , \20208 );
buf \U$15075 ( \20997 , \20208 );
buf \U$15076 ( \20998 , \20208 );
buf \U$15077 ( \20999 , \20208 );
buf \U$15078 ( \21000 , \20208 );
buf \U$15079 ( \21001 , \20208 );
buf \U$15080 ( \21002 , \20208 );
buf \U$15081 ( \21003 , \20208 );
buf \U$15082 ( \21004 , \20208 );
buf \U$15083 ( \21005 , \20208 );
buf \U$15084 ( \21006 , \20208 );
buf \U$15085 ( \21007 , \20208 );
buf \U$15086 ( \21008 , \20208 );
buf \U$15087 ( \21009 , \20208 );
buf \U$15088 ( \21010 , \20208 );
buf \U$15089 ( \21011 , \20208 );
buf \U$15090 ( \21012 , \20208 );
buf \U$15091 ( \21013 , \20208 );
buf \U$15092 ( \21014 , \20208 );
buf \U$15093 ( \21015 , \20208 );
buf \U$15094 ( \21016 , \20208 );
buf \U$15095 ( \21017 , \20208 );
buf \U$15096 ( \21018 , \20208 );
nor \U$15097 ( \21019 , \20195 , \20237 , \20238 , \20198 , \20201 , \20205 , \20208 , \20994 , \20995 , \20996 , \20997 , \20998 , \20999 , \21000 , \21001 , \21002 , \21003 , \21004 , \21005 , \21006 , \21007 , \21008 , \21009 , \21010 , \21011 , \21012 , \21013 , \21014 , \21015 , \21016 , \21017 , \21018 );
and \U$15098 ( \21020 , \8088 , \21019 );
buf \U$15099 ( \21021 , \20208 );
buf \U$15100 ( \21022 , \20208 );
buf \U$15101 ( \21023 , \20208 );
buf \U$15102 ( \21024 , \20208 );
buf \U$15103 ( \21025 , \20208 );
buf \U$15104 ( \21026 , \20208 );
buf \U$15105 ( \21027 , \20208 );
buf \U$15106 ( \21028 , \20208 );
buf \U$15107 ( \21029 , \20208 );
buf \U$15108 ( \21030 , \20208 );
buf \U$15109 ( \21031 , \20208 );
buf \U$15110 ( \21032 , \20208 );
buf \U$15111 ( \21033 , \20208 );
buf \U$15112 ( \21034 , \20208 );
buf \U$15113 ( \21035 , \20208 );
buf \U$15114 ( \21036 , \20208 );
buf \U$15115 ( \21037 , \20208 );
buf \U$15116 ( \21038 , \20208 );
buf \U$15117 ( \21039 , \20208 );
buf \U$15118 ( \21040 , \20208 );
buf \U$15119 ( \21041 , \20208 );
buf \U$15120 ( \21042 , \20208 );
buf \U$15121 ( \21043 , \20208 );
buf \U$15122 ( \21044 , \20208 );
buf \U$15123 ( \21045 , \20208 );
nor \U$15124 ( \21046 , \20236 , \20196 , \20238 , \20198 , \20201 , \20205 , \20208 , \21021 , \21022 , \21023 , \21024 , \21025 , \21026 , \21027 , \21028 , \21029 , \21030 , \21031 , \21032 , \21033 , \21034 , \21035 , \21036 , \21037 , \21038 , \21039 , \21040 , \21041 , \21042 , \21043 , \21044 , \21045 );
and \U$15125 ( \21047 , \8116 , \21046 );
buf \U$15126 ( \21048 , \20208 );
buf \U$15127 ( \21049 , \20208 );
buf \U$15128 ( \21050 , \20208 );
buf \U$15129 ( \21051 , \20208 );
buf \U$15130 ( \21052 , \20208 );
buf \U$15131 ( \21053 , \20208 );
buf \U$15132 ( \21054 , \20208 );
buf \U$15133 ( \21055 , \20208 );
buf \U$15134 ( \21056 , \20208 );
buf \U$15135 ( \21057 , \20208 );
buf \U$15136 ( \21058 , \20208 );
buf \U$15137 ( \21059 , \20208 );
buf \U$15138 ( \21060 , \20208 );
buf \U$15139 ( \21061 , \20208 );
buf \U$15140 ( \21062 , \20208 );
buf \U$15141 ( \21063 , \20208 );
buf \U$15142 ( \21064 , \20208 );
buf \U$15143 ( \21065 , \20208 );
buf \U$15144 ( \21066 , \20208 );
buf \U$15145 ( \21067 , \20208 );
buf \U$15146 ( \21068 , \20208 );
buf \U$15147 ( \21069 , \20208 );
buf \U$15148 ( \21070 , \20208 );
buf \U$15149 ( \21071 , \20208 );
buf \U$15150 ( \21072 , \20208 );
nor \U$15151 ( \21073 , \20195 , \20196 , \20238 , \20198 , \20201 , \20205 , \20208 , \21048 , \21049 , \21050 , \21051 , \21052 , \21053 , \21054 , \21055 , \21056 , \21057 , \21058 , \21059 , \21060 , \21061 , \21062 , \21063 , \21064 , \21065 , \21066 , \21067 , \21068 , \21069 , \21070 , \21071 , \21072 );
and \U$15152 ( \21074 , \8144 , \21073 );
buf \U$15153 ( \21075 , \20208 );
buf \U$15154 ( \21076 , \20208 );
buf \U$15155 ( \21077 , \20208 );
buf \U$15156 ( \21078 , \20208 );
buf \U$15157 ( \21079 , \20208 );
buf \U$15158 ( \21080 , \20208 );
buf \U$15159 ( \21081 , \20208 );
buf \U$15160 ( \21082 , \20208 );
buf \U$15161 ( \21083 , \20208 );
buf \U$15162 ( \21084 , \20208 );
buf \U$15163 ( \21085 , \20208 );
buf \U$15164 ( \21086 , \20208 );
buf \U$15165 ( \21087 , \20208 );
buf \U$15166 ( \21088 , \20208 );
buf \U$15167 ( \21089 , \20208 );
buf \U$15168 ( \21090 , \20208 );
buf \U$15169 ( \21091 , \20208 );
buf \U$15170 ( \21092 , \20208 );
buf \U$15171 ( \21093 , \20208 );
buf \U$15172 ( \21094 , \20208 );
buf \U$15173 ( \21095 , \20208 );
buf \U$15174 ( \21096 , \20208 );
buf \U$15175 ( \21097 , \20208 );
buf \U$15176 ( \21098 , \20208 );
buf \U$15177 ( \21099 , \20208 );
nor \U$15178 ( \21100 , \20236 , \20237 , \20197 , \20198 , \20201 , \20205 , \20208 , \21075 , \21076 , \21077 , \21078 , \21079 , \21080 , \21081 , \21082 , \21083 , \21084 , \21085 , \21086 , \21087 , \21088 , \21089 , \21090 , \21091 , \21092 , \21093 , \21094 , \21095 , \21096 , \21097 , \21098 , \21099 );
and \U$15179 ( \21101 , \8172 , \21100 );
buf \U$15180 ( \21102 , \20208 );
buf \U$15181 ( \21103 , \20208 );
buf \U$15182 ( \21104 , \20208 );
buf \U$15183 ( \21105 , \20208 );
buf \U$15184 ( \21106 , \20208 );
buf \U$15185 ( \21107 , \20208 );
buf \U$15186 ( \21108 , \20208 );
buf \U$15187 ( \21109 , \20208 );
buf \U$15188 ( \21110 , \20208 );
buf \U$15189 ( \21111 , \20208 );
buf \U$15190 ( \21112 , \20208 );
buf \U$15191 ( \21113 , \20208 );
buf \U$15192 ( \21114 , \20208 );
buf \U$15193 ( \21115 , \20208 );
buf \U$15194 ( \21116 , \20208 );
buf \U$15195 ( \21117 , \20208 );
buf \U$15196 ( \21118 , \20208 );
buf \U$15197 ( \21119 , \20208 );
buf \U$15198 ( \21120 , \20208 );
buf \U$15199 ( \21121 , \20208 );
buf \U$15200 ( \21122 , \20208 );
buf \U$15201 ( \21123 , \20208 );
buf \U$15202 ( \21124 , \20208 );
buf \U$15203 ( \21125 , \20208 );
buf \U$15204 ( \21126 , \20208 );
nor \U$15205 ( \21127 , \20195 , \20237 , \20197 , \20198 , \20201 , \20205 , \20208 , \21102 , \21103 , \21104 , \21105 , \21106 , \21107 , \21108 , \21109 , \21110 , \21111 , \21112 , \21113 , \21114 , \21115 , \21116 , \21117 , \21118 , \21119 , \21120 , \21121 , \21122 , \21123 , \21124 , \21125 , \21126 );
and \U$15206 ( \21128 , \8200 , \21127 );
buf \U$15207 ( \21129 , \20208 );
buf \U$15208 ( \21130 , \20208 );
buf \U$15209 ( \21131 , \20208 );
buf \U$15210 ( \21132 , \20208 );
buf \U$15211 ( \21133 , \20208 );
buf \U$15212 ( \21134 , \20208 );
buf \U$15213 ( \21135 , \20208 );
buf \U$15214 ( \21136 , \20208 );
buf \U$15215 ( \21137 , \20208 );
buf \U$15216 ( \21138 , \20208 );
buf \U$15217 ( \21139 , \20208 );
buf \U$15218 ( \21140 , \20208 );
buf \U$15219 ( \21141 , \20208 );
buf \U$15220 ( \21142 , \20208 );
buf \U$15221 ( \21143 , \20208 );
buf \U$15222 ( \21144 , \20208 );
buf \U$15223 ( \21145 , \20208 );
buf \U$15224 ( \21146 , \20208 );
buf \U$15225 ( \21147 , \20208 );
buf \U$15226 ( \21148 , \20208 );
buf \U$15227 ( \21149 , \20208 );
buf \U$15228 ( \21150 , \20208 );
buf \U$15229 ( \21151 , \20208 );
buf \U$15230 ( \21152 , \20208 );
buf \U$15231 ( \21153 , \20208 );
nor \U$15232 ( \21154 , \20236 , \20196 , \20197 , \20198 , \20201 , \20205 , \20208 , \21129 , \21130 , \21131 , \21132 , \21133 , \21134 , \21135 , \21136 , \21137 , \21138 , \21139 , \21140 , \21141 , \21142 , \21143 , \21144 , \21145 , \21146 , \21147 , \21148 , \21149 , \21150 , \21151 , \21152 , \21153 );
and \U$15233 ( \21155 , \8228 , \21154 );
or \U$15234 ( \21156 , \20750 , \20777 , \20804 , \20831 , \20858 , \20885 , \20912 , \20939 , \20966 , \20993 , \21020 , \21047 , \21074 , \21101 , \21128 , \21155 );
buf \U$15235 ( \21157 , \20208 );
not \U$15236 ( \21158 , \21157 );
buf \U$15237 ( \21159 , \20196 );
buf \U$15238 ( \21160 , \20197 );
buf \U$15239 ( \21161 , \20198 );
buf \U$15240 ( \21162 , \20201 );
buf \U$15241 ( \21163 , \20205 );
buf \U$15242 ( \21164 , \20208 );
buf \U$15243 ( \21165 , \20208 );
buf \U$15244 ( \21166 , \20208 );
buf \U$15245 ( \21167 , \20208 );
buf \U$15246 ( \21168 , \20208 );
buf \U$15247 ( \21169 , \20208 );
buf \U$15248 ( \21170 , \20208 );
buf \U$15249 ( \21171 , \20208 );
buf \U$15250 ( \21172 , \20208 );
buf \U$15251 ( \21173 , \20208 );
buf \U$15252 ( \21174 , \20208 );
buf \U$15253 ( \21175 , \20208 );
buf \U$15254 ( \21176 , \20208 );
buf \U$15255 ( \21177 , \20208 );
buf \U$15256 ( \21178 , \20208 );
buf \U$15257 ( \21179 , \20208 );
buf \U$15258 ( \21180 , \20208 );
buf \U$15259 ( \21181 , \20208 );
buf \U$15260 ( \21182 , \20208 );
buf \U$15261 ( \21183 , \20208 );
buf \U$15262 ( \21184 , \20208 );
buf \U$15263 ( \21185 , \20208 );
buf \U$15264 ( \21186 , \20208 );
buf \U$15265 ( \21187 , \20208 );
buf \U$15266 ( \21188 , \20208 );
buf \U$15267 ( \21189 , \20195 );
or \U$15268 ( \21190 , \21159 , \21160 , \21161 , \21162 , \21163 , \21164 , \21165 , \21166 , \21167 , \21168 , \21169 , \21170 , \21171 , \21172 , \21173 , \21174 , \21175 , \21176 , \21177 , \21178 , \21179 , \21180 , \21181 , \21182 , \21183 , \21184 , \21185 , \21186 , \21187 , \21188 , \21189 );
nand \U$15269 ( \21191 , \21158 , \21190 );
buf \U$15270 ( \21192 , \21191 );
buf \U$15271 ( \21193 , \20208 );
not \U$15272 ( \21194 , \21193 );
buf \U$15273 ( \21195 , \20205 );
buf \U$15274 ( \21196 , \20208 );
buf \U$15275 ( \21197 , \20208 );
buf \U$15276 ( \21198 , \20208 );
buf \U$15277 ( \21199 , \20208 );
buf \U$15278 ( \21200 , \20208 );
buf \U$15279 ( \21201 , \20208 );
buf \U$15280 ( \21202 , \20208 );
buf \U$15281 ( \21203 , \20208 );
buf \U$15282 ( \21204 , \20208 );
buf \U$15283 ( \21205 , \20208 );
buf \U$15284 ( \21206 , \20208 );
buf \U$15285 ( \21207 , \20208 );
buf \U$15286 ( \21208 , \20208 );
buf \U$15287 ( \21209 , \20208 );
buf \U$15288 ( \21210 , \20208 );
buf \U$15289 ( \21211 , \20208 );
buf \U$15290 ( \21212 , \20208 );
buf \U$15291 ( \21213 , \20208 );
buf \U$15292 ( \21214 , \20208 );
buf \U$15293 ( \21215 , \20208 );
buf \U$15294 ( \21216 , \20208 );
buf \U$15295 ( \21217 , \20208 );
buf \U$15296 ( \21218 , \20208 );
buf \U$15297 ( \21219 , \20208 );
buf \U$15298 ( \21220 , \20208 );
buf \U$15299 ( \21221 , \20201 );
buf \U$15300 ( \21222 , \20195 );
buf \U$15301 ( \21223 , \20196 );
buf \U$15302 ( \21224 , \20197 );
buf \U$15303 ( \21225 , \20198 );
or \U$15304 ( \21226 , \21222 , \21223 , \21224 , \21225 );
and \U$15305 ( \21227 , \21221 , \21226 );
or \U$15306 ( \21228 , \21195 , \21196 , \21197 , \21198 , \21199 , \21200 , \21201 , \21202 , \21203 , \21204 , \21205 , \21206 , \21207 , \21208 , \21209 , \21210 , \21211 , \21212 , \21213 , \21214 , \21215 , \21216 , \21217 , \21218 , \21219 , \21220 , \21227 );
and \U$15307 ( \21229 , \21194 , \21228 );
buf \U$15308 ( \21230 , \21229 );
or \U$15309 ( \21231 , \21192 , \21230 );
_DC g69d5 ( \21232_nG69d5 , \21156 , \21231 );
buf \U$15310 ( \21233 , \21232_nG69d5 );
xor \U$15311 ( \21234 , \20723 , \21233 );
buf \U$15312 ( \21235 , RIb7b9590_247);
and \U$15313 ( \21236 , \7126 , \20749 );
and \U$15314 ( \21237 , \7128 , \20776 );
and \U$15315 ( \21238 , \8338 , \20803 );
and \U$15316 ( \21239 , \8340 , \20830 );
and \U$15317 ( \21240 , \8342 , \20857 );
and \U$15318 ( \21241 , \8344 , \20884 );
and \U$15319 ( \21242 , \8346 , \20911 );
and \U$15320 ( \21243 , \8348 , \20938 );
and \U$15321 ( \21244 , \8350 , \20965 );
and \U$15322 ( \21245 , \8352 , \20992 );
and \U$15323 ( \21246 , \8354 , \21019 );
and \U$15324 ( \21247 , \8356 , \21046 );
and \U$15325 ( \21248 , \8358 , \21073 );
and \U$15326 ( \21249 , \8360 , \21100 );
and \U$15327 ( \21250 , \8362 , \21127 );
and \U$15328 ( \21251 , \8364 , \21154 );
or \U$15329 ( \21252 , \21236 , \21237 , \21238 , \21239 , \21240 , \21241 , \21242 , \21243 , \21244 , \21245 , \21246 , \21247 , \21248 , \21249 , \21250 , \21251 );
_DC g69ea ( \21253_nG69ea , \21252 , \21231 );
buf \U$15330 ( \21254 , \21253_nG69ea );
xor \U$15331 ( \21255 , \21235 , \21254 );
or \U$15332 ( \21256 , \21234 , \21255 );
buf \U$15333 ( \21257 , RIb7b9518_248);
and \U$15334 ( \21258 , \7136 , \20749 );
and \U$15335 ( \21259 , \7138 , \20776 );
and \U$15336 ( \21260 , \8374 , \20803 );
and \U$15337 ( \21261 , \8376 , \20830 );
and \U$15338 ( \21262 , \8378 , \20857 );
and \U$15339 ( \21263 , \8380 , \20884 );
and \U$15340 ( \21264 , \8382 , \20911 );
and \U$15341 ( \21265 , \8384 , \20938 );
and \U$15342 ( \21266 , \8386 , \20965 );
and \U$15343 ( \21267 , \8388 , \20992 );
and \U$15344 ( \21268 , \8390 , \21019 );
and \U$15345 ( \21269 , \8392 , \21046 );
and \U$15346 ( \21270 , \8394 , \21073 );
and \U$15347 ( \21271 , \8396 , \21100 );
and \U$15348 ( \21272 , \8398 , \21127 );
and \U$15349 ( \21273 , \8400 , \21154 );
or \U$15350 ( \21274 , \21258 , \21259 , \21260 , \21261 , \21262 , \21263 , \21264 , \21265 , \21266 , \21267 , \21268 , \21269 , \21270 , \21271 , \21272 , \21273 );
_DC g6a00 ( \21275_nG6a00 , \21274 , \21231 );
buf \U$15351 ( \21276 , \21275_nG6a00 );
xor \U$15352 ( \21277 , \21257 , \21276 );
or \U$15353 ( \21278 , \21256 , \21277 );
buf \U$15354 ( \21279 , RIb7b94a0_249);
and \U$15355 ( \21280 , \7146 , \20749 );
and \U$15356 ( \21281 , \7148 , \20776 );
and \U$15357 ( \21282 , \8410 , \20803 );
and \U$15358 ( \21283 , \8412 , \20830 );
and \U$15359 ( \21284 , \8414 , \20857 );
and \U$15360 ( \21285 , \8416 , \20884 );
and \U$15361 ( \21286 , \8418 , \20911 );
and \U$15362 ( \21287 , \8420 , \20938 );
and \U$15363 ( \21288 , \8422 , \20965 );
and \U$15364 ( \21289 , \8424 , \20992 );
and \U$15365 ( \21290 , \8426 , \21019 );
and \U$15366 ( \21291 , \8428 , \21046 );
and \U$15367 ( \21292 , \8430 , \21073 );
and \U$15368 ( \21293 , \8432 , \21100 );
and \U$15369 ( \21294 , \8434 , \21127 );
and \U$15370 ( \21295 , \8436 , \21154 );
or \U$15371 ( \21296 , \21280 , \21281 , \21282 , \21283 , \21284 , \21285 , \21286 , \21287 , \21288 , \21289 , \21290 , \21291 , \21292 , \21293 , \21294 , \21295 );
_DC g6a16 ( \21297_nG6a16 , \21296 , \21231 );
buf \U$15372 ( \21298 , \21297_nG6a16 );
xor \U$15373 ( \21299 , \21279 , \21298 );
or \U$15374 ( \21300 , \21278 , \21299 );
buf \U$15375 ( \21301 , RIb7b9428_250);
and \U$15376 ( \21302 , \7156 , \20749 );
and \U$15377 ( \21303 , \7158 , \20776 );
and \U$15378 ( \21304 , \8446 , \20803 );
and \U$15379 ( \21305 , \8448 , \20830 );
and \U$15380 ( \21306 , \8450 , \20857 );
and \U$15381 ( \21307 , \8452 , \20884 );
and \U$15382 ( \21308 , \8454 , \20911 );
and \U$15383 ( \21309 , \8456 , \20938 );
and \U$15384 ( \21310 , \8458 , \20965 );
and \U$15385 ( \21311 , \8460 , \20992 );
and \U$15386 ( \21312 , \8462 , \21019 );
and \U$15387 ( \21313 , \8464 , \21046 );
and \U$15388 ( \21314 , \8466 , \21073 );
and \U$15389 ( \21315 , \8468 , \21100 );
and \U$15390 ( \21316 , \8470 , \21127 );
and \U$15391 ( \21317 , \8472 , \21154 );
or \U$15392 ( \21318 , \21302 , \21303 , \21304 , \21305 , \21306 , \21307 , \21308 , \21309 , \21310 , \21311 , \21312 , \21313 , \21314 , \21315 , \21316 , \21317 );
_DC g6a2c ( \21319_nG6a2c , \21318 , \21231 );
buf \U$15393 ( \21320 , \21319_nG6a2c );
xor \U$15394 ( \21321 , \21301 , \21320 );
or \U$15395 ( \21322 , \21300 , \21321 );
buf \U$15396 ( \21323 , RIb7b93b0_251);
and \U$15397 ( \21324 , \7166 , \20749 );
and \U$15398 ( \21325 , \7168 , \20776 );
and \U$15399 ( \21326 , \8482 , \20803 );
and \U$15400 ( \21327 , \8484 , \20830 );
and \U$15401 ( \21328 , \8486 , \20857 );
and \U$15402 ( \21329 , \8488 , \20884 );
and \U$15403 ( \21330 , \8490 , \20911 );
and \U$15404 ( \21331 , \8492 , \20938 );
and \U$15405 ( \21332 , \8494 , \20965 );
and \U$15406 ( \21333 , \8496 , \20992 );
and \U$15407 ( \21334 , \8498 , \21019 );
and \U$15408 ( \21335 , \8500 , \21046 );
and \U$15409 ( \21336 , \8502 , \21073 );
and \U$15410 ( \21337 , \8504 , \21100 );
and \U$15411 ( \21338 , \8506 , \21127 );
and \U$15412 ( \21339 , \8508 , \21154 );
or \U$15413 ( \21340 , \21324 , \21325 , \21326 , \21327 , \21328 , \21329 , \21330 , \21331 , \21332 , \21333 , \21334 , \21335 , \21336 , \21337 , \21338 , \21339 );
_DC g6a42 ( \21341_nG6a42 , \21340 , \21231 );
buf \U$15414 ( \21342 , \21341_nG6a42 );
xor \U$15415 ( \21343 , \21323 , \21342 );
or \U$15416 ( \21344 , \21322 , \21343 );
buf \U$15417 ( \21345 , RIb7af720_252);
and \U$15418 ( \21346 , \7176 , \20749 );
and \U$15419 ( \21347 , \7178 , \20776 );
and \U$15420 ( \21348 , \8518 , \20803 );
and \U$15421 ( \21349 , \8520 , \20830 );
and \U$15422 ( \21350 , \8522 , \20857 );
and \U$15423 ( \21351 , \8524 , \20884 );
and \U$15424 ( \21352 , \8526 , \20911 );
and \U$15425 ( \21353 , \8528 , \20938 );
and \U$15426 ( \21354 , \8530 , \20965 );
and \U$15427 ( \21355 , \8532 , \20992 );
and \U$15428 ( \21356 , \8534 , \21019 );
and \U$15429 ( \21357 , \8536 , \21046 );
and \U$15430 ( \21358 , \8538 , \21073 );
and \U$15431 ( \21359 , \8540 , \21100 );
and \U$15432 ( \21360 , \8542 , \21127 );
and \U$15433 ( \21361 , \8544 , \21154 );
or \U$15434 ( \21362 , \21346 , \21347 , \21348 , \21349 , \21350 , \21351 , \21352 , \21353 , \21354 , \21355 , \21356 , \21357 , \21358 , \21359 , \21360 , \21361 );
_DC g6a58 ( \21363_nG6a58 , \21362 , \21231 );
buf \U$15435 ( \21364 , \21363_nG6a58 );
xor \U$15436 ( \21365 , \21345 , \21364 );
or \U$15437 ( \21366 , \21344 , \21365 );
buf \U$15438 ( \21367 , RIb7af6a8_253);
and \U$15439 ( \21368 , \7186 , \20749 );
and \U$15440 ( \21369 , \7188 , \20776 );
and \U$15441 ( \21370 , \8554 , \20803 );
and \U$15442 ( \21371 , \8556 , \20830 );
and \U$15443 ( \21372 , \8558 , \20857 );
and \U$15444 ( \21373 , \8560 , \20884 );
and \U$15445 ( \21374 , \8562 , \20911 );
and \U$15446 ( \21375 , \8564 , \20938 );
and \U$15447 ( \21376 , \8566 , \20965 );
and \U$15448 ( \21377 , \8568 , \20992 );
and \U$15449 ( \21378 , \8570 , \21019 );
and \U$15450 ( \21379 , \8572 , \21046 );
and \U$15451 ( \21380 , \8574 , \21073 );
and \U$15452 ( \21381 , \8576 , \21100 );
and \U$15453 ( \21382 , \8578 , \21127 );
and \U$15454 ( \21383 , \8580 , \21154 );
or \U$15455 ( \21384 , \21368 , \21369 , \21370 , \21371 , \21372 , \21373 , \21374 , \21375 , \21376 , \21377 , \21378 , \21379 , \21380 , \21381 , \21382 , \21383 );
_DC g6a6e ( \21385_nG6a6e , \21384 , \21231 );
buf \U$15456 ( \21386 , \21385_nG6a6e );
xor \U$15457 ( \21387 , \21367 , \21386 );
or \U$15458 ( \21388 , \21366 , \21387 );
not \U$15459 ( \21389 , \21388 );
buf \U$15460 ( \21390 , \21389 );
and \U$15461 ( \21391 , \20722 , \21390 );
buf \U$15462 ( \21392 , RIb7af630_254);
buf \U$15463 ( \21393 , \20208 );
buf \U$15464 ( \21394 , \20208 );
buf \U$15465 ( \21395 , \20208 );
buf \U$15466 ( \21396 , \20208 );
buf \U$15467 ( \21397 , \20208 );
buf \U$15468 ( \21398 , \20208 );
buf \U$15469 ( \21399 , \20208 );
buf \U$15470 ( \21400 , \20208 );
buf \U$15471 ( \21401 , \20208 );
buf \U$15472 ( \21402 , \20208 );
buf \U$15473 ( \21403 , \20208 );
buf \U$15474 ( \21404 , \20208 );
buf \U$15475 ( \21405 , \20208 );
buf \U$15476 ( \21406 , \20208 );
buf \U$15477 ( \21407 , \20208 );
buf \U$15478 ( \21408 , \20208 );
buf \U$15479 ( \21409 , \20208 );
buf \U$15480 ( \21410 , \20208 );
buf \U$15481 ( \21411 , \20208 );
buf \U$15482 ( \21412 , \20208 );
buf \U$15483 ( \21413 , \20208 );
buf \U$15484 ( \21414 , \20208 );
buf \U$15485 ( \21415 , \20208 );
buf \U$15486 ( \21416 , \20208 );
buf \U$15487 ( \21417 , \20208 );
nor \U$15488 ( \21418 , \20195 , \20196 , \20197 , \20198 , \20202 , \20205 , \20208 , \21393 , \21394 , \21395 , \21396 , \21397 , \21398 , \21399 , \21400 , \21401 , \21402 , \21403 , \21404 , \21405 , \21406 , \21407 , \21408 , \21409 , \21410 , \21411 , \21412 , \21413 , \21414 , \21415 , \21416 , \21417 );
and \U$15489 ( \21419 , \7198 , \21418 );
buf \U$15490 ( \21420 , \20208 );
buf \U$15491 ( \21421 , \20208 );
buf \U$15492 ( \21422 , \20208 );
buf \U$15493 ( \21423 , \20208 );
buf \U$15494 ( \21424 , \20208 );
buf \U$15495 ( \21425 , \20208 );
buf \U$15496 ( \21426 , \20208 );
buf \U$15497 ( \21427 , \20208 );
buf \U$15498 ( \21428 , \20208 );
buf \U$15499 ( \21429 , \20208 );
buf \U$15500 ( \21430 , \20208 );
buf \U$15501 ( \21431 , \20208 );
buf \U$15502 ( \21432 , \20208 );
buf \U$15503 ( \21433 , \20208 );
buf \U$15504 ( \21434 , \20208 );
buf \U$15505 ( \21435 , \20208 );
buf \U$15506 ( \21436 , \20208 );
buf \U$15507 ( \21437 , \20208 );
buf \U$15508 ( \21438 , \20208 );
buf \U$15509 ( \21439 , \20208 );
buf \U$15510 ( \21440 , \20208 );
buf \U$15511 ( \21441 , \20208 );
buf \U$15512 ( \21442 , \20208 );
buf \U$15513 ( \21443 , \20208 );
buf \U$15514 ( \21444 , \20208 );
nor \U$15515 ( \21445 , \20236 , \20237 , \20238 , \20239 , \20201 , \20205 , \20208 , \21420 , \21421 , \21422 , \21423 , \21424 , \21425 , \21426 , \21427 , \21428 , \21429 , \21430 , \21431 , \21432 , \21433 , \21434 , \21435 , \21436 , \21437 , \21438 , \21439 , \21440 , \21441 , \21442 , \21443 , \21444 );
and \U$15516 ( \21446 , \7200 , \21445 );
buf \U$15517 ( \21447 , \20208 );
buf \U$15518 ( \21448 , \20208 );
buf \U$15519 ( \21449 , \20208 );
buf \U$15520 ( \21450 , \20208 );
buf \U$15521 ( \21451 , \20208 );
buf \U$15522 ( \21452 , \20208 );
buf \U$15523 ( \21453 , \20208 );
buf \U$15524 ( \21454 , \20208 );
buf \U$15525 ( \21455 , \20208 );
buf \U$15526 ( \21456 , \20208 );
buf \U$15527 ( \21457 , \20208 );
buf \U$15528 ( \21458 , \20208 );
buf \U$15529 ( \21459 , \20208 );
buf \U$15530 ( \21460 , \20208 );
buf \U$15531 ( \21461 , \20208 );
buf \U$15532 ( \21462 , \20208 );
buf \U$15533 ( \21463 , \20208 );
buf \U$15534 ( \21464 , \20208 );
buf \U$15535 ( \21465 , \20208 );
buf \U$15536 ( \21466 , \20208 );
buf \U$15537 ( \21467 , \20208 );
buf \U$15538 ( \21468 , \20208 );
buf \U$15539 ( \21469 , \20208 );
buf \U$15540 ( \21470 , \20208 );
buf \U$15541 ( \21471 , \20208 );
nor \U$15542 ( \21472 , \20195 , \20237 , \20238 , \20239 , \20201 , \20205 , \20208 , \21447 , \21448 , \21449 , \21450 , \21451 , \21452 , \21453 , \21454 , \21455 , \21456 , \21457 , \21458 , \21459 , \21460 , \21461 , \21462 , \21463 , \21464 , \21465 , \21466 , \21467 , \21468 , \21469 , \21470 , \21471 );
and \U$15543 ( \21473 , \8645 , \21472 );
buf \U$15544 ( \21474 , \20208 );
buf \U$15545 ( \21475 , \20208 );
buf \U$15546 ( \21476 , \20208 );
buf \U$15547 ( \21477 , \20208 );
buf \U$15548 ( \21478 , \20208 );
buf \U$15549 ( \21479 , \20208 );
buf \U$15550 ( \21480 , \20208 );
buf \U$15551 ( \21481 , \20208 );
buf \U$15552 ( \21482 , \20208 );
buf \U$15553 ( \21483 , \20208 );
buf \U$15554 ( \21484 , \20208 );
buf \U$15555 ( \21485 , \20208 );
buf \U$15556 ( \21486 , \20208 );
buf \U$15557 ( \21487 , \20208 );
buf \U$15558 ( \21488 , \20208 );
buf \U$15559 ( \21489 , \20208 );
buf \U$15560 ( \21490 , \20208 );
buf \U$15561 ( \21491 , \20208 );
buf \U$15562 ( \21492 , \20208 );
buf \U$15563 ( \21493 , \20208 );
buf \U$15564 ( \21494 , \20208 );
buf \U$15565 ( \21495 , \20208 );
buf \U$15566 ( \21496 , \20208 );
buf \U$15567 ( \21497 , \20208 );
buf \U$15568 ( \21498 , \20208 );
nor \U$15569 ( \21499 , \20236 , \20196 , \20238 , \20239 , \20201 , \20205 , \20208 , \21474 , \21475 , \21476 , \21477 , \21478 , \21479 , \21480 , \21481 , \21482 , \21483 , \21484 , \21485 , \21486 , \21487 , \21488 , \21489 , \21490 , \21491 , \21492 , \21493 , \21494 , \21495 , \21496 , \21497 , \21498 );
and \U$15570 ( \21500 , \8673 , \21499 );
buf \U$15571 ( \21501 , \20208 );
buf \U$15572 ( \21502 , \20208 );
buf \U$15573 ( \21503 , \20208 );
buf \U$15574 ( \21504 , \20208 );
buf \U$15575 ( \21505 , \20208 );
buf \U$15576 ( \21506 , \20208 );
buf \U$15577 ( \21507 , \20208 );
buf \U$15578 ( \21508 , \20208 );
buf \U$15579 ( \21509 , \20208 );
buf \U$15580 ( \21510 , \20208 );
buf \U$15581 ( \21511 , \20208 );
buf \U$15582 ( \21512 , \20208 );
buf \U$15583 ( \21513 , \20208 );
buf \U$15584 ( \21514 , \20208 );
buf \U$15585 ( \21515 , \20208 );
buf \U$15586 ( \21516 , \20208 );
buf \U$15587 ( \21517 , \20208 );
buf \U$15588 ( \21518 , \20208 );
buf \U$15589 ( \21519 , \20208 );
buf \U$15590 ( \21520 , \20208 );
buf \U$15591 ( \21521 , \20208 );
buf \U$15592 ( \21522 , \20208 );
buf \U$15593 ( \21523 , \20208 );
buf \U$15594 ( \21524 , \20208 );
buf \U$15595 ( \21525 , \20208 );
nor \U$15596 ( \21526 , \20195 , \20196 , \20238 , \20239 , \20201 , \20205 , \20208 , \21501 , \21502 , \21503 , \21504 , \21505 , \21506 , \21507 , \21508 , \21509 , \21510 , \21511 , \21512 , \21513 , \21514 , \21515 , \21516 , \21517 , \21518 , \21519 , \21520 , \21521 , \21522 , \21523 , \21524 , \21525 );
and \U$15597 ( \21527 , \8701 , \21526 );
buf \U$15598 ( \21528 , \20208 );
buf \U$15599 ( \21529 , \20208 );
buf \U$15600 ( \21530 , \20208 );
buf \U$15601 ( \21531 , \20208 );
buf \U$15602 ( \21532 , \20208 );
buf \U$15603 ( \21533 , \20208 );
buf \U$15604 ( \21534 , \20208 );
buf \U$15605 ( \21535 , \20208 );
buf \U$15606 ( \21536 , \20208 );
buf \U$15607 ( \21537 , \20208 );
buf \U$15608 ( \21538 , \20208 );
buf \U$15609 ( \21539 , \20208 );
buf \U$15610 ( \21540 , \20208 );
buf \U$15611 ( \21541 , \20208 );
buf \U$15612 ( \21542 , \20208 );
buf \U$15613 ( \21543 , \20208 );
buf \U$15614 ( \21544 , \20208 );
buf \U$15615 ( \21545 , \20208 );
buf \U$15616 ( \21546 , \20208 );
buf \U$15617 ( \21547 , \20208 );
buf \U$15618 ( \21548 , \20208 );
buf \U$15619 ( \21549 , \20208 );
buf \U$15620 ( \21550 , \20208 );
buf \U$15621 ( \21551 , \20208 );
buf \U$15622 ( \21552 , \20208 );
nor \U$15623 ( \21553 , \20236 , \20237 , \20197 , \20239 , \20201 , \20205 , \20208 , \21528 , \21529 , \21530 , \21531 , \21532 , \21533 , \21534 , \21535 , \21536 , \21537 , \21538 , \21539 , \21540 , \21541 , \21542 , \21543 , \21544 , \21545 , \21546 , \21547 , \21548 , \21549 , \21550 , \21551 , \21552 );
and \U$15624 ( \21554 , \8729 , \21553 );
buf \U$15625 ( \21555 , \20208 );
buf \U$15626 ( \21556 , \20208 );
buf \U$15627 ( \21557 , \20208 );
buf \U$15628 ( \21558 , \20208 );
buf \U$15629 ( \21559 , \20208 );
buf \U$15630 ( \21560 , \20208 );
buf \U$15631 ( \21561 , \20208 );
buf \U$15632 ( \21562 , \20208 );
buf \U$15633 ( \21563 , \20208 );
buf \U$15634 ( \21564 , \20208 );
buf \U$15635 ( \21565 , \20208 );
buf \U$15636 ( \21566 , \20208 );
buf \U$15637 ( \21567 , \20208 );
buf \U$15638 ( \21568 , \20208 );
buf \U$15639 ( \21569 , \20208 );
buf \U$15640 ( \21570 , \20208 );
buf \U$15641 ( \21571 , \20208 );
buf \U$15642 ( \21572 , \20208 );
buf \U$15643 ( \21573 , \20208 );
buf \U$15644 ( \21574 , \20208 );
buf \U$15645 ( \21575 , \20208 );
buf \U$15646 ( \21576 , \20208 );
buf \U$15647 ( \21577 , \20208 );
buf \U$15648 ( \21578 , \20208 );
buf \U$15649 ( \21579 , \20208 );
nor \U$15650 ( \21580 , \20195 , \20237 , \20197 , \20239 , \20201 , \20205 , \20208 , \21555 , \21556 , \21557 , \21558 , \21559 , \21560 , \21561 , \21562 , \21563 , \21564 , \21565 , \21566 , \21567 , \21568 , \21569 , \21570 , \21571 , \21572 , \21573 , \21574 , \21575 , \21576 , \21577 , \21578 , \21579 );
and \U$15651 ( \21581 , \8757 , \21580 );
buf \U$15652 ( \21582 , \20208 );
buf \U$15653 ( \21583 , \20208 );
buf \U$15654 ( \21584 , \20208 );
buf \U$15655 ( \21585 , \20208 );
buf \U$15656 ( \21586 , \20208 );
buf \U$15657 ( \21587 , \20208 );
buf \U$15658 ( \21588 , \20208 );
buf \U$15659 ( \21589 , \20208 );
buf \U$15660 ( \21590 , \20208 );
buf \U$15661 ( \21591 , \20208 );
buf \U$15662 ( \21592 , \20208 );
buf \U$15663 ( \21593 , \20208 );
buf \U$15664 ( \21594 , \20208 );
buf \U$15665 ( \21595 , \20208 );
buf \U$15666 ( \21596 , \20208 );
buf \U$15667 ( \21597 , \20208 );
buf \U$15668 ( \21598 , \20208 );
buf \U$15669 ( \21599 , \20208 );
buf \U$15670 ( \21600 , \20208 );
buf \U$15671 ( \21601 , \20208 );
buf \U$15672 ( \21602 , \20208 );
buf \U$15673 ( \21603 , \20208 );
buf \U$15674 ( \21604 , \20208 );
buf \U$15675 ( \21605 , \20208 );
buf \U$15676 ( \21606 , \20208 );
nor \U$15677 ( \21607 , \20236 , \20196 , \20197 , \20239 , \20201 , \20205 , \20208 , \21582 , \21583 , \21584 , \21585 , \21586 , \21587 , \21588 , \21589 , \21590 , \21591 , \21592 , \21593 , \21594 , \21595 , \21596 , \21597 , \21598 , \21599 , \21600 , \21601 , \21602 , \21603 , \21604 , \21605 , \21606 );
and \U$15678 ( \21608 , \8785 , \21607 );
buf \U$15679 ( \21609 , \20208 );
buf \U$15680 ( \21610 , \20208 );
buf \U$15681 ( \21611 , \20208 );
buf \U$15682 ( \21612 , \20208 );
buf \U$15683 ( \21613 , \20208 );
buf \U$15684 ( \21614 , \20208 );
buf \U$15685 ( \21615 , \20208 );
buf \U$15686 ( \21616 , \20208 );
buf \U$15687 ( \21617 , \20208 );
buf \U$15688 ( \21618 , \20208 );
buf \U$15689 ( \21619 , \20208 );
buf \U$15690 ( \21620 , \20208 );
buf \U$15691 ( \21621 , \20208 );
buf \U$15692 ( \21622 , \20208 );
buf \U$15693 ( \21623 , \20208 );
buf \U$15694 ( \21624 , \20208 );
buf \U$15695 ( \21625 , \20208 );
buf \U$15696 ( \21626 , \20208 );
buf \U$15697 ( \21627 , \20208 );
buf \U$15698 ( \21628 , \20208 );
buf \U$15699 ( \21629 , \20208 );
buf \U$15700 ( \21630 , \20208 );
buf \U$15701 ( \21631 , \20208 );
buf \U$15702 ( \21632 , \20208 );
buf \U$15703 ( \21633 , \20208 );
nor \U$15704 ( \21634 , \20195 , \20196 , \20197 , \20239 , \20201 , \20205 , \20208 , \21609 , \21610 , \21611 , \21612 , \21613 , \21614 , \21615 , \21616 , \21617 , \21618 , \21619 , \21620 , \21621 , \21622 , \21623 , \21624 , \21625 , \21626 , \21627 , \21628 , \21629 , \21630 , \21631 , \21632 , \21633 );
and \U$15705 ( \21635 , \8813 , \21634 );
buf \U$15706 ( \21636 , \20208 );
buf \U$15707 ( \21637 , \20208 );
buf \U$15708 ( \21638 , \20208 );
buf \U$15709 ( \21639 , \20208 );
buf \U$15710 ( \21640 , \20208 );
buf \U$15711 ( \21641 , \20208 );
buf \U$15712 ( \21642 , \20208 );
buf \U$15713 ( \21643 , \20208 );
buf \U$15714 ( \21644 , \20208 );
buf \U$15715 ( \21645 , \20208 );
buf \U$15716 ( \21646 , \20208 );
buf \U$15717 ( \21647 , \20208 );
buf \U$15718 ( \21648 , \20208 );
buf \U$15719 ( \21649 , \20208 );
buf \U$15720 ( \21650 , \20208 );
buf \U$15721 ( \21651 , \20208 );
buf \U$15722 ( \21652 , \20208 );
buf \U$15723 ( \21653 , \20208 );
buf \U$15724 ( \21654 , \20208 );
buf \U$15725 ( \21655 , \20208 );
buf \U$15726 ( \21656 , \20208 );
buf \U$15727 ( \21657 , \20208 );
buf \U$15728 ( \21658 , \20208 );
buf \U$15729 ( \21659 , \20208 );
buf \U$15730 ( \21660 , \20208 );
nor \U$15731 ( \21661 , \20236 , \20237 , \20238 , \20198 , \20201 , \20205 , \20208 , \21636 , \21637 , \21638 , \21639 , \21640 , \21641 , \21642 , \21643 , \21644 , \21645 , \21646 , \21647 , \21648 , \21649 , \21650 , \21651 , \21652 , \21653 , \21654 , \21655 , \21656 , \21657 , \21658 , \21659 , \21660 );
and \U$15732 ( \21662 , \8841 , \21661 );
buf \U$15733 ( \21663 , \20208 );
buf \U$15734 ( \21664 , \20208 );
buf \U$15735 ( \21665 , \20208 );
buf \U$15736 ( \21666 , \20208 );
buf \U$15737 ( \21667 , \20208 );
buf \U$15738 ( \21668 , \20208 );
buf \U$15739 ( \21669 , \20208 );
buf \U$15740 ( \21670 , \20208 );
buf \U$15741 ( \21671 , \20208 );
buf \U$15742 ( \21672 , \20208 );
buf \U$15743 ( \21673 , \20208 );
buf \U$15744 ( \21674 , \20208 );
buf \U$15745 ( \21675 , \20208 );
buf \U$15746 ( \21676 , \20208 );
buf \U$15747 ( \21677 , \20208 );
buf \U$15748 ( \21678 , \20208 );
buf \U$15749 ( \21679 , \20208 );
buf \U$15750 ( \21680 , \20208 );
buf \U$15751 ( \21681 , \20208 );
buf \U$15752 ( \21682 , \20208 );
buf \U$15753 ( \21683 , \20208 );
buf \U$15754 ( \21684 , \20208 );
buf \U$15755 ( \21685 , \20208 );
buf \U$15756 ( \21686 , \20208 );
buf \U$15757 ( \21687 , \20208 );
nor \U$15758 ( \21688 , \20195 , \20237 , \20238 , \20198 , \20201 , \20205 , \20208 , \21663 , \21664 , \21665 , \21666 , \21667 , \21668 , \21669 , \21670 , \21671 , \21672 , \21673 , \21674 , \21675 , \21676 , \21677 , \21678 , \21679 , \21680 , \21681 , \21682 , \21683 , \21684 , \21685 , \21686 , \21687 );
and \U$15759 ( \21689 , \8869 , \21688 );
buf \U$15760 ( \21690 , \20208 );
buf \U$15761 ( \21691 , \20208 );
buf \U$15762 ( \21692 , \20208 );
buf \U$15763 ( \21693 , \20208 );
buf \U$15764 ( \21694 , \20208 );
buf \U$15765 ( \21695 , \20208 );
buf \U$15766 ( \21696 , \20208 );
buf \U$15767 ( \21697 , \20208 );
buf \U$15768 ( \21698 , \20208 );
buf \U$15769 ( \21699 , \20208 );
buf \U$15770 ( \21700 , \20208 );
buf \U$15771 ( \21701 , \20208 );
buf \U$15772 ( \21702 , \20208 );
buf \U$15773 ( \21703 , \20208 );
buf \U$15774 ( \21704 , \20208 );
buf \U$15775 ( \21705 , \20208 );
buf \U$15776 ( \21706 , \20208 );
buf \U$15777 ( \21707 , \20208 );
buf \U$15778 ( \21708 , \20208 );
buf \U$15779 ( \21709 , \20208 );
buf \U$15780 ( \21710 , \20208 );
buf \U$15781 ( \21711 , \20208 );
buf \U$15782 ( \21712 , \20208 );
buf \U$15783 ( \21713 , \20208 );
buf \U$15784 ( \21714 , \20208 );
nor \U$15785 ( \21715 , \20236 , \20196 , \20238 , \20198 , \20201 , \20205 , \20208 , \21690 , \21691 , \21692 , \21693 , \21694 , \21695 , \21696 , \21697 , \21698 , \21699 , \21700 , \21701 , \21702 , \21703 , \21704 , \21705 , \21706 , \21707 , \21708 , \21709 , \21710 , \21711 , \21712 , \21713 , \21714 );
and \U$15786 ( \21716 , \8897 , \21715 );
buf \U$15787 ( \21717 , \20208 );
buf \U$15788 ( \21718 , \20208 );
buf \U$15789 ( \21719 , \20208 );
buf \U$15790 ( \21720 , \20208 );
buf \U$15791 ( \21721 , \20208 );
buf \U$15792 ( \21722 , \20208 );
buf \U$15793 ( \21723 , \20208 );
buf \U$15794 ( \21724 , \20208 );
buf \U$15795 ( \21725 , \20208 );
buf \U$15796 ( \21726 , \20208 );
buf \U$15797 ( \21727 , \20208 );
buf \U$15798 ( \21728 , \20208 );
buf \U$15799 ( \21729 , \20208 );
buf \U$15800 ( \21730 , \20208 );
buf \U$15801 ( \21731 , \20208 );
buf \U$15802 ( \21732 , \20208 );
buf \U$15803 ( \21733 , \20208 );
buf \U$15804 ( \21734 , \20208 );
buf \U$15805 ( \21735 , \20208 );
buf \U$15806 ( \21736 , \20208 );
buf \U$15807 ( \21737 , \20208 );
buf \U$15808 ( \21738 , \20208 );
buf \U$15809 ( \21739 , \20208 );
buf \U$15810 ( \21740 , \20208 );
buf \U$15811 ( \21741 , \20208 );
nor \U$15812 ( \21742 , \20195 , \20196 , \20238 , \20198 , \20201 , \20205 , \20208 , \21717 , \21718 , \21719 , \21720 , \21721 , \21722 , \21723 , \21724 , \21725 , \21726 , \21727 , \21728 , \21729 , \21730 , \21731 , \21732 , \21733 , \21734 , \21735 , \21736 , \21737 , \21738 , \21739 , \21740 , \21741 );
and \U$15813 ( \21743 , \8925 , \21742 );
buf \U$15814 ( \21744 , \20208 );
buf \U$15815 ( \21745 , \20208 );
buf \U$15816 ( \21746 , \20208 );
buf \U$15817 ( \21747 , \20208 );
buf \U$15818 ( \21748 , \20208 );
buf \U$15819 ( \21749 , \20208 );
buf \U$15820 ( \21750 , \20208 );
buf \U$15821 ( \21751 , \20208 );
buf \U$15822 ( \21752 , \20208 );
buf \U$15823 ( \21753 , \20208 );
buf \U$15824 ( \21754 , \20208 );
buf \U$15825 ( \21755 , \20208 );
buf \U$15826 ( \21756 , \20208 );
buf \U$15827 ( \21757 , \20208 );
buf \U$15828 ( \21758 , \20208 );
buf \U$15829 ( \21759 , \20208 );
buf \U$15830 ( \21760 , \20208 );
buf \U$15831 ( \21761 , \20208 );
buf \U$15832 ( \21762 , \20208 );
buf \U$15833 ( \21763 , \20208 );
buf \U$15834 ( \21764 , \20208 );
buf \U$15835 ( \21765 , \20208 );
buf \U$15836 ( \21766 , \20208 );
buf \U$15837 ( \21767 , \20208 );
buf \U$15838 ( \21768 , \20208 );
nor \U$15839 ( \21769 , \20236 , \20237 , \20197 , \20198 , \20201 , \20205 , \20208 , \21744 , \21745 , \21746 , \21747 , \21748 , \21749 , \21750 , \21751 , \21752 , \21753 , \21754 , \21755 , \21756 , \21757 , \21758 , \21759 , \21760 , \21761 , \21762 , \21763 , \21764 , \21765 , \21766 , \21767 , \21768 );
and \U$15840 ( \21770 , \8953 , \21769 );
buf \U$15841 ( \21771 , \20208 );
buf \U$15842 ( \21772 , \20208 );
buf \U$15843 ( \21773 , \20208 );
buf \U$15844 ( \21774 , \20208 );
buf \U$15845 ( \21775 , \20208 );
buf \U$15846 ( \21776 , \20208 );
buf \U$15847 ( \21777 , \20208 );
buf \U$15848 ( \21778 , \20208 );
buf \U$15849 ( \21779 , \20208 );
buf \U$15850 ( \21780 , \20208 );
buf \U$15851 ( \21781 , \20208 );
buf \U$15852 ( \21782 , \20208 );
buf \U$15853 ( \21783 , \20208 );
buf \U$15854 ( \21784 , \20208 );
buf \U$15855 ( \21785 , \20208 );
buf \U$15856 ( \21786 , \20208 );
buf \U$15857 ( \21787 , \20208 );
buf \U$15858 ( \21788 , \20208 );
buf \U$15859 ( \21789 , \20208 );
buf \U$15860 ( \21790 , \20208 );
buf \U$15861 ( \21791 , \20208 );
buf \U$15862 ( \21792 , \20208 );
buf \U$15863 ( \21793 , \20208 );
buf \U$15864 ( \21794 , \20208 );
buf \U$15865 ( \21795 , \20208 );
nor \U$15866 ( \21796 , \20195 , \20237 , \20197 , \20198 , \20201 , \20205 , \20208 , \21771 , \21772 , \21773 , \21774 , \21775 , \21776 , \21777 , \21778 , \21779 , \21780 , \21781 , \21782 , \21783 , \21784 , \21785 , \21786 , \21787 , \21788 , \21789 , \21790 , \21791 , \21792 , \21793 , \21794 , \21795 );
and \U$15867 ( \21797 , \8981 , \21796 );
buf \U$15868 ( \21798 , \20208 );
buf \U$15869 ( \21799 , \20208 );
buf \U$15870 ( \21800 , \20208 );
buf \U$15871 ( \21801 , \20208 );
buf \U$15872 ( \21802 , \20208 );
buf \U$15873 ( \21803 , \20208 );
buf \U$15874 ( \21804 , \20208 );
buf \U$15875 ( \21805 , \20208 );
buf \U$15876 ( \21806 , \20208 );
buf \U$15877 ( \21807 , \20208 );
buf \U$15878 ( \21808 , \20208 );
buf \U$15879 ( \21809 , \20208 );
buf \U$15880 ( \21810 , \20208 );
buf \U$15881 ( \21811 , \20208 );
buf \U$15882 ( \21812 , \20208 );
buf \U$15883 ( \21813 , \20208 );
buf \U$15884 ( \21814 , \20208 );
buf \U$15885 ( \21815 , \20208 );
buf \U$15886 ( \21816 , \20208 );
buf \U$15887 ( \21817 , \20208 );
buf \U$15888 ( \21818 , \20208 );
buf \U$15889 ( \21819 , \20208 );
buf \U$15890 ( \21820 , \20208 );
buf \U$15891 ( \21821 , \20208 );
buf \U$15892 ( \21822 , \20208 );
nor \U$15893 ( \21823 , \20236 , \20196 , \20197 , \20198 , \20201 , \20205 , \20208 , \21798 , \21799 , \21800 , \21801 , \21802 , \21803 , \21804 , \21805 , \21806 , \21807 , \21808 , \21809 , \21810 , \21811 , \21812 , \21813 , \21814 , \21815 , \21816 , \21817 , \21818 , \21819 , \21820 , \21821 , \21822 );
and \U$15894 ( \21824 , \9009 , \21823 );
or \U$15895 ( \21825 , \21419 , \21446 , \21473 , \21500 , \21527 , \21554 , \21581 , \21608 , \21635 , \21662 , \21689 , \21716 , \21743 , \21770 , \21797 , \21824 );
buf \U$15896 ( \21826 , \20208 );
not \U$15897 ( \21827 , \21826 );
buf \U$15898 ( \21828 , \20196 );
buf \U$15899 ( \21829 , \20197 );
buf \U$15900 ( \21830 , \20198 );
buf \U$15901 ( \21831 , \20201 );
buf \U$15902 ( \21832 , \20205 );
buf \U$15903 ( \21833 , \20208 );
buf \U$15904 ( \21834 , \20208 );
buf \U$15905 ( \21835 , \20208 );
buf \U$15906 ( \21836 , \20208 );
buf \U$15907 ( \21837 , \20208 );
buf \U$15908 ( \21838 , \20208 );
buf \U$15909 ( \21839 , \20208 );
buf \U$15910 ( \21840 , \20208 );
buf \U$15911 ( \21841 , \20208 );
buf \U$15912 ( \21842 , \20208 );
buf \U$15913 ( \21843 , \20208 );
buf \U$15914 ( \21844 , \20208 );
buf \U$15915 ( \21845 , \20208 );
buf \U$15916 ( \21846 , \20208 );
buf \U$15917 ( \21847 , \20208 );
buf \U$15918 ( \21848 , \20208 );
buf \U$15919 ( \21849 , \20208 );
buf \U$15920 ( \21850 , \20208 );
buf \U$15921 ( \21851 , \20208 );
buf \U$15922 ( \21852 , \20208 );
buf \U$15923 ( \21853 , \20208 );
buf \U$15924 ( \21854 , \20208 );
buf \U$15925 ( \21855 , \20208 );
buf \U$15926 ( \21856 , \20208 );
buf \U$15927 ( \21857 , \20208 );
buf \U$15928 ( \21858 , \20195 );
or \U$15929 ( \21859 , \21828 , \21829 , \21830 , \21831 , \21832 , \21833 , \21834 , \21835 , \21836 , \21837 , \21838 , \21839 , \21840 , \21841 , \21842 , \21843 , \21844 , \21845 , \21846 , \21847 , \21848 , \21849 , \21850 , \21851 , \21852 , \21853 , \21854 , \21855 , \21856 , \21857 , \21858 );
nand \U$15930 ( \21860 , \21827 , \21859 );
buf \U$15931 ( \21861 , \21860 );
buf \U$15932 ( \21862 , \20208 );
not \U$15933 ( \21863 , \21862 );
buf \U$15934 ( \21864 , \20205 );
buf \U$15935 ( \21865 , \20208 );
buf \U$15936 ( \21866 , \20208 );
buf \U$15937 ( \21867 , \20208 );
buf \U$15938 ( \21868 , \20208 );
buf \U$15939 ( \21869 , \20208 );
buf \U$15940 ( \21870 , \20208 );
buf \U$15941 ( \21871 , \20208 );
buf \U$15942 ( \21872 , \20208 );
buf \U$15943 ( \21873 , \20208 );
buf \U$15944 ( \21874 , \20208 );
buf \U$15945 ( \21875 , \20208 );
buf \U$15946 ( \21876 , \20208 );
buf \U$15947 ( \21877 , \20208 );
buf \U$15948 ( \21878 , \20208 );
buf \U$15949 ( \21879 , \20208 );
buf \U$15950 ( \21880 , \20208 );
buf \U$15951 ( \21881 , \20208 );
buf \U$15952 ( \21882 , \20208 );
buf \U$15953 ( \21883 , \20208 );
buf \U$15954 ( \21884 , \20208 );
buf \U$15955 ( \21885 , \20208 );
buf \U$15956 ( \21886 , \20208 );
buf \U$15957 ( \21887 , \20208 );
buf \U$15958 ( \21888 , \20208 );
buf \U$15959 ( \21889 , \20208 );
buf \U$15960 ( \21890 , \20201 );
buf \U$15961 ( \21891 , \20195 );
buf \U$15962 ( \21892 , \20196 );
buf \U$15963 ( \21893 , \20197 );
buf \U$15964 ( \21894 , \20198 );
or \U$15965 ( \21895 , \21891 , \21892 , \21893 , \21894 );
and \U$15966 ( \21896 , \21890 , \21895 );
or \U$15967 ( \21897 , \21864 , \21865 , \21866 , \21867 , \21868 , \21869 , \21870 , \21871 , \21872 , \21873 , \21874 , \21875 , \21876 , \21877 , \21878 , \21879 , \21880 , \21881 , \21882 , \21883 , \21884 , \21885 , \21886 , \21887 , \21888 , \21889 , \21896 );
and \U$15968 ( \21898 , \21863 , \21897 );
buf \U$15969 ( \21899 , \21898 );
or \U$15970 ( \21900 , \21861 , \21899 );
_DC g6c72 ( \21901_nG6c72 , \21825 , \21900 );
buf \U$15971 ( \21902 , \21901_nG6c72 );
xor \U$15972 ( \21903 , \21392 , \21902 );
buf \U$15973 ( \21904 , RIb7af5b8_255);
and \U$15974 ( \21905 , \7207 , \21418 );
and \U$15975 ( \21906 , \7209 , \21445 );
and \U$15976 ( \21907 , \9119 , \21472 );
and \U$15977 ( \21908 , \9121 , \21499 );
and \U$15978 ( \21909 , \9123 , \21526 );
and \U$15979 ( \21910 , \9125 , \21553 );
and \U$15980 ( \21911 , \9127 , \21580 );
and \U$15981 ( \21912 , \9129 , \21607 );
and \U$15982 ( \21913 , \9131 , \21634 );
and \U$15983 ( \21914 , \9133 , \21661 );
and \U$15984 ( \21915 , \9135 , \21688 );
and \U$15985 ( \21916 , \9137 , \21715 );
and \U$15986 ( \21917 , \9139 , \21742 );
and \U$15987 ( \21918 , \9141 , \21769 );
and \U$15988 ( \21919 , \9143 , \21796 );
and \U$15989 ( \21920 , \9145 , \21823 );
or \U$15990 ( \21921 , \21905 , \21906 , \21907 , \21908 , \21909 , \21910 , \21911 , \21912 , \21913 , \21914 , \21915 , \21916 , \21917 , \21918 , \21919 , \21920 );
_DC g6c87 ( \21922_nG6c87 , \21921 , \21900 );
buf \U$15991 ( \21923 , \21922_nG6c87 );
xor \U$15992 ( \21924 , \21904 , \21923 );
or \U$15993 ( \21925 , \21903 , \21924 );
buf \U$15994 ( \21926 , RIb7af540_256);
and \U$15995 ( \21927 , \7217 , \21418 );
and \U$15996 ( \21928 , \7219 , \21445 );
and \U$15997 ( \21929 , \9155 , \21472 );
and \U$15998 ( \21930 , \9157 , \21499 );
and \U$15999 ( \21931 , \9159 , \21526 );
and \U$16000 ( \21932 , \9161 , \21553 );
and \U$16001 ( \21933 , \9163 , \21580 );
and \U$16002 ( \21934 , \9165 , \21607 );
and \U$16003 ( \21935 , \9167 , \21634 );
and \U$16004 ( \21936 , \9169 , \21661 );
and \U$16005 ( \21937 , \9171 , \21688 );
and \U$16006 ( \21938 , \9173 , \21715 );
and \U$16007 ( \21939 , \9175 , \21742 );
and \U$16008 ( \21940 , \9177 , \21769 );
and \U$16009 ( \21941 , \9179 , \21796 );
and \U$16010 ( \21942 , \9181 , \21823 );
or \U$16011 ( \21943 , \21927 , \21928 , \21929 , \21930 , \21931 , \21932 , \21933 , \21934 , \21935 , \21936 , \21937 , \21938 , \21939 , \21940 , \21941 , \21942 );
_DC g6c9d ( \21944_nG6c9d , \21943 , \21900 );
buf \U$16012 ( \21945 , \21944_nG6c9d );
xor \U$16013 ( \21946 , \21926 , \21945 );
or \U$16014 ( \21947 , \21925 , \21946 );
buf \U$16015 ( \21948 , RIb7af4c8_257);
and \U$16016 ( \21949 , \7227 , \21418 );
and \U$16017 ( \21950 , \7229 , \21445 );
and \U$16018 ( \21951 , \9191 , \21472 );
and \U$16019 ( \21952 , \9193 , \21499 );
and \U$16020 ( \21953 , \9195 , \21526 );
and \U$16021 ( \21954 , \9197 , \21553 );
and \U$16022 ( \21955 , \9199 , \21580 );
and \U$16023 ( \21956 , \9201 , \21607 );
and \U$16024 ( \21957 , \9203 , \21634 );
and \U$16025 ( \21958 , \9205 , \21661 );
and \U$16026 ( \21959 , \9207 , \21688 );
and \U$16027 ( \21960 , \9209 , \21715 );
and \U$16028 ( \21961 , \9211 , \21742 );
and \U$16029 ( \21962 , \9213 , \21769 );
and \U$16030 ( \21963 , \9215 , \21796 );
and \U$16031 ( \21964 , \9217 , \21823 );
or \U$16032 ( \21965 , \21949 , \21950 , \21951 , \21952 , \21953 , \21954 , \21955 , \21956 , \21957 , \21958 , \21959 , \21960 , \21961 , \21962 , \21963 , \21964 );
_DC g6cb3 ( \21966_nG6cb3 , \21965 , \21900 );
buf \U$16033 ( \21967 , \21966_nG6cb3 );
xor \U$16034 ( \21968 , \21948 , \21967 );
or \U$16035 ( \21969 , \21947 , \21968 );
buf \U$16036 ( \21970 , RIb7af450_258);
and \U$16037 ( \21971 , \7237 , \21418 );
and \U$16038 ( \21972 , \7239 , \21445 );
and \U$16039 ( \21973 , \9227 , \21472 );
and \U$16040 ( \21974 , \9229 , \21499 );
and \U$16041 ( \21975 , \9231 , \21526 );
and \U$16042 ( \21976 , \9233 , \21553 );
and \U$16043 ( \21977 , \9235 , \21580 );
and \U$16044 ( \21978 , \9237 , \21607 );
and \U$16045 ( \21979 , \9239 , \21634 );
and \U$16046 ( \21980 , \9241 , \21661 );
and \U$16047 ( \21981 , \9243 , \21688 );
and \U$16048 ( \21982 , \9245 , \21715 );
and \U$16049 ( \21983 , \9247 , \21742 );
and \U$16050 ( \21984 , \9249 , \21769 );
and \U$16051 ( \21985 , \9251 , \21796 );
and \U$16052 ( \21986 , \9253 , \21823 );
or \U$16053 ( \21987 , \21971 , \21972 , \21973 , \21974 , \21975 , \21976 , \21977 , \21978 , \21979 , \21980 , \21981 , \21982 , \21983 , \21984 , \21985 , \21986 );
_DC g6cc9 ( \21988_nG6cc9 , \21987 , \21900 );
buf \U$16054 ( \21989 , \21988_nG6cc9 );
xor \U$16055 ( \21990 , \21970 , \21989 );
or \U$16056 ( \21991 , \21969 , \21990 );
buf \U$16057 ( \21992 , RIb7af3d8_259);
and \U$16058 ( \21993 , \7247 , \21418 );
and \U$16059 ( \21994 , \7249 , \21445 );
and \U$16060 ( \21995 , \9263 , \21472 );
and \U$16061 ( \21996 , \9265 , \21499 );
and \U$16062 ( \21997 , \9267 , \21526 );
and \U$16063 ( \21998 , \9269 , \21553 );
and \U$16064 ( \21999 , \9271 , \21580 );
and \U$16065 ( \22000 , \9273 , \21607 );
and \U$16066 ( \22001 , \9275 , \21634 );
and \U$16067 ( \22002 , \9277 , \21661 );
and \U$16068 ( \22003 , \9279 , \21688 );
and \U$16069 ( \22004 , \9281 , \21715 );
and \U$16070 ( \22005 , \9283 , \21742 );
and \U$16071 ( \22006 , \9285 , \21769 );
and \U$16072 ( \22007 , \9287 , \21796 );
and \U$16073 ( \22008 , \9289 , \21823 );
or \U$16074 ( \22009 , \21993 , \21994 , \21995 , \21996 , \21997 , \21998 , \21999 , \22000 , \22001 , \22002 , \22003 , \22004 , \22005 , \22006 , \22007 , \22008 );
_DC g6cdf ( \22010_nG6cdf , \22009 , \21900 );
buf \U$16075 ( \22011 , \22010_nG6cdf );
xor \U$16076 ( \22012 , \21992 , \22011 );
or \U$16077 ( \22013 , \21991 , \22012 );
buf \U$16078 ( \22014 , RIb7a5bf8_260);
and \U$16079 ( \22015 , \7257 , \21418 );
and \U$16080 ( \22016 , \7259 , \21445 );
and \U$16081 ( \22017 , \9299 , \21472 );
and \U$16082 ( \22018 , \9301 , \21499 );
and \U$16083 ( \22019 , \9303 , \21526 );
and \U$16084 ( \22020 , \9305 , \21553 );
and \U$16085 ( \22021 , \9307 , \21580 );
and \U$16086 ( \22022 , \9309 , \21607 );
and \U$16087 ( \22023 , \9311 , \21634 );
and \U$16088 ( \22024 , \9313 , \21661 );
and \U$16089 ( \22025 , \9315 , \21688 );
and \U$16090 ( \22026 , \9317 , \21715 );
and \U$16091 ( \22027 , \9319 , \21742 );
and \U$16092 ( \22028 , \9321 , \21769 );
and \U$16093 ( \22029 , \9323 , \21796 );
and \U$16094 ( \22030 , \9325 , \21823 );
or \U$16095 ( \22031 , \22015 , \22016 , \22017 , \22018 , \22019 , \22020 , \22021 , \22022 , \22023 , \22024 , \22025 , \22026 , \22027 , \22028 , \22029 , \22030 );
_DC g6cf5 ( \22032_nG6cf5 , \22031 , \21900 );
buf \U$16096 ( \22033 , \22032_nG6cf5 );
xor \U$16097 ( \22034 , \22014 , \22033 );
or \U$16098 ( \22035 , \22013 , \22034 );
buf \U$16099 ( \22036 , RIb7a0c48_261);
and \U$16100 ( \22037 , \7267 , \21418 );
and \U$16101 ( \22038 , \7269 , \21445 );
and \U$16102 ( \22039 , \9335 , \21472 );
and \U$16103 ( \22040 , \9337 , \21499 );
and \U$16104 ( \22041 , \9339 , \21526 );
and \U$16105 ( \22042 , \9341 , \21553 );
and \U$16106 ( \22043 , \9343 , \21580 );
and \U$16107 ( \22044 , \9345 , \21607 );
and \U$16108 ( \22045 , \9347 , \21634 );
and \U$16109 ( \22046 , \9349 , \21661 );
and \U$16110 ( \22047 , \9351 , \21688 );
and \U$16111 ( \22048 , \9353 , \21715 );
and \U$16112 ( \22049 , \9355 , \21742 );
and \U$16113 ( \22050 , \9357 , \21769 );
and \U$16114 ( \22051 , \9359 , \21796 );
and \U$16115 ( \22052 , \9361 , \21823 );
or \U$16116 ( \22053 , \22037 , \22038 , \22039 , \22040 , \22041 , \22042 , \22043 , \22044 , \22045 , \22046 , \22047 , \22048 , \22049 , \22050 , \22051 , \22052 );
_DC g6d0b ( \22054_nG6d0b , \22053 , \21900 );
buf \U$16117 ( \22055 , \22054_nG6d0b );
xor \U$16118 ( \22056 , \22036 , \22055 );
or \U$16119 ( \22057 , \22035 , \22056 );
not \U$16120 ( \22058 , \22057 );
buf \U$16121 ( \22059 , \22058 );
and \U$16122 ( \22060 , \21391 , \22059 );
_HMUX g6d12 ( \22061_nG6d12 , \19910_nG64a3 , \20195 , \22060 );
buf \U$16123 ( \22062 , \19931 );
buf \U$16124 ( \22063 , \19928 );
buf \U$16125 ( \22064 , \19913 );
buf \U$16126 ( \22065 , \19916 );
buf \U$16127 ( \22066 , \19920 );
buf \U$16128 ( \22067 , \19924 );
or \U$16129 ( \22068 , \22064 , \22065 , \22066 , \22067 );
and \U$16130 ( \22069 , \22063 , \22068 );
or \U$16131 ( \22070 , \22062 , \22069 );
buf \U$16132 ( \22071 , \22070 );
_HMUX g6d1d ( \22072_nG6d1d , \20194_nG65bf , \22061_nG6d12 , \22071 );
buf \U$16133 ( \22073 , RIe5319e0_6884);
buf \U$16135 ( \22074 , \22073 );
buf \U$16136 ( \22075 , RIe549ef0_6842);
buf \U$16138 ( \22076 , \22075 );
buf \U$16139 ( \22077 , RIe549770_6843);
buf \U$16141 ( \22078 , \22077 );
buf \U$16142 ( \22079 , RIe548ff0_6844);
not \U$16143 ( \22080 , \22079 );
buf \U$16144 ( \22081 , \22080 );
buf \U$16145 ( \22082 , RIea91330_6888);
xor \U$16146 ( \22083 , \22082 , \22079 );
buf \U$16147 ( \22084 , \22083 );
not \U$16148 ( \22085 , \22084 );
and \U$16149 ( \22086 , \22082 , \22079 );
buf \U$16150 ( \22087 , \22086 );
nor \U$16151 ( \22088 , \22074 , \22076 , \22078 , \22081 , \22085 , \22087 );
and \U$16152 ( \22089 , RIe5329d0_6883, \22088 );
not \U$16153 ( \22090 , \22087 );
and \U$16154 ( \22091 , \22074 , \22076 , \22078 , \22081 , \22085 , \22090 );
and \U$16155 ( \22092 , RIeb72150_6905, \22091 );
not \U$16156 ( \22093 , \22074 );
and \U$16157 ( \22094 , \22093 , \22076 , \22078 , \22081 , \22085 , \22090 );
and \U$16158 ( \22095 , RIeab80c0_6897, \22094 );
not \U$16159 ( \22096 , \22076 );
and \U$16160 ( \22097 , \22074 , \22096 , \22078 , \22081 , \22085 , \22090 );
and \U$16161 ( \22098 , RIe5331c8_6882, \22097 );
and \U$16162 ( \22099 , \22093 , \22096 , \22078 , \22081 , \22085 , \22090 );
and \U$16163 ( \22100 , RIe5339c0_6881, \22099 );
not \U$16164 ( \22101 , \22078 );
and \U$16165 ( \22102 , \22074 , \22076 , \22101 , \22081 , \22085 , \22090 );
and \U$16166 ( \22103 , RIeab87c8_6898, \22102 );
and \U$16167 ( \22104 , \22093 , \22076 , \22101 , \22081 , \22085 , \22090 );
and \U$16168 ( \22105 , RIe5341b8_6880, \22104 );
and \U$16169 ( \22106 , \22074 , \22096 , \22101 , \22081 , \22085 , \22090 );
and \U$16170 ( \22107 , RIe5349b0_6879, \22106 );
and \U$16171 ( \22108 , \22093 , \22096 , \22101 , \22081 , \22085 , \22090 );
and \U$16172 ( \22109 , RIea94af8_6890, \22108 );
or \U$16180 ( \22110 , \22089 , \22092 , \22095 , \22098 , \22100 , \22103 , \22105 , \22107 , \22109 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
buf \U$16182 ( \22111 , \22087 );
buf \U$16183 ( \22112 , \22084 );
buf \U$16184 ( \22113 , \22074 );
buf \U$16185 ( \22114 , \22076 );
buf \U$16186 ( \22115 , \22078 );
buf \U$16187 ( \22116 , \22081 );
or \U$16188 ( \22117 , \22113 , \22114 , \22115 , \22116 );
and \U$16189 ( \22118 , \22112 , \22117 );
or \U$16190 ( \22119 , \22111 , \22118 );
buf \U$16191 ( \22120 , \22119 );
or \U$16192 ( \22121 , 1'b0 , \22120 );
_DC g6d52 ( \22122_nG6d52 , \22110 , \22121 );
not \U$16193 ( \22123 , \22122_nG6d52 );
buf \U$16194 ( \22124 , RIb7b9608_246);
and \U$16195 ( \22125 , \7117 , \22088 );
and \U$16196 ( \22126 , \7119 , \22091 );
and \U$16197 ( \22127 , \7864 , \22094 );
and \U$16198 ( \22128 , \7892 , \22097 );
and \U$16199 ( \22129 , \7920 , \22099 );
and \U$16200 ( \22130 , \7948 , \22102 );
and \U$16201 ( \22131 , \7976 , \22104 );
and \U$16202 ( \22132 , \8004 , \22106 );
and \U$16203 ( \22133 , \8032 , \22108 );
or \U$16211 ( \22134 , \22125 , \22126 , \22127 , \22128 , \22129 , \22130 , \22131 , \22132 , \22133 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6d5f ( \22135_nG6d5f , \22134 , \22121 );
buf \U$16212 ( \22136 , \22135_nG6d5f );
xor \U$16213 ( \22137 , \22124 , \22136 );
buf \U$16214 ( \22138 , RIb7b9590_247);
and \U$16215 ( \22139 , \7126 , \22088 );
and \U$16216 ( \22140 , \7128 , \22091 );
and \U$16217 ( \22141 , \8338 , \22094 );
and \U$16218 ( \22142 , \8340 , \22097 );
and \U$16219 ( \22143 , \8342 , \22099 );
and \U$16220 ( \22144 , \8344 , \22102 );
and \U$16221 ( \22145 , \8346 , \22104 );
and \U$16222 ( \22146 , \8348 , \22106 );
and \U$16223 ( \22147 , \8350 , \22108 );
or \U$16231 ( \22148 , \22139 , \22140 , \22141 , \22142 , \22143 , \22144 , \22145 , \22146 , \22147 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6d6d ( \22149_nG6d6d , \22148 , \22121 );
buf \U$16232 ( \22150 , \22149_nG6d6d );
xor \U$16233 ( \22151 , \22138 , \22150 );
or \U$16234 ( \22152 , \22137 , \22151 );
buf \U$16235 ( \22153 , RIb7b9518_248);
and \U$16236 ( \22154 , \7136 , \22088 );
and \U$16237 ( \22155 , \7138 , \22091 );
and \U$16238 ( \22156 , \8374 , \22094 );
and \U$16239 ( \22157 , \8376 , \22097 );
and \U$16240 ( \22158 , \8378 , \22099 );
and \U$16241 ( \22159 , \8380 , \22102 );
and \U$16242 ( \22160 , \8382 , \22104 );
and \U$16243 ( \22161 , \8384 , \22106 );
and \U$16244 ( \22162 , \8386 , \22108 );
or \U$16252 ( \22163 , \22154 , \22155 , \22156 , \22157 , \22158 , \22159 , \22160 , \22161 , \22162 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6d7c ( \22164_nG6d7c , \22163 , \22121 );
buf \U$16253 ( \22165 , \22164_nG6d7c );
xor \U$16254 ( \22166 , \22153 , \22165 );
or \U$16255 ( \22167 , \22152 , \22166 );
buf \U$16256 ( \22168 , RIb7b94a0_249);
and \U$16257 ( \22169 , \7146 , \22088 );
and \U$16258 ( \22170 , \7148 , \22091 );
and \U$16259 ( \22171 , \8410 , \22094 );
and \U$16260 ( \22172 , \8412 , \22097 );
and \U$16261 ( \22173 , \8414 , \22099 );
and \U$16262 ( \22174 , \8416 , \22102 );
and \U$16263 ( \22175 , \8418 , \22104 );
and \U$16264 ( \22176 , \8420 , \22106 );
and \U$16265 ( \22177 , \8422 , \22108 );
or \U$16273 ( \22178 , \22169 , \22170 , \22171 , \22172 , \22173 , \22174 , \22175 , \22176 , \22177 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6d8b ( \22179_nG6d8b , \22178 , \22121 );
buf \U$16274 ( \22180 , \22179_nG6d8b );
xor \U$16275 ( \22181 , \22168 , \22180 );
or \U$16276 ( \22182 , \22167 , \22181 );
buf \U$16277 ( \22183 , RIb7b9428_250);
and \U$16278 ( \22184 , \7156 , \22088 );
and \U$16279 ( \22185 , \7158 , \22091 );
and \U$16280 ( \22186 , \8446 , \22094 );
and \U$16281 ( \22187 , \8448 , \22097 );
and \U$16282 ( \22188 , \8450 , \22099 );
and \U$16283 ( \22189 , \8452 , \22102 );
and \U$16284 ( \22190 , \8454 , \22104 );
and \U$16285 ( \22191 , \8456 , \22106 );
and \U$16286 ( \22192 , \8458 , \22108 );
or \U$16294 ( \22193 , \22184 , \22185 , \22186 , \22187 , \22188 , \22189 , \22190 , \22191 , \22192 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6d9a ( \22194_nG6d9a , \22193 , \22121 );
buf \U$16295 ( \22195 , \22194_nG6d9a );
xor \U$16296 ( \22196 , \22183 , \22195 );
or \U$16297 ( \22197 , \22182 , \22196 );
buf \U$16298 ( \22198 , RIb7b93b0_251);
and \U$16299 ( \22199 , \7166 , \22088 );
and \U$16300 ( \22200 , \7168 , \22091 );
and \U$16301 ( \22201 , \8482 , \22094 );
and \U$16302 ( \22202 , \8484 , \22097 );
and \U$16303 ( \22203 , \8486 , \22099 );
and \U$16304 ( \22204 , \8488 , \22102 );
and \U$16305 ( \22205 , \8490 , \22104 );
and \U$16306 ( \22206 , \8492 , \22106 );
and \U$16307 ( \22207 , \8494 , \22108 );
or \U$16315 ( \22208 , \22199 , \22200 , \22201 , \22202 , \22203 , \22204 , \22205 , \22206 , \22207 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6da9 ( \22209_nG6da9 , \22208 , \22121 );
buf \U$16316 ( \22210 , \22209_nG6da9 );
xor \U$16317 ( \22211 , \22198 , \22210 );
or \U$16318 ( \22212 , \22197 , \22211 );
buf \U$16319 ( \22213 , RIb7af720_252);
and \U$16320 ( \22214 , \7176 , \22088 );
and \U$16321 ( \22215 , \7178 , \22091 );
and \U$16322 ( \22216 , \8518 , \22094 );
and \U$16323 ( \22217 , \8520 , \22097 );
and \U$16324 ( \22218 , \8522 , \22099 );
and \U$16325 ( \22219 , \8524 , \22102 );
and \U$16326 ( \22220 , \8526 , \22104 );
and \U$16327 ( \22221 , \8528 , \22106 );
and \U$16328 ( \22222 , \8530 , \22108 );
or \U$16336 ( \22223 , \22214 , \22215 , \22216 , \22217 , \22218 , \22219 , \22220 , \22221 , \22222 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6db8 ( \22224_nG6db8 , \22223 , \22121 );
buf \U$16337 ( \22225 , \22224_nG6db8 );
xor \U$16338 ( \22226 , \22213 , \22225 );
or \U$16339 ( \22227 , \22212 , \22226 );
buf \U$16340 ( \22228 , RIb7af6a8_253);
and \U$16341 ( \22229 , \7186 , \22088 );
and \U$16342 ( \22230 , \7188 , \22091 );
and \U$16343 ( \22231 , \8554 , \22094 );
and \U$16344 ( \22232 , \8556 , \22097 );
and \U$16345 ( \22233 , \8558 , \22099 );
and \U$16346 ( \22234 , \8560 , \22102 );
and \U$16347 ( \22235 , \8562 , \22104 );
and \U$16348 ( \22236 , \8564 , \22106 );
and \U$16349 ( \22237 , \8566 , \22108 );
or \U$16357 ( \22238 , \22229 , \22230 , \22231 , \22232 , \22233 , \22234 , \22235 , \22236 , \22237 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6dc7 ( \22239_nG6dc7 , \22238 , \22121 );
buf \U$16358 ( \22240 , \22239_nG6dc7 );
xor \U$16359 ( \22241 , \22228 , \22240 );
or \U$16360 ( \22242 , \22227 , \22241 );
not \U$16361 ( \22243 , \22242 );
buf \U$16362 ( \22244 , \22243 );
buf \U$16363 ( \22245 , RIb7af630_254);
and \U$16364 ( \22246 , \7198 , \22088 );
and \U$16365 ( \22247 , \7200 , \22091 );
and \U$16366 ( \22248 , \8645 , \22094 );
and \U$16367 ( \22249 , \8673 , \22097 );
and \U$16368 ( \22250 , \8701 , \22099 );
and \U$16369 ( \22251 , \8729 , \22102 );
and \U$16370 ( \22252 , \8757 , \22104 );
and \U$16371 ( \22253 , \8785 , \22106 );
and \U$16372 ( \22254 , \8813 , \22108 );
or \U$16380 ( \22255 , \22246 , \22247 , \22248 , \22249 , \22250 , \22251 , \22252 , \22253 , \22254 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6dd8 ( \22256_nG6dd8 , \22255 , \22121 );
buf \U$16381 ( \22257 , \22256_nG6dd8 );
xor \U$16382 ( \22258 , \22245 , \22257 );
buf \U$16383 ( \22259 , RIb7af5b8_255);
and \U$16384 ( \22260 , \7207 , \22088 );
and \U$16385 ( \22261 , \7209 , \22091 );
and \U$16386 ( \22262 , \9119 , \22094 );
and \U$16387 ( \22263 , \9121 , \22097 );
and \U$16388 ( \22264 , \9123 , \22099 );
and \U$16389 ( \22265 , \9125 , \22102 );
and \U$16390 ( \22266 , \9127 , \22104 );
and \U$16391 ( \22267 , \9129 , \22106 );
and \U$16392 ( \22268 , \9131 , \22108 );
or \U$16400 ( \22269 , \22260 , \22261 , \22262 , \22263 , \22264 , \22265 , \22266 , \22267 , \22268 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6de6 ( \22270_nG6de6 , \22269 , \22121 );
buf \U$16401 ( \22271 , \22270_nG6de6 );
xor \U$16402 ( \22272 , \22259 , \22271 );
or \U$16403 ( \22273 , \22258 , \22272 );
buf \U$16404 ( \22274 , RIb7af540_256);
and \U$16405 ( \22275 , \7217 , \22088 );
and \U$16406 ( \22276 , \7219 , \22091 );
and \U$16407 ( \22277 , \9155 , \22094 );
and \U$16408 ( \22278 , \9157 , \22097 );
and \U$16409 ( \22279 , \9159 , \22099 );
and \U$16410 ( \22280 , \9161 , \22102 );
and \U$16411 ( \22281 , \9163 , \22104 );
and \U$16412 ( \22282 , \9165 , \22106 );
and \U$16413 ( \22283 , \9167 , \22108 );
or \U$16421 ( \22284 , \22275 , \22276 , \22277 , \22278 , \22279 , \22280 , \22281 , \22282 , \22283 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6df5 ( \22285_nG6df5 , \22284 , \22121 );
buf \U$16422 ( \22286 , \22285_nG6df5 );
xor \U$16423 ( \22287 , \22274 , \22286 );
or \U$16424 ( \22288 , \22273 , \22287 );
buf \U$16425 ( \22289 , RIb7af4c8_257);
and \U$16426 ( \22290 , \7227 , \22088 );
and \U$16427 ( \22291 , \7229 , \22091 );
and \U$16428 ( \22292 , \9191 , \22094 );
and \U$16429 ( \22293 , \9193 , \22097 );
and \U$16430 ( \22294 , \9195 , \22099 );
and \U$16431 ( \22295 , \9197 , \22102 );
and \U$16432 ( \22296 , \9199 , \22104 );
and \U$16433 ( \22297 , \9201 , \22106 );
and \U$16434 ( \22298 , \9203 , \22108 );
or \U$16442 ( \22299 , \22290 , \22291 , \22292 , \22293 , \22294 , \22295 , \22296 , \22297 , \22298 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6e04 ( \22300_nG6e04 , \22299 , \22121 );
buf \U$16443 ( \22301 , \22300_nG6e04 );
xor \U$16444 ( \22302 , \22289 , \22301 );
or \U$16445 ( \22303 , \22288 , \22302 );
buf \U$16446 ( \22304 , RIb7af450_258);
and \U$16447 ( \22305 , \7237 , \22088 );
and \U$16448 ( \22306 , \7239 , \22091 );
and \U$16449 ( \22307 , \9227 , \22094 );
and \U$16450 ( \22308 , \9229 , \22097 );
and \U$16451 ( \22309 , \9231 , \22099 );
and \U$16452 ( \22310 , \9233 , \22102 );
and \U$16453 ( \22311 , \9235 , \22104 );
and \U$16454 ( \22312 , \9237 , \22106 );
and \U$16455 ( \22313 , \9239 , \22108 );
or \U$16463 ( \22314 , \22305 , \22306 , \22307 , \22308 , \22309 , \22310 , \22311 , \22312 , \22313 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6e13 ( \22315_nG6e13 , \22314 , \22121 );
buf \U$16464 ( \22316 , \22315_nG6e13 );
xor \U$16465 ( \22317 , \22304 , \22316 );
or \U$16466 ( \22318 , \22303 , \22317 );
buf \U$16467 ( \22319 , RIb7af3d8_259);
and \U$16468 ( \22320 , \7247 , \22088 );
and \U$16469 ( \22321 , \7249 , \22091 );
and \U$16470 ( \22322 , \9263 , \22094 );
and \U$16471 ( \22323 , \9265 , \22097 );
and \U$16472 ( \22324 , \9267 , \22099 );
and \U$16473 ( \22325 , \9269 , \22102 );
and \U$16474 ( \22326 , \9271 , \22104 );
and \U$16475 ( \22327 , \9273 , \22106 );
and \U$16476 ( \22328 , \9275 , \22108 );
or \U$16484 ( \22329 , \22320 , \22321 , \22322 , \22323 , \22324 , \22325 , \22326 , \22327 , \22328 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6e22 ( \22330_nG6e22 , \22329 , \22121 );
buf \U$16485 ( \22331 , \22330_nG6e22 );
xor \U$16486 ( \22332 , \22319 , \22331 );
or \U$16487 ( \22333 , \22318 , \22332 );
buf \U$16488 ( \22334 , RIb7a5bf8_260);
and \U$16489 ( \22335 , \7257 , \22088 );
and \U$16490 ( \22336 , \7259 , \22091 );
and \U$16491 ( \22337 , \9299 , \22094 );
and \U$16492 ( \22338 , \9301 , \22097 );
and \U$16493 ( \22339 , \9303 , \22099 );
and \U$16494 ( \22340 , \9305 , \22102 );
and \U$16495 ( \22341 , \9307 , \22104 );
and \U$16496 ( \22342 , \9309 , \22106 );
and \U$16497 ( \22343 , \9311 , \22108 );
or \U$16505 ( \22344 , \22335 , \22336 , \22337 , \22338 , \22339 , \22340 , \22341 , \22342 , \22343 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6e31 ( \22345_nG6e31 , \22344 , \22121 );
buf \U$16506 ( \22346 , \22345_nG6e31 );
xor \U$16507 ( \22347 , \22334 , \22346 );
or \U$16508 ( \22348 , \22333 , \22347 );
buf \U$16509 ( \22349 , RIb7a0c48_261);
and \U$16510 ( \22350 , \7267 , \22088 );
and \U$16511 ( \22351 , \7269 , \22091 );
and \U$16512 ( \22352 , \9335 , \22094 );
and \U$16513 ( \22353 , \9337 , \22097 );
and \U$16514 ( \22354 , \9339 , \22099 );
and \U$16515 ( \22355 , \9341 , \22102 );
and \U$16516 ( \22356 , \9343 , \22104 );
and \U$16517 ( \22357 , \9345 , \22106 );
and \U$16518 ( \22358 , \9347 , \22108 );
or \U$16526 ( \22359 , \22350 , \22351 , \22352 , \22353 , \22354 , \22355 , \22356 , \22357 , \22358 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g6e40 ( \22360_nG6e40 , \22359 , \22121 );
buf \U$16527 ( \22361 , \22360_nG6e40 );
xor \U$16528 ( \22362 , \22349 , \22361 );
or \U$16529 ( \22363 , \22348 , \22362 );
not \U$16530 ( \22364 , \22363 );
buf \U$16531 ( \22365 , \22364 );
and \U$16532 ( \22366 , \22244 , \22365 );
and \U$16533 ( \22367 , \22123 , \22366 );
_HMUX g6e48 ( \22368_nG6e48 , \22072_nG6d1d , \22074 , \22367 );
buf \U$16536 ( \22369 , \22074 );
buf \U$16539 ( \22370 , \22076 );
buf \U$16542 ( \22371 , \22078 );
buf \U$16545 ( \22372 , \22081 );
buf \U$16546 ( \22373 , \22084 );
not \U$16547 ( \22374 , \22373 );
buf \U$16548 ( \22375 , \22374 );
not \U$16549 ( \22376 , \22375 );
buf \U$16550 ( \22377 , \22087 );
xnor \U$16551 ( \22378 , \22377 , \22373 );
buf \U$16552 ( \22379 , \22378 );
or \U$16553 ( \22380 , \22377 , \22373 );
not \U$16554 ( \22381 , \22380 );
buf \U$16555 ( \22382 , \22381 );
buf \U$16556 ( \22383 , \22382 );
buf \U$16557 ( \22384 , \22382 );
buf \U$16558 ( \22385 , \22382 );
buf \U$16559 ( \22386 , \22382 );
buf \U$16560 ( \22387 , \22382 );
buf \U$16561 ( \22388 , \22382 );
buf \U$16562 ( \22389 , \22382 );
buf \U$16563 ( \22390 , \22382 );
buf \U$16564 ( \22391 , \22382 );
buf \U$16565 ( \22392 , \22382 );
buf \U$16566 ( \22393 , \22382 );
buf \U$16567 ( \22394 , \22382 );
buf \U$16568 ( \22395 , \22382 );
buf \U$16569 ( \22396 , \22382 );
buf \U$16570 ( \22397 , \22382 );
buf \U$16571 ( \22398 , \22382 );
buf \U$16572 ( \22399 , \22382 );
buf \U$16573 ( \22400 , \22382 );
buf \U$16574 ( \22401 , \22382 );
buf \U$16575 ( \22402 , \22382 );
buf \U$16576 ( \22403 , \22382 );
buf \U$16577 ( \22404 , \22382 );
buf \U$16578 ( \22405 , \22382 );
buf \U$16579 ( \22406 , \22382 );
buf \U$16580 ( \22407 , \22382 );
nor \U$16581 ( \22408 , \22369 , \22370 , \22371 , \22372 , \22376 , \22379 , \22382 , \22383 , \22384 , \22385 , \22386 , \22387 , \22388 , \22389 , \22390 , \22391 , \22392 , \22393 , \22394 , \22395 , \22396 , \22397 , \22398 , \22399 , \22400 , \22401 , \22402 , \22403 , \22404 , \22405 , \22406 , \22407 );
and \U$16582 ( \22409 , RIe5329d0_6883, \22408 );
not \U$16583 ( \22410 , \22369 );
not \U$16584 ( \22411 , \22370 );
not \U$16585 ( \22412 , \22371 );
not \U$16586 ( \22413 , \22372 );
buf \U$16587 ( \22414 , \22382 );
buf \U$16588 ( \22415 , \22382 );
buf \U$16589 ( \22416 , \22382 );
buf \U$16590 ( \22417 , \22382 );
buf \U$16591 ( \22418 , \22382 );
buf \U$16592 ( \22419 , \22382 );
buf \U$16593 ( \22420 , \22382 );
buf \U$16594 ( \22421 , \22382 );
buf \U$16595 ( \22422 , \22382 );
buf \U$16596 ( \22423 , \22382 );
buf \U$16597 ( \22424 , \22382 );
buf \U$16598 ( \22425 , \22382 );
buf \U$16599 ( \22426 , \22382 );
buf \U$16600 ( \22427 , \22382 );
buf \U$16601 ( \22428 , \22382 );
buf \U$16602 ( \22429 , \22382 );
buf \U$16603 ( \22430 , \22382 );
buf \U$16604 ( \22431 , \22382 );
buf \U$16605 ( \22432 , \22382 );
buf \U$16606 ( \22433 , \22382 );
buf \U$16607 ( \22434 , \22382 );
buf \U$16608 ( \22435 , \22382 );
buf \U$16609 ( \22436 , \22382 );
buf \U$16610 ( \22437 , \22382 );
buf \U$16611 ( \22438 , \22382 );
nor \U$16612 ( \22439 , \22410 , \22411 , \22412 , \22413 , \22375 , \22379 , \22382 , \22414 , \22415 , \22416 , \22417 , \22418 , \22419 , \22420 , \22421 , \22422 , \22423 , \22424 , \22425 , \22426 , \22427 , \22428 , \22429 , \22430 , \22431 , \22432 , \22433 , \22434 , \22435 , \22436 , \22437 , \22438 );
and \U$16613 ( \22440 , RIeb72150_6905, \22439 );
buf \U$16614 ( \22441 , \22382 );
buf \U$16615 ( \22442 , \22382 );
buf \U$16616 ( \22443 , \22382 );
buf \U$16617 ( \22444 , \22382 );
buf \U$16618 ( \22445 , \22382 );
buf \U$16619 ( \22446 , \22382 );
buf \U$16620 ( \22447 , \22382 );
buf \U$16621 ( \22448 , \22382 );
buf \U$16622 ( \22449 , \22382 );
buf \U$16623 ( \22450 , \22382 );
buf \U$16624 ( \22451 , \22382 );
buf \U$16625 ( \22452 , \22382 );
buf \U$16626 ( \22453 , \22382 );
buf \U$16627 ( \22454 , \22382 );
buf \U$16628 ( \22455 , \22382 );
buf \U$16629 ( \22456 , \22382 );
buf \U$16630 ( \22457 , \22382 );
buf \U$16631 ( \22458 , \22382 );
buf \U$16632 ( \22459 , \22382 );
buf \U$16633 ( \22460 , \22382 );
buf \U$16634 ( \22461 , \22382 );
buf \U$16635 ( \22462 , \22382 );
buf \U$16636 ( \22463 , \22382 );
buf \U$16637 ( \22464 , \22382 );
buf \U$16638 ( \22465 , \22382 );
nor \U$16639 ( \22466 , \22369 , \22411 , \22412 , \22413 , \22375 , \22379 , \22382 , \22441 , \22442 , \22443 , \22444 , \22445 , \22446 , \22447 , \22448 , \22449 , \22450 , \22451 , \22452 , \22453 , \22454 , \22455 , \22456 , \22457 , \22458 , \22459 , \22460 , \22461 , \22462 , \22463 , \22464 , \22465 );
and \U$16640 ( \22467 , RIeab80c0_6897, \22466 );
buf \U$16641 ( \22468 , \22382 );
buf \U$16642 ( \22469 , \22382 );
buf \U$16643 ( \22470 , \22382 );
buf \U$16644 ( \22471 , \22382 );
buf \U$16645 ( \22472 , \22382 );
buf \U$16646 ( \22473 , \22382 );
buf \U$16647 ( \22474 , \22382 );
buf \U$16648 ( \22475 , \22382 );
buf \U$16649 ( \22476 , \22382 );
buf \U$16650 ( \22477 , \22382 );
buf \U$16651 ( \22478 , \22382 );
buf \U$16652 ( \22479 , \22382 );
buf \U$16653 ( \22480 , \22382 );
buf \U$16654 ( \22481 , \22382 );
buf \U$16655 ( \22482 , \22382 );
buf \U$16656 ( \22483 , \22382 );
buf \U$16657 ( \22484 , \22382 );
buf \U$16658 ( \22485 , \22382 );
buf \U$16659 ( \22486 , \22382 );
buf \U$16660 ( \22487 , \22382 );
buf \U$16661 ( \22488 , \22382 );
buf \U$16662 ( \22489 , \22382 );
buf \U$16663 ( \22490 , \22382 );
buf \U$16664 ( \22491 , \22382 );
buf \U$16665 ( \22492 , \22382 );
nor \U$16666 ( \22493 , \22410 , \22370 , \22412 , \22413 , \22375 , \22379 , \22382 , \22468 , \22469 , \22470 , \22471 , \22472 , \22473 , \22474 , \22475 , \22476 , \22477 , \22478 , \22479 , \22480 , \22481 , \22482 , \22483 , \22484 , \22485 , \22486 , \22487 , \22488 , \22489 , \22490 , \22491 , \22492 );
and \U$16667 ( \22494 , RIe5331c8_6882, \22493 );
buf \U$16668 ( \22495 , \22382 );
buf \U$16669 ( \22496 , \22382 );
buf \U$16670 ( \22497 , \22382 );
buf \U$16671 ( \22498 , \22382 );
buf \U$16672 ( \22499 , \22382 );
buf \U$16673 ( \22500 , \22382 );
buf \U$16674 ( \22501 , \22382 );
buf \U$16675 ( \22502 , \22382 );
buf \U$16676 ( \22503 , \22382 );
buf \U$16677 ( \22504 , \22382 );
buf \U$16678 ( \22505 , \22382 );
buf \U$16679 ( \22506 , \22382 );
buf \U$16680 ( \22507 , \22382 );
buf \U$16681 ( \22508 , \22382 );
buf \U$16682 ( \22509 , \22382 );
buf \U$16683 ( \22510 , \22382 );
buf \U$16684 ( \22511 , \22382 );
buf \U$16685 ( \22512 , \22382 );
buf \U$16686 ( \22513 , \22382 );
buf \U$16687 ( \22514 , \22382 );
buf \U$16688 ( \22515 , \22382 );
buf \U$16689 ( \22516 , \22382 );
buf \U$16690 ( \22517 , \22382 );
buf \U$16691 ( \22518 , \22382 );
buf \U$16692 ( \22519 , \22382 );
nor \U$16693 ( \22520 , \22369 , \22370 , \22412 , \22413 , \22375 , \22379 , \22382 , \22495 , \22496 , \22497 , \22498 , \22499 , \22500 , \22501 , \22502 , \22503 , \22504 , \22505 , \22506 , \22507 , \22508 , \22509 , \22510 , \22511 , \22512 , \22513 , \22514 , \22515 , \22516 , \22517 , \22518 , \22519 );
and \U$16694 ( \22521 , RIe5339c0_6881, \22520 );
buf \U$16695 ( \22522 , \22382 );
buf \U$16696 ( \22523 , \22382 );
buf \U$16697 ( \22524 , \22382 );
buf \U$16698 ( \22525 , \22382 );
buf \U$16699 ( \22526 , \22382 );
buf \U$16700 ( \22527 , \22382 );
buf \U$16701 ( \22528 , \22382 );
buf \U$16702 ( \22529 , \22382 );
buf \U$16703 ( \22530 , \22382 );
buf \U$16704 ( \22531 , \22382 );
buf \U$16705 ( \22532 , \22382 );
buf \U$16706 ( \22533 , \22382 );
buf \U$16707 ( \22534 , \22382 );
buf \U$16708 ( \22535 , \22382 );
buf \U$16709 ( \22536 , \22382 );
buf \U$16710 ( \22537 , \22382 );
buf \U$16711 ( \22538 , \22382 );
buf \U$16712 ( \22539 , \22382 );
buf \U$16713 ( \22540 , \22382 );
buf \U$16714 ( \22541 , \22382 );
buf \U$16715 ( \22542 , \22382 );
buf \U$16716 ( \22543 , \22382 );
buf \U$16717 ( \22544 , \22382 );
buf \U$16718 ( \22545 , \22382 );
buf \U$16719 ( \22546 , \22382 );
nor \U$16720 ( \22547 , \22410 , \22411 , \22371 , \22413 , \22375 , \22379 , \22382 , \22522 , \22523 , \22524 , \22525 , \22526 , \22527 , \22528 , \22529 , \22530 , \22531 , \22532 , \22533 , \22534 , \22535 , \22536 , \22537 , \22538 , \22539 , \22540 , \22541 , \22542 , \22543 , \22544 , \22545 , \22546 );
and \U$16721 ( \22548 , RIeab87c8_6898, \22547 );
buf \U$16722 ( \22549 , \22382 );
buf \U$16723 ( \22550 , \22382 );
buf \U$16724 ( \22551 , \22382 );
buf \U$16725 ( \22552 , \22382 );
buf \U$16726 ( \22553 , \22382 );
buf \U$16727 ( \22554 , \22382 );
buf \U$16728 ( \22555 , \22382 );
buf \U$16729 ( \22556 , \22382 );
buf \U$16730 ( \22557 , \22382 );
buf \U$16731 ( \22558 , \22382 );
buf \U$16732 ( \22559 , \22382 );
buf \U$16733 ( \22560 , \22382 );
buf \U$16734 ( \22561 , \22382 );
buf \U$16735 ( \22562 , \22382 );
buf \U$16736 ( \22563 , \22382 );
buf \U$16737 ( \22564 , \22382 );
buf \U$16738 ( \22565 , \22382 );
buf \U$16739 ( \22566 , \22382 );
buf \U$16740 ( \22567 , \22382 );
buf \U$16741 ( \22568 , \22382 );
buf \U$16742 ( \22569 , \22382 );
buf \U$16743 ( \22570 , \22382 );
buf \U$16744 ( \22571 , \22382 );
buf \U$16745 ( \22572 , \22382 );
buf \U$16746 ( \22573 , \22382 );
nor \U$16747 ( \22574 , \22369 , \22411 , \22371 , \22413 , \22375 , \22379 , \22382 , \22549 , \22550 , \22551 , \22552 , \22553 , \22554 , \22555 , \22556 , \22557 , \22558 , \22559 , \22560 , \22561 , \22562 , \22563 , \22564 , \22565 , \22566 , \22567 , \22568 , \22569 , \22570 , \22571 , \22572 , \22573 );
and \U$16748 ( \22575 , RIe5341b8_6880, \22574 );
buf \U$16749 ( \22576 , \22382 );
buf \U$16750 ( \22577 , \22382 );
buf \U$16751 ( \22578 , \22382 );
buf \U$16752 ( \22579 , \22382 );
buf \U$16753 ( \22580 , \22382 );
buf \U$16754 ( \22581 , \22382 );
buf \U$16755 ( \22582 , \22382 );
buf \U$16756 ( \22583 , \22382 );
buf \U$16757 ( \22584 , \22382 );
buf \U$16758 ( \22585 , \22382 );
buf \U$16759 ( \22586 , \22382 );
buf \U$16760 ( \22587 , \22382 );
buf \U$16761 ( \22588 , \22382 );
buf \U$16762 ( \22589 , \22382 );
buf \U$16763 ( \22590 , \22382 );
buf \U$16764 ( \22591 , \22382 );
buf \U$16765 ( \22592 , \22382 );
buf \U$16766 ( \22593 , \22382 );
buf \U$16767 ( \22594 , \22382 );
buf \U$16768 ( \22595 , \22382 );
buf \U$16769 ( \22596 , \22382 );
buf \U$16770 ( \22597 , \22382 );
buf \U$16771 ( \22598 , \22382 );
buf \U$16772 ( \22599 , \22382 );
buf \U$16773 ( \22600 , \22382 );
nor \U$16774 ( \22601 , \22410 , \22370 , \22371 , \22413 , \22375 , \22379 , \22382 , \22576 , \22577 , \22578 , \22579 , \22580 , \22581 , \22582 , \22583 , \22584 , \22585 , \22586 , \22587 , \22588 , \22589 , \22590 , \22591 , \22592 , \22593 , \22594 , \22595 , \22596 , \22597 , \22598 , \22599 , \22600 );
and \U$16775 ( \22602 , RIe5349b0_6879, \22601 );
buf \U$16776 ( \22603 , \22382 );
buf \U$16777 ( \22604 , \22382 );
buf \U$16778 ( \22605 , \22382 );
buf \U$16779 ( \22606 , \22382 );
buf \U$16780 ( \22607 , \22382 );
buf \U$16781 ( \22608 , \22382 );
buf \U$16782 ( \22609 , \22382 );
buf \U$16783 ( \22610 , \22382 );
buf \U$16784 ( \22611 , \22382 );
buf \U$16785 ( \22612 , \22382 );
buf \U$16786 ( \22613 , \22382 );
buf \U$16787 ( \22614 , \22382 );
buf \U$16788 ( \22615 , \22382 );
buf \U$16789 ( \22616 , \22382 );
buf \U$16790 ( \22617 , \22382 );
buf \U$16791 ( \22618 , \22382 );
buf \U$16792 ( \22619 , \22382 );
buf \U$16793 ( \22620 , \22382 );
buf \U$16794 ( \22621 , \22382 );
buf \U$16795 ( \22622 , \22382 );
buf \U$16796 ( \22623 , \22382 );
buf \U$16797 ( \22624 , \22382 );
buf \U$16798 ( \22625 , \22382 );
buf \U$16799 ( \22626 , \22382 );
buf \U$16800 ( \22627 , \22382 );
nor \U$16801 ( \22628 , \22369 , \22370 , \22371 , \22413 , \22375 , \22379 , \22382 , \22603 , \22604 , \22605 , \22606 , \22607 , \22608 , \22609 , \22610 , \22611 , \22612 , \22613 , \22614 , \22615 , \22616 , \22617 , \22618 , \22619 , \22620 , \22621 , \22622 , \22623 , \22624 , \22625 , \22626 , \22627 );
and \U$16802 ( \22629 , RIea94af8_6890, \22628 );
buf \U$16803 ( \22630 , \22382 );
buf \U$16804 ( \22631 , \22382 );
buf \U$16805 ( \22632 , \22382 );
buf \U$16806 ( \22633 , \22382 );
buf \U$16807 ( \22634 , \22382 );
buf \U$16808 ( \22635 , \22382 );
buf \U$16809 ( \22636 , \22382 );
buf \U$16810 ( \22637 , \22382 );
buf \U$16811 ( \22638 , \22382 );
buf \U$16812 ( \22639 , \22382 );
buf \U$16813 ( \22640 , \22382 );
buf \U$16814 ( \22641 , \22382 );
buf \U$16815 ( \22642 , \22382 );
buf \U$16816 ( \22643 , \22382 );
buf \U$16817 ( \22644 , \22382 );
buf \U$16818 ( \22645 , \22382 );
buf \U$16819 ( \22646 , \22382 );
buf \U$16820 ( \22647 , \22382 );
buf \U$16821 ( \22648 , \22382 );
buf \U$16822 ( \22649 , \22382 );
buf \U$16823 ( \22650 , \22382 );
buf \U$16824 ( \22651 , \22382 );
buf \U$16825 ( \22652 , \22382 );
buf \U$16826 ( \22653 , \22382 );
buf \U$16827 ( \22654 , \22382 );
nor \U$16828 ( \22655 , \22410 , \22411 , \22412 , \22372 , \22375 , \22379 , \22382 , \22630 , \22631 , \22632 , \22633 , \22634 , \22635 , \22636 , \22637 , \22638 , \22639 , \22640 , \22641 , \22642 , \22643 , \22644 , \22645 , \22646 , \22647 , \22648 , \22649 , \22650 , \22651 , \22652 , \22653 , \22654 );
and \U$16829 ( \22656 , RIe5351a8_6878, \22655 );
buf \U$16830 ( \22657 , \22382 );
buf \U$16831 ( \22658 , \22382 );
buf \U$16832 ( \22659 , \22382 );
buf \U$16833 ( \22660 , \22382 );
buf \U$16834 ( \22661 , \22382 );
buf \U$16835 ( \22662 , \22382 );
buf \U$16836 ( \22663 , \22382 );
buf \U$16837 ( \22664 , \22382 );
buf \U$16838 ( \22665 , \22382 );
buf \U$16839 ( \22666 , \22382 );
buf \U$16840 ( \22667 , \22382 );
buf \U$16841 ( \22668 , \22382 );
buf \U$16842 ( \22669 , \22382 );
buf \U$16843 ( \22670 , \22382 );
buf \U$16844 ( \22671 , \22382 );
buf \U$16845 ( \22672 , \22382 );
buf \U$16846 ( \22673 , \22382 );
buf \U$16847 ( \22674 , \22382 );
buf \U$16848 ( \22675 , \22382 );
buf \U$16849 ( \22676 , \22382 );
buf \U$16850 ( \22677 , \22382 );
buf \U$16851 ( \22678 , \22382 );
buf \U$16852 ( \22679 , \22382 );
buf \U$16853 ( \22680 , \22382 );
buf \U$16854 ( \22681 , \22382 );
nor \U$16855 ( \22682 , \22369 , \22411 , \22412 , \22372 , \22375 , \22379 , \22382 , \22657 , \22658 , \22659 , \22660 , \22661 , \22662 , \22663 , \22664 , \22665 , \22666 , \22667 , \22668 , \22669 , \22670 , \22671 , \22672 , \22673 , \22674 , \22675 , \22676 , \22677 , \22678 , \22679 , \22680 , \22681 );
and \U$16856 ( \22683 , RIe5359a0_6877, \22682 );
buf \U$16857 ( \22684 , \22382 );
buf \U$16858 ( \22685 , \22382 );
buf \U$16859 ( \22686 , \22382 );
buf \U$16860 ( \22687 , \22382 );
buf \U$16861 ( \22688 , \22382 );
buf \U$16862 ( \22689 , \22382 );
buf \U$16863 ( \22690 , \22382 );
buf \U$16864 ( \22691 , \22382 );
buf \U$16865 ( \22692 , \22382 );
buf \U$16866 ( \22693 , \22382 );
buf \U$16867 ( \22694 , \22382 );
buf \U$16868 ( \22695 , \22382 );
buf \U$16869 ( \22696 , \22382 );
buf \U$16870 ( \22697 , \22382 );
buf \U$16871 ( \22698 , \22382 );
buf \U$16872 ( \22699 , \22382 );
buf \U$16873 ( \22700 , \22382 );
buf \U$16874 ( \22701 , \22382 );
buf \U$16875 ( \22702 , \22382 );
buf \U$16876 ( \22703 , \22382 );
buf \U$16877 ( \22704 , \22382 );
buf \U$16878 ( \22705 , \22382 );
buf \U$16879 ( \22706 , \22382 );
buf \U$16880 ( \22707 , \22382 );
buf \U$16881 ( \22708 , \22382 );
nor \U$16882 ( \22709 , \22410 , \22370 , \22412 , \22372 , \22375 , \22379 , \22382 , \22684 , \22685 , \22686 , \22687 , \22688 , \22689 , \22690 , \22691 , \22692 , \22693 , \22694 , \22695 , \22696 , \22697 , \22698 , \22699 , \22700 , \22701 , \22702 , \22703 , \22704 , \22705 , \22706 , \22707 , \22708 );
and \U$16883 ( \22710 , RIeab78c8_6895, \22709 );
buf \U$16884 ( \22711 , \22382 );
buf \U$16885 ( \22712 , \22382 );
buf \U$16886 ( \22713 , \22382 );
buf \U$16887 ( \22714 , \22382 );
buf \U$16888 ( \22715 , \22382 );
buf \U$16889 ( \22716 , \22382 );
buf \U$16890 ( \22717 , \22382 );
buf \U$16891 ( \22718 , \22382 );
buf \U$16892 ( \22719 , \22382 );
buf \U$16893 ( \22720 , \22382 );
buf \U$16894 ( \22721 , \22382 );
buf \U$16895 ( \22722 , \22382 );
buf \U$16896 ( \22723 , \22382 );
buf \U$16897 ( \22724 , \22382 );
buf \U$16898 ( \22725 , \22382 );
buf \U$16899 ( \22726 , \22382 );
buf \U$16900 ( \22727 , \22382 );
buf \U$16901 ( \22728 , \22382 );
buf \U$16902 ( \22729 , \22382 );
buf \U$16903 ( \22730 , \22382 );
buf \U$16904 ( \22731 , \22382 );
buf \U$16905 ( \22732 , \22382 );
buf \U$16906 ( \22733 , \22382 );
buf \U$16907 ( \22734 , \22382 );
buf \U$16908 ( \22735 , \22382 );
nor \U$16909 ( \22736 , \22369 , \22370 , \22412 , \22372 , \22375 , \22379 , \22382 , \22711 , \22712 , \22713 , \22714 , \22715 , \22716 , \22717 , \22718 , \22719 , \22720 , \22721 , \22722 , \22723 , \22724 , \22725 , \22726 , \22727 , \22728 , \22729 , \22730 , \22731 , \22732 , \22733 , \22734 , \22735 );
and \U$16910 ( \22737 , RIeab7d00_6896, \22736 );
buf \U$16911 ( \22738 , \22382 );
buf \U$16912 ( \22739 , \22382 );
buf \U$16913 ( \22740 , \22382 );
buf \U$16914 ( \22741 , \22382 );
buf \U$16915 ( \22742 , \22382 );
buf \U$16916 ( \22743 , \22382 );
buf \U$16917 ( \22744 , \22382 );
buf \U$16918 ( \22745 , \22382 );
buf \U$16919 ( \22746 , \22382 );
buf \U$16920 ( \22747 , \22382 );
buf \U$16921 ( \22748 , \22382 );
buf \U$16922 ( \22749 , \22382 );
buf \U$16923 ( \22750 , \22382 );
buf \U$16924 ( \22751 , \22382 );
buf \U$16925 ( \22752 , \22382 );
buf \U$16926 ( \22753 , \22382 );
buf \U$16927 ( \22754 , \22382 );
buf \U$16928 ( \22755 , \22382 );
buf \U$16929 ( \22756 , \22382 );
buf \U$16930 ( \22757 , \22382 );
buf \U$16931 ( \22758 , \22382 );
buf \U$16932 ( \22759 , \22382 );
buf \U$16933 ( \22760 , \22382 );
buf \U$16934 ( \22761 , \22382 );
buf \U$16935 ( \22762 , \22382 );
nor \U$16936 ( \22763 , \22410 , \22411 , \22371 , \22372 , \22375 , \22379 , \22382 , \22738 , \22739 , \22740 , \22741 , \22742 , \22743 , \22744 , \22745 , \22746 , \22747 , \22748 , \22749 , \22750 , \22751 , \22752 , \22753 , \22754 , \22755 , \22756 , \22757 , \22758 , \22759 , \22760 , \22761 , \22762 );
and \U$16937 ( \22764 , RIeacfa18_6902, \22763 );
buf \U$16938 ( \22765 , \22382 );
buf \U$16939 ( \22766 , \22382 );
buf \U$16940 ( \22767 , \22382 );
buf \U$16941 ( \22768 , \22382 );
buf \U$16942 ( \22769 , \22382 );
buf \U$16943 ( \22770 , \22382 );
buf \U$16944 ( \22771 , \22382 );
buf \U$16945 ( \22772 , \22382 );
buf \U$16946 ( \22773 , \22382 );
buf \U$16947 ( \22774 , \22382 );
buf \U$16948 ( \22775 , \22382 );
buf \U$16949 ( \22776 , \22382 );
buf \U$16950 ( \22777 , \22382 );
buf \U$16951 ( \22778 , \22382 );
buf \U$16952 ( \22779 , \22382 );
buf \U$16953 ( \22780 , \22382 );
buf \U$16954 ( \22781 , \22382 );
buf \U$16955 ( \22782 , \22382 );
buf \U$16956 ( \22783 , \22382 );
buf \U$16957 ( \22784 , \22382 );
buf \U$16958 ( \22785 , \22382 );
buf \U$16959 ( \22786 , \22382 );
buf \U$16960 ( \22787 , \22382 );
buf \U$16961 ( \22788 , \22382 );
buf \U$16962 ( \22789 , \22382 );
nor \U$16963 ( \22790 , \22369 , \22411 , \22371 , \22372 , \22375 , \22379 , \22382 , \22765 , \22766 , \22767 , \22768 , \22769 , \22770 , \22771 , \22772 , \22773 , \22774 , \22775 , \22776 , \22777 , \22778 , \22779 , \22780 , \22781 , \22782 , \22783 , \22784 , \22785 , \22786 , \22787 , \22788 , \22789 );
and \U$16964 ( \22791 , RIeab6518_6891, \22790 );
buf \U$16965 ( \22792 , \22382 );
buf \U$16966 ( \22793 , \22382 );
buf \U$16967 ( \22794 , \22382 );
buf \U$16968 ( \22795 , \22382 );
buf \U$16969 ( \22796 , \22382 );
buf \U$16970 ( \22797 , \22382 );
buf \U$16971 ( \22798 , \22382 );
buf \U$16972 ( \22799 , \22382 );
buf \U$16973 ( \22800 , \22382 );
buf \U$16974 ( \22801 , \22382 );
buf \U$16975 ( \22802 , \22382 );
buf \U$16976 ( \22803 , \22382 );
buf \U$16977 ( \22804 , \22382 );
buf \U$16978 ( \22805 , \22382 );
buf \U$16979 ( \22806 , \22382 );
buf \U$16980 ( \22807 , \22382 );
buf \U$16981 ( \22808 , \22382 );
buf \U$16982 ( \22809 , \22382 );
buf \U$16983 ( \22810 , \22382 );
buf \U$16984 ( \22811 , \22382 );
buf \U$16985 ( \22812 , \22382 );
buf \U$16986 ( \22813 , \22382 );
buf \U$16987 ( \22814 , \22382 );
buf \U$16988 ( \22815 , \22382 );
buf \U$16989 ( \22816 , \22382 );
nor \U$16990 ( \22817 , \22410 , \22370 , \22371 , \22372 , \22375 , \22379 , \22382 , \22792 , \22793 , \22794 , \22795 , \22796 , \22797 , \22798 , \22799 , \22800 , \22801 , \22802 , \22803 , \22804 , \22805 , \22806 , \22807 , \22808 , \22809 , \22810 , \22811 , \22812 , \22813 , \22814 , \22815 , \22816 );
and \U$16991 ( \22818 , RIeb352c8_6904, \22817 );
or \U$16992 ( \22819 , \22409 , \22440 , \22467 , \22494 , \22521 , \22548 , \22575 , \22602 , \22629 , \22656 , \22683 , \22710 , \22737 , \22764 , \22791 , \22818 );
buf \U$16993 ( \22820 , \22382 );
not \U$16994 ( \22821 , \22820 );
buf \U$16995 ( \22822 , \22370 );
buf \U$16996 ( \22823 , \22371 );
buf \U$16997 ( \22824 , \22372 );
buf \U$16998 ( \22825 , \22375 );
buf \U$16999 ( \22826 , \22379 );
buf \U$17000 ( \22827 , \22382 );
buf \U$17001 ( \22828 , \22382 );
buf \U$17002 ( \22829 , \22382 );
buf \U$17003 ( \22830 , \22382 );
buf \U$17004 ( \22831 , \22382 );
buf \U$17005 ( \22832 , \22382 );
buf \U$17006 ( \22833 , \22382 );
buf \U$17007 ( \22834 , \22382 );
buf \U$17008 ( \22835 , \22382 );
buf \U$17009 ( \22836 , \22382 );
buf \U$17010 ( \22837 , \22382 );
buf \U$17011 ( \22838 , \22382 );
buf \U$17012 ( \22839 , \22382 );
buf \U$17013 ( \22840 , \22382 );
buf \U$17014 ( \22841 , \22382 );
buf \U$17015 ( \22842 , \22382 );
buf \U$17016 ( \22843 , \22382 );
buf \U$17017 ( \22844 , \22382 );
buf \U$17018 ( \22845 , \22382 );
buf \U$17019 ( \22846 , \22382 );
buf \U$17020 ( \22847 , \22382 );
buf \U$17021 ( \22848 , \22382 );
buf \U$17022 ( \22849 , \22382 );
buf \U$17023 ( \22850 , \22382 );
buf \U$17024 ( \22851 , \22382 );
buf \U$17025 ( \22852 , \22369 );
or \U$17026 ( \22853 , \22822 , \22823 , \22824 , \22825 , \22826 , \22827 , \22828 , \22829 , \22830 , \22831 , \22832 , \22833 , \22834 , \22835 , \22836 , \22837 , \22838 , \22839 , \22840 , \22841 , \22842 , \22843 , \22844 , \22845 , \22846 , \22847 , \22848 , \22849 , \22850 , \22851 , \22852 );
nand \U$17027 ( \22854 , \22821 , \22853 );
buf \U$17028 ( \22855 , \22854 );
buf \U$17029 ( \22856 , \22382 );
not \U$17030 ( \22857 , \22856 );
buf \U$17031 ( \22858 , \22379 );
buf \U$17032 ( \22859 , \22382 );
buf \U$17033 ( \22860 , \22382 );
buf \U$17034 ( \22861 , \22382 );
buf \U$17035 ( \22862 , \22382 );
buf \U$17036 ( \22863 , \22382 );
buf \U$17037 ( \22864 , \22382 );
buf \U$17038 ( \22865 , \22382 );
buf \U$17039 ( \22866 , \22382 );
buf \U$17040 ( \22867 , \22382 );
buf \U$17041 ( \22868 , \22382 );
buf \U$17042 ( \22869 , \22382 );
buf \U$17043 ( \22870 , \22382 );
buf \U$17044 ( \22871 , \22382 );
buf \U$17045 ( \22872 , \22382 );
buf \U$17046 ( \22873 , \22382 );
buf \U$17047 ( \22874 , \22382 );
buf \U$17048 ( \22875 , \22382 );
buf \U$17049 ( \22876 , \22382 );
buf \U$17050 ( \22877 , \22382 );
buf \U$17051 ( \22878 , \22382 );
buf \U$17052 ( \22879 , \22382 );
buf \U$17053 ( \22880 , \22382 );
buf \U$17054 ( \22881 , \22382 );
buf \U$17055 ( \22882 , \22382 );
buf \U$17056 ( \22883 , \22382 );
buf \U$17057 ( \22884 , \22375 );
buf \U$17058 ( \22885 , \22369 );
buf \U$17059 ( \22886 , \22370 );
buf \U$17060 ( \22887 , \22371 );
buf \U$17061 ( \22888 , \22372 );
or \U$17062 ( \22889 , \22885 , \22886 , \22887 , \22888 );
and \U$17063 ( \22890 , \22884 , \22889 );
or \U$17064 ( \22891 , \22858 , \22859 , \22860 , \22861 , \22862 , \22863 , \22864 , \22865 , \22866 , \22867 , \22868 , \22869 , \22870 , \22871 , \22872 , \22873 , \22874 , \22875 , \22876 , \22877 , \22878 , \22879 , \22880 , \22881 , \22882 , \22883 , \22890 );
and \U$17065 ( \22892 , \22857 , \22891 );
buf \U$17066 ( \22893 , \22892 );
or \U$17067 ( \22894 , \22855 , \22893 );
_DC g705f ( \22895_nG705f , \22819 , \22894 );
not \U$17068 ( \22896 , \22895_nG705f );
buf \U$17069 ( \22897 , RIb7b9608_246);
buf \U$17070 ( \22898 , \22382 );
buf \U$17071 ( \22899 , \22382 );
buf \U$17072 ( \22900 , \22382 );
buf \U$17073 ( \22901 , \22382 );
buf \U$17074 ( \22902 , \22382 );
buf \U$17075 ( \22903 , \22382 );
buf \U$17076 ( \22904 , \22382 );
buf \U$17077 ( \22905 , \22382 );
buf \U$17078 ( \22906 , \22382 );
buf \U$17079 ( \22907 , \22382 );
buf \U$17080 ( \22908 , \22382 );
buf \U$17081 ( \22909 , \22382 );
buf \U$17082 ( \22910 , \22382 );
buf \U$17083 ( \22911 , \22382 );
buf \U$17084 ( \22912 , \22382 );
buf \U$17085 ( \22913 , \22382 );
buf \U$17086 ( \22914 , \22382 );
buf \U$17087 ( \22915 , \22382 );
buf \U$17088 ( \22916 , \22382 );
buf \U$17089 ( \22917 , \22382 );
buf \U$17090 ( \22918 , \22382 );
buf \U$17091 ( \22919 , \22382 );
buf \U$17092 ( \22920 , \22382 );
buf \U$17093 ( \22921 , \22382 );
buf \U$17094 ( \22922 , \22382 );
nor \U$17095 ( \22923 , \22369 , \22370 , \22371 , \22372 , \22376 , \22379 , \22382 , \22898 , \22899 , \22900 , \22901 , \22902 , \22903 , \22904 , \22905 , \22906 , \22907 , \22908 , \22909 , \22910 , \22911 , \22912 , \22913 , \22914 , \22915 , \22916 , \22917 , \22918 , \22919 , \22920 , \22921 , \22922 );
and \U$17096 ( \22924 , \7117 , \22923 );
buf \U$17097 ( \22925 , \22382 );
buf \U$17098 ( \22926 , \22382 );
buf \U$17099 ( \22927 , \22382 );
buf \U$17100 ( \22928 , \22382 );
buf \U$17101 ( \22929 , \22382 );
buf \U$17102 ( \22930 , \22382 );
buf \U$17103 ( \22931 , \22382 );
buf \U$17104 ( \22932 , \22382 );
buf \U$17105 ( \22933 , \22382 );
buf \U$17106 ( \22934 , \22382 );
buf \U$17107 ( \22935 , \22382 );
buf \U$17108 ( \22936 , \22382 );
buf \U$17109 ( \22937 , \22382 );
buf \U$17110 ( \22938 , \22382 );
buf \U$17111 ( \22939 , \22382 );
buf \U$17112 ( \22940 , \22382 );
buf \U$17113 ( \22941 , \22382 );
buf \U$17114 ( \22942 , \22382 );
buf \U$17115 ( \22943 , \22382 );
buf \U$17116 ( \22944 , \22382 );
buf \U$17117 ( \22945 , \22382 );
buf \U$17118 ( \22946 , \22382 );
buf \U$17119 ( \22947 , \22382 );
buf \U$17120 ( \22948 , \22382 );
buf \U$17121 ( \22949 , \22382 );
nor \U$17122 ( \22950 , \22410 , \22411 , \22412 , \22413 , \22375 , \22379 , \22382 , \22925 , \22926 , \22927 , \22928 , \22929 , \22930 , \22931 , \22932 , \22933 , \22934 , \22935 , \22936 , \22937 , \22938 , \22939 , \22940 , \22941 , \22942 , \22943 , \22944 , \22945 , \22946 , \22947 , \22948 , \22949 );
and \U$17123 ( \22951 , \7119 , \22950 );
buf \U$17124 ( \22952 , \22382 );
buf \U$17125 ( \22953 , \22382 );
buf \U$17126 ( \22954 , \22382 );
buf \U$17127 ( \22955 , \22382 );
buf \U$17128 ( \22956 , \22382 );
buf \U$17129 ( \22957 , \22382 );
buf \U$17130 ( \22958 , \22382 );
buf \U$17131 ( \22959 , \22382 );
buf \U$17132 ( \22960 , \22382 );
buf \U$17133 ( \22961 , \22382 );
buf \U$17134 ( \22962 , \22382 );
buf \U$17135 ( \22963 , \22382 );
buf \U$17136 ( \22964 , \22382 );
buf \U$17137 ( \22965 , \22382 );
buf \U$17138 ( \22966 , \22382 );
buf \U$17139 ( \22967 , \22382 );
buf \U$17140 ( \22968 , \22382 );
buf \U$17141 ( \22969 , \22382 );
buf \U$17142 ( \22970 , \22382 );
buf \U$17143 ( \22971 , \22382 );
buf \U$17144 ( \22972 , \22382 );
buf \U$17145 ( \22973 , \22382 );
buf \U$17146 ( \22974 , \22382 );
buf \U$17147 ( \22975 , \22382 );
buf \U$17148 ( \22976 , \22382 );
nor \U$17149 ( \22977 , \22369 , \22411 , \22412 , \22413 , \22375 , \22379 , \22382 , \22952 , \22953 , \22954 , \22955 , \22956 , \22957 , \22958 , \22959 , \22960 , \22961 , \22962 , \22963 , \22964 , \22965 , \22966 , \22967 , \22968 , \22969 , \22970 , \22971 , \22972 , \22973 , \22974 , \22975 , \22976 );
and \U$17150 ( \22978 , \7864 , \22977 );
buf \U$17151 ( \22979 , \22382 );
buf \U$17152 ( \22980 , \22382 );
buf \U$17153 ( \22981 , \22382 );
buf \U$17154 ( \22982 , \22382 );
buf \U$17155 ( \22983 , \22382 );
buf \U$17156 ( \22984 , \22382 );
buf \U$17157 ( \22985 , \22382 );
buf \U$17158 ( \22986 , \22382 );
buf \U$17159 ( \22987 , \22382 );
buf \U$17160 ( \22988 , \22382 );
buf \U$17161 ( \22989 , \22382 );
buf \U$17162 ( \22990 , \22382 );
buf \U$17163 ( \22991 , \22382 );
buf \U$17164 ( \22992 , \22382 );
buf \U$17165 ( \22993 , \22382 );
buf \U$17166 ( \22994 , \22382 );
buf \U$17167 ( \22995 , \22382 );
buf \U$17168 ( \22996 , \22382 );
buf \U$17169 ( \22997 , \22382 );
buf \U$17170 ( \22998 , \22382 );
buf \U$17171 ( \22999 , \22382 );
buf \U$17172 ( \23000 , \22382 );
buf \U$17173 ( \23001 , \22382 );
buf \U$17174 ( \23002 , \22382 );
buf \U$17175 ( \23003 , \22382 );
nor \U$17176 ( \23004 , \22410 , \22370 , \22412 , \22413 , \22375 , \22379 , \22382 , \22979 , \22980 , \22981 , \22982 , \22983 , \22984 , \22985 , \22986 , \22987 , \22988 , \22989 , \22990 , \22991 , \22992 , \22993 , \22994 , \22995 , \22996 , \22997 , \22998 , \22999 , \23000 , \23001 , \23002 , \23003 );
and \U$17177 ( \23005 , \7892 , \23004 );
buf \U$17178 ( \23006 , \22382 );
buf \U$17179 ( \23007 , \22382 );
buf \U$17180 ( \23008 , \22382 );
buf \U$17181 ( \23009 , \22382 );
buf \U$17182 ( \23010 , \22382 );
buf \U$17183 ( \23011 , \22382 );
buf \U$17184 ( \23012 , \22382 );
buf \U$17185 ( \23013 , \22382 );
buf \U$17186 ( \23014 , \22382 );
buf \U$17187 ( \23015 , \22382 );
buf \U$17188 ( \23016 , \22382 );
buf \U$17189 ( \23017 , \22382 );
buf \U$17190 ( \23018 , \22382 );
buf \U$17191 ( \23019 , \22382 );
buf \U$17192 ( \23020 , \22382 );
buf \U$17193 ( \23021 , \22382 );
buf \U$17194 ( \23022 , \22382 );
buf \U$17195 ( \23023 , \22382 );
buf \U$17196 ( \23024 , \22382 );
buf \U$17197 ( \23025 , \22382 );
buf \U$17198 ( \23026 , \22382 );
buf \U$17199 ( \23027 , \22382 );
buf \U$17200 ( \23028 , \22382 );
buf \U$17201 ( \23029 , \22382 );
buf \U$17202 ( \23030 , \22382 );
nor \U$17203 ( \23031 , \22369 , \22370 , \22412 , \22413 , \22375 , \22379 , \22382 , \23006 , \23007 , \23008 , \23009 , \23010 , \23011 , \23012 , \23013 , \23014 , \23015 , \23016 , \23017 , \23018 , \23019 , \23020 , \23021 , \23022 , \23023 , \23024 , \23025 , \23026 , \23027 , \23028 , \23029 , \23030 );
and \U$17204 ( \23032 , \7920 , \23031 );
buf \U$17205 ( \23033 , \22382 );
buf \U$17206 ( \23034 , \22382 );
buf \U$17207 ( \23035 , \22382 );
buf \U$17208 ( \23036 , \22382 );
buf \U$17209 ( \23037 , \22382 );
buf \U$17210 ( \23038 , \22382 );
buf \U$17211 ( \23039 , \22382 );
buf \U$17212 ( \23040 , \22382 );
buf \U$17213 ( \23041 , \22382 );
buf \U$17214 ( \23042 , \22382 );
buf \U$17215 ( \23043 , \22382 );
buf \U$17216 ( \23044 , \22382 );
buf \U$17217 ( \23045 , \22382 );
buf \U$17218 ( \23046 , \22382 );
buf \U$17219 ( \23047 , \22382 );
buf \U$17220 ( \23048 , \22382 );
buf \U$17221 ( \23049 , \22382 );
buf \U$17222 ( \23050 , \22382 );
buf \U$17223 ( \23051 , \22382 );
buf \U$17224 ( \23052 , \22382 );
buf \U$17225 ( \23053 , \22382 );
buf \U$17226 ( \23054 , \22382 );
buf \U$17227 ( \23055 , \22382 );
buf \U$17228 ( \23056 , \22382 );
buf \U$17229 ( \23057 , \22382 );
nor \U$17230 ( \23058 , \22410 , \22411 , \22371 , \22413 , \22375 , \22379 , \22382 , \23033 , \23034 , \23035 , \23036 , \23037 , \23038 , \23039 , \23040 , \23041 , \23042 , \23043 , \23044 , \23045 , \23046 , \23047 , \23048 , \23049 , \23050 , \23051 , \23052 , \23053 , \23054 , \23055 , \23056 , \23057 );
and \U$17231 ( \23059 , \7948 , \23058 );
buf \U$17232 ( \23060 , \22382 );
buf \U$17233 ( \23061 , \22382 );
buf \U$17234 ( \23062 , \22382 );
buf \U$17235 ( \23063 , \22382 );
buf \U$17236 ( \23064 , \22382 );
buf \U$17237 ( \23065 , \22382 );
buf \U$17238 ( \23066 , \22382 );
buf \U$17239 ( \23067 , \22382 );
buf \U$17240 ( \23068 , \22382 );
buf \U$17241 ( \23069 , \22382 );
buf \U$17242 ( \23070 , \22382 );
buf \U$17243 ( \23071 , \22382 );
buf \U$17244 ( \23072 , \22382 );
buf \U$17245 ( \23073 , \22382 );
buf \U$17246 ( \23074 , \22382 );
buf \U$17247 ( \23075 , \22382 );
buf \U$17248 ( \23076 , \22382 );
buf \U$17249 ( \23077 , \22382 );
buf \U$17250 ( \23078 , \22382 );
buf \U$17251 ( \23079 , \22382 );
buf \U$17252 ( \23080 , \22382 );
buf \U$17253 ( \23081 , \22382 );
buf \U$17254 ( \23082 , \22382 );
buf \U$17255 ( \23083 , \22382 );
buf \U$17256 ( \23084 , \22382 );
nor \U$17257 ( \23085 , \22369 , \22411 , \22371 , \22413 , \22375 , \22379 , \22382 , \23060 , \23061 , \23062 , \23063 , \23064 , \23065 , \23066 , \23067 , \23068 , \23069 , \23070 , \23071 , \23072 , \23073 , \23074 , \23075 , \23076 , \23077 , \23078 , \23079 , \23080 , \23081 , \23082 , \23083 , \23084 );
and \U$17258 ( \23086 , \7976 , \23085 );
buf \U$17259 ( \23087 , \22382 );
buf \U$17260 ( \23088 , \22382 );
buf \U$17261 ( \23089 , \22382 );
buf \U$17262 ( \23090 , \22382 );
buf \U$17263 ( \23091 , \22382 );
buf \U$17264 ( \23092 , \22382 );
buf \U$17265 ( \23093 , \22382 );
buf \U$17266 ( \23094 , \22382 );
buf \U$17267 ( \23095 , \22382 );
buf \U$17268 ( \23096 , \22382 );
buf \U$17269 ( \23097 , \22382 );
buf \U$17270 ( \23098 , \22382 );
buf \U$17271 ( \23099 , \22382 );
buf \U$17272 ( \23100 , \22382 );
buf \U$17273 ( \23101 , \22382 );
buf \U$17274 ( \23102 , \22382 );
buf \U$17275 ( \23103 , \22382 );
buf \U$17276 ( \23104 , \22382 );
buf \U$17277 ( \23105 , \22382 );
buf \U$17278 ( \23106 , \22382 );
buf \U$17279 ( \23107 , \22382 );
buf \U$17280 ( \23108 , \22382 );
buf \U$17281 ( \23109 , \22382 );
buf \U$17282 ( \23110 , \22382 );
buf \U$17283 ( \23111 , \22382 );
nor \U$17284 ( \23112 , \22410 , \22370 , \22371 , \22413 , \22375 , \22379 , \22382 , \23087 , \23088 , \23089 , \23090 , \23091 , \23092 , \23093 , \23094 , \23095 , \23096 , \23097 , \23098 , \23099 , \23100 , \23101 , \23102 , \23103 , \23104 , \23105 , \23106 , \23107 , \23108 , \23109 , \23110 , \23111 );
and \U$17285 ( \23113 , \8004 , \23112 );
buf \U$17286 ( \23114 , \22382 );
buf \U$17287 ( \23115 , \22382 );
buf \U$17288 ( \23116 , \22382 );
buf \U$17289 ( \23117 , \22382 );
buf \U$17290 ( \23118 , \22382 );
buf \U$17291 ( \23119 , \22382 );
buf \U$17292 ( \23120 , \22382 );
buf \U$17293 ( \23121 , \22382 );
buf \U$17294 ( \23122 , \22382 );
buf \U$17295 ( \23123 , \22382 );
buf \U$17296 ( \23124 , \22382 );
buf \U$17297 ( \23125 , \22382 );
buf \U$17298 ( \23126 , \22382 );
buf \U$17299 ( \23127 , \22382 );
buf \U$17300 ( \23128 , \22382 );
buf \U$17301 ( \23129 , \22382 );
buf \U$17302 ( \23130 , \22382 );
buf \U$17303 ( \23131 , \22382 );
buf \U$17304 ( \23132 , \22382 );
buf \U$17305 ( \23133 , \22382 );
buf \U$17306 ( \23134 , \22382 );
buf \U$17307 ( \23135 , \22382 );
buf \U$17308 ( \23136 , \22382 );
buf \U$17309 ( \23137 , \22382 );
buf \U$17310 ( \23138 , \22382 );
nor \U$17311 ( \23139 , \22369 , \22370 , \22371 , \22413 , \22375 , \22379 , \22382 , \23114 , \23115 , \23116 , \23117 , \23118 , \23119 , \23120 , \23121 , \23122 , \23123 , \23124 , \23125 , \23126 , \23127 , \23128 , \23129 , \23130 , \23131 , \23132 , \23133 , \23134 , \23135 , \23136 , \23137 , \23138 );
and \U$17312 ( \23140 , \8032 , \23139 );
buf \U$17313 ( \23141 , \22382 );
buf \U$17314 ( \23142 , \22382 );
buf \U$17315 ( \23143 , \22382 );
buf \U$17316 ( \23144 , \22382 );
buf \U$17317 ( \23145 , \22382 );
buf \U$17318 ( \23146 , \22382 );
buf \U$17319 ( \23147 , \22382 );
buf \U$17320 ( \23148 , \22382 );
buf \U$17321 ( \23149 , \22382 );
buf \U$17322 ( \23150 , \22382 );
buf \U$17323 ( \23151 , \22382 );
buf \U$17324 ( \23152 , \22382 );
buf \U$17325 ( \23153 , \22382 );
buf \U$17326 ( \23154 , \22382 );
buf \U$17327 ( \23155 , \22382 );
buf \U$17328 ( \23156 , \22382 );
buf \U$17329 ( \23157 , \22382 );
buf \U$17330 ( \23158 , \22382 );
buf \U$17331 ( \23159 , \22382 );
buf \U$17332 ( \23160 , \22382 );
buf \U$17333 ( \23161 , \22382 );
buf \U$17334 ( \23162 , \22382 );
buf \U$17335 ( \23163 , \22382 );
buf \U$17336 ( \23164 , \22382 );
buf \U$17337 ( \23165 , \22382 );
nor \U$17338 ( \23166 , \22410 , \22411 , \22412 , \22372 , \22375 , \22379 , \22382 , \23141 , \23142 , \23143 , \23144 , \23145 , \23146 , \23147 , \23148 , \23149 , \23150 , \23151 , \23152 , \23153 , \23154 , \23155 , \23156 , \23157 , \23158 , \23159 , \23160 , \23161 , \23162 , \23163 , \23164 , \23165 );
and \U$17339 ( \23167 , \8060 , \23166 );
buf \U$17340 ( \23168 , \22382 );
buf \U$17341 ( \23169 , \22382 );
buf \U$17342 ( \23170 , \22382 );
buf \U$17343 ( \23171 , \22382 );
buf \U$17344 ( \23172 , \22382 );
buf \U$17345 ( \23173 , \22382 );
buf \U$17346 ( \23174 , \22382 );
buf \U$17347 ( \23175 , \22382 );
buf \U$17348 ( \23176 , \22382 );
buf \U$17349 ( \23177 , \22382 );
buf \U$17350 ( \23178 , \22382 );
buf \U$17351 ( \23179 , \22382 );
buf \U$17352 ( \23180 , \22382 );
buf \U$17353 ( \23181 , \22382 );
buf \U$17354 ( \23182 , \22382 );
buf \U$17355 ( \23183 , \22382 );
buf \U$17356 ( \23184 , \22382 );
buf \U$17357 ( \23185 , \22382 );
buf \U$17358 ( \23186 , \22382 );
buf \U$17359 ( \23187 , \22382 );
buf \U$17360 ( \23188 , \22382 );
buf \U$17361 ( \23189 , \22382 );
buf \U$17362 ( \23190 , \22382 );
buf \U$17363 ( \23191 , \22382 );
buf \U$17364 ( \23192 , \22382 );
nor \U$17365 ( \23193 , \22369 , \22411 , \22412 , \22372 , \22375 , \22379 , \22382 , \23168 , \23169 , \23170 , \23171 , \23172 , \23173 , \23174 , \23175 , \23176 , \23177 , \23178 , \23179 , \23180 , \23181 , \23182 , \23183 , \23184 , \23185 , \23186 , \23187 , \23188 , \23189 , \23190 , \23191 , \23192 );
and \U$17366 ( \23194 , \8088 , \23193 );
buf \U$17367 ( \23195 , \22382 );
buf \U$17368 ( \23196 , \22382 );
buf \U$17369 ( \23197 , \22382 );
buf \U$17370 ( \23198 , \22382 );
buf \U$17371 ( \23199 , \22382 );
buf \U$17372 ( \23200 , \22382 );
buf \U$17373 ( \23201 , \22382 );
buf \U$17374 ( \23202 , \22382 );
buf \U$17375 ( \23203 , \22382 );
buf \U$17376 ( \23204 , \22382 );
buf \U$17377 ( \23205 , \22382 );
buf \U$17378 ( \23206 , \22382 );
buf \U$17379 ( \23207 , \22382 );
buf \U$17380 ( \23208 , \22382 );
buf \U$17381 ( \23209 , \22382 );
buf \U$17382 ( \23210 , \22382 );
buf \U$17383 ( \23211 , \22382 );
buf \U$17384 ( \23212 , \22382 );
buf \U$17385 ( \23213 , \22382 );
buf \U$17386 ( \23214 , \22382 );
buf \U$17387 ( \23215 , \22382 );
buf \U$17388 ( \23216 , \22382 );
buf \U$17389 ( \23217 , \22382 );
buf \U$17390 ( \23218 , \22382 );
buf \U$17391 ( \23219 , \22382 );
nor \U$17392 ( \23220 , \22410 , \22370 , \22412 , \22372 , \22375 , \22379 , \22382 , \23195 , \23196 , \23197 , \23198 , \23199 , \23200 , \23201 , \23202 , \23203 , \23204 , \23205 , \23206 , \23207 , \23208 , \23209 , \23210 , \23211 , \23212 , \23213 , \23214 , \23215 , \23216 , \23217 , \23218 , \23219 );
and \U$17393 ( \23221 , \8116 , \23220 );
buf \U$17394 ( \23222 , \22382 );
buf \U$17395 ( \23223 , \22382 );
buf \U$17396 ( \23224 , \22382 );
buf \U$17397 ( \23225 , \22382 );
buf \U$17398 ( \23226 , \22382 );
buf \U$17399 ( \23227 , \22382 );
buf \U$17400 ( \23228 , \22382 );
buf \U$17401 ( \23229 , \22382 );
buf \U$17402 ( \23230 , \22382 );
buf \U$17403 ( \23231 , \22382 );
buf \U$17404 ( \23232 , \22382 );
buf \U$17405 ( \23233 , \22382 );
buf \U$17406 ( \23234 , \22382 );
buf \U$17407 ( \23235 , \22382 );
buf \U$17408 ( \23236 , \22382 );
buf \U$17409 ( \23237 , \22382 );
buf \U$17410 ( \23238 , \22382 );
buf \U$17411 ( \23239 , \22382 );
buf \U$17412 ( \23240 , \22382 );
buf \U$17413 ( \23241 , \22382 );
buf \U$17414 ( \23242 , \22382 );
buf \U$17415 ( \23243 , \22382 );
buf \U$17416 ( \23244 , \22382 );
buf \U$17417 ( \23245 , \22382 );
buf \U$17418 ( \23246 , \22382 );
nor \U$17419 ( \23247 , \22369 , \22370 , \22412 , \22372 , \22375 , \22379 , \22382 , \23222 , \23223 , \23224 , \23225 , \23226 , \23227 , \23228 , \23229 , \23230 , \23231 , \23232 , \23233 , \23234 , \23235 , \23236 , \23237 , \23238 , \23239 , \23240 , \23241 , \23242 , \23243 , \23244 , \23245 , \23246 );
and \U$17420 ( \23248 , \8144 , \23247 );
buf \U$17421 ( \23249 , \22382 );
buf \U$17422 ( \23250 , \22382 );
buf \U$17423 ( \23251 , \22382 );
buf \U$17424 ( \23252 , \22382 );
buf \U$17425 ( \23253 , \22382 );
buf \U$17426 ( \23254 , \22382 );
buf \U$17427 ( \23255 , \22382 );
buf \U$17428 ( \23256 , \22382 );
buf \U$17429 ( \23257 , \22382 );
buf \U$17430 ( \23258 , \22382 );
buf \U$17431 ( \23259 , \22382 );
buf \U$17432 ( \23260 , \22382 );
buf \U$17433 ( \23261 , \22382 );
buf \U$17434 ( \23262 , \22382 );
buf \U$17435 ( \23263 , \22382 );
buf \U$17436 ( \23264 , \22382 );
buf \U$17437 ( \23265 , \22382 );
buf \U$17438 ( \23266 , \22382 );
buf \U$17439 ( \23267 , \22382 );
buf \U$17440 ( \23268 , \22382 );
buf \U$17441 ( \23269 , \22382 );
buf \U$17442 ( \23270 , \22382 );
buf \U$17443 ( \23271 , \22382 );
buf \U$17444 ( \23272 , \22382 );
buf \U$17445 ( \23273 , \22382 );
nor \U$17446 ( \23274 , \22410 , \22411 , \22371 , \22372 , \22375 , \22379 , \22382 , \23249 , \23250 , \23251 , \23252 , \23253 , \23254 , \23255 , \23256 , \23257 , \23258 , \23259 , \23260 , \23261 , \23262 , \23263 , \23264 , \23265 , \23266 , \23267 , \23268 , \23269 , \23270 , \23271 , \23272 , \23273 );
and \U$17447 ( \23275 , \8172 , \23274 );
buf \U$17448 ( \23276 , \22382 );
buf \U$17449 ( \23277 , \22382 );
buf \U$17450 ( \23278 , \22382 );
buf \U$17451 ( \23279 , \22382 );
buf \U$17452 ( \23280 , \22382 );
buf \U$17453 ( \23281 , \22382 );
buf \U$17454 ( \23282 , \22382 );
buf \U$17455 ( \23283 , \22382 );
buf \U$17456 ( \23284 , \22382 );
buf \U$17457 ( \23285 , \22382 );
buf \U$17458 ( \23286 , \22382 );
buf \U$17459 ( \23287 , \22382 );
buf \U$17460 ( \23288 , \22382 );
buf \U$17461 ( \23289 , \22382 );
buf \U$17462 ( \23290 , \22382 );
buf \U$17463 ( \23291 , \22382 );
buf \U$17464 ( \23292 , \22382 );
buf \U$17465 ( \23293 , \22382 );
buf \U$17466 ( \23294 , \22382 );
buf \U$17467 ( \23295 , \22382 );
buf \U$17468 ( \23296 , \22382 );
buf \U$17469 ( \23297 , \22382 );
buf \U$17470 ( \23298 , \22382 );
buf \U$17471 ( \23299 , \22382 );
buf \U$17472 ( \23300 , \22382 );
nor \U$17473 ( \23301 , \22369 , \22411 , \22371 , \22372 , \22375 , \22379 , \22382 , \23276 , \23277 , \23278 , \23279 , \23280 , \23281 , \23282 , \23283 , \23284 , \23285 , \23286 , \23287 , \23288 , \23289 , \23290 , \23291 , \23292 , \23293 , \23294 , \23295 , \23296 , \23297 , \23298 , \23299 , \23300 );
and \U$17474 ( \23302 , \8200 , \23301 );
buf \U$17475 ( \23303 , \22382 );
buf \U$17476 ( \23304 , \22382 );
buf \U$17477 ( \23305 , \22382 );
buf \U$17478 ( \23306 , \22382 );
buf \U$17479 ( \23307 , \22382 );
buf \U$17480 ( \23308 , \22382 );
buf \U$17481 ( \23309 , \22382 );
buf \U$17482 ( \23310 , \22382 );
buf \U$17483 ( \23311 , \22382 );
buf \U$17484 ( \23312 , \22382 );
buf \U$17485 ( \23313 , \22382 );
buf \U$17486 ( \23314 , \22382 );
buf \U$17487 ( \23315 , \22382 );
buf \U$17488 ( \23316 , \22382 );
buf \U$17489 ( \23317 , \22382 );
buf \U$17490 ( \23318 , \22382 );
buf \U$17491 ( \23319 , \22382 );
buf \U$17492 ( \23320 , \22382 );
buf \U$17493 ( \23321 , \22382 );
buf \U$17494 ( \23322 , \22382 );
buf \U$17495 ( \23323 , \22382 );
buf \U$17496 ( \23324 , \22382 );
buf \U$17497 ( \23325 , \22382 );
buf \U$17498 ( \23326 , \22382 );
buf \U$17499 ( \23327 , \22382 );
nor \U$17500 ( \23328 , \22410 , \22370 , \22371 , \22372 , \22375 , \22379 , \22382 , \23303 , \23304 , \23305 , \23306 , \23307 , \23308 , \23309 , \23310 , \23311 , \23312 , \23313 , \23314 , \23315 , \23316 , \23317 , \23318 , \23319 , \23320 , \23321 , \23322 , \23323 , \23324 , \23325 , \23326 , \23327 );
and \U$17501 ( \23329 , \8228 , \23328 );
or \U$17502 ( \23330 , \22924 , \22951 , \22978 , \23005 , \23032 , \23059 , \23086 , \23113 , \23140 , \23167 , \23194 , \23221 , \23248 , \23275 , \23302 , \23329 );
buf \U$17503 ( \23331 , \22382 );
not \U$17504 ( \23332 , \23331 );
buf \U$17505 ( \23333 , \22370 );
buf \U$17506 ( \23334 , \22371 );
buf \U$17507 ( \23335 , \22372 );
buf \U$17508 ( \23336 , \22375 );
buf \U$17509 ( \23337 , \22379 );
buf \U$17510 ( \23338 , \22382 );
buf \U$17511 ( \23339 , \22382 );
buf \U$17512 ( \23340 , \22382 );
buf \U$17513 ( \23341 , \22382 );
buf \U$17514 ( \23342 , \22382 );
buf \U$17515 ( \23343 , \22382 );
buf \U$17516 ( \23344 , \22382 );
buf \U$17517 ( \23345 , \22382 );
buf \U$17518 ( \23346 , \22382 );
buf \U$17519 ( \23347 , \22382 );
buf \U$17520 ( \23348 , \22382 );
buf \U$17521 ( \23349 , \22382 );
buf \U$17522 ( \23350 , \22382 );
buf \U$17523 ( \23351 , \22382 );
buf \U$17524 ( \23352 , \22382 );
buf \U$17525 ( \23353 , \22382 );
buf \U$17526 ( \23354 , \22382 );
buf \U$17527 ( \23355 , \22382 );
buf \U$17528 ( \23356 , \22382 );
buf \U$17529 ( \23357 , \22382 );
buf \U$17530 ( \23358 , \22382 );
buf \U$17531 ( \23359 , \22382 );
buf \U$17532 ( \23360 , \22382 );
buf \U$17533 ( \23361 , \22382 );
buf \U$17534 ( \23362 , \22382 );
buf \U$17535 ( \23363 , \22369 );
or \U$17536 ( \23364 , \23333 , \23334 , \23335 , \23336 , \23337 , \23338 , \23339 , \23340 , \23341 , \23342 , \23343 , \23344 , \23345 , \23346 , \23347 , \23348 , \23349 , \23350 , \23351 , \23352 , \23353 , \23354 , \23355 , \23356 , \23357 , \23358 , \23359 , \23360 , \23361 , \23362 , \23363 );
nand \U$17537 ( \23365 , \23332 , \23364 );
buf \U$17538 ( \23366 , \23365 );
buf \U$17539 ( \23367 , \22382 );
not \U$17540 ( \23368 , \23367 );
buf \U$17541 ( \23369 , \22379 );
buf \U$17542 ( \23370 , \22382 );
buf \U$17543 ( \23371 , \22382 );
buf \U$17544 ( \23372 , \22382 );
buf \U$17545 ( \23373 , \22382 );
buf \U$17546 ( \23374 , \22382 );
buf \U$17547 ( \23375 , \22382 );
buf \U$17548 ( \23376 , \22382 );
buf \U$17549 ( \23377 , \22382 );
buf \U$17550 ( \23378 , \22382 );
buf \U$17551 ( \23379 , \22382 );
buf \U$17552 ( \23380 , \22382 );
buf \U$17553 ( \23381 , \22382 );
buf \U$17554 ( \23382 , \22382 );
buf \U$17555 ( \23383 , \22382 );
buf \U$17556 ( \23384 , \22382 );
buf \U$17557 ( \23385 , \22382 );
buf \U$17558 ( \23386 , \22382 );
buf \U$17559 ( \23387 , \22382 );
buf \U$17560 ( \23388 , \22382 );
buf \U$17561 ( \23389 , \22382 );
buf \U$17562 ( \23390 , \22382 );
buf \U$17563 ( \23391 , \22382 );
buf \U$17564 ( \23392 , \22382 );
buf \U$17565 ( \23393 , \22382 );
buf \U$17566 ( \23394 , \22382 );
buf \U$17567 ( \23395 , \22375 );
buf \U$17568 ( \23396 , \22369 );
buf \U$17569 ( \23397 , \22370 );
buf \U$17570 ( \23398 , \22371 );
buf \U$17571 ( \23399 , \22372 );
or \U$17572 ( \23400 , \23396 , \23397 , \23398 , \23399 );
and \U$17573 ( \23401 , \23395 , \23400 );
or \U$17574 ( \23402 , \23369 , \23370 , \23371 , \23372 , \23373 , \23374 , \23375 , \23376 , \23377 , \23378 , \23379 , \23380 , \23381 , \23382 , \23383 , \23384 , \23385 , \23386 , \23387 , \23388 , \23389 , \23390 , \23391 , \23392 , \23393 , \23394 , \23401 );
and \U$17575 ( \23403 , \23368 , \23402 );
buf \U$17576 ( \23404 , \23403 );
or \U$17577 ( \23405 , \23366 , \23404 );
_DC g725e ( \23406_nG725e , \23330 , \23405 );
buf \U$17578 ( \23407 , \23406_nG725e );
xor \U$17579 ( \23408 , \22897 , \23407 );
buf \U$17580 ( \23409 , RIb7b9590_247);
and \U$17581 ( \23410 , \7126 , \22923 );
and \U$17582 ( \23411 , \7128 , \22950 );
and \U$17583 ( \23412 , \8338 , \22977 );
and \U$17584 ( \23413 , \8340 , \23004 );
and \U$17585 ( \23414 , \8342 , \23031 );
and \U$17586 ( \23415 , \8344 , \23058 );
and \U$17587 ( \23416 , \8346 , \23085 );
and \U$17588 ( \23417 , \8348 , \23112 );
and \U$17589 ( \23418 , \8350 , \23139 );
and \U$17590 ( \23419 , \8352 , \23166 );
and \U$17591 ( \23420 , \8354 , \23193 );
and \U$17592 ( \23421 , \8356 , \23220 );
and \U$17593 ( \23422 , \8358 , \23247 );
and \U$17594 ( \23423 , \8360 , \23274 );
and \U$17595 ( \23424 , \8362 , \23301 );
and \U$17596 ( \23425 , \8364 , \23328 );
or \U$17597 ( \23426 , \23410 , \23411 , \23412 , \23413 , \23414 , \23415 , \23416 , \23417 , \23418 , \23419 , \23420 , \23421 , \23422 , \23423 , \23424 , \23425 );
_DC g7273 ( \23427_nG7273 , \23426 , \23405 );
buf \U$17598 ( \23428 , \23427_nG7273 );
xor \U$17599 ( \23429 , \23409 , \23428 );
or \U$17600 ( \23430 , \23408 , \23429 );
buf \U$17601 ( \23431 , RIb7b9518_248);
and \U$17602 ( \23432 , \7136 , \22923 );
and \U$17603 ( \23433 , \7138 , \22950 );
and \U$17604 ( \23434 , \8374 , \22977 );
and \U$17605 ( \23435 , \8376 , \23004 );
and \U$17606 ( \23436 , \8378 , \23031 );
and \U$17607 ( \23437 , \8380 , \23058 );
and \U$17608 ( \23438 , \8382 , \23085 );
and \U$17609 ( \23439 , \8384 , \23112 );
and \U$17610 ( \23440 , \8386 , \23139 );
and \U$17611 ( \23441 , \8388 , \23166 );
and \U$17612 ( \23442 , \8390 , \23193 );
and \U$17613 ( \23443 , \8392 , \23220 );
and \U$17614 ( \23444 , \8394 , \23247 );
and \U$17615 ( \23445 , \8396 , \23274 );
and \U$17616 ( \23446 , \8398 , \23301 );
and \U$17617 ( \23447 , \8400 , \23328 );
or \U$17618 ( \23448 , \23432 , \23433 , \23434 , \23435 , \23436 , \23437 , \23438 , \23439 , \23440 , \23441 , \23442 , \23443 , \23444 , \23445 , \23446 , \23447 );
_DC g7289 ( \23449_nG7289 , \23448 , \23405 );
buf \U$17619 ( \23450 , \23449_nG7289 );
xor \U$17620 ( \23451 , \23431 , \23450 );
or \U$17621 ( \23452 , \23430 , \23451 );
buf \U$17622 ( \23453 , RIb7b94a0_249);
and \U$17623 ( \23454 , \7146 , \22923 );
and \U$17624 ( \23455 , \7148 , \22950 );
and \U$17625 ( \23456 , \8410 , \22977 );
and \U$17626 ( \23457 , \8412 , \23004 );
and \U$17627 ( \23458 , \8414 , \23031 );
and \U$17628 ( \23459 , \8416 , \23058 );
and \U$17629 ( \23460 , \8418 , \23085 );
and \U$17630 ( \23461 , \8420 , \23112 );
and \U$17631 ( \23462 , \8422 , \23139 );
and \U$17632 ( \23463 , \8424 , \23166 );
and \U$17633 ( \23464 , \8426 , \23193 );
and \U$17634 ( \23465 , \8428 , \23220 );
and \U$17635 ( \23466 , \8430 , \23247 );
and \U$17636 ( \23467 , \8432 , \23274 );
and \U$17637 ( \23468 , \8434 , \23301 );
and \U$17638 ( \23469 , \8436 , \23328 );
or \U$17639 ( \23470 , \23454 , \23455 , \23456 , \23457 , \23458 , \23459 , \23460 , \23461 , \23462 , \23463 , \23464 , \23465 , \23466 , \23467 , \23468 , \23469 );
_DC g729f ( \23471_nG729f , \23470 , \23405 );
buf \U$17640 ( \23472 , \23471_nG729f );
xor \U$17641 ( \23473 , \23453 , \23472 );
or \U$17642 ( \23474 , \23452 , \23473 );
buf \U$17643 ( \23475 , RIb7b9428_250);
and \U$17644 ( \23476 , \7156 , \22923 );
and \U$17645 ( \23477 , \7158 , \22950 );
and \U$17646 ( \23478 , \8446 , \22977 );
and \U$17647 ( \23479 , \8448 , \23004 );
and \U$17648 ( \23480 , \8450 , \23031 );
and \U$17649 ( \23481 , \8452 , \23058 );
and \U$17650 ( \23482 , \8454 , \23085 );
and \U$17651 ( \23483 , \8456 , \23112 );
and \U$17652 ( \23484 , \8458 , \23139 );
and \U$17653 ( \23485 , \8460 , \23166 );
and \U$17654 ( \23486 , \8462 , \23193 );
and \U$17655 ( \23487 , \8464 , \23220 );
and \U$17656 ( \23488 , \8466 , \23247 );
and \U$17657 ( \23489 , \8468 , \23274 );
and \U$17658 ( \23490 , \8470 , \23301 );
and \U$17659 ( \23491 , \8472 , \23328 );
or \U$17660 ( \23492 , \23476 , \23477 , \23478 , \23479 , \23480 , \23481 , \23482 , \23483 , \23484 , \23485 , \23486 , \23487 , \23488 , \23489 , \23490 , \23491 );
_DC g72b5 ( \23493_nG72b5 , \23492 , \23405 );
buf \U$17661 ( \23494 , \23493_nG72b5 );
xor \U$17662 ( \23495 , \23475 , \23494 );
or \U$17663 ( \23496 , \23474 , \23495 );
buf \U$17664 ( \23497 , RIb7b93b0_251);
and \U$17665 ( \23498 , \7166 , \22923 );
and \U$17666 ( \23499 , \7168 , \22950 );
and \U$17667 ( \23500 , \8482 , \22977 );
and \U$17668 ( \23501 , \8484 , \23004 );
and \U$17669 ( \23502 , \8486 , \23031 );
and \U$17670 ( \23503 , \8488 , \23058 );
and \U$17671 ( \23504 , \8490 , \23085 );
and \U$17672 ( \23505 , \8492 , \23112 );
and \U$17673 ( \23506 , \8494 , \23139 );
and \U$17674 ( \23507 , \8496 , \23166 );
and \U$17675 ( \23508 , \8498 , \23193 );
and \U$17676 ( \23509 , \8500 , \23220 );
and \U$17677 ( \23510 , \8502 , \23247 );
and \U$17678 ( \23511 , \8504 , \23274 );
and \U$17679 ( \23512 , \8506 , \23301 );
and \U$17680 ( \23513 , \8508 , \23328 );
or \U$17681 ( \23514 , \23498 , \23499 , \23500 , \23501 , \23502 , \23503 , \23504 , \23505 , \23506 , \23507 , \23508 , \23509 , \23510 , \23511 , \23512 , \23513 );
_DC g72cb ( \23515_nG72cb , \23514 , \23405 );
buf \U$17682 ( \23516 , \23515_nG72cb );
xor \U$17683 ( \23517 , \23497 , \23516 );
or \U$17684 ( \23518 , \23496 , \23517 );
buf \U$17685 ( \23519 , RIb7af720_252);
and \U$17686 ( \23520 , \7176 , \22923 );
and \U$17687 ( \23521 , \7178 , \22950 );
and \U$17688 ( \23522 , \8518 , \22977 );
and \U$17689 ( \23523 , \8520 , \23004 );
and \U$17690 ( \23524 , \8522 , \23031 );
and \U$17691 ( \23525 , \8524 , \23058 );
and \U$17692 ( \23526 , \8526 , \23085 );
and \U$17693 ( \23527 , \8528 , \23112 );
and \U$17694 ( \23528 , \8530 , \23139 );
and \U$17695 ( \23529 , \8532 , \23166 );
and \U$17696 ( \23530 , \8534 , \23193 );
and \U$17697 ( \23531 , \8536 , \23220 );
and \U$17698 ( \23532 , \8538 , \23247 );
and \U$17699 ( \23533 , \8540 , \23274 );
and \U$17700 ( \23534 , \8542 , \23301 );
and \U$17701 ( \23535 , \8544 , \23328 );
or \U$17702 ( \23536 , \23520 , \23521 , \23522 , \23523 , \23524 , \23525 , \23526 , \23527 , \23528 , \23529 , \23530 , \23531 , \23532 , \23533 , \23534 , \23535 );
_DC g72e1 ( \23537_nG72e1 , \23536 , \23405 );
buf \U$17703 ( \23538 , \23537_nG72e1 );
xor \U$17704 ( \23539 , \23519 , \23538 );
or \U$17705 ( \23540 , \23518 , \23539 );
buf \U$17706 ( \23541 , RIb7af6a8_253);
and \U$17707 ( \23542 , \7186 , \22923 );
and \U$17708 ( \23543 , \7188 , \22950 );
and \U$17709 ( \23544 , \8554 , \22977 );
and \U$17710 ( \23545 , \8556 , \23004 );
and \U$17711 ( \23546 , \8558 , \23031 );
and \U$17712 ( \23547 , \8560 , \23058 );
and \U$17713 ( \23548 , \8562 , \23085 );
and \U$17714 ( \23549 , \8564 , \23112 );
and \U$17715 ( \23550 , \8566 , \23139 );
and \U$17716 ( \23551 , \8568 , \23166 );
and \U$17717 ( \23552 , \8570 , \23193 );
and \U$17718 ( \23553 , \8572 , \23220 );
and \U$17719 ( \23554 , \8574 , \23247 );
and \U$17720 ( \23555 , \8576 , \23274 );
and \U$17721 ( \23556 , \8578 , \23301 );
and \U$17722 ( \23557 , \8580 , \23328 );
or \U$17723 ( \23558 , \23542 , \23543 , \23544 , \23545 , \23546 , \23547 , \23548 , \23549 , \23550 , \23551 , \23552 , \23553 , \23554 , \23555 , \23556 , \23557 );
_DC g72f7 ( \23559_nG72f7 , \23558 , \23405 );
buf \U$17724 ( \23560 , \23559_nG72f7 );
xor \U$17725 ( \23561 , \23541 , \23560 );
or \U$17726 ( \23562 , \23540 , \23561 );
not \U$17727 ( \23563 , \23562 );
buf \U$17728 ( \23564 , \23563 );
and \U$17729 ( \23565 , \22896 , \23564 );
buf \U$17730 ( \23566 , RIb7af630_254);
buf \U$17731 ( \23567 , \22382 );
buf \U$17732 ( \23568 , \22382 );
buf \U$17733 ( \23569 , \22382 );
buf \U$17734 ( \23570 , \22382 );
buf \U$17735 ( \23571 , \22382 );
buf \U$17736 ( \23572 , \22382 );
buf \U$17737 ( \23573 , \22382 );
buf \U$17738 ( \23574 , \22382 );
buf \U$17739 ( \23575 , \22382 );
buf \U$17740 ( \23576 , \22382 );
buf \U$17741 ( \23577 , \22382 );
buf \U$17742 ( \23578 , \22382 );
buf \U$17743 ( \23579 , \22382 );
buf \U$17744 ( \23580 , \22382 );
buf \U$17745 ( \23581 , \22382 );
buf \U$17746 ( \23582 , \22382 );
buf \U$17747 ( \23583 , \22382 );
buf \U$17748 ( \23584 , \22382 );
buf \U$17749 ( \23585 , \22382 );
buf \U$17750 ( \23586 , \22382 );
buf \U$17751 ( \23587 , \22382 );
buf \U$17752 ( \23588 , \22382 );
buf \U$17753 ( \23589 , \22382 );
buf \U$17754 ( \23590 , \22382 );
buf \U$17755 ( \23591 , \22382 );
nor \U$17756 ( \23592 , \22369 , \22370 , \22371 , \22372 , \22376 , \22379 , \22382 , \23567 , \23568 , \23569 , \23570 , \23571 , \23572 , \23573 , \23574 , \23575 , \23576 , \23577 , \23578 , \23579 , \23580 , \23581 , \23582 , \23583 , \23584 , \23585 , \23586 , \23587 , \23588 , \23589 , \23590 , \23591 );
and \U$17757 ( \23593 , \7198 , \23592 );
buf \U$17758 ( \23594 , \22382 );
buf \U$17759 ( \23595 , \22382 );
buf \U$17760 ( \23596 , \22382 );
buf \U$17761 ( \23597 , \22382 );
buf \U$17762 ( \23598 , \22382 );
buf \U$17763 ( \23599 , \22382 );
buf \U$17764 ( \23600 , \22382 );
buf \U$17765 ( \23601 , \22382 );
buf \U$17766 ( \23602 , \22382 );
buf \U$17767 ( \23603 , \22382 );
buf \U$17768 ( \23604 , \22382 );
buf \U$17769 ( \23605 , \22382 );
buf \U$17770 ( \23606 , \22382 );
buf \U$17771 ( \23607 , \22382 );
buf \U$17772 ( \23608 , \22382 );
buf \U$17773 ( \23609 , \22382 );
buf \U$17774 ( \23610 , \22382 );
buf \U$17775 ( \23611 , \22382 );
buf \U$17776 ( \23612 , \22382 );
buf \U$17777 ( \23613 , \22382 );
buf \U$17778 ( \23614 , \22382 );
buf \U$17779 ( \23615 , \22382 );
buf \U$17780 ( \23616 , \22382 );
buf \U$17781 ( \23617 , \22382 );
buf \U$17782 ( \23618 , \22382 );
nor \U$17783 ( \23619 , \22410 , \22411 , \22412 , \22413 , \22375 , \22379 , \22382 , \23594 , \23595 , \23596 , \23597 , \23598 , \23599 , \23600 , \23601 , \23602 , \23603 , \23604 , \23605 , \23606 , \23607 , \23608 , \23609 , \23610 , \23611 , \23612 , \23613 , \23614 , \23615 , \23616 , \23617 , \23618 );
and \U$17784 ( \23620 , \7200 , \23619 );
buf \U$17785 ( \23621 , \22382 );
buf \U$17786 ( \23622 , \22382 );
buf \U$17787 ( \23623 , \22382 );
buf \U$17788 ( \23624 , \22382 );
buf \U$17789 ( \23625 , \22382 );
buf \U$17790 ( \23626 , \22382 );
buf \U$17791 ( \23627 , \22382 );
buf \U$17792 ( \23628 , \22382 );
buf \U$17793 ( \23629 , \22382 );
buf \U$17794 ( \23630 , \22382 );
buf \U$17795 ( \23631 , \22382 );
buf \U$17796 ( \23632 , \22382 );
buf \U$17797 ( \23633 , \22382 );
buf \U$17798 ( \23634 , \22382 );
buf \U$17799 ( \23635 , \22382 );
buf \U$17800 ( \23636 , \22382 );
buf \U$17801 ( \23637 , \22382 );
buf \U$17802 ( \23638 , \22382 );
buf \U$17803 ( \23639 , \22382 );
buf \U$17804 ( \23640 , \22382 );
buf \U$17805 ( \23641 , \22382 );
buf \U$17806 ( \23642 , \22382 );
buf \U$17807 ( \23643 , \22382 );
buf \U$17808 ( \23644 , \22382 );
buf \U$17809 ( \23645 , \22382 );
nor \U$17810 ( \23646 , \22369 , \22411 , \22412 , \22413 , \22375 , \22379 , \22382 , \23621 , \23622 , \23623 , \23624 , \23625 , \23626 , \23627 , \23628 , \23629 , \23630 , \23631 , \23632 , \23633 , \23634 , \23635 , \23636 , \23637 , \23638 , \23639 , \23640 , \23641 , \23642 , \23643 , \23644 , \23645 );
and \U$17811 ( \23647 , \8645 , \23646 );
buf \U$17812 ( \23648 , \22382 );
buf \U$17813 ( \23649 , \22382 );
buf \U$17814 ( \23650 , \22382 );
buf \U$17815 ( \23651 , \22382 );
buf \U$17816 ( \23652 , \22382 );
buf \U$17817 ( \23653 , \22382 );
buf \U$17818 ( \23654 , \22382 );
buf \U$17819 ( \23655 , \22382 );
buf \U$17820 ( \23656 , \22382 );
buf \U$17821 ( \23657 , \22382 );
buf \U$17822 ( \23658 , \22382 );
buf \U$17823 ( \23659 , \22382 );
buf \U$17824 ( \23660 , \22382 );
buf \U$17825 ( \23661 , \22382 );
buf \U$17826 ( \23662 , \22382 );
buf \U$17827 ( \23663 , \22382 );
buf \U$17828 ( \23664 , \22382 );
buf \U$17829 ( \23665 , \22382 );
buf \U$17830 ( \23666 , \22382 );
buf \U$17831 ( \23667 , \22382 );
buf \U$17832 ( \23668 , \22382 );
buf \U$17833 ( \23669 , \22382 );
buf \U$17834 ( \23670 , \22382 );
buf \U$17835 ( \23671 , \22382 );
buf \U$17836 ( \23672 , \22382 );
nor \U$17837 ( \23673 , \22410 , \22370 , \22412 , \22413 , \22375 , \22379 , \22382 , \23648 , \23649 , \23650 , \23651 , \23652 , \23653 , \23654 , \23655 , \23656 , \23657 , \23658 , \23659 , \23660 , \23661 , \23662 , \23663 , \23664 , \23665 , \23666 , \23667 , \23668 , \23669 , \23670 , \23671 , \23672 );
and \U$17838 ( \23674 , \8673 , \23673 );
buf \U$17839 ( \23675 , \22382 );
buf \U$17840 ( \23676 , \22382 );
buf \U$17841 ( \23677 , \22382 );
buf \U$17842 ( \23678 , \22382 );
buf \U$17843 ( \23679 , \22382 );
buf \U$17844 ( \23680 , \22382 );
buf \U$17845 ( \23681 , \22382 );
buf \U$17846 ( \23682 , \22382 );
buf \U$17847 ( \23683 , \22382 );
buf \U$17848 ( \23684 , \22382 );
buf \U$17849 ( \23685 , \22382 );
buf \U$17850 ( \23686 , \22382 );
buf \U$17851 ( \23687 , \22382 );
buf \U$17852 ( \23688 , \22382 );
buf \U$17853 ( \23689 , \22382 );
buf \U$17854 ( \23690 , \22382 );
buf \U$17855 ( \23691 , \22382 );
buf \U$17856 ( \23692 , \22382 );
buf \U$17857 ( \23693 , \22382 );
buf \U$17858 ( \23694 , \22382 );
buf \U$17859 ( \23695 , \22382 );
buf \U$17860 ( \23696 , \22382 );
buf \U$17861 ( \23697 , \22382 );
buf \U$17862 ( \23698 , \22382 );
buf \U$17863 ( \23699 , \22382 );
nor \U$17864 ( \23700 , \22369 , \22370 , \22412 , \22413 , \22375 , \22379 , \22382 , \23675 , \23676 , \23677 , \23678 , \23679 , \23680 , \23681 , \23682 , \23683 , \23684 , \23685 , \23686 , \23687 , \23688 , \23689 , \23690 , \23691 , \23692 , \23693 , \23694 , \23695 , \23696 , \23697 , \23698 , \23699 );
and \U$17865 ( \23701 , \8701 , \23700 );
buf \U$17866 ( \23702 , \22382 );
buf \U$17867 ( \23703 , \22382 );
buf \U$17868 ( \23704 , \22382 );
buf \U$17869 ( \23705 , \22382 );
buf \U$17870 ( \23706 , \22382 );
buf \U$17871 ( \23707 , \22382 );
buf \U$17872 ( \23708 , \22382 );
buf \U$17873 ( \23709 , \22382 );
buf \U$17874 ( \23710 , \22382 );
buf \U$17875 ( \23711 , \22382 );
buf \U$17876 ( \23712 , \22382 );
buf \U$17877 ( \23713 , \22382 );
buf \U$17878 ( \23714 , \22382 );
buf \U$17879 ( \23715 , \22382 );
buf \U$17880 ( \23716 , \22382 );
buf \U$17881 ( \23717 , \22382 );
buf \U$17882 ( \23718 , \22382 );
buf \U$17883 ( \23719 , \22382 );
buf \U$17884 ( \23720 , \22382 );
buf \U$17885 ( \23721 , \22382 );
buf \U$17886 ( \23722 , \22382 );
buf \U$17887 ( \23723 , \22382 );
buf \U$17888 ( \23724 , \22382 );
buf \U$17889 ( \23725 , \22382 );
buf \U$17890 ( \23726 , \22382 );
nor \U$17891 ( \23727 , \22410 , \22411 , \22371 , \22413 , \22375 , \22379 , \22382 , \23702 , \23703 , \23704 , \23705 , \23706 , \23707 , \23708 , \23709 , \23710 , \23711 , \23712 , \23713 , \23714 , \23715 , \23716 , \23717 , \23718 , \23719 , \23720 , \23721 , \23722 , \23723 , \23724 , \23725 , \23726 );
and \U$17892 ( \23728 , \8729 , \23727 );
buf \U$17893 ( \23729 , \22382 );
buf \U$17894 ( \23730 , \22382 );
buf \U$17895 ( \23731 , \22382 );
buf \U$17896 ( \23732 , \22382 );
buf \U$17897 ( \23733 , \22382 );
buf \U$17898 ( \23734 , \22382 );
buf \U$17899 ( \23735 , \22382 );
buf \U$17900 ( \23736 , \22382 );
buf \U$17901 ( \23737 , \22382 );
buf \U$17902 ( \23738 , \22382 );
buf \U$17903 ( \23739 , \22382 );
buf \U$17904 ( \23740 , \22382 );
buf \U$17905 ( \23741 , \22382 );
buf \U$17906 ( \23742 , \22382 );
buf \U$17907 ( \23743 , \22382 );
buf \U$17908 ( \23744 , \22382 );
buf \U$17909 ( \23745 , \22382 );
buf \U$17910 ( \23746 , \22382 );
buf \U$17911 ( \23747 , \22382 );
buf \U$17912 ( \23748 , \22382 );
buf \U$17913 ( \23749 , \22382 );
buf \U$17914 ( \23750 , \22382 );
buf \U$17915 ( \23751 , \22382 );
buf \U$17916 ( \23752 , \22382 );
buf \U$17917 ( \23753 , \22382 );
nor \U$17918 ( \23754 , \22369 , \22411 , \22371 , \22413 , \22375 , \22379 , \22382 , \23729 , \23730 , \23731 , \23732 , \23733 , \23734 , \23735 , \23736 , \23737 , \23738 , \23739 , \23740 , \23741 , \23742 , \23743 , \23744 , \23745 , \23746 , \23747 , \23748 , \23749 , \23750 , \23751 , \23752 , \23753 );
and \U$17919 ( \23755 , \8757 , \23754 );
buf \U$17920 ( \23756 , \22382 );
buf \U$17921 ( \23757 , \22382 );
buf \U$17922 ( \23758 , \22382 );
buf \U$17923 ( \23759 , \22382 );
buf \U$17924 ( \23760 , \22382 );
buf \U$17925 ( \23761 , \22382 );
buf \U$17926 ( \23762 , \22382 );
buf \U$17927 ( \23763 , \22382 );
buf \U$17928 ( \23764 , \22382 );
buf \U$17929 ( \23765 , \22382 );
buf \U$17930 ( \23766 , \22382 );
buf \U$17931 ( \23767 , \22382 );
buf \U$17932 ( \23768 , \22382 );
buf \U$17933 ( \23769 , \22382 );
buf \U$17934 ( \23770 , \22382 );
buf \U$17935 ( \23771 , \22382 );
buf \U$17936 ( \23772 , \22382 );
buf \U$17937 ( \23773 , \22382 );
buf \U$17938 ( \23774 , \22382 );
buf \U$17939 ( \23775 , \22382 );
buf \U$17940 ( \23776 , \22382 );
buf \U$17941 ( \23777 , \22382 );
buf \U$17942 ( \23778 , \22382 );
buf \U$17943 ( \23779 , \22382 );
buf \U$17944 ( \23780 , \22382 );
nor \U$17945 ( \23781 , \22410 , \22370 , \22371 , \22413 , \22375 , \22379 , \22382 , \23756 , \23757 , \23758 , \23759 , \23760 , \23761 , \23762 , \23763 , \23764 , \23765 , \23766 , \23767 , \23768 , \23769 , \23770 , \23771 , \23772 , \23773 , \23774 , \23775 , \23776 , \23777 , \23778 , \23779 , \23780 );
and \U$17946 ( \23782 , \8785 , \23781 );
buf \U$17947 ( \23783 , \22382 );
buf \U$17948 ( \23784 , \22382 );
buf \U$17949 ( \23785 , \22382 );
buf \U$17950 ( \23786 , \22382 );
buf \U$17951 ( \23787 , \22382 );
buf \U$17952 ( \23788 , \22382 );
buf \U$17953 ( \23789 , \22382 );
buf \U$17954 ( \23790 , \22382 );
buf \U$17955 ( \23791 , \22382 );
buf \U$17956 ( \23792 , \22382 );
buf \U$17957 ( \23793 , \22382 );
buf \U$17958 ( \23794 , \22382 );
buf \U$17959 ( \23795 , \22382 );
buf \U$17960 ( \23796 , \22382 );
buf \U$17961 ( \23797 , \22382 );
buf \U$17962 ( \23798 , \22382 );
buf \U$17963 ( \23799 , \22382 );
buf \U$17964 ( \23800 , \22382 );
buf \U$17965 ( \23801 , \22382 );
buf \U$17966 ( \23802 , \22382 );
buf \U$17967 ( \23803 , \22382 );
buf \U$17968 ( \23804 , \22382 );
buf \U$17969 ( \23805 , \22382 );
buf \U$17970 ( \23806 , \22382 );
buf \U$17971 ( \23807 , \22382 );
nor \U$17972 ( \23808 , \22369 , \22370 , \22371 , \22413 , \22375 , \22379 , \22382 , \23783 , \23784 , \23785 , \23786 , \23787 , \23788 , \23789 , \23790 , \23791 , \23792 , \23793 , \23794 , \23795 , \23796 , \23797 , \23798 , \23799 , \23800 , \23801 , \23802 , \23803 , \23804 , \23805 , \23806 , \23807 );
and \U$17973 ( \23809 , \8813 , \23808 );
buf \U$17974 ( \23810 , \22382 );
buf \U$17975 ( \23811 , \22382 );
buf \U$17976 ( \23812 , \22382 );
buf \U$17977 ( \23813 , \22382 );
buf \U$17978 ( \23814 , \22382 );
buf \U$17979 ( \23815 , \22382 );
buf \U$17980 ( \23816 , \22382 );
buf \U$17981 ( \23817 , \22382 );
buf \U$17982 ( \23818 , \22382 );
buf \U$17983 ( \23819 , \22382 );
buf \U$17984 ( \23820 , \22382 );
buf \U$17985 ( \23821 , \22382 );
buf \U$17986 ( \23822 , \22382 );
buf \U$17987 ( \23823 , \22382 );
buf \U$17988 ( \23824 , \22382 );
buf \U$17989 ( \23825 , \22382 );
buf \U$17990 ( \23826 , \22382 );
buf \U$17991 ( \23827 , \22382 );
buf \U$17992 ( \23828 , \22382 );
buf \U$17993 ( \23829 , \22382 );
buf \U$17994 ( \23830 , \22382 );
buf \U$17995 ( \23831 , \22382 );
buf \U$17996 ( \23832 , \22382 );
buf \U$17997 ( \23833 , \22382 );
buf \U$17998 ( \23834 , \22382 );
nor \U$17999 ( \23835 , \22410 , \22411 , \22412 , \22372 , \22375 , \22379 , \22382 , \23810 , \23811 , \23812 , \23813 , \23814 , \23815 , \23816 , \23817 , \23818 , \23819 , \23820 , \23821 , \23822 , \23823 , \23824 , \23825 , \23826 , \23827 , \23828 , \23829 , \23830 , \23831 , \23832 , \23833 , \23834 );
and \U$18000 ( \23836 , \8841 , \23835 );
buf \U$18001 ( \23837 , \22382 );
buf \U$18002 ( \23838 , \22382 );
buf \U$18003 ( \23839 , \22382 );
buf \U$18004 ( \23840 , \22382 );
buf \U$18005 ( \23841 , \22382 );
buf \U$18006 ( \23842 , \22382 );
buf \U$18007 ( \23843 , \22382 );
buf \U$18008 ( \23844 , \22382 );
buf \U$18009 ( \23845 , \22382 );
buf \U$18010 ( \23846 , \22382 );
buf \U$18011 ( \23847 , \22382 );
buf \U$18012 ( \23848 , \22382 );
buf \U$18013 ( \23849 , \22382 );
buf \U$18014 ( \23850 , \22382 );
buf \U$18015 ( \23851 , \22382 );
buf \U$18016 ( \23852 , \22382 );
buf \U$18017 ( \23853 , \22382 );
buf \U$18018 ( \23854 , \22382 );
buf \U$18019 ( \23855 , \22382 );
buf \U$18020 ( \23856 , \22382 );
buf \U$18021 ( \23857 , \22382 );
buf \U$18022 ( \23858 , \22382 );
buf \U$18023 ( \23859 , \22382 );
buf \U$18024 ( \23860 , \22382 );
buf \U$18025 ( \23861 , \22382 );
nor \U$18026 ( \23862 , \22369 , \22411 , \22412 , \22372 , \22375 , \22379 , \22382 , \23837 , \23838 , \23839 , \23840 , \23841 , \23842 , \23843 , \23844 , \23845 , \23846 , \23847 , \23848 , \23849 , \23850 , \23851 , \23852 , \23853 , \23854 , \23855 , \23856 , \23857 , \23858 , \23859 , \23860 , \23861 );
and \U$18027 ( \23863 , \8869 , \23862 );
buf \U$18028 ( \23864 , \22382 );
buf \U$18029 ( \23865 , \22382 );
buf \U$18030 ( \23866 , \22382 );
buf \U$18031 ( \23867 , \22382 );
buf \U$18032 ( \23868 , \22382 );
buf \U$18033 ( \23869 , \22382 );
buf \U$18034 ( \23870 , \22382 );
buf \U$18035 ( \23871 , \22382 );
buf \U$18036 ( \23872 , \22382 );
buf \U$18037 ( \23873 , \22382 );
buf \U$18038 ( \23874 , \22382 );
buf \U$18039 ( \23875 , \22382 );
buf \U$18040 ( \23876 , \22382 );
buf \U$18041 ( \23877 , \22382 );
buf \U$18042 ( \23878 , \22382 );
buf \U$18043 ( \23879 , \22382 );
buf \U$18044 ( \23880 , \22382 );
buf \U$18045 ( \23881 , \22382 );
buf \U$18046 ( \23882 , \22382 );
buf \U$18047 ( \23883 , \22382 );
buf \U$18048 ( \23884 , \22382 );
buf \U$18049 ( \23885 , \22382 );
buf \U$18050 ( \23886 , \22382 );
buf \U$18051 ( \23887 , \22382 );
buf \U$18052 ( \23888 , \22382 );
nor \U$18053 ( \23889 , \22410 , \22370 , \22412 , \22372 , \22375 , \22379 , \22382 , \23864 , \23865 , \23866 , \23867 , \23868 , \23869 , \23870 , \23871 , \23872 , \23873 , \23874 , \23875 , \23876 , \23877 , \23878 , \23879 , \23880 , \23881 , \23882 , \23883 , \23884 , \23885 , \23886 , \23887 , \23888 );
and \U$18054 ( \23890 , \8897 , \23889 );
buf \U$18055 ( \23891 , \22382 );
buf \U$18056 ( \23892 , \22382 );
buf \U$18057 ( \23893 , \22382 );
buf \U$18058 ( \23894 , \22382 );
buf \U$18059 ( \23895 , \22382 );
buf \U$18060 ( \23896 , \22382 );
buf \U$18061 ( \23897 , \22382 );
buf \U$18062 ( \23898 , \22382 );
buf \U$18063 ( \23899 , \22382 );
buf \U$18064 ( \23900 , \22382 );
buf \U$18065 ( \23901 , \22382 );
buf \U$18066 ( \23902 , \22382 );
buf \U$18067 ( \23903 , \22382 );
buf \U$18068 ( \23904 , \22382 );
buf \U$18069 ( \23905 , \22382 );
buf \U$18070 ( \23906 , \22382 );
buf \U$18071 ( \23907 , \22382 );
buf \U$18072 ( \23908 , \22382 );
buf \U$18073 ( \23909 , \22382 );
buf \U$18074 ( \23910 , \22382 );
buf \U$18075 ( \23911 , \22382 );
buf \U$18076 ( \23912 , \22382 );
buf \U$18077 ( \23913 , \22382 );
buf \U$18078 ( \23914 , \22382 );
buf \U$18079 ( \23915 , \22382 );
nor \U$18080 ( \23916 , \22369 , \22370 , \22412 , \22372 , \22375 , \22379 , \22382 , \23891 , \23892 , \23893 , \23894 , \23895 , \23896 , \23897 , \23898 , \23899 , \23900 , \23901 , \23902 , \23903 , \23904 , \23905 , \23906 , \23907 , \23908 , \23909 , \23910 , \23911 , \23912 , \23913 , \23914 , \23915 );
and \U$18081 ( \23917 , \8925 , \23916 );
buf \U$18082 ( \23918 , \22382 );
buf \U$18083 ( \23919 , \22382 );
buf \U$18084 ( \23920 , \22382 );
buf \U$18085 ( \23921 , \22382 );
buf \U$18086 ( \23922 , \22382 );
buf \U$18087 ( \23923 , \22382 );
buf \U$18088 ( \23924 , \22382 );
buf \U$18089 ( \23925 , \22382 );
buf \U$18090 ( \23926 , \22382 );
buf \U$18091 ( \23927 , \22382 );
buf \U$18092 ( \23928 , \22382 );
buf \U$18093 ( \23929 , \22382 );
buf \U$18094 ( \23930 , \22382 );
buf \U$18095 ( \23931 , \22382 );
buf \U$18096 ( \23932 , \22382 );
buf \U$18097 ( \23933 , \22382 );
buf \U$18098 ( \23934 , \22382 );
buf \U$18099 ( \23935 , \22382 );
buf \U$18100 ( \23936 , \22382 );
buf \U$18101 ( \23937 , \22382 );
buf \U$18102 ( \23938 , \22382 );
buf \U$18103 ( \23939 , \22382 );
buf \U$18104 ( \23940 , \22382 );
buf \U$18105 ( \23941 , \22382 );
buf \U$18106 ( \23942 , \22382 );
nor \U$18107 ( \23943 , \22410 , \22411 , \22371 , \22372 , \22375 , \22379 , \22382 , \23918 , \23919 , \23920 , \23921 , \23922 , \23923 , \23924 , \23925 , \23926 , \23927 , \23928 , \23929 , \23930 , \23931 , \23932 , \23933 , \23934 , \23935 , \23936 , \23937 , \23938 , \23939 , \23940 , \23941 , \23942 );
and \U$18108 ( \23944 , \8953 , \23943 );
buf \U$18109 ( \23945 , \22382 );
buf \U$18110 ( \23946 , \22382 );
buf \U$18111 ( \23947 , \22382 );
buf \U$18112 ( \23948 , \22382 );
buf \U$18113 ( \23949 , \22382 );
buf \U$18114 ( \23950 , \22382 );
buf \U$18115 ( \23951 , \22382 );
buf \U$18116 ( \23952 , \22382 );
buf \U$18117 ( \23953 , \22382 );
buf \U$18118 ( \23954 , \22382 );
buf \U$18119 ( \23955 , \22382 );
buf \U$18120 ( \23956 , \22382 );
buf \U$18121 ( \23957 , \22382 );
buf \U$18122 ( \23958 , \22382 );
buf \U$18123 ( \23959 , \22382 );
buf \U$18124 ( \23960 , \22382 );
buf \U$18125 ( \23961 , \22382 );
buf \U$18126 ( \23962 , \22382 );
buf \U$18127 ( \23963 , \22382 );
buf \U$18128 ( \23964 , \22382 );
buf \U$18129 ( \23965 , \22382 );
buf \U$18130 ( \23966 , \22382 );
buf \U$18131 ( \23967 , \22382 );
buf \U$18132 ( \23968 , \22382 );
buf \U$18133 ( \23969 , \22382 );
nor \U$18134 ( \23970 , \22369 , \22411 , \22371 , \22372 , \22375 , \22379 , \22382 , \23945 , \23946 , \23947 , \23948 , \23949 , \23950 , \23951 , \23952 , \23953 , \23954 , \23955 , \23956 , \23957 , \23958 , \23959 , \23960 , \23961 , \23962 , \23963 , \23964 , \23965 , \23966 , \23967 , \23968 , \23969 );
and \U$18135 ( \23971 , \8981 , \23970 );
buf \U$18136 ( \23972 , \22382 );
buf \U$18137 ( \23973 , \22382 );
buf \U$18138 ( \23974 , \22382 );
buf \U$18139 ( \23975 , \22382 );
buf \U$18140 ( \23976 , \22382 );
buf \U$18141 ( \23977 , \22382 );
buf \U$18142 ( \23978 , \22382 );
buf \U$18143 ( \23979 , \22382 );
buf \U$18144 ( \23980 , \22382 );
buf \U$18145 ( \23981 , \22382 );
buf \U$18146 ( \23982 , \22382 );
buf \U$18147 ( \23983 , \22382 );
buf \U$18148 ( \23984 , \22382 );
buf \U$18149 ( \23985 , \22382 );
buf \U$18150 ( \23986 , \22382 );
buf \U$18151 ( \23987 , \22382 );
buf \U$18152 ( \23988 , \22382 );
buf \U$18153 ( \23989 , \22382 );
buf \U$18154 ( \23990 , \22382 );
buf \U$18155 ( \23991 , \22382 );
buf \U$18156 ( \23992 , \22382 );
buf \U$18157 ( \23993 , \22382 );
buf \U$18158 ( \23994 , \22382 );
buf \U$18159 ( \23995 , \22382 );
buf \U$18160 ( \23996 , \22382 );
nor \U$18161 ( \23997 , \22410 , \22370 , \22371 , \22372 , \22375 , \22379 , \22382 , \23972 , \23973 , \23974 , \23975 , \23976 , \23977 , \23978 , \23979 , \23980 , \23981 , \23982 , \23983 , \23984 , \23985 , \23986 , \23987 , \23988 , \23989 , \23990 , \23991 , \23992 , \23993 , \23994 , \23995 , \23996 );
and \U$18162 ( \23998 , \9009 , \23997 );
or \U$18163 ( \23999 , \23593 , \23620 , \23647 , \23674 , \23701 , \23728 , \23755 , \23782 , \23809 , \23836 , \23863 , \23890 , \23917 , \23944 , \23971 , \23998 );
buf \U$18164 ( \24000 , \22382 );
not \U$18165 ( \24001 , \24000 );
buf \U$18166 ( \24002 , \22370 );
buf \U$18167 ( \24003 , \22371 );
buf \U$18168 ( \24004 , \22372 );
buf \U$18169 ( \24005 , \22375 );
buf \U$18170 ( \24006 , \22379 );
buf \U$18171 ( \24007 , \22382 );
buf \U$18172 ( \24008 , \22382 );
buf \U$18173 ( \24009 , \22382 );
buf \U$18174 ( \24010 , \22382 );
buf \U$18175 ( \24011 , \22382 );
buf \U$18176 ( \24012 , \22382 );
buf \U$18177 ( \24013 , \22382 );
buf \U$18178 ( \24014 , \22382 );
buf \U$18179 ( \24015 , \22382 );
buf \U$18180 ( \24016 , \22382 );
buf \U$18181 ( \24017 , \22382 );
buf \U$18182 ( \24018 , \22382 );
buf \U$18183 ( \24019 , \22382 );
buf \U$18184 ( \24020 , \22382 );
buf \U$18185 ( \24021 , \22382 );
buf \U$18186 ( \24022 , \22382 );
buf \U$18187 ( \24023 , \22382 );
buf \U$18188 ( \24024 , \22382 );
buf \U$18189 ( \24025 , \22382 );
buf \U$18190 ( \24026 , \22382 );
buf \U$18191 ( \24027 , \22382 );
buf \U$18192 ( \24028 , \22382 );
buf \U$18193 ( \24029 , \22382 );
buf \U$18194 ( \24030 , \22382 );
buf \U$18195 ( \24031 , \22382 );
buf \U$18196 ( \24032 , \22369 );
or \U$18197 ( \24033 , \24002 , \24003 , \24004 , \24005 , \24006 , \24007 , \24008 , \24009 , \24010 , \24011 , \24012 , \24013 , \24014 , \24015 , \24016 , \24017 , \24018 , \24019 , \24020 , \24021 , \24022 , \24023 , \24024 , \24025 , \24026 , \24027 , \24028 , \24029 , \24030 , \24031 , \24032 );
nand \U$18198 ( \24034 , \24001 , \24033 );
buf \U$18199 ( \24035 , \24034 );
buf \U$18200 ( \24036 , \22382 );
not \U$18201 ( \24037 , \24036 );
buf \U$18202 ( \24038 , \22379 );
buf \U$18203 ( \24039 , \22382 );
buf \U$18204 ( \24040 , \22382 );
buf \U$18205 ( \24041 , \22382 );
buf \U$18206 ( \24042 , \22382 );
buf \U$18207 ( \24043 , \22382 );
buf \U$18208 ( \24044 , \22382 );
buf \U$18209 ( \24045 , \22382 );
buf \U$18210 ( \24046 , \22382 );
buf \U$18211 ( \24047 , \22382 );
buf \U$18212 ( \24048 , \22382 );
buf \U$18213 ( \24049 , \22382 );
buf \U$18214 ( \24050 , \22382 );
buf \U$18215 ( \24051 , \22382 );
buf \U$18216 ( \24052 , \22382 );
buf \U$18217 ( \24053 , \22382 );
buf \U$18218 ( \24054 , \22382 );
buf \U$18219 ( \24055 , \22382 );
buf \U$18220 ( \24056 , \22382 );
buf \U$18221 ( \24057 , \22382 );
buf \U$18222 ( \24058 , \22382 );
buf \U$18223 ( \24059 , \22382 );
buf \U$18224 ( \24060 , \22382 );
buf \U$18225 ( \24061 , \22382 );
buf \U$18226 ( \24062 , \22382 );
buf \U$18227 ( \24063 , \22382 );
buf \U$18228 ( \24064 , \22375 );
buf \U$18229 ( \24065 , \22369 );
buf \U$18230 ( \24066 , \22370 );
buf \U$18231 ( \24067 , \22371 );
buf \U$18232 ( \24068 , \22372 );
or \U$18233 ( \24069 , \24065 , \24066 , \24067 , \24068 );
and \U$18234 ( \24070 , \24064 , \24069 );
or \U$18235 ( \24071 , \24038 , \24039 , \24040 , \24041 , \24042 , \24043 , \24044 , \24045 , \24046 , \24047 , \24048 , \24049 , \24050 , \24051 , \24052 , \24053 , \24054 , \24055 , \24056 , \24057 , \24058 , \24059 , \24060 , \24061 , \24062 , \24063 , \24070 );
and \U$18236 ( \24072 , \24037 , \24071 );
buf \U$18237 ( \24073 , \24072 );
or \U$18238 ( \24074 , \24035 , \24073 );
_DC g74fb ( \24075_nG74fb , \23999 , \24074 );
buf \U$18239 ( \24076 , \24075_nG74fb );
xor \U$18240 ( \24077 , \23566 , \24076 );
buf \U$18241 ( \24078 , RIb7af5b8_255);
and \U$18242 ( \24079 , \7207 , \23592 );
and \U$18243 ( \24080 , \7209 , \23619 );
and \U$18244 ( \24081 , \9119 , \23646 );
and \U$18245 ( \24082 , \9121 , \23673 );
and \U$18246 ( \24083 , \9123 , \23700 );
and \U$18247 ( \24084 , \9125 , \23727 );
and \U$18248 ( \24085 , \9127 , \23754 );
and \U$18249 ( \24086 , \9129 , \23781 );
and \U$18250 ( \24087 , \9131 , \23808 );
and \U$18251 ( \24088 , \9133 , \23835 );
and \U$18252 ( \24089 , \9135 , \23862 );
and \U$18253 ( \24090 , \9137 , \23889 );
and \U$18254 ( \24091 , \9139 , \23916 );
and \U$18255 ( \24092 , \9141 , \23943 );
and \U$18256 ( \24093 , \9143 , \23970 );
and \U$18257 ( \24094 , \9145 , \23997 );
or \U$18258 ( \24095 , \24079 , \24080 , \24081 , \24082 , \24083 , \24084 , \24085 , \24086 , \24087 , \24088 , \24089 , \24090 , \24091 , \24092 , \24093 , \24094 );
_DC g7510 ( \24096_nG7510 , \24095 , \24074 );
buf \U$18259 ( \24097 , \24096_nG7510 );
xor \U$18260 ( \24098 , \24078 , \24097 );
or \U$18261 ( \24099 , \24077 , \24098 );
buf \U$18262 ( \24100 , RIb7af540_256);
and \U$18263 ( \24101 , \7217 , \23592 );
and \U$18264 ( \24102 , \7219 , \23619 );
and \U$18265 ( \24103 , \9155 , \23646 );
and \U$18266 ( \24104 , \9157 , \23673 );
and \U$18267 ( \24105 , \9159 , \23700 );
and \U$18268 ( \24106 , \9161 , \23727 );
and \U$18269 ( \24107 , \9163 , \23754 );
and \U$18270 ( \24108 , \9165 , \23781 );
and \U$18271 ( \24109 , \9167 , \23808 );
and \U$18272 ( \24110 , \9169 , \23835 );
and \U$18273 ( \24111 , \9171 , \23862 );
and \U$18274 ( \24112 , \9173 , \23889 );
and \U$18275 ( \24113 , \9175 , \23916 );
and \U$18276 ( \24114 , \9177 , \23943 );
and \U$18277 ( \24115 , \9179 , \23970 );
and \U$18278 ( \24116 , \9181 , \23997 );
or \U$18279 ( \24117 , \24101 , \24102 , \24103 , \24104 , \24105 , \24106 , \24107 , \24108 , \24109 , \24110 , \24111 , \24112 , \24113 , \24114 , \24115 , \24116 );
_DC g7526 ( \24118_nG7526 , \24117 , \24074 );
buf \U$18280 ( \24119 , \24118_nG7526 );
xor \U$18281 ( \24120 , \24100 , \24119 );
or \U$18282 ( \24121 , \24099 , \24120 );
buf \U$18283 ( \24122 , RIb7af4c8_257);
and \U$18284 ( \24123 , \7227 , \23592 );
and \U$18285 ( \24124 , \7229 , \23619 );
and \U$18286 ( \24125 , \9191 , \23646 );
and \U$18287 ( \24126 , \9193 , \23673 );
and \U$18288 ( \24127 , \9195 , \23700 );
and \U$18289 ( \24128 , \9197 , \23727 );
and \U$18290 ( \24129 , \9199 , \23754 );
and \U$18291 ( \24130 , \9201 , \23781 );
and \U$18292 ( \24131 , \9203 , \23808 );
and \U$18293 ( \24132 , \9205 , \23835 );
and \U$18294 ( \24133 , \9207 , \23862 );
and \U$18295 ( \24134 , \9209 , \23889 );
and \U$18296 ( \24135 , \9211 , \23916 );
and \U$18297 ( \24136 , \9213 , \23943 );
and \U$18298 ( \24137 , \9215 , \23970 );
and \U$18299 ( \24138 , \9217 , \23997 );
or \U$18300 ( \24139 , \24123 , \24124 , \24125 , \24126 , \24127 , \24128 , \24129 , \24130 , \24131 , \24132 , \24133 , \24134 , \24135 , \24136 , \24137 , \24138 );
_DC g753c ( \24140_nG753c , \24139 , \24074 );
buf \U$18301 ( \24141 , \24140_nG753c );
xor \U$18302 ( \24142 , \24122 , \24141 );
or \U$18303 ( \24143 , \24121 , \24142 );
buf \U$18304 ( \24144 , RIb7af450_258);
and \U$18305 ( \24145 , \7237 , \23592 );
and \U$18306 ( \24146 , \7239 , \23619 );
and \U$18307 ( \24147 , \9227 , \23646 );
and \U$18308 ( \24148 , \9229 , \23673 );
and \U$18309 ( \24149 , \9231 , \23700 );
and \U$18310 ( \24150 , \9233 , \23727 );
and \U$18311 ( \24151 , \9235 , \23754 );
and \U$18312 ( \24152 , \9237 , \23781 );
and \U$18313 ( \24153 , \9239 , \23808 );
and \U$18314 ( \24154 , \9241 , \23835 );
and \U$18315 ( \24155 , \9243 , \23862 );
and \U$18316 ( \24156 , \9245 , \23889 );
and \U$18317 ( \24157 , \9247 , \23916 );
and \U$18318 ( \24158 , \9249 , \23943 );
and \U$18319 ( \24159 , \9251 , \23970 );
and \U$18320 ( \24160 , \9253 , \23997 );
or \U$18321 ( \24161 , \24145 , \24146 , \24147 , \24148 , \24149 , \24150 , \24151 , \24152 , \24153 , \24154 , \24155 , \24156 , \24157 , \24158 , \24159 , \24160 );
_DC g7552 ( \24162_nG7552 , \24161 , \24074 );
buf \U$18322 ( \24163 , \24162_nG7552 );
xor \U$18323 ( \24164 , \24144 , \24163 );
or \U$18324 ( \24165 , \24143 , \24164 );
buf \U$18325 ( \24166 , RIb7af3d8_259);
and \U$18326 ( \24167 , \7247 , \23592 );
and \U$18327 ( \24168 , \7249 , \23619 );
and \U$18328 ( \24169 , \9263 , \23646 );
and \U$18329 ( \24170 , \9265 , \23673 );
and \U$18330 ( \24171 , \9267 , \23700 );
and \U$18331 ( \24172 , \9269 , \23727 );
and \U$18332 ( \24173 , \9271 , \23754 );
and \U$18333 ( \24174 , \9273 , \23781 );
and \U$18334 ( \24175 , \9275 , \23808 );
and \U$18335 ( \24176 , \9277 , \23835 );
and \U$18336 ( \24177 , \9279 , \23862 );
and \U$18337 ( \24178 , \9281 , \23889 );
and \U$18338 ( \24179 , \9283 , \23916 );
and \U$18339 ( \24180 , \9285 , \23943 );
and \U$18340 ( \24181 , \9287 , \23970 );
and \U$18341 ( \24182 , \9289 , \23997 );
or \U$18342 ( \24183 , \24167 , \24168 , \24169 , \24170 , \24171 , \24172 , \24173 , \24174 , \24175 , \24176 , \24177 , \24178 , \24179 , \24180 , \24181 , \24182 );
_DC g7568 ( \24184_nG7568 , \24183 , \24074 );
buf \U$18343 ( \24185 , \24184_nG7568 );
xor \U$18344 ( \24186 , \24166 , \24185 );
or \U$18345 ( \24187 , \24165 , \24186 );
buf \U$18346 ( \24188 , RIb7a5bf8_260);
and \U$18347 ( \24189 , \7257 , \23592 );
and \U$18348 ( \24190 , \7259 , \23619 );
and \U$18349 ( \24191 , \9299 , \23646 );
and \U$18350 ( \24192 , \9301 , \23673 );
and \U$18351 ( \24193 , \9303 , \23700 );
and \U$18352 ( \24194 , \9305 , \23727 );
and \U$18353 ( \24195 , \9307 , \23754 );
and \U$18354 ( \24196 , \9309 , \23781 );
and \U$18355 ( \24197 , \9311 , \23808 );
and \U$18356 ( \24198 , \9313 , \23835 );
and \U$18357 ( \24199 , \9315 , \23862 );
and \U$18358 ( \24200 , \9317 , \23889 );
and \U$18359 ( \24201 , \9319 , \23916 );
and \U$18360 ( \24202 , \9321 , \23943 );
and \U$18361 ( \24203 , \9323 , \23970 );
and \U$18362 ( \24204 , \9325 , \23997 );
or \U$18363 ( \24205 , \24189 , \24190 , \24191 , \24192 , \24193 , \24194 , \24195 , \24196 , \24197 , \24198 , \24199 , \24200 , \24201 , \24202 , \24203 , \24204 );
_DC g757e ( \24206_nG757e , \24205 , \24074 );
buf \U$18364 ( \24207 , \24206_nG757e );
xor \U$18365 ( \24208 , \24188 , \24207 );
or \U$18366 ( \24209 , \24187 , \24208 );
buf \U$18367 ( \24210 , RIb7a0c48_261);
and \U$18368 ( \24211 , \7267 , \23592 );
and \U$18369 ( \24212 , \7269 , \23619 );
and \U$18370 ( \24213 , \9335 , \23646 );
and \U$18371 ( \24214 , \9337 , \23673 );
and \U$18372 ( \24215 , \9339 , \23700 );
and \U$18373 ( \24216 , \9341 , \23727 );
and \U$18374 ( \24217 , \9343 , \23754 );
and \U$18375 ( \24218 , \9345 , \23781 );
and \U$18376 ( \24219 , \9347 , \23808 );
and \U$18377 ( \24220 , \9349 , \23835 );
and \U$18378 ( \24221 , \9351 , \23862 );
and \U$18379 ( \24222 , \9353 , \23889 );
and \U$18380 ( \24223 , \9355 , \23916 );
and \U$18381 ( \24224 , \9357 , \23943 );
and \U$18382 ( \24225 , \9359 , \23970 );
and \U$18383 ( \24226 , \9361 , \23997 );
or \U$18384 ( \24227 , \24211 , \24212 , \24213 , \24214 , \24215 , \24216 , \24217 , \24218 , \24219 , \24220 , \24221 , \24222 , \24223 , \24224 , \24225 , \24226 );
_DC g7594 ( \24228_nG7594 , \24227 , \24074 );
buf \U$18385 ( \24229 , \24228_nG7594 );
xor \U$18386 ( \24230 , \24210 , \24229 );
or \U$18387 ( \24231 , \24209 , \24230 );
not \U$18388 ( \24232 , \24231 );
buf \U$18389 ( \24233 , \24232 );
and \U$18390 ( \24234 , \23565 , \24233 );
_HMUX g759b ( \24235_nG759b , \22072_nG6d1d , \22369 , \24234 );
buf \U$18391 ( \24236 , \22087 );
buf \U$18392 ( \24237 , \22084 );
buf \U$18393 ( \24238 , \22074 );
buf \U$18394 ( \24239 , \22076 );
buf \U$18395 ( \24240 , \22078 );
buf \U$18396 ( \24241 , \22081 );
or \U$18397 ( \24242 , \24238 , \24239 , \24240 , \24241 );
and \U$18398 ( \24243 , \24237 , \24242 );
or \U$18399 ( \24244 , \24236 , \24243 );
buf \U$18400 ( \24245 , \24244 );
_HMUX g75a6 ( \24246_nG75a6 , \22368_nG6e48 , \24235_nG759b , \24245 );
buf \U$18401 ( \24247 , RIe5319e0_6884);
not \U$18402 ( \24248 , \24247 );
buf \U$18403 ( \24249 , \24248 );
buf \U$18404 ( \24250 , RIe549ef0_6842);
xnor \U$18405 ( \24251 , \24250 , \24247 );
buf \U$18406 ( \24252 , \24251 );
buf \U$18407 ( \24253 , RIe549770_6843);
or \U$18408 ( \24254 , \24250 , \24247 );
xnor \U$18409 ( \24255 , \24253 , \24254 );
buf \U$18410 ( \24256 , \24255 );
buf \U$18411 ( \24257 , RIe548ff0_6844);
or \U$18412 ( \24258 , \24253 , \24254 );
xor \U$18413 ( \24259 , \24257 , \24258 );
buf \U$18414 ( \24260 , \24259 );
buf \U$18415 ( \24261 , RIea91330_6888);
and \U$18416 ( \24262 , \24257 , \24258 );
xor \U$18417 ( \24263 , \24261 , \24262 );
buf \U$18418 ( \24264 , \24263 );
not \U$18419 ( \24265 , \24264 );
and \U$18420 ( \24266 , \24261 , \24262 );
buf \U$18421 ( \24267 , \24266 );
nor \U$18422 ( \24268 , \24249 , \24252 , \24256 , \24260 , \24265 , \24267 );
and \U$18423 ( \24269 , RIe5329d0_6883, \24268 );
not \U$18424 ( \24270 , \24267 );
and \U$18425 ( \24271 , \24249 , \24252 , \24256 , \24260 , \24265 , \24270 );
and \U$18426 ( \24272 , RIeb72150_6905, \24271 );
not \U$18427 ( \24273 , \24249 );
and \U$18428 ( \24274 , \24273 , \24252 , \24256 , \24260 , \24265 , \24270 );
and \U$18429 ( \24275 , RIeab80c0_6897, \24274 );
not \U$18430 ( \24276 , \24252 );
and \U$18431 ( \24277 , \24249 , \24276 , \24256 , \24260 , \24265 , \24270 );
and \U$18432 ( \24278 , RIe5331c8_6882, \24277 );
and \U$18433 ( \24279 , \24273 , \24276 , \24256 , \24260 , \24265 , \24270 );
and \U$18434 ( \24280 , RIe5339c0_6881, \24279 );
not \U$18435 ( \24281 , \24256 );
and \U$18436 ( \24282 , \24249 , \24252 , \24281 , \24260 , \24265 , \24270 );
and \U$18437 ( \24283 , RIeab87c8_6898, \24282 );
and \U$18438 ( \24284 , \24273 , \24252 , \24281 , \24260 , \24265 , \24270 );
and \U$18439 ( \24285 , RIe5341b8_6880, \24284 );
and \U$18440 ( \24286 , \24249 , \24276 , \24281 , \24260 , \24265 , \24270 );
and \U$18441 ( \24287 , RIe5349b0_6879, \24286 );
and \U$18442 ( \24288 , \24273 , \24276 , \24281 , \24260 , \24265 , \24270 );
and \U$18443 ( \24289 , RIea94af8_6890, \24288 );
nor \U$18444 ( \24290 , \24273 , \24276 , \24281 , \24260 , \24264 , \24267 );
and \U$18445 ( \24291 , RIe5351a8_6878, \24290 );
or \U$18452 ( \24292 , \24269 , \24272 , \24275 , \24278 , \24280 , \24283 , \24285 , \24287 , \24289 , \24291 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
buf \U$18454 ( \24293 , \24267 );
buf \U$18455 ( \24294 , \24264 );
buf \U$18456 ( \24295 , \24249 );
buf \U$18457 ( \24296 , \24252 );
buf \U$18458 ( \24297 , \24256 );
buf \U$18459 ( \24298 , \24260 );
or \U$18460 ( \24299 , \24295 , \24296 , \24297 , \24298 );
and \U$18461 ( \24300 , \24294 , \24299 );
or \U$18462 ( \24301 , \24293 , \24300 );
buf \U$18463 ( \24302 , \24301 );
or \U$18464 ( \24303 , 1'b0 , \24302 );
_DC g75e0 ( \24304_nG75e0 , \24292 , \24303 );
not \U$18465 ( \24305 , \24304_nG75e0 );
buf \U$18466 ( \24306 , RIb7b9608_246);
and \U$18467 ( \24307 , \7117 , \24268 );
and \U$18468 ( \24308 , \7119 , \24271 );
and \U$18469 ( \24309 , \7864 , \24274 );
and \U$18470 ( \24310 , \7892 , \24277 );
and \U$18471 ( \24311 , \7920 , \24279 );
and \U$18472 ( \24312 , \7948 , \24282 );
and \U$18473 ( \24313 , \7976 , \24284 );
and \U$18474 ( \24314 , \8004 , \24286 );
and \U$18475 ( \24315 , \8032 , \24288 );
and \U$18476 ( \24316 , \8060 , \24290 );
or \U$18483 ( \24317 , \24307 , \24308 , \24309 , \24310 , \24311 , \24312 , \24313 , \24314 , \24315 , \24316 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g75ee ( \24318_nG75ee , \24317 , \24303 );
buf \U$18484 ( \24319 , \24318_nG75ee );
xor \U$18485 ( \24320 , \24306 , \24319 );
buf \U$18486 ( \24321 , RIb7b9590_247);
and \U$18487 ( \24322 , \7126 , \24268 );
and \U$18488 ( \24323 , \7128 , \24271 );
and \U$18489 ( \24324 , \8338 , \24274 );
and \U$18490 ( \24325 , \8340 , \24277 );
and \U$18491 ( \24326 , \8342 , \24279 );
and \U$18492 ( \24327 , \8344 , \24282 );
and \U$18493 ( \24328 , \8346 , \24284 );
and \U$18494 ( \24329 , \8348 , \24286 );
and \U$18495 ( \24330 , \8350 , \24288 );
and \U$18496 ( \24331 , \8352 , \24290 );
or \U$18503 ( \24332 , \24322 , \24323 , \24324 , \24325 , \24326 , \24327 , \24328 , \24329 , \24330 , \24331 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g75fd ( \24333_nG75fd , \24332 , \24303 );
buf \U$18504 ( \24334 , \24333_nG75fd );
xor \U$18505 ( \24335 , \24321 , \24334 );
or \U$18506 ( \24336 , \24320 , \24335 );
buf \U$18507 ( \24337 , RIb7b9518_248);
and \U$18508 ( \24338 , \7136 , \24268 );
and \U$18509 ( \24339 , \7138 , \24271 );
and \U$18510 ( \24340 , \8374 , \24274 );
and \U$18511 ( \24341 , \8376 , \24277 );
and \U$18512 ( \24342 , \8378 , \24279 );
and \U$18513 ( \24343 , \8380 , \24282 );
and \U$18514 ( \24344 , \8382 , \24284 );
and \U$18515 ( \24345 , \8384 , \24286 );
and \U$18516 ( \24346 , \8386 , \24288 );
and \U$18517 ( \24347 , \8388 , \24290 );
or \U$18524 ( \24348 , \24338 , \24339 , \24340 , \24341 , \24342 , \24343 , \24344 , \24345 , \24346 , \24347 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g760d ( \24349_nG760d , \24348 , \24303 );
buf \U$18525 ( \24350 , \24349_nG760d );
xor \U$18526 ( \24351 , \24337 , \24350 );
or \U$18527 ( \24352 , \24336 , \24351 );
buf \U$18528 ( \24353 , RIb7b94a0_249);
and \U$18529 ( \24354 , \7146 , \24268 );
and \U$18530 ( \24355 , \7148 , \24271 );
and \U$18531 ( \24356 , \8410 , \24274 );
and \U$18532 ( \24357 , \8412 , \24277 );
and \U$18533 ( \24358 , \8414 , \24279 );
and \U$18534 ( \24359 , \8416 , \24282 );
and \U$18535 ( \24360 , \8418 , \24284 );
and \U$18536 ( \24361 , \8420 , \24286 );
and \U$18537 ( \24362 , \8422 , \24288 );
and \U$18538 ( \24363 , \8424 , \24290 );
or \U$18545 ( \24364 , \24354 , \24355 , \24356 , \24357 , \24358 , \24359 , \24360 , \24361 , \24362 , \24363 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g761d ( \24365_nG761d , \24364 , \24303 );
buf \U$18546 ( \24366 , \24365_nG761d );
xor \U$18547 ( \24367 , \24353 , \24366 );
or \U$18548 ( \24368 , \24352 , \24367 );
buf \U$18549 ( \24369 , RIb7b9428_250);
and \U$18550 ( \24370 , \7156 , \24268 );
and \U$18551 ( \24371 , \7158 , \24271 );
and \U$18552 ( \24372 , \8446 , \24274 );
and \U$18553 ( \24373 , \8448 , \24277 );
and \U$18554 ( \24374 , \8450 , \24279 );
and \U$18555 ( \24375 , \8452 , \24282 );
and \U$18556 ( \24376 , \8454 , \24284 );
and \U$18557 ( \24377 , \8456 , \24286 );
and \U$18558 ( \24378 , \8458 , \24288 );
and \U$18559 ( \24379 , \8460 , \24290 );
or \U$18566 ( \24380 , \24370 , \24371 , \24372 , \24373 , \24374 , \24375 , \24376 , \24377 , \24378 , \24379 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g762d ( \24381_nG762d , \24380 , \24303 );
buf \U$18567 ( \24382 , \24381_nG762d );
xor \U$18568 ( \24383 , \24369 , \24382 );
or \U$18569 ( \24384 , \24368 , \24383 );
buf \U$18570 ( \24385 , RIb7b93b0_251);
and \U$18571 ( \24386 , \7166 , \24268 );
and \U$18572 ( \24387 , \7168 , \24271 );
and \U$18573 ( \24388 , \8482 , \24274 );
and \U$18574 ( \24389 , \8484 , \24277 );
and \U$18575 ( \24390 , \8486 , \24279 );
and \U$18576 ( \24391 , \8488 , \24282 );
and \U$18577 ( \24392 , \8490 , \24284 );
and \U$18578 ( \24393 , \8492 , \24286 );
and \U$18579 ( \24394 , \8494 , \24288 );
and \U$18580 ( \24395 , \8496 , \24290 );
or \U$18587 ( \24396 , \24386 , \24387 , \24388 , \24389 , \24390 , \24391 , \24392 , \24393 , \24394 , \24395 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g763d ( \24397_nG763d , \24396 , \24303 );
buf \U$18588 ( \24398 , \24397_nG763d );
xor \U$18589 ( \24399 , \24385 , \24398 );
or \U$18590 ( \24400 , \24384 , \24399 );
buf \U$18591 ( \24401 , RIb7af720_252);
and \U$18592 ( \24402 , \7176 , \24268 );
and \U$18593 ( \24403 , \7178 , \24271 );
and \U$18594 ( \24404 , \8518 , \24274 );
and \U$18595 ( \24405 , \8520 , \24277 );
and \U$18596 ( \24406 , \8522 , \24279 );
and \U$18597 ( \24407 , \8524 , \24282 );
and \U$18598 ( \24408 , \8526 , \24284 );
and \U$18599 ( \24409 , \8528 , \24286 );
and \U$18600 ( \24410 , \8530 , \24288 );
and \U$18601 ( \24411 , \8532 , \24290 );
or \U$18608 ( \24412 , \24402 , \24403 , \24404 , \24405 , \24406 , \24407 , \24408 , \24409 , \24410 , \24411 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g764d ( \24413_nG764d , \24412 , \24303 );
buf \U$18609 ( \24414 , \24413_nG764d );
xor \U$18610 ( \24415 , \24401 , \24414 );
or \U$18611 ( \24416 , \24400 , \24415 );
buf \U$18612 ( \24417 , RIb7af6a8_253);
and \U$18613 ( \24418 , \7186 , \24268 );
and \U$18614 ( \24419 , \7188 , \24271 );
and \U$18615 ( \24420 , \8554 , \24274 );
and \U$18616 ( \24421 , \8556 , \24277 );
and \U$18617 ( \24422 , \8558 , \24279 );
and \U$18618 ( \24423 , \8560 , \24282 );
and \U$18619 ( \24424 , \8562 , \24284 );
and \U$18620 ( \24425 , \8564 , \24286 );
and \U$18621 ( \24426 , \8566 , \24288 );
and \U$18622 ( \24427 , \8568 , \24290 );
or \U$18629 ( \24428 , \24418 , \24419 , \24420 , \24421 , \24422 , \24423 , \24424 , \24425 , \24426 , \24427 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g765d ( \24429_nG765d , \24428 , \24303 );
buf \U$18630 ( \24430 , \24429_nG765d );
xor \U$18631 ( \24431 , \24417 , \24430 );
or \U$18632 ( \24432 , \24416 , \24431 );
not \U$18633 ( \24433 , \24432 );
buf \U$18634 ( \24434 , \24433 );
buf \U$18635 ( \24435 , RIb7af630_254);
and \U$18636 ( \24436 , \7198 , \24268 );
and \U$18637 ( \24437 , \7200 , \24271 );
and \U$18638 ( \24438 , \8645 , \24274 );
and \U$18639 ( \24439 , \8673 , \24277 );
and \U$18640 ( \24440 , \8701 , \24279 );
and \U$18641 ( \24441 , \8729 , \24282 );
and \U$18642 ( \24442 , \8757 , \24284 );
and \U$18643 ( \24443 , \8785 , \24286 );
and \U$18644 ( \24444 , \8813 , \24288 );
and \U$18645 ( \24445 , \8841 , \24290 );
or \U$18652 ( \24446 , \24436 , \24437 , \24438 , \24439 , \24440 , \24441 , \24442 , \24443 , \24444 , \24445 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g766f ( \24447_nG766f , \24446 , \24303 );
buf \U$18653 ( \24448 , \24447_nG766f );
xor \U$18654 ( \24449 , \24435 , \24448 );
buf \U$18655 ( \24450 , RIb7af5b8_255);
and \U$18656 ( \24451 , \7207 , \24268 );
and \U$18657 ( \24452 , \7209 , \24271 );
and \U$18658 ( \24453 , \9119 , \24274 );
and \U$18659 ( \24454 , \9121 , \24277 );
and \U$18660 ( \24455 , \9123 , \24279 );
and \U$18661 ( \24456 , \9125 , \24282 );
and \U$18662 ( \24457 , \9127 , \24284 );
and \U$18663 ( \24458 , \9129 , \24286 );
and \U$18664 ( \24459 , \9131 , \24288 );
and \U$18665 ( \24460 , \9133 , \24290 );
or \U$18672 ( \24461 , \24451 , \24452 , \24453 , \24454 , \24455 , \24456 , \24457 , \24458 , \24459 , \24460 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g767e ( \24462_nG767e , \24461 , \24303 );
buf \U$18673 ( \24463 , \24462_nG767e );
xor \U$18674 ( \24464 , \24450 , \24463 );
or \U$18675 ( \24465 , \24449 , \24464 );
buf \U$18676 ( \24466 , RIb7af540_256);
and \U$18677 ( \24467 , \7217 , \24268 );
and \U$18678 ( \24468 , \7219 , \24271 );
and \U$18679 ( \24469 , \9155 , \24274 );
and \U$18680 ( \24470 , \9157 , \24277 );
and \U$18681 ( \24471 , \9159 , \24279 );
and \U$18682 ( \24472 , \9161 , \24282 );
and \U$18683 ( \24473 , \9163 , \24284 );
and \U$18684 ( \24474 , \9165 , \24286 );
and \U$18685 ( \24475 , \9167 , \24288 );
and \U$18686 ( \24476 , \9169 , \24290 );
or \U$18693 ( \24477 , \24467 , \24468 , \24469 , \24470 , \24471 , \24472 , \24473 , \24474 , \24475 , \24476 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g768e ( \24478_nG768e , \24477 , \24303 );
buf \U$18694 ( \24479 , \24478_nG768e );
xor \U$18695 ( \24480 , \24466 , \24479 );
or \U$18696 ( \24481 , \24465 , \24480 );
buf \U$18697 ( \24482 , RIb7af4c8_257);
and \U$18698 ( \24483 , \7227 , \24268 );
and \U$18699 ( \24484 , \7229 , \24271 );
and \U$18700 ( \24485 , \9191 , \24274 );
and \U$18701 ( \24486 , \9193 , \24277 );
and \U$18702 ( \24487 , \9195 , \24279 );
and \U$18703 ( \24488 , \9197 , \24282 );
and \U$18704 ( \24489 , \9199 , \24284 );
and \U$18705 ( \24490 , \9201 , \24286 );
and \U$18706 ( \24491 , \9203 , \24288 );
and \U$18707 ( \24492 , \9205 , \24290 );
or \U$18714 ( \24493 , \24483 , \24484 , \24485 , \24486 , \24487 , \24488 , \24489 , \24490 , \24491 , \24492 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g769e ( \24494_nG769e , \24493 , \24303 );
buf \U$18715 ( \24495 , \24494_nG769e );
xor \U$18716 ( \24496 , \24482 , \24495 );
or \U$18717 ( \24497 , \24481 , \24496 );
buf \U$18718 ( \24498 , RIb7af450_258);
and \U$18719 ( \24499 , \7237 , \24268 );
and \U$18720 ( \24500 , \7239 , \24271 );
and \U$18721 ( \24501 , \9227 , \24274 );
and \U$18722 ( \24502 , \9229 , \24277 );
and \U$18723 ( \24503 , \9231 , \24279 );
and \U$18724 ( \24504 , \9233 , \24282 );
and \U$18725 ( \24505 , \9235 , \24284 );
and \U$18726 ( \24506 , \9237 , \24286 );
and \U$18727 ( \24507 , \9239 , \24288 );
and \U$18728 ( \24508 , \9241 , \24290 );
or \U$18735 ( \24509 , \24499 , \24500 , \24501 , \24502 , \24503 , \24504 , \24505 , \24506 , \24507 , \24508 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g76ae ( \24510_nG76ae , \24509 , \24303 );
buf \U$18736 ( \24511 , \24510_nG76ae );
xor \U$18737 ( \24512 , \24498 , \24511 );
or \U$18738 ( \24513 , \24497 , \24512 );
buf \U$18739 ( \24514 , RIb7af3d8_259);
and \U$18740 ( \24515 , \7247 , \24268 );
and \U$18741 ( \24516 , \7249 , \24271 );
and \U$18742 ( \24517 , \9263 , \24274 );
and \U$18743 ( \24518 , \9265 , \24277 );
and \U$18744 ( \24519 , \9267 , \24279 );
and \U$18745 ( \24520 , \9269 , \24282 );
and \U$18746 ( \24521 , \9271 , \24284 );
and \U$18747 ( \24522 , \9273 , \24286 );
and \U$18748 ( \24523 , \9275 , \24288 );
and \U$18749 ( \24524 , \9277 , \24290 );
or \U$18756 ( \24525 , \24515 , \24516 , \24517 , \24518 , \24519 , \24520 , \24521 , \24522 , \24523 , \24524 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g76be ( \24526_nG76be , \24525 , \24303 );
buf \U$18757 ( \24527 , \24526_nG76be );
xor \U$18758 ( \24528 , \24514 , \24527 );
or \U$18759 ( \24529 , \24513 , \24528 );
buf \U$18760 ( \24530 , RIb7a5bf8_260);
and \U$18761 ( \24531 , \7257 , \24268 );
and \U$18762 ( \24532 , \7259 , \24271 );
and \U$18763 ( \24533 , \9299 , \24274 );
and \U$18764 ( \24534 , \9301 , \24277 );
and \U$18765 ( \24535 , \9303 , \24279 );
and \U$18766 ( \24536 , \9305 , \24282 );
and \U$18767 ( \24537 , \9307 , \24284 );
and \U$18768 ( \24538 , \9309 , \24286 );
and \U$18769 ( \24539 , \9311 , \24288 );
and \U$18770 ( \24540 , \9313 , \24290 );
or \U$18777 ( \24541 , \24531 , \24532 , \24533 , \24534 , \24535 , \24536 , \24537 , \24538 , \24539 , \24540 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g76ce ( \24542_nG76ce , \24541 , \24303 );
buf \U$18778 ( \24543 , \24542_nG76ce );
xor \U$18779 ( \24544 , \24530 , \24543 );
or \U$18780 ( \24545 , \24529 , \24544 );
buf \U$18781 ( \24546 , RIb7a0c48_261);
and \U$18782 ( \24547 , \7267 , \24268 );
and \U$18783 ( \24548 , \7269 , \24271 );
and \U$18784 ( \24549 , \9335 , \24274 );
and \U$18785 ( \24550 , \9337 , \24277 );
and \U$18786 ( \24551 , \9339 , \24279 );
and \U$18787 ( \24552 , \9341 , \24282 );
and \U$18788 ( \24553 , \9343 , \24284 );
and \U$18789 ( \24554 , \9345 , \24286 );
and \U$18790 ( \24555 , \9347 , \24288 );
and \U$18791 ( \24556 , \9349 , \24290 );
or \U$18798 ( \24557 , \24547 , \24548 , \24549 , \24550 , \24551 , \24552 , \24553 , \24554 , \24555 , \24556 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g76de ( \24558_nG76de , \24557 , \24303 );
buf \U$18799 ( \24559 , \24558_nG76de );
xor \U$18800 ( \24560 , \24546 , \24559 );
or \U$18801 ( \24561 , \24545 , \24560 );
not \U$18802 ( \24562 , \24561 );
buf \U$18803 ( \24563 , \24562 );
and \U$18804 ( \24564 , \24434 , \24563 );
and \U$18805 ( \24565 , \24305 , \24564 );
_HMUX g76e6 ( \24566_nG76e6 , \24246_nG75a6 , \24249 , \24565 );
buf \U$18808 ( \24567 , \24249 );
buf \U$18811 ( \24568 , \24252 );
buf \U$18814 ( \24569 , \24256 );
buf \U$18817 ( \24570 , \24260 );
buf \U$18818 ( \24571 , \24264 );
not \U$18819 ( \24572 , \24571 );
buf \U$18820 ( \24573 , \24572 );
not \U$18821 ( \24574 , \24573 );
buf \U$18822 ( \24575 , \24267 );
xnor \U$18823 ( \24576 , \24575 , \24571 );
buf \U$18824 ( \24577 , \24576 );
or \U$18825 ( \24578 , \24575 , \24571 );
not \U$18826 ( \24579 , \24578 );
buf \U$18827 ( \24580 , \24579 );
buf \U$18828 ( \24581 , \24580 );
buf \U$18829 ( \24582 , \24580 );
buf \U$18830 ( \24583 , \24580 );
buf \U$18831 ( \24584 , \24580 );
buf \U$18832 ( \24585 , \24580 );
buf \U$18833 ( \24586 , \24580 );
buf \U$18834 ( \24587 , \24580 );
buf \U$18835 ( \24588 , \24580 );
buf \U$18836 ( \24589 , \24580 );
buf \U$18837 ( \24590 , \24580 );
buf \U$18838 ( \24591 , \24580 );
buf \U$18839 ( \24592 , \24580 );
buf \U$18840 ( \24593 , \24580 );
buf \U$18841 ( \24594 , \24580 );
buf \U$18842 ( \24595 , \24580 );
buf \U$18843 ( \24596 , \24580 );
buf \U$18844 ( \24597 , \24580 );
buf \U$18845 ( \24598 , \24580 );
buf \U$18846 ( \24599 , \24580 );
buf \U$18847 ( \24600 , \24580 );
buf \U$18848 ( \24601 , \24580 );
buf \U$18849 ( \24602 , \24580 );
buf \U$18850 ( \24603 , \24580 );
buf \U$18851 ( \24604 , \24580 );
buf \U$18852 ( \24605 , \24580 );
nor \U$18853 ( \24606 , \24567 , \24568 , \24569 , \24570 , \24574 , \24577 , \24580 , \24581 , \24582 , \24583 , \24584 , \24585 , \24586 , \24587 , \24588 , \24589 , \24590 , \24591 , \24592 , \24593 , \24594 , \24595 , \24596 , \24597 , \24598 , \24599 , \24600 , \24601 , \24602 , \24603 , \24604 , \24605 );
and \U$18854 ( \24607 , RIe5329d0_6883, \24606 );
not \U$18855 ( \24608 , \24567 );
not \U$18856 ( \24609 , \24568 );
not \U$18857 ( \24610 , \24569 );
not \U$18858 ( \24611 , \24570 );
buf \U$18859 ( \24612 , \24580 );
buf \U$18860 ( \24613 , \24580 );
buf \U$18861 ( \24614 , \24580 );
buf \U$18862 ( \24615 , \24580 );
buf \U$18863 ( \24616 , \24580 );
buf \U$18864 ( \24617 , \24580 );
buf \U$18865 ( \24618 , \24580 );
buf \U$18866 ( \24619 , \24580 );
buf \U$18867 ( \24620 , \24580 );
buf \U$18868 ( \24621 , \24580 );
buf \U$18869 ( \24622 , \24580 );
buf \U$18870 ( \24623 , \24580 );
buf \U$18871 ( \24624 , \24580 );
buf \U$18872 ( \24625 , \24580 );
buf \U$18873 ( \24626 , \24580 );
buf \U$18874 ( \24627 , \24580 );
buf \U$18875 ( \24628 , \24580 );
buf \U$18876 ( \24629 , \24580 );
buf \U$18877 ( \24630 , \24580 );
buf \U$18878 ( \24631 , \24580 );
buf \U$18879 ( \24632 , \24580 );
buf \U$18880 ( \24633 , \24580 );
buf \U$18881 ( \24634 , \24580 );
buf \U$18882 ( \24635 , \24580 );
buf \U$18883 ( \24636 , \24580 );
nor \U$18884 ( \24637 , \24608 , \24609 , \24610 , \24611 , \24573 , \24577 , \24580 , \24612 , \24613 , \24614 , \24615 , \24616 , \24617 , \24618 , \24619 , \24620 , \24621 , \24622 , \24623 , \24624 , \24625 , \24626 , \24627 , \24628 , \24629 , \24630 , \24631 , \24632 , \24633 , \24634 , \24635 , \24636 );
and \U$18885 ( \24638 , RIeb72150_6905, \24637 );
buf \U$18886 ( \24639 , \24580 );
buf \U$18887 ( \24640 , \24580 );
buf \U$18888 ( \24641 , \24580 );
buf \U$18889 ( \24642 , \24580 );
buf \U$18890 ( \24643 , \24580 );
buf \U$18891 ( \24644 , \24580 );
buf \U$18892 ( \24645 , \24580 );
buf \U$18893 ( \24646 , \24580 );
buf \U$18894 ( \24647 , \24580 );
buf \U$18895 ( \24648 , \24580 );
buf \U$18896 ( \24649 , \24580 );
buf \U$18897 ( \24650 , \24580 );
buf \U$18898 ( \24651 , \24580 );
buf \U$18899 ( \24652 , \24580 );
buf \U$18900 ( \24653 , \24580 );
buf \U$18901 ( \24654 , \24580 );
buf \U$18902 ( \24655 , \24580 );
buf \U$18903 ( \24656 , \24580 );
buf \U$18904 ( \24657 , \24580 );
buf \U$18905 ( \24658 , \24580 );
buf \U$18906 ( \24659 , \24580 );
buf \U$18907 ( \24660 , \24580 );
buf \U$18908 ( \24661 , \24580 );
buf \U$18909 ( \24662 , \24580 );
buf \U$18910 ( \24663 , \24580 );
nor \U$18911 ( \24664 , \24567 , \24609 , \24610 , \24611 , \24573 , \24577 , \24580 , \24639 , \24640 , \24641 , \24642 , \24643 , \24644 , \24645 , \24646 , \24647 , \24648 , \24649 , \24650 , \24651 , \24652 , \24653 , \24654 , \24655 , \24656 , \24657 , \24658 , \24659 , \24660 , \24661 , \24662 , \24663 );
and \U$18912 ( \24665 , RIeab80c0_6897, \24664 );
buf \U$18913 ( \24666 , \24580 );
buf \U$18914 ( \24667 , \24580 );
buf \U$18915 ( \24668 , \24580 );
buf \U$18916 ( \24669 , \24580 );
buf \U$18917 ( \24670 , \24580 );
buf \U$18918 ( \24671 , \24580 );
buf \U$18919 ( \24672 , \24580 );
buf \U$18920 ( \24673 , \24580 );
buf \U$18921 ( \24674 , \24580 );
buf \U$18922 ( \24675 , \24580 );
buf \U$18923 ( \24676 , \24580 );
buf \U$18924 ( \24677 , \24580 );
buf \U$18925 ( \24678 , \24580 );
buf \U$18926 ( \24679 , \24580 );
buf \U$18927 ( \24680 , \24580 );
buf \U$18928 ( \24681 , \24580 );
buf \U$18929 ( \24682 , \24580 );
buf \U$18930 ( \24683 , \24580 );
buf \U$18931 ( \24684 , \24580 );
buf \U$18932 ( \24685 , \24580 );
buf \U$18933 ( \24686 , \24580 );
buf \U$18934 ( \24687 , \24580 );
buf \U$18935 ( \24688 , \24580 );
buf \U$18936 ( \24689 , \24580 );
buf \U$18937 ( \24690 , \24580 );
nor \U$18938 ( \24691 , \24608 , \24568 , \24610 , \24611 , \24573 , \24577 , \24580 , \24666 , \24667 , \24668 , \24669 , \24670 , \24671 , \24672 , \24673 , \24674 , \24675 , \24676 , \24677 , \24678 , \24679 , \24680 , \24681 , \24682 , \24683 , \24684 , \24685 , \24686 , \24687 , \24688 , \24689 , \24690 );
and \U$18939 ( \24692 , RIe5331c8_6882, \24691 );
buf \U$18940 ( \24693 , \24580 );
buf \U$18941 ( \24694 , \24580 );
buf \U$18942 ( \24695 , \24580 );
buf \U$18943 ( \24696 , \24580 );
buf \U$18944 ( \24697 , \24580 );
buf \U$18945 ( \24698 , \24580 );
buf \U$18946 ( \24699 , \24580 );
buf \U$18947 ( \24700 , \24580 );
buf \U$18948 ( \24701 , \24580 );
buf \U$18949 ( \24702 , \24580 );
buf \U$18950 ( \24703 , \24580 );
buf \U$18951 ( \24704 , \24580 );
buf \U$18952 ( \24705 , \24580 );
buf \U$18953 ( \24706 , \24580 );
buf \U$18954 ( \24707 , \24580 );
buf \U$18955 ( \24708 , \24580 );
buf \U$18956 ( \24709 , \24580 );
buf \U$18957 ( \24710 , \24580 );
buf \U$18958 ( \24711 , \24580 );
buf \U$18959 ( \24712 , \24580 );
buf \U$18960 ( \24713 , \24580 );
buf \U$18961 ( \24714 , \24580 );
buf \U$18962 ( \24715 , \24580 );
buf \U$18963 ( \24716 , \24580 );
buf \U$18964 ( \24717 , \24580 );
nor \U$18965 ( \24718 , \24567 , \24568 , \24610 , \24611 , \24573 , \24577 , \24580 , \24693 , \24694 , \24695 , \24696 , \24697 , \24698 , \24699 , \24700 , \24701 , \24702 , \24703 , \24704 , \24705 , \24706 , \24707 , \24708 , \24709 , \24710 , \24711 , \24712 , \24713 , \24714 , \24715 , \24716 , \24717 );
and \U$18966 ( \24719 , RIe5339c0_6881, \24718 );
buf \U$18967 ( \24720 , \24580 );
buf \U$18968 ( \24721 , \24580 );
buf \U$18969 ( \24722 , \24580 );
buf \U$18970 ( \24723 , \24580 );
buf \U$18971 ( \24724 , \24580 );
buf \U$18972 ( \24725 , \24580 );
buf \U$18973 ( \24726 , \24580 );
buf \U$18974 ( \24727 , \24580 );
buf \U$18975 ( \24728 , \24580 );
buf \U$18976 ( \24729 , \24580 );
buf \U$18977 ( \24730 , \24580 );
buf \U$18978 ( \24731 , \24580 );
buf \U$18979 ( \24732 , \24580 );
buf \U$18980 ( \24733 , \24580 );
buf \U$18981 ( \24734 , \24580 );
buf \U$18982 ( \24735 , \24580 );
buf \U$18983 ( \24736 , \24580 );
buf \U$18984 ( \24737 , \24580 );
buf \U$18985 ( \24738 , \24580 );
buf \U$18986 ( \24739 , \24580 );
buf \U$18987 ( \24740 , \24580 );
buf \U$18988 ( \24741 , \24580 );
buf \U$18989 ( \24742 , \24580 );
buf \U$18990 ( \24743 , \24580 );
buf \U$18991 ( \24744 , \24580 );
nor \U$18992 ( \24745 , \24608 , \24609 , \24569 , \24611 , \24573 , \24577 , \24580 , \24720 , \24721 , \24722 , \24723 , \24724 , \24725 , \24726 , \24727 , \24728 , \24729 , \24730 , \24731 , \24732 , \24733 , \24734 , \24735 , \24736 , \24737 , \24738 , \24739 , \24740 , \24741 , \24742 , \24743 , \24744 );
and \U$18993 ( \24746 , RIeab87c8_6898, \24745 );
buf \U$18994 ( \24747 , \24580 );
buf \U$18995 ( \24748 , \24580 );
buf \U$18996 ( \24749 , \24580 );
buf \U$18997 ( \24750 , \24580 );
buf \U$18998 ( \24751 , \24580 );
buf \U$18999 ( \24752 , \24580 );
buf \U$19000 ( \24753 , \24580 );
buf \U$19001 ( \24754 , \24580 );
buf \U$19002 ( \24755 , \24580 );
buf \U$19003 ( \24756 , \24580 );
buf \U$19004 ( \24757 , \24580 );
buf \U$19005 ( \24758 , \24580 );
buf \U$19006 ( \24759 , \24580 );
buf \U$19007 ( \24760 , \24580 );
buf \U$19008 ( \24761 , \24580 );
buf \U$19009 ( \24762 , \24580 );
buf \U$19010 ( \24763 , \24580 );
buf \U$19011 ( \24764 , \24580 );
buf \U$19012 ( \24765 , \24580 );
buf \U$19013 ( \24766 , \24580 );
buf \U$19014 ( \24767 , \24580 );
buf \U$19015 ( \24768 , \24580 );
buf \U$19016 ( \24769 , \24580 );
buf \U$19017 ( \24770 , \24580 );
buf \U$19018 ( \24771 , \24580 );
nor \U$19019 ( \24772 , \24567 , \24609 , \24569 , \24611 , \24573 , \24577 , \24580 , \24747 , \24748 , \24749 , \24750 , \24751 , \24752 , \24753 , \24754 , \24755 , \24756 , \24757 , \24758 , \24759 , \24760 , \24761 , \24762 , \24763 , \24764 , \24765 , \24766 , \24767 , \24768 , \24769 , \24770 , \24771 );
and \U$19020 ( \24773 , RIe5341b8_6880, \24772 );
buf \U$19021 ( \24774 , \24580 );
buf \U$19022 ( \24775 , \24580 );
buf \U$19023 ( \24776 , \24580 );
buf \U$19024 ( \24777 , \24580 );
buf \U$19025 ( \24778 , \24580 );
buf \U$19026 ( \24779 , \24580 );
buf \U$19027 ( \24780 , \24580 );
buf \U$19028 ( \24781 , \24580 );
buf \U$19029 ( \24782 , \24580 );
buf \U$19030 ( \24783 , \24580 );
buf \U$19031 ( \24784 , \24580 );
buf \U$19032 ( \24785 , \24580 );
buf \U$19033 ( \24786 , \24580 );
buf \U$19034 ( \24787 , \24580 );
buf \U$19035 ( \24788 , \24580 );
buf \U$19036 ( \24789 , \24580 );
buf \U$19037 ( \24790 , \24580 );
buf \U$19038 ( \24791 , \24580 );
buf \U$19039 ( \24792 , \24580 );
buf \U$19040 ( \24793 , \24580 );
buf \U$19041 ( \24794 , \24580 );
buf \U$19042 ( \24795 , \24580 );
buf \U$19043 ( \24796 , \24580 );
buf \U$19044 ( \24797 , \24580 );
buf \U$19045 ( \24798 , \24580 );
nor \U$19046 ( \24799 , \24608 , \24568 , \24569 , \24611 , \24573 , \24577 , \24580 , \24774 , \24775 , \24776 , \24777 , \24778 , \24779 , \24780 , \24781 , \24782 , \24783 , \24784 , \24785 , \24786 , \24787 , \24788 , \24789 , \24790 , \24791 , \24792 , \24793 , \24794 , \24795 , \24796 , \24797 , \24798 );
and \U$19047 ( \24800 , RIe5349b0_6879, \24799 );
buf \U$19048 ( \24801 , \24580 );
buf \U$19049 ( \24802 , \24580 );
buf \U$19050 ( \24803 , \24580 );
buf \U$19051 ( \24804 , \24580 );
buf \U$19052 ( \24805 , \24580 );
buf \U$19053 ( \24806 , \24580 );
buf \U$19054 ( \24807 , \24580 );
buf \U$19055 ( \24808 , \24580 );
buf \U$19056 ( \24809 , \24580 );
buf \U$19057 ( \24810 , \24580 );
buf \U$19058 ( \24811 , \24580 );
buf \U$19059 ( \24812 , \24580 );
buf \U$19060 ( \24813 , \24580 );
buf \U$19061 ( \24814 , \24580 );
buf \U$19062 ( \24815 , \24580 );
buf \U$19063 ( \24816 , \24580 );
buf \U$19064 ( \24817 , \24580 );
buf \U$19065 ( \24818 , \24580 );
buf \U$19066 ( \24819 , \24580 );
buf \U$19067 ( \24820 , \24580 );
buf \U$19068 ( \24821 , \24580 );
buf \U$19069 ( \24822 , \24580 );
buf \U$19070 ( \24823 , \24580 );
buf \U$19071 ( \24824 , \24580 );
buf \U$19072 ( \24825 , \24580 );
nor \U$19073 ( \24826 , \24567 , \24568 , \24569 , \24611 , \24573 , \24577 , \24580 , \24801 , \24802 , \24803 , \24804 , \24805 , \24806 , \24807 , \24808 , \24809 , \24810 , \24811 , \24812 , \24813 , \24814 , \24815 , \24816 , \24817 , \24818 , \24819 , \24820 , \24821 , \24822 , \24823 , \24824 , \24825 );
and \U$19074 ( \24827 , RIea94af8_6890, \24826 );
buf \U$19075 ( \24828 , \24580 );
buf \U$19076 ( \24829 , \24580 );
buf \U$19077 ( \24830 , \24580 );
buf \U$19078 ( \24831 , \24580 );
buf \U$19079 ( \24832 , \24580 );
buf \U$19080 ( \24833 , \24580 );
buf \U$19081 ( \24834 , \24580 );
buf \U$19082 ( \24835 , \24580 );
buf \U$19083 ( \24836 , \24580 );
buf \U$19084 ( \24837 , \24580 );
buf \U$19085 ( \24838 , \24580 );
buf \U$19086 ( \24839 , \24580 );
buf \U$19087 ( \24840 , \24580 );
buf \U$19088 ( \24841 , \24580 );
buf \U$19089 ( \24842 , \24580 );
buf \U$19090 ( \24843 , \24580 );
buf \U$19091 ( \24844 , \24580 );
buf \U$19092 ( \24845 , \24580 );
buf \U$19093 ( \24846 , \24580 );
buf \U$19094 ( \24847 , \24580 );
buf \U$19095 ( \24848 , \24580 );
buf \U$19096 ( \24849 , \24580 );
buf \U$19097 ( \24850 , \24580 );
buf \U$19098 ( \24851 , \24580 );
buf \U$19099 ( \24852 , \24580 );
nor \U$19100 ( \24853 , \24608 , \24609 , \24610 , \24570 , \24573 , \24577 , \24580 , \24828 , \24829 , \24830 , \24831 , \24832 , \24833 , \24834 , \24835 , \24836 , \24837 , \24838 , \24839 , \24840 , \24841 , \24842 , \24843 , \24844 , \24845 , \24846 , \24847 , \24848 , \24849 , \24850 , \24851 , \24852 );
and \U$19101 ( \24854 , RIe5351a8_6878, \24853 );
buf \U$19102 ( \24855 , \24580 );
buf \U$19103 ( \24856 , \24580 );
buf \U$19104 ( \24857 , \24580 );
buf \U$19105 ( \24858 , \24580 );
buf \U$19106 ( \24859 , \24580 );
buf \U$19107 ( \24860 , \24580 );
buf \U$19108 ( \24861 , \24580 );
buf \U$19109 ( \24862 , \24580 );
buf \U$19110 ( \24863 , \24580 );
buf \U$19111 ( \24864 , \24580 );
buf \U$19112 ( \24865 , \24580 );
buf \U$19113 ( \24866 , \24580 );
buf \U$19114 ( \24867 , \24580 );
buf \U$19115 ( \24868 , \24580 );
buf \U$19116 ( \24869 , \24580 );
buf \U$19117 ( \24870 , \24580 );
buf \U$19118 ( \24871 , \24580 );
buf \U$19119 ( \24872 , \24580 );
buf \U$19120 ( \24873 , \24580 );
buf \U$19121 ( \24874 , \24580 );
buf \U$19122 ( \24875 , \24580 );
buf \U$19123 ( \24876 , \24580 );
buf \U$19124 ( \24877 , \24580 );
buf \U$19125 ( \24878 , \24580 );
buf \U$19126 ( \24879 , \24580 );
nor \U$19127 ( \24880 , \24567 , \24609 , \24610 , \24570 , \24573 , \24577 , \24580 , \24855 , \24856 , \24857 , \24858 , \24859 , \24860 , \24861 , \24862 , \24863 , \24864 , \24865 , \24866 , \24867 , \24868 , \24869 , \24870 , \24871 , \24872 , \24873 , \24874 , \24875 , \24876 , \24877 , \24878 , \24879 );
and \U$19128 ( \24881 , RIe5359a0_6877, \24880 );
buf \U$19129 ( \24882 , \24580 );
buf \U$19130 ( \24883 , \24580 );
buf \U$19131 ( \24884 , \24580 );
buf \U$19132 ( \24885 , \24580 );
buf \U$19133 ( \24886 , \24580 );
buf \U$19134 ( \24887 , \24580 );
buf \U$19135 ( \24888 , \24580 );
buf \U$19136 ( \24889 , \24580 );
buf \U$19137 ( \24890 , \24580 );
buf \U$19138 ( \24891 , \24580 );
buf \U$19139 ( \24892 , \24580 );
buf \U$19140 ( \24893 , \24580 );
buf \U$19141 ( \24894 , \24580 );
buf \U$19142 ( \24895 , \24580 );
buf \U$19143 ( \24896 , \24580 );
buf \U$19144 ( \24897 , \24580 );
buf \U$19145 ( \24898 , \24580 );
buf \U$19146 ( \24899 , \24580 );
buf \U$19147 ( \24900 , \24580 );
buf \U$19148 ( \24901 , \24580 );
buf \U$19149 ( \24902 , \24580 );
buf \U$19150 ( \24903 , \24580 );
buf \U$19151 ( \24904 , \24580 );
buf \U$19152 ( \24905 , \24580 );
buf \U$19153 ( \24906 , \24580 );
nor \U$19154 ( \24907 , \24608 , \24568 , \24610 , \24570 , \24573 , \24577 , \24580 , \24882 , \24883 , \24884 , \24885 , \24886 , \24887 , \24888 , \24889 , \24890 , \24891 , \24892 , \24893 , \24894 , \24895 , \24896 , \24897 , \24898 , \24899 , \24900 , \24901 , \24902 , \24903 , \24904 , \24905 , \24906 );
and \U$19155 ( \24908 , RIeab78c8_6895, \24907 );
buf \U$19156 ( \24909 , \24580 );
buf \U$19157 ( \24910 , \24580 );
buf \U$19158 ( \24911 , \24580 );
buf \U$19159 ( \24912 , \24580 );
buf \U$19160 ( \24913 , \24580 );
buf \U$19161 ( \24914 , \24580 );
buf \U$19162 ( \24915 , \24580 );
buf \U$19163 ( \24916 , \24580 );
buf \U$19164 ( \24917 , \24580 );
buf \U$19165 ( \24918 , \24580 );
buf \U$19166 ( \24919 , \24580 );
buf \U$19167 ( \24920 , \24580 );
buf \U$19168 ( \24921 , \24580 );
buf \U$19169 ( \24922 , \24580 );
buf \U$19170 ( \24923 , \24580 );
buf \U$19171 ( \24924 , \24580 );
buf \U$19172 ( \24925 , \24580 );
buf \U$19173 ( \24926 , \24580 );
buf \U$19174 ( \24927 , \24580 );
buf \U$19175 ( \24928 , \24580 );
buf \U$19176 ( \24929 , \24580 );
buf \U$19177 ( \24930 , \24580 );
buf \U$19178 ( \24931 , \24580 );
buf \U$19179 ( \24932 , \24580 );
buf \U$19180 ( \24933 , \24580 );
nor \U$19181 ( \24934 , \24567 , \24568 , \24610 , \24570 , \24573 , \24577 , \24580 , \24909 , \24910 , \24911 , \24912 , \24913 , \24914 , \24915 , \24916 , \24917 , \24918 , \24919 , \24920 , \24921 , \24922 , \24923 , \24924 , \24925 , \24926 , \24927 , \24928 , \24929 , \24930 , \24931 , \24932 , \24933 );
and \U$19182 ( \24935 , RIeab7d00_6896, \24934 );
buf \U$19183 ( \24936 , \24580 );
buf \U$19184 ( \24937 , \24580 );
buf \U$19185 ( \24938 , \24580 );
buf \U$19186 ( \24939 , \24580 );
buf \U$19187 ( \24940 , \24580 );
buf \U$19188 ( \24941 , \24580 );
buf \U$19189 ( \24942 , \24580 );
buf \U$19190 ( \24943 , \24580 );
buf \U$19191 ( \24944 , \24580 );
buf \U$19192 ( \24945 , \24580 );
buf \U$19193 ( \24946 , \24580 );
buf \U$19194 ( \24947 , \24580 );
buf \U$19195 ( \24948 , \24580 );
buf \U$19196 ( \24949 , \24580 );
buf \U$19197 ( \24950 , \24580 );
buf \U$19198 ( \24951 , \24580 );
buf \U$19199 ( \24952 , \24580 );
buf \U$19200 ( \24953 , \24580 );
buf \U$19201 ( \24954 , \24580 );
buf \U$19202 ( \24955 , \24580 );
buf \U$19203 ( \24956 , \24580 );
buf \U$19204 ( \24957 , \24580 );
buf \U$19205 ( \24958 , \24580 );
buf \U$19206 ( \24959 , \24580 );
buf \U$19207 ( \24960 , \24580 );
nor \U$19208 ( \24961 , \24608 , \24609 , \24569 , \24570 , \24573 , \24577 , \24580 , \24936 , \24937 , \24938 , \24939 , \24940 , \24941 , \24942 , \24943 , \24944 , \24945 , \24946 , \24947 , \24948 , \24949 , \24950 , \24951 , \24952 , \24953 , \24954 , \24955 , \24956 , \24957 , \24958 , \24959 , \24960 );
and \U$19209 ( \24962 , RIeacfa18_6902, \24961 );
buf \U$19210 ( \24963 , \24580 );
buf \U$19211 ( \24964 , \24580 );
buf \U$19212 ( \24965 , \24580 );
buf \U$19213 ( \24966 , \24580 );
buf \U$19214 ( \24967 , \24580 );
buf \U$19215 ( \24968 , \24580 );
buf \U$19216 ( \24969 , \24580 );
buf \U$19217 ( \24970 , \24580 );
buf \U$19218 ( \24971 , \24580 );
buf \U$19219 ( \24972 , \24580 );
buf \U$19220 ( \24973 , \24580 );
buf \U$19221 ( \24974 , \24580 );
buf \U$19222 ( \24975 , \24580 );
buf \U$19223 ( \24976 , \24580 );
buf \U$19224 ( \24977 , \24580 );
buf \U$19225 ( \24978 , \24580 );
buf \U$19226 ( \24979 , \24580 );
buf \U$19227 ( \24980 , \24580 );
buf \U$19228 ( \24981 , \24580 );
buf \U$19229 ( \24982 , \24580 );
buf \U$19230 ( \24983 , \24580 );
buf \U$19231 ( \24984 , \24580 );
buf \U$19232 ( \24985 , \24580 );
buf \U$19233 ( \24986 , \24580 );
buf \U$19234 ( \24987 , \24580 );
nor \U$19235 ( \24988 , \24567 , \24609 , \24569 , \24570 , \24573 , \24577 , \24580 , \24963 , \24964 , \24965 , \24966 , \24967 , \24968 , \24969 , \24970 , \24971 , \24972 , \24973 , \24974 , \24975 , \24976 , \24977 , \24978 , \24979 , \24980 , \24981 , \24982 , \24983 , \24984 , \24985 , \24986 , \24987 );
and \U$19236 ( \24989 , RIeab6518_6891, \24988 );
buf \U$19237 ( \24990 , \24580 );
buf \U$19238 ( \24991 , \24580 );
buf \U$19239 ( \24992 , \24580 );
buf \U$19240 ( \24993 , \24580 );
buf \U$19241 ( \24994 , \24580 );
buf \U$19242 ( \24995 , \24580 );
buf \U$19243 ( \24996 , \24580 );
buf \U$19244 ( \24997 , \24580 );
buf \U$19245 ( \24998 , \24580 );
buf \U$19246 ( \24999 , \24580 );
buf \U$19247 ( \25000 , \24580 );
buf \U$19248 ( \25001 , \24580 );
buf \U$19249 ( \25002 , \24580 );
buf \U$19250 ( \25003 , \24580 );
buf \U$19251 ( \25004 , \24580 );
buf \U$19252 ( \25005 , \24580 );
buf \U$19253 ( \25006 , \24580 );
buf \U$19254 ( \25007 , \24580 );
buf \U$19255 ( \25008 , \24580 );
buf \U$19256 ( \25009 , \24580 );
buf \U$19257 ( \25010 , \24580 );
buf \U$19258 ( \25011 , \24580 );
buf \U$19259 ( \25012 , \24580 );
buf \U$19260 ( \25013 , \24580 );
buf \U$19261 ( \25014 , \24580 );
nor \U$19262 ( \25015 , \24608 , \24568 , \24569 , \24570 , \24573 , \24577 , \24580 , \24990 , \24991 , \24992 , \24993 , \24994 , \24995 , \24996 , \24997 , \24998 , \24999 , \25000 , \25001 , \25002 , \25003 , \25004 , \25005 , \25006 , \25007 , \25008 , \25009 , \25010 , \25011 , \25012 , \25013 , \25014 );
and \U$19263 ( \25016 , RIeb352c8_6904, \25015 );
or \U$19264 ( \25017 , \24607 , \24638 , \24665 , \24692 , \24719 , \24746 , \24773 , \24800 , \24827 , \24854 , \24881 , \24908 , \24935 , \24962 , \24989 , \25016 );
buf \U$19265 ( \25018 , \24580 );
not \U$19266 ( \25019 , \25018 );
buf \U$19267 ( \25020 , \24568 );
buf \U$19268 ( \25021 , \24569 );
buf \U$19269 ( \25022 , \24570 );
buf \U$19270 ( \25023 , \24573 );
buf \U$19271 ( \25024 , \24577 );
buf \U$19272 ( \25025 , \24580 );
buf \U$19273 ( \25026 , \24580 );
buf \U$19274 ( \25027 , \24580 );
buf \U$19275 ( \25028 , \24580 );
buf \U$19276 ( \25029 , \24580 );
buf \U$19277 ( \25030 , \24580 );
buf \U$19278 ( \25031 , \24580 );
buf \U$19279 ( \25032 , \24580 );
buf \U$19280 ( \25033 , \24580 );
buf \U$19281 ( \25034 , \24580 );
buf \U$19282 ( \25035 , \24580 );
buf \U$19283 ( \25036 , \24580 );
buf \U$19284 ( \25037 , \24580 );
buf \U$19285 ( \25038 , \24580 );
buf \U$19286 ( \25039 , \24580 );
buf \U$19287 ( \25040 , \24580 );
buf \U$19288 ( \25041 , \24580 );
buf \U$19289 ( \25042 , \24580 );
buf \U$19290 ( \25043 , \24580 );
buf \U$19291 ( \25044 , \24580 );
buf \U$19292 ( \25045 , \24580 );
buf \U$19293 ( \25046 , \24580 );
buf \U$19294 ( \25047 , \24580 );
buf \U$19295 ( \25048 , \24580 );
buf \U$19296 ( \25049 , \24580 );
buf \U$19297 ( \25050 , \24567 );
or \U$19298 ( \25051 , \25020 , \25021 , \25022 , \25023 , \25024 , \25025 , \25026 , \25027 , \25028 , \25029 , \25030 , \25031 , \25032 , \25033 , \25034 , \25035 , \25036 , \25037 , \25038 , \25039 , \25040 , \25041 , \25042 , \25043 , \25044 , \25045 , \25046 , \25047 , \25048 , \25049 , \25050 );
nand \U$19299 ( \25052 , \25019 , \25051 );
buf \U$19300 ( \25053 , \25052 );
buf \U$19301 ( \25054 , \24580 );
not \U$19302 ( \25055 , \25054 );
buf \U$19303 ( \25056 , \24577 );
buf \U$19304 ( \25057 , \24580 );
buf \U$19305 ( \25058 , \24580 );
buf \U$19306 ( \25059 , \24580 );
buf \U$19307 ( \25060 , \24580 );
buf \U$19308 ( \25061 , \24580 );
buf \U$19309 ( \25062 , \24580 );
buf \U$19310 ( \25063 , \24580 );
buf \U$19311 ( \25064 , \24580 );
buf \U$19312 ( \25065 , \24580 );
buf \U$19313 ( \25066 , \24580 );
buf \U$19314 ( \25067 , \24580 );
buf \U$19315 ( \25068 , \24580 );
buf \U$19316 ( \25069 , \24580 );
buf \U$19317 ( \25070 , \24580 );
buf \U$19318 ( \25071 , \24580 );
buf \U$19319 ( \25072 , \24580 );
buf \U$19320 ( \25073 , \24580 );
buf \U$19321 ( \25074 , \24580 );
buf \U$19322 ( \25075 , \24580 );
buf \U$19323 ( \25076 , \24580 );
buf \U$19324 ( \25077 , \24580 );
buf \U$19325 ( \25078 , \24580 );
buf \U$19326 ( \25079 , \24580 );
buf \U$19327 ( \25080 , \24580 );
buf \U$19328 ( \25081 , \24580 );
buf \U$19329 ( \25082 , \24573 );
buf \U$19330 ( \25083 , \24567 );
buf \U$19331 ( \25084 , \24568 );
buf \U$19332 ( \25085 , \24569 );
buf \U$19333 ( \25086 , \24570 );
or \U$19334 ( \25087 , \25083 , \25084 , \25085 , \25086 );
and \U$19335 ( \25088 , \25082 , \25087 );
or \U$19336 ( \25089 , \25056 , \25057 , \25058 , \25059 , \25060 , \25061 , \25062 , \25063 , \25064 , \25065 , \25066 , \25067 , \25068 , \25069 , \25070 , \25071 , \25072 , \25073 , \25074 , \25075 , \25076 , \25077 , \25078 , \25079 , \25080 , \25081 , \25088 );
and \U$19337 ( \25090 , \25055 , \25089 );
buf \U$19338 ( \25091 , \25090 );
or \U$19339 ( \25092 , \25053 , \25091 );
_DC g78fd ( \25093_nG78fd , \25017 , \25092 );
not \U$19340 ( \25094 , \25093_nG78fd );
buf \U$19341 ( \25095 , RIb7b9608_246);
buf \U$19342 ( \25096 , \24580 );
buf \U$19343 ( \25097 , \24580 );
buf \U$19344 ( \25098 , \24580 );
buf \U$19345 ( \25099 , \24580 );
buf \U$19346 ( \25100 , \24580 );
buf \U$19347 ( \25101 , \24580 );
buf \U$19348 ( \25102 , \24580 );
buf \U$19349 ( \25103 , \24580 );
buf \U$19350 ( \25104 , \24580 );
buf \U$19351 ( \25105 , \24580 );
buf \U$19352 ( \25106 , \24580 );
buf \U$19353 ( \25107 , \24580 );
buf \U$19354 ( \25108 , \24580 );
buf \U$19355 ( \25109 , \24580 );
buf \U$19356 ( \25110 , \24580 );
buf \U$19357 ( \25111 , \24580 );
buf \U$19358 ( \25112 , \24580 );
buf \U$19359 ( \25113 , \24580 );
buf \U$19360 ( \25114 , \24580 );
buf \U$19361 ( \25115 , \24580 );
buf \U$19362 ( \25116 , \24580 );
buf \U$19363 ( \25117 , \24580 );
buf \U$19364 ( \25118 , \24580 );
buf \U$19365 ( \25119 , \24580 );
buf \U$19366 ( \25120 , \24580 );
nor \U$19367 ( \25121 , \24567 , \24568 , \24569 , \24570 , \24574 , \24577 , \24580 , \25096 , \25097 , \25098 , \25099 , \25100 , \25101 , \25102 , \25103 , \25104 , \25105 , \25106 , \25107 , \25108 , \25109 , \25110 , \25111 , \25112 , \25113 , \25114 , \25115 , \25116 , \25117 , \25118 , \25119 , \25120 );
and \U$19368 ( \25122 , \7117 , \25121 );
buf \U$19369 ( \25123 , \24580 );
buf \U$19370 ( \25124 , \24580 );
buf \U$19371 ( \25125 , \24580 );
buf \U$19372 ( \25126 , \24580 );
buf \U$19373 ( \25127 , \24580 );
buf \U$19374 ( \25128 , \24580 );
buf \U$19375 ( \25129 , \24580 );
buf \U$19376 ( \25130 , \24580 );
buf \U$19377 ( \25131 , \24580 );
buf \U$19378 ( \25132 , \24580 );
buf \U$19379 ( \25133 , \24580 );
buf \U$19380 ( \25134 , \24580 );
buf \U$19381 ( \25135 , \24580 );
buf \U$19382 ( \25136 , \24580 );
buf \U$19383 ( \25137 , \24580 );
buf \U$19384 ( \25138 , \24580 );
buf \U$19385 ( \25139 , \24580 );
buf \U$19386 ( \25140 , \24580 );
buf \U$19387 ( \25141 , \24580 );
buf \U$19388 ( \25142 , \24580 );
buf \U$19389 ( \25143 , \24580 );
buf \U$19390 ( \25144 , \24580 );
buf \U$19391 ( \25145 , \24580 );
buf \U$19392 ( \25146 , \24580 );
buf \U$19393 ( \25147 , \24580 );
nor \U$19394 ( \25148 , \24608 , \24609 , \24610 , \24611 , \24573 , \24577 , \24580 , \25123 , \25124 , \25125 , \25126 , \25127 , \25128 , \25129 , \25130 , \25131 , \25132 , \25133 , \25134 , \25135 , \25136 , \25137 , \25138 , \25139 , \25140 , \25141 , \25142 , \25143 , \25144 , \25145 , \25146 , \25147 );
and \U$19395 ( \25149 , \7119 , \25148 );
buf \U$19396 ( \25150 , \24580 );
buf \U$19397 ( \25151 , \24580 );
buf \U$19398 ( \25152 , \24580 );
buf \U$19399 ( \25153 , \24580 );
buf \U$19400 ( \25154 , \24580 );
buf \U$19401 ( \25155 , \24580 );
buf \U$19402 ( \25156 , \24580 );
buf \U$19403 ( \25157 , \24580 );
buf \U$19404 ( \25158 , \24580 );
buf \U$19405 ( \25159 , \24580 );
buf \U$19406 ( \25160 , \24580 );
buf \U$19407 ( \25161 , \24580 );
buf \U$19408 ( \25162 , \24580 );
buf \U$19409 ( \25163 , \24580 );
buf \U$19410 ( \25164 , \24580 );
buf \U$19411 ( \25165 , \24580 );
buf \U$19412 ( \25166 , \24580 );
buf \U$19413 ( \25167 , \24580 );
buf \U$19414 ( \25168 , \24580 );
buf \U$19415 ( \25169 , \24580 );
buf \U$19416 ( \25170 , \24580 );
buf \U$19417 ( \25171 , \24580 );
buf \U$19418 ( \25172 , \24580 );
buf \U$19419 ( \25173 , \24580 );
buf \U$19420 ( \25174 , \24580 );
nor \U$19421 ( \25175 , \24567 , \24609 , \24610 , \24611 , \24573 , \24577 , \24580 , \25150 , \25151 , \25152 , \25153 , \25154 , \25155 , \25156 , \25157 , \25158 , \25159 , \25160 , \25161 , \25162 , \25163 , \25164 , \25165 , \25166 , \25167 , \25168 , \25169 , \25170 , \25171 , \25172 , \25173 , \25174 );
and \U$19422 ( \25176 , \7864 , \25175 );
buf \U$19423 ( \25177 , \24580 );
buf \U$19424 ( \25178 , \24580 );
buf \U$19425 ( \25179 , \24580 );
buf \U$19426 ( \25180 , \24580 );
buf \U$19427 ( \25181 , \24580 );
buf \U$19428 ( \25182 , \24580 );
buf \U$19429 ( \25183 , \24580 );
buf \U$19430 ( \25184 , \24580 );
buf \U$19431 ( \25185 , \24580 );
buf \U$19432 ( \25186 , \24580 );
buf \U$19433 ( \25187 , \24580 );
buf \U$19434 ( \25188 , \24580 );
buf \U$19435 ( \25189 , \24580 );
buf \U$19436 ( \25190 , \24580 );
buf \U$19437 ( \25191 , \24580 );
buf \U$19438 ( \25192 , \24580 );
buf \U$19439 ( \25193 , \24580 );
buf \U$19440 ( \25194 , \24580 );
buf \U$19441 ( \25195 , \24580 );
buf \U$19442 ( \25196 , \24580 );
buf \U$19443 ( \25197 , \24580 );
buf \U$19444 ( \25198 , \24580 );
buf \U$19445 ( \25199 , \24580 );
buf \U$19446 ( \25200 , \24580 );
buf \U$19447 ( \25201 , \24580 );
nor \U$19448 ( \25202 , \24608 , \24568 , \24610 , \24611 , \24573 , \24577 , \24580 , \25177 , \25178 , \25179 , \25180 , \25181 , \25182 , \25183 , \25184 , \25185 , \25186 , \25187 , \25188 , \25189 , \25190 , \25191 , \25192 , \25193 , \25194 , \25195 , \25196 , \25197 , \25198 , \25199 , \25200 , \25201 );
and \U$19449 ( \25203 , \7892 , \25202 );
buf \U$19450 ( \25204 , \24580 );
buf \U$19451 ( \25205 , \24580 );
buf \U$19452 ( \25206 , \24580 );
buf \U$19453 ( \25207 , \24580 );
buf \U$19454 ( \25208 , \24580 );
buf \U$19455 ( \25209 , \24580 );
buf \U$19456 ( \25210 , \24580 );
buf \U$19457 ( \25211 , \24580 );
buf \U$19458 ( \25212 , \24580 );
buf \U$19459 ( \25213 , \24580 );
buf \U$19460 ( \25214 , \24580 );
buf \U$19461 ( \25215 , \24580 );
buf \U$19462 ( \25216 , \24580 );
buf \U$19463 ( \25217 , \24580 );
buf \U$19464 ( \25218 , \24580 );
buf \U$19465 ( \25219 , \24580 );
buf \U$19466 ( \25220 , \24580 );
buf \U$19467 ( \25221 , \24580 );
buf \U$19468 ( \25222 , \24580 );
buf \U$19469 ( \25223 , \24580 );
buf \U$19470 ( \25224 , \24580 );
buf \U$19471 ( \25225 , \24580 );
buf \U$19472 ( \25226 , \24580 );
buf \U$19473 ( \25227 , \24580 );
buf \U$19474 ( \25228 , \24580 );
nor \U$19475 ( \25229 , \24567 , \24568 , \24610 , \24611 , \24573 , \24577 , \24580 , \25204 , \25205 , \25206 , \25207 , \25208 , \25209 , \25210 , \25211 , \25212 , \25213 , \25214 , \25215 , \25216 , \25217 , \25218 , \25219 , \25220 , \25221 , \25222 , \25223 , \25224 , \25225 , \25226 , \25227 , \25228 );
and \U$19476 ( \25230 , \7920 , \25229 );
buf \U$19477 ( \25231 , \24580 );
buf \U$19478 ( \25232 , \24580 );
buf \U$19479 ( \25233 , \24580 );
buf \U$19480 ( \25234 , \24580 );
buf \U$19481 ( \25235 , \24580 );
buf \U$19482 ( \25236 , \24580 );
buf \U$19483 ( \25237 , \24580 );
buf \U$19484 ( \25238 , \24580 );
buf \U$19485 ( \25239 , \24580 );
buf \U$19486 ( \25240 , \24580 );
buf \U$19487 ( \25241 , \24580 );
buf \U$19488 ( \25242 , \24580 );
buf \U$19489 ( \25243 , \24580 );
buf \U$19490 ( \25244 , \24580 );
buf \U$19491 ( \25245 , \24580 );
buf \U$19492 ( \25246 , \24580 );
buf \U$19493 ( \25247 , \24580 );
buf \U$19494 ( \25248 , \24580 );
buf \U$19495 ( \25249 , \24580 );
buf \U$19496 ( \25250 , \24580 );
buf \U$19497 ( \25251 , \24580 );
buf \U$19498 ( \25252 , \24580 );
buf \U$19499 ( \25253 , \24580 );
buf \U$19500 ( \25254 , \24580 );
buf \U$19501 ( \25255 , \24580 );
nor \U$19502 ( \25256 , \24608 , \24609 , \24569 , \24611 , \24573 , \24577 , \24580 , \25231 , \25232 , \25233 , \25234 , \25235 , \25236 , \25237 , \25238 , \25239 , \25240 , \25241 , \25242 , \25243 , \25244 , \25245 , \25246 , \25247 , \25248 , \25249 , \25250 , \25251 , \25252 , \25253 , \25254 , \25255 );
and \U$19503 ( \25257 , \7948 , \25256 );
buf \U$19504 ( \25258 , \24580 );
buf \U$19505 ( \25259 , \24580 );
buf \U$19506 ( \25260 , \24580 );
buf \U$19507 ( \25261 , \24580 );
buf \U$19508 ( \25262 , \24580 );
buf \U$19509 ( \25263 , \24580 );
buf \U$19510 ( \25264 , \24580 );
buf \U$19511 ( \25265 , \24580 );
buf \U$19512 ( \25266 , \24580 );
buf \U$19513 ( \25267 , \24580 );
buf \U$19514 ( \25268 , \24580 );
buf \U$19515 ( \25269 , \24580 );
buf \U$19516 ( \25270 , \24580 );
buf \U$19517 ( \25271 , \24580 );
buf \U$19518 ( \25272 , \24580 );
buf \U$19519 ( \25273 , \24580 );
buf \U$19520 ( \25274 , \24580 );
buf \U$19521 ( \25275 , \24580 );
buf \U$19522 ( \25276 , \24580 );
buf \U$19523 ( \25277 , \24580 );
buf \U$19524 ( \25278 , \24580 );
buf \U$19525 ( \25279 , \24580 );
buf \U$19526 ( \25280 , \24580 );
buf \U$19527 ( \25281 , \24580 );
buf \U$19528 ( \25282 , \24580 );
nor \U$19529 ( \25283 , \24567 , \24609 , \24569 , \24611 , \24573 , \24577 , \24580 , \25258 , \25259 , \25260 , \25261 , \25262 , \25263 , \25264 , \25265 , \25266 , \25267 , \25268 , \25269 , \25270 , \25271 , \25272 , \25273 , \25274 , \25275 , \25276 , \25277 , \25278 , \25279 , \25280 , \25281 , \25282 );
and \U$19530 ( \25284 , \7976 , \25283 );
buf \U$19531 ( \25285 , \24580 );
buf \U$19532 ( \25286 , \24580 );
buf \U$19533 ( \25287 , \24580 );
buf \U$19534 ( \25288 , \24580 );
buf \U$19535 ( \25289 , \24580 );
buf \U$19536 ( \25290 , \24580 );
buf \U$19537 ( \25291 , \24580 );
buf \U$19538 ( \25292 , \24580 );
buf \U$19539 ( \25293 , \24580 );
buf \U$19540 ( \25294 , \24580 );
buf \U$19541 ( \25295 , \24580 );
buf \U$19542 ( \25296 , \24580 );
buf \U$19543 ( \25297 , \24580 );
buf \U$19544 ( \25298 , \24580 );
buf \U$19545 ( \25299 , \24580 );
buf \U$19546 ( \25300 , \24580 );
buf \U$19547 ( \25301 , \24580 );
buf \U$19548 ( \25302 , \24580 );
buf \U$19549 ( \25303 , \24580 );
buf \U$19550 ( \25304 , \24580 );
buf \U$19551 ( \25305 , \24580 );
buf \U$19552 ( \25306 , \24580 );
buf \U$19553 ( \25307 , \24580 );
buf \U$19554 ( \25308 , \24580 );
buf \U$19555 ( \25309 , \24580 );
nor \U$19556 ( \25310 , \24608 , \24568 , \24569 , \24611 , \24573 , \24577 , \24580 , \25285 , \25286 , \25287 , \25288 , \25289 , \25290 , \25291 , \25292 , \25293 , \25294 , \25295 , \25296 , \25297 , \25298 , \25299 , \25300 , \25301 , \25302 , \25303 , \25304 , \25305 , \25306 , \25307 , \25308 , \25309 );
and \U$19557 ( \25311 , \8004 , \25310 );
buf \U$19558 ( \25312 , \24580 );
buf \U$19559 ( \25313 , \24580 );
buf \U$19560 ( \25314 , \24580 );
buf \U$19561 ( \25315 , \24580 );
buf \U$19562 ( \25316 , \24580 );
buf \U$19563 ( \25317 , \24580 );
buf \U$19564 ( \25318 , \24580 );
buf \U$19565 ( \25319 , \24580 );
buf \U$19566 ( \25320 , \24580 );
buf \U$19567 ( \25321 , \24580 );
buf \U$19568 ( \25322 , \24580 );
buf \U$19569 ( \25323 , \24580 );
buf \U$19570 ( \25324 , \24580 );
buf \U$19571 ( \25325 , \24580 );
buf \U$19572 ( \25326 , \24580 );
buf \U$19573 ( \25327 , \24580 );
buf \U$19574 ( \25328 , \24580 );
buf \U$19575 ( \25329 , \24580 );
buf \U$19576 ( \25330 , \24580 );
buf \U$19577 ( \25331 , \24580 );
buf \U$19578 ( \25332 , \24580 );
buf \U$19579 ( \25333 , \24580 );
buf \U$19580 ( \25334 , \24580 );
buf \U$19581 ( \25335 , \24580 );
buf \U$19582 ( \25336 , \24580 );
nor \U$19583 ( \25337 , \24567 , \24568 , \24569 , \24611 , \24573 , \24577 , \24580 , \25312 , \25313 , \25314 , \25315 , \25316 , \25317 , \25318 , \25319 , \25320 , \25321 , \25322 , \25323 , \25324 , \25325 , \25326 , \25327 , \25328 , \25329 , \25330 , \25331 , \25332 , \25333 , \25334 , \25335 , \25336 );
and \U$19584 ( \25338 , \8032 , \25337 );
buf \U$19585 ( \25339 , \24580 );
buf \U$19586 ( \25340 , \24580 );
buf \U$19587 ( \25341 , \24580 );
buf \U$19588 ( \25342 , \24580 );
buf \U$19589 ( \25343 , \24580 );
buf \U$19590 ( \25344 , \24580 );
buf \U$19591 ( \25345 , \24580 );
buf \U$19592 ( \25346 , \24580 );
buf \U$19593 ( \25347 , \24580 );
buf \U$19594 ( \25348 , \24580 );
buf \U$19595 ( \25349 , \24580 );
buf \U$19596 ( \25350 , \24580 );
buf \U$19597 ( \25351 , \24580 );
buf \U$19598 ( \25352 , \24580 );
buf \U$19599 ( \25353 , \24580 );
buf \U$19600 ( \25354 , \24580 );
buf \U$19601 ( \25355 , \24580 );
buf \U$19602 ( \25356 , \24580 );
buf \U$19603 ( \25357 , \24580 );
buf \U$19604 ( \25358 , \24580 );
buf \U$19605 ( \25359 , \24580 );
buf \U$19606 ( \25360 , \24580 );
buf \U$19607 ( \25361 , \24580 );
buf \U$19608 ( \25362 , \24580 );
buf \U$19609 ( \25363 , \24580 );
nor \U$19610 ( \25364 , \24608 , \24609 , \24610 , \24570 , \24573 , \24577 , \24580 , \25339 , \25340 , \25341 , \25342 , \25343 , \25344 , \25345 , \25346 , \25347 , \25348 , \25349 , \25350 , \25351 , \25352 , \25353 , \25354 , \25355 , \25356 , \25357 , \25358 , \25359 , \25360 , \25361 , \25362 , \25363 );
and \U$19611 ( \25365 , \8060 , \25364 );
buf \U$19612 ( \25366 , \24580 );
buf \U$19613 ( \25367 , \24580 );
buf \U$19614 ( \25368 , \24580 );
buf \U$19615 ( \25369 , \24580 );
buf \U$19616 ( \25370 , \24580 );
buf \U$19617 ( \25371 , \24580 );
buf \U$19618 ( \25372 , \24580 );
buf \U$19619 ( \25373 , \24580 );
buf \U$19620 ( \25374 , \24580 );
buf \U$19621 ( \25375 , \24580 );
buf \U$19622 ( \25376 , \24580 );
buf \U$19623 ( \25377 , \24580 );
buf \U$19624 ( \25378 , \24580 );
buf \U$19625 ( \25379 , \24580 );
buf \U$19626 ( \25380 , \24580 );
buf \U$19627 ( \25381 , \24580 );
buf \U$19628 ( \25382 , \24580 );
buf \U$19629 ( \25383 , \24580 );
buf \U$19630 ( \25384 , \24580 );
buf \U$19631 ( \25385 , \24580 );
buf \U$19632 ( \25386 , \24580 );
buf \U$19633 ( \25387 , \24580 );
buf \U$19634 ( \25388 , \24580 );
buf \U$19635 ( \25389 , \24580 );
buf \U$19636 ( \25390 , \24580 );
nor \U$19637 ( \25391 , \24567 , \24609 , \24610 , \24570 , \24573 , \24577 , \24580 , \25366 , \25367 , \25368 , \25369 , \25370 , \25371 , \25372 , \25373 , \25374 , \25375 , \25376 , \25377 , \25378 , \25379 , \25380 , \25381 , \25382 , \25383 , \25384 , \25385 , \25386 , \25387 , \25388 , \25389 , \25390 );
and \U$19638 ( \25392 , \8088 , \25391 );
buf \U$19639 ( \25393 , \24580 );
buf \U$19640 ( \25394 , \24580 );
buf \U$19641 ( \25395 , \24580 );
buf \U$19642 ( \25396 , \24580 );
buf \U$19643 ( \25397 , \24580 );
buf \U$19644 ( \25398 , \24580 );
buf \U$19645 ( \25399 , \24580 );
buf \U$19646 ( \25400 , \24580 );
buf \U$19647 ( \25401 , \24580 );
buf \U$19648 ( \25402 , \24580 );
buf \U$19649 ( \25403 , \24580 );
buf \U$19650 ( \25404 , \24580 );
buf \U$19651 ( \25405 , \24580 );
buf \U$19652 ( \25406 , \24580 );
buf \U$19653 ( \25407 , \24580 );
buf \U$19654 ( \25408 , \24580 );
buf \U$19655 ( \25409 , \24580 );
buf \U$19656 ( \25410 , \24580 );
buf \U$19657 ( \25411 , \24580 );
buf \U$19658 ( \25412 , \24580 );
buf \U$19659 ( \25413 , \24580 );
buf \U$19660 ( \25414 , \24580 );
buf \U$19661 ( \25415 , \24580 );
buf \U$19662 ( \25416 , \24580 );
buf \U$19663 ( \25417 , \24580 );
nor \U$19664 ( \25418 , \24608 , \24568 , \24610 , \24570 , \24573 , \24577 , \24580 , \25393 , \25394 , \25395 , \25396 , \25397 , \25398 , \25399 , \25400 , \25401 , \25402 , \25403 , \25404 , \25405 , \25406 , \25407 , \25408 , \25409 , \25410 , \25411 , \25412 , \25413 , \25414 , \25415 , \25416 , \25417 );
and \U$19665 ( \25419 , \8116 , \25418 );
buf \U$19666 ( \25420 , \24580 );
buf \U$19667 ( \25421 , \24580 );
buf \U$19668 ( \25422 , \24580 );
buf \U$19669 ( \25423 , \24580 );
buf \U$19670 ( \25424 , \24580 );
buf \U$19671 ( \25425 , \24580 );
buf \U$19672 ( \25426 , \24580 );
buf \U$19673 ( \25427 , \24580 );
buf \U$19674 ( \25428 , \24580 );
buf \U$19675 ( \25429 , \24580 );
buf \U$19676 ( \25430 , \24580 );
buf \U$19677 ( \25431 , \24580 );
buf \U$19678 ( \25432 , \24580 );
buf \U$19679 ( \25433 , \24580 );
buf \U$19680 ( \25434 , \24580 );
buf \U$19681 ( \25435 , \24580 );
buf \U$19682 ( \25436 , \24580 );
buf \U$19683 ( \25437 , \24580 );
buf \U$19684 ( \25438 , \24580 );
buf \U$19685 ( \25439 , \24580 );
buf \U$19686 ( \25440 , \24580 );
buf \U$19687 ( \25441 , \24580 );
buf \U$19688 ( \25442 , \24580 );
buf \U$19689 ( \25443 , \24580 );
buf \U$19690 ( \25444 , \24580 );
nor \U$19691 ( \25445 , \24567 , \24568 , \24610 , \24570 , \24573 , \24577 , \24580 , \25420 , \25421 , \25422 , \25423 , \25424 , \25425 , \25426 , \25427 , \25428 , \25429 , \25430 , \25431 , \25432 , \25433 , \25434 , \25435 , \25436 , \25437 , \25438 , \25439 , \25440 , \25441 , \25442 , \25443 , \25444 );
and \U$19692 ( \25446 , \8144 , \25445 );
buf \U$19693 ( \25447 , \24580 );
buf \U$19694 ( \25448 , \24580 );
buf \U$19695 ( \25449 , \24580 );
buf \U$19696 ( \25450 , \24580 );
buf \U$19697 ( \25451 , \24580 );
buf \U$19698 ( \25452 , \24580 );
buf \U$19699 ( \25453 , \24580 );
buf \U$19700 ( \25454 , \24580 );
buf \U$19701 ( \25455 , \24580 );
buf \U$19702 ( \25456 , \24580 );
buf \U$19703 ( \25457 , \24580 );
buf \U$19704 ( \25458 , \24580 );
buf \U$19705 ( \25459 , \24580 );
buf \U$19706 ( \25460 , \24580 );
buf \U$19707 ( \25461 , \24580 );
buf \U$19708 ( \25462 , \24580 );
buf \U$19709 ( \25463 , \24580 );
buf \U$19710 ( \25464 , \24580 );
buf \U$19711 ( \25465 , \24580 );
buf \U$19712 ( \25466 , \24580 );
buf \U$19713 ( \25467 , \24580 );
buf \U$19714 ( \25468 , \24580 );
buf \U$19715 ( \25469 , \24580 );
buf \U$19716 ( \25470 , \24580 );
buf \U$19717 ( \25471 , \24580 );
nor \U$19718 ( \25472 , \24608 , \24609 , \24569 , \24570 , \24573 , \24577 , \24580 , \25447 , \25448 , \25449 , \25450 , \25451 , \25452 , \25453 , \25454 , \25455 , \25456 , \25457 , \25458 , \25459 , \25460 , \25461 , \25462 , \25463 , \25464 , \25465 , \25466 , \25467 , \25468 , \25469 , \25470 , \25471 );
and \U$19719 ( \25473 , \8172 , \25472 );
buf \U$19720 ( \25474 , \24580 );
buf \U$19721 ( \25475 , \24580 );
buf \U$19722 ( \25476 , \24580 );
buf \U$19723 ( \25477 , \24580 );
buf \U$19724 ( \25478 , \24580 );
buf \U$19725 ( \25479 , \24580 );
buf \U$19726 ( \25480 , \24580 );
buf \U$19727 ( \25481 , \24580 );
buf \U$19728 ( \25482 , \24580 );
buf \U$19729 ( \25483 , \24580 );
buf \U$19730 ( \25484 , \24580 );
buf \U$19731 ( \25485 , \24580 );
buf \U$19732 ( \25486 , \24580 );
buf \U$19733 ( \25487 , \24580 );
buf \U$19734 ( \25488 , \24580 );
buf \U$19735 ( \25489 , \24580 );
buf \U$19736 ( \25490 , \24580 );
buf \U$19737 ( \25491 , \24580 );
buf \U$19738 ( \25492 , \24580 );
buf \U$19739 ( \25493 , \24580 );
buf \U$19740 ( \25494 , \24580 );
buf \U$19741 ( \25495 , \24580 );
buf \U$19742 ( \25496 , \24580 );
buf \U$19743 ( \25497 , \24580 );
buf \U$19744 ( \25498 , \24580 );
nor \U$19745 ( \25499 , \24567 , \24609 , \24569 , \24570 , \24573 , \24577 , \24580 , \25474 , \25475 , \25476 , \25477 , \25478 , \25479 , \25480 , \25481 , \25482 , \25483 , \25484 , \25485 , \25486 , \25487 , \25488 , \25489 , \25490 , \25491 , \25492 , \25493 , \25494 , \25495 , \25496 , \25497 , \25498 );
and \U$19746 ( \25500 , \8200 , \25499 );
buf \U$19747 ( \25501 , \24580 );
buf \U$19748 ( \25502 , \24580 );
buf \U$19749 ( \25503 , \24580 );
buf \U$19750 ( \25504 , \24580 );
buf \U$19751 ( \25505 , \24580 );
buf \U$19752 ( \25506 , \24580 );
buf \U$19753 ( \25507 , \24580 );
buf \U$19754 ( \25508 , \24580 );
buf \U$19755 ( \25509 , \24580 );
buf \U$19756 ( \25510 , \24580 );
buf \U$19757 ( \25511 , \24580 );
buf \U$19758 ( \25512 , \24580 );
buf \U$19759 ( \25513 , \24580 );
buf \U$19760 ( \25514 , \24580 );
buf \U$19761 ( \25515 , \24580 );
buf \U$19762 ( \25516 , \24580 );
buf \U$19763 ( \25517 , \24580 );
buf \U$19764 ( \25518 , \24580 );
buf \U$19765 ( \25519 , \24580 );
buf \U$19766 ( \25520 , \24580 );
buf \U$19767 ( \25521 , \24580 );
buf \U$19768 ( \25522 , \24580 );
buf \U$19769 ( \25523 , \24580 );
buf \U$19770 ( \25524 , \24580 );
buf \U$19771 ( \25525 , \24580 );
nor \U$19772 ( \25526 , \24608 , \24568 , \24569 , \24570 , \24573 , \24577 , \24580 , \25501 , \25502 , \25503 , \25504 , \25505 , \25506 , \25507 , \25508 , \25509 , \25510 , \25511 , \25512 , \25513 , \25514 , \25515 , \25516 , \25517 , \25518 , \25519 , \25520 , \25521 , \25522 , \25523 , \25524 , \25525 );
and \U$19773 ( \25527 , \8228 , \25526 );
or \U$19774 ( \25528 , \25122 , \25149 , \25176 , \25203 , \25230 , \25257 , \25284 , \25311 , \25338 , \25365 , \25392 , \25419 , \25446 , \25473 , \25500 , \25527 );
buf \U$19775 ( \25529 , \24580 );
not \U$19776 ( \25530 , \25529 );
buf \U$19777 ( \25531 , \24568 );
buf \U$19778 ( \25532 , \24569 );
buf \U$19779 ( \25533 , \24570 );
buf \U$19780 ( \25534 , \24573 );
buf \U$19781 ( \25535 , \24577 );
buf \U$19782 ( \25536 , \24580 );
buf \U$19783 ( \25537 , \24580 );
buf \U$19784 ( \25538 , \24580 );
buf \U$19785 ( \25539 , \24580 );
buf \U$19786 ( \25540 , \24580 );
buf \U$19787 ( \25541 , \24580 );
buf \U$19788 ( \25542 , \24580 );
buf \U$19789 ( \25543 , \24580 );
buf \U$19790 ( \25544 , \24580 );
buf \U$19791 ( \25545 , \24580 );
buf \U$19792 ( \25546 , \24580 );
buf \U$19793 ( \25547 , \24580 );
buf \U$19794 ( \25548 , \24580 );
buf \U$19795 ( \25549 , \24580 );
buf \U$19796 ( \25550 , \24580 );
buf \U$19797 ( \25551 , \24580 );
buf \U$19798 ( \25552 , \24580 );
buf \U$19799 ( \25553 , \24580 );
buf \U$19800 ( \25554 , \24580 );
buf \U$19801 ( \25555 , \24580 );
buf \U$19802 ( \25556 , \24580 );
buf \U$19803 ( \25557 , \24580 );
buf \U$19804 ( \25558 , \24580 );
buf \U$19805 ( \25559 , \24580 );
buf \U$19806 ( \25560 , \24580 );
buf \U$19807 ( \25561 , \24567 );
or \U$19808 ( \25562 , \25531 , \25532 , \25533 , \25534 , \25535 , \25536 , \25537 , \25538 , \25539 , \25540 , \25541 , \25542 , \25543 , \25544 , \25545 , \25546 , \25547 , \25548 , \25549 , \25550 , \25551 , \25552 , \25553 , \25554 , \25555 , \25556 , \25557 , \25558 , \25559 , \25560 , \25561 );
nand \U$19809 ( \25563 , \25530 , \25562 );
buf \U$19810 ( \25564 , \25563 );
buf \U$19811 ( \25565 , \24580 );
not \U$19812 ( \25566 , \25565 );
buf \U$19813 ( \25567 , \24577 );
buf \U$19814 ( \25568 , \24580 );
buf \U$19815 ( \25569 , \24580 );
buf \U$19816 ( \25570 , \24580 );
buf \U$19817 ( \25571 , \24580 );
buf \U$19818 ( \25572 , \24580 );
buf \U$19819 ( \25573 , \24580 );
buf \U$19820 ( \25574 , \24580 );
buf \U$19821 ( \25575 , \24580 );
buf \U$19822 ( \25576 , \24580 );
buf \U$19823 ( \25577 , \24580 );
buf \U$19824 ( \25578 , \24580 );
buf \U$19825 ( \25579 , \24580 );
buf \U$19826 ( \25580 , \24580 );
buf \U$19827 ( \25581 , \24580 );
buf \U$19828 ( \25582 , \24580 );
buf \U$19829 ( \25583 , \24580 );
buf \U$19830 ( \25584 , \24580 );
buf \U$19831 ( \25585 , \24580 );
buf \U$19832 ( \25586 , \24580 );
buf \U$19833 ( \25587 , \24580 );
buf \U$19834 ( \25588 , \24580 );
buf \U$19835 ( \25589 , \24580 );
buf \U$19836 ( \25590 , \24580 );
buf \U$19837 ( \25591 , \24580 );
buf \U$19838 ( \25592 , \24580 );
buf \U$19839 ( \25593 , \24573 );
buf \U$19840 ( \25594 , \24567 );
buf \U$19841 ( \25595 , \24568 );
buf \U$19842 ( \25596 , \24569 );
buf \U$19843 ( \25597 , \24570 );
or \U$19844 ( \25598 , \25594 , \25595 , \25596 , \25597 );
and \U$19845 ( \25599 , \25593 , \25598 );
or \U$19846 ( \25600 , \25567 , \25568 , \25569 , \25570 , \25571 , \25572 , \25573 , \25574 , \25575 , \25576 , \25577 , \25578 , \25579 , \25580 , \25581 , \25582 , \25583 , \25584 , \25585 , \25586 , \25587 , \25588 , \25589 , \25590 , \25591 , \25592 , \25599 );
and \U$19847 ( \25601 , \25566 , \25600 );
buf \U$19848 ( \25602 , \25601 );
or \U$19849 ( \25603 , \25564 , \25602 );
_DC g7afc ( \25604_nG7afc , \25528 , \25603 );
buf \U$19850 ( \25605 , \25604_nG7afc );
xor \U$19851 ( \25606 , \25095 , \25605 );
buf \U$19852 ( \25607 , RIb7b9590_247);
and \U$19853 ( \25608 , \7126 , \25121 );
and \U$19854 ( \25609 , \7128 , \25148 );
and \U$19855 ( \25610 , \8338 , \25175 );
and \U$19856 ( \25611 , \8340 , \25202 );
and \U$19857 ( \25612 , \8342 , \25229 );
and \U$19858 ( \25613 , \8344 , \25256 );
and \U$19859 ( \25614 , \8346 , \25283 );
and \U$19860 ( \25615 , \8348 , \25310 );
and \U$19861 ( \25616 , \8350 , \25337 );
and \U$19862 ( \25617 , \8352 , \25364 );
and \U$19863 ( \25618 , \8354 , \25391 );
and \U$19864 ( \25619 , \8356 , \25418 );
and \U$19865 ( \25620 , \8358 , \25445 );
and \U$19866 ( \25621 , \8360 , \25472 );
and \U$19867 ( \25622 , \8362 , \25499 );
and \U$19868 ( \25623 , \8364 , \25526 );
or \U$19869 ( \25624 , \25608 , \25609 , \25610 , \25611 , \25612 , \25613 , \25614 , \25615 , \25616 , \25617 , \25618 , \25619 , \25620 , \25621 , \25622 , \25623 );
_DC g7b11 ( \25625_nG7b11 , \25624 , \25603 );
buf \U$19870 ( \25626 , \25625_nG7b11 );
xor \U$19871 ( \25627 , \25607 , \25626 );
or \U$19872 ( \25628 , \25606 , \25627 );
buf \U$19873 ( \25629 , RIb7b9518_248);
and \U$19874 ( \25630 , \7136 , \25121 );
and \U$19875 ( \25631 , \7138 , \25148 );
and \U$19876 ( \25632 , \8374 , \25175 );
and \U$19877 ( \25633 , \8376 , \25202 );
and \U$19878 ( \25634 , \8378 , \25229 );
and \U$19879 ( \25635 , \8380 , \25256 );
and \U$19880 ( \25636 , \8382 , \25283 );
and \U$19881 ( \25637 , \8384 , \25310 );
and \U$19882 ( \25638 , \8386 , \25337 );
and \U$19883 ( \25639 , \8388 , \25364 );
and \U$19884 ( \25640 , \8390 , \25391 );
and \U$19885 ( \25641 , \8392 , \25418 );
and \U$19886 ( \25642 , \8394 , \25445 );
and \U$19887 ( \25643 , \8396 , \25472 );
and \U$19888 ( \25644 , \8398 , \25499 );
and \U$19889 ( \25645 , \8400 , \25526 );
or \U$19890 ( \25646 , \25630 , \25631 , \25632 , \25633 , \25634 , \25635 , \25636 , \25637 , \25638 , \25639 , \25640 , \25641 , \25642 , \25643 , \25644 , \25645 );
_DC g7b27 ( \25647_nG7b27 , \25646 , \25603 );
buf \U$19891 ( \25648 , \25647_nG7b27 );
xor \U$19892 ( \25649 , \25629 , \25648 );
or \U$19893 ( \25650 , \25628 , \25649 );
buf \U$19894 ( \25651 , RIb7b94a0_249);
and \U$19895 ( \25652 , \7146 , \25121 );
and \U$19896 ( \25653 , \7148 , \25148 );
and \U$19897 ( \25654 , \8410 , \25175 );
and \U$19898 ( \25655 , \8412 , \25202 );
and \U$19899 ( \25656 , \8414 , \25229 );
and \U$19900 ( \25657 , \8416 , \25256 );
and \U$19901 ( \25658 , \8418 , \25283 );
and \U$19902 ( \25659 , \8420 , \25310 );
and \U$19903 ( \25660 , \8422 , \25337 );
and \U$19904 ( \25661 , \8424 , \25364 );
and \U$19905 ( \25662 , \8426 , \25391 );
and \U$19906 ( \25663 , \8428 , \25418 );
and \U$19907 ( \25664 , \8430 , \25445 );
and \U$19908 ( \25665 , \8432 , \25472 );
and \U$19909 ( \25666 , \8434 , \25499 );
and \U$19910 ( \25667 , \8436 , \25526 );
or \U$19911 ( \25668 , \25652 , \25653 , \25654 , \25655 , \25656 , \25657 , \25658 , \25659 , \25660 , \25661 , \25662 , \25663 , \25664 , \25665 , \25666 , \25667 );
_DC g7b3d ( \25669_nG7b3d , \25668 , \25603 );
buf \U$19912 ( \25670 , \25669_nG7b3d );
xor \U$19913 ( \25671 , \25651 , \25670 );
or \U$19914 ( \25672 , \25650 , \25671 );
buf \U$19915 ( \25673 , RIb7b9428_250);
and \U$19916 ( \25674 , \7156 , \25121 );
and \U$19917 ( \25675 , \7158 , \25148 );
and \U$19918 ( \25676 , \8446 , \25175 );
and \U$19919 ( \25677 , \8448 , \25202 );
and \U$19920 ( \25678 , \8450 , \25229 );
and \U$19921 ( \25679 , \8452 , \25256 );
and \U$19922 ( \25680 , \8454 , \25283 );
and \U$19923 ( \25681 , \8456 , \25310 );
and \U$19924 ( \25682 , \8458 , \25337 );
and \U$19925 ( \25683 , \8460 , \25364 );
and \U$19926 ( \25684 , \8462 , \25391 );
and \U$19927 ( \25685 , \8464 , \25418 );
and \U$19928 ( \25686 , \8466 , \25445 );
and \U$19929 ( \25687 , \8468 , \25472 );
and \U$19930 ( \25688 , \8470 , \25499 );
and \U$19931 ( \25689 , \8472 , \25526 );
or \U$19932 ( \25690 , \25674 , \25675 , \25676 , \25677 , \25678 , \25679 , \25680 , \25681 , \25682 , \25683 , \25684 , \25685 , \25686 , \25687 , \25688 , \25689 );
_DC g7b53 ( \25691_nG7b53 , \25690 , \25603 );
buf \U$19933 ( \25692 , \25691_nG7b53 );
xor \U$19934 ( \25693 , \25673 , \25692 );
or \U$19935 ( \25694 , \25672 , \25693 );
buf \U$19936 ( \25695 , RIb7b93b0_251);
and \U$19937 ( \25696 , \7166 , \25121 );
and \U$19938 ( \25697 , \7168 , \25148 );
and \U$19939 ( \25698 , \8482 , \25175 );
and \U$19940 ( \25699 , \8484 , \25202 );
and \U$19941 ( \25700 , \8486 , \25229 );
and \U$19942 ( \25701 , \8488 , \25256 );
and \U$19943 ( \25702 , \8490 , \25283 );
and \U$19944 ( \25703 , \8492 , \25310 );
and \U$19945 ( \25704 , \8494 , \25337 );
and \U$19946 ( \25705 , \8496 , \25364 );
and \U$19947 ( \25706 , \8498 , \25391 );
and \U$19948 ( \25707 , \8500 , \25418 );
and \U$19949 ( \25708 , \8502 , \25445 );
and \U$19950 ( \25709 , \8504 , \25472 );
and \U$19951 ( \25710 , \8506 , \25499 );
and \U$19952 ( \25711 , \8508 , \25526 );
or \U$19953 ( \25712 , \25696 , \25697 , \25698 , \25699 , \25700 , \25701 , \25702 , \25703 , \25704 , \25705 , \25706 , \25707 , \25708 , \25709 , \25710 , \25711 );
_DC g7b69 ( \25713_nG7b69 , \25712 , \25603 );
buf \U$19954 ( \25714 , \25713_nG7b69 );
xor \U$19955 ( \25715 , \25695 , \25714 );
or \U$19956 ( \25716 , \25694 , \25715 );
buf \U$19957 ( \25717 , RIb7af720_252);
and \U$19958 ( \25718 , \7176 , \25121 );
and \U$19959 ( \25719 , \7178 , \25148 );
and \U$19960 ( \25720 , \8518 , \25175 );
and \U$19961 ( \25721 , \8520 , \25202 );
and \U$19962 ( \25722 , \8522 , \25229 );
and \U$19963 ( \25723 , \8524 , \25256 );
and \U$19964 ( \25724 , \8526 , \25283 );
and \U$19965 ( \25725 , \8528 , \25310 );
and \U$19966 ( \25726 , \8530 , \25337 );
and \U$19967 ( \25727 , \8532 , \25364 );
and \U$19968 ( \25728 , \8534 , \25391 );
and \U$19969 ( \25729 , \8536 , \25418 );
and \U$19970 ( \25730 , \8538 , \25445 );
and \U$19971 ( \25731 , \8540 , \25472 );
and \U$19972 ( \25732 , \8542 , \25499 );
and \U$19973 ( \25733 , \8544 , \25526 );
or \U$19974 ( \25734 , \25718 , \25719 , \25720 , \25721 , \25722 , \25723 , \25724 , \25725 , \25726 , \25727 , \25728 , \25729 , \25730 , \25731 , \25732 , \25733 );
_DC g7b7f ( \25735_nG7b7f , \25734 , \25603 );
buf \U$19975 ( \25736 , \25735_nG7b7f );
xor \U$19976 ( \25737 , \25717 , \25736 );
or \U$19977 ( \25738 , \25716 , \25737 );
buf \U$19978 ( \25739 , RIb7af6a8_253);
and \U$19979 ( \25740 , \7186 , \25121 );
and \U$19980 ( \25741 , \7188 , \25148 );
and \U$19981 ( \25742 , \8554 , \25175 );
and \U$19982 ( \25743 , \8556 , \25202 );
and \U$19983 ( \25744 , \8558 , \25229 );
and \U$19984 ( \25745 , \8560 , \25256 );
and \U$19985 ( \25746 , \8562 , \25283 );
and \U$19986 ( \25747 , \8564 , \25310 );
and \U$19987 ( \25748 , \8566 , \25337 );
and \U$19988 ( \25749 , \8568 , \25364 );
and \U$19989 ( \25750 , \8570 , \25391 );
and \U$19990 ( \25751 , \8572 , \25418 );
and \U$19991 ( \25752 , \8574 , \25445 );
and \U$19992 ( \25753 , \8576 , \25472 );
and \U$19993 ( \25754 , \8578 , \25499 );
and \U$19994 ( \25755 , \8580 , \25526 );
or \U$19995 ( \25756 , \25740 , \25741 , \25742 , \25743 , \25744 , \25745 , \25746 , \25747 , \25748 , \25749 , \25750 , \25751 , \25752 , \25753 , \25754 , \25755 );
_DC g7b95 ( \25757_nG7b95 , \25756 , \25603 );
buf \U$19996 ( \25758 , \25757_nG7b95 );
xor \U$19997 ( \25759 , \25739 , \25758 );
or \U$19998 ( \25760 , \25738 , \25759 );
not \U$19999 ( \25761 , \25760 );
buf \U$20000 ( \25762 , \25761 );
and \U$20001 ( \25763 , \25094 , \25762 );
buf \U$20002 ( \25764 , RIb7af630_254);
buf \U$20003 ( \25765 , \24580 );
buf \U$20004 ( \25766 , \24580 );
buf \U$20005 ( \25767 , \24580 );
buf \U$20006 ( \25768 , \24580 );
buf \U$20007 ( \25769 , \24580 );
buf \U$20008 ( \25770 , \24580 );
buf \U$20009 ( \25771 , \24580 );
buf \U$20010 ( \25772 , \24580 );
buf \U$20011 ( \25773 , \24580 );
buf \U$20012 ( \25774 , \24580 );
buf \U$20013 ( \25775 , \24580 );
buf \U$20014 ( \25776 , \24580 );
buf \U$20015 ( \25777 , \24580 );
buf \U$20016 ( \25778 , \24580 );
buf \U$20017 ( \25779 , \24580 );
buf \U$20018 ( \25780 , \24580 );
buf \U$20019 ( \25781 , \24580 );
buf \U$20020 ( \25782 , \24580 );
buf \U$20021 ( \25783 , \24580 );
buf \U$20022 ( \25784 , \24580 );
buf \U$20023 ( \25785 , \24580 );
buf \U$20024 ( \25786 , \24580 );
buf \U$20025 ( \25787 , \24580 );
buf \U$20026 ( \25788 , \24580 );
buf \U$20027 ( \25789 , \24580 );
nor \U$20028 ( \25790 , \24567 , \24568 , \24569 , \24570 , \24574 , \24577 , \24580 , \25765 , \25766 , \25767 , \25768 , \25769 , \25770 , \25771 , \25772 , \25773 , \25774 , \25775 , \25776 , \25777 , \25778 , \25779 , \25780 , \25781 , \25782 , \25783 , \25784 , \25785 , \25786 , \25787 , \25788 , \25789 );
and \U$20029 ( \25791 , \7198 , \25790 );
buf \U$20030 ( \25792 , \24580 );
buf \U$20031 ( \25793 , \24580 );
buf \U$20032 ( \25794 , \24580 );
buf \U$20033 ( \25795 , \24580 );
buf \U$20034 ( \25796 , \24580 );
buf \U$20035 ( \25797 , \24580 );
buf \U$20036 ( \25798 , \24580 );
buf \U$20037 ( \25799 , \24580 );
buf \U$20038 ( \25800 , \24580 );
buf \U$20039 ( \25801 , \24580 );
buf \U$20040 ( \25802 , \24580 );
buf \U$20041 ( \25803 , \24580 );
buf \U$20042 ( \25804 , \24580 );
buf \U$20043 ( \25805 , \24580 );
buf \U$20044 ( \25806 , \24580 );
buf \U$20045 ( \25807 , \24580 );
buf \U$20046 ( \25808 , \24580 );
buf \U$20047 ( \25809 , \24580 );
buf \U$20048 ( \25810 , \24580 );
buf \U$20049 ( \25811 , \24580 );
buf \U$20050 ( \25812 , \24580 );
buf \U$20051 ( \25813 , \24580 );
buf \U$20052 ( \25814 , \24580 );
buf \U$20053 ( \25815 , \24580 );
buf \U$20054 ( \25816 , \24580 );
nor \U$20055 ( \25817 , \24608 , \24609 , \24610 , \24611 , \24573 , \24577 , \24580 , \25792 , \25793 , \25794 , \25795 , \25796 , \25797 , \25798 , \25799 , \25800 , \25801 , \25802 , \25803 , \25804 , \25805 , \25806 , \25807 , \25808 , \25809 , \25810 , \25811 , \25812 , \25813 , \25814 , \25815 , \25816 );
and \U$20056 ( \25818 , \7200 , \25817 );
buf \U$20057 ( \25819 , \24580 );
buf \U$20058 ( \25820 , \24580 );
buf \U$20059 ( \25821 , \24580 );
buf \U$20060 ( \25822 , \24580 );
buf \U$20061 ( \25823 , \24580 );
buf \U$20062 ( \25824 , \24580 );
buf \U$20063 ( \25825 , \24580 );
buf \U$20064 ( \25826 , \24580 );
buf \U$20065 ( \25827 , \24580 );
buf \U$20066 ( \25828 , \24580 );
buf \U$20067 ( \25829 , \24580 );
buf \U$20068 ( \25830 , \24580 );
buf \U$20069 ( \25831 , \24580 );
buf \U$20070 ( \25832 , \24580 );
buf \U$20071 ( \25833 , \24580 );
buf \U$20072 ( \25834 , \24580 );
buf \U$20073 ( \25835 , \24580 );
buf \U$20074 ( \25836 , \24580 );
buf \U$20075 ( \25837 , \24580 );
buf \U$20076 ( \25838 , \24580 );
buf \U$20077 ( \25839 , \24580 );
buf \U$20078 ( \25840 , \24580 );
buf \U$20079 ( \25841 , \24580 );
buf \U$20080 ( \25842 , \24580 );
buf \U$20081 ( \25843 , \24580 );
nor \U$20082 ( \25844 , \24567 , \24609 , \24610 , \24611 , \24573 , \24577 , \24580 , \25819 , \25820 , \25821 , \25822 , \25823 , \25824 , \25825 , \25826 , \25827 , \25828 , \25829 , \25830 , \25831 , \25832 , \25833 , \25834 , \25835 , \25836 , \25837 , \25838 , \25839 , \25840 , \25841 , \25842 , \25843 );
and \U$20083 ( \25845 , \8645 , \25844 );
buf \U$20084 ( \25846 , \24580 );
buf \U$20085 ( \25847 , \24580 );
buf \U$20086 ( \25848 , \24580 );
buf \U$20087 ( \25849 , \24580 );
buf \U$20088 ( \25850 , \24580 );
buf \U$20089 ( \25851 , \24580 );
buf \U$20090 ( \25852 , \24580 );
buf \U$20091 ( \25853 , \24580 );
buf \U$20092 ( \25854 , \24580 );
buf \U$20093 ( \25855 , \24580 );
buf \U$20094 ( \25856 , \24580 );
buf \U$20095 ( \25857 , \24580 );
buf \U$20096 ( \25858 , \24580 );
buf \U$20097 ( \25859 , \24580 );
buf \U$20098 ( \25860 , \24580 );
buf \U$20099 ( \25861 , \24580 );
buf \U$20100 ( \25862 , \24580 );
buf \U$20101 ( \25863 , \24580 );
buf \U$20102 ( \25864 , \24580 );
buf \U$20103 ( \25865 , \24580 );
buf \U$20104 ( \25866 , \24580 );
buf \U$20105 ( \25867 , \24580 );
buf \U$20106 ( \25868 , \24580 );
buf \U$20107 ( \25869 , \24580 );
buf \U$20108 ( \25870 , \24580 );
nor \U$20109 ( \25871 , \24608 , \24568 , \24610 , \24611 , \24573 , \24577 , \24580 , \25846 , \25847 , \25848 , \25849 , \25850 , \25851 , \25852 , \25853 , \25854 , \25855 , \25856 , \25857 , \25858 , \25859 , \25860 , \25861 , \25862 , \25863 , \25864 , \25865 , \25866 , \25867 , \25868 , \25869 , \25870 );
and \U$20110 ( \25872 , \8673 , \25871 );
buf \U$20111 ( \25873 , \24580 );
buf \U$20112 ( \25874 , \24580 );
buf \U$20113 ( \25875 , \24580 );
buf \U$20114 ( \25876 , \24580 );
buf \U$20115 ( \25877 , \24580 );
buf \U$20116 ( \25878 , \24580 );
buf \U$20117 ( \25879 , \24580 );
buf \U$20118 ( \25880 , \24580 );
buf \U$20119 ( \25881 , \24580 );
buf \U$20120 ( \25882 , \24580 );
buf \U$20121 ( \25883 , \24580 );
buf \U$20122 ( \25884 , \24580 );
buf \U$20123 ( \25885 , \24580 );
buf \U$20124 ( \25886 , \24580 );
buf \U$20125 ( \25887 , \24580 );
buf \U$20126 ( \25888 , \24580 );
buf \U$20127 ( \25889 , \24580 );
buf \U$20128 ( \25890 , \24580 );
buf \U$20129 ( \25891 , \24580 );
buf \U$20130 ( \25892 , \24580 );
buf \U$20131 ( \25893 , \24580 );
buf \U$20132 ( \25894 , \24580 );
buf \U$20133 ( \25895 , \24580 );
buf \U$20134 ( \25896 , \24580 );
buf \U$20135 ( \25897 , \24580 );
nor \U$20136 ( \25898 , \24567 , \24568 , \24610 , \24611 , \24573 , \24577 , \24580 , \25873 , \25874 , \25875 , \25876 , \25877 , \25878 , \25879 , \25880 , \25881 , \25882 , \25883 , \25884 , \25885 , \25886 , \25887 , \25888 , \25889 , \25890 , \25891 , \25892 , \25893 , \25894 , \25895 , \25896 , \25897 );
and \U$20137 ( \25899 , \8701 , \25898 );
buf \U$20138 ( \25900 , \24580 );
buf \U$20139 ( \25901 , \24580 );
buf \U$20140 ( \25902 , \24580 );
buf \U$20141 ( \25903 , \24580 );
buf \U$20142 ( \25904 , \24580 );
buf \U$20143 ( \25905 , \24580 );
buf \U$20144 ( \25906 , \24580 );
buf \U$20145 ( \25907 , \24580 );
buf \U$20146 ( \25908 , \24580 );
buf \U$20147 ( \25909 , \24580 );
buf \U$20148 ( \25910 , \24580 );
buf \U$20149 ( \25911 , \24580 );
buf \U$20150 ( \25912 , \24580 );
buf \U$20151 ( \25913 , \24580 );
buf \U$20152 ( \25914 , \24580 );
buf \U$20153 ( \25915 , \24580 );
buf \U$20154 ( \25916 , \24580 );
buf \U$20155 ( \25917 , \24580 );
buf \U$20156 ( \25918 , \24580 );
buf \U$20157 ( \25919 , \24580 );
buf \U$20158 ( \25920 , \24580 );
buf \U$20159 ( \25921 , \24580 );
buf \U$20160 ( \25922 , \24580 );
buf \U$20161 ( \25923 , \24580 );
buf \U$20162 ( \25924 , \24580 );
nor \U$20163 ( \25925 , \24608 , \24609 , \24569 , \24611 , \24573 , \24577 , \24580 , \25900 , \25901 , \25902 , \25903 , \25904 , \25905 , \25906 , \25907 , \25908 , \25909 , \25910 , \25911 , \25912 , \25913 , \25914 , \25915 , \25916 , \25917 , \25918 , \25919 , \25920 , \25921 , \25922 , \25923 , \25924 );
and \U$20164 ( \25926 , \8729 , \25925 );
buf \U$20165 ( \25927 , \24580 );
buf \U$20166 ( \25928 , \24580 );
buf \U$20167 ( \25929 , \24580 );
buf \U$20168 ( \25930 , \24580 );
buf \U$20169 ( \25931 , \24580 );
buf \U$20170 ( \25932 , \24580 );
buf \U$20171 ( \25933 , \24580 );
buf \U$20172 ( \25934 , \24580 );
buf \U$20173 ( \25935 , \24580 );
buf \U$20174 ( \25936 , \24580 );
buf \U$20175 ( \25937 , \24580 );
buf \U$20176 ( \25938 , \24580 );
buf \U$20177 ( \25939 , \24580 );
buf \U$20178 ( \25940 , \24580 );
buf \U$20179 ( \25941 , \24580 );
buf \U$20180 ( \25942 , \24580 );
buf \U$20181 ( \25943 , \24580 );
buf \U$20182 ( \25944 , \24580 );
buf \U$20183 ( \25945 , \24580 );
buf \U$20184 ( \25946 , \24580 );
buf \U$20185 ( \25947 , \24580 );
buf \U$20186 ( \25948 , \24580 );
buf \U$20187 ( \25949 , \24580 );
buf \U$20188 ( \25950 , \24580 );
buf \U$20189 ( \25951 , \24580 );
nor \U$20190 ( \25952 , \24567 , \24609 , \24569 , \24611 , \24573 , \24577 , \24580 , \25927 , \25928 , \25929 , \25930 , \25931 , \25932 , \25933 , \25934 , \25935 , \25936 , \25937 , \25938 , \25939 , \25940 , \25941 , \25942 , \25943 , \25944 , \25945 , \25946 , \25947 , \25948 , \25949 , \25950 , \25951 );
and \U$20191 ( \25953 , \8757 , \25952 );
buf \U$20192 ( \25954 , \24580 );
buf \U$20193 ( \25955 , \24580 );
buf \U$20194 ( \25956 , \24580 );
buf \U$20195 ( \25957 , \24580 );
buf \U$20196 ( \25958 , \24580 );
buf \U$20197 ( \25959 , \24580 );
buf \U$20198 ( \25960 , \24580 );
buf \U$20199 ( \25961 , \24580 );
buf \U$20200 ( \25962 , \24580 );
buf \U$20201 ( \25963 , \24580 );
buf \U$20202 ( \25964 , \24580 );
buf \U$20203 ( \25965 , \24580 );
buf \U$20204 ( \25966 , \24580 );
buf \U$20205 ( \25967 , \24580 );
buf \U$20206 ( \25968 , \24580 );
buf \U$20207 ( \25969 , \24580 );
buf \U$20208 ( \25970 , \24580 );
buf \U$20209 ( \25971 , \24580 );
buf \U$20210 ( \25972 , \24580 );
buf \U$20211 ( \25973 , \24580 );
buf \U$20212 ( \25974 , \24580 );
buf \U$20213 ( \25975 , \24580 );
buf \U$20214 ( \25976 , \24580 );
buf \U$20215 ( \25977 , \24580 );
buf \U$20216 ( \25978 , \24580 );
nor \U$20217 ( \25979 , \24608 , \24568 , \24569 , \24611 , \24573 , \24577 , \24580 , \25954 , \25955 , \25956 , \25957 , \25958 , \25959 , \25960 , \25961 , \25962 , \25963 , \25964 , \25965 , \25966 , \25967 , \25968 , \25969 , \25970 , \25971 , \25972 , \25973 , \25974 , \25975 , \25976 , \25977 , \25978 );
and \U$20218 ( \25980 , \8785 , \25979 );
buf \U$20219 ( \25981 , \24580 );
buf \U$20220 ( \25982 , \24580 );
buf \U$20221 ( \25983 , \24580 );
buf \U$20222 ( \25984 , \24580 );
buf \U$20223 ( \25985 , \24580 );
buf \U$20224 ( \25986 , \24580 );
buf \U$20225 ( \25987 , \24580 );
buf \U$20226 ( \25988 , \24580 );
buf \U$20227 ( \25989 , \24580 );
buf \U$20228 ( \25990 , \24580 );
buf \U$20229 ( \25991 , \24580 );
buf \U$20230 ( \25992 , \24580 );
buf \U$20231 ( \25993 , \24580 );
buf \U$20232 ( \25994 , \24580 );
buf \U$20233 ( \25995 , \24580 );
buf \U$20234 ( \25996 , \24580 );
buf \U$20235 ( \25997 , \24580 );
buf \U$20236 ( \25998 , \24580 );
buf \U$20237 ( \25999 , \24580 );
buf \U$20238 ( \26000 , \24580 );
buf \U$20239 ( \26001 , \24580 );
buf \U$20240 ( \26002 , \24580 );
buf \U$20241 ( \26003 , \24580 );
buf \U$20242 ( \26004 , \24580 );
buf \U$20243 ( \26005 , \24580 );
nor \U$20244 ( \26006 , \24567 , \24568 , \24569 , \24611 , \24573 , \24577 , \24580 , \25981 , \25982 , \25983 , \25984 , \25985 , \25986 , \25987 , \25988 , \25989 , \25990 , \25991 , \25992 , \25993 , \25994 , \25995 , \25996 , \25997 , \25998 , \25999 , \26000 , \26001 , \26002 , \26003 , \26004 , \26005 );
and \U$20245 ( \26007 , \8813 , \26006 );
buf \U$20246 ( \26008 , \24580 );
buf \U$20247 ( \26009 , \24580 );
buf \U$20248 ( \26010 , \24580 );
buf \U$20249 ( \26011 , \24580 );
buf \U$20250 ( \26012 , \24580 );
buf \U$20251 ( \26013 , \24580 );
buf \U$20252 ( \26014 , \24580 );
buf \U$20253 ( \26015 , \24580 );
buf \U$20254 ( \26016 , \24580 );
buf \U$20255 ( \26017 , \24580 );
buf \U$20256 ( \26018 , \24580 );
buf \U$20257 ( \26019 , \24580 );
buf \U$20258 ( \26020 , \24580 );
buf \U$20259 ( \26021 , \24580 );
buf \U$20260 ( \26022 , \24580 );
buf \U$20261 ( \26023 , \24580 );
buf \U$20262 ( \26024 , \24580 );
buf \U$20263 ( \26025 , \24580 );
buf \U$20264 ( \26026 , \24580 );
buf \U$20265 ( \26027 , \24580 );
buf \U$20266 ( \26028 , \24580 );
buf \U$20267 ( \26029 , \24580 );
buf \U$20268 ( \26030 , \24580 );
buf \U$20269 ( \26031 , \24580 );
buf \U$20270 ( \26032 , \24580 );
nor \U$20271 ( \26033 , \24608 , \24609 , \24610 , \24570 , \24573 , \24577 , \24580 , \26008 , \26009 , \26010 , \26011 , \26012 , \26013 , \26014 , \26015 , \26016 , \26017 , \26018 , \26019 , \26020 , \26021 , \26022 , \26023 , \26024 , \26025 , \26026 , \26027 , \26028 , \26029 , \26030 , \26031 , \26032 );
and \U$20272 ( \26034 , \8841 , \26033 );
buf \U$20273 ( \26035 , \24580 );
buf \U$20274 ( \26036 , \24580 );
buf \U$20275 ( \26037 , \24580 );
buf \U$20276 ( \26038 , \24580 );
buf \U$20277 ( \26039 , \24580 );
buf \U$20278 ( \26040 , \24580 );
buf \U$20279 ( \26041 , \24580 );
buf \U$20280 ( \26042 , \24580 );
buf \U$20281 ( \26043 , \24580 );
buf \U$20282 ( \26044 , \24580 );
buf \U$20283 ( \26045 , \24580 );
buf \U$20284 ( \26046 , \24580 );
buf \U$20285 ( \26047 , \24580 );
buf \U$20286 ( \26048 , \24580 );
buf \U$20287 ( \26049 , \24580 );
buf \U$20288 ( \26050 , \24580 );
buf \U$20289 ( \26051 , \24580 );
buf \U$20290 ( \26052 , \24580 );
buf \U$20291 ( \26053 , \24580 );
buf \U$20292 ( \26054 , \24580 );
buf \U$20293 ( \26055 , \24580 );
buf \U$20294 ( \26056 , \24580 );
buf \U$20295 ( \26057 , \24580 );
buf \U$20296 ( \26058 , \24580 );
buf \U$20297 ( \26059 , \24580 );
nor \U$20298 ( \26060 , \24567 , \24609 , \24610 , \24570 , \24573 , \24577 , \24580 , \26035 , \26036 , \26037 , \26038 , \26039 , \26040 , \26041 , \26042 , \26043 , \26044 , \26045 , \26046 , \26047 , \26048 , \26049 , \26050 , \26051 , \26052 , \26053 , \26054 , \26055 , \26056 , \26057 , \26058 , \26059 );
and \U$20299 ( \26061 , \8869 , \26060 );
buf \U$20300 ( \26062 , \24580 );
buf \U$20301 ( \26063 , \24580 );
buf \U$20302 ( \26064 , \24580 );
buf \U$20303 ( \26065 , \24580 );
buf \U$20304 ( \26066 , \24580 );
buf \U$20305 ( \26067 , \24580 );
buf \U$20306 ( \26068 , \24580 );
buf \U$20307 ( \26069 , \24580 );
buf \U$20308 ( \26070 , \24580 );
buf \U$20309 ( \26071 , \24580 );
buf \U$20310 ( \26072 , \24580 );
buf \U$20311 ( \26073 , \24580 );
buf \U$20312 ( \26074 , \24580 );
buf \U$20313 ( \26075 , \24580 );
buf \U$20314 ( \26076 , \24580 );
buf \U$20315 ( \26077 , \24580 );
buf \U$20316 ( \26078 , \24580 );
buf \U$20317 ( \26079 , \24580 );
buf \U$20318 ( \26080 , \24580 );
buf \U$20319 ( \26081 , \24580 );
buf \U$20320 ( \26082 , \24580 );
buf \U$20321 ( \26083 , \24580 );
buf \U$20322 ( \26084 , \24580 );
buf \U$20323 ( \26085 , \24580 );
buf \U$20324 ( \26086 , \24580 );
nor \U$20325 ( \26087 , \24608 , \24568 , \24610 , \24570 , \24573 , \24577 , \24580 , \26062 , \26063 , \26064 , \26065 , \26066 , \26067 , \26068 , \26069 , \26070 , \26071 , \26072 , \26073 , \26074 , \26075 , \26076 , \26077 , \26078 , \26079 , \26080 , \26081 , \26082 , \26083 , \26084 , \26085 , \26086 );
and \U$20326 ( \26088 , \8897 , \26087 );
buf \U$20327 ( \26089 , \24580 );
buf \U$20328 ( \26090 , \24580 );
buf \U$20329 ( \26091 , \24580 );
buf \U$20330 ( \26092 , \24580 );
buf \U$20331 ( \26093 , \24580 );
buf \U$20332 ( \26094 , \24580 );
buf \U$20333 ( \26095 , \24580 );
buf \U$20334 ( \26096 , \24580 );
buf \U$20335 ( \26097 , \24580 );
buf \U$20336 ( \26098 , \24580 );
buf \U$20337 ( \26099 , \24580 );
buf \U$20338 ( \26100 , \24580 );
buf \U$20339 ( \26101 , \24580 );
buf \U$20340 ( \26102 , \24580 );
buf \U$20341 ( \26103 , \24580 );
buf \U$20342 ( \26104 , \24580 );
buf \U$20343 ( \26105 , \24580 );
buf \U$20344 ( \26106 , \24580 );
buf \U$20345 ( \26107 , \24580 );
buf \U$20346 ( \26108 , \24580 );
buf \U$20347 ( \26109 , \24580 );
buf \U$20348 ( \26110 , \24580 );
buf \U$20349 ( \26111 , \24580 );
buf \U$20350 ( \26112 , \24580 );
buf \U$20351 ( \26113 , \24580 );
nor \U$20352 ( \26114 , \24567 , \24568 , \24610 , \24570 , \24573 , \24577 , \24580 , \26089 , \26090 , \26091 , \26092 , \26093 , \26094 , \26095 , \26096 , \26097 , \26098 , \26099 , \26100 , \26101 , \26102 , \26103 , \26104 , \26105 , \26106 , \26107 , \26108 , \26109 , \26110 , \26111 , \26112 , \26113 );
and \U$20353 ( \26115 , \8925 , \26114 );
buf \U$20354 ( \26116 , \24580 );
buf \U$20355 ( \26117 , \24580 );
buf \U$20356 ( \26118 , \24580 );
buf \U$20357 ( \26119 , \24580 );
buf \U$20358 ( \26120 , \24580 );
buf \U$20359 ( \26121 , \24580 );
buf \U$20360 ( \26122 , \24580 );
buf \U$20361 ( \26123 , \24580 );
buf \U$20362 ( \26124 , \24580 );
buf \U$20363 ( \26125 , \24580 );
buf \U$20364 ( \26126 , \24580 );
buf \U$20365 ( \26127 , \24580 );
buf \U$20366 ( \26128 , \24580 );
buf \U$20367 ( \26129 , \24580 );
buf \U$20368 ( \26130 , \24580 );
buf \U$20369 ( \26131 , \24580 );
buf \U$20370 ( \26132 , \24580 );
buf \U$20371 ( \26133 , \24580 );
buf \U$20372 ( \26134 , \24580 );
buf \U$20373 ( \26135 , \24580 );
buf \U$20374 ( \26136 , \24580 );
buf \U$20375 ( \26137 , \24580 );
buf \U$20376 ( \26138 , \24580 );
buf \U$20377 ( \26139 , \24580 );
buf \U$20378 ( \26140 , \24580 );
nor \U$20379 ( \26141 , \24608 , \24609 , \24569 , \24570 , \24573 , \24577 , \24580 , \26116 , \26117 , \26118 , \26119 , \26120 , \26121 , \26122 , \26123 , \26124 , \26125 , \26126 , \26127 , \26128 , \26129 , \26130 , \26131 , \26132 , \26133 , \26134 , \26135 , \26136 , \26137 , \26138 , \26139 , \26140 );
and \U$20380 ( \26142 , \8953 , \26141 );
buf \U$20381 ( \26143 , \24580 );
buf \U$20382 ( \26144 , \24580 );
buf \U$20383 ( \26145 , \24580 );
buf \U$20384 ( \26146 , \24580 );
buf \U$20385 ( \26147 , \24580 );
buf \U$20386 ( \26148 , \24580 );
buf \U$20387 ( \26149 , \24580 );
buf \U$20388 ( \26150 , \24580 );
buf \U$20389 ( \26151 , \24580 );
buf \U$20390 ( \26152 , \24580 );
buf \U$20391 ( \26153 , \24580 );
buf \U$20392 ( \26154 , \24580 );
buf \U$20393 ( \26155 , \24580 );
buf \U$20394 ( \26156 , \24580 );
buf \U$20395 ( \26157 , \24580 );
buf \U$20396 ( \26158 , \24580 );
buf \U$20397 ( \26159 , \24580 );
buf \U$20398 ( \26160 , \24580 );
buf \U$20399 ( \26161 , \24580 );
buf \U$20400 ( \26162 , \24580 );
buf \U$20401 ( \26163 , \24580 );
buf \U$20402 ( \26164 , \24580 );
buf \U$20403 ( \26165 , \24580 );
buf \U$20404 ( \26166 , \24580 );
buf \U$20405 ( \26167 , \24580 );
nor \U$20406 ( \26168 , \24567 , \24609 , \24569 , \24570 , \24573 , \24577 , \24580 , \26143 , \26144 , \26145 , \26146 , \26147 , \26148 , \26149 , \26150 , \26151 , \26152 , \26153 , \26154 , \26155 , \26156 , \26157 , \26158 , \26159 , \26160 , \26161 , \26162 , \26163 , \26164 , \26165 , \26166 , \26167 );
and \U$20407 ( \26169 , \8981 , \26168 );
buf \U$20408 ( \26170 , \24580 );
buf \U$20409 ( \26171 , \24580 );
buf \U$20410 ( \26172 , \24580 );
buf \U$20411 ( \26173 , \24580 );
buf \U$20412 ( \26174 , \24580 );
buf \U$20413 ( \26175 , \24580 );
buf \U$20414 ( \26176 , \24580 );
buf \U$20415 ( \26177 , \24580 );
buf \U$20416 ( \26178 , \24580 );
buf \U$20417 ( \26179 , \24580 );
buf \U$20418 ( \26180 , \24580 );
buf \U$20419 ( \26181 , \24580 );
buf \U$20420 ( \26182 , \24580 );
buf \U$20421 ( \26183 , \24580 );
buf \U$20422 ( \26184 , \24580 );
buf \U$20423 ( \26185 , \24580 );
buf \U$20424 ( \26186 , \24580 );
buf \U$20425 ( \26187 , \24580 );
buf \U$20426 ( \26188 , \24580 );
buf \U$20427 ( \26189 , \24580 );
buf \U$20428 ( \26190 , \24580 );
buf \U$20429 ( \26191 , \24580 );
buf \U$20430 ( \26192 , \24580 );
buf \U$20431 ( \26193 , \24580 );
buf \U$20432 ( \26194 , \24580 );
nor \U$20433 ( \26195 , \24608 , \24568 , \24569 , \24570 , \24573 , \24577 , \24580 , \26170 , \26171 , \26172 , \26173 , \26174 , \26175 , \26176 , \26177 , \26178 , \26179 , \26180 , \26181 , \26182 , \26183 , \26184 , \26185 , \26186 , \26187 , \26188 , \26189 , \26190 , \26191 , \26192 , \26193 , \26194 );
and \U$20434 ( \26196 , \9009 , \26195 );
or \U$20435 ( \26197 , \25791 , \25818 , \25845 , \25872 , \25899 , \25926 , \25953 , \25980 , \26007 , \26034 , \26061 , \26088 , \26115 , \26142 , \26169 , \26196 );
buf \U$20436 ( \26198 , \24580 );
not \U$20437 ( \26199 , \26198 );
buf \U$20438 ( \26200 , \24568 );
buf \U$20439 ( \26201 , \24569 );
buf \U$20440 ( \26202 , \24570 );
buf \U$20441 ( \26203 , \24573 );
buf \U$20442 ( \26204 , \24577 );
buf \U$20443 ( \26205 , \24580 );
buf \U$20444 ( \26206 , \24580 );
buf \U$20445 ( \26207 , \24580 );
buf \U$20446 ( \26208 , \24580 );
buf \U$20447 ( \26209 , \24580 );
buf \U$20448 ( \26210 , \24580 );
buf \U$20449 ( \26211 , \24580 );
buf \U$20450 ( \26212 , \24580 );
buf \U$20451 ( \26213 , \24580 );
buf \U$20452 ( \26214 , \24580 );
buf \U$20453 ( \26215 , \24580 );
buf \U$20454 ( \26216 , \24580 );
buf \U$20455 ( \26217 , \24580 );
buf \U$20456 ( \26218 , \24580 );
buf \U$20457 ( \26219 , \24580 );
buf \U$20458 ( \26220 , \24580 );
buf \U$20459 ( \26221 , \24580 );
buf \U$20460 ( \26222 , \24580 );
buf \U$20461 ( \26223 , \24580 );
buf \U$20462 ( \26224 , \24580 );
buf \U$20463 ( \26225 , \24580 );
buf \U$20464 ( \26226 , \24580 );
buf \U$20465 ( \26227 , \24580 );
buf \U$20466 ( \26228 , \24580 );
buf \U$20467 ( \26229 , \24580 );
buf \U$20468 ( \26230 , \24567 );
or \U$20469 ( \26231 , \26200 , \26201 , \26202 , \26203 , \26204 , \26205 , \26206 , \26207 , \26208 , \26209 , \26210 , \26211 , \26212 , \26213 , \26214 , \26215 , \26216 , \26217 , \26218 , \26219 , \26220 , \26221 , \26222 , \26223 , \26224 , \26225 , \26226 , \26227 , \26228 , \26229 , \26230 );
nand \U$20470 ( \26232 , \26199 , \26231 );
buf \U$20471 ( \26233 , \26232 );
buf \U$20472 ( \26234 , \24580 );
not \U$20473 ( \26235 , \26234 );
buf \U$20474 ( \26236 , \24577 );
buf \U$20475 ( \26237 , \24580 );
buf \U$20476 ( \26238 , \24580 );
buf \U$20477 ( \26239 , \24580 );
buf \U$20478 ( \26240 , \24580 );
buf \U$20479 ( \26241 , \24580 );
buf \U$20480 ( \26242 , \24580 );
buf \U$20481 ( \26243 , \24580 );
buf \U$20482 ( \26244 , \24580 );
buf \U$20483 ( \26245 , \24580 );
buf \U$20484 ( \26246 , \24580 );
buf \U$20485 ( \26247 , \24580 );
buf \U$20486 ( \26248 , \24580 );
buf \U$20487 ( \26249 , \24580 );
buf \U$20488 ( \26250 , \24580 );
buf \U$20489 ( \26251 , \24580 );
buf \U$20490 ( \26252 , \24580 );
buf \U$20491 ( \26253 , \24580 );
buf \U$20492 ( \26254 , \24580 );
buf \U$20493 ( \26255 , \24580 );
buf \U$20494 ( \26256 , \24580 );
buf \U$20495 ( \26257 , \24580 );
buf \U$20496 ( \26258 , \24580 );
buf \U$20497 ( \26259 , \24580 );
buf \U$20498 ( \26260 , \24580 );
buf \U$20499 ( \26261 , \24580 );
buf \U$20500 ( \26262 , \24573 );
buf \U$20501 ( \26263 , \24567 );
buf \U$20502 ( \26264 , \24568 );
buf \U$20503 ( \26265 , \24569 );
buf \U$20504 ( \26266 , \24570 );
or \U$20505 ( \26267 , \26263 , \26264 , \26265 , \26266 );
and \U$20506 ( \26268 , \26262 , \26267 );
or \U$20507 ( \26269 , \26236 , \26237 , \26238 , \26239 , \26240 , \26241 , \26242 , \26243 , \26244 , \26245 , \26246 , \26247 , \26248 , \26249 , \26250 , \26251 , \26252 , \26253 , \26254 , \26255 , \26256 , \26257 , \26258 , \26259 , \26260 , \26261 , \26268 );
and \U$20508 ( \26270 , \26235 , \26269 );
buf \U$20509 ( \26271 , \26270 );
or \U$20510 ( \26272 , \26233 , \26271 );
_DC g7d99 ( \26273_nG7d99 , \26197 , \26272 );
buf \U$20511 ( \26274 , \26273_nG7d99 );
xor \U$20512 ( \26275 , \25764 , \26274 );
buf \U$20513 ( \26276 , RIb7af5b8_255);
and \U$20514 ( \26277 , \7207 , \25790 );
and \U$20515 ( \26278 , \7209 , \25817 );
and \U$20516 ( \26279 , \9119 , \25844 );
and \U$20517 ( \26280 , \9121 , \25871 );
and \U$20518 ( \26281 , \9123 , \25898 );
and \U$20519 ( \26282 , \9125 , \25925 );
and \U$20520 ( \26283 , \9127 , \25952 );
and \U$20521 ( \26284 , \9129 , \25979 );
and \U$20522 ( \26285 , \9131 , \26006 );
and \U$20523 ( \26286 , \9133 , \26033 );
and \U$20524 ( \26287 , \9135 , \26060 );
and \U$20525 ( \26288 , \9137 , \26087 );
and \U$20526 ( \26289 , \9139 , \26114 );
and \U$20527 ( \26290 , \9141 , \26141 );
and \U$20528 ( \26291 , \9143 , \26168 );
and \U$20529 ( \26292 , \9145 , \26195 );
or \U$20530 ( \26293 , \26277 , \26278 , \26279 , \26280 , \26281 , \26282 , \26283 , \26284 , \26285 , \26286 , \26287 , \26288 , \26289 , \26290 , \26291 , \26292 );
_DC g7dae ( \26294_nG7dae , \26293 , \26272 );
buf \U$20531 ( \26295 , \26294_nG7dae );
xor \U$20532 ( \26296 , \26276 , \26295 );
or \U$20533 ( \26297 , \26275 , \26296 );
buf \U$20534 ( \26298 , RIb7af540_256);
and \U$20535 ( \26299 , \7217 , \25790 );
and \U$20536 ( \26300 , \7219 , \25817 );
and \U$20537 ( \26301 , \9155 , \25844 );
and \U$20538 ( \26302 , \9157 , \25871 );
and \U$20539 ( \26303 , \9159 , \25898 );
and \U$20540 ( \26304 , \9161 , \25925 );
and \U$20541 ( \26305 , \9163 , \25952 );
and \U$20542 ( \26306 , \9165 , \25979 );
and \U$20543 ( \26307 , \9167 , \26006 );
and \U$20544 ( \26308 , \9169 , \26033 );
and \U$20545 ( \26309 , \9171 , \26060 );
and \U$20546 ( \26310 , \9173 , \26087 );
and \U$20547 ( \26311 , \9175 , \26114 );
and \U$20548 ( \26312 , \9177 , \26141 );
and \U$20549 ( \26313 , \9179 , \26168 );
and \U$20550 ( \26314 , \9181 , \26195 );
or \U$20551 ( \26315 , \26299 , \26300 , \26301 , \26302 , \26303 , \26304 , \26305 , \26306 , \26307 , \26308 , \26309 , \26310 , \26311 , \26312 , \26313 , \26314 );
_DC g7dc4 ( \26316_nG7dc4 , \26315 , \26272 );
buf \U$20552 ( \26317 , \26316_nG7dc4 );
xor \U$20553 ( \26318 , \26298 , \26317 );
or \U$20554 ( \26319 , \26297 , \26318 );
buf \U$20555 ( \26320 , RIb7af4c8_257);
and \U$20556 ( \26321 , \7227 , \25790 );
and \U$20557 ( \26322 , \7229 , \25817 );
and \U$20558 ( \26323 , \9191 , \25844 );
and \U$20559 ( \26324 , \9193 , \25871 );
and \U$20560 ( \26325 , \9195 , \25898 );
and \U$20561 ( \26326 , \9197 , \25925 );
and \U$20562 ( \26327 , \9199 , \25952 );
and \U$20563 ( \26328 , \9201 , \25979 );
and \U$20564 ( \26329 , \9203 , \26006 );
and \U$20565 ( \26330 , \9205 , \26033 );
and \U$20566 ( \26331 , \9207 , \26060 );
and \U$20567 ( \26332 , \9209 , \26087 );
and \U$20568 ( \26333 , \9211 , \26114 );
and \U$20569 ( \26334 , \9213 , \26141 );
and \U$20570 ( \26335 , \9215 , \26168 );
and \U$20571 ( \26336 , \9217 , \26195 );
or \U$20572 ( \26337 , \26321 , \26322 , \26323 , \26324 , \26325 , \26326 , \26327 , \26328 , \26329 , \26330 , \26331 , \26332 , \26333 , \26334 , \26335 , \26336 );
_DC g7dda ( \26338_nG7dda , \26337 , \26272 );
buf \U$20573 ( \26339 , \26338_nG7dda );
xor \U$20574 ( \26340 , \26320 , \26339 );
or \U$20575 ( \26341 , \26319 , \26340 );
buf \U$20576 ( \26342 , RIb7af450_258);
and \U$20577 ( \26343 , \7237 , \25790 );
and \U$20578 ( \26344 , \7239 , \25817 );
and \U$20579 ( \26345 , \9227 , \25844 );
and \U$20580 ( \26346 , \9229 , \25871 );
and \U$20581 ( \26347 , \9231 , \25898 );
and \U$20582 ( \26348 , \9233 , \25925 );
and \U$20583 ( \26349 , \9235 , \25952 );
and \U$20584 ( \26350 , \9237 , \25979 );
and \U$20585 ( \26351 , \9239 , \26006 );
and \U$20586 ( \26352 , \9241 , \26033 );
and \U$20587 ( \26353 , \9243 , \26060 );
and \U$20588 ( \26354 , \9245 , \26087 );
and \U$20589 ( \26355 , \9247 , \26114 );
and \U$20590 ( \26356 , \9249 , \26141 );
and \U$20591 ( \26357 , \9251 , \26168 );
and \U$20592 ( \26358 , \9253 , \26195 );
or \U$20593 ( \26359 , \26343 , \26344 , \26345 , \26346 , \26347 , \26348 , \26349 , \26350 , \26351 , \26352 , \26353 , \26354 , \26355 , \26356 , \26357 , \26358 );
_DC g7df0 ( \26360_nG7df0 , \26359 , \26272 );
buf \U$20594 ( \26361 , \26360_nG7df0 );
xor \U$20595 ( \26362 , \26342 , \26361 );
or \U$20596 ( \26363 , \26341 , \26362 );
buf \U$20597 ( \26364 , RIb7af3d8_259);
and \U$20598 ( \26365 , \7247 , \25790 );
and \U$20599 ( \26366 , \7249 , \25817 );
and \U$20600 ( \26367 , \9263 , \25844 );
and \U$20601 ( \26368 , \9265 , \25871 );
and \U$20602 ( \26369 , \9267 , \25898 );
and \U$20603 ( \26370 , \9269 , \25925 );
and \U$20604 ( \26371 , \9271 , \25952 );
and \U$20605 ( \26372 , \9273 , \25979 );
and \U$20606 ( \26373 , \9275 , \26006 );
and \U$20607 ( \26374 , \9277 , \26033 );
and \U$20608 ( \26375 , \9279 , \26060 );
and \U$20609 ( \26376 , \9281 , \26087 );
and \U$20610 ( \26377 , \9283 , \26114 );
and \U$20611 ( \26378 , \9285 , \26141 );
and \U$20612 ( \26379 , \9287 , \26168 );
and \U$20613 ( \26380 , \9289 , \26195 );
or \U$20614 ( \26381 , \26365 , \26366 , \26367 , \26368 , \26369 , \26370 , \26371 , \26372 , \26373 , \26374 , \26375 , \26376 , \26377 , \26378 , \26379 , \26380 );
_DC g7e06 ( \26382_nG7e06 , \26381 , \26272 );
buf \U$20615 ( \26383 , \26382_nG7e06 );
xor \U$20616 ( \26384 , \26364 , \26383 );
or \U$20617 ( \26385 , \26363 , \26384 );
buf \U$20618 ( \26386 , RIb7a5bf8_260);
and \U$20619 ( \26387 , \7257 , \25790 );
and \U$20620 ( \26388 , \7259 , \25817 );
and \U$20621 ( \26389 , \9299 , \25844 );
and \U$20622 ( \26390 , \9301 , \25871 );
and \U$20623 ( \26391 , \9303 , \25898 );
and \U$20624 ( \26392 , \9305 , \25925 );
and \U$20625 ( \26393 , \9307 , \25952 );
and \U$20626 ( \26394 , \9309 , \25979 );
and \U$20627 ( \26395 , \9311 , \26006 );
and \U$20628 ( \26396 , \9313 , \26033 );
and \U$20629 ( \26397 , \9315 , \26060 );
and \U$20630 ( \26398 , \9317 , \26087 );
and \U$20631 ( \26399 , \9319 , \26114 );
and \U$20632 ( \26400 , \9321 , \26141 );
and \U$20633 ( \26401 , \9323 , \26168 );
and \U$20634 ( \26402 , \9325 , \26195 );
or \U$20635 ( \26403 , \26387 , \26388 , \26389 , \26390 , \26391 , \26392 , \26393 , \26394 , \26395 , \26396 , \26397 , \26398 , \26399 , \26400 , \26401 , \26402 );
_DC g7e1c ( \26404_nG7e1c , \26403 , \26272 );
buf \U$20636 ( \26405 , \26404_nG7e1c );
xor \U$20637 ( \26406 , \26386 , \26405 );
or \U$20638 ( \26407 , \26385 , \26406 );
buf \U$20639 ( \26408 , RIb7a0c48_261);
and \U$20640 ( \26409 , \7267 , \25790 );
and \U$20641 ( \26410 , \7269 , \25817 );
and \U$20642 ( \26411 , \9335 , \25844 );
and \U$20643 ( \26412 , \9337 , \25871 );
and \U$20644 ( \26413 , \9339 , \25898 );
and \U$20645 ( \26414 , \9341 , \25925 );
and \U$20646 ( \26415 , \9343 , \25952 );
and \U$20647 ( \26416 , \9345 , \25979 );
and \U$20648 ( \26417 , \9347 , \26006 );
and \U$20649 ( \26418 , \9349 , \26033 );
and \U$20650 ( \26419 , \9351 , \26060 );
and \U$20651 ( \26420 , \9353 , \26087 );
and \U$20652 ( \26421 , \9355 , \26114 );
and \U$20653 ( \26422 , \9357 , \26141 );
and \U$20654 ( \26423 , \9359 , \26168 );
and \U$20655 ( \26424 , \9361 , \26195 );
or \U$20656 ( \26425 , \26409 , \26410 , \26411 , \26412 , \26413 , \26414 , \26415 , \26416 , \26417 , \26418 , \26419 , \26420 , \26421 , \26422 , \26423 , \26424 );
_DC g7e32 ( \26426_nG7e32 , \26425 , \26272 );
buf \U$20657 ( \26427 , \26426_nG7e32 );
xor \U$20658 ( \26428 , \26408 , \26427 );
or \U$20659 ( \26429 , \26407 , \26428 );
not \U$20660 ( \26430 , \26429 );
buf \U$20661 ( \26431 , \26430 );
and \U$20662 ( \26432 , \25763 , \26431 );
_HMUX g7e39 ( \26433_nG7e39 , \24246_nG75a6 , \24567 , \26432 );
buf \U$20663 ( \26434 , \24267 );
buf \U$20664 ( \26435 , \24264 );
buf \U$20665 ( \26436 , \24249 );
buf \U$20666 ( \26437 , \24252 );
buf \U$20667 ( \26438 , \24256 );
buf \U$20668 ( \26439 , \24260 );
or \U$20669 ( \26440 , \26436 , \26437 , \26438 , \26439 );
and \U$20670 ( \26441 , \26435 , \26440 );
or \U$20671 ( \26442 , \26434 , \26441 );
buf \U$20672 ( \26443 , \26442 );
_HMUX g7e44 ( \26444_nG7e44 , \24566_nG76e6 , \26433_nG7e39 , \26443 );
buf \U$20673 ( \26445 , RIe5319e0_6884);
buf \U$20675 ( \26446 , \26445 );
buf \U$20676 ( \26447 , RIe549ef0_6842);
not \U$20677 ( \26448 , \26447 );
buf \U$20678 ( \26449 , \26448 );
buf \U$20679 ( \26450 , RIe549770_6843);
xnor \U$20680 ( \26451 , \26450 , \26447 );
buf \U$20681 ( \26452 , \26451 );
buf \U$20682 ( \26453 , RIe548ff0_6844);
or \U$20683 ( \26454 , \26450 , \26447 );
xor \U$20684 ( \26455 , \26453 , \26454 );
buf \U$20685 ( \26456 , \26455 );
buf \U$20686 ( \26457 , RIea91330_6888);
and \U$20687 ( \26458 , \26453 , \26454 );
xor \U$20688 ( \26459 , \26457 , \26458 );
buf \U$20689 ( \26460 , \26459 );
not \U$20690 ( \26461 , \26460 );
and \U$20691 ( \26462 , \26457 , \26458 );
buf \U$20692 ( \26463 , \26462 );
nor \U$20693 ( \26464 , \26446 , \26449 , \26452 , \26456 , \26461 , \26463 );
and \U$20694 ( \26465 , RIe5329d0_6883, \26464 );
not \U$20695 ( \26466 , \26463 );
and \U$20696 ( \26467 , \26446 , \26449 , \26452 , \26456 , \26461 , \26466 );
and \U$20697 ( \26468 , RIeb72150_6905, \26467 );
not \U$20698 ( \26469 , \26446 );
and \U$20699 ( \26470 , \26469 , \26449 , \26452 , \26456 , \26461 , \26466 );
and \U$20700 ( \26471 , RIeab80c0_6897, \26470 );
not \U$20701 ( \26472 , \26449 );
and \U$20702 ( \26473 , \26446 , \26472 , \26452 , \26456 , \26461 , \26466 );
and \U$20703 ( \26474 , RIe5331c8_6882, \26473 );
and \U$20704 ( \26475 , \26469 , \26472 , \26452 , \26456 , \26461 , \26466 );
and \U$20705 ( \26476 , RIe5339c0_6881, \26475 );
not \U$20706 ( \26477 , \26452 );
and \U$20707 ( \26478 , \26446 , \26449 , \26477 , \26456 , \26461 , \26466 );
and \U$20708 ( \26479 , RIeab87c8_6898, \26478 );
and \U$20709 ( \26480 , \26469 , \26449 , \26477 , \26456 , \26461 , \26466 );
and \U$20710 ( \26481 , RIe5341b8_6880, \26480 );
and \U$20711 ( \26482 , \26446 , \26472 , \26477 , \26456 , \26461 , \26466 );
and \U$20712 ( \26483 , RIe5349b0_6879, \26482 );
and \U$20713 ( \26484 , \26469 , \26472 , \26477 , \26456 , \26461 , \26466 );
and \U$20714 ( \26485 , RIea94af8_6890, \26484 );
nor \U$20715 ( \26486 , \26469 , \26472 , \26477 , \26456 , \26460 , \26463 );
and \U$20716 ( \26487 , RIe5351a8_6878, \26486 );
nor \U$20717 ( \26488 , \26446 , \26472 , \26477 , \26456 , \26460 , \26463 );
and \U$20718 ( \26489 , RIe5359a0_6877, \26488 );
or \U$20724 ( \26490 , \26465 , \26468 , \26471 , \26474 , \26476 , \26479 , \26481 , \26483 , \26485 , \26487 , \26489 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
buf \U$20726 ( \26491 , \26463 );
buf \U$20727 ( \26492 , \26460 );
buf \U$20728 ( \26493 , \26446 );
buf \U$20729 ( \26494 , \26449 );
buf \U$20730 ( \26495 , \26452 );
buf \U$20731 ( \26496 , \26456 );
or \U$20732 ( \26497 , \26493 , \26494 , \26495 , \26496 );
and \U$20733 ( \26498 , \26492 , \26497 );
or \U$20734 ( \26499 , \26491 , \26498 );
buf \U$20735 ( \26500 , \26499 );
or \U$20736 ( \26501 , 1'b0 , \26500 );
_DC g7e7f ( \26502_nG7e7f , \26490 , \26501 );
not \U$20737 ( \26503 , \26502_nG7e7f );
buf \U$20738 ( \26504 , RIb7b9608_246);
and \U$20739 ( \26505 , \7117 , \26464 );
and \U$20740 ( \26506 , \7119 , \26467 );
and \U$20741 ( \26507 , \7864 , \26470 );
and \U$20742 ( \26508 , \7892 , \26473 );
and \U$20743 ( \26509 , \7920 , \26475 );
and \U$20744 ( \26510 , \7948 , \26478 );
and \U$20745 ( \26511 , \7976 , \26480 );
and \U$20746 ( \26512 , \8004 , \26482 );
and \U$20747 ( \26513 , \8032 , \26484 );
and \U$20748 ( \26514 , \8060 , \26486 );
and \U$20749 ( \26515 , \8088 , \26488 );
or \U$20755 ( \26516 , \26505 , \26506 , \26507 , \26508 , \26509 , \26510 , \26511 , \26512 , \26513 , \26514 , \26515 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7e8e ( \26517_nG7e8e , \26516 , \26501 );
buf \U$20756 ( \26518 , \26517_nG7e8e );
xor \U$20757 ( \26519 , \26504 , \26518 );
buf \U$20758 ( \26520 , RIb7b9590_247);
and \U$20759 ( \26521 , \7126 , \26464 );
and \U$20760 ( \26522 , \7128 , \26467 );
and \U$20761 ( \26523 , \8338 , \26470 );
and \U$20762 ( \26524 , \8340 , \26473 );
and \U$20763 ( \26525 , \8342 , \26475 );
and \U$20764 ( \26526 , \8344 , \26478 );
and \U$20765 ( \26527 , \8346 , \26480 );
and \U$20766 ( \26528 , \8348 , \26482 );
and \U$20767 ( \26529 , \8350 , \26484 );
and \U$20768 ( \26530 , \8352 , \26486 );
and \U$20769 ( \26531 , \8354 , \26488 );
or \U$20775 ( \26532 , \26521 , \26522 , \26523 , \26524 , \26525 , \26526 , \26527 , \26528 , \26529 , \26530 , \26531 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7e9e ( \26533_nG7e9e , \26532 , \26501 );
buf \U$20776 ( \26534 , \26533_nG7e9e );
xor \U$20777 ( \26535 , \26520 , \26534 );
or \U$20778 ( \26536 , \26519 , \26535 );
buf \U$20779 ( \26537 , RIb7b9518_248);
and \U$20780 ( \26538 , \7136 , \26464 );
and \U$20781 ( \26539 , \7138 , \26467 );
and \U$20782 ( \26540 , \8374 , \26470 );
and \U$20783 ( \26541 , \8376 , \26473 );
and \U$20784 ( \26542 , \8378 , \26475 );
and \U$20785 ( \26543 , \8380 , \26478 );
and \U$20786 ( \26544 , \8382 , \26480 );
and \U$20787 ( \26545 , \8384 , \26482 );
and \U$20788 ( \26546 , \8386 , \26484 );
and \U$20789 ( \26547 , \8388 , \26486 );
and \U$20790 ( \26548 , \8390 , \26488 );
or \U$20796 ( \26549 , \26538 , \26539 , \26540 , \26541 , \26542 , \26543 , \26544 , \26545 , \26546 , \26547 , \26548 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7eaf ( \26550_nG7eaf , \26549 , \26501 );
buf \U$20797 ( \26551 , \26550_nG7eaf );
xor \U$20798 ( \26552 , \26537 , \26551 );
or \U$20799 ( \26553 , \26536 , \26552 );
buf \U$20800 ( \26554 , RIb7b94a0_249);
and \U$20801 ( \26555 , \7146 , \26464 );
and \U$20802 ( \26556 , \7148 , \26467 );
and \U$20803 ( \26557 , \8410 , \26470 );
and \U$20804 ( \26558 , \8412 , \26473 );
and \U$20805 ( \26559 , \8414 , \26475 );
and \U$20806 ( \26560 , \8416 , \26478 );
and \U$20807 ( \26561 , \8418 , \26480 );
and \U$20808 ( \26562 , \8420 , \26482 );
and \U$20809 ( \26563 , \8422 , \26484 );
and \U$20810 ( \26564 , \8424 , \26486 );
and \U$20811 ( \26565 , \8426 , \26488 );
or \U$20817 ( \26566 , \26555 , \26556 , \26557 , \26558 , \26559 , \26560 , \26561 , \26562 , \26563 , \26564 , \26565 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7ec0 ( \26567_nG7ec0 , \26566 , \26501 );
buf \U$20818 ( \26568 , \26567_nG7ec0 );
xor \U$20819 ( \26569 , \26554 , \26568 );
or \U$20820 ( \26570 , \26553 , \26569 );
buf \U$20821 ( \26571 , RIb7b9428_250);
and \U$20822 ( \26572 , \7156 , \26464 );
and \U$20823 ( \26573 , \7158 , \26467 );
and \U$20824 ( \26574 , \8446 , \26470 );
and \U$20825 ( \26575 , \8448 , \26473 );
and \U$20826 ( \26576 , \8450 , \26475 );
and \U$20827 ( \26577 , \8452 , \26478 );
and \U$20828 ( \26578 , \8454 , \26480 );
and \U$20829 ( \26579 , \8456 , \26482 );
and \U$20830 ( \26580 , \8458 , \26484 );
and \U$20831 ( \26581 , \8460 , \26486 );
and \U$20832 ( \26582 , \8462 , \26488 );
or \U$20838 ( \26583 , \26572 , \26573 , \26574 , \26575 , \26576 , \26577 , \26578 , \26579 , \26580 , \26581 , \26582 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7ed1 ( \26584_nG7ed1 , \26583 , \26501 );
buf \U$20839 ( \26585 , \26584_nG7ed1 );
xor \U$20840 ( \26586 , \26571 , \26585 );
or \U$20841 ( \26587 , \26570 , \26586 );
buf \U$20842 ( \26588 , RIb7b93b0_251);
and \U$20843 ( \26589 , \7166 , \26464 );
and \U$20844 ( \26590 , \7168 , \26467 );
and \U$20845 ( \26591 , \8482 , \26470 );
and \U$20846 ( \26592 , \8484 , \26473 );
and \U$20847 ( \26593 , \8486 , \26475 );
and \U$20848 ( \26594 , \8488 , \26478 );
and \U$20849 ( \26595 , \8490 , \26480 );
and \U$20850 ( \26596 , \8492 , \26482 );
and \U$20851 ( \26597 , \8494 , \26484 );
and \U$20852 ( \26598 , \8496 , \26486 );
and \U$20853 ( \26599 , \8498 , \26488 );
or \U$20859 ( \26600 , \26589 , \26590 , \26591 , \26592 , \26593 , \26594 , \26595 , \26596 , \26597 , \26598 , \26599 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7ee2 ( \26601_nG7ee2 , \26600 , \26501 );
buf \U$20860 ( \26602 , \26601_nG7ee2 );
xor \U$20861 ( \26603 , \26588 , \26602 );
or \U$20862 ( \26604 , \26587 , \26603 );
buf \U$20863 ( \26605 , RIb7af720_252);
and \U$20864 ( \26606 , \7176 , \26464 );
and \U$20865 ( \26607 , \7178 , \26467 );
and \U$20866 ( \26608 , \8518 , \26470 );
and \U$20867 ( \26609 , \8520 , \26473 );
and \U$20868 ( \26610 , \8522 , \26475 );
and \U$20869 ( \26611 , \8524 , \26478 );
and \U$20870 ( \26612 , \8526 , \26480 );
and \U$20871 ( \26613 , \8528 , \26482 );
and \U$20872 ( \26614 , \8530 , \26484 );
and \U$20873 ( \26615 , \8532 , \26486 );
and \U$20874 ( \26616 , \8534 , \26488 );
or \U$20880 ( \26617 , \26606 , \26607 , \26608 , \26609 , \26610 , \26611 , \26612 , \26613 , \26614 , \26615 , \26616 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7ef3 ( \26618_nG7ef3 , \26617 , \26501 );
buf \U$20881 ( \26619 , \26618_nG7ef3 );
xor \U$20882 ( \26620 , \26605 , \26619 );
or \U$20883 ( \26621 , \26604 , \26620 );
buf \U$20884 ( \26622 , RIb7af6a8_253);
and \U$20885 ( \26623 , \7186 , \26464 );
and \U$20886 ( \26624 , \7188 , \26467 );
and \U$20887 ( \26625 , \8554 , \26470 );
and \U$20888 ( \26626 , \8556 , \26473 );
and \U$20889 ( \26627 , \8558 , \26475 );
and \U$20890 ( \26628 , \8560 , \26478 );
and \U$20891 ( \26629 , \8562 , \26480 );
and \U$20892 ( \26630 , \8564 , \26482 );
and \U$20893 ( \26631 , \8566 , \26484 );
and \U$20894 ( \26632 , \8568 , \26486 );
and \U$20895 ( \26633 , \8570 , \26488 );
or \U$20901 ( \26634 , \26623 , \26624 , \26625 , \26626 , \26627 , \26628 , \26629 , \26630 , \26631 , \26632 , \26633 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7f04 ( \26635_nG7f04 , \26634 , \26501 );
buf \U$20902 ( \26636 , \26635_nG7f04 );
xor \U$20903 ( \26637 , \26622 , \26636 );
or \U$20904 ( \26638 , \26621 , \26637 );
not \U$20905 ( \26639 , \26638 );
buf \U$20906 ( \26640 , \26639 );
buf \U$20907 ( \26641 , RIb7af630_254);
and \U$20908 ( \26642 , \7198 , \26464 );
and \U$20909 ( \26643 , \7200 , \26467 );
and \U$20910 ( \26644 , \8645 , \26470 );
and \U$20911 ( \26645 , \8673 , \26473 );
and \U$20912 ( \26646 , \8701 , \26475 );
and \U$20913 ( \26647 , \8729 , \26478 );
and \U$20914 ( \26648 , \8757 , \26480 );
and \U$20915 ( \26649 , \8785 , \26482 );
and \U$20916 ( \26650 , \8813 , \26484 );
and \U$20917 ( \26651 , \8841 , \26486 );
and \U$20918 ( \26652 , \8869 , \26488 );
or \U$20924 ( \26653 , \26642 , \26643 , \26644 , \26645 , \26646 , \26647 , \26648 , \26649 , \26650 , \26651 , \26652 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7f17 ( \26654_nG7f17 , \26653 , \26501 );
buf \U$20925 ( \26655 , \26654_nG7f17 );
xor \U$20926 ( \26656 , \26641 , \26655 );
buf \U$20927 ( \26657 , RIb7af5b8_255);
and \U$20928 ( \26658 , \7207 , \26464 );
and \U$20929 ( \26659 , \7209 , \26467 );
and \U$20930 ( \26660 , \9119 , \26470 );
and \U$20931 ( \26661 , \9121 , \26473 );
and \U$20932 ( \26662 , \9123 , \26475 );
and \U$20933 ( \26663 , \9125 , \26478 );
and \U$20934 ( \26664 , \9127 , \26480 );
and \U$20935 ( \26665 , \9129 , \26482 );
and \U$20936 ( \26666 , \9131 , \26484 );
and \U$20937 ( \26667 , \9133 , \26486 );
and \U$20938 ( \26668 , \9135 , \26488 );
or \U$20944 ( \26669 , \26658 , \26659 , \26660 , \26661 , \26662 , \26663 , \26664 , \26665 , \26666 , \26667 , \26668 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7f27 ( \26670_nG7f27 , \26669 , \26501 );
buf \U$20945 ( \26671 , \26670_nG7f27 );
xor \U$20946 ( \26672 , \26657 , \26671 );
or \U$20947 ( \26673 , \26656 , \26672 );
buf \U$20948 ( \26674 , RIb7af540_256);
and \U$20949 ( \26675 , \7217 , \26464 );
and \U$20950 ( \26676 , \7219 , \26467 );
and \U$20951 ( \26677 , \9155 , \26470 );
and \U$20952 ( \26678 , \9157 , \26473 );
and \U$20953 ( \26679 , \9159 , \26475 );
and \U$20954 ( \26680 , \9161 , \26478 );
and \U$20955 ( \26681 , \9163 , \26480 );
and \U$20956 ( \26682 , \9165 , \26482 );
and \U$20957 ( \26683 , \9167 , \26484 );
and \U$20958 ( \26684 , \9169 , \26486 );
and \U$20959 ( \26685 , \9171 , \26488 );
or \U$20965 ( \26686 , \26675 , \26676 , \26677 , \26678 , \26679 , \26680 , \26681 , \26682 , \26683 , \26684 , \26685 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7f38 ( \26687_nG7f38 , \26686 , \26501 );
buf \U$20966 ( \26688 , \26687_nG7f38 );
xor \U$20967 ( \26689 , \26674 , \26688 );
or \U$20968 ( \26690 , \26673 , \26689 );
buf \U$20969 ( \26691 , RIb7af4c8_257);
and \U$20970 ( \26692 , \7227 , \26464 );
and \U$20971 ( \26693 , \7229 , \26467 );
and \U$20972 ( \26694 , \9191 , \26470 );
and \U$20973 ( \26695 , \9193 , \26473 );
and \U$20974 ( \26696 , \9195 , \26475 );
and \U$20975 ( \26697 , \9197 , \26478 );
and \U$20976 ( \26698 , \9199 , \26480 );
and \U$20977 ( \26699 , \9201 , \26482 );
and \U$20978 ( \26700 , \9203 , \26484 );
and \U$20979 ( \26701 , \9205 , \26486 );
and \U$20980 ( \26702 , \9207 , \26488 );
or \U$20986 ( \26703 , \26692 , \26693 , \26694 , \26695 , \26696 , \26697 , \26698 , \26699 , \26700 , \26701 , \26702 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7f49 ( \26704_nG7f49 , \26703 , \26501 );
buf \U$20987 ( \26705 , \26704_nG7f49 );
xor \U$20988 ( \26706 , \26691 , \26705 );
or \U$20989 ( \26707 , \26690 , \26706 );
buf \U$20990 ( \26708 , RIb7af450_258);
and \U$20991 ( \26709 , \7237 , \26464 );
and \U$20992 ( \26710 , \7239 , \26467 );
and \U$20993 ( \26711 , \9227 , \26470 );
and \U$20994 ( \26712 , \9229 , \26473 );
and \U$20995 ( \26713 , \9231 , \26475 );
and \U$20996 ( \26714 , \9233 , \26478 );
and \U$20997 ( \26715 , \9235 , \26480 );
and \U$20998 ( \26716 , \9237 , \26482 );
and \U$20999 ( \26717 , \9239 , \26484 );
and \U$21000 ( \26718 , \9241 , \26486 );
and \U$21001 ( \26719 , \9243 , \26488 );
or \U$21007 ( \26720 , \26709 , \26710 , \26711 , \26712 , \26713 , \26714 , \26715 , \26716 , \26717 , \26718 , \26719 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7f5a ( \26721_nG7f5a , \26720 , \26501 );
buf \U$21008 ( \26722 , \26721_nG7f5a );
xor \U$21009 ( \26723 , \26708 , \26722 );
or \U$21010 ( \26724 , \26707 , \26723 );
buf \U$21011 ( \26725 , RIb7af3d8_259);
and \U$21012 ( \26726 , \7247 , \26464 );
and \U$21013 ( \26727 , \7249 , \26467 );
and \U$21014 ( \26728 , \9263 , \26470 );
and \U$21015 ( \26729 , \9265 , \26473 );
and \U$21016 ( \26730 , \9267 , \26475 );
and \U$21017 ( \26731 , \9269 , \26478 );
and \U$21018 ( \26732 , \9271 , \26480 );
and \U$21019 ( \26733 , \9273 , \26482 );
and \U$21020 ( \26734 , \9275 , \26484 );
and \U$21021 ( \26735 , \9277 , \26486 );
and \U$21022 ( \26736 , \9279 , \26488 );
or \U$21028 ( \26737 , \26726 , \26727 , \26728 , \26729 , \26730 , \26731 , \26732 , \26733 , \26734 , \26735 , \26736 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7f6b ( \26738_nG7f6b , \26737 , \26501 );
buf \U$21029 ( \26739 , \26738_nG7f6b );
xor \U$21030 ( \26740 , \26725 , \26739 );
or \U$21031 ( \26741 , \26724 , \26740 );
buf \U$21032 ( \26742 , RIb7a5bf8_260);
and \U$21033 ( \26743 , \7257 , \26464 );
and \U$21034 ( \26744 , \7259 , \26467 );
and \U$21035 ( \26745 , \9299 , \26470 );
and \U$21036 ( \26746 , \9301 , \26473 );
and \U$21037 ( \26747 , \9303 , \26475 );
and \U$21038 ( \26748 , \9305 , \26478 );
and \U$21039 ( \26749 , \9307 , \26480 );
and \U$21040 ( \26750 , \9309 , \26482 );
and \U$21041 ( \26751 , \9311 , \26484 );
and \U$21042 ( \26752 , \9313 , \26486 );
and \U$21043 ( \26753 , \9315 , \26488 );
or \U$21049 ( \26754 , \26743 , \26744 , \26745 , \26746 , \26747 , \26748 , \26749 , \26750 , \26751 , \26752 , \26753 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7f7c ( \26755_nG7f7c , \26754 , \26501 );
buf \U$21050 ( \26756 , \26755_nG7f7c );
xor \U$21051 ( \26757 , \26742 , \26756 );
or \U$21052 ( \26758 , \26741 , \26757 );
buf \U$21053 ( \26759 , RIb7a0c48_261);
and \U$21054 ( \26760 , \7267 , \26464 );
and \U$21055 ( \26761 , \7269 , \26467 );
and \U$21056 ( \26762 , \9335 , \26470 );
and \U$21057 ( \26763 , \9337 , \26473 );
and \U$21058 ( \26764 , \9339 , \26475 );
and \U$21059 ( \26765 , \9341 , \26478 );
and \U$21060 ( \26766 , \9343 , \26480 );
and \U$21061 ( \26767 , \9345 , \26482 );
and \U$21062 ( \26768 , \9347 , \26484 );
and \U$21063 ( \26769 , \9349 , \26486 );
and \U$21064 ( \26770 , \9351 , \26488 );
or \U$21070 ( \26771 , \26760 , \26761 , \26762 , \26763 , \26764 , \26765 , \26766 , \26767 , \26768 , \26769 , \26770 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g7f8d ( \26772_nG7f8d , \26771 , \26501 );
buf \U$21071 ( \26773 , \26772_nG7f8d );
xor \U$21072 ( \26774 , \26759 , \26773 );
or \U$21073 ( \26775 , \26758 , \26774 );
not \U$21074 ( \26776 , \26775 );
buf \U$21075 ( \26777 , \26776 );
and \U$21076 ( \26778 , \26640 , \26777 );
and \U$21077 ( \26779 , \26503 , \26778 );
_HMUX g7f95 ( \26780_nG7f95 , \26444_nG7e44 , \26446 , \26779 );
buf \U$21080 ( \26781 , \26446 );
buf \U$21083 ( \26782 , \26449 );
buf \U$21086 ( \26783 , \26452 );
buf \U$21089 ( \26784 , \26456 );
buf \U$21090 ( \26785 , \26460 );
not \U$21091 ( \26786 , \26785 );
buf \U$21092 ( \26787 , \26786 );
not \U$21093 ( \26788 , \26787 );
buf \U$21094 ( \26789 , \26463 );
xnor \U$21095 ( \26790 , \26789 , \26785 );
buf \U$21096 ( \26791 , \26790 );
or \U$21097 ( \26792 , \26789 , \26785 );
not \U$21098 ( \26793 , \26792 );
buf \U$21099 ( \26794 , \26793 );
buf \U$21100 ( \26795 , \26794 );
buf \U$21101 ( \26796 , \26794 );
buf \U$21102 ( \26797 , \26794 );
buf \U$21103 ( \26798 , \26794 );
buf \U$21104 ( \26799 , \26794 );
buf \U$21105 ( \26800 , \26794 );
buf \U$21106 ( \26801 , \26794 );
buf \U$21107 ( \26802 , \26794 );
buf \U$21108 ( \26803 , \26794 );
buf \U$21109 ( \26804 , \26794 );
buf \U$21110 ( \26805 , \26794 );
buf \U$21111 ( \26806 , \26794 );
buf \U$21112 ( \26807 , \26794 );
buf \U$21113 ( \26808 , \26794 );
buf \U$21114 ( \26809 , \26794 );
buf \U$21115 ( \26810 , \26794 );
buf \U$21116 ( \26811 , \26794 );
buf \U$21117 ( \26812 , \26794 );
buf \U$21118 ( \26813 , \26794 );
buf \U$21119 ( \26814 , \26794 );
buf \U$21120 ( \26815 , \26794 );
buf \U$21121 ( \26816 , \26794 );
buf \U$21122 ( \26817 , \26794 );
buf \U$21123 ( \26818 , \26794 );
buf \U$21124 ( \26819 , \26794 );
nor \U$21125 ( \26820 , \26781 , \26782 , \26783 , \26784 , \26788 , \26791 , \26794 , \26795 , \26796 , \26797 , \26798 , \26799 , \26800 , \26801 , \26802 , \26803 , \26804 , \26805 , \26806 , \26807 , \26808 , \26809 , \26810 , \26811 , \26812 , \26813 , \26814 , \26815 , \26816 , \26817 , \26818 , \26819 );
and \U$21126 ( \26821 , RIe5329d0_6883, \26820 );
not \U$21127 ( \26822 , \26781 );
not \U$21128 ( \26823 , \26782 );
not \U$21129 ( \26824 , \26783 );
not \U$21130 ( \26825 , \26784 );
buf \U$21131 ( \26826 , \26794 );
buf \U$21132 ( \26827 , \26794 );
buf \U$21133 ( \26828 , \26794 );
buf \U$21134 ( \26829 , \26794 );
buf \U$21135 ( \26830 , \26794 );
buf \U$21136 ( \26831 , \26794 );
buf \U$21137 ( \26832 , \26794 );
buf \U$21138 ( \26833 , \26794 );
buf \U$21139 ( \26834 , \26794 );
buf \U$21140 ( \26835 , \26794 );
buf \U$21141 ( \26836 , \26794 );
buf \U$21142 ( \26837 , \26794 );
buf \U$21143 ( \26838 , \26794 );
buf \U$21144 ( \26839 , \26794 );
buf \U$21145 ( \26840 , \26794 );
buf \U$21146 ( \26841 , \26794 );
buf \U$21147 ( \26842 , \26794 );
buf \U$21148 ( \26843 , \26794 );
buf \U$21149 ( \26844 , \26794 );
buf \U$21150 ( \26845 , \26794 );
buf \U$21151 ( \26846 , \26794 );
buf \U$21152 ( \26847 , \26794 );
buf \U$21153 ( \26848 , \26794 );
buf \U$21154 ( \26849 , \26794 );
buf \U$21155 ( \26850 , \26794 );
nor \U$21156 ( \26851 , \26822 , \26823 , \26824 , \26825 , \26787 , \26791 , \26794 , \26826 , \26827 , \26828 , \26829 , \26830 , \26831 , \26832 , \26833 , \26834 , \26835 , \26836 , \26837 , \26838 , \26839 , \26840 , \26841 , \26842 , \26843 , \26844 , \26845 , \26846 , \26847 , \26848 , \26849 , \26850 );
and \U$21157 ( \26852 , RIeb72150_6905, \26851 );
buf \U$21158 ( \26853 , \26794 );
buf \U$21159 ( \26854 , \26794 );
buf \U$21160 ( \26855 , \26794 );
buf \U$21161 ( \26856 , \26794 );
buf \U$21162 ( \26857 , \26794 );
buf \U$21163 ( \26858 , \26794 );
buf \U$21164 ( \26859 , \26794 );
buf \U$21165 ( \26860 , \26794 );
buf \U$21166 ( \26861 , \26794 );
buf \U$21167 ( \26862 , \26794 );
buf \U$21168 ( \26863 , \26794 );
buf \U$21169 ( \26864 , \26794 );
buf \U$21170 ( \26865 , \26794 );
buf \U$21171 ( \26866 , \26794 );
buf \U$21172 ( \26867 , \26794 );
buf \U$21173 ( \26868 , \26794 );
buf \U$21174 ( \26869 , \26794 );
buf \U$21175 ( \26870 , \26794 );
buf \U$21176 ( \26871 , \26794 );
buf \U$21177 ( \26872 , \26794 );
buf \U$21178 ( \26873 , \26794 );
buf \U$21179 ( \26874 , \26794 );
buf \U$21180 ( \26875 , \26794 );
buf \U$21181 ( \26876 , \26794 );
buf \U$21182 ( \26877 , \26794 );
nor \U$21183 ( \26878 , \26781 , \26823 , \26824 , \26825 , \26787 , \26791 , \26794 , \26853 , \26854 , \26855 , \26856 , \26857 , \26858 , \26859 , \26860 , \26861 , \26862 , \26863 , \26864 , \26865 , \26866 , \26867 , \26868 , \26869 , \26870 , \26871 , \26872 , \26873 , \26874 , \26875 , \26876 , \26877 );
and \U$21184 ( \26879 , RIeab80c0_6897, \26878 );
buf \U$21185 ( \26880 , \26794 );
buf \U$21186 ( \26881 , \26794 );
buf \U$21187 ( \26882 , \26794 );
buf \U$21188 ( \26883 , \26794 );
buf \U$21189 ( \26884 , \26794 );
buf \U$21190 ( \26885 , \26794 );
buf \U$21191 ( \26886 , \26794 );
buf \U$21192 ( \26887 , \26794 );
buf \U$21193 ( \26888 , \26794 );
buf \U$21194 ( \26889 , \26794 );
buf \U$21195 ( \26890 , \26794 );
buf \U$21196 ( \26891 , \26794 );
buf \U$21197 ( \26892 , \26794 );
buf \U$21198 ( \26893 , \26794 );
buf \U$21199 ( \26894 , \26794 );
buf \U$21200 ( \26895 , \26794 );
buf \U$21201 ( \26896 , \26794 );
buf \U$21202 ( \26897 , \26794 );
buf \U$21203 ( \26898 , \26794 );
buf \U$21204 ( \26899 , \26794 );
buf \U$21205 ( \26900 , \26794 );
buf \U$21206 ( \26901 , \26794 );
buf \U$21207 ( \26902 , \26794 );
buf \U$21208 ( \26903 , \26794 );
buf \U$21209 ( \26904 , \26794 );
nor \U$21210 ( \26905 , \26822 , \26782 , \26824 , \26825 , \26787 , \26791 , \26794 , \26880 , \26881 , \26882 , \26883 , \26884 , \26885 , \26886 , \26887 , \26888 , \26889 , \26890 , \26891 , \26892 , \26893 , \26894 , \26895 , \26896 , \26897 , \26898 , \26899 , \26900 , \26901 , \26902 , \26903 , \26904 );
and \U$21211 ( \26906 , RIe5331c8_6882, \26905 );
buf \U$21212 ( \26907 , \26794 );
buf \U$21213 ( \26908 , \26794 );
buf \U$21214 ( \26909 , \26794 );
buf \U$21215 ( \26910 , \26794 );
buf \U$21216 ( \26911 , \26794 );
buf \U$21217 ( \26912 , \26794 );
buf \U$21218 ( \26913 , \26794 );
buf \U$21219 ( \26914 , \26794 );
buf \U$21220 ( \26915 , \26794 );
buf \U$21221 ( \26916 , \26794 );
buf \U$21222 ( \26917 , \26794 );
buf \U$21223 ( \26918 , \26794 );
buf \U$21224 ( \26919 , \26794 );
buf \U$21225 ( \26920 , \26794 );
buf \U$21226 ( \26921 , \26794 );
buf \U$21227 ( \26922 , \26794 );
buf \U$21228 ( \26923 , \26794 );
buf \U$21229 ( \26924 , \26794 );
buf \U$21230 ( \26925 , \26794 );
buf \U$21231 ( \26926 , \26794 );
buf \U$21232 ( \26927 , \26794 );
buf \U$21233 ( \26928 , \26794 );
buf \U$21234 ( \26929 , \26794 );
buf \U$21235 ( \26930 , \26794 );
buf \U$21236 ( \26931 , \26794 );
nor \U$21237 ( \26932 , \26781 , \26782 , \26824 , \26825 , \26787 , \26791 , \26794 , \26907 , \26908 , \26909 , \26910 , \26911 , \26912 , \26913 , \26914 , \26915 , \26916 , \26917 , \26918 , \26919 , \26920 , \26921 , \26922 , \26923 , \26924 , \26925 , \26926 , \26927 , \26928 , \26929 , \26930 , \26931 );
and \U$21238 ( \26933 , RIe5339c0_6881, \26932 );
buf \U$21239 ( \26934 , \26794 );
buf \U$21240 ( \26935 , \26794 );
buf \U$21241 ( \26936 , \26794 );
buf \U$21242 ( \26937 , \26794 );
buf \U$21243 ( \26938 , \26794 );
buf \U$21244 ( \26939 , \26794 );
buf \U$21245 ( \26940 , \26794 );
buf \U$21246 ( \26941 , \26794 );
buf \U$21247 ( \26942 , \26794 );
buf \U$21248 ( \26943 , \26794 );
buf \U$21249 ( \26944 , \26794 );
buf \U$21250 ( \26945 , \26794 );
buf \U$21251 ( \26946 , \26794 );
buf \U$21252 ( \26947 , \26794 );
buf \U$21253 ( \26948 , \26794 );
buf \U$21254 ( \26949 , \26794 );
buf \U$21255 ( \26950 , \26794 );
buf \U$21256 ( \26951 , \26794 );
buf \U$21257 ( \26952 , \26794 );
buf \U$21258 ( \26953 , \26794 );
buf \U$21259 ( \26954 , \26794 );
buf \U$21260 ( \26955 , \26794 );
buf \U$21261 ( \26956 , \26794 );
buf \U$21262 ( \26957 , \26794 );
buf \U$21263 ( \26958 , \26794 );
nor \U$21264 ( \26959 , \26822 , \26823 , \26783 , \26825 , \26787 , \26791 , \26794 , \26934 , \26935 , \26936 , \26937 , \26938 , \26939 , \26940 , \26941 , \26942 , \26943 , \26944 , \26945 , \26946 , \26947 , \26948 , \26949 , \26950 , \26951 , \26952 , \26953 , \26954 , \26955 , \26956 , \26957 , \26958 );
and \U$21265 ( \26960 , RIeab87c8_6898, \26959 );
buf \U$21266 ( \26961 , \26794 );
buf \U$21267 ( \26962 , \26794 );
buf \U$21268 ( \26963 , \26794 );
buf \U$21269 ( \26964 , \26794 );
buf \U$21270 ( \26965 , \26794 );
buf \U$21271 ( \26966 , \26794 );
buf \U$21272 ( \26967 , \26794 );
buf \U$21273 ( \26968 , \26794 );
buf \U$21274 ( \26969 , \26794 );
buf \U$21275 ( \26970 , \26794 );
buf \U$21276 ( \26971 , \26794 );
buf \U$21277 ( \26972 , \26794 );
buf \U$21278 ( \26973 , \26794 );
buf \U$21279 ( \26974 , \26794 );
buf \U$21280 ( \26975 , \26794 );
buf \U$21281 ( \26976 , \26794 );
buf \U$21282 ( \26977 , \26794 );
buf \U$21283 ( \26978 , \26794 );
buf \U$21284 ( \26979 , \26794 );
buf \U$21285 ( \26980 , \26794 );
buf \U$21286 ( \26981 , \26794 );
buf \U$21287 ( \26982 , \26794 );
buf \U$21288 ( \26983 , \26794 );
buf \U$21289 ( \26984 , \26794 );
buf \U$21290 ( \26985 , \26794 );
nor \U$21291 ( \26986 , \26781 , \26823 , \26783 , \26825 , \26787 , \26791 , \26794 , \26961 , \26962 , \26963 , \26964 , \26965 , \26966 , \26967 , \26968 , \26969 , \26970 , \26971 , \26972 , \26973 , \26974 , \26975 , \26976 , \26977 , \26978 , \26979 , \26980 , \26981 , \26982 , \26983 , \26984 , \26985 );
and \U$21292 ( \26987 , RIe5341b8_6880, \26986 );
buf \U$21293 ( \26988 , \26794 );
buf \U$21294 ( \26989 , \26794 );
buf \U$21295 ( \26990 , \26794 );
buf \U$21296 ( \26991 , \26794 );
buf \U$21297 ( \26992 , \26794 );
buf \U$21298 ( \26993 , \26794 );
buf \U$21299 ( \26994 , \26794 );
buf \U$21300 ( \26995 , \26794 );
buf \U$21301 ( \26996 , \26794 );
buf \U$21302 ( \26997 , \26794 );
buf \U$21303 ( \26998 , \26794 );
buf \U$21304 ( \26999 , \26794 );
buf \U$21305 ( \27000 , \26794 );
buf \U$21306 ( \27001 , \26794 );
buf \U$21307 ( \27002 , \26794 );
buf \U$21308 ( \27003 , \26794 );
buf \U$21309 ( \27004 , \26794 );
buf \U$21310 ( \27005 , \26794 );
buf \U$21311 ( \27006 , \26794 );
buf \U$21312 ( \27007 , \26794 );
buf \U$21313 ( \27008 , \26794 );
buf \U$21314 ( \27009 , \26794 );
buf \U$21315 ( \27010 , \26794 );
buf \U$21316 ( \27011 , \26794 );
buf \U$21317 ( \27012 , \26794 );
nor \U$21318 ( \27013 , \26822 , \26782 , \26783 , \26825 , \26787 , \26791 , \26794 , \26988 , \26989 , \26990 , \26991 , \26992 , \26993 , \26994 , \26995 , \26996 , \26997 , \26998 , \26999 , \27000 , \27001 , \27002 , \27003 , \27004 , \27005 , \27006 , \27007 , \27008 , \27009 , \27010 , \27011 , \27012 );
and \U$21319 ( \27014 , RIe5349b0_6879, \27013 );
buf \U$21320 ( \27015 , \26794 );
buf \U$21321 ( \27016 , \26794 );
buf \U$21322 ( \27017 , \26794 );
buf \U$21323 ( \27018 , \26794 );
buf \U$21324 ( \27019 , \26794 );
buf \U$21325 ( \27020 , \26794 );
buf \U$21326 ( \27021 , \26794 );
buf \U$21327 ( \27022 , \26794 );
buf \U$21328 ( \27023 , \26794 );
buf \U$21329 ( \27024 , \26794 );
buf \U$21330 ( \27025 , \26794 );
buf \U$21331 ( \27026 , \26794 );
buf \U$21332 ( \27027 , \26794 );
buf \U$21333 ( \27028 , \26794 );
buf \U$21334 ( \27029 , \26794 );
buf \U$21335 ( \27030 , \26794 );
buf \U$21336 ( \27031 , \26794 );
buf \U$21337 ( \27032 , \26794 );
buf \U$21338 ( \27033 , \26794 );
buf \U$21339 ( \27034 , \26794 );
buf \U$21340 ( \27035 , \26794 );
buf \U$21341 ( \27036 , \26794 );
buf \U$21342 ( \27037 , \26794 );
buf \U$21343 ( \27038 , \26794 );
buf \U$21344 ( \27039 , \26794 );
nor \U$21345 ( \27040 , \26781 , \26782 , \26783 , \26825 , \26787 , \26791 , \26794 , \27015 , \27016 , \27017 , \27018 , \27019 , \27020 , \27021 , \27022 , \27023 , \27024 , \27025 , \27026 , \27027 , \27028 , \27029 , \27030 , \27031 , \27032 , \27033 , \27034 , \27035 , \27036 , \27037 , \27038 , \27039 );
and \U$21346 ( \27041 , RIea94af8_6890, \27040 );
buf \U$21347 ( \27042 , \26794 );
buf \U$21348 ( \27043 , \26794 );
buf \U$21349 ( \27044 , \26794 );
buf \U$21350 ( \27045 , \26794 );
buf \U$21351 ( \27046 , \26794 );
buf \U$21352 ( \27047 , \26794 );
buf \U$21353 ( \27048 , \26794 );
buf \U$21354 ( \27049 , \26794 );
buf \U$21355 ( \27050 , \26794 );
buf \U$21356 ( \27051 , \26794 );
buf \U$21357 ( \27052 , \26794 );
buf \U$21358 ( \27053 , \26794 );
buf \U$21359 ( \27054 , \26794 );
buf \U$21360 ( \27055 , \26794 );
buf \U$21361 ( \27056 , \26794 );
buf \U$21362 ( \27057 , \26794 );
buf \U$21363 ( \27058 , \26794 );
buf \U$21364 ( \27059 , \26794 );
buf \U$21365 ( \27060 , \26794 );
buf \U$21366 ( \27061 , \26794 );
buf \U$21367 ( \27062 , \26794 );
buf \U$21368 ( \27063 , \26794 );
buf \U$21369 ( \27064 , \26794 );
buf \U$21370 ( \27065 , \26794 );
buf \U$21371 ( \27066 , \26794 );
nor \U$21372 ( \27067 , \26822 , \26823 , \26824 , \26784 , \26787 , \26791 , \26794 , \27042 , \27043 , \27044 , \27045 , \27046 , \27047 , \27048 , \27049 , \27050 , \27051 , \27052 , \27053 , \27054 , \27055 , \27056 , \27057 , \27058 , \27059 , \27060 , \27061 , \27062 , \27063 , \27064 , \27065 , \27066 );
and \U$21373 ( \27068 , RIe5351a8_6878, \27067 );
buf \U$21374 ( \27069 , \26794 );
buf \U$21375 ( \27070 , \26794 );
buf \U$21376 ( \27071 , \26794 );
buf \U$21377 ( \27072 , \26794 );
buf \U$21378 ( \27073 , \26794 );
buf \U$21379 ( \27074 , \26794 );
buf \U$21380 ( \27075 , \26794 );
buf \U$21381 ( \27076 , \26794 );
buf \U$21382 ( \27077 , \26794 );
buf \U$21383 ( \27078 , \26794 );
buf \U$21384 ( \27079 , \26794 );
buf \U$21385 ( \27080 , \26794 );
buf \U$21386 ( \27081 , \26794 );
buf \U$21387 ( \27082 , \26794 );
buf \U$21388 ( \27083 , \26794 );
buf \U$21389 ( \27084 , \26794 );
buf \U$21390 ( \27085 , \26794 );
buf \U$21391 ( \27086 , \26794 );
buf \U$21392 ( \27087 , \26794 );
buf \U$21393 ( \27088 , \26794 );
buf \U$21394 ( \27089 , \26794 );
buf \U$21395 ( \27090 , \26794 );
buf \U$21396 ( \27091 , \26794 );
buf \U$21397 ( \27092 , \26794 );
buf \U$21398 ( \27093 , \26794 );
nor \U$21399 ( \27094 , \26781 , \26823 , \26824 , \26784 , \26787 , \26791 , \26794 , \27069 , \27070 , \27071 , \27072 , \27073 , \27074 , \27075 , \27076 , \27077 , \27078 , \27079 , \27080 , \27081 , \27082 , \27083 , \27084 , \27085 , \27086 , \27087 , \27088 , \27089 , \27090 , \27091 , \27092 , \27093 );
and \U$21400 ( \27095 , RIe5359a0_6877, \27094 );
buf \U$21401 ( \27096 , \26794 );
buf \U$21402 ( \27097 , \26794 );
buf \U$21403 ( \27098 , \26794 );
buf \U$21404 ( \27099 , \26794 );
buf \U$21405 ( \27100 , \26794 );
buf \U$21406 ( \27101 , \26794 );
buf \U$21407 ( \27102 , \26794 );
buf \U$21408 ( \27103 , \26794 );
buf \U$21409 ( \27104 , \26794 );
buf \U$21410 ( \27105 , \26794 );
buf \U$21411 ( \27106 , \26794 );
buf \U$21412 ( \27107 , \26794 );
buf \U$21413 ( \27108 , \26794 );
buf \U$21414 ( \27109 , \26794 );
buf \U$21415 ( \27110 , \26794 );
buf \U$21416 ( \27111 , \26794 );
buf \U$21417 ( \27112 , \26794 );
buf \U$21418 ( \27113 , \26794 );
buf \U$21419 ( \27114 , \26794 );
buf \U$21420 ( \27115 , \26794 );
buf \U$21421 ( \27116 , \26794 );
buf \U$21422 ( \27117 , \26794 );
buf \U$21423 ( \27118 , \26794 );
buf \U$21424 ( \27119 , \26794 );
buf \U$21425 ( \27120 , \26794 );
nor \U$21426 ( \27121 , \26822 , \26782 , \26824 , \26784 , \26787 , \26791 , \26794 , \27096 , \27097 , \27098 , \27099 , \27100 , \27101 , \27102 , \27103 , \27104 , \27105 , \27106 , \27107 , \27108 , \27109 , \27110 , \27111 , \27112 , \27113 , \27114 , \27115 , \27116 , \27117 , \27118 , \27119 , \27120 );
and \U$21427 ( \27122 , RIeab78c8_6895, \27121 );
buf \U$21428 ( \27123 , \26794 );
buf \U$21429 ( \27124 , \26794 );
buf \U$21430 ( \27125 , \26794 );
buf \U$21431 ( \27126 , \26794 );
buf \U$21432 ( \27127 , \26794 );
buf \U$21433 ( \27128 , \26794 );
buf \U$21434 ( \27129 , \26794 );
buf \U$21435 ( \27130 , \26794 );
buf \U$21436 ( \27131 , \26794 );
buf \U$21437 ( \27132 , \26794 );
buf \U$21438 ( \27133 , \26794 );
buf \U$21439 ( \27134 , \26794 );
buf \U$21440 ( \27135 , \26794 );
buf \U$21441 ( \27136 , \26794 );
buf \U$21442 ( \27137 , \26794 );
buf \U$21443 ( \27138 , \26794 );
buf \U$21444 ( \27139 , \26794 );
buf \U$21445 ( \27140 , \26794 );
buf \U$21446 ( \27141 , \26794 );
buf \U$21447 ( \27142 , \26794 );
buf \U$21448 ( \27143 , \26794 );
buf \U$21449 ( \27144 , \26794 );
buf \U$21450 ( \27145 , \26794 );
buf \U$21451 ( \27146 , \26794 );
buf \U$21452 ( \27147 , \26794 );
nor \U$21453 ( \27148 , \26781 , \26782 , \26824 , \26784 , \26787 , \26791 , \26794 , \27123 , \27124 , \27125 , \27126 , \27127 , \27128 , \27129 , \27130 , \27131 , \27132 , \27133 , \27134 , \27135 , \27136 , \27137 , \27138 , \27139 , \27140 , \27141 , \27142 , \27143 , \27144 , \27145 , \27146 , \27147 );
and \U$21454 ( \27149 , RIeab7d00_6896, \27148 );
buf \U$21455 ( \27150 , \26794 );
buf \U$21456 ( \27151 , \26794 );
buf \U$21457 ( \27152 , \26794 );
buf \U$21458 ( \27153 , \26794 );
buf \U$21459 ( \27154 , \26794 );
buf \U$21460 ( \27155 , \26794 );
buf \U$21461 ( \27156 , \26794 );
buf \U$21462 ( \27157 , \26794 );
buf \U$21463 ( \27158 , \26794 );
buf \U$21464 ( \27159 , \26794 );
buf \U$21465 ( \27160 , \26794 );
buf \U$21466 ( \27161 , \26794 );
buf \U$21467 ( \27162 , \26794 );
buf \U$21468 ( \27163 , \26794 );
buf \U$21469 ( \27164 , \26794 );
buf \U$21470 ( \27165 , \26794 );
buf \U$21471 ( \27166 , \26794 );
buf \U$21472 ( \27167 , \26794 );
buf \U$21473 ( \27168 , \26794 );
buf \U$21474 ( \27169 , \26794 );
buf \U$21475 ( \27170 , \26794 );
buf \U$21476 ( \27171 , \26794 );
buf \U$21477 ( \27172 , \26794 );
buf \U$21478 ( \27173 , \26794 );
buf \U$21479 ( \27174 , \26794 );
nor \U$21480 ( \27175 , \26822 , \26823 , \26783 , \26784 , \26787 , \26791 , \26794 , \27150 , \27151 , \27152 , \27153 , \27154 , \27155 , \27156 , \27157 , \27158 , \27159 , \27160 , \27161 , \27162 , \27163 , \27164 , \27165 , \27166 , \27167 , \27168 , \27169 , \27170 , \27171 , \27172 , \27173 , \27174 );
and \U$21481 ( \27176 , RIeacfa18_6902, \27175 );
buf \U$21482 ( \27177 , \26794 );
buf \U$21483 ( \27178 , \26794 );
buf \U$21484 ( \27179 , \26794 );
buf \U$21485 ( \27180 , \26794 );
buf \U$21486 ( \27181 , \26794 );
buf \U$21487 ( \27182 , \26794 );
buf \U$21488 ( \27183 , \26794 );
buf \U$21489 ( \27184 , \26794 );
buf \U$21490 ( \27185 , \26794 );
buf \U$21491 ( \27186 , \26794 );
buf \U$21492 ( \27187 , \26794 );
buf \U$21493 ( \27188 , \26794 );
buf \U$21494 ( \27189 , \26794 );
buf \U$21495 ( \27190 , \26794 );
buf \U$21496 ( \27191 , \26794 );
buf \U$21497 ( \27192 , \26794 );
buf \U$21498 ( \27193 , \26794 );
buf \U$21499 ( \27194 , \26794 );
buf \U$21500 ( \27195 , \26794 );
buf \U$21501 ( \27196 , \26794 );
buf \U$21502 ( \27197 , \26794 );
buf \U$21503 ( \27198 , \26794 );
buf \U$21504 ( \27199 , \26794 );
buf \U$21505 ( \27200 , \26794 );
buf \U$21506 ( \27201 , \26794 );
nor \U$21507 ( \27202 , \26781 , \26823 , \26783 , \26784 , \26787 , \26791 , \26794 , \27177 , \27178 , \27179 , \27180 , \27181 , \27182 , \27183 , \27184 , \27185 , \27186 , \27187 , \27188 , \27189 , \27190 , \27191 , \27192 , \27193 , \27194 , \27195 , \27196 , \27197 , \27198 , \27199 , \27200 , \27201 );
and \U$21508 ( \27203 , RIeab6518_6891, \27202 );
buf \U$21509 ( \27204 , \26794 );
buf \U$21510 ( \27205 , \26794 );
buf \U$21511 ( \27206 , \26794 );
buf \U$21512 ( \27207 , \26794 );
buf \U$21513 ( \27208 , \26794 );
buf \U$21514 ( \27209 , \26794 );
buf \U$21515 ( \27210 , \26794 );
buf \U$21516 ( \27211 , \26794 );
buf \U$21517 ( \27212 , \26794 );
buf \U$21518 ( \27213 , \26794 );
buf \U$21519 ( \27214 , \26794 );
buf \U$21520 ( \27215 , \26794 );
buf \U$21521 ( \27216 , \26794 );
buf \U$21522 ( \27217 , \26794 );
buf \U$21523 ( \27218 , \26794 );
buf \U$21524 ( \27219 , \26794 );
buf \U$21525 ( \27220 , \26794 );
buf \U$21526 ( \27221 , \26794 );
buf \U$21527 ( \27222 , \26794 );
buf \U$21528 ( \27223 , \26794 );
buf \U$21529 ( \27224 , \26794 );
buf \U$21530 ( \27225 , \26794 );
buf \U$21531 ( \27226 , \26794 );
buf \U$21532 ( \27227 , \26794 );
buf \U$21533 ( \27228 , \26794 );
nor \U$21534 ( \27229 , \26822 , \26782 , \26783 , \26784 , \26787 , \26791 , \26794 , \27204 , \27205 , \27206 , \27207 , \27208 , \27209 , \27210 , \27211 , \27212 , \27213 , \27214 , \27215 , \27216 , \27217 , \27218 , \27219 , \27220 , \27221 , \27222 , \27223 , \27224 , \27225 , \27226 , \27227 , \27228 );
and \U$21535 ( \27230 , RIeb352c8_6904, \27229 );
or \U$21536 ( \27231 , \26821 , \26852 , \26879 , \26906 , \26933 , \26960 , \26987 , \27014 , \27041 , \27068 , \27095 , \27122 , \27149 , \27176 , \27203 , \27230 );
buf \U$21537 ( \27232 , \26794 );
not \U$21538 ( \27233 , \27232 );
buf \U$21539 ( \27234 , \26782 );
buf \U$21540 ( \27235 , \26783 );
buf \U$21541 ( \27236 , \26784 );
buf \U$21542 ( \27237 , \26787 );
buf \U$21543 ( \27238 , \26791 );
buf \U$21544 ( \27239 , \26794 );
buf \U$21545 ( \27240 , \26794 );
buf \U$21546 ( \27241 , \26794 );
buf \U$21547 ( \27242 , \26794 );
buf \U$21548 ( \27243 , \26794 );
buf \U$21549 ( \27244 , \26794 );
buf \U$21550 ( \27245 , \26794 );
buf \U$21551 ( \27246 , \26794 );
buf \U$21552 ( \27247 , \26794 );
buf \U$21553 ( \27248 , \26794 );
buf \U$21554 ( \27249 , \26794 );
buf \U$21555 ( \27250 , \26794 );
buf \U$21556 ( \27251 , \26794 );
buf \U$21557 ( \27252 , \26794 );
buf \U$21558 ( \27253 , \26794 );
buf \U$21559 ( \27254 , \26794 );
buf \U$21560 ( \27255 , \26794 );
buf \U$21561 ( \27256 , \26794 );
buf \U$21562 ( \27257 , \26794 );
buf \U$21563 ( \27258 , \26794 );
buf \U$21564 ( \27259 , \26794 );
buf \U$21565 ( \27260 , \26794 );
buf \U$21566 ( \27261 , \26794 );
buf \U$21567 ( \27262 , \26794 );
buf \U$21568 ( \27263 , \26794 );
buf \U$21569 ( \27264 , \26781 );
or \U$21570 ( \27265 , \27234 , \27235 , \27236 , \27237 , \27238 , \27239 , \27240 , \27241 , \27242 , \27243 , \27244 , \27245 , \27246 , \27247 , \27248 , \27249 , \27250 , \27251 , \27252 , \27253 , \27254 , \27255 , \27256 , \27257 , \27258 , \27259 , \27260 , \27261 , \27262 , \27263 , \27264 );
nand \U$21571 ( \27266 , \27233 , \27265 );
buf \U$21572 ( \27267 , \27266 );
buf \U$21573 ( \27268 , \26794 );
not \U$21574 ( \27269 , \27268 );
buf \U$21575 ( \27270 , \26791 );
buf \U$21576 ( \27271 , \26794 );
buf \U$21577 ( \27272 , \26794 );
buf \U$21578 ( \27273 , \26794 );
buf \U$21579 ( \27274 , \26794 );
buf \U$21580 ( \27275 , \26794 );
buf \U$21581 ( \27276 , \26794 );
buf \U$21582 ( \27277 , \26794 );
buf \U$21583 ( \27278 , \26794 );
buf \U$21584 ( \27279 , \26794 );
buf \U$21585 ( \27280 , \26794 );
buf \U$21586 ( \27281 , \26794 );
buf \U$21587 ( \27282 , \26794 );
buf \U$21588 ( \27283 , \26794 );
buf \U$21589 ( \27284 , \26794 );
buf \U$21590 ( \27285 , \26794 );
buf \U$21591 ( \27286 , \26794 );
buf \U$21592 ( \27287 , \26794 );
buf \U$21593 ( \27288 , \26794 );
buf \U$21594 ( \27289 , \26794 );
buf \U$21595 ( \27290 , \26794 );
buf \U$21596 ( \27291 , \26794 );
buf \U$21597 ( \27292 , \26794 );
buf \U$21598 ( \27293 , \26794 );
buf \U$21599 ( \27294 , \26794 );
buf \U$21600 ( \27295 , \26794 );
buf \U$21601 ( \27296 , \26787 );
buf \U$21602 ( \27297 , \26781 );
buf \U$21603 ( \27298 , \26782 );
buf \U$21604 ( \27299 , \26783 );
buf \U$21605 ( \27300 , \26784 );
or \U$21606 ( \27301 , \27297 , \27298 , \27299 , \27300 );
and \U$21607 ( \27302 , \27296 , \27301 );
or \U$21608 ( \27303 , \27270 , \27271 , \27272 , \27273 , \27274 , \27275 , \27276 , \27277 , \27278 , \27279 , \27280 , \27281 , \27282 , \27283 , \27284 , \27285 , \27286 , \27287 , \27288 , \27289 , \27290 , \27291 , \27292 , \27293 , \27294 , \27295 , \27302 );
and \U$21609 ( \27304 , \27269 , \27303 );
buf \U$21610 ( \27305 , \27304 );
or \U$21611 ( \27306 , \27267 , \27305 );
_DC g81ac ( \27307_nG81ac , \27231 , \27306 );
not \U$21612 ( \27308 , \27307_nG81ac );
buf \U$21613 ( \27309 , RIb7b9608_246);
buf \U$21614 ( \27310 , \26794 );
buf \U$21615 ( \27311 , \26794 );
buf \U$21616 ( \27312 , \26794 );
buf \U$21617 ( \27313 , \26794 );
buf \U$21618 ( \27314 , \26794 );
buf \U$21619 ( \27315 , \26794 );
buf \U$21620 ( \27316 , \26794 );
buf \U$21621 ( \27317 , \26794 );
buf \U$21622 ( \27318 , \26794 );
buf \U$21623 ( \27319 , \26794 );
buf \U$21624 ( \27320 , \26794 );
buf \U$21625 ( \27321 , \26794 );
buf \U$21626 ( \27322 , \26794 );
buf \U$21627 ( \27323 , \26794 );
buf \U$21628 ( \27324 , \26794 );
buf \U$21629 ( \27325 , \26794 );
buf \U$21630 ( \27326 , \26794 );
buf \U$21631 ( \27327 , \26794 );
buf \U$21632 ( \27328 , \26794 );
buf \U$21633 ( \27329 , \26794 );
buf \U$21634 ( \27330 , \26794 );
buf \U$21635 ( \27331 , \26794 );
buf \U$21636 ( \27332 , \26794 );
buf \U$21637 ( \27333 , \26794 );
buf \U$21638 ( \27334 , \26794 );
nor \U$21639 ( \27335 , \26781 , \26782 , \26783 , \26784 , \26788 , \26791 , \26794 , \27310 , \27311 , \27312 , \27313 , \27314 , \27315 , \27316 , \27317 , \27318 , \27319 , \27320 , \27321 , \27322 , \27323 , \27324 , \27325 , \27326 , \27327 , \27328 , \27329 , \27330 , \27331 , \27332 , \27333 , \27334 );
and \U$21640 ( \27336 , \7117 , \27335 );
buf \U$21641 ( \27337 , \26794 );
buf \U$21642 ( \27338 , \26794 );
buf \U$21643 ( \27339 , \26794 );
buf \U$21644 ( \27340 , \26794 );
buf \U$21645 ( \27341 , \26794 );
buf \U$21646 ( \27342 , \26794 );
buf \U$21647 ( \27343 , \26794 );
buf \U$21648 ( \27344 , \26794 );
buf \U$21649 ( \27345 , \26794 );
buf \U$21650 ( \27346 , \26794 );
buf \U$21651 ( \27347 , \26794 );
buf \U$21652 ( \27348 , \26794 );
buf \U$21653 ( \27349 , \26794 );
buf \U$21654 ( \27350 , \26794 );
buf \U$21655 ( \27351 , \26794 );
buf \U$21656 ( \27352 , \26794 );
buf \U$21657 ( \27353 , \26794 );
buf \U$21658 ( \27354 , \26794 );
buf \U$21659 ( \27355 , \26794 );
buf \U$21660 ( \27356 , \26794 );
buf \U$21661 ( \27357 , \26794 );
buf \U$21662 ( \27358 , \26794 );
buf \U$21663 ( \27359 , \26794 );
buf \U$21664 ( \27360 , \26794 );
buf \U$21665 ( \27361 , \26794 );
nor \U$21666 ( \27362 , \26822 , \26823 , \26824 , \26825 , \26787 , \26791 , \26794 , \27337 , \27338 , \27339 , \27340 , \27341 , \27342 , \27343 , \27344 , \27345 , \27346 , \27347 , \27348 , \27349 , \27350 , \27351 , \27352 , \27353 , \27354 , \27355 , \27356 , \27357 , \27358 , \27359 , \27360 , \27361 );
and \U$21667 ( \27363 , \7119 , \27362 );
buf \U$21668 ( \27364 , \26794 );
buf \U$21669 ( \27365 , \26794 );
buf \U$21670 ( \27366 , \26794 );
buf \U$21671 ( \27367 , \26794 );
buf \U$21672 ( \27368 , \26794 );
buf \U$21673 ( \27369 , \26794 );
buf \U$21674 ( \27370 , \26794 );
buf \U$21675 ( \27371 , \26794 );
buf \U$21676 ( \27372 , \26794 );
buf \U$21677 ( \27373 , \26794 );
buf \U$21678 ( \27374 , \26794 );
buf \U$21679 ( \27375 , \26794 );
buf \U$21680 ( \27376 , \26794 );
buf \U$21681 ( \27377 , \26794 );
buf \U$21682 ( \27378 , \26794 );
buf \U$21683 ( \27379 , \26794 );
buf \U$21684 ( \27380 , \26794 );
buf \U$21685 ( \27381 , \26794 );
buf \U$21686 ( \27382 , \26794 );
buf \U$21687 ( \27383 , \26794 );
buf \U$21688 ( \27384 , \26794 );
buf \U$21689 ( \27385 , \26794 );
buf \U$21690 ( \27386 , \26794 );
buf \U$21691 ( \27387 , \26794 );
buf \U$21692 ( \27388 , \26794 );
nor \U$21693 ( \27389 , \26781 , \26823 , \26824 , \26825 , \26787 , \26791 , \26794 , \27364 , \27365 , \27366 , \27367 , \27368 , \27369 , \27370 , \27371 , \27372 , \27373 , \27374 , \27375 , \27376 , \27377 , \27378 , \27379 , \27380 , \27381 , \27382 , \27383 , \27384 , \27385 , \27386 , \27387 , \27388 );
and \U$21694 ( \27390 , \7864 , \27389 );
buf \U$21695 ( \27391 , \26794 );
buf \U$21696 ( \27392 , \26794 );
buf \U$21697 ( \27393 , \26794 );
buf \U$21698 ( \27394 , \26794 );
buf \U$21699 ( \27395 , \26794 );
buf \U$21700 ( \27396 , \26794 );
buf \U$21701 ( \27397 , \26794 );
buf \U$21702 ( \27398 , \26794 );
buf \U$21703 ( \27399 , \26794 );
buf \U$21704 ( \27400 , \26794 );
buf \U$21705 ( \27401 , \26794 );
buf \U$21706 ( \27402 , \26794 );
buf \U$21707 ( \27403 , \26794 );
buf \U$21708 ( \27404 , \26794 );
buf \U$21709 ( \27405 , \26794 );
buf \U$21710 ( \27406 , \26794 );
buf \U$21711 ( \27407 , \26794 );
buf \U$21712 ( \27408 , \26794 );
buf \U$21713 ( \27409 , \26794 );
buf \U$21714 ( \27410 , \26794 );
buf \U$21715 ( \27411 , \26794 );
buf \U$21716 ( \27412 , \26794 );
buf \U$21717 ( \27413 , \26794 );
buf \U$21718 ( \27414 , \26794 );
buf \U$21719 ( \27415 , \26794 );
nor \U$21720 ( \27416 , \26822 , \26782 , \26824 , \26825 , \26787 , \26791 , \26794 , \27391 , \27392 , \27393 , \27394 , \27395 , \27396 , \27397 , \27398 , \27399 , \27400 , \27401 , \27402 , \27403 , \27404 , \27405 , \27406 , \27407 , \27408 , \27409 , \27410 , \27411 , \27412 , \27413 , \27414 , \27415 );
and \U$21721 ( \27417 , \7892 , \27416 );
buf \U$21722 ( \27418 , \26794 );
buf \U$21723 ( \27419 , \26794 );
buf \U$21724 ( \27420 , \26794 );
buf \U$21725 ( \27421 , \26794 );
buf \U$21726 ( \27422 , \26794 );
buf \U$21727 ( \27423 , \26794 );
buf \U$21728 ( \27424 , \26794 );
buf \U$21729 ( \27425 , \26794 );
buf \U$21730 ( \27426 , \26794 );
buf \U$21731 ( \27427 , \26794 );
buf \U$21732 ( \27428 , \26794 );
buf \U$21733 ( \27429 , \26794 );
buf \U$21734 ( \27430 , \26794 );
buf \U$21735 ( \27431 , \26794 );
buf \U$21736 ( \27432 , \26794 );
buf \U$21737 ( \27433 , \26794 );
buf \U$21738 ( \27434 , \26794 );
buf \U$21739 ( \27435 , \26794 );
buf \U$21740 ( \27436 , \26794 );
buf \U$21741 ( \27437 , \26794 );
buf \U$21742 ( \27438 , \26794 );
buf \U$21743 ( \27439 , \26794 );
buf \U$21744 ( \27440 , \26794 );
buf \U$21745 ( \27441 , \26794 );
buf \U$21746 ( \27442 , \26794 );
nor \U$21747 ( \27443 , \26781 , \26782 , \26824 , \26825 , \26787 , \26791 , \26794 , \27418 , \27419 , \27420 , \27421 , \27422 , \27423 , \27424 , \27425 , \27426 , \27427 , \27428 , \27429 , \27430 , \27431 , \27432 , \27433 , \27434 , \27435 , \27436 , \27437 , \27438 , \27439 , \27440 , \27441 , \27442 );
and \U$21748 ( \27444 , \7920 , \27443 );
buf \U$21749 ( \27445 , \26794 );
buf \U$21750 ( \27446 , \26794 );
buf \U$21751 ( \27447 , \26794 );
buf \U$21752 ( \27448 , \26794 );
buf \U$21753 ( \27449 , \26794 );
buf \U$21754 ( \27450 , \26794 );
buf \U$21755 ( \27451 , \26794 );
buf \U$21756 ( \27452 , \26794 );
buf \U$21757 ( \27453 , \26794 );
buf \U$21758 ( \27454 , \26794 );
buf \U$21759 ( \27455 , \26794 );
buf \U$21760 ( \27456 , \26794 );
buf \U$21761 ( \27457 , \26794 );
buf \U$21762 ( \27458 , \26794 );
buf \U$21763 ( \27459 , \26794 );
buf \U$21764 ( \27460 , \26794 );
buf \U$21765 ( \27461 , \26794 );
buf \U$21766 ( \27462 , \26794 );
buf \U$21767 ( \27463 , \26794 );
buf \U$21768 ( \27464 , \26794 );
buf \U$21769 ( \27465 , \26794 );
buf \U$21770 ( \27466 , \26794 );
buf \U$21771 ( \27467 , \26794 );
buf \U$21772 ( \27468 , \26794 );
buf \U$21773 ( \27469 , \26794 );
nor \U$21774 ( \27470 , \26822 , \26823 , \26783 , \26825 , \26787 , \26791 , \26794 , \27445 , \27446 , \27447 , \27448 , \27449 , \27450 , \27451 , \27452 , \27453 , \27454 , \27455 , \27456 , \27457 , \27458 , \27459 , \27460 , \27461 , \27462 , \27463 , \27464 , \27465 , \27466 , \27467 , \27468 , \27469 );
and \U$21775 ( \27471 , \7948 , \27470 );
buf \U$21776 ( \27472 , \26794 );
buf \U$21777 ( \27473 , \26794 );
buf \U$21778 ( \27474 , \26794 );
buf \U$21779 ( \27475 , \26794 );
buf \U$21780 ( \27476 , \26794 );
buf \U$21781 ( \27477 , \26794 );
buf \U$21782 ( \27478 , \26794 );
buf \U$21783 ( \27479 , \26794 );
buf \U$21784 ( \27480 , \26794 );
buf \U$21785 ( \27481 , \26794 );
buf \U$21786 ( \27482 , \26794 );
buf \U$21787 ( \27483 , \26794 );
buf \U$21788 ( \27484 , \26794 );
buf \U$21789 ( \27485 , \26794 );
buf \U$21790 ( \27486 , \26794 );
buf \U$21791 ( \27487 , \26794 );
buf \U$21792 ( \27488 , \26794 );
buf \U$21793 ( \27489 , \26794 );
buf \U$21794 ( \27490 , \26794 );
buf \U$21795 ( \27491 , \26794 );
buf \U$21796 ( \27492 , \26794 );
buf \U$21797 ( \27493 , \26794 );
buf \U$21798 ( \27494 , \26794 );
buf \U$21799 ( \27495 , \26794 );
buf \U$21800 ( \27496 , \26794 );
nor \U$21801 ( \27497 , \26781 , \26823 , \26783 , \26825 , \26787 , \26791 , \26794 , \27472 , \27473 , \27474 , \27475 , \27476 , \27477 , \27478 , \27479 , \27480 , \27481 , \27482 , \27483 , \27484 , \27485 , \27486 , \27487 , \27488 , \27489 , \27490 , \27491 , \27492 , \27493 , \27494 , \27495 , \27496 );
and \U$21802 ( \27498 , \7976 , \27497 );
buf \U$21803 ( \27499 , \26794 );
buf \U$21804 ( \27500 , \26794 );
buf \U$21805 ( \27501 , \26794 );
buf \U$21806 ( \27502 , \26794 );
buf \U$21807 ( \27503 , \26794 );
buf \U$21808 ( \27504 , \26794 );
buf \U$21809 ( \27505 , \26794 );
buf \U$21810 ( \27506 , \26794 );
buf \U$21811 ( \27507 , \26794 );
buf \U$21812 ( \27508 , \26794 );
buf \U$21813 ( \27509 , \26794 );
buf \U$21814 ( \27510 , \26794 );
buf \U$21815 ( \27511 , \26794 );
buf \U$21816 ( \27512 , \26794 );
buf \U$21817 ( \27513 , \26794 );
buf \U$21818 ( \27514 , \26794 );
buf \U$21819 ( \27515 , \26794 );
buf \U$21820 ( \27516 , \26794 );
buf \U$21821 ( \27517 , \26794 );
buf \U$21822 ( \27518 , \26794 );
buf \U$21823 ( \27519 , \26794 );
buf \U$21824 ( \27520 , \26794 );
buf \U$21825 ( \27521 , \26794 );
buf \U$21826 ( \27522 , \26794 );
buf \U$21827 ( \27523 , \26794 );
nor \U$21828 ( \27524 , \26822 , \26782 , \26783 , \26825 , \26787 , \26791 , \26794 , \27499 , \27500 , \27501 , \27502 , \27503 , \27504 , \27505 , \27506 , \27507 , \27508 , \27509 , \27510 , \27511 , \27512 , \27513 , \27514 , \27515 , \27516 , \27517 , \27518 , \27519 , \27520 , \27521 , \27522 , \27523 );
and \U$21829 ( \27525 , \8004 , \27524 );
buf \U$21830 ( \27526 , \26794 );
buf \U$21831 ( \27527 , \26794 );
buf \U$21832 ( \27528 , \26794 );
buf \U$21833 ( \27529 , \26794 );
buf \U$21834 ( \27530 , \26794 );
buf \U$21835 ( \27531 , \26794 );
buf \U$21836 ( \27532 , \26794 );
buf \U$21837 ( \27533 , \26794 );
buf \U$21838 ( \27534 , \26794 );
buf \U$21839 ( \27535 , \26794 );
buf \U$21840 ( \27536 , \26794 );
buf \U$21841 ( \27537 , \26794 );
buf \U$21842 ( \27538 , \26794 );
buf \U$21843 ( \27539 , \26794 );
buf \U$21844 ( \27540 , \26794 );
buf \U$21845 ( \27541 , \26794 );
buf \U$21846 ( \27542 , \26794 );
buf \U$21847 ( \27543 , \26794 );
buf \U$21848 ( \27544 , \26794 );
buf \U$21849 ( \27545 , \26794 );
buf \U$21850 ( \27546 , \26794 );
buf \U$21851 ( \27547 , \26794 );
buf \U$21852 ( \27548 , \26794 );
buf \U$21853 ( \27549 , \26794 );
buf \U$21854 ( \27550 , \26794 );
nor \U$21855 ( \27551 , \26781 , \26782 , \26783 , \26825 , \26787 , \26791 , \26794 , \27526 , \27527 , \27528 , \27529 , \27530 , \27531 , \27532 , \27533 , \27534 , \27535 , \27536 , \27537 , \27538 , \27539 , \27540 , \27541 , \27542 , \27543 , \27544 , \27545 , \27546 , \27547 , \27548 , \27549 , \27550 );
and \U$21856 ( \27552 , \8032 , \27551 );
buf \U$21857 ( \27553 , \26794 );
buf \U$21858 ( \27554 , \26794 );
buf \U$21859 ( \27555 , \26794 );
buf \U$21860 ( \27556 , \26794 );
buf \U$21861 ( \27557 , \26794 );
buf \U$21862 ( \27558 , \26794 );
buf \U$21863 ( \27559 , \26794 );
buf \U$21864 ( \27560 , \26794 );
buf \U$21865 ( \27561 , \26794 );
buf \U$21866 ( \27562 , \26794 );
buf \U$21867 ( \27563 , \26794 );
buf \U$21868 ( \27564 , \26794 );
buf \U$21869 ( \27565 , \26794 );
buf \U$21870 ( \27566 , \26794 );
buf \U$21871 ( \27567 , \26794 );
buf \U$21872 ( \27568 , \26794 );
buf \U$21873 ( \27569 , \26794 );
buf \U$21874 ( \27570 , \26794 );
buf \U$21875 ( \27571 , \26794 );
buf \U$21876 ( \27572 , \26794 );
buf \U$21877 ( \27573 , \26794 );
buf \U$21878 ( \27574 , \26794 );
buf \U$21879 ( \27575 , \26794 );
buf \U$21880 ( \27576 , \26794 );
buf \U$21881 ( \27577 , \26794 );
nor \U$21882 ( \27578 , \26822 , \26823 , \26824 , \26784 , \26787 , \26791 , \26794 , \27553 , \27554 , \27555 , \27556 , \27557 , \27558 , \27559 , \27560 , \27561 , \27562 , \27563 , \27564 , \27565 , \27566 , \27567 , \27568 , \27569 , \27570 , \27571 , \27572 , \27573 , \27574 , \27575 , \27576 , \27577 );
and \U$21883 ( \27579 , \8060 , \27578 );
buf \U$21884 ( \27580 , \26794 );
buf \U$21885 ( \27581 , \26794 );
buf \U$21886 ( \27582 , \26794 );
buf \U$21887 ( \27583 , \26794 );
buf \U$21888 ( \27584 , \26794 );
buf \U$21889 ( \27585 , \26794 );
buf \U$21890 ( \27586 , \26794 );
buf \U$21891 ( \27587 , \26794 );
buf \U$21892 ( \27588 , \26794 );
buf \U$21893 ( \27589 , \26794 );
buf \U$21894 ( \27590 , \26794 );
buf \U$21895 ( \27591 , \26794 );
buf \U$21896 ( \27592 , \26794 );
buf \U$21897 ( \27593 , \26794 );
buf \U$21898 ( \27594 , \26794 );
buf \U$21899 ( \27595 , \26794 );
buf \U$21900 ( \27596 , \26794 );
buf \U$21901 ( \27597 , \26794 );
buf \U$21902 ( \27598 , \26794 );
buf \U$21903 ( \27599 , \26794 );
buf \U$21904 ( \27600 , \26794 );
buf \U$21905 ( \27601 , \26794 );
buf \U$21906 ( \27602 , \26794 );
buf \U$21907 ( \27603 , \26794 );
buf \U$21908 ( \27604 , \26794 );
nor \U$21909 ( \27605 , \26781 , \26823 , \26824 , \26784 , \26787 , \26791 , \26794 , \27580 , \27581 , \27582 , \27583 , \27584 , \27585 , \27586 , \27587 , \27588 , \27589 , \27590 , \27591 , \27592 , \27593 , \27594 , \27595 , \27596 , \27597 , \27598 , \27599 , \27600 , \27601 , \27602 , \27603 , \27604 );
and \U$21910 ( \27606 , \8088 , \27605 );
buf \U$21911 ( \27607 , \26794 );
buf \U$21912 ( \27608 , \26794 );
buf \U$21913 ( \27609 , \26794 );
buf \U$21914 ( \27610 , \26794 );
buf \U$21915 ( \27611 , \26794 );
buf \U$21916 ( \27612 , \26794 );
buf \U$21917 ( \27613 , \26794 );
buf \U$21918 ( \27614 , \26794 );
buf \U$21919 ( \27615 , \26794 );
buf \U$21920 ( \27616 , \26794 );
buf \U$21921 ( \27617 , \26794 );
buf \U$21922 ( \27618 , \26794 );
buf \U$21923 ( \27619 , \26794 );
buf \U$21924 ( \27620 , \26794 );
buf \U$21925 ( \27621 , \26794 );
buf \U$21926 ( \27622 , \26794 );
buf \U$21927 ( \27623 , \26794 );
buf \U$21928 ( \27624 , \26794 );
buf \U$21929 ( \27625 , \26794 );
buf \U$21930 ( \27626 , \26794 );
buf \U$21931 ( \27627 , \26794 );
buf \U$21932 ( \27628 , \26794 );
buf \U$21933 ( \27629 , \26794 );
buf \U$21934 ( \27630 , \26794 );
buf \U$21935 ( \27631 , \26794 );
nor \U$21936 ( \27632 , \26822 , \26782 , \26824 , \26784 , \26787 , \26791 , \26794 , \27607 , \27608 , \27609 , \27610 , \27611 , \27612 , \27613 , \27614 , \27615 , \27616 , \27617 , \27618 , \27619 , \27620 , \27621 , \27622 , \27623 , \27624 , \27625 , \27626 , \27627 , \27628 , \27629 , \27630 , \27631 );
and \U$21937 ( \27633 , \8116 , \27632 );
buf \U$21938 ( \27634 , \26794 );
buf \U$21939 ( \27635 , \26794 );
buf \U$21940 ( \27636 , \26794 );
buf \U$21941 ( \27637 , \26794 );
buf \U$21942 ( \27638 , \26794 );
buf \U$21943 ( \27639 , \26794 );
buf \U$21944 ( \27640 , \26794 );
buf \U$21945 ( \27641 , \26794 );
buf \U$21946 ( \27642 , \26794 );
buf \U$21947 ( \27643 , \26794 );
buf \U$21948 ( \27644 , \26794 );
buf \U$21949 ( \27645 , \26794 );
buf \U$21950 ( \27646 , \26794 );
buf \U$21951 ( \27647 , \26794 );
buf \U$21952 ( \27648 , \26794 );
buf \U$21953 ( \27649 , \26794 );
buf \U$21954 ( \27650 , \26794 );
buf \U$21955 ( \27651 , \26794 );
buf \U$21956 ( \27652 , \26794 );
buf \U$21957 ( \27653 , \26794 );
buf \U$21958 ( \27654 , \26794 );
buf \U$21959 ( \27655 , \26794 );
buf \U$21960 ( \27656 , \26794 );
buf \U$21961 ( \27657 , \26794 );
buf \U$21962 ( \27658 , \26794 );
nor \U$21963 ( \27659 , \26781 , \26782 , \26824 , \26784 , \26787 , \26791 , \26794 , \27634 , \27635 , \27636 , \27637 , \27638 , \27639 , \27640 , \27641 , \27642 , \27643 , \27644 , \27645 , \27646 , \27647 , \27648 , \27649 , \27650 , \27651 , \27652 , \27653 , \27654 , \27655 , \27656 , \27657 , \27658 );
and \U$21964 ( \27660 , \8144 , \27659 );
buf \U$21965 ( \27661 , \26794 );
buf \U$21966 ( \27662 , \26794 );
buf \U$21967 ( \27663 , \26794 );
buf \U$21968 ( \27664 , \26794 );
buf \U$21969 ( \27665 , \26794 );
buf \U$21970 ( \27666 , \26794 );
buf \U$21971 ( \27667 , \26794 );
buf \U$21972 ( \27668 , \26794 );
buf \U$21973 ( \27669 , \26794 );
buf \U$21974 ( \27670 , \26794 );
buf \U$21975 ( \27671 , \26794 );
buf \U$21976 ( \27672 , \26794 );
buf \U$21977 ( \27673 , \26794 );
buf \U$21978 ( \27674 , \26794 );
buf \U$21979 ( \27675 , \26794 );
buf \U$21980 ( \27676 , \26794 );
buf \U$21981 ( \27677 , \26794 );
buf \U$21982 ( \27678 , \26794 );
buf \U$21983 ( \27679 , \26794 );
buf \U$21984 ( \27680 , \26794 );
buf \U$21985 ( \27681 , \26794 );
buf \U$21986 ( \27682 , \26794 );
buf \U$21987 ( \27683 , \26794 );
buf \U$21988 ( \27684 , \26794 );
buf \U$21989 ( \27685 , \26794 );
nor \U$21990 ( \27686 , \26822 , \26823 , \26783 , \26784 , \26787 , \26791 , \26794 , \27661 , \27662 , \27663 , \27664 , \27665 , \27666 , \27667 , \27668 , \27669 , \27670 , \27671 , \27672 , \27673 , \27674 , \27675 , \27676 , \27677 , \27678 , \27679 , \27680 , \27681 , \27682 , \27683 , \27684 , \27685 );
and \U$21991 ( \27687 , \8172 , \27686 );
buf \U$21992 ( \27688 , \26794 );
buf \U$21993 ( \27689 , \26794 );
buf \U$21994 ( \27690 , \26794 );
buf \U$21995 ( \27691 , \26794 );
buf \U$21996 ( \27692 , \26794 );
buf \U$21997 ( \27693 , \26794 );
buf \U$21998 ( \27694 , \26794 );
buf \U$21999 ( \27695 , \26794 );
buf \U$22000 ( \27696 , \26794 );
buf \U$22001 ( \27697 , \26794 );
buf \U$22002 ( \27698 , \26794 );
buf \U$22003 ( \27699 , \26794 );
buf \U$22004 ( \27700 , \26794 );
buf \U$22005 ( \27701 , \26794 );
buf \U$22006 ( \27702 , \26794 );
buf \U$22007 ( \27703 , \26794 );
buf \U$22008 ( \27704 , \26794 );
buf \U$22009 ( \27705 , \26794 );
buf \U$22010 ( \27706 , \26794 );
buf \U$22011 ( \27707 , \26794 );
buf \U$22012 ( \27708 , \26794 );
buf \U$22013 ( \27709 , \26794 );
buf \U$22014 ( \27710 , \26794 );
buf \U$22015 ( \27711 , \26794 );
buf \U$22016 ( \27712 , \26794 );
nor \U$22017 ( \27713 , \26781 , \26823 , \26783 , \26784 , \26787 , \26791 , \26794 , \27688 , \27689 , \27690 , \27691 , \27692 , \27693 , \27694 , \27695 , \27696 , \27697 , \27698 , \27699 , \27700 , \27701 , \27702 , \27703 , \27704 , \27705 , \27706 , \27707 , \27708 , \27709 , \27710 , \27711 , \27712 );
and \U$22018 ( \27714 , \8200 , \27713 );
buf \U$22019 ( \27715 , \26794 );
buf \U$22020 ( \27716 , \26794 );
buf \U$22021 ( \27717 , \26794 );
buf \U$22022 ( \27718 , \26794 );
buf \U$22023 ( \27719 , \26794 );
buf \U$22024 ( \27720 , \26794 );
buf \U$22025 ( \27721 , \26794 );
buf \U$22026 ( \27722 , \26794 );
buf \U$22027 ( \27723 , \26794 );
buf \U$22028 ( \27724 , \26794 );
buf \U$22029 ( \27725 , \26794 );
buf \U$22030 ( \27726 , \26794 );
buf \U$22031 ( \27727 , \26794 );
buf \U$22032 ( \27728 , \26794 );
buf \U$22033 ( \27729 , \26794 );
buf \U$22034 ( \27730 , \26794 );
buf \U$22035 ( \27731 , \26794 );
buf \U$22036 ( \27732 , \26794 );
buf \U$22037 ( \27733 , \26794 );
buf \U$22038 ( \27734 , \26794 );
buf \U$22039 ( \27735 , \26794 );
buf \U$22040 ( \27736 , \26794 );
buf \U$22041 ( \27737 , \26794 );
buf \U$22042 ( \27738 , \26794 );
buf \U$22043 ( \27739 , \26794 );
nor \U$22044 ( \27740 , \26822 , \26782 , \26783 , \26784 , \26787 , \26791 , \26794 , \27715 , \27716 , \27717 , \27718 , \27719 , \27720 , \27721 , \27722 , \27723 , \27724 , \27725 , \27726 , \27727 , \27728 , \27729 , \27730 , \27731 , \27732 , \27733 , \27734 , \27735 , \27736 , \27737 , \27738 , \27739 );
and \U$22045 ( \27741 , \8228 , \27740 );
or \U$22046 ( \27742 , \27336 , \27363 , \27390 , \27417 , \27444 , \27471 , \27498 , \27525 , \27552 , \27579 , \27606 , \27633 , \27660 , \27687 , \27714 , \27741 );
buf \U$22047 ( \27743 , \26794 );
not \U$22048 ( \27744 , \27743 );
buf \U$22049 ( \27745 , \26782 );
buf \U$22050 ( \27746 , \26783 );
buf \U$22051 ( \27747 , \26784 );
buf \U$22052 ( \27748 , \26787 );
buf \U$22053 ( \27749 , \26791 );
buf \U$22054 ( \27750 , \26794 );
buf \U$22055 ( \27751 , \26794 );
buf \U$22056 ( \27752 , \26794 );
buf \U$22057 ( \27753 , \26794 );
buf \U$22058 ( \27754 , \26794 );
buf \U$22059 ( \27755 , \26794 );
buf \U$22060 ( \27756 , \26794 );
buf \U$22061 ( \27757 , \26794 );
buf \U$22062 ( \27758 , \26794 );
buf \U$22063 ( \27759 , \26794 );
buf \U$22064 ( \27760 , \26794 );
buf \U$22065 ( \27761 , \26794 );
buf \U$22066 ( \27762 , \26794 );
buf \U$22067 ( \27763 , \26794 );
buf \U$22068 ( \27764 , \26794 );
buf \U$22069 ( \27765 , \26794 );
buf \U$22070 ( \27766 , \26794 );
buf \U$22071 ( \27767 , \26794 );
buf \U$22072 ( \27768 , \26794 );
buf \U$22073 ( \27769 , \26794 );
buf \U$22074 ( \27770 , \26794 );
buf \U$22075 ( \27771 , \26794 );
buf \U$22076 ( \27772 , \26794 );
buf \U$22077 ( \27773 , \26794 );
buf \U$22078 ( \27774 , \26794 );
buf \U$22079 ( \27775 , \26781 );
or \U$22080 ( \27776 , \27745 , \27746 , \27747 , \27748 , \27749 , \27750 , \27751 , \27752 , \27753 , \27754 , \27755 , \27756 , \27757 , \27758 , \27759 , \27760 , \27761 , \27762 , \27763 , \27764 , \27765 , \27766 , \27767 , \27768 , \27769 , \27770 , \27771 , \27772 , \27773 , \27774 , \27775 );
nand \U$22081 ( \27777 , \27744 , \27776 );
buf \U$22082 ( \27778 , \27777 );
buf \U$22083 ( \27779 , \26794 );
not \U$22084 ( \27780 , \27779 );
buf \U$22085 ( \27781 , \26791 );
buf \U$22086 ( \27782 , \26794 );
buf \U$22087 ( \27783 , \26794 );
buf \U$22088 ( \27784 , \26794 );
buf \U$22089 ( \27785 , \26794 );
buf \U$22090 ( \27786 , \26794 );
buf \U$22091 ( \27787 , \26794 );
buf \U$22092 ( \27788 , \26794 );
buf \U$22093 ( \27789 , \26794 );
buf \U$22094 ( \27790 , \26794 );
buf \U$22095 ( \27791 , \26794 );
buf \U$22096 ( \27792 , \26794 );
buf \U$22097 ( \27793 , \26794 );
buf \U$22098 ( \27794 , \26794 );
buf \U$22099 ( \27795 , \26794 );
buf \U$22100 ( \27796 , \26794 );
buf \U$22101 ( \27797 , \26794 );
buf \U$22102 ( \27798 , \26794 );
buf \U$22103 ( \27799 , \26794 );
buf \U$22104 ( \27800 , \26794 );
buf \U$22105 ( \27801 , \26794 );
buf \U$22106 ( \27802 , \26794 );
buf \U$22107 ( \27803 , \26794 );
buf \U$22108 ( \27804 , \26794 );
buf \U$22109 ( \27805 , \26794 );
buf \U$22110 ( \27806 , \26794 );
buf \U$22111 ( \27807 , \26787 );
buf \U$22112 ( \27808 , \26781 );
buf \U$22113 ( \27809 , \26782 );
buf \U$22114 ( \27810 , \26783 );
buf \U$22115 ( \27811 , \26784 );
or \U$22116 ( \27812 , \27808 , \27809 , \27810 , \27811 );
and \U$22117 ( \27813 , \27807 , \27812 );
or \U$22118 ( \27814 , \27781 , \27782 , \27783 , \27784 , \27785 , \27786 , \27787 , \27788 , \27789 , \27790 , \27791 , \27792 , \27793 , \27794 , \27795 , \27796 , \27797 , \27798 , \27799 , \27800 , \27801 , \27802 , \27803 , \27804 , \27805 , \27806 , \27813 );
and \U$22119 ( \27815 , \27780 , \27814 );
buf \U$22120 ( \27816 , \27815 );
or \U$22121 ( \27817 , \27778 , \27816 );
_DC g83ab ( \27818_nG83ab , \27742 , \27817 );
buf \U$22122 ( \27819 , \27818_nG83ab );
xor \U$22123 ( \27820 , \27309 , \27819 );
buf \U$22124 ( \27821 , RIb7b9590_247);
and \U$22125 ( \27822 , \7126 , \27335 );
and \U$22126 ( \27823 , \7128 , \27362 );
and \U$22127 ( \27824 , \8338 , \27389 );
and \U$22128 ( \27825 , \8340 , \27416 );
and \U$22129 ( \27826 , \8342 , \27443 );
and \U$22130 ( \27827 , \8344 , \27470 );
and \U$22131 ( \27828 , \8346 , \27497 );
and \U$22132 ( \27829 , \8348 , \27524 );
and \U$22133 ( \27830 , \8350 , \27551 );
and \U$22134 ( \27831 , \8352 , \27578 );
and \U$22135 ( \27832 , \8354 , \27605 );
and \U$22136 ( \27833 , \8356 , \27632 );
and \U$22137 ( \27834 , \8358 , \27659 );
and \U$22138 ( \27835 , \8360 , \27686 );
and \U$22139 ( \27836 , \8362 , \27713 );
and \U$22140 ( \27837 , \8364 , \27740 );
or \U$22141 ( \27838 , \27822 , \27823 , \27824 , \27825 , \27826 , \27827 , \27828 , \27829 , \27830 , \27831 , \27832 , \27833 , \27834 , \27835 , \27836 , \27837 );
_DC g83c0 ( \27839_nG83c0 , \27838 , \27817 );
buf \U$22142 ( \27840 , \27839_nG83c0 );
xor \U$22143 ( \27841 , \27821 , \27840 );
or \U$22144 ( \27842 , \27820 , \27841 );
buf \U$22145 ( \27843 , RIb7b9518_248);
and \U$22146 ( \27844 , \7136 , \27335 );
and \U$22147 ( \27845 , \7138 , \27362 );
and \U$22148 ( \27846 , \8374 , \27389 );
and \U$22149 ( \27847 , \8376 , \27416 );
and \U$22150 ( \27848 , \8378 , \27443 );
and \U$22151 ( \27849 , \8380 , \27470 );
and \U$22152 ( \27850 , \8382 , \27497 );
and \U$22153 ( \27851 , \8384 , \27524 );
and \U$22154 ( \27852 , \8386 , \27551 );
and \U$22155 ( \27853 , \8388 , \27578 );
and \U$22156 ( \27854 , \8390 , \27605 );
and \U$22157 ( \27855 , \8392 , \27632 );
and \U$22158 ( \27856 , \8394 , \27659 );
and \U$22159 ( \27857 , \8396 , \27686 );
and \U$22160 ( \27858 , \8398 , \27713 );
and \U$22161 ( \27859 , \8400 , \27740 );
or \U$22162 ( \27860 , \27844 , \27845 , \27846 , \27847 , \27848 , \27849 , \27850 , \27851 , \27852 , \27853 , \27854 , \27855 , \27856 , \27857 , \27858 , \27859 );
_DC g83d6 ( \27861_nG83d6 , \27860 , \27817 );
buf \U$22163 ( \27862 , \27861_nG83d6 );
xor \U$22164 ( \27863 , \27843 , \27862 );
or \U$22165 ( \27864 , \27842 , \27863 );
buf \U$22166 ( \27865 , RIb7b94a0_249);
and \U$22167 ( \27866 , \7146 , \27335 );
and \U$22168 ( \27867 , \7148 , \27362 );
and \U$22169 ( \27868 , \8410 , \27389 );
and \U$22170 ( \27869 , \8412 , \27416 );
and \U$22171 ( \27870 , \8414 , \27443 );
and \U$22172 ( \27871 , \8416 , \27470 );
and \U$22173 ( \27872 , \8418 , \27497 );
and \U$22174 ( \27873 , \8420 , \27524 );
and \U$22175 ( \27874 , \8422 , \27551 );
and \U$22176 ( \27875 , \8424 , \27578 );
and \U$22177 ( \27876 , \8426 , \27605 );
and \U$22178 ( \27877 , \8428 , \27632 );
and \U$22179 ( \27878 , \8430 , \27659 );
and \U$22180 ( \27879 , \8432 , \27686 );
and \U$22181 ( \27880 , \8434 , \27713 );
and \U$22182 ( \27881 , \8436 , \27740 );
or \U$22183 ( \27882 , \27866 , \27867 , \27868 , \27869 , \27870 , \27871 , \27872 , \27873 , \27874 , \27875 , \27876 , \27877 , \27878 , \27879 , \27880 , \27881 );
_DC g83ec ( \27883_nG83ec , \27882 , \27817 );
buf \U$22184 ( \27884 , \27883_nG83ec );
xor \U$22185 ( \27885 , \27865 , \27884 );
or \U$22186 ( \27886 , \27864 , \27885 );
buf \U$22187 ( \27887 , RIb7b9428_250);
and \U$22188 ( \27888 , \7156 , \27335 );
and \U$22189 ( \27889 , \7158 , \27362 );
and \U$22190 ( \27890 , \8446 , \27389 );
and \U$22191 ( \27891 , \8448 , \27416 );
and \U$22192 ( \27892 , \8450 , \27443 );
and \U$22193 ( \27893 , \8452 , \27470 );
and \U$22194 ( \27894 , \8454 , \27497 );
and \U$22195 ( \27895 , \8456 , \27524 );
and \U$22196 ( \27896 , \8458 , \27551 );
and \U$22197 ( \27897 , \8460 , \27578 );
and \U$22198 ( \27898 , \8462 , \27605 );
and \U$22199 ( \27899 , \8464 , \27632 );
and \U$22200 ( \27900 , \8466 , \27659 );
and \U$22201 ( \27901 , \8468 , \27686 );
and \U$22202 ( \27902 , \8470 , \27713 );
and \U$22203 ( \27903 , \8472 , \27740 );
or \U$22204 ( \27904 , \27888 , \27889 , \27890 , \27891 , \27892 , \27893 , \27894 , \27895 , \27896 , \27897 , \27898 , \27899 , \27900 , \27901 , \27902 , \27903 );
_DC g8402 ( \27905_nG8402 , \27904 , \27817 );
buf \U$22205 ( \27906 , \27905_nG8402 );
xor \U$22206 ( \27907 , \27887 , \27906 );
or \U$22207 ( \27908 , \27886 , \27907 );
buf \U$22208 ( \27909 , RIb7b93b0_251);
and \U$22209 ( \27910 , \7166 , \27335 );
and \U$22210 ( \27911 , \7168 , \27362 );
and \U$22211 ( \27912 , \8482 , \27389 );
and \U$22212 ( \27913 , \8484 , \27416 );
and \U$22213 ( \27914 , \8486 , \27443 );
and \U$22214 ( \27915 , \8488 , \27470 );
and \U$22215 ( \27916 , \8490 , \27497 );
and \U$22216 ( \27917 , \8492 , \27524 );
and \U$22217 ( \27918 , \8494 , \27551 );
and \U$22218 ( \27919 , \8496 , \27578 );
and \U$22219 ( \27920 , \8498 , \27605 );
and \U$22220 ( \27921 , \8500 , \27632 );
and \U$22221 ( \27922 , \8502 , \27659 );
and \U$22222 ( \27923 , \8504 , \27686 );
and \U$22223 ( \27924 , \8506 , \27713 );
and \U$22224 ( \27925 , \8508 , \27740 );
or \U$22225 ( \27926 , \27910 , \27911 , \27912 , \27913 , \27914 , \27915 , \27916 , \27917 , \27918 , \27919 , \27920 , \27921 , \27922 , \27923 , \27924 , \27925 );
_DC g8418 ( \27927_nG8418 , \27926 , \27817 );
buf \U$22226 ( \27928 , \27927_nG8418 );
xor \U$22227 ( \27929 , \27909 , \27928 );
or \U$22228 ( \27930 , \27908 , \27929 );
buf \U$22229 ( \27931 , RIb7af720_252);
and \U$22230 ( \27932 , \7176 , \27335 );
and \U$22231 ( \27933 , \7178 , \27362 );
and \U$22232 ( \27934 , \8518 , \27389 );
and \U$22233 ( \27935 , \8520 , \27416 );
and \U$22234 ( \27936 , \8522 , \27443 );
and \U$22235 ( \27937 , \8524 , \27470 );
and \U$22236 ( \27938 , \8526 , \27497 );
and \U$22237 ( \27939 , \8528 , \27524 );
and \U$22238 ( \27940 , \8530 , \27551 );
and \U$22239 ( \27941 , \8532 , \27578 );
and \U$22240 ( \27942 , \8534 , \27605 );
and \U$22241 ( \27943 , \8536 , \27632 );
and \U$22242 ( \27944 , \8538 , \27659 );
and \U$22243 ( \27945 , \8540 , \27686 );
and \U$22244 ( \27946 , \8542 , \27713 );
and \U$22245 ( \27947 , \8544 , \27740 );
or \U$22246 ( \27948 , \27932 , \27933 , \27934 , \27935 , \27936 , \27937 , \27938 , \27939 , \27940 , \27941 , \27942 , \27943 , \27944 , \27945 , \27946 , \27947 );
_DC g842e ( \27949_nG842e , \27948 , \27817 );
buf \U$22247 ( \27950 , \27949_nG842e );
xor \U$22248 ( \27951 , \27931 , \27950 );
or \U$22249 ( \27952 , \27930 , \27951 );
buf \U$22250 ( \27953 , RIb7af6a8_253);
and \U$22251 ( \27954 , \7186 , \27335 );
and \U$22252 ( \27955 , \7188 , \27362 );
and \U$22253 ( \27956 , \8554 , \27389 );
and \U$22254 ( \27957 , \8556 , \27416 );
and \U$22255 ( \27958 , \8558 , \27443 );
and \U$22256 ( \27959 , \8560 , \27470 );
and \U$22257 ( \27960 , \8562 , \27497 );
and \U$22258 ( \27961 , \8564 , \27524 );
and \U$22259 ( \27962 , \8566 , \27551 );
and \U$22260 ( \27963 , \8568 , \27578 );
and \U$22261 ( \27964 , \8570 , \27605 );
and \U$22262 ( \27965 , \8572 , \27632 );
and \U$22263 ( \27966 , \8574 , \27659 );
and \U$22264 ( \27967 , \8576 , \27686 );
and \U$22265 ( \27968 , \8578 , \27713 );
and \U$22266 ( \27969 , \8580 , \27740 );
or \U$22267 ( \27970 , \27954 , \27955 , \27956 , \27957 , \27958 , \27959 , \27960 , \27961 , \27962 , \27963 , \27964 , \27965 , \27966 , \27967 , \27968 , \27969 );
_DC g8444 ( \27971_nG8444 , \27970 , \27817 );
buf \U$22268 ( \27972 , \27971_nG8444 );
xor \U$22269 ( \27973 , \27953 , \27972 );
or \U$22270 ( \27974 , \27952 , \27973 );
not \U$22271 ( \27975 , \27974 );
buf \U$22272 ( \27976 , \27975 );
and \U$22273 ( \27977 , \27308 , \27976 );
buf \U$22274 ( \27978 , RIb7af630_254);
buf \U$22275 ( \27979 , \26794 );
buf \U$22276 ( \27980 , \26794 );
buf \U$22277 ( \27981 , \26794 );
buf \U$22278 ( \27982 , \26794 );
buf \U$22279 ( \27983 , \26794 );
buf \U$22280 ( \27984 , \26794 );
buf \U$22281 ( \27985 , \26794 );
buf \U$22282 ( \27986 , \26794 );
buf \U$22283 ( \27987 , \26794 );
buf \U$22284 ( \27988 , \26794 );
buf \U$22285 ( \27989 , \26794 );
buf \U$22286 ( \27990 , \26794 );
buf \U$22287 ( \27991 , \26794 );
buf \U$22288 ( \27992 , \26794 );
buf \U$22289 ( \27993 , \26794 );
buf \U$22290 ( \27994 , \26794 );
buf \U$22291 ( \27995 , \26794 );
buf \U$22292 ( \27996 , \26794 );
buf \U$22293 ( \27997 , \26794 );
buf \U$22294 ( \27998 , \26794 );
buf \U$22295 ( \27999 , \26794 );
buf \U$22296 ( \28000 , \26794 );
buf \U$22297 ( \28001 , \26794 );
buf \U$22298 ( \28002 , \26794 );
buf \U$22299 ( \28003 , \26794 );
nor \U$22300 ( \28004 , \26781 , \26782 , \26783 , \26784 , \26788 , \26791 , \26794 , \27979 , \27980 , \27981 , \27982 , \27983 , \27984 , \27985 , \27986 , \27987 , \27988 , \27989 , \27990 , \27991 , \27992 , \27993 , \27994 , \27995 , \27996 , \27997 , \27998 , \27999 , \28000 , \28001 , \28002 , \28003 );
and \U$22301 ( \28005 , \7198 , \28004 );
buf \U$22302 ( \28006 , \26794 );
buf \U$22303 ( \28007 , \26794 );
buf \U$22304 ( \28008 , \26794 );
buf \U$22305 ( \28009 , \26794 );
buf \U$22306 ( \28010 , \26794 );
buf \U$22307 ( \28011 , \26794 );
buf \U$22308 ( \28012 , \26794 );
buf \U$22309 ( \28013 , \26794 );
buf \U$22310 ( \28014 , \26794 );
buf \U$22311 ( \28015 , \26794 );
buf \U$22312 ( \28016 , \26794 );
buf \U$22313 ( \28017 , \26794 );
buf \U$22314 ( \28018 , \26794 );
buf \U$22315 ( \28019 , \26794 );
buf \U$22316 ( \28020 , \26794 );
buf \U$22317 ( \28021 , \26794 );
buf \U$22318 ( \28022 , \26794 );
buf \U$22319 ( \28023 , \26794 );
buf \U$22320 ( \28024 , \26794 );
buf \U$22321 ( \28025 , \26794 );
buf \U$22322 ( \28026 , \26794 );
buf \U$22323 ( \28027 , \26794 );
buf \U$22324 ( \28028 , \26794 );
buf \U$22325 ( \28029 , \26794 );
buf \U$22326 ( \28030 , \26794 );
nor \U$22327 ( \28031 , \26822 , \26823 , \26824 , \26825 , \26787 , \26791 , \26794 , \28006 , \28007 , \28008 , \28009 , \28010 , \28011 , \28012 , \28013 , \28014 , \28015 , \28016 , \28017 , \28018 , \28019 , \28020 , \28021 , \28022 , \28023 , \28024 , \28025 , \28026 , \28027 , \28028 , \28029 , \28030 );
and \U$22328 ( \28032 , \7200 , \28031 );
buf \U$22329 ( \28033 , \26794 );
buf \U$22330 ( \28034 , \26794 );
buf \U$22331 ( \28035 , \26794 );
buf \U$22332 ( \28036 , \26794 );
buf \U$22333 ( \28037 , \26794 );
buf \U$22334 ( \28038 , \26794 );
buf \U$22335 ( \28039 , \26794 );
buf \U$22336 ( \28040 , \26794 );
buf \U$22337 ( \28041 , \26794 );
buf \U$22338 ( \28042 , \26794 );
buf \U$22339 ( \28043 , \26794 );
buf \U$22340 ( \28044 , \26794 );
buf \U$22341 ( \28045 , \26794 );
buf \U$22342 ( \28046 , \26794 );
buf \U$22343 ( \28047 , \26794 );
buf \U$22344 ( \28048 , \26794 );
buf \U$22345 ( \28049 , \26794 );
buf \U$22346 ( \28050 , \26794 );
buf \U$22347 ( \28051 , \26794 );
buf \U$22348 ( \28052 , \26794 );
buf \U$22349 ( \28053 , \26794 );
buf \U$22350 ( \28054 , \26794 );
buf \U$22351 ( \28055 , \26794 );
buf \U$22352 ( \28056 , \26794 );
buf \U$22353 ( \28057 , \26794 );
nor \U$22354 ( \28058 , \26781 , \26823 , \26824 , \26825 , \26787 , \26791 , \26794 , \28033 , \28034 , \28035 , \28036 , \28037 , \28038 , \28039 , \28040 , \28041 , \28042 , \28043 , \28044 , \28045 , \28046 , \28047 , \28048 , \28049 , \28050 , \28051 , \28052 , \28053 , \28054 , \28055 , \28056 , \28057 );
and \U$22355 ( \28059 , \8645 , \28058 );
buf \U$22356 ( \28060 , \26794 );
buf \U$22357 ( \28061 , \26794 );
buf \U$22358 ( \28062 , \26794 );
buf \U$22359 ( \28063 , \26794 );
buf \U$22360 ( \28064 , \26794 );
buf \U$22361 ( \28065 , \26794 );
buf \U$22362 ( \28066 , \26794 );
buf \U$22363 ( \28067 , \26794 );
buf \U$22364 ( \28068 , \26794 );
buf \U$22365 ( \28069 , \26794 );
buf \U$22366 ( \28070 , \26794 );
buf \U$22367 ( \28071 , \26794 );
buf \U$22368 ( \28072 , \26794 );
buf \U$22369 ( \28073 , \26794 );
buf \U$22370 ( \28074 , \26794 );
buf \U$22371 ( \28075 , \26794 );
buf \U$22372 ( \28076 , \26794 );
buf \U$22373 ( \28077 , \26794 );
buf \U$22374 ( \28078 , \26794 );
buf \U$22375 ( \28079 , \26794 );
buf \U$22376 ( \28080 , \26794 );
buf \U$22377 ( \28081 , \26794 );
buf \U$22378 ( \28082 , \26794 );
buf \U$22379 ( \28083 , \26794 );
buf \U$22380 ( \28084 , \26794 );
nor \U$22381 ( \28085 , \26822 , \26782 , \26824 , \26825 , \26787 , \26791 , \26794 , \28060 , \28061 , \28062 , \28063 , \28064 , \28065 , \28066 , \28067 , \28068 , \28069 , \28070 , \28071 , \28072 , \28073 , \28074 , \28075 , \28076 , \28077 , \28078 , \28079 , \28080 , \28081 , \28082 , \28083 , \28084 );
and \U$22382 ( \28086 , \8673 , \28085 );
buf \U$22383 ( \28087 , \26794 );
buf \U$22384 ( \28088 , \26794 );
buf \U$22385 ( \28089 , \26794 );
buf \U$22386 ( \28090 , \26794 );
buf \U$22387 ( \28091 , \26794 );
buf \U$22388 ( \28092 , \26794 );
buf \U$22389 ( \28093 , \26794 );
buf \U$22390 ( \28094 , \26794 );
buf \U$22391 ( \28095 , \26794 );
buf \U$22392 ( \28096 , \26794 );
buf \U$22393 ( \28097 , \26794 );
buf \U$22394 ( \28098 , \26794 );
buf \U$22395 ( \28099 , \26794 );
buf \U$22396 ( \28100 , \26794 );
buf \U$22397 ( \28101 , \26794 );
buf \U$22398 ( \28102 , \26794 );
buf \U$22399 ( \28103 , \26794 );
buf \U$22400 ( \28104 , \26794 );
buf \U$22401 ( \28105 , \26794 );
buf \U$22402 ( \28106 , \26794 );
buf \U$22403 ( \28107 , \26794 );
buf \U$22404 ( \28108 , \26794 );
buf \U$22405 ( \28109 , \26794 );
buf \U$22406 ( \28110 , \26794 );
buf \U$22407 ( \28111 , \26794 );
nor \U$22408 ( \28112 , \26781 , \26782 , \26824 , \26825 , \26787 , \26791 , \26794 , \28087 , \28088 , \28089 , \28090 , \28091 , \28092 , \28093 , \28094 , \28095 , \28096 , \28097 , \28098 , \28099 , \28100 , \28101 , \28102 , \28103 , \28104 , \28105 , \28106 , \28107 , \28108 , \28109 , \28110 , \28111 );
and \U$22409 ( \28113 , \8701 , \28112 );
buf \U$22410 ( \28114 , \26794 );
buf \U$22411 ( \28115 , \26794 );
buf \U$22412 ( \28116 , \26794 );
buf \U$22413 ( \28117 , \26794 );
buf \U$22414 ( \28118 , \26794 );
buf \U$22415 ( \28119 , \26794 );
buf \U$22416 ( \28120 , \26794 );
buf \U$22417 ( \28121 , \26794 );
buf \U$22418 ( \28122 , \26794 );
buf \U$22419 ( \28123 , \26794 );
buf \U$22420 ( \28124 , \26794 );
buf \U$22421 ( \28125 , \26794 );
buf \U$22422 ( \28126 , \26794 );
buf \U$22423 ( \28127 , \26794 );
buf \U$22424 ( \28128 , \26794 );
buf \U$22425 ( \28129 , \26794 );
buf \U$22426 ( \28130 , \26794 );
buf \U$22427 ( \28131 , \26794 );
buf \U$22428 ( \28132 , \26794 );
buf \U$22429 ( \28133 , \26794 );
buf \U$22430 ( \28134 , \26794 );
buf \U$22431 ( \28135 , \26794 );
buf \U$22432 ( \28136 , \26794 );
buf \U$22433 ( \28137 , \26794 );
buf \U$22434 ( \28138 , \26794 );
nor \U$22435 ( \28139 , \26822 , \26823 , \26783 , \26825 , \26787 , \26791 , \26794 , \28114 , \28115 , \28116 , \28117 , \28118 , \28119 , \28120 , \28121 , \28122 , \28123 , \28124 , \28125 , \28126 , \28127 , \28128 , \28129 , \28130 , \28131 , \28132 , \28133 , \28134 , \28135 , \28136 , \28137 , \28138 );
and \U$22436 ( \28140 , \8729 , \28139 );
buf \U$22437 ( \28141 , \26794 );
buf \U$22438 ( \28142 , \26794 );
buf \U$22439 ( \28143 , \26794 );
buf \U$22440 ( \28144 , \26794 );
buf \U$22441 ( \28145 , \26794 );
buf \U$22442 ( \28146 , \26794 );
buf \U$22443 ( \28147 , \26794 );
buf \U$22444 ( \28148 , \26794 );
buf \U$22445 ( \28149 , \26794 );
buf \U$22446 ( \28150 , \26794 );
buf \U$22447 ( \28151 , \26794 );
buf \U$22448 ( \28152 , \26794 );
buf \U$22449 ( \28153 , \26794 );
buf \U$22450 ( \28154 , \26794 );
buf \U$22451 ( \28155 , \26794 );
buf \U$22452 ( \28156 , \26794 );
buf \U$22453 ( \28157 , \26794 );
buf \U$22454 ( \28158 , \26794 );
buf \U$22455 ( \28159 , \26794 );
buf \U$22456 ( \28160 , \26794 );
buf \U$22457 ( \28161 , \26794 );
buf \U$22458 ( \28162 , \26794 );
buf \U$22459 ( \28163 , \26794 );
buf \U$22460 ( \28164 , \26794 );
buf \U$22461 ( \28165 , \26794 );
nor \U$22462 ( \28166 , \26781 , \26823 , \26783 , \26825 , \26787 , \26791 , \26794 , \28141 , \28142 , \28143 , \28144 , \28145 , \28146 , \28147 , \28148 , \28149 , \28150 , \28151 , \28152 , \28153 , \28154 , \28155 , \28156 , \28157 , \28158 , \28159 , \28160 , \28161 , \28162 , \28163 , \28164 , \28165 );
and \U$22463 ( \28167 , \8757 , \28166 );
buf \U$22464 ( \28168 , \26794 );
buf \U$22465 ( \28169 , \26794 );
buf \U$22466 ( \28170 , \26794 );
buf \U$22467 ( \28171 , \26794 );
buf \U$22468 ( \28172 , \26794 );
buf \U$22469 ( \28173 , \26794 );
buf \U$22470 ( \28174 , \26794 );
buf \U$22471 ( \28175 , \26794 );
buf \U$22472 ( \28176 , \26794 );
buf \U$22473 ( \28177 , \26794 );
buf \U$22474 ( \28178 , \26794 );
buf \U$22475 ( \28179 , \26794 );
buf \U$22476 ( \28180 , \26794 );
buf \U$22477 ( \28181 , \26794 );
buf \U$22478 ( \28182 , \26794 );
buf \U$22479 ( \28183 , \26794 );
buf \U$22480 ( \28184 , \26794 );
buf \U$22481 ( \28185 , \26794 );
buf \U$22482 ( \28186 , \26794 );
buf \U$22483 ( \28187 , \26794 );
buf \U$22484 ( \28188 , \26794 );
buf \U$22485 ( \28189 , \26794 );
buf \U$22486 ( \28190 , \26794 );
buf \U$22487 ( \28191 , \26794 );
buf \U$22488 ( \28192 , \26794 );
nor \U$22489 ( \28193 , \26822 , \26782 , \26783 , \26825 , \26787 , \26791 , \26794 , \28168 , \28169 , \28170 , \28171 , \28172 , \28173 , \28174 , \28175 , \28176 , \28177 , \28178 , \28179 , \28180 , \28181 , \28182 , \28183 , \28184 , \28185 , \28186 , \28187 , \28188 , \28189 , \28190 , \28191 , \28192 );
and \U$22490 ( \28194 , \8785 , \28193 );
buf \U$22491 ( \28195 , \26794 );
buf \U$22492 ( \28196 , \26794 );
buf \U$22493 ( \28197 , \26794 );
buf \U$22494 ( \28198 , \26794 );
buf \U$22495 ( \28199 , \26794 );
buf \U$22496 ( \28200 , \26794 );
buf \U$22497 ( \28201 , \26794 );
buf \U$22498 ( \28202 , \26794 );
buf \U$22499 ( \28203 , \26794 );
buf \U$22500 ( \28204 , \26794 );
buf \U$22501 ( \28205 , \26794 );
buf \U$22502 ( \28206 , \26794 );
buf \U$22503 ( \28207 , \26794 );
buf \U$22504 ( \28208 , \26794 );
buf \U$22505 ( \28209 , \26794 );
buf \U$22506 ( \28210 , \26794 );
buf \U$22507 ( \28211 , \26794 );
buf \U$22508 ( \28212 , \26794 );
buf \U$22509 ( \28213 , \26794 );
buf \U$22510 ( \28214 , \26794 );
buf \U$22511 ( \28215 , \26794 );
buf \U$22512 ( \28216 , \26794 );
buf \U$22513 ( \28217 , \26794 );
buf \U$22514 ( \28218 , \26794 );
buf \U$22515 ( \28219 , \26794 );
nor \U$22516 ( \28220 , \26781 , \26782 , \26783 , \26825 , \26787 , \26791 , \26794 , \28195 , \28196 , \28197 , \28198 , \28199 , \28200 , \28201 , \28202 , \28203 , \28204 , \28205 , \28206 , \28207 , \28208 , \28209 , \28210 , \28211 , \28212 , \28213 , \28214 , \28215 , \28216 , \28217 , \28218 , \28219 );
and \U$22517 ( \28221 , \8813 , \28220 );
buf \U$22518 ( \28222 , \26794 );
buf \U$22519 ( \28223 , \26794 );
buf \U$22520 ( \28224 , \26794 );
buf \U$22521 ( \28225 , \26794 );
buf \U$22522 ( \28226 , \26794 );
buf \U$22523 ( \28227 , \26794 );
buf \U$22524 ( \28228 , \26794 );
buf \U$22525 ( \28229 , \26794 );
buf \U$22526 ( \28230 , \26794 );
buf \U$22527 ( \28231 , \26794 );
buf \U$22528 ( \28232 , \26794 );
buf \U$22529 ( \28233 , \26794 );
buf \U$22530 ( \28234 , \26794 );
buf \U$22531 ( \28235 , \26794 );
buf \U$22532 ( \28236 , \26794 );
buf \U$22533 ( \28237 , \26794 );
buf \U$22534 ( \28238 , \26794 );
buf \U$22535 ( \28239 , \26794 );
buf \U$22536 ( \28240 , \26794 );
buf \U$22537 ( \28241 , \26794 );
buf \U$22538 ( \28242 , \26794 );
buf \U$22539 ( \28243 , \26794 );
buf \U$22540 ( \28244 , \26794 );
buf \U$22541 ( \28245 , \26794 );
buf \U$22542 ( \28246 , \26794 );
nor \U$22543 ( \28247 , \26822 , \26823 , \26824 , \26784 , \26787 , \26791 , \26794 , \28222 , \28223 , \28224 , \28225 , \28226 , \28227 , \28228 , \28229 , \28230 , \28231 , \28232 , \28233 , \28234 , \28235 , \28236 , \28237 , \28238 , \28239 , \28240 , \28241 , \28242 , \28243 , \28244 , \28245 , \28246 );
and \U$22544 ( \28248 , \8841 , \28247 );
buf \U$22545 ( \28249 , \26794 );
buf \U$22546 ( \28250 , \26794 );
buf \U$22547 ( \28251 , \26794 );
buf \U$22548 ( \28252 , \26794 );
buf \U$22549 ( \28253 , \26794 );
buf \U$22550 ( \28254 , \26794 );
buf \U$22551 ( \28255 , \26794 );
buf \U$22552 ( \28256 , \26794 );
buf \U$22553 ( \28257 , \26794 );
buf \U$22554 ( \28258 , \26794 );
buf \U$22555 ( \28259 , \26794 );
buf \U$22556 ( \28260 , \26794 );
buf \U$22557 ( \28261 , \26794 );
buf \U$22558 ( \28262 , \26794 );
buf \U$22559 ( \28263 , \26794 );
buf \U$22560 ( \28264 , \26794 );
buf \U$22561 ( \28265 , \26794 );
buf \U$22562 ( \28266 , \26794 );
buf \U$22563 ( \28267 , \26794 );
buf \U$22564 ( \28268 , \26794 );
buf \U$22565 ( \28269 , \26794 );
buf \U$22566 ( \28270 , \26794 );
buf \U$22567 ( \28271 , \26794 );
buf \U$22568 ( \28272 , \26794 );
buf \U$22569 ( \28273 , \26794 );
nor \U$22570 ( \28274 , \26781 , \26823 , \26824 , \26784 , \26787 , \26791 , \26794 , \28249 , \28250 , \28251 , \28252 , \28253 , \28254 , \28255 , \28256 , \28257 , \28258 , \28259 , \28260 , \28261 , \28262 , \28263 , \28264 , \28265 , \28266 , \28267 , \28268 , \28269 , \28270 , \28271 , \28272 , \28273 );
and \U$22571 ( \28275 , \8869 , \28274 );
buf \U$22572 ( \28276 , \26794 );
buf \U$22573 ( \28277 , \26794 );
buf \U$22574 ( \28278 , \26794 );
buf \U$22575 ( \28279 , \26794 );
buf \U$22576 ( \28280 , \26794 );
buf \U$22577 ( \28281 , \26794 );
buf \U$22578 ( \28282 , \26794 );
buf \U$22579 ( \28283 , \26794 );
buf \U$22580 ( \28284 , \26794 );
buf \U$22581 ( \28285 , \26794 );
buf \U$22582 ( \28286 , \26794 );
buf \U$22583 ( \28287 , \26794 );
buf \U$22584 ( \28288 , \26794 );
buf \U$22585 ( \28289 , \26794 );
buf \U$22586 ( \28290 , \26794 );
buf \U$22587 ( \28291 , \26794 );
buf \U$22588 ( \28292 , \26794 );
buf \U$22589 ( \28293 , \26794 );
buf \U$22590 ( \28294 , \26794 );
buf \U$22591 ( \28295 , \26794 );
buf \U$22592 ( \28296 , \26794 );
buf \U$22593 ( \28297 , \26794 );
buf \U$22594 ( \28298 , \26794 );
buf \U$22595 ( \28299 , \26794 );
buf \U$22596 ( \28300 , \26794 );
nor \U$22597 ( \28301 , \26822 , \26782 , \26824 , \26784 , \26787 , \26791 , \26794 , \28276 , \28277 , \28278 , \28279 , \28280 , \28281 , \28282 , \28283 , \28284 , \28285 , \28286 , \28287 , \28288 , \28289 , \28290 , \28291 , \28292 , \28293 , \28294 , \28295 , \28296 , \28297 , \28298 , \28299 , \28300 );
and \U$22598 ( \28302 , \8897 , \28301 );
buf \U$22599 ( \28303 , \26794 );
buf \U$22600 ( \28304 , \26794 );
buf \U$22601 ( \28305 , \26794 );
buf \U$22602 ( \28306 , \26794 );
buf \U$22603 ( \28307 , \26794 );
buf \U$22604 ( \28308 , \26794 );
buf \U$22605 ( \28309 , \26794 );
buf \U$22606 ( \28310 , \26794 );
buf \U$22607 ( \28311 , \26794 );
buf \U$22608 ( \28312 , \26794 );
buf \U$22609 ( \28313 , \26794 );
buf \U$22610 ( \28314 , \26794 );
buf \U$22611 ( \28315 , \26794 );
buf \U$22612 ( \28316 , \26794 );
buf \U$22613 ( \28317 , \26794 );
buf \U$22614 ( \28318 , \26794 );
buf \U$22615 ( \28319 , \26794 );
buf \U$22616 ( \28320 , \26794 );
buf \U$22617 ( \28321 , \26794 );
buf \U$22618 ( \28322 , \26794 );
buf \U$22619 ( \28323 , \26794 );
buf \U$22620 ( \28324 , \26794 );
buf \U$22621 ( \28325 , \26794 );
buf \U$22622 ( \28326 , \26794 );
buf \U$22623 ( \28327 , \26794 );
nor \U$22624 ( \28328 , \26781 , \26782 , \26824 , \26784 , \26787 , \26791 , \26794 , \28303 , \28304 , \28305 , \28306 , \28307 , \28308 , \28309 , \28310 , \28311 , \28312 , \28313 , \28314 , \28315 , \28316 , \28317 , \28318 , \28319 , \28320 , \28321 , \28322 , \28323 , \28324 , \28325 , \28326 , \28327 );
and \U$22625 ( \28329 , \8925 , \28328 );
buf \U$22626 ( \28330 , \26794 );
buf \U$22627 ( \28331 , \26794 );
buf \U$22628 ( \28332 , \26794 );
buf \U$22629 ( \28333 , \26794 );
buf \U$22630 ( \28334 , \26794 );
buf \U$22631 ( \28335 , \26794 );
buf \U$22632 ( \28336 , \26794 );
buf \U$22633 ( \28337 , \26794 );
buf \U$22634 ( \28338 , \26794 );
buf \U$22635 ( \28339 , \26794 );
buf \U$22636 ( \28340 , \26794 );
buf \U$22637 ( \28341 , \26794 );
buf \U$22638 ( \28342 , \26794 );
buf \U$22639 ( \28343 , \26794 );
buf \U$22640 ( \28344 , \26794 );
buf \U$22641 ( \28345 , \26794 );
buf \U$22642 ( \28346 , \26794 );
buf \U$22643 ( \28347 , \26794 );
buf \U$22644 ( \28348 , \26794 );
buf \U$22645 ( \28349 , \26794 );
buf \U$22646 ( \28350 , \26794 );
buf \U$22647 ( \28351 , \26794 );
buf \U$22648 ( \28352 , \26794 );
buf \U$22649 ( \28353 , \26794 );
buf \U$22650 ( \28354 , \26794 );
nor \U$22651 ( \28355 , \26822 , \26823 , \26783 , \26784 , \26787 , \26791 , \26794 , \28330 , \28331 , \28332 , \28333 , \28334 , \28335 , \28336 , \28337 , \28338 , \28339 , \28340 , \28341 , \28342 , \28343 , \28344 , \28345 , \28346 , \28347 , \28348 , \28349 , \28350 , \28351 , \28352 , \28353 , \28354 );
and \U$22652 ( \28356 , \8953 , \28355 );
buf \U$22653 ( \28357 , \26794 );
buf \U$22654 ( \28358 , \26794 );
buf \U$22655 ( \28359 , \26794 );
buf \U$22656 ( \28360 , \26794 );
buf \U$22657 ( \28361 , \26794 );
buf \U$22658 ( \28362 , \26794 );
buf \U$22659 ( \28363 , \26794 );
buf \U$22660 ( \28364 , \26794 );
buf \U$22661 ( \28365 , \26794 );
buf \U$22662 ( \28366 , \26794 );
buf \U$22663 ( \28367 , \26794 );
buf \U$22664 ( \28368 , \26794 );
buf \U$22665 ( \28369 , \26794 );
buf \U$22666 ( \28370 , \26794 );
buf \U$22667 ( \28371 , \26794 );
buf \U$22668 ( \28372 , \26794 );
buf \U$22669 ( \28373 , \26794 );
buf \U$22670 ( \28374 , \26794 );
buf \U$22671 ( \28375 , \26794 );
buf \U$22672 ( \28376 , \26794 );
buf \U$22673 ( \28377 , \26794 );
buf \U$22674 ( \28378 , \26794 );
buf \U$22675 ( \28379 , \26794 );
buf \U$22676 ( \28380 , \26794 );
buf \U$22677 ( \28381 , \26794 );
nor \U$22678 ( \28382 , \26781 , \26823 , \26783 , \26784 , \26787 , \26791 , \26794 , \28357 , \28358 , \28359 , \28360 , \28361 , \28362 , \28363 , \28364 , \28365 , \28366 , \28367 , \28368 , \28369 , \28370 , \28371 , \28372 , \28373 , \28374 , \28375 , \28376 , \28377 , \28378 , \28379 , \28380 , \28381 );
and \U$22679 ( \28383 , \8981 , \28382 );
buf \U$22680 ( \28384 , \26794 );
buf \U$22681 ( \28385 , \26794 );
buf \U$22682 ( \28386 , \26794 );
buf \U$22683 ( \28387 , \26794 );
buf \U$22684 ( \28388 , \26794 );
buf \U$22685 ( \28389 , \26794 );
buf \U$22686 ( \28390 , \26794 );
buf \U$22687 ( \28391 , \26794 );
buf \U$22688 ( \28392 , \26794 );
buf \U$22689 ( \28393 , \26794 );
buf \U$22690 ( \28394 , \26794 );
buf \U$22691 ( \28395 , \26794 );
buf \U$22692 ( \28396 , \26794 );
buf \U$22693 ( \28397 , \26794 );
buf \U$22694 ( \28398 , \26794 );
buf \U$22695 ( \28399 , \26794 );
buf \U$22696 ( \28400 , \26794 );
buf \U$22697 ( \28401 , \26794 );
buf \U$22698 ( \28402 , \26794 );
buf \U$22699 ( \28403 , \26794 );
buf \U$22700 ( \28404 , \26794 );
buf \U$22701 ( \28405 , \26794 );
buf \U$22702 ( \28406 , \26794 );
buf \U$22703 ( \28407 , \26794 );
buf \U$22704 ( \28408 , \26794 );
nor \U$22705 ( \28409 , \26822 , \26782 , \26783 , \26784 , \26787 , \26791 , \26794 , \28384 , \28385 , \28386 , \28387 , \28388 , \28389 , \28390 , \28391 , \28392 , \28393 , \28394 , \28395 , \28396 , \28397 , \28398 , \28399 , \28400 , \28401 , \28402 , \28403 , \28404 , \28405 , \28406 , \28407 , \28408 );
and \U$22706 ( \28410 , \9009 , \28409 );
or \U$22707 ( \28411 , \28005 , \28032 , \28059 , \28086 , \28113 , \28140 , \28167 , \28194 , \28221 , \28248 , \28275 , \28302 , \28329 , \28356 , \28383 , \28410 );
buf \U$22708 ( \28412 , \26794 );
not \U$22709 ( \28413 , \28412 );
buf \U$22710 ( \28414 , \26782 );
buf \U$22711 ( \28415 , \26783 );
buf \U$22712 ( \28416 , \26784 );
buf \U$22713 ( \28417 , \26787 );
buf \U$22714 ( \28418 , \26791 );
buf \U$22715 ( \28419 , \26794 );
buf \U$22716 ( \28420 , \26794 );
buf \U$22717 ( \28421 , \26794 );
buf \U$22718 ( \28422 , \26794 );
buf \U$22719 ( \28423 , \26794 );
buf \U$22720 ( \28424 , \26794 );
buf \U$22721 ( \28425 , \26794 );
buf \U$22722 ( \28426 , \26794 );
buf \U$22723 ( \28427 , \26794 );
buf \U$22724 ( \28428 , \26794 );
buf \U$22725 ( \28429 , \26794 );
buf \U$22726 ( \28430 , \26794 );
buf \U$22727 ( \28431 , \26794 );
buf \U$22728 ( \28432 , \26794 );
buf \U$22729 ( \28433 , \26794 );
buf \U$22730 ( \28434 , \26794 );
buf \U$22731 ( \28435 , \26794 );
buf \U$22732 ( \28436 , \26794 );
buf \U$22733 ( \28437 , \26794 );
buf \U$22734 ( \28438 , \26794 );
buf \U$22735 ( \28439 , \26794 );
buf \U$22736 ( \28440 , \26794 );
buf \U$22737 ( \28441 , \26794 );
buf \U$22738 ( \28442 , \26794 );
buf \U$22739 ( \28443 , \26794 );
buf \U$22740 ( \28444 , \26781 );
or \U$22741 ( \28445 , \28414 , \28415 , \28416 , \28417 , \28418 , \28419 , \28420 , \28421 , \28422 , \28423 , \28424 , \28425 , \28426 , \28427 , \28428 , \28429 , \28430 , \28431 , \28432 , \28433 , \28434 , \28435 , \28436 , \28437 , \28438 , \28439 , \28440 , \28441 , \28442 , \28443 , \28444 );
nand \U$22742 ( \28446 , \28413 , \28445 );
buf \U$22743 ( \28447 , \28446 );
buf \U$22744 ( \28448 , \26794 );
not \U$22745 ( \28449 , \28448 );
buf \U$22746 ( \28450 , \26791 );
buf \U$22747 ( \28451 , \26794 );
buf \U$22748 ( \28452 , \26794 );
buf \U$22749 ( \28453 , \26794 );
buf \U$22750 ( \28454 , \26794 );
buf \U$22751 ( \28455 , \26794 );
buf \U$22752 ( \28456 , \26794 );
buf \U$22753 ( \28457 , \26794 );
buf \U$22754 ( \28458 , \26794 );
buf \U$22755 ( \28459 , \26794 );
buf \U$22756 ( \28460 , \26794 );
buf \U$22757 ( \28461 , \26794 );
buf \U$22758 ( \28462 , \26794 );
buf \U$22759 ( \28463 , \26794 );
buf \U$22760 ( \28464 , \26794 );
buf \U$22761 ( \28465 , \26794 );
buf \U$22762 ( \28466 , \26794 );
buf \U$22763 ( \28467 , \26794 );
buf \U$22764 ( \28468 , \26794 );
buf \U$22765 ( \28469 , \26794 );
buf \U$22766 ( \28470 , \26794 );
buf \U$22767 ( \28471 , \26794 );
buf \U$22768 ( \28472 , \26794 );
buf \U$22769 ( \28473 , \26794 );
buf \U$22770 ( \28474 , \26794 );
buf \U$22771 ( \28475 , \26794 );
buf \U$22772 ( \28476 , \26787 );
buf \U$22773 ( \28477 , \26781 );
buf \U$22774 ( \28478 , \26782 );
buf \U$22775 ( \28479 , \26783 );
buf \U$22776 ( \28480 , \26784 );
or \U$22777 ( \28481 , \28477 , \28478 , \28479 , \28480 );
and \U$22778 ( \28482 , \28476 , \28481 );
or \U$22779 ( \28483 , \28450 , \28451 , \28452 , \28453 , \28454 , \28455 , \28456 , \28457 , \28458 , \28459 , \28460 , \28461 , \28462 , \28463 , \28464 , \28465 , \28466 , \28467 , \28468 , \28469 , \28470 , \28471 , \28472 , \28473 , \28474 , \28475 , \28482 );
and \U$22780 ( \28484 , \28449 , \28483 );
buf \U$22781 ( \28485 , \28484 );
or \U$22782 ( \28486 , \28447 , \28485 );
_DC g8648 ( \28487_nG8648 , \28411 , \28486 );
buf \U$22783 ( \28488 , \28487_nG8648 );
xor \U$22784 ( \28489 , \27978 , \28488 );
buf \U$22785 ( \28490 , RIb7af5b8_255);
and \U$22786 ( \28491 , \7207 , \28004 );
and \U$22787 ( \28492 , \7209 , \28031 );
and \U$22788 ( \28493 , \9119 , \28058 );
and \U$22789 ( \28494 , \9121 , \28085 );
and \U$22790 ( \28495 , \9123 , \28112 );
and \U$22791 ( \28496 , \9125 , \28139 );
and \U$22792 ( \28497 , \9127 , \28166 );
and \U$22793 ( \28498 , \9129 , \28193 );
and \U$22794 ( \28499 , \9131 , \28220 );
and \U$22795 ( \28500 , \9133 , \28247 );
and \U$22796 ( \28501 , \9135 , \28274 );
and \U$22797 ( \28502 , \9137 , \28301 );
and \U$22798 ( \28503 , \9139 , \28328 );
and \U$22799 ( \28504 , \9141 , \28355 );
and \U$22800 ( \28505 , \9143 , \28382 );
and \U$22801 ( \28506 , \9145 , \28409 );
or \U$22802 ( \28507 , \28491 , \28492 , \28493 , \28494 , \28495 , \28496 , \28497 , \28498 , \28499 , \28500 , \28501 , \28502 , \28503 , \28504 , \28505 , \28506 );
_DC g865d ( \28508_nG865d , \28507 , \28486 );
buf \U$22803 ( \28509 , \28508_nG865d );
xor \U$22804 ( \28510 , \28490 , \28509 );
or \U$22805 ( \28511 , \28489 , \28510 );
buf \U$22806 ( \28512 , RIb7af540_256);
and \U$22807 ( \28513 , \7217 , \28004 );
and \U$22808 ( \28514 , \7219 , \28031 );
and \U$22809 ( \28515 , \9155 , \28058 );
and \U$22810 ( \28516 , \9157 , \28085 );
and \U$22811 ( \28517 , \9159 , \28112 );
and \U$22812 ( \28518 , \9161 , \28139 );
and \U$22813 ( \28519 , \9163 , \28166 );
and \U$22814 ( \28520 , \9165 , \28193 );
and \U$22815 ( \28521 , \9167 , \28220 );
and \U$22816 ( \28522 , \9169 , \28247 );
and \U$22817 ( \28523 , \9171 , \28274 );
and \U$22818 ( \28524 , \9173 , \28301 );
and \U$22819 ( \28525 , \9175 , \28328 );
and \U$22820 ( \28526 , \9177 , \28355 );
and \U$22821 ( \28527 , \9179 , \28382 );
and \U$22822 ( \28528 , \9181 , \28409 );
or \U$22823 ( \28529 , \28513 , \28514 , \28515 , \28516 , \28517 , \28518 , \28519 , \28520 , \28521 , \28522 , \28523 , \28524 , \28525 , \28526 , \28527 , \28528 );
_DC g8673 ( \28530_nG8673 , \28529 , \28486 );
buf \U$22824 ( \28531 , \28530_nG8673 );
xor \U$22825 ( \28532 , \28512 , \28531 );
or \U$22826 ( \28533 , \28511 , \28532 );
buf \U$22827 ( \28534 , RIb7af4c8_257);
and \U$22828 ( \28535 , \7227 , \28004 );
and \U$22829 ( \28536 , \7229 , \28031 );
and \U$22830 ( \28537 , \9191 , \28058 );
and \U$22831 ( \28538 , \9193 , \28085 );
and \U$22832 ( \28539 , \9195 , \28112 );
and \U$22833 ( \28540 , \9197 , \28139 );
and \U$22834 ( \28541 , \9199 , \28166 );
and \U$22835 ( \28542 , \9201 , \28193 );
and \U$22836 ( \28543 , \9203 , \28220 );
and \U$22837 ( \28544 , \9205 , \28247 );
and \U$22838 ( \28545 , \9207 , \28274 );
and \U$22839 ( \28546 , \9209 , \28301 );
and \U$22840 ( \28547 , \9211 , \28328 );
and \U$22841 ( \28548 , \9213 , \28355 );
and \U$22842 ( \28549 , \9215 , \28382 );
and \U$22843 ( \28550 , \9217 , \28409 );
or \U$22844 ( \28551 , \28535 , \28536 , \28537 , \28538 , \28539 , \28540 , \28541 , \28542 , \28543 , \28544 , \28545 , \28546 , \28547 , \28548 , \28549 , \28550 );
_DC g8689 ( \28552_nG8689 , \28551 , \28486 );
buf \U$22845 ( \28553 , \28552_nG8689 );
xor \U$22846 ( \28554 , \28534 , \28553 );
or \U$22847 ( \28555 , \28533 , \28554 );
buf \U$22848 ( \28556 , RIb7af450_258);
and \U$22849 ( \28557 , \7237 , \28004 );
and \U$22850 ( \28558 , \7239 , \28031 );
and \U$22851 ( \28559 , \9227 , \28058 );
and \U$22852 ( \28560 , \9229 , \28085 );
and \U$22853 ( \28561 , \9231 , \28112 );
and \U$22854 ( \28562 , \9233 , \28139 );
and \U$22855 ( \28563 , \9235 , \28166 );
and \U$22856 ( \28564 , \9237 , \28193 );
and \U$22857 ( \28565 , \9239 , \28220 );
and \U$22858 ( \28566 , \9241 , \28247 );
and \U$22859 ( \28567 , \9243 , \28274 );
and \U$22860 ( \28568 , \9245 , \28301 );
and \U$22861 ( \28569 , \9247 , \28328 );
and \U$22862 ( \28570 , \9249 , \28355 );
and \U$22863 ( \28571 , \9251 , \28382 );
and \U$22864 ( \28572 , \9253 , \28409 );
or \U$22865 ( \28573 , \28557 , \28558 , \28559 , \28560 , \28561 , \28562 , \28563 , \28564 , \28565 , \28566 , \28567 , \28568 , \28569 , \28570 , \28571 , \28572 );
_DC g869f ( \28574_nG869f , \28573 , \28486 );
buf \U$22866 ( \28575 , \28574_nG869f );
xor \U$22867 ( \28576 , \28556 , \28575 );
or \U$22868 ( \28577 , \28555 , \28576 );
buf \U$22869 ( \28578 , RIb7af3d8_259);
and \U$22870 ( \28579 , \7247 , \28004 );
and \U$22871 ( \28580 , \7249 , \28031 );
and \U$22872 ( \28581 , \9263 , \28058 );
and \U$22873 ( \28582 , \9265 , \28085 );
and \U$22874 ( \28583 , \9267 , \28112 );
and \U$22875 ( \28584 , \9269 , \28139 );
and \U$22876 ( \28585 , \9271 , \28166 );
and \U$22877 ( \28586 , \9273 , \28193 );
and \U$22878 ( \28587 , \9275 , \28220 );
and \U$22879 ( \28588 , \9277 , \28247 );
and \U$22880 ( \28589 , \9279 , \28274 );
and \U$22881 ( \28590 , \9281 , \28301 );
and \U$22882 ( \28591 , \9283 , \28328 );
and \U$22883 ( \28592 , \9285 , \28355 );
and \U$22884 ( \28593 , \9287 , \28382 );
and \U$22885 ( \28594 , \9289 , \28409 );
or \U$22886 ( \28595 , \28579 , \28580 , \28581 , \28582 , \28583 , \28584 , \28585 , \28586 , \28587 , \28588 , \28589 , \28590 , \28591 , \28592 , \28593 , \28594 );
_DC g86b5 ( \28596_nG86b5 , \28595 , \28486 );
buf \U$22887 ( \28597 , \28596_nG86b5 );
xor \U$22888 ( \28598 , \28578 , \28597 );
or \U$22889 ( \28599 , \28577 , \28598 );
buf \U$22890 ( \28600 , RIb7a5bf8_260);
and \U$22891 ( \28601 , \7257 , \28004 );
and \U$22892 ( \28602 , \7259 , \28031 );
and \U$22893 ( \28603 , \9299 , \28058 );
and \U$22894 ( \28604 , \9301 , \28085 );
and \U$22895 ( \28605 , \9303 , \28112 );
and \U$22896 ( \28606 , \9305 , \28139 );
and \U$22897 ( \28607 , \9307 , \28166 );
and \U$22898 ( \28608 , \9309 , \28193 );
and \U$22899 ( \28609 , \9311 , \28220 );
and \U$22900 ( \28610 , \9313 , \28247 );
and \U$22901 ( \28611 , \9315 , \28274 );
and \U$22902 ( \28612 , \9317 , \28301 );
and \U$22903 ( \28613 , \9319 , \28328 );
and \U$22904 ( \28614 , \9321 , \28355 );
and \U$22905 ( \28615 , \9323 , \28382 );
and \U$22906 ( \28616 , \9325 , \28409 );
or \U$22907 ( \28617 , \28601 , \28602 , \28603 , \28604 , \28605 , \28606 , \28607 , \28608 , \28609 , \28610 , \28611 , \28612 , \28613 , \28614 , \28615 , \28616 );
_DC g86cb ( \28618_nG86cb , \28617 , \28486 );
buf \U$22908 ( \28619 , \28618_nG86cb );
xor \U$22909 ( \28620 , \28600 , \28619 );
or \U$22910 ( \28621 , \28599 , \28620 );
buf \U$22911 ( \28622 , RIb7a0c48_261);
and \U$22912 ( \28623 , \7267 , \28004 );
and \U$22913 ( \28624 , \7269 , \28031 );
and \U$22914 ( \28625 , \9335 , \28058 );
and \U$22915 ( \28626 , \9337 , \28085 );
and \U$22916 ( \28627 , \9339 , \28112 );
and \U$22917 ( \28628 , \9341 , \28139 );
and \U$22918 ( \28629 , \9343 , \28166 );
and \U$22919 ( \28630 , \9345 , \28193 );
and \U$22920 ( \28631 , \9347 , \28220 );
and \U$22921 ( \28632 , \9349 , \28247 );
and \U$22922 ( \28633 , \9351 , \28274 );
and \U$22923 ( \28634 , \9353 , \28301 );
and \U$22924 ( \28635 , \9355 , \28328 );
and \U$22925 ( \28636 , \9357 , \28355 );
and \U$22926 ( \28637 , \9359 , \28382 );
and \U$22927 ( \28638 , \9361 , \28409 );
or \U$22928 ( \28639 , \28623 , \28624 , \28625 , \28626 , \28627 , \28628 , \28629 , \28630 , \28631 , \28632 , \28633 , \28634 , \28635 , \28636 , \28637 , \28638 );
_DC g86e1 ( \28640_nG86e1 , \28639 , \28486 );
buf \U$22929 ( \28641 , \28640_nG86e1 );
xor \U$22930 ( \28642 , \28622 , \28641 );
or \U$22931 ( \28643 , \28621 , \28642 );
not \U$22932 ( \28644 , \28643 );
buf \U$22933 ( \28645 , \28644 );
and \U$22934 ( \28646 , \27977 , \28645 );
_HMUX g86e8 ( \28647_nG86e8 , \26444_nG7e44 , \26781 , \28646 );
buf \U$22935 ( \28648 , \26463 );
buf \U$22936 ( \28649 , \26460 );
buf \U$22937 ( \28650 , \26446 );
buf \U$22938 ( \28651 , \26449 );
buf \U$22939 ( \28652 , \26452 );
buf \U$22940 ( \28653 , \26456 );
or \U$22941 ( \28654 , \28650 , \28651 , \28652 , \28653 );
and \U$22942 ( \28655 , \28649 , \28654 );
or \U$22943 ( \28656 , \28648 , \28655 );
buf \U$22944 ( \28657 , \28656 );
_HMUX g86f3 ( \28658_nG86f3 , \26780_nG7f95 , \28647_nG86e8 , \28657 );
buf \U$22945 ( \28659 , RIe5319e0_6884);
not \U$22946 ( \28660 , \28659 );
buf \U$22947 ( \28661 , \28660 );
buf \U$22948 ( \28662 , RIe549ef0_6842);
xor \U$22949 ( \28663 , \28662 , \28659 );
buf \U$22950 ( \28664 , \28663 );
buf \U$22951 ( \28665 , RIe549770_6843);
and \U$22952 ( \28666 , \28662 , \28659 );
xnor \U$22953 ( \28667 , \28665 , \28666 );
buf \U$22954 ( \28668 , \28667 );
buf \U$22955 ( \28669 , RIe548ff0_6844);
or \U$22956 ( \28670 , \28665 , \28666 );
xor \U$22957 ( \28671 , \28669 , \28670 );
buf \U$22958 ( \28672 , \28671 );
buf \U$22959 ( \28673 , RIea91330_6888);
and \U$22960 ( \28674 , \28669 , \28670 );
xor \U$22961 ( \28675 , \28673 , \28674 );
buf \U$22962 ( \28676 , \28675 );
not \U$22963 ( \28677 , \28676 );
and \U$22964 ( \28678 , \28673 , \28674 );
buf \U$22965 ( \28679 , \28678 );
nor \U$22966 ( \28680 , \28661 , \28664 , \28668 , \28672 , \28677 , \28679 );
and \U$22967 ( \28681 , RIe5329d0_6883, \28680 );
not \U$22968 ( \28682 , \28679 );
and \U$22969 ( \28683 , \28661 , \28664 , \28668 , \28672 , \28677 , \28682 );
and \U$22970 ( \28684 , RIeb72150_6905, \28683 );
not \U$22971 ( \28685 , \28661 );
and \U$22972 ( \28686 , \28685 , \28664 , \28668 , \28672 , \28677 , \28682 );
and \U$22973 ( \28687 , RIeab80c0_6897, \28686 );
not \U$22974 ( \28688 , \28664 );
and \U$22975 ( \28689 , \28661 , \28688 , \28668 , \28672 , \28677 , \28682 );
and \U$22976 ( \28690 , RIe5331c8_6882, \28689 );
and \U$22977 ( \28691 , \28685 , \28688 , \28668 , \28672 , \28677 , \28682 );
and \U$22978 ( \28692 , RIe5339c0_6881, \28691 );
not \U$22979 ( \28693 , \28668 );
and \U$22980 ( \28694 , \28661 , \28664 , \28693 , \28672 , \28677 , \28682 );
and \U$22981 ( \28695 , RIeab87c8_6898, \28694 );
and \U$22982 ( \28696 , \28685 , \28664 , \28693 , \28672 , \28677 , \28682 );
and \U$22983 ( \28697 , RIe5341b8_6880, \28696 );
and \U$22984 ( \28698 , \28661 , \28688 , \28693 , \28672 , \28677 , \28682 );
and \U$22985 ( \28699 , RIe5349b0_6879, \28698 );
and \U$22986 ( \28700 , \28685 , \28688 , \28693 , \28672 , \28677 , \28682 );
and \U$22987 ( \28701 , RIea94af8_6890, \28700 );
nor \U$22988 ( \28702 , \28685 , \28688 , \28693 , \28672 , \28676 , \28679 );
and \U$22989 ( \28703 , RIe5351a8_6878, \28702 );
nor \U$22990 ( \28704 , \28661 , \28688 , \28693 , \28672 , \28676 , \28679 );
and \U$22991 ( \28705 , RIe5359a0_6877, \28704 );
nor \U$22992 ( \28706 , \28685 , \28664 , \28693 , \28672 , \28676 , \28679 );
and \U$22993 ( \28707 , RIeab78c8_6895, \28706 );
or \U$22998 ( \28708 , \28681 , \28684 , \28687 , \28690 , \28692 , \28695 , \28697 , \28699 , \28701 , \28703 , \28705 , \28707 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
buf \U$23000 ( \28709 , \28679 );
buf \U$23001 ( \28710 , \28676 );
buf \U$23002 ( \28711 , \28661 );
buf \U$23003 ( \28712 , \28664 );
buf \U$23004 ( \28713 , \28668 );
buf \U$23005 ( \28714 , \28672 );
or \U$23006 ( \28715 , \28711 , \28712 , \28713 , \28714 );
and \U$23007 ( \28716 , \28710 , \28715 );
or \U$23008 ( \28717 , \28709 , \28716 );
buf \U$23009 ( \28718 , \28717 );
or \U$23010 ( \28719 , 1'b0 , \28718 );
_DC g8731 ( \28720_nG8731 , \28708 , \28719 );
not \U$23011 ( \28721 , \28720_nG8731 );
buf \U$23012 ( \28722 , RIb7b9608_246);
and \U$23013 ( \28723 , \7117 , \28680 );
and \U$23014 ( \28724 , \7119 , \28683 );
and \U$23015 ( \28725 , \7864 , \28686 );
and \U$23016 ( \28726 , \7892 , \28689 );
and \U$23017 ( \28727 , \7920 , \28691 );
and \U$23018 ( \28728 , \7948 , \28694 );
and \U$23019 ( \28729 , \7976 , \28696 );
and \U$23020 ( \28730 , \8004 , \28698 );
and \U$23021 ( \28731 , \8032 , \28700 );
and \U$23022 ( \28732 , \8060 , \28702 );
and \U$23023 ( \28733 , \8088 , \28704 );
and \U$23024 ( \28734 , \8116 , \28706 );
or \U$23029 ( \28735 , \28723 , \28724 , \28725 , \28726 , \28727 , \28728 , \28729 , \28730 , \28731 , \28732 , \28733 , \28734 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g8741 ( \28736_nG8741 , \28735 , \28719 );
buf \U$23030 ( \28737 , \28736_nG8741 );
xor \U$23031 ( \28738 , \28722 , \28737 );
buf \U$23032 ( \28739 , RIb7b9590_247);
and \U$23033 ( \28740 , \7126 , \28680 );
and \U$23034 ( \28741 , \7128 , \28683 );
and \U$23035 ( \28742 , \8338 , \28686 );
and \U$23036 ( \28743 , \8340 , \28689 );
and \U$23037 ( \28744 , \8342 , \28691 );
and \U$23038 ( \28745 , \8344 , \28694 );
and \U$23039 ( \28746 , \8346 , \28696 );
and \U$23040 ( \28747 , \8348 , \28698 );
and \U$23041 ( \28748 , \8350 , \28700 );
and \U$23042 ( \28749 , \8352 , \28702 );
and \U$23043 ( \28750 , \8354 , \28704 );
and \U$23044 ( \28751 , \8356 , \28706 );
or \U$23049 ( \28752 , \28740 , \28741 , \28742 , \28743 , \28744 , \28745 , \28746 , \28747 , \28748 , \28749 , \28750 , \28751 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g8752 ( \28753_nG8752 , \28752 , \28719 );
buf \U$23050 ( \28754 , \28753_nG8752 );
xor \U$23051 ( \28755 , \28739 , \28754 );
or \U$23052 ( \28756 , \28738 , \28755 );
buf \U$23053 ( \28757 , RIb7b9518_248);
and \U$23054 ( \28758 , \7136 , \28680 );
and \U$23055 ( \28759 , \7138 , \28683 );
and \U$23056 ( \28760 , \8374 , \28686 );
and \U$23057 ( \28761 , \8376 , \28689 );
and \U$23058 ( \28762 , \8378 , \28691 );
and \U$23059 ( \28763 , \8380 , \28694 );
and \U$23060 ( \28764 , \8382 , \28696 );
and \U$23061 ( \28765 , \8384 , \28698 );
and \U$23062 ( \28766 , \8386 , \28700 );
and \U$23063 ( \28767 , \8388 , \28702 );
and \U$23064 ( \28768 , \8390 , \28704 );
and \U$23065 ( \28769 , \8392 , \28706 );
or \U$23070 ( \28770 , \28758 , \28759 , \28760 , \28761 , \28762 , \28763 , \28764 , \28765 , \28766 , \28767 , \28768 , \28769 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g8764 ( \28771_nG8764 , \28770 , \28719 );
buf \U$23071 ( \28772 , \28771_nG8764 );
xor \U$23072 ( \28773 , \28757 , \28772 );
or \U$23073 ( \28774 , \28756 , \28773 );
buf \U$23074 ( \28775 , RIb7b94a0_249);
and \U$23075 ( \28776 , \7146 , \28680 );
and \U$23076 ( \28777 , \7148 , \28683 );
and \U$23077 ( \28778 , \8410 , \28686 );
and \U$23078 ( \28779 , \8412 , \28689 );
and \U$23079 ( \28780 , \8414 , \28691 );
and \U$23080 ( \28781 , \8416 , \28694 );
and \U$23081 ( \28782 , \8418 , \28696 );
and \U$23082 ( \28783 , \8420 , \28698 );
and \U$23083 ( \28784 , \8422 , \28700 );
and \U$23084 ( \28785 , \8424 , \28702 );
and \U$23085 ( \28786 , \8426 , \28704 );
and \U$23086 ( \28787 , \8428 , \28706 );
or \U$23091 ( \28788 , \28776 , \28777 , \28778 , \28779 , \28780 , \28781 , \28782 , \28783 , \28784 , \28785 , \28786 , \28787 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g8776 ( \28789_nG8776 , \28788 , \28719 );
buf \U$23092 ( \28790 , \28789_nG8776 );
xor \U$23093 ( \28791 , \28775 , \28790 );
or \U$23094 ( \28792 , \28774 , \28791 );
buf \U$23095 ( \28793 , RIb7b9428_250);
and \U$23096 ( \28794 , \7156 , \28680 );
and \U$23097 ( \28795 , \7158 , \28683 );
and \U$23098 ( \28796 , \8446 , \28686 );
and \U$23099 ( \28797 , \8448 , \28689 );
and \U$23100 ( \28798 , \8450 , \28691 );
and \U$23101 ( \28799 , \8452 , \28694 );
and \U$23102 ( \28800 , \8454 , \28696 );
and \U$23103 ( \28801 , \8456 , \28698 );
and \U$23104 ( \28802 , \8458 , \28700 );
and \U$23105 ( \28803 , \8460 , \28702 );
and \U$23106 ( \28804 , \8462 , \28704 );
and \U$23107 ( \28805 , \8464 , \28706 );
or \U$23112 ( \28806 , \28794 , \28795 , \28796 , \28797 , \28798 , \28799 , \28800 , \28801 , \28802 , \28803 , \28804 , \28805 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g8788 ( \28807_nG8788 , \28806 , \28719 );
buf \U$23113 ( \28808 , \28807_nG8788 );
xor \U$23114 ( \28809 , \28793 , \28808 );
or \U$23115 ( \28810 , \28792 , \28809 );
buf \U$23116 ( \28811 , RIb7b93b0_251);
and \U$23117 ( \28812 , \7166 , \28680 );
and \U$23118 ( \28813 , \7168 , \28683 );
and \U$23119 ( \28814 , \8482 , \28686 );
and \U$23120 ( \28815 , \8484 , \28689 );
and \U$23121 ( \28816 , \8486 , \28691 );
and \U$23122 ( \28817 , \8488 , \28694 );
and \U$23123 ( \28818 , \8490 , \28696 );
and \U$23124 ( \28819 , \8492 , \28698 );
and \U$23125 ( \28820 , \8494 , \28700 );
and \U$23126 ( \28821 , \8496 , \28702 );
and \U$23127 ( \28822 , \8498 , \28704 );
and \U$23128 ( \28823 , \8500 , \28706 );
or \U$23133 ( \28824 , \28812 , \28813 , \28814 , \28815 , \28816 , \28817 , \28818 , \28819 , \28820 , \28821 , \28822 , \28823 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g879a ( \28825_nG879a , \28824 , \28719 );
buf \U$23134 ( \28826 , \28825_nG879a );
xor \U$23135 ( \28827 , \28811 , \28826 );
or \U$23136 ( \28828 , \28810 , \28827 );
buf \U$23137 ( \28829 , RIb7af720_252);
and \U$23138 ( \28830 , \7176 , \28680 );
and \U$23139 ( \28831 , \7178 , \28683 );
and \U$23140 ( \28832 , \8518 , \28686 );
and \U$23141 ( \28833 , \8520 , \28689 );
and \U$23142 ( \28834 , \8522 , \28691 );
and \U$23143 ( \28835 , \8524 , \28694 );
and \U$23144 ( \28836 , \8526 , \28696 );
and \U$23145 ( \28837 , \8528 , \28698 );
and \U$23146 ( \28838 , \8530 , \28700 );
and \U$23147 ( \28839 , \8532 , \28702 );
and \U$23148 ( \28840 , \8534 , \28704 );
and \U$23149 ( \28841 , \8536 , \28706 );
or \U$23154 ( \28842 , \28830 , \28831 , \28832 , \28833 , \28834 , \28835 , \28836 , \28837 , \28838 , \28839 , \28840 , \28841 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g87ac ( \28843_nG87ac , \28842 , \28719 );
buf \U$23155 ( \28844 , \28843_nG87ac );
xor \U$23156 ( \28845 , \28829 , \28844 );
or \U$23157 ( \28846 , \28828 , \28845 );
buf \U$23158 ( \28847 , RIb7af6a8_253);
and \U$23159 ( \28848 , \7186 , \28680 );
and \U$23160 ( \28849 , \7188 , \28683 );
and \U$23161 ( \28850 , \8554 , \28686 );
and \U$23162 ( \28851 , \8556 , \28689 );
and \U$23163 ( \28852 , \8558 , \28691 );
and \U$23164 ( \28853 , \8560 , \28694 );
and \U$23165 ( \28854 , \8562 , \28696 );
and \U$23166 ( \28855 , \8564 , \28698 );
and \U$23167 ( \28856 , \8566 , \28700 );
and \U$23168 ( \28857 , \8568 , \28702 );
and \U$23169 ( \28858 , \8570 , \28704 );
and \U$23170 ( \28859 , \8572 , \28706 );
or \U$23175 ( \28860 , \28848 , \28849 , \28850 , \28851 , \28852 , \28853 , \28854 , \28855 , \28856 , \28857 , \28858 , \28859 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g87be ( \28861_nG87be , \28860 , \28719 );
buf \U$23176 ( \28862 , \28861_nG87be );
xor \U$23177 ( \28863 , \28847 , \28862 );
or \U$23178 ( \28864 , \28846 , \28863 );
not \U$23179 ( \28865 , \28864 );
buf \U$23180 ( \28866 , \28865 );
buf \U$23181 ( \28867 , RIb7af630_254);
and \U$23182 ( \28868 , \7198 , \28680 );
and \U$23183 ( \28869 , \7200 , \28683 );
and \U$23184 ( \28870 , \8645 , \28686 );
and \U$23185 ( \28871 , \8673 , \28689 );
and \U$23186 ( \28872 , \8701 , \28691 );
and \U$23187 ( \28873 , \8729 , \28694 );
and \U$23188 ( \28874 , \8757 , \28696 );
and \U$23189 ( \28875 , \8785 , \28698 );
and \U$23190 ( \28876 , \8813 , \28700 );
and \U$23191 ( \28877 , \8841 , \28702 );
and \U$23192 ( \28878 , \8869 , \28704 );
and \U$23193 ( \28879 , \8897 , \28706 );
or \U$23198 ( \28880 , \28868 , \28869 , \28870 , \28871 , \28872 , \28873 , \28874 , \28875 , \28876 , \28877 , \28878 , \28879 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g87d2 ( \28881_nG87d2 , \28880 , \28719 );
buf \U$23199 ( \28882 , \28881_nG87d2 );
xor \U$23200 ( \28883 , \28867 , \28882 );
buf \U$23201 ( \28884 , RIb7af5b8_255);
and \U$23202 ( \28885 , \7207 , \28680 );
and \U$23203 ( \28886 , \7209 , \28683 );
and \U$23204 ( \28887 , \9119 , \28686 );
and \U$23205 ( \28888 , \9121 , \28689 );
and \U$23206 ( \28889 , \9123 , \28691 );
and \U$23207 ( \28890 , \9125 , \28694 );
and \U$23208 ( \28891 , \9127 , \28696 );
and \U$23209 ( \28892 , \9129 , \28698 );
and \U$23210 ( \28893 , \9131 , \28700 );
and \U$23211 ( \28894 , \9133 , \28702 );
and \U$23212 ( \28895 , \9135 , \28704 );
and \U$23213 ( \28896 , \9137 , \28706 );
or \U$23218 ( \28897 , \28885 , \28886 , \28887 , \28888 , \28889 , \28890 , \28891 , \28892 , \28893 , \28894 , \28895 , \28896 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g87e3 ( \28898_nG87e3 , \28897 , \28719 );
buf \U$23219 ( \28899 , \28898_nG87e3 );
xor \U$23220 ( \28900 , \28884 , \28899 );
or \U$23221 ( \28901 , \28883 , \28900 );
buf \U$23222 ( \28902 , RIb7af540_256);
and \U$23223 ( \28903 , \7217 , \28680 );
and \U$23224 ( \28904 , \7219 , \28683 );
and \U$23225 ( \28905 , \9155 , \28686 );
and \U$23226 ( \28906 , \9157 , \28689 );
and \U$23227 ( \28907 , \9159 , \28691 );
and \U$23228 ( \28908 , \9161 , \28694 );
and \U$23229 ( \28909 , \9163 , \28696 );
and \U$23230 ( \28910 , \9165 , \28698 );
and \U$23231 ( \28911 , \9167 , \28700 );
and \U$23232 ( \28912 , \9169 , \28702 );
and \U$23233 ( \28913 , \9171 , \28704 );
and \U$23234 ( \28914 , \9173 , \28706 );
or \U$23239 ( \28915 , \28903 , \28904 , \28905 , \28906 , \28907 , \28908 , \28909 , \28910 , \28911 , \28912 , \28913 , \28914 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g87f5 ( \28916_nG87f5 , \28915 , \28719 );
buf \U$23240 ( \28917 , \28916_nG87f5 );
xor \U$23241 ( \28918 , \28902 , \28917 );
or \U$23242 ( \28919 , \28901 , \28918 );
buf \U$23243 ( \28920 , RIb7af4c8_257);
and \U$23244 ( \28921 , \7227 , \28680 );
and \U$23245 ( \28922 , \7229 , \28683 );
and \U$23246 ( \28923 , \9191 , \28686 );
and \U$23247 ( \28924 , \9193 , \28689 );
and \U$23248 ( \28925 , \9195 , \28691 );
and \U$23249 ( \28926 , \9197 , \28694 );
and \U$23250 ( \28927 , \9199 , \28696 );
and \U$23251 ( \28928 , \9201 , \28698 );
and \U$23252 ( \28929 , \9203 , \28700 );
and \U$23253 ( \28930 , \9205 , \28702 );
and \U$23254 ( \28931 , \9207 , \28704 );
and \U$23255 ( \28932 , \9209 , \28706 );
or \U$23260 ( \28933 , \28921 , \28922 , \28923 , \28924 , \28925 , \28926 , \28927 , \28928 , \28929 , \28930 , \28931 , \28932 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g8807 ( \28934_nG8807 , \28933 , \28719 );
buf \U$23261 ( \28935 , \28934_nG8807 );
xor \U$23262 ( \28936 , \28920 , \28935 );
or \U$23263 ( \28937 , \28919 , \28936 );
buf \U$23264 ( \28938 , RIb7af450_258);
and \U$23265 ( \28939 , \7237 , \28680 );
and \U$23266 ( \28940 , \7239 , \28683 );
and \U$23267 ( \28941 , \9227 , \28686 );
and \U$23268 ( \28942 , \9229 , \28689 );
and \U$23269 ( \28943 , \9231 , \28691 );
and \U$23270 ( \28944 , \9233 , \28694 );
and \U$23271 ( \28945 , \9235 , \28696 );
and \U$23272 ( \28946 , \9237 , \28698 );
and \U$23273 ( \28947 , \9239 , \28700 );
and \U$23274 ( \28948 , \9241 , \28702 );
and \U$23275 ( \28949 , \9243 , \28704 );
and \U$23276 ( \28950 , \9245 , \28706 );
or \U$23281 ( \28951 , \28939 , \28940 , \28941 , \28942 , \28943 , \28944 , \28945 , \28946 , \28947 , \28948 , \28949 , \28950 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g8819 ( \28952_nG8819 , \28951 , \28719 );
buf \U$23282 ( \28953 , \28952_nG8819 );
xor \U$23283 ( \28954 , \28938 , \28953 );
or \U$23284 ( \28955 , \28937 , \28954 );
buf \U$23285 ( \28956 , RIb7af3d8_259);
and \U$23286 ( \28957 , \7247 , \28680 );
and \U$23287 ( \28958 , \7249 , \28683 );
and \U$23288 ( \28959 , \9263 , \28686 );
and \U$23289 ( \28960 , \9265 , \28689 );
and \U$23290 ( \28961 , \9267 , \28691 );
and \U$23291 ( \28962 , \9269 , \28694 );
and \U$23292 ( \28963 , \9271 , \28696 );
and \U$23293 ( \28964 , \9273 , \28698 );
and \U$23294 ( \28965 , \9275 , \28700 );
and \U$23295 ( \28966 , \9277 , \28702 );
and \U$23296 ( \28967 , \9279 , \28704 );
and \U$23297 ( \28968 , \9281 , \28706 );
or \U$23302 ( \28969 , \28957 , \28958 , \28959 , \28960 , \28961 , \28962 , \28963 , \28964 , \28965 , \28966 , \28967 , \28968 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g882b ( \28970_nG882b , \28969 , \28719 );
buf \U$23303 ( \28971 , \28970_nG882b );
xor \U$23304 ( \28972 , \28956 , \28971 );
or \U$23305 ( \28973 , \28955 , \28972 );
buf \U$23306 ( \28974 , RIb7a5bf8_260);
and \U$23307 ( \28975 , \7257 , \28680 );
and \U$23308 ( \28976 , \7259 , \28683 );
and \U$23309 ( \28977 , \9299 , \28686 );
and \U$23310 ( \28978 , \9301 , \28689 );
and \U$23311 ( \28979 , \9303 , \28691 );
and \U$23312 ( \28980 , \9305 , \28694 );
and \U$23313 ( \28981 , \9307 , \28696 );
and \U$23314 ( \28982 , \9309 , \28698 );
and \U$23315 ( \28983 , \9311 , \28700 );
and \U$23316 ( \28984 , \9313 , \28702 );
and \U$23317 ( \28985 , \9315 , \28704 );
and \U$23318 ( \28986 , \9317 , \28706 );
or \U$23323 ( \28987 , \28975 , \28976 , \28977 , \28978 , \28979 , \28980 , \28981 , \28982 , \28983 , \28984 , \28985 , \28986 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g883d ( \28988_nG883d , \28987 , \28719 );
buf \U$23324 ( \28989 , \28988_nG883d );
xor \U$23325 ( \28990 , \28974 , \28989 );
or \U$23326 ( \28991 , \28973 , \28990 );
buf \U$23327 ( \28992 , RIb7a0c48_261);
and \U$23328 ( \28993 , \7267 , \28680 );
and \U$23329 ( \28994 , \7269 , \28683 );
and \U$23330 ( \28995 , \9335 , \28686 );
and \U$23331 ( \28996 , \9337 , \28689 );
and \U$23332 ( \28997 , \9339 , \28691 );
and \U$23333 ( \28998 , \9341 , \28694 );
and \U$23334 ( \28999 , \9343 , \28696 );
and \U$23335 ( \29000 , \9345 , \28698 );
and \U$23336 ( \29001 , \9347 , \28700 );
and \U$23337 ( \29002 , \9349 , \28702 );
and \U$23338 ( \29003 , \9351 , \28704 );
and \U$23339 ( \29004 , \9353 , \28706 );
or \U$23344 ( \29005 , \28993 , \28994 , \28995 , \28996 , \28997 , \28998 , \28999 , \29000 , \29001 , \29002 , \29003 , \29004 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
_DC g884f ( \29006_nG884f , \29005 , \28719 );
buf \U$23345 ( \29007 , \29006_nG884f );
xor \U$23346 ( \29008 , \28992 , \29007 );
or \U$23347 ( \29009 , \28991 , \29008 );
not \U$23348 ( \29010 , \29009 );
buf \U$23349 ( \29011 , \29010 );
and \U$23350 ( \29012 , \28866 , \29011 );
and \U$23351 ( \29013 , \28721 , \29012 );
_HMUX g8857 ( \29014_nG8857 , \28658_nG86f3 , \28661 , \29013 );
buf \U$23354 ( \29015 , \28661 );
buf \U$23357 ( \29016 , \28664 );
buf \U$23360 ( \29017 , \28668 );
buf \U$23363 ( \29018 , \28672 );
buf \U$23364 ( \29019 , \28676 );
not \U$23365 ( \29020 , \29019 );
buf \U$23366 ( \29021 , \29020 );
not \U$23367 ( \29022 , \29021 );
buf \U$23368 ( \29023 , \28679 );
xnor \U$23369 ( \29024 , \29023 , \29019 );
buf \U$23370 ( \29025 , \29024 );
or \U$23371 ( \29026 , \29023 , \29019 );
not \U$23372 ( \29027 , \29026 );
buf \U$23373 ( \29028 , \29027 );
buf \U$23374 ( \29029 , \29028 );
buf \U$23375 ( \29030 , \29028 );
buf \U$23376 ( \29031 , \29028 );
buf \U$23377 ( \29032 , \29028 );
buf \U$23378 ( \29033 , \29028 );
buf \U$23379 ( \29034 , \29028 );
buf \U$23380 ( \29035 , \29028 );
buf \U$23381 ( \29036 , \29028 );
buf \U$23382 ( \29037 , \29028 );
buf \U$23383 ( \29038 , \29028 );
buf \U$23384 ( \29039 , \29028 );
buf \U$23385 ( \29040 , \29028 );
buf \U$23386 ( \29041 , \29028 );
buf \U$23387 ( \29042 , \29028 );
buf \U$23388 ( \29043 , \29028 );
buf \U$23389 ( \29044 , \29028 );
buf \U$23390 ( \29045 , \29028 );
buf \U$23391 ( \29046 , \29028 );
buf \U$23392 ( \29047 , \29028 );
buf \U$23393 ( \29048 , \29028 );
buf \U$23394 ( \29049 , \29028 );
buf \U$23395 ( \29050 , \29028 );
buf \U$23396 ( \29051 , \29028 );
buf \U$23397 ( \29052 , \29028 );
buf \U$23398 ( \29053 , \29028 );
nor \U$23399 ( \29054 , \29015 , \29016 , \29017 , \29018 , \29022 , \29025 , \29028 , \29029 , \29030 , \29031 , \29032 , \29033 , \29034 , \29035 , \29036 , \29037 , \29038 , \29039 , \29040 , \29041 , \29042 , \29043 , \29044 , \29045 , \29046 , \29047 , \29048 , \29049 , \29050 , \29051 , \29052 , \29053 );
and \U$23400 ( \29055 , RIe5329d0_6883, \29054 );
not \U$23401 ( \29056 , \29015 );
not \U$23402 ( \29057 , \29016 );
not \U$23403 ( \29058 , \29017 );
not \U$23404 ( \29059 , \29018 );
buf \U$23405 ( \29060 , \29028 );
buf \U$23406 ( \29061 , \29028 );
buf \U$23407 ( \29062 , \29028 );
buf \U$23408 ( \29063 , \29028 );
buf \U$23409 ( \29064 , \29028 );
buf \U$23410 ( \29065 , \29028 );
buf \U$23411 ( \29066 , \29028 );
buf \U$23412 ( \29067 , \29028 );
buf \U$23413 ( \29068 , \29028 );
buf \U$23414 ( \29069 , \29028 );
buf \U$23415 ( \29070 , \29028 );
buf \U$23416 ( \29071 , \29028 );
buf \U$23417 ( \29072 , \29028 );
buf \U$23418 ( \29073 , \29028 );
buf \U$23419 ( \29074 , \29028 );
buf \U$23420 ( \29075 , \29028 );
buf \U$23421 ( \29076 , \29028 );
buf \U$23422 ( \29077 , \29028 );
buf \U$23423 ( \29078 , \29028 );
buf \U$23424 ( \29079 , \29028 );
buf \U$23425 ( \29080 , \29028 );
buf \U$23426 ( \29081 , \29028 );
buf \U$23427 ( \29082 , \29028 );
buf \U$23428 ( \29083 , \29028 );
buf \U$23429 ( \29084 , \29028 );
nor \U$23430 ( \29085 , \29056 , \29057 , \29058 , \29059 , \29021 , \29025 , \29028 , \29060 , \29061 , \29062 , \29063 , \29064 , \29065 , \29066 , \29067 , \29068 , \29069 , \29070 , \29071 , \29072 , \29073 , \29074 , \29075 , \29076 , \29077 , \29078 , \29079 , \29080 , \29081 , \29082 , \29083 , \29084 );
and \U$23431 ( \29086 , RIeb72150_6905, \29085 );
buf \U$23432 ( \29087 , \29028 );
buf \U$23433 ( \29088 , \29028 );
buf \U$23434 ( \29089 , \29028 );
buf \U$23435 ( \29090 , \29028 );
buf \U$23436 ( \29091 , \29028 );
buf \U$23437 ( \29092 , \29028 );
buf \U$23438 ( \29093 , \29028 );
buf \U$23439 ( \29094 , \29028 );
buf \U$23440 ( \29095 , \29028 );
buf \U$23441 ( \29096 , \29028 );
buf \U$23442 ( \29097 , \29028 );
buf \U$23443 ( \29098 , \29028 );
buf \U$23444 ( \29099 , \29028 );
buf \U$23445 ( \29100 , \29028 );
buf \U$23446 ( \29101 , \29028 );
buf \U$23447 ( \29102 , \29028 );
buf \U$23448 ( \29103 , \29028 );
buf \U$23449 ( \29104 , \29028 );
buf \U$23450 ( \29105 , \29028 );
buf \U$23451 ( \29106 , \29028 );
buf \U$23452 ( \29107 , \29028 );
buf \U$23453 ( \29108 , \29028 );
buf \U$23454 ( \29109 , \29028 );
buf \U$23455 ( \29110 , \29028 );
buf \U$23456 ( \29111 , \29028 );
nor \U$23457 ( \29112 , \29015 , \29057 , \29058 , \29059 , \29021 , \29025 , \29028 , \29087 , \29088 , \29089 , \29090 , \29091 , \29092 , \29093 , \29094 , \29095 , \29096 , \29097 , \29098 , \29099 , \29100 , \29101 , \29102 , \29103 , \29104 , \29105 , \29106 , \29107 , \29108 , \29109 , \29110 , \29111 );
and \U$23458 ( \29113 , RIeab80c0_6897, \29112 );
buf \U$23459 ( \29114 , \29028 );
buf \U$23460 ( \29115 , \29028 );
buf \U$23461 ( \29116 , \29028 );
buf \U$23462 ( \29117 , \29028 );
buf \U$23463 ( \29118 , \29028 );
buf \U$23464 ( \29119 , \29028 );
buf \U$23465 ( \29120 , \29028 );
buf \U$23466 ( \29121 , \29028 );
buf \U$23467 ( \29122 , \29028 );
buf \U$23468 ( \29123 , \29028 );
buf \U$23469 ( \29124 , \29028 );
buf \U$23470 ( \29125 , \29028 );
buf \U$23471 ( \29126 , \29028 );
buf \U$23472 ( \29127 , \29028 );
buf \U$23473 ( \29128 , \29028 );
buf \U$23474 ( \29129 , \29028 );
buf \U$23475 ( \29130 , \29028 );
buf \U$23476 ( \29131 , \29028 );
buf \U$23477 ( \29132 , \29028 );
buf \U$23478 ( \29133 , \29028 );
buf \U$23479 ( \29134 , \29028 );
buf \U$23480 ( \29135 , \29028 );
buf \U$23481 ( \29136 , \29028 );
buf \U$23482 ( \29137 , \29028 );
buf \U$23483 ( \29138 , \29028 );
nor \U$23484 ( \29139 , \29056 , \29016 , \29058 , \29059 , \29021 , \29025 , \29028 , \29114 , \29115 , \29116 , \29117 , \29118 , \29119 , \29120 , \29121 , \29122 , \29123 , \29124 , \29125 , \29126 , \29127 , \29128 , \29129 , \29130 , \29131 , \29132 , \29133 , \29134 , \29135 , \29136 , \29137 , \29138 );
and \U$23485 ( \29140 , RIe5331c8_6882, \29139 );
buf \U$23486 ( \29141 , \29028 );
buf \U$23487 ( \29142 , \29028 );
buf \U$23488 ( \29143 , \29028 );
buf \U$23489 ( \29144 , \29028 );
buf \U$23490 ( \29145 , \29028 );
buf \U$23491 ( \29146 , \29028 );
buf \U$23492 ( \29147 , \29028 );
buf \U$23493 ( \29148 , \29028 );
buf \U$23494 ( \29149 , \29028 );
buf \U$23495 ( \29150 , \29028 );
buf \U$23496 ( \29151 , \29028 );
buf \U$23497 ( \29152 , \29028 );
buf \U$23498 ( \29153 , \29028 );
buf \U$23499 ( \29154 , \29028 );
buf \U$23500 ( \29155 , \29028 );
buf \U$23501 ( \29156 , \29028 );
buf \U$23502 ( \29157 , \29028 );
buf \U$23503 ( \29158 , \29028 );
buf \U$23504 ( \29159 , \29028 );
buf \U$23505 ( \29160 , \29028 );
buf \U$23506 ( \29161 , \29028 );
buf \U$23507 ( \29162 , \29028 );
buf \U$23508 ( \29163 , \29028 );
buf \U$23509 ( \29164 , \29028 );
buf \U$23510 ( \29165 , \29028 );
nor \U$23511 ( \29166 , \29015 , \29016 , \29058 , \29059 , \29021 , \29025 , \29028 , \29141 , \29142 , \29143 , \29144 , \29145 , \29146 , \29147 , \29148 , \29149 , \29150 , \29151 , \29152 , \29153 , \29154 , \29155 , \29156 , \29157 , \29158 , \29159 , \29160 , \29161 , \29162 , \29163 , \29164 , \29165 );
and \U$23512 ( \29167 , RIe5339c0_6881, \29166 );
buf \U$23513 ( \29168 , \29028 );
buf \U$23514 ( \29169 , \29028 );
buf \U$23515 ( \29170 , \29028 );
buf \U$23516 ( \29171 , \29028 );
buf \U$23517 ( \29172 , \29028 );
buf \U$23518 ( \29173 , \29028 );
buf \U$23519 ( \29174 , \29028 );
buf \U$23520 ( \29175 , \29028 );
buf \U$23521 ( \29176 , \29028 );
buf \U$23522 ( \29177 , \29028 );
buf \U$23523 ( \29178 , \29028 );
buf \U$23524 ( \29179 , \29028 );
buf \U$23525 ( \29180 , \29028 );
buf \U$23526 ( \29181 , \29028 );
buf \U$23527 ( \29182 , \29028 );
buf \U$23528 ( \29183 , \29028 );
buf \U$23529 ( \29184 , \29028 );
buf \U$23530 ( \29185 , \29028 );
buf \U$23531 ( \29186 , \29028 );
buf \U$23532 ( \29187 , \29028 );
buf \U$23533 ( \29188 , \29028 );
buf \U$23534 ( \29189 , \29028 );
buf \U$23535 ( \29190 , \29028 );
buf \U$23536 ( \29191 , \29028 );
buf \U$23537 ( \29192 , \29028 );
nor \U$23538 ( \29193 , \29056 , \29057 , \29017 , \29059 , \29021 , \29025 , \29028 , \29168 , \29169 , \29170 , \29171 , \29172 , \29173 , \29174 , \29175 , \29176 , \29177 , \29178 , \29179 , \29180 , \29181 , \29182 , \29183 , \29184 , \29185 , \29186 , \29187 , \29188 , \29189 , \29190 , \29191 , \29192 );
and \U$23539 ( \29194 , RIeab87c8_6898, \29193 );
buf \U$23540 ( \29195 , \29028 );
buf \U$23541 ( \29196 , \29028 );
buf \U$23542 ( \29197 , \29028 );
buf \U$23543 ( \29198 , \29028 );
buf \U$23544 ( \29199 , \29028 );
buf \U$23545 ( \29200 , \29028 );
buf \U$23546 ( \29201 , \29028 );
buf \U$23547 ( \29202 , \29028 );
buf \U$23548 ( \29203 , \29028 );
buf \U$23549 ( \29204 , \29028 );
buf \U$23550 ( \29205 , \29028 );
buf \U$23551 ( \29206 , \29028 );
buf \U$23552 ( \29207 , \29028 );
buf \U$23553 ( \29208 , \29028 );
buf \U$23554 ( \29209 , \29028 );
buf \U$23555 ( \29210 , \29028 );
buf \U$23556 ( \29211 , \29028 );
buf \U$23557 ( \29212 , \29028 );
buf \U$23558 ( \29213 , \29028 );
buf \U$23559 ( \29214 , \29028 );
buf \U$23560 ( \29215 , \29028 );
buf \U$23561 ( \29216 , \29028 );
buf \U$23562 ( \29217 , \29028 );
buf \U$23563 ( \29218 , \29028 );
buf \U$23564 ( \29219 , \29028 );
nor \U$23565 ( \29220 , \29015 , \29057 , \29017 , \29059 , \29021 , \29025 , \29028 , \29195 , \29196 , \29197 , \29198 , \29199 , \29200 , \29201 , \29202 , \29203 , \29204 , \29205 , \29206 , \29207 , \29208 , \29209 , \29210 , \29211 , \29212 , \29213 , \29214 , \29215 , \29216 , \29217 , \29218 , \29219 );
and \U$23566 ( \29221 , RIe5341b8_6880, \29220 );
buf \U$23567 ( \29222 , \29028 );
buf \U$23568 ( \29223 , \29028 );
buf \U$23569 ( \29224 , \29028 );
buf \U$23570 ( \29225 , \29028 );
buf \U$23571 ( \29226 , \29028 );
buf \U$23572 ( \29227 , \29028 );
buf \U$23573 ( \29228 , \29028 );
buf \U$23574 ( \29229 , \29028 );
buf \U$23575 ( \29230 , \29028 );
buf \U$23576 ( \29231 , \29028 );
buf \U$23577 ( \29232 , \29028 );
buf \U$23578 ( \29233 , \29028 );
buf \U$23579 ( \29234 , \29028 );
buf \U$23580 ( \29235 , \29028 );
buf \U$23581 ( \29236 , \29028 );
buf \U$23582 ( \29237 , \29028 );
buf \U$23583 ( \29238 , \29028 );
buf \U$23584 ( \29239 , \29028 );
buf \U$23585 ( \29240 , \29028 );
buf \U$23586 ( \29241 , \29028 );
buf \U$23587 ( \29242 , \29028 );
buf \U$23588 ( \29243 , \29028 );
buf \U$23589 ( \29244 , \29028 );
buf \U$23590 ( \29245 , \29028 );
buf \U$23591 ( \29246 , \29028 );
nor \U$23592 ( \29247 , \29056 , \29016 , \29017 , \29059 , \29021 , \29025 , \29028 , \29222 , \29223 , \29224 , \29225 , \29226 , \29227 , \29228 , \29229 , \29230 , \29231 , \29232 , \29233 , \29234 , \29235 , \29236 , \29237 , \29238 , \29239 , \29240 , \29241 , \29242 , \29243 , \29244 , \29245 , \29246 );
and \U$23593 ( \29248 , RIe5349b0_6879, \29247 );
buf \U$23594 ( \29249 , \29028 );
buf \U$23595 ( \29250 , \29028 );
buf \U$23596 ( \29251 , \29028 );
buf \U$23597 ( \29252 , \29028 );
buf \U$23598 ( \29253 , \29028 );
buf \U$23599 ( \29254 , \29028 );
buf \U$23600 ( \29255 , \29028 );
buf \U$23601 ( \29256 , \29028 );
buf \U$23602 ( \29257 , \29028 );
buf \U$23603 ( \29258 , \29028 );
buf \U$23604 ( \29259 , \29028 );
buf \U$23605 ( \29260 , \29028 );
buf \U$23606 ( \29261 , \29028 );
buf \U$23607 ( \29262 , \29028 );
buf \U$23608 ( \29263 , \29028 );
buf \U$23609 ( \29264 , \29028 );
buf \U$23610 ( \29265 , \29028 );
buf \U$23611 ( \29266 , \29028 );
buf \U$23612 ( \29267 , \29028 );
buf \U$23613 ( \29268 , \29028 );
buf \U$23614 ( \29269 , \29028 );
buf \U$23615 ( \29270 , \29028 );
buf \U$23616 ( \29271 , \29028 );
buf \U$23617 ( \29272 , \29028 );
buf \U$23618 ( \29273 , \29028 );
nor \U$23619 ( \29274 , \29015 , \29016 , \29017 , \29059 , \29021 , \29025 , \29028 , \29249 , \29250 , \29251 , \29252 , \29253 , \29254 , \29255 , \29256 , \29257 , \29258 , \29259 , \29260 , \29261 , \29262 , \29263 , \29264 , \29265 , \29266 , \29267 , \29268 , \29269 , \29270 , \29271 , \29272 , \29273 );
and \U$23620 ( \29275 , RIea94af8_6890, \29274 );
buf \U$23621 ( \29276 , \29028 );
buf \U$23622 ( \29277 , \29028 );
buf \U$23623 ( \29278 , \29028 );
buf \U$23624 ( \29279 , \29028 );
buf \U$23625 ( \29280 , \29028 );
buf \U$23626 ( \29281 , \29028 );
buf \U$23627 ( \29282 , \29028 );
buf \U$23628 ( \29283 , \29028 );
buf \U$23629 ( \29284 , \29028 );
buf \U$23630 ( \29285 , \29028 );
buf \U$23631 ( \29286 , \29028 );
buf \U$23632 ( \29287 , \29028 );
buf \U$23633 ( \29288 , \29028 );
buf \U$23634 ( \29289 , \29028 );
buf \U$23635 ( \29290 , \29028 );
buf \U$23636 ( \29291 , \29028 );
buf \U$23637 ( \29292 , \29028 );
buf \U$23638 ( \29293 , \29028 );
buf \U$23639 ( \29294 , \29028 );
buf \U$23640 ( \29295 , \29028 );
buf \U$23641 ( \29296 , \29028 );
buf \U$23642 ( \29297 , \29028 );
buf \U$23643 ( \29298 , \29028 );
buf \U$23644 ( \29299 , \29028 );
buf \U$23645 ( \29300 , \29028 );
nor \U$23646 ( \29301 , \29056 , \29057 , \29058 , \29018 , \29021 , \29025 , \29028 , \29276 , \29277 , \29278 , \29279 , \29280 , \29281 , \29282 , \29283 , \29284 , \29285 , \29286 , \29287 , \29288 , \29289 , \29290 , \29291 , \29292 , \29293 , \29294 , \29295 , \29296 , \29297 , \29298 , \29299 , \29300 );
and \U$23647 ( \29302 , RIe5351a8_6878, \29301 );
buf \U$23648 ( \29303 , \29028 );
buf \U$23649 ( \29304 , \29028 );
buf \U$23650 ( \29305 , \29028 );
buf \U$23651 ( \29306 , \29028 );
buf \U$23652 ( \29307 , \29028 );
buf \U$23653 ( \29308 , \29028 );
buf \U$23654 ( \29309 , \29028 );
buf \U$23655 ( \29310 , \29028 );
buf \U$23656 ( \29311 , \29028 );
buf \U$23657 ( \29312 , \29028 );
buf \U$23658 ( \29313 , \29028 );
buf \U$23659 ( \29314 , \29028 );
buf \U$23660 ( \29315 , \29028 );
buf \U$23661 ( \29316 , \29028 );
buf \U$23662 ( \29317 , \29028 );
buf \U$23663 ( \29318 , \29028 );
buf \U$23664 ( \29319 , \29028 );
buf \U$23665 ( \29320 , \29028 );
buf \U$23666 ( \29321 , \29028 );
buf \U$23667 ( \29322 , \29028 );
buf \U$23668 ( \29323 , \29028 );
buf \U$23669 ( \29324 , \29028 );
buf \U$23670 ( \29325 , \29028 );
buf \U$23671 ( \29326 , \29028 );
buf \U$23672 ( \29327 , \29028 );
nor \U$23673 ( \29328 , \29015 , \29057 , \29058 , \29018 , \29021 , \29025 , \29028 , \29303 , \29304 , \29305 , \29306 , \29307 , \29308 , \29309 , \29310 , \29311 , \29312 , \29313 , \29314 , \29315 , \29316 , \29317 , \29318 , \29319 , \29320 , \29321 , \29322 , \29323 , \29324 , \29325 , \29326 , \29327 );
and \U$23674 ( \29329 , RIe5359a0_6877, \29328 );
buf \U$23675 ( \29330 , \29028 );
buf \U$23676 ( \29331 , \29028 );
buf \U$23677 ( \29332 , \29028 );
buf \U$23678 ( \29333 , \29028 );
buf \U$23679 ( \29334 , \29028 );
buf \U$23680 ( \29335 , \29028 );
buf \U$23681 ( \29336 , \29028 );
buf \U$23682 ( \29337 , \29028 );
buf \U$23683 ( \29338 , \29028 );
buf \U$23684 ( \29339 , \29028 );
buf \U$23685 ( \29340 , \29028 );
buf \U$23686 ( \29341 , \29028 );
buf \U$23687 ( \29342 , \29028 );
buf \U$23688 ( \29343 , \29028 );
buf \U$23689 ( \29344 , \29028 );
buf \U$23690 ( \29345 , \29028 );
buf \U$23691 ( \29346 , \29028 );
buf \U$23692 ( \29347 , \29028 );
buf \U$23693 ( \29348 , \29028 );
buf \U$23694 ( \29349 , \29028 );
buf \U$23695 ( \29350 , \29028 );
buf \U$23696 ( \29351 , \29028 );
buf \U$23697 ( \29352 , \29028 );
buf \U$23698 ( \29353 , \29028 );
buf \U$23699 ( \29354 , \29028 );
nor \U$23700 ( \29355 , \29056 , \29016 , \29058 , \29018 , \29021 , \29025 , \29028 , \29330 , \29331 , \29332 , \29333 , \29334 , \29335 , \29336 , \29337 , \29338 , \29339 , \29340 , \29341 , \29342 , \29343 , \29344 , \29345 , \29346 , \29347 , \29348 , \29349 , \29350 , \29351 , \29352 , \29353 , \29354 );
and \U$23701 ( \29356 , RIeab78c8_6895, \29355 );
buf \U$23702 ( \29357 , \29028 );
buf \U$23703 ( \29358 , \29028 );
buf \U$23704 ( \29359 , \29028 );
buf \U$23705 ( \29360 , \29028 );
buf \U$23706 ( \29361 , \29028 );
buf \U$23707 ( \29362 , \29028 );
buf \U$23708 ( \29363 , \29028 );
buf \U$23709 ( \29364 , \29028 );
buf \U$23710 ( \29365 , \29028 );
buf \U$23711 ( \29366 , \29028 );
buf \U$23712 ( \29367 , \29028 );
buf \U$23713 ( \29368 , \29028 );
buf \U$23714 ( \29369 , \29028 );
buf \U$23715 ( \29370 , \29028 );
buf \U$23716 ( \29371 , \29028 );
buf \U$23717 ( \29372 , \29028 );
buf \U$23718 ( \29373 , \29028 );
buf \U$23719 ( \29374 , \29028 );
buf \U$23720 ( \29375 , \29028 );
buf \U$23721 ( \29376 , \29028 );
buf \U$23722 ( \29377 , \29028 );
buf \U$23723 ( \29378 , \29028 );
buf \U$23724 ( \29379 , \29028 );
buf \U$23725 ( \29380 , \29028 );
buf \U$23726 ( \29381 , \29028 );
nor \U$23727 ( \29382 , \29015 , \29016 , \29058 , \29018 , \29021 , \29025 , \29028 , \29357 , \29358 , \29359 , \29360 , \29361 , \29362 , \29363 , \29364 , \29365 , \29366 , \29367 , \29368 , \29369 , \29370 , \29371 , \29372 , \29373 , \29374 , \29375 , \29376 , \29377 , \29378 , \29379 , \29380 , \29381 );
and \U$23728 ( \29383 , RIeab7d00_6896, \29382 );
buf \U$23729 ( \29384 , \29028 );
buf \U$23730 ( \29385 , \29028 );
buf \U$23731 ( \29386 , \29028 );
buf \U$23732 ( \29387 , \29028 );
buf \U$23733 ( \29388 , \29028 );
buf \U$23734 ( \29389 , \29028 );
buf \U$23735 ( \29390 , \29028 );
buf \U$23736 ( \29391 , \29028 );
buf \U$23737 ( \29392 , \29028 );
buf \U$23738 ( \29393 , \29028 );
buf \U$23739 ( \29394 , \29028 );
buf \U$23740 ( \29395 , \29028 );
buf \U$23741 ( \29396 , \29028 );
buf \U$23742 ( \29397 , \29028 );
buf \U$23743 ( \29398 , \29028 );
buf \U$23744 ( \29399 , \29028 );
buf \U$23745 ( \29400 , \29028 );
buf \U$23746 ( \29401 , \29028 );
buf \U$23747 ( \29402 , \29028 );
buf \U$23748 ( \29403 , \29028 );
buf \U$23749 ( \29404 , \29028 );
buf \U$23750 ( \29405 , \29028 );
buf \U$23751 ( \29406 , \29028 );
buf \U$23752 ( \29407 , \29028 );
buf \U$23753 ( \29408 , \29028 );
nor \U$23754 ( \29409 , \29056 , \29057 , \29017 , \29018 , \29021 , \29025 , \29028 , \29384 , \29385 , \29386 , \29387 , \29388 , \29389 , \29390 , \29391 , \29392 , \29393 , \29394 , \29395 , \29396 , \29397 , \29398 , \29399 , \29400 , \29401 , \29402 , \29403 , \29404 , \29405 , \29406 , \29407 , \29408 );
and \U$23755 ( \29410 , RIeacfa18_6902, \29409 );
buf \U$23756 ( \29411 , \29028 );
buf \U$23757 ( \29412 , \29028 );
buf \U$23758 ( \29413 , \29028 );
buf \U$23759 ( \29414 , \29028 );
buf \U$23760 ( \29415 , \29028 );
buf \U$23761 ( \29416 , \29028 );
buf \U$23762 ( \29417 , \29028 );
buf \U$23763 ( \29418 , \29028 );
buf \U$23764 ( \29419 , \29028 );
buf \U$23765 ( \29420 , \29028 );
buf \U$23766 ( \29421 , \29028 );
buf \U$23767 ( \29422 , \29028 );
buf \U$23768 ( \29423 , \29028 );
buf \U$23769 ( \29424 , \29028 );
buf \U$23770 ( \29425 , \29028 );
buf \U$23771 ( \29426 , \29028 );
buf \U$23772 ( \29427 , \29028 );
buf \U$23773 ( \29428 , \29028 );
buf \U$23774 ( \29429 , \29028 );
buf \U$23775 ( \29430 , \29028 );
buf \U$23776 ( \29431 , \29028 );
buf \U$23777 ( \29432 , \29028 );
buf \U$23778 ( \29433 , \29028 );
buf \U$23779 ( \29434 , \29028 );
buf \U$23780 ( \29435 , \29028 );
nor \U$23781 ( \29436 , \29015 , \29057 , \29017 , \29018 , \29021 , \29025 , \29028 , \29411 , \29412 , \29413 , \29414 , \29415 , \29416 , \29417 , \29418 , \29419 , \29420 , \29421 , \29422 , \29423 , \29424 , \29425 , \29426 , \29427 , \29428 , \29429 , \29430 , \29431 , \29432 , \29433 , \29434 , \29435 );
and \U$23782 ( \29437 , RIeab6518_6891, \29436 );
buf \U$23783 ( \29438 , \29028 );
buf \U$23784 ( \29439 , \29028 );
buf \U$23785 ( \29440 , \29028 );
buf \U$23786 ( \29441 , \29028 );
buf \U$23787 ( \29442 , \29028 );
buf \U$23788 ( \29443 , \29028 );
buf \U$23789 ( \29444 , \29028 );
buf \U$23790 ( \29445 , \29028 );
buf \U$23791 ( \29446 , \29028 );
buf \U$23792 ( \29447 , \29028 );
buf \U$23793 ( \29448 , \29028 );
buf \U$23794 ( \29449 , \29028 );
buf \U$23795 ( \29450 , \29028 );
buf \U$23796 ( \29451 , \29028 );
buf \U$23797 ( \29452 , \29028 );
buf \U$23798 ( \29453 , \29028 );
buf \U$23799 ( \29454 , \29028 );
buf \U$23800 ( \29455 , \29028 );
buf \U$23801 ( \29456 , \29028 );
buf \U$23802 ( \29457 , \29028 );
buf \U$23803 ( \29458 , \29028 );
buf \U$23804 ( \29459 , \29028 );
buf \U$23805 ( \29460 , \29028 );
buf \U$23806 ( \29461 , \29028 );
buf \U$23807 ( \29462 , \29028 );
nor \U$23808 ( \29463 , \29056 , \29016 , \29017 , \29018 , \29021 , \29025 , \29028 , \29438 , \29439 , \29440 , \29441 , \29442 , \29443 , \29444 , \29445 , \29446 , \29447 , \29448 , \29449 , \29450 , \29451 , \29452 , \29453 , \29454 , \29455 , \29456 , \29457 , \29458 , \29459 , \29460 , \29461 , \29462 );
and \U$23809 ( \29464 , RIeb352c8_6904, \29463 );
or \U$23810 ( \29465 , \29055 , \29086 , \29113 , \29140 , \29167 , \29194 , \29221 , \29248 , \29275 , \29302 , \29329 , \29356 , \29383 , \29410 , \29437 , \29464 );
buf \U$23811 ( \29466 , \29028 );
not \U$23812 ( \29467 , \29466 );
buf \U$23813 ( \29468 , \29016 );
buf \U$23814 ( \29469 , \29017 );
buf \U$23815 ( \29470 , \29018 );
buf \U$23816 ( \29471 , \29021 );
buf \U$23817 ( \29472 , \29025 );
buf \U$23818 ( \29473 , \29028 );
buf \U$23819 ( \29474 , \29028 );
buf \U$23820 ( \29475 , \29028 );
buf \U$23821 ( \29476 , \29028 );
buf \U$23822 ( \29477 , \29028 );
buf \U$23823 ( \29478 , \29028 );
buf \U$23824 ( \29479 , \29028 );
buf \U$23825 ( \29480 , \29028 );
buf \U$23826 ( \29481 , \29028 );
buf \U$23827 ( \29482 , \29028 );
buf \U$23828 ( \29483 , \29028 );
buf \U$23829 ( \29484 , \29028 );
buf \U$23830 ( \29485 , \29028 );
buf \U$23831 ( \29486 , \29028 );
buf \U$23832 ( \29487 , \29028 );
buf \U$23833 ( \29488 , \29028 );
buf \U$23834 ( \29489 , \29028 );
buf \U$23835 ( \29490 , \29028 );
buf \U$23836 ( \29491 , \29028 );
buf \U$23837 ( \29492 , \29028 );
buf \U$23838 ( \29493 , \29028 );
buf \U$23839 ( \29494 , \29028 );
buf \U$23840 ( \29495 , \29028 );
buf \U$23841 ( \29496 , \29028 );
buf \U$23842 ( \29497 , \29028 );
buf \U$23843 ( \29498 , \29015 );
or \U$23844 ( \29499 , \29468 , \29469 , \29470 , \29471 , \29472 , \29473 , \29474 , \29475 , \29476 , \29477 , \29478 , \29479 , \29480 , \29481 , \29482 , \29483 , \29484 , \29485 , \29486 , \29487 , \29488 , \29489 , \29490 , \29491 , \29492 , \29493 , \29494 , \29495 , \29496 , \29497 , \29498 );
nand \U$23845 ( \29500 , \29467 , \29499 );
buf \U$23846 ( \29501 , \29500 );
buf \U$23847 ( \29502 , \29028 );
not \U$23848 ( \29503 , \29502 );
buf \U$23849 ( \29504 , \29025 );
buf \U$23850 ( \29505 , \29028 );
buf \U$23851 ( \29506 , \29028 );
buf \U$23852 ( \29507 , \29028 );
buf \U$23853 ( \29508 , \29028 );
buf \U$23854 ( \29509 , \29028 );
buf \U$23855 ( \29510 , \29028 );
buf \U$23856 ( \29511 , \29028 );
buf \U$23857 ( \29512 , \29028 );
buf \U$23858 ( \29513 , \29028 );
buf \U$23859 ( \29514 , \29028 );
buf \U$23860 ( \29515 , \29028 );
buf \U$23861 ( \29516 , \29028 );
buf \U$23862 ( \29517 , \29028 );
buf \U$23863 ( \29518 , \29028 );
buf \U$23864 ( \29519 , \29028 );
buf \U$23865 ( \29520 , \29028 );
buf \U$23866 ( \29521 , \29028 );
buf \U$23867 ( \29522 , \29028 );
buf \U$23868 ( \29523 , \29028 );
buf \U$23869 ( \29524 , \29028 );
buf \U$23870 ( \29525 , \29028 );
buf \U$23871 ( \29526 , \29028 );
buf \U$23872 ( \29527 , \29028 );
buf \U$23873 ( \29528 , \29028 );
buf \U$23874 ( \29529 , \29028 );
buf \U$23875 ( \29530 , \29021 );
buf \U$23876 ( \29531 , \29015 );
buf \U$23877 ( \29532 , \29016 );
buf \U$23878 ( \29533 , \29017 );
buf \U$23879 ( \29534 , \29018 );
or \U$23880 ( \29535 , \29531 , \29532 , \29533 , \29534 );
and \U$23881 ( \29536 , \29530 , \29535 );
or \U$23882 ( \29537 , \29504 , \29505 , \29506 , \29507 , \29508 , \29509 , \29510 , \29511 , \29512 , \29513 , \29514 , \29515 , \29516 , \29517 , \29518 , \29519 , \29520 , \29521 , \29522 , \29523 , \29524 , \29525 , \29526 , \29527 , \29528 , \29529 , \29536 );
and \U$23883 ( \29538 , \29503 , \29537 );
buf \U$23884 ( \29539 , \29538 );
or \U$23885 ( \29540 , \29501 , \29539 );
_DC g8a6e ( \29541_nG8a6e , \29465 , \29540 );
not \U$23886 ( \29542 , \29541_nG8a6e );
buf \U$23887 ( \29543 , RIb7b9608_246);
buf \U$23888 ( \29544 , \29028 );
buf \U$23889 ( \29545 , \29028 );
buf \U$23890 ( \29546 , \29028 );
buf \U$23891 ( \29547 , \29028 );
buf \U$23892 ( \29548 , \29028 );
buf \U$23893 ( \29549 , \29028 );
buf \U$23894 ( \29550 , \29028 );
buf \U$23895 ( \29551 , \29028 );
buf \U$23896 ( \29552 , \29028 );
buf \U$23897 ( \29553 , \29028 );
buf \U$23898 ( \29554 , \29028 );
buf \U$23899 ( \29555 , \29028 );
buf \U$23900 ( \29556 , \29028 );
buf \U$23901 ( \29557 , \29028 );
buf \U$23902 ( \29558 , \29028 );
buf \U$23903 ( \29559 , \29028 );
buf \U$23904 ( \29560 , \29028 );
buf \U$23905 ( \29561 , \29028 );
buf \U$23906 ( \29562 , \29028 );
buf \U$23907 ( \29563 , \29028 );
buf \U$23908 ( \29564 , \29028 );
buf \U$23909 ( \29565 , \29028 );
buf \U$23910 ( \29566 , \29028 );
buf \U$23911 ( \29567 , \29028 );
buf \U$23912 ( \29568 , \29028 );
nor \U$23913 ( \29569 , \29015 , \29016 , \29017 , \29018 , \29022 , \29025 , \29028 , \29544 , \29545 , \29546 , \29547 , \29548 , \29549 , \29550 , \29551 , \29552 , \29553 , \29554 , \29555 , \29556 , \29557 , \29558 , \29559 , \29560 , \29561 , \29562 , \29563 , \29564 , \29565 , \29566 , \29567 , \29568 );
and \U$23914 ( \29570 , \7117 , \29569 );
buf \U$23915 ( \29571 , \29028 );
buf \U$23916 ( \29572 , \29028 );
buf \U$23917 ( \29573 , \29028 );
buf \U$23918 ( \29574 , \29028 );
buf \U$23919 ( \29575 , \29028 );
buf \U$23920 ( \29576 , \29028 );
buf \U$23921 ( \29577 , \29028 );
buf \U$23922 ( \29578 , \29028 );
buf \U$23923 ( \29579 , \29028 );
buf \U$23924 ( \29580 , \29028 );
buf \U$23925 ( \29581 , \29028 );
buf \U$23926 ( \29582 , \29028 );
buf \U$23927 ( \29583 , \29028 );
buf \U$23928 ( \29584 , \29028 );
buf \U$23929 ( \29585 , \29028 );
buf \U$23930 ( \29586 , \29028 );
buf \U$23931 ( \29587 , \29028 );
buf \U$23932 ( \29588 , \29028 );
buf \U$23933 ( \29589 , \29028 );
buf \U$23934 ( \29590 , \29028 );
buf \U$23935 ( \29591 , \29028 );
buf \U$23936 ( \29592 , \29028 );
buf \U$23937 ( \29593 , \29028 );
buf \U$23938 ( \29594 , \29028 );
buf \U$23939 ( \29595 , \29028 );
nor \U$23940 ( \29596 , \29056 , \29057 , \29058 , \29059 , \29021 , \29025 , \29028 , \29571 , \29572 , \29573 , \29574 , \29575 , \29576 , \29577 , \29578 , \29579 , \29580 , \29581 , \29582 , \29583 , \29584 , \29585 , \29586 , \29587 , \29588 , \29589 , \29590 , \29591 , \29592 , \29593 , \29594 , \29595 );
and \U$23941 ( \29597 , \7119 , \29596 );
buf \U$23942 ( \29598 , \29028 );
buf \U$23943 ( \29599 , \29028 );
buf \U$23944 ( \29600 , \29028 );
buf \U$23945 ( \29601 , \29028 );
buf \U$23946 ( \29602 , \29028 );
buf \U$23947 ( \29603 , \29028 );
buf \U$23948 ( \29604 , \29028 );
buf \U$23949 ( \29605 , \29028 );
buf \U$23950 ( \29606 , \29028 );
buf \U$23951 ( \29607 , \29028 );
buf \U$23952 ( \29608 , \29028 );
buf \U$23953 ( \29609 , \29028 );
buf \U$23954 ( \29610 , \29028 );
buf \U$23955 ( \29611 , \29028 );
buf \U$23956 ( \29612 , \29028 );
buf \U$23957 ( \29613 , \29028 );
buf \U$23958 ( \29614 , \29028 );
buf \U$23959 ( \29615 , \29028 );
buf \U$23960 ( \29616 , \29028 );
buf \U$23961 ( \29617 , \29028 );
buf \U$23962 ( \29618 , \29028 );
buf \U$23963 ( \29619 , \29028 );
buf \U$23964 ( \29620 , \29028 );
buf \U$23965 ( \29621 , \29028 );
buf \U$23966 ( \29622 , \29028 );
nor \U$23967 ( \29623 , \29015 , \29057 , \29058 , \29059 , \29021 , \29025 , \29028 , \29598 , \29599 , \29600 , \29601 , \29602 , \29603 , \29604 , \29605 , \29606 , \29607 , \29608 , \29609 , \29610 , \29611 , \29612 , \29613 , \29614 , \29615 , \29616 , \29617 , \29618 , \29619 , \29620 , \29621 , \29622 );
and \U$23968 ( \29624 , \7864 , \29623 );
buf \U$23969 ( \29625 , \29028 );
buf \U$23970 ( \29626 , \29028 );
buf \U$23971 ( \29627 , \29028 );
buf \U$23972 ( \29628 , \29028 );
buf \U$23973 ( \29629 , \29028 );
buf \U$23974 ( \29630 , \29028 );
buf \U$23975 ( \29631 , \29028 );
buf \U$23976 ( \29632 , \29028 );
buf \U$23977 ( \29633 , \29028 );
buf \U$23978 ( \29634 , \29028 );
buf \U$23979 ( \29635 , \29028 );
buf \U$23980 ( \29636 , \29028 );
buf \U$23981 ( \29637 , \29028 );
buf \U$23982 ( \29638 , \29028 );
buf \U$23983 ( \29639 , \29028 );
buf \U$23984 ( \29640 , \29028 );
buf \U$23985 ( \29641 , \29028 );
buf \U$23986 ( \29642 , \29028 );
buf \U$23987 ( \29643 , \29028 );
buf \U$23988 ( \29644 , \29028 );
buf \U$23989 ( \29645 , \29028 );
buf \U$23990 ( \29646 , \29028 );
buf \U$23991 ( \29647 , \29028 );
buf \U$23992 ( \29648 , \29028 );
buf \U$23993 ( \29649 , \29028 );
nor \U$23994 ( \29650 , \29056 , \29016 , \29058 , \29059 , \29021 , \29025 , \29028 , \29625 , \29626 , \29627 , \29628 , \29629 , \29630 , \29631 , \29632 , \29633 , \29634 , \29635 , \29636 , \29637 , \29638 , \29639 , \29640 , \29641 , \29642 , \29643 , \29644 , \29645 , \29646 , \29647 , \29648 , \29649 );
and \U$23995 ( \29651 , \7892 , \29650 );
buf \U$23996 ( \29652 , \29028 );
buf \U$23997 ( \29653 , \29028 );
buf \U$23998 ( \29654 , \29028 );
buf \U$23999 ( \29655 , \29028 );
buf \U$24000 ( \29656 , \29028 );
buf \U$24001 ( \29657 , \29028 );
buf \U$24002 ( \29658 , \29028 );
buf \U$24003 ( \29659 , \29028 );
buf \U$24004 ( \29660 , \29028 );
buf \U$24005 ( \29661 , \29028 );
buf \U$24006 ( \29662 , \29028 );
buf \U$24007 ( \29663 , \29028 );
buf \U$24008 ( \29664 , \29028 );
buf \U$24009 ( \29665 , \29028 );
buf \U$24010 ( \29666 , \29028 );
buf \U$24011 ( \29667 , \29028 );
buf \U$24012 ( \29668 , \29028 );
buf \U$24013 ( \29669 , \29028 );
buf \U$24014 ( \29670 , \29028 );
buf \U$24015 ( \29671 , \29028 );
buf \U$24016 ( \29672 , \29028 );
buf \U$24017 ( \29673 , \29028 );
buf \U$24018 ( \29674 , \29028 );
buf \U$24019 ( \29675 , \29028 );
buf \U$24020 ( \29676 , \29028 );
nor \U$24021 ( \29677 , \29015 , \29016 , \29058 , \29059 , \29021 , \29025 , \29028 , \29652 , \29653 , \29654 , \29655 , \29656 , \29657 , \29658 , \29659 , \29660 , \29661 , \29662 , \29663 , \29664 , \29665 , \29666 , \29667 , \29668 , \29669 , \29670 , \29671 , \29672 , \29673 , \29674 , \29675 , \29676 );
and \U$24022 ( \29678 , \7920 , \29677 );
buf \U$24023 ( \29679 , \29028 );
buf \U$24024 ( \29680 , \29028 );
buf \U$24025 ( \29681 , \29028 );
buf \U$24026 ( \29682 , \29028 );
buf \U$24027 ( \29683 , \29028 );
buf \U$24028 ( \29684 , \29028 );
buf \U$24029 ( \29685 , \29028 );
buf \U$24030 ( \29686 , \29028 );
buf \U$24031 ( \29687 , \29028 );
buf \U$24032 ( \29688 , \29028 );
buf \U$24033 ( \29689 , \29028 );
buf \U$24034 ( \29690 , \29028 );
buf \U$24035 ( \29691 , \29028 );
buf \U$24036 ( \29692 , \29028 );
buf \U$24037 ( \29693 , \29028 );
buf \U$24038 ( \29694 , \29028 );
buf \U$24039 ( \29695 , \29028 );
buf \U$24040 ( \29696 , \29028 );
buf \U$24041 ( \29697 , \29028 );
buf \U$24042 ( \29698 , \29028 );
buf \U$24043 ( \29699 , \29028 );
buf \U$24044 ( \29700 , \29028 );
buf \U$24045 ( \29701 , \29028 );
buf \U$24046 ( \29702 , \29028 );
buf \U$24047 ( \29703 , \29028 );
nor \U$24048 ( \29704 , \29056 , \29057 , \29017 , \29059 , \29021 , \29025 , \29028 , \29679 , \29680 , \29681 , \29682 , \29683 , \29684 , \29685 , \29686 , \29687 , \29688 , \29689 , \29690 , \29691 , \29692 , \29693 , \29694 , \29695 , \29696 , \29697 , \29698 , \29699 , \29700 , \29701 , \29702 , \29703 );
and \U$24049 ( \29705 , \7948 , \29704 );
buf \U$24050 ( \29706 , \29028 );
buf \U$24051 ( \29707 , \29028 );
buf \U$24052 ( \29708 , \29028 );
buf \U$24053 ( \29709 , \29028 );
buf \U$24054 ( \29710 , \29028 );
buf \U$24055 ( \29711 , \29028 );
buf \U$24056 ( \29712 , \29028 );
buf \U$24057 ( \29713 , \29028 );
buf \U$24058 ( \29714 , \29028 );
buf \U$24059 ( \29715 , \29028 );
buf \U$24060 ( \29716 , \29028 );
buf \U$24061 ( \29717 , \29028 );
buf \U$24062 ( \29718 , \29028 );
buf \U$24063 ( \29719 , \29028 );
buf \U$24064 ( \29720 , \29028 );
buf \U$24065 ( \29721 , \29028 );
buf \U$24066 ( \29722 , \29028 );
buf \U$24067 ( \29723 , \29028 );
buf \U$24068 ( \29724 , \29028 );
buf \U$24069 ( \29725 , \29028 );
buf \U$24070 ( \29726 , \29028 );
buf \U$24071 ( \29727 , \29028 );
buf \U$24072 ( \29728 , \29028 );
buf \U$24073 ( \29729 , \29028 );
buf \U$24074 ( \29730 , \29028 );
nor \U$24075 ( \29731 , \29015 , \29057 , \29017 , \29059 , \29021 , \29025 , \29028 , \29706 , \29707 , \29708 , \29709 , \29710 , \29711 , \29712 , \29713 , \29714 , \29715 , \29716 , \29717 , \29718 , \29719 , \29720 , \29721 , \29722 , \29723 , \29724 , \29725 , \29726 , \29727 , \29728 , \29729 , \29730 );
and \U$24076 ( \29732 , \7976 , \29731 );
buf \U$24077 ( \29733 , \29028 );
buf \U$24078 ( \29734 , \29028 );
buf \U$24079 ( \29735 , \29028 );
buf \U$24080 ( \29736 , \29028 );
buf \U$24081 ( \29737 , \29028 );
buf \U$24082 ( \29738 , \29028 );
buf \U$24083 ( \29739 , \29028 );
buf \U$24084 ( \29740 , \29028 );
buf \U$24085 ( \29741 , \29028 );
buf \U$24086 ( \29742 , \29028 );
buf \U$24087 ( \29743 , \29028 );
buf \U$24088 ( \29744 , \29028 );
buf \U$24089 ( \29745 , \29028 );
buf \U$24090 ( \29746 , \29028 );
buf \U$24091 ( \29747 , \29028 );
buf \U$24092 ( \29748 , \29028 );
buf \U$24093 ( \29749 , \29028 );
buf \U$24094 ( \29750 , \29028 );
buf \U$24095 ( \29751 , \29028 );
buf \U$24096 ( \29752 , \29028 );
buf \U$24097 ( \29753 , \29028 );
buf \U$24098 ( \29754 , \29028 );
buf \U$24099 ( \29755 , \29028 );
buf \U$24100 ( \29756 , \29028 );
buf \U$24101 ( \29757 , \29028 );
nor \U$24102 ( \29758 , \29056 , \29016 , \29017 , \29059 , \29021 , \29025 , \29028 , \29733 , \29734 , \29735 , \29736 , \29737 , \29738 , \29739 , \29740 , \29741 , \29742 , \29743 , \29744 , \29745 , \29746 , \29747 , \29748 , \29749 , \29750 , \29751 , \29752 , \29753 , \29754 , \29755 , \29756 , \29757 );
and \U$24103 ( \29759 , \8004 , \29758 );
buf \U$24104 ( \29760 , \29028 );
buf \U$24105 ( \29761 , \29028 );
buf \U$24106 ( \29762 , \29028 );
buf \U$24107 ( \29763 , \29028 );
buf \U$24108 ( \29764 , \29028 );
buf \U$24109 ( \29765 , \29028 );
buf \U$24110 ( \29766 , \29028 );
buf \U$24111 ( \29767 , \29028 );
buf \U$24112 ( \29768 , \29028 );
buf \U$24113 ( \29769 , \29028 );
buf \U$24114 ( \29770 , \29028 );
buf \U$24115 ( \29771 , \29028 );
buf \U$24116 ( \29772 , \29028 );
buf \U$24117 ( \29773 , \29028 );
buf \U$24118 ( \29774 , \29028 );
buf \U$24119 ( \29775 , \29028 );
buf \U$24120 ( \29776 , \29028 );
buf \U$24121 ( \29777 , \29028 );
buf \U$24122 ( \29778 , \29028 );
buf \U$24123 ( \29779 , \29028 );
buf \U$24124 ( \29780 , \29028 );
buf \U$24125 ( \29781 , \29028 );
buf \U$24126 ( \29782 , \29028 );
buf \U$24127 ( \29783 , \29028 );
buf \U$24128 ( \29784 , \29028 );
nor \U$24129 ( \29785 , \29015 , \29016 , \29017 , \29059 , \29021 , \29025 , \29028 , \29760 , \29761 , \29762 , \29763 , \29764 , \29765 , \29766 , \29767 , \29768 , \29769 , \29770 , \29771 , \29772 , \29773 , \29774 , \29775 , \29776 , \29777 , \29778 , \29779 , \29780 , \29781 , \29782 , \29783 , \29784 );
and \U$24130 ( \29786 , \8032 , \29785 );
buf \U$24131 ( \29787 , \29028 );
buf \U$24132 ( \29788 , \29028 );
buf \U$24133 ( \29789 , \29028 );
buf \U$24134 ( \29790 , \29028 );
buf \U$24135 ( \29791 , \29028 );
buf \U$24136 ( \29792 , \29028 );
buf \U$24137 ( \29793 , \29028 );
buf \U$24138 ( \29794 , \29028 );
buf \U$24139 ( \29795 , \29028 );
buf \U$24140 ( \29796 , \29028 );
buf \U$24141 ( \29797 , \29028 );
buf \U$24142 ( \29798 , \29028 );
buf \U$24143 ( \29799 , \29028 );
buf \U$24144 ( \29800 , \29028 );
buf \U$24145 ( \29801 , \29028 );
buf \U$24146 ( \29802 , \29028 );
buf \U$24147 ( \29803 , \29028 );
buf \U$24148 ( \29804 , \29028 );
buf \U$24149 ( \29805 , \29028 );
buf \U$24150 ( \29806 , \29028 );
buf \U$24151 ( \29807 , \29028 );
buf \U$24152 ( \29808 , \29028 );
buf \U$24153 ( \29809 , \29028 );
buf \U$24154 ( \29810 , \29028 );
buf \U$24155 ( \29811 , \29028 );
nor \U$24156 ( \29812 , \29056 , \29057 , \29058 , \29018 , \29021 , \29025 , \29028 , \29787 , \29788 , \29789 , \29790 , \29791 , \29792 , \29793 , \29794 , \29795 , \29796 , \29797 , \29798 , \29799 , \29800 , \29801 , \29802 , \29803 , \29804 , \29805 , \29806 , \29807 , \29808 , \29809 , \29810 , \29811 );
and \U$24157 ( \29813 , \8060 , \29812 );
buf \U$24158 ( \29814 , \29028 );
buf \U$24159 ( \29815 , \29028 );
buf \U$24160 ( \29816 , \29028 );
buf \U$24161 ( \29817 , \29028 );
buf \U$24162 ( \29818 , \29028 );
buf \U$24163 ( \29819 , \29028 );
buf \U$24164 ( \29820 , \29028 );
buf \U$24165 ( \29821 , \29028 );
buf \U$24166 ( \29822 , \29028 );
buf \U$24167 ( \29823 , \29028 );
buf \U$24168 ( \29824 , \29028 );
buf \U$24169 ( \29825 , \29028 );
buf \U$24170 ( \29826 , \29028 );
buf \U$24171 ( \29827 , \29028 );
buf \U$24172 ( \29828 , \29028 );
buf \U$24173 ( \29829 , \29028 );
buf \U$24174 ( \29830 , \29028 );
buf \U$24175 ( \29831 , \29028 );
buf \U$24176 ( \29832 , \29028 );
buf \U$24177 ( \29833 , \29028 );
buf \U$24178 ( \29834 , \29028 );
buf \U$24179 ( \29835 , \29028 );
buf \U$24180 ( \29836 , \29028 );
buf \U$24181 ( \29837 , \29028 );
buf \U$24182 ( \29838 , \29028 );
nor \U$24183 ( \29839 , \29015 , \29057 , \29058 , \29018 , \29021 , \29025 , \29028 , \29814 , \29815 , \29816 , \29817 , \29818 , \29819 , \29820 , \29821 , \29822 , \29823 , \29824 , \29825 , \29826 , \29827 , \29828 , \29829 , \29830 , \29831 , \29832 , \29833 , \29834 , \29835 , \29836 , \29837 , \29838 );
and \U$24184 ( \29840 , \8088 , \29839 );
buf \U$24185 ( \29841 , \29028 );
buf \U$24186 ( \29842 , \29028 );
buf \U$24187 ( \29843 , \29028 );
buf \U$24188 ( \29844 , \29028 );
buf \U$24189 ( \29845 , \29028 );
buf \U$24190 ( \29846 , \29028 );
buf \U$24191 ( \29847 , \29028 );
buf \U$24192 ( \29848 , \29028 );
buf \U$24193 ( \29849 , \29028 );
buf \U$24194 ( \29850 , \29028 );
buf \U$24195 ( \29851 , \29028 );
buf \U$24196 ( \29852 , \29028 );
buf \U$24197 ( \29853 , \29028 );
buf \U$24198 ( \29854 , \29028 );
buf \U$24199 ( \29855 , \29028 );
buf \U$24200 ( \29856 , \29028 );
buf \U$24201 ( \29857 , \29028 );
buf \U$24202 ( \29858 , \29028 );
buf \U$24203 ( \29859 , \29028 );
buf \U$24204 ( \29860 , \29028 );
buf \U$24205 ( \29861 , \29028 );
buf \U$24206 ( \29862 , \29028 );
buf \U$24207 ( \29863 , \29028 );
buf \U$24208 ( \29864 , \29028 );
buf \U$24209 ( \29865 , \29028 );
nor \U$24210 ( \29866 , \29056 , \29016 , \29058 , \29018 , \29021 , \29025 , \29028 , \29841 , \29842 , \29843 , \29844 , \29845 , \29846 , \29847 , \29848 , \29849 , \29850 , \29851 , \29852 , \29853 , \29854 , \29855 , \29856 , \29857 , \29858 , \29859 , \29860 , \29861 , \29862 , \29863 , \29864 , \29865 );
and \U$24211 ( \29867 , \8116 , \29866 );
buf \U$24212 ( \29868 , \29028 );
buf \U$24213 ( \29869 , \29028 );
buf \U$24214 ( \29870 , \29028 );
buf \U$24215 ( \29871 , \29028 );
buf \U$24216 ( \29872 , \29028 );
buf \U$24217 ( \29873 , \29028 );
buf \U$24218 ( \29874 , \29028 );
buf \U$24219 ( \29875 , \29028 );
buf \U$24220 ( \29876 , \29028 );
buf \U$24221 ( \29877 , \29028 );
buf \U$24222 ( \29878 , \29028 );
buf \U$24223 ( \29879 , \29028 );
buf \U$24224 ( \29880 , \29028 );
buf \U$24225 ( \29881 , \29028 );
buf \U$24226 ( \29882 , \29028 );
buf \U$24227 ( \29883 , \29028 );
buf \U$24228 ( \29884 , \29028 );
buf \U$24229 ( \29885 , \29028 );
buf \U$24230 ( \29886 , \29028 );
buf \U$24231 ( \29887 , \29028 );
buf \U$24232 ( \29888 , \29028 );
buf \U$24233 ( \29889 , \29028 );
buf \U$24234 ( \29890 , \29028 );
buf \U$24235 ( \29891 , \29028 );
buf \U$24236 ( \29892 , \29028 );
nor \U$24237 ( \29893 , \29015 , \29016 , \29058 , \29018 , \29021 , \29025 , \29028 , \29868 , \29869 , \29870 , \29871 , \29872 , \29873 , \29874 , \29875 , \29876 , \29877 , \29878 , \29879 , \29880 , \29881 , \29882 , \29883 , \29884 , \29885 , \29886 , \29887 , \29888 , \29889 , \29890 , \29891 , \29892 );
and \U$24238 ( \29894 , \8144 , \29893 );
buf \U$24239 ( \29895 , \29028 );
buf \U$24240 ( \29896 , \29028 );
buf \U$24241 ( \29897 , \29028 );
buf \U$24242 ( \29898 , \29028 );
buf \U$24243 ( \29899 , \29028 );
buf \U$24244 ( \29900 , \29028 );
buf \U$24245 ( \29901 , \29028 );
buf \U$24246 ( \29902 , \29028 );
buf \U$24247 ( \29903 , \29028 );
buf \U$24248 ( \29904 , \29028 );
buf \U$24249 ( \29905 , \29028 );
buf \U$24250 ( \29906 , \29028 );
buf \U$24251 ( \29907 , \29028 );
buf \U$24252 ( \29908 , \29028 );
buf \U$24253 ( \29909 , \29028 );
buf \U$24254 ( \29910 , \29028 );
buf \U$24255 ( \29911 , \29028 );
buf \U$24256 ( \29912 , \29028 );
buf \U$24257 ( \29913 , \29028 );
buf \U$24258 ( \29914 , \29028 );
buf \U$24259 ( \29915 , \29028 );
buf \U$24260 ( \29916 , \29028 );
buf \U$24261 ( \29917 , \29028 );
buf \U$24262 ( \29918 , \29028 );
buf \U$24263 ( \29919 , \29028 );
nor \U$24264 ( \29920 , \29056 , \29057 , \29017 , \29018 , \29021 , \29025 , \29028 , \29895 , \29896 , \29897 , \29898 , \29899 , \29900 , \29901 , \29902 , \29903 , \29904 , \29905 , \29906 , \29907 , \29908 , \29909 , \29910 , \29911 , \29912 , \29913 , \29914 , \29915 , \29916 , \29917 , \29918 , \29919 );
and \U$24265 ( \29921 , \8172 , \29920 );
buf \U$24266 ( \29922 , \29028 );
buf \U$24267 ( \29923 , \29028 );
buf \U$24268 ( \29924 , \29028 );
buf \U$24269 ( \29925 , \29028 );
buf \U$24270 ( \29926 , \29028 );
buf \U$24271 ( \29927 , \29028 );
buf \U$24272 ( \29928 , \29028 );
buf \U$24273 ( \29929 , \29028 );
buf \U$24274 ( \29930 , \29028 );
buf \U$24275 ( \29931 , \29028 );
buf \U$24276 ( \29932 , \29028 );
buf \U$24277 ( \29933 , \29028 );
buf \U$24278 ( \29934 , \29028 );
buf \U$24279 ( \29935 , \29028 );
buf \U$24280 ( \29936 , \29028 );
buf \U$24281 ( \29937 , \29028 );
buf \U$24282 ( \29938 , \29028 );
buf \U$24283 ( \29939 , \29028 );
buf \U$24284 ( \29940 , \29028 );
buf \U$24285 ( \29941 , \29028 );
buf \U$24286 ( \29942 , \29028 );
buf \U$24287 ( \29943 , \29028 );
buf \U$24288 ( \29944 , \29028 );
buf \U$24289 ( \29945 , \29028 );
buf \U$24290 ( \29946 , \29028 );
nor \U$24291 ( \29947 , \29015 , \29057 , \29017 , \29018 , \29021 , \29025 , \29028 , \29922 , \29923 , \29924 , \29925 , \29926 , \29927 , \29928 , \29929 , \29930 , \29931 , \29932 , \29933 , \29934 , \29935 , \29936 , \29937 , \29938 , \29939 , \29940 , \29941 , \29942 , \29943 , \29944 , \29945 , \29946 );
and \U$24292 ( \29948 , \8200 , \29947 );
buf \U$24293 ( \29949 , \29028 );
buf \U$24294 ( \29950 , \29028 );
buf \U$24295 ( \29951 , \29028 );
buf \U$24296 ( \29952 , \29028 );
buf \U$24297 ( \29953 , \29028 );
buf \U$24298 ( \29954 , \29028 );
buf \U$24299 ( \29955 , \29028 );
buf \U$24300 ( \29956 , \29028 );
buf \U$24301 ( \29957 , \29028 );
buf \U$24302 ( \29958 , \29028 );
buf \U$24303 ( \29959 , \29028 );
buf \U$24304 ( \29960 , \29028 );
buf \U$24305 ( \29961 , \29028 );
buf \U$24306 ( \29962 , \29028 );
buf \U$24307 ( \29963 , \29028 );
buf \U$24308 ( \29964 , \29028 );
buf \U$24309 ( \29965 , \29028 );
buf \U$24310 ( \29966 , \29028 );
buf \U$24311 ( \29967 , \29028 );
buf \U$24312 ( \29968 , \29028 );
buf \U$24313 ( \29969 , \29028 );
buf \U$24314 ( \29970 , \29028 );
buf \U$24315 ( \29971 , \29028 );
buf \U$24316 ( \29972 , \29028 );
buf \U$24317 ( \29973 , \29028 );
nor \U$24318 ( \29974 , \29056 , \29016 , \29017 , \29018 , \29021 , \29025 , \29028 , \29949 , \29950 , \29951 , \29952 , \29953 , \29954 , \29955 , \29956 , \29957 , \29958 , \29959 , \29960 , \29961 , \29962 , \29963 , \29964 , \29965 , \29966 , \29967 , \29968 , \29969 , \29970 , \29971 , \29972 , \29973 );
and \U$24319 ( \29975 , \8228 , \29974 );
or \U$24320 ( \29976 , \29570 , \29597 , \29624 , \29651 , \29678 , \29705 , \29732 , \29759 , \29786 , \29813 , \29840 , \29867 , \29894 , \29921 , \29948 , \29975 );
buf \U$24321 ( \29977 , \29028 );
not \U$24322 ( \29978 , \29977 );
buf \U$24323 ( \29979 , \29016 );
buf \U$24324 ( \29980 , \29017 );
buf \U$24325 ( \29981 , \29018 );
buf \U$24326 ( \29982 , \29021 );
buf \U$24327 ( \29983 , \29025 );
buf \U$24328 ( \29984 , \29028 );
buf \U$24329 ( \29985 , \29028 );
buf \U$24330 ( \29986 , \29028 );
buf \U$24331 ( \29987 , \29028 );
buf \U$24332 ( \29988 , \29028 );
buf \U$24333 ( \29989 , \29028 );
buf \U$24334 ( \29990 , \29028 );
buf \U$24335 ( \29991 , \29028 );
buf \U$24336 ( \29992 , \29028 );
buf \U$24337 ( \29993 , \29028 );
buf \U$24338 ( \29994 , \29028 );
buf \U$24339 ( \29995 , \29028 );
buf \U$24340 ( \29996 , \29028 );
buf \U$24341 ( \29997 , \29028 );
buf \U$24342 ( \29998 , \29028 );
buf \U$24343 ( \29999 , \29028 );
buf \U$24344 ( \30000 , \29028 );
buf \U$24345 ( \30001 , \29028 );
buf \U$24346 ( \30002 , \29028 );
buf \U$24347 ( \30003 , \29028 );
buf \U$24348 ( \30004 , \29028 );
buf \U$24349 ( \30005 , \29028 );
buf \U$24350 ( \30006 , \29028 );
buf \U$24351 ( \30007 , \29028 );
buf \U$24352 ( \30008 , \29028 );
buf \U$24353 ( \30009 , \29015 );
or \U$24354 ( \30010 , \29979 , \29980 , \29981 , \29982 , \29983 , \29984 , \29985 , \29986 , \29987 , \29988 , \29989 , \29990 , \29991 , \29992 , \29993 , \29994 , \29995 , \29996 , \29997 , \29998 , \29999 , \30000 , \30001 , \30002 , \30003 , \30004 , \30005 , \30006 , \30007 , \30008 , \30009 );
nand \U$24355 ( \30011 , \29978 , \30010 );
buf \U$24356 ( \30012 , \30011 );
buf \U$24357 ( \30013 , \29028 );
not \U$24358 ( \30014 , \30013 );
buf \U$24359 ( \30015 , \29025 );
buf \U$24360 ( \30016 , \29028 );
buf \U$24361 ( \30017 , \29028 );
buf \U$24362 ( \30018 , \29028 );
buf \U$24363 ( \30019 , \29028 );
buf \U$24364 ( \30020 , \29028 );
buf \U$24365 ( \30021 , \29028 );
buf \U$24366 ( \30022 , \29028 );
buf \U$24367 ( \30023 , \29028 );
buf \U$24368 ( \30024 , \29028 );
buf \U$24369 ( \30025 , \29028 );
buf \U$24370 ( \30026 , \29028 );
buf \U$24371 ( \30027 , \29028 );
buf \U$24372 ( \30028 , \29028 );
buf \U$24373 ( \30029 , \29028 );
buf \U$24374 ( \30030 , \29028 );
buf \U$24375 ( \30031 , \29028 );
buf \U$24376 ( \30032 , \29028 );
buf \U$24377 ( \30033 , \29028 );
buf \U$24378 ( \30034 , \29028 );
buf \U$24379 ( \30035 , \29028 );
buf \U$24380 ( \30036 , \29028 );
buf \U$24381 ( \30037 , \29028 );
buf \U$24382 ( \30038 , \29028 );
buf \U$24383 ( \30039 , \29028 );
buf \U$24384 ( \30040 , \29028 );
buf \U$24385 ( \30041 , \29021 );
buf \U$24386 ( \30042 , \29015 );
buf \U$24387 ( \30043 , \29016 );
buf \U$24388 ( \30044 , \29017 );
buf \U$24389 ( \30045 , \29018 );
or \U$24390 ( \30046 , \30042 , \30043 , \30044 , \30045 );
and \U$24391 ( \30047 , \30041 , \30046 );
or \U$24392 ( \30048 , \30015 , \30016 , \30017 , \30018 , \30019 , \30020 , \30021 , \30022 , \30023 , \30024 , \30025 , \30026 , \30027 , \30028 , \30029 , \30030 , \30031 , \30032 , \30033 , \30034 , \30035 , \30036 , \30037 , \30038 , \30039 , \30040 , \30047 );
and \U$24393 ( \30049 , \30014 , \30048 );
buf \U$24394 ( \30050 , \30049 );
or \U$24395 ( \30051 , \30012 , \30050 );
_DC g8c6d ( \30052_nG8c6d , \29976 , \30051 );
buf \U$24396 ( \30053 , \30052_nG8c6d );
xor \U$24397 ( \30054 , \29543 , \30053 );
buf \U$24398 ( \30055 , RIb7b9590_247);
and \U$24399 ( \30056 , \7126 , \29569 );
and \U$24400 ( \30057 , \7128 , \29596 );
and \U$24401 ( \30058 , \8338 , \29623 );
and \U$24402 ( \30059 , \8340 , \29650 );
and \U$24403 ( \30060 , \8342 , \29677 );
and \U$24404 ( \30061 , \8344 , \29704 );
and \U$24405 ( \30062 , \8346 , \29731 );
and \U$24406 ( \30063 , \8348 , \29758 );
and \U$24407 ( \30064 , \8350 , \29785 );
and \U$24408 ( \30065 , \8352 , \29812 );
and \U$24409 ( \30066 , \8354 , \29839 );
and \U$24410 ( \30067 , \8356 , \29866 );
and \U$24411 ( \30068 , \8358 , \29893 );
and \U$24412 ( \30069 , \8360 , \29920 );
and \U$24413 ( \30070 , \8362 , \29947 );
and \U$24414 ( \30071 , \8364 , \29974 );
or \U$24415 ( \30072 , \30056 , \30057 , \30058 , \30059 , \30060 , \30061 , \30062 , \30063 , \30064 , \30065 , \30066 , \30067 , \30068 , \30069 , \30070 , \30071 );
_DC g8c82 ( \30073_nG8c82 , \30072 , \30051 );
buf \U$24416 ( \30074 , \30073_nG8c82 );
xor \U$24417 ( \30075 , \30055 , \30074 );
or \U$24418 ( \30076 , \30054 , \30075 );
buf \U$24419 ( \30077 , RIb7b9518_248);
and \U$24420 ( \30078 , \7136 , \29569 );
and \U$24421 ( \30079 , \7138 , \29596 );
and \U$24422 ( \30080 , \8374 , \29623 );
and \U$24423 ( \30081 , \8376 , \29650 );
and \U$24424 ( \30082 , \8378 , \29677 );
and \U$24425 ( \30083 , \8380 , \29704 );
and \U$24426 ( \30084 , \8382 , \29731 );
and \U$24427 ( \30085 , \8384 , \29758 );
and \U$24428 ( \30086 , \8386 , \29785 );
and \U$24429 ( \30087 , \8388 , \29812 );
and \U$24430 ( \30088 , \8390 , \29839 );
and \U$24431 ( \30089 , \8392 , \29866 );
and \U$24432 ( \30090 , \8394 , \29893 );
and \U$24433 ( \30091 , \8396 , \29920 );
and \U$24434 ( \30092 , \8398 , \29947 );
and \U$24435 ( \30093 , \8400 , \29974 );
or \U$24436 ( \30094 , \30078 , \30079 , \30080 , \30081 , \30082 , \30083 , \30084 , \30085 , \30086 , \30087 , \30088 , \30089 , \30090 , \30091 , \30092 , \30093 );
_DC g8c98 ( \30095_nG8c98 , \30094 , \30051 );
buf \U$24437 ( \30096 , \30095_nG8c98 );
xor \U$24438 ( \30097 , \30077 , \30096 );
or \U$24439 ( \30098 , \30076 , \30097 );
buf \U$24440 ( \30099 , RIb7b94a0_249);
and \U$24441 ( \30100 , \7146 , \29569 );
and \U$24442 ( \30101 , \7148 , \29596 );
and \U$24443 ( \30102 , \8410 , \29623 );
and \U$24444 ( \30103 , \8412 , \29650 );
and \U$24445 ( \30104 , \8414 , \29677 );
and \U$24446 ( \30105 , \8416 , \29704 );
and \U$24447 ( \30106 , \8418 , \29731 );
and \U$24448 ( \30107 , \8420 , \29758 );
and \U$24449 ( \30108 , \8422 , \29785 );
and \U$24450 ( \30109 , \8424 , \29812 );
and \U$24451 ( \30110 , \8426 , \29839 );
and \U$24452 ( \30111 , \8428 , \29866 );
and \U$24453 ( \30112 , \8430 , \29893 );
and \U$24454 ( \30113 , \8432 , \29920 );
and \U$24455 ( \30114 , \8434 , \29947 );
and \U$24456 ( \30115 , \8436 , \29974 );
or \U$24457 ( \30116 , \30100 , \30101 , \30102 , \30103 , \30104 , \30105 , \30106 , \30107 , \30108 , \30109 , \30110 , \30111 , \30112 , \30113 , \30114 , \30115 );
_DC g8cae ( \30117_nG8cae , \30116 , \30051 );
buf \U$24458 ( \30118 , \30117_nG8cae );
xor \U$24459 ( \30119 , \30099 , \30118 );
or \U$24460 ( \30120 , \30098 , \30119 );
buf \U$24461 ( \30121 , RIb7b9428_250);
and \U$24462 ( \30122 , \7156 , \29569 );
and \U$24463 ( \30123 , \7158 , \29596 );
and \U$24464 ( \30124 , \8446 , \29623 );
and \U$24465 ( \30125 , \8448 , \29650 );
and \U$24466 ( \30126 , \8450 , \29677 );
and \U$24467 ( \30127 , \8452 , \29704 );
and \U$24468 ( \30128 , \8454 , \29731 );
and \U$24469 ( \30129 , \8456 , \29758 );
and \U$24470 ( \30130 , \8458 , \29785 );
and \U$24471 ( \30131 , \8460 , \29812 );
and \U$24472 ( \30132 , \8462 , \29839 );
and \U$24473 ( \30133 , \8464 , \29866 );
and \U$24474 ( \30134 , \8466 , \29893 );
and \U$24475 ( \30135 , \8468 , \29920 );
and \U$24476 ( \30136 , \8470 , \29947 );
and \U$24477 ( \30137 , \8472 , \29974 );
or \U$24478 ( \30138 , \30122 , \30123 , \30124 , \30125 , \30126 , \30127 , \30128 , \30129 , \30130 , \30131 , \30132 , \30133 , \30134 , \30135 , \30136 , \30137 );
_DC g8cc4 ( \30139_nG8cc4 , \30138 , \30051 );
buf \U$24479 ( \30140 , \30139_nG8cc4 );
xor \U$24480 ( \30141 , \30121 , \30140 );
or \U$24481 ( \30142 , \30120 , \30141 );
buf \U$24482 ( \30143 , RIb7b93b0_251);
and \U$24483 ( \30144 , \7166 , \29569 );
and \U$24484 ( \30145 , \7168 , \29596 );
and \U$24485 ( \30146 , \8482 , \29623 );
and \U$24486 ( \30147 , \8484 , \29650 );
and \U$24487 ( \30148 , \8486 , \29677 );
and \U$24488 ( \30149 , \8488 , \29704 );
and \U$24489 ( \30150 , \8490 , \29731 );
and \U$24490 ( \30151 , \8492 , \29758 );
and \U$24491 ( \30152 , \8494 , \29785 );
and \U$24492 ( \30153 , \8496 , \29812 );
and \U$24493 ( \30154 , \8498 , \29839 );
and \U$24494 ( \30155 , \8500 , \29866 );
and \U$24495 ( \30156 , \8502 , \29893 );
and \U$24496 ( \30157 , \8504 , \29920 );
and \U$24497 ( \30158 , \8506 , \29947 );
and \U$24498 ( \30159 , \8508 , \29974 );
or \U$24499 ( \30160 , \30144 , \30145 , \30146 , \30147 , \30148 , \30149 , \30150 , \30151 , \30152 , \30153 , \30154 , \30155 , \30156 , \30157 , \30158 , \30159 );
_DC g8cda ( \30161_nG8cda , \30160 , \30051 );
buf \U$24500 ( \30162 , \30161_nG8cda );
xor \U$24501 ( \30163 , \30143 , \30162 );
or \U$24502 ( \30164 , \30142 , \30163 );
buf \U$24503 ( \30165 , RIb7af720_252);
and \U$24504 ( \30166 , \7176 , \29569 );
and \U$24505 ( \30167 , \7178 , \29596 );
and \U$24506 ( \30168 , \8518 , \29623 );
and \U$24507 ( \30169 , \8520 , \29650 );
and \U$24508 ( \30170 , \8522 , \29677 );
and \U$24509 ( \30171 , \8524 , \29704 );
and \U$24510 ( \30172 , \8526 , \29731 );
and \U$24511 ( \30173 , \8528 , \29758 );
and \U$24512 ( \30174 , \8530 , \29785 );
and \U$24513 ( \30175 , \8532 , \29812 );
and \U$24514 ( \30176 , \8534 , \29839 );
and \U$24515 ( \30177 , \8536 , \29866 );
and \U$24516 ( \30178 , \8538 , \29893 );
and \U$24517 ( \30179 , \8540 , \29920 );
and \U$24518 ( \30180 , \8542 , \29947 );
and \U$24519 ( \30181 , \8544 , \29974 );
or \U$24520 ( \30182 , \30166 , \30167 , \30168 , \30169 , \30170 , \30171 , \30172 , \30173 , \30174 , \30175 , \30176 , \30177 , \30178 , \30179 , \30180 , \30181 );
_DC g8cf0 ( \30183_nG8cf0 , \30182 , \30051 );
buf \U$24521 ( \30184 , \30183_nG8cf0 );
xor \U$24522 ( \30185 , \30165 , \30184 );
or \U$24523 ( \30186 , \30164 , \30185 );
buf \U$24524 ( \30187 , RIb7af6a8_253);
and \U$24525 ( \30188 , \7186 , \29569 );
and \U$24526 ( \30189 , \7188 , \29596 );
and \U$24527 ( \30190 , \8554 , \29623 );
and \U$24528 ( \30191 , \8556 , \29650 );
and \U$24529 ( \30192 , \8558 , \29677 );
and \U$24530 ( \30193 , \8560 , \29704 );
and \U$24531 ( \30194 , \8562 , \29731 );
and \U$24532 ( \30195 , \8564 , \29758 );
and \U$24533 ( \30196 , \8566 , \29785 );
and \U$24534 ( \30197 , \8568 , \29812 );
and \U$24535 ( \30198 , \8570 , \29839 );
and \U$24536 ( \30199 , \8572 , \29866 );
and \U$24537 ( \30200 , \8574 , \29893 );
and \U$24538 ( \30201 , \8576 , \29920 );
and \U$24539 ( \30202 , \8578 , \29947 );
and \U$24540 ( \30203 , \8580 , \29974 );
or \U$24541 ( \30204 , \30188 , \30189 , \30190 , \30191 , \30192 , \30193 , \30194 , \30195 , \30196 , \30197 , \30198 , \30199 , \30200 , \30201 , \30202 , \30203 );
_DC g8d06 ( \30205_nG8d06 , \30204 , \30051 );
buf \U$24542 ( \30206 , \30205_nG8d06 );
xor \U$24543 ( \30207 , \30187 , \30206 );
or \U$24544 ( \30208 , \30186 , \30207 );
not \U$24545 ( \30209 , \30208 );
buf \U$24546 ( \30210 , \30209 );
and \U$24547 ( \30211 , \29542 , \30210 );
buf \U$24548 ( \30212 , RIb7af630_254);
buf \U$24549 ( \30213 , \29028 );
buf \U$24550 ( \30214 , \29028 );
buf \U$24551 ( \30215 , \29028 );
buf \U$24552 ( \30216 , \29028 );
buf \U$24553 ( \30217 , \29028 );
buf \U$24554 ( \30218 , \29028 );
buf \U$24555 ( \30219 , \29028 );
buf \U$24556 ( \30220 , \29028 );
buf \U$24557 ( \30221 , \29028 );
buf \U$24558 ( \30222 , \29028 );
buf \U$24559 ( \30223 , \29028 );
buf \U$24560 ( \30224 , \29028 );
buf \U$24561 ( \30225 , \29028 );
buf \U$24562 ( \30226 , \29028 );
buf \U$24563 ( \30227 , \29028 );
buf \U$24564 ( \30228 , \29028 );
buf \U$24565 ( \30229 , \29028 );
buf \U$24566 ( \30230 , \29028 );
buf \U$24567 ( \30231 , \29028 );
buf \U$24568 ( \30232 , \29028 );
buf \U$24569 ( \30233 , \29028 );
buf \U$24570 ( \30234 , \29028 );
buf \U$24571 ( \30235 , \29028 );
buf \U$24572 ( \30236 , \29028 );
buf \U$24573 ( \30237 , \29028 );
nor \U$24574 ( \30238 , \29015 , \29016 , \29017 , \29018 , \29022 , \29025 , \29028 , \30213 , \30214 , \30215 , \30216 , \30217 , \30218 , \30219 , \30220 , \30221 , \30222 , \30223 , \30224 , \30225 , \30226 , \30227 , \30228 , \30229 , \30230 , \30231 , \30232 , \30233 , \30234 , \30235 , \30236 , \30237 );
and \U$24575 ( \30239 , \7198 , \30238 );
buf \U$24576 ( \30240 , \29028 );
buf \U$24577 ( \30241 , \29028 );
buf \U$24578 ( \30242 , \29028 );
buf \U$24579 ( \30243 , \29028 );
buf \U$24580 ( \30244 , \29028 );
buf \U$24581 ( \30245 , \29028 );
buf \U$24582 ( \30246 , \29028 );
buf \U$24583 ( \30247 , \29028 );
buf \U$24584 ( \30248 , \29028 );
buf \U$24585 ( \30249 , \29028 );
buf \U$24586 ( \30250 , \29028 );
buf \U$24587 ( \30251 , \29028 );
buf \U$24588 ( \30252 , \29028 );
buf \U$24589 ( \30253 , \29028 );
buf \U$24590 ( \30254 , \29028 );
buf \U$24591 ( \30255 , \29028 );
buf \U$24592 ( \30256 , \29028 );
buf \U$24593 ( \30257 , \29028 );
buf \U$24594 ( \30258 , \29028 );
buf \U$24595 ( \30259 , \29028 );
buf \U$24596 ( \30260 , \29028 );
buf \U$24597 ( \30261 , \29028 );
buf \U$24598 ( \30262 , \29028 );
buf \U$24599 ( \30263 , \29028 );
buf \U$24600 ( \30264 , \29028 );
nor \U$24601 ( \30265 , \29056 , \29057 , \29058 , \29059 , \29021 , \29025 , \29028 , \30240 , \30241 , \30242 , \30243 , \30244 , \30245 , \30246 , \30247 , \30248 , \30249 , \30250 , \30251 , \30252 , \30253 , \30254 , \30255 , \30256 , \30257 , \30258 , \30259 , \30260 , \30261 , \30262 , \30263 , \30264 );
and \U$24602 ( \30266 , \7200 , \30265 );
buf \U$24603 ( \30267 , \29028 );
buf \U$24604 ( \30268 , \29028 );
buf \U$24605 ( \30269 , \29028 );
buf \U$24606 ( \30270 , \29028 );
buf \U$24607 ( \30271 , \29028 );
buf \U$24608 ( \30272 , \29028 );
buf \U$24609 ( \30273 , \29028 );
buf \U$24610 ( \30274 , \29028 );
buf \U$24611 ( \30275 , \29028 );
buf \U$24612 ( \30276 , \29028 );
buf \U$24613 ( \30277 , \29028 );
buf \U$24614 ( \30278 , \29028 );
buf \U$24615 ( \30279 , \29028 );
buf \U$24616 ( \30280 , \29028 );
buf \U$24617 ( \30281 , \29028 );
buf \U$24618 ( \30282 , \29028 );
buf \U$24619 ( \30283 , \29028 );
buf \U$24620 ( \30284 , \29028 );
buf \U$24621 ( \30285 , \29028 );
buf \U$24622 ( \30286 , \29028 );
buf \U$24623 ( \30287 , \29028 );
buf \U$24624 ( \30288 , \29028 );
buf \U$24625 ( \30289 , \29028 );
buf \U$24626 ( \30290 , \29028 );
buf \U$24627 ( \30291 , \29028 );
nor \U$24628 ( \30292 , \29015 , \29057 , \29058 , \29059 , \29021 , \29025 , \29028 , \30267 , \30268 , \30269 , \30270 , \30271 , \30272 , \30273 , \30274 , \30275 , \30276 , \30277 , \30278 , \30279 , \30280 , \30281 , \30282 , \30283 , \30284 , \30285 , \30286 , \30287 , \30288 , \30289 , \30290 , \30291 );
and \U$24629 ( \30293 , \8645 , \30292 );
buf \U$24630 ( \30294 , \29028 );
buf \U$24631 ( \30295 , \29028 );
buf \U$24632 ( \30296 , \29028 );
buf \U$24633 ( \30297 , \29028 );
buf \U$24634 ( \30298 , \29028 );
buf \U$24635 ( \30299 , \29028 );
buf \U$24636 ( \30300 , \29028 );
buf \U$24637 ( \30301 , \29028 );
buf \U$24638 ( \30302 , \29028 );
buf \U$24639 ( \30303 , \29028 );
buf \U$24640 ( \30304 , \29028 );
buf \U$24641 ( \30305 , \29028 );
buf \U$24642 ( \30306 , \29028 );
buf \U$24643 ( \30307 , \29028 );
buf \U$24644 ( \30308 , \29028 );
buf \U$24645 ( \30309 , \29028 );
buf \U$24646 ( \30310 , \29028 );
buf \U$24647 ( \30311 , \29028 );
buf \U$24648 ( \30312 , \29028 );
buf \U$24649 ( \30313 , \29028 );
buf \U$24650 ( \30314 , \29028 );
buf \U$24651 ( \30315 , \29028 );
buf \U$24652 ( \30316 , \29028 );
buf \U$24653 ( \30317 , \29028 );
buf \U$24654 ( \30318 , \29028 );
nor \U$24655 ( \30319 , \29056 , \29016 , \29058 , \29059 , \29021 , \29025 , \29028 , \30294 , \30295 , \30296 , \30297 , \30298 , \30299 , \30300 , \30301 , \30302 , \30303 , \30304 , \30305 , \30306 , \30307 , \30308 , \30309 , \30310 , \30311 , \30312 , \30313 , \30314 , \30315 , \30316 , \30317 , \30318 );
and \U$24656 ( \30320 , \8673 , \30319 );
buf \U$24657 ( \30321 , \29028 );
buf \U$24658 ( \30322 , \29028 );
buf \U$24659 ( \30323 , \29028 );
buf \U$24660 ( \30324 , \29028 );
buf \U$24661 ( \30325 , \29028 );
buf \U$24662 ( \30326 , \29028 );
buf \U$24663 ( \30327 , \29028 );
buf \U$24664 ( \30328 , \29028 );
buf \U$24665 ( \30329 , \29028 );
buf \U$24666 ( \30330 , \29028 );
buf \U$24667 ( \30331 , \29028 );
buf \U$24668 ( \30332 , \29028 );
buf \U$24669 ( \30333 , \29028 );
buf \U$24670 ( \30334 , \29028 );
buf \U$24671 ( \30335 , \29028 );
buf \U$24672 ( \30336 , \29028 );
buf \U$24673 ( \30337 , \29028 );
buf \U$24674 ( \30338 , \29028 );
buf \U$24675 ( \30339 , \29028 );
buf \U$24676 ( \30340 , \29028 );
buf \U$24677 ( \30341 , \29028 );
buf \U$24678 ( \30342 , \29028 );
buf \U$24679 ( \30343 , \29028 );
buf \U$24680 ( \30344 , \29028 );
buf \U$24681 ( \30345 , \29028 );
nor \U$24682 ( \30346 , \29015 , \29016 , \29058 , \29059 , \29021 , \29025 , \29028 , \30321 , \30322 , \30323 , \30324 , \30325 , \30326 , \30327 , \30328 , \30329 , \30330 , \30331 , \30332 , \30333 , \30334 , \30335 , \30336 , \30337 , \30338 , \30339 , \30340 , \30341 , \30342 , \30343 , \30344 , \30345 );
and \U$24683 ( \30347 , \8701 , \30346 );
buf \U$24684 ( \30348 , \29028 );
buf \U$24685 ( \30349 , \29028 );
buf \U$24686 ( \30350 , \29028 );
buf \U$24687 ( \30351 , \29028 );
buf \U$24688 ( \30352 , \29028 );
buf \U$24689 ( \30353 , \29028 );
buf \U$24690 ( \30354 , \29028 );
buf \U$24691 ( \30355 , \29028 );
buf \U$24692 ( \30356 , \29028 );
buf \U$24693 ( \30357 , \29028 );
buf \U$24694 ( \30358 , \29028 );
buf \U$24695 ( \30359 , \29028 );
buf \U$24696 ( \30360 , \29028 );
buf \U$24697 ( \30361 , \29028 );
buf \U$24698 ( \30362 , \29028 );
buf \U$24699 ( \30363 , \29028 );
buf \U$24700 ( \30364 , \29028 );
buf \U$24701 ( \30365 , \29028 );
buf \U$24702 ( \30366 , \29028 );
buf \U$24703 ( \30367 , \29028 );
buf \U$24704 ( \30368 , \29028 );
buf \U$24705 ( \30369 , \29028 );
buf \U$24706 ( \30370 , \29028 );
buf \U$24707 ( \30371 , \29028 );
buf \U$24708 ( \30372 , \29028 );
nor \U$24709 ( \30373 , \29056 , \29057 , \29017 , \29059 , \29021 , \29025 , \29028 , \30348 , \30349 , \30350 , \30351 , \30352 , \30353 , \30354 , \30355 , \30356 , \30357 , \30358 , \30359 , \30360 , \30361 , \30362 , \30363 , \30364 , \30365 , \30366 , \30367 , \30368 , \30369 , \30370 , \30371 , \30372 );
and \U$24710 ( \30374 , \8729 , \30373 );
buf \U$24711 ( \30375 , \29028 );
buf \U$24712 ( \30376 , \29028 );
buf \U$24713 ( \30377 , \29028 );
buf \U$24714 ( \30378 , \29028 );
buf \U$24715 ( \30379 , \29028 );
buf \U$24716 ( \30380 , \29028 );
buf \U$24717 ( \30381 , \29028 );
buf \U$24718 ( \30382 , \29028 );
buf \U$24719 ( \30383 , \29028 );
buf \U$24720 ( \30384 , \29028 );
buf \U$24721 ( \30385 , \29028 );
buf \U$24722 ( \30386 , \29028 );
buf \U$24723 ( \30387 , \29028 );
buf \U$24724 ( \30388 , \29028 );
buf \U$24725 ( \30389 , \29028 );
buf \U$24726 ( \30390 , \29028 );
buf \U$24727 ( \30391 , \29028 );
buf \U$24728 ( \30392 , \29028 );
buf \U$24729 ( \30393 , \29028 );
buf \U$24730 ( \30394 , \29028 );
buf \U$24731 ( \30395 , \29028 );
buf \U$24732 ( \30396 , \29028 );
buf \U$24733 ( \30397 , \29028 );
buf \U$24734 ( \30398 , \29028 );
buf \U$24735 ( \30399 , \29028 );
nor \U$24736 ( \30400 , \29015 , \29057 , \29017 , \29059 , \29021 , \29025 , \29028 , \30375 , \30376 , \30377 , \30378 , \30379 , \30380 , \30381 , \30382 , \30383 , \30384 , \30385 , \30386 , \30387 , \30388 , \30389 , \30390 , \30391 , \30392 , \30393 , \30394 , \30395 , \30396 , \30397 , \30398 , \30399 );
and \U$24737 ( \30401 , \8757 , \30400 );
buf \U$24738 ( \30402 , \29028 );
buf \U$24739 ( \30403 , \29028 );
buf \U$24740 ( \30404 , \29028 );
buf \U$24741 ( \30405 , \29028 );
buf \U$24742 ( \30406 , \29028 );
buf \U$24743 ( \30407 , \29028 );
buf \U$24744 ( \30408 , \29028 );
buf \U$24745 ( \30409 , \29028 );
buf \U$24746 ( \30410 , \29028 );
buf \U$24747 ( \30411 , \29028 );
buf \U$24748 ( \30412 , \29028 );
buf \U$24749 ( \30413 , \29028 );
buf \U$24750 ( \30414 , \29028 );
buf \U$24751 ( \30415 , \29028 );
buf \U$24752 ( \30416 , \29028 );
buf \U$24753 ( \30417 , \29028 );
buf \U$24754 ( \30418 , \29028 );
buf \U$24755 ( \30419 , \29028 );
buf \U$24756 ( \30420 , \29028 );
buf \U$24757 ( \30421 , \29028 );
buf \U$24758 ( \30422 , \29028 );
buf \U$24759 ( \30423 , \29028 );
buf \U$24760 ( \30424 , \29028 );
buf \U$24761 ( \30425 , \29028 );
buf \U$24762 ( \30426 , \29028 );
nor \U$24763 ( \30427 , \29056 , \29016 , \29017 , \29059 , \29021 , \29025 , \29028 , \30402 , \30403 , \30404 , \30405 , \30406 , \30407 , \30408 , \30409 , \30410 , \30411 , \30412 , \30413 , \30414 , \30415 , \30416 , \30417 , \30418 , \30419 , \30420 , \30421 , \30422 , \30423 , \30424 , \30425 , \30426 );
and \U$24764 ( \30428 , \8785 , \30427 );
buf \U$24765 ( \30429 , \29028 );
buf \U$24766 ( \30430 , \29028 );
buf \U$24767 ( \30431 , \29028 );
buf \U$24768 ( \30432 , \29028 );
buf \U$24769 ( \30433 , \29028 );
buf \U$24770 ( \30434 , \29028 );
buf \U$24771 ( \30435 , \29028 );
buf \U$24772 ( \30436 , \29028 );
buf \U$24773 ( \30437 , \29028 );
buf \U$24774 ( \30438 , \29028 );
buf \U$24775 ( \30439 , \29028 );
buf \U$24776 ( \30440 , \29028 );
buf \U$24777 ( \30441 , \29028 );
buf \U$24778 ( \30442 , \29028 );
buf \U$24779 ( \30443 , \29028 );
buf \U$24780 ( \30444 , \29028 );
buf \U$24781 ( \30445 , \29028 );
buf \U$24782 ( \30446 , \29028 );
buf \U$24783 ( \30447 , \29028 );
buf \U$24784 ( \30448 , \29028 );
buf \U$24785 ( \30449 , \29028 );
buf \U$24786 ( \30450 , \29028 );
buf \U$24787 ( \30451 , \29028 );
buf \U$24788 ( \30452 , \29028 );
buf \U$24789 ( \30453 , \29028 );
nor \U$24790 ( \30454 , \29015 , \29016 , \29017 , \29059 , \29021 , \29025 , \29028 , \30429 , \30430 , \30431 , \30432 , \30433 , \30434 , \30435 , \30436 , \30437 , \30438 , \30439 , \30440 , \30441 , \30442 , \30443 , \30444 , \30445 , \30446 , \30447 , \30448 , \30449 , \30450 , \30451 , \30452 , \30453 );
and \U$24791 ( \30455 , \8813 , \30454 );
buf \U$24792 ( \30456 , \29028 );
buf \U$24793 ( \30457 , \29028 );
buf \U$24794 ( \30458 , \29028 );
buf \U$24795 ( \30459 , \29028 );
buf \U$24796 ( \30460 , \29028 );
buf \U$24797 ( \30461 , \29028 );
buf \U$24798 ( \30462 , \29028 );
buf \U$24799 ( \30463 , \29028 );
buf \U$24800 ( \30464 , \29028 );
buf \U$24801 ( \30465 , \29028 );
buf \U$24802 ( \30466 , \29028 );
buf \U$24803 ( \30467 , \29028 );
buf \U$24804 ( \30468 , \29028 );
buf \U$24805 ( \30469 , \29028 );
buf \U$24806 ( \30470 , \29028 );
buf \U$24807 ( \30471 , \29028 );
buf \U$24808 ( \30472 , \29028 );
buf \U$24809 ( \30473 , \29028 );
buf \U$24810 ( \30474 , \29028 );
buf \U$24811 ( \30475 , \29028 );
buf \U$24812 ( \30476 , \29028 );
buf \U$24813 ( \30477 , \29028 );
buf \U$24814 ( \30478 , \29028 );
buf \U$24815 ( \30479 , \29028 );
buf \U$24816 ( \30480 , \29028 );
nor \U$24817 ( \30481 , \29056 , \29057 , \29058 , \29018 , \29021 , \29025 , \29028 , \30456 , \30457 , \30458 , \30459 , \30460 , \30461 , \30462 , \30463 , \30464 , \30465 , \30466 , \30467 , \30468 , \30469 , \30470 , \30471 , \30472 , \30473 , \30474 , \30475 , \30476 , \30477 , \30478 , \30479 , \30480 );
and \U$24818 ( \30482 , \8841 , \30481 );
buf \U$24819 ( \30483 , \29028 );
buf \U$24820 ( \30484 , \29028 );
buf \U$24821 ( \30485 , \29028 );
buf \U$24822 ( \30486 , \29028 );
buf \U$24823 ( \30487 , \29028 );
buf \U$24824 ( \30488 , \29028 );
buf \U$24825 ( \30489 , \29028 );
buf \U$24826 ( \30490 , \29028 );
buf \U$24827 ( \30491 , \29028 );
buf \U$24828 ( \30492 , \29028 );
buf \U$24829 ( \30493 , \29028 );
buf \U$24830 ( \30494 , \29028 );
buf \U$24831 ( \30495 , \29028 );
buf \U$24832 ( \30496 , \29028 );
buf \U$24833 ( \30497 , \29028 );
buf \U$24834 ( \30498 , \29028 );
buf \U$24835 ( \30499 , \29028 );
buf \U$24836 ( \30500 , \29028 );
buf \U$24837 ( \30501 , \29028 );
buf \U$24838 ( \30502 , \29028 );
buf \U$24839 ( \30503 , \29028 );
buf \U$24840 ( \30504 , \29028 );
buf \U$24841 ( \30505 , \29028 );
buf \U$24842 ( \30506 , \29028 );
buf \U$24843 ( \30507 , \29028 );
nor \U$24844 ( \30508 , \29015 , \29057 , \29058 , \29018 , \29021 , \29025 , \29028 , \30483 , \30484 , \30485 , \30486 , \30487 , \30488 , \30489 , \30490 , \30491 , \30492 , \30493 , \30494 , \30495 , \30496 , \30497 , \30498 , \30499 , \30500 , \30501 , \30502 , \30503 , \30504 , \30505 , \30506 , \30507 );
and \U$24845 ( \30509 , \8869 , \30508 );
buf \U$24846 ( \30510 , \29028 );
buf \U$24847 ( \30511 , \29028 );
buf \U$24848 ( \30512 , \29028 );
buf \U$24849 ( \30513 , \29028 );
buf \U$24850 ( \30514 , \29028 );
buf \U$24851 ( \30515 , \29028 );
buf \U$24852 ( \30516 , \29028 );
buf \U$24853 ( \30517 , \29028 );
buf \U$24854 ( \30518 , \29028 );
buf \U$24855 ( \30519 , \29028 );
buf \U$24856 ( \30520 , \29028 );
buf \U$24857 ( \30521 , \29028 );
buf \U$24858 ( \30522 , \29028 );
buf \U$24859 ( \30523 , \29028 );
buf \U$24860 ( \30524 , \29028 );
buf \U$24861 ( \30525 , \29028 );
buf \U$24862 ( \30526 , \29028 );
buf \U$24863 ( \30527 , \29028 );
buf \U$24864 ( \30528 , \29028 );
buf \U$24865 ( \30529 , \29028 );
buf \U$24866 ( \30530 , \29028 );
buf \U$24867 ( \30531 , \29028 );
buf \U$24868 ( \30532 , \29028 );
buf \U$24869 ( \30533 , \29028 );
buf \U$24870 ( \30534 , \29028 );
nor \U$24871 ( \30535 , \29056 , \29016 , \29058 , \29018 , \29021 , \29025 , \29028 , \30510 , \30511 , \30512 , \30513 , \30514 , \30515 , \30516 , \30517 , \30518 , \30519 , \30520 , \30521 , \30522 , \30523 , \30524 , \30525 , \30526 , \30527 , \30528 , \30529 , \30530 , \30531 , \30532 , \30533 , \30534 );
and \U$24872 ( \30536 , \8897 , \30535 );
buf \U$24873 ( \30537 , \29028 );
buf \U$24874 ( \30538 , \29028 );
buf \U$24875 ( \30539 , \29028 );
buf \U$24876 ( \30540 , \29028 );
buf \U$24877 ( \30541 , \29028 );
buf \U$24878 ( \30542 , \29028 );
buf \U$24879 ( \30543 , \29028 );
buf \U$24880 ( \30544 , \29028 );
buf \U$24881 ( \30545 , \29028 );
buf \U$24882 ( \30546 , \29028 );
buf \U$24883 ( \30547 , \29028 );
buf \U$24884 ( \30548 , \29028 );
buf \U$24885 ( \30549 , \29028 );
buf \U$24886 ( \30550 , \29028 );
buf \U$24887 ( \30551 , \29028 );
buf \U$24888 ( \30552 , \29028 );
buf \U$24889 ( \30553 , \29028 );
buf \U$24890 ( \30554 , \29028 );
buf \U$24891 ( \30555 , \29028 );
buf \U$24892 ( \30556 , \29028 );
buf \U$24893 ( \30557 , \29028 );
buf \U$24894 ( \30558 , \29028 );
buf \U$24895 ( \30559 , \29028 );
buf \U$24896 ( \30560 , \29028 );
buf \U$24897 ( \30561 , \29028 );
nor \U$24898 ( \30562 , \29015 , \29016 , \29058 , \29018 , \29021 , \29025 , \29028 , \30537 , \30538 , \30539 , \30540 , \30541 , \30542 , \30543 , \30544 , \30545 , \30546 , \30547 , \30548 , \30549 , \30550 , \30551 , \30552 , \30553 , \30554 , \30555 , \30556 , \30557 , \30558 , \30559 , \30560 , \30561 );
and \U$24899 ( \30563 , \8925 , \30562 );
buf \U$24900 ( \30564 , \29028 );
buf \U$24901 ( \30565 , \29028 );
buf \U$24902 ( \30566 , \29028 );
buf \U$24903 ( \30567 , \29028 );
buf \U$24904 ( \30568 , \29028 );
buf \U$24905 ( \30569 , \29028 );
buf \U$24906 ( \30570 , \29028 );
buf \U$24907 ( \30571 , \29028 );
buf \U$24908 ( \30572 , \29028 );
buf \U$24909 ( \30573 , \29028 );
buf \U$24910 ( \30574 , \29028 );
buf \U$24911 ( \30575 , \29028 );
buf \U$24912 ( \30576 , \29028 );
buf \U$24913 ( \30577 , \29028 );
buf \U$24914 ( \30578 , \29028 );
buf \U$24915 ( \30579 , \29028 );
buf \U$24916 ( \30580 , \29028 );
buf \U$24917 ( \30581 , \29028 );
buf \U$24918 ( \30582 , \29028 );
buf \U$24919 ( \30583 , \29028 );
buf \U$24920 ( \30584 , \29028 );
buf \U$24921 ( \30585 , \29028 );
buf \U$24922 ( \30586 , \29028 );
buf \U$24923 ( \30587 , \29028 );
buf \U$24924 ( \30588 , \29028 );
nor \U$24925 ( \30589 , \29056 , \29057 , \29017 , \29018 , \29021 , \29025 , \29028 , \30564 , \30565 , \30566 , \30567 , \30568 , \30569 , \30570 , \30571 , \30572 , \30573 , \30574 , \30575 , \30576 , \30577 , \30578 , \30579 , \30580 , \30581 , \30582 , \30583 , \30584 , \30585 , \30586 , \30587 , \30588 );
and \U$24926 ( \30590 , \8953 , \30589 );
buf \U$24927 ( \30591 , \29028 );
buf \U$24928 ( \30592 , \29028 );
buf \U$24929 ( \30593 , \29028 );
buf \U$24930 ( \30594 , \29028 );
buf \U$24931 ( \30595 , \29028 );
buf \U$24932 ( \30596 , \29028 );
buf \U$24933 ( \30597 , \29028 );
buf \U$24934 ( \30598 , \29028 );
buf \U$24935 ( \30599 , \29028 );
buf \U$24936 ( \30600 , \29028 );
buf \U$24937 ( \30601 , \29028 );
buf \U$24938 ( \30602 , \29028 );
buf \U$24939 ( \30603 , \29028 );
buf \U$24940 ( \30604 , \29028 );
buf \U$24941 ( \30605 , \29028 );
buf \U$24942 ( \30606 , \29028 );
buf \U$24943 ( \30607 , \29028 );
buf \U$24944 ( \30608 , \29028 );
buf \U$24945 ( \30609 , \29028 );
buf \U$24946 ( \30610 , \29028 );
buf \U$24947 ( \30611 , \29028 );
buf \U$24948 ( \30612 , \29028 );
buf \U$24949 ( \30613 , \29028 );
buf \U$24950 ( \30614 , \29028 );
buf \U$24951 ( \30615 , \29028 );
nor \U$24952 ( \30616 , \29015 , \29057 , \29017 , \29018 , \29021 , \29025 , \29028 , \30591 , \30592 , \30593 , \30594 , \30595 , \30596 , \30597 , \30598 , \30599 , \30600 , \30601 , \30602 , \30603 , \30604 , \30605 , \30606 , \30607 , \30608 , \30609 , \30610 , \30611 , \30612 , \30613 , \30614 , \30615 );
and \U$24953 ( \30617 , \8981 , \30616 );
buf \U$24954 ( \30618 , \29028 );
buf \U$24955 ( \30619 , \29028 );
buf \U$24956 ( \30620 , \29028 );
buf \U$24957 ( \30621 , \29028 );
buf \U$24958 ( \30622 , \29028 );
buf \U$24959 ( \30623 , \29028 );
buf \U$24960 ( \30624 , \29028 );
buf \U$24961 ( \30625 , \29028 );
buf \U$24962 ( \30626 , \29028 );
buf \U$24963 ( \30627 , \29028 );
buf \U$24964 ( \30628 , \29028 );
buf \U$24965 ( \30629 , \29028 );
buf \U$24966 ( \30630 , \29028 );
buf \U$24967 ( \30631 , \29028 );
buf \U$24968 ( \30632 , \29028 );
buf \U$24969 ( \30633 , \29028 );
buf \U$24970 ( \30634 , \29028 );
buf \U$24971 ( \30635 , \29028 );
buf \U$24972 ( \30636 , \29028 );
buf \U$24973 ( \30637 , \29028 );
buf \U$24974 ( \30638 , \29028 );
buf \U$24975 ( \30639 , \29028 );
buf \U$24976 ( \30640 , \29028 );
buf \U$24977 ( \30641 , \29028 );
buf \U$24978 ( \30642 , \29028 );
nor \U$24979 ( \30643 , \29056 , \29016 , \29017 , \29018 , \29021 , \29025 , \29028 , \30618 , \30619 , \30620 , \30621 , \30622 , \30623 , \30624 , \30625 , \30626 , \30627 , \30628 , \30629 , \30630 , \30631 , \30632 , \30633 , \30634 , \30635 , \30636 , \30637 , \30638 , \30639 , \30640 , \30641 , \30642 );
and \U$24980 ( \30644 , \9009 , \30643 );
or \U$24981 ( \30645 , \30239 , \30266 , \30293 , \30320 , \30347 , \30374 , \30401 , \30428 , \30455 , \30482 , \30509 , \30536 , \30563 , \30590 , \30617 , \30644 );
buf \U$24982 ( \30646 , \29028 );
not \U$24983 ( \30647 , \30646 );
buf \U$24984 ( \30648 , \29016 );
buf \U$24985 ( \30649 , \29017 );
buf \U$24986 ( \30650 , \29018 );
buf \U$24987 ( \30651 , \29021 );
buf \U$24988 ( \30652 , \29025 );
buf \U$24989 ( \30653 , \29028 );
buf \U$24990 ( \30654 , \29028 );
buf \U$24991 ( \30655 , \29028 );
buf \U$24992 ( \30656 , \29028 );
buf \U$24993 ( \30657 , \29028 );
buf \U$24994 ( \30658 , \29028 );
buf \U$24995 ( \30659 , \29028 );
buf \U$24996 ( \30660 , \29028 );
buf \U$24997 ( \30661 , \29028 );
buf \U$24998 ( \30662 , \29028 );
buf \U$24999 ( \30663 , \29028 );
buf \U$25000 ( \30664 , \29028 );
buf \U$25001 ( \30665 , \29028 );
buf \U$25002 ( \30666 , \29028 );
buf \U$25003 ( \30667 , \29028 );
buf \U$25004 ( \30668 , \29028 );
buf \U$25005 ( \30669 , \29028 );
buf \U$25006 ( \30670 , \29028 );
buf \U$25007 ( \30671 , \29028 );
buf \U$25008 ( \30672 , \29028 );
buf \U$25009 ( \30673 , \29028 );
buf \U$25010 ( \30674 , \29028 );
buf \U$25011 ( \30675 , \29028 );
buf \U$25012 ( \30676 , \29028 );
buf \U$25013 ( \30677 , \29028 );
buf \U$25014 ( \30678 , \29015 );
or \U$25015 ( \30679 , \30648 , \30649 , \30650 , \30651 , \30652 , \30653 , \30654 , \30655 , \30656 , \30657 , \30658 , \30659 , \30660 , \30661 , \30662 , \30663 , \30664 , \30665 , \30666 , \30667 , \30668 , \30669 , \30670 , \30671 , \30672 , \30673 , \30674 , \30675 , \30676 , \30677 , \30678 );
nand \U$25016 ( \30680 , \30647 , \30679 );
buf \U$25017 ( \30681 , \30680 );
buf \U$25018 ( \30682 , \29028 );
not \U$25019 ( \30683 , \30682 );
buf \U$25020 ( \30684 , \29025 );
buf \U$25021 ( \30685 , \29028 );
buf \U$25022 ( \30686 , \29028 );
buf \U$25023 ( \30687 , \29028 );
buf \U$25024 ( \30688 , \29028 );
buf \U$25025 ( \30689 , \29028 );
buf \U$25026 ( \30690 , \29028 );
buf \U$25027 ( \30691 , \29028 );
buf \U$25028 ( \30692 , \29028 );
buf \U$25029 ( \30693 , \29028 );
buf \U$25030 ( \30694 , \29028 );
buf \U$25031 ( \30695 , \29028 );
buf \U$25032 ( \30696 , \29028 );
buf \U$25033 ( \30697 , \29028 );
buf \U$25034 ( \30698 , \29028 );
buf \U$25035 ( \30699 , \29028 );
buf \U$25036 ( \30700 , \29028 );
buf \U$25037 ( \30701 , \29028 );
buf \U$25038 ( \30702 , \29028 );
buf \U$25039 ( \30703 , \29028 );
buf \U$25040 ( \30704 , \29028 );
buf \U$25041 ( \30705 , \29028 );
buf \U$25042 ( \30706 , \29028 );
buf \U$25043 ( \30707 , \29028 );
buf \U$25044 ( \30708 , \29028 );
buf \U$25045 ( \30709 , \29028 );
buf \U$25046 ( \30710 , \29021 );
buf \U$25047 ( \30711 , \29015 );
buf \U$25048 ( \30712 , \29016 );
buf \U$25049 ( \30713 , \29017 );
buf \U$25050 ( \30714 , \29018 );
or \U$25051 ( \30715 , \30711 , \30712 , \30713 , \30714 );
and \U$25052 ( \30716 , \30710 , \30715 );
or \U$25053 ( \30717 , \30684 , \30685 , \30686 , \30687 , \30688 , \30689 , \30690 , \30691 , \30692 , \30693 , \30694 , \30695 , \30696 , \30697 , \30698 , \30699 , \30700 , \30701 , \30702 , \30703 , \30704 , \30705 , \30706 , \30707 , \30708 , \30709 , \30716 );
and \U$25054 ( \30718 , \30683 , \30717 );
buf \U$25055 ( \30719 , \30718 );
or \U$25056 ( \30720 , \30681 , \30719 );
_DC g8f0a ( \30721_nG8f0a , \30645 , \30720 );
buf \U$25057 ( \30722 , \30721_nG8f0a );
xor \U$25058 ( \30723 , \30212 , \30722 );
buf \U$25059 ( \30724 , RIb7af5b8_255);
and \U$25060 ( \30725 , \7207 , \30238 );
and \U$25061 ( \30726 , \7209 , \30265 );
and \U$25062 ( \30727 , \9119 , \30292 );
and \U$25063 ( \30728 , \9121 , \30319 );
and \U$25064 ( \30729 , \9123 , \30346 );
and \U$25065 ( \30730 , \9125 , \30373 );
and \U$25066 ( \30731 , \9127 , \30400 );
and \U$25067 ( \30732 , \9129 , \30427 );
and \U$25068 ( \30733 , \9131 , \30454 );
and \U$25069 ( \30734 , \9133 , \30481 );
and \U$25070 ( \30735 , \9135 , \30508 );
and \U$25071 ( \30736 , \9137 , \30535 );
and \U$25072 ( \30737 , \9139 , \30562 );
and \U$25073 ( \30738 , \9141 , \30589 );
and \U$25074 ( \30739 , \9143 , \30616 );
and \U$25075 ( \30740 , \9145 , \30643 );
or \U$25076 ( \30741 , \30725 , \30726 , \30727 , \30728 , \30729 , \30730 , \30731 , \30732 , \30733 , \30734 , \30735 , \30736 , \30737 , \30738 , \30739 , \30740 );
_DC g8f1f ( \30742_nG8f1f , \30741 , \30720 );
buf \U$25077 ( \30743 , \30742_nG8f1f );
xor \U$25078 ( \30744 , \30724 , \30743 );
or \U$25079 ( \30745 , \30723 , \30744 );
buf \U$25080 ( \30746 , RIb7af540_256);
and \U$25081 ( \30747 , \7217 , \30238 );
and \U$25082 ( \30748 , \7219 , \30265 );
and \U$25083 ( \30749 , \9155 , \30292 );
and \U$25084 ( \30750 , \9157 , \30319 );
and \U$25085 ( \30751 , \9159 , \30346 );
and \U$25086 ( \30752 , \9161 , \30373 );
and \U$25087 ( \30753 , \9163 , \30400 );
and \U$25088 ( \30754 , \9165 , \30427 );
and \U$25089 ( \30755 , \9167 , \30454 );
and \U$25090 ( \30756 , \9169 , \30481 );
and \U$25091 ( \30757 , \9171 , \30508 );
and \U$25092 ( \30758 , \9173 , \30535 );
and \U$25093 ( \30759 , \9175 , \30562 );
and \U$25094 ( \30760 , \9177 , \30589 );
and \U$25095 ( \30761 , \9179 , \30616 );
and \U$25096 ( \30762 , \9181 , \30643 );
or \U$25097 ( \30763 , \30747 , \30748 , \30749 , \30750 , \30751 , \30752 , \30753 , \30754 , \30755 , \30756 , \30757 , \30758 , \30759 , \30760 , \30761 , \30762 );
_DC g8f35 ( \30764_nG8f35 , \30763 , \30720 );
buf \U$25098 ( \30765 , \30764_nG8f35 );
xor \U$25099 ( \30766 , \30746 , \30765 );
or \U$25100 ( \30767 , \30745 , \30766 );
buf \U$25101 ( \30768 , RIb7af4c8_257);
and \U$25102 ( \30769 , \7227 , \30238 );
and \U$25103 ( \30770 , \7229 , \30265 );
and \U$25104 ( \30771 , \9191 , \30292 );
and \U$25105 ( \30772 , \9193 , \30319 );
and \U$25106 ( \30773 , \9195 , \30346 );
and \U$25107 ( \30774 , \9197 , \30373 );
and \U$25108 ( \30775 , \9199 , \30400 );
and \U$25109 ( \30776 , \9201 , \30427 );
and \U$25110 ( \30777 , \9203 , \30454 );
and \U$25111 ( \30778 , \9205 , \30481 );
and \U$25112 ( \30779 , \9207 , \30508 );
and \U$25113 ( \30780 , \9209 , \30535 );
and \U$25114 ( \30781 , \9211 , \30562 );
and \U$25115 ( \30782 , \9213 , \30589 );
and \U$25116 ( \30783 , \9215 , \30616 );
and \U$25117 ( \30784 , \9217 , \30643 );
or \U$25118 ( \30785 , \30769 , \30770 , \30771 , \30772 , \30773 , \30774 , \30775 , \30776 , \30777 , \30778 , \30779 , \30780 , \30781 , \30782 , \30783 , \30784 );
_DC g8f4b ( \30786_nG8f4b , \30785 , \30720 );
buf \U$25119 ( \30787 , \30786_nG8f4b );
xor \U$25120 ( \30788 , \30768 , \30787 );
or \U$25121 ( \30789 , \30767 , \30788 );
buf \U$25122 ( \30790 , RIb7af450_258);
and \U$25123 ( \30791 , \7237 , \30238 );
and \U$25124 ( \30792 , \7239 , \30265 );
and \U$25125 ( \30793 , \9227 , \30292 );
and \U$25126 ( \30794 , \9229 , \30319 );
and \U$25127 ( \30795 , \9231 , \30346 );
and \U$25128 ( \30796 , \9233 , \30373 );
and \U$25129 ( \30797 , \9235 , \30400 );
and \U$25130 ( \30798 , \9237 , \30427 );
and \U$25131 ( \30799 , \9239 , \30454 );
and \U$25132 ( \30800 , \9241 , \30481 );
and \U$25133 ( \30801 , \9243 , \30508 );
and \U$25134 ( \30802 , \9245 , \30535 );
and \U$25135 ( \30803 , \9247 , \30562 );
and \U$25136 ( \30804 , \9249 , \30589 );
and \U$25137 ( \30805 , \9251 , \30616 );
and \U$25138 ( \30806 , \9253 , \30643 );
or \U$25139 ( \30807 , \30791 , \30792 , \30793 , \30794 , \30795 , \30796 , \30797 , \30798 , \30799 , \30800 , \30801 , \30802 , \30803 , \30804 , \30805 , \30806 );
_DC g8f61 ( \30808_nG8f61 , \30807 , \30720 );
buf \U$25140 ( \30809 , \30808_nG8f61 );
xor \U$25141 ( \30810 , \30790 , \30809 );
or \U$25142 ( \30811 , \30789 , \30810 );
buf \U$25143 ( \30812 , RIb7af3d8_259);
and \U$25144 ( \30813 , \7247 , \30238 );
and \U$25145 ( \30814 , \7249 , \30265 );
and \U$25146 ( \30815 , \9263 , \30292 );
and \U$25147 ( \30816 , \9265 , \30319 );
and \U$25148 ( \30817 , \9267 , \30346 );
and \U$25149 ( \30818 , \9269 , \30373 );
and \U$25150 ( \30819 , \9271 , \30400 );
and \U$25151 ( \30820 , \9273 , \30427 );
and \U$25152 ( \30821 , \9275 , \30454 );
and \U$25153 ( \30822 , \9277 , \30481 );
and \U$25154 ( \30823 , \9279 , \30508 );
and \U$25155 ( \30824 , \9281 , \30535 );
and \U$25156 ( \30825 , \9283 , \30562 );
and \U$25157 ( \30826 , \9285 , \30589 );
and \U$25158 ( \30827 , \9287 , \30616 );
and \U$25159 ( \30828 , \9289 , \30643 );
or \U$25160 ( \30829 , \30813 , \30814 , \30815 , \30816 , \30817 , \30818 , \30819 , \30820 , \30821 , \30822 , \30823 , \30824 , \30825 , \30826 , \30827 , \30828 );
_DC g8f77 ( \30830_nG8f77 , \30829 , \30720 );
buf \U$25161 ( \30831 , \30830_nG8f77 );
xor \U$25162 ( \30832 , \30812 , \30831 );
or \U$25163 ( \30833 , \30811 , \30832 );
buf \U$25164 ( \30834 , RIb7a5bf8_260);
and \U$25165 ( \30835 , \7257 , \30238 );
and \U$25166 ( \30836 , \7259 , \30265 );
and \U$25167 ( \30837 , \9299 , \30292 );
and \U$25168 ( \30838 , \9301 , \30319 );
and \U$25169 ( \30839 , \9303 , \30346 );
and \U$25170 ( \30840 , \9305 , \30373 );
and \U$25171 ( \30841 , \9307 , \30400 );
and \U$25172 ( \30842 , \9309 , \30427 );
and \U$25173 ( \30843 , \9311 , \30454 );
and \U$25174 ( \30844 , \9313 , \30481 );
and \U$25175 ( \30845 , \9315 , \30508 );
and \U$25176 ( \30846 , \9317 , \30535 );
and \U$25177 ( \30847 , \9319 , \30562 );
and \U$25178 ( \30848 , \9321 , \30589 );
and \U$25179 ( \30849 , \9323 , \30616 );
and \U$25180 ( \30850 , \9325 , \30643 );
or \U$25181 ( \30851 , \30835 , \30836 , \30837 , \30838 , \30839 , \30840 , \30841 , \30842 , \30843 , \30844 , \30845 , \30846 , \30847 , \30848 , \30849 , \30850 );
_DC g8f8d ( \30852_nG8f8d , \30851 , \30720 );
buf \U$25182 ( \30853 , \30852_nG8f8d );
xor \U$25183 ( \30854 , \30834 , \30853 );
or \U$25184 ( \30855 , \30833 , \30854 );
buf \U$25185 ( \30856 , RIb7a0c48_261);
and \U$25186 ( \30857 , \7267 , \30238 );
and \U$25187 ( \30858 , \7269 , \30265 );
and \U$25188 ( \30859 , \9335 , \30292 );
and \U$25189 ( \30860 , \9337 , \30319 );
and \U$25190 ( \30861 , \9339 , \30346 );
and \U$25191 ( \30862 , \9341 , \30373 );
and \U$25192 ( \30863 , \9343 , \30400 );
and \U$25193 ( \30864 , \9345 , \30427 );
and \U$25194 ( \30865 , \9347 , \30454 );
and \U$25195 ( \30866 , \9349 , \30481 );
and \U$25196 ( \30867 , \9351 , \30508 );
and \U$25197 ( \30868 , \9353 , \30535 );
and \U$25198 ( \30869 , \9355 , \30562 );
and \U$25199 ( \30870 , \9357 , \30589 );
and \U$25200 ( \30871 , \9359 , \30616 );
and \U$25201 ( \30872 , \9361 , \30643 );
or \U$25202 ( \30873 , \30857 , \30858 , \30859 , \30860 , \30861 , \30862 , \30863 , \30864 , \30865 , \30866 , \30867 , \30868 , \30869 , \30870 , \30871 , \30872 );
_DC g8fa3 ( \30874_nG8fa3 , \30873 , \30720 );
buf \U$25203 ( \30875 , \30874_nG8fa3 );
xor \U$25204 ( \30876 , \30856 , \30875 );
or \U$25205 ( \30877 , \30855 , \30876 );
not \U$25206 ( \30878 , \30877 );
buf \U$25207 ( \30879 , \30878 );
and \U$25208 ( \30880 , \30211 , \30879 );
_HMUX g8faa ( \30881_nG8faa , \28658_nG86f3 , \29015 , \30880 );
buf \U$25209 ( \30882 , \28679 );
buf \U$25210 ( \30883 , \28676 );
buf \U$25211 ( \30884 , \28661 );
buf \U$25212 ( \30885 , \28664 );
buf \U$25213 ( \30886 , \28668 );
buf \U$25214 ( \30887 , \28672 );
or \U$25215 ( \30888 , \30884 , \30885 , \30886 , \30887 );
and \U$25216 ( \30889 , \30883 , \30888 );
or \U$25217 ( \30890 , \30882 , \30889 );
buf \U$25218 ( \30891 , \30890 );
_HMUX g8fb5 ( \30892_nG8fb5 , \29014_nG8857 , \30881_nG8faa , \30891 );
buf \U$25219 ( \30893 , RIe5319e0_6884);
buf \U$25221 ( \30894 , \30893 );
buf \U$25222 ( \30895 , RIe549ef0_6842);
buf \U$25224 ( \30896 , \30895 );
buf \U$25225 ( \30897 , RIe549770_6843);
not \U$25226 ( \30898 , \30897 );
buf \U$25227 ( \30899 , \30898 );
buf \U$25228 ( \30900 , RIe548ff0_6844);
xor \U$25229 ( \30901 , \30900 , \30897 );
buf \U$25230 ( \30902 , \30901 );
buf \U$25231 ( \30903 , RIea91330_6888);
and \U$25232 ( \30904 , \30900 , \30897 );
xor \U$25233 ( \30905 , \30903 , \30904 );
buf \U$25234 ( \30906 , \30905 );
not \U$25235 ( \30907 , \30906 );
and \U$25236 ( \30908 , \30903 , \30904 );
buf \U$25237 ( \30909 , \30908 );
nor \U$25238 ( \30910 , \30894 , \30896 , \30899 , \30902 , \30907 , \30909 );
and \U$25239 ( \30911 , RIe5329d0_6883, \30910 );
not \U$25240 ( \30912 , \30909 );
and \U$25241 ( \30913 , \30894 , \30896 , \30899 , \30902 , \30907 , \30912 );
and \U$25242 ( \30914 , RIeb72150_6905, \30913 );
not \U$25243 ( \30915 , \30894 );
and \U$25244 ( \30916 , \30915 , \30896 , \30899 , \30902 , \30907 , \30912 );
and \U$25245 ( \30917 , RIeab80c0_6897, \30916 );
not \U$25246 ( \30918 , \30896 );
and \U$25247 ( \30919 , \30894 , \30918 , \30899 , \30902 , \30907 , \30912 );
and \U$25248 ( \30920 , RIe5331c8_6882, \30919 );
and \U$25249 ( \30921 , \30915 , \30918 , \30899 , \30902 , \30907 , \30912 );
and \U$25250 ( \30922 , RIe5339c0_6881, \30921 );
not \U$25251 ( \30923 , \30899 );
and \U$25252 ( \30924 , \30894 , \30896 , \30923 , \30902 , \30907 , \30912 );
and \U$25253 ( \30925 , RIeab87c8_6898, \30924 );
and \U$25254 ( \30926 , \30915 , \30896 , \30923 , \30902 , \30907 , \30912 );
and \U$25255 ( \30927 , RIe5341b8_6880, \30926 );
and \U$25256 ( \30928 , \30894 , \30918 , \30923 , \30902 , \30907 , \30912 );
and \U$25257 ( \30929 , RIe5349b0_6879, \30928 );
and \U$25258 ( \30930 , \30915 , \30918 , \30923 , \30902 , \30907 , \30912 );
and \U$25259 ( \30931 , RIea94af8_6890, \30930 );
nor \U$25260 ( \30932 , \30915 , \30918 , \30923 , \30902 , \30906 , \30909 );
and \U$25261 ( \30933 , RIe5351a8_6878, \30932 );
nor \U$25262 ( \30934 , \30894 , \30918 , \30923 , \30902 , \30906 , \30909 );
and \U$25263 ( \30935 , RIe5359a0_6877, \30934 );
nor \U$25264 ( \30936 , \30915 , \30896 , \30923 , \30902 , \30906 , \30909 );
and \U$25265 ( \30937 , RIeab78c8_6895, \30936 );
nor \U$25266 ( \30938 , \30894 , \30896 , \30923 , \30902 , \30906 , \30909 );
and \U$25267 ( \30939 , RIeab7d00_6896, \30938 );
or \U$25271 ( \30940 , \30911 , \30914 , \30917 , \30920 , \30922 , \30925 , \30927 , \30929 , \30931 , \30933 , \30935 , \30937 , \30939 , 1'b0 , 1'b0 , 1'b0 );
buf \U$25273 ( \30941 , \30909 );
buf \U$25274 ( \30942 , \30906 );
buf \U$25275 ( \30943 , \30894 );
buf \U$25276 ( \30944 , \30896 );
buf \U$25277 ( \30945 , \30899 );
buf \U$25278 ( \30946 , \30902 );
or \U$25279 ( \30947 , \30943 , \30944 , \30945 , \30946 );
and \U$25280 ( \30948 , \30942 , \30947 );
or \U$25281 ( \30949 , \30941 , \30948 );
buf \U$25282 ( \30950 , \30949 );
or \U$25283 ( \30951 , 1'b0 , \30950 );
_DC g8ff3 ( \30952_nG8ff3 , \30940 , \30951 );
not \U$25284 ( \30953 , \30952_nG8ff3 );
buf \U$25285 ( \30954 , RIb7b9608_246);
and \U$25286 ( \30955 , \7117 , \30910 );
and \U$25287 ( \30956 , \7119 , \30913 );
and \U$25288 ( \30957 , \7864 , \30916 );
and \U$25289 ( \30958 , \7892 , \30919 );
and \U$25290 ( \30959 , \7920 , \30921 );
and \U$25291 ( \30960 , \7948 , \30924 );
and \U$25292 ( \30961 , \7976 , \30926 );
and \U$25293 ( \30962 , \8004 , \30928 );
and \U$25294 ( \30963 , \8032 , \30930 );
and \U$25295 ( \30964 , \8060 , \30932 );
and \U$25296 ( \30965 , \8088 , \30934 );
and \U$25297 ( \30966 , \8116 , \30936 );
and \U$25298 ( \30967 , \8144 , \30938 );
or \U$25302 ( \30968 , \30955 , \30956 , \30957 , \30958 , \30959 , \30960 , \30961 , \30962 , \30963 , \30964 , \30965 , \30966 , \30967 , 1'b0 , 1'b0 , 1'b0 );
_DC g9004 ( \30969_nG9004 , \30968 , \30951 );
buf \U$25303 ( \30970 , \30969_nG9004 );
xor \U$25304 ( \30971 , \30954 , \30970 );
buf \U$25305 ( \30972 , RIb7b9590_247);
and \U$25306 ( \30973 , \7126 , \30910 );
and \U$25307 ( \30974 , \7128 , \30913 );
and \U$25308 ( \30975 , \8338 , \30916 );
and \U$25309 ( \30976 , \8340 , \30919 );
and \U$25310 ( \30977 , \8342 , \30921 );
and \U$25311 ( \30978 , \8344 , \30924 );
and \U$25312 ( \30979 , \8346 , \30926 );
and \U$25313 ( \30980 , \8348 , \30928 );
and \U$25314 ( \30981 , \8350 , \30930 );
and \U$25315 ( \30982 , \8352 , \30932 );
and \U$25316 ( \30983 , \8354 , \30934 );
and \U$25317 ( \30984 , \8356 , \30936 );
and \U$25318 ( \30985 , \8358 , \30938 );
or \U$25322 ( \30986 , \30973 , \30974 , \30975 , \30976 , \30977 , \30978 , \30979 , \30980 , \30981 , \30982 , \30983 , \30984 , \30985 , 1'b0 , 1'b0 , 1'b0 );
_DC g9016 ( \30987_nG9016 , \30986 , \30951 );
buf \U$25323 ( \30988 , \30987_nG9016 );
xor \U$25324 ( \30989 , \30972 , \30988 );
or \U$25325 ( \30990 , \30971 , \30989 );
buf \U$25326 ( \30991 , RIb7b9518_248);
and \U$25327 ( \30992 , \7136 , \30910 );
and \U$25328 ( \30993 , \7138 , \30913 );
and \U$25329 ( \30994 , \8374 , \30916 );
and \U$25330 ( \30995 , \8376 , \30919 );
and \U$25331 ( \30996 , \8378 , \30921 );
and \U$25332 ( \30997 , \8380 , \30924 );
and \U$25333 ( \30998 , \8382 , \30926 );
and \U$25334 ( \30999 , \8384 , \30928 );
and \U$25335 ( \31000 , \8386 , \30930 );
and \U$25336 ( \31001 , \8388 , \30932 );
and \U$25337 ( \31002 , \8390 , \30934 );
and \U$25338 ( \31003 , \8392 , \30936 );
and \U$25339 ( \31004 , \8394 , \30938 );
or \U$25343 ( \31005 , \30992 , \30993 , \30994 , \30995 , \30996 , \30997 , \30998 , \30999 , \31000 , \31001 , \31002 , \31003 , \31004 , 1'b0 , 1'b0 , 1'b0 );
_DC g9029 ( \31006_nG9029 , \31005 , \30951 );
buf \U$25344 ( \31007 , \31006_nG9029 );
xor \U$25345 ( \31008 , \30991 , \31007 );
or \U$25346 ( \31009 , \30990 , \31008 );
buf \U$25347 ( \31010 , RIb7b94a0_249);
and \U$25348 ( \31011 , \7146 , \30910 );
and \U$25349 ( \31012 , \7148 , \30913 );
and \U$25350 ( \31013 , \8410 , \30916 );
and \U$25351 ( \31014 , \8412 , \30919 );
and \U$25352 ( \31015 , \8414 , \30921 );
and \U$25353 ( \31016 , \8416 , \30924 );
and \U$25354 ( \31017 , \8418 , \30926 );
and \U$25355 ( \31018 , \8420 , \30928 );
and \U$25356 ( \31019 , \8422 , \30930 );
and \U$25357 ( \31020 , \8424 , \30932 );
and \U$25358 ( \31021 , \8426 , \30934 );
and \U$25359 ( \31022 , \8428 , \30936 );
and \U$25360 ( \31023 , \8430 , \30938 );
or \U$25364 ( \31024 , \31011 , \31012 , \31013 , \31014 , \31015 , \31016 , \31017 , \31018 , \31019 , \31020 , \31021 , \31022 , \31023 , 1'b0 , 1'b0 , 1'b0 );
_DC g903c ( \31025_nG903c , \31024 , \30951 );
buf \U$25365 ( \31026 , \31025_nG903c );
xor \U$25366 ( \31027 , \31010 , \31026 );
or \U$25367 ( \31028 , \31009 , \31027 );
buf \U$25368 ( \31029 , RIb7b9428_250);
and \U$25369 ( \31030 , \7156 , \30910 );
and \U$25370 ( \31031 , \7158 , \30913 );
and \U$25371 ( \31032 , \8446 , \30916 );
and \U$25372 ( \31033 , \8448 , \30919 );
and \U$25373 ( \31034 , \8450 , \30921 );
and \U$25374 ( \31035 , \8452 , \30924 );
and \U$25375 ( \31036 , \8454 , \30926 );
and \U$25376 ( \31037 , \8456 , \30928 );
and \U$25377 ( \31038 , \8458 , \30930 );
and \U$25378 ( \31039 , \8460 , \30932 );
and \U$25379 ( \31040 , \8462 , \30934 );
and \U$25380 ( \31041 , \8464 , \30936 );
and \U$25381 ( \31042 , \8466 , \30938 );
or \U$25385 ( \31043 , \31030 , \31031 , \31032 , \31033 , \31034 , \31035 , \31036 , \31037 , \31038 , \31039 , \31040 , \31041 , \31042 , 1'b0 , 1'b0 , 1'b0 );
_DC g904f ( \31044_nG904f , \31043 , \30951 );
buf \U$25386 ( \31045 , \31044_nG904f );
xor \U$25387 ( \31046 , \31029 , \31045 );
or \U$25388 ( \31047 , \31028 , \31046 );
buf \U$25389 ( \31048 , RIb7b93b0_251);
and \U$25390 ( \31049 , \7166 , \30910 );
and \U$25391 ( \31050 , \7168 , \30913 );
and \U$25392 ( \31051 , \8482 , \30916 );
and \U$25393 ( \31052 , \8484 , \30919 );
and \U$25394 ( \31053 , \8486 , \30921 );
and \U$25395 ( \31054 , \8488 , \30924 );
and \U$25396 ( \31055 , \8490 , \30926 );
and \U$25397 ( \31056 , \8492 , \30928 );
and \U$25398 ( \31057 , \8494 , \30930 );
and \U$25399 ( \31058 , \8496 , \30932 );
and \U$25400 ( \31059 , \8498 , \30934 );
and \U$25401 ( \31060 , \8500 , \30936 );
and \U$25402 ( \31061 , \8502 , \30938 );
or \U$25406 ( \31062 , \31049 , \31050 , \31051 , \31052 , \31053 , \31054 , \31055 , \31056 , \31057 , \31058 , \31059 , \31060 , \31061 , 1'b0 , 1'b0 , 1'b0 );
_DC g9062 ( \31063_nG9062 , \31062 , \30951 );
buf \U$25407 ( \31064 , \31063_nG9062 );
xor \U$25408 ( \31065 , \31048 , \31064 );
or \U$25409 ( \31066 , \31047 , \31065 );
buf \U$25410 ( \31067 , RIb7af720_252);
and \U$25411 ( \31068 , \7176 , \30910 );
and \U$25412 ( \31069 , \7178 , \30913 );
and \U$25413 ( \31070 , \8518 , \30916 );
and \U$25414 ( \31071 , \8520 , \30919 );
and \U$25415 ( \31072 , \8522 , \30921 );
and \U$25416 ( \31073 , \8524 , \30924 );
and \U$25417 ( \31074 , \8526 , \30926 );
and \U$25418 ( \31075 , \8528 , \30928 );
and \U$25419 ( \31076 , \8530 , \30930 );
and \U$25420 ( \31077 , \8532 , \30932 );
and \U$25421 ( \31078 , \8534 , \30934 );
and \U$25422 ( \31079 , \8536 , \30936 );
and \U$25423 ( \31080 , \8538 , \30938 );
or \U$25427 ( \31081 , \31068 , \31069 , \31070 , \31071 , \31072 , \31073 , \31074 , \31075 , \31076 , \31077 , \31078 , \31079 , \31080 , 1'b0 , 1'b0 , 1'b0 );
_DC g9075 ( \31082_nG9075 , \31081 , \30951 );
buf \U$25428 ( \31083 , \31082_nG9075 );
xor \U$25429 ( \31084 , \31067 , \31083 );
or \U$25430 ( \31085 , \31066 , \31084 );
buf \U$25431 ( \31086 , RIb7af6a8_253);
and \U$25432 ( \31087 , \7186 , \30910 );
and \U$25433 ( \31088 , \7188 , \30913 );
and \U$25434 ( \31089 , \8554 , \30916 );
and \U$25435 ( \31090 , \8556 , \30919 );
and \U$25436 ( \31091 , \8558 , \30921 );
and \U$25437 ( \31092 , \8560 , \30924 );
and \U$25438 ( \31093 , \8562 , \30926 );
and \U$25439 ( \31094 , \8564 , \30928 );
and \U$25440 ( \31095 , \8566 , \30930 );
and \U$25441 ( \31096 , \8568 , \30932 );
and \U$25442 ( \31097 , \8570 , \30934 );
and \U$25443 ( \31098 , \8572 , \30936 );
and \U$25444 ( \31099 , \8574 , \30938 );
or \U$25448 ( \31100 , \31087 , \31088 , \31089 , \31090 , \31091 , \31092 , \31093 , \31094 , \31095 , \31096 , \31097 , \31098 , \31099 , 1'b0 , 1'b0 , 1'b0 );
_DC g9088 ( \31101_nG9088 , \31100 , \30951 );
buf \U$25449 ( \31102 , \31101_nG9088 );
xor \U$25450 ( \31103 , \31086 , \31102 );
or \U$25451 ( \31104 , \31085 , \31103 );
not \U$25452 ( \31105 , \31104 );
buf \U$25453 ( \31106 , \31105 );
buf \U$25454 ( \31107 , RIb7af630_254);
and \U$25455 ( \31108 , \7198 , \30910 );
and \U$25456 ( \31109 , \7200 , \30913 );
and \U$25457 ( \31110 , \8645 , \30916 );
and \U$25458 ( \31111 , \8673 , \30919 );
and \U$25459 ( \31112 , \8701 , \30921 );
and \U$25460 ( \31113 , \8729 , \30924 );
and \U$25461 ( \31114 , \8757 , \30926 );
and \U$25462 ( \31115 , \8785 , \30928 );
and \U$25463 ( \31116 , \8813 , \30930 );
and \U$25464 ( \31117 , \8841 , \30932 );
and \U$25465 ( \31118 , \8869 , \30934 );
and \U$25466 ( \31119 , \8897 , \30936 );
and \U$25467 ( \31120 , \8925 , \30938 );
or \U$25471 ( \31121 , \31108 , \31109 , \31110 , \31111 , \31112 , \31113 , \31114 , \31115 , \31116 , \31117 , \31118 , \31119 , \31120 , 1'b0 , 1'b0 , 1'b0 );
_DC g909d ( \31122_nG909d , \31121 , \30951 );
buf \U$25472 ( \31123 , \31122_nG909d );
xor \U$25473 ( \31124 , \31107 , \31123 );
buf \U$25474 ( \31125 , RIb7af5b8_255);
and \U$25475 ( \31126 , \7207 , \30910 );
and \U$25476 ( \31127 , \7209 , \30913 );
and \U$25477 ( \31128 , \9119 , \30916 );
and \U$25478 ( \31129 , \9121 , \30919 );
and \U$25479 ( \31130 , \9123 , \30921 );
and \U$25480 ( \31131 , \9125 , \30924 );
and \U$25481 ( \31132 , \9127 , \30926 );
and \U$25482 ( \31133 , \9129 , \30928 );
and \U$25483 ( \31134 , \9131 , \30930 );
and \U$25484 ( \31135 , \9133 , \30932 );
and \U$25485 ( \31136 , \9135 , \30934 );
and \U$25486 ( \31137 , \9137 , \30936 );
and \U$25487 ( \31138 , \9139 , \30938 );
or \U$25491 ( \31139 , \31126 , \31127 , \31128 , \31129 , \31130 , \31131 , \31132 , \31133 , \31134 , \31135 , \31136 , \31137 , \31138 , 1'b0 , 1'b0 , 1'b0 );
_DC g90af ( \31140_nG90af , \31139 , \30951 );
buf \U$25492 ( \31141 , \31140_nG90af );
xor \U$25493 ( \31142 , \31125 , \31141 );
or \U$25494 ( \31143 , \31124 , \31142 );
buf \U$25495 ( \31144 , RIb7af540_256);
and \U$25496 ( \31145 , \7217 , \30910 );
and \U$25497 ( \31146 , \7219 , \30913 );
and \U$25498 ( \31147 , \9155 , \30916 );
and \U$25499 ( \31148 , \9157 , \30919 );
and \U$25500 ( \31149 , \9159 , \30921 );
and \U$25501 ( \31150 , \9161 , \30924 );
and \U$25502 ( \31151 , \9163 , \30926 );
and \U$25503 ( \31152 , \9165 , \30928 );
and \U$25504 ( \31153 , \9167 , \30930 );
and \U$25505 ( \31154 , \9169 , \30932 );
and \U$25506 ( \31155 , \9171 , \30934 );
and \U$25507 ( \31156 , \9173 , \30936 );
and \U$25508 ( \31157 , \9175 , \30938 );
or \U$25512 ( \31158 , \31145 , \31146 , \31147 , \31148 , \31149 , \31150 , \31151 , \31152 , \31153 , \31154 , \31155 , \31156 , \31157 , 1'b0 , 1'b0 , 1'b0 );
_DC g90c2 ( \31159_nG90c2 , \31158 , \30951 );
buf \U$25513 ( \31160 , \31159_nG90c2 );
xor \U$25514 ( \31161 , \31144 , \31160 );
or \U$25515 ( \31162 , \31143 , \31161 );
buf \U$25516 ( \31163 , RIb7af4c8_257);
and \U$25517 ( \31164 , \7227 , \30910 );
and \U$25518 ( \31165 , \7229 , \30913 );
and \U$25519 ( \31166 , \9191 , \30916 );
and \U$25520 ( \31167 , \9193 , \30919 );
and \U$25521 ( \31168 , \9195 , \30921 );
and \U$25522 ( \31169 , \9197 , \30924 );
and \U$25523 ( \31170 , \9199 , \30926 );
and \U$25524 ( \31171 , \9201 , \30928 );
and \U$25525 ( \31172 , \9203 , \30930 );
and \U$25526 ( \31173 , \9205 , \30932 );
and \U$25527 ( \31174 , \9207 , \30934 );
and \U$25528 ( \31175 , \9209 , \30936 );
and \U$25529 ( \31176 , \9211 , \30938 );
or \U$25533 ( \31177 , \31164 , \31165 , \31166 , \31167 , \31168 , \31169 , \31170 , \31171 , \31172 , \31173 , \31174 , \31175 , \31176 , 1'b0 , 1'b0 , 1'b0 );
_DC g90d5 ( \31178_nG90d5 , \31177 , \30951 );
buf \U$25534 ( \31179 , \31178_nG90d5 );
xor \U$25535 ( \31180 , \31163 , \31179 );
or \U$25536 ( \31181 , \31162 , \31180 );
buf \U$25537 ( \31182 , RIb7af450_258);
and \U$25538 ( \31183 , \7237 , \30910 );
and \U$25539 ( \31184 , \7239 , \30913 );
and \U$25540 ( \31185 , \9227 , \30916 );
and \U$25541 ( \31186 , \9229 , \30919 );
and \U$25542 ( \31187 , \9231 , \30921 );
and \U$25543 ( \31188 , \9233 , \30924 );
and \U$25544 ( \31189 , \9235 , \30926 );
and \U$25545 ( \31190 , \9237 , \30928 );
and \U$25546 ( \31191 , \9239 , \30930 );
and \U$25547 ( \31192 , \9241 , \30932 );
and \U$25548 ( \31193 , \9243 , \30934 );
and \U$25549 ( \31194 , \9245 , \30936 );
and \U$25550 ( \31195 , \9247 , \30938 );
or \U$25554 ( \31196 , \31183 , \31184 , \31185 , \31186 , \31187 , \31188 , \31189 , \31190 , \31191 , \31192 , \31193 , \31194 , \31195 , 1'b0 , 1'b0 , 1'b0 );
_DC g90e8 ( \31197_nG90e8 , \31196 , \30951 );
buf \U$25555 ( \31198 , \31197_nG90e8 );
xor \U$25556 ( \31199 , \31182 , \31198 );
or \U$25557 ( \31200 , \31181 , \31199 );
buf \U$25558 ( \31201 , RIb7af3d8_259);
and \U$25559 ( \31202 , \7247 , \30910 );
and \U$25560 ( \31203 , \7249 , \30913 );
and \U$25561 ( \31204 , \9263 , \30916 );
and \U$25562 ( \31205 , \9265 , \30919 );
and \U$25563 ( \31206 , \9267 , \30921 );
and \U$25564 ( \31207 , \9269 , \30924 );
and \U$25565 ( \31208 , \9271 , \30926 );
and \U$25566 ( \31209 , \9273 , \30928 );
and \U$25567 ( \31210 , \9275 , \30930 );
and \U$25568 ( \31211 , \9277 , \30932 );
and \U$25569 ( \31212 , \9279 , \30934 );
and \U$25570 ( \31213 , \9281 , \30936 );
and \U$25571 ( \31214 , \9283 , \30938 );
or \U$25575 ( \31215 , \31202 , \31203 , \31204 , \31205 , \31206 , \31207 , \31208 , \31209 , \31210 , \31211 , \31212 , \31213 , \31214 , 1'b0 , 1'b0 , 1'b0 );
_DC g90fb ( \31216_nG90fb , \31215 , \30951 );
buf \U$25576 ( \31217 , \31216_nG90fb );
xor \U$25577 ( \31218 , \31201 , \31217 );
or \U$25578 ( \31219 , \31200 , \31218 );
buf \U$25579 ( \31220 , RIb7a5bf8_260);
and \U$25580 ( \31221 , \7257 , \30910 );
and \U$25581 ( \31222 , \7259 , \30913 );
and \U$25582 ( \31223 , \9299 , \30916 );
and \U$25583 ( \31224 , \9301 , \30919 );
and \U$25584 ( \31225 , \9303 , \30921 );
and \U$25585 ( \31226 , \9305 , \30924 );
and \U$25586 ( \31227 , \9307 , \30926 );
and \U$25587 ( \31228 , \9309 , \30928 );
and \U$25588 ( \31229 , \9311 , \30930 );
and \U$25589 ( \31230 , \9313 , \30932 );
and \U$25590 ( \31231 , \9315 , \30934 );
and \U$25591 ( \31232 , \9317 , \30936 );
and \U$25592 ( \31233 , \9319 , \30938 );
or \U$25596 ( \31234 , \31221 , \31222 , \31223 , \31224 , \31225 , \31226 , \31227 , \31228 , \31229 , \31230 , \31231 , \31232 , \31233 , 1'b0 , 1'b0 , 1'b0 );
_DC g910e ( \31235_nG910e , \31234 , \30951 );
buf \U$25597 ( \31236 , \31235_nG910e );
xor \U$25598 ( \31237 , \31220 , \31236 );
or \U$25599 ( \31238 , \31219 , \31237 );
buf \U$25600 ( \31239 , RIb7a0c48_261);
and \U$25601 ( \31240 , \7267 , \30910 );
and \U$25602 ( \31241 , \7269 , \30913 );
and \U$25603 ( \31242 , \9335 , \30916 );
and \U$25604 ( \31243 , \9337 , \30919 );
and \U$25605 ( \31244 , \9339 , \30921 );
and \U$25606 ( \31245 , \9341 , \30924 );
and \U$25607 ( \31246 , \9343 , \30926 );
and \U$25608 ( \31247 , \9345 , \30928 );
and \U$25609 ( \31248 , \9347 , \30930 );
and \U$25610 ( \31249 , \9349 , \30932 );
and \U$25611 ( \31250 , \9351 , \30934 );
and \U$25612 ( \31251 , \9353 , \30936 );
and \U$25613 ( \31252 , \9355 , \30938 );
or \U$25617 ( \31253 , \31240 , \31241 , \31242 , \31243 , \31244 , \31245 , \31246 , \31247 , \31248 , \31249 , \31250 , \31251 , \31252 , 1'b0 , 1'b0 , 1'b0 );
_DC g9121 ( \31254_nG9121 , \31253 , \30951 );
buf \U$25618 ( \31255 , \31254_nG9121 );
xor \U$25619 ( \31256 , \31239 , \31255 );
or \U$25620 ( \31257 , \31238 , \31256 );
not \U$25621 ( \31258 , \31257 );
buf \U$25622 ( \31259 , \31258 );
and \U$25623 ( \31260 , \31106 , \31259 );
and \U$25624 ( \31261 , \30953 , \31260 );
_HMUX g9129 ( \31262_nG9129 , \30892_nG8fb5 , \30894 , \31261 );
buf \U$25627 ( \31263 , \30894 );
buf \U$25630 ( \31264 , \30896 );
buf \U$25633 ( \31265 , \30899 );
buf \U$25636 ( \31266 , \30902 );
buf \U$25637 ( \31267 , \30906 );
not \U$25638 ( \31268 , \31267 );
buf \U$25639 ( \31269 , \31268 );
not \U$25640 ( \31270 , \31269 );
buf \U$25641 ( \31271 , \30909 );
xnor \U$25642 ( \31272 , \31271 , \31267 );
buf \U$25643 ( \31273 , \31272 );
or \U$25644 ( \31274 , \31271 , \31267 );
not \U$25645 ( \31275 , \31274 );
buf \U$25646 ( \31276 , \31275 );
buf \U$25647 ( \31277 , \31276 );
buf \U$25648 ( \31278 , \31276 );
buf \U$25649 ( \31279 , \31276 );
buf \U$25650 ( \31280 , \31276 );
buf \U$25651 ( \31281 , \31276 );
buf \U$25652 ( \31282 , \31276 );
buf \U$25653 ( \31283 , \31276 );
buf \U$25654 ( \31284 , \31276 );
buf \U$25655 ( \31285 , \31276 );
buf \U$25656 ( \31286 , \31276 );
buf \U$25657 ( \31287 , \31276 );
buf \U$25658 ( \31288 , \31276 );
buf \U$25659 ( \31289 , \31276 );
buf \U$25660 ( \31290 , \31276 );
buf \U$25661 ( \31291 , \31276 );
buf \U$25662 ( \31292 , \31276 );
buf \U$25663 ( \31293 , \31276 );
buf \U$25664 ( \31294 , \31276 );
buf \U$25665 ( \31295 , \31276 );
buf \U$25666 ( \31296 , \31276 );
buf \U$25667 ( \31297 , \31276 );
buf \U$25668 ( \31298 , \31276 );
buf \U$25669 ( \31299 , \31276 );
buf \U$25670 ( \31300 , \31276 );
buf \U$25671 ( \31301 , \31276 );
nor \U$25672 ( \31302 , \31263 , \31264 , \31265 , \31266 , \31270 , \31273 , \31276 , \31277 , \31278 , \31279 , \31280 , \31281 , \31282 , \31283 , \31284 , \31285 , \31286 , \31287 , \31288 , \31289 , \31290 , \31291 , \31292 , \31293 , \31294 , \31295 , \31296 , \31297 , \31298 , \31299 , \31300 , \31301 );
and \U$25673 ( \31303 , RIe5329d0_6883, \31302 );
not \U$25674 ( \31304 , \31263 );
not \U$25675 ( \31305 , \31264 );
not \U$25676 ( \31306 , \31265 );
not \U$25677 ( \31307 , \31266 );
buf \U$25678 ( \31308 , \31276 );
buf \U$25679 ( \31309 , \31276 );
buf \U$25680 ( \31310 , \31276 );
buf \U$25681 ( \31311 , \31276 );
buf \U$25682 ( \31312 , \31276 );
buf \U$25683 ( \31313 , \31276 );
buf \U$25684 ( \31314 , \31276 );
buf \U$25685 ( \31315 , \31276 );
buf \U$25686 ( \31316 , \31276 );
buf \U$25687 ( \31317 , \31276 );
buf \U$25688 ( \31318 , \31276 );
buf \U$25689 ( \31319 , \31276 );
buf \U$25690 ( \31320 , \31276 );
buf \U$25691 ( \31321 , \31276 );
buf \U$25692 ( \31322 , \31276 );
buf \U$25693 ( \31323 , \31276 );
buf \U$25694 ( \31324 , \31276 );
buf \U$25695 ( \31325 , \31276 );
buf \U$25696 ( \31326 , \31276 );
buf \U$25697 ( \31327 , \31276 );
buf \U$25698 ( \31328 , \31276 );
buf \U$25699 ( \31329 , \31276 );
buf \U$25700 ( \31330 , \31276 );
buf \U$25701 ( \31331 , \31276 );
buf \U$25702 ( \31332 , \31276 );
nor \U$25703 ( \31333 , \31304 , \31305 , \31306 , \31307 , \31269 , \31273 , \31276 , \31308 , \31309 , \31310 , \31311 , \31312 , \31313 , \31314 , \31315 , \31316 , \31317 , \31318 , \31319 , \31320 , \31321 , \31322 , \31323 , \31324 , \31325 , \31326 , \31327 , \31328 , \31329 , \31330 , \31331 , \31332 );
and \U$25704 ( \31334 , RIeb72150_6905, \31333 );
buf \U$25705 ( \31335 , \31276 );
buf \U$25706 ( \31336 , \31276 );
buf \U$25707 ( \31337 , \31276 );
buf \U$25708 ( \31338 , \31276 );
buf \U$25709 ( \31339 , \31276 );
buf \U$25710 ( \31340 , \31276 );
buf \U$25711 ( \31341 , \31276 );
buf \U$25712 ( \31342 , \31276 );
buf \U$25713 ( \31343 , \31276 );
buf \U$25714 ( \31344 , \31276 );
buf \U$25715 ( \31345 , \31276 );
buf \U$25716 ( \31346 , \31276 );
buf \U$25717 ( \31347 , \31276 );
buf \U$25718 ( \31348 , \31276 );
buf \U$25719 ( \31349 , \31276 );
buf \U$25720 ( \31350 , \31276 );
buf \U$25721 ( \31351 , \31276 );
buf \U$25722 ( \31352 , \31276 );
buf \U$25723 ( \31353 , \31276 );
buf \U$25724 ( \31354 , \31276 );
buf \U$25725 ( \31355 , \31276 );
buf \U$25726 ( \31356 , \31276 );
buf \U$25727 ( \31357 , \31276 );
buf \U$25728 ( \31358 , \31276 );
buf \U$25729 ( \31359 , \31276 );
nor \U$25730 ( \31360 , \31263 , \31305 , \31306 , \31307 , \31269 , \31273 , \31276 , \31335 , \31336 , \31337 , \31338 , \31339 , \31340 , \31341 , \31342 , \31343 , \31344 , \31345 , \31346 , \31347 , \31348 , \31349 , \31350 , \31351 , \31352 , \31353 , \31354 , \31355 , \31356 , \31357 , \31358 , \31359 );
and \U$25731 ( \31361 , RIeab80c0_6897, \31360 );
buf \U$25732 ( \31362 , \31276 );
buf \U$25733 ( \31363 , \31276 );
buf \U$25734 ( \31364 , \31276 );
buf \U$25735 ( \31365 , \31276 );
buf \U$25736 ( \31366 , \31276 );
buf \U$25737 ( \31367 , \31276 );
buf \U$25738 ( \31368 , \31276 );
buf \U$25739 ( \31369 , \31276 );
buf \U$25740 ( \31370 , \31276 );
buf \U$25741 ( \31371 , \31276 );
buf \U$25742 ( \31372 , \31276 );
buf \U$25743 ( \31373 , \31276 );
buf \U$25744 ( \31374 , \31276 );
buf \U$25745 ( \31375 , \31276 );
buf \U$25746 ( \31376 , \31276 );
buf \U$25747 ( \31377 , \31276 );
buf \U$25748 ( \31378 , \31276 );
buf \U$25749 ( \31379 , \31276 );
buf \U$25750 ( \31380 , \31276 );
buf \U$25751 ( \31381 , \31276 );
buf \U$25752 ( \31382 , \31276 );
buf \U$25753 ( \31383 , \31276 );
buf \U$25754 ( \31384 , \31276 );
buf \U$25755 ( \31385 , \31276 );
buf \U$25756 ( \31386 , \31276 );
nor \U$25757 ( \31387 , \31304 , \31264 , \31306 , \31307 , \31269 , \31273 , \31276 , \31362 , \31363 , \31364 , \31365 , \31366 , \31367 , \31368 , \31369 , \31370 , \31371 , \31372 , \31373 , \31374 , \31375 , \31376 , \31377 , \31378 , \31379 , \31380 , \31381 , \31382 , \31383 , \31384 , \31385 , \31386 );
and \U$25758 ( \31388 , RIe5331c8_6882, \31387 );
buf \U$25759 ( \31389 , \31276 );
buf \U$25760 ( \31390 , \31276 );
buf \U$25761 ( \31391 , \31276 );
buf \U$25762 ( \31392 , \31276 );
buf \U$25763 ( \31393 , \31276 );
buf \U$25764 ( \31394 , \31276 );
buf \U$25765 ( \31395 , \31276 );
buf \U$25766 ( \31396 , \31276 );
buf \U$25767 ( \31397 , \31276 );
buf \U$25768 ( \31398 , \31276 );
buf \U$25769 ( \31399 , \31276 );
buf \U$25770 ( \31400 , \31276 );
buf \U$25771 ( \31401 , \31276 );
buf \U$25772 ( \31402 , \31276 );
buf \U$25773 ( \31403 , \31276 );
buf \U$25774 ( \31404 , \31276 );
buf \U$25775 ( \31405 , \31276 );
buf \U$25776 ( \31406 , \31276 );
buf \U$25777 ( \31407 , \31276 );
buf \U$25778 ( \31408 , \31276 );
buf \U$25779 ( \31409 , \31276 );
buf \U$25780 ( \31410 , \31276 );
buf \U$25781 ( \31411 , \31276 );
buf \U$25782 ( \31412 , \31276 );
buf \U$25783 ( \31413 , \31276 );
nor \U$25784 ( \31414 , \31263 , \31264 , \31306 , \31307 , \31269 , \31273 , \31276 , \31389 , \31390 , \31391 , \31392 , \31393 , \31394 , \31395 , \31396 , \31397 , \31398 , \31399 , \31400 , \31401 , \31402 , \31403 , \31404 , \31405 , \31406 , \31407 , \31408 , \31409 , \31410 , \31411 , \31412 , \31413 );
and \U$25785 ( \31415 , RIe5339c0_6881, \31414 );
buf \U$25786 ( \31416 , \31276 );
buf \U$25787 ( \31417 , \31276 );
buf \U$25788 ( \31418 , \31276 );
buf \U$25789 ( \31419 , \31276 );
buf \U$25790 ( \31420 , \31276 );
buf \U$25791 ( \31421 , \31276 );
buf \U$25792 ( \31422 , \31276 );
buf \U$25793 ( \31423 , \31276 );
buf \U$25794 ( \31424 , \31276 );
buf \U$25795 ( \31425 , \31276 );
buf \U$25796 ( \31426 , \31276 );
buf \U$25797 ( \31427 , \31276 );
buf \U$25798 ( \31428 , \31276 );
buf \U$25799 ( \31429 , \31276 );
buf \U$25800 ( \31430 , \31276 );
buf \U$25801 ( \31431 , \31276 );
buf \U$25802 ( \31432 , \31276 );
buf \U$25803 ( \31433 , \31276 );
buf \U$25804 ( \31434 , \31276 );
buf \U$25805 ( \31435 , \31276 );
buf \U$25806 ( \31436 , \31276 );
buf \U$25807 ( \31437 , \31276 );
buf \U$25808 ( \31438 , \31276 );
buf \U$25809 ( \31439 , \31276 );
buf \U$25810 ( \31440 , \31276 );
nor \U$25811 ( \31441 , \31304 , \31305 , \31265 , \31307 , \31269 , \31273 , \31276 , \31416 , \31417 , \31418 , \31419 , \31420 , \31421 , \31422 , \31423 , \31424 , \31425 , \31426 , \31427 , \31428 , \31429 , \31430 , \31431 , \31432 , \31433 , \31434 , \31435 , \31436 , \31437 , \31438 , \31439 , \31440 );
and \U$25812 ( \31442 , RIeab87c8_6898, \31441 );
buf \U$25813 ( \31443 , \31276 );
buf \U$25814 ( \31444 , \31276 );
buf \U$25815 ( \31445 , \31276 );
buf \U$25816 ( \31446 , \31276 );
buf \U$25817 ( \31447 , \31276 );
buf \U$25818 ( \31448 , \31276 );
buf \U$25819 ( \31449 , \31276 );
buf \U$25820 ( \31450 , \31276 );
buf \U$25821 ( \31451 , \31276 );
buf \U$25822 ( \31452 , \31276 );
buf \U$25823 ( \31453 , \31276 );
buf \U$25824 ( \31454 , \31276 );
buf \U$25825 ( \31455 , \31276 );
buf \U$25826 ( \31456 , \31276 );
buf \U$25827 ( \31457 , \31276 );
buf \U$25828 ( \31458 , \31276 );
buf \U$25829 ( \31459 , \31276 );
buf \U$25830 ( \31460 , \31276 );
buf \U$25831 ( \31461 , \31276 );
buf \U$25832 ( \31462 , \31276 );
buf \U$25833 ( \31463 , \31276 );
buf \U$25834 ( \31464 , \31276 );
buf \U$25835 ( \31465 , \31276 );
buf \U$25836 ( \31466 , \31276 );
buf \U$25837 ( \31467 , \31276 );
nor \U$25838 ( \31468 , \31263 , \31305 , \31265 , \31307 , \31269 , \31273 , \31276 , \31443 , \31444 , \31445 , \31446 , \31447 , \31448 , \31449 , \31450 , \31451 , \31452 , \31453 , \31454 , \31455 , \31456 , \31457 , \31458 , \31459 , \31460 , \31461 , \31462 , \31463 , \31464 , \31465 , \31466 , \31467 );
and \U$25839 ( \31469 , RIe5341b8_6880, \31468 );
buf \U$25840 ( \31470 , \31276 );
buf \U$25841 ( \31471 , \31276 );
buf \U$25842 ( \31472 , \31276 );
buf \U$25843 ( \31473 , \31276 );
buf \U$25844 ( \31474 , \31276 );
buf \U$25845 ( \31475 , \31276 );
buf \U$25846 ( \31476 , \31276 );
buf \U$25847 ( \31477 , \31276 );
buf \U$25848 ( \31478 , \31276 );
buf \U$25849 ( \31479 , \31276 );
buf \U$25850 ( \31480 , \31276 );
buf \U$25851 ( \31481 , \31276 );
buf \U$25852 ( \31482 , \31276 );
buf \U$25853 ( \31483 , \31276 );
buf \U$25854 ( \31484 , \31276 );
buf \U$25855 ( \31485 , \31276 );
buf \U$25856 ( \31486 , \31276 );
buf \U$25857 ( \31487 , \31276 );
buf \U$25858 ( \31488 , \31276 );
buf \U$25859 ( \31489 , \31276 );
buf \U$25860 ( \31490 , \31276 );
buf \U$25861 ( \31491 , \31276 );
buf \U$25862 ( \31492 , \31276 );
buf \U$25863 ( \31493 , \31276 );
buf \U$25864 ( \31494 , \31276 );
nor \U$25865 ( \31495 , \31304 , \31264 , \31265 , \31307 , \31269 , \31273 , \31276 , \31470 , \31471 , \31472 , \31473 , \31474 , \31475 , \31476 , \31477 , \31478 , \31479 , \31480 , \31481 , \31482 , \31483 , \31484 , \31485 , \31486 , \31487 , \31488 , \31489 , \31490 , \31491 , \31492 , \31493 , \31494 );
and \U$25866 ( \31496 , RIe5349b0_6879, \31495 );
buf \U$25867 ( \31497 , \31276 );
buf \U$25868 ( \31498 , \31276 );
buf \U$25869 ( \31499 , \31276 );
buf \U$25870 ( \31500 , \31276 );
buf \U$25871 ( \31501 , \31276 );
buf \U$25872 ( \31502 , \31276 );
buf \U$25873 ( \31503 , \31276 );
buf \U$25874 ( \31504 , \31276 );
buf \U$25875 ( \31505 , \31276 );
buf \U$25876 ( \31506 , \31276 );
buf \U$25877 ( \31507 , \31276 );
buf \U$25878 ( \31508 , \31276 );
buf \U$25879 ( \31509 , \31276 );
buf \U$25880 ( \31510 , \31276 );
buf \U$25881 ( \31511 , \31276 );
buf \U$25882 ( \31512 , \31276 );
buf \U$25883 ( \31513 , \31276 );
buf \U$25884 ( \31514 , \31276 );
buf \U$25885 ( \31515 , \31276 );
buf \U$25886 ( \31516 , \31276 );
buf \U$25887 ( \31517 , \31276 );
buf \U$25888 ( \31518 , \31276 );
buf \U$25889 ( \31519 , \31276 );
buf \U$25890 ( \31520 , \31276 );
buf \U$25891 ( \31521 , \31276 );
nor \U$25892 ( \31522 , \31263 , \31264 , \31265 , \31307 , \31269 , \31273 , \31276 , \31497 , \31498 , \31499 , \31500 , \31501 , \31502 , \31503 , \31504 , \31505 , \31506 , \31507 , \31508 , \31509 , \31510 , \31511 , \31512 , \31513 , \31514 , \31515 , \31516 , \31517 , \31518 , \31519 , \31520 , \31521 );
and \U$25893 ( \31523 , RIea94af8_6890, \31522 );
buf \U$25894 ( \31524 , \31276 );
buf \U$25895 ( \31525 , \31276 );
buf \U$25896 ( \31526 , \31276 );
buf \U$25897 ( \31527 , \31276 );
buf \U$25898 ( \31528 , \31276 );
buf \U$25899 ( \31529 , \31276 );
buf \U$25900 ( \31530 , \31276 );
buf \U$25901 ( \31531 , \31276 );
buf \U$25902 ( \31532 , \31276 );
buf \U$25903 ( \31533 , \31276 );
buf \U$25904 ( \31534 , \31276 );
buf \U$25905 ( \31535 , \31276 );
buf \U$25906 ( \31536 , \31276 );
buf \U$25907 ( \31537 , \31276 );
buf \U$25908 ( \31538 , \31276 );
buf \U$25909 ( \31539 , \31276 );
buf \U$25910 ( \31540 , \31276 );
buf \U$25911 ( \31541 , \31276 );
buf \U$25912 ( \31542 , \31276 );
buf \U$25913 ( \31543 , \31276 );
buf \U$25914 ( \31544 , \31276 );
buf \U$25915 ( \31545 , \31276 );
buf \U$25916 ( \31546 , \31276 );
buf \U$25917 ( \31547 , \31276 );
buf \U$25918 ( \31548 , \31276 );
nor \U$25919 ( \31549 , \31304 , \31305 , \31306 , \31266 , \31269 , \31273 , \31276 , \31524 , \31525 , \31526 , \31527 , \31528 , \31529 , \31530 , \31531 , \31532 , \31533 , \31534 , \31535 , \31536 , \31537 , \31538 , \31539 , \31540 , \31541 , \31542 , \31543 , \31544 , \31545 , \31546 , \31547 , \31548 );
and \U$25920 ( \31550 , RIe5351a8_6878, \31549 );
buf \U$25921 ( \31551 , \31276 );
buf \U$25922 ( \31552 , \31276 );
buf \U$25923 ( \31553 , \31276 );
buf \U$25924 ( \31554 , \31276 );
buf \U$25925 ( \31555 , \31276 );
buf \U$25926 ( \31556 , \31276 );
buf \U$25927 ( \31557 , \31276 );
buf \U$25928 ( \31558 , \31276 );
buf \U$25929 ( \31559 , \31276 );
buf \U$25930 ( \31560 , \31276 );
buf \U$25931 ( \31561 , \31276 );
buf \U$25932 ( \31562 , \31276 );
buf \U$25933 ( \31563 , \31276 );
buf \U$25934 ( \31564 , \31276 );
buf \U$25935 ( \31565 , \31276 );
buf \U$25936 ( \31566 , \31276 );
buf \U$25937 ( \31567 , \31276 );
buf \U$25938 ( \31568 , \31276 );
buf \U$25939 ( \31569 , \31276 );
buf \U$25940 ( \31570 , \31276 );
buf \U$25941 ( \31571 , \31276 );
buf \U$25942 ( \31572 , \31276 );
buf \U$25943 ( \31573 , \31276 );
buf \U$25944 ( \31574 , \31276 );
buf \U$25945 ( \31575 , \31276 );
nor \U$25946 ( \31576 , \31263 , \31305 , \31306 , \31266 , \31269 , \31273 , \31276 , \31551 , \31552 , \31553 , \31554 , \31555 , \31556 , \31557 , \31558 , \31559 , \31560 , \31561 , \31562 , \31563 , \31564 , \31565 , \31566 , \31567 , \31568 , \31569 , \31570 , \31571 , \31572 , \31573 , \31574 , \31575 );
and \U$25947 ( \31577 , RIe5359a0_6877, \31576 );
buf \U$25948 ( \31578 , \31276 );
buf \U$25949 ( \31579 , \31276 );
buf \U$25950 ( \31580 , \31276 );
buf \U$25951 ( \31581 , \31276 );
buf \U$25952 ( \31582 , \31276 );
buf \U$25953 ( \31583 , \31276 );
buf \U$25954 ( \31584 , \31276 );
buf \U$25955 ( \31585 , \31276 );
buf \U$25956 ( \31586 , \31276 );
buf \U$25957 ( \31587 , \31276 );
buf \U$25958 ( \31588 , \31276 );
buf \U$25959 ( \31589 , \31276 );
buf \U$25960 ( \31590 , \31276 );
buf \U$25961 ( \31591 , \31276 );
buf \U$25962 ( \31592 , \31276 );
buf \U$25963 ( \31593 , \31276 );
buf \U$25964 ( \31594 , \31276 );
buf \U$25965 ( \31595 , \31276 );
buf \U$25966 ( \31596 , \31276 );
buf \U$25967 ( \31597 , \31276 );
buf \U$25968 ( \31598 , \31276 );
buf \U$25969 ( \31599 , \31276 );
buf \U$25970 ( \31600 , \31276 );
buf \U$25971 ( \31601 , \31276 );
buf \U$25972 ( \31602 , \31276 );
nor \U$25973 ( \31603 , \31304 , \31264 , \31306 , \31266 , \31269 , \31273 , \31276 , \31578 , \31579 , \31580 , \31581 , \31582 , \31583 , \31584 , \31585 , \31586 , \31587 , \31588 , \31589 , \31590 , \31591 , \31592 , \31593 , \31594 , \31595 , \31596 , \31597 , \31598 , \31599 , \31600 , \31601 , \31602 );
and \U$25974 ( \31604 , RIeab78c8_6895, \31603 );
buf \U$25975 ( \31605 , \31276 );
buf \U$25976 ( \31606 , \31276 );
buf \U$25977 ( \31607 , \31276 );
buf \U$25978 ( \31608 , \31276 );
buf \U$25979 ( \31609 , \31276 );
buf \U$25980 ( \31610 , \31276 );
buf \U$25981 ( \31611 , \31276 );
buf \U$25982 ( \31612 , \31276 );
buf \U$25983 ( \31613 , \31276 );
buf \U$25984 ( \31614 , \31276 );
buf \U$25985 ( \31615 , \31276 );
buf \U$25986 ( \31616 , \31276 );
buf \U$25987 ( \31617 , \31276 );
buf \U$25988 ( \31618 , \31276 );
buf \U$25989 ( \31619 , \31276 );
buf \U$25990 ( \31620 , \31276 );
buf \U$25991 ( \31621 , \31276 );
buf \U$25992 ( \31622 , \31276 );
buf \U$25993 ( \31623 , \31276 );
buf \U$25994 ( \31624 , \31276 );
buf \U$25995 ( \31625 , \31276 );
buf \U$25996 ( \31626 , \31276 );
buf \U$25997 ( \31627 , \31276 );
buf \U$25998 ( \31628 , \31276 );
buf \U$25999 ( \31629 , \31276 );
nor \U$26000 ( \31630 , \31263 , \31264 , \31306 , \31266 , \31269 , \31273 , \31276 , \31605 , \31606 , \31607 , \31608 , \31609 , \31610 , \31611 , \31612 , \31613 , \31614 , \31615 , \31616 , \31617 , \31618 , \31619 , \31620 , \31621 , \31622 , \31623 , \31624 , \31625 , \31626 , \31627 , \31628 , \31629 );
and \U$26001 ( \31631 , RIeab7d00_6896, \31630 );
buf \U$26002 ( \31632 , \31276 );
buf \U$26003 ( \31633 , \31276 );
buf \U$26004 ( \31634 , \31276 );
buf \U$26005 ( \31635 , \31276 );
buf \U$26006 ( \31636 , \31276 );
buf \U$26007 ( \31637 , \31276 );
buf \U$26008 ( \31638 , \31276 );
buf \U$26009 ( \31639 , \31276 );
buf \U$26010 ( \31640 , \31276 );
buf \U$26011 ( \31641 , \31276 );
buf \U$26012 ( \31642 , \31276 );
buf \U$26013 ( \31643 , \31276 );
buf \U$26014 ( \31644 , \31276 );
buf \U$26015 ( \31645 , \31276 );
buf \U$26016 ( \31646 , \31276 );
buf \U$26017 ( \31647 , \31276 );
buf \U$26018 ( \31648 , \31276 );
buf \U$26019 ( \31649 , \31276 );
buf \U$26020 ( \31650 , \31276 );
buf \U$26021 ( \31651 , \31276 );
buf \U$26022 ( \31652 , \31276 );
buf \U$26023 ( \31653 , \31276 );
buf \U$26024 ( \31654 , \31276 );
buf \U$26025 ( \31655 , \31276 );
buf \U$26026 ( \31656 , \31276 );
nor \U$26027 ( \31657 , \31304 , \31305 , \31265 , \31266 , \31269 , \31273 , \31276 , \31632 , \31633 , \31634 , \31635 , \31636 , \31637 , \31638 , \31639 , \31640 , \31641 , \31642 , \31643 , \31644 , \31645 , \31646 , \31647 , \31648 , \31649 , \31650 , \31651 , \31652 , \31653 , \31654 , \31655 , \31656 );
and \U$26028 ( \31658 , RIeacfa18_6902, \31657 );
buf \U$26029 ( \31659 , \31276 );
buf \U$26030 ( \31660 , \31276 );
buf \U$26031 ( \31661 , \31276 );
buf \U$26032 ( \31662 , \31276 );
buf \U$26033 ( \31663 , \31276 );
buf \U$26034 ( \31664 , \31276 );
buf \U$26035 ( \31665 , \31276 );
buf \U$26036 ( \31666 , \31276 );
buf \U$26037 ( \31667 , \31276 );
buf \U$26038 ( \31668 , \31276 );
buf \U$26039 ( \31669 , \31276 );
buf \U$26040 ( \31670 , \31276 );
buf \U$26041 ( \31671 , \31276 );
buf \U$26042 ( \31672 , \31276 );
buf \U$26043 ( \31673 , \31276 );
buf \U$26044 ( \31674 , \31276 );
buf \U$26045 ( \31675 , \31276 );
buf \U$26046 ( \31676 , \31276 );
buf \U$26047 ( \31677 , \31276 );
buf \U$26048 ( \31678 , \31276 );
buf \U$26049 ( \31679 , \31276 );
buf \U$26050 ( \31680 , \31276 );
buf \U$26051 ( \31681 , \31276 );
buf \U$26052 ( \31682 , \31276 );
buf \U$26053 ( \31683 , \31276 );
nor \U$26054 ( \31684 , \31263 , \31305 , \31265 , \31266 , \31269 , \31273 , \31276 , \31659 , \31660 , \31661 , \31662 , \31663 , \31664 , \31665 , \31666 , \31667 , \31668 , \31669 , \31670 , \31671 , \31672 , \31673 , \31674 , \31675 , \31676 , \31677 , \31678 , \31679 , \31680 , \31681 , \31682 , \31683 );
and \U$26055 ( \31685 , RIeab6518_6891, \31684 );
buf \U$26056 ( \31686 , \31276 );
buf \U$26057 ( \31687 , \31276 );
buf \U$26058 ( \31688 , \31276 );
buf \U$26059 ( \31689 , \31276 );
buf \U$26060 ( \31690 , \31276 );
buf \U$26061 ( \31691 , \31276 );
buf \U$26062 ( \31692 , \31276 );
buf \U$26063 ( \31693 , \31276 );
buf \U$26064 ( \31694 , \31276 );
buf \U$26065 ( \31695 , \31276 );
buf \U$26066 ( \31696 , \31276 );
buf \U$26067 ( \31697 , \31276 );
buf \U$26068 ( \31698 , \31276 );
buf \U$26069 ( \31699 , \31276 );
buf \U$26070 ( \31700 , \31276 );
buf \U$26071 ( \31701 , \31276 );
buf \U$26072 ( \31702 , \31276 );
buf \U$26073 ( \31703 , \31276 );
buf \U$26074 ( \31704 , \31276 );
buf \U$26075 ( \31705 , \31276 );
buf \U$26076 ( \31706 , \31276 );
buf \U$26077 ( \31707 , \31276 );
buf \U$26078 ( \31708 , \31276 );
buf \U$26079 ( \31709 , \31276 );
buf \U$26080 ( \31710 , \31276 );
nor \U$26081 ( \31711 , \31304 , \31264 , \31265 , \31266 , \31269 , \31273 , \31276 , \31686 , \31687 , \31688 , \31689 , \31690 , \31691 , \31692 , \31693 , \31694 , \31695 , \31696 , \31697 , \31698 , \31699 , \31700 , \31701 , \31702 , \31703 , \31704 , \31705 , \31706 , \31707 , \31708 , \31709 , \31710 );
and \U$26082 ( \31712 , RIeb352c8_6904, \31711 );
or \U$26083 ( \31713 , \31303 , \31334 , \31361 , \31388 , \31415 , \31442 , \31469 , \31496 , \31523 , \31550 , \31577 , \31604 , \31631 , \31658 , \31685 , \31712 );
buf \U$26084 ( \31714 , \31276 );
not \U$26085 ( \31715 , \31714 );
buf \U$26086 ( \31716 , \31264 );
buf \U$26087 ( \31717 , \31265 );
buf \U$26088 ( \31718 , \31266 );
buf \U$26089 ( \31719 , \31269 );
buf \U$26090 ( \31720 , \31273 );
buf \U$26091 ( \31721 , \31276 );
buf \U$26092 ( \31722 , \31276 );
buf \U$26093 ( \31723 , \31276 );
buf \U$26094 ( \31724 , \31276 );
buf \U$26095 ( \31725 , \31276 );
buf \U$26096 ( \31726 , \31276 );
buf \U$26097 ( \31727 , \31276 );
buf \U$26098 ( \31728 , \31276 );
buf \U$26099 ( \31729 , \31276 );
buf \U$26100 ( \31730 , \31276 );
buf \U$26101 ( \31731 , \31276 );
buf \U$26102 ( \31732 , \31276 );
buf \U$26103 ( \31733 , \31276 );
buf \U$26104 ( \31734 , \31276 );
buf \U$26105 ( \31735 , \31276 );
buf \U$26106 ( \31736 , \31276 );
buf \U$26107 ( \31737 , \31276 );
buf \U$26108 ( \31738 , \31276 );
buf \U$26109 ( \31739 , \31276 );
buf \U$26110 ( \31740 , \31276 );
buf \U$26111 ( \31741 , \31276 );
buf \U$26112 ( \31742 , \31276 );
buf \U$26113 ( \31743 , \31276 );
buf \U$26114 ( \31744 , \31276 );
buf \U$26115 ( \31745 , \31276 );
buf \U$26116 ( \31746 , \31263 );
or \U$26117 ( \31747 , \31716 , \31717 , \31718 , \31719 , \31720 , \31721 , \31722 , \31723 , \31724 , \31725 , \31726 , \31727 , \31728 , \31729 , \31730 , \31731 , \31732 , \31733 , \31734 , \31735 , \31736 , \31737 , \31738 , \31739 , \31740 , \31741 , \31742 , \31743 , \31744 , \31745 , \31746 );
nand \U$26118 ( \31748 , \31715 , \31747 );
buf \U$26119 ( \31749 , \31748 );
buf \U$26120 ( \31750 , \31276 );
not \U$26121 ( \31751 , \31750 );
buf \U$26122 ( \31752 , \31273 );
buf \U$26123 ( \31753 , \31276 );
buf \U$26124 ( \31754 , \31276 );
buf \U$26125 ( \31755 , \31276 );
buf \U$26126 ( \31756 , \31276 );
buf \U$26127 ( \31757 , \31276 );
buf \U$26128 ( \31758 , \31276 );
buf \U$26129 ( \31759 , \31276 );
buf \U$26130 ( \31760 , \31276 );
buf \U$26131 ( \31761 , \31276 );
buf \U$26132 ( \31762 , \31276 );
buf \U$26133 ( \31763 , \31276 );
buf \U$26134 ( \31764 , \31276 );
buf \U$26135 ( \31765 , \31276 );
buf \U$26136 ( \31766 , \31276 );
buf \U$26137 ( \31767 , \31276 );
buf \U$26138 ( \31768 , \31276 );
buf \U$26139 ( \31769 , \31276 );
buf \U$26140 ( \31770 , \31276 );
buf \U$26141 ( \31771 , \31276 );
buf \U$26142 ( \31772 , \31276 );
buf \U$26143 ( \31773 , \31276 );
buf \U$26144 ( \31774 , \31276 );
buf \U$26145 ( \31775 , \31276 );
buf \U$26146 ( \31776 , \31276 );
buf \U$26147 ( \31777 , \31276 );
buf \U$26148 ( \31778 , \31269 );
buf \U$26149 ( \31779 , \31263 );
buf \U$26150 ( \31780 , \31264 );
buf \U$26151 ( \31781 , \31265 );
buf \U$26152 ( \31782 , \31266 );
or \U$26153 ( \31783 , \31779 , \31780 , \31781 , \31782 );
and \U$26154 ( \31784 , \31778 , \31783 );
or \U$26155 ( \31785 , \31752 , \31753 , \31754 , \31755 , \31756 , \31757 , \31758 , \31759 , \31760 , \31761 , \31762 , \31763 , \31764 , \31765 , \31766 , \31767 , \31768 , \31769 , \31770 , \31771 , \31772 , \31773 , \31774 , \31775 , \31776 , \31777 , \31784 );
and \U$26156 ( \31786 , \31751 , \31785 );
buf \U$26157 ( \31787 , \31786 );
or \U$26158 ( \31788 , \31749 , \31787 );
_DC g9340 ( \31789_nG9340 , \31713 , \31788 );
not \U$26159 ( \31790 , \31789_nG9340 );
buf \U$26160 ( \31791 , RIb7b9608_246);
buf \U$26161 ( \31792 , \31276 );
buf \U$26162 ( \31793 , \31276 );
buf \U$26163 ( \31794 , \31276 );
buf \U$26164 ( \31795 , \31276 );
buf \U$26165 ( \31796 , \31276 );
buf \U$26166 ( \31797 , \31276 );
buf \U$26167 ( \31798 , \31276 );
buf \U$26168 ( \31799 , \31276 );
buf \U$26169 ( \31800 , \31276 );
buf \U$26170 ( \31801 , \31276 );
buf \U$26171 ( \31802 , \31276 );
buf \U$26172 ( \31803 , \31276 );
buf \U$26173 ( \31804 , \31276 );
buf \U$26174 ( \31805 , \31276 );
buf \U$26175 ( \31806 , \31276 );
buf \U$26176 ( \31807 , \31276 );
buf \U$26177 ( \31808 , \31276 );
buf \U$26178 ( \31809 , \31276 );
buf \U$26179 ( \31810 , \31276 );
buf \U$26180 ( \31811 , \31276 );
buf \U$26181 ( \31812 , \31276 );
buf \U$26182 ( \31813 , \31276 );
buf \U$26183 ( \31814 , \31276 );
buf \U$26184 ( \31815 , \31276 );
buf \U$26185 ( \31816 , \31276 );
nor \U$26186 ( \31817 , \31263 , \31264 , \31265 , \31266 , \31270 , \31273 , \31276 , \31792 , \31793 , \31794 , \31795 , \31796 , \31797 , \31798 , \31799 , \31800 , \31801 , \31802 , \31803 , \31804 , \31805 , \31806 , \31807 , \31808 , \31809 , \31810 , \31811 , \31812 , \31813 , \31814 , \31815 , \31816 );
and \U$26187 ( \31818 , \7117 , \31817 );
buf \U$26188 ( \31819 , \31276 );
buf \U$26189 ( \31820 , \31276 );
buf \U$26190 ( \31821 , \31276 );
buf \U$26191 ( \31822 , \31276 );
buf \U$26192 ( \31823 , \31276 );
buf \U$26193 ( \31824 , \31276 );
buf \U$26194 ( \31825 , \31276 );
buf \U$26195 ( \31826 , \31276 );
buf \U$26196 ( \31827 , \31276 );
buf \U$26197 ( \31828 , \31276 );
buf \U$26198 ( \31829 , \31276 );
buf \U$26199 ( \31830 , \31276 );
buf \U$26200 ( \31831 , \31276 );
buf \U$26201 ( \31832 , \31276 );
buf \U$26202 ( \31833 , \31276 );
buf \U$26203 ( \31834 , \31276 );
buf \U$26204 ( \31835 , \31276 );
buf \U$26205 ( \31836 , \31276 );
buf \U$26206 ( \31837 , \31276 );
buf \U$26207 ( \31838 , \31276 );
buf \U$26208 ( \31839 , \31276 );
buf \U$26209 ( \31840 , \31276 );
buf \U$26210 ( \31841 , \31276 );
buf \U$26211 ( \31842 , \31276 );
buf \U$26212 ( \31843 , \31276 );
nor \U$26213 ( \31844 , \31304 , \31305 , \31306 , \31307 , \31269 , \31273 , \31276 , \31819 , \31820 , \31821 , \31822 , \31823 , \31824 , \31825 , \31826 , \31827 , \31828 , \31829 , \31830 , \31831 , \31832 , \31833 , \31834 , \31835 , \31836 , \31837 , \31838 , \31839 , \31840 , \31841 , \31842 , \31843 );
and \U$26214 ( \31845 , \7119 , \31844 );
buf \U$26215 ( \31846 , \31276 );
buf \U$26216 ( \31847 , \31276 );
buf \U$26217 ( \31848 , \31276 );
buf \U$26218 ( \31849 , \31276 );
buf \U$26219 ( \31850 , \31276 );
buf \U$26220 ( \31851 , \31276 );
buf \U$26221 ( \31852 , \31276 );
buf \U$26222 ( \31853 , \31276 );
buf \U$26223 ( \31854 , \31276 );
buf \U$26224 ( \31855 , \31276 );
buf \U$26225 ( \31856 , \31276 );
buf \U$26226 ( \31857 , \31276 );
buf \U$26227 ( \31858 , \31276 );
buf \U$26228 ( \31859 , \31276 );
buf \U$26229 ( \31860 , \31276 );
buf \U$26230 ( \31861 , \31276 );
buf \U$26231 ( \31862 , \31276 );
buf \U$26232 ( \31863 , \31276 );
buf \U$26233 ( \31864 , \31276 );
buf \U$26234 ( \31865 , \31276 );
buf \U$26235 ( \31866 , \31276 );
buf \U$26236 ( \31867 , \31276 );
buf \U$26237 ( \31868 , \31276 );
buf \U$26238 ( \31869 , \31276 );
buf \U$26239 ( \31870 , \31276 );
nor \U$26240 ( \31871 , \31263 , \31305 , \31306 , \31307 , \31269 , \31273 , \31276 , \31846 , \31847 , \31848 , \31849 , \31850 , \31851 , \31852 , \31853 , \31854 , \31855 , \31856 , \31857 , \31858 , \31859 , \31860 , \31861 , \31862 , \31863 , \31864 , \31865 , \31866 , \31867 , \31868 , \31869 , \31870 );
and \U$26241 ( \31872 , \7864 , \31871 );
buf \U$26242 ( \31873 , \31276 );
buf \U$26243 ( \31874 , \31276 );
buf \U$26244 ( \31875 , \31276 );
buf \U$26245 ( \31876 , \31276 );
buf \U$26246 ( \31877 , \31276 );
buf \U$26247 ( \31878 , \31276 );
buf \U$26248 ( \31879 , \31276 );
buf \U$26249 ( \31880 , \31276 );
buf \U$26250 ( \31881 , \31276 );
buf \U$26251 ( \31882 , \31276 );
buf \U$26252 ( \31883 , \31276 );
buf \U$26253 ( \31884 , \31276 );
buf \U$26254 ( \31885 , \31276 );
buf \U$26255 ( \31886 , \31276 );
buf \U$26256 ( \31887 , \31276 );
buf \U$26257 ( \31888 , \31276 );
buf \U$26258 ( \31889 , \31276 );
buf \U$26259 ( \31890 , \31276 );
buf \U$26260 ( \31891 , \31276 );
buf \U$26261 ( \31892 , \31276 );
buf \U$26262 ( \31893 , \31276 );
buf \U$26263 ( \31894 , \31276 );
buf \U$26264 ( \31895 , \31276 );
buf \U$26265 ( \31896 , \31276 );
buf \U$26266 ( \31897 , \31276 );
nor \U$26267 ( \31898 , \31304 , \31264 , \31306 , \31307 , \31269 , \31273 , \31276 , \31873 , \31874 , \31875 , \31876 , \31877 , \31878 , \31879 , \31880 , \31881 , \31882 , \31883 , \31884 , \31885 , \31886 , \31887 , \31888 , \31889 , \31890 , \31891 , \31892 , \31893 , \31894 , \31895 , \31896 , \31897 );
and \U$26268 ( \31899 , \7892 , \31898 );
buf \U$26269 ( \31900 , \31276 );
buf \U$26270 ( \31901 , \31276 );
buf \U$26271 ( \31902 , \31276 );
buf \U$26272 ( \31903 , \31276 );
buf \U$26273 ( \31904 , \31276 );
buf \U$26274 ( \31905 , \31276 );
buf \U$26275 ( \31906 , \31276 );
buf \U$26276 ( \31907 , \31276 );
buf \U$26277 ( \31908 , \31276 );
buf \U$26278 ( \31909 , \31276 );
buf \U$26279 ( \31910 , \31276 );
buf \U$26280 ( \31911 , \31276 );
buf \U$26281 ( \31912 , \31276 );
buf \U$26282 ( \31913 , \31276 );
buf \U$26283 ( \31914 , \31276 );
buf \U$26284 ( \31915 , \31276 );
buf \U$26285 ( \31916 , \31276 );
buf \U$26286 ( \31917 , \31276 );
buf \U$26287 ( \31918 , \31276 );
buf \U$26288 ( \31919 , \31276 );
buf \U$26289 ( \31920 , \31276 );
buf \U$26290 ( \31921 , \31276 );
buf \U$26291 ( \31922 , \31276 );
buf \U$26292 ( \31923 , \31276 );
buf \U$26293 ( \31924 , \31276 );
nor \U$26294 ( \31925 , \31263 , \31264 , \31306 , \31307 , \31269 , \31273 , \31276 , \31900 , \31901 , \31902 , \31903 , \31904 , \31905 , \31906 , \31907 , \31908 , \31909 , \31910 , \31911 , \31912 , \31913 , \31914 , \31915 , \31916 , \31917 , \31918 , \31919 , \31920 , \31921 , \31922 , \31923 , \31924 );
and \U$26295 ( \31926 , \7920 , \31925 );
buf \U$26296 ( \31927 , \31276 );
buf \U$26297 ( \31928 , \31276 );
buf \U$26298 ( \31929 , \31276 );
buf \U$26299 ( \31930 , \31276 );
buf \U$26300 ( \31931 , \31276 );
buf \U$26301 ( \31932 , \31276 );
buf \U$26302 ( \31933 , \31276 );
buf \U$26303 ( \31934 , \31276 );
buf \U$26304 ( \31935 , \31276 );
buf \U$26305 ( \31936 , \31276 );
buf \U$26306 ( \31937 , \31276 );
buf \U$26307 ( \31938 , \31276 );
buf \U$26308 ( \31939 , \31276 );
buf \U$26309 ( \31940 , \31276 );
buf \U$26310 ( \31941 , \31276 );
buf \U$26311 ( \31942 , \31276 );
buf \U$26312 ( \31943 , \31276 );
buf \U$26313 ( \31944 , \31276 );
buf \U$26314 ( \31945 , \31276 );
buf \U$26315 ( \31946 , \31276 );
buf \U$26316 ( \31947 , \31276 );
buf \U$26317 ( \31948 , \31276 );
buf \U$26318 ( \31949 , \31276 );
buf \U$26319 ( \31950 , \31276 );
buf \U$26320 ( \31951 , \31276 );
nor \U$26321 ( \31952 , \31304 , \31305 , \31265 , \31307 , \31269 , \31273 , \31276 , \31927 , \31928 , \31929 , \31930 , \31931 , \31932 , \31933 , \31934 , \31935 , \31936 , \31937 , \31938 , \31939 , \31940 , \31941 , \31942 , \31943 , \31944 , \31945 , \31946 , \31947 , \31948 , \31949 , \31950 , \31951 );
and \U$26322 ( \31953 , \7948 , \31952 );
buf \U$26323 ( \31954 , \31276 );
buf \U$26324 ( \31955 , \31276 );
buf \U$26325 ( \31956 , \31276 );
buf \U$26326 ( \31957 , \31276 );
buf \U$26327 ( \31958 , \31276 );
buf \U$26328 ( \31959 , \31276 );
buf \U$26329 ( \31960 , \31276 );
buf \U$26330 ( \31961 , \31276 );
buf \U$26331 ( \31962 , \31276 );
buf \U$26332 ( \31963 , \31276 );
buf \U$26333 ( \31964 , \31276 );
buf \U$26334 ( \31965 , \31276 );
buf \U$26335 ( \31966 , \31276 );
buf \U$26336 ( \31967 , \31276 );
buf \U$26337 ( \31968 , \31276 );
buf \U$26338 ( \31969 , \31276 );
buf \U$26339 ( \31970 , \31276 );
buf \U$26340 ( \31971 , \31276 );
buf \U$26341 ( \31972 , \31276 );
buf \U$26342 ( \31973 , \31276 );
buf \U$26343 ( \31974 , \31276 );
buf \U$26344 ( \31975 , \31276 );
buf \U$26345 ( \31976 , \31276 );
buf \U$26346 ( \31977 , \31276 );
buf \U$26347 ( \31978 , \31276 );
nor \U$26348 ( \31979 , \31263 , \31305 , \31265 , \31307 , \31269 , \31273 , \31276 , \31954 , \31955 , \31956 , \31957 , \31958 , \31959 , \31960 , \31961 , \31962 , \31963 , \31964 , \31965 , \31966 , \31967 , \31968 , \31969 , \31970 , \31971 , \31972 , \31973 , \31974 , \31975 , \31976 , \31977 , \31978 );
and \U$26349 ( \31980 , \7976 , \31979 );
buf \U$26350 ( \31981 , \31276 );
buf \U$26351 ( \31982 , \31276 );
buf \U$26352 ( \31983 , \31276 );
buf \U$26353 ( \31984 , \31276 );
buf \U$26354 ( \31985 , \31276 );
buf \U$26355 ( \31986 , \31276 );
buf \U$26356 ( \31987 , \31276 );
buf \U$26357 ( \31988 , \31276 );
buf \U$26358 ( \31989 , \31276 );
buf \U$26359 ( \31990 , \31276 );
buf \U$26360 ( \31991 , \31276 );
buf \U$26361 ( \31992 , \31276 );
buf \U$26362 ( \31993 , \31276 );
buf \U$26363 ( \31994 , \31276 );
buf \U$26364 ( \31995 , \31276 );
buf \U$26365 ( \31996 , \31276 );
buf \U$26366 ( \31997 , \31276 );
buf \U$26367 ( \31998 , \31276 );
buf \U$26368 ( \31999 , \31276 );
buf \U$26369 ( \32000 , \31276 );
buf \U$26370 ( \32001 , \31276 );
buf \U$26371 ( \32002 , \31276 );
buf \U$26372 ( \32003 , \31276 );
buf \U$26373 ( \32004 , \31276 );
buf \U$26374 ( \32005 , \31276 );
nor \U$26375 ( \32006 , \31304 , \31264 , \31265 , \31307 , \31269 , \31273 , \31276 , \31981 , \31982 , \31983 , \31984 , \31985 , \31986 , \31987 , \31988 , \31989 , \31990 , \31991 , \31992 , \31993 , \31994 , \31995 , \31996 , \31997 , \31998 , \31999 , \32000 , \32001 , \32002 , \32003 , \32004 , \32005 );
and \U$26376 ( \32007 , \8004 , \32006 );
buf \U$26377 ( \32008 , \31276 );
buf \U$26378 ( \32009 , \31276 );
buf \U$26379 ( \32010 , \31276 );
buf \U$26380 ( \32011 , \31276 );
buf \U$26381 ( \32012 , \31276 );
buf \U$26382 ( \32013 , \31276 );
buf \U$26383 ( \32014 , \31276 );
buf \U$26384 ( \32015 , \31276 );
buf \U$26385 ( \32016 , \31276 );
buf \U$26386 ( \32017 , \31276 );
buf \U$26387 ( \32018 , \31276 );
buf \U$26388 ( \32019 , \31276 );
buf \U$26389 ( \32020 , \31276 );
buf \U$26390 ( \32021 , \31276 );
buf \U$26391 ( \32022 , \31276 );
buf \U$26392 ( \32023 , \31276 );
buf \U$26393 ( \32024 , \31276 );
buf \U$26394 ( \32025 , \31276 );
buf \U$26395 ( \32026 , \31276 );
buf \U$26396 ( \32027 , \31276 );
buf \U$26397 ( \32028 , \31276 );
buf \U$26398 ( \32029 , \31276 );
buf \U$26399 ( \32030 , \31276 );
buf \U$26400 ( \32031 , \31276 );
buf \U$26401 ( \32032 , \31276 );
nor \U$26402 ( \32033 , \31263 , \31264 , \31265 , \31307 , \31269 , \31273 , \31276 , \32008 , \32009 , \32010 , \32011 , \32012 , \32013 , \32014 , \32015 , \32016 , \32017 , \32018 , \32019 , \32020 , \32021 , \32022 , \32023 , \32024 , \32025 , \32026 , \32027 , \32028 , \32029 , \32030 , \32031 , \32032 );
and \U$26403 ( \32034 , \8032 , \32033 );
buf \U$26404 ( \32035 , \31276 );
buf \U$26405 ( \32036 , \31276 );
buf \U$26406 ( \32037 , \31276 );
buf \U$26407 ( \32038 , \31276 );
buf \U$26408 ( \32039 , \31276 );
buf \U$26409 ( \32040 , \31276 );
buf \U$26410 ( \32041 , \31276 );
buf \U$26411 ( \32042 , \31276 );
buf \U$26412 ( \32043 , \31276 );
buf \U$26413 ( \32044 , \31276 );
buf \U$26414 ( \32045 , \31276 );
buf \U$26415 ( \32046 , \31276 );
buf \U$26416 ( \32047 , \31276 );
buf \U$26417 ( \32048 , \31276 );
buf \U$26418 ( \32049 , \31276 );
buf \U$26419 ( \32050 , \31276 );
buf \U$26420 ( \32051 , \31276 );
buf \U$26421 ( \32052 , \31276 );
buf \U$26422 ( \32053 , \31276 );
buf \U$26423 ( \32054 , \31276 );
buf \U$26424 ( \32055 , \31276 );
buf \U$26425 ( \32056 , \31276 );
buf \U$26426 ( \32057 , \31276 );
buf \U$26427 ( \32058 , \31276 );
buf \U$26428 ( \32059 , \31276 );
nor \U$26429 ( \32060 , \31304 , \31305 , \31306 , \31266 , \31269 , \31273 , \31276 , \32035 , \32036 , \32037 , \32038 , \32039 , \32040 , \32041 , \32042 , \32043 , \32044 , \32045 , \32046 , \32047 , \32048 , \32049 , \32050 , \32051 , \32052 , \32053 , \32054 , \32055 , \32056 , \32057 , \32058 , \32059 );
and \U$26430 ( \32061 , \8060 , \32060 );
buf \U$26431 ( \32062 , \31276 );
buf \U$26432 ( \32063 , \31276 );
buf \U$26433 ( \32064 , \31276 );
buf \U$26434 ( \32065 , \31276 );
buf \U$26435 ( \32066 , \31276 );
buf \U$26436 ( \32067 , \31276 );
buf \U$26437 ( \32068 , \31276 );
buf \U$26438 ( \32069 , \31276 );
buf \U$26439 ( \32070 , \31276 );
buf \U$26440 ( \32071 , \31276 );
buf \U$26441 ( \32072 , \31276 );
buf \U$26442 ( \32073 , \31276 );
buf \U$26443 ( \32074 , \31276 );
buf \U$26444 ( \32075 , \31276 );
buf \U$26445 ( \32076 , \31276 );
buf \U$26446 ( \32077 , \31276 );
buf \U$26447 ( \32078 , \31276 );
buf \U$26448 ( \32079 , \31276 );
buf \U$26449 ( \32080 , \31276 );
buf \U$26450 ( \32081 , \31276 );
buf \U$26451 ( \32082 , \31276 );
buf \U$26452 ( \32083 , \31276 );
buf \U$26453 ( \32084 , \31276 );
buf \U$26454 ( \32085 , \31276 );
buf \U$26455 ( \32086 , \31276 );
nor \U$26456 ( \32087 , \31263 , \31305 , \31306 , \31266 , \31269 , \31273 , \31276 , \32062 , \32063 , \32064 , \32065 , \32066 , \32067 , \32068 , \32069 , \32070 , \32071 , \32072 , \32073 , \32074 , \32075 , \32076 , \32077 , \32078 , \32079 , \32080 , \32081 , \32082 , \32083 , \32084 , \32085 , \32086 );
and \U$26457 ( \32088 , \8088 , \32087 );
buf \U$26458 ( \32089 , \31276 );
buf \U$26459 ( \32090 , \31276 );
buf \U$26460 ( \32091 , \31276 );
buf \U$26461 ( \32092 , \31276 );
buf \U$26462 ( \32093 , \31276 );
buf \U$26463 ( \32094 , \31276 );
buf \U$26464 ( \32095 , \31276 );
buf \U$26465 ( \32096 , \31276 );
buf \U$26466 ( \32097 , \31276 );
buf \U$26467 ( \32098 , \31276 );
buf \U$26468 ( \32099 , \31276 );
buf \U$26469 ( \32100 , \31276 );
buf \U$26470 ( \32101 , \31276 );
buf \U$26471 ( \32102 , \31276 );
buf \U$26472 ( \32103 , \31276 );
buf \U$26473 ( \32104 , \31276 );
buf \U$26474 ( \32105 , \31276 );
buf \U$26475 ( \32106 , \31276 );
buf \U$26476 ( \32107 , \31276 );
buf \U$26477 ( \32108 , \31276 );
buf \U$26478 ( \32109 , \31276 );
buf \U$26479 ( \32110 , \31276 );
buf \U$26480 ( \32111 , \31276 );
buf \U$26481 ( \32112 , \31276 );
buf \U$26482 ( \32113 , \31276 );
nor \U$26483 ( \32114 , \31304 , \31264 , \31306 , \31266 , \31269 , \31273 , \31276 , \32089 , \32090 , \32091 , \32092 , \32093 , \32094 , \32095 , \32096 , \32097 , \32098 , \32099 , \32100 , \32101 , \32102 , \32103 , \32104 , \32105 , \32106 , \32107 , \32108 , \32109 , \32110 , \32111 , \32112 , \32113 );
and \U$26484 ( \32115 , \8116 , \32114 );
buf \U$26485 ( \32116 , \31276 );
buf \U$26486 ( \32117 , \31276 );
buf \U$26487 ( \32118 , \31276 );
buf \U$26488 ( \32119 , \31276 );
buf \U$26489 ( \32120 , \31276 );
buf \U$26490 ( \32121 , \31276 );
buf \U$26491 ( \32122 , \31276 );
buf \U$26492 ( \32123 , \31276 );
buf \U$26493 ( \32124 , \31276 );
buf \U$26494 ( \32125 , \31276 );
buf \U$26495 ( \32126 , \31276 );
buf \U$26496 ( \32127 , \31276 );
buf \U$26497 ( \32128 , \31276 );
buf \U$26498 ( \32129 , \31276 );
buf \U$26499 ( \32130 , \31276 );
buf \U$26500 ( \32131 , \31276 );
buf \U$26501 ( \32132 , \31276 );
buf \U$26502 ( \32133 , \31276 );
buf \U$26503 ( \32134 , \31276 );
buf \U$26504 ( \32135 , \31276 );
buf \U$26505 ( \32136 , \31276 );
buf \U$26506 ( \32137 , \31276 );
buf \U$26507 ( \32138 , \31276 );
buf \U$26508 ( \32139 , \31276 );
buf \U$26509 ( \32140 , \31276 );
nor \U$26510 ( \32141 , \31263 , \31264 , \31306 , \31266 , \31269 , \31273 , \31276 , \32116 , \32117 , \32118 , \32119 , \32120 , \32121 , \32122 , \32123 , \32124 , \32125 , \32126 , \32127 , \32128 , \32129 , \32130 , \32131 , \32132 , \32133 , \32134 , \32135 , \32136 , \32137 , \32138 , \32139 , \32140 );
and \U$26511 ( \32142 , \8144 , \32141 );
buf \U$26512 ( \32143 , \31276 );
buf \U$26513 ( \32144 , \31276 );
buf \U$26514 ( \32145 , \31276 );
buf \U$26515 ( \32146 , \31276 );
buf \U$26516 ( \32147 , \31276 );
buf \U$26517 ( \32148 , \31276 );
buf \U$26518 ( \32149 , \31276 );
buf \U$26519 ( \32150 , \31276 );
buf \U$26520 ( \32151 , \31276 );
buf \U$26521 ( \32152 , \31276 );
buf \U$26522 ( \32153 , \31276 );
buf \U$26523 ( \32154 , \31276 );
buf \U$26524 ( \32155 , \31276 );
buf \U$26525 ( \32156 , \31276 );
buf \U$26526 ( \32157 , \31276 );
buf \U$26527 ( \32158 , \31276 );
buf \U$26528 ( \32159 , \31276 );
buf \U$26529 ( \32160 , \31276 );
buf \U$26530 ( \32161 , \31276 );
buf \U$26531 ( \32162 , \31276 );
buf \U$26532 ( \32163 , \31276 );
buf \U$26533 ( \32164 , \31276 );
buf \U$26534 ( \32165 , \31276 );
buf \U$26535 ( \32166 , \31276 );
buf \U$26536 ( \32167 , \31276 );
nor \U$26537 ( \32168 , \31304 , \31305 , \31265 , \31266 , \31269 , \31273 , \31276 , \32143 , \32144 , \32145 , \32146 , \32147 , \32148 , \32149 , \32150 , \32151 , \32152 , \32153 , \32154 , \32155 , \32156 , \32157 , \32158 , \32159 , \32160 , \32161 , \32162 , \32163 , \32164 , \32165 , \32166 , \32167 );
and \U$26538 ( \32169 , \8172 , \32168 );
buf \U$26539 ( \32170 , \31276 );
buf \U$26540 ( \32171 , \31276 );
buf \U$26541 ( \32172 , \31276 );
buf \U$26542 ( \32173 , \31276 );
buf \U$26543 ( \32174 , \31276 );
buf \U$26544 ( \32175 , \31276 );
buf \U$26545 ( \32176 , \31276 );
buf \U$26546 ( \32177 , \31276 );
buf \U$26547 ( \32178 , \31276 );
buf \U$26548 ( \32179 , \31276 );
buf \U$26549 ( \32180 , \31276 );
buf \U$26550 ( \32181 , \31276 );
buf \U$26551 ( \32182 , \31276 );
buf \U$26552 ( \32183 , \31276 );
buf \U$26553 ( \32184 , \31276 );
buf \U$26554 ( \32185 , \31276 );
buf \U$26555 ( \32186 , \31276 );
buf \U$26556 ( \32187 , \31276 );
buf \U$26557 ( \32188 , \31276 );
buf \U$26558 ( \32189 , \31276 );
buf \U$26559 ( \32190 , \31276 );
buf \U$26560 ( \32191 , \31276 );
buf \U$26561 ( \32192 , \31276 );
buf \U$26562 ( \32193 , \31276 );
buf \U$26563 ( \32194 , \31276 );
nor \U$26564 ( \32195 , \31263 , \31305 , \31265 , \31266 , \31269 , \31273 , \31276 , \32170 , \32171 , \32172 , \32173 , \32174 , \32175 , \32176 , \32177 , \32178 , \32179 , \32180 , \32181 , \32182 , \32183 , \32184 , \32185 , \32186 , \32187 , \32188 , \32189 , \32190 , \32191 , \32192 , \32193 , \32194 );
and \U$26565 ( \32196 , \8200 , \32195 );
buf \U$26566 ( \32197 , \31276 );
buf \U$26567 ( \32198 , \31276 );
buf \U$26568 ( \32199 , \31276 );
buf \U$26569 ( \32200 , \31276 );
buf \U$26570 ( \32201 , \31276 );
buf \U$26571 ( \32202 , \31276 );
buf \U$26572 ( \32203 , \31276 );
buf \U$26573 ( \32204 , \31276 );
buf \U$26574 ( \32205 , \31276 );
buf \U$26575 ( \32206 , \31276 );
buf \U$26576 ( \32207 , \31276 );
buf \U$26577 ( \32208 , \31276 );
buf \U$26578 ( \32209 , \31276 );
buf \U$26579 ( \32210 , \31276 );
buf \U$26580 ( \32211 , \31276 );
buf \U$26581 ( \32212 , \31276 );
buf \U$26582 ( \32213 , \31276 );
buf \U$26583 ( \32214 , \31276 );
buf \U$26584 ( \32215 , \31276 );
buf \U$26585 ( \32216 , \31276 );
buf \U$26586 ( \32217 , \31276 );
buf \U$26587 ( \32218 , \31276 );
buf \U$26588 ( \32219 , \31276 );
buf \U$26589 ( \32220 , \31276 );
buf \U$26590 ( \32221 , \31276 );
nor \U$26591 ( \32222 , \31304 , \31264 , \31265 , \31266 , \31269 , \31273 , \31276 , \32197 , \32198 , \32199 , \32200 , \32201 , \32202 , \32203 , \32204 , \32205 , \32206 , \32207 , \32208 , \32209 , \32210 , \32211 , \32212 , \32213 , \32214 , \32215 , \32216 , \32217 , \32218 , \32219 , \32220 , \32221 );
and \U$26592 ( \32223 , \8228 , \32222 );
or \U$26593 ( \32224 , \31818 , \31845 , \31872 , \31899 , \31926 , \31953 , \31980 , \32007 , \32034 , \32061 , \32088 , \32115 , \32142 , \32169 , \32196 , \32223 );
buf \U$26594 ( \32225 , \31276 );
not \U$26595 ( \32226 , \32225 );
buf \U$26596 ( \32227 , \31264 );
buf \U$26597 ( \32228 , \31265 );
buf \U$26598 ( \32229 , \31266 );
buf \U$26599 ( \32230 , \31269 );
buf \U$26600 ( \32231 , \31273 );
buf \U$26601 ( \32232 , \31276 );
buf \U$26602 ( \32233 , \31276 );
buf \U$26603 ( \32234 , \31276 );
buf \U$26604 ( \32235 , \31276 );
buf \U$26605 ( \32236 , \31276 );
buf \U$26606 ( \32237 , \31276 );
buf \U$26607 ( \32238 , \31276 );
buf \U$26608 ( \32239 , \31276 );
buf \U$26609 ( \32240 , \31276 );
buf \U$26610 ( \32241 , \31276 );
buf \U$26611 ( \32242 , \31276 );
buf \U$26612 ( \32243 , \31276 );
buf \U$26613 ( \32244 , \31276 );
buf \U$26614 ( \32245 , \31276 );
buf \U$26615 ( \32246 , \31276 );
buf \U$26616 ( \32247 , \31276 );
buf \U$26617 ( \32248 , \31276 );
buf \U$26618 ( \32249 , \31276 );
buf \U$26619 ( \32250 , \31276 );
buf \U$26620 ( \32251 , \31276 );
buf \U$26621 ( \32252 , \31276 );
buf \U$26622 ( \32253 , \31276 );
buf \U$26623 ( \32254 , \31276 );
buf \U$26624 ( \32255 , \31276 );
buf \U$26625 ( \32256 , \31276 );
buf \U$26626 ( \32257 , \31263 );
or \U$26627 ( \32258 , \32227 , \32228 , \32229 , \32230 , \32231 , \32232 , \32233 , \32234 , \32235 , \32236 , \32237 , \32238 , \32239 , \32240 , \32241 , \32242 , \32243 , \32244 , \32245 , \32246 , \32247 , \32248 , \32249 , \32250 , \32251 , \32252 , \32253 , \32254 , \32255 , \32256 , \32257 );
nand \U$26628 ( \32259 , \32226 , \32258 );
buf \U$26629 ( \32260 , \32259 );
buf \U$26630 ( \32261 , \31276 );
not \U$26631 ( \32262 , \32261 );
buf \U$26632 ( \32263 , \31273 );
buf \U$26633 ( \32264 , \31276 );
buf \U$26634 ( \32265 , \31276 );
buf \U$26635 ( \32266 , \31276 );
buf \U$26636 ( \32267 , \31276 );
buf \U$26637 ( \32268 , \31276 );
buf \U$26638 ( \32269 , \31276 );
buf \U$26639 ( \32270 , \31276 );
buf \U$26640 ( \32271 , \31276 );
buf \U$26641 ( \32272 , \31276 );
buf \U$26642 ( \32273 , \31276 );
buf \U$26643 ( \32274 , \31276 );
buf \U$26644 ( \32275 , \31276 );
buf \U$26645 ( \32276 , \31276 );
buf \U$26646 ( \32277 , \31276 );
buf \U$26647 ( \32278 , \31276 );
buf \U$26648 ( \32279 , \31276 );
buf \U$26649 ( \32280 , \31276 );
buf \U$26650 ( \32281 , \31276 );
buf \U$26651 ( \32282 , \31276 );
buf \U$26652 ( \32283 , \31276 );
buf \U$26653 ( \32284 , \31276 );
buf \U$26654 ( \32285 , \31276 );
buf \U$26655 ( \32286 , \31276 );
buf \U$26656 ( \32287 , \31276 );
buf \U$26657 ( \32288 , \31276 );
buf \U$26658 ( \32289 , \31269 );
buf \U$26659 ( \32290 , \31263 );
buf \U$26660 ( \32291 , \31264 );
buf \U$26661 ( \32292 , \31265 );
buf \U$26662 ( \32293 , \31266 );
or \U$26663 ( \32294 , \32290 , \32291 , \32292 , \32293 );
and \U$26664 ( \32295 , \32289 , \32294 );
or \U$26665 ( \32296 , \32263 , \32264 , \32265 , \32266 , \32267 , \32268 , \32269 , \32270 , \32271 , \32272 , \32273 , \32274 , \32275 , \32276 , \32277 , \32278 , \32279 , \32280 , \32281 , \32282 , \32283 , \32284 , \32285 , \32286 , \32287 , \32288 , \32295 );
and \U$26666 ( \32297 , \32262 , \32296 );
buf \U$26667 ( \32298 , \32297 );
or \U$26668 ( \32299 , \32260 , \32298 );
_DC g953f ( \32300_nG953f , \32224 , \32299 );
buf \U$26669 ( \32301 , \32300_nG953f );
xor \U$26670 ( \32302 , \31791 , \32301 );
buf \U$26671 ( \32303 , RIb7b9590_247);
and \U$26672 ( \32304 , \7126 , \31817 );
and \U$26673 ( \32305 , \7128 , \31844 );
and \U$26674 ( \32306 , \8338 , \31871 );
and \U$26675 ( \32307 , \8340 , \31898 );
and \U$26676 ( \32308 , \8342 , \31925 );
and \U$26677 ( \32309 , \8344 , \31952 );
and \U$26678 ( \32310 , \8346 , \31979 );
and \U$26679 ( \32311 , \8348 , \32006 );
and \U$26680 ( \32312 , \8350 , \32033 );
and \U$26681 ( \32313 , \8352 , \32060 );
and \U$26682 ( \32314 , \8354 , \32087 );
and \U$26683 ( \32315 , \8356 , \32114 );
and \U$26684 ( \32316 , \8358 , \32141 );
and \U$26685 ( \32317 , \8360 , \32168 );
and \U$26686 ( \32318 , \8362 , \32195 );
and \U$26687 ( \32319 , \8364 , \32222 );
or \U$26688 ( \32320 , \32304 , \32305 , \32306 , \32307 , \32308 , \32309 , \32310 , \32311 , \32312 , \32313 , \32314 , \32315 , \32316 , \32317 , \32318 , \32319 );
_DC g9554 ( \32321_nG9554 , \32320 , \32299 );
buf \U$26689 ( \32322 , \32321_nG9554 );
xor \U$26690 ( \32323 , \32303 , \32322 );
or \U$26691 ( \32324 , \32302 , \32323 );
buf \U$26692 ( \32325 , RIb7b9518_248);
and \U$26693 ( \32326 , \7136 , \31817 );
and \U$26694 ( \32327 , \7138 , \31844 );
and \U$26695 ( \32328 , \8374 , \31871 );
and \U$26696 ( \32329 , \8376 , \31898 );
and \U$26697 ( \32330 , \8378 , \31925 );
and \U$26698 ( \32331 , \8380 , \31952 );
and \U$26699 ( \32332 , \8382 , \31979 );
and \U$26700 ( \32333 , \8384 , \32006 );
and \U$26701 ( \32334 , \8386 , \32033 );
and \U$26702 ( \32335 , \8388 , \32060 );
and \U$26703 ( \32336 , \8390 , \32087 );
and \U$26704 ( \32337 , \8392 , \32114 );
and \U$26705 ( \32338 , \8394 , \32141 );
and \U$26706 ( \32339 , \8396 , \32168 );
and \U$26707 ( \32340 , \8398 , \32195 );
and \U$26708 ( \32341 , \8400 , \32222 );
or \U$26709 ( \32342 , \32326 , \32327 , \32328 , \32329 , \32330 , \32331 , \32332 , \32333 , \32334 , \32335 , \32336 , \32337 , \32338 , \32339 , \32340 , \32341 );
_DC g956a ( \32343_nG956a , \32342 , \32299 );
buf \U$26710 ( \32344 , \32343_nG956a );
xor \U$26711 ( \32345 , \32325 , \32344 );
or \U$26712 ( \32346 , \32324 , \32345 );
buf \U$26713 ( \32347 , RIb7b94a0_249);
and \U$26714 ( \32348 , \7146 , \31817 );
and \U$26715 ( \32349 , \7148 , \31844 );
and \U$26716 ( \32350 , \8410 , \31871 );
and \U$26717 ( \32351 , \8412 , \31898 );
and \U$26718 ( \32352 , \8414 , \31925 );
and \U$26719 ( \32353 , \8416 , \31952 );
and \U$26720 ( \32354 , \8418 , \31979 );
and \U$26721 ( \32355 , \8420 , \32006 );
and \U$26722 ( \32356 , \8422 , \32033 );
and \U$26723 ( \32357 , \8424 , \32060 );
and \U$26724 ( \32358 , \8426 , \32087 );
and \U$26725 ( \32359 , \8428 , \32114 );
and \U$26726 ( \32360 , \8430 , \32141 );
and \U$26727 ( \32361 , \8432 , \32168 );
and \U$26728 ( \32362 , \8434 , \32195 );
and \U$26729 ( \32363 , \8436 , \32222 );
or \U$26730 ( \32364 , \32348 , \32349 , \32350 , \32351 , \32352 , \32353 , \32354 , \32355 , \32356 , \32357 , \32358 , \32359 , \32360 , \32361 , \32362 , \32363 );
_DC g9580 ( \32365_nG9580 , \32364 , \32299 );
buf \U$26731 ( \32366 , \32365_nG9580 );
xor \U$26732 ( \32367 , \32347 , \32366 );
or \U$26733 ( \32368 , \32346 , \32367 );
buf \U$26734 ( \32369 , RIb7b9428_250);
and \U$26735 ( \32370 , \7156 , \31817 );
and \U$26736 ( \32371 , \7158 , \31844 );
and \U$26737 ( \32372 , \8446 , \31871 );
and \U$26738 ( \32373 , \8448 , \31898 );
and \U$26739 ( \32374 , \8450 , \31925 );
and \U$26740 ( \32375 , \8452 , \31952 );
and \U$26741 ( \32376 , \8454 , \31979 );
and \U$26742 ( \32377 , \8456 , \32006 );
and \U$26743 ( \32378 , \8458 , \32033 );
and \U$26744 ( \32379 , \8460 , \32060 );
and \U$26745 ( \32380 , \8462 , \32087 );
and \U$26746 ( \32381 , \8464 , \32114 );
and \U$26747 ( \32382 , \8466 , \32141 );
and \U$26748 ( \32383 , \8468 , \32168 );
and \U$26749 ( \32384 , \8470 , \32195 );
and \U$26750 ( \32385 , \8472 , \32222 );
or \U$26751 ( \32386 , \32370 , \32371 , \32372 , \32373 , \32374 , \32375 , \32376 , \32377 , \32378 , \32379 , \32380 , \32381 , \32382 , \32383 , \32384 , \32385 );
_DC g9596 ( \32387_nG9596 , \32386 , \32299 );
buf \U$26752 ( \32388 , \32387_nG9596 );
xor \U$26753 ( \32389 , \32369 , \32388 );
or \U$26754 ( \32390 , \32368 , \32389 );
buf \U$26755 ( \32391 , RIb7b93b0_251);
and \U$26756 ( \32392 , \7166 , \31817 );
and \U$26757 ( \32393 , \7168 , \31844 );
and \U$26758 ( \32394 , \8482 , \31871 );
and \U$26759 ( \32395 , \8484 , \31898 );
and \U$26760 ( \32396 , \8486 , \31925 );
and \U$26761 ( \32397 , \8488 , \31952 );
and \U$26762 ( \32398 , \8490 , \31979 );
and \U$26763 ( \32399 , \8492 , \32006 );
and \U$26764 ( \32400 , \8494 , \32033 );
and \U$26765 ( \32401 , \8496 , \32060 );
and \U$26766 ( \32402 , \8498 , \32087 );
and \U$26767 ( \32403 , \8500 , \32114 );
and \U$26768 ( \32404 , \8502 , \32141 );
and \U$26769 ( \32405 , \8504 , \32168 );
and \U$26770 ( \32406 , \8506 , \32195 );
and \U$26771 ( \32407 , \8508 , \32222 );
or \U$26772 ( \32408 , \32392 , \32393 , \32394 , \32395 , \32396 , \32397 , \32398 , \32399 , \32400 , \32401 , \32402 , \32403 , \32404 , \32405 , \32406 , \32407 );
_DC g95ac ( \32409_nG95ac , \32408 , \32299 );
buf \U$26773 ( \32410 , \32409_nG95ac );
xor \U$26774 ( \32411 , \32391 , \32410 );
or \U$26775 ( \32412 , \32390 , \32411 );
buf \U$26776 ( \32413 , RIb7af720_252);
and \U$26777 ( \32414 , \7176 , \31817 );
and \U$26778 ( \32415 , \7178 , \31844 );
and \U$26779 ( \32416 , \8518 , \31871 );
and \U$26780 ( \32417 , \8520 , \31898 );
and \U$26781 ( \32418 , \8522 , \31925 );
and \U$26782 ( \32419 , \8524 , \31952 );
and \U$26783 ( \32420 , \8526 , \31979 );
and \U$26784 ( \32421 , \8528 , \32006 );
and \U$26785 ( \32422 , \8530 , \32033 );
and \U$26786 ( \32423 , \8532 , \32060 );
and \U$26787 ( \32424 , \8534 , \32087 );
and \U$26788 ( \32425 , \8536 , \32114 );
and \U$26789 ( \32426 , \8538 , \32141 );
and \U$26790 ( \32427 , \8540 , \32168 );
and \U$26791 ( \32428 , \8542 , \32195 );
and \U$26792 ( \32429 , \8544 , \32222 );
or \U$26793 ( \32430 , \32414 , \32415 , \32416 , \32417 , \32418 , \32419 , \32420 , \32421 , \32422 , \32423 , \32424 , \32425 , \32426 , \32427 , \32428 , \32429 );
_DC g95c2 ( \32431_nG95c2 , \32430 , \32299 );
buf \U$26794 ( \32432 , \32431_nG95c2 );
xor \U$26795 ( \32433 , \32413 , \32432 );
or \U$26796 ( \32434 , \32412 , \32433 );
buf \U$26797 ( \32435 , RIb7af6a8_253);
and \U$26798 ( \32436 , \7186 , \31817 );
and \U$26799 ( \32437 , \7188 , \31844 );
and \U$26800 ( \32438 , \8554 , \31871 );
and \U$26801 ( \32439 , \8556 , \31898 );
and \U$26802 ( \32440 , \8558 , \31925 );
and \U$26803 ( \32441 , \8560 , \31952 );
and \U$26804 ( \32442 , \8562 , \31979 );
and \U$26805 ( \32443 , \8564 , \32006 );
and \U$26806 ( \32444 , \8566 , \32033 );
and \U$26807 ( \32445 , \8568 , \32060 );
and \U$26808 ( \32446 , \8570 , \32087 );
and \U$26809 ( \32447 , \8572 , \32114 );
and \U$26810 ( \32448 , \8574 , \32141 );
and \U$26811 ( \32449 , \8576 , \32168 );
and \U$26812 ( \32450 , \8578 , \32195 );
and \U$26813 ( \32451 , \8580 , \32222 );
or \U$26814 ( \32452 , \32436 , \32437 , \32438 , \32439 , \32440 , \32441 , \32442 , \32443 , \32444 , \32445 , \32446 , \32447 , \32448 , \32449 , \32450 , \32451 );
_DC g95d8 ( \32453_nG95d8 , \32452 , \32299 );
buf \U$26815 ( \32454 , \32453_nG95d8 );
xor \U$26816 ( \32455 , \32435 , \32454 );
or \U$26817 ( \32456 , \32434 , \32455 );
not \U$26818 ( \32457 , \32456 );
buf \U$26819 ( \32458 , \32457 );
and \U$26820 ( \32459 , \31790 , \32458 );
buf \U$26821 ( \32460 , RIb7af630_254);
buf \U$26822 ( \32461 , \31276 );
buf \U$26823 ( \32462 , \31276 );
buf \U$26824 ( \32463 , \31276 );
buf \U$26825 ( \32464 , \31276 );
buf \U$26826 ( \32465 , \31276 );
buf \U$26827 ( \32466 , \31276 );
buf \U$26828 ( \32467 , \31276 );
buf \U$26829 ( \32468 , \31276 );
buf \U$26830 ( \32469 , \31276 );
buf \U$26831 ( \32470 , \31276 );
buf \U$26832 ( \32471 , \31276 );
buf \U$26833 ( \32472 , \31276 );
buf \U$26834 ( \32473 , \31276 );
buf \U$26835 ( \32474 , \31276 );
buf \U$26836 ( \32475 , \31276 );
buf \U$26837 ( \32476 , \31276 );
buf \U$26838 ( \32477 , \31276 );
buf \U$26839 ( \32478 , \31276 );
buf \U$26840 ( \32479 , \31276 );
buf \U$26841 ( \32480 , \31276 );
buf \U$26842 ( \32481 , \31276 );
buf \U$26843 ( \32482 , \31276 );
buf \U$26844 ( \32483 , \31276 );
buf \U$26845 ( \32484 , \31276 );
buf \U$26846 ( \32485 , \31276 );
nor \U$26847 ( \32486 , \31263 , \31264 , \31265 , \31266 , \31270 , \31273 , \31276 , \32461 , \32462 , \32463 , \32464 , \32465 , \32466 , \32467 , \32468 , \32469 , \32470 , \32471 , \32472 , \32473 , \32474 , \32475 , \32476 , \32477 , \32478 , \32479 , \32480 , \32481 , \32482 , \32483 , \32484 , \32485 );
and \U$26848 ( \32487 , \7198 , \32486 );
buf \U$26849 ( \32488 , \31276 );
buf \U$26850 ( \32489 , \31276 );
buf \U$26851 ( \32490 , \31276 );
buf \U$26852 ( \32491 , \31276 );
buf \U$26853 ( \32492 , \31276 );
buf \U$26854 ( \32493 , \31276 );
buf \U$26855 ( \32494 , \31276 );
buf \U$26856 ( \32495 , \31276 );
buf \U$26857 ( \32496 , \31276 );
buf \U$26858 ( \32497 , \31276 );
buf \U$26859 ( \32498 , \31276 );
buf \U$26860 ( \32499 , \31276 );
buf \U$26861 ( \32500 , \31276 );
buf \U$26862 ( \32501 , \31276 );
buf \U$26863 ( \32502 , \31276 );
buf \U$26864 ( \32503 , \31276 );
buf \U$26865 ( \32504 , \31276 );
buf \U$26866 ( \32505 , \31276 );
buf \U$26867 ( \32506 , \31276 );
buf \U$26868 ( \32507 , \31276 );
buf \U$26869 ( \32508 , \31276 );
buf \U$26870 ( \32509 , \31276 );
buf \U$26871 ( \32510 , \31276 );
buf \U$26872 ( \32511 , \31276 );
buf \U$26873 ( \32512 , \31276 );
nor \U$26874 ( \32513 , \31304 , \31305 , \31306 , \31307 , \31269 , \31273 , \31276 , \32488 , \32489 , \32490 , \32491 , \32492 , \32493 , \32494 , \32495 , \32496 , \32497 , \32498 , \32499 , \32500 , \32501 , \32502 , \32503 , \32504 , \32505 , \32506 , \32507 , \32508 , \32509 , \32510 , \32511 , \32512 );
and \U$26875 ( \32514 , \7200 , \32513 );
buf \U$26876 ( \32515 , \31276 );
buf \U$26877 ( \32516 , \31276 );
buf \U$26878 ( \32517 , \31276 );
buf \U$26879 ( \32518 , \31276 );
buf \U$26880 ( \32519 , \31276 );
buf \U$26881 ( \32520 , \31276 );
buf \U$26882 ( \32521 , \31276 );
buf \U$26883 ( \32522 , \31276 );
buf \U$26884 ( \32523 , \31276 );
buf \U$26885 ( \32524 , \31276 );
buf \U$26886 ( \32525 , \31276 );
buf \U$26887 ( \32526 , \31276 );
buf \U$26888 ( \32527 , \31276 );
buf \U$26889 ( \32528 , \31276 );
buf \U$26890 ( \32529 , \31276 );
buf \U$26891 ( \32530 , \31276 );
buf \U$26892 ( \32531 , \31276 );
buf \U$26893 ( \32532 , \31276 );
buf \U$26894 ( \32533 , \31276 );
buf \U$26895 ( \32534 , \31276 );
buf \U$26896 ( \32535 , \31276 );
buf \U$26897 ( \32536 , \31276 );
buf \U$26898 ( \32537 , \31276 );
buf \U$26899 ( \32538 , \31276 );
buf \U$26900 ( \32539 , \31276 );
nor \U$26901 ( \32540 , \31263 , \31305 , \31306 , \31307 , \31269 , \31273 , \31276 , \32515 , \32516 , \32517 , \32518 , \32519 , \32520 , \32521 , \32522 , \32523 , \32524 , \32525 , \32526 , \32527 , \32528 , \32529 , \32530 , \32531 , \32532 , \32533 , \32534 , \32535 , \32536 , \32537 , \32538 , \32539 );
and \U$26902 ( \32541 , \8645 , \32540 );
buf \U$26903 ( \32542 , \31276 );
buf \U$26904 ( \32543 , \31276 );
buf \U$26905 ( \32544 , \31276 );
buf \U$26906 ( \32545 , \31276 );
buf \U$26907 ( \32546 , \31276 );
buf \U$26908 ( \32547 , \31276 );
buf \U$26909 ( \32548 , \31276 );
buf \U$26910 ( \32549 , \31276 );
buf \U$26911 ( \32550 , \31276 );
buf \U$26912 ( \32551 , \31276 );
buf \U$26913 ( \32552 , \31276 );
buf \U$26914 ( \32553 , \31276 );
buf \U$26915 ( \32554 , \31276 );
buf \U$26916 ( \32555 , \31276 );
buf \U$26917 ( \32556 , \31276 );
buf \U$26918 ( \32557 , \31276 );
buf \U$26919 ( \32558 , \31276 );
buf \U$26920 ( \32559 , \31276 );
buf \U$26921 ( \32560 , \31276 );
buf \U$26922 ( \32561 , \31276 );
buf \U$26923 ( \32562 , \31276 );
buf \U$26924 ( \32563 , \31276 );
buf \U$26925 ( \32564 , \31276 );
buf \U$26926 ( \32565 , \31276 );
buf \U$26927 ( \32566 , \31276 );
nor \U$26928 ( \32567 , \31304 , \31264 , \31306 , \31307 , \31269 , \31273 , \31276 , \32542 , \32543 , \32544 , \32545 , \32546 , \32547 , \32548 , \32549 , \32550 , \32551 , \32552 , \32553 , \32554 , \32555 , \32556 , \32557 , \32558 , \32559 , \32560 , \32561 , \32562 , \32563 , \32564 , \32565 , \32566 );
and \U$26929 ( \32568 , \8673 , \32567 );
buf \U$26930 ( \32569 , \31276 );
buf \U$26931 ( \32570 , \31276 );
buf \U$26932 ( \32571 , \31276 );
buf \U$26933 ( \32572 , \31276 );
buf \U$26934 ( \32573 , \31276 );
buf \U$26935 ( \32574 , \31276 );
buf \U$26936 ( \32575 , \31276 );
buf \U$26937 ( \32576 , \31276 );
buf \U$26938 ( \32577 , \31276 );
buf \U$26939 ( \32578 , \31276 );
buf \U$26940 ( \32579 , \31276 );
buf \U$26941 ( \32580 , \31276 );
buf \U$26942 ( \32581 , \31276 );
buf \U$26943 ( \32582 , \31276 );
buf \U$26944 ( \32583 , \31276 );
buf \U$26945 ( \32584 , \31276 );
buf \U$26946 ( \32585 , \31276 );
buf \U$26947 ( \32586 , \31276 );
buf \U$26948 ( \32587 , \31276 );
buf \U$26949 ( \32588 , \31276 );
buf \U$26950 ( \32589 , \31276 );
buf \U$26951 ( \32590 , \31276 );
buf \U$26952 ( \32591 , \31276 );
buf \U$26953 ( \32592 , \31276 );
buf \U$26954 ( \32593 , \31276 );
nor \U$26955 ( \32594 , \31263 , \31264 , \31306 , \31307 , \31269 , \31273 , \31276 , \32569 , \32570 , \32571 , \32572 , \32573 , \32574 , \32575 , \32576 , \32577 , \32578 , \32579 , \32580 , \32581 , \32582 , \32583 , \32584 , \32585 , \32586 , \32587 , \32588 , \32589 , \32590 , \32591 , \32592 , \32593 );
and \U$26956 ( \32595 , \8701 , \32594 );
buf \U$26957 ( \32596 , \31276 );
buf \U$26958 ( \32597 , \31276 );
buf \U$26959 ( \32598 , \31276 );
buf \U$26960 ( \32599 , \31276 );
buf \U$26961 ( \32600 , \31276 );
buf \U$26962 ( \32601 , \31276 );
buf \U$26963 ( \32602 , \31276 );
buf \U$26964 ( \32603 , \31276 );
buf \U$26965 ( \32604 , \31276 );
buf \U$26966 ( \32605 , \31276 );
buf \U$26967 ( \32606 , \31276 );
buf \U$26968 ( \32607 , \31276 );
buf \U$26969 ( \32608 , \31276 );
buf \U$26970 ( \32609 , \31276 );
buf \U$26971 ( \32610 , \31276 );
buf \U$26972 ( \32611 , \31276 );
buf \U$26973 ( \32612 , \31276 );
buf \U$26974 ( \32613 , \31276 );
buf \U$26975 ( \32614 , \31276 );
buf \U$26976 ( \32615 , \31276 );
buf \U$26977 ( \32616 , \31276 );
buf \U$26978 ( \32617 , \31276 );
buf \U$26979 ( \32618 , \31276 );
buf \U$26980 ( \32619 , \31276 );
buf \U$26981 ( \32620 , \31276 );
nor \U$26982 ( \32621 , \31304 , \31305 , \31265 , \31307 , \31269 , \31273 , \31276 , \32596 , \32597 , \32598 , \32599 , \32600 , \32601 , \32602 , \32603 , \32604 , \32605 , \32606 , \32607 , \32608 , \32609 , \32610 , \32611 , \32612 , \32613 , \32614 , \32615 , \32616 , \32617 , \32618 , \32619 , \32620 );
and \U$26983 ( \32622 , \8729 , \32621 );
buf \U$26984 ( \32623 , \31276 );
buf \U$26985 ( \32624 , \31276 );
buf \U$26986 ( \32625 , \31276 );
buf \U$26987 ( \32626 , \31276 );
buf \U$26988 ( \32627 , \31276 );
buf \U$26989 ( \32628 , \31276 );
buf \U$26990 ( \32629 , \31276 );
buf \U$26991 ( \32630 , \31276 );
buf \U$26992 ( \32631 , \31276 );
buf \U$26993 ( \32632 , \31276 );
buf \U$26994 ( \32633 , \31276 );
buf \U$26995 ( \32634 , \31276 );
buf \U$26996 ( \32635 , \31276 );
buf \U$26997 ( \32636 , \31276 );
buf \U$26998 ( \32637 , \31276 );
buf \U$26999 ( \32638 , \31276 );
buf \U$27000 ( \32639 , \31276 );
buf \U$27001 ( \32640 , \31276 );
buf \U$27002 ( \32641 , \31276 );
buf \U$27003 ( \32642 , \31276 );
buf \U$27004 ( \32643 , \31276 );
buf \U$27005 ( \32644 , \31276 );
buf \U$27006 ( \32645 , \31276 );
buf \U$27007 ( \32646 , \31276 );
buf \U$27008 ( \32647 , \31276 );
nor \U$27009 ( \32648 , \31263 , \31305 , \31265 , \31307 , \31269 , \31273 , \31276 , \32623 , \32624 , \32625 , \32626 , \32627 , \32628 , \32629 , \32630 , \32631 , \32632 , \32633 , \32634 , \32635 , \32636 , \32637 , \32638 , \32639 , \32640 , \32641 , \32642 , \32643 , \32644 , \32645 , \32646 , \32647 );
and \U$27010 ( \32649 , \8757 , \32648 );
buf \U$27011 ( \32650 , \31276 );
buf \U$27012 ( \32651 , \31276 );
buf \U$27013 ( \32652 , \31276 );
buf \U$27014 ( \32653 , \31276 );
buf \U$27015 ( \32654 , \31276 );
buf \U$27016 ( \32655 , \31276 );
buf \U$27017 ( \32656 , \31276 );
buf \U$27018 ( \32657 , \31276 );
buf \U$27019 ( \32658 , \31276 );
buf \U$27020 ( \32659 , \31276 );
buf \U$27021 ( \32660 , \31276 );
buf \U$27022 ( \32661 , \31276 );
buf \U$27023 ( \32662 , \31276 );
buf \U$27024 ( \32663 , \31276 );
buf \U$27025 ( \32664 , \31276 );
buf \U$27026 ( \32665 , \31276 );
buf \U$27027 ( \32666 , \31276 );
buf \U$27028 ( \32667 , \31276 );
buf \U$27029 ( \32668 , \31276 );
buf \U$27030 ( \32669 , \31276 );
buf \U$27031 ( \32670 , \31276 );
buf \U$27032 ( \32671 , \31276 );
buf \U$27033 ( \32672 , \31276 );
buf \U$27034 ( \32673 , \31276 );
buf \U$27035 ( \32674 , \31276 );
nor \U$27036 ( \32675 , \31304 , \31264 , \31265 , \31307 , \31269 , \31273 , \31276 , \32650 , \32651 , \32652 , \32653 , \32654 , \32655 , \32656 , \32657 , \32658 , \32659 , \32660 , \32661 , \32662 , \32663 , \32664 , \32665 , \32666 , \32667 , \32668 , \32669 , \32670 , \32671 , \32672 , \32673 , \32674 );
and \U$27037 ( \32676 , \8785 , \32675 );
buf \U$27038 ( \32677 , \31276 );
buf \U$27039 ( \32678 , \31276 );
buf \U$27040 ( \32679 , \31276 );
buf \U$27041 ( \32680 , \31276 );
buf \U$27042 ( \32681 , \31276 );
buf \U$27043 ( \32682 , \31276 );
buf \U$27044 ( \32683 , \31276 );
buf \U$27045 ( \32684 , \31276 );
buf \U$27046 ( \32685 , \31276 );
buf \U$27047 ( \32686 , \31276 );
buf \U$27048 ( \32687 , \31276 );
buf \U$27049 ( \32688 , \31276 );
buf \U$27050 ( \32689 , \31276 );
buf \U$27051 ( \32690 , \31276 );
buf \U$27052 ( \32691 , \31276 );
buf \U$27053 ( \32692 , \31276 );
buf \U$27054 ( \32693 , \31276 );
buf \U$27055 ( \32694 , \31276 );
buf \U$27056 ( \32695 , \31276 );
buf \U$27057 ( \32696 , \31276 );
buf \U$27058 ( \32697 , \31276 );
buf \U$27059 ( \32698 , \31276 );
buf \U$27060 ( \32699 , \31276 );
buf \U$27061 ( \32700 , \31276 );
buf \U$27062 ( \32701 , \31276 );
nor \U$27063 ( \32702 , \31263 , \31264 , \31265 , \31307 , \31269 , \31273 , \31276 , \32677 , \32678 , \32679 , \32680 , \32681 , \32682 , \32683 , \32684 , \32685 , \32686 , \32687 , \32688 , \32689 , \32690 , \32691 , \32692 , \32693 , \32694 , \32695 , \32696 , \32697 , \32698 , \32699 , \32700 , \32701 );
and \U$27064 ( \32703 , \8813 , \32702 );
buf \U$27065 ( \32704 , \31276 );
buf \U$27066 ( \32705 , \31276 );
buf \U$27067 ( \32706 , \31276 );
buf \U$27068 ( \32707 , \31276 );
buf \U$27069 ( \32708 , \31276 );
buf \U$27070 ( \32709 , \31276 );
buf \U$27071 ( \32710 , \31276 );
buf \U$27072 ( \32711 , \31276 );
buf \U$27073 ( \32712 , \31276 );
buf \U$27074 ( \32713 , \31276 );
buf \U$27075 ( \32714 , \31276 );
buf \U$27076 ( \32715 , \31276 );
buf \U$27077 ( \32716 , \31276 );
buf \U$27078 ( \32717 , \31276 );
buf \U$27079 ( \32718 , \31276 );
buf \U$27080 ( \32719 , \31276 );
buf \U$27081 ( \32720 , \31276 );
buf \U$27082 ( \32721 , \31276 );
buf \U$27083 ( \32722 , \31276 );
buf \U$27084 ( \32723 , \31276 );
buf \U$27085 ( \32724 , \31276 );
buf \U$27086 ( \32725 , \31276 );
buf \U$27087 ( \32726 , \31276 );
buf \U$27088 ( \32727 , \31276 );
buf \U$27089 ( \32728 , \31276 );
nor \U$27090 ( \32729 , \31304 , \31305 , \31306 , \31266 , \31269 , \31273 , \31276 , \32704 , \32705 , \32706 , \32707 , \32708 , \32709 , \32710 , \32711 , \32712 , \32713 , \32714 , \32715 , \32716 , \32717 , \32718 , \32719 , \32720 , \32721 , \32722 , \32723 , \32724 , \32725 , \32726 , \32727 , \32728 );
and \U$27091 ( \32730 , \8841 , \32729 );
buf \U$27092 ( \32731 , \31276 );
buf \U$27093 ( \32732 , \31276 );
buf \U$27094 ( \32733 , \31276 );
buf \U$27095 ( \32734 , \31276 );
buf \U$27096 ( \32735 , \31276 );
buf \U$27097 ( \32736 , \31276 );
buf \U$27098 ( \32737 , \31276 );
buf \U$27099 ( \32738 , \31276 );
buf \U$27100 ( \32739 , \31276 );
buf \U$27101 ( \32740 , \31276 );
buf \U$27102 ( \32741 , \31276 );
buf \U$27103 ( \32742 , \31276 );
buf \U$27104 ( \32743 , \31276 );
buf \U$27105 ( \32744 , \31276 );
buf \U$27106 ( \32745 , \31276 );
buf \U$27107 ( \32746 , \31276 );
buf \U$27108 ( \32747 , \31276 );
buf \U$27109 ( \32748 , \31276 );
buf \U$27110 ( \32749 , \31276 );
buf \U$27111 ( \32750 , \31276 );
buf \U$27112 ( \32751 , \31276 );
buf \U$27113 ( \32752 , \31276 );
buf \U$27114 ( \32753 , \31276 );
buf \U$27115 ( \32754 , \31276 );
buf \U$27116 ( \32755 , \31276 );
nor \U$27117 ( \32756 , \31263 , \31305 , \31306 , \31266 , \31269 , \31273 , \31276 , \32731 , \32732 , \32733 , \32734 , \32735 , \32736 , \32737 , \32738 , \32739 , \32740 , \32741 , \32742 , \32743 , \32744 , \32745 , \32746 , \32747 , \32748 , \32749 , \32750 , \32751 , \32752 , \32753 , \32754 , \32755 );
and \U$27118 ( \32757 , \8869 , \32756 );
buf \U$27119 ( \32758 , \31276 );
buf \U$27120 ( \32759 , \31276 );
buf \U$27121 ( \32760 , \31276 );
buf \U$27122 ( \32761 , \31276 );
buf \U$27123 ( \32762 , \31276 );
buf \U$27124 ( \32763 , \31276 );
buf \U$27125 ( \32764 , \31276 );
buf \U$27126 ( \32765 , \31276 );
buf \U$27127 ( \32766 , \31276 );
buf \U$27128 ( \32767 , \31276 );
buf \U$27129 ( \32768 , \31276 );
buf \U$27130 ( \32769 , \31276 );
buf \U$27131 ( \32770 , \31276 );
buf \U$27132 ( \32771 , \31276 );
buf \U$27133 ( \32772 , \31276 );
buf \U$27134 ( \32773 , \31276 );
buf \U$27135 ( \32774 , \31276 );
buf \U$27136 ( \32775 , \31276 );
buf \U$27137 ( \32776 , \31276 );
buf \U$27138 ( \32777 , \31276 );
buf \U$27139 ( \32778 , \31276 );
buf \U$27140 ( \32779 , \31276 );
buf \U$27141 ( \32780 , \31276 );
buf \U$27142 ( \32781 , \31276 );
buf \U$27143 ( \32782 , \31276 );
nor \U$27144 ( \32783 , \31304 , \31264 , \31306 , \31266 , \31269 , \31273 , \31276 , \32758 , \32759 , \32760 , \32761 , \32762 , \32763 , \32764 , \32765 , \32766 , \32767 , \32768 , \32769 , \32770 , \32771 , \32772 , \32773 , \32774 , \32775 , \32776 , \32777 , \32778 , \32779 , \32780 , \32781 , \32782 );
and \U$27145 ( \32784 , \8897 , \32783 );
buf \U$27146 ( \32785 , \31276 );
buf \U$27147 ( \32786 , \31276 );
buf \U$27148 ( \32787 , \31276 );
buf \U$27149 ( \32788 , \31276 );
buf \U$27150 ( \32789 , \31276 );
buf \U$27151 ( \32790 , \31276 );
buf \U$27152 ( \32791 , \31276 );
buf \U$27153 ( \32792 , \31276 );
buf \U$27154 ( \32793 , \31276 );
buf \U$27155 ( \32794 , \31276 );
buf \U$27156 ( \32795 , \31276 );
buf \U$27157 ( \32796 , \31276 );
buf \U$27158 ( \32797 , \31276 );
buf \U$27159 ( \32798 , \31276 );
buf \U$27160 ( \32799 , \31276 );
buf \U$27161 ( \32800 , \31276 );
buf \U$27162 ( \32801 , \31276 );
buf \U$27163 ( \32802 , \31276 );
buf \U$27164 ( \32803 , \31276 );
buf \U$27165 ( \32804 , \31276 );
buf \U$27166 ( \32805 , \31276 );
buf \U$27167 ( \32806 , \31276 );
buf \U$27168 ( \32807 , \31276 );
buf \U$27169 ( \32808 , \31276 );
buf \U$27170 ( \32809 , \31276 );
nor \U$27171 ( \32810 , \31263 , \31264 , \31306 , \31266 , \31269 , \31273 , \31276 , \32785 , \32786 , \32787 , \32788 , \32789 , \32790 , \32791 , \32792 , \32793 , \32794 , \32795 , \32796 , \32797 , \32798 , \32799 , \32800 , \32801 , \32802 , \32803 , \32804 , \32805 , \32806 , \32807 , \32808 , \32809 );
and \U$27172 ( \32811 , \8925 , \32810 );
buf \U$27173 ( \32812 , \31276 );
buf \U$27174 ( \32813 , \31276 );
buf \U$27175 ( \32814 , \31276 );
buf \U$27176 ( \32815 , \31276 );
buf \U$27177 ( \32816 , \31276 );
buf \U$27178 ( \32817 , \31276 );
buf \U$27179 ( \32818 , \31276 );
buf \U$27180 ( \32819 , \31276 );
buf \U$27181 ( \32820 , \31276 );
buf \U$27182 ( \32821 , \31276 );
buf \U$27183 ( \32822 , \31276 );
buf \U$27184 ( \32823 , \31276 );
buf \U$27185 ( \32824 , \31276 );
buf \U$27186 ( \32825 , \31276 );
buf \U$27187 ( \32826 , \31276 );
buf \U$27188 ( \32827 , \31276 );
buf \U$27189 ( \32828 , \31276 );
buf \U$27190 ( \32829 , \31276 );
buf \U$27191 ( \32830 , \31276 );
buf \U$27192 ( \32831 , \31276 );
buf \U$27193 ( \32832 , \31276 );
buf \U$27194 ( \32833 , \31276 );
buf \U$27195 ( \32834 , \31276 );
buf \U$27196 ( \32835 , \31276 );
buf \U$27197 ( \32836 , \31276 );
nor \U$27198 ( \32837 , \31304 , \31305 , \31265 , \31266 , \31269 , \31273 , \31276 , \32812 , \32813 , \32814 , \32815 , \32816 , \32817 , \32818 , \32819 , \32820 , \32821 , \32822 , \32823 , \32824 , \32825 , \32826 , \32827 , \32828 , \32829 , \32830 , \32831 , \32832 , \32833 , \32834 , \32835 , \32836 );
and \U$27199 ( \32838 , \8953 , \32837 );
buf \U$27200 ( \32839 , \31276 );
buf \U$27201 ( \32840 , \31276 );
buf \U$27202 ( \32841 , \31276 );
buf \U$27203 ( \32842 , \31276 );
buf \U$27204 ( \32843 , \31276 );
buf \U$27205 ( \32844 , \31276 );
buf \U$27206 ( \32845 , \31276 );
buf \U$27207 ( \32846 , \31276 );
buf \U$27208 ( \32847 , \31276 );
buf \U$27209 ( \32848 , \31276 );
buf \U$27210 ( \32849 , \31276 );
buf \U$27211 ( \32850 , \31276 );
buf \U$27212 ( \32851 , \31276 );
buf \U$27213 ( \32852 , \31276 );
buf \U$27214 ( \32853 , \31276 );
buf \U$27215 ( \32854 , \31276 );
buf \U$27216 ( \32855 , \31276 );
buf \U$27217 ( \32856 , \31276 );
buf \U$27218 ( \32857 , \31276 );
buf \U$27219 ( \32858 , \31276 );
buf \U$27220 ( \32859 , \31276 );
buf \U$27221 ( \32860 , \31276 );
buf \U$27222 ( \32861 , \31276 );
buf \U$27223 ( \32862 , \31276 );
buf \U$27224 ( \32863 , \31276 );
nor \U$27225 ( \32864 , \31263 , \31305 , \31265 , \31266 , \31269 , \31273 , \31276 , \32839 , \32840 , \32841 , \32842 , \32843 , \32844 , \32845 , \32846 , \32847 , \32848 , \32849 , \32850 , \32851 , \32852 , \32853 , \32854 , \32855 , \32856 , \32857 , \32858 , \32859 , \32860 , \32861 , \32862 , \32863 );
and \U$27226 ( \32865 , \8981 , \32864 );
buf \U$27227 ( \32866 , \31276 );
buf \U$27228 ( \32867 , \31276 );
buf \U$27229 ( \32868 , \31276 );
buf \U$27230 ( \32869 , \31276 );
buf \U$27231 ( \32870 , \31276 );
buf \U$27232 ( \32871 , \31276 );
buf \U$27233 ( \32872 , \31276 );
buf \U$27234 ( \32873 , \31276 );
buf \U$27235 ( \32874 , \31276 );
buf \U$27236 ( \32875 , \31276 );
buf \U$27237 ( \32876 , \31276 );
buf \U$27238 ( \32877 , \31276 );
buf \U$27239 ( \32878 , \31276 );
buf \U$27240 ( \32879 , \31276 );
buf \U$27241 ( \32880 , \31276 );
buf \U$27242 ( \32881 , \31276 );
buf \U$27243 ( \32882 , \31276 );
buf \U$27244 ( \32883 , \31276 );
buf \U$27245 ( \32884 , \31276 );
buf \U$27246 ( \32885 , \31276 );
buf \U$27247 ( \32886 , \31276 );
buf \U$27248 ( \32887 , \31276 );
buf \U$27249 ( \32888 , \31276 );
buf \U$27250 ( \32889 , \31276 );
buf \U$27251 ( \32890 , \31276 );
nor \U$27252 ( \32891 , \31304 , \31264 , \31265 , \31266 , \31269 , \31273 , \31276 , \32866 , \32867 , \32868 , \32869 , \32870 , \32871 , \32872 , \32873 , \32874 , \32875 , \32876 , \32877 , \32878 , \32879 , \32880 , \32881 , \32882 , \32883 , \32884 , \32885 , \32886 , \32887 , \32888 , \32889 , \32890 );
and \U$27253 ( \32892 , \9009 , \32891 );
or \U$27254 ( \32893 , \32487 , \32514 , \32541 , \32568 , \32595 , \32622 , \32649 , \32676 , \32703 , \32730 , \32757 , \32784 , \32811 , \32838 , \32865 , \32892 );
buf \U$27255 ( \32894 , \31276 );
not \U$27256 ( \32895 , \32894 );
buf \U$27257 ( \32896 , \31264 );
buf \U$27258 ( \32897 , \31265 );
buf \U$27259 ( \32898 , \31266 );
buf \U$27260 ( \32899 , \31269 );
buf \U$27261 ( \32900 , \31273 );
buf \U$27262 ( \32901 , \31276 );
buf \U$27263 ( \32902 , \31276 );
buf \U$27264 ( \32903 , \31276 );
buf \U$27265 ( \32904 , \31276 );
buf \U$27266 ( \32905 , \31276 );
buf \U$27267 ( \32906 , \31276 );
buf \U$27268 ( \32907 , \31276 );
buf \U$27269 ( \32908 , \31276 );
buf \U$27270 ( \32909 , \31276 );
buf \U$27271 ( \32910 , \31276 );
buf \U$27272 ( \32911 , \31276 );
buf \U$27273 ( \32912 , \31276 );
buf \U$27274 ( \32913 , \31276 );
buf \U$27275 ( \32914 , \31276 );
buf \U$27276 ( \32915 , \31276 );
buf \U$27277 ( \32916 , \31276 );
buf \U$27278 ( \32917 , \31276 );
buf \U$27279 ( \32918 , \31276 );
buf \U$27280 ( \32919 , \31276 );
buf \U$27281 ( \32920 , \31276 );
buf \U$27282 ( \32921 , \31276 );
buf \U$27283 ( \32922 , \31276 );
buf \U$27284 ( \32923 , \31276 );
buf \U$27285 ( \32924 , \31276 );
buf \U$27286 ( \32925 , \31276 );
buf \U$27287 ( \32926 , \31263 );
or \U$27288 ( \32927 , \32896 , \32897 , \32898 , \32899 , \32900 , \32901 , \32902 , \32903 , \32904 , \32905 , \32906 , \32907 , \32908 , \32909 , \32910 , \32911 , \32912 , \32913 , \32914 , \32915 , \32916 , \32917 , \32918 , \32919 , \32920 , \32921 , \32922 , \32923 , \32924 , \32925 , \32926 );
nand \U$27289 ( \32928 , \32895 , \32927 );
buf \U$27290 ( \32929 , \32928 );
buf \U$27291 ( \32930 , \31276 );
not \U$27292 ( \32931 , \32930 );
buf \U$27293 ( \32932 , \31273 );
buf \U$27294 ( \32933 , \31276 );
buf \U$27295 ( \32934 , \31276 );
buf \U$27296 ( \32935 , \31276 );
buf \U$27297 ( \32936 , \31276 );
buf \U$27298 ( \32937 , \31276 );
buf \U$27299 ( \32938 , \31276 );
buf \U$27300 ( \32939 , \31276 );
buf \U$27301 ( \32940 , \31276 );
buf \U$27302 ( \32941 , \31276 );
buf \U$27303 ( \32942 , \31276 );
buf \U$27304 ( \32943 , \31276 );
buf \U$27305 ( \32944 , \31276 );
buf \U$27306 ( \32945 , \31276 );
buf \U$27307 ( \32946 , \31276 );
buf \U$27308 ( \32947 , \31276 );
buf \U$27309 ( \32948 , \31276 );
buf \U$27310 ( \32949 , \31276 );
buf \U$27311 ( \32950 , \31276 );
buf \U$27312 ( \32951 , \31276 );
buf \U$27313 ( \32952 , \31276 );
buf \U$27314 ( \32953 , \31276 );
buf \U$27315 ( \32954 , \31276 );
buf \U$27316 ( \32955 , \31276 );
buf \U$27317 ( \32956 , \31276 );
buf \U$27318 ( \32957 , \31276 );
buf \U$27319 ( \32958 , \31269 );
buf \U$27320 ( \32959 , \31263 );
buf \U$27321 ( \32960 , \31264 );
buf \U$27322 ( \32961 , \31265 );
buf \U$27323 ( \32962 , \31266 );
or \U$27324 ( \32963 , \32959 , \32960 , \32961 , \32962 );
and \U$27325 ( \32964 , \32958 , \32963 );
or \U$27326 ( \32965 , \32932 , \32933 , \32934 , \32935 , \32936 , \32937 , \32938 , \32939 , \32940 , \32941 , \32942 , \32943 , \32944 , \32945 , \32946 , \32947 , \32948 , \32949 , \32950 , \32951 , \32952 , \32953 , \32954 , \32955 , \32956 , \32957 , \32964 );
and \U$27327 ( \32966 , \32931 , \32965 );
buf \U$27328 ( \32967 , \32966 );
or \U$27329 ( \32968 , \32929 , \32967 );
_DC g97dc ( \32969_nG97dc , \32893 , \32968 );
buf \U$27330 ( \32970 , \32969_nG97dc );
xor \U$27331 ( \32971 , \32460 , \32970 );
buf \U$27332 ( \32972 , RIb7af5b8_255);
and \U$27333 ( \32973 , \7207 , \32486 );
and \U$27334 ( \32974 , \7209 , \32513 );
and \U$27335 ( \32975 , \9119 , \32540 );
and \U$27336 ( \32976 , \9121 , \32567 );
and \U$27337 ( \32977 , \9123 , \32594 );
and \U$27338 ( \32978 , \9125 , \32621 );
and \U$27339 ( \32979 , \9127 , \32648 );
and \U$27340 ( \32980 , \9129 , \32675 );
and \U$27341 ( \32981 , \9131 , \32702 );
and \U$27342 ( \32982 , \9133 , \32729 );
and \U$27343 ( \32983 , \9135 , \32756 );
and \U$27344 ( \32984 , \9137 , \32783 );
and \U$27345 ( \32985 , \9139 , \32810 );
and \U$27346 ( \32986 , \9141 , \32837 );
and \U$27347 ( \32987 , \9143 , \32864 );
and \U$27348 ( \32988 , \9145 , \32891 );
or \U$27349 ( \32989 , \32973 , \32974 , \32975 , \32976 , \32977 , \32978 , \32979 , \32980 , \32981 , \32982 , \32983 , \32984 , \32985 , \32986 , \32987 , \32988 );
_DC g97f1 ( \32990_nG97f1 , \32989 , \32968 );
buf \U$27350 ( \32991 , \32990_nG97f1 );
xor \U$27351 ( \32992 , \32972 , \32991 );
or \U$27352 ( \32993 , \32971 , \32992 );
buf \U$27353 ( \32994 , RIb7af540_256);
and \U$27354 ( \32995 , \7217 , \32486 );
and \U$27355 ( \32996 , \7219 , \32513 );
and \U$27356 ( \32997 , \9155 , \32540 );
and \U$27357 ( \32998 , \9157 , \32567 );
and \U$27358 ( \32999 , \9159 , \32594 );
and \U$27359 ( \33000 , \9161 , \32621 );
and \U$27360 ( \33001 , \9163 , \32648 );
and \U$27361 ( \33002 , \9165 , \32675 );
and \U$27362 ( \33003 , \9167 , \32702 );
and \U$27363 ( \33004 , \9169 , \32729 );
and \U$27364 ( \33005 , \9171 , \32756 );
and \U$27365 ( \33006 , \9173 , \32783 );
and \U$27366 ( \33007 , \9175 , \32810 );
and \U$27367 ( \33008 , \9177 , \32837 );
and \U$27368 ( \33009 , \9179 , \32864 );
and \U$27369 ( \33010 , \9181 , \32891 );
or \U$27370 ( \33011 , \32995 , \32996 , \32997 , \32998 , \32999 , \33000 , \33001 , \33002 , \33003 , \33004 , \33005 , \33006 , \33007 , \33008 , \33009 , \33010 );
_DC g9807 ( \33012_nG9807 , \33011 , \32968 );
buf \U$27371 ( \33013 , \33012_nG9807 );
xor \U$27372 ( \33014 , \32994 , \33013 );
or \U$27373 ( \33015 , \32993 , \33014 );
buf \U$27374 ( \33016 , RIb7af4c8_257);
and \U$27375 ( \33017 , \7227 , \32486 );
and \U$27376 ( \33018 , \7229 , \32513 );
and \U$27377 ( \33019 , \9191 , \32540 );
and \U$27378 ( \33020 , \9193 , \32567 );
and \U$27379 ( \33021 , \9195 , \32594 );
and \U$27380 ( \33022 , \9197 , \32621 );
and \U$27381 ( \33023 , \9199 , \32648 );
and \U$27382 ( \33024 , \9201 , \32675 );
and \U$27383 ( \33025 , \9203 , \32702 );
and \U$27384 ( \33026 , \9205 , \32729 );
and \U$27385 ( \33027 , \9207 , \32756 );
and \U$27386 ( \33028 , \9209 , \32783 );
and \U$27387 ( \33029 , \9211 , \32810 );
and \U$27388 ( \33030 , \9213 , \32837 );
and \U$27389 ( \33031 , \9215 , \32864 );
and \U$27390 ( \33032 , \9217 , \32891 );
or \U$27391 ( \33033 , \33017 , \33018 , \33019 , \33020 , \33021 , \33022 , \33023 , \33024 , \33025 , \33026 , \33027 , \33028 , \33029 , \33030 , \33031 , \33032 );
_DC g981d ( \33034_nG981d , \33033 , \32968 );
buf \U$27392 ( \33035 , \33034_nG981d );
xor \U$27393 ( \33036 , \33016 , \33035 );
or \U$27394 ( \33037 , \33015 , \33036 );
buf \U$27395 ( \33038 , RIb7af450_258);
and \U$27396 ( \33039 , \7237 , \32486 );
and \U$27397 ( \33040 , \7239 , \32513 );
and \U$27398 ( \33041 , \9227 , \32540 );
and \U$27399 ( \33042 , \9229 , \32567 );
and \U$27400 ( \33043 , \9231 , \32594 );
and \U$27401 ( \33044 , \9233 , \32621 );
and \U$27402 ( \33045 , \9235 , \32648 );
and \U$27403 ( \33046 , \9237 , \32675 );
and \U$27404 ( \33047 , \9239 , \32702 );
and \U$27405 ( \33048 , \9241 , \32729 );
and \U$27406 ( \33049 , \9243 , \32756 );
and \U$27407 ( \33050 , \9245 , \32783 );
and \U$27408 ( \33051 , \9247 , \32810 );
and \U$27409 ( \33052 , \9249 , \32837 );
and \U$27410 ( \33053 , \9251 , \32864 );
and \U$27411 ( \33054 , \9253 , \32891 );
or \U$27412 ( \33055 , \33039 , \33040 , \33041 , \33042 , \33043 , \33044 , \33045 , \33046 , \33047 , \33048 , \33049 , \33050 , \33051 , \33052 , \33053 , \33054 );
_DC g9833 ( \33056_nG9833 , \33055 , \32968 );
buf \U$27413 ( \33057 , \33056_nG9833 );
xor \U$27414 ( \33058 , \33038 , \33057 );
or \U$27415 ( \33059 , \33037 , \33058 );
buf \U$27416 ( \33060 , RIb7af3d8_259);
and \U$27417 ( \33061 , \7247 , \32486 );
and \U$27418 ( \33062 , \7249 , \32513 );
and \U$27419 ( \33063 , \9263 , \32540 );
and \U$27420 ( \33064 , \9265 , \32567 );
and \U$27421 ( \33065 , \9267 , \32594 );
and \U$27422 ( \33066 , \9269 , \32621 );
and \U$27423 ( \33067 , \9271 , \32648 );
and \U$27424 ( \33068 , \9273 , \32675 );
and \U$27425 ( \33069 , \9275 , \32702 );
and \U$27426 ( \33070 , \9277 , \32729 );
and \U$27427 ( \33071 , \9279 , \32756 );
and \U$27428 ( \33072 , \9281 , \32783 );
and \U$27429 ( \33073 , \9283 , \32810 );
and \U$27430 ( \33074 , \9285 , \32837 );
and \U$27431 ( \33075 , \9287 , \32864 );
and \U$27432 ( \33076 , \9289 , \32891 );
or \U$27433 ( \33077 , \33061 , \33062 , \33063 , \33064 , \33065 , \33066 , \33067 , \33068 , \33069 , \33070 , \33071 , \33072 , \33073 , \33074 , \33075 , \33076 );
_DC g9849 ( \33078_nG9849 , \33077 , \32968 );
buf \U$27434 ( \33079 , \33078_nG9849 );
xor \U$27435 ( \33080 , \33060 , \33079 );
or \U$27436 ( \33081 , \33059 , \33080 );
buf \U$27437 ( \33082 , RIb7a5bf8_260);
and \U$27438 ( \33083 , \7257 , \32486 );
and \U$27439 ( \33084 , \7259 , \32513 );
and \U$27440 ( \33085 , \9299 , \32540 );
and \U$27441 ( \33086 , \9301 , \32567 );
and \U$27442 ( \33087 , \9303 , \32594 );
and \U$27443 ( \33088 , \9305 , \32621 );
and \U$27444 ( \33089 , \9307 , \32648 );
and \U$27445 ( \33090 , \9309 , \32675 );
and \U$27446 ( \33091 , \9311 , \32702 );
and \U$27447 ( \33092 , \9313 , \32729 );
and \U$27448 ( \33093 , \9315 , \32756 );
and \U$27449 ( \33094 , \9317 , \32783 );
and \U$27450 ( \33095 , \9319 , \32810 );
and \U$27451 ( \33096 , \9321 , \32837 );
and \U$27452 ( \33097 , \9323 , \32864 );
and \U$27453 ( \33098 , \9325 , \32891 );
or \U$27454 ( \33099 , \33083 , \33084 , \33085 , \33086 , \33087 , \33088 , \33089 , \33090 , \33091 , \33092 , \33093 , \33094 , \33095 , \33096 , \33097 , \33098 );
_DC g985f ( \33100_nG985f , \33099 , \32968 );
buf \U$27455 ( \33101 , \33100_nG985f );
xor \U$27456 ( \33102 , \33082 , \33101 );
or \U$27457 ( \33103 , \33081 , \33102 );
buf \U$27458 ( \33104 , RIb7a0c48_261);
and \U$27459 ( \33105 , \7267 , \32486 );
and \U$27460 ( \33106 , \7269 , \32513 );
and \U$27461 ( \33107 , \9335 , \32540 );
and \U$27462 ( \33108 , \9337 , \32567 );
and \U$27463 ( \33109 , \9339 , \32594 );
and \U$27464 ( \33110 , \9341 , \32621 );
and \U$27465 ( \33111 , \9343 , \32648 );
and \U$27466 ( \33112 , \9345 , \32675 );
and \U$27467 ( \33113 , \9347 , \32702 );
and \U$27468 ( \33114 , \9349 , \32729 );
and \U$27469 ( \33115 , \9351 , \32756 );
and \U$27470 ( \33116 , \9353 , \32783 );
and \U$27471 ( \33117 , \9355 , \32810 );
and \U$27472 ( \33118 , \9357 , \32837 );
and \U$27473 ( \33119 , \9359 , \32864 );
and \U$27474 ( \33120 , \9361 , \32891 );
or \U$27475 ( \33121 , \33105 , \33106 , \33107 , \33108 , \33109 , \33110 , \33111 , \33112 , \33113 , \33114 , \33115 , \33116 , \33117 , \33118 , \33119 , \33120 );
_DC g9875 ( \33122_nG9875 , \33121 , \32968 );
buf \U$27476 ( \33123 , \33122_nG9875 );
xor \U$27477 ( \33124 , \33104 , \33123 );
or \U$27478 ( \33125 , \33103 , \33124 );
not \U$27479 ( \33126 , \33125 );
buf \U$27480 ( \33127 , \33126 );
and \U$27481 ( \33128 , \32459 , \33127 );
_HMUX g987c ( \33129_nG987c , \30892_nG8fb5 , \31263 , \33128 );
buf \U$27482 ( \33130 , \30909 );
buf \U$27483 ( \33131 , \30906 );
buf \U$27484 ( \33132 , \30894 );
buf \U$27485 ( \33133 , \30896 );
buf \U$27486 ( \33134 , \30899 );
buf \U$27487 ( \33135 , \30902 );
or \U$27488 ( \33136 , \33132 , \33133 , \33134 , \33135 );
and \U$27489 ( \33137 , \33131 , \33136 );
or \U$27490 ( \33138 , \33130 , \33137 );
buf \U$27491 ( \33139 , \33138 );
_HMUX g9887 ( \33140_nG9887 , \31262_nG9129 , \33129_nG987c , \33139 );
buf \U$27492 ( \33141 , RIe5319e0_6884);
not \U$27493 ( \33142 , \33141 );
buf \U$27494 ( \33143 , \33142 );
buf \U$27495 ( \33144 , RIe549ef0_6842);
xnor \U$27496 ( \33145 , \33144 , \33141 );
buf \U$27497 ( \33146 , \33145 );
buf \U$27498 ( \33147 , RIe549770_6843);
or \U$27499 ( \33148 , \33144 , \33141 );
xor \U$27500 ( \33149 , \33147 , \33148 );
buf \U$27501 ( \33150 , \33149 );
buf \U$27502 ( \33151 , RIe548ff0_6844);
and \U$27503 ( \33152 , \33147 , \33148 );
xor \U$27504 ( \33153 , \33151 , \33152 );
buf \U$27505 ( \33154 , \33153 );
buf \U$27506 ( \33155 , RIea91330_6888);
and \U$27507 ( \33156 , \33151 , \33152 );
xor \U$27508 ( \33157 , \33155 , \33156 );
buf \U$27509 ( \33158 , \33157 );
not \U$27510 ( \33159 , \33158 );
and \U$27511 ( \33160 , \33155 , \33156 );
buf \U$27512 ( \33161 , \33160 );
nor \U$27513 ( \33162 , \33143 , \33146 , \33150 , \33154 , \33159 , \33161 );
and \U$27514 ( \33163 , RIe5329d0_6883, \33162 );
not \U$27515 ( \33164 , \33161 );
and \U$27516 ( \33165 , \33143 , \33146 , \33150 , \33154 , \33159 , \33164 );
and \U$27517 ( \33166 , RIeb72150_6905, \33165 );
not \U$27518 ( \33167 , \33143 );
and \U$27519 ( \33168 , \33167 , \33146 , \33150 , \33154 , \33159 , \33164 );
and \U$27520 ( \33169 , RIeab80c0_6897, \33168 );
not \U$27521 ( \33170 , \33146 );
and \U$27522 ( \33171 , \33143 , \33170 , \33150 , \33154 , \33159 , \33164 );
and \U$27523 ( \33172 , RIe5331c8_6882, \33171 );
and \U$27524 ( \33173 , \33167 , \33170 , \33150 , \33154 , \33159 , \33164 );
and \U$27525 ( \33174 , RIe5339c0_6881, \33173 );
not \U$27526 ( \33175 , \33150 );
and \U$27527 ( \33176 , \33143 , \33146 , \33175 , \33154 , \33159 , \33164 );
and \U$27528 ( \33177 , RIeab87c8_6898, \33176 );
and \U$27529 ( \33178 , \33167 , \33146 , \33175 , \33154 , \33159 , \33164 );
and \U$27530 ( \33179 , RIe5341b8_6880, \33178 );
and \U$27531 ( \33180 , \33143 , \33170 , \33175 , \33154 , \33159 , \33164 );
and \U$27532 ( \33181 , RIe5349b0_6879, \33180 );
and \U$27533 ( \33182 , \33167 , \33170 , \33175 , \33154 , \33159 , \33164 );
and \U$27534 ( \33183 , RIea94af8_6890, \33182 );
nor \U$27535 ( \33184 , \33167 , \33170 , \33175 , \33154 , \33158 , \33161 );
and \U$27536 ( \33185 , RIe5351a8_6878, \33184 );
nor \U$27537 ( \33186 , \33143 , \33170 , \33175 , \33154 , \33158 , \33161 );
and \U$27538 ( \33187 , RIe5359a0_6877, \33186 );
nor \U$27539 ( \33188 , \33167 , \33146 , \33175 , \33154 , \33158 , \33161 );
and \U$27540 ( \33189 , RIeab78c8_6895, \33188 );
nor \U$27541 ( \33190 , \33143 , \33146 , \33175 , \33154 , \33158 , \33161 );
and \U$27542 ( \33191 , RIeab7d00_6896, \33190 );
nor \U$27543 ( \33192 , \33167 , \33170 , \33150 , \33154 , \33158 , \33161 );
and \U$27544 ( \33193 , RIeacfa18_6902, \33192 );
or \U$27547 ( \33194 , \33163 , \33166 , \33169 , \33172 , \33174 , \33177 , \33179 , \33181 , \33183 , \33185 , \33187 , \33189 , \33191 , \33193 , 1'b0 , 1'b0 );
buf \U$27549 ( \33195 , \33161 );
buf \U$27550 ( \33196 , \33158 );
buf \U$27551 ( \33197 , \33143 );
buf \U$27552 ( \33198 , \33146 );
buf \U$27553 ( \33199 , \33150 );
buf \U$27554 ( \33200 , \33154 );
or \U$27555 ( \33201 , \33197 , \33198 , \33199 , \33200 );
and \U$27556 ( \33202 , \33196 , \33201 );
or \U$27557 ( \33203 , \33195 , \33202 );
buf \U$27558 ( \33204 , \33203 );
or \U$27559 ( \33205 , 1'b0 , \33204 );
_DC g98c9 ( \33206_nG98c9 , \33194 , \33205 );
not \U$27560 ( \33207 , \33206_nG98c9 );
buf \U$27561 ( \33208 , RIb7b9608_246);
and \U$27562 ( \33209 , \7117 , \33162 );
and \U$27563 ( \33210 , \7119 , \33165 );
and \U$27564 ( \33211 , \7864 , \33168 );
and \U$27565 ( \33212 , \7892 , \33171 );
and \U$27566 ( \33213 , \7920 , \33173 );
and \U$27567 ( \33214 , \7948 , \33176 );
and \U$27568 ( \33215 , \7976 , \33178 );
and \U$27569 ( \33216 , \8004 , \33180 );
and \U$27570 ( \33217 , \8032 , \33182 );
and \U$27571 ( \33218 , \8060 , \33184 );
and \U$27572 ( \33219 , \8088 , \33186 );
and \U$27573 ( \33220 , \8116 , \33188 );
and \U$27574 ( \33221 , \8144 , \33190 );
and \U$27575 ( \33222 , \8172 , \33192 );
or \U$27578 ( \33223 , \33209 , \33210 , \33211 , \33212 , \33213 , \33214 , \33215 , \33216 , \33217 , \33218 , \33219 , \33220 , \33221 , \33222 , 1'b0 , 1'b0 );
_DC g98db ( \33224_nG98db , \33223 , \33205 );
buf \U$27579 ( \33225 , \33224_nG98db );
xor \U$27580 ( \33226 , \33208 , \33225 );
buf \U$27581 ( \33227 , RIb7b9590_247);
and \U$27582 ( \33228 , \7126 , \33162 );
and \U$27583 ( \33229 , \7128 , \33165 );
and \U$27584 ( \33230 , \8338 , \33168 );
and \U$27585 ( \33231 , \8340 , \33171 );
and \U$27586 ( \33232 , \8342 , \33173 );
and \U$27587 ( \33233 , \8344 , \33176 );
and \U$27588 ( \33234 , \8346 , \33178 );
and \U$27589 ( \33235 , \8348 , \33180 );
and \U$27590 ( \33236 , \8350 , \33182 );
and \U$27591 ( \33237 , \8352 , \33184 );
and \U$27592 ( \33238 , \8354 , \33186 );
and \U$27593 ( \33239 , \8356 , \33188 );
and \U$27594 ( \33240 , \8358 , \33190 );
and \U$27595 ( \33241 , \8360 , \33192 );
or \U$27598 ( \33242 , \33228 , \33229 , \33230 , \33231 , \33232 , \33233 , \33234 , \33235 , \33236 , \33237 , \33238 , \33239 , \33240 , \33241 , 1'b0 , 1'b0 );
_DC g98ee ( \33243_nG98ee , \33242 , \33205 );
buf \U$27599 ( \33244 , \33243_nG98ee );
xor \U$27600 ( \33245 , \33227 , \33244 );
or \U$27601 ( \33246 , \33226 , \33245 );
buf \U$27602 ( \33247 , RIb7b9518_248);
and \U$27603 ( \33248 , \7136 , \33162 );
and \U$27604 ( \33249 , \7138 , \33165 );
and \U$27605 ( \33250 , \8374 , \33168 );
and \U$27606 ( \33251 , \8376 , \33171 );
and \U$27607 ( \33252 , \8378 , \33173 );
and \U$27608 ( \33253 , \8380 , \33176 );
and \U$27609 ( \33254 , \8382 , \33178 );
and \U$27610 ( \33255 , \8384 , \33180 );
and \U$27611 ( \33256 , \8386 , \33182 );
and \U$27612 ( \33257 , \8388 , \33184 );
and \U$27613 ( \33258 , \8390 , \33186 );
and \U$27614 ( \33259 , \8392 , \33188 );
and \U$27615 ( \33260 , \8394 , \33190 );
and \U$27616 ( \33261 , \8396 , \33192 );
or \U$27619 ( \33262 , \33248 , \33249 , \33250 , \33251 , \33252 , \33253 , \33254 , \33255 , \33256 , \33257 , \33258 , \33259 , \33260 , \33261 , 1'b0 , 1'b0 );
_DC g9902 ( \33263_nG9902 , \33262 , \33205 );
buf \U$27620 ( \33264 , \33263_nG9902 );
xor \U$27621 ( \33265 , \33247 , \33264 );
or \U$27622 ( \33266 , \33246 , \33265 );
buf \U$27623 ( \33267 , RIb7b94a0_249);
and \U$27624 ( \33268 , \7146 , \33162 );
and \U$27625 ( \33269 , \7148 , \33165 );
and \U$27626 ( \33270 , \8410 , \33168 );
and \U$27627 ( \33271 , \8412 , \33171 );
and \U$27628 ( \33272 , \8414 , \33173 );
and \U$27629 ( \33273 , \8416 , \33176 );
and \U$27630 ( \33274 , \8418 , \33178 );
and \U$27631 ( \33275 , \8420 , \33180 );
and \U$27632 ( \33276 , \8422 , \33182 );
and \U$27633 ( \33277 , \8424 , \33184 );
and \U$27634 ( \33278 , \8426 , \33186 );
and \U$27635 ( \33279 , \8428 , \33188 );
and \U$27636 ( \33280 , \8430 , \33190 );
and \U$27637 ( \33281 , \8432 , \33192 );
or \U$27640 ( \33282 , \33268 , \33269 , \33270 , \33271 , \33272 , \33273 , \33274 , \33275 , \33276 , \33277 , \33278 , \33279 , \33280 , \33281 , 1'b0 , 1'b0 );
_DC g9916 ( \33283_nG9916 , \33282 , \33205 );
buf \U$27641 ( \33284 , \33283_nG9916 );
xor \U$27642 ( \33285 , \33267 , \33284 );
or \U$27643 ( \33286 , \33266 , \33285 );
buf \U$27644 ( \33287 , RIb7b9428_250);
and \U$27645 ( \33288 , \7156 , \33162 );
and \U$27646 ( \33289 , \7158 , \33165 );
and \U$27647 ( \33290 , \8446 , \33168 );
and \U$27648 ( \33291 , \8448 , \33171 );
and \U$27649 ( \33292 , \8450 , \33173 );
and \U$27650 ( \33293 , \8452 , \33176 );
and \U$27651 ( \33294 , \8454 , \33178 );
and \U$27652 ( \33295 , \8456 , \33180 );
and \U$27653 ( \33296 , \8458 , \33182 );
and \U$27654 ( \33297 , \8460 , \33184 );
and \U$27655 ( \33298 , \8462 , \33186 );
and \U$27656 ( \33299 , \8464 , \33188 );
and \U$27657 ( \33300 , \8466 , \33190 );
and \U$27658 ( \33301 , \8468 , \33192 );
or \U$27661 ( \33302 , \33288 , \33289 , \33290 , \33291 , \33292 , \33293 , \33294 , \33295 , \33296 , \33297 , \33298 , \33299 , \33300 , \33301 , 1'b0 , 1'b0 );
_DC g992a ( \33303_nG992a , \33302 , \33205 );
buf \U$27662 ( \33304 , \33303_nG992a );
xor \U$27663 ( \33305 , \33287 , \33304 );
or \U$27664 ( \33306 , \33286 , \33305 );
buf \U$27665 ( \33307 , RIb7b93b0_251);
and \U$27666 ( \33308 , \7166 , \33162 );
and \U$27667 ( \33309 , \7168 , \33165 );
and \U$27668 ( \33310 , \8482 , \33168 );
and \U$27669 ( \33311 , \8484 , \33171 );
and \U$27670 ( \33312 , \8486 , \33173 );
and \U$27671 ( \33313 , \8488 , \33176 );
and \U$27672 ( \33314 , \8490 , \33178 );
and \U$27673 ( \33315 , \8492 , \33180 );
and \U$27674 ( \33316 , \8494 , \33182 );
and \U$27675 ( \33317 , \8496 , \33184 );
and \U$27676 ( \33318 , \8498 , \33186 );
and \U$27677 ( \33319 , \8500 , \33188 );
and \U$27678 ( \33320 , \8502 , \33190 );
and \U$27679 ( \33321 , \8504 , \33192 );
or \U$27682 ( \33322 , \33308 , \33309 , \33310 , \33311 , \33312 , \33313 , \33314 , \33315 , \33316 , \33317 , \33318 , \33319 , \33320 , \33321 , 1'b0 , 1'b0 );
_DC g993e ( \33323_nG993e , \33322 , \33205 );
buf \U$27683 ( \33324 , \33323_nG993e );
xor \U$27684 ( \33325 , \33307 , \33324 );
or \U$27685 ( \33326 , \33306 , \33325 );
buf \U$27686 ( \33327 , RIb7af720_252);
and \U$27687 ( \33328 , \7176 , \33162 );
and \U$27688 ( \33329 , \7178 , \33165 );
and \U$27689 ( \33330 , \8518 , \33168 );
and \U$27690 ( \33331 , \8520 , \33171 );
and \U$27691 ( \33332 , \8522 , \33173 );
and \U$27692 ( \33333 , \8524 , \33176 );
and \U$27693 ( \33334 , \8526 , \33178 );
and \U$27694 ( \33335 , \8528 , \33180 );
and \U$27695 ( \33336 , \8530 , \33182 );
and \U$27696 ( \33337 , \8532 , \33184 );
and \U$27697 ( \33338 , \8534 , \33186 );
and \U$27698 ( \33339 , \8536 , \33188 );
and \U$27699 ( \33340 , \8538 , \33190 );
and \U$27700 ( \33341 , \8540 , \33192 );
or \U$27703 ( \33342 , \33328 , \33329 , \33330 , \33331 , \33332 , \33333 , \33334 , \33335 , \33336 , \33337 , \33338 , \33339 , \33340 , \33341 , 1'b0 , 1'b0 );
_DC g9952 ( \33343_nG9952 , \33342 , \33205 );
buf \U$27704 ( \33344 , \33343_nG9952 );
xor \U$27705 ( \33345 , \33327 , \33344 );
or \U$27706 ( \33346 , \33326 , \33345 );
buf \U$27707 ( \33347 , RIb7af6a8_253);
and \U$27708 ( \33348 , \7186 , \33162 );
and \U$27709 ( \33349 , \7188 , \33165 );
and \U$27710 ( \33350 , \8554 , \33168 );
and \U$27711 ( \33351 , \8556 , \33171 );
and \U$27712 ( \33352 , \8558 , \33173 );
and \U$27713 ( \33353 , \8560 , \33176 );
and \U$27714 ( \33354 , \8562 , \33178 );
and \U$27715 ( \33355 , \8564 , \33180 );
and \U$27716 ( \33356 , \8566 , \33182 );
and \U$27717 ( \33357 , \8568 , \33184 );
and \U$27718 ( \33358 , \8570 , \33186 );
and \U$27719 ( \33359 , \8572 , \33188 );
and \U$27720 ( \33360 , \8574 , \33190 );
and \U$27721 ( \33361 , \8576 , \33192 );
or \U$27724 ( \33362 , \33348 , \33349 , \33350 , \33351 , \33352 , \33353 , \33354 , \33355 , \33356 , \33357 , \33358 , \33359 , \33360 , \33361 , 1'b0 , 1'b0 );
_DC g9966 ( \33363_nG9966 , \33362 , \33205 );
buf \U$27725 ( \33364 , \33363_nG9966 );
xor \U$27726 ( \33365 , \33347 , \33364 );
or \U$27727 ( \33366 , \33346 , \33365 );
not \U$27728 ( \33367 , \33366 );
buf \U$27729 ( \33368 , \33367 );
buf \U$27730 ( \33369 , RIb7af630_254);
and \U$27731 ( \33370 , \7198 , \33162 );
and \U$27732 ( \33371 , \7200 , \33165 );
and \U$27733 ( \33372 , \8645 , \33168 );
and \U$27734 ( \33373 , \8673 , \33171 );
and \U$27735 ( \33374 , \8701 , \33173 );
and \U$27736 ( \33375 , \8729 , \33176 );
and \U$27737 ( \33376 , \8757 , \33178 );
and \U$27738 ( \33377 , \8785 , \33180 );
and \U$27739 ( \33378 , \8813 , \33182 );
and \U$27740 ( \33379 , \8841 , \33184 );
and \U$27741 ( \33380 , \8869 , \33186 );
and \U$27742 ( \33381 , \8897 , \33188 );
and \U$27743 ( \33382 , \8925 , \33190 );
and \U$27744 ( \33383 , \8953 , \33192 );
or \U$27747 ( \33384 , \33370 , \33371 , \33372 , \33373 , \33374 , \33375 , \33376 , \33377 , \33378 , \33379 , \33380 , \33381 , \33382 , \33383 , 1'b0 , 1'b0 );
_DC g997c ( \33385_nG997c , \33384 , \33205 );
buf \U$27748 ( \33386 , \33385_nG997c );
xor \U$27749 ( \33387 , \33369 , \33386 );
buf \U$27750 ( \33388 , RIb7af5b8_255);
and \U$27751 ( \33389 , \7207 , \33162 );
and \U$27752 ( \33390 , \7209 , \33165 );
and \U$27753 ( \33391 , \9119 , \33168 );
and \U$27754 ( \33392 , \9121 , \33171 );
and \U$27755 ( \33393 , \9123 , \33173 );
and \U$27756 ( \33394 , \9125 , \33176 );
and \U$27757 ( \33395 , \9127 , \33178 );
and \U$27758 ( \33396 , \9129 , \33180 );
and \U$27759 ( \33397 , \9131 , \33182 );
and \U$27760 ( \33398 , \9133 , \33184 );
and \U$27761 ( \33399 , \9135 , \33186 );
and \U$27762 ( \33400 , \9137 , \33188 );
and \U$27763 ( \33401 , \9139 , \33190 );
and \U$27764 ( \33402 , \9141 , \33192 );
or \U$27767 ( \33403 , \33389 , \33390 , \33391 , \33392 , \33393 , \33394 , \33395 , \33396 , \33397 , \33398 , \33399 , \33400 , \33401 , \33402 , 1'b0 , 1'b0 );
_DC g998f ( \33404_nG998f , \33403 , \33205 );
buf \U$27768 ( \33405 , \33404_nG998f );
xor \U$27769 ( \33406 , \33388 , \33405 );
or \U$27770 ( \33407 , \33387 , \33406 );
buf \U$27771 ( \33408 , RIb7af540_256);
and \U$27772 ( \33409 , \7217 , \33162 );
and \U$27773 ( \33410 , \7219 , \33165 );
and \U$27774 ( \33411 , \9155 , \33168 );
and \U$27775 ( \33412 , \9157 , \33171 );
and \U$27776 ( \33413 , \9159 , \33173 );
and \U$27777 ( \33414 , \9161 , \33176 );
and \U$27778 ( \33415 , \9163 , \33178 );
and \U$27779 ( \33416 , \9165 , \33180 );
and \U$27780 ( \33417 , \9167 , \33182 );
and \U$27781 ( \33418 , \9169 , \33184 );
and \U$27782 ( \33419 , \9171 , \33186 );
and \U$27783 ( \33420 , \9173 , \33188 );
and \U$27784 ( \33421 , \9175 , \33190 );
and \U$27785 ( \33422 , \9177 , \33192 );
or \U$27788 ( \33423 , \33409 , \33410 , \33411 , \33412 , \33413 , \33414 , \33415 , \33416 , \33417 , \33418 , \33419 , \33420 , \33421 , \33422 , 1'b0 , 1'b0 );
_DC g99a3 ( \33424_nG99a3 , \33423 , \33205 );
buf \U$27789 ( \33425 , \33424_nG99a3 );
xor \U$27790 ( \33426 , \33408 , \33425 );
or \U$27791 ( \33427 , \33407 , \33426 );
buf \U$27792 ( \33428 , RIb7af4c8_257);
and \U$27793 ( \33429 , \7227 , \33162 );
and \U$27794 ( \33430 , \7229 , \33165 );
and \U$27795 ( \33431 , \9191 , \33168 );
and \U$27796 ( \33432 , \9193 , \33171 );
and \U$27797 ( \33433 , \9195 , \33173 );
and \U$27798 ( \33434 , \9197 , \33176 );
and \U$27799 ( \33435 , \9199 , \33178 );
and \U$27800 ( \33436 , \9201 , \33180 );
and \U$27801 ( \33437 , \9203 , \33182 );
and \U$27802 ( \33438 , \9205 , \33184 );
and \U$27803 ( \33439 , \9207 , \33186 );
and \U$27804 ( \33440 , \9209 , \33188 );
and \U$27805 ( \33441 , \9211 , \33190 );
and \U$27806 ( \33442 , \9213 , \33192 );
or \U$27809 ( \33443 , \33429 , \33430 , \33431 , \33432 , \33433 , \33434 , \33435 , \33436 , \33437 , \33438 , \33439 , \33440 , \33441 , \33442 , 1'b0 , 1'b0 );
_DC g99b7 ( \33444_nG99b7 , \33443 , \33205 );
buf \U$27810 ( \33445 , \33444_nG99b7 );
xor \U$27811 ( \33446 , \33428 , \33445 );
or \U$27812 ( \33447 , \33427 , \33446 );
buf \U$27813 ( \33448 , RIb7af450_258);
and \U$27814 ( \33449 , \7237 , \33162 );
and \U$27815 ( \33450 , \7239 , \33165 );
and \U$27816 ( \33451 , \9227 , \33168 );
and \U$27817 ( \33452 , \9229 , \33171 );
and \U$27818 ( \33453 , \9231 , \33173 );
and \U$27819 ( \33454 , \9233 , \33176 );
and \U$27820 ( \33455 , \9235 , \33178 );
and \U$27821 ( \33456 , \9237 , \33180 );
and \U$27822 ( \33457 , \9239 , \33182 );
and \U$27823 ( \33458 , \9241 , \33184 );
and \U$27824 ( \33459 , \9243 , \33186 );
and \U$27825 ( \33460 , \9245 , \33188 );
and \U$27826 ( \33461 , \9247 , \33190 );
and \U$27827 ( \33462 , \9249 , \33192 );
or \U$27830 ( \33463 , \33449 , \33450 , \33451 , \33452 , \33453 , \33454 , \33455 , \33456 , \33457 , \33458 , \33459 , \33460 , \33461 , \33462 , 1'b0 , 1'b0 );
_DC g99cb ( \33464_nG99cb , \33463 , \33205 );
buf \U$27831 ( \33465 , \33464_nG99cb );
xor \U$27832 ( \33466 , \33448 , \33465 );
or \U$27833 ( \33467 , \33447 , \33466 );
buf \U$27834 ( \33468 , RIb7af3d8_259);
and \U$27835 ( \33469 , \7247 , \33162 );
and \U$27836 ( \33470 , \7249 , \33165 );
and \U$27837 ( \33471 , \9263 , \33168 );
and \U$27838 ( \33472 , \9265 , \33171 );
and \U$27839 ( \33473 , \9267 , \33173 );
and \U$27840 ( \33474 , \9269 , \33176 );
and \U$27841 ( \33475 , \9271 , \33178 );
and \U$27842 ( \33476 , \9273 , \33180 );
and \U$27843 ( \33477 , \9275 , \33182 );
and \U$27844 ( \33478 , \9277 , \33184 );
and \U$27845 ( \33479 , \9279 , \33186 );
and \U$27846 ( \33480 , \9281 , \33188 );
and \U$27847 ( \33481 , \9283 , \33190 );
and \U$27848 ( \33482 , \9285 , \33192 );
or \U$27851 ( \33483 , \33469 , \33470 , \33471 , \33472 , \33473 , \33474 , \33475 , \33476 , \33477 , \33478 , \33479 , \33480 , \33481 , \33482 , 1'b0 , 1'b0 );
_DC g99df ( \33484_nG99df , \33483 , \33205 );
buf \U$27852 ( \33485 , \33484_nG99df );
xor \U$27853 ( \33486 , \33468 , \33485 );
or \U$27854 ( \33487 , \33467 , \33486 );
buf \U$27855 ( \33488 , RIb7a5bf8_260);
and \U$27856 ( \33489 , \7257 , \33162 );
and \U$27857 ( \33490 , \7259 , \33165 );
and \U$27858 ( \33491 , \9299 , \33168 );
and \U$27859 ( \33492 , \9301 , \33171 );
and \U$27860 ( \33493 , \9303 , \33173 );
and \U$27861 ( \33494 , \9305 , \33176 );
and \U$27862 ( \33495 , \9307 , \33178 );
and \U$27863 ( \33496 , \9309 , \33180 );
and \U$27864 ( \33497 , \9311 , \33182 );
and \U$27865 ( \33498 , \9313 , \33184 );
and \U$27866 ( \33499 , \9315 , \33186 );
and \U$27867 ( \33500 , \9317 , \33188 );
and \U$27868 ( \33501 , \9319 , \33190 );
and \U$27869 ( \33502 , \9321 , \33192 );
or \U$27872 ( \33503 , \33489 , \33490 , \33491 , \33492 , \33493 , \33494 , \33495 , \33496 , \33497 , \33498 , \33499 , \33500 , \33501 , \33502 , 1'b0 , 1'b0 );
_DC g99f3 ( \33504_nG99f3 , \33503 , \33205 );
buf \U$27873 ( \33505 , \33504_nG99f3 );
xor \U$27874 ( \33506 , \33488 , \33505 );
or \U$27875 ( \33507 , \33487 , \33506 );
buf \U$27876 ( \33508 , RIb7a0c48_261);
and \U$27877 ( \33509 , \7267 , \33162 );
and \U$27878 ( \33510 , \7269 , \33165 );
and \U$27879 ( \33511 , \9335 , \33168 );
and \U$27880 ( \33512 , \9337 , \33171 );
and \U$27881 ( \33513 , \9339 , \33173 );
and \U$27882 ( \33514 , \9341 , \33176 );
and \U$27883 ( \33515 , \9343 , \33178 );
and \U$27884 ( \33516 , \9345 , \33180 );
and \U$27885 ( \33517 , \9347 , \33182 );
and \U$27886 ( \33518 , \9349 , \33184 );
and \U$27887 ( \33519 , \9351 , \33186 );
and \U$27888 ( \33520 , \9353 , \33188 );
and \U$27889 ( \33521 , \9355 , \33190 );
and \U$27890 ( \33522 , \9357 , \33192 );
or \U$27893 ( \33523 , \33509 , \33510 , \33511 , \33512 , \33513 , \33514 , \33515 , \33516 , \33517 , \33518 , \33519 , \33520 , \33521 , \33522 , 1'b0 , 1'b0 );
_DC g9a07 ( \33524_nG9a07 , \33523 , \33205 );
buf \U$27894 ( \33525 , \33524_nG9a07 );
xor \U$27895 ( \33526 , \33508 , \33525 );
or \U$27896 ( \33527 , \33507 , \33526 );
not \U$27897 ( \33528 , \33527 );
buf \U$27898 ( \33529 , \33528 );
and \U$27899 ( \33530 , \33368 , \33529 );
and \U$27900 ( \33531 , \33207 , \33530 );
_HMUX g9a0f ( \33532_nG9a0f , \33140_nG9887 , \33143 , \33531 );
buf \U$27903 ( \33533 , \33143 );
buf \U$27906 ( \33534 , \33146 );
buf \U$27909 ( \33535 , \33150 );
buf \U$27912 ( \33536 , \33154 );
buf \U$27913 ( \33537 , \33158 );
not \U$27914 ( \33538 , \33537 );
buf \U$27915 ( \33539 , \33538 );
not \U$27916 ( \33540 , \33539 );
buf \U$27917 ( \33541 , \33161 );
xnor \U$27918 ( \33542 , \33541 , \33537 );
buf \U$27919 ( \33543 , \33542 );
or \U$27920 ( \33544 , \33541 , \33537 );
not \U$27921 ( \33545 , \33544 );
buf \U$27922 ( \33546 , \33545 );
buf \U$27923 ( \33547 , \33546 );
buf \U$27924 ( \33548 , \33546 );
buf \U$27925 ( \33549 , \33546 );
buf \U$27926 ( \33550 , \33546 );
buf \U$27927 ( \33551 , \33546 );
buf \U$27928 ( \33552 , \33546 );
buf \U$27929 ( \33553 , \33546 );
buf \U$27930 ( \33554 , \33546 );
buf \U$27931 ( \33555 , \33546 );
buf \U$27932 ( \33556 , \33546 );
buf \U$27933 ( \33557 , \33546 );
buf \U$27934 ( \33558 , \33546 );
buf \U$27935 ( \33559 , \33546 );
buf \U$27936 ( \33560 , \33546 );
buf \U$27937 ( \33561 , \33546 );
buf \U$27938 ( \33562 , \33546 );
buf \U$27939 ( \33563 , \33546 );
buf \U$27940 ( \33564 , \33546 );
buf \U$27941 ( \33565 , \33546 );
buf \U$27942 ( \33566 , \33546 );
buf \U$27943 ( \33567 , \33546 );
buf \U$27944 ( \33568 , \33546 );
buf \U$27945 ( \33569 , \33546 );
buf \U$27946 ( \33570 , \33546 );
buf \U$27947 ( \33571 , \33546 );
nor \U$27948 ( \33572 , \33533 , \33534 , \33535 , \33536 , \33540 , \33543 , \33546 , \33547 , \33548 , \33549 , \33550 , \33551 , \33552 , \33553 , \33554 , \33555 , \33556 , \33557 , \33558 , \33559 , \33560 , \33561 , \33562 , \33563 , \33564 , \33565 , \33566 , \33567 , \33568 , \33569 , \33570 , \33571 );
and \U$27949 ( \33573 , RIe5329d0_6883, \33572 );
not \U$27950 ( \33574 , \33533 );
not \U$27951 ( \33575 , \33534 );
not \U$27952 ( \33576 , \33535 );
not \U$27953 ( \33577 , \33536 );
buf \U$27954 ( \33578 , \33546 );
buf \U$27955 ( \33579 , \33546 );
buf \U$27956 ( \33580 , \33546 );
buf \U$27957 ( \33581 , \33546 );
buf \U$27958 ( \33582 , \33546 );
buf \U$27959 ( \33583 , \33546 );
buf \U$27960 ( \33584 , \33546 );
buf \U$27961 ( \33585 , \33546 );
buf \U$27962 ( \33586 , \33546 );
buf \U$27963 ( \33587 , \33546 );
buf \U$27964 ( \33588 , \33546 );
buf \U$27965 ( \33589 , \33546 );
buf \U$27966 ( \33590 , \33546 );
buf \U$27967 ( \33591 , \33546 );
buf \U$27968 ( \33592 , \33546 );
buf \U$27969 ( \33593 , \33546 );
buf \U$27970 ( \33594 , \33546 );
buf \U$27971 ( \33595 , \33546 );
buf \U$27972 ( \33596 , \33546 );
buf \U$27973 ( \33597 , \33546 );
buf \U$27974 ( \33598 , \33546 );
buf \U$27975 ( \33599 , \33546 );
buf \U$27976 ( \33600 , \33546 );
buf \U$27977 ( \33601 , \33546 );
buf \U$27978 ( \33602 , \33546 );
nor \U$27979 ( \33603 , \33574 , \33575 , \33576 , \33577 , \33539 , \33543 , \33546 , \33578 , \33579 , \33580 , \33581 , \33582 , \33583 , \33584 , \33585 , \33586 , \33587 , \33588 , \33589 , \33590 , \33591 , \33592 , \33593 , \33594 , \33595 , \33596 , \33597 , \33598 , \33599 , \33600 , \33601 , \33602 );
and \U$27980 ( \33604 , RIeb72150_6905, \33603 );
buf \U$27981 ( \33605 , \33546 );
buf \U$27982 ( \33606 , \33546 );
buf \U$27983 ( \33607 , \33546 );
buf \U$27984 ( \33608 , \33546 );
buf \U$27985 ( \33609 , \33546 );
buf \U$27986 ( \33610 , \33546 );
buf \U$27987 ( \33611 , \33546 );
buf \U$27988 ( \33612 , \33546 );
buf \U$27989 ( \33613 , \33546 );
buf \U$27990 ( \33614 , \33546 );
buf \U$27991 ( \33615 , \33546 );
buf \U$27992 ( \33616 , \33546 );
buf \U$27993 ( \33617 , \33546 );
buf \U$27994 ( \33618 , \33546 );
buf \U$27995 ( \33619 , \33546 );
buf \U$27996 ( \33620 , \33546 );
buf \U$27997 ( \33621 , \33546 );
buf \U$27998 ( \33622 , \33546 );
buf \U$27999 ( \33623 , \33546 );
buf \U$28000 ( \33624 , \33546 );
buf \U$28001 ( \33625 , \33546 );
buf \U$28002 ( \33626 , \33546 );
buf \U$28003 ( \33627 , \33546 );
buf \U$28004 ( \33628 , \33546 );
buf \U$28005 ( \33629 , \33546 );
nor \U$28006 ( \33630 , \33533 , \33575 , \33576 , \33577 , \33539 , \33543 , \33546 , \33605 , \33606 , \33607 , \33608 , \33609 , \33610 , \33611 , \33612 , \33613 , \33614 , \33615 , \33616 , \33617 , \33618 , \33619 , \33620 , \33621 , \33622 , \33623 , \33624 , \33625 , \33626 , \33627 , \33628 , \33629 );
and \U$28007 ( \33631 , RIeab80c0_6897, \33630 );
buf \U$28008 ( \33632 , \33546 );
buf \U$28009 ( \33633 , \33546 );
buf \U$28010 ( \33634 , \33546 );
buf \U$28011 ( \33635 , \33546 );
buf \U$28012 ( \33636 , \33546 );
buf \U$28013 ( \33637 , \33546 );
buf \U$28014 ( \33638 , \33546 );
buf \U$28015 ( \33639 , \33546 );
buf \U$28016 ( \33640 , \33546 );
buf \U$28017 ( \33641 , \33546 );
buf \U$28018 ( \33642 , \33546 );
buf \U$28019 ( \33643 , \33546 );
buf \U$28020 ( \33644 , \33546 );
buf \U$28021 ( \33645 , \33546 );
buf \U$28022 ( \33646 , \33546 );
buf \U$28023 ( \33647 , \33546 );
buf \U$28024 ( \33648 , \33546 );
buf \U$28025 ( \33649 , \33546 );
buf \U$28026 ( \33650 , \33546 );
buf \U$28027 ( \33651 , \33546 );
buf \U$28028 ( \33652 , \33546 );
buf \U$28029 ( \33653 , \33546 );
buf \U$28030 ( \33654 , \33546 );
buf \U$28031 ( \33655 , \33546 );
buf \U$28032 ( \33656 , \33546 );
nor \U$28033 ( \33657 , \33574 , \33534 , \33576 , \33577 , \33539 , \33543 , \33546 , \33632 , \33633 , \33634 , \33635 , \33636 , \33637 , \33638 , \33639 , \33640 , \33641 , \33642 , \33643 , \33644 , \33645 , \33646 , \33647 , \33648 , \33649 , \33650 , \33651 , \33652 , \33653 , \33654 , \33655 , \33656 );
and \U$28034 ( \33658 , RIe5331c8_6882, \33657 );
buf \U$28035 ( \33659 , \33546 );
buf \U$28036 ( \33660 , \33546 );
buf \U$28037 ( \33661 , \33546 );
buf \U$28038 ( \33662 , \33546 );
buf \U$28039 ( \33663 , \33546 );
buf \U$28040 ( \33664 , \33546 );
buf \U$28041 ( \33665 , \33546 );
buf \U$28042 ( \33666 , \33546 );
buf \U$28043 ( \33667 , \33546 );
buf \U$28044 ( \33668 , \33546 );
buf \U$28045 ( \33669 , \33546 );
buf \U$28046 ( \33670 , \33546 );
buf \U$28047 ( \33671 , \33546 );
buf \U$28048 ( \33672 , \33546 );
buf \U$28049 ( \33673 , \33546 );
buf \U$28050 ( \33674 , \33546 );
buf \U$28051 ( \33675 , \33546 );
buf \U$28052 ( \33676 , \33546 );
buf \U$28053 ( \33677 , \33546 );
buf \U$28054 ( \33678 , \33546 );
buf \U$28055 ( \33679 , \33546 );
buf \U$28056 ( \33680 , \33546 );
buf \U$28057 ( \33681 , \33546 );
buf \U$28058 ( \33682 , \33546 );
buf \U$28059 ( \33683 , \33546 );
nor \U$28060 ( \33684 , \33533 , \33534 , \33576 , \33577 , \33539 , \33543 , \33546 , \33659 , \33660 , \33661 , \33662 , \33663 , \33664 , \33665 , \33666 , \33667 , \33668 , \33669 , \33670 , \33671 , \33672 , \33673 , \33674 , \33675 , \33676 , \33677 , \33678 , \33679 , \33680 , \33681 , \33682 , \33683 );
and \U$28061 ( \33685 , RIe5339c0_6881, \33684 );
buf \U$28062 ( \33686 , \33546 );
buf \U$28063 ( \33687 , \33546 );
buf \U$28064 ( \33688 , \33546 );
buf \U$28065 ( \33689 , \33546 );
buf \U$28066 ( \33690 , \33546 );
buf \U$28067 ( \33691 , \33546 );
buf \U$28068 ( \33692 , \33546 );
buf \U$28069 ( \33693 , \33546 );
buf \U$28070 ( \33694 , \33546 );
buf \U$28071 ( \33695 , \33546 );
buf \U$28072 ( \33696 , \33546 );
buf \U$28073 ( \33697 , \33546 );
buf \U$28074 ( \33698 , \33546 );
buf \U$28075 ( \33699 , \33546 );
buf \U$28076 ( \33700 , \33546 );
buf \U$28077 ( \33701 , \33546 );
buf \U$28078 ( \33702 , \33546 );
buf \U$28079 ( \33703 , \33546 );
buf \U$28080 ( \33704 , \33546 );
buf \U$28081 ( \33705 , \33546 );
buf \U$28082 ( \33706 , \33546 );
buf \U$28083 ( \33707 , \33546 );
buf \U$28084 ( \33708 , \33546 );
buf \U$28085 ( \33709 , \33546 );
buf \U$28086 ( \33710 , \33546 );
nor \U$28087 ( \33711 , \33574 , \33575 , \33535 , \33577 , \33539 , \33543 , \33546 , \33686 , \33687 , \33688 , \33689 , \33690 , \33691 , \33692 , \33693 , \33694 , \33695 , \33696 , \33697 , \33698 , \33699 , \33700 , \33701 , \33702 , \33703 , \33704 , \33705 , \33706 , \33707 , \33708 , \33709 , \33710 );
and \U$28088 ( \33712 , RIeab87c8_6898, \33711 );
buf \U$28089 ( \33713 , \33546 );
buf \U$28090 ( \33714 , \33546 );
buf \U$28091 ( \33715 , \33546 );
buf \U$28092 ( \33716 , \33546 );
buf \U$28093 ( \33717 , \33546 );
buf \U$28094 ( \33718 , \33546 );
buf \U$28095 ( \33719 , \33546 );
buf \U$28096 ( \33720 , \33546 );
buf \U$28097 ( \33721 , \33546 );
buf \U$28098 ( \33722 , \33546 );
buf \U$28099 ( \33723 , \33546 );
buf \U$28100 ( \33724 , \33546 );
buf \U$28101 ( \33725 , \33546 );
buf \U$28102 ( \33726 , \33546 );
buf \U$28103 ( \33727 , \33546 );
buf \U$28104 ( \33728 , \33546 );
buf \U$28105 ( \33729 , \33546 );
buf \U$28106 ( \33730 , \33546 );
buf \U$28107 ( \33731 , \33546 );
buf \U$28108 ( \33732 , \33546 );
buf \U$28109 ( \33733 , \33546 );
buf \U$28110 ( \33734 , \33546 );
buf \U$28111 ( \33735 , \33546 );
buf \U$28112 ( \33736 , \33546 );
buf \U$28113 ( \33737 , \33546 );
nor \U$28114 ( \33738 , \33533 , \33575 , \33535 , \33577 , \33539 , \33543 , \33546 , \33713 , \33714 , \33715 , \33716 , \33717 , \33718 , \33719 , \33720 , \33721 , \33722 , \33723 , \33724 , \33725 , \33726 , \33727 , \33728 , \33729 , \33730 , \33731 , \33732 , \33733 , \33734 , \33735 , \33736 , \33737 );
and \U$28115 ( \33739 , RIe5341b8_6880, \33738 );
buf \U$28116 ( \33740 , \33546 );
buf \U$28117 ( \33741 , \33546 );
buf \U$28118 ( \33742 , \33546 );
buf \U$28119 ( \33743 , \33546 );
buf \U$28120 ( \33744 , \33546 );
buf \U$28121 ( \33745 , \33546 );
buf \U$28122 ( \33746 , \33546 );
buf \U$28123 ( \33747 , \33546 );
buf \U$28124 ( \33748 , \33546 );
buf \U$28125 ( \33749 , \33546 );
buf \U$28126 ( \33750 , \33546 );
buf \U$28127 ( \33751 , \33546 );
buf \U$28128 ( \33752 , \33546 );
buf \U$28129 ( \33753 , \33546 );
buf \U$28130 ( \33754 , \33546 );
buf \U$28131 ( \33755 , \33546 );
buf \U$28132 ( \33756 , \33546 );
buf \U$28133 ( \33757 , \33546 );
buf \U$28134 ( \33758 , \33546 );
buf \U$28135 ( \33759 , \33546 );
buf \U$28136 ( \33760 , \33546 );
buf \U$28137 ( \33761 , \33546 );
buf \U$28138 ( \33762 , \33546 );
buf \U$28139 ( \33763 , \33546 );
buf \U$28140 ( \33764 , \33546 );
nor \U$28141 ( \33765 , \33574 , \33534 , \33535 , \33577 , \33539 , \33543 , \33546 , \33740 , \33741 , \33742 , \33743 , \33744 , \33745 , \33746 , \33747 , \33748 , \33749 , \33750 , \33751 , \33752 , \33753 , \33754 , \33755 , \33756 , \33757 , \33758 , \33759 , \33760 , \33761 , \33762 , \33763 , \33764 );
and \U$28142 ( \33766 , RIe5349b0_6879, \33765 );
buf \U$28143 ( \33767 , \33546 );
buf \U$28144 ( \33768 , \33546 );
buf \U$28145 ( \33769 , \33546 );
buf \U$28146 ( \33770 , \33546 );
buf \U$28147 ( \33771 , \33546 );
buf \U$28148 ( \33772 , \33546 );
buf \U$28149 ( \33773 , \33546 );
buf \U$28150 ( \33774 , \33546 );
buf \U$28151 ( \33775 , \33546 );
buf \U$28152 ( \33776 , \33546 );
buf \U$28153 ( \33777 , \33546 );
buf \U$28154 ( \33778 , \33546 );
buf \U$28155 ( \33779 , \33546 );
buf \U$28156 ( \33780 , \33546 );
buf \U$28157 ( \33781 , \33546 );
buf \U$28158 ( \33782 , \33546 );
buf \U$28159 ( \33783 , \33546 );
buf \U$28160 ( \33784 , \33546 );
buf \U$28161 ( \33785 , \33546 );
buf \U$28162 ( \33786 , \33546 );
buf \U$28163 ( \33787 , \33546 );
buf \U$28164 ( \33788 , \33546 );
buf \U$28165 ( \33789 , \33546 );
buf \U$28166 ( \33790 , \33546 );
buf \U$28167 ( \33791 , \33546 );
nor \U$28168 ( \33792 , \33533 , \33534 , \33535 , \33577 , \33539 , \33543 , \33546 , \33767 , \33768 , \33769 , \33770 , \33771 , \33772 , \33773 , \33774 , \33775 , \33776 , \33777 , \33778 , \33779 , \33780 , \33781 , \33782 , \33783 , \33784 , \33785 , \33786 , \33787 , \33788 , \33789 , \33790 , \33791 );
and \U$28169 ( \33793 , RIea94af8_6890, \33792 );
buf \U$28170 ( \33794 , \33546 );
buf \U$28171 ( \33795 , \33546 );
buf \U$28172 ( \33796 , \33546 );
buf \U$28173 ( \33797 , \33546 );
buf \U$28174 ( \33798 , \33546 );
buf \U$28175 ( \33799 , \33546 );
buf \U$28176 ( \33800 , \33546 );
buf \U$28177 ( \33801 , \33546 );
buf \U$28178 ( \33802 , \33546 );
buf \U$28179 ( \33803 , \33546 );
buf \U$28180 ( \33804 , \33546 );
buf \U$28181 ( \33805 , \33546 );
buf \U$28182 ( \33806 , \33546 );
buf \U$28183 ( \33807 , \33546 );
buf \U$28184 ( \33808 , \33546 );
buf \U$28185 ( \33809 , \33546 );
buf \U$28186 ( \33810 , \33546 );
buf \U$28187 ( \33811 , \33546 );
buf \U$28188 ( \33812 , \33546 );
buf \U$28189 ( \33813 , \33546 );
buf \U$28190 ( \33814 , \33546 );
buf \U$28191 ( \33815 , \33546 );
buf \U$28192 ( \33816 , \33546 );
buf \U$28193 ( \33817 , \33546 );
buf \U$28194 ( \33818 , \33546 );
nor \U$28195 ( \33819 , \33574 , \33575 , \33576 , \33536 , \33539 , \33543 , \33546 , \33794 , \33795 , \33796 , \33797 , \33798 , \33799 , \33800 , \33801 , \33802 , \33803 , \33804 , \33805 , \33806 , \33807 , \33808 , \33809 , \33810 , \33811 , \33812 , \33813 , \33814 , \33815 , \33816 , \33817 , \33818 );
and \U$28196 ( \33820 , RIe5351a8_6878, \33819 );
buf \U$28197 ( \33821 , \33546 );
buf \U$28198 ( \33822 , \33546 );
buf \U$28199 ( \33823 , \33546 );
buf \U$28200 ( \33824 , \33546 );
buf \U$28201 ( \33825 , \33546 );
buf \U$28202 ( \33826 , \33546 );
buf \U$28203 ( \33827 , \33546 );
buf \U$28204 ( \33828 , \33546 );
buf \U$28205 ( \33829 , \33546 );
buf \U$28206 ( \33830 , \33546 );
buf \U$28207 ( \33831 , \33546 );
buf \U$28208 ( \33832 , \33546 );
buf \U$28209 ( \33833 , \33546 );
buf \U$28210 ( \33834 , \33546 );
buf \U$28211 ( \33835 , \33546 );
buf \U$28212 ( \33836 , \33546 );
buf \U$28213 ( \33837 , \33546 );
buf \U$28214 ( \33838 , \33546 );
buf \U$28215 ( \33839 , \33546 );
buf \U$28216 ( \33840 , \33546 );
buf \U$28217 ( \33841 , \33546 );
buf \U$28218 ( \33842 , \33546 );
buf \U$28219 ( \33843 , \33546 );
buf \U$28220 ( \33844 , \33546 );
buf \U$28221 ( \33845 , \33546 );
nor \U$28222 ( \33846 , \33533 , \33575 , \33576 , \33536 , \33539 , \33543 , \33546 , \33821 , \33822 , \33823 , \33824 , \33825 , \33826 , \33827 , \33828 , \33829 , \33830 , \33831 , \33832 , \33833 , \33834 , \33835 , \33836 , \33837 , \33838 , \33839 , \33840 , \33841 , \33842 , \33843 , \33844 , \33845 );
and \U$28223 ( \33847 , RIe5359a0_6877, \33846 );
buf \U$28224 ( \33848 , \33546 );
buf \U$28225 ( \33849 , \33546 );
buf \U$28226 ( \33850 , \33546 );
buf \U$28227 ( \33851 , \33546 );
buf \U$28228 ( \33852 , \33546 );
buf \U$28229 ( \33853 , \33546 );
buf \U$28230 ( \33854 , \33546 );
buf \U$28231 ( \33855 , \33546 );
buf \U$28232 ( \33856 , \33546 );
buf \U$28233 ( \33857 , \33546 );
buf \U$28234 ( \33858 , \33546 );
buf \U$28235 ( \33859 , \33546 );
buf \U$28236 ( \33860 , \33546 );
buf \U$28237 ( \33861 , \33546 );
buf \U$28238 ( \33862 , \33546 );
buf \U$28239 ( \33863 , \33546 );
buf \U$28240 ( \33864 , \33546 );
buf \U$28241 ( \33865 , \33546 );
buf \U$28242 ( \33866 , \33546 );
buf \U$28243 ( \33867 , \33546 );
buf \U$28244 ( \33868 , \33546 );
buf \U$28245 ( \33869 , \33546 );
buf \U$28246 ( \33870 , \33546 );
buf \U$28247 ( \33871 , \33546 );
buf \U$28248 ( \33872 , \33546 );
nor \U$28249 ( \33873 , \33574 , \33534 , \33576 , \33536 , \33539 , \33543 , \33546 , \33848 , \33849 , \33850 , \33851 , \33852 , \33853 , \33854 , \33855 , \33856 , \33857 , \33858 , \33859 , \33860 , \33861 , \33862 , \33863 , \33864 , \33865 , \33866 , \33867 , \33868 , \33869 , \33870 , \33871 , \33872 );
and \U$28250 ( \33874 , RIeab78c8_6895, \33873 );
buf \U$28251 ( \33875 , \33546 );
buf \U$28252 ( \33876 , \33546 );
buf \U$28253 ( \33877 , \33546 );
buf \U$28254 ( \33878 , \33546 );
buf \U$28255 ( \33879 , \33546 );
buf \U$28256 ( \33880 , \33546 );
buf \U$28257 ( \33881 , \33546 );
buf \U$28258 ( \33882 , \33546 );
buf \U$28259 ( \33883 , \33546 );
buf \U$28260 ( \33884 , \33546 );
buf \U$28261 ( \33885 , \33546 );
buf \U$28262 ( \33886 , \33546 );
buf \U$28263 ( \33887 , \33546 );
buf \U$28264 ( \33888 , \33546 );
buf \U$28265 ( \33889 , \33546 );
buf \U$28266 ( \33890 , \33546 );
buf \U$28267 ( \33891 , \33546 );
buf \U$28268 ( \33892 , \33546 );
buf \U$28269 ( \33893 , \33546 );
buf \U$28270 ( \33894 , \33546 );
buf \U$28271 ( \33895 , \33546 );
buf \U$28272 ( \33896 , \33546 );
buf \U$28273 ( \33897 , \33546 );
buf \U$28274 ( \33898 , \33546 );
buf \U$28275 ( \33899 , \33546 );
nor \U$28276 ( \33900 , \33533 , \33534 , \33576 , \33536 , \33539 , \33543 , \33546 , \33875 , \33876 , \33877 , \33878 , \33879 , \33880 , \33881 , \33882 , \33883 , \33884 , \33885 , \33886 , \33887 , \33888 , \33889 , \33890 , \33891 , \33892 , \33893 , \33894 , \33895 , \33896 , \33897 , \33898 , \33899 );
and \U$28277 ( \33901 , RIeab7d00_6896, \33900 );
buf \U$28278 ( \33902 , \33546 );
buf \U$28279 ( \33903 , \33546 );
buf \U$28280 ( \33904 , \33546 );
buf \U$28281 ( \33905 , \33546 );
buf \U$28282 ( \33906 , \33546 );
buf \U$28283 ( \33907 , \33546 );
buf \U$28284 ( \33908 , \33546 );
buf \U$28285 ( \33909 , \33546 );
buf \U$28286 ( \33910 , \33546 );
buf \U$28287 ( \33911 , \33546 );
buf \U$28288 ( \33912 , \33546 );
buf \U$28289 ( \33913 , \33546 );
buf \U$28290 ( \33914 , \33546 );
buf \U$28291 ( \33915 , \33546 );
buf \U$28292 ( \33916 , \33546 );
buf \U$28293 ( \33917 , \33546 );
buf \U$28294 ( \33918 , \33546 );
buf \U$28295 ( \33919 , \33546 );
buf \U$28296 ( \33920 , \33546 );
buf \U$28297 ( \33921 , \33546 );
buf \U$28298 ( \33922 , \33546 );
buf \U$28299 ( \33923 , \33546 );
buf \U$28300 ( \33924 , \33546 );
buf \U$28301 ( \33925 , \33546 );
buf \U$28302 ( \33926 , \33546 );
nor \U$28303 ( \33927 , \33574 , \33575 , \33535 , \33536 , \33539 , \33543 , \33546 , \33902 , \33903 , \33904 , \33905 , \33906 , \33907 , \33908 , \33909 , \33910 , \33911 , \33912 , \33913 , \33914 , \33915 , \33916 , \33917 , \33918 , \33919 , \33920 , \33921 , \33922 , \33923 , \33924 , \33925 , \33926 );
and \U$28304 ( \33928 , RIeacfa18_6902, \33927 );
buf \U$28305 ( \33929 , \33546 );
buf \U$28306 ( \33930 , \33546 );
buf \U$28307 ( \33931 , \33546 );
buf \U$28308 ( \33932 , \33546 );
buf \U$28309 ( \33933 , \33546 );
buf \U$28310 ( \33934 , \33546 );
buf \U$28311 ( \33935 , \33546 );
buf \U$28312 ( \33936 , \33546 );
buf \U$28313 ( \33937 , \33546 );
buf \U$28314 ( \33938 , \33546 );
buf \U$28315 ( \33939 , \33546 );
buf \U$28316 ( \33940 , \33546 );
buf \U$28317 ( \33941 , \33546 );
buf \U$28318 ( \33942 , \33546 );
buf \U$28319 ( \33943 , \33546 );
buf \U$28320 ( \33944 , \33546 );
buf \U$28321 ( \33945 , \33546 );
buf \U$28322 ( \33946 , \33546 );
buf \U$28323 ( \33947 , \33546 );
buf \U$28324 ( \33948 , \33546 );
buf \U$28325 ( \33949 , \33546 );
buf \U$28326 ( \33950 , \33546 );
buf \U$28327 ( \33951 , \33546 );
buf \U$28328 ( \33952 , \33546 );
buf \U$28329 ( \33953 , \33546 );
nor \U$28330 ( \33954 , \33533 , \33575 , \33535 , \33536 , \33539 , \33543 , \33546 , \33929 , \33930 , \33931 , \33932 , \33933 , \33934 , \33935 , \33936 , \33937 , \33938 , \33939 , \33940 , \33941 , \33942 , \33943 , \33944 , \33945 , \33946 , \33947 , \33948 , \33949 , \33950 , \33951 , \33952 , \33953 );
and \U$28331 ( \33955 , RIeab6518_6891, \33954 );
buf \U$28332 ( \33956 , \33546 );
buf \U$28333 ( \33957 , \33546 );
buf \U$28334 ( \33958 , \33546 );
buf \U$28335 ( \33959 , \33546 );
buf \U$28336 ( \33960 , \33546 );
buf \U$28337 ( \33961 , \33546 );
buf \U$28338 ( \33962 , \33546 );
buf \U$28339 ( \33963 , \33546 );
buf \U$28340 ( \33964 , \33546 );
buf \U$28341 ( \33965 , \33546 );
buf \U$28342 ( \33966 , \33546 );
buf \U$28343 ( \33967 , \33546 );
buf \U$28344 ( \33968 , \33546 );
buf \U$28345 ( \33969 , \33546 );
buf \U$28346 ( \33970 , \33546 );
buf \U$28347 ( \33971 , \33546 );
buf \U$28348 ( \33972 , \33546 );
buf \U$28349 ( \33973 , \33546 );
buf \U$28350 ( \33974 , \33546 );
buf \U$28351 ( \33975 , \33546 );
buf \U$28352 ( \33976 , \33546 );
buf \U$28353 ( \33977 , \33546 );
buf \U$28354 ( \33978 , \33546 );
buf \U$28355 ( \33979 , \33546 );
buf \U$28356 ( \33980 , \33546 );
nor \U$28357 ( \33981 , \33574 , \33534 , \33535 , \33536 , \33539 , \33543 , \33546 , \33956 , \33957 , \33958 , \33959 , \33960 , \33961 , \33962 , \33963 , \33964 , \33965 , \33966 , \33967 , \33968 , \33969 , \33970 , \33971 , \33972 , \33973 , \33974 , \33975 , \33976 , \33977 , \33978 , \33979 , \33980 );
and \U$28358 ( \33982 , RIeb352c8_6904, \33981 );
or \U$28359 ( \33983 , \33573 , \33604 , \33631 , \33658 , \33685 , \33712 , \33739 , \33766 , \33793 , \33820 , \33847 , \33874 , \33901 , \33928 , \33955 , \33982 );
buf \U$28360 ( \33984 , \33546 );
not \U$28361 ( \33985 , \33984 );
buf \U$28362 ( \33986 , \33534 );
buf \U$28363 ( \33987 , \33535 );
buf \U$28364 ( \33988 , \33536 );
buf \U$28365 ( \33989 , \33539 );
buf \U$28366 ( \33990 , \33543 );
buf \U$28367 ( \33991 , \33546 );
buf \U$28368 ( \33992 , \33546 );
buf \U$28369 ( \33993 , \33546 );
buf \U$28370 ( \33994 , \33546 );
buf \U$28371 ( \33995 , \33546 );
buf \U$28372 ( \33996 , \33546 );
buf \U$28373 ( \33997 , \33546 );
buf \U$28374 ( \33998 , \33546 );
buf \U$28375 ( \33999 , \33546 );
buf \U$28376 ( \34000 , \33546 );
buf \U$28377 ( \34001 , \33546 );
buf \U$28378 ( \34002 , \33546 );
buf \U$28379 ( \34003 , \33546 );
buf \U$28380 ( \34004 , \33546 );
buf \U$28381 ( \34005 , \33546 );
buf \U$28382 ( \34006 , \33546 );
buf \U$28383 ( \34007 , \33546 );
buf \U$28384 ( \34008 , \33546 );
buf \U$28385 ( \34009 , \33546 );
buf \U$28386 ( \34010 , \33546 );
buf \U$28387 ( \34011 , \33546 );
buf \U$28388 ( \34012 , \33546 );
buf \U$28389 ( \34013 , \33546 );
buf \U$28390 ( \34014 , \33546 );
buf \U$28391 ( \34015 , \33546 );
buf \U$28392 ( \34016 , \33533 );
or \U$28393 ( \34017 , \33986 , \33987 , \33988 , \33989 , \33990 , \33991 , \33992 , \33993 , \33994 , \33995 , \33996 , \33997 , \33998 , \33999 , \34000 , \34001 , \34002 , \34003 , \34004 , \34005 , \34006 , \34007 , \34008 , \34009 , \34010 , \34011 , \34012 , \34013 , \34014 , \34015 , \34016 );
nand \U$28394 ( \34018 , \33985 , \34017 );
buf \U$28395 ( \34019 , \34018 );
buf \U$28396 ( \34020 , \33546 );
not \U$28397 ( \34021 , \34020 );
buf \U$28398 ( \34022 , \33543 );
buf \U$28399 ( \34023 , \33546 );
buf \U$28400 ( \34024 , \33546 );
buf \U$28401 ( \34025 , \33546 );
buf \U$28402 ( \34026 , \33546 );
buf \U$28403 ( \34027 , \33546 );
buf \U$28404 ( \34028 , \33546 );
buf \U$28405 ( \34029 , \33546 );
buf \U$28406 ( \34030 , \33546 );
buf \U$28407 ( \34031 , \33546 );
buf \U$28408 ( \34032 , \33546 );
buf \U$28409 ( \34033 , \33546 );
buf \U$28410 ( \34034 , \33546 );
buf \U$28411 ( \34035 , \33546 );
buf \U$28412 ( \34036 , \33546 );
buf \U$28413 ( \34037 , \33546 );
buf \U$28414 ( \34038 , \33546 );
buf \U$28415 ( \34039 , \33546 );
buf \U$28416 ( \34040 , \33546 );
buf \U$28417 ( \34041 , \33546 );
buf \U$28418 ( \34042 , \33546 );
buf \U$28419 ( \34043 , \33546 );
buf \U$28420 ( \34044 , \33546 );
buf \U$28421 ( \34045 , \33546 );
buf \U$28422 ( \34046 , \33546 );
buf \U$28423 ( \34047 , \33546 );
buf \U$28424 ( \34048 , \33539 );
buf \U$28425 ( \34049 , \33533 );
buf \U$28426 ( \34050 , \33534 );
buf \U$28427 ( \34051 , \33535 );
buf \U$28428 ( \34052 , \33536 );
or \U$28429 ( \34053 , \34049 , \34050 , \34051 , \34052 );
and \U$28430 ( \34054 , \34048 , \34053 );
or \U$28431 ( \34055 , \34022 , \34023 , \34024 , \34025 , \34026 , \34027 , \34028 , \34029 , \34030 , \34031 , \34032 , \34033 , \34034 , \34035 , \34036 , \34037 , \34038 , \34039 , \34040 , \34041 , \34042 , \34043 , \34044 , \34045 , \34046 , \34047 , \34054 );
and \U$28432 ( \34056 , \34021 , \34055 );
buf \U$28433 ( \34057 , \34056 );
or \U$28434 ( \34058 , \34019 , \34057 );
_DC g9c26 ( \34059_nG9c26 , \33983 , \34058 );
not \U$28435 ( \34060 , \34059_nG9c26 );
buf \U$28436 ( \34061 , RIb7b9608_246);
buf \U$28437 ( \34062 , \33546 );
buf \U$28438 ( \34063 , \33546 );
buf \U$28439 ( \34064 , \33546 );
buf \U$28440 ( \34065 , \33546 );
buf \U$28441 ( \34066 , \33546 );
buf \U$28442 ( \34067 , \33546 );
buf \U$28443 ( \34068 , \33546 );
buf \U$28444 ( \34069 , \33546 );
buf \U$28445 ( \34070 , \33546 );
buf \U$28446 ( \34071 , \33546 );
buf \U$28447 ( \34072 , \33546 );
buf \U$28448 ( \34073 , \33546 );
buf \U$28449 ( \34074 , \33546 );
buf \U$28450 ( \34075 , \33546 );
buf \U$28451 ( \34076 , \33546 );
buf \U$28452 ( \34077 , \33546 );
buf \U$28453 ( \34078 , \33546 );
buf \U$28454 ( \34079 , \33546 );
buf \U$28455 ( \34080 , \33546 );
buf \U$28456 ( \34081 , \33546 );
buf \U$28457 ( \34082 , \33546 );
buf \U$28458 ( \34083 , \33546 );
buf \U$28459 ( \34084 , \33546 );
buf \U$28460 ( \34085 , \33546 );
buf \U$28461 ( \34086 , \33546 );
nor \U$28462 ( \34087 , \33533 , \33534 , \33535 , \33536 , \33540 , \33543 , \33546 , \34062 , \34063 , \34064 , \34065 , \34066 , \34067 , \34068 , \34069 , \34070 , \34071 , \34072 , \34073 , \34074 , \34075 , \34076 , \34077 , \34078 , \34079 , \34080 , \34081 , \34082 , \34083 , \34084 , \34085 , \34086 );
and \U$28463 ( \34088 , \7117 , \34087 );
buf \U$28464 ( \34089 , \33546 );
buf \U$28465 ( \34090 , \33546 );
buf \U$28466 ( \34091 , \33546 );
buf \U$28467 ( \34092 , \33546 );
buf \U$28468 ( \34093 , \33546 );
buf \U$28469 ( \34094 , \33546 );
buf \U$28470 ( \34095 , \33546 );
buf \U$28471 ( \34096 , \33546 );
buf \U$28472 ( \34097 , \33546 );
buf \U$28473 ( \34098 , \33546 );
buf \U$28474 ( \34099 , \33546 );
buf \U$28475 ( \34100 , \33546 );
buf \U$28476 ( \34101 , \33546 );
buf \U$28477 ( \34102 , \33546 );
buf \U$28478 ( \34103 , \33546 );
buf \U$28479 ( \34104 , \33546 );
buf \U$28480 ( \34105 , \33546 );
buf \U$28481 ( \34106 , \33546 );
buf \U$28482 ( \34107 , \33546 );
buf \U$28483 ( \34108 , \33546 );
buf \U$28484 ( \34109 , \33546 );
buf \U$28485 ( \34110 , \33546 );
buf \U$28486 ( \34111 , \33546 );
buf \U$28487 ( \34112 , \33546 );
buf \U$28488 ( \34113 , \33546 );
nor \U$28489 ( \34114 , \33574 , \33575 , \33576 , \33577 , \33539 , \33543 , \33546 , \34089 , \34090 , \34091 , \34092 , \34093 , \34094 , \34095 , \34096 , \34097 , \34098 , \34099 , \34100 , \34101 , \34102 , \34103 , \34104 , \34105 , \34106 , \34107 , \34108 , \34109 , \34110 , \34111 , \34112 , \34113 );
and \U$28490 ( \34115 , \7119 , \34114 );
buf \U$28491 ( \34116 , \33546 );
buf \U$28492 ( \34117 , \33546 );
buf \U$28493 ( \34118 , \33546 );
buf \U$28494 ( \34119 , \33546 );
buf \U$28495 ( \34120 , \33546 );
buf \U$28496 ( \34121 , \33546 );
buf \U$28497 ( \34122 , \33546 );
buf \U$28498 ( \34123 , \33546 );
buf \U$28499 ( \34124 , \33546 );
buf \U$28500 ( \34125 , \33546 );
buf \U$28501 ( \34126 , \33546 );
buf \U$28502 ( \34127 , \33546 );
buf \U$28503 ( \34128 , \33546 );
buf \U$28504 ( \34129 , \33546 );
buf \U$28505 ( \34130 , \33546 );
buf \U$28506 ( \34131 , \33546 );
buf \U$28507 ( \34132 , \33546 );
buf \U$28508 ( \34133 , \33546 );
buf \U$28509 ( \34134 , \33546 );
buf \U$28510 ( \34135 , \33546 );
buf \U$28511 ( \34136 , \33546 );
buf \U$28512 ( \34137 , \33546 );
buf \U$28513 ( \34138 , \33546 );
buf \U$28514 ( \34139 , \33546 );
buf \U$28515 ( \34140 , \33546 );
nor \U$28516 ( \34141 , \33533 , \33575 , \33576 , \33577 , \33539 , \33543 , \33546 , \34116 , \34117 , \34118 , \34119 , \34120 , \34121 , \34122 , \34123 , \34124 , \34125 , \34126 , \34127 , \34128 , \34129 , \34130 , \34131 , \34132 , \34133 , \34134 , \34135 , \34136 , \34137 , \34138 , \34139 , \34140 );
and \U$28517 ( \34142 , \7864 , \34141 );
buf \U$28518 ( \34143 , \33546 );
buf \U$28519 ( \34144 , \33546 );
buf \U$28520 ( \34145 , \33546 );
buf \U$28521 ( \34146 , \33546 );
buf \U$28522 ( \34147 , \33546 );
buf \U$28523 ( \34148 , \33546 );
buf \U$28524 ( \34149 , \33546 );
buf \U$28525 ( \34150 , \33546 );
buf \U$28526 ( \34151 , \33546 );
buf \U$28527 ( \34152 , \33546 );
buf \U$28528 ( \34153 , \33546 );
buf \U$28529 ( \34154 , \33546 );
buf \U$28530 ( \34155 , \33546 );
buf \U$28531 ( \34156 , \33546 );
buf \U$28532 ( \34157 , \33546 );
buf \U$28533 ( \34158 , \33546 );
buf \U$28534 ( \34159 , \33546 );
buf \U$28535 ( \34160 , \33546 );
buf \U$28536 ( \34161 , \33546 );
buf \U$28537 ( \34162 , \33546 );
buf \U$28538 ( \34163 , \33546 );
buf \U$28539 ( \34164 , \33546 );
buf \U$28540 ( \34165 , \33546 );
buf \U$28541 ( \34166 , \33546 );
buf \U$28542 ( \34167 , \33546 );
nor \U$28543 ( \34168 , \33574 , \33534 , \33576 , \33577 , \33539 , \33543 , \33546 , \34143 , \34144 , \34145 , \34146 , \34147 , \34148 , \34149 , \34150 , \34151 , \34152 , \34153 , \34154 , \34155 , \34156 , \34157 , \34158 , \34159 , \34160 , \34161 , \34162 , \34163 , \34164 , \34165 , \34166 , \34167 );
and \U$28544 ( \34169 , \7892 , \34168 );
buf \U$28545 ( \34170 , \33546 );
buf \U$28546 ( \34171 , \33546 );
buf \U$28547 ( \34172 , \33546 );
buf \U$28548 ( \34173 , \33546 );
buf \U$28549 ( \34174 , \33546 );
buf \U$28550 ( \34175 , \33546 );
buf \U$28551 ( \34176 , \33546 );
buf \U$28552 ( \34177 , \33546 );
buf \U$28553 ( \34178 , \33546 );
buf \U$28554 ( \34179 , \33546 );
buf \U$28555 ( \34180 , \33546 );
buf \U$28556 ( \34181 , \33546 );
buf \U$28557 ( \34182 , \33546 );
buf \U$28558 ( \34183 , \33546 );
buf \U$28559 ( \34184 , \33546 );
buf \U$28560 ( \34185 , \33546 );
buf \U$28561 ( \34186 , \33546 );
buf \U$28562 ( \34187 , \33546 );
buf \U$28563 ( \34188 , \33546 );
buf \U$28564 ( \34189 , \33546 );
buf \U$28565 ( \34190 , \33546 );
buf \U$28566 ( \34191 , \33546 );
buf \U$28567 ( \34192 , \33546 );
buf \U$28568 ( \34193 , \33546 );
buf \U$28569 ( \34194 , \33546 );
nor \U$28570 ( \34195 , \33533 , \33534 , \33576 , \33577 , \33539 , \33543 , \33546 , \34170 , \34171 , \34172 , \34173 , \34174 , \34175 , \34176 , \34177 , \34178 , \34179 , \34180 , \34181 , \34182 , \34183 , \34184 , \34185 , \34186 , \34187 , \34188 , \34189 , \34190 , \34191 , \34192 , \34193 , \34194 );
and \U$28571 ( \34196 , \7920 , \34195 );
buf \U$28572 ( \34197 , \33546 );
buf \U$28573 ( \34198 , \33546 );
buf \U$28574 ( \34199 , \33546 );
buf \U$28575 ( \34200 , \33546 );
buf \U$28576 ( \34201 , \33546 );
buf \U$28577 ( \34202 , \33546 );
buf \U$28578 ( \34203 , \33546 );
buf \U$28579 ( \34204 , \33546 );
buf \U$28580 ( \34205 , \33546 );
buf \U$28581 ( \34206 , \33546 );
buf \U$28582 ( \34207 , \33546 );
buf \U$28583 ( \34208 , \33546 );
buf \U$28584 ( \34209 , \33546 );
buf \U$28585 ( \34210 , \33546 );
buf \U$28586 ( \34211 , \33546 );
buf \U$28587 ( \34212 , \33546 );
buf \U$28588 ( \34213 , \33546 );
buf \U$28589 ( \34214 , \33546 );
buf \U$28590 ( \34215 , \33546 );
buf \U$28591 ( \34216 , \33546 );
buf \U$28592 ( \34217 , \33546 );
buf \U$28593 ( \34218 , \33546 );
buf \U$28594 ( \34219 , \33546 );
buf \U$28595 ( \34220 , \33546 );
buf \U$28596 ( \34221 , \33546 );
nor \U$28597 ( \34222 , \33574 , \33575 , \33535 , \33577 , \33539 , \33543 , \33546 , \34197 , \34198 , \34199 , \34200 , \34201 , \34202 , \34203 , \34204 , \34205 , \34206 , \34207 , \34208 , \34209 , \34210 , \34211 , \34212 , \34213 , \34214 , \34215 , \34216 , \34217 , \34218 , \34219 , \34220 , \34221 );
and \U$28598 ( \34223 , \7948 , \34222 );
buf \U$28599 ( \34224 , \33546 );
buf \U$28600 ( \34225 , \33546 );
buf \U$28601 ( \34226 , \33546 );
buf \U$28602 ( \34227 , \33546 );
buf \U$28603 ( \34228 , \33546 );
buf \U$28604 ( \34229 , \33546 );
buf \U$28605 ( \34230 , \33546 );
buf \U$28606 ( \34231 , \33546 );
buf \U$28607 ( \34232 , \33546 );
buf \U$28608 ( \34233 , \33546 );
buf \U$28609 ( \34234 , \33546 );
buf \U$28610 ( \34235 , \33546 );
buf \U$28611 ( \34236 , \33546 );
buf \U$28612 ( \34237 , \33546 );
buf \U$28613 ( \34238 , \33546 );
buf \U$28614 ( \34239 , \33546 );
buf \U$28615 ( \34240 , \33546 );
buf \U$28616 ( \34241 , \33546 );
buf \U$28617 ( \34242 , \33546 );
buf \U$28618 ( \34243 , \33546 );
buf \U$28619 ( \34244 , \33546 );
buf \U$28620 ( \34245 , \33546 );
buf \U$28621 ( \34246 , \33546 );
buf \U$28622 ( \34247 , \33546 );
buf \U$28623 ( \34248 , \33546 );
nor \U$28624 ( \34249 , \33533 , \33575 , \33535 , \33577 , \33539 , \33543 , \33546 , \34224 , \34225 , \34226 , \34227 , \34228 , \34229 , \34230 , \34231 , \34232 , \34233 , \34234 , \34235 , \34236 , \34237 , \34238 , \34239 , \34240 , \34241 , \34242 , \34243 , \34244 , \34245 , \34246 , \34247 , \34248 );
and \U$28625 ( \34250 , \7976 , \34249 );
buf \U$28626 ( \34251 , \33546 );
buf \U$28627 ( \34252 , \33546 );
buf \U$28628 ( \34253 , \33546 );
buf \U$28629 ( \34254 , \33546 );
buf \U$28630 ( \34255 , \33546 );
buf \U$28631 ( \34256 , \33546 );
buf \U$28632 ( \34257 , \33546 );
buf \U$28633 ( \34258 , \33546 );
buf \U$28634 ( \34259 , \33546 );
buf \U$28635 ( \34260 , \33546 );
buf \U$28636 ( \34261 , \33546 );
buf \U$28637 ( \34262 , \33546 );
buf \U$28638 ( \34263 , \33546 );
buf \U$28639 ( \34264 , \33546 );
buf \U$28640 ( \34265 , \33546 );
buf \U$28641 ( \34266 , \33546 );
buf \U$28642 ( \34267 , \33546 );
buf \U$28643 ( \34268 , \33546 );
buf \U$28644 ( \34269 , \33546 );
buf \U$28645 ( \34270 , \33546 );
buf \U$28646 ( \34271 , \33546 );
buf \U$28647 ( \34272 , \33546 );
buf \U$28648 ( \34273 , \33546 );
buf \U$28649 ( \34274 , \33546 );
buf \U$28650 ( \34275 , \33546 );
nor \U$28651 ( \34276 , \33574 , \33534 , \33535 , \33577 , \33539 , \33543 , \33546 , \34251 , \34252 , \34253 , \34254 , \34255 , \34256 , \34257 , \34258 , \34259 , \34260 , \34261 , \34262 , \34263 , \34264 , \34265 , \34266 , \34267 , \34268 , \34269 , \34270 , \34271 , \34272 , \34273 , \34274 , \34275 );
and \U$28652 ( \34277 , \8004 , \34276 );
buf \U$28653 ( \34278 , \33546 );
buf \U$28654 ( \34279 , \33546 );
buf \U$28655 ( \34280 , \33546 );
buf \U$28656 ( \34281 , \33546 );
buf \U$28657 ( \34282 , \33546 );
buf \U$28658 ( \34283 , \33546 );
buf \U$28659 ( \34284 , \33546 );
buf \U$28660 ( \34285 , \33546 );
buf \U$28661 ( \34286 , \33546 );
buf \U$28662 ( \34287 , \33546 );
buf \U$28663 ( \34288 , \33546 );
buf \U$28664 ( \34289 , \33546 );
buf \U$28665 ( \34290 , \33546 );
buf \U$28666 ( \34291 , \33546 );
buf \U$28667 ( \34292 , \33546 );
buf \U$28668 ( \34293 , \33546 );
buf \U$28669 ( \34294 , \33546 );
buf \U$28670 ( \34295 , \33546 );
buf \U$28671 ( \34296 , \33546 );
buf \U$28672 ( \34297 , \33546 );
buf \U$28673 ( \34298 , \33546 );
buf \U$28674 ( \34299 , \33546 );
buf \U$28675 ( \34300 , \33546 );
buf \U$28676 ( \34301 , \33546 );
buf \U$28677 ( \34302 , \33546 );
nor \U$28678 ( \34303 , \33533 , \33534 , \33535 , \33577 , \33539 , \33543 , \33546 , \34278 , \34279 , \34280 , \34281 , \34282 , \34283 , \34284 , \34285 , \34286 , \34287 , \34288 , \34289 , \34290 , \34291 , \34292 , \34293 , \34294 , \34295 , \34296 , \34297 , \34298 , \34299 , \34300 , \34301 , \34302 );
and \U$28679 ( \34304 , \8032 , \34303 );
buf \U$28680 ( \34305 , \33546 );
buf \U$28681 ( \34306 , \33546 );
buf \U$28682 ( \34307 , \33546 );
buf \U$28683 ( \34308 , \33546 );
buf \U$28684 ( \34309 , \33546 );
buf \U$28685 ( \34310 , \33546 );
buf \U$28686 ( \34311 , \33546 );
buf \U$28687 ( \34312 , \33546 );
buf \U$28688 ( \34313 , \33546 );
buf \U$28689 ( \34314 , \33546 );
buf \U$28690 ( \34315 , \33546 );
buf \U$28691 ( \34316 , \33546 );
buf \U$28692 ( \34317 , \33546 );
buf \U$28693 ( \34318 , \33546 );
buf \U$28694 ( \34319 , \33546 );
buf \U$28695 ( \34320 , \33546 );
buf \U$28696 ( \34321 , \33546 );
buf \U$28697 ( \34322 , \33546 );
buf \U$28698 ( \34323 , \33546 );
buf \U$28699 ( \34324 , \33546 );
buf \U$28700 ( \34325 , \33546 );
buf \U$28701 ( \34326 , \33546 );
buf \U$28702 ( \34327 , \33546 );
buf \U$28703 ( \34328 , \33546 );
buf \U$28704 ( \34329 , \33546 );
nor \U$28705 ( \34330 , \33574 , \33575 , \33576 , \33536 , \33539 , \33543 , \33546 , \34305 , \34306 , \34307 , \34308 , \34309 , \34310 , \34311 , \34312 , \34313 , \34314 , \34315 , \34316 , \34317 , \34318 , \34319 , \34320 , \34321 , \34322 , \34323 , \34324 , \34325 , \34326 , \34327 , \34328 , \34329 );
and \U$28706 ( \34331 , \8060 , \34330 );
buf \U$28707 ( \34332 , \33546 );
buf \U$28708 ( \34333 , \33546 );
buf \U$28709 ( \34334 , \33546 );
buf \U$28710 ( \34335 , \33546 );
buf \U$28711 ( \34336 , \33546 );
buf \U$28712 ( \34337 , \33546 );
buf \U$28713 ( \34338 , \33546 );
buf \U$28714 ( \34339 , \33546 );
buf \U$28715 ( \34340 , \33546 );
buf \U$28716 ( \34341 , \33546 );
buf \U$28717 ( \34342 , \33546 );
buf \U$28718 ( \34343 , \33546 );
buf \U$28719 ( \34344 , \33546 );
buf \U$28720 ( \34345 , \33546 );
buf \U$28721 ( \34346 , \33546 );
buf \U$28722 ( \34347 , \33546 );
buf \U$28723 ( \34348 , \33546 );
buf \U$28724 ( \34349 , \33546 );
buf \U$28725 ( \34350 , \33546 );
buf \U$28726 ( \34351 , \33546 );
buf \U$28727 ( \34352 , \33546 );
buf \U$28728 ( \34353 , \33546 );
buf \U$28729 ( \34354 , \33546 );
buf \U$28730 ( \34355 , \33546 );
buf \U$28731 ( \34356 , \33546 );
nor \U$28732 ( \34357 , \33533 , \33575 , \33576 , \33536 , \33539 , \33543 , \33546 , \34332 , \34333 , \34334 , \34335 , \34336 , \34337 , \34338 , \34339 , \34340 , \34341 , \34342 , \34343 , \34344 , \34345 , \34346 , \34347 , \34348 , \34349 , \34350 , \34351 , \34352 , \34353 , \34354 , \34355 , \34356 );
and \U$28733 ( \34358 , \8088 , \34357 );
buf \U$28734 ( \34359 , \33546 );
buf \U$28735 ( \34360 , \33546 );
buf \U$28736 ( \34361 , \33546 );
buf \U$28737 ( \34362 , \33546 );
buf \U$28738 ( \34363 , \33546 );
buf \U$28739 ( \34364 , \33546 );
buf \U$28740 ( \34365 , \33546 );
buf \U$28741 ( \34366 , \33546 );
buf \U$28742 ( \34367 , \33546 );
buf \U$28743 ( \34368 , \33546 );
buf \U$28744 ( \34369 , \33546 );
buf \U$28745 ( \34370 , \33546 );
buf \U$28746 ( \34371 , \33546 );
buf \U$28747 ( \34372 , \33546 );
buf \U$28748 ( \34373 , \33546 );
buf \U$28749 ( \34374 , \33546 );
buf \U$28750 ( \34375 , \33546 );
buf \U$28751 ( \34376 , \33546 );
buf \U$28752 ( \34377 , \33546 );
buf \U$28753 ( \34378 , \33546 );
buf \U$28754 ( \34379 , \33546 );
buf \U$28755 ( \34380 , \33546 );
buf \U$28756 ( \34381 , \33546 );
buf \U$28757 ( \34382 , \33546 );
buf \U$28758 ( \34383 , \33546 );
nor \U$28759 ( \34384 , \33574 , \33534 , \33576 , \33536 , \33539 , \33543 , \33546 , \34359 , \34360 , \34361 , \34362 , \34363 , \34364 , \34365 , \34366 , \34367 , \34368 , \34369 , \34370 , \34371 , \34372 , \34373 , \34374 , \34375 , \34376 , \34377 , \34378 , \34379 , \34380 , \34381 , \34382 , \34383 );
and \U$28760 ( \34385 , \8116 , \34384 );
buf \U$28761 ( \34386 , \33546 );
buf \U$28762 ( \34387 , \33546 );
buf \U$28763 ( \34388 , \33546 );
buf \U$28764 ( \34389 , \33546 );
buf \U$28765 ( \34390 , \33546 );
buf \U$28766 ( \34391 , \33546 );
buf \U$28767 ( \34392 , \33546 );
buf \U$28768 ( \34393 , \33546 );
buf \U$28769 ( \34394 , \33546 );
buf \U$28770 ( \34395 , \33546 );
buf \U$28771 ( \34396 , \33546 );
buf \U$28772 ( \34397 , \33546 );
buf \U$28773 ( \34398 , \33546 );
buf \U$28774 ( \34399 , \33546 );
buf \U$28775 ( \34400 , \33546 );
buf \U$28776 ( \34401 , \33546 );
buf \U$28777 ( \34402 , \33546 );
buf \U$28778 ( \34403 , \33546 );
buf \U$28779 ( \34404 , \33546 );
buf \U$28780 ( \34405 , \33546 );
buf \U$28781 ( \34406 , \33546 );
buf \U$28782 ( \34407 , \33546 );
buf \U$28783 ( \34408 , \33546 );
buf \U$28784 ( \34409 , \33546 );
buf \U$28785 ( \34410 , \33546 );
nor \U$28786 ( \34411 , \33533 , \33534 , \33576 , \33536 , \33539 , \33543 , \33546 , \34386 , \34387 , \34388 , \34389 , \34390 , \34391 , \34392 , \34393 , \34394 , \34395 , \34396 , \34397 , \34398 , \34399 , \34400 , \34401 , \34402 , \34403 , \34404 , \34405 , \34406 , \34407 , \34408 , \34409 , \34410 );
and \U$28787 ( \34412 , \8144 , \34411 );
buf \U$28788 ( \34413 , \33546 );
buf \U$28789 ( \34414 , \33546 );
buf \U$28790 ( \34415 , \33546 );
buf \U$28791 ( \34416 , \33546 );
buf \U$28792 ( \34417 , \33546 );
buf \U$28793 ( \34418 , \33546 );
buf \U$28794 ( \34419 , \33546 );
buf \U$28795 ( \34420 , \33546 );
buf \U$28796 ( \34421 , \33546 );
buf \U$28797 ( \34422 , \33546 );
buf \U$28798 ( \34423 , \33546 );
buf \U$28799 ( \34424 , \33546 );
buf \U$28800 ( \34425 , \33546 );
buf \U$28801 ( \34426 , \33546 );
buf \U$28802 ( \34427 , \33546 );
buf \U$28803 ( \34428 , \33546 );
buf \U$28804 ( \34429 , \33546 );
buf \U$28805 ( \34430 , \33546 );
buf \U$28806 ( \34431 , \33546 );
buf \U$28807 ( \34432 , \33546 );
buf \U$28808 ( \34433 , \33546 );
buf \U$28809 ( \34434 , \33546 );
buf \U$28810 ( \34435 , \33546 );
buf \U$28811 ( \34436 , \33546 );
buf \U$28812 ( \34437 , \33546 );
nor \U$28813 ( \34438 , \33574 , \33575 , \33535 , \33536 , \33539 , \33543 , \33546 , \34413 , \34414 , \34415 , \34416 , \34417 , \34418 , \34419 , \34420 , \34421 , \34422 , \34423 , \34424 , \34425 , \34426 , \34427 , \34428 , \34429 , \34430 , \34431 , \34432 , \34433 , \34434 , \34435 , \34436 , \34437 );
and \U$28814 ( \34439 , \8172 , \34438 );
buf \U$28815 ( \34440 , \33546 );
buf \U$28816 ( \34441 , \33546 );
buf \U$28817 ( \34442 , \33546 );
buf \U$28818 ( \34443 , \33546 );
buf \U$28819 ( \34444 , \33546 );
buf \U$28820 ( \34445 , \33546 );
buf \U$28821 ( \34446 , \33546 );
buf \U$28822 ( \34447 , \33546 );
buf \U$28823 ( \34448 , \33546 );
buf \U$28824 ( \34449 , \33546 );
buf \U$28825 ( \34450 , \33546 );
buf \U$28826 ( \34451 , \33546 );
buf \U$28827 ( \34452 , \33546 );
buf \U$28828 ( \34453 , \33546 );
buf \U$28829 ( \34454 , \33546 );
buf \U$28830 ( \34455 , \33546 );
buf \U$28831 ( \34456 , \33546 );
buf \U$28832 ( \34457 , \33546 );
buf \U$28833 ( \34458 , \33546 );
buf \U$28834 ( \34459 , \33546 );
buf \U$28835 ( \34460 , \33546 );
buf \U$28836 ( \34461 , \33546 );
buf \U$28837 ( \34462 , \33546 );
buf \U$28838 ( \34463 , \33546 );
buf \U$28839 ( \34464 , \33546 );
nor \U$28840 ( \34465 , \33533 , \33575 , \33535 , \33536 , \33539 , \33543 , \33546 , \34440 , \34441 , \34442 , \34443 , \34444 , \34445 , \34446 , \34447 , \34448 , \34449 , \34450 , \34451 , \34452 , \34453 , \34454 , \34455 , \34456 , \34457 , \34458 , \34459 , \34460 , \34461 , \34462 , \34463 , \34464 );
and \U$28841 ( \34466 , \8200 , \34465 );
buf \U$28842 ( \34467 , \33546 );
buf \U$28843 ( \34468 , \33546 );
buf \U$28844 ( \34469 , \33546 );
buf \U$28845 ( \34470 , \33546 );
buf \U$28846 ( \34471 , \33546 );
buf \U$28847 ( \34472 , \33546 );
buf \U$28848 ( \34473 , \33546 );
buf \U$28849 ( \34474 , \33546 );
buf \U$28850 ( \34475 , \33546 );
buf \U$28851 ( \34476 , \33546 );
buf \U$28852 ( \34477 , \33546 );
buf \U$28853 ( \34478 , \33546 );
buf \U$28854 ( \34479 , \33546 );
buf \U$28855 ( \34480 , \33546 );
buf \U$28856 ( \34481 , \33546 );
buf \U$28857 ( \34482 , \33546 );
buf \U$28858 ( \34483 , \33546 );
buf \U$28859 ( \34484 , \33546 );
buf \U$28860 ( \34485 , \33546 );
buf \U$28861 ( \34486 , \33546 );
buf \U$28862 ( \34487 , \33546 );
buf \U$28863 ( \34488 , \33546 );
buf \U$28864 ( \34489 , \33546 );
buf \U$28865 ( \34490 , \33546 );
buf \U$28866 ( \34491 , \33546 );
nor \U$28867 ( \34492 , \33574 , \33534 , \33535 , \33536 , \33539 , \33543 , \33546 , \34467 , \34468 , \34469 , \34470 , \34471 , \34472 , \34473 , \34474 , \34475 , \34476 , \34477 , \34478 , \34479 , \34480 , \34481 , \34482 , \34483 , \34484 , \34485 , \34486 , \34487 , \34488 , \34489 , \34490 , \34491 );
and \U$28868 ( \34493 , \8228 , \34492 );
or \U$28869 ( \34494 , \34088 , \34115 , \34142 , \34169 , \34196 , \34223 , \34250 , \34277 , \34304 , \34331 , \34358 , \34385 , \34412 , \34439 , \34466 , \34493 );
buf \U$28870 ( \34495 , \33546 );
not \U$28871 ( \34496 , \34495 );
buf \U$28872 ( \34497 , \33534 );
buf \U$28873 ( \34498 , \33535 );
buf \U$28874 ( \34499 , \33536 );
buf \U$28875 ( \34500 , \33539 );
buf \U$28876 ( \34501 , \33543 );
buf \U$28877 ( \34502 , \33546 );
buf \U$28878 ( \34503 , \33546 );
buf \U$28879 ( \34504 , \33546 );
buf \U$28880 ( \34505 , \33546 );
buf \U$28881 ( \34506 , \33546 );
buf \U$28882 ( \34507 , \33546 );
buf \U$28883 ( \34508 , \33546 );
buf \U$28884 ( \34509 , \33546 );
buf \U$28885 ( \34510 , \33546 );
buf \U$28886 ( \34511 , \33546 );
buf \U$28887 ( \34512 , \33546 );
buf \U$28888 ( \34513 , \33546 );
buf \U$28889 ( \34514 , \33546 );
buf \U$28890 ( \34515 , \33546 );
buf \U$28891 ( \34516 , \33546 );
buf \U$28892 ( \34517 , \33546 );
buf \U$28893 ( \34518 , \33546 );
buf \U$28894 ( \34519 , \33546 );
buf \U$28895 ( \34520 , \33546 );
buf \U$28896 ( \34521 , \33546 );
buf \U$28897 ( \34522 , \33546 );
buf \U$28898 ( \34523 , \33546 );
buf \U$28899 ( \34524 , \33546 );
buf \U$28900 ( \34525 , \33546 );
buf \U$28901 ( \34526 , \33546 );
buf \U$28902 ( \34527 , \33533 );
or \U$28903 ( \34528 , \34497 , \34498 , \34499 , \34500 , \34501 , \34502 , \34503 , \34504 , \34505 , \34506 , \34507 , \34508 , \34509 , \34510 , \34511 , \34512 , \34513 , \34514 , \34515 , \34516 , \34517 , \34518 , \34519 , \34520 , \34521 , \34522 , \34523 , \34524 , \34525 , \34526 , \34527 );
nand \U$28904 ( \34529 , \34496 , \34528 );
buf \U$28905 ( \34530 , \34529 );
buf \U$28906 ( \34531 , \33546 );
not \U$28907 ( \34532 , \34531 );
buf \U$28908 ( \34533 , \33543 );
buf \U$28909 ( \34534 , \33546 );
buf \U$28910 ( \34535 , \33546 );
buf \U$28911 ( \34536 , \33546 );
buf \U$28912 ( \34537 , \33546 );
buf \U$28913 ( \34538 , \33546 );
buf \U$28914 ( \34539 , \33546 );
buf \U$28915 ( \34540 , \33546 );
buf \U$28916 ( \34541 , \33546 );
buf \U$28917 ( \34542 , \33546 );
buf \U$28918 ( \34543 , \33546 );
buf \U$28919 ( \34544 , \33546 );
buf \U$28920 ( \34545 , \33546 );
buf \U$28921 ( \34546 , \33546 );
buf \U$28922 ( \34547 , \33546 );
buf \U$28923 ( \34548 , \33546 );
buf \U$28924 ( \34549 , \33546 );
buf \U$28925 ( \34550 , \33546 );
buf \U$28926 ( \34551 , \33546 );
buf \U$28927 ( \34552 , \33546 );
buf \U$28928 ( \34553 , \33546 );
buf \U$28929 ( \34554 , \33546 );
buf \U$28930 ( \34555 , \33546 );
buf \U$28931 ( \34556 , \33546 );
buf \U$28932 ( \34557 , \33546 );
buf \U$28933 ( \34558 , \33546 );
buf \U$28934 ( \34559 , \33539 );
buf \U$28935 ( \34560 , \33533 );
buf \U$28936 ( \34561 , \33534 );
buf \U$28937 ( \34562 , \33535 );
buf \U$28938 ( \34563 , \33536 );
or \U$28939 ( \34564 , \34560 , \34561 , \34562 , \34563 );
and \U$28940 ( \34565 , \34559 , \34564 );
or \U$28941 ( \34566 , \34533 , \34534 , \34535 , \34536 , \34537 , \34538 , \34539 , \34540 , \34541 , \34542 , \34543 , \34544 , \34545 , \34546 , \34547 , \34548 , \34549 , \34550 , \34551 , \34552 , \34553 , \34554 , \34555 , \34556 , \34557 , \34558 , \34565 );
and \U$28942 ( \34567 , \34532 , \34566 );
buf \U$28943 ( \34568 , \34567 );
or \U$28944 ( \34569 , \34530 , \34568 );
_DC g9e25 ( \34570_nG9e25 , \34494 , \34569 );
buf \U$28945 ( \34571 , \34570_nG9e25 );
xor \U$28946 ( \34572 , \34061 , \34571 );
buf \U$28947 ( \34573 , RIb7b9590_247);
and \U$28948 ( \34574 , \7126 , \34087 );
and \U$28949 ( \34575 , \7128 , \34114 );
and \U$28950 ( \34576 , \8338 , \34141 );
and \U$28951 ( \34577 , \8340 , \34168 );
and \U$28952 ( \34578 , \8342 , \34195 );
and \U$28953 ( \34579 , \8344 , \34222 );
and \U$28954 ( \34580 , \8346 , \34249 );
and \U$28955 ( \34581 , \8348 , \34276 );
and \U$28956 ( \34582 , \8350 , \34303 );
and \U$28957 ( \34583 , \8352 , \34330 );
and \U$28958 ( \34584 , \8354 , \34357 );
and \U$28959 ( \34585 , \8356 , \34384 );
and \U$28960 ( \34586 , \8358 , \34411 );
and \U$28961 ( \34587 , \8360 , \34438 );
and \U$28962 ( \34588 , \8362 , \34465 );
and \U$28963 ( \34589 , \8364 , \34492 );
or \U$28964 ( \34590 , \34574 , \34575 , \34576 , \34577 , \34578 , \34579 , \34580 , \34581 , \34582 , \34583 , \34584 , \34585 , \34586 , \34587 , \34588 , \34589 );
_DC g9e3a ( \34591_nG9e3a , \34590 , \34569 );
buf \U$28965 ( \34592 , \34591_nG9e3a );
xor \U$28966 ( \34593 , \34573 , \34592 );
or \U$28967 ( \34594 , \34572 , \34593 );
buf \U$28968 ( \34595 , RIb7b9518_248);
and \U$28969 ( \34596 , \7136 , \34087 );
and \U$28970 ( \34597 , \7138 , \34114 );
and \U$28971 ( \34598 , \8374 , \34141 );
and \U$28972 ( \34599 , \8376 , \34168 );
and \U$28973 ( \34600 , \8378 , \34195 );
and \U$28974 ( \34601 , \8380 , \34222 );
and \U$28975 ( \34602 , \8382 , \34249 );
and \U$28976 ( \34603 , \8384 , \34276 );
and \U$28977 ( \34604 , \8386 , \34303 );
and \U$28978 ( \34605 , \8388 , \34330 );
and \U$28979 ( \34606 , \8390 , \34357 );
and \U$28980 ( \34607 , \8392 , \34384 );
and \U$28981 ( \34608 , \8394 , \34411 );
and \U$28982 ( \34609 , \8396 , \34438 );
and \U$28983 ( \34610 , \8398 , \34465 );
and \U$28984 ( \34611 , \8400 , \34492 );
or \U$28985 ( \34612 , \34596 , \34597 , \34598 , \34599 , \34600 , \34601 , \34602 , \34603 , \34604 , \34605 , \34606 , \34607 , \34608 , \34609 , \34610 , \34611 );
_DC g9e50 ( \34613_nG9e50 , \34612 , \34569 );
buf \U$28986 ( \34614 , \34613_nG9e50 );
xor \U$28987 ( \34615 , \34595 , \34614 );
or \U$28988 ( \34616 , \34594 , \34615 );
buf \U$28989 ( \34617 , RIb7b94a0_249);
and \U$28990 ( \34618 , \7146 , \34087 );
and \U$28991 ( \34619 , \7148 , \34114 );
and \U$28992 ( \34620 , \8410 , \34141 );
and \U$28993 ( \34621 , \8412 , \34168 );
and \U$28994 ( \34622 , \8414 , \34195 );
and \U$28995 ( \34623 , \8416 , \34222 );
and \U$28996 ( \34624 , \8418 , \34249 );
and \U$28997 ( \34625 , \8420 , \34276 );
and \U$28998 ( \34626 , \8422 , \34303 );
and \U$28999 ( \34627 , \8424 , \34330 );
and \U$29000 ( \34628 , \8426 , \34357 );
and \U$29001 ( \34629 , \8428 , \34384 );
and \U$29002 ( \34630 , \8430 , \34411 );
and \U$29003 ( \34631 , \8432 , \34438 );
and \U$29004 ( \34632 , \8434 , \34465 );
and \U$29005 ( \34633 , \8436 , \34492 );
or \U$29006 ( \34634 , \34618 , \34619 , \34620 , \34621 , \34622 , \34623 , \34624 , \34625 , \34626 , \34627 , \34628 , \34629 , \34630 , \34631 , \34632 , \34633 );
_DC g9e66 ( \34635_nG9e66 , \34634 , \34569 );
buf \U$29007 ( \34636 , \34635_nG9e66 );
xor \U$29008 ( \34637 , \34617 , \34636 );
or \U$29009 ( \34638 , \34616 , \34637 );
buf \U$29010 ( \34639 , RIb7b9428_250);
and \U$29011 ( \34640 , \7156 , \34087 );
and \U$29012 ( \34641 , \7158 , \34114 );
and \U$29013 ( \34642 , \8446 , \34141 );
and \U$29014 ( \34643 , \8448 , \34168 );
and \U$29015 ( \34644 , \8450 , \34195 );
and \U$29016 ( \34645 , \8452 , \34222 );
and \U$29017 ( \34646 , \8454 , \34249 );
and \U$29018 ( \34647 , \8456 , \34276 );
and \U$29019 ( \34648 , \8458 , \34303 );
and \U$29020 ( \34649 , \8460 , \34330 );
and \U$29021 ( \34650 , \8462 , \34357 );
and \U$29022 ( \34651 , \8464 , \34384 );
and \U$29023 ( \34652 , \8466 , \34411 );
and \U$29024 ( \34653 , \8468 , \34438 );
and \U$29025 ( \34654 , \8470 , \34465 );
and \U$29026 ( \34655 , \8472 , \34492 );
or \U$29027 ( \34656 , \34640 , \34641 , \34642 , \34643 , \34644 , \34645 , \34646 , \34647 , \34648 , \34649 , \34650 , \34651 , \34652 , \34653 , \34654 , \34655 );
_DC g9e7c ( \34657_nG9e7c , \34656 , \34569 );
buf \U$29028 ( \34658 , \34657_nG9e7c );
xor \U$29029 ( \34659 , \34639 , \34658 );
or \U$29030 ( \34660 , \34638 , \34659 );
buf \U$29031 ( \34661 , RIb7b93b0_251);
and \U$29032 ( \34662 , \7166 , \34087 );
and \U$29033 ( \34663 , \7168 , \34114 );
and \U$29034 ( \34664 , \8482 , \34141 );
and \U$29035 ( \34665 , \8484 , \34168 );
and \U$29036 ( \34666 , \8486 , \34195 );
and \U$29037 ( \34667 , \8488 , \34222 );
and \U$29038 ( \34668 , \8490 , \34249 );
and \U$29039 ( \34669 , \8492 , \34276 );
and \U$29040 ( \34670 , \8494 , \34303 );
and \U$29041 ( \34671 , \8496 , \34330 );
and \U$29042 ( \34672 , \8498 , \34357 );
and \U$29043 ( \34673 , \8500 , \34384 );
and \U$29044 ( \34674 , \8502 , \34411 );
and \U$29045 ( \34675 , \8504 , \34438 );
and \U$29046 ( \34676 , \8506 , \34465 );
and \U$29047 ( \34677 , \8508 , \34492 );
or \U$29048 ( \34678 , \34662 , \34663 , \34664 , \34665 , \34666 , \34667 , \34668 , \34669 , \34670 , \34671 , \34672 , \34673 , \34674 , \34675 , \34676 , \34677 );
_DC g9e92 ( \34679_nG9e92 , \34678 , \34569 );
buf \U$29049 ( \34680 , \34679_nG9e92 );
xor \U$29050 ( \34681 , \34661 , \34680 );
or \U$29051 ( \34682 , \34660 , \34681 );
buf \U$29052 ( \34683 , RIb7af720_252);
and \U$29053 ( \34684 , \7176 , \34087 );
and \U$29054 ( \34685 , \7178 , \34114 );
and \U$29055 ( \34686 , \8518 , \34141 );
and \U$29056 ( \34687 , \8520 , \34168 );
and \U$29057 ( \34688 , \8522 , \34195 );
and \U$29058 ( \34689 , \8524 , \34222 );
and \U$29059 ( \34690 , \8526 , \34249 );
and \U$29060 ( \34691 , \8528 , \34276 );
and \U$29061 ( \34692 , \8530 , \34303 );
and \U$29062 ( \34693 , \8532 , \34330 );
and \U$29063 ( \34694 , \8534 , \34357 );
and \U$29064 ( \34695 , \8536 , \34384 );
and \U$29065 ( \34696 , \8538 , \34411 );
and \U$29066 ( \34697 , \8540 , \34438 );
and \U$29067 ( \34698 , \8542 , \34465 );
and \U$29068 ( \34699 , \8544 , \34492 );
or \U$29069 ( \34700 , \34684 , \34685 , \34686 , \34687 , \34688 , \34689 , \34690 , \34691 , \34692 , \34693 , \34694 , \34695 , \34696 , \34697 , \34698 , \34699 );
_DC g9ea8 ( \34701_nG9ea8 , \34700 , \34569 );
buf \U$29070 ( \34702 , \34701_nG9ea8 );
xor \U$29071 ( \34703 , \34683 , \34702 );
or \U$29072 ( \34704 , \34682 , \34703 );
buf \U$29073 ( \34705 , RIb7af6a8_253);
and \U$29074 ( \34706 , \7186 , \34087 );
and \U$29075 ( \34707 , \7188 , \34114 );
and \U$29076 ( \34708 , \8554 , \34141 );
and \U$29077 ( \34709 , \8556 , \34168 );
and \U$29078 ( \34710 , \8558 , \34195 );
and \U$29079 ( \34711 , \8560 , \34222 );
and \U$29080 ( \34712 , \8562 , \34249 );
and \U$29081 ( \34713 , \8564 , \34276 );
and \U$29082 ( \34714 , \8566 , \34303 );
and \U$29083 ( \34715 , \8568 , \34330 );
and \U$29084 ( \34716 , \8570 , \34357 );
and \U$29085 ( \34717 , \8572 , \34384 );
and \U$29086 ( \34718 , \8574 , \34411 );
and \U$29087 ( \34719 , \8576 , \34438 );
and \U$29088 ( \34720 , \8578 , \34465 );
and \U$29089 ( \34721 , \8580 , \34492 );
or \U$29090 ( \34722 , \34706 , \34707 , \34708 , \34709 , \34710 , \34711 , \34712 , \34713 , \34714 , \34715 , \34716 , \34717 , \34718 , \34719 , \34720 , \34721 );
_DC g9ebe ( \34723_nG9ebe , \34722 , \34569 );
buf \U$29091 ( \34724 , \34723_nG9ebe );
xor \U$29092 ( \34725 , \34705 , \34724 );
or \U$29093 ( \34726 , \34704 , \34725 );
not \U$29094 ( \34727 , \34726 );
buf \U$29095 ( \34728 , \34727 );
and \U$29096 ( \34729 , \34060 , \34728 );
buf \U$29097 ( \34730 , RIb7af630_254);
buf \U$29098 ( \34731 , \33546 );
buf \U$29099 ( \34732 , \33546 );
buf \U$29100 ( \34733 , \33546 );
buf \U$29101 ( \34734 , \33546 );
buf \U$29102 ( \34735 , \33546 );
buf \U$29103 ( \34736 , \33546 );
buf \U$29104 ( \34737 , \33546 );
buf \U$29105 ( \34738 , \33546 );
buf \U$29106 ( \34739 , \33546 );
buf \U$29107 ( \34740 , \33546 );
buf \U$29108 ( \34741 , \33546 );
buf \U$29109 ( \34742 , \33546 );
buf \U$29110 ( \34743 , \33546 );
buf \U$29111 ( \34744 , \33546 );
buf \U$29112 ( \34745 , \33546 );
buf \U$29113 ( \34746 , \33546 );
buf \U$29114 ( \34747 , \33546 );
buf \U$29115 ( \34748 , \33546 );
buf \U$29116 ( \34749 , \33546 );
buf \U$29117 ( \34750 , \33546 );
buf \U$29118 ( \34751 , \33546 );
buf \U$29119 ( \34752 , \33546 );
buf \U$29120 ( \34753 , \33546 );
buf \U$29121 ( \34754 , \33546 );
buf \U$29122 ( \34755 , \33546 );
nor \U$29123 ( \34756 , \33533 , \33534 , \33535 , \33536 , \33540 , \33543 , \33546 , \34731 , \34732 , \34733 , \34734 , \34735 , \34736 , \34737 , \34738 , \34739 , \34740 , \34741 , \34742 , \34743 , \34744 , \34745 , \34746 , \34747 , \34748 , \34749 , \34750 , \34751 , \34752 , \34753 , \34754 , \34755 );
and \U$29124 ( \34757 , \7198 , \34756 );
buf \U$29125 ( \34758 , \33546 );
buf \U$29126 ( \34759 , \33546 );
buf \U$29127 ( \34760 , \33546 );
buf \U$29128 ( \34761 , \33546 );
buf \U$29129 ( \34762 , \33546 );
buf \U$29130 ( \34763 , \33546 );
buf \U$29131 ( \34764 , \33546 );
buf \U$29132 ( \34765 , \33546 );
buf \U$29133 ( \34766 , \33546 );
buf \U$29134 ( \34767 , \33546 );
buf \U$29135 ( \34768 , \33546 );
buf \U$29136 ( \34769 , \33546 );
buf \U$29137 ( \34770 , \33546 );
buf \U$29138 ( \34771 , \33546 );
buf \U$29139 ( \34772 , \33546 );
buf \U$29140 ( \34773 , \33546 );
buf \U$29141 ( \34774 , \33546 );
buf \U$29142 ( \34775 , \33546 );
buf \U$29143 ( \34776 , \33546 );
buf \U$29144 ( \34777 , \33546 );
buf \U$29145 ( \34778 , \33546 );
buf \U$29146 ( \34779 , \33546 );
buf \U$29147 ( \34780 , \33546 );
buf \U$29148 ( \34781 , \33546 );
buf \U$29149 ( \34782 , \33546 );
nor \U$29150 ( \34783 , \33574 , \33575 , \33576 , \33577 , \33539 , \33543 , \33546 , \34758 , \34759 , \34760 , \34761 , \34762 , \34763 , \34764 , \34765 , \34766 , \34767 , \34768 , \34769 , \34770 , \34771 , \34772 , \34773 , \34774 , \34775 , \34776 , \34777 , \34778 , \34779 , \34780 , \34781 , \34782 );
and \U$29151 ( \34784 , \7200 , \34783 );
buf \U$29152 ( \34785 , \33546 );
buf \U$29153 ( \34786 , \33546 );
buf \U$29154 ( \34787 , \33546 );
buf \U$29155 ( \34788 , \33546 );
buf \U$29156 ( \34789 , \33546 );
buf \U$29157 ( \34790 , \33546 );
buf \U$29158 ( \34791 , \33546 );
buf \U$29159 ( \34792 , \33546 );
buf \U$29160 ( \34793 , \33546 );
buf \U$29161 ( \34794 , \33546 );
buf \U$29162 ( \34795 , \33546 );
buf \U$29163 ( \34796 , \33546 );
buf \U$29164 ( \34797 , \33546 );
buf \U$29165 ( \34798 , \33546 );
buf \U$29166 ( \34799 , \33546 );
buf \U$29167 ( \34800 , \33546 );
buf \U$29168 ( \34801 , \33546 );
buf \U$29169 ( \34802 , \33546 );
buf \U$29170 ( \34803 , \33546 );
buf \U$29171 ( \34804 , \33546 );
buf \U$29172 ( \34805 , \33546 );
buf \U$29173 ( \34806 , \33546 );
buf \U$29174 ( \34807 , \33546 );
buf \U$29175 ( \34808 , \33546 );
buf \U$29176 ( \34809 , \33546 );
nor \U$29177 ( \34810 , \33533 , \33575 , \33576 , \33577 , \33539 , \33543 , \33546 , \34785 , \34786 , \34787 , \34788 , \34789 , \34790 , \34791 , \34792 , \34793 , \34794 , \34795 , \34796 , \34797 , \34798 , \34799 , \34800 , \34801 , \34802 , \34803 , \34804 , \34805 , \34806 , \34807 , \34808 , \34809 );
and \U$29178 ( \34811 , \8645 , \34810 );
buf \U$29179 ( \34812 , \33546 );
buf \U$29180 ( \34813 , \33546 );
buf \U$29181 ( \34814 , \33546 );
buf \U$29182 ( \34815 , \33546 );
buf \U$29183 ( \34816 , \33546 );
buf \U$29184 ( \34817 , \33546 );
buf \U$29185 ( \34818 , \33546 );
buf \U$29186 ( \34819 , \33546 );
buf \U$29187 ( \34820 , \33546 );
buf \U$29188 ( \34821 , \33546 );
buf \U$29189 ( \34822 , \33546 );
buf \U$29190 ( \34823 , \33546 );
buf \U$29191 ( \34824 , \33546 );
buf \U$29192 ( \34825 , \33546 );
buf \U$29193 ( \34826 , \33546 );
buf \U$29194 ( \34827 , \33546 );
buf \U$29195 ( \34828 , \33546 );
buf \U$29196 ( \34829 , \33546 );
buf \U$29197 ( \34830 , \33546 );
buf \U$29198 ( \34831 , \33546 );
buf \U$29199 ( \34832 , \33546 );
buf \U$29200 ( \34833 , \33546 );
buf \U$29201 ( \34834 , \33546 );
buf \U$29202 ( \34835 , \33546 );
buf \U$29203 ( \34836 , \33546 );
nor \U$29204 ( \34837 , \33574 , \33534 , \33576 , \33577 , \33539 , \33543 , \33546 , \34812 , \34813 , \34814 , \34815 , \34816 , \34817 , \34818 , \34819 , \34820 , \34821 , \34822 , \34823 , \34824 , \34825 , \34826 , \34827 , \34828 , \34829 , \34830 , \34831 , \34832 , \34833 , \34834 , \34835 , \34836 );
and \U$29205 ( \34838 , \8673 , \34837 );
buf \U$29206 ( \34839 , \33546 );
buf \U$29207 ( \34840 , \33546 );
buf \U$29208 ( \34841 , \33546 );
buf \U$29209 ( \34842 , \33546 );
buf \U$29210 ( \34843 , \33546 );
buf \U$29211 ( \34844 , \33546 );
buf \U$29212 ( \34845 , \33546 );
buf \U$29213 ( \34846 , \33546 );
buf \U$29214 ( \34847 , \33546 );
buf \U$29215 ( \34848 , \33546 );
buf \U$29216 ( \34849 , \33546 );
buf \U$29217 ( \34850 , \33546 );
buf \U$29218 ( \34851 , \33546 );
buf \U$29219 ( \34852 , \33546 );
buf \U$29220 ( \34853 , \33546 );
buf \U$29221 ( \34854 , \33546 );
buf \U$29222 ( \34855 , \33546 );
buf \U$29223 ( \34856 , \33546 );
buf \U$29224 ( \34857 , \33546 );
buf \U$29225 ( \34858 , \33546 );
buf \U$29226 ( \34859 , \33546 );
buf \U$29227 ( \34860 , \33546 );
buf \U$29228 ( \34861 , \33546 );
buf \U$29229 ( \34862 , \33546 );
buf \U$29230 ( \34863 , \33546 );
nor \U$29231 ( \34864 , \33533 , \33534 , \33576 , \33577 , \33539 , \33543 , \33546 , \34839 , \34840 , \34841 , \34842 , \34843 , \34844 , \34845 , \34846 , \34847 , \34848 , \34849 , \34850 , \34851 , \34852 , \34853 , \34854 , \34855 , \34856 , \34857 , \34858 , \34859 , \34860 , \34861 , \34862 , \34863 );
and \U$29232 ( \34865 , \8701 , \34864 );
buf \U$29233 ( \34866 , \33546 );
buf \U$29234 ( \34867 , \33546 );
buf \U$29235 ( \34868 , \33546 );
buf \U$29236 ( \34869 , \33546 );
buf \U$29237 ( \34870 , \33546 );
buf \U$29238 ( \34871 , \33546 );
buf \U$29239 ( \34872 , \33546 );
buf \U$29240 ( \34873 , \33546 );
buf \U$29241 ( \34874 , \33546 );
buf \U$29242 ( \34875 , \33546 );
buf \U$29243 ( \34876 , \33546 );
buf \U$29244 ( \34877 , \33546 );
buf \U$29245 ( \34878 , \33546 );
buf \U$29246 ( \34879 , \33546 );
buf \U$29247 ( \34880 , \33546 );
buf \U$29248 ( \34881 , \33546 );
buf \U$29249 ( \34882 , \33546 );
buf \U$29250 ( \34883 , \33546 );
buf \U$29251 ( \34884 , \33546 );
buf \U$29252 ( \34885 , \33546 );
buf \U$29253 ( \34886 , \33546 );
buf \U$29254 ( \34887 , \33546 );
buf \U$29255 ( \34888 , \33546 );
buf \U$29256 ( \34889 , \33546 );
buf \U$29257 ( \34890 , \33546 );
nor \U$29258 ( \34891 , \33574 , \33575 , \33535 , \33577 , \33539 , \33543 , \33546 , \34866 , \34867 , \34868 , \34869 , \34870 , \34871 , \34872 , \34873 , \34874 , \34875 , \34876 , \34877 , \34878 , \34879 , \34880 , \34881 , \34882 , \34883 , \34884 , \34885 , \34886 , \34887 , \34888 , \34889 , \34890 );
and \U$29259 ( \34892 , \8729 , \34891 );
buf \U$29260 ( \34893 , \33546 );
buf \U$29261 ( \34894 , \33546 );
buf \U$29262 ( \34895 , \33546 );
buf \U$29263 ( \34896 , \33546 );
buf \U$29264 ( \34897 , \33546 );
buf \U$29265 ( \34898 , \33546 );
buf \U$29266 ( \34899 , \33546 );
buf \U$29267 ( \34900 , \33546 );
buf \U$29268 ( \34901 , \33546 );
buf \U$29269 ( \34902 , \33546 );
buf \U$29270 ( \34903 , \33546 );
buf \U$29271 ( \34904 , \33546 );
buf \U$29272 ( \34905 , \33546 );
buf \U$29273 ( \34906 , \33546 );
buf \U$29274 ( \34907 , \33546 );
buf \U$29275 ( \34908 , \33546 );
buf \U$29276 ( \34909 , \33546 );
buf \U$29277 ( \34910 , \33546 );
buf \U$29278 ( \34911 , \33546 );
buf \U$29279 ( \34912 , \33546 );
buf \U$29280 ( \34913 , \33546 );
buf \U$29281 ( \34914 , \33546 );
buf \U$29282 ( \34915 , \33546 );
buf \U$29283 ( \34916 , \33546 );
buf \U$29284 ( \34917 , \33546 );
nor \U$29285 ( \34918 , \33533 , \33575 , \33535 , \33577 , \33539 , \33543 , \33546 , \34893 , \34894 , \34895 , \34896 , \34897 , \34898 , \34899 , \34900 , \34901 , \34902 , \34903 , \34904 , \34905 , \34906 , \34907 , \34908 , \34909 , \34910 , \34911 , \34912 , \34913 , \34914 , \34915 , \34916 , \34917 );
and \U$29286 ( \34919 , \8757 , \34918 );
buf \U$29287 ( \34920 , \33546 );
buf \U$29288 ( \34921 , \33546 );
buf \U$29289 ( \34922 , \33546 );
buf \U$29290 ( \34923 , \33546 );
buf \U$29291 ( \34924 , \33546 );
buf \U$29292 ( \34925 , \33546 );
buf \U$29293 ( \34926 , \33546 );
buf \U$29294 ( \34927 , \33546 );
buf \U$29295 ( \34928 , \33546 );
buf \U$29296 ( \34929 , \33546 );
buf \U$29297 ( \34930 , \33546 );
buf \U$29298 ( \34931 , \33546 );
buf \U$29299 ( \34932 , \33546 );
buf \U$29300 ( \34933 , \33546 );
buf \U$29301 ( \34934 , \33546 );
buf \U$29302 ( \34935 , \33546 );
buf \U$29303 ( \34936 , \33546 );
buf \U$29304 ( \34937 , \33546 );
buf \U$29305 ( \34938 , \33546 );
buf \U$29306 ( \34939 , \33546 );
buf \U$29307 ( \34940 , \33546 );
buf \U$29308 ( \34941 , \33546 );
buf \U$29309 ( \34942 , \33546 );
buf \U$29310 ( \34943 , \33546 );
buf \U$29311 ( \34944 , \33546 );
nor \U$29312 ( \34945 , \33574 , \33534 , \33535 , \33577 , \33539 , \33543 , \33546 , \34920 , \34921 , \34922 , \34923 , \34924 , \34925 , \34926 , \34927 , \34928 , \34929 , \34930 , \34931 , \34932 , \34933 , \34934 , \34935 , \34936 , \34937 , \34938 , \34939 , \34940 , \34941 , \34942 , \34943 , \34944 );
and \U$29313 ( \34946 , \8785 , \34945 );
buf \U$29314 ( \34947 , \33546 );
buf \U$29315 ( \34948 , \33546 );
buf \U$29316 ( \34949 , \33546 );
buf \U$29317 ( \34950 , \33546 );
buf \U$29318 ( \34951 , \33546 );
buf \U$29319 ( \34952 , \33546 );
buf \U$29320 ( \34953 , \33546 );
buf \U$29321 ( \34954 , \33546 );
buf \U$29322 ( \34955 , \33546 );
buf \U$29323 ( \34956 , \33546 );
buf \U$29324 ( \34957 , \33546 );
buf \U$29325 ( \34958 , \33546 );
buf \U$29326 ( \34959 , \33546 );
buf \U$29327 ( \34960 , \33546 );
buf \U$29328 ( \34961 , \33546 );
buf \U$29329 ( \34962 , \33546 );
buf \U$29330 ( \34963 , \33546 );
buf \U$29331 ( \34964 , \33546 );
buf \U$29332 ( \34965 , \33546 );
buf \U$29333 ( \34966 , \33546 );
buf \U$29334 ( \34967 , \33546 );
buf \U$29335 ( \34968 , \33546 );
buf \U$29336 ( \34969 , \33546 );
buf \U$29337 ( \34970 , \33546 );
buf \U$29338 ( \34971 , \33546 );
nor \U$29339 ( \34972 , \33533 , \33534 , \33535 , \33577 , \33539 , \33543 , \33546 , \34947 , \34948 , \34949 , \34950 , \34951 , \34952 , \34953 , \34954 , \34955 , \34956 , \34957 , \34958 , \34959 , \34960 , \34961 , \34962 , \34963 , \34964 , \34965 , \34966 , \34967 , \34968 , \34969 , \34970 , \34971 );
and \U$29340 ( \34973 , \8813 , \34972 );
buf \U$29341 ( \34974 , \33546 );
buf \U$29342 ( \34975 , \33546 );
buf \U$29343 ( \34976 , \33546 );
buf \U$29344 ( \34977 , \33546 );
buf \U$29345 ( \34978 , \33546 );
buf \U$29346 ( \34979 , \33546 );
buf \U$29347 ( \34980 , \33546 );
buf \U$29348 ( \34981 , \33546 );
buf \U$29349 ( \34982 , \33546 );
buf \U$29350 ( \34983 , \33546 );
buf \U$29351 ( \34984 , \33546 );
buf \U$29352 ( \34985 , \33546 );
buf \U$29353 ( \34986 , \33546 );
buf \U$29354 ( \34987 , \33546 );
buf \U$29355 ( \34988 , \33546 );
buf \U$29356 ( \34989 , \33546 );
buf \U$29357 ( \34990 , \33546 );
buf \U$29358 ( \34991 , \33546 );
buf \U$29359 ( \34992 , \33546 );
buf \U$29360 ( \34993 , \33546 );
buf \U$29361 ( \34994 , \33546 );
buf \U$29362 ( \34995 , \33546 );
buf \U$29363 ( \34996 , \33546 );
buf \U$29364 ( \34997 , \33546 );
buf \U$29365 ( \34998 , \33546 );
nor \U$29366 ( \34999 , \33574 , \33575 , \33576 , \33536 , \33539 , \33543 , \33546 , \34974 , \34975 , \34976 , \34977 , \34978 , \34979 , \34980 , \34981 , \34982 , \34983 , \34984 , \34985 , \34986 , \34987 , \34988 , \34989 , \34990 , \34991 , \34992 , \34993 , \34994 , \34995 , \34996 , \34997 , \34998 );
and \U$29367 ( \35000 , \8841 , \34999 );
buf \U$29368 ( \35001 , \33546 );
buf \U$29369 ( \35002 , \33546 );
buf \U$29370 ( \35003 , \33546 );
buf \U$29371 ( \35004 , \33546 );
buf \U$29372 ( \35005 , \33546 );
buf \U$29373 ( \35006 , \33546 );
buf \U$29374 ( \35007 , \33546 );
buf \U$29375 ( \35008 , \33546 );
buf \U$29376 ( \35009 , \33546 );
buf \U$29377 ( \35010 , \33546 );
buf \U$29378 ( \35011 , \33546 );
buf \U$29379 ( \35012 , \33546 );
buf \U$29380 ( \35013 , \33546 );
buf \U$29381 ( \35014 , \33546 );
buf \U$29382 ( \35015 , \33546 );
buf \U$29383 ( \35016 , \33546 );
buf \U$29384 ( \35017 , \33546 );
buf \U$29385 ( \35018 , \33546 );
buf \U$29386 ( \35019 , \33546 );
buf \U$29387 ( \35020 , \33546 );
buf \U$29388 ( \35021 , \33546 );
buf \U$29389 ( \35022 , \33546 );
buf \U$29390 ( \35023 , \33546 );
buf \U$29391 ( \35024 , \33546 );
buf \U$29392 ( \35025 , \33546 );
nor \U$29393 ( \35026 , \33533 , \33575 , \33576 , \33536 , \33539 , \33543 , \33546 , \35001 , \35002 , \35003 , \35004 , \35005 , \35006 , \35007 , \35008 , \35009 , \35010 , \35011 , \35012 , \35013 , \35014 , \35015 , \35016 , \35017 , \35018 , \35019 , \35020 , \35021 , \35022 , \35023 , \35024 , \35025 );
and \U$29394 ( \35027 , \8869 , \35026 );
buf \U$29395 ( \35028 , \33546 );
buf \U$29396 ( \35029 , \33546 );
buf \U$29397 ( \35030 , \33546 );
buf \U$29398 ( \35031 , \33546 );
buf \U$29399 ( \35032 , \33546 );
buf \U$29400 ( \35033 , \33546 );
buf \U$29401 ( \35034 , \33546 );
buf \U$29402 ( \35035 , \33546 );
buf \U$29403 ( \35036 , \33546 );
buf \U$29404 ( \35037 , \33546 );
buf \U$29405 ( \35038 , \33546 );
buf \U$29406 ( \35039 , \33546 );
buf \U$29407 ( \35040 , \33546 );
buf \U$29408 ( \35041 , \33546 );
buf \U$29409 ( \35042 , \33546 );
buf \U$29410 ( \35043 , \33546 );
buf \U$29411 ( \35044 , \33546 );
buf \U$29412 ( \35045 , \33546 );
buf \U$29413 ( \35046 , \33546 );
buf \U$29414 ( \35047 , \33546 );
buf \U$29415 ( \35048 , \33546 );
buf \U$29416 ( \35049 , \33546 );
buf \U$29417 ( \35050 , \33546 );
buf \U$29418 ( \35051 , \33546 );
buf \U$29419 ( \35052 , \33546 );
nor \U$29420 ( \35053 , \33574 , \33534 , \33576 , \33536 , \33539 , \33543 , \33546 , \35028 , \35029 , \35030 , \35031 , \35032 , \35033 , \35034 , \35035 , \35036 , \35037 , \35038 , \35039 , \35040 , \35041 , \35042 , \35043 , \35044 , \35045 , \35046 , \35047 , \35048 , \35049 , \35050 , \35051 , \35052 );
and \U$29421 ( \35054 , \8897 , \35053 );
buf \U$29422 ( \35055 , \33546 );
buf \U$29423 ( \35056 , \33546 );
buf \U$29424 ( \35057 , \33546 );
buf \U$29425 ( \35058 , \33546 );
buf \U$29426 ( \35059 , \33546 );
buf \U$29427 ( \35060 , \33546 );
buf \U$29428 ( \35061 , \33546 );
buf \U$29429 ( \35062 , \33546 );
buf \U$29430 ( \35063 , \33546 );
buf \U$29431 ( \35064 , \33546 );
buf \U$29432 ( \35065 , \33546 );
buf \U$29433 ( \35066 , \33546 );
buf \U$29434 ( \35067 , \33546 );
buf \U$29435 ( \35068 , \33546 );
buf \U$29436 ( \35069 , \33546 );
buf \U$29437 ( \35070 , \33546 );
buf \U$29438 ( \35071 , \33546 );
buf \U$29439 ( \35072 , \33546 );
buf \U$29440 ( \35073 , \33546 );
buf \U$29441 ( \35074 , \33546 );
buf \U$29442 ( \35075 , \33546 );
buf \U$29443 ( \35076 , \33546 );
buf \U$29444 ( \35077 , \33546 );
buf \U$29445 ( \35078 , \33546 );
buf \U$29446 ( \35079 , \33546 );
nor \U$29447 ( \35080 , \33533 , \33534 , \33576 , \33536 , \33539 , \33543 , \33546 , \35055 , \35056 , \35057 , \35058 , \35059 , \35060 , \35061 , \35062 , \35063 , \35064 , \35065 , \35066 , \35067 , \35068 , \35069 , \35070 , \35071 , \35072 , \35073 , \35074 , \35075 , \35076 , \35077 , \35078 , \35079 );
and \U$29448 ( \35081 , \8925 , \35080 );
buf \U$29449 ( \35082 , \33546 );
buf \U$29450 ( \35083 , \33546 );
buf \U$29451 ( \35084 , \33546 );
buf \U$29452 ( \35085 , \33546 );
buf \U$29453 ( \35086 , \33546 );
buf \U$29454 ( \35087 , \33546 );
buf \U$29455 ( \35088 , \33546 );
buf \U$29456 ( \35089 , \33546 );
buf \U$29457 ( \35090 , \33546 );
buf \U$29458 ( \35091 , \33546 );
buf \U$29459 ( \35092 , \33546 );
buf \U$29460 ( \35093 , \33546 );
buf \U$29461 ( \35094 , \33546 );
buf \U$29462 ( \35095 , \33546 );
buf \U$29463 ( \35096 , \33546 );
buf \U$29464 ( \35097 , \33546 );
buf \U$29465 ( \35098 , \33546 );
buf \U$29466 ( \35099 , \33546 );
buf \U$29467 ( \35100 , \33546 );
buf \U$29468 ( \35101 , \33546 );
buf \U$29469 ( \35102 , \33546 );
buf \U$29470 ( \35103 , \33546 );
buf \U$29471 ( \35104 , \33546 );
buf \U$29472 ( \35105 , \33546 );
buf \U$29473 ( \35106 , \33546 );
nor \U$29474 ( \35107 , \33574 , \33575 , \33535 , \33536 , \33539 , \33543 , \33546 , \35082 , \35083 , \35084 , \35085 , \35086 , \35087 , \35088 , \35089 , \35090 , \35091 , \35092 , \35093 , \35094 , \35095 , \35096 , \35097 , \35098 , \35099 , \35100 , \35101 , \35102 , \35103 , \35104 , \35105 , \35106 );
and \U$29475 ( \35108 , \8953 , \35107 );
buf \U$29476 ( \35109 , \33546 );
buf \U$29477 ( \35110 , \33546 );
buf \U$29478 ( \35111 , \33546 );
buf \U$29479 ( \35112 , \33546 );
buf \U$29480 ( \35113 , \33546 );
buf \U$29481 ( \35114 , \33546 );
buf \U$29482 ( \35115 , \33546 );
buf \U$29483 ( \35116 , \33546 );
buf \U$29484 ( \35117 , \33546 );
buf \U$29485 ( \35118 , \33546 );
buf \U$29486 ( \35119 , \33546 );
buf \U$29487 ( \35120 , \33546 );
buf \U$29488 ( \35121 , \33546 );
buf \U$29489 ( \35122 , \33546 );
buf \U$29490 ( \35123 , \33546 );
buf \U$29491 ( \35124 , \33546 );
buf \U$29492 ( \35125 , \33546 );
buf \U$29493 ( \35126 , \33546 );
buf \U$29494 ( \35127 , \33546 );
buf \U$29495 ( \35128 , \33546 );
buf \U$29496 ( \35129 , \33546 );
buf \U$29497 ( \35130 , \33546 );
buf \U$29498 ( \35131 , \33546 );
buf \U$29499 ( \35132 , \33546 );
buf \U$29500 ( \35133 , \33546 );
nor \U$29501 ( \35134 , \33533 , \33575 , \33535 , \33536 , \33539 , \33543 , \33546 , \35109 , \35110 , \35111 , \35112 , \35113 , \35114 , \35115 , \35116 , \35117 , \35118 , \35119 , \35120 , \35121 , \35122 , \35123 , \35124 , \35125 , \35126 , \35127 , \35128 , \35129 , \35130 , \35131 , \35132 , \35133 );
and \U$29502 ( \35135 , \8981 , \35134 );
buf \U$29503 ( \35136 , \33546 );
buf \U$29504 ( \35137 , \33546 );
buf \U$29505 ( \35138 , \33546 );
buf \U$29506 ( \35139 , \33546 );
buf \U$29507 ( \35140 , \33546 );
buf \U$29508 ( \35141 , \33546 );
buf \U$29509 ( \35142 , \33546 );
buf \U$29510 ( \35143 , \33546 );
buf \U$29511 ( \35144 , \33546 );
buf \U$29512 ( \35145 , \33546 );
buf \U$29513 ( \35146 , \33546 );
buf \U$29514 ( \35147 , \33546 );
buf \U$29515 ( \35148 , \33546 );
buf \U$29516 ( \35149 , \33546 );
buf \U$29517 ( \35150 , \33546 );
buf \U$29518 ( \35151 , \33546 );
buf \U$29519 ( \35152 , \33546 );
buf \U$29520 ( \35153 , \33546 );
buf \U$29521 ( \35154 , \33546 );
buf \U$29522 ( \35155 , \33546 );
buf \U$29523 ( \35156 , \33546 );
buf \U$29524 ( \35157 , \33546 );
buf \U$29525 ( \35158 , \33546 );
buf \U$29526 ( \35159 , \33546 );
buf \U$29527 ( \35160 , \33546 );
nor \U$29528 ( \35161 , \33574 , \33534 , \33535 , \33536 , \33539 , \33543 , \33546 , \35136 , \35137 , \35138 , \35139 , \35140 , \35141 , \35142 , \35143 , \35144 , \35145 , \35146 , \35147 , \35148 , \35149 , \35150 , \35151 , \35152 , \35153 , \35154 , \35155 , \35156 , \35157 , \35158 , \35159 , \35160 );
and \U$29529 ( \35162 , \9009 , \35161 );
or \U$29530 ( \35163 , \34757 , \34784 , \34811 , \34838 , \34865 , \34892 , \34919 , \34946 , \34973 , \35000 , \35027 , \35054 , \35081 , \35108 , \35135 , \35162 );
buf \U$29531 ( \35164 , \33546 );
not \U$29532 ( \35165 , \35164 );
buf \U$29533 ( \35166 , \33534 );
buf \U$29534 ( \35167 , \33535 );
buf \U$29535 ( \35168 , \33536 );
buf \U$29536 ( \35169 , \33539 );
buf \U$29537 ( \35170 , \33543 );
buf \U$29538 ( \35171 , \33546 );
buf \U$29539 ( \35172 , \33546 );
buf \U$29540 ( \35173 , \33546 );
buf \U$29541 ( \35174 , \33546 );
buf \U$29542 ( \35175 , \33546 );
buf \U$29543 ( \35176 , \33546 );
buf \U$29544 ( \35177 , \33546 );
buf \U$29545 ( \35178 , \33546 );
buf \U$29546 ( \35179 , \33546 );
buf \U$29547 ( \35180 , \33546 );
buf \U$29548 ( \35181 , \33546 );
buf \U$29549 ( \35182 , \33546 );
buf \U$29550 ( \35183 , \33546 );
buf \U$29551 ( \35184 , \33546 );
buf \U$29552 ( \35185 , \33546 );
buf \U$29553 ( \35186 , \33546 );
buf \U$29554 ( \35187 , \33546 );
buf \U$29555 ( \35188 , \33546 );
buf \U$29556 ( \35189 , \33546 );
buf \U$29557 ( \35190 , \33546 );
buf \U$29558 ( \35191 , \33546 );
buf \U$29559 ( \35192 , \33546 );
buf \U$29560 ( \35193 , \33546 );
buf \U$29561 ( \35194 , \33546 );
buf \U$29562 ( \35195 , \33546 );
buf \U$29563 ( \35196 , \33533 );
or \U$29564 ( \35197 , \35166 , \35167 , \35168 , \35169 , \35170 , \35171 , \35172 , \35173 , \35174 , \35175 , \35176 , \35177 , \35178 , \35179 , \35180 , \35181 , \35182 , \35183 , \35184 , \35185 , \35186 , \35187 , \35188 , \35189 , \35190 , \35191 , \35192 , \35193 , \35194 , \35195 , \35196 );
nand \U$29565 ( \35198 , \35165 , \35197 );
buf \U$29566 ( \35199 , \35198 );
buf \U$29567 ( \35200 , \33546 );
not \U$29568 ( \35201 , \35200 );
buf \U$29569 ( \35202 , \33543 );
buf \U$29570 ( \35203 , \33546 );
buf \U$29571 ( \35204 , \33546 );
buf \U$29572 ( \35205 , \33546 );
buf \U$29573 ( \35206 , \33546 );
buf \U$29574 ( \35207 , \33546 );
buf \U$29575 ( \35208 , \33546 );
buf \U$29576 ( \35209 , \33546 );
buf \U$29577 ( \35210 , \33546 );
buf \U$29578 ( \35211 , \33546 );
buf \U$29579 ( \35212 , \33546 );
buf \U$29580 ( \35213 , \33546 );
buf \U$29581 ( \35214 , \33546 );
buf \U$29582 ( \35215 , \33546 );
buf \U$29583 ( \35216 , \33546 );
buf \U$29584 ( \35217 , \33546 );
buf \U$29585 ( \35218 , \33546 );
buf \U$29586 ( \35219 , \33546 );
buf \U$29587 ( \35220 , \33546 );
buf \U$29588 ( \35221 , \33546 );
buf \U$29589 ( \35222 , \33546 );
buf \U$29590 ( \35223 , \33546 );
buf \U$29591 ( \35224 , \33546 );
buf \U$29592 ( \35225 , \33546 );
buf \U$29593 ( \35226 , \33546 );
buf \U$29594 ( \35227 , \33546 );
buf \U$29595 ( \35228 , \33539 );
buf \U$29596 ( \35229 , \33533 );
buf \U$29597 ( \35230 , \33534 );
buf \U$29598 ( \35231 , \33535 );
buf \U$29599 ( \35232 , \33536 );
or \U$29600 ( \35233 , \35229 , \35230 , \35231 , \35232 );
and \U$29601 ( \35234 , \35228 , \35233 );
or \U$29602 ( \35235 , \35202 , \35203 , \35204 , \35205 , \35206 , \35207 , \35208 , \35209 , \35210 , \35211 , \35212 , \35213 , \35214 , \35215 , \35216 , \35217 , \35218 , \35219 , \35220 , \35221 , \35222 , \35223 , \35224 , \35225 , \35226 , \35227 , \35234 );
and \U$29603 ( \35236 , \35201 , \35235 );
buf \U$29604 ( \35237 , \35236 );
or \U$29605 ( \35238 , \35199 , \35237 );
_DC ga0c2 ( \35239_nGa0c2 , \35163 , \35238 );
buf \U$29606 ( \35240 , \35239_nGa0c2 );
xor \U$29607 ( \35241 , \34730 , \35240 );
buf \U$29608 ( \35242 , RIb7af5b8_255);
and \U$29609 ( \35243 , \7207 , \34756 );
and \U$29610 ( \35244 , \7209 , \34783 );
and \U$29611 ( \35245 , \9119 , \34810 );
and \U$29612 ( \35246 , \9121 , \34837 );
and \U$29613 ( \35247 , \9123 , \34864 );
and \U$29614 ( \35248 , \9125 , \34891 );
and \U$29615 ( \35249 , \9127 , \34918 );
and \U$29616 ( \35250 , \9129 , \34945 );
and \U$29617 ( \35251 , \9131 , \34972 );
and \U$29618 ( \35252 , \9133 , \34999 );
and \U$29619 ( \35253 , \9135 , \35026 );
and \U$29620 ( \35254 , \9137 , \35053 );
and \U$29621 ( \35255 , \9139 , \35080 );
and \U$29622 ( \35256 , \9141 , \35107 );
and \U$29623 ( \35257 , \9143 , \35134 );
and \U$29624 ( \35258 , \9145 , \35161 );
or \U$29625 ( \35259 , \35243 , \35244 , \35245 , \35246 , \35247 , \35248 , \35249 , \35250 , \35251 , \35252 , \35253 , \35254 , \35255 , \35256 , \35257 , \35258 );
_DC ga0d7 ( \35260_nGa0d7 , \35259 , \35238 );
buf \U$29626 ( \35261 , \35260_nGa0d7 );
xor \U$29627 ( \35262 , \35242 , \35261 );
or \U$29628 ( \35263 , \35241 , \35262 );
buf \U$29629 ( \35264 , RIb7af540_256);
and \U$29630 ( \35265 , \7217 , \34756 );
and \U$29631 ( \35266 , \7219 , \34783 );
and \U$29632 ( \35267 , \9155 , \34810 );
and \U$29633 ( \35268 , \9157 , \34837 );
and \U$29634 ( \35269 , \9159 , \34864 );
and \U$29635 ( \35270 , \9161 , \34891 );
and \U$29636 ( \35271 , \9163 , \34918 );
and \U$29637 ( \35272 , \9165 , \34945 );
and \U$29638 ( \35273 , \9167 , \34972 );
and \U$29639 ( \35274 , \9169 , \34999 );
and \U$29640 ( \35275 , \9171 , \35026 );
and \U$29641 ( \35276 , \9173 , \35053 );
and \U$29642 ( \35277 , \9175 , \35080 );
and \U$29643 ( \35278 , \9177 , \35107 );
and \U$29644 ( \35279 , \9179 , \35134 );
and \U$29645 ( \35280 , \9181 , \35161 );
or \U$29646 ( \35281 , \35265 , \35266 , \35267 , \35268 , \35269 , \35270 , \35271 , \35272 , \35273 , \35274 , \35275 , \35276 , \35277 , \35278 , \35279 , \35280 );
_DC ga0ed ( \35282_nGa0ed , \35281 , \35238 );
buf \U$29647 ( \35283 , \35282_nGa0ed );
xor \U$29648 ( \35284 , \35264 , \35283 );
or \U$29649 ( \35285 , \35263 , \35284 );
buf \U$29650 ( \35286 , RIb7af4c8_257);
and \U$29651 ( \35287 , \7227 , \34756 );
and \U$29652 ( \35288 , \7229 , \34783 );
and \U$29653 ( \35289 , \9191 , \34810 );
and \U$29654 ( \35290 , \9193 , \34837 );
and \U$29655 ( \35291 , \9195 , \34864 );
and \U$29656 ( \35292 , \9197 , \34891 );
and \U$29657 ( \35293 , \9199 , \34918 );
and \U$29658 ( \35294 , \9201 , \34945 );
and \U$29659 ( \35295 , \9203 , \34972 );
and \U$29660 ( \35296 , \9205 , \34999 );
and \U$29661 ( \35297 , \9207 , \35026 );
and \U$29662 ( \35298 , \9209 , \35053 );
and \U$29663 ( \35299 , \9211 , \35080 );
and \U$29664 ( \35300 , \9213 , \35107 );
and \U$29665 ( \35301 , \9215 , \35134 );
and \U$29666 ( \35302 , \9217 , \35161 );
or \U$29667 ( \35303 , \35287 , \35288 , \35289 , \35290 , \35291 , \35292 , \35293 , \35294 , \35295 , \35296 , \35297 , \35298 , \35299 , \35300 , \35301 , \35302 );
_DC ga103 ( \35304_nGa103 , \35303 , \35238 );
buf \U$29668 ( \35305 , \35304_nGa103 );
xor \U$29669 ( \35306 , \35286 , \35305 );
or \U$29670 ( \35307 , \35285 , \35306 );
buf \U$29671 ( \35308 , RIb7af450_258);
and \U$29672 ( \35309 , \7237 , \34756 );
and \U$29673 ( \35310 , \7239 , \34783 );
and \U$29674 ( \35311 , \9227 , \34810 );
and \U$29675 ( \35312 , \9229 , \34837 );
and \U$29676 ( \35313 , \9231 , \34864 );
and \U$29677 ( \35314 , \9233 , \34891 );
and \U$29678 ( \35315 , \9235 , \34918 );
and \U$29679 ( \35316 , \9237 , \34945 );
and \U$29680 ( \35317 , \9239 , \34972 );
and \U$29681 ( \35318 , \9241 , \34999 );
and \U$29682 ( \35319 , \9243 , \35026 );
and \U$29683 ( \35320 , \9245 , \35053 );
and \U$29684 ( \35321 , \9247 , \35080 );
and \U$29685 ( \35322 , \9249 , \35107 );
and \U$29686 ( \35323 , \9251 , \35134 );
and \U$29687 ( \35324 , \9253 , \35161 );
or \U$29688 ( \35325 , \35309 , \35310 , \35311 , \35312 , \35313 , \35314 , \35315 , \35316 , \35317 , \35318 , \35319 , \35320 , \35321 , \35322 , \35323 , \35324 );
_DC ga119 ( \35326_nGa119 , \35325 , \35238 );
buf \U$29689 ( \35327 , \35326_nGa119 );
xor \U$29690 ( \35328 , \35308 , \35327 );
or \U$29691 ( \35329 , \35307 , \35328 );
buf \U$29692 ( \35330 , RIb7af3d8_259);
and \U$29693 ( \35331 , \7247 , \34756 );
and \U$29694 ( \35332 , \7249 , \34783 );
and \U$29695 ( \35333 , \9263 , \34810 );
and \U$29696 ( \35334 , \9265 , \34837 );
and \U$29697 ( \35335 , \9267 , \34864 );
and \U$29698 ( \35336 , \9269 , \34891 );
and \U$29699 ( \35337 , \9271 , \34918 );
and \U$29700 ( \35338 , \9273 , \34945 );
and \U$29701 ( \35339 , \9275 , \34972 );
and \U$29702 ( \35340 , \9277 , \34999 );
and \U$29703 ( \35341 , \9279 , \35026 );
and \U$29704 ( \35342 , \9281 , \35053 );
and \U$29705 ( \35343 , \9283 , \35080 );
and \U$29706 ( \35344 , \9285 , \35107 );
and \U$29707 ( \35345 , \9287 , \35134 );
and \U$29708 ( \35346 , \9289 , \35161 );
or \U$29709 ( \35347 , \35331 , \35332 , \35333 , \35334 , \35335 , \35336 , \35337 , \35338 , \35339 , \35340 , \35341 , \35342 , \35343 , \35344 , \35345 , \35346 );
_DC ga12f ( \35348_nGa12f , \35347 , \35238 );
buf \U$29710 ( \35349 , \35348_nGa12f );
xor \U$29711 ( \35350 , \35330 , \35349 );
or \U$29712 ( \35351 , \35329 , \35350 );
buf \U$29713 ( \35352 , RIb7a5bf8_260);
and \U$29714 ( \35353 , \7257 , \34756 );
and \U$29715 ( \35354 , \7259 , \34783 );
and \U$29716 ( \35355 , \9299 , \34810 );
and \U$29717 ( \35356 , \9301 , \34837 );
and \U$29718 ( \35357 , \9303 , \34864 );
and \U$29719 ( \35358 , \9305 , \34891 );
and \U$29720 ( \35359 , \9307 , \34918 );
and \U$29721 ( \35360 , \9309 , \34945 );
and \U$29722 ( \35361 , \9311 , \34972 );
and \U$29723 ( \35362 , \9313 , \34999 );
and \U$29724 ( \35363 , \9315 , \35026 );
and \U$29725 ( \35364 , \9317 , \35053 );
and \U$29726 ( \35365 , \9319 , \35080 );
and \U$29727 ( \35366 , \9321 , \35107 );
and \U$29728 ( \35367 , \9323 , \35134 );
and \U$29729 ( \35368 , \9325 , \35161 );
or \U$29730 ( \35369 , \35353 , \35354 , \35355 , \35356 , \35357 , \35358 , \35359 , \35360 , \35361 , \35362 , \35363 , \35364 , \35365 , \35366 , \35367 , \35368 );
_DC ga145 ( \35370_nGa145 , \35369 , \35238 );
buf \U$29731 ( \35371 , \35370_nGa145 );
xor \U$29732 ( \35372 , \35352 , \35371 );
or \U$29733 ( \35373 , \35351 , \35372 );
buf \U$29734 ( \35374 , RIb7a0c48_261);
and \U$29735 ( \35375 , \7267 , \34756 );
and \U$29736 ( \35376 , \7269 , \34783 );
and \U$29737 ( \35377 , \9335 , \34810 );
and \U$29738 ( \35378 , \9337 , \34837 );
and \U$29739 ( \35379 , \9339 , \34864 );
and \U$29740 ( \35380 , \9341 , \34891 );
and \U$29741 ( \35381 , \9343 , \34918 );
and \U$29742 ( \35382 , \9345 , \34945 );
and \U$29743 ( \35383 , \9347 , \34972 );
and \U$29744 ( \35384 , \9349 , \34999 );
and \U$29745 ( \35385 , \9351 , \35026 );
and \U$29746 ( \35386 , \9353 , \35053 );
and \U$29747 ( \35387 , \9355 , \35080 );
and \U$29748 ( \35388 , \9357 , \35107 );
and \U$29749 ( \35389 , \9359 , \35134 );
and \U$29750 ( \35390 , \9361 , \35161 );
or \U$29751 ( \35391 , \35375 , \35376 , \35377 , \35378 , \35379 , \35380 , \35381 , \35382 , \35383 , \35384 , \35385 , \35386 , \35387 , \35388 , \35389 , \35390 );
_DC ga15b ( \35392_nGa15b , \35391 , \35238 );
buf \U$29752 ( \35393 , \35392_nGa15b );
xor \U$29753 ( \35394 , \35374 , \35393 );
or \U$29754 ( \35395 , \35373 , \35394 );
not \U$29755 ( \35396 , \35395 );
buf \U$29756 ( \35397 , \35396 );
and \U$29757 ( \35398 , \34729 , \35397 );
_HMUX ga162 ( \35399_nGa162 , \33140_nG9887 , \33533 , \35398 );
buf \U$29758 ( \35400 , \33161 );
buf \U$29759 ( \35401 , \33158 );
buf \U$29760 ( \35402 , \33143 );
buf \U$29761 ( \35403 , \33146 );
buf \U$29762 ( \35404 , \33150 );
buf \U$29763 ( \35405 , \33154 );
or \U$29764 ( \35406 , \35402 , \35403 , \35404 , \35405 );
and \U$29765 ( \35407 , \35401 , \35406 );
or \U$29766 ( \35408 , \35400 , \35407 );
buf \U$29767 ( \35409 , \35408 );
_HMUX ga16d ( \35410_nGa16d , \33532_nG9a0f , \35399_nGa162 , \35409 );
buf \U$29768 ( \35411 , RIe5319e0_6884);
buf \U$29770 ( \35412 , \35411 );
buf \U$29771 ( \35413 , RIe549ef0_6842);
not \U$29772 ( \35414 , \35413 );
buf \U$29773 ( \35415 , \35414 );
buf \U$29774 ( \35416 , RIe549770_6843);
xor \U$29775 ( \35417 , \35416 , \35413 );
buf \U$29776 ( \35418 , \35417 );
buf \U$29777 ( \35419 , RIe548ff0_6844);
and \U$29778 ( \35420 , \35416 , \35413 );
xor \U$29779 ( \35421 , \35419 , \35420 );
buf \U$29780 ( \35422 , \35421 );
buf \U$29781 ( \35423 , RIea91330_6888);
and \U$29782 ( \35424 , \35419 , \35420 );
xor \U$29783 ( \35425 , \35423 , \35424 );
buf \U$29784 ( \35426 , \35425 );
not \U$29785 ( \35427 , \35426 );
and \U$29786 ( \35428 , \35423 , \35424 );
buf \U$29787 ( \35429 , \35428 );
nor \U$29788 ( \35430 , \35412 , \35415 , \35418 , \35422 , \35427 , \35429 );
and \U$29789 ( \35431 , RIe5329d0_6883, \35430 );
not \U$29790 ( \35432 , \35429 );
and \U$29791 ( \35433 , \35412 , \35415 , \35418 , \35422 , \35427 , \35432 );
and \U$29792 ( \35434 , RIeb72150_6905, \35433 );
not \U$29793 ( \35435 , \35412 );
and \U$29794 ( \35436 , \35435 , \35415 , \35418 , \35422 , \35427 , \35432 );
and \U$29795 ( \35437 , RIeab80c0_6897, \35436 );
not \U$29796 ( \35438 , \35415 );
and \U$29797 ( \35439 , \35412 , \35438 , \35418 , \35422 , \35427 , \35432 );
and \U$29798 ( \35440 , RIe5331c8_6882, \35439 );
and \U$29799 ( \35441 , \35435 , \35438 , \35418 , \35422 , \35427 , \35432 );
and \U$29800 ( \35442 , RIe5339c0_6881, \35441 );
not \U$29801 ( \35443 , \35418 );
and \U$29802 ( \35444 , \35412 , \35415 , \35443 , \35422 , \35427 , \35432 );
and \U$29803 ( \35445 , RIeab87c8_6898, \35444 );
and \U$29804 ( \35446 , \35435 , \35415 , \35443 , \35422 , \35427 , \35432 );
and \U$29805 ( \35447 , RIe5341b8_6880, \35446 );
and \U$29806 ( \35448 , \35412 , \35438 , \35443 , \35422 , \35427 , \35432 );
and \U$29807 ( \35449 , RIe5349b0_6879, \35448 );
and \U$29808 ( \35450 , \35435 , \35438 , \35443 , \35422 , \35427 , \35432 );
and \U$29809 ( \35451 , RIea94af8_6890, \35450 );
nor \U$29810 ( \35452 , \35435 , \35438 , \35443 , \35422 , \35426 , \35429 );
and \U$29811 ( \35453 , RIe5351a8_6878, \35452 );
nor \U$29812 ( \35454 , \35412 , \35438 , \35443 , \35422 , \35426 , \35429 );
and \U$29813 ( \35455 , RIe5359a0_6877, \35454 );
nor \U$29814 ( \35456 , \35435 , \35415 , \35443 , \35422 , \35426 , \35429 );
and \U$29815 ( \35457 , RIeab78c8_6895, \35456 );
nor \U$29816 ( \35458 , \35412 , \35415 , \35443 , \35422 , \35426 , \35429 );
and \U$29817 ( \35459 , RIeab7d00_6896, \35458 );
nor \U$29818 ( \35460 , \35435 , \35438 , \35418 , \35422 , \35426 , \35429 );
and \U$29819 ( \35461 , RIeacfa18_6902, \35460 );
nor \U$29820 ( \35462 , \35412 , \35438 , \35418 , \35422 , \35426 , \35429 );
and \U$29821 ( \35463 , RIeab6518_6891, \35462 );
or \U$29823 ( \35464 , \35431 , \35434 , \35437 , \35440 , \35442 , \35445 , \35447 , \35449 , \35451 , \35453 , \35455 , \35457 , \35459 , \35461 , \35463 , 1'b0 );
buf \U$29825 ( \35465 , \35429 );
buf \U$29826 ( \35466 , \35426 );
buf \U$29827 ( \35467 , \35412 );
buf \U$29828 ( \35468 , \35415 );
buf \U$29829 ( \35469 , \35418 );
buf \U$29830 ( \35470 , \35422 );
or \U$29831 ( \35471 , \35467 , \35468 , \35469 , \35470 );
and \U$29832 ( \35472 , \35466 , \35471 );
or \U$29833 ( \35473 , \35465 , \35472 );
buf \U$29834 ( \35474 , \35473 );
or \U$29835 ( \35475 , 1'b0 , \35474 );
_DC ga1b0 ( \35476_nGa1b0 , \35464 , \35475 );
not \U$29836 ( \35477 , \35476_nGa1b0 );
buf \U$29837 ( \35478 , RIb7b9608_246);
and \U$29838 ( \35479 , \7117 , \35430 );
and \U$29839 ( \35480 , \7119 , \35433 );
and \U$29840 ( \35481 , \7864 , \35436 );
and \U$29841 ( \35482 , \7892 , \35439 );
and \U$29842 ( \35483 , \7920 , \35441 );
and \U$29843 ( \35484 , \7948 , \35444 );
and \U$29844 ( \35485 , \7976 , \35446 );
and \U$29845 ( \35486 , \8004 , \35448 );
and \U$29846 ( \35487 , \8032 , \35450 );
and \U$29847 ( \35488 , \8060 , \35452 );
and \U$29848 ( \35489 , \8088 , \35454 );
and \U$29849 ( \35490 , \8116 , \35456 );
and \U$29850 ( \35491 , \8144 , \35458 );
and \U$29851 ( \35492 , \8172 , \35460 );
and \U$29852 ( \35493 , \8200 , \35462 );
or \U$29854 ( \35494 , \35479 , \35480 , \35481 , \35482 , \35483 , \35484 , \35485 , \35486 , \35487 , \35488 , \35489 , \35490 , \35491 , \35492 , \35493 , 1'b0 );
_DC ga1c3 ( \35495_nGa1c3 , \35494 , \35475 );
buf \U$29855 ( \35496 , \35495_nGa1c3 );
xor \U$29856 ( \35497 , \35478 , \35496 );
buf \U$29857 ( \35498 , RIb7b9590_247);
and \U$29858 ( \35499 , \7126 , \35430 );
and \U$29859 ( \35500 , \7128 , \35433 );
and \U$29860 ( \35501 , \8338 , \35436 );
and \U$29861 ( \35502 , \8340 , \35439 );
and \U$29862 ( \35503 , \8342 , \35441 );
and \U$29863 ( \35504 , \8344 , \35444 );
and \U$29864 ( \35505 , \8346 , \35446 );
and \U$29865 ( \35506 , \8348 , \35448 );
and \U$29866 ( \35507 , \8350 , \35450 );
and \U$29867 ( \35508 , \8352 , \35452 );
and \U$29868 ( \35509 , \8354 , \35454 );
and \U$29869 ( \35510 , \8356 , \35456 );
and \U$29870 ( \35511 , \8358 , \35458 );
and \U$29871 ( \35512 , \8360 , \35460 );
and \U$29872 ( \35513 , \8362 , \35462 );
or \U$29874 ( \35514 , \35499 , \35500 , \35501 , \35502 , \35503 , \35504 , \35505 , \35506 , \35507 , \35508 , \35509 , \35510 , \35511 , \35512 , \35513 , 1'b0 );
_DC ga1d7 ( \35515_nGa1d7 , \35514 , \35475 );
buf \U$29875 ( \35516 , \35515_nGa1d7 );
xor \U$29876 ( \35517 , \35498 , \35516 );
or \U$29877 ( \35518 , \35497 , \35517 );
buf \U$29878 ( \35519 , RIb7b9518_248);
and \U$29879 ( \35520 , \7136 , \35430 );
and \U$29880 ( \35521 , \7138 , \35433 );
and \U$29881 ( \35522 , \8374 , \35436 );
and \U$29882 ( \35523 , \8376 , \35439 );
and \U$29883 ( \35524 , \8378 , \35441 );
and \U$29884 ( \35525 , \8380 , \35444 );
and \U$29885 ( \35526 , \8382 , \35446 );
and \U$29886 ( \35527 , \8384 , \35448 );
and \U$29887 ( \35528 , \8386 , \35450 );
and \U$29888 ( \35529 , \8388 , \35452 );
and \U$29889 ( \35530 , \8390 , \35454 );
and \U$29890 ( \35531 , \8392 , \35456 );
and \U$29891 ( \35532 , \8394 , \35458 );
and \U$29892 ( \35533 , \8396 , \35460 );
and \U$29893 ( \35534 , \8398 , \35462 );
or \U$29895 ( \35535 , \35520 , \35521 , \35522 , \35523 , \35524 , \35525 , \35526 , \35527 , \35528 , \35529 , \35530 , \35531 , \35532 , \35533 , \35534 , 1'b0 );
_DC ga1ec ( \35536_nGa1ec , \35535 , \35475 );
buf \U$29896 ( \35537 , \35536_nGa1ec );
xor \U$29897 ( \35538 , \35519 , \35537 );
or \U$29898 ( \35539 , \35518 , \35538 );
buf \U$29899 ( \35540 , RIb7b94a0_249);
and \U$29900 ( \35541 , \7146 , \35430 );
and \U$29901 ( \35542 , \7148 , \35433 );
and \U$29902 ( \35543 , \8410 , \35436 );
and \U$29903 ( \35544 , \8412 , \35439 );
and \U$29904 ( \35545 , \8414 , \35441 );
and \U$29905 ( \35546 , \8416 , \35444 );
and \U$29906 ( \35547 , \8418 , \35446 );
and \U$29907 ( \35548 , \8420 , \35448 );
and \U$29908 ( \35549 , \8422 , \35450 );
and \U$29909 ( \35550 , \8424 , \35452 );
and \U$29910 ( \35551 , \8426 , \35454 );
and \U$29911 ( \35552 , \8428 , \35456 );
and \U$29912 ( \35553 , \8430 , \35458 );
and \U$29913 ( \35554 , \8432 , \35460 );
and \U$29914 ( \35555 , \8434 , \35462 );
or \U$29916 ( \35556 , \35541 , \35542 , \35543 , \35544 , \35545 , \35546 , \35547 , \35548 , \35549 , \35550 , \35551 , \35552 , \35553 , \35554 , \35555 , 1'b0 );
_DC ga201 ( \35557_nGa201 , \35556 , \35475 );
buf \U$29917 ( \35558 , \35557_nGa201 );
xor \U$29918 ( \35559 , \35540 , \35558 );
or \U$29919 ( \35560 , \35539 , \35559 );
buf \U$29920 ( \35561 , RIb7b9428_250);
and \U$29921 ( \35562 , \7156 , \35430 );
and \U$29922 ( \35563 , \7158 , \35433 );
and \U$29923 ( \35564 , \8446 , \35436 );
and \U$29924 ( \35565 , \8448 , \35439 );
and \U$29925 ( \35566 , \8450 , \35441 );
and \U$29926 ( \35567 , \8452 , \35444 );
and \U$29927 ( \35568 , \8454 , \35446 );
and \U$29928 ( \35569 , \8456 , \35448 );
and \U$29929 ( \35570 , \8458 , \35450 );
and \U$29930 ( \35571 , \8460 , \35452 );
and \U$29931 ( \35572 , \8462 , \35454 );
and \U$29932 ( \35573 , \8464 , \35456 );
and \U$29933 ( \35574 , \8466 , \35458 );
and \U$29934 ( \35575 , \8468 , \35460 );
and \U$29935 ( \35576 , \8470 , \35462 );
or \U$29937 ( \35577 , \35562 , \35563 , \35564 , \35565 , \35566 , \35567 , \35568 , \35569 , \35570 , \35571 , \35572 , \35573 , \35574 , \35575 , \35576 , 1'b0 );
_DC ga216 ( \35578_nGa216 , \35577 , \35475 );
buf \U$29938 ( \35579 , \35578_nGa216 );
xor \U$29939 ( \35580 , \35561 , \35579 );
or \U$29940 ( \35581 , \35560 , \35580 );
buf \U$29941 ( \35582 , RIb7b93b0_251);
and \U$29942 ( \35583 , \7166 , \35430 );
and \U$29943 ( \35584 , \7168 , \35433 );
and \U$29944 ( \35585 , \8482 , \35436 );
and \U$29945 ( \35586 , \8484 , \35439 );
and \U$29946 ( \35587 , \8486 , \35441 );
and \U$29947 ( \35588 , \8488 , \35444 );
and \U$29948 ( \35589 , \8490 , \35446 );
and \U$29949 ( \35590 , \8492 , \35448 );
and \U$29950 ( \35591 , \8494 , \35450 );
and \U$29951 ( \35592 , \8496 , \35452 );
and \U$29952 ( \35593 , \8498 , \35454 );
and \U$29953 ( \35594 , \8500 , \35456 );
and \U$29954 ( \35595 , \8502 , \35458 );
and \U$29955 ( \35596 , \8504 , \35460 );
and \U$29956 ( \35597 , \8506 , \35462 );
or \U$29958 ( \35598 , \35583 , \35584 , \35585 , \35586 , \35587 , \35588 , \35589 , \35590 , \35591 , \35592 , \35593 , \35594 , \35595 , \35596 , \35597 , 1'b0 );
_DC ga22b ( \35599_nGa22b , \35598 , \35475 );
buf \U$29959 ( \35600 , \35599_nGa22b );
xor \U$29960 ( \35601 , \35582 , \35600 );
or \U$29961 ( \35602 , \35581 , \35601 );
buf \U$29962 ( \35603 , RIb7af720_252);
and \U$29963 ( \35604 , \7176 , \35430 );
and \U$29964 ( \35605 , \7178 , \35433 );
and \U$29965 ( \35606 , \8518 , \35436 );
and \U$29966 ( \35607 , \8520 , \35439 );
and \U$29967 ( \35608 , \8522 , \35441 );
and \U$29968 ( \35609 , \8524 , \35444 );
and \U$29969 ( \35610 , \8526 , \35446 );
and \U$29970 ( \35611 , \8528 , \35448 );
and \U$29971 ( \35612 , \8530 , \35450 );
and \U$29972 ( \35613 , \8532 , \35452 );
and \U$29973 ( \35614 , \8534 , \35454 );
and \U$29974 ( \35615 , \8536 , \35456 );
and \U$29975 ( \35616 , \8538 , \35458 );
and \U$29976 ( \35617 , \8540 , \35460 );
and \U$29977 ( \35618 , \8542 , \35462 );
or \U$29979 ( \35619 , \35604 , \35605 , \35606 , \35607 , \35608 , \35609 , \35610 , \35611 , \35612 , \35613 , \35614 , \35615 , \35616 , \35617 , \35618 , 1'b0 );
_DC ga240 ( \35620_nGa240 , \35619 , \35475 );
buf \U$29980 ( \35621 , \35620_nGa240 );
xor \U$29981 ( \35622 , \35603 , \35621 );
or \U$29982 ( \35623 , \35602 , \35622 );
buf \U$29983 ( \35624 , RIb7af6a8_253);
and \U$29984 ( \35625 , \7186 , \35430 );
and \U$29985 ( \35626 , \7188 , \35433 );
and \U$29986 ( \35627 , \8554 , \35436 );
and \U$29987 ( \35628 , \8556 , \35439 );
and \U$29988 ( \35629 , \8558 , \35441 );
and \U$29989 ( \35630 , \8560 , \35444 );
and \U$29990 ( \35631 , \8562 , \35446 );
and \U$29991 ( \35632 , \8564 , \35448 );
and \U$29992 ( \35633 , \8566 , \35450 );
and \U$29993 ( \35634 , \8568 , \35452 );
and \U$29994 ( \35635 , \8570 , \35454 );
and \U$29995 ( \35636 , \8572 , \35456 );
and \U$29996 ( \35637 , \8574 , \35458 );
and \U$29997 ( \35638 , \8576 , \35460 );
and \U$29998 ( \35639 , \8578 , \35462 );
or \U$30000 ( \35640 , \35625 , \35626 , \35627 , \35628 , \35629 , \35630 , \35631 , \35632 , \35633 , \35634 , \35635 , \35636 , \35637 , \35638 , \35639 , 1'b0 );
_DC ga255 ( \35641_nGa255 , \35640 , \35475 );
buf \U$30001 ( \35642 , \35641_nGa255 );
xor \U$30002 ( \35643 , \35624 , \35642 );
or \U$30003 ( \35644 , \35623 , \35643 );
not \U$30004 ( \35645 , \35644 );
buf \U$30005 ( \35646 , \35645 );
buf \U$30006 ( \35647 , RIb7af630_254);
and \U$30007 ( \35648 , \7198 , \35430 );
and \U$30008 ( \35649 , \7200 , \35433 );
and \U$30009 ( \35650 , \8645 , \35436 );
and \U$30010 ( \35651 , \8673 , \35439 );
and \U$30011 ( \35652 , \8701 , \35441 );
and \U$30012 ( \35653 , \8729 , \35444 );
and \U$30013 ( \35654 , \8757 , \35446 );
and \U$30014 ( \35655 , \8785 , \35448 );
and \U$30015 ( \35656 , \8813 , \35450 );
and \U$30016 ( \35657 , \8841 , \35452 );
and \U$30017 ( \35658 , \8869 , \35454 );
and \U$30018 ( \35659 , \8897 , \35456 );
and \U$30019 ( \35660 , \8925 , \35458 );
and \U$30020 ( \35661 , \8953 , \35460 );
and \U$30021 ( \35662 , \8981 , \35462 );
or \U$30023 ( \35663 , \35648 , \35649 , \35650 , \35651 , \35652 , \35653 , \35654 , \35655 , \35656 , \35657 , \35658 , \35659 , \35660 , \35661 , \35662 , 1'b0 );
_DC ga26c ( \35664_nGa26c , \35663 , \35475 );
buf \U$30024 ( \35665 , \35664_nGa26c );
xor \U$30025 ( \35666 , \35647 , \35665 );
buf \U$30026 ( \35667 , RIb7af5b8_255);
and \U$30027 ( \35668 , \7207 , \35430 );
and \U$30028 ( \35669 , \7209 , \35433 );
and \U$30029 ( \35670 , \9119 , \35436 );
and \U$30030 ( \35671 , \9121 , \35439 );
and \U$30031 ( \35672 , \9123 , \35441 );
and \U$30032 ( \35673 , \9125 , \35444 );
and \U$30033 ( \35674 , \9127 , \35446 );
and \U$30034 ( \35675 , \9129 , \35448 );
and \U$30035 ( \35676 , \9131 , \35450 );
and \U$30036 ( \35677 , \9133 , \35452 );
and \U$30037 ( \35678 , \9135 , \35454 );
and \U$30038 ( \35679 , \9137 , \35456 );
and \U$30039 ( \35680 , \9139 , \35458 );
and \U$30040 ( \35681 , \9141 , \35460 );
and \U$30041 ( \35682 , \9143 , \35462 );
or \U$30043 ( \35683 , \35668 , \35669 , \35670 , \35671 , \35672 , \35673 , \35674 , \35675 , \35676 , \35677 , \35678 , \35679 , \35680 , \35681 , \35682 , 1'b0 );
_DC ga280 ( \35684_nGa280 , \35683 , \35475 );
buf \U$30044 ( \35685 , \35684_nGa280 );
xor \U$30045 ( \35686 , \35667 , \35685 );
or \U$30046 ( \35687 , \35666 , \35686 );
buf \U$30047 ( \35688 , RIb7af540_256);
and \U$30048 ( \35689 , \7217 , \35430 );
and \U$30049 ( \35690 , \7219 , \35433 );
and \U$30050 ( \35691 , \9155 , \35436 );
and \U$30051 ( \35692 , \9157 , \35439 );
and \U$30052 ( \35693 , \9159 , \35441 );
and \U$30053 ( \35694 , \9161 , \35444 );
and \U$30054 ( \35695 , \9163 , \35446 );
and \U$30055 ( \35696 , \9165 , \35448 );
and \U$30056 ( \35697 , \9167 , \35450 );
and \U$30057 ( \35698 , \9169 , \35452 );
and \U$30058 ( \35699 , \9171 , \35454 );
and \U$30059 ( \35700 , \9173 , \35456 );
and \U$30060 ( \35701 , \9175 , \35458 );
and \U$30061 ( \35702 , \9177 , \35460 );
and \U$30062 ( \35703 , \9179 , \35462 );
or \U$30064 ( \35704 , \35689 , \35690 , \35691 , \35692 , \35693 , \35694 , \35695 , \35696 , \35697 , \35698 , \35699 , \35700 , \35701 , \35702 , \35703 , 1'b0 );
_DC ga295 ( \35705_nGa295 , \35704 , \35475 );
buf \U$30065 ( \35706 , \35705_nGa295 );
xor \U$30066 ( \35707 , \35688 , \35706 );
or \U$30067 ( \35708 , \35687 , \35707 );
buf \U$30068 ( \35709 , RIb7af4c8_257);
and \U$30069 ( \35710 , \7227 , \35430 );
and \U$30070 ( \35711 , \7229 , \35433 );
and \U$30071 ( \35712 , \9191 , \35436 );
and \U$30072 ( \35713 , \9193 , \35439 );
and \U$30073 ( \35714 , \9195 , \35441 );
and \U$30074 ( \35715 , \9197 , \35444 );
and \U$30075 ( \35716 , \9199 , \35446 );
and \U$30076 ( \35717 , \9201 , \35448 );
and \U$30077 ( \35718 , \9203 , \35450 );
and \U$30078 ( \35719 , \9205 , \35452 );
and \U$30079 ( \35720 , \9207 , \35454 );
and \U$30080 ( \35721 , \9209 , \35456 );
and \U$30081 ( \35722 , \9211 , \35458 );
and \U$30082 ( \35723 , \9213 , \35460 );
and \U$30083 ( \35724 , \9215 , \35462 );
or \U$30085 ( \35725 , \35710 , \35711 , \35712 , \35713 , \35714 , \35715 , \35716 , \35717 , \35718 , \35719 , \35720 , \35721 , \35722 , \35723 , \35724 , 1'b0 );
_DC ga2aa ( \35726_nGa2aa , \35725 , \35475 );
buf \U$30086 ( \35727 , \35726_nGa2aa );
xor \U$30087 ( \35728 , \35709 , \35727 );
or \U$30088 ( \35729 , \35708 , \35728 );
buf \U$30089 ( \35730 , RIb7af450_258);
and \U$30090 ( \35731 , \7237 , \35430 );
and \U$30091 ( \35732 , \7239 , \35433 );
and \U$30092 ( \35733 , \9227 , \35436 );
and \U$30093 ( \35734 , \9229 , \35439 );
and \U$30094 ( \35735 , \9231 , \35441 );
and \U$30095 ( \35736 , \9233 , \35444 );
and \U$30096 ( \35737 , \9235 , \35446 );
and \U$30097 ( \35738 , \9237 , \35448 );
and \U$30098 ( \35739 , \9239 , \35450 );
and \U$30099 ( \35740 , \9241 , \35452 );
and \U$30100 ( \35741 , \9243 , \35454 );
and \U$30101 ( \35742 , \9245 , \35456 );
and \U$30102 ( \35743 , \9247 , \35458 );
and \U$30103 ( \35744 , \9249 , \35460 );
and \U$30104 ( \35745 , \9251 , \35462 );
or \U$30106 ( \35746 , \35731 , \35732 , \35733 , \35734 , \35735 , \35736 , \35737 , \35738 , \35739 , \35740 , \35741 , \35742 , \35743 , \35744 , \35745 , 1'b0 );
_DC ga2bf ( \35747_nGa2bf , \35746 , \35475 );
buf \U$30107 ( \35748 , \35747_nGa2bf );
xor \U$30108 ( \35749 , \35730 , \35748 );
or \U$30109 ( \35750 , \35729 , \35749 );
buf \U$30110 ( \35751 , RIb7af3d8_259);
and \U$30111 ( \35752 , \7247 , \35430 );
and \U$30112 ( \35753 , \7249 , \35433 );
and \U$30113 ( \35754 , \9263 , \35436 );
and \U$30114 ( \35755 , \9265 , \35439 );
and \U$30115 ( \35756 , \9267 , \35441 );
and \U$30116 ( \35757 , \9269 , \35444 );
and \U$30117 ( \35758 , \9271 , \35446 );
and \U$30118 ( \35759 , \9273 , \35448 );
and \U$30119 ( \35760 , \9275 , \35450 );
and \U$30120 ( \35761 , \9277 , \35452 );
and \U$30121 ( \35762 , \9279 , \35454 );
and \U$30122 ( \35763 , \9281 , \35456 );
and \U$30123 ( \35764 , \9283 , \35458 );
and \U$30124 ( \35765 , \9285 , \35460 );
and \U$30125 ( \35766 , \9287 , \35462 );
or \U$30127 ( \35767 , \35752 , \35753 , \35754 , \35755 , \35756 , \35757 , \35758 , \35759 , \35760 , \35761 , \35762 , \35763 , \35764 , \35765 , \35766 , 1'b0 );
_DC ga2d4 ( \35768_nGa2d4 , \35767 , \35475 );
buf \U$30128 ( \35769 , \35768_nGa2d4 );
xor \U$30129 ( \35770 , \35751 , \35769 );
or \U$30130 ( \35771 , \35750 , \35770 );
buf \U$30131 ( \35772 , RIb7a5bf8_260);
and \U$30132 ( \35773 , \7257 , \35430 );
and \U$30133 ( \35774 , \7259 , \35433 );
and \U$30134 ( \35775 , \9299 , \35436 );
and \U$30135 ( \35776 , \9301 , \35439 );
and \U$30136 ( \35777 , \9303 , \35441 );
and \U$30137 ( \35778 , \9305 , \35444 );
and \U$30138 ( \35779 , \9307 , \35446 );
and \U$30139 ( \35780 , \9309 , \35448 );
and \U$30140 ( \35781 , \9311 , \35450 );
and \U$30141 ( \35782 , \9313 , \35452 );
and \U$30142 ( \35783 , \9315 , \35454 );
and \U$30143 ( \35784 , \9317 , \35456 );
and \U$30144 ( \35785 , \9319 , \35458 );
and \U$30145 ( \35786 , \9321 , \35460 );
and \U$30146 ( \35787 , \9323 , \35462 );
or \U$30148 ( \35788 , \35773 , \35774 , \35775 , \35776 , \35777 , \35778 , \35779 , \35780 , \35781 , \35782 , \35783 , \35784 , \35785 , \35786 , \35787 , 1'b0 );
_DC ga2e9 ( \35789_nGa2e9 , \35788 , \35475 );
buf \U$30149 ( \35790 , \35789_nGa2e9 );
xor \U$30150 ( \35791 , \35772 , \35790 );
or \U$30151 ( \35792 , \35771 , \35791 );
buf \U$30152 ( \35793 , RIb7a0c48_261);
and \U$30153 ( \35794 , \7267 , \35430 );
and \U$30154 ( \35795 , \7269 , \35433 );
and \U$30155 ( \35796 , \9335 , \35436 );
and \U$30156 ( \35797 , \9337 , \35439 );
and \U$30157 ( \35798 , \9339 , \35441 );
and \U$30158 ( \35799 , \9341 , \35444 );
and \U$30159 ( \35800 , \9343 , \35446 );
and \U$30160 ( \35801 , \9345 , \35448 );
and \U$30161 ( \35802 , \9347 , \35450 );
and \U$30162 ( \35803 , \9349 , \35452 );
and \U$30163 ( \35804 , \9351 , \35454 );
and \U$30164 ( \35805 , \9353 , \35456 );
and \U$30165 ( \35806 , \9355 , \35458 );
and \U$30166 ( \35807 , \9357 , \35460 );
and \U$30167 ( \35808 , \9359 , \35462 );
or \U$30169 ( \35809 , \35794 , \35795 , \35796 , \35797 , \35798 , \35799 , \35800 , \35801 , \35802 , \35803 , \35804 , \35805 , \35806 , \35807 , \35808 , 1'b0 );
_DC ga2fe ( \35810_nGa2fe , \35809 , \35475 );
buf \U$30170 ( \35811 , \35810_nGa2fe );
xor \U$30171 ( \35812 , \35793 , \35811 );
or \U$30172 ( \35813 , \35792 , \35812 );
not \U$30173 ( \35814 , \35813 );
buf \U$30174 ( \35815 , \35814 );
and \U$30175 ( \35816 , \35646 , \35815 );
and \U$30176 ( \35817 , \35477 , \35816 );
_HMUX ga306 ( \35818_nGa306 , \35410_nGa16d , \35412 , \35817 );
buf \U$30179 ( \35819 , \35412 );
buf \U$30182 ( \35820 , \35415 );
buf \U$30185 ( \35821 , \35418 );
buf \U$30188 ( \35822 , \35422 );
buf \U$30189 ( \35823 , \35426 );
not \U$30190 ( \35824 , \35823 );
buf \U$30191 ( \35825 , \35824 );
not \U$30192 ( \35826 , \35825 );
buf \U$30193 ( \35827 , \35429 );
xnor \U$30194 ( \35828 , \35827 , \35823 );
buf \U$30195 ( \35829 , \35828 );
or \U$30196 ( \35830 , \35827 , \35823 );
not \U$30197 ( \35831 , \35830 );
buf \U$30198 ( \35832 , \35831 );
buf \U$30199 ( \35833 , \35832 );
buf \U$30200 ( \35834 , \35832 );
buf \U$30201 ( \35835 , \35832 );
buf \U$30202 ( \35836 , \35832 );
buf \U$30203 ( \35837 , \35832 );
buf \U$30204 ( \35838 , \35832 );
buf \U$30205 ( \35839 , \35832 );
buf \U$30206 ( \35840 , \35832 );
buf \U$30207 ( \35841 , \35832 );
buf \U$30208 ( \35842 , \35832 );
buf \U$30209 ( \35843 , \35832 );
buf \U$30210 ( \35844 , \35832 );
buf \U$30211 ( \35845 , \35832 );
buf \U$30212 ( \35846 , \35832 );
buf \U$30213 ( \35847 , \35832 );
buf \U$30214 ( \35848 , \35832 );
buf \U$30215 ( \35849 , \35832 );
buf \U$30216 ( \35850 , \35832 );
buf \U$30217 ( \35851 , \35832 );
buf \U$30218 ( \35852 , \35832 );
buf \U$30219 ( \35853 , \35832 );
buf \U$30220 ( \35854 , \35832 );
buf \U$30221 ( \35855 , \35832 );
buf \U$30222 ( \35856 , \35832 );
buf \U$30223 ( \35857 , \35832 );
nor \U$30224 ( \35858 , \35819 , \35820 , \35821 , \35822 , \35826 , \35829 , \35832 , \35833 , \35834 , \35835 , \35836 , \35837 , \35838 , \35839 , \35840 , \35841 , \35842 , \35843 , \35844 , \35845 , \35846 , \35847 , \35848 , \35849 , \35850 , \35851 , \35852 , \35853 , \35854 , \35855 , \35856 , \35857 );
and \U$30225 ( \35859 , RIe5329d0_6883, \35858 );
not \U$30226 ( \35860 , \35819 );
not \U$30227 ( \35861 , \35820 );
not \U$30228 ( \35862 , \35821 );
not \U$30229 ( \35863 , \35822 );
buf \U$30230 ( \35864 , \35832 );
buf \U$30231 ( \35865 , \35832 );
buf \U$30232 ( \35866 , \35832 );
buf \U$30233 ( \35867 , \35832 );
buf \U$30234 ( \35868 , \35832 );
buf \U$30235 ( \35869 , \35832 );
buf \U$30236 ( \35870 , \35832 );
buf \U$30237 ( \35871 , \35832 );
buf \U$30238 ( \35872 , \35832 );
buf \U$30239 ( \35873 , \35832 );
buf \U$30240 ( \35874 , \35832 );
buf \U$30241 ( \35875 , \35832 );
buf \U$30242 ( \35876 , \35832 );
buf \U$30243 ( \35877 , \35832 );
buf \U$30244 ( \35878 , \35832 );
buf \U$30245 ( \35879 , \35832 );
buf \U$30246 ( \35880 , \35832 );
buf \U$30247 ( \35881 , \35832 );
buf \U$30248 ( \35882 , \35832 );
buf \U$30249 ( \35883 , \35832 );
buf \U$30250 ( \35884 , \35832 );
buf \U$30251 ( \35885 , \35832 );
buf \U$30252 ( \35886 , \35832 );
buf \U$30253 ( \35887 , \35832 );
buf \U$30254 ( \35888 , \35832 );
nor \U$30255 ( \35889 , \35860 , \35861 , \35862 , \35863 , \35825 , \35829 , \35832 , \35864 , \35865 , \35866 , \35867 , \35868 , \35869 , \35870 , \35871 , \35872 , \35873 , \35874 , \35875 , \35876 , \35877 , \35878 , \35879 , \35880 , \35881 , \35882 , \35883 , \35884 , \35885 , \35886 , \35887 , \35888 );
and \U$30256 ( \35890 , RIeb72150_6905, \35889 );
buf \U$30257 ( \35891 , \35832 );
buf \U$30258 ( \35892 , \35832 );
buf \U$30259 ( \35893 , \35832 );
buf \U$30260 ( \35894 , \35832 );
buf \U$30261 ( \35895 , \35832 );
buf \U$30262 ( \35896 , \35832 );
buf \U$30263 ( \35897 , \35832 );
buf \U$30264 ( \35898 , \35832 );
buf \U$30265 ( \35899 , \35832 );
buf \U$30266 ( \35900 , \35832 );
buf \U$30267 ( \35901 , \35832 );
buf \U$30268 ( \35902 , \35832 );
buf \U$30269 ( \35903 , \35832 );
buf \U$30270 ( \35904 , \35832 );
buf \U$30271 ( \35905 , \35832 );
buf \U$30272 ( \35906 , \35832 );
buf \U$30273 ( \35907 , \35832 );
buf \U$30274 ( \35908 , \35832 );
buf \U$30275 ( \35909 , \35832 );
buf \U$30276 ( \35910 , \35832 );
buf \U$30277 ( \35911 , \35832 );
buf \U$30278 ( \35912 , \35832 );
buf \U$30279 ( \35913 , \35832 );
buf \U$30280 ( \35914 , \35832 );
buf \U$30281 ( \35915 , \35832 );
nor \U$30282 ( \35916 , \35819 , \35861 , \35862 , \35863 , \35825 , \35829 , \35832 , \35891 , \35892 , \35893 , \35894 , \35895 , \35896 , \35897 , \35898 , \35899 , \35900 , \35901 , \35902 , \35903 , \35904 , \35905 , \35906 , \35907 , \35908 , \35909 , \35910 , \35911 , \35912 , \35913 , \35914 , \35915 );
and \U$30283 ( \35917 , RIeab80c0_6897, \35916 );
buf \U$30284 ( \35918 , \35832 );
buf \U$30285 ( \35919 , \35832 );
buf \U$30286 ( \35920 , \35832 );
buf \U$30287 ( \35921 , \35832 );
buf \U$30288 ( \35922 , \35832 );
buf \U$30289 ( \35923 , \35832 );
buf \U$30290 ( \35924 , \35832 );
buf \U$30291 ( \35925 , \35832 );
buf \U$30292 ( \35926 , \35832 );
buf \U$30293 ( \35927 , \35832 );
buf \U$30294 ( \35928 , \35832 );
buf \U$30295 ( \35929 , \35832 );
buf \U$30296 ( \35930 , \35832 );
buf \U$30297 ( \35931 , \35832 );
buf \U$30298 ( \35932 , \35832 );
buf \U$30299 ( \35933 , \35832 );
buf \U$30300 ( \35934 , \35832 );
buf \U$30301 ( \35935 , \35832 );
buf \U$30302 ( \35936 , \35832 );
buf \U$30303 ( \35937 , \35832 );
buf \U$30304 ( \35938 , \35832 );
buf \U$30305 ( \35939 , \35832 );
buf \U$30306 ( \35940 , \35832 );
buf \U$30307 ( \35941 , \35832 );
buf \U$30308 ( \35942 , \35832 );
nor \U$30309 ( \35943 , \35860 , \35820 , \35862 , \35863 , \35825 , \35829 , \35832 , \35918 , \35919 , \35920 , \35921 , \35922 , \35923 , \35924 , \35925 , \35926 , \35927 , \35928 , \35929 , \35930 , \35931 , \35932 , \35933 , \35934 , \35935 , \35936 , \35937 , \35938 , \35939 , \35940 , \35941 , \35942 );
and \U$30310 ( \35944 , RIe5331c8_6882, \35943 );
buf \U$30311 ( \35945 , \35832 );
buf \U$30312 ( \35946 , \35832 );
buf \U$30313 ( \35947 , \35832 );
buf \U$30314 ( \35948 , \35832 );
buf \U$30315 ( \35949 , \35832 );
buf \U$30316 ( \35950 , \35832 );
buf \U$30317 ( \35951 , \35832 );
buf \U$30318 ( \35952 , \35832 );
buf \U$30319 ( \35953 , \35832 );
buf \U$30320 ( \35954 , \35832 );
buf \U$30321 ( \35955 , \35832 );
buf \U$30322 ( \35956 , \35832 );
buf \U$30323 ( \35957 , \35832 );
buf \U$30324 ( \35958 , \35832 );
buf \U$30325 ( \35959 , \35832 );
buf \U$30326 ( \35960 , \35832 );
buf \U$30327 ( \35961 , \35832 );
buf \U$30328 ( \35962 , \35832 );
buf \U$30329 ( \35963 , \35832 );
buf \U$30330 ( \35964 , \35832 );
buf \U$30331 ( \35965 , \35832 );
buf \U$30332 ( \35966 , \35832 );
buf \U$30333 ( \35967 , \35832 );
buf \U$30334 ( \35968 , \35832 );
buf \U$30335 ( \35969 , \35832 );
nor \U$30336 ( \35970 , \35819 , \35820 , \35862 , \35863 , \35825 , \35829 , \35832 , \35945 , \35946 , \35947 , \35948 , \35949 , \35950 , \35951 , \35952 , \35953 , \35954 , \35955 , \35956 , \35957 , \35958 , \35959 , \35960 , \35961 , \35962 , \35963 , \35964 , \35965 , \35966 , \35967 , \35968 , \35969 );
and \U$30337 ( \35971 , RIe5339c0_6881, \35970 );
buf \U$30338 ( \35972 , \35832 );
buf \U$30339 ( \35973 , \35832 );
buf \U$30340 ( \35974 , \35832 );
buf \U$30341 ( \35975 , \35832 );
buf \U$30342 ( \35976 , \35832 );
buf \U$30343 ( \35977 , \35832 );
buf \U$30344 ( \35978 , \35832 );
buf \U$30345 ( \35979 , \35832 );
buf \U$30346 ( \35980 , \35832 );
buf \U$30347 ( \35981 , \35832 );
buf \U$30348 ( \35982 , \35832 );
buf \U$30349 ( \35983 , \35832 );
buf \U$30350 ( \35984 , \35832 );
buf \U$30351 ( \35985 , \35832 );
buf \U$30352 ( \35986 , \35832 );
buf \U$30353 ( \35987 , \35832 );
buf \U$30354 ( \35988 , \35832 );
buf \U$30355 ( \35989 , \35832 );
buf \U$30356 ( \35990 , \35832 );
buf \U$30357 ( \35991 , \35832 );
buf \U$30358 ( \35992 , \35832 );
buf \U$30359 ( \35993 , \35832 );
buf \U$30360 ( \35994 , \35832 );
buf \U$30361 ( \35995 , \35832 );
buf \U$30362 ( \35996 , \35832 );
nor \U$30363 ( \35997 , \35860 , \35861 , \35821 , \35863 , \35825 , \35829 , \35832 , \35972 , \35973 , \35974 , \35975 , \35976 , \35977 , \35978 , \35979 , \35980 , \35981 , \35982 , \35983 , \35984 , \35985 , \35986 , \35987 , \35988 , \35989 , \35990 , \35991 , \35992 , \35993 , \35994 , \35995 , \35996 );
and \U$30364 ( \35998 , RIeab87c8_6898, \35997 );
buf \U$30365 ( \35999 , \35832 );
buf \U$30366 ( \36000 , \35832 );
buf \U$30367 ( \36001 , \35832 );
buf \U$30368 ( \36002 , \35832 );
buf \U$30369 ( \36003 , \35832 );
buf \U$30370 ( \36004 , \35832 );
buf \U$30371 ( \36005 , \35832 );
buf \U$30372 ( \36006 , \35832 );
buf \U$30373 ( \36007 , \35832 );
buf \U$30374 ( \36008 , \35832 );
buf \U$30375 ( \36009 , \35832 );
buf \U$30376 ( \36010 , \35832 );
buf \U$30377 ( \36011 , \35832 );
buf \U$30378 ( \36012 , \35832 );
buf \U$30379 ( \36013 , \35832 );
buf \U$30380 ( \36014 , \35832 );
buf \U$30381 ( \36015 , \35832 );
buf \U$30382 ( \36016 , \35832 );
buf \U$30383 ( \36017 , \35832 );
buf \U$30384 ( \36018 , \35832 );
buf \U$30385 ( \36019 , \35832 );
buf \U$30386 ( \36020 , \35832 );
buf \U$30387 ( \36021 , \35832 );
buf \U$30388 ( \36022 , \35832 );
buf \U$30389 ( \36023 , \35832 );
nor \U$30390 ( \36024 , \35819 , \35861 , \35821 , \35863 , \35825 , \35829 , \35832 , \35999 , \36000 , \36001 , \36002 , \36003 , \36004 , \36005 , \36006 , \36007 , \36008 , \36009 , \36010 , \36011 , \36012 , \36013 , \36014 , \36015 , \36016 , \36017 , \36018 , \36019 , \36020 , \36021 , \36022 , \36023 );
and \U$30391 ( \36025 , RIe5341b8_6880, \36024 );
buf \U$30392 ( \36026 , \35832 );
buf \U$30393 ( \36027 , \35832 );
buf \U$30394 ( \36028 , \35832 );
buf \U$30395 ( \36029 , \35832 );
buf \U$30396 ( \36030 , \35832 );
buf \U$30397 ( \36031 , \35832 );
buf \U$30398 ( \36032 , \35832 );
buf \U$30399 ( \36033 , \35832 );
buf \U$30400 ( \36034 , \35832 );
buf \U$30401 ( \36035 , \35832 );
buf \U$30402 ( \36036 , \35832 );
buf \U$30403 ( \36037 , \35832 );
buf \U$30404 ( \36038 , \35832 );
buf \U$30405 ( \36039 , \35832 );
buf \U$30406 ( \36040 , \35832 );
buf \U$30407 ( \36041 , \35832 );
buf \U$30408 ( \36042 , \35832 );
buf \U$30409 ( \36043 , \35832 );
buf \U$30410 ( \36044 , \35832 );
buf \U$30411 ( \36045 , \35832 );
buf \U$30412 ( \36046 , \35832 );
buf \U$30413 ( \36047 , \35832 );
buf \U$30414 ( \36048 , \35832 );
buf \U$30415 ( \36049 , \35832 );
buf \U$30416 ( \36050 , \35832 );
nor \U$30417 ( \36051 , \35860 , \35820 , \35821 , \35863 , \35825 , \35829 , \35832 , \36026 , \36027 , \36028 , \36029 , \36030 , \36031 , \36032 , \36033 , \36034 , \36035 , \36036 , \36037 , \36038 , \36039 , \36040 , \36041 , \36042 , \36043 , \36044 , \36045 , \36046 , \36047 , \36048 , \36049 , \36050 );
and \U$30418 ( \36052 , RIe5349b0_6879, \36051 );
buf \U$30419 ( \36053 , \35832 );
buf \U$30420 ( \36054 , \35832 );
buf \U$30421 ( \36055 , \35832 );
buf \U$30422 ( \36056 , \35832 );
buf \U$30423 ( \36057 , \35832 );
buf \U$30424 ( \36058 , \35832 );
buf \U$30425 ( \36059 , \35832 );
buf \U$30426 ( \36060 , \35832 );
buf \U$30427 ( \36061 , \35832 );
buf \U$30428 ( \36062 , \35832 );
buf \U$30429 ( \36063 , \35832 );
buf \U$30430 ( \36064 , \35832 );
buf \U$30431 ( \36065 , \35832 );
buf \U$30432 ( \36066 , \35832 );
buf \U$30433 ( \36067 , \35832 );
buf \U$30434 ( \36068 , \35832 );
buf \U$30435 ( \36069 , \35832 );
buf \U$30436 ( \36070 , \35832 );
buf \U$30437 ( \36071 , \35832 );
buf \U$30438 ( \36072 , \35832 );
buf \U$30439 ( \36073 , \35832 );
buf \U$30440 ( \36074 , \35832 );
buf \U$30441 ( \36075 , \35832 );
buf \U$30442 ( \36076 , \35832 );
buf \U$30443 ( \36077 , \35832 );
nor \U$30444 ( \36078 , \35819 , \35820 , \35821 , \35863 , \35825 , \35829 , \35832 , \36053 , \36054 , \36055 , \36056 , \36057 , \36058 , \36059 , \36060 , \36061 , \36062 , \36063 , \36064 , \36065 , \36066 , \36067 , \36068 , \36069 , \36070 , \36071 , \36072 , \36073 , \36074 , \36075 , \36076 , \36077 );
and \U$30445 ( \36079 , RIea94af8_6890, \36078 );
buf \U$30446 ( \36080 , \35832 );
buf \U$30447 ( \36081 , \35832 );
buf \U$30448 ( \36082 , \35832 );
buf \U$30449 ( \36083 , \35832 );
buf \U$30450 ( \36084 , \35832 );
buf \U$30451 ( \36085 , \35832 );
buf \U$30452 ( \36086 , \35832 );
buf \U$30453 ( \36087 , \35832 );
buf \U$30454 ( \36088 , \35832 );
buf \U$30455 ( \36089 , \35832 );
buf \U$30456 ( \36090 , \35832 );
buf \U$30457 ( \36091 , \35832 );
buf \U$30458 ( \36092 , \35832 );
buf \U$30459 ( \36093 , \35832 );
buf \U$30460 ( \36094 , \35832 );
buf \U$30461 ( \36095 , \35832 );
buf \U$30462 ( \36096 , \35832 );
buf \U$30463 ( \36097 , \35832 );
buf \U$30464 ( \36098 , \35832 );
buf \U$30465 ( \36099 , \35832 );
buf \U$30466 ( \36100 , \35832 );
buf \U$30467 ( \36101 , \35832 );
buf \U$30468 ( \36102 , \35832 );
buf \U$30469 ( \36103 , \35832 );
buf \U$30470 ( \36104 , \35832 );
nor \U$30471 ( \36105 , \35860 , \35861 , \35862 , \35822 , \35825 , \35829 , \35832 , \36080 , \36081 , \36082 , \36083 , \36084 , \36085 , \36086 , \36087 , \36088 , \36089 , \36090 , \36091 , \36092 , \36093 , \36094 , \36095 , \36096 , \36097 , \36098 , \36099 , \36100 , \36101 , \36102 , \36103 , \36104 );
and \U$30472 ( \36106 , RIe5351a8_6878, \36105 );
buf \U$30473 ( \36107 , \35832 );
buf \U$30474 ( \36108 , \35832 );
buf \U$30475 ( \36109 , \35832 );
buf \U$30476 ( \36110 , \35832 );
buf \U$30477 ( \36111 , \35832 );
buf \U$30478 ( \36112 , \35832 );
buf \U$30479 ( \36113 , \35832 );
buf \U$30480 ( \36114 , \35832 );
buf \U$30481 ( \36115 , \35832 );
buf \U$30482 ( \36116 , \35832 );
buf \U$30483 ( \36117 , \35832 );
buf \U$30484 ( \36118 , \35832 );
buf \U$30485 ( \36119 , \35832 );
buf \U$30486 ( \36120 , \35832 );
buf \U$30487 ( \36121 , \35832 );
buf \U$30488 ( \36122 , \35832 );
buf \U$30489 ( \36123 , \35832 );
buf \U$30490 ( \36124 , \35832 );
buf \U$30491 ( \36125 , \35832 );
buf \U$30492 ( \36126 , \35832 );
buf \U$30493 ( \36127 , \35832 );
buf \U$30494 ( \36128 , \35832 );
buf \U$30495 ( \36129 , \35832 );
buf \U$30496 ( \36130 , \35832 );
buf \U$30497 ( \36131 , \35832 );
nor \U$30498 ( \36132 , \35819 , \35861 , \35862 , \35822 , \35825 , \35829 , \35832 , \36107 , \36108 , \36109 , \36110 , \36111 , \36112 , \36113 , \36114 , \36115 , \36116 , \36117 , \36118 , \36119 , \36120 , \36121 , \36122 , \36123 , \36124 , \36125 , \36126 , \36127 , \36128 , \36129 , \36130 , \36131 );
and \U$30499 ( \36133 , RIe5359a0_6877, \36132 );
buf \U$30500 ( \36134 , \35832 );
buf \U$30501 ( \36135 , \35832 );
buf \U$30502 ( \36136 , \35832 );
buf \U$30503 ( \36137 , \35832 );
buf \U$30504 ( \36138 , \35832 );
buf \U$30505 ( \36139 , \35832 );
buf \U$30506 ( \36140 , \35832 );
buf \U$30507 ( \36141 , \35832 );
buf \U$30508 ( \36142 , \35832 );
buf \U$30509 ( \36143 , \35832 );
buf \U$30510 ( \36144 , \35832 );
buf \U$30511 ( \36145 , \35832 );
buf \U$30512 ( \36146 , \35832 );
buf \U$30513 ( \36147 , \35832 );
buf \U$30514 ( \36148 , \35832 );
buf \U$30515 ( \36149 , \35832 );
buf \U$30516 ( \36150 , \35832 );
buf \U$30517 ( \36151 , \35832 );
buf \U$30518 ( \36152 , \35832 );
buf \U$30519 ( \36153 , \35832 );
buf \U$30520 ( \36154 , \35832 );
buf \U$30521 ( \36155 , \35832 );
buf \U$30522 ( \36156 , \35832 );
buf \U$30523 ( \36157 , \35832 );
buf \U$30524 ( \36158 , \35832 );
nor \U$30525 ( \36159 , \35860 , \35820 , \35862 , \35822 , \35825 , \35829 , \35832 , \36134 , \36135 , \36136 , \36137 , \36138 , \36139 , \36140 , \36141 , \36142 , \36143 , \36144 , \36145 , \36146 , \36147 , \36148 , \36149 , \36150 , \36151 , \36152 , \36153 , \36154 , \36155 , \36156 , \36157 , \36158 );
and \U$30526 ( \36160 , RIeab78c8_6895, \36159 );
buf \U$30527 ( \36161 , \35832 );
buf \U$30528 ( \36162 , \35832 );
buf \U$30529 ( \36163 , \35832 );
buf \U$30530 ( \36164 , \35832 );
buf \U$30531 ( \36165 , \35832 );
buf \U$30532 ( \36166 , \35832 );
buf \U$30533 ( \36167 , \35832 );
buf \U$30534 ( \36168 , \35832 );
buf \U$30535 ( \36169 , \35832 );
buf \U$30536 ( \36170 , \35832 );
buf \U$30537 ( \36171 , \35832 );
buf \U$30538 ( \36172 , \35832 );
buf \U$30539 ( \36173 , \35832 );
buf \U$30540 ( \36174 , \35832 );
buf \U$30541 ( \36175 , \35832 );
buf \U$30542 ( \36176 , \35832 );
buf \U$30543 ( \36177 , \35832 );
buf \U$30544 ( \36178 , \35832 );
buf \U$30545 ( \36179 , \35832 );
buf \U$30546 ( \36180 , \35832 );
buf \U$30547 ( \36181 , \35832 );
buf \U$30548 ( \36182 , \35832 );
buf \U$30549 ( \36183 , \35832 );
buf \U$30550 ( \36184 , \35832 );
buf \U$30551 ( \36185 , \35832 );
nor \U$30552 ( \36186 , \35819 , \35820 , \35862 , \35822 , \35825 , \35829 , \35832 , \36161 , \36162 , \36163 , \36164 , \36165 , \36166 , \36167 , \36168 , \36169 , \36170 , \36171 , \36172 , \36173 , \36174 , \36175 , \36176 , \36177 , \36178 , \36179 , \36180 , \36181 , \36182 , \36183 , \36184 , \36185 );
and \U$30553 ( \36187 , RIeab7d00_6896, \36186 );
buf \U$30554 ( \36188 , \35832 );
buf \U$30555 ( \36189 , \35832 );
buf \U$30556 ( \36190 , \35832 );
buf \U$30557 ( \36191 , \35832 );
buf \U$30558 ( \36192 , \35832 );
buf \U$30559 ( \36193 , \35832 );
buf \U$30560 ( \36194 , \35832 );
buf \U$30561 ( \36195 , \35832 );
buf \U$30562 ( \36196 , \35832 );
buf \U$30563 ( \36197 , \35832 );
buf \U$30564 ( \36198 , \35832 );
buf \U$30565 ( \36199 , \35832 );
buf \U$30566 ( \36200 , \35832 );
buf \U$30567 ( \36201 , \35832 );
buf \U$30568 ( \36202 , \35832 );
buf \U$30569 ( \36203 , \35832 );
buf \U$30570 ( \36204 , \35832 );
buf \U$30571 ( \36205 , \35832 );
buf \U$30572 ( \36206 , \35832 );
buf \U$30573 ( \36207 , \35832 );
buf \U$30574 ( \36208 , \35832 );
buf \U$30575 ( \36209 , \35832 );
buf \U$30576 ( \36210 , \35832 );
buf \U$30577 ( \36211 , \35832 );
buf \U$30578 ( \36212 , \35832 );
nor \U$30579 ( \36213 , \35860 , \35861 , \35821 , \35822 , \35825 , \35829 , \35832 , \36188 , \36189 , \36190 , \36191 , \36192 , \36193 , \36194 , \36195 , \36196 , \36197 , \36198 , \36199 , \36200 , \36201 , \36202 , \36203 , \36204 , \36205 , \36206 , \36207 , \36208 , \36209 , \36210 , \36211 , \36212 );
and \U$30580 ( \36214 , RIeacfa18_6902, \36213 );
buf \U$30581 ( \36215 , \35832 );
buf \U$30582 ( \36216 , \35832 );
buf \U$30583 ( \36217 , \35832 );
buf \U$30584 ( \36218 , \35832 );
buf \U$30585 ( \36219 , \35832 );
buf \U$30586 ( \36220 , \35832 );
buf \U$30587 ( \36221 , \35832 );
buf \U$30588 ( \36222 , \35832 );
buf \U$30589 ( \36223 , \35832 );
buf \U$30590 ( \36224 , \35832 );
buf \U$30591 ( \36225 , \35832 );
buf \U$30592 ( \36226 , \35832 );
buf \U$30593 ( \36227 , \35832 );
buf \U$30594 ( \36228 , \35832 );
buf \U$30595 ( \36229 , \35832 );
buf \U$30596 ( \36230 , \35832 );
buf \U$30597 ( \36231 , \35832 );
buf \U$30598 ( \36232 , \35832 );
buf \U$30599 ( \36233 , \35832 );
buf \U$30600 ( \36234 , \35832 );
buf \U$30601 ( \36235 , \35832 );
buf \U$30602 ( \36236 , \35832 );
buf \U$30603 ( \36237 , \35832 );
buf \U$30604 ( \36238 , \35832 );
buf \U$30605 ( \36239 , \35832 );
nor \U$30606 ( \36240 , \35819 , \35861 , \35821 , \35822 , \35825 , \35829 , \35832 , \36215 , \36216 , \36217 , \36218 , \36219 , \36220 , \36221 , \36222 , \36223 , \36224 , \36225 , \36226 , \36227 , \36228 , \36229 , \36230 , \36231 , \36232 , \36233 , \36234 , \36235 , \36236 , \36237 , \36238 , \36239 );
and \U$30607 ( \36241 , RIeab6518_6891, \36240 );
buf \U$30608 ( \36242 , \35832 );
buf \U$30609 ( \36243 , \35832 );
buf \U$30610 ( \36244 , \35832 );
buf \U$30611 ( \36245 , \35832 );
buf \U$30612 ( \36246 , \35832 );
buf \U$30613 ( \36247 , \35832 );
buf \U$30614 ( \36248 , \35832 );
buf \U$30615 ( \36249 , \35832 );
buf \U$30616 ( \36250 , \35832 );
buf \U$30617 ( \36251 , \35832 );
buf \U$30618 ( \36252 , \35832 );
buf \U$30619 ( \36253 , \35832 );
buf \U$30620 ( \36254 , \35832 );
buf \U$30621 ( \36255 , \35832 );
buf \U$30622 ( \36256 , \35832 );
buf \U$30623 ( \36257 , \35832 );
buf \U$30624 ( \36258 , \35832 );
buf \U$30625 ( \36259 , \35832 );
buf \U$30626 ( \36260 , \35832 );
buf \U$30627 ( \36261 , \35832 );
buf \U$30628 ( \36262 , \35832 );
buf \U$30629 ( \36263 , \35832 );
buf \U$30630 ( \36264 , \35832 );
buf \U$30631 ( \36265 , \35832 );
buf \U$30632 ( \36266 , \35832 );
nor \U$30633 ( \36267 , \35860 , \35820 , \35821 , \35822 , \35825 , \35829 , \35832 , \36242 , \36243 , \36244 , \36245 , \36246 , \36247 , \36248 , \36249 , \36250 , \36251 , \36252 , \36253 , \36254 , \36255 , \36256 , \36257 , \36258 , \36259 , \36260 , \36261 , \36262 , \36263 , \36264 , \36265 , \36266 );
and \U$30634 ( \36268 , RIeb352c8_6904, \36267 );
or \U$30635 ( \36269 , \35859 , \35890 , \35917 , \35944 , \35971 , \35998 , \36025 , \36052 , \36079 , \36106 , \36133 , \36160 , \36187 , \36214 , \36241 , \36268 );
buf \U$30636 ( \36270 , \35832 );
not \U$30637 ( \36271 , \36270 );
buf \U$30638 ( \36272 , \35820 );
buf \U$30639 ( \36273 , \35821 );
buf \U$30640 ( \36274 , \35822 );
buf \U$30641 ( \36275 , \35825 );
buf \U$30642 ( \36276 , \35829 );
buf \U$30643 ( \36277 , \35832 );
buf \U$30644 ( \36278 , \35832 );
buf \U$30645 ( \36279 , \35832 );
buf \U$30646 ( \36280 , \35832 );
buf \U$30647 ( \36281 , \35832 );
buf \U$30648 ( \36282 , \35832 );
buf \U$30649 ( \36283 , \35832 );
buf \U$30650 ( \36284 , \35832 );
buf \U$30651 ( \36285 , \35832 );
buf \U$30652 ( \36286 , \35832 );
buf \U$30653 ( \36287 , \35832 );
buf \U$30654 ( \36288 , \35832 );
buf \U$30655 ( \36289 , \35832 );
buf \U$30656 ( \36290 , \35832 );
buf \U$30657 ( \36291 , \35832 );
buf \U$30658 ( \36292 , \35832 );
buf \U$30659 ( \36293 , \35832 );
buf \U$30660 ( \36294 , \35832 );
buf \U$30661 ( \36295 , \35832 );
buf \U$30662 ( \36296 , \35832 );
buf \U$30663 ( \36297 , \35832 );
buf \U$30664 ( \36298 , \35832 );
buf \U$30665 ( \36299 , \35832 );
buf \U$30666 ( \36300 , \35832 );
buf \U$30667 ( \36301 , \35832 );
buf \U$30668 ( \36302 , \35819 );
or \U$30669 ( \36303 , \36272 , \36273 , \36274 , \36275 , \36276 , \36277 , \36278 , \36279 , \36280 , \36281 , \36282 , \36283 , \36284 , \36285 , \36286 , \36287 , \36288 , \36289 , \36290 , \36291 , \36292 , \36293 , \36294 , \36295 , \36296 , \36297 , \36298 , \36299 , \36300 , \36301 , \36302 );
nand \U$30670 ( \36304 , \36271 , \36303 );
buf \U$30671 ( \36305 , \36304 );
buf \U$30672 ( \36306 , \35832 );
not \U$30673 ( \36307 , \36306 );
buf \U$30674 ( \36308 , \35829 );
buf \U$30675 ( \36309 , \35832 );
buf \U$30676 ( \36310 , \35832 );
buf \U$30677 ( \36311 , \35832 );
buf \U$30678 ( \36312 , \35832 );
buf \U$30679 ( \36313 , \35832 );
buf \U$30680 ( \36314 , \35832 );
buf \U$30681 ( \36315 , \35832 );
buf \U$30682 ( \36316 , \35832 );
buf \U$30683 ( \36317 , \35832 );
buf \U$30684 ( \36318 , \35832 );
buf \U$30685 ( \36319 , \35832 );
buf \U$30686 ( \36320 , \35832 );
buf \U$30687 ( \36321 , \35832 );
buf \U$30688 ( \36322 , \35832 );
buf \U$30689 ( \36323 , \35832 );
buf \U$30690 ( \36324 , \35832 );
buf \U$30691 ( \36325 , \35832 );
buf \U$30692 ( \36326 , \35832 );
buf \U$30693 ( \36327 , \35832 );
buf \U$30694 ( \36328 , \35832 );
buf \U$30695 ( \36329 , \35832 );
buf \U$30696 ( \36330 , \35832 );
buf \U$30697 ( \36331 , \35832 );
buf \U$30698 ( \36332 , \35832 );
buf \U$30699 ( \36333 , \35832 );
buf \U$30700 ( \36334 , \35825 );
buf \U$30701 ( \36335 , \35819 );
buf \U$30702 ( \36336 , \35820 );
buf \U$30703 ( \36337 , \35821 );
buf \U$30704 ( \36338 , \35822 );
or \U$30705 ( \36339 , \36335 , \36336 , \36337 , \36338 );
and \U$30706 ( \36340 , \36334 , \36339 );
or \U$30707 ( \36341 , \36308 , \36309 , \36310 , \36311 , \36312 , \36313 , \36314 , \36315 , \36316 , \36317 , \36318 , \36319 , \36320 , \36321 , \36322 , \36323 , \36324 , \36325 , \36326 , \36327 , \36328 , \36329 , \36330 , \36331 , \36332 , \36333 , \36340 );
and \U$30708 ( \36342 , \36307 , \36341 );
buf \U$30709 ( \36343 , \36342 );
or \U$30710 ( \36344 , \36305 , \36343 );
_DC ga51d ( \36345_nGa51d , \36269 , \36344 );
not \U$30711 ( \36346 , \36345_nGa51d );
buf \U$30712 ( \36347 , RIb7b9608_246);
buf \U$30713 ( \36348 , \35832 );
buf \U$30714 ( \36349 , \35832 );
buf \U$30715 ( \36350 , \35832 );
buf \U$30716 ( \36351 , \35832 );
buf \U$30717 ( \36352 , \35832 );
buf \U$30718 ( \36353 , \35832 );
buf \U$30719 ( \36354 , \35832 );
buf \U$30720 ( \36355 , \35832 );
buf \U$30721 ( \36356 , \35832 );
buf \U$30722 ( \36357 , \35832 );
buf \U$30723 ( \36358 , \35832 );
buf \U$30724 ( \36359 , \35832 );
buf \U$30725 ( \36360 , \35832 );
buf \U$30726 ( \36361 , \35832 );
buf \U$30727 ( \36362 , \35832 );
buf \U$30728 ( \36363 , \35832 );
buf \U$30729 ( \36364 , \35832 );
buf \U$30730 ( \36365 , \35832 );
buf \U$30731 ( \36366 , \35832 );
buf \U$30732 ( \36367 , \35832 );
buf \U$30733 ( \36368 , \35832 );
buf \U$30734 ( \36369 , \35832 );
buf \U$30735 ( \36370 , \35832 );
buf \U$30736 ( \36371 , \35832 );
buf \U$30737 ( \36372 , \35832 );
nor \U$30738 ( \36373 , \35819 , \35820 , \35821 , \35822 , \35826 , \35829 , \35832 , \36348 , \36349 , \36350 , \36351 , \36352 , \36353 , \36354 , \36355 , \36356 , \36357 , \36358 , \36359 , \36360 , \36361 , \36362 , \36363 , \36364 , \36365 , \36366 , \36367 , \36368 , \36369 , \36370 , \36371 , \36372 );
and \U$30739 ( \36374 , \7117 , \36373 );
buf \U$30740 ( \36375 , \35832 );
buf \U$30741 ( \36376 , \35832 );
buf \U$30742 ( \36377 , \35832 );
buf \U$30743 ( \36378 , \35832 );
buf \U$30744 ( \36379 , \35832 );
buf \U$30745 ( \36380 , \35832 );
buf \U$30746 ( \36381 , \35832 );
buf \U$30747 ( \36382 , \35832 );
buf \U$30748 ( \36383 , \35832 );
buf \U$30749 ( \36384 , \35832 );
buf \U$30750 ( \36385 , \35832 );
buf \U$30751 ( \36386 , \35832 );
buf \U$30752 ( \36387 , \35832 );
buf \U$30753 ( \36388 , \35832 );
buf \U$30754 ( \36389 , \35832 );
buf \U$30755 ( \36390 , \35832 );
buf \U$30756 ( \36391 , \35832 );
buf \U$30757 ( \36392 , \35832 );
buf \U$30758 ( \36393 , \35832 );
buf \U$30759 ( \36394 , \35832 );
buf \U$30760 ( \36395 , \35832 );
buf \U$30761 ( \36396 , \35832 );
buf \U$30762 ( \36397 , \35832 );
buf \U$30763 ( \36398 , \35832 );
buf \U$30764 ( \36399 , \35832 );
nor \U$30765 ( \36400 , \35860 , \35861 , \35862 , \35863 , \35825 , \35829 , \35832 , \36375 , \36376 , \36377 , \36378 , \36379 , \36380 , \36381 , \36382 , \36383 , \36384 , \36385 , \36386 , \36387 , \36388 , \36389 , \36390 , \36391 , \36392 , \36393 , \36394 , \36395 , \36396 , \36397 , \36398 , \36399 );
and \U$30766 ( \36401 , \7119 , \36400 );
buf \U$30767 ( \36402 , \35832 );
buf \U$30768 ( \36403 , \35832 );
buf \U$30769 ( \36404 , \35832 );
buf \U$30770 ( \36405 , \35832 );
buf \U$30771 ( \36406 , \35832 );
buf \U$30772 ( \36407 , \35832 );
buf \U$30773 ( \36408 , \35832 );
buf \U$30774 ( \36409 , \35832 );
buf \U$30775 ( \36410 , \35832 );
buf \U$30776 ( \36411 , \35832 );
buf \U$30777 ( \36412 , \35832 );
buf \U$30778 ( \36413 , \35832 );
buf \U$30779 ( \36414 , \35832 );
buf \U$30780 ( \36415 , \35832 );
buf \U$30781 ( \36416 , \35832 );
buf \U$30782 ( \36417 , \35832 );
buf \U$30783 ( \36418 , \35832 );
buf \U$30784 ( \36419 , \35832 );
buf \U$30785 ( \36420 , \35832 );
buf \U$30786 ( \36421 , \35832 );
buf \U$30787 ( \36422 , \35832 );
buf \U$30788 ( \36423 , \35832 );
buf \U$30789 ( \36424 , \35832 );
buf \U$30790 ( \36425 , \35832 );
buf \U$30791 ( \36426 , \35832 );
nor \U$30792 ( \36427 , \35819 , \35861 , \35862 , \35863 , \35825 , \35829 , \35832 , \36402 , \36403 , \36404 , \36405 , \36406 , \36407 , \36408 , \36409 , \36410 , \36411 , \36412 , \36413 , \36414 , \36415 , \36416 , \36417 , \36418 , \36419 , \36420 , \36421 , \36422 , \36423 , \36424 , \36425 , \36426 );
and \U$30793 ( \36428 , \7864 , \36427 );
buf \U$30794 ( \36429 , \35832 );
buf \U$30795 ( \36430 , \35832 );
buf \U$30796 ( \36431 , \35832 );
buf \U$30797 ( \36432 , \35832 );
buf \U$30798 ( \36433 , \35832 );
buf \U$30799 ( \36434 , \35832 );
buf \U$30800 ( \36435 , \35832 );
buf \U$30801 ( \36436 , \35832 );
buf \U$30802 ( \36437 , \35832 );
buf \U$30803 ( \36438 , \35832 );
buf \U$30804 ( \36439 , \35832 );
buf \U$30805 ( \36440 , \35832 );
buf \U$30806 ( \36441 , \35832 );
buf \U$30807 ( \36442 , \35832 );
buf \U$30808 ( \36443 , \35832 );
buf \U$30809 ( \36444 , \35832 );
buf \U$30810 ( \36445 , \35832 );
buf \U$30811 ( \36446 , \35832 );
buf \U$30812 ( \36447 , \35832 );
buf \U$30813 ( \36448 , \35832 );
buf \U$30814 ( \36449 , \35832 );
buf \U$30815 ( \36450 , \35832 );
buf \U$30816 ( \36451 , \35832 );
buf \U$30817 ( \36452 , \35832 );
buf \U$30818 ( \36453 , \35832 );
nor \U$30819 ( \36454 , \35860 , \35820 , \35862 , \35863 , \35825 , \35829 , \35832 , \36429 , \36430 , \36431 , \36432 , \36433 , \36434 , \36435 , \36436 , \36437 , \36438 , \36439 , \36440 , \36441 , \36442 , \36443 , \36444 , \36445 , \36446 , \36447 , \36448 , \36449 , \36450 , \36451 , \36452 , \36453 );
and \U$30820 ( \36455 , \7892 , \36454 );
buf \U$30821 ( \36456 , \35832 );
buf \U$30822 ( \36457 , \35832 );
buf \U$30823 ( \36458 , \35832 );
buf \U$30824 ( \36459 , \35832 );
buf \U$30825 ( \36460 , \35832 );
buf \U$30826 ( \36461 , \35832 );
buf \U$30827 ( \36462 , \35832 );
buf \U$30828 ( \36463 , \35832 );
buf \U$30829 ( \36464 , \35832 );
buf \U$30830 ( \36465 , \35832 );
buf \U$30831 ( \36466 , \35832 );
buf \U$30832 ( \36467 , \35832 );
buf \U$30833 ( \36468 , \35832 );
buf \U$30834 ( \36469 , \35832 );
buf \U$30835 ( \36470 , \35832 );
buf \U$30836 ( \36471 , \35832 );
buf \U$30837 ( \36472 , \35832 );
buf \U$30838 ( \36473 , \35832 );
buf \U$30839 ( \36474 , \35832 );
buf \U$30840 ( \36475 , \35832 );
buf \U$30841 ( \36476 , \35832 );
buf \U$30842 ( \36477 , \35832 );
buf \U$30843 ( \36478 , \35832 );
buf \U$30844 ( \36479 , \35832 );
buf \U$30845 ( \36480 , \35832 );
nor \U$30846 ( \36481 , \35819 , \35820 , \35862 , \35863 , \35825 , \35829 , \35832 , \36456 , \36457 , \36458 , \36459 , \36460 , \36461 , \36462 , \36463 , \36464 , \36465 , \36466 , \36467 , \36468 , \36469 , \36470 , \36471 , \36472 , \36473 , \36474 , \36475 , \36476 , \36477 , \36478 , \36479 , \36480 );
and \U$30847 ( \36482 , \7920 , \36481 );
buf \U$30848 ( \36483 , \35832 );
buf \U$30849 ( \36484 , \35832 );
buf \U$30850 ( \36485 , \35832 );
buf \U$30851 ( \36486 , \35832 );
buf \U$30852 ( \36487 , \35832 );
buf \U$30853 ( \36488 , \35832 );
buf \U$30854 ( \36489 , \35832 );
buf \U$30855 ( \36490 , \35832 );
buf \U$30856 ( \36491 , \35832 );
buf \U$30857 ( \36492 , \35832 );
buf \U$30858 ( \36493 , \35832 );
buf \U$30859 ( \36494 , \35832 );
buf \U$30860 ( \36495 , \35832 );
buf \U$30861 ( \36496 , \35832 );
buf \U$30862 ( \36497 , \35832 );
buf \U$30863 ( \36498 , \35832 );
buf \U$30864 ( \36499 , \35832 );
buf \U$30865 ( \36500 , \35832 );
buf \U$30866 ( \36501 , \35832 );
buf \U$30867 ( \36502 , \35832 );
buf \U$30868 ( \36503 , \35832 );
buf \U$30869 ( \36504 , \35832 );
buf \U$30870 ( \36505 , \35832 );
buf \U$30871 ( \36506 , \35832 );
buf \U$30872 ( \36507 , \35832 );
nor \U$30873 ( \36508 , \35860 , \35861 , \35821 , \35863 , \35825 , \35829 , \35832 , \36483 , \36484 , \36485 , \36486 , \36487 , \36488 , \36489 , \36490 , \36491 , \36492 , \36493 , \36494 , \36495 , \36496 , \36497 , \36498 , \36499 , \36500 , \36501 , \36502 , \36503 , \36504 , \36505 , \36506 , \36507 );
and \U$30874 ( \36509 , \7948 , \36508 );
buf \U$30875 ( \36510 , \35832 );
buf \U$30876 ( \36511 , \35832 );
buf \U$30877 ( \36512 , \35832 );
buf \U$30878 ( \36513 , \35832 );
buf \U$30879 ( \36514 , \35832 );
buf \U$30880 ( \36515 , \35832 );
buf \U$30881 ( \36516 , \35832 );
buf \U$30882 ( \36517 , \35832 );
buf \U$30883 ( \36518 , \35832 );
buf \U$30884 ( \36519 , \35832 );
buf \U$30885 ( \36520 , \35832 );
buf \U$30886 ( \36521 , \35832 );
buf \U$30887 ( \36522 , \35832 );
buf \U$30888 ( \36523 , \35832 );
buf \U$30889 ( \36524 , \35832 );
buf \U$30890 ( \36525 , \35832 );
buf \U$30891 ( \36526 , \35832 );
buf \U$30892 ( \36527 , \35832 );
buf \U$30893 ( \36528 , \35832 );
buf \U$30894 ( \36529 , \35832 );
buf \U$30895 ( \36530 , \35832 );
buf \U$30896 ( \36531 , \35832 );
buf \U$30897 ( \36532 , \35832 );
buf \U$30898 ( \36533 , \35832 );
buf \U$30899 ( \36534 , \35832 );
nor \U$30900 ( \36535 , \35819 , \35861 , \35821 , \35863 , \35825 , \35829 , \35832 , \36510 , \36511 , \36512 , \36513 , \36514 , \36515 , \36516 , \36517 , \36518 , \36519 , \36520 , \36521 , \36522 , \36523 , \36524 , \36525 , \36526 , \36527 , \36528 , \36529 , \36530 , \36531 , \36532 , \36533 , \36534 );
and \U$30901 ( \36536 , \7976 , \36535 );
buf \U$30902 ( \36537 , \35832 );
buf \U$30903 ( \36538 , \35832 );
buf \U$30904 ( \36539 , \35832 );
buf \U$30905 ( \36540 , \35832 );
buf \U$30906 ( \36541 , \35832 );
buf \U$30907 ( \36542 , \35832 );
buf \U$30908 ( \36543 , \35832 );
buf \U$30909 ( \36544 , \35832 );
buf \U$30910 ( \36545 , \35832 );
buf \U$30911 ( \36546 , \35832 );
buf \U$30912 ( \36547 , \35832 );
buf \U$30913 ( \36548 , \35832 );
buf \U$30914 ( \36549 , \35832 );
buf \U$30915 ( \36550 , \35832 );
buf \U$30916 ( \36551 , \35832 );
buf \U$30917 ( \36552 , \35832 );
buf \U$30918 ( \36553 , \35832 );
buf \U$30919 ( \36554 , \35832 );
buf \U$30920 ( \36555 , \35832 );
buf \U$30921 ( \36556 , \35832 );
buf \U$30922 ( \36557 , \35832 );
buf \U$30923 ( \36558 , \35832 );
buf \U$30924 ( \36559 , \35832 );
buf \U$30925 ( \36560 , \35832 );
buf \U$30926 ( \36561 , \35832 );
nor \U$30927 ( \36562 , \35860 , \35820 , \35821 , \35863 , \35825 , \35829 , \35832 , \36537 , \36538 , \36539 , \36540 , \36541 , \36542 , \36543 , \36544 , \36545 , \36546 , \36547 , \36548 , \36549 , \36550 , \36551 , \36552 , \36553 , \36554 , \36555 , \36556 , \36557 , \36558 , \36559 , \36560 , \36561 );
and \U$30928 ( \36563 , \8004 , \36562 );
buf \U$30929 ( \36564 , \35832 );
buf \U$30930 ( \36565 , \35832 );
buf \U$30931 ( \36566 , \35832 );
buf \U$30932 ( \36567 , \35832 );
buf \U$30933 ( \36568 , \35832 );
buf \U$30934 ( \36569 , \35832 );
buf \U$30935 ( \36570 , \35832 );
buf \U$30936 ( \36571 , \35832 );
buf \U$30937 ( \36572 , \35832 );
buf \U$30938 ( \36573 , \35832 );
buf \U$30939 ( \36574 , \35832 );
buf \U$30940 ( \36575 , \35832 );
buf \U$30941 ( \36576 , \35832 );
buf \U$30942 ( \36577 , \35832 );
buf \U$30943 ( \36578 , \35832 );
buf \U$30944 ( \36579 , \35832 );
buf \U$30945 ( \36580 , \35832 );
buf \U$30946 ( \36581 , \35832 );
buf \U$30947 ( \36582 , \35832 );
buf \U$30948 ( \36583 , \35832 );
buf \U$30949 ( \36584 , \35832 );
buf \U$30950 ( \36585 , \35832 );
buf \U$30951 ( \36586 , \35832 );
buf \U$30952 ( \36587 , \35832 );
buf \U$30953 ( \36588 , \35832 );
nor \U$30954 ( \36589 , \35819 , \35820 , \35821 , \35863 , \35825 , \35829 , \35832 , \36564 , \36565 , \36566 , \36567 , \36568 , \36569 , \36570 , \36571 , \36572 , \36573 , \36574 , \36575 , \36576 , \36577 , \36578 , \36579 , \36580 , \36581 , \36582 , \36583 , \36584 , \36585 , \36586 , \36587 , \36588 );
and \U$30955 ( \36590 , \8032 , \36589 );
buf \U$30956 ( \36591 , \35832 );
buf \U$30957 ( \36592 , \35832 );
buf \U$30958 ( \36593 , \35832 );
buf \U$30959 ( \36594 , \35832 );
buf \U$30960 ( \36595 , \35832 );
buf \U$30961 ( \36596 , \35832 );
buf \U$30962 ( \36597 , \35832 );
buf \U$30963 ( \36598 , \35832 );
buf \U$30964 ( \36599 , \35832 );
buf \U$30965 ( \36600 , \35832 );
buf \U$30966 ( \36601 , \35832 );
buf \U$30967 ( \36602 , \35832 );
buf \U$30968 ( \36603 , \35832 );
buf \U$30969 ( \36604 , \35832 );
buf \U$30970 ( \36605 , \35832 );
buf \U$30971 ( \36606 , \35832 );
buf \U$30972 ( \36607 , \35832 );
buf \U$30973 ( \36608 , \35832 );
buf \U$30974 ( \36609 , \35832 );
buf \U$30975 ( \36610 , \35832 );
buf \U$30976 ( \36611 , \35832 );
buf \U$30977 ( \36612 , \35832 );
buf \U$30978 ( \36613 , \35832 );
buf \U$30979 ( \36614 , \35832 );
buf \U$30980 ( \36615 , \35832 );
nor \U$30981 ( \36616 , \35860 , \35861 , \35862 , \35822 , \35825 , \35829 , \35832 , \36591 , \36592 , \36593 , \36594 , \36595 , \36596 , \36597 , \36598 , \36599 , \36600 , \36601 , \36602 , \36603 , \36604 , \36605 , \36606 , \36607 , \36608 , \36609 , \36610 , \36611 , \36612 , \36613 , \36614 , \36615 );
and \U$30982 ( \36617 , \8060 , \36616 );
buf \U$30983 ( \36618 , \35832 );
buf \U$30984 ( \36619 , \35832 );
buf \U$30985 ( \36620 , \35832 );
buf \U$30986 ( \36621 , \35832 );
buf \U$30987 ( \36622 , \35832 );
buf \U$30988 ( \36623 , \35832 );
buf \U$30989 ( \36624 , \35832 );
buf \U$30990 ( \36625 , \35832 );
buf \U$30991 ( \36626 , \35832 );
buf \U$30992 ( \36627 , \35832 );
buf \U$30993 ( \36628 , \35832 );
buf \U$30994 ( \36629 , \35832 );
buf \U$30995 ( \36630 , \35832 );
buf \U$30996 ( \36631 , \35832 );
buf \U$30997 ( \36632 , \35832 );
buf \U$30998 ( \36633 , \35832 );
buf \U$30999 ( \36634 , \35832 );
buf \U$31000 ( \36635 , \35832 );
buf \U$31001 ( \36636 , \35832 );
buf \U$31002 ( \36637 , \35832 );
buf \U$31003 ( \36638 , \35832 );
buf \U$31004 ( \36639 , \35832 );
buf \U$31005 ( \36640 , \35832 );
buf \U$31006 ( \36641 , \35832 );
buf \U$31007 ( \36642 , \35832 );
nor \U$31008 ( \36643 , \35819 , \35861 , \35862 , \35822 , \35825 , \35829 , \35832 , \36618 , \36619 , \36620 , \36621 , \36622 , \36623 , \36624 , \36625 , \36626 , \36627 , \36628 , \36629 , \36630 , \36631 , \36632 , \36633 , \36634 , \36635 , \36636 , \36637 , \36638 , \36639 , \36640 , \36641 , \36642 );
and \U$31009 ( \36644 , \8088 , \36643 );
buf \U$31010 ( \36645 , \35832 );
buf \U$31011 ( \36646 , \35832 );
buf \U$31012 ( \36647 , \35832 );
buf \U$31013 ( \36648 , \35832 );
buf \U$31014 ( \36649 , \35832 );
buf \U$31015 ( \36650 , \35832 );
buf \U$31016 ( \36651 , \35832 );
buf \U$31017 ( \36652 , \35832 );
buf \U$31018 ( \36653 , \35832 );
buf \U$31019 ( \36654 , \35832 );
buf \U$31020 ( \36655 , \35832 );
buf \U$31021 ( \36656 , \35832 );
buf \U$31022 ( \36657 , \35832 );
buf \U$31023 ( \36658 , \35832 );
buf \U$31024 ( \36659 , \35832 );
buf \U$31025 ( \36660 , \35832 );
buf \U$31026 ( \36661 , \35832 );
buf \U$31027 ( \36662 , \35832 );
buf \U$31028 ( \36663 , \35832 );
buf \U$31029 ( \36664 , \35832 );
buf \U$31030 ( \36665 , \35832 );
buf \U$31031 ( \36666 , \35832 );
buf \U$31032 ( \36667 , \35832 );
buf \U$31033 ( \36668 , \35832 );
buf \U$31034 ( \36669 , \35832 );
nor \U$31035 ( \36670 , \35860 , \35820 , \35862 , \35822 , \35825 , \35829 , \35832 , \36645 , \36646 , \36647 , \36648 , \36649 , \36650 , \36651 , \36652 , \36653 , \36654 , \36655 , \36656 , \36657 , \36658 , \36659 , \36660 , \36661 , \36662 , \36663 , \36664 , \36665 , \36666 , \36667 , \36668 , \36669 );
and \U$31036 ( \36671 , \8116 , \36670 );
buf \U$31037 ( \36672 , \35832 );
buf \U$31038 ( \36673 , \35832 );
buf \U$31039 ( \36674 , \35832 );
buf \U$31040 ( \36675 , \35832 );
buf \U$31041 ( \36676 , \35832 );
buf \U$31042 ( \36677 , \35832 );
buf \U$31043 ( \36678 , \35832 );
buf \U$31044 ( \36679 , \35832 );
buf \U$31045 ( \36680 , \35832 );
buf \U$31046 ( \36681 , \35832 );
buf \U$31047 ( \36682 , \35832 );
buf \U$31048 ( \36683 , \35832 );
buf \U$31049 ( \36684 , \35832 );
buf \U$31050 ( \36685 , \35832 );
buf \U$31051 ( \36686 , \35832 );
buf \U$31052 ( \36687 , \35832 );
buf \U$31053 ( \36688 , \35832 );
buf \U$31054 ( \36689 , \35832 );
buf \U$31055 ( \36690 , \35832 );
buf \U$31056 ( \36691 , \35832 );
buf \U$31057 ( \36692 , \35832 );
buf \U$31058 ( \36693 , \35832 );
buf \U$31059 ( \36694 , \35832 );
buf \U$31060 ( \36695 , \35832 );
buf \U$31061 ( \36696 , \35832 );
nor \U$31062 ( \36697 , \35819 , \35820 , \35862 , \35822 , \35825 , \35829 , \35832 , \36672 , \36673 , \36674 , \36675 , \36676 , \36677 , \36678 , \36679 , \36680 , \36681 , \36682 , \36683 , \36684 , \36685 , \36686 , \36687 , \36688 , \36689 , \36690 , \36691 , \36692 , \36693 , \36694 , \36695 , \36696 );
and \U$31063 ( \36698 , \8144 , \36697 );
buf \U$31064 ( \36699 , \35832 );
buf \U$31065 ( \36700 , \35832 );
buf \U$31066 ( \36701 , \35832 );
buf \U$31067 ( \36702 , \35832 );
buf \U$31068 ( \36703 , \35832 );
buf \U$31069 ( \36704 , \35832 );
buf \U$31070 ( \36705 , \35832 );
buf \U$31071 ( \36706 , \35832 );
buf \U$31072 ( \36707 , \35832 );
buf \U$31073 ( \36708 , \35832 );
buf \U$31074 ( \36709 , \35832 );
buf \U$31075 ( \36710 , \35832 );
buf \U$31076 ( \36711 , \35832 );
buf \U$31077 ( \36712 , \35832 );
buf \U$31078 ( \36713 , \35832 );
buf \U$31079 ( \36714 , \35832 );
buf \U$31080 ( \36715 , \35832 );
buf \U$31081 ( \36716 , \35832 );
buf \U$31082 ( \36717 , \35832 );
buf \U$31083 ( \36718 , \35832 );
buf \U$31084 ( \36719 , \35832 );
buf \U$31085 ( \36720 , \35832 );
buf \U$31086 ( \36721 , \35832 );
buf \U$31087 ( \36722 , \35832 );
buf \U$31088 ( \36723 , \35832 );
nor \U$31089 ( \36724 , \35860 , \35861 , \35821 , \35822 , \35825 , \35829 , \35832 , \36699 , \36700 , \36701 , \36702 , \36703 , \36704 , \36705 , \36706 , \36707 , \36708 , \36709 , \36710 , \36711 , \36712 , \36713 , \36714 , \36715 , \36716 , \36717 , \36718 , \36719 , \36720 , \36721 , \36722 , \36723 );
and \U$31090 ( \36725 , \8172 , \36724 );
buf \U$31091 ( \36726 , \35832 );
buf \U$31092 ( \36727 , \35832 );
buf \U$31093 ( \36728 , \35832 );
buf \U$31094 ( \36729 , \35832 );
buf \U$31095 ( \36730 , \35832 );
buf \U$31096 ( \36731 , \35832 );
buf \U$31097 ( \36732 , \35832 );
buf \U$31098 ( \36733 , \35832 );
buf \U$31099 ( \36734 , \35832 );
buf \U$31100 ( \36735 , \35832 );
buf \U$31101 ( \36736 , \35832 );
buf \U$31102 ( \36737 , \35832 );
buf \U$31103 ( \36738 , \35832 );
buf \U$31104 ( \36739 , \35832 );
buf \U$31105 ( \36740 , \35832 );
buf \U$31106 ( \36741 , \35832 );
buf \U$31107 ( \36742 , \35832 );
buf \U$31108 ( \36743 , \35832 );
buf \U$31109 ( \36744 , \35832 );
buf \U$31110 ( \36745 , \35832 );
buf \U$31111 ( \36746 , \35832 );
buf \U$31112 ( \36747 , \35832 );
buf \U$31113 ( \36748 , \35832 );
buf \U$31114 ( \36749 , \35832 );
buf \U$31115 ( \36750 , \35832 );
nor \U$31116 ( \36751 , \35819 , \35861 , \35821 , \35822 , \35825 , \35829 , \35832 , \36726 , \36727 , \36728 , \36729 , \36730 , \36731 , \36732 , \36733 , \36734 , \36735 , \36736 , \36737 , \36738 , \36739 , \36740 , \36741 , \36742 , \36743 , \36744 , \36745 , \36746 , \36747 , \36748 , \36749 , \36750 );
and \U$31117 ( \36752 , \8200 , \36751 );
buf \U$31118 ( \36753 , \35832 );
buf \U$31119 ( \36754 , \35832 );
buf \U$31120 ( \36755 , \35832 );
buf \U$31121 ( \36756 , \35832 );
buf \U$31122 ( \36757 , \35832 );
buf \U$31123 ( \36758 , \35832 );
buf \U$31124 ( \36759 , \35832 );
buf \U$31125 ( \36760 , \35832 );
buf \U$31126 ( \36761 , \35832 );
buf \U$31127 ( \36762 , \35832 );
buf \U$31128 ( \36763 , \35832 );
buf \U$31129 ( \36764 , \35832 );
buf \U$31130 ( \36765 , \35832 );
buf \U$31131 ( \36766 , \35832 );
buf \U$31132 ( \36767 , \35832 );
buf \U$31133 ( \36768 , \35832 );
buf \U$31134 ( \36769 , \35832 );
buf \U$31135 ( \36770 , \35832 );
buf \U$31136 ( \36771 , \35832 );
buf \U$31137 ( \36772 , \35832 );
buf \U$31138 ( \36773 , \35832 );
buf \U$31139 ( \36774 , \35832 );
buf \U$31140 ( \36775 , \35832 );
buf \U$31141 ( \36776 , \35832 );
buf \U$31142 ( \36777 , \35832 );
nor \U$31143 ( \36778 , \35860 , \35820 , \35821 , \35822 , \35825 , \35829 , \35832 , \36753 , \36754 , \36755 , \36756 , \36757 , \36758 , \36759 , \36760 , \36761 , \36762 , \36763 , \36764 , \36765 , \36766 , \36767 , \36768 , \36769 , \36770 , \36771 , \36772 , \36773 , \36774 , \36775 , \36776 , \36777 );
and \U$31144 ( \36779 , \8228 , \36778 );
or \U$31145 ( \36780 , \36374 , \36401 , \36428 , \36455 , \36482 , \36509 , \36536 , \36563 , \36590 , \36617 , \36644 , \36671 , \36698 , \36725 , \36752 , \36779 );
buf \U$31146 ( \36781 , \35832 );
not \U$31147 ( \36782 , \36781 );
buf \U$31148 ( \36783 , \35820 );
buf \U$31149 ( \36784 , \35821 );
buf \U$31150 ( \36785 , \35822 );
buf \U$31151 ( \36786 , \35825 );
buf \U$31152 ( \36787 , \35829 );
buf \U$31153 ( \36788 , \35832 );
buf \U$31154 ( \36789 , \35832 );
buf \U$31155 ( \36790 , \35832 );
buf \U$31156 ( \36791 , \35832 );
buf \U$31157 ( \36792 , \35832 );
buf \U$31158 ( \36793 , \35832 );
buf \U$31159 ( \36794 , \35832 );
buf \U$31160 ( \36795 , \35832 );
buf \U$31161 ( \36796 , \35832 );
buf \U$31162 ( \36797 , \35832 );
buf \U$31163 ( \36798 , \35832 );
buf \U$31164 ( \36799 , \35832 );
buf \U$31165 ( \36800 , \35832 );
buf \U$31166 ( \36801 , \35832 );
buf \U$31167 ( \36802 , \35832 );
buf \U$31168 ( \36803 , \35832 );
buf \U$31169 ( \36804 , \35832 );
buf \U$31170 ( \36805 , \35832 );
buf \U$31171 ( \36806 , \35832 );
buf \U$31172 ( \36807 , \35832 );
buf \U$31173 ( \36808 , \35832 );
buf \U$31174 ( \36809 , \35832 );
buf \U$31175 ( \36810 , \35832 );
buf \U$31176 ( \36811 , \35832 );
buf \U$31177 ( \36812 , \35832 );
buf \U$31178 ( \36813 , \35819 );
or \U$31179 ( \36814 , \36783 , \36784 , \36785 , \36786 , \36787 , \36788 , \36789 , \36790 , \36791 , \36792 , \36793 , \36794 , \36795 , \36796 , \36797 , \36798 , \36799 , \36800 , \36801 , \36802 , \36803 , \36804 , \36805 , \36806 , \36807 , \36808 , \36809 , \36810 , \36811 , \36812 , \36813 );
nand \U$31180 ( \36815 , \36782 , \36814 );
buf \U$31181 ( \36816 , \36815 );
buf \U$31182 ( \36817 , \35832 );
not \U$31183 ( \36818 , \36817 );
buf \U$31184 ( \36819 , \35829 );
buf \U$31185 ( \36820 , \35832 );
buf \U$31186 ( \36821 , \35832 );
buf \U$31187 ( \36822 , \35832 );
buf \U$31188 ( \36823 , \35832 );
buf \U$31189 ( \36824 , \35832 );
buf \U$31190 ( \36825 , \35832 );
buf \U$31191 ( \36826 , \35832 );
buf \U$31192 ( \36827 , \35832 );
buf \U$31193 ( \36828 , \35832 );
buf \U$31194 ( \36829 , \35832 );
buf \U$31195 ( \36830 , \35832 );
buf \U$31196 ( \36831 , \35832 );
buf \U$31197 ( \36832 , \35832 );
buf \U$31198 ( \36833 , \35832 );
buf \U$31199 ( \36834 , \35832 );
buf \U$31200 ( \36835 , \35832 );
buf \U$31201 ( \36836 , \35832 );
buf \U$31202 ( \36837 , \35832 );
buf \U$31203 ( \36838 , \35832 );
buf \U$31204 ( \36839 , \35832 );
buf \U$31205 ( \36840 , \35832 );
buf \U$31206 ( \36841 , \35832 );
buf \U$31207 ( \36842 , \35832 );
buf \U$31208 ( \36843 , \35832 );
buf \U$31209 ( \36844 , \35832 );
buf \U$31210 ( \36845 , \35825 );
buf \U$31211 ( \36846 , \35819 );
buf \U$31212 ( \36847 , \35820 );
buf \U$31213 ( \36848 , \35821 );
buf \U$31214 ( \36849 , \35822 );
or \U$31215 ( \36850 , \36846 , \36847 , \36848 , \36849 );
and \U$31216 ( \36851 , \36845 , \36850 );
or \U$31217 ( \36852 , \36819 , \36820 , \36821 , \36822 , \36823 , \36824 , \36825 , \36826 , \36827 , \36828 , \36829 , \36830 , \36831 , \36832 , \36833 , \36834 , \36835 , \36836 , \36837 , \36838 , \36839 , \36840 , \36841 , \36842 , \36843 , \36844 , \36851 );
and \U$31218 ( \36853 , \36818 , \36852 );
buf \U$31219 ( \36854 , \36853 );
or \U$31220 ( \36855 , \36816 , \36854 );
_DC ga71c ( \36856_nGa71c , \36780 , \36855 );
buf \U$31221 ( \36857 , \36856_nGa71c );
xor \U$31222 ( \36858 , \36347 , \36857 );
buf \U$31223 ( \36859 , RIb7b9590_247);
and \U$31224 ( \36860 , \7126 , \36373 );
and \U$31225 ( \36861 , \7128 , \36400 );
and \U$31226 ( \36862 , \8338 , \36427 );
and \U$31227 ( \36863 , \8340 , \36454 );
and \U$31228 ( \36864 , \8342 , \36481 );
and \U$31229 ( \36865 , \8344 , \36508 );
and \U$31230 ( \36866 , \8346 , \36535 );
and \U$31231 ( \36867 , \8348 , \36562 );
and \U$31232 ( \36868 , \8350 , \36589 );
and \U$31233 ( \36869 , \8352 , \36616 );
and \U$31234 ( \36870 , \8354 , \36643 );
and \U$31235 ( \36871 , \8356 , \36670 );
and \U$31236 ( \36872 , \8358 , \36697 );
and \U$31237 ( \36873 , \8360 , \36724 );
and \U$31238 ( \36874 , \8362 , \36751 );
and \U$31239 ( \36875 , \8364 , \36778 );
or \U$31240 ( \36876 , \36860 , \36861 , \36862 , \36863 , \36864 , \36865 , \36866 , \36867 , \36868 , \36869 , \36870 , \36871 , \36872 , \36873 , \36874 , \36875 );
_DC ga731 ( \36877_nGa731 , \36876 , \36855 );
buf \U$31241 ( \36878 , \36877_nGa731 );
xor \U$31242 ( \36879 , \36859 , \36878 );
or \U$31243 ( \36880 , \36858 , \36879 );
buf \U$31244 ( \36881 , RIb7b9518_248);
and \U$31245 ( \36882 , \7136 , \36373 );
and \U$31246 ( \36883 , \7138 , \36400 );
and \U$31247 ( \36884 , \8374 , \36427 );
and \U$31248 ( \36885 , \8376 , \36454 );
and \U$31249 ( \36886 , \8378 , \36481 );
and \U$31250 ( \36887 , \8380 , \36508 );
and \U$31251 ( \36888 , \8382 , \36535 );
and \U$31252 ( \36889 , \8384 , \36562 );
and \U$31253 ( \36890 , \8386 , \36589 );
and \U$31254 ( \36891 , \8388 , \36616 );
and \U$31255 ( \36892 , \8390 , \36643 );
and \U$31256 ( \36893 , \8392 , \36670 );
and \U$31257 ( \36894 , \8394 , \36697 );
and \U$31258 ( \36895 , \8396 , \36724 );
and \U$31259 ( \36896 , \8398 , \36751 );
and \U$31260 ( \36897 , \8400 , \36778 );
or \U$31261 ( \36898 , \36882 , \36883 , \36884 , \36885 , \36886 , \36887 , \36888 , \36889 , \36890 , \36891 , \36892 , \36893 , \36894 , \36895 , \36896 , \36897 );
_DC ga747 ( \36899_nGa747 , \36898 , \36855 );
buf \U$31262 ( \36900 , \36899_nGa747 );
xor \U$31263 ( \36901 , \36881 , \36900 );
or \U$31264 ( \36902 , \36880 , \36901 );
buf \U$31265 ( \36903 , RIb7b94a0_249);
and \U$31266 ( \36904 , \7146 , \36373 );
and \U$31267 ( \36905 , \7148 , \36400 );
and \U$31268 ( \36906 , \8410 , \36427 );
and \U$31269 ( \36907 , \8412 , \36454 );
and \U$31270 ( \36908 , \8414 , \36481 );
and \U$31271 ( \36909 , \8416 , \36508 );
and \U$31272 ( \36910 , \8418 , \36535 );
and \U$31273 ( \36911 , \8420 , \36562 );
and \U$31274 ( \36912 , \8422 , \36589 );
and \U$31275 ( \36913 , \8424 , \36616 );
and \U$31276 ( \36914 , \8426 , \36643 );
and \U$31277 ( \36915 , \8428 , \36670 );
and \U$31278 ( \36916 , \8430 , \36697 );
and \U$31279 ( \36917 , \8432 , \36724 );
and \U$31280 ( \36918 , \8434 , \36751 );
and \U$31281 ( \36919 , \8436 , \36778 );
or \U$31282 ( \36920 , \36904 , \36905 , \36906 , \36907 , \36908 , \36909 , \36910 , \36911 , \36912 , \36913 , \36914 , \36915 , \36916 , \36917 , \36918 , \36919 );
_DC ga75d ( \36921_nGa75d , \36920 , \36855 );
buf \U$31283 ( \36922 , \36921_nGa75d );
xor \U$31284 ( \36923 , \36903 , \36922 );
or \U$31285 ( \36924 , \36902 , \36923 );
buf \U$31286 ( \36925 , RIb7b9428_250);
and \U$31287 ( \36926 , \7156 , \36373 );
and \U$31288 ( \36927 , \7158 , \36400 );
and \U$31289 ( \36928 , \8446 , \36427 );
and \U$31290 ( \36929 , \8448 , \36454 );
and \U$31291 ( \36930 , \8450 , \36481 );
and \U$31292 ( \36931 , \8452 , \36508 );
and \U$31293 ( \36932 , \8454 , \36535 );
and \U$31294 ( \36933 , \8456 , \36562 );
and \U$31295 ( \36934 , \8458 , \36589 );
and \U$31296 ( \36935 , \8460 , \36616 );
and \U$31297 ( \36936 , \8462 , \36643 );
and \U$31298 ( \36937 , \8464 , \36670 );
and \U$31299 ( \36938 , \8466 , \36697 );
and \U$31300 ( \36939 , \8468 , \36724 );
and \U$31301 ( \36940 , \8470 , \36751 );
and \U$31302 ( \36941 , \8472 , \36778 );
or \U$31303 ( \36942 , \36926 , \36927 , \36928 , \36929 , \36930 , \36931 , \36932 , \36933 , \36934 , \36935 , \36936 , \36937 , \36938 , \36939 , \36940 , \36941 );
_DC ga773 ( \36943_nGa773 , \36942 , \36855 );
buf \U$31304 ( \36944 , \36943_nGa773 );
xor \U$31305 ( \36945 , \36925 , \36944 );
or \U$31306 ( \36946 , \36924 , \36945 );
buf \U$31307 ( \36947 , RIb7b93b0_251);
and \U$31308 ( \36948 , \7166 , \36373 );
and \U$31309 ( \36949 , \7168 , \36400 );
and \U$31310 ( \36950 , \8482 , \36427 );
and \U$31311 ( \36951 , \8484 , \36454 );
and \U$31312 ( \36952 , \8486 , \36481 );
and \U$31313 ( \36953 , \8488 , \36508 );
and \U$31314 ( \36954 , \8490 , \36535 );
and \U$31315 ( \36955 , \8492 , \36562 );
and \U$31316 ( \36956 , \8494 , \36589 );
and \U$31317 ( \36957 , \8496 , \36616 );
and \U$31318 ( \36958 , \8498 , \36643 );
and \U$31319 ( \36959 , \8500 , \36670 );
and \U$31320 ( \36960 , \8502 , \36697 );
and \U$31321 ( \36961 , \8504 , \36724 );
and \U$31322 ( \36962 , \8506 , \36751 );
and \U$31323 ( \36963 , \8508 , \36778 );
or \U$31324 ( \36964 , \36948 , \36949 , \36950 , \36951 , \36952 , \36953 , \36954 , \36955 , \36956 , \36957 , \36958 , \36959 , \36960 , \36961 , \36962 , \36963 );
_DC ga789 ( \36965_nGa789 , \36964 , \36855 );
buf \U$31325 ( \36966 , \36965_nGa789 );
xor \U$31326 ( \36967 , \36947 , \36966 );
or \U$31327 ( \36968 , \36946 , \36967 );
buf \U$31328 ( \36969 , RIb7af720_252);
and \U$31329 ( \36970 , \7176 , \36373 );
and \U$31330 ( \36971 , \7178 , \36400 );
and \U$31331 ( \36972 , \8518 , \36427 );
and \U$31332 ( \36973 , \8520 , \36454 );
and \U$31333 ( \36974 , \8522 , \36481 );
and \U$31334 ( \36975 , \8524 , \36508 );
and \U$31335 ( \36976 , \8526 , \36535 );
and \U$31336 ( \36977 , \8528 , \36562 );
and \U$31337 ( \36978 , \8530 , \36589 );
and \U$31338 ( \36979 , \8532 , \36616 );
and \U$31339 ( \36980 , \8534 , \36643 );
and \U$31340 ( \36981 , \8536 , \36670 );
and \U$31341 ( \36982 , \8538 , \36697 );
and \U$31342 ( \36983 , \8540 , \36724 );
and \U$31343 ( \36984 , \8542 , \36751 );
and \U$31344 ( \36985 , \8544 , \36778 );
or \U$31345 ( \36986 , \36970 , \36971 , \36972 , \36973 , \36974 , \36975 , \36976 , \36977 , \36978 , \36979 , \36980 , \36981 , \36982 , \36983 , \36984 , \36985 );
_DC ga79f ( \36987_nGa79f , \36986 , \36855 );
buf \U$31346 ( \36988 , \36987_nGa79f );
xor \U$31347 ( \36989 , \36969 , \36988 );
or \U$31348 ( \36990 , \36968 , \36989 );
buf \U$31349 ( \36991 , RIb7af6a8_253);
and \U$31350 ( \36992 , \7186 , \36373 );
and \U$31351 ( \36993 , \7188 , \36400 );
and \U$31352 ( \36994 , \8554 , \36427 );
and \U$31353 ( \36995 , \8556 , \36454 );
and \U$31354 ( \36996 , \8558 , \36481 );
and \U$31355 ( \36997 , \8560 , \36508 );
and \U$31356 ( \36998 , \8562 , \36535 );
and \U$31357 ( \36999 , \8564 , \36562 );
and \U$31358 ( \37000 , \8566 , \36589 );
and \U$31359 ( \37001 , \8568 , \36616 );
and \U$31360 ( \37002 , \8570 , \36643 );
and \U$31361 ( \37003 , \8572 , \36670 );
and \U$31362 ( \37004 , \8574 , \36697 );
and \U$31363 ( \37005 , \8576 , \36724 );
and \U$31364 ( \37006 , \8578 , \36751 );
and \U$31365 ( \37007 , \8580 , \36778 );
or \U$31366 ( \37008 , \36992 , \36993 , \36994 , \36995 , \36996 , \36997 , \36998 , \36999 , \37000 , \37001 , \37002 , \37003 , \37004 , \37005 , \37006 , \37007 );
_DC ga7b5 ( \37009_nGa7b5 , \37008 , \36855 );
buf \U$31367 ( \37010 , \37009_nGa7b5 );
xor \U$31368 ( \37011 , \36991 , \37010 );
or \U$31369 ( \37012 , \36990 , \37011 );
not \U$31370 ( \37013 , \37012 );
buf \U$31371 ( \37014 , \37013 );
and \U$31372 ( \37015 , \36346 , \37014 );
buf \U$31373 ( \37016 , RIb7af630_254);
buf \U$31374 ( \37017 , \35832 );
buf \U$31375 ( \37018 , \35832 );
buf \U$31376 ( \37019 , \35832 );
buf \U$31377 ( \37020 , \35832 );
buf \U$31378 ( \37021 , \35832 );
buf \U$31379 ( \37022 , \35832 );
buf \U$31380 ( \37023 , \35832 );
buf \U$31381 ( \37024 , \35832 );
buf \U$31382 ( \37025 , \35832 );
buf \U$31383 ( \37026 , \35832 );
buf \U$31384 ( \37027 , \35832 );
buf \U$31385 ( \37028 , \35832 );
buf \U$31386 ( \37029 , \35832 );
buf \U$31387 ( \37030 , \35832 );
buf \U$31388 ( \37031 , \35832 );
buf \U$31389 ( \37032 , \35832 );
buf \U$31390 ( \37033 , \35832 );
buf \U$31391 ( \37034 , \35832 );
buf \U$31392 ( \37035 , \35832 );
buf \U$31393 ( \37036 , \35832 );
buf \U$31394 ( \37037 , \35832 );
buf \U$31395 ( \37038 , \35832 );
buf \U$31396 ( \37039 , \35832 );
buf \U$31397 ( \37040 , \35832 );
buf \U$31398 ( \37041 , \35832 );
nor \U$31399 ( \37042 , \35819 , \35820 , \35821 , \35822 , \35826 , \35829 , \35832 , \37017 , \37018 , \37019 , \37020 , \37021 , \37022 , \37023 , \37024 , \37025 , \37026 , \37027 , \37028 , \37029 , \37030 , \37031 , \37032 , \37033 , \37034 , \37035 , \37036 , \37037 , \37038 , \37039 , \37040 , \37041 );
and \U$31400 ( \37043 , \7198 , \37042 );
buf \U$31401 ( \37044 , \35832 );
buf \U$31402 ( \37045 , \35832 );
buf \U$31403 ( \37046 , \35832 );
buf \U$31404 ( \37047 , \35832 );
buf \U$31405 ( \37048 , \35832 );
buf \U$31406 ( \37049 , \35832 );
buf \U$31407 ( \37050 , \35832 );
buf \U$31408 ( \37051 , \35832 );
buf \U$31409 ( \37052 , \35832 );
buf \U$31410 ( \37053 , \35832 );
buf \U$31411 ( \37054 , \35832 );
buf \U$31412 ( \37055 , \35832 );
buf \U$31413 ( \37056 , \35832 );
buf \U$31414 ( \37057 , \35832 );
buf \U$31415 ( \37058 , \35832 );
buf \U$31416 ( \37059 , \35832 );
buf \U$31417 ( \37060 , \35832 );
buf \U$31418 ( \37061 , \35832 );
buf \U$31419 ( \37062 , \35832 );
buf \U$31420 ( \37063 , \35832 );
buf \U$31421 ( \37064 , \35832 );
buf \U$31422 ( \37065 , \35832 );
buf \U$31423 ( \37066 , \35832 );
buf \U$31424 ( \37067 , \35832 );
buf \U$31425 ( \37068 , \35832 );
nor \U$31426 ( \37069 , \35860 , \35861 , \35862 , \35863 , \35825 , \35829 , \35832 , \37044 , \37045 , \37046 , \37047 , \37048 , \37049 , \37050 , \37051 , \37052 , \37053 , \37054 , \37055 , \37056 , \37057 , \37058 , \37059 , \37060 , \37061 , \37062 , \37063 , \37064 , \37065 , \37066 , \37067 , \37068 );
and \U$31427 ( \37070 , \7200 , \37069 );
buf \U$31428 ( \37071 , \35832 );
buf \U$31429 ( \37072 , \35832 );
buf \U$31430 ( \37073 , \35832 );
buf \U$31431 ( \37074 , \35832 );
buf \U$31432 ( \37075 , \35832 );
buf \U$31433 ( \37076 , \35832 );
buf \U$31434 ( \37077 , \35832 );
buf \U$31435 ( \37078 , \35832 );
buf \U$31436 ( \37079 , \35832 );
buf \U$31437 ( \37080 , \35832 );
buf \U$31438 ( \37081 , \35832 );
buf \U$31439 ( \37082 , \35832 );
buf \U$31440 ( \37083 , \35832 );
buf \U$31441 ( \37084 , \35832 );
buf \U$31442 ( \37085 , \35832 );
buf \U$31443 ( \37086 , \35832 );
buf \U$31444 ( \37087 , \35832 );
buf \U$31445 ( \37088 , \35832 );
buf \U$31446 ( \37089 , \35832 );
buf \U$31447 ( \37090 , \35832 );
buf \U$31448 ( \37091 , \35832 );
buf \U$31449 ( \37092 , \35832 );
buf \U$31450 ( \37093 , \35832 );
buf \U$31451 ( \37094 , \35832 );
buf \U$31452 ( \37095 , \35832 );
nor \U$31453 ( \37096 , \35819 , \35861 , \35862 , \35863 , \35825 , \35829 , \35832 , \37071 , \37072 , \37073 , \37074 , \37075 , \37076 , \37077 , \37078 , \37079 , \37080 , \37081 , \37082 , \37083 , \37084 , \37085 , \37086 , \37087 , \37088 , \37089 , \37090 , \37091 , \37092 , \37093 , \37094 , \37095 );
and \U$31454 ( \37097 , \8645 , \37096 );
buf \U$31455 ( \37098 , \35832 );
buf \U$31456 ( \37099 , \35832 );
buf \U$31457 ( \37100 , \35832 );
buf \U$31458 ( \37101 , \35832 );
buf \U$31459 ( \37102 , \35832 );
buf \U$31460 ( \37103 , \35832 );
buf \U$31461 ( \37104 , \35832 );
buf \U$31462 ( \37105 , \35832 );
buf \U$31463 ( \37106 , \35832 );
buf \U$31464 ( \37107 , \35832 );
buf \U$31465 ( \37108 , \35832 );
buf \U$31466 ( \37109 , \35832 );
buf \U$31467 ( \37110 , \35832 );
buf \U$31468 ( \37111 , \35832 );
buf \U$31469 ( \37112 , \35832 );
buf \U$31470 ( \37113 , \35832 );
buf \U$31471 ( \37114 , \35832 );
buf \U$31472 ( \37115 , \35832 );
buf \U$31473 ( \37116 , \35832 );
buf \U$31474 ( \37117 , \35832 );
buf \U$31475 ( \37118 , \35832 );
buf \U$31476 ( \37119 , \35832 );
buf \U$31477 ( \37120 , \35832 );
buf \U$31478 ( \37121 , \35832 );
buf \U$31479 ( \37122 , \35832 );
nor \U$31480 ( \37123 , \35860 , \35820 , \35862 , \35863 , \35825 , \35829 , \35832 , \37098 , \37099 , \37100 , \37101 , \37102 , \37103 , \37104 , \37105 , \37106 , \37107 , \37108 , \37109 , \37110 , \37111 , \37112 , \37113 , \37114 , \37115 , \37116 , \37117 , \37118 , \37119 , \37120 , \37121 , \37122 );
and \U$31481 ( \37124 , \8673 , \37123 );
buf \U$31482 ( \37125 , \35832 );
buf \U$31483 ( \37126 , \35832 );
buf \U$31484 ( \37127 , \35832 );
buf \U$31485 ( \37128 , \35832 );
buf \U$31486 ( \37129 , \35832 );
buf \U$31487 ( \37130 , \35832 );
buf \U$31488 ( \37131 , \35832 );
buf \U$31489 ( \37132 , \35832 );
buf \U$31490 ( \37133 , \35832 );
buf \U$31491 ( \37134 , \35832 );
buf \U$31492 ( \37135 , \35832 );
buf \U$31493 ( \37136 , \35832 );
buf \U$31494 ( \37137 , \35832 );
buf \U$31495 ( \37138 , \35832 );
buf \U$31496 ( \37139 , \35832 );
buf \U$31497 ( \37140 , \35832 );
buf \U$31498 ( \37141 , \35832 );
buf \U$31499 ( \37142 , \35832 );
buf \U$31500 ( \37143 , \35832 );
buf \U$31501 ( \37144 , \35832 );
buf \U$31502 ( \37145 , \35832 );
buf \U$31503 ( \37146 , \35832 );
buf \U$31504 ( \37147 , \35832 );
buf \U$31505 ( \37148 , \35832 );
buf \U$31506 ( \37149 , \35832 );
nor \U$31507 ( \37150 , \35819 , \35820 , \35862 , \35863 , \35825 , \35829 , \35832 , \37125 , \37126 , \37127 , \37128 , \37129 , \37130 , \37131 , \37132 , \37133 , \37134 , \37135 , \37136 , \37137 , \37138 , \37139 , \37140 , \37141 , \37142 , \37143 , \37144 , \37145 , \37146 , \37147 , \37148 , \37149 );
and \U$31508 ( \37151 , \8701 , \37150 );
buf \U$31509 ( \37152 , \35832 );
buf \U$31510 ( \37153 , \35832 );
buf \U$31511 ( \37154 , \35832 );
buf \U$31512 ( \37155 , \35832 );
buf \U$31513 ( \37156 , \35832 );
buf \U$31514 ( \37157 , \35832 );
buf \U$31515 ( \37158 , \35832 );
buf \U$31516 ( \37159 , \35832 );
buf \U$31517 ( \37160 , \35832 );
buf \U$31518 ( \37161 , \35832 );
buf \U$31519 ( \37162 , \35832 );
buf \U$31520 ( \37163 , \35832 );
buf \U$31521 ( \37164 , \35832 );
buf \U$31522 ( \37165 , \35832 );
buf \U$31523 ( \37166 , \35832 );
buf \U$31524 ( \37167 , \35832 );
buf \U$31525 ( \37168 , \35832 );
buf \U$31526 ( \37169 , \35832 );
buf \U$31527 ( \37170 , \35832 );
buf \U$31528 ( \37171 , \35832 );
buf \U$31529 ( \37172 , \35832 );
buf \U$31530 ( \37173 , \35832 );
buf \U$31531 ( \37174 , \35832 );
buf \U$31532 ( \37175 , \35832 );
buf \U$31533 ( \37176 , \35832 );
nor \U$31534 ( \37177 , \35860 , \35861 , \35821 , \35863 , \35825 , \35829 , \35832 , \37152 , \37153 , \37154 , \37155 , \37156 , \37157 , \37158 , \37159 , \37160 , \37161 , \37162 , \37163 , \37164 , \37165 , \37166 , \37167 , \37168 , \37169 , \37170 , \37171 , \37172 , \37173 , \37174 , \37175 , \37176 );
and \U$31535 ( \37178 , \8729 , \37177 );
buf \U$31536 ( \37179 , \35832 );
buf \U$31537 ( \37180 , \35832 );
buf \U$31538 ( \37181 , \35832 );
buf \U$31539 ( \37182 , \35832 );
buf \U$31540 ( \37183 , \35832 );
buf \U$31541 ( \37184 , \35832 );
buf \U$31542 ( \37185 , \35832 );
buf \U$31543 ( \37186 , \35832 );
buf \U$31544 ( \37187 , \35832 );
buf \U$31545 ( \37188 , \35832 );
buf \U$31546 ( \37189 , \35832 );
buf \U$31547 ( \37190 , \35832 );
buf \U$31548 ( \37191 , \35832 );
buf \U$31549 ( \37192 , \35832 );
buf \U$31550 ( \37193 , \35832 );
buf \U$31551 ( \37194 , \35832 );
buf \U$31552 ( \37195 , \35832 );
buf \U$31553 ( \37196 , \35832 );
buf \U$31554 ( \37197 , \35832 );
buf \U$31555 ( \37198 , \35832 );
buf \U$31556 ( \37199 , \35832 );
buf \U$31557 ( \37200 , \35832 );
buf \U$31558 ( \37201 , \35832 );
buf \U$31559 ( \37202 , \35832 );
buf \U$31560 ( \37203 , \35832 );
nor \U$31561 ( \37204 , \35819 , \35861 , \35821 , \35863 , \35825 , \35829 , \35832 , \37179 , \37180 , \37181 , \37182 , \37183 , \37184 , \37185 , \37186 , \37187 , \37188 , \37189 , \37190 , \37191 , \37192 , \37193 , \37194 , \37195 , \37196 , \37197 , \37198 , \37199 , \37200 , \37201 , \37202 , \37203 );
and \U$31562 ( \37205 , \8757 , \37204 );
buf \U$31563 ( \37206 , \35832 );
buf \U$31564 ( \37207 , \35832 );
buf \U$31565 ( \37208 , \35832 );
buf \U$31566 ( \37209 , \35832 );
buf \U$31567 ( \37210 , \35832 );
buf \U$31568 ( \37211 , \35832 );
buf \U$31569 ( \37212 , \35832 );
buf \U$31570 ( \37213 , \35832 );
buf \U$31571 ( \37214 , \35832 );
buf \U$31572 ( \37215 , \35832 );
buf \U$31573 ( \37216 , \35832 );
buf \U$31574 ( \37217 , \35832 );
buf \U$31575 ( \37218 , \35832 );
buf \U$31576 ( \37219 , \35832 );
buf \U$31577 ( \37220 , \35832 );
buf \U$31578 ( \37221 , \35832 );
buf \U$31579 ( \37222 , \35832 );
buf \U$31580 ( \37223 , \35832 );
buf \U$31581 ( \37224 , \35832 );
buf \U$31582 ( \37225 , \35832 );
buf \U$31583 ( \37226 , \35832 );
buf \U$31584 ( \37227 , \35832 );
buf \U$31585 ( \37228 , \35832 );
buf \U$31586 ( \37229 , \35832 );
buf \U$31587 ( \37230 , \35832 );
nor \U$31588 ( \37231 , \35860 , \35820 , \35821 , \35863 , \35825 , \35829 , \35832 , \37206 , \37207 , \37208 , \37209 , \37210 , \37211 , \37212 , \37213 , \37214 , \37215 , \37216 , \37217 , \37218 , \37219 , \37220 , \37221 , \37222 , \37223 , \37224 , \37225 , \37226 , \37227 , \37228 , \37229 , \37230 );
and \U$31589 ( \37232 , \8785 , \37231 );
buf \U$31590 ( \37233 , \35832 );
buf \U$31591 ( \37234 , \35832 );
buf \U$31592 ( \37235 , \35832 );
buf \U$31593 ( \37236 , \35832 );
buf \U$31594 ( \37237 , \35832 );
buf \U$31595 ( \37238 , \35832 );
buf \U$31596 ( \37239 , \35832 );
buf \U$31597 ( \37240 , \35832 );
buf \U$31598 ( \37241 , \35832 );
buf \U$31599 ( \37242 , \35832 );
buf \U$31600 ( \37243 , \35832 );
buf \U$31601 ( \37244 , \35832 );
buf \U$31602 ( \37245 , \35832 );
buf \U$31603 ( \37246 , \35832 );
buf \U$31604 ( \37247 , \35832 );
buf \U$31605 ( \37248 , \35832 );
buf \U$31606 ( \37249 , \35832 );
buf \U$31607 ( \37250 , \35832 );
buf \U$31608 ( \37251 , \35832 );
buf \U$31609 ( \37252 , \35832 );
buf \U$31610 ( \37253 , \35832 );
buf \U$31611 ( \37254 , \35832 );
buf \U$31612 ( \37255 , \35832 );
buf \U$31613 ( \37256 , \35832 );
buf \U$31614 ( \37257 , \35832 );
nor \U$31615 ( \37258 , \35819 , \35820 , \35821 , \35863 , \35825 , \35829 , \35832 , \37233 , \37234 , \37235 , \37236 , \37237 , \37238 , \37239 , \37240 , \37241 , \37242 , \37243 , \37244 , \37245 , \37246 , \37247 , \37248 , \37249 , \37250 , \37251 , \37252 , \37253 , \37254 , \37255 , \37256 , \37257 );
and \U$31616 ( \37259 , \8813 , \37258 );
buf \U$31617 ( \37260 , \35832 );
buf \U$31618 ( \37261 , \35832 );
buf \U$31619 ( \37262 , \35832 );
buf \U$31620 ( \37263 , \35832 );
buf \U$31621 ( \37264 , \35832 );
buf \U$31622 ( \37265 , \35832 );
buf \U$31623 ( \37266 , \35832 );
buf \U$31624 ( \37267 , \35832 );
buf \U$31625 ( \37268 , \35832 );
buf \U$31626 ( \37269 , \35832 );
buf \U$31627 ( \37270 , \35832 );
buf \U$31628 ( \37271 , \35832 );
buf \U$31629 ( \37272 , \35832 );
buf \U$31630 ( \37273 , \35832 );
buf \U$31631 ( \37274 , \35832 );
buf \U$31632 ( \37275 , \35832 );
buf \U$31633 ( \37276 , \35832 );
buf \U$31634 ( \37277 , \35832 );
buf \U$31635 ( \37278 , \35832 );
buf \U$31636 ( \37279 , \35832 );
buf \U$31637 ( \37280 , \35832 );
buf \U$31638 ( \37281 , \35832 );
buf \U$31639 ( \37282 , \35832 );
buf \U$31640 ( \37283 , \35832 );
buf \U$31641 ( \37284 , \35832 );
nor \U$31642 ( \37285 , \35860 , \35861 , \35862 , \35822 , \35825 , \35829 , \35832 , \37260 , \37261 , \37262 , \37263 , \37264 , \37265 , \37266 , \37267 , \37268 , \37269 , \37270 , \37271 , \37272 , \37273 , \37274 , \37275 , \37276 , \37277 , \37278 , \37279 , \37280 , \37281 , \37282 , \37283 , \37284 );
and \U$31643 ( \37286 , \8841 , \37285 );
buf \U$31644 ( \37287 , \35832 );
buf \U$31645 ( \37288 , \35832 );
buf \U$31646 ( \37289 , \35832 );
buf \U$31647 ( \37290 , \35832 );
buf \U$31648 ( \37291 , \35832 );
buf \U$31649 ( \37292 , \35832 );
buf \U$31650 ( \37293 , \35832 );
buf \U$31651 ( \37294 , \35832 );
buf \U$31652 ( \37295 , \35832 );
buf \U$31653 ( \37296 , \35832 );
buf \U$31654 ( \37297 , \35832 );
buf \U$31655 ( \37298 , \35832 );
buf \U$31656 ( \37299 , \35832 );
buf \U$31657 ( \37300 , \35832 );
buf \U$31658 ( \37301 , \35832 );
buf \U$31659 ( \37302 , \35832 );
buf \U$31660 ( \37303 , \35832 );
buf \U$31661 ( \37304 , \35832 );
buf \U$31662 ( \37305 , \35832 );
buf \U$31663 ( \37306 , \35832 );
buf \U$31664 ( \37307 , \35832 );
buf \U$31665 ( \37308 , \35832 );
buf \U$31666 ( \37309 , \35832 );
buf \U$31667 ( \37310 , \35832 );
buf \U$31668 ( \37311 , \35832 );
nor \U$31669 ( \37312 , \35819 , \35861 , \35862 , \35822 , \35825 , \35829 , \35832 , \37287 , \37288 , \37289 , \37290 , \37291 , \37292 , \37293 , \37294 , \37295 , \37296 , \37297 , \37298 , \37299 , \37300 , \37301 , \37302 , \37303 , \37304 , \37305 , \37306 , \37307 , \37308 , \37309 , \37310 , \37311 );
and \U$31670 ( \37313 , \8869 , \37312 );
buf \U$31671 ( \37314 , \35832 );
buf \U$31672 ( \37315 , \35832 );
buf \U$31673 ( \37316 , \35832 );
buf \U$31674 ( \37317 , \35832 );
buf \U$31675 ( \37318 , \35832 );
buf \U$31676 ( \37319 , \35832 );
buf \U$31677 ( \37320 , \35832 );
buf \U$31678 ( \37321 , \35832 );
buf \U$31679 ( \37322 , \35832 );
buf \U$31680 ( \37323 , \35832 );
buf \U$31681 ( \37324 , \35832 );
buf \U$31682 ( \37325 , \35832 );
buf \U$31683 ( \37326 , \35832 );
buf \U$31684 ( \37327 , \35832 );
buf \U$31685 ( \37328 , \35832 );
buf \U$31686 ( \37329 , \35832 );
buf \U$31687 ( \37330 , \35832 );
buf \U$31688 ( \37331 , \35832 );
buf \U$31689 ( \37332 , \35832 );
buf \U$31690 ( \37333 , \35832 );
buf \U$31691 ( \37334 , \35832 );
buf \U$31692 ( \37335 , \35832 );
buf \U$31693 ( \37336 , \35832 );
buf \U$31694 ( \37337 , \35832 );
buf \U$31695 ( \37338 , \35832 );
nor \U$31696 ( \37339 , \35860 , \35820 , \35862 , \35822 , \35825 , \35829 , \35832 , \37314 , \37315 , \37316 , \37317 , \37318 , \37319 , \37320 , \37321 , \37322 , \37323 , \37324 , \37325 , \37326 , \37327 , \37328 , \37329 , \37330 , \37331 , \37332 , \37333 , \37334 , \37335 , \37336 , \37337 , \37338 );
and \U$31697 ( \37340 , \8897 , \37339 );
buf \U$31698 ( \37341 , \35832 );
buf \U$31699 ( \37342 , \35832 );
buf \U$31700 ( \37343 , \35832 );
buf \U$31701 ( \37344 , \35832 );
buf \U$31702 ( \37345 , \35832 );
buf \U$31703 ( \37346 , \35832 );
buf \U$31704 ( \37347 , \35832 );
buf \U$31705 ( \37348 , \35832 );
buf \U$31706 ( \37349 , \35832 );
buf \U$31707 ( \37350 , \35832 );
buf \U$31708 ( \37351 , \35832 );
buf \U$31709 ( \37352 , \35832 );
buf \U$31710 ( \37353 , \35832 );
buf \U$31711 ( \37354 , \35832 );
buf \U$31712 ( \37355 , \35832 );
buf \U$31713 ( \37356 , \35832 );
buf \U$31714 ( \37357 , \35832 );
buf \U$31715 ( \37358 , \35832 );
buf \U$31716 ( \37359 , \35832 );
buf \U$31717 ( \37360 , \35832 );
buf \U$31718 ( \37361 , \35832 );
buf \U$31719 ( \37362 , \35832 );
buf \U$31720 ( \37363 , \35832 );
buf \U$31721 ( \37364 , \35832 );
buf \U$31722 ( \37365 , \35832 );
nor \U$31723 ( \37366 , \35819 , \35820 , \35862 , \35822 , \35825 , \35829 , \35832 , \37341 , \37342 , \37343 , \37344 , \37345 , \37346 , \37347 , \37348 , \37349 , \37350 , \37351 , \37352 , \37353 , \37354 , \37355 , \37356 , \37357 , \37358 , \37359 , \37360 , \37361 , \37362 , \37363 , \37364 , \37365 );
and \U$31724 ( \37367 , \8925 , \37366 );
buf \U$31725 ( \37368 , \35832 );
buf \U$31726 ( \37369 , \35832 );
buf \U$31727 ( \37370 , \35832 );
buf \U$31728 ( \37371 , \35832 );
buf \U$31729 ( \37372 , \35832 );
buf \U$31730 ( \37373 , \35832 );
buf \U$31731 ( \37374 , \35832 );
buf \U$31732 ( \37375 , \35832 );
buf \U$31733 ( \37376 , \35832 );
buf \U$31734 ( \37377 , \35832 );
buf \U$31735 ( \37378 , \35832 );
buf \U$31736 ( \37379 , \35832 );
buf \U$31737 ( \37380 , \35832 );
buf \U$31738 ( \37381 , \35832 );
buf \U$31739 ( \37382 , \35832 );
buf \U$31740 ( \37383 , \35832 );
buf \U$31741 ( \37384 , \35832 );
buf \U$31742 ( \37385 , \35832 );
buf \U$31743 ( \37386 , \35832 );
buf \U$31744 ( \37387 , \35832 );
buf \U$31745 ( \37388 , \35832 );
buf \U$31746 ( \37389 , \35832 );
buf \U$31747 ( \37390 , \35832 );
buf \U$31748 ( \37391 , \35832 );
buf \U$31749 ( \37392 , \35832 );
nor \U$31750 ( \37393 , \35860 , \35861 , \35821 , \35822 , \35825 , \35829 , \35832 , \37368 , \37369 , \37370 , \37371 , \37372 , \37373 , \37374 , \37375 , \37376 , \37377 , \37378 , \37379 , \37380 , \37381 , \37382 , \37383 , \37384 , \37385 , \37386 , \37387 , \37388 , \37389 , \37390 , \37391 , \37392 );
and \U$31751 ( \37394 , \8953 , \37393 );
buf \U$31752 ( \37395 , \35832 );
buf \U$31753 ( \37396 , \35832 );
buf \U$31754 ( \37397 , \35832 );
buf \U$31755 ( \37398 , \35832 );
buf \U$31756 ( \37399 , \35832 );
buf \U$31757 ( \37400 , \35832 );
buf \U$31758 ( \37401 , \35832 );
buf \U$31759 ( \37402 , \35832 );
buf \U$31760 ( \37403 , \35832 );
buf \U$31761 ( \37404 , \35832 );
buf \U$31762 ( \37405 , \35832 );
buf \U$31763 ( \37406 , \35832 );
buf \U$31764 ( \37407 , \35832 );
buf \U$31765 ( \37408 , \35832 );
buf \U$31766 ( \37409 , \35832 );
buf \U$31767 ( \37410 , \35832 );
buf \U$31768 ( \37411 , \35832 );
buf \U$31769 ( \37412 , \35832 );
buf \U$31770 ( \37413 , \35832 );
buf \U$31771 ( \37414 , \35832 );
buf \U$31772 ( \37415 , \35832 );
buf \U$31773 ( \37416 , \35832 );
buf \U$31774 ( \37417 , \35832 );
buf \U$31775 ( \37418 , \35832 );
buf \U$31776 ( \37419 , \35832 );
nor \U$31777 ( \37420 , \35819 , \35861 , \35821 , \35822 , \35825 , \35829 , \35832 , \37395 , \37396 , \37397 , \37398 , \37399 , \37400 , \37401 , \37402 , \37403 , \37404 , \37405 , \37406 , \37407 , \37408 , \37409 , \37410 , \37411 , \37412 , \37413 , \37414 , \37415 , \37416 , \37417 , \37418 , \37419 );
and \U$31778 ( \37421 , \8981 , \37420 );
buf \U$31779 ( \37422 , \35832 );
buf \U$31780 ( \37423 , \35832 );
buf \U$31781 ( \37424 , \35832 );
buf \U$31782 ( \37425 , \35832 );
buf \U$31783 ( \37426 , \35832 );
buf \U$31784 ( \37427 , \35832 );
buf \U$31785 ( \37428 , \35832 );
buf \U$31786 ( \37429 , \35832 );
buf \U$31787 ( \37430 , \35832 );
buf \U$31788 ( \37431 , \35832 );
buf \U$31789 ( \37432 , \35832 );
buf \U$31790 ( \37433 , \35832 );
buf \U$31791 ( \37434 , \35832 );
buf \U$31792 ( \37435 , \35832 );
buf \U$31793 ( \37436 , \35832 );
buf \U$31794 ( \37437 , \35832 );
buf \U$31795 ( \37438 , \35832 );
buf \U$31796 ( \37439 , \35832 );
buf \U$31797 ( \37440 , \35832 );
buf \U$31798 ( \37441 , \35832 );
buf \U$31799 ( \37442 , \35832 );
buf \U$31800 ( \37443 , \35832 );
buf \U$31801 ( \37444 , \35832 );
buf \U$31802 ( \37445 , \35832 );
buf \U$31803 ( \37446 , \35832 );
nor \U$31804 ( \37447 , \35860 , \35820 , \35821 , \35822 , \35825 , \35829 , \35832 , \37422 , \37423 , \37424 , \37425 , \37426 , \37427 , \37428 , \37429 , \37430 , \37431 , \37432 , \37433 , \37434 , \37435 , \37436 , \37437 , \37438 , \37439 , \37440 , \37441 , \37442 , \37443 , \37444 , \37445 , \37446 );
and \U$31805 ( \37448 , \9009 , \37447 );
or \U$31806 ( \37449 , \37043 , \37070 , \37097 , \37124 , \37151 , \37178 , \37205 , \37232 , \37259 , \37286 , \37313 , \37340 , \37367 , \37394 , \37421 , \37448 );
buf \U$31807 ( \37450 , \35832 );
not \U$31808 ( \37451 , \37450 );
buf \U$31809 ( \37452 , \35820 );
buf \U$31810 ( \37453 , \35821 );
buf \U$31811 ( \37454 , \35822 );
buf \U$31812 ( \37455 , \35825 );
buf \U$31813 ( \37456 , \35829 );
buf \U$31814 ( \37457 , \35832 );
buf \U$31815 ( \37458 , \35832 );
buf \U$31816 ( \37459 , \35832 );
buf \U$31817 ( \37460 , \35832 );
buf \U$31818 ( \37461 , \35832 );
buf \U$31819 ( \37462 , \35832 );
buf \U$31820 ( \37463 , \35832 );
buf \U$31821 ( \37464 , \35832 );
buf \U$31822 ( \37465 , \35832 );
buf \U$31823 ( \37466 , \35832 );
buf \U$31824 ( \37467 , \35832 );
buf \U$31825 ( \37468 , \35832 );
buf \U$31826 ( \37469 , \35832 );
buf \U$31827 ( \37470 , \35832 );
buf \U$31828 ( \37471 , \35832 );
buf \U$31829 ( \37472 , \35832 );
buf \U$31830 ( \37473 , \35832 );
buf \U$31831 ( \37474 , \35832 );
buf \U$31832 ( \37475 , \35832 );
buf \U$31833 ( \37476 , \35832 );
buf \U$31834 ( \37477 , \35832 );
buf \U$31835 ( \37478 , \35832 );
buf \U$31836 ( \37479 , \35832 );
buf \U$31837 ( \37480 , \35832 );
buf \U$31838 ( \37481 , \35832 );
buf \U$31839 ( \37482 , \35819 );
or \U$31840 ( \37483 , \37452 , \37453 , \37454 , \37455 , \37456 , \37457 , \37458 , \37459 , \37460 , \37461 , \37462 , \37463 , \37464 , \37465 , \37466 , \37467 , \37468 , \37469 , \37470 , \37471 , \37472 , \37473 , \37474 , \37475 , \37476 , \37477 , \37478 , \37479 , \37480 , \37481 , \37482 );
nand \U$31841 ( \37484 , \37451 , \37483 );
buf \U$31842 ( \37485 , \37484 );
buf \U$31843 ( \37486 , \35832 );
not \U$31844 ( \37487 , \37486 );
buf \U$31845 ( \37488 , \35829 );
buf \U$31846 ( \37489 , \35832 );
buf \U$31847 ( \37490 , \35832 );
buf \U$31848 ( \37491 , \35832 );
buf \U$31849 ( \37492 , \35832 );
buf \U$31850 ( \37493 , \35832 );
buf \U$31851 ( \37494 , \35832 );
buf \U$31852 ( \37495 , \35832 );
buf \U$31853 ( \37496 , \35832 );
buf \U$31854 ( \37497 , \35832 );
buf \U$31855 ( \37498 , \35832 );
buf \U$31856 ( \37499 , \35832 );
buf \U$31857 ( \37500 , \35832 );
buf \U$31858 ( \37501 , \35832 );
buf \U$31859 ( \37502 , \35832 );
buf \U$31860 ( \37503 , \35832 );
buf \U$31861 ( \37504 , \35832 );
buf \U$31862 ( \37505 , \35832 );
buf \U$31863 ( \37506 , \35832 );
buf \U$31864 ( \37507 , \35832 );
buf \U$31865 ( \37508 , \35832 );
buf \U$31866 ( \37509 , \35832 );
buf \U$31867 ( \37510 , \35832 );
buf \U$31868 ( \37511 , \35832 );
buf \U$31869 ( \37512 , \35832 );
buf \U$31870 ( \37513 , \35832 );
buf \U$31871 ( \37514 , \35825 );
buf \U$31872 ( \37515 , \35819 );
buf \U$31873 ( \37516 , \35820 );
buf \U$31874 ( \37517 , \35821 );
buf \U$31875 ( \37518 , \35822 );
or \U$31876 ( \37519 , \37515 , \37516 , \37517 , \37518 );
and \U$31877 ( \37520 , \37514 , \37519 );
or \U$31878 ( \37521 , \37488 , \37489 , \37490 , \37491 , \37492 , \37493 , \37494 , \37495 , \37496 , \37497 , \37498 , \37499 , \37500 , \37501 , \37502 , \37503 , \37504 , \37505 , \37506 , \37507 , \37508 , \37509 , \37510 , \37511 , \37512 , \37513 , \37520 );
and \U$31879 ( \37522 , \37487 , \37521 );
buf \U$31880 ( \37523 , \37522 );
or \U$31881 ( \37524 , \37485 , \37523 );
_DC ga9b9 ( \37525_nGa9b9 , \37449 , \37524 );
buf \U$31882 ( \37526 , \37525_nGa9b9 );
xor \U$31883 ( \37527 , \37016 , \37526 );
buf \U$31884 ( \37528 , RIb7af5b8_255);
and \U$31885 ( \37529 , \7207 , \37042 );
and \U$31886 ( \37530 , \7209 , \37069 );
and \U$31887 ( \37531 , \9119 , \37096 );
and \U$31888 ( \37532 , \9121 , \37123 );
and \U$31889 ( \37533 , \9123 , \37150 );
and \U$31890 ( \37534 , \9125 , \37177 );
and \U$31891 ( \37535 , \9127 , \37204 );
and \U$31892 ( \37536 , \9129 , \37231 );
and \U$31893 ( \37537 , \9131 , \37258 );
and \U$31894 ( \37538 , \9133 , \37285 );
and \U$31895 ( \37539 , \9135 , \37312 );
and \U$31896 ( \37540 , \9137 , \37339 );
and \U$31897 ( \37541 , \9139 , \37366 );
and \U$31898 ( \37542 , \9141 , \37393 );
and \U$31899 ( \37543 , \9143 , \37420 );
and \U$31900 ( \37544 , \9145 , \37447 );
or \U$31901 ( \37545 , \37529 , \37530 , \37531 , \37532 , \37533 , \37534 , \37535 , \37536 , \37537 , \37538 , \37539 , \37540 , \37541 , \37542 , \37543 , \37544 );
_DC ga9ce ( \37546_nGa9ce , \37545 , \37524 );
buf \U$31902 ( \37547 , \37546_nGa9ce );
xor \U$31903 ( \37548 , \37528 , \37547 );
or \U$31904 ( \37549 , \37527 , \37548 );
buf \U$31905 ( \37550 , RIb7af540_256);
and \U$31906 ( \37551 , \7217 , \37042 );
and \U$31907 ( \37552 , \7219 , \37069 );
and \U$31908 ( \37553 , \9155 , \37096 );
and \U$31909 ( \37554 , \9157 , \37123 );
and \U$31910 ( \37555 , \9159 , \37150 );
and \U$31911 ( \37556 , \9161 , \37177 );
and \U$31912 ( \37557 , \9163 , \37204 );
and \U$31913 ( \37558 , \9165 , \37231 );
and \U$31914 ( \37559 , \9167 , \37258 );
and \U$31915 ( \37560 , \9169 , \37285 );
and \U$31916 ( \37561 , \9171 , \37312 );
and \U$31917 ( \37562 , \9173 , \37339 );
and \U$31918 ( \37563 , \9175 , \37366 );
and \U$31919 ( \37564 , \9177 , \37393 );
and \U$31920 ( \37565 , \9179 , \37420 );
and \U$31921 ( \37566 , \9181 , \37447 );
or \U$31922 ( \37567 , \37551 , \37552 , \37553 , \37554 , \37555 , \37556 , \37557 , \37558 , \37559 , \37560 , \37561 , \37562 , \37563 , \37564 , \37565 , \37566 );
_DC ga9e4 ( \37568_nGa9e4 , \37567 , \37524 );
buf \U$31923 ( \37569 , \37568_nGa9e4 );
xor \U$31924 ( \37570 , \37550 , \37569 );
or \U$31925 ( \37571 , \37549 , \37570 );
buf \U$31926 ( \37572 , RIb7af4c8_257);
and \U$31927 ( \37573 , \7227 , \37042 );
and \U$31928 ( \37574 , \7229 , \37069 );
and \U$31929 ( \37575 , \9191 , \37096 );
and \U$31930 ( \37576 , \9193 , \37123 );
and \U$31931 ( \37577 , \9195 , \37150 );
and \U$31932 ( \37578 , \9197 , \37177 );
and \U$31933 ( \37579 , \9199 , \37204 );
and \U$31934 ( \37580 , \9201 , \37231 );
and \U$31935 ( \37581 , \9203 , \37258 );
and \U$31936 ( \37582 , \9205 , \37285 );
and \U$31937 ( \37583 , \9207 , \37312 );
and \U$31938 ( \37584 , \9209 , \37339 );
and \U$31939 ( \37585 , \9211 , \37366 );
and \U$31940 ( \37586 , \9213 , \37393 );
and \U$31941 ( \37587 , \9215 , \37420 );
and \U$31942 ( \37588 , \9217 , \37447 );
or \U$31943 ( \37589 , \37573 , \37574 , \37575 , \37576 , \37577 , \37578 , \37579 , \37580 , \37581 , \37582 , \37583 , \37584 , \37585 , \37586 , \37587 , \37588 );
_DC ga9fa ( \37590_nGa9fa , \37589 , \37524 );
buf \U$31944 ( \37591 , \37590_nGa9fa );
xor \U$31945 ( \37592 , \37572 , \37591 );
or \U$31946 ( \37593 , \37571 , \37592 );
buf \U$31947 ( \37594 , RIb7af450_258);
and \U$31948 ( \37595 , \7237 , \37042 );
and \U$31949 ( \37596 , \7239 , \37069 );
and \U$31950 ( \37597 , \9227 , \37096 );
and \U$31951 ( \37598 , \9229 , \37123 );
and \U$31952 ( \37599 , \9231 , \37150 );
and \U$31953 ( \37600 , \9233 , \37177 );
and \U$31954 ( \37601 , \9235 , \37204 );
and \U$31955 ( \37602 , \9237 , \37231 );
and \U$31956 ( \37603 , \9239 , \37258 );
and \U$31957 ( \37604 , \9241 , \37285 );
and \U$31958 ( \37605 , \9243 , \37312 );
and \U$31959 ( \37606 , \9245 , \37339 );
and \U$31960 ( \37607 , \9247 , \37366 );
and \U$31961 ( \37608 , \9249 , \37393 );
and \U$31962 ( \37609 , \9251 , \37420 );
and \U$31963 ( \37610 , \9253 , \37447 );
or \U$31964 ( \37611 , \37595 , \37596 , \37597 , \37598 , \37599 , \37600 , \37601 , \37602 , \37603 , \37604 , \37605 , \37606 , \37607 , \37608 , \37609 , \37610 );
_DC gaa10 ( \37612_nGaa10 , \37611 , \37524 );
buf \U$31965 ( \37613 , \37612_nGaa10 );
xor \U$31966 ( \37614 , \37594 , \37613 );
or \U$31967 ( \37615 , \37593 , \37614 );
buf \U$31968 ( \37616 , RIb7af3d8_259);
and \U$31969 ( \37617 , \7247 , \37042 );
and \U$31970 ( \37618 , \7249 , \37069 );
and \U$31971 ( \37619 , \9263 , \37096 );
and \U$31972 ( \37620 , \9265 , \37123 );
and \U$31973 ( \37621 , \9267 , \37150 );
and \U$31974 ( \37622 , \9269 , \37177 );
and \U$31975 ( \37623 , \9271 , \37204 );
and \U$31976 ( \37624 , \9273 , \37231 );
and \U$31977 ( \37625 , \9275 , \37258 );
and \U$31978 ( \37626 , \9277 , \37285 );
and \U$31979 ( \37627 , \9279 , \37312 );
and \U$31980 ( \37628 , \9281 , \37339 );
and \U$31981 ( \37629 , \9283 , \37366 );
and \U$31982 ( \37630 , \9285 , \37393 );
and \U$31983 ( \37631 , \9287 , \37420 );
and \U$31984 ( \37632 , \9289 , \37447 );
or \U$31985 ( \37633 , \37617 , \37618 , \37619 , \37620 , \37621 , \37622 , \37623 , \37624 , \37625 , \37626 , \37627 , \37628 , \37629 , \37630 , \37631 , \37632 );
_DC gaa26 ( \37634_nGaa26 , \37633 , \37524 );
buf \U$31986 ( \37635 , \37634_nGaa26 );
xor \U$31987 ( \37636 , \37616 , \37635 );
or \U$31988 ( \37637 , \37615 , \37636 );
buf \U$31989 ( \37638 , RIb7a5bf8_260);
and \U$31990 ( \37639 , \7257 , \37042 );
and \U$31991 ( \37640 , \7259 , \37069 );
and \U$31992 ( \37641 , \9299 , \37096 );
and \U$31993 ( \37642 , \9301 , \37123 );
and \U$31994 ( \37643 , \9303 , \37150 );
and \U$31995 ( \37644 , \9305 , \37177 );
and \U$31996 ( \37645 , \9307 , \37204 );
and \U$31997 ( \37646 , \9309 , \37231 );
and \U$31998 ( \37647 , \9311 , \37258 );
and \U$31999 ( \37648 , \9313 , \37285 );
and \U$32000 ( \37649 , \9315 , \37312 );
and \U$32001 ( \37650 , \9317 , \37339 );
and \U$32002 ( \37651 , \9319 , \37366 );
and \U$32003 ( \37652 , \9321 , \37393 );
and \U$32004 ( \37653 , \9323 , \37420 );
and \U$32005 ( \37654 , \9325 , \37447 );
or \U$32006 ( \37655 , \37639 , \37640 , \37641 , \37642 , \37643 , \37644 , \37645 , \37646 , \37647 , \37648 , \37649 , \37650 , \37651 , \37652 , \37653 , \37654 );
_DC gaa3c ( \37656_nGaa3c , \37655 , \37524 );
buf \U$32007 ( \37657 , \37656_nGaa3c );
xor \U$32008 ( \37658 , \37638 , \37657 );
or \U$32009 ( \37659 , \37637 , \37658 );
buf \U$32010 ( \37660 , RIb7a0c48_261);
and \U$32011 ( \37661 , \7267 , \37042 );
and \U$32012 ( \37662 , \7269 , \37069 );
and \U$32013 ( \37663 , \9335 , \37096 );
and \U$32014 ( \37664 , \9337 , \37123 );
and \U$32015 ( \37665 , \9339 , \37150 );
and \U$32016 ( \37666 , \9341 , \37177 );
and \U$32017 ( \37667 , \9343 , \37204 );
and \U$32018 ( \37668 , \9345 , \37231 );
and \U$32019 ( \37669 , \9347 , \37258 );
and \U$32020 ( \37670 , \9349 , \37285 );
and \U$32021 ( \37671 , \9351 , \37312 );
and \U$32022 ( \37672 , \9353 , \37339 );
and \U$32023 ( \37673 , \9355 , \37366 );
and \U$32024 ( \37674 , \9357 , \37393 );
and \U$32025 ( \37675 , \9359 , \37420 );
and \U$32026 ( \37676 , \9361 , \37447 );
or \U$32027 ( \37677 , \37661 , \37662 , \37663 , \37664 , \37665 , \37666 , \37667 , \37668 , \37669 , \37670 , \37671 , \37672 , \37673 , \37674 , \37675 , \37676 );
_DC gaa52 ( \37678_nGaa52 , \37677 , \37524 );
buf \U$32028 ( \37679 , \37678_nGaa52 );
xor \U$32029 ( \37680 , \37660 , \37679 );
or \U$32030 ( \37681 , \37659 , \37680 );
not \U$32031 ( \37682 , \37681 );
buf \U$32032 ( \37683 , \37682 );
and \U$32033 ( \37684 , \37015 , \37683 );
_HMUX gaa59 ( \37685_nGaa59 , \35410_nGa16d , \35819 , \37684 );
buf \U$32034 ( \37686 , \35429 );
buf \U$32035 ( \37687 , \35426 );
buf \U$32036 ( \37688 , \35412 );
buf \U$32037 ( \37689 , \35415 );
buf \U$32038 ( \37690 , \35418 );
buf \U$32039 ( \37691 , \35422 );
or \U$32040 ( \37692 , \37688 , \37689 , \37690 , \37691 );
and \U$32041 ( \37693 , \37687 , \37692 );
or \U$32042 ( \37694 , \37686 , \37693 );
buf \U$32043 ( \37695 , \37694 );
_HMUX gaa64 ( \37696_nGaa64 , \35818_nGa306 , \37685_nGaa59 , \37695 );
buf \U$32044 ( \37697 , RIe5319e0_6884);
not \U$32045 ( \37698 , \37697 );
buf \U$32046 ( \37699 , \37698 );
buf \U$32047 ( \37700 , RIe549ef0_6842);
xor \U$32048 ( \37701 , \37700 , \37697 );
buf \U$32049 ( \37702 , \37701 );
buf \U$32050 ( \37703 , RIe549770_6843);
and \U$32051 ( \37704 , \37700 , \37697 );
xor \U$32052 ( \37705 , \37703 , \37704 );
buf \U$32053 ( \37706 , \37705 );
buf \U$32054 ( \37707 , RIe548ff0_6844);
and \U$32055 ( \37708 , \37703 , \37704 );
xor \U$32056 ( \37709 , \37707 , \37708 );
buf \U$32057 ( \37710 , \37709 );
buf \U$32058 ( \37711 , RIea91330_6888);
and \U$32059 ( \37712 , \37707 , \37708 );
xor \U$32060 ( \37713 , \37711 , \37712 );
buf \U$32061 ( \37714 , \37713 );
not \U$32062 ( \37715 , \37714 );
and \U$32063 ( \37716 , \37711 , \37712 );
buf \U$32064 ( \37717 , \37716 );
nor \U$32065 ( \37718 , \37699 , \37702 , \37706 , \37710 , \37715 , \37717 );
and \U$32066 ( \37719 , RIe5329d0_6883, \37718 );
not \U$32067 ( \37720 , \37717 );
and \U$32068 ( \37721 , \37699 , \37702 , \37706 , \37710 , \37715 , \37720 );
and \U$32069 ( \37722 , RIeb72150_6905, \37721 );
not \U$32070 ( \37723 , \37699 );
and \U$32071 ( \37724 , \37723 , \37702 , \37706 , \37710 , \37715 , \37720 );
and \U$32072 ( \37725 , RIeab80c0_6897, \37724 );
not \U$32073 ( \37726 , \37702 );
and \U$32074 ( \37727 , \37699 , \37726 , \37706 , \37710 , \37715 , \37720 );
and \U$32075 ( \37728 , RIe5331c8_6882, \37727 );
and \U$32076 ( \37729 , \37723 , \37726 , \37706 , \37710 , \37715 , \37720 );
and \U$32077 ( \37730 , RIe5339c0_6881, \37729 );
not \U$32078 ( \37731 , \37706 );
and \U$32079 ( \37732 , \37699 , \37702 , \37731 , \37710 , \37715 , \37720 );
and \U$32080 ( \37733 , RIeab87c8_6898, \37732 );
and \U$32081 ( \37734 , \37723 , \37702 , \37731 , \37710 , \37715 , \37720 );
and \U$32082 ( \37735 , RIe5341b8_6880, \37734 );
and \U$32083 ( \37736 , \37699 , \37726 , \37731 , \37710 , \37715 , \37720 );
and \U$32084 ( \37737 , RIe5349b0_6879, \37736 );
and \U$32085 ( \37738 , \37723 , \37726 , \37731 , \37710 , \37715 , \37720 );
and \U$32086 ( \37739 , RIea94af8_6890, \37738 );
nor \U$32087 ( \37740 , \37723 , \37726 , \37731 , \37710 , \37714 , \37717 );
and \U$32088 ( \37741 , RIe5351a8_6878, \37740 );
nor \U$32089 ( \37742 , \37699 , \37726 , \37731 , \37710 , \37714 , \37717 );
and \U$32090 ( \37743 , RIe5359a0_6877, \37742 );
nor \U$32091 ( \37744 , \37723 , \37702 , \37731 , \37710 , \37714 , \37717 );
and \U$32092 ( \37745 , RIeab78c8_6895, \37744 );
nor \U$32093 ( \37746 , \37699 , \37702 , \37731 , \37710 , \37714 , \37717 );
and \U$32094 ( \37747 , RIeab7d00_6896, \37746 );
nor \U$32095 ( \37748 , \37723 , \37726 , \37706 , \37710 , \37714 , \37717 );
and \U$32096 ( \37749 , RIeacfa18_6902, \37748 );
nor \U$32097 ( \37750 , \37699 , \37726 , \37706 , \37710 , \37714 , \37717 );
and \U$32098 ( \37751 , RIeab6518_6891, \37750 );
nor \U$32099 ( \37752 , \37723 , \37702 , \37706 , \37710 , \37714 , \37717 );
and \U$32100 ( \37753 , RIeb352c8_6904, \37752 );
or \U$32101 ( \37754 , \37719 , \37722 , \37725 , \37728 , \37730 , \37733 , \37735 , \37737 , \37739 , \37741 , \37743 , \37745 , \37747 , \37749 , \37751 , \37753 );
buf \U$32103 ( \37755 , \37717 );
buf \U$32104 ( \37756 , \37714 );
buf \U$32105 ( \37757 , \37699 );
buf \U$32106 ( \37758 , \37702 );
buf \U$32107 ( \37759 , \37706 );
buf \U$32108 ( \37760 , \37710 );
or \U$32109 ( \37761 , \37757 , \37758 , \37759 , \37760 );
and \U$32110 ( \37762 , \37756 , \37761 );
or \U$32111 ( \37763 , \37755 , \37762 );
buf \U$32112 ( \37764 , \37763 );
or \U$32113 ( \37765 , 1'b0 , \37764 );
_DC gaaaa ( \37766_nGaaaa , \37754 , \37765 );
not \U$32114 ( \37767 , \37766_nGaaaa );
buf \U$32115 ( \37768 , RIb7b9608_246);
and \U$32116 ( \37769 , \7117 , \37718 );
and \U$32117 ( \37770 , \7119 , \37721 );
and \U$32118 ( \37771 , \7864 , \37724 );
and \U$32119 ( \37772 , \7892 , \37727 );
and \U$32120 ( \37773 , \7920 , \37729 );
and \U$32121 ( \37774 , \7948 , \37732 );
and \U$32122 ( \37775 , \7976 , \37734 );
and \U$32123 ( \37776 , \8004 , \37736 );
and \U$32124 ( \37777 , \8032 , \37738 );
and \U$32125 ( \37778 , \8060 , \37740 );
and \U$32126 ( \37779 , \8088 , \37742 );
and \U$32127 ( \37780 , \8116 , \37744 );
and \U$32128 ( \37781 , \8144 , \37746 );
and \U$32129 ( \37782 , \8172 , \37748 );
and \U$32130 ( \37783 , \8200 , \37750 );
and \U$32131 ( \37784 , \8228 , \37752 );
or \U$32132 ( \37785 , \37769 , \37770 , \37771 , \37772 , \37773 , \37774 , \37775 , \37776 , \37777 , \37778 , \37779 , \37780 , \37781 , \37782 , \37783 , \37784 );
_DC gaabe ( \37786_nGaabe , \37785 , \37765 );
buf \U$32133 ( \37787 , \37786_nGaabe );
xor \U$32134 ( \37788 , \37768 , \37787 );
buf \U$32135 ( \37789 , RIb7b9590_247);
and \U$32136 ( \37790 , \7126 , \37718 );
and \U$32137 ( \37791 , \7128 , \37721 );
and \U$32138 ( \37792 , \8338 , \37724 );
and \U$32139 ( \37793 , \8340 , \37727 );
and \U$32140 ( \37794 , \8342 , \37729 );
and \U$32141 ( \37795 , \8344 , \37732 );
and \U$32142 ( \37796 , \8346 , \37734 );
and \U$32143 ( \37797 , \8348 , \37736 );
and \U$32144 ( \37798 , \8350 , \37738 );
and \U$32145 ( \37799 , \8352 , \37740 );
and \U$32146 ( \37800 , \8354 , \37742 );
and \U$32147 ( \37801 , \8356 , \37744 );
and \U$32148 ( \37802 , \8358 , \37746 );
and \U$32149 ( \37803 , \8360 , \37748 );
and \U$32150 ( \37804 , \8362 , \37750 );
and \U$32151 ( \37805 , \8364 , \37752 );
or \U$32152 ( \37806 , \37790 , \37791 , \37792 , \37793 , \37794 , \37795 , \37796 , \37797 , \37798 , \37799 , \37800 , \37801 , \37802 , \37803 , \37804 , \37805 );
_DC gaad3 ( \37807_nGaad3 , \37806 , \37765 );
buf \U$32153 ( \37808 , \37807_nGaad3 );
xor \U$32154 ( \37809 , \37789 , \37808 );
or \U$32155 ( \37810 , \37788 , \37809 );
buf \U$32156 ( \37811 , RIb7b9518_248);
and \U$32157 ( \37812 , \7136 , \37718 );
and \U$32158 ( \37813 , \7138 , \37721 );
and \U$32159 ( \37814 , \8374 , \37724 );
and \U$32160 ( \37815 , \8376 , \37727 );
and \U$32161 ( \37816 , \8378 , \37729 );
and \U$32162 ( \37817 , \8380 , \37732 );
and \U$32163 ( \37818 , \8382 , \37734 );
and \U$32164 ( \37819 , \8384 , \37736 );
and \U$32165 ( \37820 , \8386 , \37738 );
and \U$32166 ( \37821 , \8388 , \37740 );
and \U$32167 ( \37822 , \8390 , \37742 );
and \U$32168 ( \37823 , \8392 , \37744 );
and \U$32169 ( \37824 , \8394 , \37746 );
and \U$32170 ( \37825 , \8396 , \37748 );
and \U$32171 ( \37826 , \8398 , \37750 );
and \U$32172 ( \37827 , \8400 , \37752 );
or \U$32173 ( \37828 , \37812 , \37813 , \37814 , \37815 , \37816 , \37817 , \37818 , \37819 , \37820 , \37821 , \37822 , \37823 , \37824 , \37825 , \37826 , \37827 );
_DC gaae9 ( \37829_nGaae9 , \37828 , \37765 );
buf \U$32174 ( \37830 , \37829_nGaae9 );
xor \U$32175 ( \37831 , \37811 , \37830 );
or \U$32176 ( \37832 , \37810 , \37831 );
buf \U$32177 ( \37833 , RIb7b94a0_249);
and \U$32178 ( \37834 , \7146 , \37718 );
and \U$32179 ( \37835 , \7148 , \37721 );
and \U$32180 ( \37836 , \8410 , \37724 );
and \U$32181 ( \37837 , \8412 , \37727 );
and \U$32182 ( \37838 , \8414 , \37729 );
and \U$32183 ( \37839 , \8416 , \37732 );
and \U$32184 ( \37840 , \8418 , \37734 );
and \U$32185 ( \37841 , \8420 , \37736 );
and \U$32186 ( \37842 , \8422 , \37738 );
and \U$32187 ( \37843 , \8424 , \37740 );
and \U$32188 ( \37844 , \8426 , \37742 );
and \U$32189 ( \37845 , \8428 , \37744 );
and \U$32190 ( \37846 , \8430 , \37746 );
and \U$32191 ( \37847 , \8432 , \37748 );
and \U$32192 ( \37848 , \8434 , \37750 );
and \U$32193 ( \37849 , \8436 , \37752 );
or \U$32194 ( \37850 , \37834 , \37835 , \37836 , \37837 , \37838 , \37839 , \37840 , \37841 , \37842 , \37843 , \37844 , \37845 , \37846 , \37847 , \37848 , \37849 );
_DC gaaff ( \37851_nGaaff , \37850 , \37765 );
buf \U$32195 ( \37852 , \37851_nGaaff );
xor \U$32196 ( \37853 , \37833 , \37852 );
or \U$32197 ( \37854 , \37832 , \37853 );
buf \U$32198 ( \37855 , RIb7b9428_250);
and \U$32199 ( \37856 , \7156 , \37718 );
and \U$32200 ( \37857 , \7158 , \37721 );
and \U$32201 ( \37858 , \8446 , \37724 );
and \U$32202 ( \37859 , \8448 , \37727 );
and \U$32203 ( \37860 , \8450 , \37729 );
and \U$32204 ( \37861 , \8452 , \37732 );
and \U$32205 ( \37862 , \8454 , \37734 );
and \U$32206 ( \37863 , \8456 , \37736 );
and \U$32207 ( \37864 , \8458 , \37738 );
and \U$32208 ( \37865 , \8460 , \37740 );
and \U$32209 ( \37866 , \8462 , \37742 );
and \U$32210 ( \37867 , \8464 , \37744 );
and \U$32211 ( \37868 , \8466 , \37746 );
and \U$32212 ( \37869 , \8468 , \37748 );
and \U$32213 ( \37870 , \8470 , \37750 );
and \U$32214 ( \37871 , \8472 , \37752 );
or \U$32215 ( \37872 , \37856 , \37857 , \37858 , \37859 , \37860 , \37861 , \37862 , \37863 , \37864 , \37865 , \37866 , \37867 , \37868 , \37869 , \37870 , \37871 );
_DC gab15 ( \37873_nGab15 , \37872 , \37765 );
buf \U$32216 ( \37874 , \37873_nGab15 );
xor \U$32217 ( \37875 , \37855 , \37874 );
or \U$32218 ( \37876 , \37854 , \37875 );
buf \U$32219 ( \37877 , RIb7b93b0_251);
and \U$32220 ( \37878 , \7166 , \37718 );
and \U$32221 ( \37879 , \7168 , \37721 );
and \U$32222 ( \37880 , \8482 , \37724 );
and \U$32223 ( \37881 , \8484 , \37727 );
and \U$32224 ( \37882 , \8486 , \37729 );
and \U$32225 ( \37883 , \8488 , \37732 );
and \U$32226 ( \37884 , \8490 , \37734 );
and \U$32227 ( \37885 , \8492 , \37736 );
and \U$32228 ( \37886 , \8494 , \37738 );
and \U$32229 ( \37887 , \8496 , \37740 );
and \U$32230 ( \37888 , \8498 , \37742 );
and \U$32231 ( \37889 , \8500 , \37744 );
and \U$32232 ( \37890 , \8502 , \37746 );
and \U$32233 ( \37891 , \8504 , \37748 );
and \U$32234 ( \37892 , \8506 , \37750 );
and \U$32235 ( \37893 , \8508 , \37752 );
or \U$32236 ( \37894 , \37878 , \37879 , \37880 , \37881 , \37882 , \37883 , \37884 , \37885 , \37886 , \37887 , \37888 , \37889 , \37890 , \37891 , \37892 , \37893 );
_DC gab2b ( \37895_nGab2b , \37894 , \37765 );
buf \U$32237 ( \37896 , \37895_nGab2b );
xor \U$32238 ( \37897 , \37877 , \37896 );
or \U$32239 ( \37898 , \37876 , \37897 );
buf \U$32240 ( \37899 , RIb7af720_252);
and \U$32241 ( \37900 , \7176 , \37718 );
and \U$32242 ( \37901 , \7178 , \37721 );
and \U$32243 ( \37902 , \8518 , \37724 );
and \U$32244 ( \37903 , \8520 , \37727 );
and \U$32245 ( \37904 , \8522 , \37729 );
and \U$32246 ( \37905 , \8524 , \37732 );
and \U$32247 ( \37906 , \8526 , \37734 );
and \U$32248 ( \37907 , \8528 , \37736 );
and \U$32249 ( \37908 , \8530 , \37738 );
and \U$32250 ( \37909 , \8532 , \37740 );
and \U$32251 ( \37910 , \8534 , \37742 );
and \U$32252 ( \37911 , \8536 , \37744 );
and \U$32253 ( \37912 , \8538 , \37746 );
and \U$32254 ( \37913 , \8540 , \37748 );
and \U$32255 ( \37914 , \8542 , \37750 );
and \U$32256 ( \37915 , \8544 , \37752 );
or \U$32257 ( \37916 , \37900 , \37901 , \37902 , \37903 , \37904 , \37905 , \37906 , \37907 , \37908 , \37909 , \37910 , \37911 , \37912 , \37913 , \37914 , \37915 );
_DC gab41 ( \37917_nGab41 , \37916 , \37765 );
buf \U$32258 ( \37918 , \37917_nGab41 );
xor \U$32259 ( \37919 , \37899 , \37918 );
or \U$32260 ( \37920 , \37898 , \37919 );
buf \U$32261 ( \37921 , RIb7af6a8_253);
and \U$32262 ( \37922 , \7186 , \37718 );
and \U$32263 ( \37923 , \7188 , \37721 );
and \U$32264 ( \37924 , \8554 , \37724 );
and \U$32265 ( \37925 , \8556 , \37727 );
and \U$32266 ( \37926 , \8558 , \37729 );
and \U$32267 ( \37927 , \8560 , \37732 );
and \U$32268 ( \37928 , \8562 , \37734 );
and \U$32269 ( \37929 , \8564 , \37736 );
and \U$32270 ( \37930 , \8566 , \37738 );
and \U$32271 ( \37931 , \8568 , \37740 );
and \U$32272 ( \37932 , \8570 , \37742 );
and \U$32273 ( \37933 , \8572 , \37744 );
and \U$32274 ( \37934 , \8574 , \37746 );
and \U$32275 ( \37935 , \8576 , \37748 );
and \U$32276 ( \37936 , \8578 , \37750 );
and \U$32277 ( \37937 , \8580 , \37752 );
or \U$32278 ( \37938 , \37922 , \37923 , \37924 , \37925 , \37926 , \37927 , \37928 , \37929 , \37930 , \37931 , \37932 , \37933 , \37934 , \37935 , \37936 , \37937 );
_DC gab57 ( \37939_nGab57 , \37938 , \37765 );
buf \U$32279 ( \37940 , \37939_nGab57 );
xor \U$32280 ( \37941 , \37921 , \37940 );
or \U$32281 ( \37942 , \37920 , \37941 );
not \U$32282 ( \37943 , \37942 );
buf \U$32283 ( \37944 , \37943 );
buf \U$32284 ( \37945 , RIb7af630_254);
and \U$32285 ( \37946 , \7198 , \37718 );
and \U$32286 ( \37947 , \7200 , \37721 );
and \U$32287 ( \37948 , \8645 , \37724 );
and \U$32288 ( \37949 , \8673 , \37727 );
and \U$32289 ( \37950 , \8701 , \37729 );
and \U$32290 ( \37951 , \8729 , \37732 );
and \U$32291 ( \37952 , \8757 , \37734 );
and \U$32292 ( \37953 , \8785 , \37736 );
and \U$32293 ( \37954 , \8813 , \37738 );
and \U$32294 ( \37955 , \8841 , \37740 );
and \U$32295 ( \37956 , \8869 , \37742 );
and \U$32296 ( \37957 , \8897 , \37744 );
and \U$32297 ( \37958 , \8925 , \37746 );
and \U$32298 ( \37959 , \8953 , \37748 );
and \U$32299 ( \37960 , \8981 , \37750 );
and \U$32300 ( \37961 , \9009 , \37752 );
or \U$32301 ( \37962 , \37946 , \37947 , \37948 , \37949 , \37950 , \37951 , \37952 , \37953 , \37954 , \37955 , \37956 , \37957 , \37958 , \37959 , \37960 , \37961 );
_DC gab6f ( \37963_nGab6f , \37962 , \37765 );
buf \U$32302 ( \37964 , \37963_nGab6f );
xor \U$32303 ( \37965 , \37945 , \37964 );
buf \U$32304 ( \37966 , RIb7af5b8_255);
and \U$32305 ( \37967 , \7207 , \37718 );
and \U$32306 ( \37968 , \7209 , \37721 );
and \U$32307 ( \37969 , \9119 , \37724 );
and \U$32308 ( \37970 , \9121 , \37727 );
and \U$32309 ( \37971 , \9123 , \37729 );
and \U$32310 ( \37972 , \9125 , \37732 );
and \U$32311 ( \37973 , \9127 , \37734 );
and \U$32312 ( \37974 , \9129 , \37736 );
and \U$32313 ( \37975 , \9131 , \37738 );
and \U$32314 ( \37976 , \9133 , \37740 );
and \U$32315 ( \37977 , \9135 , \37742 );
and \U$32316 ( \37978 , \9137 , \37744 );
and \U$32317 ( \37979 , \9139 , \37746 );
and \U$32318 ( \37980 , \9141 , \37748 );
and \U$32319 ( \37981 , \9143 , \37750 );
and \U$32320 ( \37982 , \9145 , \37752 );
or \U$32321 ( \37983 , \37967 , \37968 , \37969 , \37970 , \37971 , \37972 , \37973 , \37974 , \37975 , \37976 , \37977 , \37978 , \37979 , \37980 , \37981 , \37982 );
_DC gab84 ( \37984_nGab84 , \37983 , \37765 );
buf \U$32322 ( \37985 , \37984_nGab84 );
xor \U$32323 ( \37986 , \37966 , \37985 );
or \U$32324 ( \37987 , \37965 , \37986 );
buf \U$32325 ( \37988 , RIb7af540_256);
and \U$32326 ( \37989 , \7217 , \37718 );
and \U$32327 ( \37990 , \7219 , \37721 );
and \U$32328 ( \37991 , \9155 , \37724 );
and \U$32329 ( \37992 , \9157 , \37727 );
and \U$32330 ( \37993 , \9159 , \37729 );
and \U$32331 ( \37994 , \9161 , \37732 );
and \U$32332 ( \37995 , \9163 , \37734 );
and \U$32333 ( \37996 , \9165 , \37736 );
and \U$32334 ( \37997 , \9167 , \37738 );
and \U$32335 ( \37998 , \9169 , \37740 );
and \U$32336 ( \37999 , \9171 , \37742 );
and \U$32337 ( \38000 , \9173 , \37744 );
and \U$32338 ( \38001 , \9175 , \37746 );
and \U$32339 ( \38002 , \9177 , \37748 );
and \U$32340 ( \38003 , \9179 , \37750 );
and \U$32341 ( \38004 , \9181 , \37752 );
or \U$32342 ( \38005 , \37989 , \37990 , \37991 , \37992 , \37993 , \37994 , \37995 , \37996 , \37997 , \37998 , \37999 , \38000 , \38001 , \38002 , \38003 , \38004 );
_DC gab9a ( \38006_nGab9a , \38005 , \37765 );
buf \U$32343 ( \38007 , \38006_nGab9a );
xor \U$32344 ( \38008 , \37988 , \38007 );
or \U$32345 ( \38009 , \37987 , \38008 );
buf \U$32346 ( \38010 , RIb7af4c8_257);
and \U$32347 ( \38011 , \7227 , \37718 );
and \U$32348 ( \38012 , \7229 , \37721 );
and \U$32349 ( \38013 , \9191 , \37724 );
and \U$32350 ( \38014 , \9193 , \37727 );
and \U$32351 ( \38015 , \9195 , \37729 );
and \U$32352 ( \38016 , \9197 , \37732 );
and \U$32353 ( \38017 , \9199 , \37734 );
and \U$32354 ( \38018 , \9201 , \37736 );
and \U$32355 ( \38019 , \9203 , \37738 );
and \U$32356 ( \38020 , \9205 , \37740 );
and \U$32357 ( \38021 , \9207 , \37742 );
and \U$32358 ( \38022 , \9209 , \37744 );
and \U$32359 ( \38023 , \9211 , \37746 );
and \U$32360 ( \38024 , \9213 , \37748 );
and \U$32361 ( \38025 , \9215 , \37750 );
and \U$32362 ( \38026 , \9217 , \37752 );
or \U$32363 ( \38027 , \38011 , \38012 , \38013 , \38014 , \38015 , \38016 , \38017 , \38018 , \38019 , \38020 , \38021 , \38022 , \38023 , \38024 , \38025 , \38026 );
_DC gabb0 ( \38028_nGabb0 , \38027 , \37765 );
buf \U$32364 ( \38029 , \38028_nGabb0 );
xor \U$32365 ( \38030 , \38010 , \38029 );
or \U$32366 ( \38031 , \38009 , \38030 );
buf \U$32367 ( \38032 , RIb7af450_258);
and \U$32368 ( \38033 , \7237 , \37718 );
and \U$32369 ( \38034 , \7239 , \37721 );
and \U$32370 ( \38035 , \9227 , \37724 );
and \U$32371 ( \38036 , \9229 , \37727 );
and \U$32372 ( \38037 , \9231 , \37729 );
and \U$32373 ( \38038 , \9233 , \37732 );
and \U$32374 ( \38039 , \9235 , \37734 );
and \U$32375 ( \38040 , \9237 , \37736 );
and \U$32376 ( \38041 , \9239 , \37738 );
and \U$32377 ( \38042 , \9241 , \37740 );
and \U$32378 ( \38043 , \9243 , \37742 );
and \U$32379 ( \38044 , \9245 , \37744 );
and \U$32380 ( \38045 , \9247 , \37746 );
and \U$32381 ( \38046 , \9249 , \37748 );
and \U$32382 ( \38047 , \9251 , \37750 );
and \U$32383 ( \38048 , \9253 , \37752 );
or \U$32384 ( \38049 , \38033 , \38034 , \38035 , \38036 , \38037 , \38038 , \38039 , \38040 , \38041 , \38042 , \38043 , \38044 , \38045 , \38046 , \38047 , \38048 );
_DC gabc6 ( \38050_nGabc6 , \38049 , \37765 );
buf \U$32385 ( \38051 , \38050_nGabc6 );
xor \U$32386 ( \38052 , \38032 , \38051 );
or \U$32387 ( \38053 , \38031 , \38052 );
buf \U$32388 ( \38054 , RIb7af3d8_259);
and \U$32389 ( \38055 , \7247 , \37718 );
and \U$32390 ( \38056 , \7249 , \37721 );
and \U$32391 ( \38057 , \9263 , \37724 );
and \U$32392 ( \38058 , \9265 , \37727 );
and \U$32393 ( \38059 , \9267 , \37729 );
and \U$32394 ( \38060 , \9269 , \37732 );
and \U$32395 ( \38061 , \9271 , \37734 );
and \U$32396 ( \38062 , \9273 , \37736 );
and \U$32397 ( \38063 , \9275 , \37738 );
and \U$32398 ( \38064 , \9277 , \37740 );
and \U$32399 ( \38065 , \9279 , \37742 );
and \U$32400 ( \38066 , \9281 , \37744 );
and \U$32401 ( \38067 , \9283 , \37746 );
and \U$32402 ( \38068 , \9285 , \37748 );
and \U$32403 ( \38069 , \9287 , \37750 );
and \U$32404 ( \38070 , \9289 , \37752 );
or \U$32405 ( \38071 , \38055 , \38056 , \38057 , \38058 , \38059 , \38060 , \38061 , \38062 , \38063 , \38064 , \38065 , \38066 , \38067 , \38068 , \38069 , \38070 );
_DC gabdc ( \38072_nGabdc , \38071 , \37765 );
buf \U$32406 ( \38073 , \38072_nGabdc );
xor \U$32407 ( \38074 , \38054 , \38073 );
or \U$32408 ( \38075 , \38053 , \38074 );
buf \U$32409 ( \38076 , RIb7a5bf8_260);
and \U$32410 ( \38077 , \7257 , \37718 );
and \U$32411 ( \38078 , \7259 , \37721 );
and \U$32412 ( \38079 , \9299 , \37724 );
and \U$32413 ( \38080 , \9301 , \37727 );
and \U$32414 ( \38081 , \9303 , \37729 );
and \U$32415 ( \38082 , \9305 , \37732 );
and \U$32416 ( \38083 , \9307 , \37734 );
and \U$32417 ( \38084 , \9309 , \37736 );
and \U$32418 ( \38085 , \9311 , \37738 );
and \U$32419 ( \38086 , \9313 , \37740 );
and \U$32420 ( \38087 , \9315 , \37742 );
and \U$32421 ( \38088 , \9317 , \37744 );
and \U$32422 ( \38089 , \9319 , \37746 );
and \U$32423 ( \38090 , \9321 , \37748 );
and \U$32424 ( \38091 , \9323 , \37750 );
and \U$32425 ( \38092 , \9325 , \37752 );
or \U$32426 ( \38093 , \38077 , \38078 , \38079 , \38080 , \38081 , \38082 , \38083 , \38084 , \38085 , \38086 , \38087 , \38088 , \38089 , \38090 , \38091 , \38092 );
_DC gabf2 ( \38094_nGabf2 , \38093 , \37765 );
buf \U$32427 ( \38095 , \38094_nGabf2 );
xor \U$32428 ( \38096 , \38076 , \38095 );
or \U$32429 ( \38097 , \38075 , \38096 );
buf \U$32430 ( \38098 , RIb7a0c48_261);
and \U$32431 ( \38099 , \7267 , \37718 );
and \U$32432 ( \38100 , \7269 , \37721 );
and \U$32433 ( \38101 , \9335 , \37724 );
and \U$32434 ( \38102 , \9337 , \37727 );
and \U$32435 ( \38103 , \9339 , \37729 );
and \U$32436 ( \38104 , \9341 , \37732 );
and \U$32437 ( \38105 , \9343 , \37734 );
and \U$32438 ( \38106 , \9345 , \37736 );
and \U$32439 ( \38107 , \9347 , \37738 );
and \U$32440 ( \38108 , \9349 , \37740 );
and \U$32441 ( \38109 , \9351 , \37742 );
and \U$32442 ( \38110 , \9353 , \37744 );
and \U$32443 ( \38111 , \9355 , \37746 );
and \U$32444 ( \38112 , \9357 , \37748 );
and \U$32445 ( \38113 , \9359 , \37750 );
and \U$32446 ( \38114 , \9361 , \37752 );
or \U$32447 ( \38115 , \38099 , \38100 , \38101 , \38102 , \38103 , \38104 , \38105 , \38106 , \38107 , \38108 , \38109 , \38110 , \38111 , \38112 , \38113 , \38114 );
_DC gac08 ( \38116_nGac08 , \38115 , \37765 );
buf \U$32448 ( \38117 , \38116_nGac08 );
xor \U$32449 ( \38118 , \38098 , \38117 );
or \U$32450 ( \38119 , \38097 , \38118 );
not \U$32451 ( \38120 , \38119 );
buf \U$32452 ( \38121 , \38120 );
and \U$32453 ( \38122 , \37944 , \38121 );
and \U$32454 ( \38123 , \37767 , \38122 );
_HMUX gac10 ( \38124_nGac10 , \37696_nGaa64 , \37699 , \38123 );
buf \U$32457 ( \38125 , \37699 );
buf \U$32460 ( \38126 , \37702 );
buf \U$32463 ( \38127 , \37706 );
buf \U$32466 ( \38128 , \37710 );
buf \U$32467 ( \38129 , \37714 );
not \U$32468 ( \38130 , \38129 );
buf \U$32469 ( \38131 , \38130 );
not \U$32470 ( \38132 , \38131 );
buf \U$32471 ( \38133 , \37717 );
xnor \U$32472 ( \38134 , \38133 , \38129 );
buf \U$32473 ( \38135 , \38134 );
or \U$32474 ( \38136 , \38133 , \38129 );
not \U$32475 ( \38137 , \38136 );
buf \U$32476 ( \38138 , \38137 );
buf \U$32477 ( \38139 , \38138 );
buf \U$32478 ( \38140 , \38138 );
buf \U$32479 ( \38141 , \38138 );
buf \U$32480 ( \38142 , \38138 );
buf \U$32481 ( \38143 , \38138 );
buf \U$32482 ( \38144 , \38138 );
buf \U$32483 ( \38145 , \38138 );
buf \U$32484 ( \38146 , \38138 );
buf \U$32485 ( \38147 , \38138 );
buf \U$32486 ( \38148 , \38138 );
buf \U$32487 ( \38149 , \38138 );
buf \U$32488 ( \38150 , \38138 );
buf \U$32489 ( \38151 , \38138 );
buf \U$32490 ( \38152 , \38138 );
buf \U$32491 ( \38153 , \38138 );
buf \U$32492 ( \38154 , \38138 );
buf \U$32493 ( \38155 , \38138 );
buf \U$32494 ( \38156 , \38138 );
buf \U$32495 ( \38157 , \38138 );
buf \U$32496 ( \38158 , \38138 );
buf \U$32497 ( \38159 , \38138 );
buf \U$32498 ( \38160 , \38138 );
buf \U$32499 ( \38161 , \38138 );
buf \U$32500 ( \38162 , \38138 );
buf \U$32501 ( \38163 , \38138 );
nor \U$32502 ( \38164 , \38125 , \38126 , \38127 , \38128 , \38132 , \38135 , \38138 , \38139 , \38140 , \38141 , \38142 , \38143 , \38144 , \38145 , \38146 , \38147 , \38148 , \38149 , \38150 , \38151 , \38152 , \38153 , \38154 , \38155 , \38156 , \38157 , \38158 , \38159 , \38160 , \38161 , \38162 , \38163 );
and \U$32503 ( \38165 , RIe5329d0_6883, \38164 );
not \U$32504 ( \38166 , \38125 );
not \U$32505 ( \38167 , \38126 );
not \U$32506 ( \38168 , \38127 );
not \U$32507 ( \38169 , \38128 );
buf \U$32508 ( \38170 , \38138 );
buf \U$32509 ( \38171 , \38138 );
buf \U$32510 ( \38172 , \38138 );
buf \U$32511 ( \38173 , \38138 );
buf \U$32512 ( \38174 , \38138 );
buf \U$32513 ( \38175 , \38138 );
buf \U$32514 ( \38176 , \38138 );
buf \U$32515 ( \38177 , \38138 );
buf \U$32516 ( \38178 , \38138 );
buf \U$32517 ( \38179 , \38138 );
buf \U$32518 ( \38180 , \38138 );
buf \U$32519 ( \38181 , \38138 );
buf \U$32520 ( \38182 , \38138 );
buf \U$32521 ( \38183 , \38138 );
buf \U$32522 ( \38184 , \38138 );
buf \U$32523 ( \38185 , \38138 );
buf \U$32524 ( \38186 , \38138 );
buf \U$32525 ( \38187 , \38138 );
buf \U$32526 ( \38188 , \38138 );
buf \U$32527 ( \38189 , \38138 );
buf \U$32528 ( \38190 , \38138 );
buf \U$32529 ( \38191 , \38138 );
buf \U$32530 ( \38192 , \38138 );
buf \U$32531 ( \38193 , \38138 );
buf \U$32532 ( \38194 , \38138 );
nor \U$32533 ( \38195 , \38166 , \38167 , \38168 , \38169 , \38131 , \38135 , \38138 , \38170 , \38171 , \38172 , \38173 , \38174 , \38175 , \38176 , \38177 , \38178 , \38179 , \38180 , \38181 , \38182 , \38183 , \38184 , \38185 , \38186 , \38187 , \38188 , \38189 , \38190 , \38191 , \38192 , \38193 , \38194 );
and \U$32534 ( \38196 , RIeb72150_6905, \38195 );
buf \U$32535 ( \38197 , \38138 );
buf \U$32536 ( \38198 , \38138 );
buf \U$32537 ( \38199 , \38138 );
buf \U$32538 ( \38200 , \38138 );
buf \U$32539 ( \38201 , \38138 );
buf \U$32540 ( \38202 , \38138 );
buf \U$32541 ( \38203 , \38138 );
buf \U$32542 ( \38204 , \38138 );
buf \U$32543 ( \38205 , \38138 );
buf \U$32544 ( \38206 , \38138 );
buf \U$32545 ( \38207 , \38138 );
buf \U$32546 ( \38208 , \38138 );
buf \U$32547 ( \38209 , \38138 );
buf \U$32548 ( \38210 , \38138 );
buf \U$32549 ( \38211 , \38138 );
buf \U$32550 ( \38212 , \38138 );
buf \U$32551 ( \38213 , \38138 );
buf \U$32552 ( \38214 , \38138 );
buf \U$32553 ( \38215 , \38138 );
buf \U$32554 ( \38216 , \38138 );
buf \U$32555 ( \38217 , \38138 );
buf \U$32556 ( \38218 , \38138 );
buf \U$32557 ( \38219 , \38138 );
buf \U$32558 ( \38220 , \38138 );
buf \U$32559 ( \38221 , \38138 );
nor \U$32560 ( \38222 , \38125 , \38167 , \38168 , \38169 , \38131 , \38135 , \38138 , \38197 , \38198 , \38199 , \38200 , \38201 , \38202 , \38203 , \38204 , \38205 , \38206 , \38207 , \38208 , \38209 , \38210 , \38211 , \38212 , \38213 , \38214 , \38215 , \38216 , \38217 , \38218 , \38219 , \38220 , \38221 );
and \U$32561 ( \38223 , RIeab80c0_6897, \38222 );
buf \U$32562 ( \38224 , \38138 );
buf \U$32563 ( \38225 , \38138 );
buf \U$32564 ( \38226 , \38138 );
buf \U$32565 ( \38227 , \38138 );
buf \U$32566 ( \38228 , \38138 );
buf \U$32567 ( \38229 , \38138 );
buf \U$32568 ( \38230 , \38138 );
buf \U$32569 ( \38231 , \38138 );
buf \U$32570 ( \38232 , \38138 );
buf \U$32571 ( \38233 , \38138 );
buf \U$32572 ( \38234 , \38138 );
buf \U$32573 ( \38235 , \38138 );
buf \U$32574 ( \38236 , \38138 );
buf \U$32575 ( \38237 , \38138 );
buf \U$32576 ( \38238 , \38138 );
buf \U$32577 ( \38239 , \38138 );
buf \U$32578 ( \38240 , \38138 );
buf \U$32579 ( \38241 , \38138 );
buf \U$32580 ( \38242 , \38138 );
buf \U$32581 ( \38243 , \38138 );
buf \U$32582 ( \38244 , \38138 );
buf \U$32583 ( \38245 , \38138 );
buf \U$32584 ( \38246 , \38138 );
buf \U$32585 ( \38247 , \38138 );
buf \U$32586 ( \38248 , \38138 );
nor \U$32587 ( \38249 , \38166 , \38126 , \38168 , \38169 , \38131 , \38135 , \38138 , \38224 , \38225 , \38226 , \38227 , \38228 , \38229 , \38230 , \38231 , \38232 , \38233 , \38234 , \38235 , \38236 , \38237 , \38238 , \38239 , \38240 , \38241 , \38242 , \38243 , \38244 , \38245 , \38246 , \38247 , \38248 );
and \U$32588 ( \38250 , RIe5331c8_6882, \38249 );
buf \U$32589 ( \38251 , \38138 );
buf \U$32590 ( \38252 , \38138 );
buf \U$32591 ( \38253 , \38138 );
buf \U$32592 ( \38254 , \38138 );
buf \U$32593 ( \38255 , \38138 );
buf \U$32594 ( \38256 , \38138 );
buf \U$32595 ( \38257 , \38138 );
buf \U$32596 ( \38258 , \38138 );
buf \U$32597 ( \38259 , \38138 );
buf \U$32598 ( \38260 , \38138 );
buf \U$32599 ( \38261 , \38138 );
buf \U$32600 ( \38262 , \38138 );
buf \U$32601 ( \38263 , \38138 );
buf \U$32602 ( \38264 , \38138 );
buf \U$32603 ( \38265 , \38138 );
buf \U$32604 ( \38266 , \38138 );
buf \U$32605 ( \38267 , \38138 );
buf \U$32606 ( \38268 , \38138 );
buf \U$32607 ( \38269 , \38138 );
buf \U$32608 ( \38270 , \38138 );
buf \U$32609 ( \38271 , \38138 );
buf \U$32610 ( \38272 , \38138 );
buf \U$32611 ( \38273 , \38138 );
buf \U$32612 ( \38274 , \38138 );
buf \U$32613 ( \38275 , \38138 );
nor \U$32614 ( \38276 , \38125 , \38126 , \38168 , \38169 , \38131 , \38135 , \38138 , \38251 , \38252 , \38253 , \38254 , \38255 , \38256 , \38257 , \38258 , \38259 , \38260 , \38261 , \38262 , \38263 , \38264 , \38265 , \38266 , \38267 , \38268 , \38269 , \38270 , \38271 , \38272 , \38273 , \38274 , \38275 );
and \U$32615 ( \38277 , RIe5339c0_6881, \38276 );
buf \U$32616 ( \38278 , \38138 );
buf \U$32617 ( \38279 , \38138 );
buf \U$32618 ( \38280 , \38138 );
buf \U$32619 ( \38281 , \38138 );
buf \U$32620 ( \38282 , \38138 );
buf \U$32621 ( \38283 , \38138 );
buf \U$32622 ( \38284 , \38138 );
buf \U$32623 ( \38285 , \38138 );
buf \U$32624 ( \38286 , \38138 );
buf \U$32625 ( \38287 , \38138 );
buf \U$32626 ( \38288 , \38138 );
buf \U$32627 ( \38289 , \38138 );
buf \U$32628 ( \38290 , \38138 );
buf \U$32629 ( \38291 , \38138 );
buf \U$32630 ( \38292 , \38138 );
buf \U$32631 ( \38293 , \38138 );
buf \U$32632 ( \38294 , \38138 );
buf \U$32633 ( \38295 , \38138 );
buf \U$32634 ( \38296 , \38138 );
buf \U$32635 ( \38297 , \38138 );
buf \U$32636 ( \38298 , \38138 );
buf \U$32637 ( \38299 , \38138 );
buf \U$32638 ( \38300 , \38138 );
buf \U$32639 ( \38301 , \38138 );
buf \U$32640 ( \38302 , \38138 );
nor \U$32641 ( \38303 , \38166 , \38167 , \38127 , \38169 , \38131 , \38135 , \38138 , \38278 , \38279 , \38280 , \38281 , \38282 , \38283 , \38284 , \38285 , \38286 , \38287 , \38288 , \38289 , \38290 , \38291 , \38292 , \38293 , \38294 , \38295 , \38296 , \38297 , \38298 , \38299 , \38300 , \38301 , \38302 );
and \U$32642 ( \38304 , RIeab87c8_6898, \38303 );
buf \U$32643 ( \38305 , \38138 );
buf \U$32644 ( \38306 , \38138 );
buf \U$32645 ( \38307 , \38138 );
buf \U$32646 ( \38308 , \38138 );
buf \U$32647 ( \38309 , \38138 );
buf \U$32648 ( \38310 , \38138 );
buf \U$32649 ( \38311 , \38138 );
buf \U$32650 ( \38312 , \38138 );
buf \U$32651 ( \38313 , \38138 );
buf \U$32652 ( \38314 , \38138 );
buf \U$32653 ( \38315 , \38138 );
buf \U$32654 ( \38316 , \38138 );
buf \U$32655 ( \38317 , \38138 );
buf \U$32656 ( \38318 , \38138 );
buf \U$32657 ( \38319 , \38138 );
buf \U$32658 ( \38320 , \38138 );
buf \U$32659 ( \38321 , \38138 );
buf \U$32660 ( \38322 , \38138 );
buf \U$32661 ( \38323 , \38138 );
buf \U$32662 ( \38324 , \38138 );
buf \U$32663 ( \38325 , \38138 );
buf \U$32664 ( \38326 , \38138 );
buf \U$32665 ( \38327 , \38138 );
buf \U$32666 ( \38328 , \38138 );
buf \U$32667 ( \38329 , \38138 );
nor \U$32668 ( \38330 , \38125 , \38167 , \38127 , \38169 , \38131 , \38135 , \38138 , \38305 , \38306 , \38307 , \38308 , \38309 , \38310 , \38311 , \38312 , \38313 , \38314 , \38315 , \38316 , \38317 , \38318 , \38319 , \38320 , \38321 , \38322 , \38323 , \38324 , \38325 , \38326 , \38327 , \38328 , \38329 );
and \U$32669 ( \38331 , RIe5341b8_6880, \38330 );
buf \U$32670 ( \38332 , \38138 );
buf \U$32671 ( \38333 , \38138 );
buf \U$32672 ( \38334 , \38138 );
buf \U$32673 ( \38335 , \38138 );
buf \U$32674 ( \38336 , \38138 );
buf \U$32675 ( \38337 , \38138 );
buf \U$32676 ( \38338 , \38138 );
buf \U$32677 ( \38339 , \38138 );
buf \U$32678 ( \38340 , \38138 );
buf \U$32679 ( \38341 , \38138 );
buf \U$32680 ( \38342 , \38138 );
buf \U$32681 ( \38343 , \38138 );
buf \U$32682 ( \38344 , \38138 );
buf \U$32683 ( \38345 , \38138 );
buf \U$32684 ( \38346 , \38138 );
buf \U$32685 ( \38347 , \38138 );
buf \U$32686 ( \38348 , \38138 );
buf \U$32687 ( \38349 , \38138 );
buf \U$32688 ( \38350 , \38138 );
buf \U$32689 ( \38351 , \38138 );
buf \U$32690 ( \38352 , \38138 );
buf \U$32691 ( \38353 , \38138 );
buf \U$32692 ( \38354 , \38138 );
buf \U$32693 ( \38355 , \38138 );
buf \U$32694 ( \38356 , \38138 );
nor \U$32695 ( \38357 , \38166 , \38126 , \38127 , \38169 , \38131 , \38135 , \38138 , \38332 , \38333 , \38334 , \38335 , \38336 , \38337 , \38338 , \38339 , \38340 , \38341 , \38342 , \38343 , \38344 , \38345 , \38346 , \38347 , \38348 , \38349 , \38350 , \38351 , \38352 , \38353 , \38354 , \38355 , \38356 );
and \U$32696 ( \38358 , RIe5349b0_6879, \38357 );
buf \U$32697 ( \38359 , \38138 );
buf \U$32698 ( \38360 , \38138 );
buf \U$32699 ( \38361 , \38138 );
buf \U$32700 ( \38362 , \38138 );
buf \U$32701 ( \38363 , \38138 );
buf \U$32702 ( \38364 , \38138 );
buf \U$32703 ( \38365 , \38138 );
buf \U$32704 ( \38366 , \38138 );
buf \U$32705 ( \38367 , \38138 );
buf \U$32706 ( \38368 , \38138 );
buf \U$32707 ( \38369 , \38138 );
buf \U$32708 ( \38370 , \38138 );
buf \U$32709 ( \38371 , \38138 );
buf \U$32710 ( \38372 , \38138 );
buf \U$32711 ( \38373 , \38138 );
buf \U$32712 ( \38374 , \38138 );
buf \U$32713 ( \38375 , \38138 );
buf \U$32714 ( \38376 , \38138 );
buf \U$32715 ( \38377 , \38138 );
buf \U$32716 ( \38378 , \38138 );
buf \U$32717 ( \38379 , \38138 );
buf \U$32718 ( \38380 , \38138 );
buf \U$32719 ( \38381 , \38138 );
buf \U$32720 ( \38382 , \38138 );
buf \U$32721 ( \38383 , \38138 );
nor \U$32722 ( \38384 , \38125 , \38126 , \38127 , \38169 , \38131 , \38135 , \38138 , \38359 , \38360 , \38361 , \38362 , \38363 , \38364 , \38365 , \38366 , \38367 , \38368 , \38369 , \38370 , \38371 , \38372 , \38373 , \38374 , \38375 , \38376 , \38377 , \38378 , \38379 , \38380 , \38381 , \38382 , \38383 );
and \U$32723 ( \38385 , RIea94af8_6890, \38384 );
buf \U$32724 ( \38386 , \38138 );
buf \U$32725 ( \38387 , \38138 );
buf \U$32726 ( \38388 , \38138 );
buf \U$32727 ( \38389 , \38138 );
buf \U$32728 ( \38390 , \38138 );
buf \U$32729 ( \38391 , \38138 );
buf \U$32730 ( \38392 , \38138 );
buf \U$32731 ( \38393 , \38138 );
buf \U$32732 ( \38394 , \38138 );
buf \U$32733 ( \38395 , \38138 );
buf \U$32734 ( \38396 , \38138 );
buf \U$32735 ( \38397 , \38138 );
buf \U$32736 ( \38398 , \38138 );
buf \U$32737 ( \38399 , \38138 );
buf \U$32738 ( \38400 , \38138 );
buf \U$32739 ( \38401 , \38138 );
buf \U$32740 ( \38402 , \38138 );
buf \U$32741 ( \38403 , \38138 );
buf \U$32742 ( \38404 , \38138 );
buf \U$32743 ( \38405 , \38138 );
buf \U$32744 ( \38406 , \38138 );
buf \U$32745 ( \38407 , \38138 );
buf \U$32746 ( \38408 , \38138 );
buf \U$32747 ( \38409 , \38138 );
buf \U$32748 ( \38410 , \38138 );
nor \U$32749 ( \38411 , \38166 , \38167 , \38168 , \38128 , \38131 , \38135 , \38138 , \38386 , \38387 , \38388 , \38389 , \38390 , \38391 , \38392 , \38393 , \38394 , \38395 , \38396 , \38397 , \38398 , \38399 , \38400 , \38401 , \38402 , \38403 , \38404 , \38405 , \38406 , \38407 , \38408 , \38409 , \38410 );
and \U$32750 ( \38412 , RIe5351a8_6878, \38411 );
buf \U$32751 ( \38413 , \38138 );
buf \U$32752 ( \38414 , \38138 );
buf \U$32753 ( \38415 , \38138 );
buf \U$32754 ( \38416 , \38138 );
buf \U$32755 ( \38417 , \38138 );
buf \U$32756 ( \38418 , \38138 );
buf \U$32757 ( \38419 , \38138 );
buf \U$32758 ( \38420 , \38138 );
buf \U$32759 ( \38421 , \38138 );
buf \U$32760 ( \38422 , \38138 );
buf \U$32761 ( \38423 , \38138 );
buf \U$32762 ( \38424 , \38138 );
buf \U$32763 ( \38425 , \38138 );
buf \U$32764 ( \38426 , \38138 );
buf \U$32765 ( \38427 , \38138 );
buf \U$32766 ( \38428 , \38138 );
buf \U$32767 ( \38429 , \38138 );
buf \U$32768 ( \38430 , \38138 );
buf \U$32769 ( \38431 , \38138 );
buf \U$32770 ( \38432 , \38138 );
buf \U$32771 ( \38433 , \38138 );
buf \U$32772 ( \38434 , \38138 );
buf \U$32773 ( \38435 , \38138 );
buf \U$32774 ( \38436 , \38138 );
buf \U$32775 ( \38437 , \38138 );
nor \U$32776 ( \38438 , \38125 , \38167 , \38168 , \38128 , \38131 , \38135 , \38138 , \38413 , \38414 , \38415 , \38416 , \38417 , \38418 , \38419 , \38420 , \38421 , \38422 , \38423 , \38424 , \38425 , \38426 , \38427 , \38428 , \38429 , \38430 , \38431 , \38432 , \38433 , \38434 , \38435 , \38436 , \38437 );
and \U$32777 ( \38439 , RIe5359a0_6877, \38438 );
buf \U$32778 ( \38440 , \38138 );
buf \U$32779 ( \38441 , \38138 );
buf \U$32780 ( \38442 , \38138 );
buf \U$32781 ( \38443 , \38138 );
buf \U$32782 ( \38444 , \38138 );
buf \U$32783 ( \38445 , \38138 );
buf \U$32784 ( \38446 , \38138 );
buf \U$32785 ( \38447 , \38138 );
buf \U$32786 ( \38448 , \38138 );
buf \U$32787 ( \38449 , \38138 );
buf \U$32788 ( \38450 , \38138 );
buf \U$32789 ( \38451 , \38138 );
buf \U$32790 ( \38452 , \38138 );
buf \U$32791 ( \38453 , \38138 );
buf \U$32792 ( \38454 , \38138 );
buf \U$32793 ( \38455 , \38138 );
buf \U$32794 ( \38456 , \38138 );
buf \U$32795 ( \38457 , \38138 );
buf \U$32796 ( \38458 , \38138 );
buf \U$32797 ( \38459 , \38138 );
buf \U$32798 ( \38460 , \38138 );
buf \U$32799 ( \38461 , \38138 );
buf \U$32800 ( \38462 , \38138 );
buf \U$32801 ( \38463 , \38138 );
buf \U$32802 ( \38464 , \38138 );
nor \U$32803 ( \38465 , \38166 , \38126 , \38168 , \38128 , \38131 , \38135 , \38138 , \38440 , \38441 , \38442 , \38443 , \38444 , \38445 , \38446 , \38447 , \38448 , \38449 , \38450 , \38451 , \38452 , \38453 , \38454 , \38455 , \38456 , \38457 , \38458 , \38459 , \38460 , \38461 , \38462 , \38463 , \38464 );
and \U$32804 ( \38466 , RIeab78c8_6895, \38465 );
buf \U$32805 ( \38467 , \38138 );
buf \U$32806 ( \38468 , \38138 );
buf \U$32807 ( \38469 , \38138 );
buf \U$32808 ( \38470 , \38138 );
buf \U$32809 ( \38471 , \38138 );
buf \U$32810 ( \38472 , \38138 );
buf \U$32811 ( \38473 , \38138 );
buf \U$32812 ( \38474 , \38138 );
buf \U$32813 ( \38475 , \38138 );
buf \U$32814 ( \38476 , \38138 );
buf \U$32815 ( \38477 , \38138 );
buf \U$32816 ( \38478 , \38138 );
buf \U$32817 ( \38479 , \38138 );
buf \U$32818 ( \38480 , \38138 );
buf \U$32819 ( \38481 , \38138 );
buf \U$32820 ( \38482 , \38138 );
buf \U$32821 ( \38483 , \38138 );
buf \U$32822 ( \38484 , \38138 );
buf \U$32823 ( \38485 , \38138 );
buf \U$32824 ( \38486 , \38138 );
buf \U$32825 ( \38487 , \38138 );
buf \U$32826 ( \38488 , \38138 );
buf \U$32827 ( \38489 , \38138 );
buf \U$32828 ( \38490 , \38138 );
buf \U$32829 ( \38491 , \38138 );
nor \U$32830 ( \38492 , \38125 , \38126 , \38168 , \38128 , \38131 , \38135 , \38138 , \38467 , \38468 , \38469 , \38470 , \38471 , \38472 , \38473 , \38474 , \38475 , \38476 , \38477 , \38478 , \38479 , \38480 , \38481 , \38482 , \38483 , \38484 , \38485 , \38486 , \38487 , \38488 , \38489 , \38490 , \38491 );
and \U$32831 ( \38493 , RIeab7d00_6896, \38492 );
buf \U$32832 ( \38494 , \38138 );
buf \U$32833 ( \38495 , \38138 );
buf \U$32834 ( \38496 , \38138 );
buf \U$32835 ( \38497 , \38138 );
buf \U$32836 ( \38498 , \38138 );
buf \U$32837 ( \38499 , \38138 );
buf \U$32838 ( \38500 , \38138 );
buf \U$32839 ( \38501 , \38138 );
buf \U$32840 ( \38502 , \38138 );
buf \U$32841 ( \38503 , \38138 );
buf \U$32842 ( \38504 , \38138 );
buf \U$32843 ( \38505 , \38138 );
buf \U$32844 ( \38506 , \38138 );
buf \U$32845 ( \38507 , \38138 );
buf \U$32846 ( \38508 , \38138 );
buf \U$32847 ( \38509 , \38138 );
buf \U$32848 ( \38510 , \38138 );
buf \U$32849 ( \38511 , \38138 );
buf \U$32850 ( \38512 , \38138 );
buf \U$32851 ( \38513 , \38138 );
buf \U$32852 ( \38514 , \38138 );
buf \U$32853 ( \38515 , \38138 );
buf \U$32854 ( \38516 , \38138 );
buf \U$32855 ( \38517 , \38138 );
buf \U$32856 ( \38518 , \38138 );
nor \U$32857 ( \38519 , \38166 , \38167 , \38127 , \38128 , \38131 , \38135 , \38138 , \38494 , \38495 , \38496 , \38497 , \38498 , \38499 , \38500 , \38501 , \38502 , \38503 , \38504 , \38505 , \38506 , \38507 , \38508 , \38509 , \38510 , \38511 , \38512 , \38513 , \38514 , \38515 , \38516 , \38517 , \38518 );
and \U$32858 ( \38520 , RIeacfa18_6902, \38519 );
buf \U$32859 ( \38521 , \38138 );
buf \U$32860 ( \38522 , \38138 );
buf \U$32861 ( \38523 , \38138 );
buf \U$32862 ( \38524 , \38138 );
buf \U$32863 ( \38525 , \38138 );
buf \U$32864 ( \38526 , \38138 );
buf \U$32865 ( \38527 , \38138 );
buf \U$32866 ( \38528 , \38138 );
buf \U$32867 ( \38529 , \38138 );
buf \U$32868 ( \38530 , \38138 );
buf \U$32869 ( \38531 , \38138 );
buf \U$32870 ( \38532 , \38138 );
buf \U$32871 ( \38533 , \38138 );
buf \U$32872 ( \38534 , \38138 );
buf \U$32873 ( \38535 , \38138 );
buf \U$32874 ( \38536 , \38138 );
buf \U$32875 ( \38537 , \38138 );
buf \U$32876 ( \38538 , \38138 );
buf \U$32877 ( \38539 , \38138 );
buf \U$32878 ( \38540 , \38138 );
buf \U$32879 ( \38541 , \38138 );
buf \U$32880 ( \38542 , \38138 );
buf \U$32881 ( \38543 , \38138 );
buf \U$32882 ( \38544 , \38138 );
buf \U$32883 ( \38545 , \38138 );
nor \U$32884 ( \38546 , \38125 , \38167 , \38127 , \38128 , \38131 , \38135 , \38138 , \38521 , \38522 , \38523 , \38524 , \38525 , \38526 , \38527 , \38528 , \38529 , \38530 , \38531 , \38532 , \38533 , \38534 , \38535 , \38536 , \38537 , \38538 , \38539 , \38540 , \38541 , \38542 , \38543 , \38544 , \38545 );
and \U$32885 ( \38547 , RIeab6518_6891, \38546 );
buf \U$32886 ( \38548 , \38138 );
buf \U$32887 ( \38549 , \38138 );
buf \U$32888 ( \38550 , \38138 );
buf \U$32889 ( \38551 , \38138 );
buf \U$32890 ( \38552 , \38138 );
buf \U$32891 ( \38553 , \38138 );
buf \U$32892 ( \38554 , \38138 );
buf \U$32893 ( \38555 , \38138 );
buf \U$32894 ( \38556 , \38138 );
buf \U$32895 ( \38557 , \38138 );
buf \U$32896 ( \38558 , \38138 );
buf \U$32897 ( \38559 , \38138 );
buf \U$32898 ( \38560 , \38138 );
buf \U$32899 ( \38561 , \38138 );
buf \U$32900 ( \38562 , \38138 );
buf \U$32901 ( \38563 , \38138 );
buf \U$32902 ( \38564 , \38138 );
buf \U$32903 ( \38565 , \38138 );
buf \U$32904 ( \38566 , \38138 );
buf \U$32905 ( \38567 , \38138 );
buf \U$32906 ( \38568 , \38138 );
buf \U$32907 ( \38569 , \38138 );
buf \U$32908 ( \38570 , \38138 );
buf \U$32909 ( \38571 , \38138 );
buf \U$32910 ( \38572 , \38138 );
nor \U$32911 ( \38573 , \38166 , \38126 , \38127 , \38128 , \38131 , \38135 , \38138 , \38548 , \38549 , \38550 , \38551 , \38552 , \38553 , \38554 , \38555 , \38556 , \38557 , \38558 , \38559 , \38560 , \38561 , \38562 , \38563 , \38564 , \38565 , \38566 , \38567 , \38568 , \38569 , \38570 , \38571 , \38572 );
and \U$32912 ( \38574 , RIeb352c8_6904, \38573 );
or \U$32913 ( \38575 , \38165 , \38196 , \38223 , \38250 , \38277 , \38304 , \38331 , \38358 , \38385 , \38412 , \38439 , \38466 , \38493 , \38520 , \38547 , \38574 );
buf \U$32914 ( \38576 , \38138 );
not \U$32915 ( \38577 , \38576 );
buf \U$32916 ( \38578 , \38126 );
buf \U$32917 ( \38579 , \38127 );
buf \U$32918 ( \38580 , \38128 );
buf \U$32919 ( \38581 , \38131 );
buf \U$32920 ( \38582 , \38135 );
buf \U$32921 ( \38583 , \38138 );
buf \U$32922 ( \38584 , \38138 );
buf \U$32923 ( \38585 , \38138 );
buf \U$32924 ( \38586 , \38138 );
buf \U$32925 ( \38587 , \38138 );
buf \U$32926 ( \38588 , \38138 );
buf \U$32927 ( \38589 , \38138 );
buf \U$32928 ( \38590 , \38138 );
buf \U$32929 ( \38591 , \38138 );
buf \U$32930 ( \38592 , \38138 );
buf \U$32931 ( \38593 , \38138 );
buf \U$32932 ( \38594 , \38138 );
buf \U$32933 ( \38595 , \38138 );
buf \U$32934 ( \38596 , \38138 );
buf \U$32935 ( \38597 , \38138 );
buf \U$32936 ( \38598 , \38138 );
buf \U$32937 ( \38599 , \38138 );
buf \U$32938 ( \38600 , \38138 );
buf \U$32939 ( \38601 , \38138 );
buf \U$32940 ( \38602 , \38138 );
buf \U$32941 ( \38603 , \38138 );
buf \U$32942 ( \38604 , \38138 );
buf \U$32943 ( \38605 , \38138 );
buf \U$32944 ( \38606 , \38138 );
buf \U$32945 ( \38607 , \38138 );
buf \U$32946 ( \38608 , \38125 );
or \U$32947 ( \38609 , \38578 , \38579 , \38580 , \38581 , \38582 , \38583 , \38584 , \38585 , \38586 , \38587 , \38588 , \38589 , \38590 , \38591 , \38592 , \38593 , \38594 , \38595 , \38596 , \38597 , \38598 , \38599 , \38600 , \38601 , \38602 , \38603 , \38604 , \38605 , \38606 , \38607 , \38608 );
nand \U$32948 ( \38610 , \38577 , \38609 );
buf \U$32949 ( \38611 , \38610 );
buf \U$32950 ( \38612 , \38138 );
not \U$32951 ( \38613 , \38612 );
buf \U$32952 ( \38614 , \38135 );
buf \U$32953 ( \38615 , \38138 );
buf \U$32954 ( \38616 , \38138 );
buf \U$32955 ( \38617 , \38138 );
buf \U$32956 ( \38618 , \38138 );
buf \U$32957 ( \38619 , \38138 );
buf \U$32958 ( \38620 , \38138 );
buf \U$32959 ( \38621 , \38138 );
buf \U$32960 ( \38622 , \38138 );
buf \U$32961 ( \38623 , \38138 );
buf \U$32962 ( \38624 , \38138 );
buf \U$32963 ( \38625 , \38138 );
buf \U$32964 ( \38626 , \38138 );
buf \U$32965 ( \38627 , \38138 );
buf \U$32966 ( \38628 , \38138 );
buf \U$32967 ( \38629 , \38138 );
buf \U$32968 ( \38630 , \38138 );
buf \U$32969 ( \38631 , \38138 );
buf \U$32970 ( \38632 , \38138 );
buf \U$32971 ( \38633 , \38138 );
buf \U$32972 ( \38634 , \38138 );
buf \U$32973 ( \38635 , \38138 );
buf \U$32974 ( \38636 , \38138 );
buf \U$32975 ( \38637 , \38138 );
buf \U$32976 ( \38638 , \38138 );
buf \U$32977 ( \38639 , \38138 );
buf \U$32978 ( \38640 , \38131 );
buf \U$32979 ( \38641 , \38125 );
buf \U$32980 ( \38642 , \38126 );
buf \U$32981 ( \38643 , \38127 );
buf \U$32982 ( \38644 , \38128 );
or \U$32983 ( \38645 , \38641 , \38642 , \38643 , \38644 );
and \U$32984 ( \38646 , \38640 , \38645 );
or \U$32985 ( \38647 , \38614 , \38615 , \38616 , \38617 , \38618 , \38619 , \38620 , \38621 , \38622 , \38623 , \38624 , \38625 , \38626 , \38627 , \38628 , \38629 , \38630 , \38631 , \38632 , \38633 , \38634 , \38635 , \38636 , \38637 , \38638 , \38639 , \38646 );
and \U$32986 ( \38648 , \38613 , \38647 );
buf \U$32987 ( \38649 , \38648 );
or \U$32988 ( \38650 , \38611 , \38649 );
_DC gae27 ( \38651_nGae27 , \38575 , \38650 );
not \U$32989 ( \38652 , \38651_nGae27 );
buf \U$32990 ( \38653 , RIb7b9608_246);
buf \U$32991 ( \38654 , \38138 );
buf \U$32992 ( \38655 , \38138 );
buf \U$32993 ( \38656 , \38138 );
buf \U$32994 ( \38657 , \38138 );
buf \U$32995 ( \38658 , \38138 );
buf \U$32996 ( \38659 , \38138 );
buf \U$32997 ( \38660 , \38138 );
buf \U$32998 ( \38661 , \38138 );
buf \U$32999 ( \38662 , \38138 );
buf \U$33000 ( \38663 , \38138 );
buf \U$33001 ( \38664 , \38138 );
buf \U$33002 ( \38665 , \38138 );
buf \U$33003 ( \38666 , \38138 );
buf \U$33004 ( \38667 , \38138 );
buf \U$33005 ( \38668 , \38138 );
buf \U$33006 ( \38669 , \38138 );
buf \U$33007 ( \38670 , \38138 );
buf \U$33008 ( \38671 , \38138 );
buf \U$33009 ( \38672 , \38138 );
buf \U$33010 ( \38673 , \38138 );
buf \U$33011 ( \38674 , \38138 );
buf \U$33012 ( \38675 , \38138 );
buf \U$33013 ( \38676 , \38138 );
buf \U$33014 ( \38677 , \38138 );
buf \U$33015 ( \38678 , \38138 );
nor \U$33016 ( \38679 , \38125 , \38126 , \38127 , \38128 , \38132 , \38135 , \38138 , \38654 , \38655 , \38656 , \38657 , \38658 , \38659 , \38660 , \38661 , \38662 , \38663 , \38664 , \38665 , \38666 , \38667 , \38668 , \38669 , \38670 , \38671 , \38672 , \38673 , \38674 , \38675 , \38676 , \38677 , \38678 );
and \U$33017 ( \38680 , \7117 , \38679 );
buf \U$33018 ( \38681 , \38138 );
buf \U$33019 ( \38682 , \38138 );
buf \U$33020 ( \38683 , \38138 );
buf \U$33021 ( \38684 , \38138 );
buf \U$33022 ( \38685 , \38138 );
buf \U$33023 ( \38686 , \38138 );
buf \U$33024 ( \38687 , \38138 );
buf \U$33025 ( \38688 , \38138 );
buf \U$33026 ( \38689 , \38138 );
buf \U$33027 ( \38690 , \38138 );
buf \U$33028 ( \38691 , \38138 );
buf \U$33029 ( \38692 , \38138 );
buf \U$33030 ( \38693 , \38138 );
buf \U$33031 ( \38694 , \38138 );
buf \U$33032 ( \38695 , \38138 );
buf \U$33033 ( \38696 , \38138 );
buf \U$33034 ( \38697 , \38138 );
buf \U$33035 ( \38698 , \38138 );
buf \U$33036 ( \38699 , \38138 );
buf \U$33037 ( \38700 , \38138 );
buf \U$33038 ( \38701 , \38138 );
buf \U$33039 ( \38702 , \38138 );
buf \U$33040 ( \38703 , \38138 );
buf \U$33041 ( \38704 , \38138 );
buf \U$33042 ( \38705 , \38138 );
nor \U$33043 ( \38706 , \38166 , \38167 , \38168 , \38169 , \38131 , \38135 , \38138 , \38681 , \38682 , \38683 , \38684 , \38685 , \38686 , \38687 , \38688 , \38689 , \38690 , \38691 , \38692 , \38693 , \38694 , \38695 , \38696 , \38697 , \38698 , \38699 , \38700 , \38701 , \38702 , \38703 , \38704 , \38705 );
and \U$33044 ( \38707 , \7119 , \38706 );
buf \U$33045 ( \38708 , \38138 );
buf \U$33046 ( \38709 , \38138 );
buf \U$33047 ( \38710 , \38138 );
buf \U$33048 ( \38711 , \38138 );
buf \U$33049 ( \38712 , \38138 );
buf \U$33050 ( \38713 , \38138 );
buf \U$33051 ( \38714 , \38138 );
buf \U$33052 ( \38715 , \38138 );
buf \U$33053 ( \38716 , \38138 );
buf \U$33054 ( \38717 , \38138 );
buf \U$33055 ( \38718 , \38138 );
buf \U$33056 ( \38719 , \38138 );
buf \U$33057 ( \38720 , \38138 );
buf \U$33058 ( \38721 , \38138 );
buf \U$33059 ( \38722 , \38138 );
buf \U$33060 ( \38723 , \38138 );
buf \U$33061 ( \38724 , \38138 );
buf \U$33062 ( \38725 , \38138 );
buf \U$33063 ( \38726 , \38138 );
buf \U$33064 ( \38727 , \38138 );
buf \U$33065 ( \38728 , \38138 );
buf \U$33066 ( \38729 , \38138 );
buf \U$33067 ( \38730 , \38138 );
buf \U$33068 ( \38731 , \38138 );
buf \U$33069 ( \38732 , \38138 );
nor \U$33070 ( \38733 , \38125 , \38167 , \38168 , \38169 , \38131 , \38135 , \38138 , \38708 , \38709 , \38710 , \38711 , \38712 , \38713 , \38714 , \38715 , \38716 , \38717 , \38718 , \38719 , \38720 , \38721 , \38722 , \38723 , \38724 , \38725 , \38726 , \38727 , \38728 , \38729 , \38730 , \38731 , \38732 );
and \U$33071 ( \38734 , \7864 , \38733 );
buf \U$33072 ( \38735 , \38138 );
buf \U$33073 ( \38736 , \38138 );
buf \U$33074 ( \38737 , \38138 );
buf \U$33075 ( \38738 , \38138 );
buf \U$33076 ( \38739 , \38138 );
buf \U$33077 ( \38740 , \38138 );
buf \U$33078 ( \38741 , \38138 );
buf \U$33079 ( \38742 , \38138 );
buf \U$33080 ( \38743 , \38138 );
buf \U$33081 ( \38744 , \38138 );
buf \U$33082 ( \38745 , \38138 );
buf \U$33083 ( \38746 , \38138 );
buf \U$33084 ( \38747 , \38138 );
buf \U$33085 ( \38748 , \38138 );
buf \U$33086 ( \38749 , \38138 );
buf \U$33087 ( \38750 , \38138 );
buf \U$33088 ( \38751 , \38138 );
buf \U$33089 ( \38752 , \38138 );
buf \U$33090 ( \38753 , \38138 );
buf \U$33091 ( \38754 , \38138 );
buf \U$33092 ( \38755 , \38138 );
buf \U$33093 ( \38756 , \38138 );
buf \U$33094 ( \38757 , \38138 );
buf \U$33095 ( \38758 , \38138 );
buf \U$33096 ( \38759 , \38138 );
nor \U$33097 ( \38760 , \38166 , \38126 , \38168 , \38169 , \38131 , \38135 , \38138 , \38735 , \38736 , \38737 , \38738 , \38739 , \38740 , \38741 , \38742 , \38743 , \38744 , \38745 , \38746 , \38747 , \38748 , \38749 , \38750 , \38751 , \38752 , \38753 , \38754 , \38755 , \38756 , \38757 , \38758 , \38759 );
and \U$33098 ( \38761 , \7892 , \38760 );
buf \U$33099 ( \38762 , \38138 );
buf \U$33100 ( \38763 , \38138 );
buf \U$33101 ( \38764 , \38138 );
buf \U$33102 ( \38765 , \38138 );
buf \U$33103 ( \38766 , \38138 );
buf \U$33104 ( \38767 , \38138 );
buf \U$33105 ( \38768 , \38138 );
buf \U$33106 ( \38769 , \38138 );
buf \U$33107 ( \38770 , \38138 );
buf \U$33108 ( \38771 , \38138 );
buf \U$33109 ( \38772 , \38138 );
buf \U$33110 ( \38773 , \38138 );
buf \U$33111 ( \38774 , \38138 );
buf \U$33112 ( \38775 , \38138 );
buf \U$33113 ( \38776 , \38138 );
buf \U$33114 ( \38777 , \38138 );
buf \U$33115 ( \38778 , \38138 );
buf \U$33116 ( \38779 , \38138 );
buf \U$33117 ( \38780 , \38138 );
buf \U$33118 ( \38781 , \38138 );
buf \U$33119 ( \38782 , \38138 );
buf \U$33120 ( \38783 , \38138 );
buf \U$33121 ( \38784 , \38138 );
buf \U$33122 ( \38785 , \38138 );
buf \U$33123 ( \38786 , \38138 );
nor \U$33124 ( \38787 , \38125 , \38126 , \38168 , \38169 , \38131 , \38135 , \38138 , \38762 , \38763 , \38764 , \38765 , \38766 , \38767 , \38768 , \38769 , \38770 , \38771 , \38772 , \38773 , \38774 , \38775 , \38776 , \38777 , \38778 , \38779 , \38780 , \38781 , \38782 , \38783 , \38784 , \38785 , \38786 );
and \U$33125 ( \38788 , \7920 , \38787 );
buf \U$33126 ( \38789 , \38138 );
buf \U$33127 ( \38790 , \38138 );
buf \U$33128 ( \38791 , \38138 );
buf \U$33129 ( \38792 , \38138 );
buf \U$33130 ( \38793 , \38138 );
buf \U$33131 ( \38794 , \38138 );
buf \U$33132 ( \38795 , \38138 );
buf \U$33133 ( \38796 , \38138 );
buf \U$33134 ( \38797 , \38138 );
buf \U$33135 ( \38798 , \38138 );
buf \U$33136 ( \38799 , \38138 );
buf \U$33137 ( \38800 , \38138 );
buf \U$33138 ( \38801 , \38138 );
buf \U$33139 ( \38802 , \38138 );
buf \U$33140 ( \38803 , \38138 );
buf \U$33141 ( \38804 , \38138 );
buf \U$33142 ( \38805 , \38138 );
buf \U$33143 ( \38806 , \38138 );
buf \U$33144 ( \38807 , \38138 );
buf \U$33145 ( \38808 , \38138 );
buf \U$33146 ( \38809 , \38138 );
buf \U$33147 ( \38810 , \38138 );
buf \U$33148 ( \38811 , \38138 );
buf \U$33149 ( \38812 , \38138 );
buf \U$33150 ( \38813 , \38138 );
nor \U$33151 ( \38814 , \38166 , \38167 , \38127 , \38169 , \38131 , \38135 , \38138 , \38789 , \38790 , \38791 , \38792 , \38793 , \38794 , \38795 , \38796 , \38797 , \38798 , \38799 , \38800 , \38801 , \38802 , \38803 , \38804 , \38805 , \38806 , \38807 , \38808 , \38809 , \38810 , \38811 , \38812 , \38813 );
and \U$33152 ( \38815 , \7948 , \38814 );
buf \U$33153 ( \38816 , \38138 );
buf \U$33154 ( \38817 , \38138 );
buf \U$33155 ( \38818 , \38138 );
buf \U$33156 ( \38819 , \38138 );
buf \U$33157 ( \38820 , \38138 );
buf \U$33158 ( \38821 , \38138 );
buf \U$33159 ( \38822 , \38138 );
buf \U$33160 ( \38823 , \38138 );
buf \U$33161 ( \38824 , \38138 );
buf \U$33162 ( \38825 , \38138 );
buf \U$33163 ( \38826 , \38138 );
buf \U$33164 ( \38827 , \38138 );
buf \U$33165 ( \38828 , \38138 );
buf \U$33166 ( \38829 , \38138 );
buf \U$33167 ( \38830 , \38138 );
buf \U$33168 ( \38831 , \38138 );
buf \U$33169 ( \38832 , \38138 );
buf \U$33170 ( \38833 , \38138 );
buf \U$33171 ( \38834 , \38138 );
buf \U$33172 ( \38835 , \38138 );
buf \U$33173 ( \38836 , \38138 );
buf \U$33174 ( \38837 , \38138 );
buf \U$33175 ( \38838 , \38138 );
buf \U$33176 ( \38839 , \38138 );
buf \U$33177 ( \38840 , \38138 );
nor \U$33178 ( \38841 , \38125 , \38167 , \38127 , \38169 , \38131 , \38135 , \38138 , \38816 , \38817 , \38818 , \38819 , \38820 , \38821 , \38822 , \38823 , \38824 , \38825 , \38826 , \38827 , \38828 , \38829 , \38830 , \38831 , \38832 , \38833 , \38834 , \38835 , \38836 , \38837 , \38838 , \38839 , \38840 );
and \U$33179 ( \38842 , \7976 , \38841 );
buf \U$33180 ( \38843 , \38138 );
buf \U$33181 ( \38844 , \38138 );
buf \U$33182 ( \38845 , \38138 );
buf \U$33183 ( \38846 , \38138 );
buf \U$33184 ( \38847 , \38138 );
buf \U$33185 ( \38848 , \38138 );
buf \U$33186 ( \38849 , \38138 );
buf \U$33187 ( \38850 , \38138 );
buf \U$33188 ( \38851 , \38138 );
buf \U$33189 ( \38852 , \38138 );
buf \U$33190 ( \38853 , \38138 );
buf \U$33191 ( \38854 , \38138 );
buf \U$33192 ( \38855 , \38138 );
buf \U$33193 ( \38856 , \38138 );
buf \U$33194 ( \38857 , \38138 );
buf \U$33195 ( \38858 , \38138 );
buf \U$33196 ( \38859 , \38138 );
buf \U$33197 ( \38860 , \38138 );
buf \U$33198 ( \38861 , \38138 );
buf \U$33199 ( \38862 , \38138 );
buf \U$33200 ( \38863 , \38138 );
buf \U$33201 ( \38864 , \38138 );
buf \U$33202 ( \38865 , \38138 );
buf \U$33203 ( \38866 , \38138 );
buf \U$33204 ( \38867 , \38138 );
nor \U$33205 ( \38868 , \38166 , \38126 , \38127 , \38169 , \38131 , \38135 , \38138 , \38843 , \38844 , \38845 , \38846 , \38847 , \38848 , \38849 , \38850 , \38851 , \38852 , \38853 , \38854 , \38855 , \38856 , \38857 , \38858 , \38859 , \38860 , \38861 , \38862 , \38863 , \38864 , \38865 , \38866 , \38867 );
and \U$33206 ( \38869 , \8004 , \38868 );
buf \U$33207 ( \38870 , \38138 );
buf \U$33208 ( \38871 , \38138 );
buf \U$33209 ( \38872 , \38138 );
buf \U$33210 ( \38873 , \38138 );
buf \U$33211 ( \38874 , \38138 );
buf \U$33212 ( \38875 , \38138 );
buf \U$33213 ( \38876 , \38138 );
buf \U$33214 ( \38877 , \38138 );
buf \U$33215 ( \38878 , \38138 );
buf \U$33216 ( \38879 , \38138 );
buf \U$33217 ( \38880 , \38138 );
buf \U$33218 ( \38881 , \38138 );
buf \U$33219 ( \38882 , \38138 );
buf \U$33220 ( \38883 , \38138 );
buf \U$33221 ( \38884 , \38138 );
buf \U$33222 ( \38885 , \38138 );
buf \U$33223 ( \38886 , \38138 );
buf \U$33224 ( \38887 , \38138 );
buf \U$33225 ( \38888 , \38138 );
buf \U$33226 ( \38889 , \38138 );
buf \U$33227 ( \38890 , \38138 );
buf \U$33228 ( \38891 , \38138 );
buf \U$33229 ( \38892 , \38138 );
buf \U$33230 ( \38893 , \38138 );
buf \U$33231 ( \38894 , \38138 );
nor \U$33232 ( \38895 , \38125 , \38126 , \38127 , \38169 , \38131 , \38135 , \38138 , \38870 , \38871 , \38872 , \38873 , \38874 , \38875 , \38876 , \38877 , \38878 , \38879 , \38880 , \38881 , \38882 , \38883 , \38884 , \38885 , \38886 , \38887 , \38888 , \38889 , \38890 , \38891 , \38892 , \38893 , \38894 );
and \U$33233 ( \38896 , \8032 , \38895 );
buf \U$33234 ( \38897 , \38138 );
buf \U$33235 ( \38898 , \38138 );
buf \U$33236 ( \38899 , \38138 );
buf \U$33237 ( \38900 , \38138 );
buf \U$33238 ( \38901 , \38138 );
buf \U$33239 ( \38902 , \38138 );
buf \U$33240 ( \38903 , \38138 );
buf \U$33241 ( \38904 , \38138 );
buf \U$33242 ( \38905 , \38138 );
buf \U$33243 ( \38906 , \38138 );
buf \U$33244 ( \38907 , \38138 );
buf \U$33245 ( \38908 , \38138 );
buf \U$33246 ( \38909 , \38138 );
buf \U$33247 ( \38910 , \38138 );
buf \U$33248 ( \38911 , \38138 );
buf \U$33249 ( \38912 , \38138 );
buf \U$33250 ( \38913 , \38138 );
buf \U$33251 ( \38914 , \38138 );
buf \U$33252 ( \38915 , \38138 );
buf \U$33253 ( \38916 , \38138 );
buf \U$33254 ( \38917 , \38138 );
buf \U$33255 ( \38918 , \38138 );
buf \U$33256 ( \38919 , \38138 );
buf \U$33257 ( \38920 , \38138 );
buf \U$33258 ( \38921 , \38138 );
nor \U$33259 ( \38922 , \38166 , \38167 , \38168 , \38128 , \38131 , \38135 , \38138 , \38897 , \38898 , \38899 , \38900 , \38901 , \38902 , \38903 , \38904 , \38905 , \38906 , \38907 , \38908 , \38909 , \38910 , \38911 , \38912 , \38913 , \38914 , \38915 , \38916 , \38917 , \38918 , \38919 , \38920 , \38921 );
and \U$33260 ( \38923 , \8060 , \38922 );
buf \U$33261 ( \38924 , \38138 );
buf \U$33262 ( \38925 , \38138 );
buf \U$33263 ( \38926 , \38138 );
buf \U$33264 ( \38927 , \38138 );
buf \U$33265 ( \38928 , \38138 );
buf \U$33266 ( \38929 , \38138 );
buf \U$33267 ( \38930 , \38138 );
buf \U$33268 ( \38931 , \38138 );
buf \U$33269 ( \38932 , \38138 );
buf \U$33270 ( \38933 , \38138 );
buf \U$33271 ( \38934 , \38138 );
buf \U$33272 ( \38935 , \38138 );
buf \U$33273 ( \38936 , \38138 );
buf \U$33274 ( \38937 , \38138 );
buf \U$33275 ( \38938 , \38138 );
buf \U$33276 ( \38939 , \38138 );
buf \U$33277 ( \38940 , \38138 );
buf \U$33278 ( \38941 , \38138 );
buf \U$33279 ( \38942 , \38138 );
buf \U$33280 ( \38943 , \38138 );
buf \U$33281 ( \38944 , \38138 );
buf \U$33282 ( \38945 , \38138 );
buf \U$33283 ( \38946 , \38138 );
buf \U$33284 ( \38947 , \38138 );
buf \U$33285 ( \38948 , \38138 );
nor \U$33286 ( \38949 , \38125 , \38167 , \38168 , \38128 , \38131 , \38135 , \38138 , \38924 , \38925 , \38926 , \38927 , \38928 , \38929 , \38930 , \38931 , \38932 , \38933 , \38934 , \38935 , \38936 , \38937 , \38938 , \38939 , \38940 , \38941 , \38942 , \38943 , \38944 , \38945 , \38946 , \38947 , \38948 );
and \U$33287 ( \38950 , \8088 , \38949 );
buf \U$33288 ( \38951 , \38138 );
buf \U$33289 ( \38952 , \38138 );
buf \U$33290 ( \38953 , \38138 );
buf \U$33291 ( \38954 , \38138 );
buf \U$33292 ( \38955 , \38138 );
buf \U$33293 ( \38956 , \38138 );
buf \U$33294 ( \38957 , \38138 );
buf \U$33295 ( \38958 , \38138 );
buf \U$33296 ( \38959 , \38138 );
buf \U$33297 ( \38960 , \38138 );
buf \U$33298 ( \38961 , \38138 );
buf \U$33299 ( \38962 , \38138 );
buf \U$33300 ( \38963 , \38138 );
buf \U$33301 ( \38964 , \38138 );
buf \U$33302 ( \38965 , \38138 );
buf \U$33303 ( \38966 , \38138 );
buf \U$33304 ( \38967 , \38138 );
buf \U$33305 ( \38968 , \38138 );
buf \U$33306 ( \38969 , \38138 );
buf \U$33307 ( \38970 , \38138 );
buf \U$33308 ( \38971 , \38138 );
buf \U$33309 ( \38972 , \38138 );
buf \U$33310 ( \38973 , \38138 );
buf \U$33311 ( \38974 , \38138 );
buf \U$33312 ( \38975 , \38138 );
nor \U$33313 ( \38976 , \38166 , \38126 , \38168 , \38128 , \38131 , \38135 , \38138 , \38951 , \38952 , \38953 , \38954 , \38955 , \38956 , \38957 , \38958 , \38959 , \38960 , \38961 , \38962 , \38963 , \38964 , \38965 , \38966 , \38967 , \38968 , \38969 , \38970 , \38971 , \38972 , \38973 , \38974 , \38975 );
and \U$33314 ( \38977 , \8116 , \38976 );
buf \U$33315 ( \38978 , \38138 );
buf \U$33316 ( \38979 , \38138 );
buf \U$33317 ( \38980 , \38138 );
buf \U$33318 ( \38981 , \38138 );
buf \U$33319 ( \38982 , \38138 );
buf \U$33320 ( \38983 , \38138 );
buf \U$33321 ( \38984 , \38138 );
buf \U$33322 ( \38985 , \38138 );
buf \U$33323 ( \38986 , \38138 );
buf \U$33324 ( \38987 , \38138 );
buf \U$33325 ( \38988 , \38138 );
buf \U$33326 ( \38989 , \38138 );
buf \U$33327 ( \38990 , \38138 );
buf \U$33328 ( \38991 , \38138 );
buf \U$33329 ( \38992 , \38138 );
buf \U$33330 ( \38993 , \38138 );
buf \U$33331 ( \38994 , \38138 );
buf \U$33332 ( \38995 , \38138 );
buf \U$33333 ( \38996 , \38138 );
buf \U$33334 ( \38997 , \38138 );
buf \U$33335 ( \38998 , \38138 );
buf \U$33336 ( \38999 , \38138 );
buf \U$33337 ( \39000 , \38138 );
buf \U$33338 ( \39001 , \38138 );
buf \U$33339 ( \39002 , \38138 );
nor \U$33340 ( \39003 , \38125 , \38126 , \38168 , \38128 , \38131 , \38135 , \38138 , \38978 , \38979 , \38980 , \38981 , \38982 , \38983 , \38984 , \38985 , \38986 , \38987 , \38988 , \38989 , \38990 , \38991 , \38992 , \38993 , \38994 , \38995 , \38996 , \38997 , \38998 , \38999 , \39000 , \39001 , \39002 );
and \U$33341 ( \39004 , \8144 , \39003 );
buf \U$33342 ( \39005 , \38138 );
buf \U$33343 ( \39006 , \38138 );
buf \U$33344 ( \39007 , \38138 );
buf \U$33345 ( \39008 , \38138 );
buf \U$33346 ( \39009 , \38138 );
buf \U$33347 ( \39010 , \38138 );
buf \U$33348 ( \39011 , \38138 );
buf \U$33349 ( \39012 , \38138 );
buf \U$33350 ( \39013 , \38138 );
buf \U$33351 ( \39014 , \38138 );
buf \U$33352 ( \39015 , \38138 );
buf \U$33353 ( \39016 , \38138 );
buf \U$33354 ( \39017 , \38138 );
buf \U$33355 ( \39018 , \38138 );
buf \U$33356 ( \39019 , \38138 );
buf \U$33357 ( \39020 , \38138 );
buf \U$33358 ( \39021 , \38138 );
buf \U$33359 ( \39022 , \38138 );
buf \U$33360 ( \39023 , \38138 );
buf \U$33361 ( \39024 , \38138 );
buf \U$33362 ( \39025 , \38138 );
buf \U$33363 ( \39026 , \38138 );
buf \U$33364 ( \39027 , \38138 );
buf \U$33365 ( \39028 , \38138 );
buf \U$33366 ( \39029 , \38138 );
nor \U$33367 ( \39030 , \38166 , \38167 , \38127 , \38128 , \38131 , \38135 , \38138 , \39005 , \39006 , \39007 , \39008 , \39009 , \39010 , \39011 , \39012 , \39013 , \39014 , \39015 , \39016 , \39017 , \39018 , \39019 , \39020 , \39021 , \39022 , \39023 , \39024 , \39025 , \39026 , \39027 , \39028 , \39029 );
and \U$33368 ( \39031 , \8172 , \39030 );
buf \U$33369 ( \39032 , \38138 );
buf \U$33370 ( \39033 , \38138 );
buf \U$33371 ( \39034 , \38138 );
buf \U$33372 ( \39035 , \38138 );
buf \U$33373 ( \39036 , \38138 );
buf \U$33374 ( \39037 , \38138 );
buf \U$33375 ( \39038 , \38138 );
buf \U$33376 ( \39039 , \38138 );
buf \U$33377 ( \39040 , \38138 );
buf \U$33378 ( \39041 , \38138 );
buf \U$33379 ( \39042 , \38138 );
buf \U$33380 ( \39043 , \38138 );
buf \U$33381 ( \39044 , \38138 );
buf \U$33382 ( \39045 , \38138 );
buf \U$33383 ( \39046 , \38138 );
buf \U$33384 ( \39047 , \38138 );
buf \U$33385 ( \39048 , \38138 );
buf \U$33386 ( \39049 , \38138 );
buf \U$33387 ( \39050 , \38138 );
buf \U$33388 ( \39051 , \38138 );
buf \U$33389 ( \39052 , \38138 );
buf \U$33390 ( \39053 , \38138 );
buf \U$33391 ( \39054 , \38138 );
buf \U$33392 ( \39055 , \38138 );
buf \U$33393 ( \39056 , \38138 );
nor \U$33394 ( \39057 , \38125 , \38167 , \38127 , \38128 , \38131 , \38135 , \38138 , \39032 , \39033 , \39034 , \39035 , \39036 , \39037 , \39038 , \39039 , \39040 , \39041 , \39042 , \39043 , \39044 , \39045 , \39046 , \39047 , \39048 , \39049 , \39050 , \39051 , \39052 , \39053 , \39054 , \39055 , \39056 );
and \U$33395 ( \39058 , \8200 , \39057 );
buf \U$33396 ( \39059 , \38138 );
buf \U$33397 ( \39060 , \38138 );
buf \U$33398 ( \39061 , \38138 );
buf \U$33399 ( \39062 , \38138 );
buf \U$33400 ( \39063 , \38138 );
buf \U$33401 ( \39064 , \38138 );
buf \U$33402 ( \39065 , \38138 );
buf \U$33403 ( \39066 , \38138 );
buf \U$33404 ( \39067 , \38138 );
buf \U$33405 ( \39068 , \38138 );
buf \U$33406 ( \39069 , \38138 );
buf \U$33407 ( \39070 , \38138 );
buf \U$33408 ( \39071 , \38138 );
buf \U$33409 ( \39072 , \38138 );
buf \U$33410 ( \39073 , \38138 );
buf \U$33411 ( \39074 , \38138 );
buf \U$33412 ( \39075 , \38138 );
buf \U$33413 ( \39076 , \38138 );
buf \U$33414 ( \39077 , \38138 );
buf \U$33415 ( \39078 , \38138 );
buf \U$33416 ( \39079 , \38138 );
buf \U$33417 ( \39080 , \38138 );
buf \U$33418 ( \39081 , \38138 );
buf \U$33419 ( \39082 , \38138 );
buf \U$33420 ( \39083 , \38138 );
nor \U$33421 ( \39084 , \38166 , \38126 , \38127 , \38128 , \38131 , \38135 , \38138 , \39059 , \39060 , \39061 , \39062 , \39063 , \39064 , \39065 , \39066 , \39067 , \39068 , \39069 , \39070 , \39071 , \39072 , \39073 , \39074 , \39075 , \39076 , \39077 , \39078 , \39079 , \39080 , \39081 , \39082 , \39083 );
and \U$33422 ( \39085 , \8228 , \39084 );
or \U$33423 ( \39086 , \38680 , \38707 , \38734 , \38761 , \38788 , \38815 , \38842 , \38869 , \38896 , \38923 , \38950 , \38977 , \39004 , \39031 , \39058 , \39085 );
buf \U$33424 ( \39087 , \38138 );
not \U$33425 ( \39088 , \39087 );
buf \U$33426 ( \39089 , \38126 );
buf \U$33427 ( \39090 , \38127 );
buf \U$33428 ( \39091 , \38128 );
buf \U$33429 ( \39092 , \38131 );
buf \U$33430 ( \39093 , \38135 );
buf \U$33431 ( \39094 , \38138 );
buf \U$33432 ( \39095 , \38138 );
buf \U$33433 ( \39096 , \38138 );
buf \U$33434 ( \39097 , \38138 );
buf \U$33435 ( \39098 , \38138 );
buf \U$33436 ( \39099 , \38138 );
buf \U$33437 ( \39100 , \38138 );
buf \U$33438 ( \39101 , \38138 );
buf \U$33439 ( \39102 , \38138 );
buf \U$33440 ( \39103 , \38138 );
buf \U$33441 ( \39104 , \38138 );
buf \U$33442 ( \39105 , \38138 );
buf \U$33443 ( \39106 , \38138 );
buf \U$33444 ( \39107 , \38138 );
buf \U$33445 ( \39108 , \38138 );
buf \U$33446 ( \39109 , \38138 );
buf \U$33447 ( \39110 , \38138 );
buf \U$33448 ( \39111 , \38138 );
buf \U$33449 ( \39112 , \38138 );
buf \U$33450 ( \39113 , \38138 );
buf \U$33451 ( \39114 , \38138 );
buf \U$33452 ( \39115 , \38138 );
buf \U$33453 ( \39116 , \38138 );
buf \U$33454 ( \39117 , \38138 );
buf \U$33455 ( \39118 , \38138 );
buf \U$33456 ( \39119 , \38125 );
or \U$33457 ( \39120 , \39089 , \39090 , \39091 , \39092 , \39093 , \39094 , \39095 , \39096 , \39097 , \39098 , \39099 , \39100 , \39101 , \39102 , \39103 , \39104 , \39105 , \39106 , \39107 , \39108 , \39109 , \39110 , \39111 , \39112 , \39113 , \39114 , \39115 , \39116 , \39117 , \39118 , \39119 );
nand \U$33458 ( \39121 , \39088 , \39120 );
buf \U$33459 ( \39122 , \39121 );
buf \U$33460 ( \39123 , \38138 );
not \U$33461 ( \39124 , \39123 );
buf \U$33462 ( \39125 , \38135 );
buf \U$33463 ( \39126 , \38138 );
buf \U$33464 ( \39127 , \38138 );
buf \U$33465 ( \39128 , \38138 );
buf \U$33466 ( \39129 , \38138 );
buf \U$33467 ( \39130 , \38138 );
buf \U$33468 ( \39131 , \38138 );
buf \U$33469 ( \39132 , \38138 );
buf \U$33470 ( \39133 , \38138 );
buf \U$33471 ( \39134 , \38138 );
buf \U$33472 ( \39135 , \38138 );
buf \U$33473 ( \39136 , \38138 );
buf \U$33474 ( \39137 , \38138 );
buf \U$33475 ( \39138 , \38138 );
buf \U$33476 ( \39139 , \38138 );
buf \U$33477 ( \39140 , \38138 );
buf \U$33478 ( \39141 , \38138 );
buf \U$33479 ( \39142 , \38138 );
buf \U$33480 ( \39143 , \38138 );
buf \U$33481 ( \39144 , \38138 );
buf \U$33482 ( \39145 , \38138 );
buf \U$33483 ( \39146 , \38138 );
buf \U$33484 ( \39147 , \38138 );
buf \U$33485 ( \39148 , \38138 );
buf \U$33486 ( \39149 , \38138 );
buf \U$33487 ( \39150 , \38138 );
buf \U$33488 ( \39151 , \38131 );
buf \U$33489 ( \39152 , \38125 );
buf \U$33490 ( \39153 , \38126 );
buf \U$33491 ( \39154 , \38127 );
buf \U$33492 ( \39155 , \38128 );
or \U$33493 ( \39156 , \39152 , \39153 , \39154 , \39155 );
and \U$33494 ( \39157 , \39151 , \39156 );
or \U$33495 ( \39158 , \39125 , \39126 , \39127 , \39128 , \39129 , \39130 , \39131 , \39132 , \39133 , \39134 , \39135 , \39136 , \39137 , \39138 , \39139 , \39140 , \39141 , \39142 , \39143 , \39144 , \39145 , \39146 , \39147 , \39148 , \39149 , \39150 , \39157 );
and \U$33496 ( \39159 , \39124 , \39158 );
buf \U$33497 ( \39160 , \39159 );
or \U$33498 ( \39161 , \39122 , \39160 );
_DC gb026 ( \39162_nGb026 , \39086 , \39161 );
buf \U$33499 ( \39163 , \39162_nGb026 );
xor \U$33500 ( \39164 , \38653 , \39163 );
buf \U$33501 ( \39165 , RIb7b9590_247);
and \U$33502 ( \39166 , \7126 , \38679 );
and \U$33503 ( \39167 , \7128 , \38706 );
and \U$33504 ( \39168 , \8338 , \38733 );
and \U$33505 ( \39169 , \8340 , \38760 );
and \U$33506 ( \39170 , \8342 , \38787 );
and \U$33507 ( \39171 , \8344 , \38814 );
and \U$33508 ( \39172 , \8346 , \38841 );
and \U$33509 ( \39173 , \8348 , \38868 );
and \U$33510 ( \39174 , \8350 , \38895 );
and \U$33511 ( \39175 , \8352 , \38922 );
and \U$33512 ( \39176 , \8354 , \38949 );
and \U$33513 ( \39177 , \8356 , \38976 );
and \U$33514 ( \39178 , \8358 , \39003 );
and \U$33515 ( \39179 , \8360 , \39030 );
and \U$33516 ( \39180 , \8362 , \39057 );
and \U$33517 ( \39181 , \8364 , \39084 );
or \U$33518 ( \39182 , \39166 , \39167 , \39168 , \39169 , \39170 , \39171 , \39172 , \39173 , \39174 , \39175 , \39176 , \39177 , \39178 , \39179 , \39180 , \39181 );
_DC gb03b ( \39183_nGb03b , \39182 , \39161 );
buf \U$33519 ( \39184 , \39183_nGb03b );
xor \U$33520 ( \39185 , \39165 , \39184 );
or \U$33521 ( \39186 , \39164 , \39185 );
buf \U$33522 ( \39187 , RIb7b9518_248);
and \U$33523 ( \39188 , \7136 , \38679 );
and \U$33524 ( \39189 , \7138 , \38706 );
and \U$33525 ( \39190 , \8374 , \38733 );
and \U$33526 ( \39191 , \8376 , \38760 );
and \U$33527 ( \39192 , \8378 , \38787 );
and \U$33528 ( \39193 , \8380 , \38814 );
and \U$33529 ( \39194 , \8382 , \38841 );
and \U$33530 ( \39195 , \8384 , \38868 );
and \U$33531 ( \39196 , \8386 , \38895 );
and \U$33532 ( \39197 , \8388 , \38922 );
and \U$33533 ( \39198 , \8390 , \38949 );
and \U$33534 ( \39199 , \8392 , \38976 );
and \U$33535 ( \39200 , \8394 , \39003 );
and \U$33536 ( \39201 , \8396 , \39030 );
and \U$33537 ( \39202 , \8398 , \39057 );
and \U$33538 ( \39203 , \8400 , \39084 );
or \U$33539 ( \39204 , \39188 , \39189 , \39190 , \39191 , \39192 , \39193 , \39194 , \39195 , \39196 , \39197 , \39198 , \39199 , \39200 , \39201 , \39202 , \39203 );
_DC gb051 ( \39205_nGb051 , \39204 , \39161 );
buf \U$33540 ( \39206 , \39205_nGb051 );
xor \U$33541 ( \39207 , \39187 , \39206 );
or \U$33542 ( \39208 , \39186 , \39207 );
buf \U$33543 ( \39209 , RIb7b94a0_249);
and \U$33544 ( \39210 , \7146 , \38679 );
and \U$33545 ( \39211 , \7148 , \38706 );
and \U$33546 ( \39212 , \8410 , \38733 );
and \U$33547 ( \39213 , \8412 , \38760 );
and \U$33548 ( \39214 , \8414 , \38787 );
and \U$33549 ( \39215 , \8416 , \38814 );
and \U$33550 ( \39216 , \8418 , \38841 );
and \U$33551 ( \39217 , \8420 , \38868 );
and \U$33552 ( \39218 , \8422 , \38895 );
and \U$33553 ( \39219 , \8424 , \38922 );
and \U$33554 ( \39220 , \8426 , \38949 );
and \U$33555 ( \39221 , \8428 , \38976 );
and \U$33556 ( \39222 , \8430 , \39003 );
and \U$33557 ( \39223 , \8432 , \39030 );
and \U$33558 ( \39224 , \8434 , \39057 );
and \U$33559 ( \39225 , \8436 , \39084 );
or \U$33560 ( \39226 , \39210 , \39211 , \39212 , \39213 , \39214 , \39215 , \39216 , \39217 , \39218 , \39219 , \39220 , \39221 , \39222 , \39223 , \39224 , \39225 );
_DC gb067 ( \39227_nGb067 , \39226 , \39161 );
buf \U$33561 ( \39228 , \39227_nGb067 );
xor \U$33562 ( \39229 , \39209 , \39228 );
or \U$33563 ( \39230 , \39208 , \39229 );
buf \U$33564 ( \39231 , RIb7b9428_250);
and \U$33565 ( \39232 , \7156 , \38679 );
and \U$33566 ( \39233 , \7158 , \38706 );
and \U$33567 ( \39234 , \8446 , \38733 );
and \U$33568 ( \39235 , \8448 , \38760 );
and \U$33569 ( \39236 , \8450 , \38787 );
and \U$33570 ( \39237 , \8452 , \38814 );
and \U$33571 ( \39238 , \8454 , \38841 );
and \U$33572 ( \39239 , \8456 , \38868 );
and \U$33573 ( \39240 , \8458 , \38895 );
and \U$33574 ( \39241 , \8460 , \38922 );
and \U$33575 ( \39242 , \8462 , \38949 );
and \U$33576 ( \39243 , \8464 , \38976 );
and \U$33577 ( \39244 , \8466 , \39003 );
and \U$33578 ( \39245 , \8468 , \39030 );
and \U$33579 ( \39246 , \8470 , \39057 );
and \U$33580 ( \39247 , \8472 , \39084 );
or \U$33581 ( \39248 , \39232 , \39233 , \39234 , \39235 , \39236 , \39237 , \39238 , \39239 , \39240 , \39241 , \39242 , \39243 , \39244 , \39245 , \39246 , \39247 );
_DC gb07d ( \39249_nGb07d , \39248 , \39161 );
buf \U$33582 ( \39250 , \39249_nGb07d );
xor \U$33583 ( \39251 , \39231 , \39250 );
or \U$33584 ( \39252 , \39230 , \39251 );
buf \U$33585 ( \39253 , RIb7b93b0_251);
and \U$33586 ( \39254 , \7166 , \38679 );
and \U$33587 ( \39255 , \7168 , \38706 );
and \U$33588 ( \39256 , \8482 , \38733 );
and \U$33589 ( \39257 , \8484 , \38760 );
and \U$33590 ( \39258 , \8486 , \38787 );
and \U$33591 ( \39259 , \8488 , \38814 );
and \U$33592 ( \39260 , \8490 , \38841 );
and \U$33593 ( \39261 , \8492 , \38868 );
and \U$33594 ( \39262 , \8494 , \38895 );
and \U$33595 ( \39263 , \8496 , \38922 );
and \U$33596 ( \39264 , \8498 , \38949 );
and \U$33597 ( \39265 , \8500 , \38976 );
and \U$33598 ( \39266 , \8502 , \39003 );
and \U$33599 ( \39267 , \8504 , \39030 );
and \U$33600 ( \39268 , \8506 , \39057 );
and \U$33601 ( \39269 , \8508 , \39084 );
or \U$33602 ( \39270 , \39254 , \39255 , \39256 , \39257 , \39258 , \39259 , \39260 , \39261 , \39262 , \39263 , \39264 , \39265 , \39266 , \39267 , \39268 , \39269 );
_DC gb093 ( \39271_nGb093 , \39270 , \39161 );
buf \U$33603 ( \39272 , \39271_nGb093 );
xor \U$33604 ( \39273 , \39253 , \39272 );
or \U$33605 ( \39274 , \39252 , \39273 );
buf \U$33606 ( \39275 , RIb7af720_252);
and \U$33607 ( \39276 , \7176 , \38679 );
and \U$33608 ( \39277 , \7178 , \38706 );
and \U$33609 ( \39278 , \8518 , \38733 );
and \U$33610 ( \39279 , \8520 , \38760 );
and \U$33611 ( \39280 , \8522 , \38787 );
and \U$33612 ( \39281 , \8524 , \38814 );
and \U$33613 ( \39282 , \8526 , \38841 );
and \U$33614 ( \39283 , \8528 , \38868 );
and \U$33615 ( \39284 , \8530 , \38895 );
and \U$33616 ( \39285 , \8532 , \38922 );
and \U$33617 ( \39286 , \8534 , \38949 );
and \U$33618 ( \39287 , \8536 , \38976 );
and \U$33619 ( \39288 , \8538 , \39003 );
and \U$33620 ( \39289 , \8540 , \39030 );
and \U$33621 ( \39290 , \8542 , \39057 );
and \U$33622 ( \39291 , \8544 , \39084 );
or \U$33623 ( \39292 , \39276 , \39277 , \39278 , \39279 , \39280 , \39281 , \39282 , \39283 , \39284 , \39285 , \39286 , \39287 , \39288 , \39289 , \39290 , \39291 );
_DC gb0a9 ( \39293_nGb0a9 , \39292 , \39161 );
buf \U$33624 ( \39294 , \39293_nGb0a9 );
xor \U$33625 ( \39295 , \39275 , \39294 );
or \U$33626 ( \39296 , \39274 , \39295 );
buf \U$33627 ( \39297 , RIb7af6a8_253);
and \U$33628 ( \39298 , \7186 , \38679 );
and \U$33629 ( \39299 , \7188 , \38706 );
and \U$33630 ( \39300 , \8554 , \38733 );
and \U$33631 ( \39301 , \8556 , \38760 );
and \U$33632 ( \39302 , \8558 , \38787 );
and \U$33633 ( \39303 , \8560 , \38814 );
and \U$33634 ( \39304 , \8562 , \38841 );
and \U$33635 ( \39305 , \8564 , \38868 );
and \U$33636 ( \39306 , \8566 , \38895 );
and \U$33637 ( \39307 , \8568 , \38922 );
and \U$33638 ( \39308 , \8570 , \38949 );
and \U$33639 ( \39309 , \8572 , \38976 );
and \U$33640 ( \39310 , \8574 , \39003 );
and \U$33641 ( \39311 , \8576 , \39030 );
and \U$33642 ( \39312 , \8578 , \39057 );
and \U$33643 ( \39313 , \8580 , \39084 );
or \U$33644 ( \39314 , \39298 , \39299 , \39300 , \39301 , \39302 , \39303 , \39304 , \39305 , \39306 , \39307 , \39308 , \39309 , \39310 , \39311 , \39312 , \39313 );
_DC gb0bf ( \39315_nGb0bf , \39314 , \39161 );
buf \U$33645 ( \39316 , \39315_nGb0bf );
xor \U$33646 ( \39317 , \39297 , \39316 );
or \U$33647 ( \39318 , \39296 , \39317 );
not \U$33648 ( \39319 , \39318 );
buf \U$33649 ( \39320 , \39319 );
and \U$33650 ( \39321 , \38652 , \39320 );
buf \U$33651 ( \39322 , RIb7af630_254);
buf \U$33652 ( \39323 , \38138 );
buf \U$33653 ( \39324 , \38138 );
buf \U$33654 ( \39325 , \38138 );
buf \U$33655 ( \39326 , \38138 );
buf \U$33656 ( \39327 , \38138 );
buf \U$33657 ( \39328 , \38138 );
buf \U$33658 ( \39329 , \38138 );
buf \U$33659 ( \39330 , \38138 );
buf \U$33660 ( \39331 , \38138 );
buf \U$33661 ( \39332 , \38138 );
buf \U$33662 ( \39333 , \38138 );
buf \U$33663 ( \39334 , \38138 );
buf \U$33664 ( \39335 , \38138 );
buf \U$33665 ( \39336 , \38138 );
buf \U$33666 ( \39337 , \38138 );
buf \U$33667 ( \39338 , \38138 );
buf \U$33668 ( \39339 , \38138 );
buf \U$33669 ( \39340 , \38138 );
buf \U$33670 ( \39341 , \38138 );
buf \U$33671 ( \39342 , \38138 );
buf \U$33672 ( \39343 , \38138 );
buf \U$33673 ( \39344 , \38138 );
buf \U$33674 ( \39345 , \38138 );
buf \U$33675 ( \39346 , \38138 );
buf \U$33676 ( \39347 , \38138 );
nor \U$33677 ( \39348 , \38125 , \38126 , \38127 , \38128 , \38132 , \38135 , \38138 , \39323 , \39324 , \39325 , \39326 , \39327 , \39328 , \39329 , \39330 , \39331 , \39332 , \39333 , \39334 , \39335 , \39336 , \39337 , \39338 , \39339 , \39340 , \39341 , \39342 , \39343 , \39344 , \39345 , \39346 , \39347 );
and \U$33678 ( \39349 , \7198 , \39348 );
buf \U$33679 ( \39350 , \38138 );
buf \U$33680 ( \39351 , \38138 );
buf \U$33681 ( \39352 , \38138 );
buf \U$33682 ( \39353 , \38138 );
buf \U$33683 ( \39354 , \38138 );
buf \U$33684 ( \39355 , \38138 );
buf \U$33685 ( \39356 , \38138 );
buf \U$33686 ( \39357 , \38138 );
buf \U$33687 ( \39358 , \38138 );
buf \U$33688 ( \39359 , \38138 );
buf \U$33689 ( \39360 , \38138 );
buf \U$33690 ( \39361 , \38138 );
buf \U$33691 ( \39362 , \38138 );
buf \U$33692 ( \39363 , \38138 );
buf \U$33693 ( \39364 , \38138 );
buf \U$33694 ( \39365 , \38138 );
buf \U$33695 ( \39366 , \38138 );
buf \U$33696 ( \39367 , \38138 );
buf \U$33697 ( \39368 , \38138 );
buf \U$33698 ( \39369 , \38138 );
buf \U$33699 ( \39370 , \38138 );
buf \U$33700 ( \39371 , \38138 );
buf \U$33701 ( \39372 , \38138 );
buf \U$33702 ( \39373 , \38138 );
buf \U$33703 ( \39374 , \38138 );
nor \U$33704 ( \39375 , \38166 , \38167 , \38168 , \38169 , \38131 , \38135 , \38138 , \39350 , \39351 , \39352 , \39353 , \39354 , \39355 , \39356 , \39357 , \39358 , \39359 , \39360 , \39361 , \39362 , \39363 , \39364 , \39365 , \39366 , \39367 , \39368 , \39369 , \39370 , \39371 , \39372 , \39373 , \39374 );
and \U$33705 ( \39376 , \7200 , \39375 );
buf \U$33706 ( \39377 , \38138 );
buf \U$33707 ( \39378 , \38138 );
buf \U$33708 ( \39379 , \38138 );
buf \U$33709 ( \39380 , \38138 );
buf \U$33710 ( \39381 , \38138 );
buf \U$33711 ( \39382 , \38138 );
buf \U$33712 ( \39383 , \38138 );
buf \U$33713 ( \39384 , \38138 );
buf \U$33714 ( \39385 , \38138 );
buf \U$33715 ( \39386 , \38138 );
buf \U$33716 ( \39387 , \38138 );
buf \U$33717 ( \39388 , \38138 );
buf \U$33718 ( \39389 , \38138 );
buf \U$33719 ( \39390 , \38138 );
buf \U$33720 ( \39391 , \38138 );
buf \U$33721 ( \39392 , \38138 );
buf \U$33722 ( \39393 , \38138 );
buf \U$33723 ( \39394 , \38138 );
buf \U$33724 ( \39395 , \38138 );
buf \U$33725 ( \39396 , \38138 );
buf \U$33726 ( \39397 , \38138 );
buf \U$33727 ( \39398 , \38138 );
buf \U$33728 ( \39399 , \38138 );
buf \U$33729 ( \39400 , \38138 );
buf \U$33730 ( \39401 , \38138 );
nor \U$33731 ( \39402 , \38125 , \38167 , \38168 , \38169 , \38131 , \38135 , \38138 , \39377 , \39378 , \39379 , \39380 , \39381 , \39382 , \39383 , \39384 , \39385 , \39386 , \39387 , \39388 , \39389 , \39390 , \39391 , \39392 , \39393 , \39394 , \39395 , \39396 , \39397 , \39398 , \39399 , \39400 , \39401 );
and \U$33732 ( \39403 , \8645 , \39402 );
buf \U$33733 ( \39404 , \38138 );
buf \U$33734 ( \39405 , \38138 );
buf \U$33735 ( \39406 , \38138 );
buf \U$33736 ( \39407 , \38138 );
buf \U$33737 ( \39408 , \38138 );
buf \U$33738 ( \39409 , \38138 );
buf \U$33739 ( \39410 , \38138 );
buf \U$33740 ( \39411 , \38138 );
buf \U$33741 ( \39412 , \38138 );
buf \U$33742 ( \39413 , \38138 );
buf \U$33743 ( \39414 , \38138 );
buf \U$33744 ( \39415 , \38138 );
buf \U$33745 ( \39416 , \38138 );
buf \U$33746 ( \39417 , \38138 );
buf \U$33747 ( \39418 , \38138 );
buf \U$33748 ( \39419 , \38138 );
buf \U$33749 ( \39420 , \38138 );
buf \U$33750 ( \39421 , \38138 );
buf \U$33751 ( \39422 , \38138 );
buf \U$33752 ( \39423 , \38138 );
buf \U$33753 ( \39424 , \38138 );
buf \U$33754 ( \39425 , \38138 );
buf \U$33755 ( \39426 , \38138 );
buf \U$33756 ( \39427 , \38138 );
buf \U$33757 ( \39428 , \38138 );
nor \U$33758 ( \39429 , \38166 , \38126 , \38168 , \38169 , \38131 , \38135 , \38138 , \39404 , \39405 , \39406 , \39407 , \39408 , \39409 , \39410 , \39411 , \39412 , \39413 , \39414 , \39415 , \39416 , \39417 , \39418 , \39419 , \39420 , \39421 , \39422 , \39423 , \39424 , \39425 , \39426 , \39427 , \39428 );
and \U$33759 ( \39430 , \8673 , \39429 );
buf \U$33760 ( \39431 , \38138 );
buf \U$33761 ( \39432 , \38138 );
buf \U$33762 ( \39433 , \38138 );
buf \U$33763 ( \39434 , \38138 );
buf \U$33764 ( \39435 , \38138 );
buf \U$33765 ( \39436 , \38138 );
buf \U$33766 ( \39437 , \38138 );
buf \U$33767 ( \39438 , \38138 );
buf \U$33768 ( \39439 , \38138 );
buf \U$33769 ( \39440 , \38138 );
buf \U$33770 ( \39441 , \38138 );
buf \U$33771 ( \39442 , \38138 );
buf \U$33772 ( \39443 , \38138 );
buf \U$33773 ( \39444 , \38138 );
buf \U$33774 ( \39445 , \38138 );
buf \U$33775 ( \39446 , \38138 );
buf \U$33776 ( \39447 , \38138 );
buf \U$33777 ( \39448 , \38138 );
buf \U$33778 ( \39449 , \38138 );
buf \U$33779 ( \39450 , \38138 );
buf \U$33780 ( \39451 , \38138 );
buf \U$33781 ( \39452 , \38138 );
buf \U$33782 ( \39453 , \38138 );
buf \U$33783 ( \39454 , \38138 );
buf \U$33784 ( \39455 , \38138 );
nor \U$33785 ( \39456 , \38125 , \38126 , \38168 , \38169 , \38131 , \38135 , \38138 , \39431 , \39432 , \39433 , \39434 , \39435 , \39436 , \39437 , \39438 , \39439 , \39440 , \39441 , \39442 , \39443 , \39444 , \39445 , \39446 , \39447 , \39448 , \39449 , \39450 , \39451 , \39452 , \39453 , \39454 , \39455 );
and \U$33786 ( \39457 , \8701 , \39456 );
buf \U$33787 ( \39458 , \38138 );
buf \U$33788 ( \39459 , \38138 );
buf \U$33789 ( \39460 , \38138 );
buf \U$33790 ( \39461 , \38138 );
buf \U$33791 ( \39462 , \38138 );
buf \U$33792 ( \39463 , \38138 );
buf \U$33793 ( \39464 , \38138 );
buf \U$33794 ( \39465 , \38138 );
buf \U$33795 ( \39466 , \38138 );
buf \U$33796 ( \39467 , \38138 );
buf \U$33797 ( \39468 , \38138 );
buf \U$33798 ( \39469 , \38138 );
buf \U$33799 ( \39470 , \38138 );
buf \U$33800 ( \39471 , \38138 );
buf \U$33801 ( \39472 , \38138 );
buf \U$33802 ( \39473 , \38138 );
buf \U$33803 ( \39474 , \38138 );
buf \U$33804 ( \39475 , \38138 );
buf \U$33805 ( \39476 , \38138 );
buf \U$33806 ( \39477 , \38138 );
buf \U$33807 ( \39478 , \38138 );
buf \U$33808 ( \39479 , \38138 );
buf \U$33809 ( \39480 , \38138 );
buf \U$33810 ( \39481 , \38138 );
buf \U$33811 ( \39482 , \38138 );
nor \U$33812 ( \39483 , \38166 , \38167 , \38127 , \38169 , \38131 , \38135 , \38138 , \39458 , \39459 , \39460 , \39461 , \39462 , \39463 , \39464 , \39465 , \39466 , \39467 , \39468 , \39469 , \39470 , \39471 , \39472 , \39473 , \39474 , \39475 , \39476 , \39477 , \39478 , \39479 , \39480 , \39481 , \39482 );
and \U$33813 ( \39484 , \8729 , \39483 );
buf \U$33814 ( \39485 , \38138 );
buf \U$33815 ( \39486 , \38138 );
buf \U$33816 ( \39487 , \38138 );
buf \U$33817 ( \39488 , \38138 );
buf \U$33818 ( \39489 , \38138 );
buf \U$33819 ( \39490 , \38138 );
buf \U$33820 ( \39491 , \38138 );
buf \U$33821 ( \39492 , \38138 );
buf \U$33822 ( \39493 , \38138 );
buf \U$33823 ( \39494 , \38138 );
buf \U$33824 ( \39495 , \38138 );
buf \U$33825 ( \39496 , \38138 );
buf \U$33826 ( \39497 , \38138 );
buf \U$33827 ( \39498 , \38138 );
buf \U$33828 ( \39499 , \38138 );
buf \U$33829 ( \39500 , \38138 );
buf \U$33830 ( \39501 , \38138 );
buf \U$33831 ( \39502 , \38138 );
buf \U$33832 ( \39503 , \38138 );
buf \U$33833 ( \39504 , \38138 );
buf \U$33834 ( \39505 , \38138 );
buf \U$33835 ( \39506 , \38138 );
buf \U$33836 ( \39507 , \38138 );
buf \U$33837 ( \39508 , \38138 );
buf \U$33838 ( \39509 , \38138 );
nor \U$33839 ( \39510 , \38125 , \38167 , \38127 , \38169 , \38131 , \38135 , \38138 , \39485 , \39486 , \39487 , \39488 , \39489 , \39490 , \39491 , \39492 , \39493 , \39494 , \39495 , \39496 , \39497 , \39498 , \39499 , \39500 , \39501 , \39502 , \39503 , \39504 , \39505 , \39506 , \39507 , \39508 , \39509 );
and \U$33840 ( \39511 , \8757 , \39510 );
buf \U$33841 ( \39512 , \38138 );
buf \U$33842 ( \39513 , \38138 );
buf \U$33843 ( \39514 , \38138 );
buf \U$33844 ( \39515 , \38138 );
buf \U$33845 ( \39516 , \38138 );
buf \U$33846 ( \39517 , \38138 );
buf \U$33847 ( \39518 , \38138 );
buf \U$33848 ( \39519 , \38138 );
buf \U$33849 ( \39520 , \38138 );
buf \U$33850 ( \39521 , \38138 );
buf \U$33851 ( \39522 , \38138 );
buf \U$33852 ( \39523 , \38138 );
buf \U$33853 ( \39524 , \38138 );
buf \U$33854 ( \39525 , \38138 );
buf \U$33855 ( \39526 , \38138 );
buf \U$33856 ( \39527 , \38138 );
buf \U$33857 ( \39528 , \38138 );
buf \U$33858 ( \39529 , \38138 );
buf \U$33859 ( \39530 , \38138 );
buf \U$33860 ( \39531 , \38138 );
buf \U$33861 ( \39532 , \38138 );
buf \U$33862 ( \39533 , \38138 );
buf \U$33863 ( \39534 , \38138 );
buf \U$33864 ( \39535 , \38138 );
buf \U$33865 ( \39536 , \38138 );
nor \U$33866 ( \39537 , \38166 , \38126 , \38127 , \38169 , \38131 , \38135 , \38138 , \39512 , \39513 , \39514 , \39515 , \39516 , \39517 , \39518 , \39519 , \39520 , \39521 , \39522 , \39523 , \39524 , \39525 , \39526 , \39527 , \39528 , \39529 , \39530 , \39531 , \39532 , \39533 , \39534 , \39535 , \39536 );
and \U$33867 ( \39538 , \8785 , \39537 );
buf \U$33868 ( \39539 , \38138 );
buf \U$33869 ( \39540 , \38138 );
buf \U$33870 ( \39541 , \38138 );
buf \U$33871 ( \39542 , \38138 );
buf \U$33872 ( \39543 , \38138 );
buf \U$33873 ( \39544 , \38138 );
buf \U$33874 ( \39545 , \38138 );
buf \U$33875 ( \39546 , \38138 );
buf \U$33876 ( \39547 , \38138 );
buf \U$33877 ( \39548 , \38138 );
buf \U$33878 ( \39549 , \38138 );
buf \U$33879 ( \39550 , \38138 );
buf \U$33880 ( \39551 , \38138 );
buf \U$33881 ( \39552 , \38138 );
buf \U$33882 ( \39553 , \38138 );
buf \U$33883 ( \39554 , \38138 );
buf \U$33884 ( \39555 , \38138 );
buf \U$33885 ( \39556 , \38138 );
buf \U$33886 ( \39557 , \38138 );
buf \U$33887 ( \39558 , \38138 );
buf \U$33888 ( \39559 , \38138 );
buf \U$33889 ( \39560 , \38138 );
buf \U$33890 ( \39561 , \38138 );
buf \U$33891 ( \39562 , \38138 );
buf \U$33892 ( \39563 , \38138 );
nor \U$33893 ( \39564 , \38125 , \38126 , \38127 , \38169 , \38131 , \38135 , \38138 , \39539 , \39540 , \39541 , \39542 , \39543 , \39544 , \39545 , \39546 , \39547 , \39548 , \39549 , \39550 , \39551 , \39552 , \39553 , \39554 , \39555 , \39556 , \39557 , \39558 , \39559 , \39560 , \39561 , \39562 , \39563 );
and \U$33894 ( \39565 , \8813 , \39564 );
buf \U$33895 ( \39566 , \38138 );
buf \U$33896 ( \39567 , \38138 );
buf \U$33897 ( \39568 , \38138 );
buf \U$33898 ( \39569 , \38138 );
buf \U$33899 ( \39570 , \38138 );
buf \U$33900 ( \39571 , \38138 );
buf \U$33901 ( \39572 , \38138 );
buf \U$33902 ( \39573 , \38138 );
buf \U$33903 ( \39574 , \38138 );
buf \U$33904 ( \39575 , \38138 );
buf \U$33905 ( \39576 , \38138 );
buf \U$33906 ( \39577 , \38138 );
buf \U$33907 ( \39578 , \38138 );
buf \U$33908 ( \39579 , \38138 );
buf \U$33909 ( \39580 , \38138 );
buf \U$33910 ( \39581 , \38138 );
buf \U$33911 ( \39582 , \38138 );
buf \U$33912 ( \39583 , \38138 );
buf \U$33913 ( \39584 , \38138 );
buf \U$33914 ( \39585 , \38138 );
buf \U$33915 ( \39586 , \38138 );
buf \U$33916 ( \39587 , \38138 );
buf \U$33917 ( \39588 , \38138 );
buf \U$33918 ( \39589 , \38138 );
buf \U$33919 ( \39590 , \38138 );
nor \U$33920 ( \39591 , \38166 , \38167 , \38168 , \38128 , \38131 , \38135 , \38138 , \39566 , \39567 , \39568 , \39569 , \39570 , \39571 , \39572 , \39573 , \39574 , \39575 , \39576 , \39577 , \39578 , \39579 , \39580 , \39581 , \39582 , \39583 , \39584 , \39585 , \39586 , \39587 , \39588 , \39589 , \39590 );
and \U$33921 ( \39592 , \8841 , \39591 );
buf \U$33922 ( \39593 , \38138 );
buf \U$33923 ( \39594 , \38138 );
buf \U$33924 ( \39595 , \38138 );
buf \U$33925 ( \39596 , \38138 );
buf \U$33926 ( \39597 , \38138 );
buf \U$33927 ( \39598 , \38138 );
buf \U$33928 ( \39599 , \38138 );
buf \U$33929 ( \39600 , \38138 );
buf \U$33930 ( \39601 , \38138 );
buf \U$33931 ( \39602 , \38138 );
buf \U$33932 ( \39603 , \38138 );
buf \U$33933 ( \39604 , \38138 );
buf \U$33934 ( \39605 , \38138 );
buf \U$33935 ( \39606 , \38138 );
buf \U$33936 ( \39607 , \38138 );
buf \U$33937 ( \39608 , \38138 );
buf \U$33938 ( \39609 , \38138 );
buf \U$33939 ( \39610 , \38138 );
buf \U$33940 ( \39611 , \38138 );
buf \U$33941 ( \39612 , \38138 );
buf \U$33942 ( \39613 , \38138 );
buf \U$33943 ( \39614 , \38138 );
buf \U$33944 ( \39615 , \38138 );
buf \U$33945 ( \39616 , \38138 );
buf \U$33946 ( \39617 , \38138 );
nor \U$33947 ( \39618 , \38125 , \38167 , \38168 , \38128 , \38131 , \38135 , \38138 , \39593 , \39594 , \39595 , \39596 , \39597 , \39598 , \39599 , \39600 , \39601 , \39602 , \39603 , \39604 , \39605 , \39606 , \39607 , \39608 , \39609 , \39610 , \39611 , \39612 , \39613 , \39614 , \39615 , \39616 , \39617 );
and \U$33948 ( \39619 , \8869 , \39618 );
buf \U$33949 ( \39620 , \38138 );
buf \U$33950 ( \39621 , \38138 );
buf \U$33951 ( \39622 , \38138 );
buf \U$33952 ( \39623 , \38138 );
buf \U$33953 ( \39624 , \38138 );
buf \U$33954 ( \39625 , \38138 );
buf \U$33955 ( \39626 , \38138 );
buf \U$33956 ( \39627 , \38138 );
buf \U$33957 ( \39628 , \38138 );
buf \U$33958 ( \39629 , \38138 );
buf \U$33959 ( \39630 , \38138 );
buf \U$33960 ( \39631 , \38138 );
buf \U$33961 ( \39632 , \38138 );
buf \U$33962 ( \39633 , \38138 );
buf \U$33963 ( \39634 , \38138 );
buf \U$33964 ( \39635 , \38138 );
buf \U$33965 ( \39636 , \38138 );
buf \U$33966 ( \39637 , \38138 );
buf \U$33967 ( \39638 , \38138 );
buf \U$33968 ( \39639 , \38138 );
buf \U$33969 ( \39640 , \38138 );
buf \U$33970 ( \39641 , \38138 );
buf \U$33971 ( \39642 , \38138 );
buf \U$33972 ( \39643 , \38138 );
buf \U$33973 ( \39644 , \38138 );
nor \U$33974 ( \39645 , \38166 , \38126 , \38168 , \38128 , \38131 , \38135 , \38138 , \39620 , \39621 , \39622 , \39623 , \39624 , \39625 , \39626 , \39627 , \39628 , \39629 , \39630 , \39631 , \39632 , \39633 , \39634 , \39635 , \39636 , \39637 , \39638 , \39639 , \39640 , \39641 , \39642 , \39643 , \39644 );
and \U$33975 ( \39646 , \8897 , \39645 );
buf \U$33976 ( \39647 , \38138 );
buf \U$33977 ( \39648 , \38138 );
buf \U$33978 ( \39649 , \38138 );
buf \U$33979 ( \39650 , \38138 );
buf \U$33980 ( \39651 , \38138 );
buf \U$33981 ( \39652 , \38138 );
buf \U$33982 ( \39653 , \38138 );
buf \U$33983 ( \39654 , \38138 );
buf \U$33984 ( \39655 , \38138 );
buf \U$33985 ( \39656 , \38138 );
buf \U$33986 ( \39657 , \38138 );
buf \U$33987 ( \39658 , \38138 );
buf \U$33988 ( \39659 , \38138 );
buf \U$33989 ( \39660 , \38138 );
buf \U$33990 ( \39661 , \38138 );
buf \U$33991 ( \39662 , \38138 );
buf \U$33992 ( \39663 , \38138 );
buf \U$33993 ( \39664 , \38138 );
buf \U$33994 ( \39665 , \38138 );
buf \U$33995 ( \39666 , \38138 );
buf \U$33996 ( \39667 , \38138 );
buf \U$33997 ( \39668 , \38138 );
buf \U$33998 ( \39669 , \38138 );
buf \U$33999 ( \39670 , \38138 );
buf \U$34000 ( \39671 , \38138 );
nor \U$34001 ( \39672 , \38125 , \38126 , \38168 , \38128 , \38131 , \38135 , \38138 , \39647 , \39648 , \39649 , \39650 , \39651 , \39652 , \39653 , \39654 , \39655 , \39656 , \39657 , \39658 , \39659 , \39660 , \39661 , \39662 , \39663 , \39664 , \39665 , \39666 , \39667 , \39668 , \39669 , \39670 , \39671 );
and \U$34002 ( \39673 , \8925 , \39672 );
buf \U$34003 ( \39674 , \38138 );
buf \U$34004 ( \39675 , \38138 );
buf \U$34005 ( \39676 , \38138 );
buf \U$34006 ( \39677 , \38138 );
buf \U$34007 ( \39678 , \38138 );
buf \U$34008 ( \39679 , \38138 );
buf \U$34009 ( \39680 , \38138 );
buf \U$34010 ( \39681 , \38138 );
buf \U$34011 ( \39682 , \38138 );
buf \U$34012 ( \39683 , \38138 );
buf \U$34013 ( \39684 , \38138 );
buf \U$34014 ( \39685 , \38138 );
buf \U$34015 ( \39686 , \38138 );
buf \U$34016 ( \39687 , \38138 );
buf \U$34017 ( \39688 , \38138 );
buf \U$34018 ( \39689 , \38138 );
buf \U$34019 ( \39690 , \38138 );
buf \U$34020 ( \39691 , \38138 );
buf \U$34021 ( \39692 , \38138 );
buf \U$34022 ( \39693 , \38138 );
buf \U$34023 ( \39694 , \38138 );
buf \U$34024 ( \39695 , \38138 );
buf \U$34025 ( \39696 , \38138 );
buf \U$34026 ( \39697 , \38138 );
buf \U$34027 ( \39698 , \38138 );
nor \U$34028 ( \39699 , \38166 , \38167 , \38127 , \38128 , \38131 , \38135 , \38138 , \39674 , \39675 , \39676 , \39677 , \39678 , \39679 , \39680 , \39681 , \39682 , \39683 , \39684 , \39685 , \39686 , \39687 , \39688 , \39689 , \39690 , \39691 , \39692 , \39693 , \39694 , \39695 , \39696 , \39697 , \39698 );
and \U$34029 ( \39700 , \8953 , \39699 );
buf \U$34030 ( \39701 , \38138 );
buf \U$34031 ( \39702 , \38138 );
buf \U$34032 ( \39703 , \38138 );
buf \U$34033 ( \39704 , \38138 );
buf \U$34034 ( \39705 , \38138 );
buf \U$34035 ( \39706 , \38138 );
buf \U$34036 ( \39707 , \38138 );
buf \U$34037 ( \39708 , \38138 );
buf \U$34038 ( \39709 , \38138 );
buf \U$34039 ( \39710 , \38138 );
buf \U$34040 ( \39711 , \38138 );
buf \U$34041 ( \39712 , \38138 );
buf \U$34042 ( \39713 , \38138 );
buf \U$34043 ( \39714 , \38138 );
buf \U$34044 ( \39715 , \38138 );
buf \U$34045 ( \39716 , \38138 );
buf \U$34046 ( \39717 , \38138 );
buf \U$34047 ( \39718 , \38138 );
buf \U$34048 ( \39719 , \38138 );
buf \U$34049 ( \39720 , \38138 );
buf \U$34050 ( \39721 , \38138 );
buf \U$34051 ( \39722 , \38138 );
buf \U$34052 ( \39723 , \38138 );
buf \U$34053 ( \39724 , \38138 );
buf \U$34054 ( \39725 , \38138 );
nor \U$34055 ( \39726 , \38125 , \38167 , \38127 , \38128 , \38131 , \38135 , \38138 , \39701 , \39702 , \39703 , \39704 , \39705 , \39706 , \39707 , \39708 , \39709 , \39710 , \39711 , \39712 , \39713 , \39714 , \39715 , \39716 , \39717 , \39718 , \39719 , \39720 , \39721 , \39722 , \39723 , \39724 , \39725 );
and \U$34056 ( \39727 , \8981 , \39726 );
buf \U$34057 ( \39728 , \38138 );
buf \U$34058 ( \39729 , \38138 );
buf \U$34059 ( \39730 , \38138 );
buf \U$34060 ( \39731 , \38138 );
buf \U$34061 ( \39732 , \38138 );
buf \U$34062 ( \39733 , \38138 );
buf \U$34063 ( \39734 , \38138 );
buf \U$34064 ( \39735 , \38138 );
buf \U$34065 ( \39736 , \38138 );
buf \U$34066 ( \39737 , \38138 );
buf \U$34067 ( \39738 , \38138 );
buf \U$34068 ( \39739 , \38138 );
buf \U$34069 ( \39740 , \38138 );
buf \U$34070 ( \39741 , \38138 );
buf \U$34071 ( \39742 , \38138 );
buf \U$34072 ( \39743 , \38138 );
buf \U$34073 ( \39744 , \38138 );
buf \U$34074 ( \39745 , \38138 );
buf \U$34075 ( \39746 , \38138 );
buf \U$34076 ( \39747 , \38138 );
buf \U$34077 ( \39748 , \38138 );
buf \U$34078 ( \39749 , \38138 );
buf \U$34079 ( \39750 , \38138 );
buf \U$34080 ( \39751 , \38138 );
buf \U$34081 ( \39752 , \38138 );
nor \U$34082 ( \39753 , \38166 , \38126 , \38127 , \38128 , \38131 , \38135 , \38138 , \39728 , \39729 , \39730 , \39731 , \39732 , \39733 , \39734 , \39735 , \39736 , \39737 , \39738 , \39739 , \39740 , \39741 , \39742 , \39743 , \39744 , \39745 , \39746 , \39747 , \39748 , \39749 , \39750 , \39751 , \39752 );
and \U$34083 ( \39754 , \9009 , \39753 );
or \U$34084 ( \39755 , \39349 , \39376 , \39403 , \39430 , \39457 , \39484 , \39511 , \39538 , \39565 , \39592 , \39619 , \39646 , \39673 , \39700 , \39727 , \39754 );
buf \U$34085 ( \39756 , \38138 );
not \U$34086 ( \39757 , \39756 );
buf \U$34087 ( \39758 , \38126 );
buf \U$34088 ( \39759 , \38127 );
buf \U$34089 ( \39760 , \38128 );
buf \U$34090 ( \39761 , \38131 );
buf \U$34091 ( \39762 , \38135 );
buf \U$34092 ( \39763 , \38138 );
buf \U$34093 ( \39764 , \38138 );
buf \U$34094 ( \39765 , \38138 );
buf \U$34095 ( \39766 , \38138 );
buf \U$34096 ( \39767 , \38138 );
buf \U$34097 ( \39768 , \38138 );
buf \U$34098 ( \39769 , \38138 );
buf \U$34099 ( \39770 , \38138 );
buf \U$34100 ( \39771 , \38138 );
buf \U$34101 ( \39772 , \38138 );
buf \U$34102 ( \39773 , \38138 );
buf \U$34103 ( \39774 , \38138 );
buf \U$34104 ( \39775 , \38138 );
buf \U$34105 ( \39776 , \38138 );
buf \U$34106 ( \39777 , \38138 );
buf \U$34107 ( \39778 , \38138 );
buf \U$34108 ( \39779 , \38138 );
buf \U$34109 ( \39780 , \38138 );
buf \U$34110 ( \39781 , \38138 );
buf \U$34111 ( \39782 , \38138 );
buf \U$34112 ( \39783 , \38138 );
buf \U$34113 ( \39784 , \38138 );
buf \U$34114 ( \39785 , \38138 );
buf \U$34115 ( \39786 , \38138 );
buf \U$34116 ( \39787 , \38138 );
buf \U$34117 ( \39788 , \38125 );
or \U$34118 ( \39789 , \39758 , \39759 , \39760 , \39761 , \39762 , \39763 , \39764 , \39765 , \39766 , \39767 , \39768 , \39769 , \39770 , \39771 , \39772 , \39773 , \39774 , \39775 , \39776 , \39777 , \39778 , \39779 , \39780 , \39781 , \39782 , \39783 , \39784 , \39785 , \39786 , \39787 , \39788 );
nand \U$34119 ( \39790 , \39757 , \39789 );
buf \U$34120 ( \39791 , \39790 );
buf \U$34121 ( \39792 , \38138 );
not \U$34122 ( \39793 , \39792 );
buf \U$34123 ( \39794 , \38135 );
buf \U$34124 ( \39795 , \38138 );
buf \U$34125 ( \39796 , \38138 );
buf \U$34126 ( \39797 , \38138 );
buf \U$34127 ( \39798 , \38138 );
buf \U$34128 ( \39799 , \38138 );
buf \U$34129 ( \39800 , \38138 );
buf \U$34130 ( \39801 , \38138 );
buf \U$34131 ( \39802 , \38138 );
buf \U$34132 ( \39803 , \38138 );
buf \U$34133 ( \39804 , \38138 );
buf \U$34134 ( \39805 , \38138 );
buf \U$34135 ( \39806 , \38138 );
buf \U$34136 ( \39807 , \38138 );
buf \U$34137 ( \39808 , \38138 );
buf \U$34138 ( \39809 , \38138 );
buf \U$34139 ( \39810 , \38138 );
buf \U$34140 ( \39811 , \38138 );
buf \U$34141 ( \39812 , \38138 );
buf \U$34142 ( \39813 , \38138 );
buf \U$34143 ( \39814 , \38138 );
buf \U$34144 ( \39815 , \38138 );
buf \U$34145 ( \39816 , \38138 );
buf \U$34146 ( \39817 , \38138 );
buf \U$34147 ( \39818 , \38138 );
buf \U$34148 ( \39819 , \38138 );
buf \U$34149 ( \39820 , \38131 );
buf \U$34150 ( \39821 , \38125 );
buf \U$34151 ( \39822 , \38126 );
buf \U$34152 ( \39823 , \38127 );
buf \U$34153 ( \39824 , \38128 );
or \U$34154 ( \39825 , \39821 , \39822 , \39823 , \39824 );
and \U$34155 ( \39826 , \39820 , \39825 );
or \U$34156 ( \39827 , \39794 , \39795 , \39796 , \39797 , \39798 , \39799 , \39800 , \39801 , \39802 , \39803 , \39804 , \39805 , \39806 , \39807 , \39808 , \39809 , \39810 , \39811 , \39812 , \39813 , \39814 , \39815 , \39816 , \39817 , \39818 , \39819 , \39826 );
and \U$34157 ( \39828 , \39793 , \39827 );
buf \U$34158 ( \39829 , \39828 );
or \U$34159 ( \39830 , \39791 , \39829 );
_DC gb2c3 ( \39831_nGb2c3 , \39755 , \39830 );
buf \U$34160 ( \39832 , \39831_nGb2c3 );
xor \U$34161 ( \39833 , \39322 , \39832 );
buf \U$34162 ( \39834 , RIb7af5b8_255);
and \U$34163 ( \39835 , \7207 , \39348 );
and \U$34164 ( \39836 , \7209 , \39375 );
and \U$34165 ( \39837 , \9119 , \39402 );
and \U$34166 ( \39838 , \9121 , \39429 );
and \U$34167 ( \39839 , \9123 , \39456 );
and \U$34168 ( \39840 , \9125 , \39483 );
and \U$34169 ( \39841 , \9127 , \39510 );
and \U$34170 ( \39842 , \9129 , \39537 );
and \U$34171 ( \39843 , \9131 , \39564 );
and \U$34172 ( \39844 , \9133 , \39591 );
and \U$34173 ( \39845 , \9135 , \39618 );
and \U$34174 ( \39846 , \9137 , \39645 );
and \U$34175 ( \39847 , \9139 , \39672 );
and \U$34176 ( \39848 , \9141 , \39699 );
and \U$34177 ( \39849 , \9143 , \39726 );
and \U$34178 ( \39850 , \9145 , \39753 );
or \U$34179 ( \39851 , \39835 , \39836 , \39837 , \39838 , \39839 , \39840 , \39841 , \39842 , \39843 , \39844 , \39845 , \39846 , \39847 , \39848 , \39849 , \39850 );
_DC gb2d8 ( \39852_nGb2d8 , \39851 , \39830 );
buf \U$34180 ( \39853 , \39852_nGb2d8 );
xor \U$34181 ( \39854 , \39834 , \39853 );
or \U$34182 ( \39855 , \39833 , \39854 );
buf \U$34183 ( \39856 , RIb7af540_256);
and \U$34184 ( \39857 , \7217 , \39348 );
and \U$34185 ( \39858 , \7219 , \39375 );
and \U$34186 ( \39859 , \9155 , \39402 );
and \U$34187 ( \39860 , \9157 , \39429 );
and \U$34188 ( \39861 , \9159 , \39456 );
and \U$34189 ( \39862 , \9161 , \39483 );
and \U$34190 ( \39863 , \9163 , \39510 );
and \U$34191 ( \39864 , \9165 , \39537 );
and \U$34192 ( \39865 , \9167 , \39564 );
and \U$34193 ( \39866 , \9169 , \39591 );
and \U$34194 ( \39867 , \9171 , \39618 );
and \U$34195 ( \39868 , \9173 , \39645 );
and \U$34196 ( \39869 , \9175 , \39672 );
and \U$34197 ( \39870 , \9177 , \39699 );
and \U$34198 ( \39871 , \9179 , \39726 );
and \U$34199 ( \39872 , \9181 , \39753 );
or \U$34200 ( \39873 , \39857 , \39858 , \39859 , \39860 , \39861 , \39862 , \39863 , \39864 , \39865 , \39866 , \39867 , \39868 , \39869 , \39870 , \39871 , \39872 );
_DC gb2ee ( \39874_nGb2ee , \39873 , \39830 );
buf \U$34201 ( \39875 , \39874_nGb2ee );
xor \U$34202 ( \39876 , \39856 , \39875 );
or \U$34203 ( \39877 , \39855 , \39876 );
buf \U$34204 ( \39878 , RIb7af4c8_257);
and \U$34205 ( \39879 , \7227 , \39348 );
and \U$34206 ( \39880 , \7229 , \39375 );
and \U$34207 ( \39881 , \9191 , \39402 );
and \U$34208 ( \39882 , \9193 , \39429 );
and \U$34209 ( \39883 , \9195 , \39456 );
and \U$34210 ( \39884 , \9197 , \39483 );
and \U$34211 ( \39885 , \9199 , \39510 );
and \U$34212 ( \39886 , \9201 , \39537 );
and \U$34213 ( \39887 , \9203 , \39564 );
and \U$34214 ( \39888 , \9205 , \39591 );
and \U$34215 ( \39889 , \9207 , \39618 );
and \U$34216 ( \39890 , \9209 , \39645 );
and \U$34217 ( \39891 , \9211 , \39672 );
and \U$34218 ( \39892 , \9213 , \39699 );
and \U$34219 ( \39893 , \9215 , \39726 );
and \U$34220 ( \39894 , \9217 , \39753 );
or \U$34221 ( \39895 , \39879 , \39880 , \39881 , \39882 , \39883 , \39884 , \39885 , \39886 , \39887 , \39888 , \39889 , \39890 , \39891 , \39892 , \39893 , \39894 );
_DC gb304 ( \39896_nGb304 , \39895 , \39830 );
buf \U$34222 ( \39897 , \39896_nGb304 );
xor \U$34223 ( \39898 , \39878 , \39897 );
or \U$34224 ( \39899 , \39877 , \39898 );
buf \U$34225 ( \39900 , RIb7af450_258);
and \U$34226 ( \39901 , \7237 , \39348 );
and \U$34227 ( \39902 , \7239 , \39375 );
and \U$34228 ( \39903 , \9227 , \39402 );
and \U$34229 ( \39904 , \9229 , \39429 );
and \U$34230 ( \39905 , \9231 , \39456 );
and \U$34231 ( \39906 , \9233 , \39483 );
and \U$34232 ( \39907 , \9235 , \39510 );
and \U$34233 ( \39908 , \9237 , \39537 );
and \U$34234 ( \39909 , \9239 , \39564 );
and \U$34235 ( \39910 , \9241 , \39591 );
and \U$34236 ( \39911 , \9243 , \39618 );
and \U$34237 ( \39912 , \9245 , \39645 );
and \U$34238 ( \39913 , \9247 , \39672 );
and \U$34239 ( \39914 , \9249 , \39699 );
and \U$34240 ( \39915 , \9251 , \39726 );
and \U$34241 ( \39916 , \9253 , \39753 );
or \U$34242 ( \39917 , \39901 , \39902 , \39903 , \39904 , \39905 , \39906 , \39907 , \39908 , \39909 , \39910 , \39911 , \39912 , \39913 , \39914 , \39915 , \39916 );
_DC gb31a ( \39918_nGb31a , \39917 , \39830 );
buf \U$34243 ( \39919 , \39918_nGb31a );
xor \U$34244 ( \39920 , \39900 , \39919 );
or \U$34245 ( \39921 , \39899 , \39920 );
buf \U$34246 ( \39922 , RIb7af3d8_259);
and \U$34247 ( \39923 , \7247 , \39348 );
and \U$34248 ( \39924 , \7249 , \39375 );
and \U$34249 ( \39925 , \9263 , \39402 );
and \U$34250 ( \39926 , \9265 , \39429 );
and \U$34251 ( \39927 , \9267 , \39456 );
and \U$34252 ( \39928 , \9269 , \39483 );
and \U$34253 ( \39929 , \9271 , \39510 );
and \U$34254 ( \39930 , \9273 , \39537 );
and \U$34255 ( \39931 , \9275 , \39564 );
and \U$34256 ( \39932 , \9277 , \39591 );
and \U$34257 ( \39933 , \9279 , \39618 );
and \U$34258 ( \39934 , \9281 , \39645 );
and \U$34259 ( \39935 , \9283 , \39672 );
and \U$34260 ( \39936 , \9285 , \39699 );
and \U$34261 ( \39937 , \9287 , \39726 );
and \U$34262 ( \39938 , \9289 , \39753 );
or \U$34263 ( \39939 , \39923 , \39924 , \39925 , \39926 , \39927 , \39928 , \39929 , \39930 , \39931 , \39932 , \39933 , \39934 , \39935 , \39936 , \39937 , \39938 );
_DC gb330 ( \39940_nGb330 , \39939 , \39830 );
buf \U$34264 ( \39941 , \39940_nGb330 );
xor \U$34265 ( \39942 , \39922 , \39941 );
or \U$34266 ( \39943 , \39921 , \39942 );
buf \U$34267 ( \39944 , RIb7a5bf8_260);
and \U$34268 ( \39945 , \7257 , \39348 );
and \U$34269 ( \39946 , \7259 , \39375 );
and \U$34270 ( \39947 , \9299 , \39402 );
and \U$34271 ( \39948 , \9301 , \39429 );
and \U$34272 ( \39949 , \9303 , \39456 );
and \U$34273 ( \39950 , \9305 , \39483 );
and \U$34274 ( \39951 , \9307 , \39510 );
and \U$34275 ( \39952 , \9309 , \39537 );
and \U$34276 ( \39953 , \9311 , \39564 );
and \U$34277 ( \39954 , \9313 , \39591 );
and \U$34278 ( \39955 , \9315 , \39618 );
and \U$34279 ( \39956 , \9317 , \39645 );
and \U$34280 ( \39957 , \9319 , \39672 );
and \U$34281 ( \39958 , \9321 , \39699 );
and \U$34282 ( \39959 , \9323 , \39726 );
and \U$34283 ( \39960 , \9325 , \39753 );
or \U$34284 ( \39961 , \39945 , \39946 , \39947 , \39948 , \39949 , \39950 , \39951 , \39952 , \39953 , \39954 , \39955 , \39956 , \39957 , \39958 , \39959 , \39960 );
_DC gb346 ( \39962_nGb346 , \39961 , \39830 );
buf \U$34285 ( \39963 , \39962_nGb346 );
xor \U$34286 ( \39964 , \39944 , \39963 );
or \U$34287 ( \39965 , \39943 , \39964 );
buf \U$34288 ( \39966 , RIb7a0c48_261);
and \U$34289 ( \39967 , \7267 , \39348 );
and \U$34290 ( \39968 , \7269 , \39375 );
and \U$34291 ( \39969 , \9335 , \39402 );
and \U$34292 ( \39970 , \9337 , \39429 );
and \U$34293 ( \39971 , \9339 , \39456 );
and \U$34294 ( \39972 , \9341 , \39483 );
and \U$34295 ( \39973 , \9343 , \39510 );
and \U$34296 ( \39974 , \9345 , \39537 );
and \U$34297 ( \39975 , \9347 , \39564 );
and \U$34298 ( \39976 , \9349 , \39591 );
and \U$34299 ( \39977 , \9351 , \39618 );
and \U$34300 ( \39978 , \9353 , \39645 );
and \U$34301 ( \39979 , \9355 , \39672 );
and \U$34302 ( \39980 , \9357 , \39699 );
and \U$34303 ( \39981 , \9359 , \39726 );
and \U$34304 ( \39982 , \9361 , \39753 );
or \U$34305 ( \39983 , \39967 , \39968 , \39969 , \39970 , \39971 , \39972 , \39973 , \39974 , \39975 , \39976 , \39977 , \39978 , \39979 , \39980 , \39981 , \39982 );
_DC gb35c ( \39984_nGb35c , \39983 , \39830 );
buf \U$34306 ( \39985 , \39984_nGb35c );
xor \U$34307 ( \39986 , \39966 , \39985 );
or \U$34308 ( \39987 , \39965 , \39986 );
not \U$34309 ( \39988 , \39987 );
buf \U$34310 ( \39989 , \39988 );
and \U$34311 ( \39990 , \39321 , \39989 );
_HMUX gb363 ( \39991_nGb363 , \37696_nGaa64 , \38125 , \39990 );
buf \U$34312 ( \39992 , \37717 );
buf \U$34313 ( \39993 , \37714 );
buf \U$34314 ( \39994 , \37699 );
buf \U$34315 ( \39995 , \37702 );
buf \U$34316 ( \39996 , \37706 );
buf \U$34317 ( \39997 , \37710 );
or \U$34318 ( \39998 , \39994 , \39995 , \39996 , \39997 );
and \U$34319 ( \39999 , \39993 , \39998 );
or \U$34320 ( \40000 , \39992 , \39999 );
buf \U$34321 ( \40001 , \40000 );
_HMUX gb36e ( \40002_nGb36e , \38124_nGac10 , \39991_nGb363 , \40001 );
nor \U$34322 ( \40003 , RIe5319e0_6884, RIe549ef0_6842, RIe549770_6843, RIe548ff0_6844, \7063 );
and \U$34323 ( \40004 , RIe5329d0_6883, \40003 );
and \U$34324 ( \40005 , RIe5319e0_6884, RIe549ef0_6842, RIe549770_6843, RIe548ff0_6844, \7063 );
and \U$34325 ( \40006 , RIeb72150_6905, \40005 );
not \U$34326 ( \40007 , RIe5319e0_6884);
and \U$34327 ( \40008 , \40007 , RIe549ef0_6842, RIe549770_6843, RIe548ff0_6844, \7063 );
and \U$34328 ( \40009 , RIeab80c0_6897, \40008 );
and \U$34329 ( \40010 , RIe5319e0_6884, \7061 , RIe549770_6843, RIe548ff0_6844, \7063 );
and \U$34330 ( \40011 , RIe5331c8_6882, \40010 );
and \U$34331 ( \40012 , \40007 , \7061 , RIe549770_6843, RIe548ff0_6844, \7063 );
and \U$34332 ( \40013 , RIe5339c0_6881, \40012 );
and \U$34333 ( \40014 , RIe5319e0_6884, RIe549ef0_6842, \7062 , RIe548ff0_6844, \7063 );
and \U$34334 ( \40015 , RIeab87c8_6898, \40014 );
and \U$34335 ( \40016 , \40007 , RIe549ef0_6842, \7062 , RIe548ff0_6844, \7063 );
and \U$34336 ( \40017 , RIe5341b8_6880, \40016 );
and \U$34337 ( \40018 , RIe5319e0_6884, \7061 , \7062 , RIe548ff0_6844, \7063 );
and \U$34338 ( \40019 , RIe5349b0_6879, \40018 );
and \U$34339 ( \40020 , \40007 , \7061 , \7062 , RIe548ff0_6844, \7063 );
and \U$34340 ( \40021 , RIea94af8_6890, \40020 );
nor \U$34341 ( \40022 , \40007 , \7061 , \7062 , RIe548ff0_6844, RIea91330_6888);
and \U$34342 ( \40023 , RIe5351a8_6878, \40022 );
nor \U$34343 ( \40024 , RIe5319e0_6884, \7061 , \7062 , RIe548ff0_6844, RIea91330_6888);
and \U$34344 ( \40025 , RIe5359a0_6877, \40024 );
nor \U$34345 ( \40026 , \40007 , RIe549ef0_6842, \7062 , RIe548ff0_6844, RIea91330_6888);
and \U$34346 ( \40027 , RIeab78c8_6895, \40026 );
nor \U$34347 ( \40028 , RIe5319e0_6884, RIe549ef0_6842, \7062 , RIe548ff0_6844, RIea91330_6888);
and \U$34348 ( \40029 , RIeab7d00_6896, \40028 );
nor \U$34349 ( \40030 , \40007 , \7061 , RIe549770_6843, RIe548ff0_6844, RIea91330_6888);
and \U$34350 ( \40031 , RIeacfa18_6902, \40030 );
nor \U$34351 ( \40032 , RIe5319e0_6884, \7061 , RIe549770_6843, RIe548ff0_6844, RIea91330_6888);
and \U$34352 ( \40033 , RIeab6518_6891, \40032 );
nor \U$34353 ( \40034 , \40007 , RIe549ef0_6842, RIe549770_6843, RIe548ff0_6844, RIea91330_6888);
and \U$34354 ( \40035 , RIeb352c8_6904, \40034 );
or \U$34355 ( \40036 , \40004 , \40006 , \40009 , \40011 , \40013 , \40015 , \40017 , \40019 , \40021 , \40023 , \40025 , \40027 , \40029 , \40031 , \40033 , \40035 );
buf \U$34356 ( \40037 , RIe549ef0_6842);
buf \U$34357 ( \40038 , RIe549770_6843);
buf \U$34358 ( \40039 , RIe548ff0_6844);
buf \U$34359 ( \40040 , RIea91330_6888);
buf \U$34360 ( \40041 , RIe5319e0_6884);
nor \U$34361 ( \40042 , \40037 , \40038 , \40039 , \40040 , \40041 );
buf \U$34362 ( \40043 , \40042 );
buf \U$34363 ( \40044 , RIea91330_6888);
buf \U$34364 ( \40045 , RIe5319e0_6884);
buf \U$34365 ( \40046 , RIe549ef0_6842);
buf \U$34366 ( \40047 , RIe549770_6843);
buf \U$34367 ( \40048 , RIe548ff0_6844);
or \U$34368 ( \40049 , \40045 , \40046 , \40047 , \40048 );
and \U$34369 ( \40050 , \40044 , \40049 );
buf \U$34370 ( \40051 , \40050 );
or \U$34371 ( \40052 , \40043 , \40051 );
_DC gb3a4 ( \40053_nGb3a4 , \40036 , \40052 );
not \U$34372 ( \40054 , \40053_nGb3a4 );
buf \U$34373 ( \40055 , RIb7b9608_246);
and \U$34374 ( \40056 , \7117 , \40003 );
and \U$34375 ( \40057 , \7119 , \40005 );
and \U$34376 ( \40058 , \7864 , \40008 );
and \U$34377 ( \40059 , \7892 , \40010 );
and \U$34378 ( \40060 , \7920 , \40012 );
and \U$34379 ( \40061 , \7948 , \40014 );
and \U$34380 ( \40062 , \7976 , \40016 );
and \U$34381 ( \40063 , \8004 , \40018 );
and \U$34382 ( \40064 , \8032 , \40020 );
and \U$34383 ( \40065 , \8060 , \40022 );
and \U$34384 ( \40066 , \8088 , \40024 );
and \U$34385 ( \40067 , \8116 , \40026 );
and \U$34386 ( \40068 , \8144 , \40028 );
and \U$34387 ( \40069 , \8172 , \40030 );
and \U$34388 ( \40070 , \8200 , \40032 );
and \U$34389 ( \40071 , \8228 , \40034 );
or \U$34390 ( \40072 , \40056 , \40057 , \40058 , \40059 , \40060 , \40061 , \40062 , \40063 , \40064 , \40065 , \40066 , \40067 , \40068 , \40069 , \40070 , \40071 );
_DC gb3b8 ( \40073_nGb3b8 , \40072 , \40052 );
buf \U$34391 ( \40074 , \40073_nGb3b8 );
xor \U$34392 ( \40075 , \40055 , \40074 );
buf \U$34393 ( \40076 , RIb7b9590_247);
and \U$34394 ( \40077 , \7126 , \40003 );
and \U$34395 ( \40078 , \7128 , \40005 );
and \U$34396 ( \40079 , \8338 , \40008 );
and \U$34397 ( \40080 , \8340 , \40010 );
and \U$34398 ( \40081 , \8342 , \40012 );
and \U$34399 ( \40082 , \8344 , \40014 );
and \U$34400 ( \40083 , \8346 , \40016 );
and \U$34401 ( \40084 , \8348 , \40018 );
and \U$34402 ( \40085 , \8350 , \40020 );
and \U$34403 ( \40086 , \8352 , \40022 );
and \U$34404 ( \40087 , \8354 , \40024 );
and \U$34405 ( \40088 , \8356 , \40026 );
and \U$34406 ( \40089 , \8358 , \40028 );
and \U$34407 ( \40090 , \8360 , \40030 );
and \U$34408 ( \40091 , \8362 , \40032 );
and \U$34409 ( \40092 , \8364 , \40034 );
or \U$34410 ( \40093 , \40077 , \40078 , \40079 , \40080 , \40081 , \40082 , \40083 , \40084 , \40085 , \40086 , \40087 , \40088 , \40089 , \40090 , \40091 , \40092 );
_DC gb3cd ( \40094_nGb3cd , \40093 , \40052 );
buf \U$34411 ( \40095 , \40094_nGb3cd );
xor \U$34412 ( \40096 , \40076 , \40095 );
or \U$34413 ( \40097 , \40075 , \40096 );
buf \U$34414 ( \40098 , RIb7b9518_248);
and \U$34415 ( \40099 , \7136 , \40003 );
and \U$34416 ( \40100 , \7138 , \40005 );
and \U$34417 ( \40101 , \8374 , \40008 );
and \U$34418 ( \40102 , \8376 , \40010 );
and \U$34419 ( \40103 , \8378 , \40012 );
and \U$34420 ( \40104 , \8380 , \40014 );
and \U$34421 ( \40105 , \8382 , \40016 );
and \U$34422 ( \40106 , \8384 , \40018 );
and \U$34423 ( \40107 , \8386 , \40020 );
and \U$34424 ( \40108 , \8388 , \40022 );
and \U$34425 ( \40109 , \8390 , \40024 );
and \U$34426 ( \40110 , \8392 , \40026 );
and \U$34427 ( \40111 , \8394 , \40028 );
and \U$34428 ( \40112 , \8396 , \40030 );
and \U$34429 ( \40113 , \8398 , \40032 );
and \U$34430 ( \40114 , \8400 , \40034 );
or \U$34431 ( \40115 , \40099 , \40100 , \40101 , \40102 , \40103 , \40104 , \40105 , \40106 , \40107 , \40108 , \40109 , \40110 , \40111 , \40112 , \40113 , \40114 );
_DC gb3e3 ( \40116_nGb3e3 , \40115 , \40052 );
buf \U$34432 ( \40117 , \40116_nGb3e3 );
xor \U$34433 ( \40118 , \40098 , \40117 );
or \U$34434 ( \40119 , \40097 , \40118 );
buf \U$34435 ( \40120 , RIb7b94a0_249);
and \U$34436 ( \40121 , \7146 , \40003 );
and \U$34437 ( \40122 , \7148 , \40005 );
and \U$34438 ( \40123 , \8410 , \40008 );
and \U$34439 ( \40124 , \8412 , \40010 );
and \U$34440 ( \40125 , \8414 , \40012 );
and \U$34441 ( \40126 , \8416 , \40014 );
and \U$34442 ( \40127 , \8418 , \40016 );
and \U$34443 ( \40128 , \8420 , \40018 );
and \U$34444 ( \40129 , \8422 , \40020 );
and \U$34445 ( \40130 , \8424 , \40022 );
and \U$34446 ( \40131 , \8426 , \40024 );
and \U$34447 ( \40132 , \8428 , \40026 );
and \U$34448 ( \40133 , \8430 , \40028 );
and \U$34449 ( \40134 , \8432 , \40030 );
and \U$34450 ( \40135 , \8434 , \40032 );
and \U$34451 ( \40136 , \8436 , \40034 );
or \U$34452 ( \40137 , \40121 , \40122 , \40123 , \40124 , \40125 , \40126 , \40127 , \40128 , \40129 , \40130 , \40131 , \40132 , \40133 , \40134 , \40135 , \40136 );
_DC gb3f9 ( \40138_nGb3f9 , \40137 , \40052 );
buf \U$34453 ( \40139 , \40138_nGb3f9 );
xor \U$34454 ( \40140 , \40120 , \40139 );
or \U$34455 ( \40141 , \40119 , \40140 );
buf \U$34456 ( \40142 , RIb7b9428_250);
and \U$34457 ( \40143 , \7156 , \40003 );
and \U$34458 ( \40144 , \7158 , \40005 );
and \U$34459 ( \40145 , \8446 , \40008 );
and \U$34460 ( \40146 , \8448 , \40010 );
and \U$34461 ( \40147 , \8450 , \40012 );
and \U$34462 ( \40148 , \8452 , \40014 );
and \U$34463 ( \40149 , \8454 , \40016 );
and \U$34464 ( \40150 , \8456 , \40018 );
and \U$34465 ( \40151 , \8458 , \40020 );
and \U$34466 ( \40152 , \8460 , \40022 );
and \U$34467 ( \40153 , \8462 , \40024 );
and \U$34468 ( \40154 , \8464 , \40026 );
and \U$34469 ( \40155 , \8466 , \40028 );
and \U$34470 ( \40156 , \8468 , \40030 );
and \U$34471 ( \40157 , \8470 , \40032 );
and \U$34472 ( \40158 , \8472 , \40034 );
or \U$34473 ( \40159 , \40143 , \40144 , \40145 , \40146 , \40147 , \40148 , \40149 , \40150 , \40151 , \40152 , \40153 , \40154 , \40155 , \40156 , \40157 , \40158 );
_DC gb40f ( \40160_nGb40f , \40159 , \40052 );
buf \U$34474 ( \40161 , \40160_nGb40f );
xor \U$34475 ( \40162 , \40142 , \40161 );
or \U$34476 ( \40163 , \40141 , \40162 );
buf \U$34477 ( \40164 , RIb7b93b0_251);
and \U$34478 ( \40165 , \7166 , \40003 );
and \U$34479 ( \40166 , \7168 , \40005 );
and \U$34480 ( \40167 , \8482 , \40008 );
and \U$34481 ( \40168 , \8484 , \40010 );
and \U$34482 ( \40169 , \8486 , \40012 );
and \U$34483 ( \40170 , \8488 , \40014 );
and \U$34484 ( \40171 , \8490 , \40016 );
and \U$34485 ( \40172 , \8492 , \40018 );
and \U$34486 ( \40173 , \8494 , \40020 );
and \U$34487 ( \40174 , \8496 , \40022 );
and \U$34488 ( \40175 , \8498 , \40024 );
and \U$34489 ( \40176 , \8500 , \40026 );
and \U$34490 ( \40177 , \8502 , \40028 );
and \U$34491 ( \40178 , \8504 , \40030 );
and \U$34492 ( \40179 , \8506 , \40032 );
and \U$34493 ( \40180 , \8508 , \40034 );
or \U$34494 ( \40181 , \40165 , \40166 , \40167 , \40168 , \40169 , \40170 , \40171 , \40172 , \40173 , \40174 , \40175 , \40176 , \40177 , \40178 , \40179 , \40180 );
_DC gb425 ( \40182_nGb425 , \40181 , \40052 );
buf \U$34495 ( \40183 , \40182_nGb425 );
xor \U$34496 ( \40184 , \40164 , \40183 );
or \U$34497 ( \40185 , \40163 , \40184 );
buf \U$34498 ( \40186 , RIb7af720_252);
and \U$34499 ( \40187 , \7176 , \40003 );
and \U$34500 ( \40188 , \7178 , \40005 );
and \U$34501 ( \40189 , \8518 , \40008 );
and \U$34502 ( \40190 , \8520 , \40010 );
and \U$34503 ( \40191 , \8522 , \40012 );
and \U$34504 ( \40192 , \8524 , \40014 );
and \U$34505 ( \40193 , \8526 , \40016 );
and \U$34506 ( \40194 , \8528 , \40018 );
and \U$34507 ( \40195 , \8530 , \40020 );
and \U$34508 ( \40196 , \8532 , \40022 );
and \U$34509 ( \40197 , \8534 , \40024 );
and \U$34510 ( \40198 , \8536 , \40026 );
and \U$34511 ( \40199 , \8538 , \40028 );
and \U$34512 ( \40200 , \8540 , \40030 );
and \U$34513 ( \40201 , \8542 , \40032 );
and \U$34514 ( \40202 , \8544 , \40034 );
or \U$34515 ( \40203 , \40187 , \40188 , \40189 , \40190 , \40191 , \40192 , \40193 , \40194 , \40195 , \40196 , \40197 , \40198 , \40199 , \40200 , \40201 , \40202 );
_DC gb43b ( \40204_nGb43b , \40203 , \40052 );
buf \U$34516 ( \40205 , \40204_nGb43b );
xor \U$34517 ( \40206 , \40186 , \40205 );
or \U$34518 ( \40207 , \40185 , \40206 );
buf \U$34519 ( \40208 , RIb7af6a8_253);
and \U$34520 ( \40209 , \7186 , \40003 );
and \U$34521 ( \40210 , \7188 , \40005 );
and \U$34522 ( \40211 , \8554 , \40008 );
and \U$34523 ( \40212 , \8556 , \40010 );
and \U$34524 ( \40213 , \8558 , \40012 );
and \U$34525 ( \40214 , \8560 , \40014 );
and \U$34526 ( \40215 , \8562 , \40016 );
and \U$34527 ( \40216 , \8564 , \40018 );
and \U$34528 ( \40217 , \8566 , \40020 );
and \U$34529 ( \40218 , \8568 , \40022 );
and \U$34530 ( \40219 , \8570 , \40024 );
and \U$34531 ( \40220 , \8572 , \40026 );
and \U$34532 ( \40221 , \8574 , \40028 );
and \U$34533 ( \40222 , \8576 , \40030 );
and \U$34534 ( \40223 , \8578 , \40032 );
and \U$34535 ( \40224 , \8580 , \40034 );
or \U$34536 ( \40225 , \40209 , \40210 , \40211 , \40212 , \40213 , \40214 , \40215 , \40216 , \40217 , \40218 , \40219 , \40220 , \40221 , \40222 , \40223 , \40224 );
_DC gb451 ( \40226_nGb451 , \40225 , \40052 );
buf \U$34537 ( \40227 , \40226_nGb451 );
xor \U$34538 ( \40228 , \40208 , \40227 );
or \U$34539 ( \40229 , \40207 , \40228 );
not \U$34540 ( \40230 , \40229 );
buf \U$34541 ( \40231 , \40230 );
buf \U$34542 ( \40232 , RIb7af630_254);
and \U$34543 ( \40233 , \7198 , \40003 );
and \U$34544 ( \40234 , \7200 , \40005 );
and \U$34545 ( \40235 , \8645 , \40008 );
and \U$34546 ( \40236 , \8673 , \40010 );
and \U$34547 ( \40237 , \8701 , \40012 );
and \U$34548 ( \40238 , \8729 , \40014 );
and \U$34549 ( \40239 , \8757 , \40016 );
and \U$34550 ( \40240 , \8785 , \40018 );
and \U$34551 ( \40241 , \8813 , \40020 );
and \U$34552 ( \40242 , \8841 , \40022 );
and \U$34553 ( \40243 , \8869 , \40024 );
and \U$34554 ( \40244 , \8897 , \40026 );
and \U$34555 ( \40245 , \8925 , \40028 );
and \U$34556 ( \40246 , \8953 , \40030 );
and \U$34557 ( \40247 , \8981 , \40032 );
and \U$34558 ( \40248 , \9009 , \40034 );
or \U$34559 ( \40249 , \40233 , \40234 , \40235 , \40236 , \40237 , \40238 , \40239 , \40240 , \40241 , \40242 , \40243 , \40244 , \40245 , \40246 , \40247 , \40248 );
_DC gb469 ( \40250_nGb469 , \40249 , \40052 );
buf \U$34560 ( \40251 , \40250_nGb469 );
xor \U$34561 ( \40252 , \40232 , \40251 );
buf \U$34562 ( \40253 , RIb7af5b8_255);
and \U$34563 ( \40254 , \7207 , \40003 );
and \U$34564 ( \40255 , \7209 , \40005 );
and \U$34565 ( \40256 , \9119 , \40008 );
and \U$34566 ( \40257 , \9121 , \40010 );
and \U$34567 ( \40258 , \9123 , \40012 );
and \U$34568 ( \40259 , \9125 , \40014 );
and \U$34569 ( \40260 , \9127 , \40016 );
and \U$34570 ( \40261 , \9129 , \40018 );
and \U$34571 ( \40262 , \9131 , \40020 );
and \U$34572 ( \40263 , \9133 , \40022 );
and \U$34573 ( \40264 , \9135 , \40024 );
and \U$34574 ( \40265 , \9137 , \40026 );
and \U$34575 ( \40266 , \9139 , \40028 );
and \U$34576 ( \40267 , \9141 , \40030 );
and \U$34577 ( \40268 , \9143 , \40032 );
and \U$34578 ( \40269 , \9145 , \40034 );
or \U$34579 ( \40270 , \40254 , \40255 , \40256 , \40257 , \40258 , \40259 , \40260 , \40261 , \40262 , \40263 , \40264 , \40265 , \40266 , \40267 , \40268 , \40269 );
_DC gb47e ( \40271_nGb47e , \40270 , \40052 );
buf \U$34580 ( \40272 , \40271_nGb47e );
xor \U$34581 ( \40273 , \40253 , \40272 );
or \U$34582 ( \40274 , \40252 , \40273 );
buf \U$34583 ( \40275 , RIb7af540_256);
and \U$34584 ( \40276 , \7217 , \40003 );
and \U$34585 ( \40277 , \7219 , \40005 );
and \U$34586 ( \40278 , \9155 , \40008 );
and \U$34587 ( \40279 , \9157 , \40010 );
and \U$34588 ( \40280 , \9159 , \40012 );
and \U$34589 ( \40281 , \9161 , \40014 );
and \U$34590 ( \40282 , \9163 , \40016 );
and \U$34591 ( \40283 , \9165 , \40018 );
and \U$34592 ( \40284 , \9167 , \40020 );
and \U$34593 ( \40285 , \9169 , \40022 );
and \U$34594 ( \40286 , \9171 , \40024 );
and \U$34595 ( \40287 , \9173 , \40026 );
and \U$34596 ( \40288 , \9175 , \40028 );
and \U$34597 ( \40289 , \9177 , \40030 );
and \U$34598 ( \40290 , \9179 , \40032 );
and \U$34599 ( \40291 , \9181 , \40034 );
or \U$34600 ( \40292 , \40276 , \40277 , \40278 , \40279 , \40280 , \40281 , \40282 , \40283 , \40284 , \40285 , \40286 , \40287 , \40288 , \40289 , \40290 , \40291 );
_DC gb494 ( \40293_nGb494 , \40292 , \40052 );
buf \U$34601 ( \40294 , \40293_nGb494 );
xor \U$34602 ( \40295 , \40275 , \40294 );
or \U$34603 ( \40296 , \40274 , \40295 );
buf \U$34604 ( \40297 , RIb7af4c8_257);
and \U$34605 ( \40298 , \7227 , \40003 );
and \U$34606 ( \40299 , \7229 , \40005 );
and \U$34607 ( \40300 , \9191 , \40008 );
and \U$34608 ( \40301 , \9193 , \40010 );
and \U$34609 ( \40302 , \9195 , \40012 );
and \U$34610 ( \40303 , \9197 , \40014 );
and \U$34611 ( \40304 , \9199 , \40016 );
and \U$34612 ( \40305 , \9201 , \40018 );
and \U$34613 ( \40306 , \9203 , \40020 );
and \U$34614 ( \40307 , \9205 , \40022 );
and \U$34615 ( \40308 , \9207 , \40024 );
and \U$34616 ( \40309 , \9209 , \40026 );
and \U$34617 ( \40310 , \9211 , \40028 );
and \U$34618 ( \40311 , \9213 , \40030 );
and \U$34619 ( \40312 , \9215 , \40032 );
and \U$34620 ( \40313 , \9217 , \40034 );
or \U$34621 ( \40314 , \40298 , \40299 , \40300 , \40301 , \40302 , \40303 , \40304 , \40305 , \40306 , \40307 , \40308 , \40309 , \40310 , \40311 , \40312 , \40313 );
_DC gb4aa ( \40315_nGb4aa , \40314 , \40052 );
buf \U$34622 ( \40316 , \40315_nGb4aa );
xor \U$34623 ( \40317 , \40297 , \40316 );
or \U$34624 ( \40318 , \40296 , \40317 );
buf \U$34625 ( \40319 , RIb7af450_258);
and \U$34626 ( \40320 , \7237 , \40003 );
and \U$34627 ( \40321 , \7239 , \40005 );
and \U$34628 ( \40322 , \9227 , \40008 );
and \U$34629 ( \40323 , \9229 , \40010 );
and \U$34630 ( \40324 , \9231 , \40012 );
and \U$34631 ( \40325 , \9233 , \40014 );
and \U$34632 ( \40326 , \9235 , \40016 );
and \U$34633 ( \40327 , \9237 , \40018 );
and \U$34634 ( \40328 , \9239 , \40020 );
and \U$34635 ( \40329 , \9241 , \40022 );
and \U$34636 ( \40330 , \9243 , \40024 );
and \U$34637 ( \40331 , \9245 , \40026 );
and \U$34638 ( \40332 , \9247 , \40028 );
and \U$34639 ( \40333 , \9249 , \40030 );
and \U$34640 ( \40334 , \9251 , \40032 );
and \U$34641 ( \40335 , \9253 , \40034 );
or \U$34642 ( \40336 , \40320 , \40321 , \40322 , \40323 , \40324 , \40325 , \40326 , \40327 , \40328 , \40329 , \40330 , \40331 , \40332 , \40333 , \40334 , \40335 );
_DC gb4c0 ( \40337_nGb4c0 , \40336 , \40052 );
buf \U$34643 ( \40338 , \40337_nGb4c0 );
xor \U$34644 ( \40339 , \40319 , \40338 );
or \U$34645 ( \40340 , \40318 , \40339 );
buf \U$34646 ( \40341 , RIb7af3d8_259);
and \U$34647 ( \40342 , \7247 , \40003 );
and \U$34648 ( \40343 , \7249 , \40005 );
and \U$34649 ( \40344 , \9263 , \40008 );
and \U$34650 ( \40345 , \9265 , \40010 );
and \U$34651 ( \40346 , \9267 , \40012 );
and \U$34652 ( \40347 , \9269 , \40014 );
and \U$34653 ( \40348 , \9271 , \40016 );
and \U$34654 ( \40349 , \9273 , \40018 );
and \U$34655 ( \40350 , \9275 , \40020 );
and \U$34656 ( \40351 , \9277 , \40022 );
and \U$34657 ( \40352 , \9279 , \40024 );
and \U$34658 ( \40353 , \9281 , \40026 );
and \U$34659 ( \40354 , \9283 , \40028 );
and \U$34660 ( \40355 , \9285 , \40030 );
and \U$34661 ( \40356 , \9287 , \40032 );
and \U$34662 ( \40357 , \9289 , \40034 );
or \U$34663 ( \40358 , \40342 , \40343 , \40344 , \40345 , \40346 , \40347 , \40348 , \40349 , \40350 , \40351 , \40352 , \40353 , \40354 , \40355 , \40356 , \40357 );
_DC gb4d6 ( \40359_nGb4d6 , \40358 , \40052 );
buf \U$34664 ( \40360 , \40359_nGb4d6 );
xor \U$34665 ( \40361 , \40341 , \40360 );
or \U$34666 ( \40362 , \40340 , \40361 );
buf \U$34667 ( \40363 , RIb7a5bf8_260);
and \U$34668 ( \40364 , \7257 , \40003 );
and \U$34669 ( \40365 , \7259 , \40005 );
and \U$34670 ( \40366 , \9299 , \40008 );
and \U$34671 ( \40367 , \9301 , \40010 );
and \U$34672 ( \40368 , \9303 , \40012 );
and \U$34673 ( \40369 , \9305 , \40014 );
and \U$34674 ( \40370 , \9307 , \40016 );
and \U$34675 ( \40371 , \9309 , \40018 );
and \U$34676 ( \40372 , \9311 , \40020 );
and \U$34677 ( \40373 , \9313 , \40022 );
and \U$34678 ( \40374 , \9315 , \40024 );
and \U$34679 ( \40375 , \9317 , \40026 );
and \U$34680 ( \40376 , \9319 , \40028 );
and \U$34681 ( \40377 , \9321 , \40030 );
and \U$34682 ( \40378 , \9323 , \40032 );
and \U$34683 ( \40379 , \9325 , \40034 );
or \U$34684 ( \40380 , \40364 , \40365 , \40366 , \40367 , \40368 , \40369 , \40370 , \40371 , \40372 , \40373 , \40374 , \40375 , \40376 , \40377 , \40378 , \40379 );
_DC gb4ec ( \40381_nGb4ec , \40380 , \40052 );
buf \U$34685 ( \40382 , \40381_nGb4ec );
xor \U$34686 ( \40383 , \40363 , \40382 );
or \U$34687 ( \40384 , \40362 , \40383 );
buf \U$34688 ( \40385 , RIb7a0c48_261);
and \U$34689 ( \40386 , \7267 , \40003 );
and \U$34690 ( \40387 , \7269 , \40005 );
and \U$34691 ( \40388 , \9335 , \40008 );
and \U$34692 ( \40389 , \9337 , \40010 );
and \U$34693 ( \40390 , \9339 , \40012 );
and \U$34694 ( \40391 , \9341 , \40014 );
and \U$34695 ( \40392 , \9343 , \40016 );
and \U$34696 ( \40393 , \9345 , \40018 );
and \U$34697 ( \40394 , \9347 , \40020 );
and \U$34698 ( \40395 , \9349 , \40022 );
and \U$34699 ( \40396 , \9351 , \40024 );
and \U$34700 ( \40397 , \9353 , \40026 );
and \U$34701 ( \40398 , \9355 , \40028 );
and \U$34702 ( \40399 , \9357 , \40030 );
and \U$34703 ( \40400 , \9359 , \40032 );
and \U$34704 ( \40401 , \9361 , \40034 );
or \U$34705 ( \40402 , \40386 , \40387 , \40388 , \40389 , \40390 , \40391 , \40392 , \40393 , \40394 , \40395 , \40396 , \40397 , \40398 , \40399 , \40400 , \40401 );
_DC gb502 ( \40403_nGb502 , \40402 , \40052 );
buf \U$34706 ( \40404 , \40403_nGb502 );
xor \U$34707 ( \40405 , \40385 , \40404 );
or \U$34708 ( \40406 , \40384 , \40405 );
not \U$34709 ( \40407 , \40406 );
buf \U$34710 ( \40408 , \40407 );
and \U$34711 ( \40409 , \40231 , \40408 );
and \U$34712 ( \40410 , \40054 , \40409 );
_HMUX gb50a ( \40411_nGb50a , \40002_nGb36e , RIe5319e0_6884 , \40410 );
buf \U$34713 ( \40412 , RIe5319e0_6884);
buf \U$34715 ( \40413 , \40412 );
not \U$34717 ( \40414 , \40413 );
buf \U$34718 ( \40415 , RIe549ef0_6842);
buf \U$34720 ( \40416 , \40415 );
not \U$34721 ( \40417 , \40416 );
buf \U$34722 ( \40418 , RIe549770_6843);
buf \U$34724 ( \40419 , \40418 );
not \U$34725 ( \40420 , \40419 );
buf \U$34726 ( \40421 , RIe548ff0_6844);
buf \U$34728 ( \40422 , \40421 );
not \U$34729 ( \40423 , \40422 );
buf \U$34730 ( \40424 , RIea91330_6888);
not \U$34731 ( \40425 , \40424 );
buf \U$34732 ( \40426 , \40425 );
buf \U$34733 ( \40427 , \40425 );
buf \U$34734 ( \40428 , \40427 );
buf \U$34735 ( \40429 , \40427 );
buf \U$34736 ( \40430 , \40427 );
buf \U$34737 ( \40431 , \40427 );
buf \U$34738 ( \40432 , \40427 );
buf \U$34739 ( \40433 , \40427 );
buf \U$34740 ( \40434 , \40427 );
buf \U$34741 ( \40435 , \40427 );
buf \U$34742 ( \40436 , \40427 );
buf \U$34743 ( \40437 , \40427 );
buf \U$34744 ( \40438 , \40427 );
buf \U$34745 ( \40439 , \40427 );
buf \U$34746 ( \40440 , \40427 );
buf \U$34747 ( \40441 , \40427 );
buf \U$34748 ( \40442 , \40427 );
buf \U$34749 ( \40443 , \40427 );
buf \U$34750 ( \40444 , \40427 );
buf \U$34751 ( \40445 , \40427 );
buf \U$34752 ( \40446 , \40427 );
buf \U$34753 ( \40447 , \40427 );
buf \U$34754 ( \40448 , \40427 );
buf \U$34755 ( \40449 , \40427 );
buf \U$34756 ( \40450 , \40427 );
buf \U$34757 ( \40451 , \40427 );
buf \U$34758 ( \40452 , \40427 );
buf \U$34759 ( \40453 , \40427 );
nor \U$34760 ( \40454 , \40414 , \40417 , \40420 , \40423 , \40426 , \40427 , \40428 , \40429 , \40430 , \40431 , \40432 , \40433 , \40434 , \40435 , \40436 , \40437 , \40438 , \40439 , \40440 , \40441 , \40442 , \40443 , \40444 , \40445 , \40446 , \40447 , \40448 , \40449 , \40450 , \40451 , \40452 , \40453 );
and \U$34761 ( \40455 , RIeb72150_6905, \40454 );
buf \U$34762 ( \40456 , \40427 );
buf \U$34763 ( \40457 , \40427 );
buf \U$34764 ( \40458 , \40427 );
buf \U$34765 ( \40459 , \40427 );
buf \U$34766 ( \40460 , \40427 );
buf \U$34767 ( \40461 , \40427 );
buf \U$34768 ( \40462 , \40427 );
buf \U$34769 ( \40463 , \40427 );
buf \U$34770 ( \40464 , \40427 );
buf \U$34771 ( \40465 , \40427 );
buf \U$34772 ( \40466 , \40427 );
buf \U$34773 ( \40467 , \40427 );
buf \U$34774 ( \40468 , \40427 );
buf \U$34775 ( \40469 , \40427 );
buf \U$34776 ( \40470 , \40427 );
buf \U$34777 ( \40471 , \40427 );
buf \U$34778 ( \40472 , \40427 );
buf \U$34779 ( \40473 , \40427 );
buf \U$34780 ( \40474 , \40427 );
buf \U$34781 ( \40475 , \40427 );
buf \U$34782 ( \40476 , \40427 );
buf \U$34783 ( \40477 , \40427 );
buf \U$34784 ( \40478 , \40427 );
buf \U$34785 ( \40479 , \40427 );
buf \U$34786 ( \40480 , \40427 );
buf \U$34787 ( \40481 , \40427 );
nor \U$34788 ( \40482 , \40413 , \40417 , \40420 , \40423 , \40426 , \40427 , \40456 , \40457 , \40458 , \40459 , \40460 , \40461 , \40462 , \40463 , \40464 , \40465 , \40466 , \40467 , \40468 , \40469 , \40470 , \40471 , \40472 , \40473 , \40474 , \40475 , \40476 , \40477 , \40478 , \40479 , \40480 , \40481 );
and \U$34789 ( \40483 , RIeab80c0_6897, \40482 );
buf \U$34790 ( \40484 , \40427 );
buf \U$34791 ( \40485 , \40427 );
buf \U$34792 ( \40486 , \40427 );
buf \U$34793 ( \40487 , \40427 );
buf \U$34794 ( \40488 , \40427 );
buf \U$34795 ( \40489 , \40427 );
buf \U$34796 ( \40490 , \40427 );
buf \U$34797 ( \40491 , \40427 );
buf \U$34798 ( \40492 , \40427 );
buf \U$34799 ( \40493 , \40427 );
buf \U$34800 ( \40494 , \40427 );
buf \U$34801 ( \40495 , \40427 );
buf \U$34802 ( \40496 , \40427 );
buf \U$34803 ( \40497 , \40427 );
buf \U$34804 ( \40498 , \40427 );
buf \U$34805 ( \40499 , \40427 );
buf \U$34806 ( \40500 , \40427 );
buf \U$34807 ( \40501 , \40427 );
buf \U$34808 ( \40502 , \40427 );
buf \U$34809 ( \40503 , \40427 );
buf \U$34810 ( \40504 , \40427 );
buf \U$34811 ( \40505 , \40427 );
buf \U$34812 ( \40506 , \40427 );
buf \U$34813 ( \40507 , \40427 );
buf \U$34814 ( \40508 , \40427 );
buf \U$34815 ( \40509 , \40427 );
nor \U$34816 ( \40510 , \40414 , \40416 , \40420 , \40423 , \40426 , \40427 , \40484 , \40485 , \40486 , \40487 , \40488 , \40489 , \40490 , \40491 , \40492 , \40493 , \40494 , \40495 , \40496 , \40497 , \40498 , \40499 , \40500 , \40501 , \40502 , \40503 , \40504 , \40505 , \40506 , \40507 , \40508 , \40509 );
and \U$34817 ( \40511 , RIe5331c8_6882, \40510 );
buf \U$34818 ( \40512 , \40427 );
buf \U$34819 ( \40513 , \40427 );
buf \U$34820 ( \40514 , \40427 );
buf \U$34821 ( \40515 , \40427 );
buf \U$34822 ( \40516 , \40427 );
buf \U$34823 ( \40517 , \40427 );
buf \U$34824 ( \40518 , \40427 );
buf \U$34825 ( \40519 , \40427 );
buf \U$34826 ( \40520 , \40427 );
buf \U$34827 ( \40521 , \40427 );
buf \U$34828 ( \40522 , \40427 );
buf \U$34829 ( \40523 , \40427 );
buf \U$34830 ( \40524 , \40427 );
buf \U$34831 ( \40525 , \40427 );
buf \U$34832 ( \40526 , \40427 );
buf \U$34833 ( \40527 , \40427 );
buf \U$34834 ( \40528 , \40427 );
buf \U$34835 ( \40529 , \40427 );
buf \U$34836 ( \40530 , \40427 );
buf \U$34837 ( \40531 , \40427 );
buf \U$34838 ( \40532 , \40427 );
buf \U$34839 ( \40533 , \40427 );
buf \U$34840 ( \40534 , \40427 );
buf \U$34841 ( \40535 , \40427 );
buf \U$34842 ( \40536 , \40427 );
buf \U$34843 ( \40537 , \40427 );
nor \U$34844 ( \40538 , \40413 , \40416 , \40420 , \40423 , \40426 , \40427 , \40512 , \40513 , \40514 , \40515 , \40516 , \40517 , \40518 , \40519 , \40520 , \40521 , \40522 , \40523 , \40524 , \40525 , \40526 , \40527 , \40528 , \40529 , \40530 , \40531 , \40532 , \40533 , \40534 , \40535 , \40536 , \40537 );
and \U$34845 ( \40539 , RIe5339c0_6881, \40538 );
buf \U$34846 ( \40540 , \40427 );
buf \U$34847 ( \40541 , \40427 );
buf \U$34848 ( \40542 , \40427 );
buf \U$34849 ( \40543 , \40427 );
buf \U$34850 ( \40544 , \40427 );
buf \U$34851 ( \40545 , \40427 );
buf \U$34852 ( \40546 , \40427 );
buf \U$34853 ( \40547 , \40427 );
buf \U$34854 ( \40548 , \40427 );
buf \U$34855 ( \40549 , \40427 );
buf \U$34856 ( \40550 , \40427 );
buf \U$34857 ( \40551 , \40427 );
buf \U$34858 ( \40552 , \40427 );
buf \U$34859 ( \40553 , \40427 );
buf \U$34860 ( \40554 , \40427 );
buf \U$34861 ( \40555 , \40427 );
buf \U$34862 ( \40556 , \40427 );
buf \U$34863 ( \40557 , \40427 );
buf \U$34864 ( \40558 , \40427 );
buf \U$34865 ( \40559 , \40427 );
buf \U$34866 ( \40560 , \40427 );
buf \U$34867 ( \40561 , \40427 );
buf \U$34868 ( \40562 , \40427 );
buf \U$34869 ( \40563 , \40427 );
buf \U$34870 ( \40564 , \40427 );
buf \U$34871 ( \40565 , \40427 );
nor \U$34872 ( \40566 , \40414 , \40417 , \40419 , \40423 , \40426 , \40427 , \40540 , \40541 , \40542 , \40543 , \40544 , \40545 , \40546 , \40547 , \40548 , \40549 , \40550 , \40551 , \40552 , \40553 , \40554 , \40555 , \40556 , \40557 , \40558 , \40559 , \40560 , \40561 , \40562 , \40563 , \40564 , \40565 );
and \U$34873 ( \40567 , RIeab87c8_6898, \40566 );
buf \U$34874 ( \40568 , \40427 );
buf \U$34875 ( \40569 , \40427 );
buf \U$34876 ( \40570 , \40427 );
buf \U$34877 ( \40571 , \40427 );
buf \U$34878 ( \40572 , \40427 );
buf \U$34879 ( \40573 , \40427 );
buf \U$34880 ( \40574 , \40427 );
buf \U$34881 ( \40575 , \40427 );
buf \U$34882 ( \40576 , \40427 );
buf \U$34883 ( \40577 , \40427 );
buf \U$34884 ( \40578 , \40427 );
buf \U$34885 ( \40579 , \40427 );
buf \U$34886 ( \40580 , \40427 );
buf \U$34887 ( \40581 , \40427 );
buf \U$34888 ( \40582 , \40427 );
buf \U$34889 ( \40583 , \40427 );
buf \U$34890 ( \40584 , \40427 );
buf \U$34891 ( \40585 , \40427 );
buf \U$34892 ( \40586 , \40427 );
buf \U$34893 ( \40587 , \40427 );
buf \U$34894 ( \40588 , \40427 );
buf \U$34895 ( \40589 , \40427 );
buf \U$34896 ( \40590 , \40427 );
buf \U$34897 ( \40591 , \40427 );
buf \U$34898 ( \40592 , \40427 );
buf \U$34899 ( \40593 , \40427 );
nor \U$34900 ( \40594 , \40413 , \40417 , \40419 , \40423 , \40426 , \40427 , \40568 , \40569 , \40570 , \40571 , \40572 , \40573 , \40574 , \40575 , \40576 , \40577 , \40578 , \40579 , \40580 , \40581 , \40582 , \40583 , \40584 , \40585 , \40586 , \40587 , \40588 , \40589 , \40590 , \40591 , \40592 , \40593 );
and \U$34901 ( \40595 , RIe5341b8_6880, \40594 );
buf \U$34902 ( \40596 , \40427 );
buf \U$34903 ( \40597 , \40427 );
buf \U$34904 ( \40598 , \40427 );
buf \U$34905 ( \40599 , \40427 );
buf \U$34906 ( \40600 , \40427 );
buf \U$34907 ( \40601 , \40427 );
buf \U$34908 ( \40602 , \40427 );
buf \U$34909 ( \40603 , \40427 );
buf \U$34910 ( \40604 , \40427 );
buf \U$34911 ( \40605 , \40427 );
buf \U$34912 ( \40606 , \40427 );
buf \U$34913 ( \40607 , \40427 );
buf \U$34914 ( \40608 , \40427 );
buf \U$34915 ( \40609 , \40427 );
buf \U$34916 ( \40610 , \40427 );
buf \U$34917 ( \40611 , \40427 );
buf \U$34918 ( \40612 , \40427 );
buf \U$34919 ( \40613 , \40427 );
buf \U$34920 ( \40614 , \40427 );
buf \U$34921 ( \40615 , \40427 );
buf \U$34922 ( \40616 , \40427 );
buf \U$34923 ( \40617 , \40427 );
buf \U$34924 ( \40618 , \40427 );
buf \U$34925 ( \40619 , \40427 );
buf \U$34926 ( \40620 , \40427 );
buf \U$34927 ( \40621 , \40427 );
nor \U$34928 ( \40622 , \40414 , \40416 , \40419 , \40423 , \40426 , \40427 , \40596 , \40597 , \40598 , \40599 , \40600 , \40601 , \40602 , \40603 , \40604 , \40605 , \40606 , \40607 , \40608 , \40609 , \40610 , \40611 , \40612 , \40613 , \40614 , \40615 , \40616 , \40617 , \40618 , \40619 , \40620 , \40621 );
and \U$34929 ( \40623 , RIe5349b0_6879, \40622 );
buf \U$34930 ( \40624 , \40427 );
buf \U$34931 ( \40625 , \40427 );
buf \U$34932 ( \40626 , \40427 );
buf \U$34933 ( \40627 , \40427 );
buf \U$34934 ( \40628 , \40427 );
buf \U$34935 ( \40629 , \40427 );
buf \U$34936 ( \40630 , \40427 );
buf \U$34937 ( \40631 , \40427 );
buf \U$34938 ( \40632 , \40427 );
buf \U$34939 ( \40633 , \40427 );
buf \U$34940 ( \40634 , \40427 );
buf \U$34941 ( \40635 , \40427 );
buf \U$34942 ( \40636 , \40427 );
buf \U$34943 ( \40637 , \40427 );
buf \U$34944 ( \40638 , \40427 );
buf \U$34945 ( \40639 , \40427 );
buf \U$34946 ( \40640 , \40427 );
buf \U$34947 ( \40641 , \40427 );
buf \U$34948 ( \40642 , \40427 );
buf \U$34949 ( \40643 , \40427 );
buf \U$34950 ( \40644 , \40427 );
buf \U$34951 ( \40645 , \40427 );
buf \U$34952 ( \40646 , \40427 );
buf \U$34953 ( \40647 , \40427 );
buf \U$34954 ( \40648 , \40427 );
buf \U$34955 ( \40649 , \40427 );
nor \U$34956 ( \40650 , \40413 , \40416 , \40419 , \40423 , \40426 , \40427 , \40624 , \40625 , \40626 , \40627 , \40628 , \40629 , \40630 , \40631 , \40632 , \40633 , \40634 , \40635 , \40636 , \40637 , \40638 , \40639 , \40640 , \40641 , \40642 , \40643 , \40644 , \40645 , \40646 , \40647 , \40648 , \40649 );
and \U$34957 ( \40651 , RIea94af8_6890, \40650 );
buf \U$34958 ( \40652 , \40427 );
buf \U$34959 ( \40653 , \40427 );
buf \U$34960 ( \40654 , \40427 );
buf \U$34961 ( \40655 , \40427 );
buf \U$34962 ( \40656 , \40427 );
buf \U$34963 ( \40657 , \40427 );
buf \U$34964 ( \40658 , \40427 );
buf \U$34965 ( \40659 , \40427 );
buf \U$34966 ( \40660 , \40427 );
buf \U$34967 ( \40661 , \40427 );
buf \U$34968 ( \40662 , \40427 );
buf \U$34969 ( \40663 , \40427 );
buf \U$34970 ( \40664 , \40427 );
buf \U$34971 ( \40665 , \40427 );
buf \U$34972 ( \40666 , \40427 );
buf \U$34973 ( \40667 , \40427 );
buf \U$34974 ( \40668 , \40427 );
buf \U$34975 ( \40669 , \40427 );
buf \U$34976 ( \40670 , \40427 );
buf \U$34977 ( \40671 , \40427 );
buf \U$34978 ( \40672 , \40427 );
buf \U$34979 ( \40673 , \40427 );
buf \U$34980 ( \40674 , \40427 );
buf \U$34981 ( \40675 , \40427 );
buf \U$34982 ( \40676 , \40427 );
buf \U$34983 ( \40677 , \40427 );
nor \U$34984 ( \40678 , \40414 , \40417 , \40420 , \40422 , \40426 , \40427 , \40652 , \40653 , \40654 , \40655 , \40656 , \40657 , \40658 , \40659 , \40660 , \40661 , \40662 , \40663 , \40664 , \40665 , \40666 , \40667 , \40668 , \40669 , \40670 , \40671 , \40672 , \40673 , \40674 , \40675 , \40676 , \40677 );
and \U$34985 ( \40679 , RIe5351a8_6878, \40678 );
buf \U$34986 ( \40680 , \40427 );
buf \U$34987 ( \40681 , \40427 );
buf \U$34988 ( \40682 , \40427 );
buf \U$34989 ( \40683 , \40427 );
buf \U$34990 ( \40684 , \40427 );
buf \U$34991 ( \40685 , \40427 );
buf \U$34992 ( \40686 , \40427 );
buf \U$34993 ( \40687 , \40427 );
buf \U$34994 ( \40688 , \40427 );
buf \U$34995 ( \40689 , \40427 );
buf \U$34996 ( \40690 , \40427 );
buf \U$34997 ( \40691 , \40427 );
buf \U$34998 ( \40692 , \40427 );
buf \U$34999 ( \40693 , \40427 );
buf \U$35000 ( \40694 , \40427 );
buf \U$35001 ( \40695 , \40427 );
buf \U$35002 ( \40696 , \40427 );
buf \U$35003 ( \40697 , \40427 );
buf \U$35004 ( \40698 , \40427 );
buf \U$35005 ( \40699 , \40427 );
buf \U$35006 ( \40700 , \40427 );
buf \U$35007 ( \40701 , \40427 );
buf \U$35008 ( \40702 , \40427 );
buf \U$35009 ( \40703 , \40427 );
buf \U$35010 ( \40704 , \40427 );
buf \U$35011 ( \40705 , \40427 );
nor \U$35012 ( \40706 , \40413 , \40417 , \40420 , \40422 , \40426 , \40427 , \40680 , \40681 , \40682 , \40683 , \40684 , \40685 , \40686 , \40687 , \40688 , \40689 , \40690 , \40691 , \40692 , \40693 , \40694 , \40695 , \40696 , \40697 , \40698 , \40699 , \40700 , \40701 , \40702 , \40703 , \40704 , \40705 );
and \U$35013 ( \40707 , RIe5359a0_6877, \40706 );
buf \U$35014 ( \40708 , \40427 );
buf \U$35015 ( \40709 , \40427 );
buf \U$35016 ( \40710 , \40427 );
buf \U$35017 ( \40711 , \40427 );
buf \U$35018 ( \40712 , \40427 );
buf \U$35019 ( \40713 , \40427 );
buf \U$35020 ( \40714 , \40427 );
buf \U$35021 ( \40715 , \40427 );
buf \U$35022 ( \40716 , \40427 );
buf \U$35023 ( \40717 , \40427 );
buf \U$35024 ( \40718 , \40427 );
buf \U$35025 ( \40719 , \40427 );
buf \U$35026 ( \40720 , \40427 );
buf \U$35027 ( \40721 , \40427 );
buf \U$35028 ( \40722 , \40427 );
buf \U$35029 ( \40723 , \40427 );
buf \U$35030 ( \40724 , \40427 );
buf \U$35031 ( \40725 , \40427 );
buf \U$35032 ( \40726 , \40427 );
buf \U$35033 ( \40727 , \40427 );
buf \U$35034 ( \40728 , \40427 );
buf \U$35035 ( \40729 , \40427 );
buf \U$35036 ( \40730 , \40427 );
buf \U$35037 ( \40731 , \40427 );
buf \U$35038 ( \40732 , \40427 );
buf \U$35039 ( \40733 , \40427 );
nor \U$35040 ( \40734 , \40414 , \40416 , \40420 , \40422 , \40426 , \40427 , \40708 , \40709 , \40710 , \40711 , \40712 , \40713 , \40714 , \40715 , \40716 , \40717 , \40718 , \40719 , \40720 , \40721 , \40722 , \40723 , \40724 , \40725 , \40726 , \40727 , \40728 , \40729 , \40730 , \40731 , \40732 , \40733 );
and \U$35041 ( \40735 , RIeab78c8_6895, \40734 );
buf \U$35042 ( \40736 , \40427 );
buf \U$35043 ( \40737 , \40427 );
buf \U$35044 ( \40738 , \40427 );
buf \U$35045 ( \40739 , \40427 );
buf \U$35046 ( \40740 , \40427 );
buf \U$35047 ( \40741 , \40427 );
buf \U$35048 ( \40742 , \40427 );
buf \U$35049 ( \40743 , \40427 );
buf \U$35050 ( \40744 , \40427 );
buf \U$35051 ( \40745 , \40427 );
buf \U$35052 ( \40746 , \40427 );
buf \U$35053 ( \40747 , \40427 );
buf \U$35054 ( \40748 , \40427 );
buf \U$35055 ( \40749 , \40427 );
buf \U$35056 ( \40750 , \40427 );
buf \U$35057 ( \40751 , \40427 );
buf \U$35058 ( \40752 , \40427 );
buf \U$35059 ( \40753 , \40427 );
buf \U$35060 ( \40754 , \40427 );
buf \U$35061 ( \40755 , \40427 );
buf \U$35062 ( \40756 , \40427 );
buf \U$35063 ( \40757 , \40427 );
buf \U$35064 ( \40758 , \40427 );
buf \U$35065 ( \40759 , \40427 );
buf \U$35066 ( \40760 , \40427 );
buf \U$35067 ( \40761 , \40427 );
nor \U$35068 ( \40762 , \40413 , \40416 , \40420 , \40422 , \40426 , \40427 , \40736 , \40737 , \40738 , \40739 , \40740 , \40741 , \40742 , \40743 , \40744 , \40745 , \40746 , \40747 , \40748 , \40749 , \40750 , \40751 , \40752 , \40753 , \40754 , \40755 , \40756 , \40757 , \40758 , \40759 , \40760 , \40761 );
and \U$35069 ( \40763 , RIeab7d00_6896, \40762 );
buf \U$35070 ( \40764 , \40427 );
buf \U$35071 ( \40765 , \40427 );
buf \U$35072 ( \40766 , \40427 );
buf \U$35073 ( \40767 , \40427 );
buf \U$35074 ( \40768 , \40427 );
buf \U$35075 ( \40769 , \40427 );
buf \U$35076 ( \40770 , \40427 );
buf \U$35077 ( \40771 , \40427 );
buf \U$35078 ( \40772 , \40427 );
buf \U$35079 ( \40773 , \40427 );
buf \U$35080 ( \40774 , \40427 );
buf \U$35081 ( \40775 , \40427 );
buf \U$35082 ( \40776 , \40427 );
buf \U$35083 ( \40777 , \40427 );
buf \U$35084 ( \40778 , \40427 );
buf \U$35085 ( \40779 , \40427 );
buf \U$35086 ( \40780 , \40427 );
buf \U$35087 ( \40781 , \40427 );
buf \U$35088 ( \40782 , \40427 );
buf \U$35089 ( \40783 , \40427 );
buf \U$35090 ( \40784 , \40427 );
buf \U$35091 ( \40785 , \40427 );
buf \U$35092 ( \40786 , \40427 );
buf \U$35093 ( \40787 , \40427 );
buf \U$35094 ( \40788 , \40427 );
buf \U$35095 ( \40789 , \40427 );
nor \U$35096 ( \40790 , \40414 , \40417 , \40419 , \40422 , \40426 , \40427 , \40764 , \40765 , \40766 , \40767 , \40768 , \40769 , \40770 , \40771 , \40772 , \40773 , \40774 , \40775 , \40776 , \40777 , \40778 , \40779 , \40780 , \40781 , \40782 , \40783 , \40784 , \40785 , \40786 , \40787 , \40788 , \40789 );
and \U$35097 ( \40791 , RIeacfa18_6902, \40790 );
buf \U$35098 ( \40792 , \40427 );
buf \U$35099 ( \40793 , \40427 );
buf \U$35100 ( \40794 , \40427 );
buf \U$35101 ( \40795 , \40427 );
buf \U$35102 ( \40796 , \40427 );
buf \U$35103 ( \40797 , \40427 );
buf \U$35104 ( \40798 , \40427 );
buf \U$35105 ( \40799 , \40427 );
buf \U$35106 ( \40800 , \40427 );
buf \U$35107 ( \40801 , \40427 );
buf \U$35108 ( \40802 , \40427 );
buf \U$35109 ( \40803 , \40427 );
buf \U$35110 ( \40804 , \40427 );
buf \U$35111 ( \40805 , \40427 );
buf \U$35112 ( \40806 , \40427 );
buf \U$35113 ( \40807 , \40427 );
buf \U$35114 ( \40808 , \40427 );
buf \U$35115 ( \40809 , \40427 );
buf \U$35116 ( \40810 , \40427 );
buf \U$35117 ( \40811 , \40427 );
buf \U$35118 ( \40812 , \40427 );
buf \U$35119 ( \40813 , \40427 );
buf \U$35120 ( \40814 , \40427 );
buf \U$35121 ( \40815 , \40427 );
buf \U$35122 ( \40816 , \40427 );
buf \U$35123 ( \40817 , \40427 );
nor \U$35124 ( \40818 , \40413 , \40417 , \40419 , \40422 , \40426 , \40427 , \40792 , \40793 , \40794 , \40795 , \40796 , \40797 , \40798 , \40799 , \40800 , \40801 , \40802 , \40803 , \40804 , \40805 , \40806 , \40807 , \40808 , \40809 , \40810 , \40811 , \40812 , \40813 , \40814 , \40815 , \40816 , \40817 );
and \U$35125 ( \40819 , RIeab6518_6891, \40818 );
buf \U$35126 ( \40820 , \40427 );
buf \U$35127 ( \40821 , \40427 );
buf \U$35128 ( \40822 , \40427 );
buf \U$35129 ( \40823 , \40427 );
buf \U$35130 ( \40824 , \40427 );
buf \U$35131 ( \40825 , \40427 );
buf \U$35132 ( \40826 , \40427 );
buf \U$35133 ( \40827 , \40427 );
buf \U$35134 ( \40828 , \40427 );
buf \U$35135 ( \40829 , \40427 );
buf \U$35136 ( \40830 , \40427 );
buf \U$35137 ( \40831 , \40427 );
buf \U$35138 ( \40832 , \40427 );
buf \U$35139 ( \40833 , \40427 );
buf \U$35140 ( \40834 , \40427 );
buf \U$35141 ( \40835 , \40427 );
buf \U$35142 ( \40836 , \40427 );
buf \U$35143 ( \40837 , \40427 );
buf \U$35144 ( \40838 , \40427 );
buf \U$35145 ( \40839 , \40427 );
buf \U$35146 ( \40840 , \40427 );
buf \U$35147 ( \40841 , \40427 );
buf \U$35148 ( \40842 , \40427 );
buf \U$35149 ( \40843 , \40427 );
buf \U$35150 ( \40844 , \40427 );
buf \U$35151 ( \40845 , \40427 );
nor \U$35152 ( \40846 , \40414 , \40416 , \40419 , \40422 , \40426 , \40427 , \40820 , \40821 , \40822 , \40823 , \40824 , \40825 , \40826 , \40827 , \40828 , \40829 , \40830 , \40831 , \40832 , \40833 , \40834 , \40835 , \40836 , \40837 , \40838 , \40839 , \40840 , \40841 , \40842 , \40843 , \40844 , \40845 );
and \U$35153 ( \40847 , RIeb352c8_6904, \40846 );
or \U$35154 ( \40848 , 1'b0 , \40455 , \40483 , \40511 , \40539 , \40567 , \40595 , \40623 , \40651 , \40679 , \40707 , \40735 , \40763 , \40791 , \40819 , \40847 );
buf \U$35155 ( \40849 , \40427 );
not \U$35156 ( \40850 , \40849 );
buf \U$35157 ( \40851 , \40416 );
buf \U$35158 ( \40852 , \40419 );
buf \U$35159 ( \40853 , \40422 );
buf \U$35160 ( \40854 , \40426 );
buf \U$35161 ( \40855 , \40427 );
buf \U$35162 ( \40856 , \40427 );
buf \U$35163 ( \40857 , \40427 );
buf \U$35164 ( \40858 , \40427 );
buf \U$35165 ( \40859 , \40427 );
buf \U$35166 ( \40860 , \40427 );
buf \U$35167 ( \40861 , \40427 );
buf \U$35168 ( \40862 , \40427 );
buf \U$35169 ( \40863 , \40427 );
buf \U$35170 ( \40864 , \40427 );
buf \U$35171 ( \40865 , \40427 );
buf \U$35172 ( \40866 , \40427 );
buf \U$35173 ( \40867 , \40427 );
buf \U$35174 ( \40868 , \40427 );
buf \U$35175 ( \40869 , \40427 );
buf \U$35176 ( \40870 , \40427 );
buf \U$35177 ( \40871 , \40427 );
buf \U$35178 ( \40872 , \40427 );
buf \U$35179 ( \40873 , \40427 );
buf \U$35180 ( \40874 , \40427 );
buf \U$35181 ( \40875 , \40427 );
buf \U$35182 ( \40876 , \40427 );
buf \U$35183 ( \40877 , \40427 );
buf \U$35184 ( \40878 , \40427 );
buf \U$35185 ( \40879 , \40427 );
buf \U$35186 ( \40880 , \40427 );
buf \U$35187 ( \40881 , \40413 );
or \U$35188 ( \40882 , \40851 , \40852 , \40853 , \40854 , \40855 , \40856 , \40857 , \40858 , \40859 , \40860 , \40861 , \40862 , \40863 , \40864 , \40865 , \40866 , \40867 , \40868 , \40869 , \40870 , \40871 , \40872 , \40873 , \40874 , \40875 , \40876 , \40877 , \40878 , \40879 , \40880 , \40881 );
nand \U$35189 ( \40883 , \40850 , \40882 );
buf \U$35190 ( \40884 , \40883 );
or \U$35192 ( \40885 , \40884 , 1'b0 );
_DC gb6e9 ( \40886_nGb6e9 , \40848 , \40885 );
not \U$35193 ( \40887 , \40886_nGb6e9 );
buf \U$35194 ( \40888 , RIb7b9608_246);
buf \U$35196 ( \40889 , \40427 );
buf \U$35197 ( \40890 , \40427 );
buf \U$35198 ( \40891 , \40427 );
buf \U$35199 ( \40892 , \40427 );
buf \U$35200 ( \40893 , \40427 );
buf \U$35201 ( \40894 , \40427 );
buf \U$35202 ( \40895 , \40427 );
buf \U$35203 ( \40896 , \40427 );
buf \U$35204 ( \40897 , \40427 );
buf \U$35205 ( \40898 , \40427 );
buf \U$35206 ( \40899 , \40427 );
buf \U$35207 ( \40900 , \40427 );
buf \U$35208 ( \40901 , \40427 );
buf \U$35209 ( \40902 , \40427 );
buf \U$35210 ( \40903 , \40427 );
buf \U$35211 ( \40904 , \40427 );
buf \U$35212 ( \40905 , \40427 );
buf \U$35213 ( \40906 , \40427 );
buf \U$35214 ( \40907 , \40427 );
buf \U$35215 ( \40908 , \40427 );
buf \U$35216 ( \40909 , \40427 );
buf \U$35217 ( \40910 , \40427 );
buf \U$35218 ( \40911 , \40427 );
buf \U$35219 ( \40912 , \40427 );
buf \U$35220 ( \40913 , \40427 );
buf \U$35221 ( \40914 , \40427 );
nor \U$35222 ( \40915 , \40414 , \40417 , \40420 , \40423 , \40426 , \40427 , \40889 , \40890 , \40891 , \40892 , \40893 , \40894 , \40895 , \40896 , \40897 , \40898 , \40899 , \40900 , \40901 , \40902 , \40903 , \40904 , \40905 , \40906 , \40907 , \40908 , \40909 , \40910 , \40911 , \40912 , \40913 , \40914 );
and \U$35223 ( \40916 , \7119 , \40915 );
buf \U$35224 ( \40917 , \40427 );
buf \U$35225 ( \40918 , \40427 );
buf \U$35226 ( \40919 , \40427 );
buf \U$35227 ( \40920 , \40427 );
buf \U$35228 ( \40921 , \40427 );
buf \U$35229 ( \40922 , \40427 );
buf \U$35230 ( \40923 , \40427 );
buf \U$35231 ( \40924 , \40427 );
buf \U$35232 ( \40925 , \40427 );
buf \U$35233 ( \40926 , \40427 );
buf \U$35234 ( \40927 , \40427 );
buf \U$35235 ( \40928 , \40427 );
buf \U$35236 ( \40929 , \40427 );
buf \U$35237 ( \40930 , \40427 );
buf \U$35238 ( \40931 , \40427 );
buf \U$35239 ( \40932 , \40427 );
buf \U$35240 ( \40933 , \40427 );
buf \U$35241 ( \40934 , \40427 );
buf \U$35242 ( \40935 , \40427 );
buf \U$35243 ( \40936 , \40427 );
buf \U$35244 ( \40937 , \40427 );
buf \U$35245 ( \40938 , \40427 );
buf \U$35246 ( \40939 , \40427 );
buf \U$35247 ( \40940 , \40427 );
buf \U$35248 ( \40941 , \40427 );
buf \U$35249 ( \40942 , \40427 );
nor \U$35250 ( \40943 , \40413 , \40417 , \40420 , \40423 , \40426 , \40427 , \40917 , \40918 , \40919 , \40920 , \40921 , \40922 , \40923 , \40924 , \40925 , \40926 , \40927 , \40928 , \40929 , \40930 , \40931 , \40932 , \40933 , \40934 , \40935 , \40936 , \40937 , \40938 , \40939 , \40940 , \40941 , \40942 );
and \U$35251 ( \40944 , \7864 , \40943 );
buf \U$35252 ( \40945 , \40427 );
buf \U$35253 ( \40946 , \40427 );
buf \U$35254 ( \40947 , \40427 );
buf \U$35255 ( \40948 , \40427 );
buf \U$35256 ( \40949 , \40427 );
buf \U$35257 ( \40950 , \40427 );
buf \U$35258 ( \40951 , \40427 );
buf \U$35259 ( \40952 , \40427 );
buf \U$35260 ( \40953 , \40427 );
buf \U$35261 ( \40954 , \40427 );
buf \U$35262 ( \40955 , \40427 );
buf \U$35263 ( \40956 , \40427 );
buf \U$35264 ( \40957 , \40427 );
buf \U$35265 ( \40958 , \40427 );
buf \U$35266 ( \40959 , \40427 );
buf \U$35267 ( \40960 , \40427 );
buf \U$35268 ( \40961 , \40427 );
buf \U$35269 ( \40962 , \40427 );
buf \U$35270 ( \40963 , \40427 );
buf \U$35271 ( \40964 , \40427 );
buf \U$35272 ( \40965 , \40427 );
buf \U$35273 ( \40966 , \40427 );
buf \U$35274 ( \40967 , \40427 );
buf \U$35275 ( \40968 , \40427 );
buf \U$35276 ( \40969 , \40427 );
buf \U$35277 ( \40970 , \40427 );
nor \U$35278 ( \40971 , \40414 , \40416 , \40420 , \40423 , \40426 , \40427 , \40945 , \40946 , \40947 , \40948 , \40949 , \40950 , \40951 , \40952 , \40953 , \40954 , \40955 , \40956 , \40957 , \40958 , \40959 , \40960 , \40961 , \40962 , \40963 , \40964 , \40965 , \40966 , \40967 , \40968 , \40969 , \40970 );
and \U$35279 ( \40972 , \7892 , \40971 );
buf \U$35280 ( \40973 , \40427 );
buf \U$35281 ( \40974 , \40427 );
buf \U$35282 ( \40975 , \40427 );
buf \U$35283 ( \40976 , \40427 );
buf \U$35284 ( \40977 , \40427 );
buf \U$35285 ( \40978 , \40427 );
buf \U$35286 ( \40979 , \40427 );
buf \U$35287 ( \40980 , \40427 );
buf \U$35288 ( \40981 , \40427 );
buf \U$35289 ( \40982 , \40427 );
buf \U$35290 ( \40983 , \40427 );
buf \U$35291 ( \40984 , \40427 );
buf \U$35292 ( \40985 , \40427 );
buf \U$35293 ( \40986 , \40427 );
buf \U$35294 ( \40987 , \40427 );
buf \U$35295 ( \40988 , \40427 );
buf \U$35296 ( \40989 , \40427 );
buf \U$35297 ( \40990 , \40427 );
buf \U$35298 ( \40991 , \40427 );
buf \U$35299 ( \40992 , \40427 );
buf \U$35300 ( \40993 , \40427 );
buf \U$35301 ( \40994 , \40427 );
buf \U$35302 ( \40995 , \40427 );
buf \U$35303 ( \40996 , \40427 );
buf \U$35304 ( \40997 , \40427 );
buf \U$35305 ( \40998 , \40427 );
nor \U$35306 ( \40999 , \40413 , \40416 , \40420 , \40423 , \40426 , \40427 , \40973 , \40974 , \40975 , \40976 , \40977 , \40978 , \40979 , \40980 , \40981 , \40982 , \40983 , \40984 , \40985 , \40986 , \40987 , \40988 , \40989 , \40990 , \40991 , \40992 , \40993 , \40994 , \40995 , \40996 , \40997 , \40998 );
and \U$35307 ( \41000 , \7920 , \40999 );
buf \U$35308 ( \41001 , \40427 );
buf \U$35309 ( \41002 , \40427 );
buf \U$35310 ( \41003 , \40427 );
buf \U$35311 ( \41004 , \40427 );
buf \U$35312 ( \41005 , \40427 );
buf \U$35313 ( \41006 , \40427 );
buf \U$35314 ( \41007 , \40427 );
buf \U$35315 ( \41008 , \40427 );
buf \U$35316 ( \41009 , \40427 );
buf \U$35317 ( \41010 , \40427 );
buf \U$35318 ( \41011 , \40427 );
buf \U$35319 ( \41012 , \40427 );
buf \U$35320 ( \41013 , \40427 );
buf \U$35321 ( \41014 , \40427 );
buf \U$35322 ( \41015 , \40427 );
buf \U$35323 ( \41016 , \40427 );
buf \U$35324 ( \41017 , \40427 );
buf \U$35325 ( \41018 , \40427 );
buf \U$35326 ( \41019 , \40427 );
buf \U$35327 ( \41020 , \40427 );
buf \U$35328 ( \41021 , \40427 );
buf \U$35329 ( \41022 , \40427 );
buf \U$35330 ( \41023 , \40427 );
buf \U$35331 ( \41024 , \40427 );
buf \U$35332 ( \41025 , \40427 );
buf \U$35333 ( \41026 , \40427 );
nor \U$35334 ( \41027 , \40414 , \40417 , \40419 , \40423 , \40426 , \40427 , \41001 , \41002 , \41003 , \41004 , \41005 , \41006 , \41007 , \41008 , \41009 , \41010 , \41011 , \41012 , \41013 , \41014 , \41015 , \41016 , \41017 , \41018 , \41019 , \41020 , \41021 , \41022 , \41023 , \41024 , \41025 , \41026 );
and \U$35335 ( \41028 , \7948 , \41027 );
buf \U$35336 ( \41029 , \40427 );
buf \U$35337 ( \41030 , \40427 );
buf \U$35338 ( \41031 , \40427 );
buf \U$35339 ( \41032 , \40427 );
buf \U$35340 ( \41033 , \40427 );
buf \U$35341 ( \41034 , \40427 );
buf \U$35342 ( \41035 , \40427 );
buf \U$35343 ( \41036 , \40427 );
buf \U$35344 ( \41037 , \40427 );
buf \U$35345 ( \41038 , \40427 );
buf \U$35346 ( \41039 , \40427 );
buf \U$35347 ( \41040 , \40427 );
buf \U$35348 ( \41041 , \40427 );
buf \U$35349 ( \41042 , \40427 );
buf \U$35350 ( \41043 , \40427 );
buf \U$35351 ( \41044 , \40427 );
buf \U$35352 ( \41045 , \40427 );
buf \U$35353 ( \41046 , \40427 );
buf \U$35354 ( \41047 , \40427 );
buf \U$35355 ( \41048 , \40427 );
buf \U$35356 ( \41049 , \40427 );
buf \U$35357 ( \41050 , \40427 );
buf \U$35358 ( \41051 , \40427 );
buf \U$35359 ( \41052 , \40427 );
buf \U$35360 ( \41053 , \40427 );
buf \U$35361 ( \41054 , \40427 );
nor \U$35362 ( \41055 , \40413 , \40417 , \40419 , \40423 , \40426 , \40427 , \41029 , \41030 , \41031 , \41032 , \41033 , \41034 , \41035 , \41036 , \41037 , \41038 , \41039 , \41040 , \41041 , \41042 , \41043 , \41044 , \41045 , \41046 , \41047 , \41048 , \41049 , \41050 , \41051 , \41052 , \41053 , \41054 );
and \U$35363 ( \41056 , \7976 , \41055 );
buf \U$35364 ( \41057 , \40427 );
buf \U$35365 ( \41058 , \40427 );
buf \U$35366 ( \41059 , \40427 );
buf \U$35367 ( \41060 , \40427 );
buf \U$35368 ( \41061 , \40427 );
buf \U$35369 ( \41062 , \40427 );
buf \U$35370 ( \41063 , \40427 );
buf \U$35371 ( \41064 , \40427 );
buf \U$35372 ( \41065 , \40427 );
buf \U$35373 ( \41066 , \40427 );
buf \U$35374 ( \41067 , \40427 );
buf \U$35375 ( \41068 , \40427 );
buf \U$35376 ( \41069 , \40427 );
buf \U$35377 ( \41070 , \40427 );
buf \U$35378 ( \41071 , \40427 );
buf \U$35379 ( \41072 , \40427 );
buf \U$35380 ( \41073 , \40427 );
buf \U$35381 ( \41074 , \40427 );
buf \U$35382 ( \41075 , \40427 );
buf \U$35383 ( \41076 , \40427 );
buf \U$35384 ( \41077 , \40427 );
buf \U$35385 ( \41078 , \40427 );
buf \U$35386 ( \41079 , \40427 );
buf \U$35387 ( \41080 , \40427 );
buf \U$35388 ( \41081 , \40427 );
buf \U$35389 ( \41082 , \40427 );
nor \U$35390 ( \41083 , \40414 , \40416 , \40419 , \40423 , \40426 , \40427 , \41057 , \41058 , \41059 , \41060 , \41061 , \41062 , \41063 , \41064 , \41065 , \41066 , \41067 , \41068 , \41069 , \41070 , \41071 , \41072 , \41073 , \41074 , \41075 , \41076 , \41077 , \41078 , \41079 , \41080 , \41081 , \41082 );
and \U$35391 ( \41084 , \8004 , \41083 );
buf \U$35392 ( \41085 , \40427 );
buf \U$35393 ( \41086 , \40427 );
buf \U$35394 ( \41087 , \40427 );
buf \U$35395 ( \41088 , \40427 );
buf \U$35396 ( \41089 , \40427 );
buf \U$35397 ( \41090 , \40427 );
buf \U$35398 ( \41091 , \40427 );
buf \U$35399 ( \41092 , \40427 );
buf \U$35400 ( \41093 , \40427 );
buf \U$35401 ( \41094 , \40427 );
buf \U$35402 ( \41095 , \40427 );
buf \U$35403 ( \41096 , \40427 );
buf \U$35404 ( \41097 , \40427 );
buf \U$35405 ( \41098 , \40427 );
buf \U$35406 ( \41099 , \40427 );
buf \U$35407 ( \41100 , \40427 );
buf \U$35408 ( \41101 , \40427 );
buf \U$35409 ( \41102 , \40427 );
buf \U$35410 ( \41103 , \40427 );
buf \U$35411 ( \41104 , \40427 );
buf \U$35412 ( \41105 , \40427 );
buf \U$35413 ( \41106 , \40427 );
buf \U$35414 ( \41107 , \40427 );
buf \U$35415 ( \41108 , \40427 );
buf \U$35416 ( \41109 , \40427 );
buf \U$35417 ( \41110 , \40427 );
nor \U$35418 ( \41111 , \40413 , \40416 , \40419 , \40423 , \40426 , \40427 , \41085 , \41086 , \41087 , \41088 , \41089 , \41090 , \41091 , \41092 , \41093 , \41094 , \41095 , \41096 , \41097 , \41098 , \41099 , \41100 , \41101 , \41102 , \41103 , \41104 , \41105 , \41106 , \41107 , \41108 , \41109 , \41110 );
and \U$35419 ( \41112 , \8032 , \41111 );
buf \U$35420 ( \41113 , \40427 );
buf \U$35421 ( \41114 , \40427 );
buf \U$35422 ( \41115 , \40427 );
buf \U$35423 ( \41116 , \40427 );
buf \U$35424 ( \41117 , \40427 );
buf \U$35425 ( \41118 , \40427 );
buf \U$35426 ( \41119 , \40427 );
buf \U$35427 ( \41120 , \40427 );
buf \U$35428 ( \41121 , \40427 );
buf \U$35429 ( \41122 , \40427 );
buf \U$35430 ( \41123 , \40427 );
buf \U$35431 ( \41124 , \40427 );
buf \U$35432 ( \41125 , \40427 );
buf \U$35433 ( \41126 , \40427 );
buf \U$35434 ( \41127 , \40427 );
buf \U$35435 ( \41128 , \40427 );
buf \U$35436 ( \41129 , \40427 );
buf \U$35437 ( \41130 , \40427 );
buf \U$35438 ( \41131 , \40427 );
buf \U$35439 ( \41132 , \40427 );
buf \U$35440 ( \41133 , \40427 );
buf \U$35441 ( \41134 , \40427 );
buf \U$35442 ( \41135 , \40427 );
buf \U$35443 ( \41136 , \40427 );
buf \U$35444 ( \41137 , \40427 );
buf \U$35445 ( \41138 , \40427 );
nor \U$35446 ( \41139 , \40414 , \40417 , \40420 , \40422 , \40426 , \40427 , \41113 , \41114 , \41115 , \41116 , \41117 , \41118 , \41119 , \41120 , \41121 , \41122 , \41123 , \41124 , \41125 , \41126 , \41127 , \41128 , \41129 , \41130 , \41131 , \41132 , \41133 , \41134 , \41135 , \41136 , \41137 , \41138 );
and \U$35447 ( \41140 , \8060 , \41139 );
buf \U$35448 ( \41141 , \40427 );
buf \U$35449 ( \41142 , \40427 );
buf \U$35450 ( \41143 , \40427 );
buf \U$35451 ( \41144 , \40427 );
buf \U$35452 ( \41145 , \40427 );
buf \U$35453 ( \41146 , \40427 );
buf \U$35454 ( \41147 , \40427 );
buf \U$35455 ( \41148 , \40427 );
buf \U$35456 ( \41149 , \40427 );
buf \U$35457 ( \41150 , \40427 );
buf \U$35458 ( \41151 , \40427 );
buf \U$35459 ( \41152 , \40427 );
buf \U$35460 ( \41153 , \40427 );
buf \U$35461 ( \41154 , \40427 );
buf \U$35462 ( \41155 , \40427 );
buf \U$35463 ( \41156 , \40427 );
buf \U$35464 ( \41157 , \40427 );
buf \U$35465 ( \41158 , \40427 );
buf \U$35466 ( \41159 , \40427 );
buf \U$35467 ( \41160 , \40427 );
buf \U$35468 ( \41161 , \40427 );
buf \U$35469 ( \41162 , \40427 );
buf \U$35470 ( \41163 , \40427 );
buf \U$35471 ( \41164 , \40427 );
buf \U$35472 ( \41165 , \40427 );
buf \U$35473 ( \41166 , \40427 );
nor \U$35474 ( \41167 , \40413 , \40417 , \40420 , \40422 , \40426 , \40427 , \41141 , \41142 , \41143 , \41144 , \41145 , \41146 , \41147 , \41148 , \41149 , \41150 , \41151 , \41152 , \41153 , \41154 , \41155 , \41156 , \41157 , \41158 , \41159 , \41160 , \41161 , \41162 , \41163 , \41164 , \41165 , \41166 );
and \U$35475 ( \41168 , \8088 , \41167 );
buf \U$35476 ( \41169 , \40427 );
buf \U$35477 ( \41170 , \40427 );
buf \U$35478 ( \41171 , \40427 );
buf \U$35479 ( \41172 , \40427 );
buf \U$35480 ( \41173 , \40427 );
buf \U$35481 ( \41174 , \40427 );
buf \U$35482 ( \41175 , \40427 );
buf \U$35483 ( \41176 , \40427 );
buf \U$35484 ( \41177 , \40427 );
buf \U$35485 ( \41178 , \40427 );
buf \U$35486 ( \41179 , \40427 );
buf \U$35487 ( \41180 , \40427 );
buf \U$35488 ( \41181 , \40427 );
buf \U$35489 ( \41182 , \40427 );
buf \U$35490 ( \41183 , \40427 );
buf \U$35491 ( \41184 , \40427 );
buf \U$35492 ( \41185 , \40427 );
buf \U$35493 ( \41186 , \40427 );
buf \U$35494 ( \41187 , \40427 );
buf \U$35495 ( \41188 , \40427 );
buf \U$35496 ( \41189 , \40427 );
buf \U$35497 ( \41190 , \40427 );
buf \U$35498 ( \41191 , \40427 );
buf \U$35499 ( \41192 , \40427 );
buf \U$35500 ( \41193 , \40427 );
buf \U$35501 ( \41194 , \40427 );
nor \U$35502 ( \41195 , \40414 , \40416 , \40420 , \40422 , \40426 , \40427 , \41169 , \41170 , \41171 , \41172 , \41173 , \41174 , \41175 , \41176 , \41177 , \41178 , \41179 , \41180 , \41181 , \41182 , \41183 , \41184 , \41185 , \41186 , \41187 , \41188 , \41189 , \41190 , \41191 , \41192 , \41193 , \41194 );
and \U$35503 ( \41196 , \8116 , \41195 );
buf \U$35504 ( \41197 , \40427 );
buf \U$35505 ( \41198 , \40427 );
buf \U$35506 ( \41199 , \40427 );
buf \U$35507 ( \41200 , \40427 );
buf \U$35508 ( \41201 , \40427 );
buf \U$35509 ( \41202 , \40427 );
buf \U$35510 ( \41203 , \40427 );
buf \U$35511 ( \41204 , \40427 );
buf \U$35512 ( \41205 , \40427 );
buf \U$35513 ( \41206 , \40427 );
buf \U$35514 ( \41207 , \40427 );
buf \U$35515 ( \41208 , \40427 );
buf \U$35516 ( \41209 , \40427 );
buf \U$35517 ( \41210 , \40427 );
buf \U$35518 ( \41211 , \40427 );
buf \U$35519 ( \41212 , \40427 );
buf \U$35520 ( \41213 , \40427 );
buf \U$35521 ( \41214 , \40427 );
buf \U$35522 ( \41215 , \40427 );
buf \U$35523 ( \41216 , \40427 );
buf \U$35524 ( \41217 , \40427 );
buf \U$35525 ( \41218 , \40427 );
buf \U$35526 ( \41219 , \40427 );
buf \U$35527 ( \41220 , \40427 );
buf \U$35528 ( \41221 , \40427 );
buf \U$35529 ( \41222 , \40427 );
nor \U$35530 ( \41223 , \40413 , \40416 , \40420 , \40422 , \40426 , \40427 , \41197 , \41198 , \41199 , \41200 , \41201 , \41202 , \41203 , \41204 , \41205 , \41206 , \41207 , \41208 , \41209 , \41210 , \41211 , \41212 , \41213 , \41214 , \41215 , \41216 , \41217 , \41218 , \41219 , \41220 , \41221 , \41222 );
and \U$35531 ( \41224 , \8144 , \41223 );
buf \U$35532 ( \41225 , \40427 );
buf \U$35533 ( \41226 , \40427 );
buf \U$35534 ( \41227 , \40427 );
buf \U$35535 ( \41228 , \40427 );
buf \U$35536 ( \41229 , \40427 );
buf \U$35537 ( \41230 , \40427 );
buf \U$35538 ( \41231 , \40427 );
buf \U$35539 ( \41232 , \40427 );
buf \U$35540 ( \41233 , \40427 );
buf \U$35541 ( \41234 , \40427 );
buf \U$35542 ( \41235 , \40427 );
buf \U$35543 ( \41236 , \40427 );
buf \U$35544 ( \41237 , \40427 );
buf \U$35545 ( \41238 , \40427 );
buf \U$35546 ( \41239 , \40427 );
buf \U$35547 ( \41240 , \40427 );
buf \U$35548 ( \41241 , \40427 );
buf \U$35549 ( \41242 , \40427 );
buf \U$35550 ( \41243 , \40427 );
buf \U$35551 ( \41244 , \40427 );
buf \U$35552 ( \41245 , \40427 );
buf \U$35553 ( \41246 , \40427 );
buf \U$35554 ( \41247 , \40427 );
buf \U$35555 ( \41248 , \40427 );
buf \U$35556 ( \41249 , \40427 );
buf \U$35557 ( \41250 , \40427 );
nor \U$35558 ( \41251 , \40414 , \40417 , \40419 , \40422 , \40426 , \40427 , \41225 , \41226 , \41227 , \41228 , \41229 , \41230 , \41231 , \41232 , \41233 , \41234 , \41235 , \41236 , \41237 , \41238 , \41239 , \41240 , \41241 , \41242 , \41243 , \41244 , \41245 , \41246 , \41247 , \41248 , \41249 , \41250 );
and \U$35559 ( \41252 , \8172 , \41251 );
buf \U$35560 ( \41253 , \40427 );
buf \U$35561 ( \41254 , \40427 );
buf \U$35562 ( \41255 , \40427 );
buf \U$35563 ( \41256 , \40427 );
buf \U$35564 ( \41257 , \40427 );
buf \U$35565 ( \41258 , \40427 );
buf \U$35566 ( \41259 , \40427 );
buf \U$35567 ( \41260 , \40427 );
buf \U$35568 ( \41261 , \40427 );
buf \U$35569 ( \41262 , \40427 );
buf \U$35570 ( \41263 , \40427 );
buf \U$35571 ( \41264 , \40427 );
buf \U$35572 ( \41265 , \40427 );
buf \U$35573 ( \41266 , \40427 );
buf \U$35574 ( \41267 , \40427 );
buf \U$35575 ( \41268 , \40427 );
buf \U$35576 ( \41269 , \40427 );
buf \U$35577 ( \41270 , \40427 );
buf \U$35578 ( \41271 , \40427 );
buf \U$35579 ( \41272 , \40427 );
buf \U$35580 ( \41273 , \40427 );
buf \U$35581 ( \41274 , \40427 );
buf \U$35582 ( \41275 , \40427 );
buf \U$35583 ( \41276 , \40427 );
buf \U$35584 ( \41277 , \40427 );
buf \U$35585 ( \41278 , \40427 );
nor \U$35586 ( \41279 , \40413 , \40417 , \40419 , \40422 , \40426 , \40427 , \41253 , \41254 , \41255 , \41256 , \41257 , \41258 , \41259 , \41260 , \41261 , \41262 , \41263 , \41264 , \41265 , \41266 , \41267 , \41268 , \41269 , \41270 , \41271 , \41272 , \41273 , \41274 , \41275 , \41276 , \41277 , \41278 );
and \U$35587 ( \41280 , \8200 , \41279 );
buf \U$35588 ( \41281 , \40427 );
buf \U$35589 ( \41282 , \40427 );
buf \U$35590 ( \41283 , \40427 );
buf \U$35591 ( \41284 , \40427 );
buf \U$35592 ( \41285 , \40427 );
buf \U$35593 ( \41286 , \40427 );
buf \U$35594 ( \41287 , \40427 );
buf \U$35595 ( \41288 , \40427 );
buf \U$35596 ( \41289 , \40427 );
buf \U$35597 ( \41290 , \40427 );
buf \U$35598 ( \41291 , \40427 );
buf \U$35599 ( \41292 , \40427 );
buf \U$35600 ( \41293 , \40427 );
buf \U$35601 ( \41294 , \40427 );
buf \U$35602 ( \41295 , \40427 );
buf \U$35603 ( \41296 , \40427 );
buf \U$35604 ( \41297 , \40427 );
buf \U$35605 ( \41298 , \40427 );
buf \U$35606 ( \41299 , \40427 );
buf \U$35607 ( \41300 , \40427 );
buf \U$35608 ( \41301 , \40427 );
buf \U$35609 ( \41302 , \40427 );
buf \U$35610 ( \41303 , \40427 );
buf \U$35611 ( \41304 , \40427 );
buf \U$35612 ( \41305 , \40427 );
buf \U$35613 ( \41306 , \40427 );
nor \U$35614 ( \41307 , \40414 , \40416 , \40419 , \40422 , \40426 , \40427 , \41281 , \41282 , \41283 , \41284 , \41285 , \41286 , \41287 , \41288 , \41289 , \41290 , \41291 , \41292 , \41293 , \41294 , \41295 , \41296 , \41297 , \41298 , \41299 , \41300 , \41301 , \41302 , \41303 , \41304 , \41305 , \41306 );
and \U$35615 ( \41308 , \8228 , \41307 );
or \U$35616 ( \41309 , 1'b0 , \40916 , \40944 , \40972 , \41000 , \41028 , \41056 , \41084 , \41112 , \41140 , \41168 , \41196 , \41224 , \41252 , \41280 , \41308 );
buf \U$35617 ( \41310 , \40427 );
not \U$35618 ( \41311 , \41310 );
buf \U$35619 ( \41312 , \40416 );
buf \U$35620 ( \41313 , \40419 );
buf \U$35621 ( \41314 , \40422 );
buf \U$35622 ( \41315 , \40426 );
buf \U$35623 ( \41316 , \40427 );
buf \U$35624 ( \41317 , \40427 );
buf \U$35625 ( \41318 , \40427 );
buf \U$35626 ( \41319 , \40427 );
buf \U$35627 ( \41320 , \40427 );
buf \U$35628 ( \41321 , \40427 );
buf \U$35629 ( \41322 , \40427 );
buf \U$35630 ( \41323 , \40427 );
buf \U$35631 ( \41324 , \40427 );
buf \U$35632 ( \41325 , \40427 );
buf \U$35633 ( \41326 , \40427 );
buf \U$35634 ( \41327 , \40427 );
buf \U$35635 ( \41328 , \40427 );
buf \U$35636 ( \41329 , \40427 );
buf \U$35637 ( \41330 , \40427 );
buf \U$35638 ( \41331 , \40427 );
buf \U$35639 ( \41332 , \40427 );
buf \U$35640 ( \41333 , \40427 );
buf \U$35641 ( \41334 , \40427 );
buf \U$35642 ( \41335 , \40427 );
buf \U$35643 ( \41336 , \40427 );
buf \U$35644 ( \41337 , \40427 );
buf \U$35645 ( \41338 , \40427 );
buf \U$35646 ( \41339 , \40427 );
buf \U$35647 ( \41340 , \40427 );
buf \U$35648 ( \41341 , \40427 );
buf \U$35649 ( \41342 , \40413 );
or \U$35650 ( \41343 , \41312 , \41313 , \41314 , \41315 , \41316 , \41317 , \41318 , \41319 , \41320 , \41321 , \41322 , \41323 , \41324 , \41325 , \41326 , \41327 , \41328 , \41329 , \41330 , \41331 , \41332 , \41333 , \41334 , \41335 , \41336 , \41337 , \41338 , \41339 , \41340 , \41341 , \41342 );
nand \U$35651 ( \41344 , \41311 , \41343 );
buf \U$35652 ( \41345 , \41344 );
or \U$35654 ( \41346 , \41345 , 1'b0 );
_DC gb8b6 ( \41347_nGb8b6 , \41309 , \41346 );
buf \U$35655 ( \41348 , \41347_nGb8b6 );
xor \U$35656 ( \41349 , \40888 , \41348 );
buf \U$35657 ( \41350 , RIb7b9590_247);
and \U$35659 ( \41351 , \7128 , \40915 );
and \U$35660 ( \41352 , \8338 , \40943 );
and \U$35661 ( \41353 , \8340 , \40971 );
and \U$35662 ( \41354 , \8342 , \40999 );
and \U$35663 ( \41355 , \8344 , \41027 );
and \U$35664 ( \41356 , \8346 , \41055 );
and \U$35665 ( \41357 , \8348 , \41083 );
and \U$35666 ( \41358 , \8350 , \41111 );
and \U$35667 ( \41359 , \8352 , \41139 );
and \U$35668 ( \41360 , \8354 , \41167 );
and \U$35669 ( \41361 , \8356 , \41195 );
and \U$35670 ( \41362 , \8358 , \41223 );
and \U$35671 ( \41363 , \8360 , \41251 );
and \U$35672 ( \41364 , \8362 , \41279 );
and \U$35673 ( \41365 , \8364 , \41307 );
or \U$35674 ( \41366 , 1'b0 , \41351 , \41352 , \41353 , \41354 , \41355 , \41356 , \41357 , \41358 , \41359 , \41360 , \41361 , \41362 , \41363 , \41364 , \41365 );
_DC gb8ca ( \41367_nGb8ca , \41366 , \41346 );
buf \U$35675 ( \41368 , \41367_nGb8ca );
xor \U$35676 ( \41369 , \41350 , \41368 );
or \U$35677 ( \41370 , \41349 , \41369 );
buf \U$35678 ( \41371 , RIb7b9518_248);
and \U$35680 ( \41372 , \7138 , \40915 );
and \U$35681 ( \41373 , \8374 , \40943 );
and \U$35682 ( \41374 , \8376 , \40971 );
and \U$35683 ( \41375 , \8378 , \40999 );
and \U$35684 ( \41376 , \8380 , \41027 );
and \U$35685 ( \41377 , \8382 , \41055 );
and \U$35686 ( \41378 , \8384 , \41083 );
and \U$35687 ( \41379 , \8386 , \41111 );
and \U$35688 ( \41380 , \8388 , \41139 );
and \U$35689 ( \41381 , \8390 , \41167 );
and \U$35690 ( \41382 , \8392 , \41195 );
and \U$35691 ( \41383 , \8394 , \41223 );
and \U$35692 ( \41384 , \8396 , \41251 );
and \U$35693 ( \41385 , \8398 , \41279 );
and \U$35694 ( \41386 , \8400 , \41307 );
or \U$35695 ( \41387 , 1'b0 , \41372 , \41373 , \41374 , \41375 , \41376 , \41377 , \41378 , \41379 , \41380 , \41381 , \41382 , \41383 , \41384 , \41385 , \41386 );
_DC gb8df ( \41388_nGb8df , \41387 , \41346 );
buf \U$35696 ( \41389 , \41388_nGb8df );
xor \U$35697 ( \41390 , \41371 , \41389 );
or \U$35698 ( \41391 , \41370 , \41390 );
buf \U$35699 ( \41392 , RIb7b94a0_249);
and \U$35701 ( \41393 , \7148 , \40915 );
and \U$35702 ( \41394 , \8410 , \40943 );
and \U$35703 ( \41395 , \8412 , \40971 );
and \U$35704 ( \41396 , \8414 , \40999 );
and \U$35705 ( \41397 , \8416 , \41027 );
and \U$35706 ( \41398 , \8418 , \41055 );
and \U$35707 ( \41399 , \8420 , \41083 );
and \U$35708 ( \41400 , \8422 , \41111 );
and \U$35709 ( \41401 , \8424 , \41139 );
and \U$35710 ( \41402 , \8426 , \41167 );
and \U$35711 ( \41403 , \8428 , \41195 );
and \U$35712 ( \41404 , \8430 , \41223 );
and \U$35713 ( \41405 , \8432 , \41251 );
and \U$35714 ( \41406 , \8434 , \41279 );
and \U$35715 ( \41407 , \8436 , \41307 );
or \U$35716 ( \41408 , 1'b0 , \41393 , \41394 , \41395 , \41396 , \41397 , \41398 , \41399 , \41400 , \41401 , \41402 , \41403 , \41404 , \41405 , \41406 , \41407 );
_DC gb8f4 ( \41409_nGb8f4 , \41408 , \41346 );
buf \U$35717 ( \41410 , \41409_nGb8f4 );
xor \U$35718 ( \41411 , \41392 , \41410 );
or \U$35719 ( \41412 , \41391 , \41411 );
buf \U$35720 ( \41413 , RIb7b9428_250);
and \U$35722 ( \41414 , \7158 , \40915 );
and \U$35723 ( \41415 , \8446 , \40943 );
and \U$35724 ( \41416 , \8448 , \40971 );
and \U$35725 ( \41417 , \8450 , \40999 );
and \U$35726 ( \41418 , \8452 , \41027 );
and \U$35727 ( \41419 , \8454 , \41055 );
and \U$35728 ( \41420 , \8456 , \41083 );
and \U$35729 ( \41421 , \8458 , \41111 );
and \U$35730 ( \41422 , \8460 , \41139 );
and \U$35731 ( \41423 , \8462 , \41167 );
and \U$35732 ( \41424 , \8464 , \41195 );
and \U$35733 ( \41425 , \8466 , \41223 );
and \U$35734 ( \41426 , \8468 , \41251 );
and \U$35735 ( \41427 , \8470 , \41279 );
and \U$35736 ( \41428 , \8472 , \41307 );
or \U$35737 ( \41429 , 1'b0 , \41414 , \41415 , \41416 , \41417 , \41418 , \41419 , \41420 , \41421 , \41422 , \41423 , \41424 , \41425 , \41426 , \41427 , \41428 );
_DC gb909 ( \41430_nGb909 , \41429 , \41346 );
buf \U$35738 ( \41431 , \41430_nGb909 );
xor \U$35739 ( \41432 , \41413 , \41431 );
or \U$35740 ( \41433 , \41412 , \41432 );
buf \U$35741 ( \41434 , RIb7b93b0_251);
and \U$35743 ( \41435 , \7168 , \40915 );
and \U$35744 ( \41436 , \8482 , \40943 );
and \U$35745 ( \41437 , \8484 , \40971 );
and \U$35746 ( \41438 , \8486 , \40999 );
and \U$35747 ( \41439 , \8488 , \41027 );
and \U$35748 ( \41440 , \8490 , \41055 );
and \U$35749 ( \41441 , \8492 , \41083 );
and \U$35750 ( \41442 , \8494 , \41111 );
and \U$35751 ( \41443 , \8496 , \41139 );
and \U$35752 ( \41444 , \8498 , \41167 );
and \U$35753 ( \41445 , \8500 , \41195 );
and \U$35754 ( \41446 , \8502 , \41223 );
and \U$35755 ( \41447 , \8504 , \41251 );
and \U$35756 ( \41448 , \8506 , \41279 );
and \U$35757 ( \41449 , \8508 , \41307 );
or \U$35758 ( \41450 , 1'b0 , \41435 , \41436 , \41437 , \41438 , \41439 , \41440 , \41441 , \41442 , \41443 , \41444 , \41445 , \41446 , \41447 , \41448 , \41449 );
_DC gb91e ( \41451_nGb91e , \41450 , \41346 );
buf \U$35759 ( \41452 , \41451_nGb91e );
xor \U$35760 ( \41453 , \41434 , \41452 );
or \U$35761 ( \41454 , \41433 , \41453 );
buf \U$35762 ( \41455 , RIb7af720_252);
and \U$35764 ( \41456 , \7178 , \40915 );
and \U$35765 ( \41457 , \8518 , \40943 );
and \U$35766 ( \41458 , \8520 , \40971 );
and \U$35767 ( \41459 , \8522 , \40999 );
and \U$35768 ( \41460 , \8524 , \41027 );
and \U$35769 ( \41461 , \8526 , \41055 );
and \U$35770 ( \41462 , \8528 , \41083 );
and \U$35771 ( \41463 , \8530 , \41111 );
and \U$35772 ( \41464 , \8532 , \41139 );
and \U$35773 ( \41465 , \8534 , \41167 );
and \U$35774 ( \41466 , \8536 , \41195 );
and \U$35775 ( \41467 , \8538 , \41223 );
and \U$35776 ( \41468 , \8540 , \41251 );
and \U$35777 ( \41469 , \8542 , \41279 );
and \U$35778 ( \41470 , \8544 , \41307 );
or \U$35779 ( \41471 , 1'b0 , \41456 , \41457 , \41458 , \41459 , \41460 , \41461 , \41462 , \41463 , \41464 , \41465 , \41466 , \41467 , \41468 , \41469 , \41470 );
_DC gb933 ( \41472_nGb933 , \41471 , \41346 );
buf \U$35780 ( \41473 , \41472_nGb933 );
xor \U$35781 ( \41474 , \41455 , \41473 );
or \U$35782 ( \41475 , \41454 , \41474 );
buf \U$35783 ( \41476 , RIb7af6a8_253);
and \U$35785 ( \41477 , \7188 , \40915 );
and \U$35786 ( \41478 , \8554 , \40943 );
and \U$35787 ( \41479 , \8556 , \40971 );
and \U$35788 ( \41480 , \8558 , \40999 );
and \U$35789 ( \41481 , \8560 , \41027 );
and \U$35790 ( \41482 , \8562 , \41055 );
and \U$35791 ( \41483 , \8564 , \41083 );
and \U$35792 ( \41484 , \8566 , \41111 );
and \U$35793 ( \41485 , \8568 , \41139 );
and \U$35794 ( \41486 , \8570 , \41167 );
and \U$35795 ( \41487 , \8572 , \41195 );
and \U$35796 ( \41488 , \8574 , \41223 );
and \U$35797 ( \41489 , \8576 , \41251 );
and \U$35798 ( \41490 , \8578 , \41279 );
and \U$35799 ( \41491 , \8580 , \41307 );
or \U$35800 ( \41492 , 1'b0 , \41477 , \41478 , \41479 , \41480 , \41481 , \41482 , \41483 , \41484 , \41485 , \41486 , \41487 , \41488 , \41489 , \41490 , \41491 );
_DC gb948 ( \41493_nGb948 , \41492 , \41346 );
buf \U$35801 ( \41494 , \41493_nGb948 );
xor \U$35802 ( \41495 , \41476 , \41494 );
or \U$35803 ( \41496 , \41475 , \41495 );
not \U$35804 ( \41497 , \41496 );
buf \U$35805 ( \41498 , \41497 );
and \U$35806 ( \41499 , \40887 , \41498 );
buf \U$35807 ( \41500 , RIb7af630_254);
buf \U$35809 ( \41501 , \40427 );
buf \U$35810 ( \41502 , \40427 );
buf \U$35811 ( \41503 , \40427 );
buf \U$35812 ( \41504 , \40427 );
buf \U$35813 ( \41505 , \40427 );
buf \U$35814 ( \41506 , \40427 );
buf \U$35815 ( \41507 , \40427 );
buf \U$35816 ( \41508 , \40427 );
buf \U$35817 ( \41509 , \40427 );
buf \U$35818 ( \41510 , \40427 );
buf \U$35819 ( \41511 , \40427 );
buf \U$35820 ( \41512 , \40427 );
buf \U$35821 ( \41513 , \40427 );
buf \U$35822 ( \41514 , \40427 );
buf \U$35823 ( \41515 , \40427 );
buf \U$35824 ( \41516 , \40427 );
buf \U$35825 ( \41517 , \40427 );
buf \U$35826 ( \41518 , \40427 );
buf \U$35827 ( \41519 , \40427 );
buf \U$35828 ( \41520 , \40427 );
buf \U$35829 ( \41521 , \40427 );
buf \U$35830 ( \41522 , \40427 );
buf \U$35831 ( \41523 , \40427 );
buf \U$35832 ( \41524 , \40427 );
buf \U$35833 ( \41525 , \40427 );
buf \U$35834 ( \41526 , \40427 );
nor \U$35835 ( \41527 , \40414 , \40417 , \40420 , \40423 , \40426 , \40427 , \41501 , \41502 , \41503 , \41504 , \41505 , \41506 , \41507 , \41508 , \41509 , \41510 , \41511 , \41512 , \41513 , \41514 , \41515 , \41516 , \41517 , \41518 , \41519 , \41520 , \41521 , \41522 , \41523 , \41524 , \41525 , \41526 );
and \U$35836 ( \41528 , \7200 , \41527 );
buf \U$35837 ( \41529 , \40427 );
buf \U$35838 ( \41530 , \40427 );
buf \U$35839 ( \41531 , \40427 );
buf \U$35840 ( \41532 , \40427 );
buf \U$35841 ( \41533 , \40427 );
buf \U$35842 ( \41534 , \40427 );
buf \U$35843 ( \41535 , \40427 );
buf \U$35844 ( \41536 , \40427 );
buf \U$35845 ( \41537 , \40427 );
buf \U$35846 ( \41538 , \40427 );
buf \U$35847 ( \41539 , \40427 );
buf \U$35848 ( \41540 , \40427 );
buf \U$35849 ( \41541 , \40427 );
buf \U$35850 ( \41542 , \40427 );
buf \U$35851 ( \41543 , \40427 );
buf \U$35852 ( \41544 , \40427 );
buf \U$35853 ( \41545 , \40427 );
buf \U$35854 ( \41546 , \40427 );
buf \U$35855 ( \41547 , \40427 );
buf \U$35856 ( \41548 , \40427 );
buf \U$35857 ( \41549 , \40427 );
buf \U$35858 ( \41550 , \40427 );
buf \U$35859 ( \41551 , \40427 );
buf \U$35860 ( \41552 , \40427 );
buf \U$35861 ( \41553 , \40427 );
buf \U$35862 ( \41554 , \40427 );
nor \U$35863 ( \41555 , \40413 , \40417 , \40420 , \40423 , \40426 , \40427 , \41529 , \41530 , \41531 , \41532 , \41533 , \41534 , \41535 , \41536 , \41537 , \41538 , \41539 , \41540 , \41541 , \41542 , \41543 , \41544 , \41545 , \41546 , \41547 , \41548 , \41549 , \41550 , \41551 , \41552 , \41553 , \41554 );
and \U$35864 ( \41556 , \8645 , \41555 );
buf \U$35865 ( \41557 , \40427 );
buf \U$35866 ( \41558 , \40427 );
buf \U$35867 ( \41559 , \40427 );
buf \U$35868 ( \41560 , \40427 );
buf \U$35869 ( \41561 , \40427 );
buf \U$35870 ( \41562 , \40427 );
buf \U$35871 ( \41563 , \40427 );
buf \U$35872 ( \41564 , \40427 );
buf \U$35873 ( \41565 , \40427 );
buf \U$35874 ( \41566 , \40427 );
buf \U$35875 ( \41567 , \40427 );
buf \U$35876 ( \41568 , \40427 );
buf \U$35877 ( \41569 , \40427 );
buf \U$35878 ( \41570 , \40427 );
buf \U$35879 ( \41571 , \40427 );
buf \U$35880 ( \41572 , \40427 );
buf \U$35881 ( \41573 , \40427 );
buf \U$35882 ( \41574 , \40427 );
buf \U$35883 ( \41575 , \40427 );
buf \U$35884 ( \41576 , \40427 );
buf \U$35885 ( \41577 , \40427 );
buf \U$35886 ( \41578 , \40427 );
buf \U$35887 ( \41579 , \40427 );
buf \U$35888 ( \41580 , \40427 );
buf \U$35889 ( \41581 , \40427 );
buf \U$35890 ( \41582 , \40427 );
nor \U$35891 ( \41583 , \40414 , \40416 , \40420 , \40423 , \40426 , \40427 , \41557 , \41558 , \41559 , \41560 , \41561 , \41562 , \41563 , \41564 , \41565 , \41566 , \41567 , \41568 , \41569 , \41570 , \41571 , \41572 , \41573 , \41574 , \41575 , \41576 , \41577 , \41578 , \41579 , \41580 , \41581 , \41582 );
and \U$35892 ( \41584 , \8673 , \41583 );
buf \U$35893 ( \41585 , \40427 );
buf \U$35894 ( \41586 , \40427 );
buf \U$35895 ( \41587 , \40427 );
buf \U$35896 ( \41588 , \40427 );
buf \U$35897 ( \41589 , \40427 );
buf \U$35898 ( \41590 , \40427 );
buf \U$35899 ( \41591 , \40427 );
buf \U$35900 ( \41592 , \40427 );
buf \U$35901 ( \41593 , \40427 );
buf \U$35902 ( \41594 , \40427 );
buf \U$35903 ( \41595 , \40427 );
buf \U$35904 ( \41596 , \40427 );
buf \U$35905 ( \41597 , \40427 );
buf \U$35906 ( \41598 , \40427 );
buf \U$35907 ( \41599 , \40427 );
buf \U$35908 ( \41600 , \40427 );
buf \U$35909 ( \41601 , \40427 );
buf \U$35910 ( \41602 , \40427 );
buf \U$35911 ( \41603 , \40427 );
buf \U$35912 ( \41604 , \40427 );
buf \U$35913 ( \41605 , \40427 );
buf \U$35914 ( \41606 , \40427 );
buf \U$35915 ( \41607 , \40427 );
buf \U$35916 ( \41608 , \40427 );
buf \U$35917 ( \41609 , \40427 );
buf \U$35918 ( \41610 , \40427 );
nor \U$35919 ( \41611 , \40413 , \40416 , \40420 , \40423 , \40426 , \40427 , \41585 , \41586 , \41587 , \41588 , \41589 , \41590 , \41591 , \41592 , \41593 , \41594 , \41595 , \41596 , \41597 , \41598 , \41599 , \41600 , \41601 , \41602 , \41603 , \41604 , \41605 , \41606 , \41607 , \41608 , \41609 , \41610 );
and \U$35920 ( \41612 , \8701 , \41611 );
buf \U$35921 ( \41613 , \40427 );
buf \U$35922 ( \41614 , \40427 );
buf \U$35923 ( \41615 , \40427 );
buf \U$35924 ( \41616 , \40427 );
buf \U$35925 ( \41617 , \40427 );
buf \U$35926 ( \41618 , \40427 );
buf \U$35927 ( \41619 , \40427 );
buf \U$35928 ( \41620 , \40427 );
buf \U$35929 ( \41621 , \40427 );
buf \U$35930 ( \41622 , \40427 );
buf \U$35931 ( \41623 , \40427 );
buf \U$35932 ( \41624 , \40427 );
buf \U$35933 ( \41625 , \40427 );
buf \U$35934 ( \41626 , \40427 );
buf \U$35935 ( \41627 , \40427 );
buf \U$35936 ( \41628 , \40427 );
buf \U$35937 ( \41629 , \40427 );
buf \U$35938 ( \41630 , \40427 );
buf \U$35939 ( \41631 , \40427 );
buf \U$35940 ( \41632 , \40427 );
buf \U$35941 ( \41633 , \40427 );
buf \U$35942 ( \41634 , \40427 );
buf \U$35943 ( \41635 , \40427 );
buf \U$35944 ( \41636 , \40427 );
buf \U$35945 ( \41637 , \40427 );
buf \U$35946 ( \41638 , \40427 );
nor \U$35947 ( \41639 , \40414 , \40417 , \40419 , \40423 , \40426 , \40427 , \41613 , \41614 , \41615 , \41616 , \41617 , \41618 , \41619 , \41620 , \41621 , \41622 , \41623 , \41624 , \41625 , \41626 , \41627 , \41628 , \41629 , \41630 , \41631 , \41632 , \41633 , \41634 , \41635 , \41636 , \41637 , \41638 );
and \U$35948 ( \41640 , \8729 , \41639 );
buf \U$35949 ( \41641 , \40427 );
buf \U$35950 ( \41642 , \40427 );
buf \U$35951 ( \41643 , \40427 );
buf \U$35952 ( \41644 , \40427 );
buf \U$35953 ( \41645 , \40427 );
buf \U$35954 ( \41646 , \40427 );
buf \U$35955 ( \41647 , \40427 );
buf \U$35956 ( \41648 , \40427 );
buf \U$35957 ( \41649 , \40427 );
buf \U$35958 ( \41650 , \40427 );
buf \U$35959 ( \41651 , \40427 );
buf \U$35960 ( \41652 , \40427 );
buf \U$35961 ( \41653 , \40427 );
buf \U$35962 ( \41654 , \40427 );
buf \U$35963 ( \41655 , \40427 );
buf \U$35964 ( \41656 , \40427 );
buf \U$35965 ( \41657 , \40427 );
buf \U$35966 ( \41658 , \40427 );
buf \U$35967 ( \41659 , \40427 );
buf \U$35968 ( \41660 , \40427 );
buf \U$35969 ( \41661 , \40427 );
buf \U$35970 ( \41662 , \40427 );
buf \U$35971 ( \41663 , \40427 );
buf \U$35972 ( \41664 , \40427 );
buf \U$35973 ( \41665 , \40427 );
buf \U$35974 ( \41666 , \40427 );
nor \U$35975 ( \41667 , \40413 , \40417 , \40419 , \40423 , \40426 , \40427 , \41641 , \41642 , \41643 , \41644 , \41645 , \41646 , \41647 , \41648 , \41649 , \41650 , \41651 , \41652 , \41653 , \41654 , \41655 , \41656 , \41657 , \41658 , \41659 , \41660 , \41661 , \41662 , \41663 , \41664 , \41665 , \41666 );
and \U$35976 ( \41668 , \8757 , \41667 );
buf \U$35977 ( \41669 , \40427 );
buf \U$35978 ( \41670 , \40427 );
buf \U$35979 ( \41671 , \40427 );
buf \U$35980 ( \41672 , \40427 );
buf \U$35981 ( \41673 , \40427 );
buf \U$35982 ( \41674 , \40427 );
buf \U$35983 ( \41675 , \40427 );
buf \U$35984 ( \41676 , \40427 );
buf \U$35985 ( \41677 , \40427 );
buf \U$35986 ( \41678 , \40427 );
buf \U$35987 ( \41679 , \40427 );
buf \U$35988 ( \41680 , \40427 );
buf \U$35989 ( \41681 , \40427 );
buf \U$35990 ( \41682 , \40427 );
buf \U$35991 ( \41683 , \40427 );
buf \U$35992 ( \41684 , \40427 );
buf \U$35993 ( \41685 , \40427 );
buf \U$35994 ( \41686 , \40427 );
buf \U$35995 ( \41687 , \40427 );
buf \U$35996 ( \41688 , \40427 );
buf \U$35997 ( \41689 , \40427 );
buf \U$35998 ( \41690 , \40427 );
buf \U$35999 ( \41691 , \40427 );
buf \U$36000 ( \41692 , \40427 );
buf \U$36001 ( \41693 , \40427 );
buf \U$36002 ( \41694 , \40427 );
nor \U$36003 ( \41695 , \40414 , \40416 , \40419 , \40423 , \40426 , \40427 , \41669 , \41670 , \41671 , \41672 , \41673 , \41674 , \41675 , \41676 , \41677 , \41678 , \41679 , \41680 , \41681 , \41682 , \41683 , \41684 , \41685 , \41686 , \41687 , \41688 , \41689 , \41690 , \41691 , \41692 , \41693 , \41694 );
and \U$36004 ( \41696 , \8785 , \41695 );
buf \U$36005 ( \41697 , \40427 );
buf \U$36006 ( \41698 , \40427 );
buf \U$36007 ( \41699 , \40427 );
buf \U$36008 ( \41700 , \40427 );
buf \U$36009 ( \41701 , \40427 );
buf \U$36010 ( \41702 , \40427 );
buf \U$36011 ( \41703 , \40427 );
buf \U$36012 ( \41704 , \40427 );
buf \U$36013 ( \41705 , \40427 );
buf \U$36014 ( \41706 , \40427 );
buf \U$36015 ( \41707 , \40427 );
buf \U$36016 ( \41708 , \40427 );
buf \U$36017 ( \41709 , \40427 );
buf \U$36018 ( \41710 , \40427 );
buf \U$36019 ( \41711 , \40427 );
buf \U$36020 ( \41712 , \40427 );
buf \U$36021 ( \41713 , \40427 );
buf \U$36022 ( \41714 , \40427 );
buf \U$36023 ( \41715 , \40427 );
buf \U$36024 ( \41716 , \40427 );
buf \U$36025 ( \41717 , \40427 );
buf \U$36026 ( \41718 , \40427 );
buf \U$36027 ( \41719 , \40427 );
buf \U$36028 ( \41720 , \40427 );
buf \U$36029 ( \41721 , \40427 );
buf \U$36030 ( \41722 , \40427 );
nor \U$36031 ( \41723 , \40413 , \40416 , \40419 , \40423 , \40426 , \40427 , \41697 , \41698 , \41699 , \41700 , \41701 , \41702 , \41703 , \41704 , \41705 , \41706 , \41707 , \41708 , \41709 , \41710 , \41711 , \41712 , \41713 , \41714 , \41715 , \41716 , \41717 , \41718 , \41719 , \41720 , \41721 , \41722 );
and \U$36032 ( \41724 , \8813 , \41723 );
buf \U$36033 ( \41725 , \40427 );
buf \U$36034 ( \41726 , \40427 );
buf \U$36035 ( \41727 , \40427 );
buf \U$36036 ( \41728 , \40427 );
buf \U$36037 ( \41729 , \40427 );
buf \U$36038 ( \41730 , \40427 );
buf \U$36039 ( \41731 , \40427 );
buf \U$36040 ( \41732 , \40427 );
buf \U$36041 ( \41733 , \40427 );
buf \U$36042 ( \41734 , \40427 );
buf \U$36043 ( \41735 , \40427 );
buf \U$36044 ( \41736 , \40427 );
buf \U$36045 ( \41737 , \40427 );
buf \U$36046 ( \41738 , \40427 );
buf \U$36047 ( \41739 , \40427 );
buf \U$36048 ( \41740 , \40427 );
buf \U$36049 ( \41741 , \40427 );
buf \U$36050 ( \41742 , \40427 );
buf \U$36051 ( \41743 , \40427 );
buf \U$36052 ( \41744 , \40427 );
buf \U$36053 ( \41745 , \40427 );
buf \U$36054 ( \41746 , \40427 );
buf \U$36055 ( \41747 , \40427 );
buf \U$36056 ( \41748 , \40427 );
buf \U$36057 ( \41749 , \40427 );
buf \U$36058 ( \41750 , \40427 );
nor \U$36059 ( \41751 , \40414 , \40417 , \40420 , \40422 , \40426 , \40427 , \41725 , \41726 , \41727 , \41728 , \41729 , \41730 , \41731 , \41732 , \41733 , \41734 , \41735 , \41736 , \41737 , \41738 , \41739 , \41740 , \41741 , \41742 , \41743 , \41744 , \41745 , \41746 , \41747 , \41748 , \41749 , \41750 );
and \U$36060 ( \41752 , \8841 , \41751 );
buf \U$36061 ( \41753 , \40427 );
buf \U$36062 ( \41754 , \40427 );
buf \U$36063 ( \41755 , \40427 );
buf \U$36064 ( \41756 , \40427 );
buf \U$36065 ( \41757 , \40427 );
buf \U$36066 ( \41758 , \40427 );
buf \U$36067 ( \41759 , \40427 );
buf \U$36068 ( \41760 , \40427 );
buf \U$36069 ( \41761 , \40427 );
buf \U$36070 ( \41762 , \40427 );
buf \U$36071 ( \41763 , \40427 );
buf \U$36072 ( \41764 , \40427 );
buf \U$36073 ( \41765 , \40427 );
buf \U$36074 ( \41766 , \40427 );
buf \U$36075 ( \41767 , \40427 );
buf \U$36076 ( \41768 , \40427 );
buf \U$36077 ( \41769 , \40427 );
buf \U$36078 ( \41770 , \40427 );
buf \U$36079 ( \41771 , \40427 );
buf \U$36080 ( \41772 , \40427 );
buf \U$36081 ( \41773 , \40427 );
buf \U$36082 ( \41774 , \40427 );
buf \U$36083 ( \41775 , \40427 );
buf \U$36084 ( \41776 , \40427 );
buf \U$36085 ( \41777 , \40427 );
buf \U$36086 ( \41778 , \40427 );
nor \U$36087 ( \41779 , \40413 , \40417 , \40420 , \40422 , \40426 , \40427 , \41753 , \41754 , \41755 , \41756 , \41757 , \41758 , \41759 , \41760 , \41761 , \41762 , \41763 , \41764 , \41765 , \41766 , \41767 , \41768 , \41769 , \41770 , \41771 , \41772 , \41773 , \41774 , \41775 , \41776 , \41777 , \41778 );
and \U$36088 ( \41780 , \8869 , \41779 );
buf \U$36089 ( \41781 , \40427 );
buf \U$36090 ( \41782 , \40427 );
buf \U$36091 ( \41783 , \40427 );
buf \U$36092 ( \41784 , \40427 );
buf \U$36093 ( \41785 , \40427 );
buf \U$36094 ( \41786 , \40427 );
buf \U$36095 ( \41787 , \40427 );
buf \U$36096 ( \41788 , \40427 );
buf \U$36097 ( \41789 , \40427 );
buf \U$36098 ( \41790 , \40427 );
buf \U$36099 ( \41791 , \40427 );
buf \U$36100 ( \41792 , \40427 );
buf \U$36101 ( \41793 , \40427 );
buf \U$36102 ( \41794 , \40427 );
buf \U$36103 ( \41795 , \40427 );
buf \U$36104 ( \41796 , \40427 );
buf \U$36105 ( \41797 , \40427 );
buf \U$36106 ( \41798 , \40427 );
buf \U$36107 ( \41799 , \40427 );
buf \U$36108 ( \41800 , \40427 );
buf \U$36109 ( \41801 , \40427 );
buf \U$36110 ( \41802 , \40427 );
buf \U$36111 ( \41803 , \40427 );
buf \U$36112 ( \41804 , \40427 );
buf \U$36113 ( \41805 , \40427 );
buf \U$36114 ( \41806 , \40427 );
nor \U$36115 ( \41807 , \40414 , \40416 , \40420 , \40422 , \40426 , \40427 , \41781 , \41782 , \41783 , \41784 , \41785 , \41786 , \41787 , \41788 , \41789 , \41790 , \41791 , \41792 , \41793 , \41794 , \41795 , \41796 , \41797 , \41798 , \41799 , \41800 , \41801 , \41802 , \41803 , \41804 , \41805 , \41806 );
and \U$36116 ( \41808 , \8897 , \41807 );
buf \U$36117 ( \41809 , \40427 );
buf \U$36118 ( \41810 , \40427 );
buf \U$36119 ( \41811 , \40427 );
buf \U$36120 ( \41812 , \40427 );
buf \U$36121 ( \41813 , \40427 );
buf \U$36122 ( \41814 , \40427 );
buf \U$36123 ( \41815 , \40427 );
buf \U$36124 ( \41816 , \40427 );
buf \U$36125 ( \41817 , \40427 );
buf \U$36126 ( \41818 , \40427 );
buf \U$36127 ( \41819 , \40427 );
buf \U$36128 ( \41820 , \40427 );
buf \U$36129 ( \41821 , \40427 );
buf \U$36130 ( \41822 , \40427 );
buf \U$36131 ( \41823 , \40427 );
buf \U$36132 ( \41824 , \40427 );
buf \U$36133 ( \41825 , \40427 );
buf \U$36134 ( \41826 , \40427 );
buf \U$36135 ( \41827 , \40427 );
buf \U$36136 ( \41828 , \40427 );
buf \U$36137 ( \41829 , \40427 );
buf \U$36138 ( \41830 , \40427 );
buf \U$36139 ( \41831 , \40427 );
buf \U$36140 ( \41832 , \40427 );
buf \U$36141 ( \41833 , \40427 );
buf \U$36142 ( \41834 , \40427 );
nor \U$36143 ( \41835 , \40413 , \40416 , \40420 , \40422 , \40426 , \40427 , \41809 , \41810 , \41811 , \41812 , \41813 , \41814 , \41815 , \41816 , \41817 , \41818 , \41819 , \41820 , \41821 , \41822 , \41823 , \41824 , \41825 , \41826 , \41827 , \41828 , \41829 , \41830 , \41831 , \41832 , \41833 , \41834 );
and \U$36144 ( \41836 , \8925 , \41835 );
buf \U$36145 ( \41837 , \40427 );
buf \U$36146 ( \41838 , \40427 );
buf \U$36147 ( \41839 , \40427 );
buf \U$36148 ( \41840 , \40427 );
buf \U$36149 ( \41841 , \40427 );
buf \U$36150 ( \41842 , \40427 );
buf \U$36151 ( \41843 , \40427 );
buf \U$36152 ( \41844 , \40427 );
buf \U$36153 ( \41845 , \40427 );
buf \U$36154 ( \41846 , \40427 );
buf \U$36155 ( \41847 , \40427 );
buf \U$36156 ( \41848 , \40427 );
buf \U$36157 ( \41849 , \40427 );
buf \U$36158 ( \41850 , \40427 );
buf \U$36159 ( \41851 , \40427 );
buf \U$36160 ( \41852 , \40427 );
buf \U$36161 ( \41853 , \40427 );
buf \U$36162 ( \41854 , \40427 );
buf \U$36163 ( \41855 , \40427 );
buf \U$36164 ( \41856 , \40427 );
buf \U$36165 ( \41857 , \40427 );
buf \U$36166 ( \41858 , \40427 );
buf \U$36167 ( \41859 , \40427 );
buf \U$36168 ( \41860 , \40427 );
buf \U$36169 ( \41861 , \40427 );
buf \U$36170 ( \41862 , \40427 );
nor \U$36171 ( \41863 , \40414 , \40417 , \40419 , \40422 , \40426 , \40427 , \41837 , \41838 , \41839 , \41840 , \41841 , \41842 , \41843 , \41844 , \41845 , \41846 , \41847 , \41848 , \41849 , \41850 , \41851 , \41852 , \41853 , \41854 , \41855 , \41856 , \41857 , \41858 , \41859 , \41860 , \41861 , \41862 );
and \U$36172 ( \41864 , \8953 , \41863 );
buf \U$36173 ( \41865 , \40427 );
buf \U$36174 ( \41866 , \40427 );
buf \U$36175 ( \41867 , \40427 );
buf \U$36176 ( \41868 , \40427 );
buf \U$36177 ( \41869 , \40427 );
buf \U$36178 ( \41870 , \40427 );
buf \U$36179 ( \41871 , \40427 );
buf \U$36180 ( \41872 , \40427 );
buf \U$36181 ( \41873 , \40427 );
buf \U$36182 ( \41874 , \40427 );
buf \U$36183 ( \41875 , \40427 );
buf \U$36184 ( \41876 , \40427 );
buf \U$36185 ( \41877 , \40427 );
buf \U$36186 ( \41878 , \40427 );
buf \U$36187 ( \41879 , \40427 );
buf \U$36188 ( \41880 , \40427 );
buf \U$36189 ( \41881 , \40427 );
buf \U$36190 ( \41882 , \40427 );
buf \U$36191 ( \41883 , \40427 );
buf \U$36192 ( \41884 , \40427 );
buf \U$36193 ( \41885 , \40427 );
buf \U$36194 ( \41886 , \40427 );
buf \U$36195 ( \41887 , \40427 );
buf \U$36196 ( \41888 , \40427 );
buf \U$36197 ( \41889 , \40427 );
buf \U$36198 ( \41890 , \40427 );
nor \U$36199 ( \41891 , \40413 , \40417 , \40419 , \40422 , \40426 , \40427 , \41865 , \41866 , \41867 , \41868 , \41869 , \41870 , \41871 , \41872 , \41873 , \41874 , \41875 , \41876 , \41877 , \41878 , \41879 , \41880 , \41881 , \41882 , \41883 , \41884 , \41885 , \41886 , \41887 , \41888 , \41889 , \41890 );
and \U$36200 ( \41892 , \8981 , \41891 );
buf \U$36201 ( \41893 , \40427 );
buf \U$36202 ( \41894 , \40427 );
buf \U$36203 ( \41895 , \40427 );
buf \U$36204 ( \41896 , \40427 );
buf \U$36205 ( \41897 , \40427 );
buf \U$36206 ( \41898 , \40427 );
buf \U$36207 ( \41899 , \40427 );
buf \U$36208 ( \41900 , \40427 );
buf \U$36209 ( \41901 , \40427 );
buf \U$36210 ( \41902 , \40427 );
buf \U$36211 ( \41903 , \40427 );
buf \U$36212 ( \41904 , \40427 );
buf \U$36213 ( \41905 , \40427 );
buf \U$36214 ( \41906 , \40427 );
buf \U$36215 ( \41907 , \40427 );
buf \U$36216 ( \41908 , \40427 );
buf \U$36217 ( \41909 , \40427 );
buf \U$36218 ( \41910 , \40427 );
buf \U$36219 ( \41911 , \40427 );
buf \U$36220 ( \41912 , \40427 );
buf \U$36221 ( \41913 , \40427 );
buf \U$36222 ( \41914 , \40427 );
buf \U$36223 ( \41915 , \40427 );
buf \U$36224 ( \41916 , \40427 );
buf \U$36225 ( \41917 , \40427 );
buf \U$36226 ( \41918 , \40427 );
nor \U$36227 ( \41919 , \40414 , \40416 , \40419 , \40422 , \40426 , \40427 , \41893 , \41894 , \41895 , \41896 , \41897 , \41898 , \41899 , \41900 , \41901 , \41902 , \41903 , \41904 , \41905 , \41906 , \41907 , \41908 , \41909 , \41910 , \41911 , \41912 , \41913 , \41914 , \41915 , \41916 , \41917 , \41918 );
and \U$36228 ( \41920 , \9009 , \41919 );
or \U$36229 ( \41921 , 1'b0 , \41528 , \41556 , \41584 , \41612 , \41640 , \41668 , \41696 , \41724 , \41752 , \41780 , \41808 , \41836 , \41864 , \41892 , \41920 );
buf \U$36230 ( \41922 , \40427 );
not \U$36231 ( \41923 , \41922 );
buf \U$36232 ( \41924 , \40416 );
buf \U$36233 ( \41925 , \40419 );
buf \U$36234 ( \41926 , \40422 );
buf \U$36235 ( \41927 , \40426 );
buf \U$36236 ( \41928 , \40427 );
buf \U$36237 ( \41929 , \40427 );
buf \U$36238 ( \41930 , \40427 );
buf \U$36239 ( \41931 , \40427 );
buf \U$36240 ( \41932 , \40427 );
buf \U$36241 ( \41933 , \40427 );
buf \U$36242 ( \41934 , \40427 );
buf \U$36243 ( \41935 , \40427 );
buf \U$36244 ( \41936 , \40427 );
buf \U$36245 ( \41937 , \40427 );
buf \U$36246 ( \41938 , \40427 );
buf \U$36247 ( \41939 , \40427 );
buf \U$36248 ( \41940 , \40427 );
buf \U$36249 ( \41941 , \40427 );
buf \U$36250 ( \41942 , \40427 );
buf \U$36251 ( \41943 , \40427 );
buf \U$36252 ( \41944 , \40427 );
buf \U$36253 ( \41945 , \40427 );
buf \U$36254 ( \41946 , \40427 );
buf \U$36255 ( \41947 , \40427 );
buf \U$36256 ( \41948 , \40427 );
buf \U$36257 ( \41949 , \40427 );
buf \U$36258 ( \41950 , \40427 );
buf \U$36259 ( \41951 , \40427 );
buf \U$36260 ( \41952 , \40427 );
buf \U$36261 ( \41953 , \40427 );
buf \U$36262 ( \41954 , \40413 );
or \U$36263 ( \41955 , \41924 , \41925 , \41926 , \41927 , \41928 , \41929 , \41930 , \41931 , \41932 , \41933 , \41934 , \41935 , \41936 , \41937 , \41938 , \41939 , \41940 , \41941 , \41942 , \41943 , \41944 , \41945 , \41946 , \41947 , \41948 , \41949 , \41950 , \41951 , \41952 , \41953 , \41954 );
nand \U$36264 ( \41956 , \41923 , \41955 );
buf \U$36265 ( \41957 , \41956 );
or \U$36267 ( \41958 , \41957 , 1'b0 );
_DC gbb1a ( \41959_nGbb1a , \41921 , \41958 );
buf \U$36268 ( \41960 , \41959_nGbb1a );
xor \U$36269 ( \41961 , \41500 , \41960 );
buf \U$36270 ( \41962 , RIb7af5b8_255);
and \U$36272 ( \41963 , \7209 , \41527 );
and \U$36273 ( \41964 , \9119 , \41555 );
and \U$36274 ( \41965 , \9121 , \41583 );
and \U$36275 ( \41966 , \9123 , \41611 );
and \U$36276 ( \41967 , \9125 , \41639 );
and \U$36277 ( \41968 , \9127 , \41667 );
and \U$36278 ( \41969 , \9129 , \41695 );
and \U$36279 ( \41970 , \9131 , \41723 );
and \U$36280 ( \41971 , \9133 , \41751 );
and \U$36281 ( \41972 , \9135 , \41779 );
and \U$36282 ( \41973 , \9137 , \41807 );
and \U$36283 ( \41974 , \9139 , \41835 );
and \U$36284 ( \41975 , \9141 , \41863 );
and \U$36285 ( \41976 , \9143 , \41891 );
and \U$36286 ( \41977 , \9145 , \41919 );
or \U$36287 ( \41978 , 1'b0 , \41963 , \41964 , \41965 , \41966 , \41967 , \41968 , \41969 , \41970 , \41971 , \41972 , \41973 , \41974 , \41975 , \41976 , \41977 );
_DC gbb2e ( \41979_nGbb2e , \41978 , \41958 );
buf \U$36288 ( \41980 , \41979_nGbb2e );
xor \U$36289 ( \41981 , \41962 , \41980 );
or \U$36290 ( \41982 , \41961 , \41981 );
buf \U$36291 ( \41983 , RIb7af540_256);
and \U$36293 ( \41984 , \7219 , \41527 );
and \U$36294 ( \41985 , \9155 , \41555 );
and \U$36295 ( \41986 , \9157 , \41583 );
and \U$36296 ( \41987 , \9159 , \41611 );
and \U$36297 ( \41988 , \9161 , \41639 );
and \U$36298 ( \41989 , \9163 , \41667 );
and \U$36299 ( \41990 , \9165 , \41695 );
and \U$36300 ( \41991 , \9167 , \41723 );
and \U$36301 ( \41992 , \9169 , \41751 );
and \U$36302 ( \41993 , \9171 , \41779 );
and \U$36303 ( \41994 , \9173 , \41807 );
and \U$36304 ( \41995 , \9175 , \41835 );
and \U$36305 ( \41996 , \9177 , \41863 );
and \U$36306 ( \41997 , \9179 , \41891 );
and \U$36307 ( \41998 , \9181 , \41919 );
or \U$36308 ( \41999 , 1'b0 , \41984 , \41985 , \41986 , \41987 , \41988 , \41989 , \41990 , \41991 , \41992 , \41993 , \41994 , \41995 , \41996 , \41997 , \41998 );
_DC gbb43 ( \42000_nGbb43 , \41999 , \41958 );
buf \U$36309 ( \42001 , \42000_nGbb43 );
xor \U$36310 ( \42002 , \41983 , \42001 );
or \U$36311 ( \42003 , \41982 , \42002 );
buf \U$36312 ( \42004 , RIb7af4c8_257);
and \U$36314 ( \42005 , \7229 , \41527 );
and \U$36315 ( \42006 , \9191 , \41555 );
and \U$36316 ( \42007 , \9193 , \41583 );
and \U$36317 ( \42008 , \9195 , \41611 );
and \U$36318 ( \42009 , \9197 , \41639 );
and \U$36319 ( \42010 , \9199 , \41667 );
and \U$36320 ( \42011 , \9201 , \41695 );
and \U$36321 ( \42012 , \9203 , \41723 );
and \U$36322 ( \42013 , \9205 , \41751 );
and \U$36323 ( \42014 , \9207 , \41779 );
and \U$36324 ( \42015 , \9209 , \41807 );
and \U$36325 ( \42016 , \9211 , \41835 );
and \U$36326 ( \42017 , \9213 , \41863 );
and \U$36327 ( \42018 , \9215 , \41891 );
and \U$36328 ( \42019 , \9217 , \41919 );
or \U$36329 ( \42020 , 1'b0 , \42005 , \42006 , \42007 , \42008 , \42009 , \42010 , \42011 , \42012 , \42013 , \42014 , \42015 , \42016 , \42017 , \42018 , \42019 );
_DC gbb58 ( \42021_nGbb58 , \42020 , \41958 );
buf \U$36330 ( \42022 , \42021_nGbb58 );
xor \U$36331 ( \42023 , \42004 , \42022 );
or \U$36332 ( \42024 , \42003 , \42023 );
buf \U$36333 ( \42025 , RIb7af450_258);
and \U$36335 ( \42026 , \7239 , \41527 );
and \U$36336 ( \42027 , \9227 , \41555 );
and \U$36337 ( \42028 , \9229 , \41583 );
and \U$36338 ( \42029 , \9231 , \41611 );
and \U$36339 ( \42030 , \9233 , \41639 );
and \U$36340 ( \42031 , \9235 , \41667 );
and \U$36341 ( \42032 , \9237 , \41695 );
and \U$36342 ( \42033 , \9239 , \41723 );
and \U$36343 ( \42034 , \9241 , \41751 );
and \U$36344 ( \42035 , \9243 , \41779 );
and \U$36345 ( \42036 , \9245 , \41807 );
and \U$36346 ( \42037 , \9247 , \41835 );
and \U$36347 ( \42038 , \9249 , \41863 );
and \U$36348 ( \42039 , \9251 , \41891 );
and \U$36349 ( \42040 , \9253 , \41919 );
or \U$36350 ( \42041 , 1'b0 , \42026 , \42027 , \42028 , \42029 , \42030 , \42031 , \42032 , \42033 , \42034 , \42035 , \42036 , \42037 , \42038 , \42039 , \42040 );
_DC gbb6d ( \42042_nGbb6d , \42041 , \41958 );
buf \U$36351 ( \42043 , \42042_nGbb6d );
xor \U$36352 ( \42044 , \42025 , \42043 );
or \U$36353 ( \42045 , \42024 , \42044 );
buf \U$36354 ( \42046 , RIb7af3d8_259);
and \U$36356 ( \42047 , \7249 , \41527 );
and \U$36357 ( \42048 , \9263 , \41555 );
and \U$36358 ( \42049 , \9265 , \41583 );
and \U$36359 ( \42050 , \9267 , \41611 );
and \U$36360 ( \42051 , \9269 , \41639 );
and \U$36361 ( \42052 , \9271 , \41667 );
and \U$36362 ( \42053 , \9273 , \41695 );
and \U$36363 ( \42054 , \9275 , \41723 );
and \U$36364 ( \42055 , \9277 , \41751 );
and \U$36365 ( \42056 , \9279 , \41779 );
and \U$36366 ( \42057 , \9281 , \41807 );
and \U$36367 ( \42058 , \9283 , \41835 );
and \U$36368 ( \42059 , \9285 , \41863 );
and \U$36369 ( \42060 , \9287 , \41891 );
and \U$36370 ( \42061 , \9289 , \41919 );
or \U$36371 ( \42062 , 1'b0 , \42047 , \42048 , \42049 , \42050 , \42051 , \42052 , \42053 , \42054 , \42055 , \42056 , \42057 , \42058 , \42059 , \42060 , \42061 );
_DC gbb82 ( \42063_nGbb82 , \42062 , \41958 );
buf \U$36372 ( \42064 , \42063_nGbb82 );
xor \U$36373 ( \42065 , \42046 , \42064 );
or \U$36374 ( \42066 , \42045 , \42065 );
buf \U$36375 ( \42067 , RIb7a5bf8_260);
and \U$36377 ( \42068 , \7259 , \41527 );
and \U$36378 ( \42069 , \9299 , \41555 );
and \U$36379 ( \42070 , \9301 , \41583 );
and \U$36380 ( \42071 , \9303 , \41611 );
and \U$36381 ( \42072 , \9305 , \41639 );
and \U$36382 ( \42073 , \9307 , \41667 );
and \U$36383 ( \42074 , \9309 , \41695 );
and \U$36384 ( \42075 , \9311 , \41723 );
and \U$36385 ( \42076 , \9313 , \41751 );
and \U$36386 ( \42077 , \9315 , \41779 );
and \U$36387 ( \42078 , \9317 , \41807 );
and \U$36388 ( \42079 , \9319 , \41835 );
and \U$36389 ( \42080 , \9321 , \41863 );
and \U$36390 ( \42081 , \9323 , \41891 );
and \U$36391 ( \42082 , \9325 , \41919 );
or \U$36392 ( \42083 , 1'b0 , \42068 , \42069 , \42070 , \42071 , \42072 , \42073 , \42074 , \42075 , \42076 , \42077 , \42078 , \42079 , \42080 , \42081 , \42082 );
_DC gbb97 ( \42084_nGbb97 , \42083 , \41958 );
buf \U$36393 ( \42085 , \42084_nGbb97 );
xor \U$36394 ( \42086 , \42067 , \42085 );
or \U$36395 ( \42087 , \42066 , \42086 );
buf \U$36396 ( \42088 , RIb7a0c48_261);
and \U$36398 ( \42089 , \7269 , \41527 );
and \U$36399 ( \42090 , \9335 , \41555 );
and \U$36400 ( \42091 , \9337 , \41583 );
and \U$36401 ( \42092 , \9339 , \41611 );
and \U$36402 ( \42093 , \9341 , \41639 );
and \U$36403 ( \42094 , \9343 , \41667 );
and \U$36404 ( \42095 , \9345 , \41695 );
and \U$36405 ( \42096 , \9347 , \41723 );
and \U$36406 ( \42097 , \9349 , \41751 );
and \U$36407 ( \42098 , \9351 , \41779 );
and \U$36408 ( \42099 , \9353 , \41807 );
and \U$36409 ( \42100 , \9355 , \41835 );
and \U$36410 ( \42101 , \9357 , \41863 );
and \U$36411 ( \42102 , \9359 , \41891 );
and \U$36412 ( \42103 , \9361 , \41919 );
or \U$36413 ( \42104 , 1'b0 , \42089 , \42090 , \42091 , \42092 , \42093 , \42094 , \42095 , \42096 , \42097 , \42098 , \42099 , \42100 , \42101 , \42102 , \42103 );
_DC gbbac ( \42105_nGbbac , \42104 , \41958 );
buf \U$36414 ( \42106 , \42105_nGbbac );
xor \U$36415 ( \42107 , \42088 , \42106 );
or \U$36416 ( \42108 , \42087 , \42107 );
not \U$36417 ( \42109 , \42108 );
buf \U$36418 ( \42110 , \42109 );
and \U$36419 ( \42111 , \41499 , \42110 );
_HMUX gbbb3 ( \42112_nGbbb3 , \40002_nGb36e , \40413 , \42111 );
buf \U$36420 ( \42113 , RIea91330_6888);
buf \U$36421 ( \42114 , RIe5319e0_6884);
buf \U$36422 ( \42115 , RIe549ef0_6842);
buf \U$36423 ( \42116 , RIe549770_6843);
buf \U$36424 ( \42117 , RIe548ff0_6844);
or \U$36425 ( \42118 , \42114 , \42115 , \42116 , \42117 );
and \U$36426 ( \42119 , \42113 , \42118 );
buf \U$36427 ( \42120 , \42119 );
_HMUX gbbbc ( \42121_nGbbbc , \40411_nGb50a , \42112_nGbbb3 , \42120 );
_HMUX gbbbd ( \42122_nGbbbd , RIe549ef0_6842 , \7081 , \7279 );
_HMUX gbbbe ( \42123_nGbbbe , RIe549ef0_6842 , \7282 , \9370 );
_HMUX gbbbf ( \42124_nGbbbf , \42122_nGbbbd , \42123_nGbbbe , \9381 );
_HMUX gbbc0 ( \42125_nGbbc0 , \42124_nGbbbf , \9387 , \9571 );
_HMUX gbbc1 ( \42126_nGbbc1 , \42124_nGbbbf , \9574 , \11438 );
_HMUX gbbc2 ( \42127_nGbbc2 , \42125_nGbbc0 , \42126_nGbbc1 , \11449 );
_HMUX gbbc3 ( \42128_nGbbc3 , \42127_nGbbc2 , \11456 , \11660 );
_HMUX gbbc4 ( \42129_nGbbc4 , \42127_nGbbc2 , \11663 , \13527 );
_HMUX gbbc5 ( \42130_nGbbc5 , \42128_nGbbc3 , \42129_nGbbc4 , \13538 );
_HMUX gbbc6 ( \42131_nGbbc6 , \42130_nGbbc5 , \13543 , \13763 );
_HMUX gbbc7 ( \42132_nGbbc7 , \42130_nGbbc5 , \13766 , \15630 );
_HMUX gbbc8 ( \42133_nGbbc8 , \42131_nGbbc6 , \42132_nGbbc7 , \15641 );
_HMUX gbbc9 ( \42134_nGbbc9 , \42133_nGbbc8 , \15648 , \15889 );
_HMUX gbbca ( \42135_nGbbca , \42133_nGbbc8 , \15892 , \17756 );
_HMUX gbbcb ( \42136_nGbbcb , \42134_nGbbc9 , \42135_nGbbca , \17767 );
_HMUX gbbcc ( \42137_nGbbcc , \42136_nGbbcb , \17773 , \18031 );
_HMUX gbbcd ( \42138_nGbbcd , \42136_nGbbcb , \18034 , \19898 );
_HMUX gbbce ( \42139_nGbbce , \42137_nGbbcc , \42138_nGbbcd , \19909 );
_HMUX gbbcf ( \42140_nGbbcf , \42139_nGbbce , \19916 , \20193 );
_HMUX gbbd0 ( \42141_nGbbd0 , \42139_nGbbce , \20196 , \22060 );
_HMUX gbbd1 ( \42142_nGbbd1 , \42140_nGbbcf , \42141_nGbbd0 , \22071 );
_HMUX gbbd2 ( \42143_nGbbd2 , \42142_nGbbd1 , \22076 , \22367 );
_HMUX gbbd3 ( \42144_nGbbd3 , \42142_nGbbd1 , \22370 , \24234 );
_HMUX gbbd4 ( \42145_nGbbd4 , \42143_nGbbd2 , \42144_nGbbd3 , \24245 );
_HMUX gbbd5 ( \42146_nGbbd5 , \42145_nGbbd4 , \24252 , \24565 );
_HMUX gbbd6 ( \42147_nGbbd6 , \42145_nGbbd4 , \24568 , \26432 );
_HMUX gbbd7 ( \42148_nGbbd7 , \42146_nGbbd5 , \42147_nGbbd6 , \26443 );
_HMUX gbbd8 ( \42149_nGbbd8 , \42148_nGbbd7 , \26449 , \26779 );
_HMUX gbbd9 ( \42150_nGbbd9 , \42148_nGbbd7 , \26782 , \28646 );
_HMUX gbbda ( \42151_nGbbda , \42149_nGbbd8 , \42150_nGbbd9 , \28657 );
_HMUX gbbdb ( \42152_nGbbdb , \42151_nGbbda , \28664 , \29013 );
_HMUX gbbdc ( \42153_nGbbdc , \42151_nGbbda , \29016 , \30880 );
_HMUX gbbdd ( \42154_nGbbdd , \42152_nGbbdb , \42153_nGbbdc , \30891 );
_HMUX gbbde ( \42155_nGbbde , \42154_nGbbdd , \30896 , \31261 );
_HMUX gbbdf ( \42156_nGbbdf , \42154_nGbbdd , \31264 , \33128 );
_HMUX gbbe0 ( \42157_nGbbe0 , \42155_nGbbde , \42156_nGbbdf , \33139 );
_HMUX gbbe1 ( \42158_nGbbe1 , \42157_nGbbe0 , \33146 , \33531 );
_HMUX gbbe2 ( \42159_nGbbe2 , \42157_nGbbe0 , \33534 , \35398 );
_HMUX gbbe3 ( \42160_nGbbe3 , \42158_nGbbe1 , \42159_nGbbe2 , \35409 );
_HMUX gbbe4 ( \42161_nGbbe4 , \42160_nGbbe3 , \35415 , \35817 );
_HMUX gbbe5 ( \42162_nGbbe5 , \42160_nGbbe3 , \35820 , \37684 );
_HMUX gbbe6 ( \42163_nGbbe6 , \42161_nGbbe4 , \42162_nGbbe5 , \37695 );
_HMUX gbbe7 ( \42164_nGbbe7 , \42163_nGbbe6 , \37702 , \38123 );
_HMUX gbbe8 ( \42165_nGbbe8 , \42163_nGbbe6 , \38126 , \39990 );
_HMUX gbbe9 ( \42166_nGbbe9 , \42164_nGbbe7 , \42165_nGbbe8 , \40001 );
_HMUX gbbea ( \42167_nGbbea , \42166_nGbbe9 , RIe549ef0_6842 , \40410 );
_HMUX gbbeb ( \42168_nGbbeb , \42166_nGbbe9 , \40416 , \42111 );
_HMUX gbbec ( \42169_nGbbec , \42167_nGbbea , \42168_nGbbeb , \42120 );
not \U$36428 ( \42170 , \42169_nGbbec );
_HMUX gbbed ( \42171_nGbbed , RIe549770_6843 , \7085 , \7279 );
_HMUX gbbee ( \42172_nGbbee , RIe549770_6843 , \7283 , \9370 );
_HMUX gbbef ( \42173_nGbbef , \42171_nGbbed , \42172_nGbbee , \9381 );
_HMUX gbbf0 ( \42174_nGbbf0 , \42173_nGbbef , \9390 , \9571 );
_HMUX gbbf1 ( \42175_nGbbf1 , \42173_nGbbef , \9575 , \11438 );
_HMUX gbbf2 ( \42176_nGbbf2 , \42174_nGbbf0 , \42175_nGbbf1 , \11449 );
_HMUX gbbf3 ( \42177_nGbbf3 , \42176_nGbbf2 , \11460 , \11660 );
_HMUX gbbf4 ( \42178_nGbbf4 , \42176_nGbbf2 , \11664 , \13527 );
_HMUX gbbf5 ( \42179_nGbbf5 , \42177_nGbbf3 , \42178_nGbbf4 , \13538 );
_HMUX gbbf6 ( \42180_nGbbf6 , \42179_nGbbf5 , \13546 , \13763 );
_HMUX gbbf7 ( \42181_nGbbf7 , \42179_nGbbf5 , \13767 , \15630 );
_HMUX gbbf8 ( \42182_nGbbf8 , \42180_nGbbf6 , \42181_nGbbf7 , \15641 );
_HMUX gbbf9 ( \42183_nGbbf9 , \42182_nGbbf8 , \15652 , \15889 );
_HMUX gbbfa ( \42184_nGbbfa , \42182_nGbbf8 , \15893 , \17756 );
_HMUX gbbfb ( \42185_nGbbfb , \42183_nGbbf9 , \42184_nGbbfa , \17767 );
_HMUX gbbfc ( \42186_nGbbfc , \42185_nGbbfb , \17776 , \18031 );
_HMUX gbbfd ( \42187_nGbbfd , \42185_nGbbfb , \18035 , \19898 );
_HMUX gbbfe ( \42188_nGbbfe , \42186_nGbbfc , \42187_nGbbfd , \19909 );
_HMUX gbbff ( \42189_nGbbff , \42188_nGbbfe , \19920 , \20193 );
_HMUX gbc00 ( \42190_nGbc00 , \42188_nGbbfe , \20197 , \22060 );
_HMUX gbc01 ( \42191_nGbc01 , \42189_nGbbff , \42190_nGbc00 , \22071 );
_HMUX gbc02 ( \42192_nGbc02 , \42191_nGbc01 , \22078 , \22367 );
_HMUX gbc03 ( \42193_nGbc03 , \42191_nGbc01 , \22371 , \24234 );
_HMUX gbc04 ( \42194_nGbc04 , \42192_nGbc02 , \42193_nGbc03 , \24245 );
_HMUX gbc05 ( \42195_nGbc05 , \42194_nGbc04 , \24256 , \24565 );
_HMUX gbc06 ( \42196_nGbc06 , \42194_nGbc04 , \24569 , \26432 );
_HMUX gbc07 ( \42197_nGbc07 , \42195_nGbc05 , \42196_nGbc06 , \26443 );
_HMUX gbc08 ( \42198_nGbc08 , \42197_nGbc07 , \26452 , \26779 );
_HMUX gbc09 ( \42199_nGbc09 , \42197_nGbc07 , \26783 , \28646 );
_HMUX gbc0a ( \42200_nGbc0a , \42198_nGbc08 , \42199_nGbc09 , \28657 );
_HMUX gbc0b ( \42201_nGbc0b , \42200_nGbc0a , \28668 , \29013 );
_HMUX gbc0c ( \42202_nGbc0c , \42200_nGbc0a , \29017 , \30880 );
_HMUX gbc0d ( \42203_nGbc0d , \42201_nGbc0b , \42202_nGbc0c , \30891 );
_HMUX gbc0e ( \42204_nGbc0e , \42203_nGbc0d , \30899 , \31261 );
_HMUX gbc0f ( \42205_nGbc0f , \42203_nGbc0d , \31265 , \33128 );
_HMUX gbc10 ( \42206_nGbc10 , \42204_nGbc0e , \42205_nGbc0f , \33139 );
_HMUX gbc11 ( \42207_nGbc11 , \42206_nGbc10 , \33150 , \33531 );
_HMUX gbc12 ( \42208_nGbc12 , \42206_nGbc10 , \33535 , \35398 );
_HMUX gbc13 ( \42209_nGbc13 , \42207_nGbc11 , \42208_nGbc12 , \35409 );
_HMUX gbc14 ( \42210_nGbc14 , \42209_nGbc13 , \35418 , \35817 );
_HMUX gbc15 ( \42211_nGbc15 , \42209_nGbc13 , \35821 , \37684 );
_HMUX gbc16 ( \42212_nGbc16 , \42210_nGbc14 , \42211_nGbc15 , \37695 );
_HMUX gbc17 ( \42213_nGbc17 , \42212_nGbc16 , \37706 , \38123 );
_HMUX gbc18 ( \42214_nGbc18 , \42212_nGbc16 , \38127 , \39990 );
_HMUX gbc19 ( \42215_nGbc19 , \42213_nGbc17 , \42214_nGbc18 , \40001 );
_HMUX gbc1a ( \42216_nGbc1a , \42215_nGbc19 , RIe549770_6843 , \40410 );
_HMUX gbc1b ( \42217_nGbc1b , \42215_nGbc19 , \40419 , \42111 );
_HMUX gbc1c ( \42218_nGbc1c , \42216_nGbc1a , \42217_nGbc1b , \42120 );
not \U$36429 ( \42219 , \42218_nGbc1c );
_HMUX gbc1d ( \42220_nGbc1d , RIe548ff0_6844 , \7089 , \7279 );
_HMUX gbc1e ( \42221_nGbc1e , RIe548ff0_6844 , \7284 , \9370 );
_HMUX gbc1f ( \42222_nGbc1f , \42220_nGbc1d , \42221_nGbc1e , \9381 );
_HMUX gbc20 ( \42223_nGbc20 , \42222_nGbc1f , \9394 , \9571 );
_HMUX gbc21 ( \42224_nGbc21 , \42222_nGbc1f , \9576 , \11438 );
_HMUX gbc22 ( \42225_nGbc22 , \42223_nGbc20 , \42224_nGbc21 , \11449 );
_HMUX gbc23 ( \42226_nGbc23 , \42225_nGbc22 , \11464 , \11660 );
_HMUX gbc24 ( \42227_nGbc24 , \42225_nGbc22 , \11665 , \13527 );
_HMUX gbc25 ( \42228_nGbc25 , \42226_nGbc23 , \42227_nGbc24 , \13538 );
_HMUX gbc26 ( \42229_nGbc26 , \42228_nGbc25 , \13549 , \13763 );
_HMUX gbc27 ( \42230_nGbc27 , \42228_nGbc25 , \13768 , \15630 );
_HMUX gbc28 ( \42231_nGbc28 , \42229_nGbc26 , \42230_nGbc27 , \15641 );
_HMUX gbc29 ( \42232_nGbc29 , \42231_nGbc28 , \15656 , \15889 );
_HMUX gbc2a ( \42233_nGbc2a , \42231_nGbc28 , \15894 , \17756 );
_HMUX gbc2b ( \42234_nGbc2b , \42232_nGbc29 , \42233_nGbc2a , \17767 );
_HMUX gbc2c ( \42235_nGbc2c , \42234_nGbc2b , \17780 , \18031 );
_HMUX gbc2d ( \42236_nGbc2d , \42234_nGbc2b , \18036 , \19898 );
_HMUX gbc2e ( \42237_nGbc2e , \42235_nGbc2c , \42236_nGbc2d , \19909 );
_HMUX gbc2f ( \42238_nGbc2f , \42237_nGbc2e , \19924 , \20193 );
_HMUX gbc30 ( \42239_nGbc30 , \42237_nGbc2e , \20198 , \22060 );
_HMUX gbc31 ( \42240_nGbc31 , \42238_nGbc2f , \42239_nGbc30 , \22071 );
_HMUX gbc32 ( \42241_nGbc32 , \42240_nGbc31 , \22081 , \22367 );
_HMUX gbc33 ( \42242_nGbc33 , \42240_nGbc31 , \22372 , \24234 );
_HMUX gbc34 ( \42243_nGbc34 , \42241_nGbc32 , \42242_nGbc33 , \24245 );
_HMUX gbc35 ( \42244_nGbc35 , \42243_nGbc34 , \24260 , \24565 );
_HMUX gbc36 ( \42245_nGbc36 , \42243_nGbc34 , \24570 , \26432 );
_HMUX gbc37 ( \42246_nGbc37 , \42244_nGbc35 , \42245_nGbc36 , \26443 );
_HMUX gbc38 ( \42247_nGbc38 , \42246_nGbc37 , \26456 , \26779 );
_HMUX gbc39 ( \42248_nGbc39 , \42246_nGbc37 , \26784 , \28646 );
_HMUX gbc3a ( \42249_nGbc3a , \42247_nGbc38 , \42248_nGbc39 , \28657 );
_HMUX gbc3b ( \42250_nGbc3b , \42249_nGbc3a , \28672 , \29013 );
_HMUX gbc3c ( \42251_nGbc3c , \42249_nGbc3a , \29018 , \30880 );
_HMUX gbc3d ( \42252_nGbc3d , \42250_nGbc3b , \42251_nGbc3c , \30891 );
_HMUX gbc3e ( \42253_nGbc3e , \42252_nGbc3d , \30902 , \31261 );
_HMUX gbc3f ( \42254_nGbc3f , \42252_nGbc3d , \31266 , \33128 );
_HMUX gbc40 ( \42255_nGbc40 , \42253_nGbc3e , \42254_nGbc3f , \33139 );
_HMUX gbc41 ( \42256_nGbc41 , \42255_nGbc40 , \33154 , \33531 );
_HMUX gbc42 ( \42257_nGbc42 , \42255_nGbc40 , \33536 , \35398 );
_HMUX gbc43 ( \42258_nGbc43 , \42256_nGbc41 , \42257_nGbc42 , \35409 );
_HMUX gbc44 ( \42259_nGbc44 , \42258_nGbc43 , \35422 , \35817 );
_HMUX gbc45 ( \42260_nGbc45 , \42258_nGbc43 , \35822 , \37684 );
_HMUX gbc46 ( \42261_nGbc46 , \42259_nGbc44 , \42260_nGbc45 , \37695 );
_HMUX gbc47 ( \42262_nGbc47 , \42261_nGbc46 , \37710 , \38123 );
_HMUX gbc48 ( \42263_nGbc48 , \42261_nGbc46 , \38128 , \39990 );
_HMUX gbc49 ( \42264_nGbc49 , \42262_nGbc47 , \42263_nGbc48 , \40001 );
_HMUX gbc4a ( \42265_nGbc4a , \42264_nGbc49 , RIe548ff0_6844 , \40410 );
_HMUX gbc4b ( \42266_nGbc4b , \42264_nGbc49 , \40422 , \42111 );
_HMUX gbc4c ( \42267_nGbc4c , \42265_nGbc4a , \42266_nGbc4b , \42120 );
_HMUX gbc4d ( \42268_nGbc4d , RIea91330_6888 , \7093 , \7279 );
_HMUX gbc4e ( \42269_nGbc4e , RIea91330_6888 , \7287 , \9370 );
_HMUX gbc4f ( \42270_nGbc4f , \42268_nGbc4d , \42269_nGbc4e , \9381 );
_HMUX gbc50 ( \42271_nGbc50 , \42270_nGbc4f , \9398 , \9571 );
_HMUX gbc51 ( \42272_nGbc51 , \42270_nGbc4f , \9579 , \11438 );
_HMUX gbc52 ( \42273_nGbc52 , \42271_nGbc50 , \42272_nGbc51 , \11449 );
_HMUX gbc53 ( \42274_nGbc53 , \42273_nGbc52 , \11468 , \11660 );
_HMUX gbc54 ( \42275_nGbc54 , \42273_nGbc52 , \11668 , \13527 );
_HMUX gbc55 ( \42276_nGbc55 , \42274_nGbc53 , \42275_nGbc54 , \13538 );
_HMUX gbc56 ( \42277_nGbc56 , \42276_nGbc55 , \13553 , \13763 );
_HMUX gbc57 ( \42278_nGbc57 , \42276_nGbc55 , \13771 , \15630 );
_HMUX gbc58 ( \42279_nGbc58 , \42277_nGbc56 , \42278_nGbc57 , \15641 );
_HMUX gbc59 ( \42280_nGbc59 , \42279_nGbc58 , \15660 , \15889 );
_HMUX gbc5a ( \42281_nGbc5a , \42279_nGbc58 , \15897 , \17756 );
_HMUX gbc5b ( \42282_nGbc5b , \42280_nGbc59 , \42281_nGbc5a , \17767 );
_HMUX gbc5c ( \42283_nGbc5c , \42282_nGbc5b , \17784 , \18031 );
_HMUX gbc5d ( \42284_nGbc5d , \42282_nGbc5b , \18039 , \19898 );
_HMUX gbc5e ( \42285_nGbc5e , \42283_nGbc5c , \42284_nGbc5d , \19909 );
_HMUX gbc5f ( \42286_nGbc5f , \42285_nGbc5e , \19928 , \20193 );
_HMUX gbc60 ( \42287_nGbc60 , \42285_nGbc5e , \20201 , \22060 );
_HMUX gbc61 ( \42288_nGbc61 , \42286_nGbc5f , \42287_nGbc60 , \22071 );
_HMUX gbc62 ( \42289_nGbc62 , \42288_nGbc61 , \22084 , \22367 );
_HMUX gbc63 ( \42290_nGbc63 , \42288_nGbc61 , \22375 , \24234 );
_HMUX gbc64 ( \42291_nGbc64 , \42289_nGbc62 , \42290_nGbc63 , \24245 );
_HMUX gbc65 ( \42292_nGbc65 , \42291_nGbc64 , \24264 , \24565 );
_HMUX gbc66 ( \42293_nGbc66 , \42291_nGbc64 , \24573 , \26432 );
_HMUX gbc67 ( \42294_nGbc67 , \42292_nGbc65 , \42293_nGbc66 , \26443 );
_HMUX gbc68 ( \42295_nGbc68 , \42294_nGbc67 , \26460 , \26779 );
_HMUX gbc69 ( \42296_nGbc69 , \42294_nGbc67 , \26787 , \28646 );
_HMUX gbc6a ( \42297_nGbc6a , \42295_nGbc68 , \42296_nGbc69 , \28657 );
_HMUX gbc6b ( \42298_nGbc6b , \42297_nGbc6a , \28676 , \29013 );
_HMUX gbc6c ( \42299_nGbc6c , \42297_nGbc6a , \29021 , \30880 );
_HMUX gbc6d ( \42300_nGbc6d , \42298_nGbc6b , \42299_nGbc6c , \30891 );
_HMUX gbc6e ( \42301_nGbc6e , \42300_nGbc6d , \30906 , \31261 );
_HMUX gbc6f ( \42302_nGbc6f , \42300_nGbc6d , \31269 , \33128 );
_HMUX gbc70 ( \42303_nGbc70 , \42301_nGbc6e , \42302_nGbc6f , \33139 );
_HMUX gbc71 ( \42304_nGbc71 , \42303_nGbc70 , \33158 , \33531 );
_HMUX gbc72 ( \42305_nGbc72 , \42303_nGbc70 , \33539 , \35398 );
_HMUX gbc73 ( \42306_nGbc73 , \42304_nGbc71 , \42305_nGbc72 , \35409 );
_HMUX gbc74 ( \42307_nGbc74 , \42306_nGbc73 , \35426 , \35817 );
_HMUX gbc75 ( \42308_nGbc75 , \42306_nGbc73 , \35825 , \37684 );
_HMUX gbc76 ( \42309_nGbc76 , \42307_nGbc74 , \42308_nGbc75 , \37695 );
_HMUX gbc77 ( \42310_nGbc77 , \42309_nGbc76 , \37714 , \38123 );
_HMUX gbc78 ( \42311_nGbc78 , \42309_nGbc76 , \38131 , \39990 );
_HMUX gbc79 ( \42312_nGbc79 , \42310_nGbc77 , \42311_nGbc78 , \40001 );
_HMUX gbc7a ( \42313_nGbc7a , \42312_nGbc79 , RIea91330_6888 , \40410 );
_HMUX gbc7b ( \42314_nGbc7b , \42312_nGbc79 , \40426 , \42111 );
_HMUX gbc7c ( \42315_nGbc7c , \42313_nGbc7a , \42314_nGbc7b , \42120 );
not \U$36430 ( \42316 , \42315_nGbc7c );
and \U$36431 ( \42317 , \42121_nGbbbc , \42170 , \42219 , \42267_nGbc4c , \42316 );
buf \U$36432 ( \42318 , \42317 );
and \U$36433 ( \42319 , \7075 , \42318 );
_HMUX g1489b ( \42320_nG1489b , \7068_nG14891 , \7074_nG14897 , \42319 );
and \U$36434 ( \42321 , \42319 , \7066 );
and \U$36435 ( \42322 , \42321 , \7065 );
_HMUX g1489e ( \42323_nG1489e , \42320_nG1489b , RIde67cd8_3982 , \42322 );
not \U$36436 ( \42324 , RIde4ec88_4006);
buf \U$36437 ( \42325 , RIb7b9680_245);
and \U$36438 ( \42326 , RIde4ec88_4006, \42325 );
or \U$36439 ( \42327 , \42324 , \42326 );
and \U$36440 ( \42328 , \42327 , \7075 );
and \U$36441 ( \42329 , \42328 , \42318 );
_HMUX g148a5 ( \42330_nG148a5 , \42323_nG1489e , RIde5fec0_3994 , \42329 );
buf \U$36443 ( \42331 , RIb79b338_274);
and \U$36444 ( \42332 , \7065 , \42331 );
_HMUX g148a6 ( \42333_nG148a6 , \42330_nG148a5 , 1'b0 , \42332 );
buf \U$36445 ( \42334 , \42333_nG148a6 );
buf \U$36446 ( \42335 , RIde68638_3981);
xnor \U$36447 ( \42336 , \42335 , \7056 );
buf \U$36448 ( \42337 , \42336 );
_HMUX g148aa ( \42338_nG148aa , \42337 , 1'b0 , \7059 );
_HMUX g148ab ( \42339_nG148ab , RIde68638_3981 , \42338_nG148aa , \7067 );
buf \U$36450 ( \42340 , RIde68638_3981);
xor \U$36451 ( \42341 , \42340 , \7069 );
buf \U$36452 ( \42342 , \42341 );
_HMUX g148af ( \42343_nG148af , \42342 , RIde68638_3981 , \7073 );
_HMUX g148b0 ( \42344_nG148b0 , \42339_nG148ab , \42343_nG148af , \42319 );
_HMUX g148b1 ( \42345_nG148b1 , \42344_nG148b0 , RIde68638_3981 , \42322 );
_HMUX g148b2 ( \42346_nG148b2 , \42345_nG148b1 , RIde60988_3993 , \42329 );
_HMUX g148b3 ( \42347_nG148b3 , \42346_nG148b2 , 1'b0 , \42332 );
buf \U$36454 ( \42348 , \42347_nG148b3 );
buf \U$36455 ( \42349 , RIde68f20_3980);
or \U$36456 ( \42350 , \42335 , \7056 );
xnor \U$36457 ( \42351 , \42349 , \42350 );
buf \U$36458 ( \42352 , \42351 );
_HMUX g148b8 ( \42353_nG148b8 , \42352 , 1'b0 , \7059 );
_HMUX g148b9 ( \42354_nG148b9 , RIde68f20_3980 , \42353_nG148b8 , \7067 );
buf \U$36460 ( \42355 , RIde68f20_3980);
and \U$36461 ( \42356 , \42340 , \7069 );
xor \U$36462 ( \42357 , \42355 , \42356 );
buf \U$36463 ( \42358 , \42357 );
_HMUX g148be ( \42359_nG148be , \42358 , RIde68f20_3980 , \7073 );
_HMUX g148bf ( \42360_nG148bf , \42354_nG148b9 , \42359_nG148be , \42319 );
_HMUX g148c0 ( \42361_nG148c0 , \42360_nG148bf , RIde68f20_3980 , \42322 );
_HMUX g148c1 ( \42362_nG148c1 , \42361_nG148c0 , RIde612e8_3992 , \42329 );
_HMUX g148c2 ( \42363_nG148c2 , \42362_nG148c1 , 1'b0 , \42332 );
buf \U$36465 ( \42364 , \42363_nG148c2 );
or \U$36466 ( \42365 , \42334 , \42348 , \42364 );
buf \U$36467 ( \42366 , \42365 );
buf \U$36468 ( \42367 , RIde6ad98_3977);
buf \U$36469 ( \42368 , RIde6a2d0_3978);
buf \U$36470 ( \42369 , RIde69970_3979);
and \U$36471 ( \42370 , \42368 , \42369 );
xor \U$36472 ( \42371 , \42367 , \42370 );
buf \U$36473 ( \42372 , \42371 );
not \U$36474 ( \42373 , RIde6ad98_3977);
nor \U$36475 ( \42374 , RIde69970_3979, RIde6a2d0_3978, \42373 );
not \U$36476 ( \42375 , \42374 );
and \U$36477 ( \42376 , \7067 , \42375 );
_HMUX g14887 ( \42377_nG14887 , RIde6ad98_3977 , \42372 , \42376 );
_HMUX g14888 ( \42378_nG14888 , \42377_nG14887 , 1'b0 , \42332 );
buf \U$36479 ( \42379 , \42378_nG14888 );
not \U$36480 ( \42380 , \42379 );
buf \U$36481 ( \42381 , RIde63250_3989);
buf \U$36482 ( \42382 , RIde62878_3990);
buf \U$36483 ( \42383 , RIde61e28_3991);
and \U$36484 ( \42384 , \42382 , \42383 );
xor \U$36485 ( \42385 , \42381 , \42384 );
buf \U$36486 ( \42386 , \42385 );
not \U$36487 ( \42387 , RIe546890_6849);
not \U$36488 ( \42388 , RIe546098_6850);
not \U$36489 ( \42389 , RIe545648_6852);
and \U$36490 ( \42390 , RIea90778_6887, \42387 , \42388 , RIe545dc8_6851, \42389 );
buf \U$36491 ( \42391 , \42390 );
buf \U$36492 ( \42392 , RIb839848_152);
and \U$36493 ( \42393 , \42391 , \42392 );
not \U$36494 ( \42394 , RIde62878_3990);
and \U$36495 ( \42395 , RIde61e28_3991, \42394 , RIde63250_3989);
not \U$36496 ( \42396 , \42395 );
and \U$36497 ( \42397 , \42393 , \42396 );
_HMUX g14945 ( \42398_nG14945 , RIde63250_3989 , \42386 , \42397 );
buf \U$36498 ( \42399 , RIde63250_3989);
buf \U$36499 ( \42400 , RIde62878_3990);
xor \U$36500 ( \42401 , \42399 , \42400 );
buf \U$36501 ( \42402 , \42401 );
not \U$36502 ( \42403 , RIde61e28_3991);
and \U$36503 ( \42404 , \42403 , \42394 , RIde63250_3989);
or \U$36504 ( \42405 , \42404 , \42395 );
_HMUX g14949 ( \42406_nG14949 , \42402 , RIde63250_3989 , \42405 );
buf \U$36505 ( \42407 , RIb839668_156);
and \U$36506 ( \42408 , \42391 , \42407 );
_HMUX g1494a ( \42409_nG1494a , \42398_nG14945 , \42406_nG14949 , \42408 );
buf \U$36508 ( \42410 , RIb8396e0_155);
and \U$36509 ( \42411 , \42391 , \42410 );
_HMUX g1494b ( \42412_nG1494b , \42409_nG1494a , 1'b0 , \42411 );
and \U$36511 ( \42413 , \42411 , \42407 );
_HMUX g1494c ( \42414_nG1494c , \42412_nG1494b , 1'b0 , \42413 );
buf \U$36512 ( \42415 , \42414_nG1494c );
and \U$36513 ( \42416 , \42380 , \42415 );
xor \U$36514 ( \42417 , \42368 , \42369 );
buf \U$36515 ( \42418 , \42417 );
_HMUX g14881 ( \42419_nG14881 , RIde6a2d0_3978 , \42418 , \42376 );
_HMUX g14882 ( \42420_nG14882 , \42419_nG14881 , 1'b0 , \42332 );
buf \U$36517 ( \42421 , \42420_nG14882 );
not \U$36518 ( \42422 , \42421 );
xor \U$36519 ( \42423 , \42382 , \42383 );
buf \U$36520 ( \42424 , \42423 );
_HMUX g14936 ( \42425_nG14936 , RIde62878_3990 , \42424 , \42397 );
not \U$36521 ( \42426 , \42400 );
buf \U$36522 ( \42427 , \42426 );
_HMUX g1493d ( \42428_nG1493d , \42427 , RIde62878_3990 , \42405 );
_HMUX g1493e ( \42429_nG1493e , \42425_nG14936 , \42428_nG1493d , \42408 );
_HMUX g1493f ( \42430_nG1493f , \42429_nG1493e , 1'b0 , \42411 );
_HMUX g14940 ( \42431_nG14940 , \42430_nG1493f , 1'b1 , \42413 );
buf \U$36525 ( \42432 , \42431_nG14940 );
and \U$36526 ( \42433 , \42422 , \42432 );
not \U$36527 ( \42434 , \42369 );
buf \U$36528 ( \42435 , \42434 );
_HMUX g1487a ( \42436_nG1487a , RIde69970_3979 , \42435 , \42376 );
_HMUX g1487d ( \42437_nG1487d , \42436_nG1487a , 1'b0 , \42332 );
buf \U$36530 ( \42438 , \42437_nG1487d );
not \U$36531 ( \42439 , \42438 );
not \U$36532 ( \42440 , \42383 );
buf \U$36533 ( \42441 , \42440 );
_HMUX g14926 ( \42442_nG14926 , RIde61e28_3991 , \42441 , \42397 );
buf \U$36534 ( \42443 , RIde61e28_3991);
buf g1492a( \42444_nG1492a , \42443 );
_HMUX g1492d ( \42445_nG1492d , \42442_nG14926 , \42444_nG1492a , \42408 );
_HMUX g14930 ( \42446_nG14930 , \42445_nG1492d , 1'b1 , \42411 );
_HMUX g14932 ( \42447_nG14932 , \42446_nG14930 , 1'b0 , \42413 );
buf \U$36539 ( \42448 , \42447_nG14932 );
and \U$36540 ( \42449 , \42439 , \42448 );
xnor \U$36541 ( \42450 , \42432 , \42421 );
and \U$36542 ( \42451 , \42449 , \42450 );
or \U$36543 ( \42452 , \42433 , \42451 );
xnor \U$36544 ( \42453 , \42415 , \42379 );
and \U$36545 ( \42454 , \42452 , \42453 );
or \U$36546 ( \42455 , \42416 , \42454 );
buf \U$36547 ( \42456 , \42455 );
and \U$36548 ( \42457 , \42366 , \42456 );
buf \U$36550 ( \42458 , RIb79b3b0_273);
and \U$36551 ( \42459 , \42318 , \42458 );
_HMUX g149bd ( \42460_nG149bd , RIde5f3f8_3995 , \42325 , \42459 );
not \U$36552 ( \42461 , \42460_nG149bd );
or \U$36553 ( \42462 , \42461 , \42324 );
and \U$36554 ( \42463 , \42366 , \42462 );
_HMUX g149c1 ( \42464_nG149c1 , \42457 , 1'b1 , \42463 );
buf \U$36555 ( \42465 , \42464_nG149c1 );
not \U$36556 ( \42466 , RIe5319e0_6884);
nor \U$36557 ( \42467 , \42466 , RIe549ef0_6842, RIe549770_6843, RIe548ff0_6844, RIea91330_6888);
not \U$36558 ( \42468 , RIe549ef0_6842);
nor \U$36559 ( \42469 , RIe5319e0_6884, \42468 , RIe549770_6843, RIe548ff0_6844, RIea91330_6888);
or \U$36560 ( \42470 , \42467 , \42469 );
nor \U$36561 ( \42471 , \42466 , \42468 , RIe549770_6843, RIe548ff0_6844, RIea91330_6888);
or \U$36562 ( \42472 , \42470 , \42471 );
not \U$36563 ( \42473 , RIe548ff0_6844);
not \U$36564 ( \42474 , RIea91330_6888);
and \U$36565 ( \42475 , \42466 , \42468 , RIe549770_6843, \42473 , \42474 );
or \U$36566 ( \42476 , \42472 , \42475 );
and \U$36567 ( \42477 , RIe5319e0_6884, \42468 , RIe549770_6843, \42473 , \42474 );
or \U$36568 ( \42478 , \42476 , \42477 );
and \U$36569 ( \42479 , \42466 , RIe549ef0_6842, RIe549770_6843, \42473 , \42474 );
or \U$36570 ( \42480 , \42478 , \42479 );
and \U$36571 ( \42481 , RIe5319e0_6884, RIe549ef0_6842, RIe549770_6843, \42473 , \42474 );
or \U$36572 ( \42482 , \42480 , \42481 );
nor \U$36573 ( \42483 , RIe5319e0_6884, RIe549ef0_6842, RIe549770_6843, \42473 , RIea91330_6888);
or \U$36574 ( \42484 , \42482 , \42483 );
nor \U$36575 ( \42485 , \42466 , RIe549ef0_6842, RIe549770_6843, \42473 , RIea91330_6888);
or \U$36576 ( \42486 , \42484 , \42485 );
nor \U$36577 ( \42487 , RIe5319e0_6884, \42468 , RIe549770_6843, \42473 , RIea91330_6888);
or \U$36578 ( \42488 , \42486 , \42487 );
nor \U$36579 ( \42489 , \42466 , \42468 , RIe549770_6843, \42473 , RIea91330_6888);
or \U$36580 ( \42490 , \42488 , \42489 );
and \U$36581 ( \42491 , \42466 , \42468 , RIe549770_6843, RIe548ff0_6844, \42474 );
or \U$36582 ( \42492 , \42490 , \42491 );
and \U$36583 ( \42493 , RIe5319e0_6884, \42468 , RIe549770_6843, RIe548ff0_6844, \42474 );
or \U$36584 ( \42494 , \42492 , \42493 );
and \U$36585 ( \42495 , \42466 , RIe549ef0_6842, RIe549770_6843, RIe548ff0_6844, \42474 );
or \U$36586 ( \42496 , \42494 , \42495 );
and \U$36587 ( \42497 , RIe5319e0_6884, RIe549ef0_6842, RIe549770_6843, RIe548ff0_6844, \42474 );
or \U$36588 ( \42498 , \42496 , \42497 );
nor \U$36589 ( \42499 , RIe5319e0_6884, RIe549ef0_6842, RIe549770_6843, RIe548ff0_6844, \42474 );
or \U$36590 ( \42500 , \42498 , \42499 );
buf \U$36591 ( \42501 , \42500 );
not \U$36592 ( \42502 , \42501 );
buf \U$36593 ( \42503 , \42502 );
_DC g1a9a6_GF_IsGateDCbyConstraint ( \42504_nG1a9a6 , \42465 , \42503 );
buf \U$36594 ( \42505 , \42504_nG1a9a6 );
buf \U$36595 ( \42506 , \42333_nG148a6 );
_DC g1abf3_GF_IsGateDCbyConstraint ( \42507_nG1abf3 , \42506 , \42503 );
buf \U$36596 ( \42508 , \42507_nG1abf3 );
buf \U$36597 ( \42509 , \42347_nG148b3 );
_DC g1abf4_GF_IsGateDCbyConstraint ( \42510_nG1abf4 , \42509 , \42503 );
buf \U$36598 ( \42511 , \42510_nG1abf4 );
buf \U$36599 ( \42512 , \42363_nG148c2 );
_DC g1abf5_GF_IsGateDCbyConstraint ( \42513_nG1abf5 , \42512 , \42503 );
buf \U$36600 ( \42514 , \42513_nG1abf5 );
buf \U$36601 ( \42515 , \42460_nG149bd );
_DC g1abef_GF_IsGateDCbyConstraint ( \42516_nG1abef , \42515 , \42503 );
buf \U$36602 ( \42517 , \42516_nG1abef );
buf \U$36603 ( \42518 , RIb7b96f8_244);
_HMUX g14a2a ( \42519_nG14a2a , RIde4c8e8_4009 , \42518 , \42459 );
buf \U$36604 ( \42520 , \42519_nG14a2a );
_DC g1a98c_GF_IsGateDCbyConstraint ( \42521_nG1a98c , \42520 , \42503 );
buf \U$36605 ( \42522 , \42521_nG1a98c );
buf \U$36606 ( \42523 , RIb7c20c8_243);
_HMUX g14a2c ( \42524_nG14a2c , RIde4d6f8_4008 , \42523 , \42459 );
buf \U$36607 ( \42525 , \42524_nG14a2c );
_DC g1a98e_GF_IsGateDCbyConstraint ( \42526_nG1a98e , \42525 , \42503 );
buf \U$36608 ( \42527 , \42526_nG1a98e );
buf \U$36609 ( \42528 , RIb7c5728_242);
_HMUX g14a2e ( \42529_nG14a2e , RIde431f8_4020 , \42528 , \42459 );
buf \U$36610 ( \42530 , \42529_nG14a2e );
_DC g1a990_GF_IsGateDCbyConstraint ( \42531_nG1a990 , \42530 , \42503 );
buf \U$36611 ( \42532 , \42531_nG1a990 );
buf \U$36612 ( \42533 , RIb7c57a0_241);
_HMUX g14a30 ( \42534_nG14a30 , RIde43f90_4019 , \42533 , \42459 );
buf \U$36613 ( \42535 , \42534_nG14a30 );
_DC g1a992_GF_IsGateDCbyConstraint ( \42536_nG1a992 , \42535 , \42503 );
buf \U$36614 ( \42537 , \42536_nG1a992 );
buf \U$36615 ( \42538 , RIb7c5818_240);
_HMUX g14a32 ( \42539_nG14a32 , RIde44da0_4018 , \42538 , \42459 );
buf \U$36616 ( \42540 , \42539_nG14a32 );
_DC g1a994_GF_IsGateDCbyConstraint ( \42541_nG1a994 , \42540 , \42503 );
buf \U$36617 ( \42542 , \42541_nG1a994 );
buf \U$36618 ( \42543 , RIb7c5890_239);
_HMUX g14a34 ( \42544_nG14a34 , RIde45ac0_4017 , \42543 , \42459 );
buf \U$36619 ( \42545 , \42544_nG14a34 );
_DC g1a996_GF_IsGateDCbyConstraint ( \42546_nG1a996 , \42545 , \42503 );
buf \U$36620 ( \42547 , \42546_nG1a996 );
buf \U$36621 ( \42548 , RIb7c5908_238);
_HMUX g14a36 ( \42549_nG14a36 , RIde468d0_4016 , \42548 , \42459 );
buf \U$36622 ( \42550 , \42549_nG14a36 );
_DC g1a998_GF_IsGateDCbyConstraint ( \42551_nG1a998 , \42550 , \42503 );
buf \U$36623 ( \42552 , \42551_nG1a998 );
buf \U$36624 ( \42553 , RIb7a09f0_266);
_HMUX g14a28 ( \42554_nG14a28 , RIde4fb10_4005 , \42553 , \42459 );
buf \U$36625 ( \42555 , \42554_nG14a28 );
_DC g1a98a_GF_IsGateDCbyConstraint ( \42556_nG1a98a , \42555 , \42503 );
buf \U$36626 ( \42557 , \42556_nG1a98a );
buf \U$36627 ( \42558 , RIb7a0a68_265);
_HMUX g14a20 ( \42559_nG14a20 , RIde49300_4013 , \42558 , \42459 );
buf \U$36628 ( \42560 , \42559_nG14a20 );
_DC g1a982_GF_IsGateDCbyConstraint ( \42561_nG1a982 , \42560 , \42503 );
buf \U$36629 ( \42562 , \42561_nG1a982 );
buf \U$36630 ( \42563 , RIb7a0ae0_264);
_HMUX g14a22 ( \42564_nG14a22 , RIde4a020_4012 , \42563 , \42459 );
buf \U$36631 ( \42565 , \42564_nG14a22 );
_DC g1a984_GF_IsGateDCbyConstraint ( \42566_nG1a984 , \42565 , \42503 );
buf \U$36632 ( \42567 , \42566_nG1a984 );
buf \U$36633 ( \42568 , RIb7a0b58_263);
_HMUX g14a24 ( \42569_nG14a24 , RIde4ae30_4011 , \42568 , \42459 );
buf \U$36634 ( \42570 , \42569_nG14a24 );
_DC g1a986_GF_IsGateDCbyConstraint ( \42571_nG1a986 , \42570 , \42503 );
buf \U$36635 ( \42572 , \42571_nG1a986 );
buf \U$36636 ( \42573 , RIb7a0bd0_262);
_HMUX g14a26 ( \42574_nG14a26 , RIde4bb50_4010 , \42573 , \42459 );
buf \U$36637 ( \42575 , \42574_nG14a26 );
_DC g1a988_GF_IsGateDCbyConstraint ( \42576_nG1a988 , \42575 , \42503 );
buf \U$36638 ( \42577 , \42576_nG1a988 );
buf \U$36639 ( \42578 , RIb87eb00_69);
buf \U$36640 ( \42579 , RIe667bb0_6885);
buf \U$36641 ( \42580 , RIe667f70_6886);
nor \U$36642 ( \42581 , \42579 , \42580 );
_HMUX g14ebe ( \42582_nG14ebe , RIdbee210_3713 , \42578 , \42581 );
buf \U$36643 ( \42583 , \42391 );
not \U$36644 ( \42584 , RIb839b90_145);
and \U$36645 ( \42585 , RIb839848_152, \42584 );
and \U$36646 ( \42586 , RIb8396e0_155, RIb839b90_145);
or \U$36647 ( \42587 , \42585 , \42586 );
buf \U$36648 ( \42588 , \42587 );
buf \U$36649 ( \42589 , \42588 );
and \U$36650 ( \42590 , \42583 , \42589 );
_HMUX g14ebf ( \42591_nG14ebf , RIdbee210_3713 , \42582_nG14ebe , \42590 );
buf \U$36651 ( \42592 , RIb7c5980_237);
buf \U$36652 ( \42593 , RIeab7058_6894);
buf \U$36653 ( \42594 , RIea91768_6889);
nor \U$36654 ( \42595 , \42593 , \42594 );
_HMUX g14ec1 ( \42596_nG14ec1 , RIdbee210_3713 , \42592 , \42595 );
buf \U$36655 ( \42597 , \42318 );
buf \U$36656 ( \42598 , \7075 );
and \U$36657 ( \42599 , \42597 , \42598 );
_HMUX g14ec2 ( \42600_nG14ec2 , \42591_nG14ebf , \42596_nG14ec1 , \42599 );
buf \U$36658 ( \42601 , \42600_nG14ec2 );
_DC g1ab60_GF_IsGateDCbyConstraint ( \42602_nG1ab60 , \42601 , \42503 );
buf \U$36659 ( \42603 , \42602_nG1ab60 );
buf \U$36660 ( \42604 , RIb87eb78_68);
_HMUX g14ec3 ( \42605_nG14ec3 , RIdbecc08_3714 , \42604 , \42581 );
_HMUX g14ec4 ( \42606_nG14ec4 , RIdbecc08_3714 , \42605_nG14ec3 , \42590 );
buf \U$36661 ( \42607 , RIb7c59f8_236);
_HMUX g14ec5 ( \42608_nG14ec5 , RIdbecc08_3714 , \42607 , \42595 );
_HMUX g14ec6 ( \42609_nG14ec6 , \42606_nG14ec4 , \42608_nG14ec5 , \42599 );
buf \U$36662 ( \42610 , \42609_nG14ec6 );
_DC g1ab76_GF_IsGateDCbyConstraint ( \42611_nG1ab76 , \42610 , \42503 );
buf \U$36663 ( \42612 , \42611_nG1ab76 );
buf \U$36664 ( \42613 , RIb87ebf0_67);
_HMUX g14ec7 ( \42614_nG14ec7 , RIdbebab0_3715 , \42613 , \42581 );
_HMUX g14ec8 ( \42615_nG14ec8 , RIdbebab0_3715 , \42614_nG14ec7 , \42590 );
buf \U$36665 ( \42616 , RIb7c5a70_235);
_HMUX g14ec9 ( \42617_nG14ec9 , RIdbebab0_3715 , \42616 , \42595 );
_HMUX g14eca ( \42618_nG14eca , \42615_nG14ec8 , \42617_nG14ec9 , \42599 );
buf \U$36666 ( \42619 , \42618_nG14eca );
_DC g1ab8c_GF_IsGateDCbyConstraint ( \42620_nG1ab8c , \42619 , \42503 );
buf \U$36667 ( \42621 , \42620_nG1ab8c );
buf \U$36668 ( \42622 , RIb882ca0_66);
_HMUX g14ecb ( \42623_nG14ecb , RIdbea4a8_3716 , \42622 , \42581 );
_HMUX g14ecc ( \42624_nG14ecc , RIdbea4a8_3716 , \42623_nG14ecb , \42590 );
buf \U$36669 ( \42625 , RIb7cade0_234);
_HMUX g14ecd ( \42626_nG14ecd , RIdbea4a8_3716 , \42625 , \42595 );
_HMUX g14ece ( \42627_nG14ece , \42624_nG14ecc , \42626_nG14ecd , \42599 );
buf \U$36670 ( \42628 , \42627_nG14ece );
_DC g1aba2_GF_IsGateDCbyConstraint ( \42629_nG1aba2 , \42628 , \42503 );
buf \U$36671 ( \42630 , \42629_nG1aba2 );
buf \U$36672 ( \42631 , RIb885310_65);
_HMUX g14ecf ( \42632_nG14ecf , RIdbe9350_3717 , \42631 , \42581 );
_HMUX g14ed0 ( \42633_nG14ed0 , RIdbe9350_3717 , \42632_nG14ecf , \42590 );
buf \U$36673 ( \42634 , RIb7cae58_233);
_HMUX g14ed1 ( \42635_nG14ed1 , RIdbe9350_3717 , \42634 , \42595 );
_HMUX g14ed2 ( \42636_nG14ed2 , \42633_nG14ed0 , \42635_nG14ed1 , \42599 );
buf \U$36674 ( \42637 , \42636_nG14ed2 );
_DC g1abb8_GF_IsGateDCbyConstraint ( \42638_nG1abb8 , \42637 , \42503 );
buf \U$36675 ( \42639 , \42638_nG1abb8 );
buf \U$36676 ( \42640 , RIb885388_64);
_HMUX g14ed3 ( \42641_nG14ed3 , RIdbe7d48_3718 , \42640 , \42581 );
_HMUX g14ed4 ( \42642_nG14ed4 , RIdbe7d48_3718 , \42641_nG14ed3 , \42590 );
buf \U$36677 ( \42643 , RIb7caed0_232);
_HMUX g14ed5 ( \42644_nG14ed5 , RIdbe7d48_3718 , \42643 , \42595 );
_HMUX g14ed6 ( \42645_nG14ed6 , \42642_nG14ed4 , \42644_nG14ed5 , \42599 );
buf \U$36678 ( \42646 , \42645_nG14ed6 );
_DC g1abce_GF_IsGateDCbyConstraint ( \42647_nG1abce , \42646 , \42503 );
buf \U$36679 ( \42648 , \42647_nG1abce );
buf \U$36680 ( \42649 , RIb885400_63);
_HMUX g14ed7 ( \42650_nG14ed7 , RIdbe6bf0_3719 , \42649 , \42581 );
_HMUX g14ed8 ( \42651_nG14ed8 , RIdbe6bf0_3719 , \42650_nG14ed7 , \42590 );
buf \U$36681 ( \42652 , RIb7caf48_231);
_HMUX g14ed9 ( \42653_nG14ed9 , RIdbe6bf0_3719 , \42652 , \42595 );
_HMUX g14eda ( \42654_nG14eda , \42651_nG14ed8 , \42653_nG14ed9 , \42599 );
buf \U$36682 ( \42655 , \42654_nG14eda );
_DC g1abda_GF_IsGateDCbyConstraint ( \42656_nG1abda , \42655 , \42503 );
buf \U$36683 ( \42657 , \42656_nG1abda );
buf \U$36684 ( \42658 , RIb885478_62);
_HMUX g14edb ( \42659_nG14edb , RIdbe5a98_3720 , \42658 , \42581 );
_HMUX g14edc ( \42660_nG14edc , RIdbe5a98_3720 , \42659_nG14edb , \42590 );
buf \U$36685 ( \42661 , RIb7cafc0_230);
_HMUX g14edd ( \42662_nG14edd , RIdbe5a98_3720 , \42661 , \42595 );
_HMUX g14ede ( \42663_nG14ede , \42660_nG14edc , \42662_nG14edd , \42599 );
buf \U$36686 ( \42664 , \42663_nG14ede );
_DC g1abdc_GF_IsGateDCbyConstraint ( \42665_nG1abdc , \42664 , \42503 );
buf \U$36687 ( \42666 , \42665_nG1abdc );
buf \U$36688 ( \42667 , RIb8854f0_61);
_HMUX g14edf ( \42668_nG14edf , RIdbe4490_3721 , \42667 , \42581 );
_HMUX g14ee0 ( \42669_nG14ee0 , RIdbe4490_3721 , \42668_nG14edf , \42590 );
buf \U$36689 ( \42670 , RIb7cb038_229);
_HMUX g14ee1 ( \42671_nG14ee1 , RIdbe4490_3721 , \42670 , \42595 );
_HMUX g14ee2 ( \42672_nG14ee2 , \42669_nG14ee0 , \42671_nG14ee1 , \42599 );
buf \U$36690 ( \42673 , \42672_nG14ee2 );
_DC g1abde_GF_IsGateDCbyConstraint ( \42674_nG1abde , \42673 , \42503 );
buf \U$36691 ( \42675 , \42674_nG1abde );
buf \U$36692 ( \42676 , RIb885568_60);
_HMUX g14ee3 ( \42677_nG14ee3 , RIdbe3338_3722 , \42676 , \42581 );
_HMUX g14ee4 ( \42678_nG14ee4 , RIdbe3338_3722 , \42677_nG14ee3 , \42590 );
buf \U$36693 ( \42679 , RIb7cb0b0_228);
_HMUX g14ee5 ( \42680_nG14ee5 , RIdbe3338_3722 , \42679 , \42595 );
_HMUX g14ee6 ( \42681_nG14ee6 , \42678_nG14ee4 , \42680_nG14ee5 , \42599 );
buf \U$36694 ( \42682 , \42681_nG14ee6 );
_DC g1ab62_GF_IsGateDCbyConstraint ( \42683_nG1ab62 , \42682 , \42503 );
buf \U$36695 ( \42684 , \42683_nG1ab62 );
buf \U$36696 ( \42685 , RIb8855e0_59);
_HMUX g14ee7 ( \42686_nG14ee7 , RIdbe1d30_3723 , \42685 , \42581 );
_HMUX g14ee8 ( \42687_nG14ee8 , RIdbe1d30_3723 , \42686_nG14ee7 , \42590 );
buf \U$36697 ( \42688 , RIb7cb128_227);
_HMUX g14ee9 ( \42689_nG14ee9 , RIdbe1d30_3723 , \42688 , \42595 );
_HMUX g14eea ( \42690_nG14eea , \42687_nG14ee8 , \42689_nG14ee9 , \42599 );
buf \U$36698 ( \42691 , \42690_nG14eea );
_DC g1ab64_GF_IsGateDCbyConstraint ( \42692_nG1ab64 , \42691 , \42503 );
buf \U$36699 ( \42693 , \42692_nG1ab64 );
buf \U$36700 ( \42694 , RIb885658_58);
_HMUX g14eeb ( \42695_nG14eeb , RIdbe0bd8_3724 , \42694 , \42581 );
_HMUX g14eec ( \42696_nG14eec , RIdbe0bd8_3724 , \42695_nG14eeb , \42590 );
buf \U$36701 ( \42697 , RIb7d00d8_226);
_HMUX g14eed ( \42698_nG14eed , RIdbe0bd8_3724 , \42697 , \42595 );
_HMUX g14eee ( \42699_nG14eee , \42696_nG14eec , \42698_nG14eed , \42599 );
buf \U$36702 ( \42700 , \42699_nG14eee );
_DC g1ab66_GF_IsGateDCbyConstraint ( \42701_nG1ab66 , \42700 , \42503 );
buf \U$36703 ( \42702 , \42701_nG1ab66 );
buf \U$36704 ( \42703 , RIb8856d0_57);
_HMUX g14eef ( \42704_nG14eef , RIdaab098_3725 , \42703 , \42581 );
_HMUX g14ef0 ( \42705_nG14ef0 , RIdaab098_3725 , \42704_nG14eef , \42590 );
buf \U$36705 ( \42706 , RIb8263d8_225);
_HMUX g14ef1 ( \42707_nG14ef1 , RIdaab098_3725 , \42706 , \42595 );
_HMUX g14ef2 ( \42708_nG14ef2 , \42705_nG14ef0 , \42707_nG14ef1 , \42599 );
buf \U$36706 ( \42709 , \42708_nG14ef2 );
_DC g1ab68_GF_IsGateDCbyConstraint ( \42710_nG1ab68 , \42709 , \42503 );
buf \U$36707 ( \42711 , \42710_nG1ab68 );
buf \U$36708 ( \42712 , RIb885748_56);
_HMUX g14ef3 ( \42713_nG14ef3 , RIdaaf0d0_3726 , \42712 , \42581 );
_HMUX g14ef4 ( \42714_nG14ef4 , RIdaaf0d0_3726 , \42713_nG14ef3 , \42590 );
buf \U$36709 ( \42715 , RIb826e28_224);
_HMUX g14ef5 ( \42716_nG14ef5 , RIdaaf0d0_3726 , \42715 , \42595 );
_HMUX g14ef6 ( \42717_nG14ef6 , \42714_nG14ef4 , \42716_nG14ef5 , \42599 );
buf \U$36710 ( \42718 , \42717_nG14ef6 );
_DC g1ab6a_GF_IsGateDCbyConstraint ( \42719_nG1ab6a , \42718 , \42503 );
buf \U$36711 ( \42720 , \42719_nG1ab6a );
buf \U$36712 ( \42721 , RIb8857c0_55);
_HMUX g14ef7 ( \42722_nG14ef7 , RIdab2fa0_3727 , \42721 , \42581 );
_HMUX g14ef8 ( \42723_nG14ef8 , RIdab2fa0_3727 , \42722_nG14ef7 , \42590 );
buf \U$36713 ( \42724 , RIb826ea0_223);
_HMUX g14ef9 ( \42725_nG14ef9 , RIdab2fa0_3727 , \42724 , \42595 );
_HMUX g14efa ( \42726_nG14efa , \42723_nG14ef8 , \42725_nG14ef9 , \42599 );
buf \U$36714 ( \42727 , \42726_nG14efa );
_DC g1ab6c_GF_IsGateDCbyConstraint ( \42728_nG1ab6c , \42727 , \42503 );
buf \U$36715 ( \42729 , \42728_nG1ab6c );
buf \U$36716 ( \42730 , RIb885838_54);
_HMUX g14efb ( \42731_nG14efb , RIdab8e50_3728 , \42730 , \42581 );
_HMUX g14efc ( \42732_nG14efc , RIdab8e50_3728 , \42731_nG14efb , \42590 );
buf \U$36717 ( \42733 , RIb826f18_222);
_HMUX g14efd ( \42734_nG14efd , RIdab8e50_3728 , \42733 , \42595 );
_HMUX g14efe ( \42735_nG14efe , \42732_nG14efc , \42734_nG14efd , \42599 );
buf \U$36718 ( \42736 , \42735_nG14efe );
_DC g1ab6e_GF_IsGateDCbyConstraint ( \42737_nG1ab6e , \42736 , \42503 );
buf \U$36719 ( \42738 , \42737_nG1ab6e );
buf \U$36720 ( \42739 , RIb8858b0_53);
_HMUX g14eff ( \42740_nG14eff , RIdabcf00_3729 , \42739 , \42581 );
_HMUX g14f00 ( \42741_nG14f00 , RIdabcf00_3729 , \42740_nG14eff , \42590 );
buf \U$36721 ( \42742 , RIb826f90_221);
_HMUX g14f01 ( \42743_nG14f01 , RIdabcf00_3729 , \42742 , \42595 );
_HMUX g14f02 ( \42744_nG14f02 , \42741_nG14f00 , \42743_nG14f01 , \42599 );
buf \U$36722 ( \42745 , \42744_nG14f02 );
_DC g1ab70_GF_IsGateDCbyConstraint ( \42746_nG1ab70 , \42745 , \42503 );
buf \U$36723 ( \42747 , \42746_nG1ab70 );
buf \U$36724 ( \42748 , RIb885928_52);
_HMUX g14f03 ( \42749_nG14f03 , RIdac3788_3730 , \42748 , \42581 );
_HMUX g14f04 ( \42750_nG14f04 , RIdac3788_3730 , \42749_nG14f03 , \42590 );
buf \U$36725 ( \42751 , RIb8293a8_220);
_HMUX g14f05 ( \42752_nG14f05 , RIdac3788_3730 , \42751 , \42595 );
_HMUX g14f06 ( \42753_nG14f06 , \42750_nG14f04 , \42752_nG14f05 , \42599 );
buf \U$36726 ( \42754 , \42753_nG14f06 );
_DC g1ab72_GF_IsGateDCbyConstraint ( \42755_nG1ab72 , \42754 , \42503 );
buf \U$36727 ( \42756 , \42755_nG1ab72 );
buf \U$36728 ( \42757 , RIb8859a0_51);
_HMUX g14f07 ( \42758_nG14f07 , RIdac8eb8_3731 , \42757 , \42581 );
_HMUX g14f08 ( \42759_nG14f08 , RIdac8eb8_3731 , \42758_nG14f07 , \42590 );
buf \U$36729 ( \42760 , RIb829420_219);
_HMUX g14f09 ( \42761_nG14f09 , RIdac8eb8_3731 , \42760 , \42595 );
_HMUX g14f0a ( \42762_nG14f0a , \42759_nG14f08 , \42761_nG14f09 , \42599 );
buf \U$36730 ( \42763 , \42762_nG14f0a );
_DC g1ab74_GF_IsGateDCbyConstraint ( \42764_nG1ab74 , \42763 , \42503 );
buf \U$36731 ( \42765 , \42764_nG1ab74 );
buf \U$36732 ( \42766 , RIb885a18_50);
_HMUX g14f0b ( \42767_nG14f0b , RIdacf650_3732 , \42766 , \42581 );
_HMUX g14f0c ( \42768_nG14f0c , RIdacf650_3732 , \42767_nG14f0b , \42590 );
buf \U$36733 ( \42769 , RIb829498_218);
_HMUX g14f0d ( \42770_nG14f0d , RIdacf650_3732 , \42769 , \42595 );
_HMUX g14f0e ( \42771_nG14f0e , \42768_nG14f0c , \42770_nG14f0d , \42599 );
buf \U$36734 ( \42772 , \42771_nG14f0e );
_DC g1ab78_GF_IsGateDCbyConstraint ( \42773_nG1ab78 , \42772 , \42503 );
buf \U$36735 ( \42774 , \42773_nG1ab78 );
buf \U$36736 ( \42775 , RIb885a90_49);
_HMUX g14f0f ( \42776_nG14f0f , RIdad4fd8_3733 , \42775 , \42581 );
_HMUX g14f10 ( \42777_nG14f10 , RIdad4fd8_3733 , \42776_nG14f0f , \42590 );
buf \U$36737 ( \42778 , RIb829510_217);
_HMUX g14f11 ( \42779_nG14f11 , RIdad4fd8_3733 , \42778 , \42595 );
_HMUX g14f12 ( \42780_nG14f12 , \42777_nG14f10 , \42779_nG14f11 , \42599 );
buf \U$36738 ( \42781 , \42780_nG14f12 );
_DC g1ab7a_GF_IsGateDCbyConstraint ( \42782_nG1ab7a , \42781 , \42503 );
buf \U$36739 ( \42783 , \42782_nG1ab7a );
buf \U$36740 ( \42784 , RIb885b08_48);
_HMUX g14f13 ( \42785_nG14f13 , RIdadaf00_3734 , \42784 , \42581 );
_HMUX g14f14 ( \42786_nG14f14 , RIdadaf00_3734 , \42785_nG14f13 , \42590 );
buf \U$36741 ( \42787 , RIb829588_216);
_HMUX g14f15 ( \42788_nG14f15 , RIdadaf00_3734 , \42787 , \42595 );
_HMUX g14f16 ( \42789_nG14f16 , \42786_nG14f14 , \42788_nG14f15 , \42599 );
buf \U$36742 ( \42790 , \42789_nG14f16 );
_DC g1ab7c_GF_IsGateDCbyConstraint ( \42791_nG1ab7c , \42790 , \42503 );
buf \U$36743 ( \42792 , \42791_nG1ab7c );
buf \U$36744 ( \42793 , RIb885b80_47);
_HMUX g14f17 ( \42794_nG14f17 , RIdae2610_3735 , \42793 , \42581 );
_HMUX g14f18 ( \42795_nG14f18 , RIdae2610_3735 , \42794_nG14f17 , \42590 );
buf \U$36745 ( \42796 , RIb829600_215);
_HMUX g14f19 ( \42797_nG14f19 , RIdae2610_3735 , \42796 , \42595 );
_HMUX g14f1a ( \42798_nG14f1a , \42795_nG14f18 , \42797_nG14f19 , \42599 );
buf \U$36746 ( \42799 , \42798_nG14f1a );
_DC g1ab7e_GF_IsGateDCbyConstraint ( \42800_nG1ab7e , \42799 , \42503 );
buf \U$36747 ( \42801 , \42800_nG1ab7e );
buf \U$36748 ( \42802 , RIb885bf8_46);
_HMUX g14f1b ( \42803_nG14f1b , RIdae8268_3736 , \42802 , \42581 );
_HMUX g14f1c ( \42804_nG14f1c , RIdae8268_3736 , \42803_nG14f1b , \42590 );
buf \U$36749 ( \42805 , RIb829678_214);
_HMUX g14f1d ( \42806_nG14f1d , RIdae8268_3736 , \42805 , \42595 );
_HMUX g14f1e ( \42807_nG14f1e , \42804_nG14f1c , \42806_nG14f1d , \42599 );
buf \U$36750 ( \42808 , \42807_nG14f1e );
_DC g1ab80_GF_IsGateDCbyConstraint ( \42809_nG1ab80 , \42808 , \42503 );
buf \U$36751 ( \42810 , \42809_nG1ab80 );
buf \U$36752 ( \42811 , RIb885c70_45);
_HMUX g14f1f ( \42812_nG14f1f , RIdaef720_3737 , \42811 , \42581 );
_HMUX g14f20 ( \42813_nG14f20 , RIdaef720_3737 , \42812_nG14f1f , \42590 );
buf \U$36753 ( \42814 , RIb8296f0_213);
_HMUX g14f21 ( \42815_nG14f21 , RIdaef720_3737 , \42814 , \42595 );
_HMUX g14f22 ( \42816_nG14f22 , \42813_nG14f20 , \42815_nG14f21 , \42599 );
buf \U$36754 ( \42817 , \42816_nG14f22 );
_DC g1ab82_GF_IsGateDCbyConstraint ( \42818_nG1ab82 , \42817 , \42503 );
buf \U$36755 ( \42819 , \42818_nG1ab82 );
buf \U$36756 ( \42820 , RIb885ce8_44);
_HMUX g14f23 ( \42821_nG14f23 , RIdaf4e50_3738 , \42820 , \42581 );
_HMUX g14f24 ( \42822_nG14f24 , RIdaf4e50_3738 , \42821_nG14f23 , \42590 );
buf \U$36757 ( \42823 , RIb82dae8_212);
_HMUX g14f25 ( \42824_nG14f25 , RIdaf4e50_3738 , \42823 , \42595 );
_HMUX g14f26 ( \42825_nG14f26 , \42822_nG14f24 , \42824_nG14f25 , \42599 );
buf \U$36758 ( \42826 , \42825_nG14f26 );
_DC g1ab84_GF_IsGateDCbyConstraint ( \42827_nG1ab84 , \42826 , \42503 );
buf \U$36759 ( \42828 , \42827_nG1ab84 );
buf \U$36760 ( \42829 , RIb885d60_43);
_HMUX g14f27 ( \42830_nG14f27 , RIdafa508_3739 , \42829 , \42581 );
_HMUX g14f28 ( \42831_nG14f28 , RIdafa508_3739 , \42830_nG14f27 , \42590 );
buf \U$36761 ( \42832 , RIb82db60_211);
_HMUX g14f29 ( \42833_nG14f29 , RIdafa508_3739 , \42832 , \42595 );
_HMUX g14f2a ( \42834_nG14f2a , \42831_nG14f28 , \42833_nG14f29 , \42599 );
buf \U$36762 ( \42835 , \42834_nG14f2a );
_DC g1ab86_GF_IsGateDCbyConstraint ( \42836_nG1ab86 , \42835 , \42503 );
buf \U$36763 ( \42837 , \42836_nG1ab86 );
buf \U$36764 ( \42838 , RIb885dd8_42);
_HMUX g14f2b ( \42839_nG14f2b , RIdafe630_3740 , \42838 , \42581 );
_HMUX g14f2c ( \42840_nG14f2c , RIdafe630_3740 , \42839_nG14f2b , \42590 );
buf \U$36765 ( \42841 , RIb82dbd8_210);
_HMUX g14f2d ( \42842_nG14f2d , RIdafe630_3740 , \42841 , \42595 );
_HMUX g14f2e ( \42843_nG14f2e , \42840_nG14f2c , \42842_nG14f2d , \42599 );
buf \U$36766 ( \42844 , \42843_nG14f2e );
_DC g1ab88_GF_IsGateDCbyConstraint ( \42845_nG1ab88 , \42844 , \42503 );
buf \U$36767 ( \42846 , \42845_nG1ab88 );
buf \U$36768 ( \42847 , RIb885e50_41);
_HMUX g14f2f ( \42848_nG14f2f , RIdb03b08_3741 , \42847 , \42581 );
_HMUX g14f30 ( \42849_nG14f30 , RIdb03b08_3741 , \42848_nG14f2f , \42590 );
buf \U$36769 ( \42850 , RIb82dc50_209);
_HMUX g14f31 ( \42851_nG14f31 , RIdb03b08_3741 , \42850 , \42595 );
_HMUX g14f32 ( \42852_nG14f32 , \42849_nG14f30 , \42851_nG14f31 , \42599 );
buf \U$36770 ( \42853 , \42852_nG14f32 );
_DC g1ab8a_GF_IsGateDCbyConstraint ( \42854_nG1ab8a , \42853 , \42503 );
buf \U$36771 ( \42855 , \42854_nG1ab8a );
buf \U$36772 ( \42856 , RIb885ec8_40);
_HMUX g14f33 ( \42857_nG14f33 , RIdb09d00_3742 , \42856 , \42581 );
_HMUX g14f34 ( \42858_nG14f34 , RIdb09d00_3742 , \42857_nG14f33 , \42590 );
buf \U$36773 ( \42859 , RIb82dcc8_208);
_HMUX g14f35 ( \42860_nG14f35 , RIdb09d00_3742 , \42859 , \42595 );
_HMUX g14f36 ( \42861_nG14f36 , \42858_nG14f34 , \42860_nG14f35 , \42599 );
buf \U$36774 ( \42862 , \42861_nG14f36 );
_DC g1ab8e_GF_IsGateDCbyConstraint ( \42863_nG1ab8e , \42862 , \42503 );
buf \U$36775 ( \42864 , \42863_nG1ab8e );
buf \U$36776 ( \42865 , RIb885f40_39);
_HMUX g14f37 ( \42866_nG14f37 , RIdb0e440_3743 , \42865 , \42581 );
_HMUX g14f38 ( \42867_nG14f38 , RIdb0e440_3743 , \42866_nG14f37 , \42590 );
buf \U$36777 ( \42868 , RIb82dd40_207);
_HMUX g14f39 ( \42869_nG14f39 , RIdb0e440_3743 , \42868 , \42595 );
_HMUX g14f3a ( \42870_nG14f3a , \42867_nG14f38 , \42869_nG14f39 , \42599 );
buf \U$36778 ( \42871 , \42870_nG14f3a );
_DC g1ab90_GF_IsGateDCbyConstraint ( \42872_nG1ab90 , \42871 , \42503 );
buf \U$36779 ( \42873 , \42872_nG1ab90 );
buf \U$36780 ( \42874 , RIb885fb8_38);
_HMUX g14f3b ( \42875_nG14f3b , RIdb13468_3744 , \42874 , \42581 );
_HMUX g14f3c ( \42876_nG14f3c , RIdb13468_3744 , \42875_nG14f3b , \42590 );
buf \U$36781 ( \42877 , RIb82ddb8_206);
_HMUX g14f3d ( \42878_nG14f3d , RIdb13468_3744 , \42877 , \42595 );
_HMUX g14f3e ( \42879_nG14f3e , \42876_nG14f3c , \42878_nG14f3d , \42599 );
buf \U$36782 ( \42880 , \42879_nG14f3e );
_DC g1ab92_GF_IsGateDCbyConstraint ( \42881_nG1ab92 , \42880 , \42503 );
buf \U$36783 ( \42882 , \42881_nG1ab92 );
buf \U$36784 ( \42883 , RIb886030_37);
_HMUX g14f3f ( \42884_nG14f3f , RId9d7370_3745 , \42883 , \42581 );
_HMUX g14f40 ( \42885_nG14f40 , RId9d7370_3745 , \42884_nG14f3f , \42590 );
buf \U$36785 ( \42886 , RIb82de30_205);
_HMUX g14f41 ( \42887_nG14f41 , RId9d7370_3745 , \42886 , \42595 );
_HMUX g14f42 ( \42888_nG14f42 , \42885_nG14f40 , \42887_nG14f41 , \42599 );
buf \U$36786 ( \42889 , \42888_nG14f42 );
_DC g1ab94_GF_IsGateDCbyConstraint ( \42890_nG1ab94 , \42889 , \42503 );
buf \U$36787 ( \42891 , \42890_nG1ab94 );
buf \U$36788 ( \42892 , RIb8860a8_36);
_HMUX g14f43 ( \42893_nG14f43 , RId9d25a0_3746 , \42892 , \42581 );
_HMUX g14f44 ( \42894_nG14f44 , RId9d25a0_3746 , \42893_nG14f43 , \42590 );
buf \U$36789 ( \42895 , RIb832228_204);
_HMUX g14f45 ( \42896_nG14f45 , RId9d25a0_3746 , \42895 , \42595 );
_HMUX g14f46 ( \42897_nG14f46 , \42894_nG14f44 , \42896_nG14f45 , \42599 );
buf \U$36790 ( \42898 , \42897_nG14f46 );
_DC g1ab96_GF_IsGateDCbyConstraint ( \42899_nG1ab96 , \42898 , \42503 );
buf \U$36791 ( \42900 , \42899_nG1ab96 );
buf \U$36792 ( \42901 , RIb886120_35);
_HMUX g14f47 ( \42902_nG14f47 , RId9cd0c8_3747 , \42901 , \42581 );
_HMUX g14f48 ( \42903_nG14f48 , RId9cd0c8_3747 , \42902_nG14f47 , \42590 );
buf \U$36793 ( \42904 , RIb8322a0_203);
_HMUX g14f49 ( \42905_nG14f49 , RId9cd0c8_3747 , \42904 , \42595 );
_HMUX g14f4a ( \42906_nG14f4a , \42903_nG14f48 , \42905_nG14f49 , \42599 );
buf \U$36794 ( \42907 , \42906_nG14f4a );
_DC g1ab98_GF_IsGateDCbyConstraint ( \42908_nG1ab98 , \42907 , \42503 );
buf \U$36795 ( \42909 , \42908_nG1ab98 );
buf \U$36796 ( \42910 , RIb886198_34);
_HMUX g14f4b ( \42911_nG14f4b , RId9c86b8_3748 , \42910 , \42581 );
_HMUX g14f4c ( \42912_nG14f4c , RId9c86b8_3748 , \42911_nG14f4b , \42590 );
buf \U$36797 ( \42913 , RIb832318_202);
_HMUX g14f4d ( \42914_nG14f4d , RId9c86b8_3748 , \42913 , \42595 );
_HMUX g14f4e ( \42915_nG14f4e , \42912_nG14f4c , \42914_nG14f4d , \42599 );
buf \U$36798 ( \42916 , \42915_nG14f4e );
_DC g1ab9a_GF_IsGateDCbyConstraint ( \42917_nG1ab9a , \42916 , \42503 );
buf \U$36799 ( \42918 , \42917_nG1ab9a );
buf \U$36800 ( \42919 , RIb886210_33);
_HMUX g14f4f ( \42920_nG14f4f , RIda940a0_3749 , \42919 , \42581 );
_HMUX g14f50 ( \42921_nG14f50 , RIda940a0_3749 , \42920_nG14f4f , \42590 );
buf \U$36801 ( \42922 , RIb832390_201);
_HMUX g14f51 ( \42923_nG14f51 , RIda940a0_3749 , \42922 , \42595 );
_HMUX g14f52 ( \42924_nG14f52 , \42921_nG14f50 , \42923_nG14f51 , \42599 );
buf \U$36802 ( \42925 , \42924_nG14f52 );
_DC g1ab9c_GF_IsGateDCbyConstraint ( \42926_nG1ab9c , \42925 , \42503 );
buf \U$36803 ( \42927 , \42926_nG1ab9c );
buf \U$36804 ( \42928 , RIb886288_32);
_HMUX g14f53 ( \42929_nG14f53 , RIda91850_3750 , \42928 , \42581 );
_HMUX g14f54 ( \42930_nG14f54 , RIda91850_3750 , \42929_nG14f53 , \42590 );
buf \U$36805 ( \42931 , RIb832408_200);
_HMUX g14f55 ( \42932_nG14f55 , RIda91850_3750 , \42931 , \42595 );
_HMUX g14f56 ( \42933_nG14f56 , \42930_nG14f54 , \42932_nG14f55 , \42599 );
buf \U$36806 ( \42934 , \42933_nG14f56 );
_DC g1ab9e_GF_IsGateDCbyConstraint ( \42935_nG1ab9e , \42934 , \42503 );
buf \U$36807 ( \42936 , \42935_nG1ab9e );
buf \U$36808 ( \42937 , RIb886300_31);
_HMUX g14f57 ( \42938_nG14f57 , RIda8dbd8_3751 , \42937 , \42581 );
_HMUX g14f58 ( \42939_nG14f58 , RIda8dbd8_3751 , \42938_nG14f57 , \42590 );
buf \U$36809 ( \42940 , RIb832480_199);
_HMUX g14f59 ( \42941_nG14f59 , RIda8dbd8_3751 , \42940 , \42595 );
_HMUX g14f5a ( \42942_nG14f5a , \42939_nG14f58 , \42941_nG14f59 , \42599 );
buf \U$36810 ( \42943 , \42942_nG14f5a );
_DC g1aba0_GF_IsGateDCbyConstraint ( \42944_nG1aba0 , \42943 , \42503 );
buf \U$36811 ( \42945 , \42944_nG1aba0 );
buf \U$36812 ( \42946 , RIb886378_30);
_HMUX g14f5b ( \42947_nG14f5b , RIda8a7d0_3752 , \42946 , \42581 );
_HMUX g14f5c ( \42948_nG14f5c , RIda8a7d0_3752 , \42947_nG14f5b , \42590 );
buf \U$36813 ( \42949 , RIb8324f8_198);
_HMUX g14f5d ( \42950_nG14f5d , RIda8a7d0_3752 , \42949 , \42595 );
_HMUX g14f5e ( \42951_nG14f5e , \42948_nG14f5c , \42950_nG14f5d , \42599 );
buf \U$36814 ( \42952 , \42951_nG14f5e );
_DC g1aba4_GF_IsGateDCbyConstraint ( \42953_nG1aba4 , \42952 , \42503 );
buf \U$36815 ( \42954 , \42953_nG1aba4 );
buf \U$36816 ( \42955 , RIb8863f0_29);
_HMUX g14f5f ( \42956_nG14f5f , RIda86978_3753 , \42955 , \42581 );
_HMUX g14f60 ( \42957_nG14f60 , RIda86978_3753 , \42956_nG14f5f , \42590 );
buf \U$36817 ( \42958 , RIb832570_197);
_HMUX g14f61 ( \42959_nG14f61 , RIda86978_3753 , \42958 , \42595 );
_HMUX g14f62 ( \42960_nG14f62 , \42957_nG14f60 , \42959_nG14f61 , \42599 );
buf \U$36818 ( \42961 , \42960_nG14f62 );
_DC g1aba6_GF_IsGateDCbyConstraint ( \42962_nG1aba6 , \42961 , \42503 );
buf \U$36819 ( \42963 , \42962_nG1aba6 );
buf \U$36820 ( \42964 , RIb886468_28);
_HMUX g14f63 ( \42965_nG14f63 , RIda835e8_3754 , \42964 , \42581 );
_HMUX g14f64 ( \42966_nG14f64 , RIda835e8_3754 , \42965_nG14f63 , \42590 );
buf \U$36821 ( \42967 , RIb8383a8_196);
_HMUX g14f65 ( \42968_nG14f65 , RIda835e8_3754 , \42967 , \42595 );
_HMUX g14f66 ( \42969_nG14f66 , \42966_nG14f64 , \42968_nG14f65 , \42599 );
buf \U$36822 ( \42970 , \42969_nG14f66 );
_DC g1aba8_GF_IsGateDCbyConstraint ( \42971_nG1aba8 , \42970 , \42503 );
buf \U$36823 ( \42972 , \42971_nG1aba8 );
buf \U$36824 ( \42973 , RIb8864e0_27);
_HMUX g14f67 ( \42974_nG14f67 , RIda80f00_3755 , \42973 , \42581 );
_HMUX g14f68 ( \42975_nG14f68 , RIda80f00_3755 , \42974_nG14f67 , \42590 );
buf \U$36825 ( \42976 , RIb838420_195);
_HMUX g14f69 ( \42977_nG14f69 , RIda80f00_3755 , \42976 , \42595 );
_HMUX g14f6a ( \42978_nG14f6a , \42975_nG14f68 , \42977_nG14f69 , \42599 );
buf \U$36826 ( \42979 , \42978_nG14f6a );
_DC g1abaa_GF_IsGateDCbyConstraint ( \42980_nG1abaa , \42979 , \42503 );
buf \U$36827 ( \42981 , \42980_nG1abaa );
buf \U$36828 ( \42982 , RIb886558_26);
_HMUX g14f6b ( \42983_nG14f6b , RIda7daf8_3756 , \42982 , \42581 );
_HMUX g14f6c ( \42984_nG14f6c , RIda7daf8_3756 , \42983_nG14f6b , \42590 );
buf \U$36829 ( \42985 , RIb838498_194);
_HMUX g14f6d ( \42986_nG14f6d , RIda7daf8_3756 , \42985 , \42595 );
_HMUX g14f6e ( \42987_nG14f6e , \42984_nG14f6c , \42986_nG14f6d , \42599 );
buf \U$36830 ( \42988 , \42987_nG14f6e );
_DC g1abac_GF_IsGateDCbyConstraint ( \42989_nG1abac , \42988 , \42503 );
buf \U$36831 ( \42990 , \42989_nG1abac );
buf \U$36832 ( \42991 , RIb8865d0_25);
_HMUX g14f6f ( \42992_nG14f6f , RIda7a7e0_3757 , \42991 , \42581 );
_HMUX g14f70 ( \42993_nG14f70 , RIda7a7e0_3757 , \42992_nG14f6f , \42590 );
buf \U$36833 ( \42994 , RIb838510_193);
_HMUX g14f71 ( \42995_nG14f71 , RIda7a7e0_3757 , \42994 , \42595 );
_HMUX g14f72 ( \42996_nG14f72 , \42993_nG14f70 , \42995_nG14f71 , \42599 );
buf \U$36834 ( \42997 , \42996_nG14f72 );
_DC g1abae_GF_IsGateDCbyConstraint ( \42998_nG1abae , \42997 , \42503 );
buf \U$36835 ( \42999 , \42998_nG1abae );
buf \U$36836 ( \43000 , RIb886648_24);
_HMUX g14f73 ( \43001_nG14f73 , RIda745e8_3758 , \43000 , \42581 );
_HMUX g14f74 ( \43002_nG14f74 , RIda745e8_3758 , \43001_nG14f73 , \42590 );
buf \U$36837 ( \43003 , RIb838588_192);
_HMUX g14f75 ( \43004_nG14f75 , RIda745e8_3758 , \43003 , \42595 );
_HMUX g14f76 ( \43005_nG14f76 , \43002_nG14f74 , \43004_nG14f75 , \42599 );
buf \U$36838 ( \43006 , \43005_nG14f76 );
_DC g1abb0_GF_IsGateDCbyConstraint ( \43007_nG1abb0 , \43006 , \42503 );
buf \U$36839 ( \43008 , \43007_nG1abb0 );
buf \U$36840 ( \43009 , RIb8866c0_23);
_HMUX g14f77 ( \43010_nG14f77 , RIda6e018_3759 , \43009 , \42581 );
_HMUX g14f78 ( \43011_nG14f78 , RIda6e018_3759 , \43010_nG14f77 , \42590 );
buf \U$36841 ( \43012 , RIb838600_191);
_HMUX g14f79 ( \43013_nG14f79 , RIda6e018_3759 , \43012 , \42595 );
_HMUX g14f7a ( \43014_nG14f7a , \43011_nG14f78 , \43013_nG14f79 , \42599 );
buf \U$36842 ( \43015 , \43014_nG14f7a );
_DC g1abb2_GF_IsGateDCbyConstraint ( \43016_nG1abb2 , \43015 , \42503 );
buf \U$36843 ( \43017 , \43016_nG1abb2 );
buf \U$36844 ( \43018 , RIb886738_22);
_HMUX g14f7b ( \43019_nG14f7b , RIda65e40_3760 , \43018 , \42581 );
_HMUX g14f7c ( \43020_nG14f7c , RIda65e40_3760 , \43019_nG14f7b , \42590 );
buf \U$36845 ( \43021 , RIb838678_190);
_HMUX g14f7d ( \43022_nG14f7d , RIda65e40_3760 , \43021 , \42595 );
_HMUX g14f7e ( \43023_nG14f7e , \43020_nG14f7c , \43022_nG14f7d , \42599 );
buf \U$36846 ( \43024 , \43023_nG14f7e );
_DC g1abb4_GF_IsGateDCbyConstraint ( \43025_nG1abb4 , \43024 , \42503 );
buf \U$36847 ( \43026 , \43025_nG1abb4 );
buf \U$36848 ( \43027 , RIb8867b0_21);
_HMUX g14f7f ( \43028_nG14f7f , RIda5f888_3761 , \43027 , \42581 );
_HMUX g14f80 ( \43029_nG14f80 , RIda5f888_3761 , \43028_nG14f7f , \42590 );
buf \U$36849 ( \43030 , RIb8386f0_189);
_HMUX g14f81 ( \43031_nG14f81 , RIda5f888_3761 , \43030 , \42595 );
_HMUX g14f82 ( \43032_nG14f82 , \43029_nG14f80 , \43031_nG14f81 , \42599 );
buf \U$36850 ( \43033 , \43032_nG14f82 );
_DC g1abb6_GF_IsGateDCbyConstraint ( \43034_nG1abb6 , \43033 , \42503 );
buf \U$36851 ( \43035 , \43034_nG1abb6 );
buf \U$36852 ( \43036 , RIb886828_20);
_HMUX g14f83 ( \43037_nG14f83 , RIda59780_3762 , \43036 , \42581 );
_HMUX g14f84 ( \43038_nG14f84 , RIda59780_3762 , \43037_nG14f83 , \42590 );
buf \U$36853 ( \43039 , RIb838768_188);
_HMUX g14f85 ( \43040_nG14f85 , RIda59780_3762 , \43039 , \42595 );
_HMUX g14f86 ( \43041_nG14f86 , \43038_nG14f84 , \43040_nG14f85 , \42599 );
buf \U$36854 ( \43042 , \43041_nG14f86 );
_DC g1abba_GF_IsGateDCbyConstraint ( \43043_nG1abba , \43042 , \42503 );
buf \U$36855 ( \43044 , \43043_nG1abba );
buf \U$36856 ( \43045 , RIb8868a0_19);
_HMUX g14f87 ( \43046_nG14f87 , RIda510f8_3763 , \43045 , \42581 );
_HMUX g14f88 ( \43047_nG14f88 , RIda510f8_3763 , \43046_nG14f87 , \42590 );
buf \U$36857 ( \43048 , RIb8387e0_187);
_HMUX g14f89 ( \43049_nG14f89 , RIda510f8_3763 , \43048 , \42595 );
_HMUX g14f8a ( \43050_nG14f8a , \43047_nG14f88 , \43049_nG14f89 , \42599 );
buf \U$36858 ( \43051 , \43050_nG14f8a );
_DC g1abbc_GF_IsGateDCbyConstraint ( \43052_nG1abbc , \43051 , \42503 );
buf \U$36859 ( \43053 , \43052_nG1abbc );
buf \U$36860 ( \43054 , RIb886918_18);
_HMUX g14f8b ( \43055_nG14f8b , RIda4aff0_3764 , \43054 , \42581 );
_HMUX g14f8c ( \43056_nG14f8c , RIda4aff0_3764 , \43055_nG14f8b , \42590 );
buf \U$36861 ( \43057 , RIb838858_186);
_HMUX g14f8d ( \43058_nG14f8d , RIda4aff0_3764 , \43057 , \42595 );
_HMUX g14f8e ( \43059_nG14f8e , \43056_nG14f8c , \43058_nG14f8d , \42599 );
buf \U$36862 ( \43060 , \43059_nG14f8e );
_DC g1abbe_GF_IsGateDCbyConstraint ( \43061_nG1abbe , \43060 , \42503 );
buf \U$36863 ( \43062 , \43061_nG1abbe );
buf \U$36864 ( \43063 , RIb886990_17);
_HMUX g14f8f ( \43064_nG14f8f , RId927408_3765 , \43063 , \42581 );
_HMUX g14f90 ( \43065_nG14f90 , RId927408_3765 , \43064_nG14f8f , \42590 );
buf \U$36865 ( \43066 , RIb8388d0_185);
_HMUX g14f91 ( \43067_nG14f91 , RId927408_3765 , \43066 , \42595 );
_HMUX g14f92 ( \43068_nG14f92 , \43065_nG14f90 , \43067_nG14f91 , \42599 );
buf \U$36866 ( \43069 , \43068_nG14f92 );
_DC g1abc0_GF_IsGateDCbyConstraint ( \43070_nG1abc0 , \43069 , \42503 );
buf \U$36867 ( \43071 , \43070_nG1abc0 );
buf \U$36868 ( \43072 , RIb886a08_16);
_HMUX g14f93 ( \43073_nG14f93 , RId943680_3766 , \43072 , \42581 );
_HMUX g14f94 ( \43074_nG14f94 , RId943680_3766 , \43073_nG14f93 , \42590 );
buf \U$36869 ( \43075 , RIb838948_184);
_HMUX g14f95 ( \43076_nG14f95 , RId943680_3766 , \43075 , \42595 );
_HMUX g14f96 ( \43077_nG14f96 , \43074_nG14f94 , \43076_nG14f95 , \42599 );
buf \U$36870 ( \43078 , \43077_nG14f96 );
_DC g1abc2_GF_IsGateDCbyConstraint ( \43079_nG1abc2 , \43078 , \42503 );
buf \U$36871 ( \43080 , \43079_nG1abc2 );
buf \U$36872 ( \43081 , RIb886a80_15);
_HMUX g14f97 ( \43082_nG14f97 , RId96ccd8_3767 , \43081 , \42581 );
_HMUX g14f98 ( \43083_nG14f98 , RId96ccd8_3767 , \43082_nG14f97 , \42590 );
buf \U$36873 ( \43084 , RIb8389c0_183);
_HMUX g14f99 ( \43085_nG14f99 , RId96ccd8_3767 , \43084 , \42595 );
_HMUX g14f9a ( \43086_nG14f9a , \43083_nG14f98 , \43085_nG14f99 , \42599 );
buf \U$36874 ( \43087 , \43086_nG14f9a );
_DC g1abc4_GF_IsGateDCbyConstraint ( \43088_nG1abc4 , \43087 , \42503 );
buf \U$36875 ( \43089 , \43088_nG1abc4 );
buf \U$36876 ( \43090 , RIb886af8_14);
_HMUX g14f9b ( \43091_nG14f9b , RId988b30_3768 , \43090 , \42581 );
_HMUX g14f9c ( \43092_nG14f9c , RId988b30_3768 , \43091_nG14f9b , \42590 );
buf \U$36877 ( \43093 , RIb838a38_182);
_HMUX g14f9d ( \43094_nG14f9d , RId988b30_3768 , \43093 , \42595 );
_HMUX g14f9e ( \43095_nG14f9e , \43092_nG14f9c , \43094_nG14f9d , \42599 );
buf \U$36878 ( \43096 , \43095_nG14f9e );
_DC g1abc6_GF_IsGateDCbyConstraint ( \43097_nG1abc6 , \43096 , \42503 );
buf \U$36879 ( \43098 , \43097_nG1abc6 );
buf \U$36880 ( \43099 , RIb886b70_13);
_HMUX g14f9f ( \43100_nG14f9f , RId90bb68_3769 , \43099 , \42581 );
_HMUX g14fa0 ( \43101_nG14fa0 , RId90bb68_3769 , \43100_nG14f9f , \42590 );
buf \U$36881 ( \43102 , RIb838ab0_181);
_HMUX g14fa1 ( \43103_nG14fa1 , RId90bb68_3769 , \43102 , \42595 );
_HMUX g14fa2 ( \43104_nG14fa2 , \43101_nG14fa0 , \43103_nG14fa1 , \42599 );
buf \U$36882 ( \43105 , \43104_nG14fa2 );
_DC g1abc8_GF_IsGateDCbyConstraint ( \43106_nG1abc8 , \43105 , \42503 );
buf \U$36883 ( \43107 , \43106_nG1abc8 );
buf \U$36884 ( \43108 , RIb886be8_12);
_HMUX g14fa3 ( \43109_nG14fa3 , RId8f7438_3770 , \43108 , \42581 );
_HMUX g14fa4 ( \43110_nG14fa4 , RId8f7438_3770 , \43109_nG14fa3 , \42590 );
buf \U$36885 ( \43111 , RIb838b28_180);
_HMUX g14fa5 ( \43112_nG14fa5 , RId8f7438_3770 , \43111 , \42595 );
_HMUX g14fa6 ( \43113_nG14fa6 , \43110_nG14fa4 , \43112_nG14fa5 , \42599 );
buf \U$36886 ( \43114 , \43113_nG14fa6 );
_DC g1abca_GF_IsGateDCbyConstraint ( \43115_nG1abca , \43114 , \42503 );
buf \U$36887 ( \43116 , \43115_nG1abca );
buf \U$36888 ( \43117 , RIb886c60_11);
_HMUX g14fa7 ( \43118_nG14fa7 , RId8d6dc8_3771 , \43117 , \42581 );
_HMUX g14fa8 ( \43119_nG14fa8 , RId8d6dc8_3771 , \43118_nG14fa7 , \42590 );
buf \U$36889 ( \43120 , RIb838ba0_179);
_HMUX g14fa9 ( \43121_nG14fa9 , RId8d6dc8_3771 , \43120 , \42595 );
_HMUX g14faa ( \43122_nG14faa , \43119_nG14fa8 , \43121_nG14fa9 , \42599 );
buf \U$36890 ( \43123 , \43122_nG14faa );
_DC g1abcc_GF_IsGateDCbyConstraint ( \43124_nG1abcc , \43123 , \42503 );
buf \U$36891 ( \43125 , \43124_nG1abcc );
buf \U$36892 ( \43126 , RIb886cd8_10);
_HMUX g14fab ( \43127_nG14fab , RId6c4d70_3772 , \43126 , \42581 );
_HMUX g14fac ( \43128_nG14fac , RId6c4d70_3772 , \43127_nG14fab , \42590 );
buf \U$36893 ( \43129 , RIb838c18_178);
_HMUX g14fad ( \43130_nG14fad , RId6c4d70_3772 , \43129 , \42595 );
_HMUX g14fae ( \43131_nG14fae , \43128_nG14fac , \43130_nG14fad , \42599 );
buf \U$36894 ( \43132 , \43131_nG14fae );
_DC g1abd0_GF_IsGateDCbyConstraint ( \43133_nG1abd0 , \43132 , \42503 );
buf \U$36895 ( \43134 , \43133_nG1abd0 );
buf \U$36896 ( \43135 , RIb886d50_9);
_HMUX g14faf ( \43136_nG14faf , RId6ae7c8_3773 , \43135 , \42581 );
_HMUX g14fb0 ( \43137_nG14fb0 , RId6ae7c8_3773 , \43136_nG14faf , \42590 );
buf \U$36897 ( \43138 , RIb838c90_177);
_HMUX g14fb1 ( \43139_nG14fb1 , RId6ae7c8_3773 , \43138 , \42595 );
_HMUX g14fb2 ( \43140_nG14fb2 , \43137_nG14fb0 , \43139_nG14fb1 , \42599 );
buf \U$36898 ( \43141 , \43140_nG14fb2 );
_DC g1abd2_GF_IsGateDCbyConstraint ( \43142_nG1abd2 , \43141 , \42503 );
buf \U$36899 ( \43143 , \43142_nG1abd2 );
buf \U$36900 ( \43144 , RIb886dc8_8);
_HMUX g14fb3 ( \43145_nG14fb3 , RId835578_3774 , \43144 , \42581 );
_HMUX g14fb4 ( \43146_nG14fb4 , RId835578_3774 , \43145_nG14fb3 , \42590 );
buf \U$36901 ( \43147 , RIb838d08_176);
_HMUX g14fb5 ( \43148_nG14fb5 , RId835578_3774 , \43147 , \42595 );
_HMUX g14fb6 ( \43149_nG14fb6 , \43146_nG14fb4 , \43148_nG14fb5 , \42599 );
buf \U$36902 ( \43150 , \43149_nG14fb6 );
_DC g1abd4_GF_IsGateDCbyConstraint ( \43151_nG1abd4 , \43150 , \42503 );
buf \U$36903 ( \43152 , \43151_nG1abd4 );
buf \U$36904 ( \43153 , RIb886e40_7);
_HMUX g14fb7 ( \43154_nG14fb7 , RId8a9d50_3775 , \43153 , \42581 );
_HMUX g14fb8 ( \43155_nG14fb8 , RId8a9d50_3775 , \43154_nG14fb7 , \42590 );
buf \U$36905 ( \43156 , RIb838d80_175);
_HMUX g14fb9 ( \43157_nG14fb9 , RId8a9d50_3775 , \43156 , \42595 );
_HMUX g14fba ( \43158_nG14fba , \43155_nG14fb8 , \43157_nG14fb9 , \42599 );
buf \U$36906 ( \43159 , \43158_nG14fba );
_DC g1abd6_GF_IsGateDCbyConstraint ( \43160_nG1abd6 , \43159 , \42503 );
buf \U$36907 ( \43161 , \43160_nG1abd6 );
buf \U$36908 ( \43162 , RIb886eb8_6);
_HMUX g14fbb ( \43163_nG14fbb , RId862aa0_3776 , \43162 , \42581 );
_HMUX g14fbc ( \43164_nG14fbc , RId862aa0_3776 , \43163_nG14fbb , \42590 );
buf \U$36909 ( \43165 , RIb838df8_174);
_HMUX g14fbd ( \43166_nG14fbd , RId862aa0_3776 , \43165 , \42595 );
_HMUX g14fbe ( \43167_nG14fbe , \43164_nG14fbc , \43166_nG14fbd , \42599 );
buf \U$36910 ( \43168 , \43167_nG14fbe );
_DC g1abd8_GF_IsGateDCbyConstraint ( \43169_nG1abd8 , \43168 , \42503 );
buf \U$36911 ( \43170 , \43169_nG1abd8 );
not \U$36912 ( \43171 , \42580 );
and \U$36913 ( \43172 , \42579 , \43171 );
_HMUX g14dbd ( \43173_nG14dbd , RId99e778_3777 , \42578 , \43172 );
_HMUX g14dbe ( \43174_nG14dbe , RId99e778_3777 , \43173_nG14dbd , \42590 );
not \U$36914 ( \43175 , \42594 );
and \U$36915 ( \43176 , \42593 , \43175 );
_HMUX g14dc0 ( \43177_nG14dc0 , RId99e778_3777 , \42592 , \43176 );
_HMUX g14dc1 ( \43178_nG14dc1 , \43174_nG14dbe , \43177_nG14dc0 , \42599 );
buf \U$36916 ( \43179 , \43178_nG14dc1 );
_DC g1aae0_GF_IsGateDCbyConstraint ( \43180_nG1aae0 , \43179 , \42503 );
buf \U$36917 ( \43181 , \43180_nG1aae0 );
_HMUX g14dc2 ( \43182_nG14dc2 , RId9ac620_3778 , \42604 , \43172 );
_HMUX g14dc3 ( \43183_nG14dc3 , RId9ac620_3778 , \43182_nG14dc2 , \42590 );
_HMUX g14dc4 ( \43184_nG14dc4 , RId9ac620_3778 , \42607 , \43176 );
_HMUX g14dc5 ( \43185_nG14dc5 , \43183_nG14dc3 , \43184_nG14dc4 , \42599 );
buf \U$36918 ( \43186 , \43185_nG14dc5 );
_DC g1aaf6_GF_IsGateDCbyConstraint ( \43187_nG1aaf6 , \43186 , \42503 );
buf \U$36919 ( \43188 , \43187_nG1aaf6 );
_HMUX g14dc6 ( \43189_nG14dc6 , RId9b8290_3779 , \42613 , \43172 );
_HMUX g14dc7 ( \43190_nG14dc7 , RId9b8290_3779 , \43189_nG14dc6 , \42590 );
_HMUX g14dc8 ( \43191_nG14dc8 , RId9b8290_3779 , \42616 , \43176 );
_HMUX g14dc9 ( \43192_nG14dc9 , \43190_nG14dc7 , \43191_nG14dc8 , \42599 );
buf \U$36920 ( \43193 , \43192_nG14dc9 );
_DC g1ab0c_GF_IsGateDCbyConstraint ( \43194_nG1ab0c , \43193 , \42503 );
buf \U$36921 ( \43195 , \43194_nG1ab0c );
_HMUX g14dca ( \43196_nG14dca , RId9bdfd8_3780 , \42622 , \43172 );
_HMUX g14dcb ( \43197_nG14dcb , RId9bdfd8_3780 , \43196_nG14dca , \42590 );
_HMUX g14dcc ( \43198_nG14dcc , RId9bdfd8_3780 , \42625 , \43176 );
_HMUX g14dcd ( \43199_nG14dcd , \43197_nG14dcb , \43198_nG14dcc , \42599 );
buf \U$36922 ( \43200 , \43199_nG14dcd );
_DC g1ab22_GF_IsGateDCbyConstraint ( \43201_nG1ab22 , \43200 , \42503 );
buf \U$36923 ( \43202 , \43201_nG1ab22 );
_HMUX g14dce ( \43203_nG14dce , RId90fe70_3781 , \42631 , \43172 );
_HMUX g14dcf ( \43204_nG14dcf , RId90fe70_3781 , \43203_nG14dce , \42590 );
_HMUX g14dd0 ( \43205_nG14dd0 , RId90fe70_3781 , \42634 , \43176 );
_HMUX g14dd1 ( \43206_nG14dd1 , \43204_nG14dcf , \43205_nG14dd0 , \42599 );
buf \U$36924 ( \43207 , \43206_nG14dd1 );
_DC g1ab38_GF_IsGateDCbyConstraint ( \43208_nG1ab38 , \43207 , \42503 );
buf \U$36925 ( \43209 , \43208_nG1ab38 );
_HMUX g14dd2 ( \43210_nG14dd2 , RId918b10_3782 , \42640 , \43172 );
_HMUX g14dd3 ( \43211_nG14dd3 , RId918b10_3782 , \43210_nG14dd2 , \42590 );
_HMUX g14dd4 ( \43212_nG14dd4 , RId918b10_3782 , \42643 , \43176 );
_HMUX g14dd5 ( \43213_nG14dd5 , \43211_nG14dd3 , \43212_nG14dd4 , \42599 );
buf \U$36926 ( \43214 , \43213_nG14dd5 );
_DC g1ab4e_GF_IsGateDCbyConstraint ( \43215_nG1ab4e , \43214 , \42503 );
buf \U$36927 ( \43216 , \43215_nG1ab4e );
_HMUX g14dd6 ( \43217_nG14dd6 , RIda42698_3783 , \42649 , \43172 );
_HMUX g14dd7 ( \43218_nG14dd7 , RIda42698_3783 , \43217_nG14dd6 , \42590 );
_HMUX g14dd8 ( \43219_nG14dd8 , RIda42698_3783 , \42652 , \43176 );
_HMUX g14dd9 ( \43220_nG14dd9 , \43218_nG14dd7 , \43219_nG14dd8 , \42599 );
buf \U$36928 ( \43221 , \43220_nG14dd9 );
_DC g1ab5a_GF_IsGateDCbyConstraint ( \43222_nG1ab5a , \43221 , \42503 );
buf \U$36929 ( \43223 , \43222_nG1ab5a );
_HMUX g14dda ( \43224_nG14dda , RIda33a58_3784 , \42658 , \43172 );
_HMUX g14ddb ( \43225_nG14ddb , RIda33a58_3784 , \43224_nG14dda , \42590 );
_HMUX g14ddc ( \43226_nG14ddc , RIda33a58_3784 , \42661 , \43176 );
_HMUX g14ddd ( \43227_nG14ddd , \43225_nG14ddb , \43226_nG14ddc , \42599 );
buf \U$36930 ( \43228 , \43227_nG14ddd );
_DC g1ab5c_GF_IsGateDCbyConstraint ( \43229_nG1ab5c , \43228 , \42503 );
buf \U$36931 ( \43230 , \43229_nG1ab5c );
_HMUX g14dde ( \43231_nG14dde , RIda28b08_3785 , \42667 , \43172 );
_HMUX g14ddf ( \43232_nG14ddf , RIda28b08_3785 , \43231_nG14dde , \42590 );
_HMUX g14de0 ( \43233_nG14de0 , RIda28b08_3785 , \42670 , \43176 );
_HMUX g14de1 ( \43234_nG14de1 , \43232_nG14ddf , \43233_nG14de0 , \42599 );
buf \U$36932 ( \43235 , \43234_nG14de1 );
_DC g1ab5e_GF_IsGateDCbyConstraint ( \43236_nG1ab5e , \43235 , \42503 );
buf \U$36933 ( \43237 , \43236_nG1ab5e );
_HMUX g14de2 ( \43238_nG14de2 , RIda18aa0_3786 , \42676 , \43172 );
_HMUX g14de3 ( \43239_nG14de3 , RIda18aa0_3786 , \43238_nG14de2 , \42590 );
_HMUX g14de4 ( \43240_nG14de4 , RIda18aa0_3786 , \42679 , \43176 );
_HMUX g14de5 ( \43241_nG14de5 , \43239_nG14de3 , \43240_nG14de4 , \42599 );
buf \U$36934 ( \43242 , \43241_nG14de5 );
_DC g1aae2_GF_IsGateDCbyConstraint ( \43243_nG1aae2 , \43242 , \42503 );
buf \U$36935 ( \43244 , \43243_nG1aae2 );
_HMUX g14de6 ( \43245_nG14de6 , RIda0b288_3787 , \42685 , \43172 );
_HMUX g14de7 ( \43246_nG14de7 , RIda0b288_3787 , \43245_nG14de6 , \42590 );
_HMUX g14de8 ( \43247_nG14de8 , RIda0b288_3787 , \42688 , \43176 );
_HMUX g14de9 ( \43248_nG14de9 , \43246_nG14de7 , \43247_nG14de8 , \42599 );
buf \U$36936 ( \43249 , \43248_nG14de9 );
_DC g1aae4_GF_IsGateDCbyConstraint ( \43250_nG1aae4 , \43249 , \42503 );
buf \U$36937 ( \43251 , \43250_nG1aae4 );
_HMUX g14dea ( \43252_nG14dea , RId9f8d18_3788 , \42694 , \43172 );
_HMUX g14deb ( \43253_nG14deb , RId9f8d18_3788 , \43252_nG14dea , \42590 );
_HMUX g14dec ( \43254_nG14dec , RId9f8d18_3788 , \42697 , \43176 );
_HMUX g14ded ( \43255_nG14ded , \43253_nG14deb , \43254_nG14dec , \42599 );
buf \U$36938 ( \43256 , \43255_nG14ded );
_DC g1aae6_GF_IsGateDCbyConstraint ( \43257_nG1aae6 , \43256 , \42503 );
buf \U$36939 ( \43258 , \43257_nG1aae6 );
_HMUX g14dee ( \43259_nG14dee , RId9ec9a0_3789 , \42703 , \43172 );
_HMUX g14def ( \43260_nG14def , RId9ec9a0_3789 , \43259_nG14dee , \42590 );
_HMUX g14df0 ( \43261_nG14df0 , RId9ec9a0_3789 , \42706 , \43176 );
_HMUX g14df1 ( \43262_nG14df1 , \43260_nG14def , \43261_nG14df0 , \42599 );
buf \U$36940 ( \43263 , \43262_nG14df1 );
_DC g1aae8_GF_IsGateDCbyConstraint ( \43264_nG1aae8 , \43263 , \42503 );
buf \U$36941 ( \43265 , \43264_nG1aae8 );
_HMUX g14df2 ( \43266_nG14df2 , RId9e3418_3790 , \42712 , \43172 );
_HMUX g14df3 ( \43267_nG14df3 , RId9e3418_3790 , \43266_nG14df2 , \42590 );
_HMUX g14df4 ( \43268_nG14df4 , RId9e3418_3790 , \42715 , \43176 );
_HMUX g14df5 ( \43269_nG14df5 , \43267_nG14df3 , \43268_nG14df4 , \42599 );
buf \U$36942 ( \43270 , \43269_nG14df5 );
_DC g1aaea_GF_IsGateDCbyConstraint ( \43271_nG1aaea , \43270 , \42503 );
buf \U$36943 ( \43272 , \43271_nG1aaea );
_HMUX g14df6 ( \43273_nG14df6 , RIdb156a0_3791 , \42721 , \43172 );
_HMUX g14df7 ( \43274_nG14df7 , RIdb156a0_3791 , \43273_nG14df6 , \42590 );
_HMUX g14df8 ( \43275_nG14df8 , RIdb156a0_3791 , \42724 , \43176 );
_HMUX g14df9 ( \43276_nG14df9 , \43274_nG14df7 , \43275_nG14df8 , \42599 );
buf \U$36944 ( \43277 , \43276_nG14df9 );
_DC g1aaec_GF_IsGateDCbyConstraint ( \43278_nG1aaec , \43277 , \42503 );
buf \U$36945 ( \43279 , \43278_nG1aaec );
_HMUX g14dfa ( \43280_nG14dfa , RIdb17f68_3792 , \42730 , \43172 );
_HMUX g14dfb ( \43281_nG14dfb , RIdb17f68_3792 , \43280_nG14dfa , \42590 );
_HMUX g14dfc ( \43282_nG14dfc , RIdb17f68_3792 , \42733 , \43176 );
_HMUX g14dfd ( \43283_nG14dfd , \43281_nG14dfb , \43282_nG14dfc , \42599 );
buf \U$36946 ( \43284 , \43283_nG14dfd );
_DC g1aaee_GF_IsGateDCbyConstraint ( \43285_nG1aaee , \43284 , \42503 );
buf \U$36947 ( \43286 , \43285_nG1aaee );
_HMUX g14dfe ( \43287_nG14dfe , RIdb1b640_3793 , \42739 , \43172 );
_HMUX g14dff ( \43288_nG14dff , RIdb1b640_3793 , \43287_nG14dfe , \42590 );
_HMUX g14e00 ( \43289_nG14e00 , RIdb1b640_3793 , \42742 , \43176 );
_HMUX g14e01 ( \43290_nG14e01 , \43288_nG14dff , \43289_nG14e00 , \42599 );
buf \U$36948 ( \43291 , \43290_nG14e01 );
_DC g1aaf0_GF_IsGateDCbyConstraint ( \43292_nG1aaf0 , \43291 , \42503 );
buf \U$36949 ( \43293 , \43292_nG1aaf0 );
_HMUX g14e02 ( \43294_nG14e02 , RIdb1df08_3794 , \42748 , \43172 );
_HMUX g14e03 ( \43295_nG14e03 , RIdb1df08_3794 , \43294_nG14e02 , \42590 );
_HMUX g14e04 ( \43296_nG14e04 , RIdb1df08_3794 , \42751 , \43176 );
_HMUX g14e05 ( \43297_nG14e05 , \43295_nG14e03 , \43296_nG14e04 , \42599 );
buf \U$36950 ( \43298 , \43297_nG14e05 );
_DC g1aaf2_GF_IsGateDCbyConstraint ( \43299_nG1aaf2 , \43298 , \42503 );
buf \U$36951 ( \43300 , \43299_nG1aaf2 );
_HMUX g14e06 ( \43301_nG14e06 , RIdb215e0_3795 , \42757 , \43172 );
_HMUX g14e07 ( \43302_nG14e07 , RIdb215e0_3795 , \43301_nG14e06 , \42590 );
_HMUX g14e08 ( \43303_nG14e08 , RIdb215e0_3795 , \42760 , \43176 );
_HMUX g14e09 ( \43304_nG14e09 , \43302_nG14e07 , \43303_nG14e08 , \42599 );
buf \U$36952 ( \43305 , \43304_nG14e09 );
_DC g1aaf4_GF_IsGateDCbyConstraint ( \43306_nG1aaf4 , \43305 , \42503 );
buf \U$36953 ( \43307 , \43306_nG1aaf4 );
_HMUX g14e0a ( \43308_nG14e0a , RIdb23ea8_3796 , \42766 , \43172 );
_HMUX g14e0b ( \43309_nG14e0b , RIdb23ea8_3796 , \43308_nG14e0a , \42590 );
_HMUX g14e0c ( \43310_nG14e0c , RIdb23ea8_3796 , \42769 , \43176 );
_HMUX g14e0d ( \43311_nG14e0d , \43309_nG14e0b , \43310_nG14e0c , \42599 );
buf \U$36954 ( \43312 , \43311_nG14e0d );
_DC g1aaf8_GF_IsGateDCbyConstraint ( \43313_nG1aaf8 , \43312 , \42503 );
buf \U$36955 ( \43314 , \43313_nG1aaf8 );
_HMUX g14e0e ( \43315_nG14e0e , RIdb26c20_3797 , \42775 , \43172 );
_HMUX g14e0f ( \43316_nG14e0f , RIdb26c20_3797 , \43315_nG14e0e , \42590 );
_HMUX g14e10 ( \43317_nG14e10 , RIdb26c20_3797 , \42778 , \43176 );
_HMUX g14e11 ( \43318_nG14e11 , \43316_nG14e0f , \43317_nG14e10 , \42599 );
buf \U$36956 ( \43319 , \43318_nG14e11 );
_DC g1aafa_GF_IsGateDCbyConstraint ( \43320_nG1aafa , \43319 , \42503 );
buf \U$36957 ( \43321 , \43320_nG1aafa );
_HMUX g14e12 ( \43322_nG14e12 , RIdb29e48_3798 , \42784 , \43172 );
_HMUX g14e13 ( \43323_nG14e13 , RIdb29e48_3798 , \43322_nG14e12 , \42590 );
_HMUX g14e14 ( \43324_nG14e14 , RIdb29e48_3798 , \42787 , \43176 );
_HMUX g14e15 ( \43325_nG14e15 , \43323_nG14e13 , \43324_nG14e14 , \42599 );
buf \U$36958 ( \43326 , \43325_nG14e15 );
_DC g1aafc_GF_IsGateDCbyConstraint ( \43327_nG1aafc , \43326 , \42503 );
buf \U$36959 ( \43328 , \43327_nG1aafc );
_HMUX g14e16 ( \43329_nG14e16 , RIdb2cbc0_3799 , \42793 , \43172 );
_HMUX g14e17 ( \43330_nG14e17 , RIdb2cbc0_3799 , \43329_nG14e16 , \42590 );
_HMUX g14e18 ( \43331_nG14e18 , RIdb2cbc0_3799 , \42796 , \43176 );
_HMUX g14e19 ( \43332_nG14e19 , \43330_nG14e17 , \43331_nG14e18 , \42599 );
buf \U$36960 ( \43333 , \43332_nG14e19 );
_DC g1aafe_GF_IsGateDCbyConstraint ( \43334_nG1aafe , \43333 , \42503 );
buf \U$36961 ( \43335 , \43334_nG1aafe );
_HMUX g14e1a ( \43336_nG14e1a , RIdb2fde8_3800 , \42802 , \43172 );
_HMUX g14e1b ( \43337_nG14e1b , RIdb2fde8_3800 , \43336_nG14e1a , \42590 );
_HMUX g14e1c ( \43338_nG14e1c , RIdb2fde8_3800 , \42805 , \43176 );
_HMUX g14e1d ( \43339_nG14e1d , \43337_nG14e1b , \43338_nG14e1c , \42599 );
buf \U$36962 ( \43340 , \43339_nG14e1d );
_DC g1ab00_GF_IsGateDCbyConstraint ( \43341_nG1ab00 , \43340 , \42503 );
buf \U$36963 ( \43342 , \43341_nG1ab00 );
_HMUX g14e1e ( \43343_nG14e1e , RIdb32b60_3801 , \42811 , \43172 );
_HMUX g14e1f ( \43344_nG14e1f , RIdb32b60_3801 , \43343_nG14e1e , \42590 );
_HMUX g14e20 ( \43345_nG14e20 , RIdb32b60_3801 , \42814 , \43176 );
_HMUX g14e21 ( \43346_nG14e21 , \43344_nG14e1f , \43345_nG14e20 , \42599 );
buf \U$36964 ( \43347 , \43346_nG14e21 );
_DC g1ab02_GF_IsGateDCbyConstraint ( \43348_nG1ab02 , \43347 , \42503 );
buf \U$36965 ( \43349 , \43348_nG1ab02 );
_HMUX g14e22 ( \43350_nG14e22 , RIdb35d88_3802 , \42820 , \43172 );
_HMUX g14e23 ( \43351_nG14e23 , RIdb35d88_3802 , \43350_nG14e22 , \42590 );
_HMUX g14e24 ( \43352_nG14e24 , RIdb35d88_3802 , \42823 , \43176 );
_HMUX g14e25 ( \43353_nG14e25 , \43351_nG14e23 , \43352_nG14e24 , \42599 );
buf \U$36966 ( \43354 , \43353_nG14e25 );
_DC g1ab04_GF_IsGateDCbyConstraint ( \43355_nG1ab04 , \43354 , \42503 );
buf \U$36967 ( \43356 , \43355_nG1ab04 );
_HMUX g14e26 ( \43357_nG14e26 , RIdb38b00_3803 , \42829 , \43172 );
_HMUX g14e27 ( \43358_nG14e27 , RIdb38b00_3803 , \43357_nG14e26 , \42590 );
_HMUX g14e28 ( \43359_nG14e28 , RIdb38b00_3803 , \42832 , \43176 );
_HMUX g14e29 ( \43360_nG14e29 , \43358_nG14e27 , \43359_nG14e28 , \42599 );
buf \U$36968 ( \43361 , \43360_nG14e29 );
_DC g1ab06_GF_IsGateDCbyConstraint ( \43362_nG1ab06 , \43361 , \42503 );
buf \U$36969 ( \43363 , \43362_nG1ab06 );
_HMUX g14e2a ( \43364_nG14e2a , RIdb3b3c8_3804 , \42838 , \43172 );
_HMUX g14e2b ( \43365_nG14e2b , RIdb3b3c8_3804 , \43364_nG14e2a , \42590 );
_HMUX g14e2c ( \43366_nG14e2c , RIdb3b3c8_3804 , \42841 , \43176 );
_HMUX g14e2d ( \43367_nG14e2d , \43365_nG14e2b , \43366_nG14e2c , \42599 );
buf \U$36970 ( \43368 , \43367_nG14e2d );
_DC g1ab08_GF_IsGateDCbyConstraint ( \43369_nG1ab08 , \43368 , \42503 );
buf \U$36971 ( \43370 , \43369_nG1ab08 );
_HMUX g14e2e ( \43371_nG14e2e , RIdb3eaa0_3805 , \42847 , \43172 );
_HMUX g14e2f ( \43372_nG14e2f , RIdb3eaa0_3805 , \43371_nG14e2e , \42590 );
_HMUX g14e30 ( \43373_nG14e30 , RIdb3eaa0_3805 , \42850 , \43176 );
_HMUX g14e31 ( \43374_nG14e31 , \43372_nG14e2f , \43373_nG14e30 , \42599 );
buf \U$36972 ( \43375 , \43374_nG14e31 );
_DC g1ab0a_GF_IsGateDCbyConstraint ( \43376_nG1ab0a , \43375 , \42503 );
buf \U$36973 ( \43377 , \43376_nG1ab0a );
_HMUX g14e32 ( \43378_nG14e32 , RIdb404e0_3806 , \42856 , \43172 );
_HMUX g14e33 ( \43379_nG14e33 , RIdb404e0_3806 , \43378_nG14e32 , \42590 );
_HMUX g14e34 ( \43380_nG14e34 , RIdb404e0_3806 , \42859 , \43176 );
_HMUX g14e35 ( \43381_nG14e35 , \43379_nG14e33 , \43380_nG14e34 , \42599 );
buf \U$36974 ( \43382 , \43381_nG14e35 );
_DC g1ab0e_GF_IsGateDCbyConstraint ( \43383_nG1ab0e , \43382 , \42503 );
buf \U$36975 ( \43384 , \43383_nG1ab0e );
_HMUX g14e36 ( \43385_nG14e36 , RIdb422e0_3807 , \42865 , \43172 );
_HMUX g14e37 ( \43386_nG14e37 , RIdb422e0_3807 , \43385_nG14e36 , \42590 );
_HMUX g14e38 ( \43387_nG14e38 , RIdb422e0_3807 , \42868 , \43176 );
_HMUX g14e39 ( \43388_nG14e39 , \43386_nG14e37 , \43387_nG14e38 , \42599 );
buf \U$36976 ( \43389 , \43388_nG14e39 );
_DC g1ab10_GF_IsGateDCbyConstraint ( \43390_nG1ab10 , \43389 , \42503 );
buf \U$36977 ( \43391 , \43390_nG1ab10 );
_HMUX g14e3a ( \43392_nG14e3a , RIdb43ac8_3808 , \42874 , \43172 );
_HMUX g14e3b ( \43393_nG14e3b , RIdb43ac8_3808 , \43392_nG14e3a , \42590 );
_HMUX g14e3c ( \43394_nG14e3c , RIdb43ac8_3808 , \42877 , \43176 );
_HMUX g14e3d ( \43395_nG14e3d , \43393_nG14e3b , \43394_nG14e3c , \42599 );
buf \U$36978 ( \43396 , \43395_nG14e3d );
_DC g1ab12_GF_IsGateDCbyConstraint ( \43397_nG1ab12 , \43396 , \42503 );
buf \U$36979 ( \43398 , \43397_nG1ab12 );
_HMUX g14e3e ( \43399_nG14e3e , RIdb45850_3809 , \42883 , \43172 );
_HMUX g14e3f ( \43400_nG14e3f , RIdb45850_3809 , \43399_nG14e3e , \42590 );
_HMUX g14e40 ( \43401_nG14e40 , RIdb45850_3809 , \42886 , \43176 );
_HMUX g14e41 ( \43402_nG14e41 , \43400_nG14e3f , \43401_nG14e40 , \42599 );
buf \U$36980 ( \43403 , \43402_nG14e41 );
_DC g1ab14_GF_IsGateDCbyConstraint ( \43404_nG1ab14 , \43403 , \42503 );
buf \U$36981 ( \43405 , \43404_nG1ab14 );
_HMUX g14e42 ( \43406_nG14e42 , RIdb47128_3810 , \42892 , \43172 );
_HMUX g14e43 ( \43407_nG14e43 , RIdb47128_3810 , \43406_nG14e42 , \42590 );
_HMUX g14e44 ( \43408_nG14e44 , RIdb47128_3810 , \42895 , \43176 );
_HMUX g14e45 ( \43409_nG14e45 , \43407_nG14e43 , \43408_nG14e44 , \42599 );
buf \U$36982 ( \43410 , \43409_nG14e45 );
_DC g1ab16_GF_IsGateDCbyConstraint ( \43411_nG1ab16 , \43410 , \42503 );
buf \U$36983 ( \43412 , \43411_nG1ab16 );
_HMUX g14e46 ( \43413_nG14e46 , RIdb483e8_3811 , \42901 , \43172 );
_HMUX g14e47 ( \43414_nG14e47 , RIdb483e8_3811 , \43413_nG14e46 , \42590 );
_HMUX g14e48 ( \43415_nG14e48 , RIdb483e8_3811 , \42904 , \43176 );
_HMUX g14e49 ( \43416_nG14e49 , \43414_nG14e47 , \43415_nG14e48 , \42599 );
buf \U$36984 ( \43417 , \43416_nG14e49 );
_DC g1ab18_GF_IsGateDCbyConstraint ( \43418_nG1ab18 , \43417 , \42503 );
buf \U$36985 ( \43419 , \43418_nG1ab18 );
_HMUX g14e4a ( \43420_nG14e4a , RIdb49888_3812 , \42910 , \43172 );
_HMUX g14e4b ( \43421_nG14e4b , RIdb49888_3812 , \43420_nG14e4a , \42590 );
_HMUX g14e4c ( \43422_nG14e4c , RIdb49888_3812 , \42913 , \43176 );
_HMUX g14e4d ( \43423_nG14e4d , \43421_nG14e4b , \43422_nG14e4c , \42599 );
buf \U$36986 ( \43424 , \43423_nG14e4d );
_DC g1ab1a_GF_IsGateDCbyConstraint ( \43425_nG1ab1a , \43424 , \42503 );
buf \U$36987 ( \43426 , \43425_nG1ab1a );
_HMUX g14e4e ( \43427_nG14e4e , RIdb4abc0_3813 , \42919 , \43172 );
_HMUX g14e4f ( \43428_nG14e4f , RIdb4abc0_3813 , \43427_nG14e4e , \42590 );
_HMUX g14e50 ( \43429_nG14e50 , RIdb4abc0_3813 , \42922 , \43176 );
_HMUX g14e51 ( \43430_nG14e51 , \43428_nG14e4f , \43429_nG14e50 , \42599 );
buf \U$36988 ( \43431 , \43430_nG14e51 );
_DC g1ab1c_GF_IsGateDCbyConstraint ( \43432_nG1ab1c , \43431 , \42503 );
buf \U$36989 ( \43433 , \43432_nG1ab1c );
_HMUX g14e52 ( \43434_nG14e52 , RIdb4c330_3814 , \42928 , \43172 );
_HMUX g14e53 ( \43435_nG14e53 , RIdb4c330_3814 , \43434_nG14e52 , \42590 );
_HMUX g14e54 ( \43436_nG14e54 , RIdb4c330_3814 , \42931 , \43176 );
_HMUX g14e55 ( \43437_nG14e55 , \43435_nG14e53 , \43436_nG14e54 , \42599 );
buf \U$36990 ( \43438 , \43437_nG14e55 );
_DC g1ab1e_GF_IsGateDCbyConstraint ( \43439_nG1ab1e , \43438 , \42503 );
buf \U$36991 ( \43440 , \43439_nG1ab1e );
_HMUX g14e56 ( \43441_nG14e56 , RIdb4d410_3815 , \42937 , \43172 );
_HMUX g14e57 ( \43442_nG14e57 , RIdb4d410_3815 , \43441_nG14e56 , \42590 );
_HMUX g14e58 ( \43443_nG14e58 , RIdb4d410_3815 , \42940 , \43176 );
_HMUX g14e59 ( \43444_nG14e59 , \43442_nG14e57 , \43443_nG14e58 , \42599 );
buf \U$36992 ( \43445 , \43444_nG14e59 );
_DC g1ab20_GF_IsGateDCbyConstraint ( \43446_nG1ab20 , \43445 , \42503 );
buf \U$36993 ( \43447 , \43446_nG1ab20 );
_HMUX g14e5a ( \43448_nG14e5a , RIdb4e5e0_3816 , \42946 , \43172 );
_HMUX g14e5b ( \43449_nG14e5b , RIdb4e5e0_3816 , \43448_nG14e5a , \42590 );
_HMUX g14e5c ( \43450_nG14e5c , RIdb4e5e0_3816 , \42949 , \43176 );
_HMUX g14e5d ( \43451_nG14e5d , \43449_nG14e5b , \43450_nG14e5c , \42599 );
buf \U$36994 ( \43452 , \43451_nG14e5d );
_DC g1ab24_GF_IsGateDCbyConstraint ( \43453_nG1ab24 , \43452 , \42503 );
buf \U$36995 ( \43454 , \43453_nG1ab24 );
_HMUX g14e5e ( \43455_nG14e5e , RIdb4fa08_3817 , \42955 , \43172 );
_HMUX g14e5f ( \43456_nG14e5f , RIdb4fa08_3817 , \43455_nG14e5e , \42590 );
_HMUX g14e60 ( \43457_nG14e60 , RIdb4fa08_3817 , \42958 , \43176 );
_HMUX g14e61 ( \43458_nG14e61 , \43456_nG14e5f , \43457_nG14e60 , \42599 );
buf \U$36996 ( \43459 , \43458_nG14e61 );
_DC g1ab26_GF_IsGateDCbyConstraint ( \43460_nG1ab26 , \43459 , \42503 );
buf \U$36997 ( \43461 , \43460_nG1ab26 );
_HMUX g14e62 ( \43462_nG14e62 , RIdb51100_3818 , \42964 , \43172 );
_HMUX g14e63 ( \43463_nG14e63 , RIdb51100_3818 , \43462_nG14e62 , \42590 );
_HMUX g14e64 ( \43464_nG14e64 , RIdb51100_3818 , \42967 , \43176 );
_HMUX g14e65 ( \43465_nG14e65 , \43463_nG14e63 , \43464_nG14e64 , \42599 );
buf \U$36998 ( \43466 , \43465_nG14e65 );
_DC g1ab28_GF_IsGateDCbyConstraint ( \43467_nG1ab28 , \43466 , \42503 );
buf \U$36999 ( \43468 , \43467_nG1ab28 );
_HMUX g14e66 ( \43469_nG14e66 , RIdb52c30_3819 , \42973 , \43172 );
_HMUX g14e67 ( \43470_nG14e67 , RIdb52c30_3819 , \43469_nG14e66 , \42590 );
_HMUX g14e68 ( \43471_nG14e68 , RIdb52c30_3819 , \42976 , \43176 );
_HMUX g14e69 ( \43472_nG14e69 , \43470_nG14e67 , \43471_nG14e68 , \42599 );
buf \U$37000 ( \43473 , \43472_nG14e69 );
_DC g1ab2a_GF_IsGateDCbyConstraint ( \43474_nG1ab2a , \43473 , \42503 );
buf \U$37001 ( \43475 , \43474_nG1ab2a );
_HMUX g14e6a ( \43476_nG14e6a , RIdb541c0_3820 , \42982 , \43172 );
_HMUX g14e6b ( \43477_nG14e6b , RIdb541c0_3820 , \43476_nG14e6a , \42590 );
_HMUX g14e6c ( \43478_nG14e6c , RIdb541c0_3820 , \42985 , \43176 );
_HMUX g14e6d ( \43479_nG14e6d , \43477_nG14e6b , \43478_nG14e6c , \42599 );
buf \U$37002 ( \43480 , \43479_nG14e6d );
_DC g1ab2c_GF_IsGateDCbyConstraint ( \43481_nG1ab2c , \43480 , \42503 );
buf \U$37003 ( \43482 , \43481_nG1ab2c );
_HMUX g14e6e ( \43483_nG14e6e , RIdb559a8_3821 , \42991 , \43172 );
_HMUX g14e6f ( \43484_nG14e6f , RIdb559a8_3821 , \43483_nG14e6e , \42590 );
_HMUX g14e70 ( \43485_nG14e70 , RIdb559a8_3821 , \42994 , \43176 );
_HMUX g14e71 ( \43486_nG14e71 , \43484_nG14e6f , \43485_nG14e70 , \42599 );
buf \U$37004 ( \43487 , \43486_nG14e71 );
_DC g1ab2e_GF_IsGateDCbyConstraint ( \43488_nG1ab2e , \43487 , \42503 );
buf \U$37005 ( \43489 , \43488_nG1ab2e );
_HMUX g14e72 ( \43490_nG14e72 , RIdb56e48_3822 , \43000 , \43172 );
_HMUX g14e73 ( \43491_nG14e73 , RIdb56e48_3822 , \43490_nG14e72 , \42590 );
_HMUX g14e74 ( \43492_nG14e74 , RIdb56e48_3822 , \43003 , \43176 );
_HMUX g14e75 ( \43493_nG14e75 , \43491_nG14e73 , \43492_nG14e74 , \42599 );
buf \U$37006 ( \43494 , \43493_nG14e75 );
_DC g1ab30_GF_IsGateDCbyConstraint ( \43495_nG1ab30 , \43494 , \42503 );
buf \U$37007 ( \43496 , \43495_nG1ab30 );
_HMUX g14e76 ( \43497_nG14e76 , RIdb58900_3823 , \43009 , \43172 );
_HMUX g14e77 ( \43498_nG14e77 , RIdb58900_3823 , \43497_nG14e76 , \42590 );
_HMUX g14e78 ( \43499_nG14e78 , RIdb58900_3823 , \43012 , \43176 );
_HMUX g14e79 ( \43500_nG14e79 , \43498_nG14e77 , \43499_nG14e78 , \42599 );
buf \U$37008 ( \43501 , \43500_nG14e79 );
_DC g1ab32_GF_IsGateDCbyConstraint ( \43502_nG1ab32 , \43501 , \42503 );
buf \U$37009 ( \43503 , \43502_nG1ab32 );
_HMUX g14e7a ( \43504_nG14e7a , RIdb5a070_3824 , \43018 , \43172 );
_HMUX g14e7b ( \43505_nG14e7b , RIdb5a070_3824 , \43504_nG14e7a , \42590 );
_HMUX g14e7c ( \43506_nG14e7c , RIdb5a070_3824 , \43021 , \43176 );
_HMUX g14e7d ( \43507_nG14e7d , \43505_nG14e7b , \43506_nG14e7c , \42599 );
buf \U$37010 ( \43508 , \43507_nG14e7d );
_DC g1ab34_GF_IsGateDCbyConstraint ( \43509_nG1ab34 , \43508 , \42503 );
buf \U$37011 ( \43510 , \43509_nG1ab34 );
_HMUX g14e7e ( \43511_nG14e7e , RIdb5b588_3825 , \43027 , \43172 );
_HMUX g14e7f ( \43512_nG14e7f , RIdb5b588_3825 , \43511_nG14e7e , \42590 );
_HMUX g14e80 ( \43513_nG14e80 , RIdb5b588_3825 , \43030 , \43176 );
_HMUX g14e81 ( \43514_nG14e81 , \43512_nG14e7f , \43513_nG14e80 , \42599 );
buf \U$37012 ( \43515 , \43514_nG14e81 );
_DC g1ab36_GF_IsGateDCbyConstraint ( \43516_nG1ab36 , \43515 , \42503 );
buf \U$37013 ( \43517 , \43516_nG1ab36 );
_HMUX g14e82 ( \43518_nG14e82 , RIdb5d0b8_3826 , \43036 , \43172 );
_HMUX g14e83 ( \43519_nG14e83 , RIdb5d0b8_3826 , \43518_nG14e82 , \42590 );
_HMUX g14e84 ( \43520_nG14e84 , RIdb5d0b8_3826 , \43039 , \43176 );
_HMUX g14e85 ( \43521_nG14e85 , \43519_nG14e83 , \43520_nG14e84 , \42599 );
buf \U$37014 ( \43522 , \43521_nG14e85 );
_DC g1ab3a_GF_IsGateDCbyConstraint ( \43523_nG1ab3a , \43522 , \42503 );
buf \U$37015 ( \43524 , \43523_nG1ab3a );
_HMUX g14e86 ( \43525_nG14e86 , RIdb5e3f0_3827 , \43045 , \43172 );
_HMUX g14e87 ( \43526_nG14e87 , RIdb5e3f0_3827 , \43525_nG14e86 , \42590 );
_HMUX g14e88 ( \43527_nG14e88 , RIdb5e3f0_3827 , \43048 , \43176 );
_HMUX g14e89 ( \43528_nG14e89 , \43526_nG14e87 , \43527_nG14e88 , \42599 );
buf \U$37016 ( \43529 , \43528_nG14e89 );
_DC g1ab3c_GF_IsGateDCbyConstraint ( \43530_nG1ab3c , \43529 , \42503 );
buf \U$37017 ( \43531 , \43530_nG1ab3c );
_HMUX g14e8a ( \43532_nG14e8a , RIda95720_3828 , \43054 , \43172 );
_HMUX g14e8b ( \43533_nG14e8b , RIda95720_3828 , \43532_nG14e8a , \42590 );
_HMUX g14e8c ( \43534_nG14e8c , RIda95720_3828 , \43057 , \43176 );
_HMUX g14e8d ( \43535_nG14e8d , \43533_nG14e8b , \43534_nG14e8c , \42599 );
buf \U$37018 ( \43536 , \43535_nG14e8d );
_DC g1ab3e_GF_IsGateDCbyConstraint ( \43537_nG1ab3e , \43536 , \42503 );
buf \U$37019 ( \43538 , \43537_nG1ab3e );
_HMUX g14e8e ( \43539_nG14e8e , RIda97598_3829 , \43063 , \43172 );
_HMUX g14e8f ( \43540_nG14e8f , RIda97598_3829 , \43539_nG14e8e , \42590 );
_HMUX g14e90 ( \43541_nG14e90 , RIda97598_3829 , \43066 , \43176 );
_HMUX g14e91 ( \43542_nG14e91 , \43540_nG14e8f , \43541_nG14e90 , \42599 );
buf \U$37020 ( \43543 , \43542_nG14e91 );
_DC g1ab40_GF_IsGateDCbyConstraint ( \43544_nG1ab40 , \43543 , \42503 );
buf \U$37021 ( \43545 , \43544_nG1ab40 );
_HMUX g14e92 ( \43546_nG14e92 , RIda99a28_3830 , \43072 , \43172 );
_HMUX g14e93 ( \43547_nG14e93 , RIda99a28_3830 , \43546_nG14e92 , \42590 );
_HMUX g14e94 ( \43548_nG14e94 , RIda99a28_3830 , \43075 , \43176 );
_HMUX g14e95 ( \43549_nG14e95 , \43547_nG14e93 , \43548_nG14e94 , \42599 );
buf \U$37022 ( \43550 , \43549_nG14e95 );
_DC g1ab42_GF_IsGateDCbyConstraint ( \43551_nG1ab42 , \43550 , \42503 );
buf \U$37023 ( \43552 , \43551_nG1ab42 );
_HMUX g14e96 ( \43553_nG14e96 , RIda9bd50_3831 , \43081 , \43172 );
_HMUX g14e97 ( \43554_nG14e97 , RIda9bd50_3831 , \43553_nG14e96 , \42590 );
_HMUX g14e98 ( \43555_nG14e98 , RIda9bd50_3831 , \43084 , \43176 );
_HMUX g14e99 ( \43556_nG14e99 , \43554_nG14e97 , \43555_nG14e98 , \42599 );
buf \U$37024 ( \43557 , \43556_nG14e99 );
_DC g1ab44_GF_IsGateDCbyConstraint ( \43558_nG1ab44 , \43557 , \42503 );
buf \U$37025 ( \43559 , \43558_nG1ab44 );
_HMUX g14e9a ( \43560_nG14e9a , RIda9df10_3832 , \43090 , \43172 );
_HMUX g14e9b ( \43561_nG14e9b , RIda9df10_3832 , \43560_nG14e9a , \42590 );
_HMUX g14e9c ( \43562_nG14e9c , RIda9df10_3832 , \43093 , \43176 );
_HMUX g14e9d ( \43563_nG14e9d , \43561_nG14e9b , \43562_nG14e9c , \42599 );
buf \U$37026 ( \43564 , \43563_nG14e9d );
_DC g1ab46_GF_IsGateDCbyConstraint ( \43565_nG1ab46 , \43564 , \42503 );
buf \U$37027 ( \43566 , \43565_nG1ab46 );
_HMUX g14e9e ( \43567_nG14e9e , RIda9f4a0_3833 , \43099 , \43172 );
_HMUX g14e9f ( \43568_nG14e9f , RIda9f4a0_3833 , \43567_nG14e9e , \42590 );
_HMUX g14ea0 ( \43569_nG14ea0 , RIda9f4a0_3833 , \43102 , \43176 );
_HMUX g14ea1 ( \43570_nG14ea1 , \43568_nG14e9f , \43569_nG14ea0 , \42599 );
buf \U$37028 ( \43571 , \43570_nG14ea1 );
_DC g1ab48_GF_IsGateDCbyConstraint ( \43572_nG1ab48 , \43571 , \42503 );
buf \U$37029 ( \43573 , \43572_nG1ab48 );
_HMUX g14ea2 ( \43574_nG14ea2 , RIdaa1228_3834 , \43108 , \43172 );
_HMUX g14ea3 ( \43575_nG14ea3 , RIdaa1228_3834 , \43574_nG14ea2 , \42590 );
_HMUX g14ea4 ( \43576_nG14ea4 , RIdaa1228_3834 , \43111 , \43176 );
_HMUX g14ea5 ( \43577_nG14ea5 , \43575_nG14ea3 , \43576_nG14ea4 , \42599 );
buf \U$37030 ( \43578 , \43577_nG14ea5 );
_DC g1ab4a_GF_IsGateDCbyConstraint ( \43579_nG1ab4a , \43578 , \42503 );
buf \U$37031 ( \43580 , \43579_nG1ab4a );
_HMUX g14ea6 ( \43581_nG14ea6 , RIdaa2d58_3835 , \43117 , \43172 );
_HMUX g14ea7 ( \43582_nG14ea7 , RIdaa2d58_3835 , \43581_nG14ea6 , \42590 );
_HMUX g14ea8 ( \43583_nG14ea8 , RIdaa2d58_3835 , \43120 , \43176 );
_HMUX g14ea9 ( \43584_nG14ea9 , \43582_nG14ea7 , \43583_nG14ea8 , \42599 );
buf \U$37032 ( \43585 , \43584_nG14ea9 );
_DC g1ab4c_GF_IsGateDCbyConstraint ( \43586_nG1ab4c , \43585 , \42503 );
buf \U$37033 ( \43587 , \43586_nG1ab4c );
_HMUX g14eaa ( \43588_nG14eaa , RIdaa4a68_3836 , \43126 , \43172 );
_HMUX g14eab ( \43589_nG14eab , RIdaa4a68_3836 , \43588_nG14eaa , \42590 );
_HMUX g14eac ( \43590_nG14eac , RIdaa4a68_3836 , \43129 , \43176 );
_HMUX g14ead ( \43591_nG14ead , \43589_nG14eab , \43590_nG14eac , \42599 );
buf \U$37034 ( \43592 , \43591_nG14ead );
_DC g1ab50_GF_IsGateDCbyConstraint ( \43593_nG1ab50 , \43592 , \42503 );
buf \U$37035 ( \43594 , \43593_nG1ab50 );
_HMUX g14eae ( \43595_nG14eae , RIdaa6b38_3837 , \43135 , \43172 );
_HMUX g14eaf ( \43596_nG14eaf , RIdaa6b38_3837 , \43595_nG14eae , \42590 );
_HMUX g14eb0 ( \43597_nG14eb0 , RIdaa6b38_3837 , \43138 , \43176 );
_HMUX g14eb1 ( \43598_nG14eb1 , \43596_nG14eaf , \43597_nG14eb0 , \42599 );
buf \U$37036 ( \43599 , \43598_nG14eb1 );
_DC g1ab52_GF_IsGateDCbyConstraint ( \43600_nG1ab52 , \43599 , \42503 );
buf \U$37037 ( \43601 , \43600_nG1ab52 );
_HMUX g14eb2 ( \43602_nG14eb2 , RIdaa89b0_3838 , \43144 , \43172 );
_HMUX g14eb3 ( \43603_nG14eb3 , RIdaa89b0_3838 , \43602_nG14eb2 , \42590 );
_HMUX g14eb4 ( \43604_nG14eb4 , RIdaa89b0_3838 , \43147 , \43176 );
_HMUX g14eb5 ( \43605_nG14eb5 , \43603_nG14eb3 , \43604_nG14eb4 , \42599 );
buf \U$37038 ( \43606 , \43605_nG14eb5 );
_DC g1ab54_GF_IsGateDCbyConstraint ( \43607_nG1ab54 , \43606 , \42503 );
buf \U$37039 ( \43608 , \43607_nG1ab54 );
_HMUX g14eb6 ( \43609_nG14eb6 , RIdbdf030_3839 , \43153 , \43172 );
_HMUX g14eb7 ( \43610_nG14eb7 , RIdbdf030_3839 , \43609_nG14eb6 , \42590 );
_HMUX g14eb8 ( \43611_nG14eb8 , RIdbdf030_3839 , \43156 , \43176 );
_HMUX g14eb9 ( \43612_nG14eb9 , \43610_nG14eb7 , \43611_nG14eb8 , \42599 );
buf \U$37040 ( \43613 , \43612_nG14eb9 );
_DC g1ab56_GF_IsGateDCbyConstraint ( \43614_nG1ab56 , \43613 , \42503 );
buf \U$37041 ( \43615 , \43614_nG1ab56 );
_HMUX g14eba ( \43616_nG14eba , RIdbdcd80_3840 , \43162 , \43172 );
_HMUX g14ebb ( \43617_nG14ebb , RIdbdcd80_3840 , \43616_nG14eba , \42590 );
_HMUX g14ebc ( \43618_nG14ebc , RIdbdcd80_3840 , \43165 , \43176 );
_HMUX g14ebd ( \43619_nG14ebd , \43617_nG14ebb , \43618_nG14ebc , \42599 );
buf \U$37042 ( \43620 , \43619_nG14ebd );
_DC g1ab58_GF_IsGateDCbyConstraint ( \43621_nG1ab58 , \43620 , \42503 );
buf \U$37043 ( \43622 , \43621_nG1ab58 );
nor \U$37044 ( \43623 , \42579 , \43171 );
_HMUX g14cbb ( \43624_nG14cbb , RIdbdaff8_3841 , \42578 , \43623 );
_HMUX g14cbc ( \43625_nG14cbc , RIdbdaff8_3841 , \43624_nG14cbb , \42590 );
nor \U$37045 ( \43626 , \42593 , \43175 );
_HMUX g14cbf ( \43627_nG14cbf , RIdbdaff8_3841 , \42592 , \43626 );
_HMUX g14cc0 ( \43628_nG14cc0 , \43625_nG14cbc , \43627_nG14cbf , \42599 );
buf \U$37046 ( \43629 , \43628_nG14cc0 );
_DC g1aa60_GF_IsGateDCbyConstraint ( \43630_nG1aa60 , \43629 , \42503 );
buf \U$37047 ( \43631 , \43630_nG1aa60 );
_HMUX g14cc1 ( \43632_nG14cc1 , RIdbd9540_3842 , \42604 , \43623 );
_HMUX g14cc2 ( \43633_nG14cc2 , RIdbd9540_3842 , \43632_nG14cc1 , \42590 );
_HMUX g14cc3 ( \43634_nG14cc3 , RIdbd9540_3842 , \42607 , \43626 );
_HMUX g14cc4 ( \43635_nG14cc4 , \43633_nG14cc2 , \43634_nG14cc3 , \42599 );
buf \U$37048 ( \43636 , \43635_nG14cc4 );
_DC g1aa76_GF_IsGateDCbyConstraint ( \43637_nG1aa76 , \43636 , \42503 );
buf \U$37049 ( \43638 , \43637_nG1aa76 );
_HMUX g14cc5 ( \43639_nG14cc5 , RIdbd6e58_3843 , \42613 , \43623 );
_HMUX g14cc6 ( \43640_nG14cc6 , RIdbd6e58_3843 , \43639_nG14cc5 , \42590 );
_HMUX g14cc7 ( \43641_nG14cc7 , RIdbd6e58_3843 , \42616 , \43626 );
_HMUX g14cc8 ( \43642_nG14cc8 , \43640_nG14cc6 , \43641_nG14cc7 , \42599 );
buf \U$37050 ( \43643 , \43642_nG14cc8 );
_DC g1aa8c_GF_IsGateDCbyConstraint ( \43644_nG1aa8c , \43643 , \42503 );
buf \U$37051 ( \43645 , \43644_nG1aa8c );
_HMUX g14cc9 ( \43646_nG14cc9 , RIdbd4860_3844 , \42622 , \43623 );
_HMUX g14cca ( \43647_nG14cca , RIdbd4860_3844 , \43646_nG14cc9 , \42590 );
_HMUX g14ccb ( \43648_nG14ccb , RIdbd4860_3844 , \42625 , \43626 );
_HMUX g14ccc ( \43649_nG14ccc , \43647_nG14cca , \43648_nG14ccb , \42599 );
buf \U$37052 ( \43650 , \43649_nG14ccc );
_DC g1aaa2_GF_IsGateDCbyConstraint ( \43651_nG1aaa2 , \43650 , \42503 );
buf \U$37053 ( \43652 , \43651_nG1aaa2 );
_HMUX g14ccd ( \43653_nG14ccd , RIdbd25b0_3845 , \42631 , \43623 );
_HMUX g14cce ( \43654_nG14cce , RIdbd25b0_3845 , \43653_nG14ccd , \42590 );
_HMUX g14ccf ( \43655_nG14ccf , RIdbd25b0_3845 , \42634 , \43626 );
_HMUX g14cd0 ( \43656_nG14cd0 , \43654_nG14cce , \43655_nG14ccf , \42599 );
buf \U$37054 ( \43657 , \43656_nG14cd0 );
_DC g1aab8_GF_IsGateDCbyConstraint ( \43658_nG1aab8 , \43657 , \42503 );
buf \U$37055 ( \43659 , \43658_nG1aab8 );
_HMUX g14cd1 ( \43660_nG14cd1 , RIdbd0030_3846 , \42640 , \43623 );
_HMUX g14cd2 ( \43661_nG14cd2 , RIdbd0030_3846 , \43660_nG14cd1 , \42590 );
_HMUX g14cd3 ( \43662_nG14cd3 , RIdbd0030_3846 , \42643 , \43626 );
_HMUX g14cd4 ( \43663_nG14cd4 , \43661_nG14cd2 , \43662_nG14cd3 , \42599 );
buf \U$37056 ( \43664 , \43663_nG14cd4 );
_DC g1aace_GF_IsGateDCbyConstraint ( \43665_nG1aace , \43664 , \42503 );
buf \U$37057 ( \43666 , \43665_nG1aace );
_HMUX g14cd5 ( \43667_nG14cd5 , RIdbcdc18_3847 , \42649 , \43623 );
_HMUX g14cd6 ( \43668_nG14cd6 , RIdbcdc18_3847 , \43667_nG14cd5 , \42590 );
_HMUX g14cd7 ( \43669_nG14cd7 , RIdbcdc18_3847 , \42652 , \43626 );
_HMUX g14cd8 ( \43670_nG14cd8 , \43668_nG14cd6 , \43669_nG14cd7 , \42599 );
buf \U$37058 ( \43671 , \43670_nG14cd8 );
_DC g1aada_GF_IsGateDCbyConstraint ( \43672_nG1aada , \43671 , \42503 );
buf \U$37059 ( \43673 , \43672_nG1aada );
_HMUX g14cd9 ( \43674_nG14cd9 , RIdbcb800_3848 , \42658 , \43623 );
_HMUX g14cda ( \43675_nG14cda , RIdbcb800_3848 , \43674_nG14cd9 , \42590 );
_HMUX g14cdb ( \43676_nG14cdb , RIdbcb800_3848 , \42661 , \43626 );
_HMUX g14cdc ( \43677_nG14cdc , \43675_nG14cda , \43676_nG14cdb , \42599 );
buf \U$37060 ( \43678 , \43677_nG14cdc );
_DC g1aadc_GF_IsGateDCbyConstraint ( \43679_nG1aadc , \43678 , \42503 );
buf \U$37061 ( \43680 , \43679_nG1aadc );
_HMUX g14cdd ( \43681_nG14cdd , RIdbc9730_3849 , \42667 , \43623 );
_HMUX g14cde ( \43682_nG14cde , RIdbc9730_3849 , \43681_nG14cdd , \42590 );
_HMUX g14cdf ( \43683_nG14cdf , RIdbc9730_3849 , \42670 , \43626 );
_HMUX g14ce0 ( \43684_nG14ce0 , \43682_nG14cde , \43683_nG14cdf , \42599 );
buf \U$37062 ( \43685 , \43684_nG14ce0 );
_DC g1aade_GF_IsGateDCbyConstraint ( \43686_nG1aade , \43685 , \42503 );
buf \U$37063 ( \43687 , \43686_nG1aade );
_HMUX g14ce1 ( \43688_nG14ce1 , RIdbc7a20_3850 , \42676 , \43623 );
_HMUX g14ce2 ( \43689_nG14ce2 , RIdbc7a20_3850 , \43688_nG14ce1 , \42590 );
_HMUX g14ce3 ( \43690_nG14ce3 , RIdbc7a20_3850 , \42679 , \43626 );
_HMUX g14ce4 ( \43691_nG14ce4 , \43689_nG14ce2 , \43690_nG14ce3 , \42599 );
buf \U$37064 ( \43692 , \43691_nG14ce4 );
_DC g1aa62_GF_IsGateDCbyConstraint ( \43693_nG1aa62 , \43692 , \42503 );
buf \U$37065 ( \43694 , \43693_nG1aa62 );
_HMUX g14ce5 ( \43695_nG14ce5 , RIdbc5e78_3851 , \42685 , \43623 );
_HMUX g14ce6 ( \43696_nG14ce6 , RIdbc5e78_3851 , \43695_nG14ce5 , \42590 );
_HMUX g14ce7 ( \43697_nG14ce7 , RIdbc5e78_3851 , \42688 , \43626 );
_HMUX g14ce8 ( \43698_nG14ce8 , \43696_nG14ce6 , \43697_nG14ce7 , \42599 );
buf \U$37066 ( \43699 , \43698_nG14ce8 );
_DC g1aa64_GF_IsGateDCbyConstraint ( \43700_nG1aa64 , \43699 , \42503 );
buf \U$37067 ( \43701 , \43700_nG1aa64 );
_HMUX g14ce9 ( \43702_nG14ce9 , RIdbc40f0_3852 , \42694 , \43623 );
_HMUX g14cea ( \43703_nG14cea , RIdbc40f0_3852 , \43702_nG14ce9 , \42590 );
_HMUX g14ceb ( \43704_nG14ceb , RIdbc40f0_3852 , \42697 , \43626 );
_HMUX g14cec ( \43705_nG14cec , \43703_nG14cea , \43704_nG14ceb , \42599 );
buf \U$37068 ( \43706 , \43705_nG14cec );
_DC g1aa66_GF_IsGateDCbyConstraint ( \43707_nG1aa66 , \43706 , \42503 );
buf \U$37069 ( \43708 , \43707_nG1aa66 );
_HMUX g14ced ( \43709_nG14ced , RIdbc1f30_3853 , \42703 , \43623 );
_HMUX g14cee ( \43710_nG14cee , RIdbc1f30_3853 , \43709_nG14ced , \42590 );
_HMUX g14cef ( \43711_nG14cef , RIdbc1f30_3853 , \42706 , \43626 );
_HMUX g14cf0 ( \43712_nG14cf0 , \43710_nG14cee , \43711_nG14cef , \42599 );
buf \U$37070 ( \43713 , \43712_nG14cf0 );
_DC g1aa68_GF_IsGateDCbyConstraint ( \43714_nG1aa68 , \43713 , \42503 );
buf \U$37071 ( \43715 , \43714_nG1aa68 );
_HMUX g14cf1 ( \43716_nG14cf1 , RIdbbf938_3854 , \42712 , \43623 );
_HMUX g14cf2 ( \43717_nG14cf2 , RIdbbf938_3854 , \43716_nG14cf1 , \42590 );
_HMUX g14cf3 ( \43718_nG14cf3 , RIdbbf938_3854 , \42715 , \43626 );
_HMUX g14cf4 ( \43719_nG14cf4 , \43717_nG14cf2 , \43718_nG14cf3 , \42599 );
buf \U$37072 ( \43720 , \43719_nG14cf4 );
_DC g1aa6a_GF_IsGateDCbyConstraint ( \43721_nG1aa6a , \43720 , \42503 );
buf \U$37073 ( \43722 , \43721_nG1aa6a );
_HMUX g14cf5 ( \43723_nG14cf5 , RIdbbd4a8_3855 , \42721 , \43623 );
_HMUX g14cf6 ( \43724_nG14cf6 , RIdbbd4a8_3855 , \43723_nG14cf5 , \42590 );
_HMUX g14cf7 ( \43725_nG14cf7 , RIdbbd4a8_3855 , \42724 , \43626 );
_HMUX g14cf8 ( \43726_nG14cf8 , \43724_nG14cf6 , \43725_nG14cf7 , \42599 );
buf \U$37074 ( \43727 , \43726_nG14cf8 );
_DC g1aa6c_GF_IsGateDCbyConstraint ( \43728_nG1aa6c , \43727 , \42503 );
buf \U$37075 ( \43729 , \43728_nG1aa6c );
_HMUX g14cf9 ( \43730_nG14cf9 , RIdbba910_3856 , \42730 , \43623 );
_HMUX g14cfa ( \43731_nG14cfa , RIdbba910_3856 , \43730_nG14cf9 , \42590 );
_HMUX g14cfb ( \43732_nG14cfb , RIdbba910_3856 , \42733 , \43626 );
_HMUX g14cfc ( \43733_nG14cfc , \43731_nG14cfa , \43732_nG14cfb , \42599 );
buf \U$37076 ( \43734 , \43733_nG14cfc );
_DC g1aa6e_GF_IsGateDCbyConstraint ( \43735_nG1aa6e , \43734 , \42503 );
buf \U$37077 ( \43736 , \43735_nG1aa6e );
_HMUX g14cfd ( \43737_nG14cfd , RIdbb8480_3857 , \42739 , \43623 );
_HMUX g14cfe ( \43738_nG14cfe , RIdbb8480_3857 , \43737_nG14cfd , \42590 );
_HMUX g14cff ( \43739_nG14cff , RIdbb8480_3857 , \42742 , \43626 );
_HMUX g14d00 ( \43740_nG14d00 , \43738_nG14cfe , \43739_nG14cff , \42599 );
buf \U$37078 ( \43741 , \43740_nG14d00 );
_DC g1aa70_GF_IsGateDCbyConstraint ( \43742_nG1aa70 , \43741 , \42503 );
buf \U$37079 ( \43743 , \43742_nG1aa70 );
_HMUX g14d01 ( \43744_nG14d01 , RIdbb58e8_3858 , \42748 , \43623 );
_HMUX g14d02 ( \43745_nG14d02 , RIdbb58e8_3858 , \43744_nG14d01 , \42590 );
_HMUX g14d03 ( \43746_nG14d03 , RIdbb58e8_3858 , \42751 , \43626 );
_HMUX g14d04 ( \43747_nG14d04 , \43745_nG14d02 , \43746_nG14d03 , \42599 );
buf \U$37080 ( \43748 , \43747_nG14d04 );
_DC g1aa72_GF_IsGateDCbyConstraint ( \43749_nG1aa72 , \43748 , \42503 );
buf \U$37081 ( \43750 , \43749_nG1aa72 );
_HMUX g14d05 ( \43751_nG14d05 , RIdbb2648_3859 , \42757 , \43623 );
_HMUX g14d06 ( \43752_nG14d06 , RIdbb2648_3859 , \43751_nG14d05 , \42590 );
_HMUX g14d07 ( \43753_nG14d07 , RIdbb2648_3859 , \42760 , \43626 );
_HMUX g14d08 ( \43754_nG14d08 , \43752_nG14d06 , \43753_nG14d07 , \42599 );
buf \U$37082 ( \43755 , \43754_nG14d08 );
_DC g1aa74_GF_IsGateDCbyConstraint ( \43756_nG1aa74 , \43755 , \42503 );
buf \U$37083 ( \43757 , \43756_nG1aa74 );
_HMUX g14d09 ( \43758_nG14d09 , RIdbb0758_3860 , \42766 , \43623 );
_HMUX g14d0a ( \43759_nG14d0a , RIdbb0758_3860 , \43758_nG14d09 , \42590 );
_HMUX g14d0b ( \43760_nG14d0b , RIdbb0758_3860 , \42769 , \43626 );
_HMUX g14d0c ( \43761_nG14d0c , \43759_nG14d0a , \43760_nG14d0b , \42599 );
buf \U$37084 ( \43762 , \43761_nG14d0c );
_DC g1aa78_GF_IsGateDCbyConstraint ( \43763_nG1aa78 , \43762 , \42503 );
buf \U$37085 ( \43764 , \43763_nG1aa78 );
_HMUX g14d0d ( \43765_nG14d0d , RIdbad788_3861 , \42775 , \43623 );
_HMUX g14d0e ( \43766_nG14d0e , RIdbad788_3861 , \43765_nG14d0d , \42590 );
_HMUX g14d0f ( \43767_nG14d0f , RIdbad788_3861 , \42778 , \43626 );
_HMUX g14d10 ( \43768_nG14d10 , \43766_nG14d0e , \43767_nG14d0f , \42599 );
buf \U$37086 ( \43769 , \43768_nG14d10 );
_DC g1aa7a_GF_IsGateDCbyConstraint ( \43770_nG1aa7a , \43769 , \42503 );
buf \U$37087 ( \43771 , \43770_nG1aa7a );
_HMUX g14d11 ( \43772_nG14d11 , RIdbaad58_3862 , \42784 , \43623 );
_HMUX g14d12 ( \43773_nG14d12 , RIdbaad58_3862 , \43772_nG14d11 , \42590 );
_HMUX g14d13 ( \43774_nG14d13 , RIdbaad58_3862 , \42787 , \43626 );
_HMUX g14d14 ( \43775_nG14d14 , \43773_nG14d12 , \43774_nG14d13 , \42599 );
buf \U$37088 ( \43776 , \43775_nG14d14 );
_DC g1aa7c_GF_IsGateDCbyConstraint ( \43777_nG1aa7c , \43776 , \42503 );
buf \U$37089 ( \43778 , \43777_nG1aa7c );
_HMUX g14d15 ( \43779_nG14d15 , RIdba7d88_3863 , \42793 , \43623 );
_HMUX g14d16 ( \43780_nG14d16 , RIdba7d88_3863 , \43779_nG14d15 , \42590 );
_HMUX g14d17 ( \43781_nG14d17 , RIdba7d88_3863 , \42796 , \43626 );
_HMUX g14d18 ( \43782_nG14d18 , \43780_nG14d16 , \43781_nG14d17 , \42599 );
buf \U$37090 ( \43783 , \43782_nG14d18 );
_DC g1aa7e_GF_IsGateDCbyConstraint ( \43784_nG1aa7e , \43783 , \42503 );
buf \U$37091 ( \43785 , \43784_nG1aa7e );
_HMUX g14d19 ( \43786_nG14d19 , RIdba55b0_3864 , \42802 , \43623 );
_HMUX g14d1a ( \43787_nG14d1a , RIdba55b0_3864 , \43786_nG14d19 , \42590 );
_HMUX g14d1b ( \43788_nG14d1b , RIdba55b0_3864 , \42805 , \43626 );
_HMUX g14d1c ( \43789_nG14d1c , \43787_nG14d1a , \43788_nG14d1b , \42599 );
buf \U$37092 ( \43790 , \43789_nG14d1c );
_DC g1aa80_GF_IsGateDCbyConstraint ( \43791_nG1aa80 , \43790 , \42503 );
buf \U$37093 ( \43792 , \43791_nG1aa80 );
_HMUX g14d1d ( \43793_nG14d1d , RIdba2ce8_3865 , \42811 , \43623 );
_HMUX g14d1e ( \43794_nG14d1e , RIdba2ce8_3865 , \43793_nG14d1d , \42590 );
_HMUX g14d1f ( \43795_nG14d1f , RIdba2ce8_3865 , \42814 , \43626 );
_HMUX g14d20 ( \43796_nG14d20 , \43794_nG14d1e , \43795_nG14d1f , \42599 );
buf \U$37094 ( \43797 , \43796_nG14d20 );
_DC g1aa82_GF_IsGateDCbyConstraint ( \43798_nG1aa82 , \43797 , \42503 );
buf \U$37095 ( \43799 , \43798_nG1aa82 );
_HMUX g14d21 ( \43800_nG14d21 , RIdb9fe80_3866 , \42820 , \43623 );
_HMUX g14d22 ( \43801_nG14d22 , RIdb9fe80_3866 , \43800_nG14d21 , \42590 );
_HMUX g14d23 ( \43802_nG14d23 , RIdb9fe80_3866 , \42823 , \43626 );
_HMUX g14d24 ( \43803_nG14d24 , \43801_nG14d22 , \43802_nG14d23 , \42599 );
buf \U$37096 ( \43804 , \43803_nG14d24 );
_DC g1aa84_GF_IsGateDCbyConstraint ( \43805_nG1aa84 , \43804 , \42503 );
buf \U$37097 ( \43806 , \43805_nG1aa84 );
_HMUX g14d25 ( \43807_nG14d25 , RIdb9d4c8_3867 , \42829 , \43623 );
_HMUX g14d26 ( \43808_nG14d26 , RIdb9d4c8_3867 , \43807_nG14d25 , \42590 );
_HMUX g14d27 ( \43809_nG14d27 , RIdb9d4c8_3867 , \42832 , \43626 );
_HMUX g14d28 ( \43810_nG14d28 , \43808_nG14d26 , \43809_nG14d27 , \42599 );
buf \U$37098 ( \43811 , \43810_nG14d28 );
_DC g1aa86_GF_IsGateDCbyConstraint ( \43812_nG1aa86 , \43811 , \42503 );
buf \U$37099 ( \43813 , \43812_nG1aa86 );
_HMUX g14d29 ( \43814_nG14d29 , RIdb9acf0_3868 , \42838 , \43623 );
_HMUX g14d2a ( \43815_nG14d2a , RIdb9acf0_3868 , \43814_nG14d29 , \42590 );
_HMUX g14d2b ( \43816_nG14d2b , RIdb9acf0_3868 , \42841 , \43626 );
_HMUX g14d2c ( \43817_nG14d2c , \43815_nG14d2a , \43816_nG14d2b , \42599 );
buf \U$37100 ( \43818 , \43817_nG14d2c );
_DC g1aa88_GF_IsGateDCbyConstraint ( \43819_nG1aa88 , \43818 , \42503 );
buf \U$37101 ( \43820 , \43819_nG1aa88 );
_HMUX g14d2d ( \43821_nG14d2d , RIdb98c20_3869 , \42847 , \43623 );
_HMUX g14d2e ( \43822_nG14d2e , RIdb98c20_3869 , \43821_nG14d2d , \42590 );
_HMUX g14d2f ( \43823_nG14d2f , RIdb98c20_3869 , \42850 , \43626 );
_HMUX g14d30 ( \43824_nG14d30 , \43822_nG14d2e , \43823_nG14d2f , \42599 );
buf \U$37102 ( \43825 , \43824_nG14d30 );
_DC g1aa8a_GF_IsGateDCbyConstraint ( \43826_nG1aa8a , \43825 , \42503 );
buf \U$37103 ( \43827 , \43826_nG1aa8a );
_HMUX g14d31 ( \43828_nG14d31 , RIdb96178_3870 , \42856 , \43623 );
_HMUX g14d32 ( \43829_nG14d32 , RIdb96178_3870 , \43828_nG14d31 , \42590 );
_HMUX g14d33 ( \43830_nG14d33 , RIdb96178_3870 , \42859 , \43626 );
_HMUX g14d34 ( \43831_nG14d34 , \43829_nG14d32 , \43830_nG14d33 , \42599 );
buf \U$37104 ( \43832 , \43831_nG14d34 );
_DC g1aa8e_GF_IsGateDCbyConstraint ( \43833_nG1aa8e , \43832 , \42503 );
buf \U$37105 ( \43834 , \43833_nG1aa8e );
_HMUX g14d35 ( \43835_nG14d35 , RIdb93ce8_3871 , \42865 , \43623 );
_HMUX g14d36 ( \43836_nG14d36 , RIdb93ce8_3871 , \43835_nG14d35 , \42590 );
_HMUX g14d37 ( \43837_nG14d37 , RIdb93ce8_3871 , \42868 , \43626 );
_HMUX g14d38 ( \43838_nG14d38 , \43836_nG14d36 , \43837_nG14d37 , \42599 );
buf \U$37106 ( \43839 , \43838_nG14d38 );
_DC g1aa90_GF_IsGateDCbyConstraint ( \43840_nG1aa90 , \43839 , \42503 );
buf \U$37107 ( \43841 , \43840_nG1aa90 );
_HMUX g14d39 ( \43842_nG14d39 , RIdb916f0_3872 , \42874 , \43623 );
_HMUX g14d3a ( \43843_nG14d3a , RIdb916f0_3872 , \43842_nG14d39 , \42590 );
_HMUX g14d3b ( \43844_nG14d3b , RIdb916f0_3872 , \42877 , \43626 );
_HMUX g14d3c ( \43845_nG14d3c , \43843_nG14d3a , \43844_nG14d3b , \42599 );
buf \U$37108 ( \43846 , \43845_nG14d3c );
_DC g1aa92_GF_IsGateDCbyConstraint ( \43847_nG1aa92 , \43846 , \42503 );
buf \U$37109 ( \43848 , \43847_nG1aa92 );
_HMUX g14d3d ( \43849_nG14d3d , RIdb8e2e8_3873 , \42883 , \43623 );
_HMUX g14d3e ( \43850_nG14d3e , RIdb8e2e8_3873 , \43849_nG14d3d , \42590 );
_HMUX g14d3f ( \43851_nG14d3f , RIdb8e2e8_3873 , \42886 , \43626 );
_HMUX g14d40 ( \43852_nG14d40 , \43850_nG14d3e , \43851_nG14d3f , \42599 );
buf \U$37110 ( \43853 , \43852_nG14d40 );
_DC g1aa94_GF_IsGateDCbyConstraint ( \43854_nG1aa94 , \43853 , \42503 );
buf \U$37111 ( \43855 , \43854_nG1aa94 );
_HMUX g14d41 ( \43856_nG14d41 , RIdb8b840_3874 , \42892 , \43623 );
_HMUX g14d42 ( \43857_nG14d42 , RIdb8b840_3874 , \43856_nG14d41 , \42590 );
_HMUX g14d43 ( \43858_nG14d43 , RIdb8b840_3874 , \42895 , \43626 );
_HMUX g14d44 ( \43859_nG14d44 , \43857_nG14d42 , \43858_nG14d43 , \42599 );
buf \U$37112 ( \43860 , \43859_nG14d44 );
_DC g1aa96_GF_IsGateDCbyConstraint ( \43861_nG1aa96 , \43860 , \42503 );
buf \U$37113 ( \43862 , \43861_nG1aa96 );
_HMUX g14d45 ( \43863_nG14d45 , RIdb890e0_3875 , \42901 , \43623 );
_HMUX g14d46 ( \43864_nG14d46 , RIdb890e0_3875 , \43863_nG14d45 , \42590 );
_HMUX g14d47 ( \43865_nG14d47 , RIdb890e0_3875 , \42904 , \43626 );
_HMUX g14d48 ( \43866_nG14d48 , \43864_nG14d46 , \43865_nG14d47 , \42599 );
buf \U$37114 ( \43867 , \43866_nG14d48 );
_DC g1aa98_GF_IsGateDCbyConstraint ( \43868_nG1aa98 , \43867 , \42503 );
buf \U$37115 ( \43869 , \43868_nG1aa98 );
_HMUX g14d49 ( \43870_nG14d49 , RIdb86cc8_3876 , \42910 , \43623 );
_HMUX g14d4a ( \43871_nG14d4a , RIdb86cc8_3876 , \43870_nG14d49 , \42590 );
_HMUX g14d4b ( \43872_nG14d4b , RIdb86cc8_3876 , \42913 , \43626 );
_HMUX g14d4c ( \43873_nG14d4c , \43871_nG14d4a , \43872_nG14d4b , \42599 );
buf \U$37116 ( \43874 , \43873_nG14d4c );
_DC g1aa9a_GF_IsGateDCbyConstraint ( \43875_nG1aa9a , \43874 , \42503 );
buf \U$37117 ( \43876 , \43875_nG1aa9a );
_HMUX g14d4d ( \43877_nG14d4d , RIdb84ec8_3877 , \42919 , \43623 );
_HMUX g14d4e ( \43878_nG14d4e , RIdb84ec8_3877 , \43877_nG14d4d , \42590 );
_HMUX g14d4f ( \43879_nG14d4f , RIdb84ec8_3877 , \42922 , \43626 );
_HMUX g14d50 ( \43880_nG14d50 , \43878_nG14d4e , \43879_nG14d4f , \42599 );
buf \U$37118 ( \43881 , \43880_nG14d50 );
_DC g1aa9c_GF_IsGateDCbyConstraint ( \43882_nG1aa9c , \43881 , \42503 );
buf \U$37119 ( \43883 , \43882_nG1aa9c );
_HMUX g14d51 ( \43884_nG14d51 , RIdb83410_3878 , \42928 , \43623 );
_HMUX g14d52 ( \43885_nG14d52 , RIdb83410_3878 , \43884_nG14d51 , \42590 );
_HMUX g14d53 ( \43886_nG14d53 , RIdb83410_3878 , \42931 , \43626 );
_HMUX g14d54 ( \43887_nG14d54 , \43885_nG14d52 , \43886_nG14d53 , \42599 );
buf \U$37120 ( \43888 , \43887_nG14d54 );
_DC g1aa9e_GF_IsGateDCbyConstraint ( \43889_nG1aa9e , \43888 , \42503 );
buf \U$37121 ( \43890 , \43889_nG1aa9e );
_HMUX g14d55 ( \43891_nG14d55 , RIdb81700_3879 , \42937 , \43623 );
_HMUX g14d56 ( \43892_nG14d56 , RIdb81700_3879 , \43891_nG14d55 , \42590 );
_HMUX g14d57 ( \43893_nG14d57 , RIdb81700_3879 , \42940 , \43626 );
_HMUX g14d58 ( \43894_nG14d58 , \43892_nG14d56 , \43893_nG14d57 , \42599 );
buf \U$37122 ( \43895 , \43894_nG14d58 );
_DC g1aaa0_GF_IsGateDCbyConstraint ( \43896_nG1aaa0 , \43895 , \42503 );
buf \U$37123 ( \43897 , \43896_nG1aaa0 );
_HMUX g14d59 ( \43898_nG14d59 , RIdb7fa68_3880 , \42946 , \43623 );
_HMUX g14d5a ( \43899_nG14d5a , RIdb7fa68_3880 , \43898_nG14d59 , \42590 );
_HMUX g14d5b ( \43900_nG14d5b , RIdb7fa68_3880 , \42949 , \43626 );
_HMUX g14d5c ( \43901_nG14d5c , \43899_nG14d5a , \43900_nG14d5b , \42599 );
buf \U$37124 ( \43902 , \43901_nG14d5c );
_DC g1aaa4_GF_IsGateDCbyConstraint ( \43903_nG1aaa4 , \43902 , \42503 );
buf \U$37125 ( \43904 , \43903_nG1aaa4 );
_HMUX g14d5d ( \43905_nG14d5d , RIdb7db78_3881 , \42955 , \43623 );
_HMUX g14d5e ( \43906_nG14d5e , RIdb7db78_3881 , \43905_nG14d5d , \42590 );
_HMUX g14d5f ( \43907_nG14d5f , RIdb7db78_3881 , \42958 , \43626 );
_HMUX g14d60 ( \43908_nG14d60 , \43906_nG14d5e , \43907_nG14d5f , \42599 );
buf \U$37126 ( \43909 , \43908_nG14d60 );
_DC g1aaa6_GF_IsGateDCbyConstraint ( \43910_nG1aaa6 , \43909 , \42503 );
buf \U$37127 ( \43911 , \43910_nG1aaa6 );
_HMUX g14d61 ( \43912_nG14d61 , RIdb7bb98_3882 , \42964 , \43623 );
_HMUX g14d62 ( \43913_nG14d62 , RIdb7bb98_3882 , \43912_nG14d61 , \42590 );
_HMUX g14d63 ( \43914_nG14d63 , RIdb7bb98_3882 , \42967 , \43626 );
_HMUX g14d64 ( \43915_nG14d64 , \43913_nG14d62 , \43914_nG14d63 , \42599 );
buf \U$37128 ( \43916 , \43915_nG14d64 );
_DC g1aaa8_GF_IsGateDCbyConstraint ( \43917_nG1aaa8 , \43916 , \42503 );
buf \U$37129 ( \43918 , \43917_nG1aaa8 );
_HMUX g14d65 ( \43919_nG14d65 , RIdb79e10_3883 , \42973 , \43623 );
_HMUX g14d66 ( \43920_nG14d66 , RIdb79e10_3883 , \43919_nG14d65 , \42590 );
_HMUX g14d67 ( \43921_nG14d67 , RIdb79e10_3883 , \42976 , \43626 );
_HMUX g14d68 ( \43922_nG14d68 , \43920_nG14d66 , \43921_nG14d67 , \42599 );
buf \U$37130 ( \43923 , \43922_nG14d68 );
_DC g1aaaa_GF_IsGateDCbyConstraint ( \43924_nG1aaaa , \43923 , \42503 );
buf \U$37131 ( \43925 , \43924_nG1aaaa );
_HMUX g14d69 ( \43926_nG14d69 , RIdb78268_3884 , \42982 , \43623 );
_HMUX g14d6a ( \43927_nG14d6a , RIdb78268_3884 , \43926_nG14d69 , \42590 );
_HMUX g14d6b ( \43928_nG14d6b , RIdb78268_3884 , \42985 , \43626 );
_HMUX g14d6c ( \43929_nG14d6c , \43927_nG14d6a , \43928_nG14d6b , \42599 );
buf \U$37132 ( \43930 , \43929_nG14d6c );
_DC g1aaac_GF_IsGateDCbyConstraint ( \43931_nG1aaac , \43930 , \42503 );
buf \U$37133 ( \43932 , \43931_nG1aaac );
_HMUX g14d6d ( \43933_nG14d6d , RIdb76828_3885 , \42991 , \43623 );
_HMUX g14d6e ( \43934_nG14d6e , RIdb76828_3885 , \43933_nG14d6d , \42590 );
_HMUX g14d6f ( \43935_nG14d6f , RIdb76828_3885 , \42994 , \43626 );
_HMUX g14d70 ( \43936_nG14d70 , \43934_nG14d6e , \43935_nG14d6f , \42599 );
buf \U$37134 ( \43937 , \43936_nG14d70 );
_DC g1aaae_GF_IsGateDCbyConstraint ( \43938_nG1aaae , \43937 , \42503 );
buf \U$37135 ( \43939 , \43938_nG1aaae );
_HMUX g14d71 ( \43940_nG14d71 , RIdb746e0_3886 , \43000 , \43623 );
_HMUX g14d72 ( \43941_nG14d72 , RIdb746e0_3886 , \43940_nG14d71 , \42590 );
_HMUX g14d73 ( \43942_nG14d73 , RIdb746e0_3886 , \43003 , \43626 );
_HMUX g14d74 ( \43943_nG14d74 , \43941_nG14d72 , \43942_nG14d73 , \42599 );
buf \U$37136 ( \43944 , \43943_nG14d74 );
_DC g1aab0_GF_IsGateDCbyConstraint ( \43945_nG1aab0 , \43944 , \42503 );
buf \U$37137 ( \43946 , \43945_nG1aab0 );
_HMUX g14d75 ( \43947_nG14d75 , RIdda9490_3887 , \43009 , \43623 );
_HMUX g14d76 ( \43948_nG14d76 , RIdda9490_3887 , \43947_nG14d75 , \42590 );
_HMUX g14d77 ( \43949_nG14d77 , RIdda9490_3887 , \43012 , \43626 );
_HMUX g14d78 ( \43950_nG14d78 , \43948_nG14d76 , \43949_nG14d77 , \42599 );
buf \U$37138 ( \43951 , \43950_nG14d78 );
_DC g1aab2_GF_IsGateDCbyConstraint ( \43952_nG1aab2 , \43951 , \42503 );
buf \U$37139 ( \43953 , \43952_nG1aab2 );
_HMUX g14d79 ( \43954_nG14d79 , RIdda9c88_3888 , \43018 , \43623 );
_HMUX g14d7a ( \43955_nG14d7a , RIdda9c88_3888 , \43954_nG14d79 , \42590 );
_HMUX g14d7b ( \43956_nG14d7b , RIdda9c88_3888 , \43021 , \43626 );
_HMUX g14d7c ( \43957_nG14d7c , \43955_nG14d7a , \43956_nG14d7b , \42599 );
buf \U$37140 ( \43958 , \43957_nG14d7c );
_DC g1aab4_GF_IsGateDCbyConstraint ( \43959_nG1aab4 , \43958 , \42503 );
buf \U$37141 ( \43960 , \43959_nG1aab4 );
_HMUX g14d7d ( \43961_nG14d7d , RIddaa480_3889 , \43027 , \43623 );
_HMUX g14d7e ( \43962_nG14d7e , RIddaa480_3889 , \43961_nG14d7d , \42590 );
_HMUX g14d7f ( \43963_nG14d7f , RIddaa480_3889 , \43030 , \43626 );
_HMUX g14d80 ( \43964_nG14d80 , \43962_nG14d7e , \43963_nG14d7f , \42599 );
buf \U$37142 ( \43965 , \43964_nG14d80 );
_DC g1aab6_GF_IsGateDCbyConstraint ( \43966_nG1aab6 , \43965 , \42503 );
buf \U$37143 ( \43967 , \43966_nG1aab6 );
_HMUX g14d81 ( \43968_nG14d81 , RIddaac78_3890 , \43036 , \43623 );
_HMUX g14d82 ( \43969_nG14d82 , RIddaac78_3890 , \43968_nG14d81 , \42590 );
_HMUX g14d83 ( \43970_nG14d83 , RIddaac78_3890 , \43039 , \43626 );
_HMUX g14d84 ( \43971_nG14d84 , \43969_nG14d82 , \43970_nG14d83 , \42599 );
buf \U$37144 ( \43972 , \43971_nG14d84 );
_DC g1aaba_GF_IsGateDCbyConstraint ( \43973_nG1aaba , \43972 , \42503 );
buf \U$37145 ( \43974 , \43973_nG1aaba );
_HMUX g14d85 ( \43975_nG14d85 , RIddab470_3891 , \43045 , \43623 );
_HMUX g14d86 ( \43976_nG14d86 , RIddab470_3891 , \43975_nG14d85 , \42590 );
_HMUX g14d87 ( \43977_nG14d87 , RIddab470_3891 , \43048 , \43626 );
_HMUX g14d88 ( \43978_nG14d88 , \43976_nG14d86 , \43977_nG14d87 , \42599 );
buf \U$37146 ( \43979 , \43978_nG14d88 );
_DC g1aabc_GF_IsGateDCbyConstraint ( \43980_nG1aabc , \43979 , \42503 );
buf \U$37147 ( \43981 , \43980_nG1aabc );
_HMUX g14d89 ( \43982_nG14d89 , RIddabc68_3892 , \43054 , \43623 );
_HMUX g14d8a ( \43983_nG14d8a , RIddabc68_3892 , \43982_nG14d89 , \42590 );
_HMUX g14d8b ( \43984_nG14d8b , RIddabc68_3892 , \43057 , \43626 );
_HMUX g14d8c ( \43985_nG14d8c , \43983_nG14d8a , \43984_nG14d8b , \42599 );
buf \U$37148 ( \43986 , \43985_nG14d8c );
_DC g1aabe_GF_IsGateDCbyConstraint ( \43987_nG1aabe , \43986 , \42503 );
buf \U$37149 ( \43988 , \43987_nG1aabe );
_HMUX g14d8d ( \43989_nG14d8d , RIddac460_3893 , \43063 , \43623 );
_HMUX g14d8e ( \43990_nG14d8e , RIddac460_3893 , \43989_nG14d8d , \42590 );
_HMUX g14d8f ( \43991_nG14d8f , RIddac460_3893 , \43066 , \43626 );
_HMUX g14d90 ( \43992_nG14d90 , \43990_nG14d8e , \43991_nG14d8f , \42599 );
buf \U$37150 ( \43993 , \43992_nG14d90 );
_DC g1aac0_GF_IsGateDCbyConstraint ( \43994_nG1aac0 , \43993 , \42503 );
buf \U$37151 ( \43995 , \43994_nG1aac0 );
_HMUX g14d91 ( \43996_nG14d91 , RIddacc58_3894 , \43072 , \43623 );
_HMUX g14d92 ( \43997_nG14d92 , RIddacc58_3894 , \43996_nG14d91 , \42590 );
_HMUX g14d93 ( \43998_nG14d93 , RIddacc58_3894 , \43075 , \43626 );
_HMUX g14d94 ( \43999_nG14d94 , \43997_nG14d92 , \43998_nG14d93 , \42599 );
buf \U$37152 ( \44000 , \43999_nG14d94 );
_DC g1aac2_GF_IsGateDCbyConstraint ( \44001_nG1aac2 , \44000 , \42503 );
buf \U$37153 ( \44002 , \44001_nG1aac2 );
_HMUX g14d95 ( \44003_nG14d95 , RIddad450_3895 , \43081 , \43623 );
_HMUX g14d96 ( \44004_nG14d96 , RIddad450_3895 , \44003_nG14d95 , \42590 );
_HMUX g14d97 ( \44005_nG14d97 , RIddad450_3895 , \43084 , \43626 );
_HMUX g14d98 ( \44006_nG14d98 , \44004_nG14d96 , \44005_nG14d97 , \42599 );
buf \U$37154 ( \44007 , \44006_nG14d98 );
_DC g1aac4_GF_IsGateDCbyConstraint ( \44008_nG1aac4 , \44007 , \42503 );
buf \U$37155 ( \44009 , \44008_nG1aac4 );
_HMUX g14d99 ( \44010_nG14d99 , RIddadc48_3896 , \43090 , \43623 );
_HMUX g14d9a ( \44011_nG14d9a , RIddadc48_3896 , \44010_nG14d99 , \42590 );
_HMUX g14d9b ( \44012_nG14d9b , RIddadc48_3896 , \43093 , \43626 );
_HMUX g14d9c ( \44013_nG14d9c , \44011_nG14d9a , \44012_nG14d9b , \42599 );
buf \U$37156 ( \44014 , \44013_nG14d9c );
_DC g1aac6_GF_IsGateDCbyConstraint ( \44015_nG1aac6 , \44014 , \42503 );
buf \U$37157 ( \44016 , \44015_nG1aac6 );
_HMUX g14d9d ( \44017_nG14d9d , RIddae440_3897 , \43099 , \43623 );
_HMUX g14d9e ( \44018_nG14d9e , RIddae440_3897 , \44017_nG14d9d , \42590 );
_HMUX g14d9f ( \44019_nG14d9f , RIddae440_3897 , \43102 , \43626 );
_HMUX g14da0 ( \44020_nG14da0 , \44018_nG14d9e , \44019_nG14d9f , \42599 );
buf \U$37158 ( \44021 , \44020_nG14da0 );
_DC g1aac8_GF_IsGateDCbyConstraint ( \44022_nG1aac8 , \44021 , \42503 );
buf \U$37159 ( \44023 , \44022_nG1aac8 );
_HMUX g14da1 ( \44024_nG14da1 , RIddaec38_3898 , \43108 , \43623 );
_HMUX g14da2 ( \44025_nG14da2 , RIddaec38_3898 , \44024_nG14da1 , \42590 );
_HMUX g14da3 ( \44026_nG14da3 , RIddaec38_3898 , \43111 , \43626 );
_HMUX g14da4 ( \44027_nG14da4 , \44025_nG14da2 , \44026_nG14da3 , \42599 );
buf \U$37160 ( \44028 , \44027_nG14da4 );
_DC g1aaca_GF_IsGateDCbyConstraint ( \44029_nG1aaca , \44028 , \42503 );
buf \U$37161 ( \44030 , \44029_nG1aaca );
_HMUX g14da5 ( \44031_nG14da5 , RIddaf430_3899 , \43117 , \43623 );
_HMUX g14da6 ( \44032_nG14da6 , RIddaf430_3899 , \44031_nG14da5 , \42590 );
_HMUX g14da7 ( \44033_nG14da7 , RIddaf430_3899 , \43120 , \43626 );
_HMUX g14da8 ( \44034_nG14da8 , \44032_nG14da6 , \44033_nG14da7 , \42599 );
buf \U$37162 ( \44035 , \44034_nG14da8 );
_DC g1aacc_GF_IsGateDCbyConstraint ( \44036_nG1aacc , \44035 , \42503 );
buf \U$37163 ( \44037 , \44036_nG1aacc );
_HMUX g14da9 ( \44038_nG14da9 , RIddafc28_3900 , \43126 , \43623 );
_HMUX g14daa ( \44039_nG14daa , RIddafc28_3900 , \44038_nG14da9 , \42590 );
_HMUX g14dab ( \44040_nG14dab , RIddafc28_3900 , \43129 , \43626 );
_HMUX g14dac ( \44041_nG14dac , \44039_nG14daa , \44040_nG14dab , \42599 );
buf \U$37164 ( \44042 , \44041_nG14dac );
_DC g1aad0_GF_IsGateDCbyConstraint ( \44043_nG1aad0 , \44042 , \42503 );
buf \U$37165 ( \44044 , \44043_nG1aad0 );
_HMUX g14dad ( \44045_nG14dad , RIddb0420_3901 , \43135 , \43623 );
_HMUX g14dae ( \44046_nG14dae , RIddb0420_3901 , \44045_nG14dad , \42590 );
_HMUX g14daf ( \44047_nG14daf , RIddb0420_3901 , \43138 , \43626 );
_HMUX g14db0 ( \44048_nG14db0 , \44046_nG14dae , \44047_nG14daf , \42599 );
buf \U$37166 ( \44049 , \44048_nG14db0 );
_DC g1aad2_GF_IsGateDCbyConstraint ( \44050_nG1aad2 , \44049 , \42503 );
buf \U$37167 ( \44051 , \44050_nG1aad2 );
_HMUX g14db1 ( \44052_nG14db1 , RIddb0c18_3902 , \43144 , \43623 );
_HMUX g14db2 ( \44053_nG14db2 , RIddb0c18_3902 , \44052_nG14db1 , \42590 );
_HMUX g14db3 ( \44054_nG14db3 , RIddb0c18_3902 , \43147 , \43626 );
_HMUX g14db4 ( \44055_nG14db4 , \44053_nG14db2 , \44054_nG14db3 , \42599 );
buf \U$37168 ( \44056 , \44055_nG14db4 );
_DC g1aad4_GF_IsGateDCbyConstraint ( \44057_nG1aad4 , \44056 , \42503 );
buf \U$37169 ( \44058 , \44057_nG1aad4 );
_HMUX g14db5 ( \44059_nG14db5 , RIddb1410_3903 , \43153 , \43623 );
_HMUX g14db6 ( \44060_nG14db6 , RIddb1410_3903 , \44059_nG14db5 , \42590 );
_HMUX g14db7 ( \44061_nG14db7 , RIddb1410_3903 , \43156 , \43626 );
_HMUX g14db8 ( \44062_nG14db8 , \44060_nG14db6 , \44061_nG14db7 , \42599 );
buf \U$37170 ( \44063 , \44062_nG14db8 );
_DC g1aad6_GF_IsGateDCbyConstraint ( \44064_nG1aad6 , \44063 , \42503 );
buf \U$37171 ( \44065 , \44064_nG1aad6 );
_HMUX g14db9 ( \44066_nG14db9 , RIddb1c08_3904 , \43162 , \43623 );
_HMUX g14dba ( \44067_nG14dba , RIddb1c08_3904 , \44066_nG14db9 , \42590 );
_HMUX g14dbb ( \44068_nG14dbb , RIddb1c08_3904 , \43165 , \43626 );
_HMUX g14dbc ( \44069_nG14dbc , \44067_nG14dba , \44068_nG14dbb , \42599 );
buf \U$37172 ( \44070 , \44069_nG14dbc );
_DC g1aad8_GF_IsGateDCbyConstraint ( \44071_nG1aad8 , \44070 , \42503 );
buf \U$37173 ( \44072 , \44071_nG1aad8 );
and \U$37174 ( \44073 , \42579 , \42580 );
_HMUX g14b39 ( \44074_nG14b39 , RIddb2400_3905 , \42578 , \44073 );
_HMUX g14b3a ( \44075_nG14b3a , RIddb2400_3905 , \44074_nG14b39 , \42590 );
and \U$37175 ( \44076 , \42593 , \42594 );
_HMUX g14b3f ( \44077_nG14b3f , RIddb2400_3905 , \42592 , \44076 );
_HMUX g14b40 ( \44078_nG14b40 , \44075_nG14b3a , \44077_nG14b3f , \42599 );
buf \U$37176 ( \44079 , \44078_nG14b40 );
_DC g1a9e0_GF_IsGateDCbyConstraint ( \44080_nG1a9e0 , \44079 , \42503 );
buf \U$37177 ( \44081 , \44080_nG1a9e0 );
_HMUX g14b42 ( \44082_nG14b42 , RIddb2bf8_3906 , \42604 , \44073 );
_HMUX g14b43 ( \44083_nG14b43 , RIddb2bf8_3906 , \44082_nG14b42 , \42590 );
_HMUX g14b45 ( \44084_nG14b45 , RIddb2bf8_3906 , \42607 , \44076 );
_HMUX g14b46 ( \44085_nG14b46 , \44083_nG14b43 , \44084_nG14b45 , \42599 );
buf \U$37178 ( \44086 , \44085_nG14b46 );
_DC g1a9f6_GF_IsGateDCbyConstraint ( \44087_nG1a9f6 , \44086 , \42503 );
buf \U$37179 ( \44088 , \44087_nG1a9f6 );
_HMUX g14b48 ( \44089_nG14b48 , RIddb33f0_3907 , \42613 , \44073 );
_HMUX g14b49 ( \44090_nG14b49 , RIddb33f0_3907 , \44089_nG14b48 , \42590 );
_HMUX g14b4b ( \44091_nG14b4b , RIddb33f0_3907 , \42616 , \44076 );
_HMUX g14b4c ( \44092_nG14b4c , \44090_nG14b49 , \44091_nG14b4b , \42599 );
buf \U$37180 ( \44093 , \44092_nG14b4c );
_DC g1aa0c_GF_IsGateDCbyConstraint ( \44094_nG1aa0c , \44093 , \42503 );
buf \U$37181 ( \44095 , \44094_nG1aa0c );
_HMUX g14b4e ( \44096_nG14b4e , RIddb3be8_3908 , \42622 , \44073 );
_HMUX g14b4f ( \44097_nG14b4f , RIddb3be8_3908 , \44096_nG14b4e , \42590 );
_HMUX g14b51 ( \44098_nG14b51 , RIddb3be8_3908 , \42625 , \44076 );
_HMUX g14b52 ( \44099_nG14b52 , \44097_nG14b4f , \44098_nG14b51 , \42599 );
buf \U$37182 ( \44100 , \44099_nG14b52 );
_DC g1aa22_GF_IsGateDCbyConstraint ( \44101_nG1aa22 , \44100 , \42503 );
buf \U$37183 ( \44102 , \44101_nG1aa22 );
_HMUX g14b54 ( \44103_nG14b54 , RIddb43e0_3909 , \42631 , \44073 );
_HMUX g14b55 ( \44104_nG14b55 , RIddb43e0_3909 , \44103_nG14b54 , \42590 );
_HMUX g14b57 ( \44105_nG14b57 , RIddb43e0_3909 , \42634 , \44076 );
_HMUX g14b58 ( \44106_nG14b58 , \44104_nG14b55 , \44105_nG14b57 , \42599 );
buf \U$37184 ( \44107 , \44106_nG14b58 );
_DC g1aa38_GF_IsGateDCbyConstraint ( \44108_nG1aa38 , \44107 , \42503 );
buf \U$37185 ( \44109 , \44108_nG1aa38 );
_HMUX g14b5a ( \44110_nG14b5a , RIddb4bd8_3910 , \42640 , \44073 );
_HMUX g14b5b ( \44111_nG14b5b , RIddb4bd8_3910 , \44110_nG14b5a , \42590 );
_HMUX g14b5d ( \44112_nG14b5d , RIddb4bd8_3910 , \42643 , \44076 );
_HMUX g14b5e ( \44113_nG14b5e , \44111_nG14b5b , \44112_nG14b5d , \42599 );
buf \U$37186 ( \44114 , \44113_nG14b5e );
_DC g1aa4e_GF_IsGateDCbyConstraint ( \44115_nG1aa4e , \44114 , \42503 );
buf \U$37187 ( \44116 , \44115_nG1aa4e );
_HMUX g14b60 ( \44117_nG14b60 , RIddb53d0_3911 , \42649 , \44073 );
_HMUX g14b61 ( \44118_nG14b61 , RIddb53d0_3911 , \44117_nG14b60 , \42590 );
_HMUX g14b63 ( \44119_nG14b63 , RIddb53d0_3911 , \42652 , \44076 );
_HMUX g14b64 ( \44120_nG14b64 , \44118_nG14b61 , \44119_nG14b63 , \42599 );
buf \U$37188 ( \44121 , \44120_nG14b64 );
_DC g1aa5a_GF_IsGateDCbyConstraint ( \44122_nG1aa5a , \44121 , \42503 );
buf \U$37189 ( \44123 , \44122_nG1aa5a );
_HMUX g14b66 ( \44124_nG14b66 , RIddb5bc8_3912 , \42658 , \44073 );
_HMUX g14b67 ( \44125_nG14b67 , RIddb5bc8_3912 , \44124_nG14b66 , \42590 );
_HMUX g14b69 ( \44126_nG14b69 , RIddb5bc8_3912 , \42661 , \44076 );
_HMUX g14b6a ( \44127_nG14b6a , \44125_nG14b67 , \44126_nG14b69 , \42599 );
buf \U$37190 ( \44128 , \44127_nG14b6a );
_DC g1aa5c_GF_IsGateDCbyConstraint ( \44129_nG1aa5c , \44128 , \42503 );
buf \U$37191 ( \44130 , \44129_nG1aa5c );
_HMUX g14b6c ( \44131_nG14b6c , RIddb63c0_3913 , \42667 , \44073 );
_HMUX g14b6d ( \44132_nG14b6d , RIddb63c0_3913 , \44131_nG14b6c , \42590 );
_HMUX g14b6f ( \44133_nG14b6f , RIddb63c0_3913 , \42670 , \44076 );
_HMUX g14b70 ( \44134_nG14b70 , \44132_nG14b6d , \44133_nG14b6f , \42599 );
buf \U$37192 ( \44135 , \44134_nG14b70 );
_DC g1aa5e_GF_IsGateDCbyConstraint ( \44136_nG1aa5e , \44135 , \42503 );
buf \U$37193 ( \44137 , \44136_nG1aa5e );
_HMUX g14b72 ( \44138_nG14b72 , RIddb6bb8_3914 , \42676 , \44073 );
_HMUX g14b73 ( \44139_nG14b73 , RIddb6bb8_3914 , \44138_nG14b72 , \42590 );
_HMUX g14b75 ( \44140_nG14b75 , RIddb6bb8_3914 , \42679 , \44076 );
_HMUX g14b76 ( \44141_nG14b76 , \44139_nG14b73 , \44140_nG14b75 , \42599 );
buf \U$37194 ( \44142 , \44141_nG14b76 );
_DC g1a9e2_GF_IsGateDCbyConstraint ( \44143_nG1a9e2 , \44142 , \42503 );
buf \U$37195 ( \44144 , \44143_nG1a9e2 );
_HMUX g14b78 ( \44145_nG14b78 , RIddb73b0_3915 , \42685 , \44073 );
_HMUX g14b79 ( \44146_nG14b79 , RIddb73b0_3915 , \44145_nG14b78 , \42590 );
_HMUX g14b7b ( \44147_nG14b7b , RIddb73b0_3915 , \42688 , \44076 );
_HMUX g14b7c ( \44148_nG14b7c , \44146_nG14b79 , \44147_nG14b7b , \42599 );
buf \U$37196 ( \44149 , \44148_nG14b7c );
_DC g1a9e4_GF_IsGateDCbyConstraint ( \44150_nG1a9e4 , \44149 , \42503 );
buf \U$37197 ( \44151 , \44150_nG1a9e4 );
_HMUX g14b7e ( \44152_nG14b7e , RIddb7ba8_3916 , \42694 , \44073 );
_HMUX g14b7f ( \44153_nG14b7f , RIddb7ba8_3916 , \44152_nG14b7e , \42590 );
_HMUX g14b81 ( \44154_nG14b81 , RIddb7ba8_3916 , \42697 , \44076 );
_HMUX g14b82 ( \44155_nG14b82 , \44153_nG14b7f , \44154_nG14b81 , \42599 );
buf \U$37198 ( \44156 , \44155_nG14b82 );
_DC g1a9e6_GF_IsGateDCbyConstraint ( \44157_nG1a9e6 , \44156 , \42503 );
buf \U$37199 ( \44158 , \44157_nG1a9e6 );
_HMUX g14b84 ( \44159_nG14b84 , RIddb83a0_3917 , \42703 , \44073 );
_HMUX g14b85 ( \44160_nG14b85 , RIddb83a0_3917 , \44159_nG14b84 , \42590 );
_HMUX g14b87 ( \44161_nG14b87 , RIddb83a0_3917 , \42706 , \44076 );
_HMUX g14b88 ( \44162_nG14b88 , \44160_nG14b85 , \44161_nG14b87 , \42599 );
buf \U$37200 ( \44163 , \44162_nG14b88 );
_DC g1a9e8_GF_IsGateDCbyConstraint ( \44164_nG1a9e8 , \44163 , \42503 );
buf \U$37201 ( \44165 , \44164_nG1a9e8 );
_HMUX g14b8a ( \44166_nG14b8a , RIddb8b98_3918 , \42712 , \44073 );
_HMUX g14b8b ( \44167_nG14b8b , RIddb8b98_3918 , \44166_nG14b8a , \42590 );
_HMUX g14b8d ( \44168_nG14b8d , RIddb8b98_3918 , \42715 , \44076 );
_HMUX g14b8e ( \44169_nG14b8e , \44167_nG14b8b , \44168_nG14b8d , \42599 );
buf \U$37202 ( \44170 , \44169_nG14b8e );
_DC g1a9ea_GF_IsGateDCbyConstraint ( \44171_nG1a9ea , \44170 , \42503 );
buf \U$37203 ( \44172 , \44171_nG1a9ea );
_HMUX g14b90 ( \44173_nG14b90 , RIddb9390_3919 , \42721 , \44073 );
_HMUX g14b91 ( \44174_nG14b91 , RIddb9390_3919 , \44173_nG14b90 , \42590 );
_HMUX g14b93 ( \44175_nG14b93 , RIddb9390_3919 , \42724 , \44076 );
_HMUX g14b94 ( \44176_nG14b94 , \44174_nG14b91 , \44175_nG14b93 , \42599 );
buf \U$37204 ( \44177 , \44176_nG14b94 );
_DC g1a9ec_GF_IsGateDCbyConstraint ( \44178_nG1a9ec , \44177 , \42503 );
buf \U$37205 ( \44179 , \44178_nG1a9ec );
_HMUX g14b96 ( \44180_nG14b96 , RIddb9b88_3920 , \42730 , \44073 );
_HMUX g14b97 ( \44181_nG14b97 , RIddb9b88_3920 , \44180_nG14b96 , \42590 );
_HMUX g14b99 ( \44182_nG14b99 , RIddb9b88_3920 , \42733 , \44076 );
_HMUX g14b9a ( \44183_nG14b9a , \44181_nG14b97 , \44182_nG14b99 , \42599 );
buf \U$37206 ( \44184 , \44183_nG14b9a );
_DC g1a9ee_GF_IsGateDCbyConstraint ( \44185_nG1a9ee , \44184 , \42503 );
buf \U$37207 ( \44186 , \44185_nG1a9ee );
_HMUX g14b9c ( \44187_nG14b9c , RIddba380_3921 , \42739 , \44073 );
_HMUX g14b9d ( \44188_nG14b9d , RIddba380_3921 , \44187_nG14b9c , \42590 );
_HMUX g14b9f ( \44189_nG14b9f , RIddba380_3921 , \42742 , \44076 );
_HMUX g14ba0 ( \44190_nG14ba0 , \44188_nG14b9d , \44189_nG14b9f , \42599 );
buf \U$37208 ( \44191 , \44190_nG14ba0 );
_DC g1a9f0_GF_IsGateDCbyConstraint ( \44192_nG1a9f0 , \44191 , \42503 );
buf \U$37209 ( \44193 , \44192_nG1a9f0 );
_HMUX g14ba2 ( \44194_nG14ba2 , RIddbab78_3922 , \42748 , \44073 );
_HMUX g14ba3 ( \44195_nG14ba3 , RIddbab78_3922 , \44194_nG14ba2 , \42590 );
_HMUX g14ba5 ( \44196_nG14ba5 , RIddbab78_3922 , \42751 , \44076 );
_HMUX g14ba6 ( \44197_nG14ba6 , \44195_nG14ba3 , \44196_nG14ba5 , \42599 );
buf \U$37210 ( \44198 , \44197_nG14ba6 );
_DC g1a9f2_GF_IsGateDCbyConstraint ( \44199_nG1a9f2 , \44198 , \42503 );
buf \U$37211 ( \44200 , \44199_nG1a9f2 );
_HMUX g14ba8 ( \44201_nG14ba8 , RIddbb370_3923 , \42757 , \44073 );
_HMUX g14ba9 ( \44202_nG14ba9 , RIddbb370_3923 , \44201_nG14ba8 , \42590 );
_HMUX g14bab ( \44203_nG14bab , RIddbb370_3923 , \42760 , \44076 );
_HMUX g14bac ( \44204_nG14bac , \44202_nG14ba9 , \44203_nG14bab , \42599 );
buf \U$37212 ( \44205 , \44204_nG14bac );
_DC g1a9f4_GF_IsGateDCbyConstraint ( \44206_nG1a9f4 , \44205 , \42503 );
buf \U$37213 ( \44207 , \44206_nG1a9f4 );
_HMUX g14bae ( \44208_nG14bae , RIddbbb68_3924 , \42766 , \44073 );
_HMUX g14baf ( \44209_nG14baf , RIddbbb68_3924 , \44208_nG14bae , \42590 );
_HMUX g14bb1 ( \44210_nG14bb1 , RIddbbb68_3924 , \42769 , \44076 );
_HMUX g14bb2 ( \44211_nG14bb2 , \44209_nG14baf , \44210_nG14bb1 , \42599 );
buf \U$37214 ( \44212 , \44211_nG14bb2 );
_DC g1a9f8_GF_IsGateDCbyConstraint ( \44213_nG1a9f8 , \44212 , \42503 );
buf \U$37215 ( \44214 , \44213_nG1a9f8 );
_HMUX g14bb4 ( \44215_nG14bb4 , RIddbc360_3925 , \42775 , \44073 );
_HMUX g14bb5 ( \44216_nG14bb5 , RIddbc360_3925 , \44215_nG14bb4 , \42590 );
_HMUX g14bb7 ( \44217_nG14bb7 , RIddbc360_3925 , \42778 , \44076 );
_HMUX g14bb8 ( \44218_nG14bb8 , \44216_nG14bb5 , \44217_nG14bb7 , \42599 );
buf \U$37216 ( \44219 , \44218_nG14bb8 );
_DC g1a9fa_GF_IsGateDCbyConstraint ( \44220_nG1a9fa , \44219 , \42503 );
buf \U$37217 ( \44221 , \44220_nG1a9fa );
_HMUX g14bba ( \44222_nG14bba , RIddbcb58_3926 , \42784 , \44073 );
_HMUX g14bbb ( \44223_nG14bbb , RIddbcb58_3926 , \44222_nG14bba , \42590 );
_HMUX g14bbd ( \44224_nG14bbd , RIddbcb58_3926 , \42787 , \44076 );
_HMUX g14bbe ( \44225_nG14bbe , \44223_nG14bbb , \44224_nG14bbd , \42599 );
buf \U$37218 ( \44226 , \44225_nG14bbe );
_DC g1a9fc_GF_IsGateDCbyConstraint ( \44227_nG1a9fc , \44226 , \42503 );
buf \U$37219 ( \44228 , \44227_nG1a9fc );
_HMUX g14bc0 ( \44229_nG14bc0 , RIddbd350_3927 , \42793 , \44073 );
_HMUX g14bc1 ( \44230_nG14bc1 , RIddbd350_3927 , \44229_nG14bc0 , \42590 );
_HMUX g14bc3 ( \44231_nG14bc3 , RIddbd350_3927 , \42796 , \44076 );
_HMUX g14bc4 ( \44232_nG14bc4 , \44230_nG14bc1 , \44231_nG14bc3 , \42599 );
buf \U$37220 ( \44233 , \44232_nG14bc4 );
_DC g1a9fe_GF_IsGateDCbyConstraint ( \44234_nG1a9fe , \44233 , \42503 );
buf \U$37221 ( \44235 , \44234_nG1a9fe );
_HMUX g14bc6 ( \44236_nG14bc6 , RIddbdb48_3928 , \42802 , \44073 );
_HMUX g14bc7 ( \44237_nG14bc7 , RIddbdb48_3928 , \44236_nG14bc6 , \42590 );
_HMUX g14bc9 ( \44238_nG14bc9 , RIddbdb48_3928 , \42805 , \44076 );
_HMUX g14bca ( \44239_nG14bca , \44237_nG14bc7 , \44238_nG14bc9 , \42599 );
buf \U$37222 ( \44240 , \44239_nG14bca );
_DC g1aa00_GF_IsGateDCbyConstraint ( \44241_nG1aa00 , \44240 , \42503 );
buf \U$37223 ( \44242 , \44241_nG1aa00 );
_HMUX g14bcc ( \44243_nG14bcc , RIddbe340_3929 , \42811 , \44073 );
_HMUX g14bcd ( \44244_nG14bcd , RIddbe340_3929 , \44243_nG14bcc , \42590 );
_HMUX g14bcf ( \44245_nG14bcf , RIddbe340_3929 , \42814 , \44076 );
_HMUX g14bd0 ( \44246_nG14bd0 , \44244_nG14bcd , \44245_nG14bcf , \42599 );
buf \U$37224 ( \44247 , \44246_nG14bd0 );
_DC g1aa02_GF_IsGateDCbyConstraint ( \44248_nG1aa02 , \44247 , \42503 );
buf \U$37225 ( \44249 , \44248_nG1aa02 );
_HMUX g14bd2 ( \44250_nG14bd2 , RIddbeb38_3930 , \42820 , \44073 );
_HMUX g14bd3 ( \44251_nG14bd3 , RIddbeb38_3930 , \44250_nG14bd2 , \42590 );
_HMUX g14bd5 ( \44252_nG14bd5 , RIddbeb38_3930 , \42823 , \44076 );
_HMUX g14bd6 ( \44253_nG14bd6 , \44251_nG14bd3 , \44252_nG14bd5 , \42599 );
buf \U$37226 ( \44254 , \44253_nG14bd6 );
_DC g1aa04_GF_IsGateDCbyConstraint ( \44255_nG1aa04 , \44254 , \42503 );
buf \U$37227 ( \44256 , \44255_nG1aa04 );
_HMUX g14bd8 ( \44257_nG14bd8 , RIddbf330_3931 , \42829 , \44073 );
_HMUX g14bd9 ( \44258_nG14bd9 , RIddbf330_3931 , \44257_nG14bd8 , \42590 );
_HMUX g14bdb ( \44259_nG14bdb , RIddbf330_3931 , \42832 , \44076 );
_HMUX g14bdc ( \44260_nG14bdc , \44258_nG14bd9 , \44259_nG14bdb , \42599 );
buf \U$37228 ( \44261 , \44260_nG14bdc );
_DC g1aa06_GF_IsGateDCbyConstraint ( \44262_nG1aa06 , \44261 , \42503 );
buf \U$37229 ( \44263 , \44262_nG1aa06 );
_HMUX g14bde ( \44264_nG14bde , RIddbfb28_3932 , \42838 , \44073 );
_HMUX g14bdf ( \44265_nG14bdf , RIddbfb28_3932 , \44264_nG14bde , \42590 );
_HMUX g14be1 ( \44266_nG14be1 , RIddbfb28_3932 , \42841 , \44076 );
_HMUX g14be2 ( \44267_nG14be2 , \44265_nG14bdf , \44266_nG14be1 , \42599 );
buf \U$37230 ( \44268 , \44267_nG14be2 );
_DC g1aa08_GF_IsGateDCbyConstraint ( \44269_nG1aa08 , \44268 , \42503 );
buf \U$37231 ( \44270 , \44269_nG1aa08 );
_HMUX g14be4 ( \44271_nG14be4 , RIddc0320_3933 , \42847 , \44073 );
_HMUX g14be5 ( \44272_nG14be5 , RIddc0320_3933 , \44271_nG14be4 , \42590 );
_HMUX g14be7 ( \44273_nG14be7 , RIddc0320_3933 , \42850 , \44076 );
_HMUX g14be8 ( \44274_nG14be8 , \44272_nG14be5 , \44273_nG14be7 , \42599 );
buf \U$37232 ( \44275 , \44274_nG14be8 );
_DC g1aa0a_GF_IsGateDCbyConstraint ( \44276_nG1aa0a , \44275 , \42503 );
buf \U$37233 ( \44277 , \44276_nG1aa0a );
_HMUX g14bea ( \44278_nG14bea , RIddc0b18_3934 , \42856 , \44073 );
_HMUX g14beb ( \44279_nG14beb , RIddc0b18_3934 , \44278_nG14bea , \42590 );
_HMUX g14bed ( \44280_nG14bed , RIddc0b18_3934 , \42859 , \44076 );
_HMUX g14bee ( \44281_nG14bee , \44279_nG14beb , \44280_nG14bed , \42599 );
buf \U$37234 ( \44282 , \44281_nG14bee );
_DC g1aa0e_GF_IsGateDCbyConstraint ( \44283_nG1aa0e , \44282 , \42503 );
buf \U$37235 ( \44284 , \44283_nG1aa0e );
_HMUX g14bf0 ( \44285_nG14bf0 , RIddc1310_3935 , \42865 , \44073 );
_HMUX g14bf1 ( \44286_nG14bf1 , RIddc1310_3935 , \44285_nG14bf0 , \42590 );
_HMUX g14bf3 ( \44287_nG14bf3 , RIddc1310_3935 , \42868 , \44076 );
_HMUX g14bf4 ( \44288_nG14bf4 , \44286_nG14bf1 , \44287_nG14bf3 , \42599 );
buf \U$37236 ( \44289 , \44288_nG14bf4 );
_DC g1aa10_GF_IsGateDCbyConstraint ( \44290_nG1aa10 , \44289 , \42503 );
buf \U$37237 ( \44291 , \44290_nG1aa10 );
_HMUX g14bf6 ( \44292_nG14bf6 , RIddc1b08_3936 , \42874 , \44073 );
_HMUX g14bf7 ( \44293_nG14bf7 , RIddc1b08_3936 , \44292_nG14bf6 , \42590 );
_HMUX g14bf9 ( \44294_nG14bf9 , RIddc1b08_3936 , \42877 , \44076 );
_HMUX g14bfa ( \44295_nG14bfa , \44293_nG14bf7 , \44294_nG14bf9 , \42599 );
buf \U$37238 ( \44296 , \44295_nG14bfa );
_DC g1aa12_GF_IsGateDCbyConstraint ( \44297_nG1aa12 , \44296 , \42503 );
buf \U$37239 ( \44298 , \44297_nG1aa12 );
_HMUX g14bfc ( \44299_nG14bfc , RIddc2300_3937 , \42883 , \44073 );
_HMUX g14bfd ( \44300_nG14bfd , RIddc2300_3937 , \44299_nG14bfc , \42590 );
_HMUX g14bff ( \44301_nG14bff , RIddc2300_3937 , \42886 , \44076 );
_HMUX g14c00 ( \44302_nG14c00 , \44300_nG14bfd , \44301_nG14bff , \42599 );
buf \U$37240 ( \44303 , \44302_nG14c00 );
_DC g1aa14_GF_IsGateDCbyConstraint ( \44304_nG1aa14 , \44303 , \42503 );
buf \U$37241 ( \44305 , \44304_nG1aa14 );
_HMUX g14c02 ( \44306_nG14c02 , RIddc2af8_3938 , \42892 , \44073 );
_HMUX g14c03 ( \44307_nG14c03 , RIddc2af8_3938 , \44306_nG14c02 , \42590 );
_HMUX g14c05 ( \44308_nG14c05 , RIddc2af8_3938 , \42895 , \44076 );
_HMUX g14c06 ( \44309_nG14c06 , \44307_nG14c03 , \44308_nG14c05 , \42599 );
buf \U$37242 ( \44310 , \44309_nG14c06 );
_DC g1aa16_GF_IsGateDCbyConstraint ( \44311_nG1aa16 , \44310 , \42503 );
buf \U$37243 ( \44312 , \44311_nG1aa16 );
_HMUX g14c08 ( \44313_nG14c08 , RIddc32f0_3939 , \42901 , \44073 );
_HMUX g14c09 ( \44314_nG14c09 , RIddc32f0_3939 , \44313_nG14c08 , \42590 );
_HMUX g14c0b ( \44315_nG14c0b , RIddc32f0_3939 , \42904 , \44076 );
_HMUX g14c0c ( \44316_nG14c0c , \44314_nG14c09 , \44315_nG14c0b , \42599 );
buf \U$37244 ( \44317 , \44316_nG14c0c );
_DC g1aa18_GF_IsGateDCbyConstraint ( \44318_nG1aa18 , \44317 , \42503 );
buf \U$37245 ( \44319 , \44318_nG1aa18 );
_HMUX g14c0e ( \44320_nG14c0e , RIddc3ae8_3940 , \42910 , \44073 );
_HMUX g14c0f ( \44321_nG14c0f , RIddc3ae8_3940 , \44320_nG14c0e , \42590 );
_HMUX g14c11 ( \44322_nG14c11 , RIddc3ae8_3940 , \42913 , \44076 );
_HMUX g14c12 ( \44323_nG14c12 , \44321_nG14c0f , \44322_nG14c11 , \42599 );
buf \U$37246 ( \44324 , \44323_nG14c12 );
_DC g1aa1a_GF_IsGateDCbyConstraint ( \44325_nG1aa1a , \44324 , \42503 );
buf \U$37247 ( \44326 , \44325_nG1aa1a );
_HMUX g14c14 ( \44327_nG14c14 , RIddc42e0_3941 , \42919 , \44073 );
_HMUX g14c15 ( \44328_nG14c15 , RIddc42e0_3941 , \44327_nG14c14 , \42590 );
_HMUX g14c17 ( \44329_nG14c17 , RIddc42e0_3941 , \42922 , \44076 );
_HMUX g14c18 ( \44330_nG14c18 , \44328_nG14c15 , \44329_nG14c17 , \42599 );
buf \U$37248 ( \44331 , \44330_nG14c18 );
_DC g1aa1c_GF_IsGateDCbyConstraint ( \44332_nG1aa1c , \44331 , \42503 );
buf \U$37249 ( \44333 , \44332_nG1aa1c );
_HMUX g14c1a ( \44334_nG14c1a , RIddc4ad8_3942 , \42928 , \44073 );
_HMUX g14c1b ( \44335_nG14c1b , RIddc4ad8_3942 , \44334_nG14c1a , \42590 );
_HMUX g14c1d ( \44336_nG14c1d , RIddc4ad8_3942 , \42931 , \44076 );
_HMUX g14c1e ( \44337_nG14c1e , \44335_nG14c1b , \44336_nG14c1d , \42599 );
buf \U$37250 ( \44338 , \44337_nG14c1e );
_DC g1aa1e_GF_IsGateDCbyConstraint ( \44339_nG1aa1e , \44338 , \42503 );
buf \U$37251 ( \44340 , \44339_nG1aa1e );
_HMUX g14c20 ( \44341_nG14c20 , RIddc52d0_3943 , \42937 , \44073 );
_HMUX g14c21 ( \44342_nG14c21 , RIddc52d0_3943 , \44341_nG14c20 , \42590 );
_HMUX g14c23 ( \44343_nG14c23 , RIddc52d0_3943 , \42940 , \44076 );
_HMUX g14c24 ( \44344_nG14c24 , \44342_nG14c21 , \44343_nG14c23 , \42599 );
buf \U$37252 ( \44345 , \44344_nG14c24 );
_DC g1aa20_GF_IsGateDCbyConstraint ( \44346_nG1aa20 , \44345 , \42503 );
buf \U$37253 ( \44347 , \44346_nG1aa20 );
_HMUX g14c26 ( \44348_nG14c26 , RIddc5ac8_3944 , \42946 , \44073 );
_HMUX g14c27 ( \44349_nG14c27 , RIddc5ac8_3944 , \44348_nG14c26 , \42590 );
_HMUX g14c29 ( \44350_nG14c29 , RIddc5ac8_3944 , \42949 , \44076 );
_HMUX g14c2a ( \44351_nG14c2a , \44349_nG14c27 , \44350_nG14c29 , \42599 );
buf \U$37254 ( \44352 , \44351_nG14c2a );
_DC g1aa24_GF_IsGateDCbyConstraint ( \44353_nG1aa24 , \44352 , \42503 );
buf \U$37255 ( \44354 , \44353_nG1aa24 );
_HMUX g14c2c ( \44355_nG14c2c , RIddc62c0_3945 , \42955 , \44073 );
_HMUX g14c2d ( \44356_nG14c2d , RIddc62c0_3945 , \44355_nG14c2c , \42590 );
_HMUX g14c2f ( \44357_nG14c2f , RIddc62c0_3945 , \42958 , \44076 );
_HMUX g14c30 ( \44358_nG14c30 , \44356_nG14c2d , \44357_nG14c2f , \42599 );
buf \U$37256 ( \44359 , \44358_nG14c30 );
_DC g1aa26_GF_IsGateDCbyConstraint ( \44360_nG1aa26 , \44359 , \42503 );
buf \U$37257 ( \44361 , \44360_nG1aa26 );
_HMUX g14c32 ( \44362_nG14c32 , RIddc6ab8_3946 , \42964 , \44073 );
_HMUX g14c33 ( \44363_nG14c33 , RIddc6ab8_3946 , \44362_nG14c32 , \42590 );
_HMUX g14c35 ( \44364_nG14c35 , RIddc6ab8_3946 , \42967 , \44076 );
_HMUX g14c36 ( \44365_nG14c36 , \44363_nG14c33 , \44364_nG14c35 , \42599 );
buf \U$37258 ( \44366 , \44365_nG14c36 );
_DC g1aa28_GF_IsGateDCbyConstraint ( \44367_nG1aa28 , \44366 , \42503 );
buf \U$37259 ( \44368 , \44367_nG1aa28 );
_HMUX g14c38 ( \44369_nG14c38 , RIddc72b0_3947 , \42973 , \44073 );
_HMUX g14c39 ( \44370_nG14c39 , RIddc72b0_3947 , \44369_nG14c38 , \42590 );
_HMUX g14c3b ( \44371_nG14c3b , RIddc72b0_3947 , \42976 , \44076 );
_HMUX g14c3c ( \44372_nG14c3c , \44370_nG14c39 , \44371_nG14c3b , \42599 );
buf \U$37260 ( \44373 , \44372_nG14c3c );
_DC g1aa2a_GF_IsGateDCbyConstraint ( \44374_nG1aa2a , \44373 , \42503 );
buf \U$37261 ( \44375 , \44374_nG1aa2a );
_HMUX g14c3e ( \44376_nG14c3e , RIddc7aa8_3948 , \42982 , \44073 );
_HMUX g14c3f ( \44377_nG14c3f , RIddc7aa8_3948 , \44376_nG14c3e , \42590 );
_HMUX g14c41 ( \44378_nG14c41 , RIddc7aa8_3948 , \42985 , \44076 );
_HMUX g14c42 ( \44379_nG14c42 , \44377_nG14c3f , \44378_nG14c41 , \42599 );
buf \U$37262 ( \44380 , \44379_nG14c42 );
_DC g1aa2c_GF_IsGateDCbyConstraint ( \44381_nG1aa2c , \44380 , \42503 );
buf \U$37263 ( \44382 , \44381_nG1aa2c );
_HMUX g14c44 ( \44383_nG14c44 , RIddc82a0_3949 , \42991 , \44073 );
_HMUX g14c45 ( \44384_nG14c45 , RIddc82a0_3949 , \44383_nG14c44 , \42590 );
_HMUX g14c47 ( \44385_nG14c47 , RIddc82a0_3949 , \42994 , \44076 );
_HMUX g14c48 ( \44386_nG14c48 , \44384_nG14c45 , \44385_nG14c47 , \42599 );
buf \U$37264 ( \44387 , \44386_nG14c48 );
_DC g1aa2e_GF_IsGateDCbyConstraint ( \44388_nG1aa2e , \44387 , \42503 );
buf \U$37265 ( \44389 , \44388_nG1aa2e );
_HMUX g14c4a ( \44390_nG14c4a , RIddc8a98_3950 , \43000 , \44073 );
_HMUX g14c4b ( \44391_nG14c4b , RIddc8a98_3950 , \44390_nG14c4a , \42590 );
_HMUX g14c4d ( \44392_nG14c4d , RIddc8a98_3950 , \43003 , \44076 );
_HMUX g14c4e ( \44393_nG14c4e , \44391_nG14c4b , \44392_nG14c4d , \42599 );
buf \U$37266 ( \44394 , \44393_nG14c4e );
_DC g1aa30_GF_IsGateDCbyConstraint ( \44395_nG1aa30 , \44394 , \42503 );
buf \U$37267 ( \44396 , \44395_nG1aa30 );
_HMUX g14c50 ( \44397_nG14c50 , RIddc9290_3951 , \43009 , \44073 );
_HMUX g14c51 ( \44398_nG14c51 , RIddc9290_3951 , \44397_nG14c50 , \42590 );
_HMUX g14c53 ( \44399_nG14c53 , RIddc9290_3951 , \43012 , \44076 );
_HMUX g14c54 ( \44400_nG14c54 , \44398_nG14c51 , \44399_nG14c53 , \42599 );
buf \U$37268 ( \44401 , \44400_nG14c54 );
_DC g1aa32_GF_IsGateDCbyConstraint ( \44402_nG1aa32 , \44401 , \42503 );
buf \U$37269 ( \44403 , \44402_nG1aa32 );
_HMUX g14c56 ( \44404_nG14c56 , RIddc9a88_3952 , \43018 , \44073 );
_HMUX g14c57 ( \44405_nG14c57 , RIddc9a88_3952 , \44404_nG14c56 , \42590 );
_HMUX g14c59 ( \44406_nG14c59 , RIddc9a88_3952 , \43021 , \44076 );
_HMUX g14c5a ( \44407_nG14c5a , \44405_nG14c57 , \44406_nG14c59 , \42599 );
buf \U$37270 ( \44408 , \44407_nG14c5a );
_DC g1aa34_GF_IsGateDCbyConstraint ( \44409_nG1aa34 , \44408 , \42503 );
buf \U$37271 ( \44410 , \44409_nG1aa34 );
_HMUX g14c5c ( \44411_nG14c5c , RIddca280_3953 , \43027 , \44073 );
_HMUX g14c5d ( \44412_nG14c5d , RIddca280_3953 , \44411_nG14c5c , \42590 );
_HMUX g14c5f ( \44413_nG14c5f , RIddca280_3953 , \43030 , \44076 );
_HMUX g14c60 ( \44414_nG14c60 , \44412_nG14c5d , \44413_nG14c5f , \42599 );
buf \U$37272 ( \44415 , \44414_nG14c60 );
_DC g1aa36_GF_IsGateDCbyConstraint ( \44416_nG1aa36 , \44415 , \42503 );
buf \U$37273 ( \44417 , \44416_nG1aa36 );
_HMUX g14c62 ( \44418_nG14c62 , RIddcaa78_3954 , \43036 , \44073 );
_HMUX g14c63 ( \44419_nG14c63 , RIddcaa78_3954 , \44418_nG14c62 , \42590 );
_HMUX g14c65 ( \44420_nG14c65 , RIddcaa78_3954 , \43039 , \44076 );
_HMUX g14c66 ( \44421_nG14c66 , \44419_nG14c63 , \44420_nG14c65 , \42599 );
buf \U$37274 ( \44422 , \44421_nG14c66 );
_DC g1aa3a_GF_IsGateDCbyConstraint ( \44423_nG1aa3a , \44422 , \42503 );
buf \U$37275 ( \44424 , \44423_nG1aa3a );
_HMUX g14c68 ( \44425_nG14c68 , RIddcb270_3955 , \43045 , \44073 );
_HMUX g14c69 ( \44426_nG14c69 , RIddcb270_3955 , \44425_nG14c68 , \42590 );
_HMUX g14c6b ( \44427_nG14c6b , RIddcb270_3955 , \43048 , \44076 );
_HMUX g14c6c ( \44428_nG14c6c , \44426_nG14c69 , \44427_nG14c6b , \42599 );
buf \U$37276 ( \44429 , \44428_nG14c6c );
_DC g1aa3c_GF_IsGateDCbyConstraint ( \44430_nG1aa3c , \44429 , \42503 );
buf \U$37277 ( \44431 , \44430_nG1aa3c );
_HMUX g14c6e ( \44432_nG14c6e , RIddcba68_3956 , \43054 , \44073 );
_HMUX g14c6f ( \44433_nG14c6f , RIddcba68_3956 , \44432_nG14c6e , \42590 );
_HMUX g14c71 ( \44434_nG14c71 , RIddcba68_3956 , \43057 , \44076 );
_HMUX g14c72 ( \44435_nG14c72 , \44433_nG14c6f , \44434_nG14c71 , \42599 );
buf \U$37278 ( \44436 , \44435_nG14c72 );
_DC g1aa3e_GF_IsGateDCbyConstraint ( \44437_nG1aa3e , \44436 , \42503 );
buf \U$37279 ( \44438 , \44437_nG1aa3e );
_HMUX g14c74 ( \44439_nG14c74 , RIddcc260_3957 , \43063 , \44073 );
_HMUX g14c75 ( \44440_nG14c75 , RIddcc260_3957 , \44439_nG14c74 , \42590 );
_HMUX g14c77 ( \44441_nG14c77 , RIddcc260_3957 , \43066 , \44076 );
_HMUX g14c78 ( \44442_nG14c78 , \44440_nG14c75 , \44441_nG14c77 , \42599 );
buf \U$37280 ( \44443 , \44442_nG14c78 );
_DC g1aa40_GF_IsGateDCbyConstraint ( \44444_nG1aa40 , \44443 , \42503 );
buf \U$37281 ( \44445 , \44444_nG1aa40 );
_HMUX g14c7a ( \44446_nG14c7a , RIddcca58_3958 , \43072 , \44073 );
_HMUX g14c7b ( \44447_nG14c7b , RIddcca58_3958 , \44446_nG14c7a , \42590 );
_HMUX g14c7d ( \44448_nG14c7d , RIddcca58_3958 , \43075 , \44076 );
_HMUX g14c7e ( \44449_nG14c7e , \44447_nG14c7b , \44448_nG14c7d , \42599 );
buf \U$37282 ( \44450 , \44449_nG14c7e );
_DC g1aa42_GF_IsGateDCbyConstraint ( \44451_nG1aa42 , \44450 , \42503 );
buf \U$37283 ( \44452 , \44451_nG1aa42 );
_HMUX g14c80 ( \44453_nG14c80 , RIddcd250_3959 , \43081 , \44073 );
_HMUX g14c81 ( \44454_nG14c81 , RIddcd250_3959 , \44453_nG14c80 , \42590 );
_HMUX g14c83 ( \44455_nG14c83 , RIddcd250_3959 , \43084 , \44076 );
_HMUX g14c84 ( \44456_nG14c84 , \44454_nG14c81 , \44455_nG14c83 , \42599 );
buf \U$37284 ( \44457 , \44456_nG14c84 );
_DC g1aa44_GF_IsGateDCbyConstraint ( \44458_nG1aa44 , \44457 , \42503 );
buf \U$37285 ( \44459 , \44458_nG1aa44 );
_HMUX g14c86 ( \44460_nG14c86 , RIddcda48_3960 , \43090 , \44073 );
_HMUX g14c87 ( \44461_nG14c87 , RIddcda48_3960 , \44460_nG14c86 , \42590 );
_HMUX g14c89 ( \44462_nG14c89 , RIddcda48_3960 , \43093 , \44076 );
_HMUX g14c8a ( \44463_nG14c8a , \44461_nG14c87 , \44462_nG14c89 , \42599 );
buf \U$37286 ( \44464 , \44463_nG14c8a );
_DC g1aa46_GF_IsGateDCbyConstraint ( \44465_nG1aa46 , \44464 , \42503 );
buf \U$37287 ( \44466 , \44465_nG1aa46 );
_HMUX g14c8c ( \44467_nG14c8c , RIddce240_3961 , \43099 , \44073 );
_HMUX g14c8d ( \44468_nG14c8d , RIddce240_3961 , \44467_nG14c8c , \42590 );
_HMUX g14c8f ( \44469_nG14c8f , RIddce240_3961 , \43102 , \44076 );
_HMUX g14c90 ( \44470_nG14c90 , \44468_nG14c8d , \44469_nG14c8f , \42599 );
buf \U$37288 ( \44471 , \44470_nG14c90 );
_DC g1aa48_GF_IsGateDCbyConstraint ( \44472_nG1aa48 , \44471 , \42503 );
buf \U$37289 ( \44473 , \44472_nG1aa48 );
_HMUX g14c92 ( \44474_nG14c92 , RIddcea38_3962 , \43108 , \44073 );
_HMUX g14c93 ( \44475_nG14c93 , RIddcea38_3962 , \44474_nG14c92 , \42590 );
_HMUX g14c95 ( \44476_nG14c95 , RIddcea38_3962 , \43111 , \44076 );
_HMUX g14c96 ( \44477_nG14c96 , \44475_nG14c93 , \44476_nG14c95 , \42599 );
buf \U$37290 ( \44478 , \44477_nG14c96 );
_DC g1aa4a_GF_IsGateDCbyConstraint ( \44479_nG1aa4a , \44478 , \42503 );
buf \U$37291 ( \44480 , \44479_nG1aa4a );
_HMUX g14c98 ( \44481_nG14c98 , RIddcf230_3963 , \43117 , \44073 );
_HMUX g14c99 ( \44482_nG14c99 , RIddcf230_3963 , \44481_nG14c98 , \42590 );
_HMUX g14c9b ( \44483_nG14c9b , RIddcf230_3963 , \43120 , \44076 );
_HMUX g14c9c ( \44484_nG14c9c , \44482_nG14c99 , \44483_nG14c9b , \42599 );
buf \U$37292 ( \44485 , \44484_nG14c9c );
_DC g1aa4c_GF_IsGateDCbyConstraint ( \44486_nG1aa4c , \44485 , \42503 );
buf \U$37293 ( \44487 , \44486_nG1aa4c );
_HMUX g14c9e ( \44488_nG14c9e , RIddcfa28_3964 , \43126 , \44073 );
_HMUX g14c9f ( \44489_nG14c9f , RIddcfa28_3964 , \44488_nG14c9e , \42590 );
_HMUX g14ca1 ( \44490_nG14ca1 , RIddcfa28_3964 , \43129 , \44076 );
_HMUX g14ca2 ( \44491_nG14ca2 , \44489_nG14c9f , \44490_nG14ca1 , \42599 );
buf \U$37294 ( \44492 , \44491_nG14ca2 );
_DC g1aa50_GF_IsGateDCbyConstraint ( \44493_nG1aa50 , \44492 , \42503 );
buf \U$37295 ( \44494 , \44493_nG1aa50 );
_HMUX g14ca4 ( \44495_nG14ca4 , RIddd0220_3965 , \43135 , \44073 );
_HMUX g14ca5 ( \44496_nG14ca5 , RIddd0220_3965 , \44495_nG14ca4 , \42590 );
_HMUX g14ca7 ( \44497_nG14ca7 , RIddd0220_3965 , \43138 , \44076 );
_HMUX g14ca8 ( \44498_nG14ca8 , \44496_nG14ca5 , \44497_nG14ca7 , \42599 );
buf \U$37296 ( \44499 , \44498_nG14ca8 );
_DC g1aa52_GF_IsGateDCbyConstraint ( \44500_nG1aa52 , \44499 , \42503 );
buf \U$37297 ( \44501 , \44500_nG1aa52 );
_HMUX g14caa ( \44502_nG14caa , RIddd0a18_3966 , \43144 , \44073 );
_HMUX g14cab ( \44503_nG14cab , RIddd0a18_3966 , \44502_nG14caa , \42590 );
_HMUX g14cad ( \44504_nG14cad , RIddd0a18_3966 , \43147 , \44076 );
_HMUX g14cae ( \44505_nG14cae , \44503_nG14cab , \44504_nG14cad , \42599 );
buf \U$37298 ( \44506 , \44505_nG14cae );
_DC g1aa54_GF_IsGateDCbyConstraint ( \44507_nG1aa54 , \44506 , \42503 );
buf \U$37299 ( \44508 , \44507_nG1aa54 );
_HMUX g14cb0 ( \44509_nG14cb0 , RIddd1210_3967 , \43153 , \44073 );
_HMUX g14cb1 ( \44510_nG14cb1 , RIddd1210_3967 , \44509_nG14cb0 , \42590 );
_HMUX g14cb3 ( \44511_nG14cb3 , RIddd1210_3967 , \43156 , \44076 );
_HMUX g14cb4 ( \44512_nG14cb4 , \44510_nG14cb1 , \44511_nG14cb3 , \42599 );
buf \U$37300 ( \44513 , \44512_nG14cb4 );
_DC g1aa56_GF_IsGateDCbyConstraint ( \44514_nG1aa56 , \44513 , \42503 );
buf \U$37301 ( \44515 , \44514_nG1aa56 );
_HMUX g14cb6 ( \44516_nG14cb6 , RIddd1a08_3968 , \43162 , \44073 );
_HMUX g14cb7 ( \44517_nG14cb7 , RIddd1a08_3968 , \44516_nG14cb6 , \42590 );
_HMUX g14cb9 ( \44518_nG14cb9 , RIddd1a08_3968 , \43165 , \44076 );
_HMUX g14cba ( \44519_nG14cba , \44517_nG14cb7 , \44518_nG14cb9 , \42599 );
buf \U$37302 ( \44520 , \44519_nG14cba );
_DC g1aa58_GF_IsGateDCbyConstraint ( \44521_nG1aa58 , \44520 , \42503 );
buf \U$37303 ( \44522 , \44521_nG1aa58 );
buf \U$37304 ( \44523 , RIb86fc68_77);
_HMUX g14b0b ( \44524_nG14b0b , RIdc0fbb8_3681 , \44523 , \42581 );
not \U$37305 ( \44525 , \42590 );
or \U$37306 ( \44526 , \42599 , \44525 );
_HMUX g14b0c ( \44527_nG14b0c , \44524_nG14b0b , RIdc0fbb8_3681 , \44526 );
buf \U$37307 ( \44528 , \44527_nG14b0c );
_DC g1a9c8_GF_IsGateDCbyConstraint ( \44529_nG1a9c8 , \44528 , \42503 );
buf \U$37308 ( \44530 , \44529_nG1a9c8 );
buf \U$37309 ( \44531 , RIb86fce0_76);
_HMUX g14b0d ( \44532_nG14b0d , RIdc0f0f0_3682 , \44531 , \42581 );
_HMUX g14b0e ( \44533_nG14b0e , \44532_nG14b0d , RIdc0f0f0_3682 , \44526 );
buf \U$37310 ( \44534 , \44533_nG14b0e );
_DC g1a9ca_GF_IsGateDCbyConstraint ( \44535_nG1a9ca , \44534 , \42503 );
buf \U$37311 ( \44536 , \44535_nG1a9ca );
buf \U$37312 ( \44537 , RIb86fd58_75);
_HMUX g14b0f ( \44538_nG14b0f , RIdc0e5b0_3683 , \44537 , \42581 );
_HMUX g14b10 ( \44539_nG14b10 , \44538_nG14b0f , RIdc0e5b0_3683 , \44526 );
buf \U$37313 ( \44540 , \44539_nG14b10 );
_DC g1a9cc_GF_IsGateDCbyConstraint ( \44541_nG1a9cc , \44540 , \42503 );
buf \U$37314 ( \44542 , \44541_nG1a9cc );
buf \U$37315 ( \44543 , RIb87e8a8_74);
_HMUX g14b11 ( \44544_nG14b11 , RIdc0dae8_3684 , \44543 , \42581 );
_HMUX g14b12 ( \44545_nG14b12 , \44544_nG14b11 , RIdc0dae8_3684 , \44526 );
buf \U$37316 ( \44546 , \44545_nG14b12 );
_DC g1a9ce_GF_IsGateDCbyConstraint ( \44547_nG1a9ce , \44546 , \42503 );
buf \U$37317 ( \44548 , \44547_nG1a9ce );
buf \U$37318 ( \44549 , RIb87e920_73);
_HMUX g14b13 ( \44550_nG14b13 , RIdc0cfa8_3685 , \44549 , \42581 );
_HMUX g14b14 ( \44551_nG14b14 , \44550_nG14b13 , RIdc0cfa8_3685 , \44526 );
buf \U$37319 ( \44552 , \44551_nG14b14 );
_DC g1a9d0_GF_IsGateDCbyConstraint ( \44553_nG1a9d0 , \44552 , \42503 );
buf \U$37320 ( \44554 , \44553_nG1a9d0 );
buf \U$37321 ( \44555 , RIb87e998_72);
_HMUX g14b15 ( \44556_nG14b15 , RIdc0c3f0_3686 , \44555 , \42581 );
_HMUX g14b16 ( \44557_nG14b16 , \44556_nG14b15 , RIdc0c3f0_3686 , \44526 );
buf \U$37322 ( \44558 , \44557_nG14b16 );
_DC g1a9d2_GF_IsGateDCbyConstraint ( \44559_nG1a9d2 , \44558 , \42503 );
buf \U$37323 ( \44560 , \44559_nG1a9d2 );
buf \U$37324 ( \44561 , RIb87ea10_71);
_HMUX g14b17 ( \44562_nG14b17 , RIdc0b7c0_3687 , \44561 , \42581 );
_HMUX g14b18 ( \44563_nG14b18 , \44562_nG14b17 , RIdc0b7c0_3687 , \44526 );
buf \U$37325 ( \44564 , \44563_nG14b18 );
_DC g1a9d4_GF_IsGateDCbyConstraint ( \44565_nG1a9d4 , \44564 , \42503 );
buf \U$37326 ( \44566 , \44565_nG1a9d4 );
buf \U$37327 ( \44567 , RIb87ea88_70);
_HMUX g14b19 ( \44568_nG14b19 , RIdc0ac08_3688 , \44567 , \42581 );
_HMUX g14b1a ( \44569_nG14b1a , \44568_nG14b19 , RIdc0ac08_3688 , \44526 );
buf \U$37328 ( \44570 , \44569_nG14b1a );
_DC g1a9d6_GF_IsGateDCbyConstraint ( \44571_nG1a9d6 , \44570 , \42503 );
buf \U$37329 ( \44572 , \44571_nG1a9d6 );
_HMUX g14afa ( \44573_nG14afa , RIdc09f60_3689 , \44523 , \43172 );
_HMUX g14afb ( \44574_nG14afb , \44573_nG14afa , RIdc09f60_3689 , \44526 );
buf \U$37330 ( \44575 , \44574_nG14afb );
_DC g1a9b8_GF_IsGateDCbyConstraint ( \44576_nG1a9b8 , \44575 , \42503 );
buf \U$37331 ( \44577 , \44576_nG1a9b8 );
_HMUX g14afc ( \44578_nG14afc , RIdc093a8_3690 , \44531 , \43172 );
_HMUX g14afd ( \44579_nG14afd , \44578_nG14afc , RIdc093a8_3690 , \44526 );
buf \U$37332 ( \44580 , \44579_nG14afd );
_DC g1a9ba_GF_IsGateDCbyConstraint ( \44581_nG1a9ba , \44580 , \42503 );
buf \U$37333 ( \44582 , \44581_nG1a9ba );
_HMUX g14afe ( \44583_nG14afe , RIdc08700_3691 , \44537 , \43172 );
_HMUX g14aff ( \44584_nG14aff , \44583_nG14afe , RIdc08700_3691 , \44526 );
buf \U$37334 ( \44585 , \44584_nG14aff );
_DC g1a9bc_GF_IsGateDCbyConstraint ( \44586_nG1a9bc , \44585 , \42503 );
buf \U$37335 ( \44587 , \44586_nG1a9bc );
_HMUX g14b00 ( \44588_nG14b00 , RIdc07878_3692 , \44543 , \43172 );
_HMUX g14b01 ( \44589_nG14b01 , \44588_nG14b00 , RIdc07878_3692 , \44526 );
buf \U$37336 ( \44590 , \44589_nG14b01 );
_DC g1a9be_GF_IsGateDCbyConstraint ( \44591_nG1a9be , \44590 , \42503 );
buf \U$37337 ( \44592 , \44591_nG1a9be );
_HMUX g14b02 ( \44593_nG14b02 , RIdc06270_3693 , \44549 , \43172 );
_HMUX g14b03 ( \44594_nG14b03 , \44593_nG14b02 , RIdc06270_3693 , \44526 );
buf \U$37338 ( \44595 , \44594_nG14b03 );
_DC g1a9c0_GF_IsGateDCbyConstraint ( \44596_nG1a9c0 , \44595 , \42503 );
buf \U$37339 ( \44597 , \44596_nG1a9c0 );
_HMUX g14b04 ( \44598_nG14b04 , RIdc05118_3694 , \44555 , \43172 );
_HMUX g14b05 ( \44599_nG14b05 , \44598_nG14b04 , RIdc05118_3694 , \44526 );
buf \U$37340 ( \44600 , \44599_nG14b05 );
_DC g1a9c2_GF_IsGateDCbyConstraint ( \44601_nG1a9c2 , \44600 , \42503 );
buf \U$37341 ( \44602 , \44601_nG1a9c2 );
_HMUX g14b06 ( \44603_nG14b06 , RIdc03b10_3695 , \44561 , \43172 );
_HMUX g14b07 ( \44604_nG14b07 , \44603_nG14b06 , RIdc03b10_3695 , \44526 );
buf \U$37342 ( \44605 , \44604_nG14b07 );
_DC g1a9c4_GF_IsGateDCbyConstraint ( \44606_nG1a9c4 , \44605 , \42503 );
buf \U$37343 ( \44607 , \44606_nG1a9c4 );
_HMUX g14b08 ( \44608_nG14b08 , RIdc029b8_3696 , \44567 , \43172 );
_HMUX g14b09 ( \44609_nG14b09 , \44608_nG14b08 , RIdc029b8_3696 , \44526 );
buf \U$37344 ( \44610 , \44609_nG14b09 );
_DC g1a9c6_GF_IsGateDCbyConstraint ( \44611_nG1a9c6 , \44610 , \42503 );
buf \U$37345 ( \44612 , \44611_nG1a9c6 );
_HMUX g14ae9 ( \44613_nG14ae9 , RIdc013b0_3697 , \44523 , \43623 );
_HMUX g14aea ( \44614_nG14aea , \44613_nG14ae9 , RIdc013b0_3697 , \44526 );
buf \U$37346 ( \44615 , \44614_nG14aea );
_DC g1a9a8_GF_IsGateDCbyConstraint ( \44616_nG1a9a8 , \44615 , \42503 );
buf \U$37347 ( \44617 , \44616_nG1a9a8 );
_HMUX g14aeb ( \44618_nG14aeb , RIdc00258_3698 , \44531 , \43623 );
_HMUX g14aec ( \44619_nG14aec , \44618_nG14aeb , RIdc00258_3698 , \44526 );
buf \U$37348 ( \44620 , \44619_nG14aec );
_DC g1a9aa_GF_IsGateDCbyConstraint ( \44621_nG1a9aa , \44620 , \42503 );
buf \U$37349 ( \44622 , \44621_nG1a9aa );
_HMUX g14aed ( \44623_nG14aed , RIdbff100_3699 , \44537 , \43623 );
_HMUX g14aee ( \44624_nG14aee , \44623_nG14aed , RIdbff100_3699 , \44526 );
buf \U$37350 ( \44625 , \44624_nG14aee );
_DC g1a9ac_GF_IsGateDCbyConstraint ( \44626_nG1a9ac , \44625 , \42503 );
buf \U$37351 ( \44627 , \44626_nG1a9ac );
_HMUX g14aef ( \44628_nG14aef , RIdbfdaf8_3700 , \44543 , \43623 );
_HMUX g14af0 ( \44629_nG14af0 , \44628_nG14aef , RIdbfdaf8_3700 , \44526 );
buf \U$37352 ( \44630 , \44629_nG14af0 );
_DC g1a9ae_GF_IsGateDCbyConstraint ( \44631_nG1a9ae , \44630 , \42503 );
buf \U$37353 ( \44632 , \44631_nG1a9ae );
_HMUX g14af1 ( \44633_nG14af1 , RIdbfc9a0_3701 , \44549 , \43623 );
_HMUX g14af2 ( \44634_nG14af2 , \44633_nG14af1 , RIdbfc9a0_3701 , \44526 );
buf \U$37354 ( \44635 , \44634_nG14af2 );
_DC g1a9b0_GF_IsGateDCbyConstraint ( \44636_nG1a9b0 , \44635 , \42503 );
buf \U$37355 ( \44637 , \44636_nG1a9b0 );
_HMUX g14af3 ( \44638_nG14af3 , RIdbfb398_3702 , \44555 , \43623 );
_HMUX g14af4 ( \44639_nG14af4 , \44638_nG14af3 , RIdbfb398_3702 , \44526 );
buf \U$37356 ( \44640 , \44639_nG14af4 );
_DC g1a9b2_GF_IsGateDCbyConstraint ( \44641_nG1a9b2 , \44640 , \42503 );
buf \U$37357 ( \44642 , \44641_nG1a9b2 );
_HMUX g14af5 ( \44643_nG14af5 , RIdbfa240_3703 , \44561 , \43623 );
_HMUX g14af6 ( \44644_nG14af6 , \44643_nG14af5 , RIdbfa240_3703 , \44526 );
buf \U$37358 ( \44645 , \44644_nG14af6 );
_DC g1a9b4_GF_IsGateDCbyConstraint ( \44646_nG1a9b4 , \44645 , \42503 );
buf \U$37359 ( \44647 , \44646_nG1a9b4 );
_HMUX g14af7 ( \44648_nG14af7 , RIdbf8c38_3704 , \44567 , \43623 );
_HMUX g14af8 ( \44649_nG14af8 , \44648_nG14af7 , RIdbf8c38_3704 , \44526 );
buf \U$37360 ( \44650 , \44649_nG14af8 );
_DC g1a9b6_GF_IsGateDCbyConstraint ( \44651_nG1a9b6 , \44650 , \42503 );
buf \U$37361 ( \44652 , \44651_nG1a9b6 );
_HMUX g14ac8 ( \44653_nG14ac8 , RIdbf7ae0_3705 , \44523 , \44073 );
_HMUX g14ad1 ( \44654_nG14ad1 , \44653_nG14ac8 , RIdbf7ae0_3705 , \44526 );
buf \U$37362 ( \44655 , \44654_nG14ad1 );
_DC g1abe0_GF_IsGateDCbyConstraint ( \44656_nG1abe0 , \44655 , \42503 );
buf \U$37363 ( \44657 , \44656_nG1abe0 );
_HMUX g14ad3 ( \44658_nG14ad3 , RIdbf6988_3706 , \44531 , \44073 );
_HMUX g14ad4 ( \44659_nG14ad4 , \44658_nG14ad3 , RIdbf6988_3706 , \44526 );
buf \U$37364 ( \44660 , \44659_nG14ad4 );
_DC g1abe2_GF_IsGateDCbyConstraint ( \44661_nG1abe2 , \44660 , \42503 );
buf \U$37365 ( \44662 , \44661_nG1abe2 );
_HMUX g14ad6 ( \44663_nG14ad6 , RIdbf5380_3707 , \44537 , \44073 );
_HMUX g14ad7 ( \44664_nG14ad7 , \44663_nG14ad6 , RIdbf5380_3707 , \44526 );
buf \U$37366 ( \44665 , \44664_nG14ad7 );
_DC g1abe4_GF_IsGateDCbyConstraint ( \44666_nG1abe4 , \44665 , \42503 );
buf \U$37367 ( \44667 , \44666_nG1abe4 );
_HMUX g14ad9 ( \44668_nG14ad9 , RIdbf4228_3708 , \44543 , \44073 );
_HMUX g14ada ( \44669_nG14ada , \44668_nG14ad9 , RIdbf4228_3708 , \44526 );
buf \U$37368 ( \44670 , \44669_nG14ada );
_DC g1abe6_GF_IsGateDCbyConstraint ( \44671_nG1abe6 , \44670 , \42503 );
buf \U$37369 ( \44672 , \44671_nG1abe6 );
_HMUX g14adc ( \44673_nG14adc , RIdbf2c20_3709 , \44549 , \44073 );
_HMUX g14add ( \44674_nG14add , \44673_nG14adc , RIdbf2c20_3709 , \44526 );
buf \U$37370 ( \44675 , \44674_nG14add );
_DC g1abe8_GF_IsGateDCbyConstraint ( \44676_nG1abe8 , \44675 , \42503 );
buf \U$37371 ( \44677 , \44676_nG1abe8 );
_HMUX g14adf ( \44678_nG14adf , RIdbf1ac8_3710 , \44555 , \44073 );
_HMUX g14ae0 ( \44679_nG14ae0 , \44678_nG14adf , RIdbf1ac8_3710 , \44526 );
buf \U$37372 ( \44680 , \44679_nG14ae0 );
_DC g1abea_GF_IsGateDCbyConstraint ( \44681_nG1abea , \44680 , \42503 );
buf \U$37373 ( \44682 , \44681_nG1abea );
_HMUX g14ae2 ( \44683_nG14ae2 , RIdbf04c0_3711 , \44561 , \44073 );
_HMUX g14ae3 ( \44684_nG14ae3 , \44683_nG14ae2 , RIdbf04c0_3711 , \44526 );
buf \U$37374 ( \44685 , \44684_nG14ae3 );
_DC g1abec_GF_IsGateDCbyConstraint ( \44686_nG1abec , \44685 , \42503 );
buf \U$37375 ( \44687 , \44686_nG1abec );
_HMUX g14ae5 ( \44688_nG14ae5 , RIdbef368_3712 , \44567 , \44073 );
_HMUX g14ae6 ( \44689_nG14ae6 , \44688_nG14ae5 , RIdbef368_3712 , \44526 );
buf \U$37376 ( \44690 , \44689_nG14ae6 );
_DC g1abee_GF_IsGateDCbyConstraint ( \44691_nG1abee , \44690 , \42503 );
buf \U$37377 ( \44692 , \44691_nG1abee );
and \U$37379 ( \44693 , \42317 , RIb79b428_272);
_HMUX gbcb6 ( \44694_nGbcb6 , RIe5349b0_6879 , 1'b1 , \44693 );
and \U$37380 ( \44695 , \42390 , RIb8396e0_155);
not \U$37381 ( \44696 , \44695 );
and \U$37382 ( \44697 , \44694_nGbcb6 , \44696 );
_DC g1ac03_GF_IsGateDCbyConstraint ( \44698_nG1ac03 , \44697 , \42503 );
buf \U$37383 ( \44699 , \44698_nG1ac03 );
buf \U$37384 ( \44700 , RIe5efc28_6741);
nor \U$37385 ( \44701 , \42121_nGbbbc , \42169_nGbbec , \42218_nGbc1c , \42267_nGbc4c , \42316 );
and \U$37386 ( \44702 , \44700 , \44701 );
buf \U$37387 ( \44703 , RIe527288_6346);
and \U$37388 ( \44704 , \42121_nGbbbc , \42169_nGbbec , \42218_nGbc1c , \42267_nGbc4c , \42316 );
and \U$37389 ( \44705 , \44703 , \44704 );
buf \U$37390 ( \44706 , RIe45e528_5951);
not \U$37391 ( \44707 , \42121_nGbbbc );
and \U$37392 ( \44708 , \44707 , \42169_nGbbec , \42218_nGbc1c , \42267_nGbc4c , \42316 );
and \U$37393 ( \44709 , \44706 , \44708 );
buf \U$37394 ( \44710 , RIe395df8_5556);
and \U$37395 ( \44711 , \42121_nGbbbc , \42170 , \42218_nGbc1c , \42267_nGbc4c , \42316 );
and \U$37396 ( \44712 , \44710 , \44711 );
buf \U$37397 ( \44713 , RIe1ca840_5161);
and \U$37398 ( \44714 , \44707 , \42170 , \42218_nGbc1c , \42267_nGbc4c , \42316 );
and \U$37399 ( \44715 , \44713 , \44714 );
buf \U$37400 ( \44716 , RIe100460_4766);
and \U$37401 ( \44717 , \42121_nGbbbc , \42169_nGbbec , \42219 , \42267_nGbc4c , \42316 );
and \U$37402 ( \44718 , \44716 , \44717 );
buf \U$37403 ( \44719 , RIe036f80_4371);
and \U$37404 ( \44720 , \44707 , \42169_nGbbec , \42219 , \42267_nGbc4c , \42316 );
and \U$37405 ( \44721 , \44719 , \44720 );
buf \U$37406 ( \44722 , RIde6b9c8_3976);
and \U$37407 ( \44723 , \42121_nGbbbc , \42170 , \42219 , \42267_nGbc4c , \42316 );
and \U$37408 ( \44724 , \44722 , \44723 );
buf \U$37409 ( \44725 , RIdda31a8_3581);
and \U$37410 ( \44726 , \44707 , \42170 , \42219 , \42267_nGbc4c , \42316 );
and \U$37411 ( \44727 , \44725 , \44726 );
buf \U$37412 ( \44728 , RIdbd9c48_3186);
nor \U$37413 ( \44729 , \44707 , \42170 , \42219 , \42267_nGbc4c , \42315_nGbc7c );
and \U$37414 ( \44730 , \44728 , \44729 );
buf \U$37415 ( \44731 , RIdb0e968_2791);
nor \U$37416 ( \44732 , \42121_nGbbbc , \42170 , \42219 , \42267_nGbc4c , \42315_nGbc7c );
and \U$37417 ( \44733 , \44731 , \44732 );
buf \U$37418 ( \44734 , RIda3bc30_2396);
nor \U$37419 ( \44735 , \44707 , \42169_nGbbec , \42219 , \42267_nGbc4c , \42315_nGbc7c );
and \U$37420 ( \44736 , \44734 , \44735 );
buf \U$37421 ( \44737 , RId987e10_2001);
nor \U$37422 ( \44738 , \42121_nGbbbc , \42169_nGbbec , \42219 , \42267_nGbc4c , \42315_nGbc7c );
and \U$37423 ( \44739 , \44737 , \44738 );
buf \U$37424 ( \44740 , RId8bc950_1606);
nor \U$37425 ( \44741 , \44707 , \42170 , \42218_nGbc1c , \42267_nGbc4c , \42315_nGbc7c );
and \U$37426 ( \44742 , \44740 , \44741 );
buf \U$37427 ( \44743 , RId7f4028_1211);
nor \U$37428 ( \44744 , \42121_nGbbbc , \42170 , \42218_nGbc1c , \42267_nGbc4c , \42315_nGbc7c );
and \U$37429 ( \44745 , \44743 , \44744 );
buf \U$37430 ( \44746 , RId72b4a8_816);
nor \U$37431 ( \44747 , \44707 , \42169_nGbbec , \42218_nGbc1c , \42267_nGbc4c , \42315_nGbc7c );
and \U$37432 ( \44748 , \44746 , \44747 );
or \U$37433 ( \44749 , \44702 , \44705 , \44709 , \44712 , \44715 , \44718 , \44721 , \44724 , \44727 , \44730 , \44733 , \44736 , \44739 , \44742 , \44745 , \44748 );
buf \U$37434 ( \44750 , \42169_nGbbec );
buf \U$37435 ( \44751 , \42218_nGbc1c );
buf \U$37436 ( \44752 , \42267_nGbc4c );
buf \U$37437 ( \44753 , \42315_nGbc7c );
buf \U$37438 ( \44754 , \42121_nGbbbc );
nor \U$37439 ( \44755 , \44750 , \44751 , \44752 , \44753 , \44754 );
buf \U$37440 ( \44756 , \44755 );
buf \U$37441 ( \44757 , \42315_nGbc7c );
buf \U$37442 ( \44758 , \42121_nGbbbc );
buf \U$37443 ( \44759 , \42169_nGbbec );
buf \U$37444 ( \44760 , \42218_nGbc1c );
buf \U$37445 ( \44761 , \42267_nGbc4c );
or \U$37446 ( \44762 , \44758 , \44759 , \44760 , \44761 );
and \U$37447 ( \44763 , \44757 , \44762 );
buf \U$37448 ( \44764 , \44763 );
or \U$37449 ( \44765 , \44756 , \44764 );
_DC ge706 ( \44766_nGe706 , \44749 , \44765 );
buf \U$37450 ( \44767 , \44766_nGe706 );
_DC g1ade5_GF_IsGateDCbyConstraint ( \44768_nG1ade5 , \44767 , \42503 );
buf \U$37451 ( \44769 , \44768_nG1ade5 );
buf \U$37452 ( \44770 , RIe5d6d40_6768);
and \U$37453 ( \44771 , \44770 , \44701 );
buf \U$37454 ( \44772 , RIe5117a8_6369);
and \U$37455 ( \44773 , \44772 , \44704 );
buf \U$37456 ( \44774 , RIe444fb0_5975);
and \U$37457 ( \44775 , \44774 , \44708 );
buf \U$37458 ( \44776 , RIe37f9b8_5584);
and \U$37459 ( \44777 , \44776 , \44711 );
buf \U$37460 ( \44778 , RIe1ac2a0_5191);
and \U$37461 ( \44779 , \44778 , \44714 );
buf \U$37462 ( \44780 , RIe0e8ec8_4791);
and \U$37463 ( \44781 , \44780 , \44717 );
buf \U$37464 ( \44782 , RIe022a30_4393);
and \U$37465 ( \44783 , \44782 , \44720 );
buf \U$37466 ( \44784 , RIde4ec88_4006);
and \U$37467 ( \44785 , \44784 , \44723 );
buf \U$37468 ( \44786 , RIdd8ba30_3609);
and \U$37469 ( \44787 , \44786 , \44726 );
buf \U$37470 ( \44788 , RIdbc4870_3212);
and \U$37471 ( \44789 , \44788 , \44729 );
buf \U$37472 ( \44790 , RIdaf5f30_2820);
and \U$37473 ( \44791 , \44790 , \44732 );
buf \U$37474 ( \44792 , RIda25c28_2423);
and \U$37475 ( \44793 , \44792 , \44735 );
buf \U$37476 ( \44794 , RId96d278_2032);
and \U$37477 ( \44795 , \44794 , \44738 );
buf \U$37478 ( \44796 , RId8aa728_1632);
and \U$37479 ( \44797 , \44796 , \44741 );
buf \U$37480 ( \44798 , RId7dcb80_1235);
and \U$37481 ( \44799 , \44798 , \44744 );
buf \U$37482 ( \44800 , RId710748_846);
and \U$37483 ( \44801 , \44800 , \44747 );
or \U$37484 ( \44802 , \44771 , \44773 , \44775 , \44777 , \44779 , \44781 , \44783 , \44785 , \44787 , \44789 , \44791 , \44793 , \44795 , \44797 , \44799 , \44801 );
_DC ge728 ( \44803_nGe728 , \44802 , \44765 );
not \U$37485 ( \44804 , \44803_nGe728 );
_DC g1ac11_GF_IsGateDCbyConstraint ( \44805_nG1ac11 , \44804 , \42503 );
buf \U$37486 ( \44806 , \44805_nG1ac11 );
buf \U$37487 ( \44807 , RIb87eb00_69);
buf \U$37488 ( \44808 , RIe667bb0_6885);
buf \U$37489 ( \44809 , RIe667f70_6886);
nor \U$37490 ( \44810 , \44808 , \44809 );
_HMUX g17ab0 ( \44811_nG17ab0 , RIe3ac2b0_6083 , \44807 , \44810 );
and \U$37491 ( \44812 , RIea90778_6887, RIe546890_6849, RIe546098_6850, RIe545dc8_6851, \42389 );
buf \U$37492 ( \44813 , \44812 );
buf \U$37493 ( \44814 , \44813 );
buf \U$37494 ( \44815 , \42587 );
buf \U$37495 ( \44816 , \44815 );
and \U$37496 ( \44817 , \44814 , \44816 );
_HMUX g17ab1 ( \44818_nG17ab1 , RIe3ac2b0_6083 , \44811_nG17ab0 , \44817 );
buf \U$37497 ( \44819 , RIb7c5980_237);
buf \U$37498 ( \44820 , RIeab7058_6894);
buf \U$37499 ( \44821 , RIea91768_6889);
nor \U$37500 ( \44822 , \44820 , \44821 );
_HMUX g17ab3 ( \44823_nG17ab3 , RIe3ac2b0_6083 , \44819 , \44822 );
and \U$37501 ( \44824 , \42121_nGbbbc , \42169_nGbbec , \42218_nGbc1c , \42267_nGbc4c , \42316 );
buf \U$37502 ( \44825 , \44824 );
buf \U$37503 ( \44826 , \44825 );
buf \U$37504 ( \44827 , RIb79b518_270);
buf \U$37505 ( \44828 , \44827 );
and \U$37506 ( \44829 , \44826 , \44828 );
_HMUX g17ab4 ( \44830_nG17ab4 , \44818_nG17ab1 , \44823_nG17ab3 , \44829 );
buf \U$37507 ( \44831 , \44830_nG17ab4 );
_DC g1927e_GF_IsGateDCbyConstraint ( \44832_nG1927e , \44831 , \42503 );
buf \U$37508 ( \44833 , \44832_nG1927e );
buf \U$37509 ( \44834 , RIb87eb78_68);
_HMUX g17ab5 ( \44835_nG17ab5 , RIe3aaca8_6084 , \44834 , \44810 );
_HMUX g17ab6 ( \44836_nG17ab6 , RIe3aaca8_6084 , \44835_nG17ab5 , \44817 );
buf \U$37510 ( \44837 , RIb7c59f8_236);
_HMUX g17ab7 ( \44838_nG17ab7 , RIe3aaca8_6084 , \44837 , \44822 );
_HMUX g17ab8 ( \44839_nG17ab8 , \44836_nG17ab6 , \44838_nG17ab7 , \44829 );
buf \U$37511 ( \44840 , \44839_nG17ab8 );
_DC g19294_GF_IsGateDCbyConstraint ( \44841_nG19294 , \44840 , \42503 );
buf \U$37512 ( \44842 , \44841_nG19294 );
buf \U$37513 ( \44843 , RIb87ebf0_67);
_HMUX g17ab9 ( \44844_nG17ab9 , RIe3a9b50_6085 , \44843 , \44810 );
_HMUX g17aba ( \44845_nG17aba , RIe3a9b50_6085 , \44844_nG17ab9 , \44817 );
buf \U$37514 ( \44846 , RIb7c5a70_235);
_HMUX g17abb ( \44847_nG17abb , RIe3a9b50_6085 , \44846 , \44822 );
_HMUX g17abc ( \44848_nG17abc , \44845_nG17aba , \44847_nG17abb , \44829 );
buf \U$37515 ( \44849 , \44848_nG17abc );
_DC g192aa_GF_IsGateDCbyConstraint ( \44850_nG192aa , \44849 , \42503 );
buf \U$37516 ( \44851 , \44850_nG192aa );
buf \U$37517 ( \44852 , RIb882ca0_66);
_HMUX g17abd ( \44853_nG17abd , RIe3a8548_6086 , \44852 , \44810 );
_HMUX g17abe ( \44854_nG17abe , RIe3a8548_6086 , \44853_nG17abd , \44817 );
buf \U$37518 ( \44855 , RIb7cade0_234);
_HMUX g17abf ( \44856_nG17abf , RIe3a8548_6086 , \44855 , \44822 );
_HMUX g17ac0 ( \44857_nG17ac0 , \44854_nG17abe , \44856_nG17abf , \44829 );
buf \U$37519 ( \44858 , \44857_nG17ac0 );
_DC g192c0_GF_IsGateDCbyConstraint ( \44859_nG192c0 , \44858 , \42503 );
buf \U$37520 ( \44860 , \44859_nG192c0 );
buf \U$37521 ( \44861 , RIb885310_65);
_HMUX g17ac1 ( \44862_nG17ac1 , RIe3a73f0_6087 , \44861 , \44810 );
_HMUX g17ac2 ( \44863_nG17ac2 , RIe3a73f0_6087 , \44862_nG17ac1 , \44817 );
buf \U$37522 ( \44864 , RIb7cae58_233);
_HMUX g17ac3 ( \44865_nG17ac3 , RIe3a73f0_6087 , \44864 , \44822 );
_HMUX g17ac4 ( \44866_nG17ac4 , \44863_nG17ac2 , \44865_nG17ac3 , \44829 );
buf \U$37523 ( \44867 , \44866_nG17ac4 );
_DC g192d6_GF_IsGateDCbyConstraint ( \44868_nG192d6 , \44867 , \42503 );
buf \U$37524 ( \44869 , \44868_nG192d6 );
buf \U$37525 ( \44870 , RIb885388_64);
_HMUX g17ac5 ( \44871_nG17ac5 , RIe3a6298_6088 , \44870 , \44810 );
_HMUX g17ac6 ( \44872_nG17ac6 , RIe3a6298_6088 , \44871_nG17ac5 , \44817 );
buf \U$37526 ( \44873 , RIb7caed0_232);
_HMUX g17ac7 ( \44874_nG17ac7 , RIe3a6298_6088 , \44873 , \44822 );
_HMUX g17ac8 ( \44875_nG17ac8 , \44872_nG17ac6 , \44874_nG17ac7 , \44829 );
buf \U$37527 ( \44876 , \44875_nG17ac8 );
_DC g192ec_GF_IsGateDCbyConstraint ( \44877_nG192ec , \44876 , \42503 );
buf \U$37528 ( \44878 , \44877_nG192ec );
buf \U$37529 ( \44879 , RIb885400_63);
_HMUX g17ac9 ( \44880_nG17ac9 , RIe3a4c90_6089 , \44879 , \44810 );
_HMUX g17aca ( \44881_nG17aca , RIe3a4c90_6089 , \44880_nG17ac9 , \44817 );
buf \U$37530 ( \44882 , RIb7caf48_231);
_HMUX g17acb ( \44883_nG17acb , RIe3a4c90_6089 , \44882 , \44822 );
_HMUX g17acc ( \44884_nG17acc , \44881_nG17aca , \44883_nG17acb , \44829 );
buf \U$37531 ( \44885 , \44884_nG17acc );
_DC g192f8_GF_IsGateDCbyConstraint ( \44886_nG192f8 , \44885 , \42503 );
buf \U$37532 ( \44887 , \44886_nG192f8 );
buf \U$37533 ( \44888 , RIb885478_62);
_HMUX g17acd ( \44889_nG17acd , RIe3a3b38_6090 , \44888 , \44810 );
_HMUX g17ace ( \44890_nG17ace , RIe3a3b38_6090 , \44889_nG17acd , \44817 );
buf \U$37534 ( \44891 , RIb7cafc0_230);
_HMUX g17acf ( \44892_nG17acf , RIe3a3b38_6090 , \44891 , \44822 );
_HMUX g17ad0 ( \44893_nG17ad0 , \44890_nG17ace , \44892_nG17acf , \44829 );
buf \U$37535 ( \44894 , \44893_nG17ad0 );
_DC g192fa_GF_IsGateDCbyConstraint ( \44895_nG192fa , \44894 , \42503 );
buf \U$37536 ( \44896 , \44895_nG192fa );
buf \U$37537 ( \44897 , RIb8854f0_61);
_HMUX g17ad1 ( \44898_nG17ad1 , RIe3a2530_6091 , \44897 , \44810 );
_HMUX g17ad2 ( \44899_nG17ad2 , RIe3a2530_6091 , \44898_nG17ad1 , \44817 );
buf \U$37538 ( \44900 , RIb7cb038_229);
_HMUX g17ad3 ( \44901_nG17ad3 , RIe3a2530_6091 , \44900 , \44822 );
_HMUX g17ad4 ( \44902_nG17ad4 , \44899_nG17ad2 , \44901_nG17ad3 , \44829 );
buf \U$37539 ( \44903 , \44902_nG17ad4 );
_DC g192fc_GF_IsGateDCbyConstraint ( \44904_nG192fc , \44903 , \42503 );
buf \U$37540 ( \44905 , \44904_nG192fc );
buf \U$37541 ( \44906 , RIb885568_60);
_HMUX g17ad5 ( \44907_nG17ad5 , RIe3a13d8_6092 , \44906 , \44810 );
_HMUX g17ad6 ( \44908_nG17ad6 , RIe3a13d8_6092 , \44907_nG17ad5 , \44817 );
buf \U$37542 ( \44909 , RIb7cb0b0_228);
_HMUX g17ad7 ( \44910_nG17ad7 , RIe3a13d8_6092 , \44909 , \44822 );
_HMUX g17ad8 ( \44911_nG17ad8 , \44908_nG17ad6 , \44910_nG17ad7 , \44829 );
buf \U$37543 ( \44912 , \44911_nG17ad8 );
_DC g19280_GF_IsGateDCbyConstraint ( \44913_nG19280 , \44912 , \42503 );
buf \U$37544 ( \44914 , \44913_nG19280 );
buf \U$37545 ( \44915 , RIb8855e0_59);
_HMUX g17ad9 ( \44916_nG17ad9 , RIe39fdd0_6093 , \44915 , \44810 );
_HMUX g17ada ( \44917_nG17ada , RIe39fdd0_6093 , \44916_nG17ad9 , \44817 );
buf \U$37546 ( \44918 , RIb7cb128_227);
_HMUX g17adb ( \44919_nG17adb , RIe39fdd0_6093 , \44918 , \44822 );
_HMUX g17adc ( \44920_nG17adc , \44917_nG17ada , \44919_nG17adb , \44829 );
buf \U$37547 ( \44921 , \44920_nG17adc );
_DC g19282_GF_IsGateDCbyConstraint ( \44922_nG19282 , \44921 , \42503 );
buf \U$37548 ( \44923 , \44922_nG19282 );
buf \U$37549 ( \44924 , RIb885658_58);
_HMUX g17add ( \44925_nG17add , RIe39ec78_6094 , \44924 , \44810 );
_HMUX g17ade ( \44926_nG17ade , RIe39ec78_6094 , \44925_nG17add , \44817 );
buf \U$37550 ( \44927 , RIb7d00d8_226);
_HMUX g17adf ( \44928_nG17adf , RIe39ec78_6094 , \44927 , \44822 );
_HMUX g17ae0 ( \44929_nG17ae0 , \44926_nG17ade , \44928_nG17adf , \44829 );
buf \U$37551 ( \44930 , \44929_nG17ae0 );
_DC g19284_GF_IsGateDCbyConstraint ( \44931_nG19284 , \44930 , \42503 );
buf \U$37552 ( \44932 , \44931_nG19284 );
buf \U$37553 ( \44933 , RIb8856d0_57);
_HMUX g17ae1 ( \44934_nG17ae1 , RIe39db20_6095 , \44933 , \44810 );
_HMUX g17ae2 ( \44935_nG17ae2 , RIe39db20_6095 , \44934_nG17ae1 , \44817 );
buf \U$37554 ( \44936 , RIb8263d8_225);
_HMUX g17ae3 ( \44937_nG17ae3 , RIe39db20_6095 , \44936 , \44822 );
_HMUX g17ae4 ( \44938_nG17ae4 , \44935_nG17ae2 , \44937_nG17ae3 , \44829 );
buf \U$37555 ( \44939 , \44938_nG17ae4 );
_DC g19286_GF_IsGateDCbyConstraint ( \44940_nG19286 , \44939 , \42503 );
buf \U$37556 ( \44941 , \44940_nG19286 );
buf \U$37557 ( \44942 , RIb885748_56);
_HMUX g17ae5 ( \44943_nG17ae5 , RIe39c518_6096 , \44942 , \44810 );
_HMUX g17ae6 ( \44944_nG17ae6 , RIe39c518_6096 , \44943_nG17ae5 , \44817 );
buf \U$37558 ( \44945 , RIb826e28_224);
_HMUX g17ae7 ( \44946_nG17ae7 , RIe39c518_6096 , \44945 , \44822 );
_HMUX g17ae8 ( \44947_nG17ae8 , \44944_nG17ae6 , \44946_nG17ae7 , \44829 );
buf \U$37559 ( \44948 , \44947_nG17ae8 );
_DC g19288_GF_IsGateDCbyConstraint ( \44949_nG19288 , \44948 , \42503 );
buf \U$37560 ( \44950 , \44949_nG19288 );
buf \U$37561 ( \44951 , RIb8857c0_55);
_HMUX g17ae9 ( \44952_nG17ae9 , RIe1694d8_6097 , \44951 , \44810 );
_HMUX g17aea ( \44953_nG17aea , RIe1694d8_6097 , \44952_nG17ae9 , \44817 );
buf \U$37562 ( \44954 , RIb826ea0_223);
_HMUX g17aeb ( \44955_nG17aeb , RIe1694d8_6097 , \44954 , \44822 );
_HMUX g17aec ( \44956_nG17aec , \44953_nG17aea , \44955_nG17aeb , \44829 );
buf \U$37563 ( \44957 , \44956_nG17aec );
_DC g1928a_GF_IsGateDCbyConstraint ( \44958_nG1928a , \44957 , \42503 );
buf \U$37564 ( \44959 , \44958_nG1928a );
buf \U$37565 ( \44960 , RIb885838_54);
_HMUX g17aed ( \44961_nG17aed , RIe16e398_6098 , \44960 , \44810 );
_HMUX g17aee ( \44962_nG17aee , RIe16e398_6098 , \44961_nG17aed , \44817 );
buf \U$37566 ( \44963 , RIb826f18_222);
_HMUX g17aef ( \44964_nG17aef , RIe16e398_6098 , \44963 , \44822 );
_HMUX g17af0 ( \44965_nG17af0 , \44962_nG17aee , \44964_nG17aef , \44829 );
buf \U$37567 ( \44966 , \44965_nG17af0 );
_DC g1928c_GF_IsGateDCbyConstraint ( \44967_nG1928c , \44966 , \42503 );
buf \U$37568 ( \44968 , \44967_nG1928c );
buf \U$37569 ( \44969 , RIb8858b0_53);
_HMUX g17af1 ( \44970_nG17af1 , RIe173270_6099 , \44969 , \44810 );
_HMUX g17af2 ( \44971_nG17af2 , RIe173270_6099 , \44970_nG17af1 , \44817 );
buf \U$37570 ( \44972 , RIb826f90_221);
_HMUX g17af3 ( \44973_nG17af3 , RIe173270_6099 , \44972 , \44822 );
_HMUX g17af4 ( \44974_nG17af4 , \44971_nG17af2 , \44973_nG17af3 , \44829 );
buf \U$37571 ( \44975 , \44974_nG17af4 );
_DC g1928e_GF_IsGateDCbyConstraint ( \44976_nG1928e , \44975 , \42503 );
buf \U$37572 ( \44977 , \44976_nG1928e );
buf \U$37573 ( \44978 , RIb885928_52);
_HMUX g17af5 ( \44979_nG17af5 , RIe178388_6100 , \44978 , \44810 );
_HMUX g17af6 ( \44980_nG17af6 , RIe178388_6100 , \44979_nG17af5 , \44817 );
buf \U$37574 ( \44981 , RIb8293a8_220);
_HMUX g17af7 ( \44982_nG17af7 , RIe178388_6100 , \44981 , \44822 );
_HMUX g17af8 ( \44983_nG17af8 , \44980_nG17af6 , \44982_nG17af7 , \44829 );
buf \U$37575 ( \44984 , \44983_nG17af8 );
_DC g19290_GF_IsGateDCbyConstraint ( \44985_nG19290 , \44984 , \42503 );
buf \U$37576 ( \44986 , \44985_nG19290 );
buf \U$37577 ( \44987 , RIb8859a0_51);
_HMUX g17af9 ( \44988_nG17af9 , RIe17c780_6101 , \44987 , \44810 );
_HMUX g17afa ( \44989_nG17afa , RIe17c780_6101 , \44988_nG17af9 , \44817 );
buf \U$37578 ( \44990 , RIb829420_219);
_HMUX g17afb ( \44991_nG17afb , RIe17c780_6101 , \44990 , \44822 );
_HMUX g17afc ( \44992_nG17afc , \44989_nG17afa , \44991_nG17afb , \44829 );
buf \U$37579 ( \44993 , \44992_nG17afc );
_DC g19292_GF_IsGateDCbyConstraint ( \44994_nG19292 , \44993 , \42503 );
buf \U$37580 ( \44995 , \44994_nG19292 );
buf \U$37581 ( \44996 , RIb885a18_50);
_HMUX g17afd ( \44997_nG17afd , RIe1805d8_6102 , \44996 , \44810 );
_HMUX g17afe ( \44998_nG17afe , RIe1805d8_6102 , \44997_nG17afd , \44817 );
buf \U$37582 ( \44999 , RIb829498_218);
_HMUX g17aff ( \45000_nG17aff , RIe1805d8_6102 , \44999 , \44822 );
_HMUX g17b00 ( \45001_nG17b00 , \44998_nG17afe , \45000_nG17aff , \44829 );
buf \U$37583 ( \45002 , \45001_nG17b00 );
_DC g19296_GF_IsGateDCbyConstraint ( \45003_nG19296 , \45002 , \42503 );
buf \U$37584 ( \45004 , \45003_nG19296 );
buf \U$37585 ( \45005 , RIb885a90_49);
_HMUX g17b01 ( \45006_nG17b01 , RIe1877c0_6103 , \45005 , \44810 );
_HMUX g17b02 ( \45007_nG17b02 , RIe1877c0_6103 , \45006_nG17b01 , \44817 );
buf \U$37586 ( \45008 , RIb829510_217);
_HMUX g17b03 ( \45009_nG17b03 , RIe1877c0_6103 , \45008 , \44822 );
_HMUX g17b04 ( \45010_nG17b04 , \45007_nG17b02 , \45009_nG17b03 , \44829 );
buf \U$37587 ( \45011 , \45010_nG17b04 );
_DC g19298_GF_IsGateDCbyConstraint ( \45012_nG19298 , \45011 , \42503 );
buf \U$37588 ( \45013 , \45012_nG19298 );
buf \U$37589 ( \45014 , RIb885b08_48);
_HMUX g17b05 ( \45015_nG17b05 , RIe18c9c8_6104 , \45014 , \44810 );
_HMUX g17b06 ( \45016_nG17b06 , RIe18c9c8_6104 , \45015_nG17b05 , \44817 );
buf \U$37590 ( \45017 , RIb829588_216);
_HMUX g17b07 ( \45018_nG17b07 , RIe18c9c8_6104 , \45017 , \44822 );
_HMUX g17b08 ( \45019_nG17b08 , \45016_nG17b06 , \45018_nG17b07 , \44829 );
buf \U$37591 ( \45020 , \45019_nG17b08 );
_DC g1929a_GF_IsGateDCbyConstraint ( \45021_nG1929a , \45020 , \42503 );
buf \U$37592 ( \45022 , \45021_nG1929a );
buf \U$37593 ( \45023 , RIb885b80_47);
_HMUX g17b09 ( \45024_nG17b09 , RIe192ff8_6105 , \45023 , \44810 );
_HMUX g17b0a ( \45025_nG17b0a , RIe192ff8_6105 , \45024_nG17b09 , \44817 );
buf \U$37594 ( \45026 , RIb829600_215);
_HMUX g17b0b ( \45027_nG17b0b , RIe192ff8_6105 , \45026 , \44822 );
_HMUX g17b0c ( \45028_nG17b0c , \45025_nG17b0a , \45027_nG17b0b , \44829 );
buf \U$37595 ( \45029 , \45028_nG17b0c );
_DC g1929c_GF_IsGateDCbyConstraint ( \45030_nG1929c , \45029 , \42503 );
buf \U$37596 ( \45031 , \45030_nG1929c );
buf \U$37597 ( \45032 , RIb885bf8_46);
_HMUX g17b0d ( \45033_nG17b0d , RIe198cc8_6106 , \45032 , \44810 );
_HMUX g17b0e ( \45034_nG17b0e , RIe198cc8_6106 , \45033_nG17b0d , \44817 );
buf \U$37598 ( \45035 , RIb829678_214);
_HMUX g17b0f ( \45036_nG17b0f , RIe198cc8_6106 , \45035 , \44822 );
_HMUX g17b10 ( \45037_nG17b10 , \45034_nG17b0e , \45036_nG17b0f , \44829 );
buf \U$37599 ( \45038 , \45037_nG17b10 );
_DC g1929e_GF_IsGateDCbyConstraint ( \45039_nG1929e , \45038 , \42503 );
buf \U$37600 ( \45040 , \45039_nG1929e );
buf \U$37601 ( \45041 , RIb885c70_45);
_HMUX g17b11 ( \45042_nG17b11 , RIe1a05b8_6107 , \45041 , \44810 );
_HMUX g17b12 ( \45043_nG17b12 , RIe1a05b8_6107 , \45042_nG17b11 , \44817 );
buf \U$37602 ( \45044 , RIb8296f0_213);
_HMUX g17b13 ( \45045_nG17b13 , RIe1a05b8_6107 , \45044 , \44822 );
_HMUX g17b14 ( \45046_nG17b14 , \45043_nG17b12 , \45045_nG17b13 , \44829 );
buf \U$37603 ( \45047 , \45046_nG17b14 );
_DC g192a0_GF_IsGateDCbyConstraint ( \45048_nG192a0 , \45047 , \42503 );
buf \U$37604 ( \45049 , \45048_nG192a0 );
buf \U$37605 ( \45050 , RIb885ce8_44);
_HMUX g17b15 ( \45051_nG17b15 , RIe1a6300_6108 , \45050 , \44810 );
_HMUX g17b16 ( \45052_nG17b16 , RIe1a6300_6108 , \45051_nG17b15 , \44817 );
buf \U$37606 ( \45053 , RIb82dae8_212);
_HMUX g17b17 ( \45054_nG17b17 , RIe1a6300_6108 , \45053 , \44822 );
_HMUX g17b18 ( \45055_nG17b18 , \45052_nG17b16 , \45054_nG17b17 , \44829 );
buf \U$37607 ( \45056 , \45055_nG17b18 );
_DC g192a2_GF_IsGateDCbyConstraint ( \45057_nG192a2 , \45056 , \42503 );
buf \U$37608 ( \45058 , \45057_nG192a2 );
buf \U$37609 ( \45059 , RIb885d60_43);
_HMUX g17b19 ( \45060_nG17b19 , RIe1ac318_6109 , \45059 , \44810 );
_HMUX g17b1a ( \45061_nG17b1a , RIe1ac318_6109 , \45060_nG17b19 , \44817 );
buf \U$37610 ( \45062 , RIb82db60_211);
_HMUX g17b1b ( \45063_nG17b1b , RIe1ac318_6109 , \45062 , \44822 );
_HMUX g17b1c ( \45064_nG17b1c , \45061_nG17b1a , \45063_nG17b1b , \44829 );
buf \U$37611 ( \45065 , \45064_nG17b1c );
_DC g192a4_GF_IsGateDCbyConstraint ( \45066_nG192a4 , \45065 , \42503 );
buf \U$37612 ( \45067 , \45066_nG192a4 );
buf \U$37613 ( \45068 , RIb885dd8_42);
_HMUX g17b1d ( \45069_nG17b1d , RIe1b2420_6110 , \45068 , \44810 );
_HMUX g17b1e ( \45070_nG17b1e , RIe1b2420_6110 , \45069_nG17b1d , \44817 );
buf \U$37614 ( \45071 , RIb82dbd8_210);
_HMUX g17b1f ( \45072_nG17b1f , RIe1b2420_6110 , \45071 , \44822 );
_HMUX g17b20 ( \45073_nG17b20 , \45070_nG17b1e , \45072_nG17b1f , \44829 );
buf \U$37615 ( \45074 , \45073_nG17b20 );
_DC g192a6_GF_IsGateDCbyConstraint ( \45075_nG192a6 , \45074 , \42503 );
buf \U$37616 ( \45076 , \45075_nG192a6 );
buf \U$37617 ( \45077 , RIb885e50_41);
_HMUX g17b21 ( \45078_nG17b21 , RIe1b7970_6111 , \45077 , \44810 );
_HMUX g17b22 ( \45079_nG17b22 , RIe1b7970_6111 , \45078_nG17b21 , \44817 );
buf \U$37618 ( \45080 , RIb82dc50_209);
_HMUX g17b23 ( \45081_nG17b23 , RIe1b7970_6111 , \45080 , \44822 );
_HMUX g17b24 ( \45082_nG17b24 , \45079_nG17b22 , \45081_nG17b23 , \44829 );
buf \U$37619 ( \45083 , \45082_nG17b24 );
_DC g192a8_GF_IsGateDCbyConstraint ( \45084_nG192a8 , \45083 , \42503 );
buf \U$37620 ( \45085 , \45084_nG192a8 );
buf \U$37621 ( \45086 , RIb885ec8_40);
_HMUX g17b25 ( \45087_nG17b25 , RIe1bce48_6112 , \45086 , \44810 );
_HMUX g17b26 ( \45088_nG17b26 , RIe1bce48_6112 , \45087_nG17b25 , \44817 );
buf \U$37622 ( \45089 , RIb82dcc8_208);
_HMUX g17b27 ( \45090_nG17b27 , RIe1bce48_6112 , \45089 , \44822 );
_HMUX g17b28 ( \45091_nG17b28 , \45088_nG17b26 , \45090_nG17b27 , \44829 );
buf \U$37623 ( \45092 , \45091_nG17b28 );
_DC g192ac_GF_IsGateDCbyConstraint ( \45093_nG192ac , \45092 , \42503 );
buf \U$37624 ( \45094 , \45093_nG192ac );
buf \U$37625 ( \45095 , RIb885f40_39);
_HMUX g17b29 ( \45096_nG17b29 , RIe1c12b8_6113 , \45095 , \44810 );
_HMUX g17b2a ( \45097_nG17b2a , RIe1c12b8_6113 , \45096_nG17b29 , \44817 );
buf \U$37626 ( \45098 , RIb82dd40_207);
_HMUX g17b2b ( \45099_nG17b2b , RIe1c12b8_6113 , \45098 , \44822 );
_HMUX g17b2c ( \45100_nG17b2c , \45097_nG17b2a , \45099_nG17b2b , \44829 );
buf \U$37627 ( \45101 , \45100_nG17b2c );
_DC g192ae_GF_IsGateDCbyConstraint ( \45102_nG192ae , \45101 , \42503 );
buf \U$37628 ( \45103 , \45102_nG192ae );
buf \U$37629 ( \45104 , RIb885fb8_38);
_HMUX g17b2d ( \45105_nG17b2d , RIe1c7960_6114 , \45104 , \44810 );
_HMUX g17b2e ( \45106_nG17b2e , RIe1c7960_6114 , \45105_nG17b2d , \44817 );
buf \U$37630 ( \45107 , RIb82ddb8_206);
_HMUX g17b2f ( \45108_nG17b2f , RIe1c7960_6114 , \45107 , \44822 );
_HMUX g17b30 ( \45109_nG17b30 , \45106_nG17b2e , \45108_nG17b2f , \44829 );
buf \U$37631 ( \45110 , \45109_nG17b30 );
_DC g192b0_GF_IsGateDCbyConstraint ( \45111_nG192b0 , \45110 , \42503 );
buf \U$37632 ( \45112 , \45111_nG192b0 );
buf \U$37633 ( \45113 , RIb886030_37);
_HMUX g17b31 ( \45114_nG17b31 , RIe1cc820_6115 , \45113 , \44810 );
_HMUX g17b32 ( \45115_nG17b32 , RIe1cc820_6115 , \45114_nG17b31 , \44817 );
buf \U$37634 ( \45116 , RIb82de30_205);
_HMUX g17b33 ( \45117_nG17b33 , RIe1cc820_6115 , \45116 , \44822 );
_HMUX g17b34 ( \45118_nG17b34 , \45115_nG17b32 , \45117_nG17b33 , \44829 );
buf \U$37635 ( \45119 , \45118_nG17b34 );
_DC g192b2_GF_IsGateDCbyConstraint ( \45120_nG192b2 , \45119 , \42503 );
buf \U$37636 ( \45121 , \45120_nG192b2 );
buf \U$37637 ( \45122 , RIb8860a8_36);
_HMUX g17b35 ( \45123_nG17b35 , RIe1d0fd8_6116 , \45122 , \44810 );
_HMUX g17b36 ( \45124_nG17b36 , RIe1d0fd8_6116 , \45123_nG17b35 , \44817 );
buf \U$37638 ( \45125 , RIb832228_204);
_HMUX g17b37 ( \45126_nG17b37 , RIe1d0fd8_6116 , \45125 , \44822 );
_HMUX g17b38 ( \45127_nG17b38 , \45124_nG17b36 , \45126_nG17b37 , \44829 );
buf \U$37639 ( \45128 , \45127_nG17b38 );
_DC g192b4_GF_IsGateDCbyConstraint ( \45129_nG192b4 , \45128 , \42503 );
buf \U$37640 ( \45130 , \45129_nG192b4 );
buf \U$37641 ( \45131 , RIb886120_35);
_HMUX g17b39 ( \45132_nG17b39 , RIe094940_6117 , \45131 , \44810 );
_HMUX g17b3a ( \45133_nG17b3a , RIe094940_6117 , \45132_nG17b39 , \44817 );
buf \U$37642 ( \45134 , RIb8322a0_203);
_HMUX g17b3b ( \45135_nG17b3b , RIe094940_6117 , \45134 , \44822 );
_HMUX g17b3c ( \45136_nG17b3c , \45133_nG17b3a , \45135_nG17b3b , \44829 );
buf \U$37643 ( \45137 , \45136_nG17b3c );
_DC g192b6_GF_IsGateDCbyConstraint ( \45138_nG192b6 , \45137 , \42503 );
buf \U$37644 ( \45139 , \45138_nG192b6 );
buf \U$37645 ( \45140 , RIb886198_34);
_HMUX g17b3d ( \45141_nG17b3d , RIe090368_6118 , \45140 , \44810 );
_HMUX g17b3e ( \45142_nG17b3e , RIe090368_6118 , \45141_nG17b3d , \44817 );
buf \U$37646 ( \45143 , RIb832318_202);
_HMUX g17b3f ( \45144_nG17b3f , RIe090368_6118 , \45143 , \44822 );
_HMUX g17b40 ( \45145_nG17b40 , \45142_nG17b3e , \45144_nG17b3f , \44829 );
buf \U$37647 ( \45146 , \45145_nG17b40 );
_DC g192b8_GF_IsGateDCbyConstraint ( \45147_nG192b8 , \45146 , \42503 );
buf \U$37648 ( \45148 , \45147_nG192b8 );
buf \U$37649 ( \45149 , RIb886210_33);
_HMUX g17b41 ( \45150_nG17b41 , RIe08b700_6119 , \45149 , \44810 );
_HMUX g17b42 ( \45151_nG17b42 , RIe08b700_6119 , \45150_nG17b41 , \44817 );
buf \U$37650 ( \45152 , RIb832390_201);
_HMUX g17b43 ( \45153_nG17b43 , RIe08b700_6119 , \45152 , \44822 );
_HMUX g17b44 ( \45154_nG17b44 , \45151_nG17b42 , \45153_nG17b43 , \44829 );
buf \U$37651 ( \45155 , \45154_nG17b44 );
_DC g192ba_GF_IsGateDCbyConstraint ( \45156_nG192ba , \45155 , \42503 );
buf \U$37652 ( \45157 , \45156_nG192ba );
buf \U$37653 ( \45158 , RIb886288_32);
_HMUX g17b45 ( \45159_nG17b45 , RIe087a10_6120 , \45158 , \44810 );
_HMUX g17b46 ( \45160_nG17b46 , RIe087a10_6120 , \45159_nG17b45 , \44817 );
buf \U$37654 ( \45161 , RIb832408_200);
_HMUX g17b47 ( \45162_nG17b47 , RIe087a10_6120 , \45161 , \44822 );
_HMUX g17b48 ( \45163_nG17b48 , \45160_nG17b46 , \45162_nG17b47 , \44829 );
buf \U$37655 ( \45164 , \45163_nG17b48 );
_DC g192bc_GF_IsGateDCbyConstraint ( \45165_nG192bc , \45164 , \42503 );
buf \U$37656 ( \45166 , \45165_nG192bc );
buf \U$37657 ( \45167 , RIb886300_31);
_HMUX g17b49 ( \45168_nG17b49 , RIe14c9f0_6121 , \45167 , \44810 );
_HMUX g17b4a ( \45169_nG17b4a , RIe14c9f0_6121 , \45168_nG17b49 , \44817 );
buf \U$37658 ( \45170 , RIb832480_199);
_HMUX g17b4b ( \45171_nG17b4b , RIe14c9f0_6121 , \45170 , \44822 );
_HMUX g17b4c ( \45172_nG17b4c , \45169_nG17b4a , \45171_nG17b4b , \44829 );
buf \U$37659 ( \45173 , \45172_nG17b4c );
_DC g192be_GF_IsGateDCbyConstraint ( \45174_nG192be , \45173 , \42503 );
buf \U$37660 ( \45175 , \45174_nG192be );
buf \U$37661 ( \45176 , RIb886378_30);
_HMUX g17b4d ( \45177_nG17b4d , RIe1495e8_6122 , \45176 , \44810 );
_HMUX g17b4e ( \45178_nG17b4e , RIe1495e8_6122 , \45177_nG17b4d , \44817 );
buf \U$37662 ( \45179 , RIb8324f8_198);
_HMUX g17b4f ( \45180_nG17b4f , RIe1495e8_6122 , \45179 , \44822 );
_HMUX g17b50 ( \45181_nG17b50 , \45178_nG17b4e , \45180_nG17b4f , \44829 );
buf \U$37663 ( \45182 , \45181_nG17b50 );
_DC g192c2_GF_IsGateDCbyConstraint ( \45183_nG192c2 , \45182 , \42503 );
buf \U$37664 ( \45184 , \45183_nG192c2 );
buf \U$37665 ( \45185 , RIb8863f0_29);
_HMUX g17b51 ( \45186_nG17b51 , RIe146348_6123 , \45185 , \44810 );
_HMUX g17b52 ( \45187_nG17b52 , RIe146348_6123 , \45186_nG17b51 , \44817 );
buf \U$37666 ( \45188 , RIb832570_197);
_HMUX g17b53 ( \45189_nG17b53 , RIe146348_6123 , \45188 , \44822 );
_HMUX g17b54 ( \45190_nG17b54 , \45187_nG17b52 , \45189_nG17b53 , \44829 );
buf \U$37667 ( \45191 , \45190_nG17b54 );
_DC g192c4_GF_IsGateDCbyConstraint ( \45192_nG192c4 , \45191 , \42503 );
buf \U$37668 ( \45193 , \45192_nG192c4 );
buf \U$37669 ( \45194 , RIb886468_28);
_HMUX g17b55 ( \45195_nG17b55 , RIe143210_6124 , \45194 , \44810 );
_HMUX g17b56 ( \45196_nG17b56 , RIe143210_6124 , \45195_nG17b55 , \44817 );
buf \U$37670 ( \45197 , RIb8383a8_196);
_HMUX g17b57 ( \45198_nG17b57 , RIe143210_6124 , \45197 , \44822 );
_HMUX g17b58 ( \45199_nG17b58 , \45196_nG17b56 , \45198_nG17b57 , \44829 );
buf \U$37671 ( \45200 , \45199_nG17b58 );
_DC g192c6_GF_IsGateDCbyConstraint ( \45201_nG192c6 , \45200 , \42503 );
buf \U$37672 ( \45202 , \45201_nG192c6 );
buf \U$37673 ( \45203 , RIb8864e0_27);
_HMUX g17b59 ( \45204_nG17b59 , RIe140a38_6125 , \45203 , \44810 );
_HMUX g17b5a ( \45205_nG17b5a , RIe140a38_6125 , \45204_nG17b59 , \44817 );
buf \U$37674 ( \45206 , RIb838420_195);
_HMUX g17b5b ( \45207_nG17b5b , RIe140a38_6125 , \45206 , \44822 );
_HMUX g17b5c ( \45208_nG17b5c , \45205_nG17b5a , \45207_nG17b5b , \44829 );
buf \U$37675 ( \45209 , \45208_nG17b5c );
_DC g192c8_GF_IsGateDCbyConstraint ( \45210_nG192c8 , \45209 , \42503 );
buf \U$37676 ( \45211 , \45210_nG192c8 );
buf \U$37677 ( \45212 , RIb886558_26);
_HMUX g17b5d ( \45213_nG17b5d , RIe13d4c8_6126 , \45212 , \44810 );
_HMUX g17b5e ( \45214_nG17b5e , RIe13d4c8_6126 , \45213_nG17b5d , \44817 );
buf \U$37678 ( \45215 , RIb838498_194);
_HMUX g17b5f ( \45216_nG17b5f , RIe13d4c8_6126 , \45215 , \44822 );
_HMUX g17b60 ( \45217_nG17b60 , \45214_nG17b5e , \45216_nG17b5f , \44829 );
buf \U$37679 ( \45218 , \45217_nG17b60 );
_DC g192ca_GF_IsGateDCbyConstraint ( \45219_nG192ca , \45218 , \42503 );
buf \U$37680 ( \45220 , \45219_nG192ca );
buf \U$37681 ( \45221 , RIb8865d0_25);
_HMUX g17b61 ( \45222_nG17b61 , RIe13a660_6127 , \45221 , \44810 );
_HMUX g17b62 ( \45223_nG17b62 , RIe13a660_6127 , \45222_nG17b61 , \44817 );
buf \U$37682 ( \45224 , RIb838510_193);
_HMUX g17b63 ( \45225_nG17b63 , RIe13a660_6127 , \45224 , \44822 );
_HMUX g17b64 ( \45226_nG17b64 , \45223_nG17b62 , \45225_nG17b63 , \44829 );
buf \U$37683 ( \45227 , \45226_nG17b64 );
_DC g192cc_GF_IsGateDCbyConstraint ( \45228_nG192cc , \45227 , \42503 );
buf \U$37684 ( \45229 , \45228_nG192cc );
buf \U$37685 ( \45230 , RIb886648_24);
_HMUX g17b65 ( \45231_nG17b65 , RIe137168_6128 , \45230 , \44810 );
_HMUX g17b66 ( \45232_nG17b66 , RIe137168_6128 , \45231_nG17b65 , \44817 );
buf \U$37686 ( \45233 , RIb838588_192);
_HMUX g17b67 ( \45234_nG17b67 , RIe137168_6128 , \45233 , \44822 );
_HMUX g17b68 ( \45235_nG17b68 , \45232_nG17b66 , \45234_nG17b67 , \44829 );
buf \U$37687 ( \45236 , \45235_nG17b68 );
_DC g192ce_GF_IsGateDCbyConstraint ( \45237_nG192ce , \45236 , \42503 );
buf \U$37688 ( \45238 , \45237_nG192ce );
buf \U$37689 ( \45239 , RIb8866c0_23);
_HMUX g17b69 ( \45240_nG17b69 , RIe133a18_6129 , \45239 , \44810 );
_HMUX g17b6a ( \45241_nG17b6a , RIe133a18_6129 , \45240_nG17b69 , \44817 );
buf \U$37690 ( \45242 , RIb838600_191);
_HMUX g17b6b ( \45243_nG17b6b , RIe133a18_6129 , \45242 , \44822 );
_HMUX g17b6c ( \45244_nG17b6c , \45241_nG17b6a , \45243_nG17b6b , \44829 );
buf \U$37691 ( \45245 , \45244_nG17b6c );
_DC g192d0_GF_IsGateDCbyConstraint ( \45246_nG192d0 , \45245 , \42503 );
buf \U$37692 ( \45247 , \45246_nG192d0 );
buf \U$37693 ( \45248 , RIb886738_22);
_HMUX g17b6d ( \45249_nG17b6d , RIe12fda0_6130 , \45248 , \44810 );
_HMUX g17b6e ( \45250_nG17b6e , RIe12fda0_6130 , \45249_nG17b6d , \44817 );
buf \U$37694 ( \45251 , RIb838678_190);
_HMUX g17b6f ( \45252_nG17b6f , RIe12fda0_6130 , \45251 , \44822 );
_HMUX g17b70 ( \45253_nG17b70 , \45250_nG17b6e , \45252_nG17b6f , \44829 );
buf \U$37695 ( \45254 , \45253_nG17b70 );
_DC g192d2_GF_IsGateDCbyConstraint ( \45255_nG192d2 , \45254 , \42503 );
buf \U$37696 ( \45256 , \45255_nG192d2 );
buf \U$37697 ( \45257 , RIb8867b0_21);
_HMUX g17b71 ( \45258_nG17b71 , RIe1280f0_6131 , \45257 , \44810 );
_HMUX g17b72 ( \45259_nG17b72 , RIe1280f0_6131 , \45258_nG17b71 , \44817 );
buf \U$37698 ( \45260 , RIb8386f0_189);
_HMUX g17b73 ( \45261_nG17b73 , RIe1280f0_6131 , \45260 , \44822 );
_HMUX g17b74 ( \45262_nG17b74 , \45259_nG17b72 , \45261_nG17b73 , \44829 );
buf \U$37699 ( \45263 , \45262_nG17b74 );
_DC g192d4_GF_IsGateDCbyConstraint ( \45264_nG192d4 , \45263 , \42503 );
buf \U$37700 ( \45265 , \45264_nG192d4 );
buf \U$37701 ( \45266 , RIb886828_20);
_HMUX g17b75 ( \45267_nG17b75 , RIe121b38_6132 , \45266 , \44810 );
_HMUX g17b76 ( \45268_nG17b76 , RIe121b38_6132 , \45267_nG17b75 , \44817 );
buf \U$37702 ( \45269 , RIb838768_188);
_HMUX g17b77 ( \45270_nG17b77 , RIe121b38_6132 , \45269 , \44822 );
_HMUX g17b78 ( \45271_nG17b78 , \45268_nG17b76 , \45270_nG17b77 , \44829 );
buf \U$37703 ( \45272 , \45271_nG17b78 );
_DC g192d8_GF_IsGateDCbyConstraint ( \45273_nG192d8 , \45272 , \42503 );
buf \U$37704 ( \45274 , \45273_nG192d8 );
buf \U$37705 ( \45275 , RIb8868a0_19);
_HMUX g17b79 ( \45276_nG17b79 , RIe1194b0_6133 , \45275 , \44810 );
_HMUX g17b7a ( \45277_nG17b7a , RIe1194b0_6133 , \45276_nG17b79 , \44817 );
buf \U$37706 ( \45278 , RIb8387e0_187);
_HMUX g17b7b ( \45279_nG17b7b , RIe1194b0_6133 , \45278 , \44822 );
_HMUX g17b7c ( \45280_nG17b7c , \45277_nG17b7a , \45279_nG17b7b , \44829 );
buf \U$37707 ( \45281 , \45280_nG17b7c );
_DC g192da_GF_IsGateDCbyConstraint ( \45282_nG192da , \45281 , \42503 );
buf \U$37708 ( \45283 , \45282_nG192da );
buf \U$37709 ( \45284 , RIb886918_18);
_HMUX g17b7d ( \45285_nG17b7d , RIe1133a8_6134 , \45284 , \44810 );
_HMUX g17b7e ( \45286_nG17b7e , RIe1133a8_6134 , \45285_nG17b7d , \44817 );
buf \U$37710 ( \45287 , RIb838858_186);
_HMUX g17b7f ( \45288_nG17b7f , RIe1133a8_6134 , \45287 , \44822 );
_HMUX g17b80 ( \45289_nG17b80 , \45286_nG17b7e , \45288_nG17b7f , \44829 );
buf \U$37711 ( \45290 , \45289_nG17b80 );
_DC g192dc_GF_IsGateDCbyConstraint ( \45291_nG192dc , \45290 , \42503 );
buf \U$37712 ( \45292 , \45291_nG192dc );
buf \U$37713 ( \45293 , RIb886990_17);
_HMUX g17b81 ( \45294_nG17b81 , RIe10ad20_6135 , \45293 , \44810 );
_HMUX g17b82 ( \45295_nG17b82 , RIe10ad20_6135 , \45294_nG17b81 , \44817 );
buf \U$37714 ( \45296 , RIb8388d0_185);
_HMUX g17b83 ( \45297_nG17b83 , RIe10ad20_6135 , \45296 , \44822 );
_HMUX g17b84 ( \45298_nG17b84 , \45295_nG17b82 , \45297_nG17b83 , \44829 );
buf \U$37715 ( \45299 , \45298_nG17b84 );
_DC g192de_GF_IsGateDCbyConstraint ( \45300_nG192de , \45299 , \42503 );
buf \U$37716 ( \45301 , \45300_nG192de );
buf \U$37717 ( \45302 , RIb886a08_16);
_HMUX g17b85 ( \45303_nG17b85 , RIdfd70d0_6136 , \45302 , \44810 );
_HMUX g17b86 ( \45304_nG17b86 , RIdfd70d0_6136 , \45303_nG17b85 , \44817 );
buf \U$37718 ( \45305 , RIb838948_184);
_HMUX g17b87 ( \45306_nG17b87 , RIdfd70d0_6136 , \45305 , \44822 );
_HMUX g17b88 ( \45307_nG17b88 , \45304_nG17b86 , \45306_nG17b87 , \44829 );
buf \U$37719 ( \45308 , \45307_nG17b88 );
_DC g192e0_GF_IsGateDCbyConstraint ( \45309_nG192e0 , \45308 , \42503 );
buf \U$37720 ( \45310 , \45309_nG192e0 );
buf \U$37721 ( \45311 , RIb886a80_15);
_HMUX g17b89 ( \45312_nG17b89 , RIdff52b0_6137 , \45311 , \44810 );
_HMUX g17b8a ( \45313_nG17b8a , RIdff52b0_6137 , \45312_nG17b89 , \44817 );
buf \U$37722 ( \45314 , RIb8389c0_183);
_HMUX g17b8b ( \45315_nG17b8b , RIdff52b0_6137 , \45314 , \44822 );
_HMUX g17b8c ( \45316_nG17b8c , \45313_nG17b8a , \45315_nG17b8b , \44829 );
buf \U$37723 ( \45317 , \45316_nG17b8c );
_DC g192e2_GF_IsGateDCbyConstraint ( \45318_nG192e2 , \45317 , \42503 );
buf \U$37724 ( \45319 , \45318_nG192e2 );
buf \U$37725 ( \45320 , RIb886af8_14);
_HMUX g17b8d ( \45321_nG17b8d , RIe01ea70_6138 , \45320 , \44810 );
_HMUX g17b8e ( \45322_nG17b8e , RIe01ea70_6138 , \45321_nG17b8d , \44817 );
buf \U$37726 ( \45323 , RIb838a38_182);
_HMUX g17b8f ( \45324_nG17b8f , RIe01ea70_6138 , \45323 , \44822 );
_HMUX g17b90 ( \45325_nG17b90 , \45322_nG17b8e , \45324_nG17b8f , \44829 );
buf \U$37727 ( \45326 , \45325_nG17b90 );
_DC g192e4_GF_IsGateDCbyConstraint ( \45327_nG192e4 , \45326 , \42503 );
buf \U$37728 ( \45328 , \45327_nG192e4 );
buf \U$37729 ( \45329 , RIb886b70_13);
_HMUX g17b91 ( \45330_nG17b91 , RIe03a5e0_6139 , \45329 , \44810 );
_HMUX g17b92 ( \45331_nG17b92 , RIe03a5e0_6139 , \45330_nG17b91 , \44817 );
buf \U$37730 ( \45332 , RIb838ab0_181);
_HMUX g17b93 ( \45333_nG17b93 , RIe03a5e0_6139 , \45332 , \44822 );
_HMUX g17b94 ( \45334_nG17b94 , \45331_nG17b92 , \45333_nG17b93 , \44829 );
buf \U$37731 ( \45335 , \45334_nG17b94 );
_DC g192e6_GF_IsGateDCbyConstraint ( \45336_nG192e6 , \45335 , \42503 );
buf \U$37732 ( \45337 , \45336_nG192e6 );
buf \U$37733 ( \45338 , RIb886be8_12);
_HMUX g17b95 ( \45339_nG17b95 , RIdfb6cb8_6140 , \45338 , \44810 );
_HMUX g17b96 ( \45340_nG17b96 , RIdfb6cb8_6140 , \45339_nG17b95 , \44817 );
buf \U$37734 ( \45341 , RIb838b28_180);
_HMUX g17b97 ( \45342_nG17b97 , RIdfb6cb8_6140 , \45341 , \44822 );
_HMUX g17b98 ( \45343_nG17b98 , \45340_nG17b96 , \45342_nG17b97 , \44829 );
buf \U$37735 ( \45344 , \45343_nG17b98 );
_DC g192e8_GF_IsGateDCbyConstraint ( \45345_nG192e8 , \45344 , \42503 );
buf \U$37736 ( \45346 , \45345_nG192e8 );
buf \U$37737 ( \45347 , RIb886c60_11);
_HMUX g17b99 ( \45348_nG17b99 , RIdfa46d0_6141 , \45347 , \44810 );
_HMUX g17b9a ( \45349_nG17b9a , RIdfa46d0_6141 , \45348_nG17b99 , \44817 );
buf \U$37738 ( \45350 , RIb838ba0_179);
_HMUX g17b9b ( \45351_nG17b9b , RIdfa46d0_6141 , \45350 , \44822 );
_HMUX g17b9c ( \45352_nG17b9c , \45349_nG17b9a , \45351_nG17b9b , \44829 );
buf \U$37739 ( \45353 , \45352_nG17b9c );
_DC g192ea_GF_IsGateDCbyConstraint ( \45354_nG192ea , \45353 , \42503 );
buf \U$37740 ( \45355 , \45354_nG192ea );
buf \U$37741 ( \45356 , RIb886cd8_10);
_HMUX g17b9d ( \45357_nG17b9d , RIdf7c7e8_6142 , \45356 , \44810 );
_HMUX g17b9e ( \45358_nG17b9e , RIdf7c7e8_6142 , \45357_nG17b9d , \44817 );
buf \U$37742 ( \45359 , RIb838c18_178);
_HMUX g17b9f ( \45360_nG17b9f , RIdf7c7e8_6142 , \45359 , \44822 );
_HMUX g17ba0 ( \45361_nG17ba0 , \45358_nG17b9e , \45360_nG17b9f , \44829 );
buf \U$37743 ( \45362 , \45361_nG17ba0 );
_DC g192ee_GF_IsGateDCbyConstraint ( \45363_nG192ee , \45362 , \42503 );
buf \U$37744 ( \45364 , \45363_nG192ee );
buf \U$37745 ( \45365 , RIb886d50_9);
_HMUX g17ba1 ( \45366_nG17ba1 , RIdc22218_6143 , \45365 , \44810 );
_HMUX g17ba2 ( \45367_nG17ba2 , RIdc22218_6143 , \45366_nG17ba1 , \44817 );
buf \U$37746 ( \45368 , RIb838c90_177);
_HMUX g17ba3 ( \45369_nG17ba3 , RIdc22218_6143 , \45368 , \44822 );
_HMUX g17ba4 ( \45370_nG17ba4 , \45367_nG17ba2 , \45369_nG17ba3 , \44829 );
buf \U$37747 ( \45371 , \45370_nG17ba4 );
_DC g192f0_GF_IsGateDCbyConstraint ( \45372_nG192f0 , \45371 , \42503 );
buf \U$37748 ( \45373 , \45372_nG192f0 );
buf \U$37749 ( \45374 , RIb886dc8_8);
_HMUX g17ba5 ( \45375_nG17ba5 , RIda953d8_6144 , \45374 , \44810 );
_HMUX g17ba6 ( \45376_nG17ba6 , RIda953d8_6144 , \45375_nG17ba5 , \44817 );
buf \U$37750 ( \45377 , RIb838d08_176);
_HMUX g17ba7 ( \45378_nG17ba7 , RIda953d8_6144 , \45377 , \44822 );
_HMUX g17ba8 ( \45379_nG17ba8 , \45376_nG17ba6 , \45378_nG17ba7 , \44829 );
buf \U$37751 ( \45380 , \45379_nG17ba8 );
_DC g192f2_GF_IsGateDCbyConstraint ( \45381_nG192f2 , \45380 , \42503 );
buf \U$37752 ( \45382 , \45381_nG192f2 );
buf \U$37753 ( \45383 , RIb886e40_7);
_HMUX g17ba9 ( \45384_nG17ba9 , RIddeaf80_6145 , \45383 , \44810 );
_HMUX g17baa ( \45385_nG17baa , RIddeaf80_6145 , \45384_nG17ba9 , \44817 );
buf \U$37754 ( \45386 , RIb838d80_175);
_HMUX g17bab ( \45387_nG17bab , RIddeaf80_6145 , \45386 , \44822 );
_HMUX g17bac ( \45388_nG17bac , \45385_nG17baa , \45387_nG17bab , \44829 );
buf \U$37755 ( \45389 , \45388_nG17bac );
_DC g192f4_GF_IsGateDCbyConstraint ( \45390_nG192f4 , \45389 , \42503 );
buf \U$37756 ( \45391 , \45390_nG192f4 );
buf \U$37757 ( \45392 , RIb886eb8_6);
_HMUX g17bad ( \45393_nG17bad , RIde58a80_6146 , \45392 , \44810 );
_HMUX g17bae ( \45394_nG17bae , RIde58a80_6146 , \45393_nG17bad , \44817 );
buf \U$37758 ( \45395 , RIb838df8_174);
_HMUX g17baf ( \45396_nG17baf , RIde58a80_6146 , \45395 , \44822 );
_HMUX g17bb0 ( \45397_nG17bb0 , \45394_nG17bae , \45396_nG17baf , \44829 );
buf \U$37759 ( \45398 , \45397_nG17bb0 );
_DC g192f6_GF_IsGateDCbyConstraint ( \45399_nG192f6 , \45398 , \42503 );
buf \U$37760 ( \45400 , \45399_nG192f6 );
not \U$37761 ( \45401 , \44809 );
and \U$37762 ( \45402 , \44808 , \45401 );
_HMUX g179af ( \45403_nG179af , RIe03fa40_6147 , \44807 , \45402 );
_HMUX g179b0 ( \45404_nG179b0 , RIe03fa40_6147 , \45403_nG179af , \44817 );
not \U$37763 ( \45405 , \44821 );
and \U$37764 ( \45406 , \44820 , \45405 );
_HMUX g179b2 ( \45407_nG179b2 , RIe03fa40_6147 , \44819 , \45406 );
_HMUX g179b3 ( \45408_nG179b3 , \45404_nG179b0 , \45407_nG179b2 , \44829 );
buf \U$37765 ( \45409 , \45408_nG179b3 );
_DC g191fe_GF_IsGateDCbyConstraint ( \45410_nG191fe , \45409 , \42503 );
buf \U$37766 ( \45411 , \45410_nG191fe );
_HMUX g179b4 ( \45412_nG179b4 , RIe04e338_6148 , \44834 , \45402 );
_HMUX g179b5 ( \45413_nG179b5 , RIe04e338_6148 , \45412_nG179b4 , \44817 );
_HMUX g179b6 ( \45414_nG179b6 , RIe04e338_6148 , \44837 , \45406 );
_HMUX g179b7 ( \45415_nG179b7 , \45413_nG179b5 , \45414_nG179b6 , \44829 );
buf \U$37767 ( \45416 , \45415_nG179b7 );
_DC g19214_GF_IsGateDCbyConstraint ( \45417_nG19214 , \45416 , \42503 );
buf \U$37768 ( \45418 , \45417_nG19214 );
_HMUX g179b8 ( \45419_nG179b8 , RIe0629f0_6149 , \44843 , \45402 );
_HMUX g179b9 ( \45420_nG179b9 , RIe0629f0_6149 , \45419_nG179b8 , \44817 );
_HMUX g179ba ( \45421_nG179ba , RIe0629f0_6149 , \44846 , \45406 );
_HMUX g179bb ( \45422_nG179bb , \45420_nG179b9 , \45421_nG179ba , \44829 );
buf \U$37769 ( \45423 , \45422_nG179bb );
_DC g1922a_GF_IsGateDCbyConstraint ( \45424_nG1922a , \45423 , \42503 );
buf \U$37770 ( \45425 , \45424_nG1922a );
_HMUX g179bc ( \45426_nG179bc , RIe06c608_6150 , \44852 , \45402 );
_HMUX g179bd ( \45427_nG179bd , RIe06c608_6150 , \45426_nG179bc , \44817 );
_HMUX g179be ( \45428_nG179be , RIe06c608_6150 , \44855 , \45406 );
_HMUX g179bf ( \45429_nG179bf , \45427_nG179bd , \45428_nG179be , \44829 );
buf \U$37771 ( \45430 , \45429_nG179bf );
_DC g19240_GF_IsGateDCbyConstraint ( \45431_nG19240 , \45430 , \42503 );
buf \U$37772 ( \45432 , \45431_nG19240 );
_HMUX g179c0 ( \45433_nG179c0 , RIe0732e0_6151 , \44861 , \45402 );
_HMUX g179c1 ( \45434_nG179c1 , RIe0732e0_6151 , \45433_nG179c0 , \44817 );
_HMUX g179c2 ( \45435_nG179c2 , RIe0732e0_6151 , \44864 , \45406 );
_HMUX g179c3 ( \45436_nG179c3 , \45434_nG179c1 , \45435_nG179c2 , \44829 );
buf \U$37773 ( \45437 , \45436_nG179c3 );
_DC g19256_GF_IsGateDCbyConstraint ( \45438_nG19256 , \45437 , \42503 );
buf \U$37774 ( \45439 , \45438_nG19256 );
_HMUX g179c4 ( \45440_nG179c4 , RIe07d0d8_6152 , \44870 , \45402 );
_HMUX g179c5 ( \45441_nG179c5 , RIe07d0d8_6152 , \45440_nG179c4 , \44817 );
_HMUX g179c6 ( \45442_nG179c6 , RIe07d0d8_6152 , \44873 , \45406 );
_HMUX g179c7 ( \45443_nG179c7 , \45441_nG179c5 , \45442_nG179c6 , \44829 );
buf \U$37775 ( \45444 , \45443_nG179c7 );
_DC g1926c_GF_IsGateDCbyConstraint ( \45445_nG1926c , \45444 , \42503 );
buf \U$37776 ( \45446 , \45445_nG1926c );
_HMUX g179c8 ( \45447_nG179c8 , RIe084158_6153 , \44879 , \45402 );
_HMUX g179c9 ( \45448_nG179c9 , RIe084158_6153 , \45447_nG179c8 , \44817 );
_HMUX g179ca ( \45449_nG179ca , RIe084158_6153 , \44882 , \45406 );
_HMUX g179cb ( \45450_nG179cb , \45448_nG179c9 , \45449_nG179ca , \44829 );
buf \U$37777 ( \45451 , \45450_nG179cb );
_DC g19278_GF_IsGateDCbyConstraint ( \45452_nG19278 , \45451 , \42503 );
buf \U$37778 ( \45453 , \45452_nG19278 );
_HMUX g179cc ( \45454_nG179cc , RIdfc61e0_6154 , \44888 , \45402 );
_HMUX g179cd ( \45455_nG179cd , RIdfc61e0_6154 , \45454_nG179cc , \44817 );
_HMUX g179ce ( \45456_nG179ce , RIdfc61e0_6154 , \44891 , \45406 );
_HMUX g179cf ( \45457_nG179cf , \45455_nG179cd , \45456_nG179ce , \44829 );
buf \U$37779 ( \45458 , \45457_nG179cf );
_DC g1927a_GF_IsGateDCbyConstraint ( \45459_nG1927a , \45458 , \42503 );
buf \U$37780 ( \45460 , \45459_nG1927a );
_HMUX g179d0 ( \45461_nG179d0 , RIe106838_6155 , \44897 , \45402 );
_HMUX g179d1 ( \45462_nG179d1 , RIe106838_6155 , \45461_nG179d0 , \44817 );
_HMUX g179d2 ( \45463_nG179d2 , RIe106838_6155 , \44900 , \45406 );
_HMUX g179d3 ( \45464_nG179d3 , \45462_nG179d1 , \45463_nG179d2 , \44829 );
buf \U$37781 ( \45465 , \45464_nG179d3 );
_DC g1927c_GF_IsGateDCbyConstraint ( \45466_nG1927c , \45465 , \42503 );
buf \U$37782 ( \45467 , \45466_nG1927c );
_HMUX g179d4 ( \45468_nG179d4 , RIe0f8198_6156 , \44906 , \45402 );
_HMUX g179d5 ( \45469_nG179d5 , RIe0f8198_6156 , \45468_nG179d4 , \44817 );
_HMUX g179d6 ( \45470_nG179d6 , RIe0f8198_6156 , \44909 , \45406 );
_HMUX g179d7 ( \45471_nG179d7 , \45469_nG179d5 , \45470_nG179d6 , \44829 );
buf \U$37783 ( \45472 , \45471_nG179d7 );
_DC g19200_GF_IsGateDCbyConstraint ( \45473_nG19200 , \45472 , \42503 );
buf \U$37784 ( \45474 , \45473_nG19200 );
_HMUX g179d8 ( \45475_nG179d8 , RIe0eed00_6157 , \44915 , \45402 );
_HMUX g179d9 ( \45476_nG179d9 , RIe0eed00_6157 , \45475_nG179d8 , \44817 );
_HMUX g179da ( \45477_nG179da , RIe0eed00_6157 , \44918 , \45406 );
_HMUX g179db ( \45478_nG179db , \45476_nG179d9 , \45477_nG179da , \44829 );
buf \U$37785 ( \45479 , \45478_nG179db );
_DC g19202_GF_IsGateDCbyConstraint ( \45480_nG19202 , \45479 , \42503 );
buf \U$37786 ( \45481 , \45480_nG19202 );
_HMUX g179dc ( \45482_nG179dc , RIe0e2b68_6158 , \44924 , \45402 );
_HMUX g179dd ( \45483_nG179dd , RIe0e2b68_6158 , \45482_nG179dc , \44817 );
_HMUX g179de ( \45484_nG179de , RIe0e2b68_6158 , \44927 , \45406 );
_HMUX g179df ( \45485_nG179df , \45483_nG179dd , \45484_nG179de , \44829 );
buf \U$37787 ( \45486 , \45485_nG179df );
_DC g19204_GF_IsGateDCbyConstraint ( \45487_nG19204 , \45486 , \42503 );
buf \U$37788 ( \45488 , \45487_nG19204 );
_HMUX g179e0 ( \45489_nG179e0 , RIe0d0b98_6159 , \44933 , \45402 );
_HMUX g179e1 ( \45490_nG179e1 , RIe0d0b98_6159 , \45489_nG179e0 , \44817 );
_HMUX g179e2 ( \45491_nG179e2 , RIe0d0b98_6159 , \44936 , \45406 );
_HMUX g179e3 ( \45492_nG179e3 , \45490_nG179e1 , \45491_nG179e2 , \44829 );
buf \U$37789 ( \45493 , \45492_nG179e3 );
_DC g19206_GF_IsGateDCbyConstraint ( \45494_nG19206 , \45493 , \42503 );
buf \U$37790 ( \45495 , \45494_nG19206 );
_HMUX g179e4 ( \45496_nG179e4 , RIe0c3998_6160 , \44942 , \45402 );
_HMUX g179e5 ( \45497_nG179e5 , RIe0c3998_6160 , \45496_nG179e4 , \44817 );
_HMUX g179e6 ( \45498_nG179e6 , RIe0c3998_6160 , \44945 , \45406 );
_HMUX g179e7 ( \45499_nG179e7 , \45497_nG179e5 , \45498_nG179e6 , \44829 );
buf \U$37791 ( \45500 , \45499_nG179e7 );
_DC g19208_GF_IsGateDCbyConstraint ( \45501_nG19208 , \45500 , \42503 );
buf \U$37792 ( \45502 , \45501_nG19208 );
_HMUX g179e8 ( \45503_nG179e8 , RIe0b0960_6161 , \44951 , \45402 );
_HMUX g179e9 ( \45504_nG179e9 , RIe0b0960_6161 , \45503_nG179e8 , \44817 );
_HMUX g179ea ( \45505_nG179ea , RIe0b0960_6161 , \44954 , \45406 );
_HMUX g179eb ( \45506_nG179eb , \45504_nG179e9 , \45505_nG179ea , \44829 );
buf \U$37793 ( \45507 , \45506_nG179eb );
_DC g1920a_GF_IsGateDCbyConstraint ( \45508_nG1920a , \45507 , \42503 );
buf \U$37794 ( \45509 , \45508_nG1920a );
_HMUX g179ec ( \45510_nG179ec , RIe0a6988_6162 , \44960 , \45402 );
_HMUX g179ed ( \45511_nG179ed , RIe0a6988_6162 , \45510_nG179ec , \44817 );
_HMUX g179ee ( \45512_nG179ee , RIe0a6988_6162 , \44963 , \45406 );
_HMUX g179ef ( \45513_nG179ef , \45511_nG179ed , \45512_nG179ee , \44829 );
buf \U$37795 ( \45514 , \45513_nG179ef );
_DC g1920c_GF_IsGateDCbyConstraint ( \45515_nG1920c , \45514 , \42503 );
buf \U$37796 ( \45516 , \45515_nG1920c );
_HMUX g179f0 ( \45517_nG179f0 , RIe099440_6163 , \44969 , \45402 );
_HMUX g179f1 ( \45518_nG179f1 , RIe099440_6163 , \45517_nG179f0 , \44817 );
_HMUX g179f2 ( \45519_nG179f2 , RIe099440_6163 , \44972 , \45406 );
_HMUX g179f3 ( \45520_nG179f3 , \45518_nG179f1 , \45519_nG179f2 , \44829 );
buf \U$37797 ( \45521 , \45520_nG179f3 );
_DC g1920e_GF_IsGateDCbyConstraint ( \45522_nG1920e , \45521 , \42503 );
buf \U$37798 ( \45523 , \45522_nG1920e );
_HMUX g179f4 ( \45524_nG179f4 , RIe1d3c60_6164 , \44978 , \45402 );
_HMUX g179f5 ( \45525_nG179f5 , RIe1d3c60_6164 , \45524_nG179f4 , \44817 );
_HMUX g179f6 ( \45526_nG179f6 , RIe1d3c60_6164 , \44981 , \45406 );
_HMUX g179f7 ( \45527_nG179f7 , \45525_nG179f5 , \45526_nG179f6 , \44829 );
buf \U$37799 ( \45528 , \45527_nG179f7 );
_DC g19210_GF_IsGateDCbyConstraint ( \45529_nG19210 , \45528 , \42503 );
buf \U$37800 ( \45530 , \45529_nG19210 );
_HMUX g179f8 ( \45531_nG179f8 , RIe1d69d8_6165 , \44987 , \45402 );
_HMUX g179f9 ( \45532_nG179f9 , RIe1d69d8_6165 , \45531_nG179f8 , \44817 );
_HMUX g179fa ( \45533_nG179fa , RIe1d69d8_6165 , \44990 , \45406 );
_HMUX g179fb ( \45534_nG179fb , \45532_nG179f9 , \45533_nG179fa , \44829 );
buf \U$37801 ( \45535 , \45534_nG179fb );
_DC g19212_GF_IsGateDCbyConstraint ( \45536_nG19212 , \45535 , \42503 );
buf \U$37802 ( \45537 , \45536_nG19212 );
_HMUX g179fc ( \45538_nG179fc , RIe1d9c00_6166 , \44996 , \45402 );
_HMUX g179fd ( \45539_nG179fd , RIe1d9c00_6166 , \45538_nG179fc , \44817 );
_HMUX g179fe ( \45540_nG179fe , RIe1d9c00_6166 , \44999 , \45406 );
_HMUX g179ff ( \45541_nG179ff , \45539_nG179fd , \45540_nG179fe , \44829 );
buf \U$37803 ( \45542 , \45541_nG179ff );
_DC g19216_GF_IsGateDCbyConstraint ( \45543_nG19216 , \45542 , \42503 );
buf \U$37804 ( \45544 , \45543_nG19216 );
_HMUX g17a00 ( \45545_nG17a00 , RIe1dc978_6167 , \45005 , \45402 );
_HMUX g17a01 ( \45546_nG17a01 , RIe1dc978_6167 , \45545_nG17a00 , \44817 );
_HMUX g17a02 ( \45547_nG17a02 , RIe1dc978_6167 , \45008 , \45406 );
_HMUX g17a03 ( \45548_nG17a03 , \45546_nG17a01 , \45547_nG17a02 , \44829 );
buf \U$37805 ( \45549 , \45548_nG17a03 );
_DC g19218_GF_IsGateDCbyConstraint ( \45550_nG19218 , \45549 , \42503 );
buf \U$37806 ( \45551 , \45550_nG19218 );
_HMUX g17a04 ( \45552_nG17a04 , RIe1dfba0_6168 , \45014 , \45402 );
_HMUX g17a05 ( \45553_nG17a05 , RIe1dfba0_6168 , \45552_nG17a04 , \44817 );
_HMUX g17a06 ( \45554_nG17a06 , RIe1dfba0_6168 , \45017 , \45406 );
_HMUX g17a07 ( \45555_nG17a07 , \45553_nG17a05 , \45554_nG17a06 , \44829 );
buf \U$37807 ( \45556 , \45555_nG17a07 );
_DC g1921a_GF_IsGateDCbyConstraint ( \45557_nG1921a , \45556 , \42503 );
buf \U$37808 ( \45558 , \45557_nG1921a );
_HMUX g17a08 ( \45559_nG17a08 , RIe1e2918_6169 , \45023 , \45402 );
_HMUX g17a09 ( \45560_nG17a09 , RIe1e2918_6169 , \45559_nG17a08 , \44817 );
_HMUX g17a0a ( \45561_nG17a0a , RIe1e2918_6169 , \45026 , \45406 );
_HMUX g17a0b ( \45562_nG17a0b , \45560_nG17a09 , \45561_nG17a0a , \44829 );
buf \U$37809 ( \45563 , \45562_nG17a0b );
_DC g1921c_GF_IsGateDCbyConstraint ( \45564_nG1921c , \45563 , \42503 );
buf \U$37810 ( \45565 , \45564_nG1921c );
_HMUX g17a0c ( \45566_nG17a0c , RIe1e5b40_6170 , \45032 , \45402 );
_HMUX g17a0d ( \45567_nG17a0d , RIe1e5b40_6170 , \45566_nG17a0c , \44817 );
_HMUX g17a0e ( \45568_nG17a0e , RIe1e5b40_6170 , \45035 , \45406 );
_HMUX g17a0f ( \45569_nG17a0f , \45567_nG17a0d , \45568_nG17a0e , \44829 );
buf \U$37811 ( \45570 , \45569_nG17a0f );
_DC g1921e_GF_IsGateDCbyConstraint ( \45571_nG1921e , \45570 , \42503 );
buf \U$37812 ( \45572 , \45571_nG1921e );
_HMUX g17a10 ( \45573_nG17a10 , RIe1e88b8_6171 , \45041 , \45402 );
_HMUX g17a11 ( \45574_nG17a11 , RIe1e88b8_6171 , \45573_nG17a10 , \44817 );
_HMUX g17a12 ( \45575_nG17a12 , RIe1e88b8_6171 , \45044 , \45406 );
_HMUX g17a13 ( \45576_nG17a13 , \45574_nG17a11 , \45575_nG17a12 , \44829 );
buf \U$37813 ( \45577 , \45576_nG17a13 );
_DC g19220_GF_IsGateDCbyConstraint ( \45578_nG19220 , \45577 , \42503 );
buf \U$37814 ( \45579 , \45578_nG19220 );
_HMUX g17a14 ( \45580_nG17a14 , RIe1eb180_6172 , \45050 , \45402 );
_HMUX g17a15 ( \45581_nG17a15 , RIe1eb180_6172 , \45580_nG17a14 , \44817 );
_HMUX g17a16 ( \45582_nG17a16 , RIe1eb180_6172 , \45053 , \45406 );
_HMUX g17a17 ( \45583_nG17a17 , \45581_nG17a15 , \45582_nG17a16 , \44829 );
buf \U$37815 ( \45584 , \45583_nG17a17 );
_DC g19222_GF_IsGateDCbyConstraint ( \45585_nG19222 , \45584 , \42503 );
buf \U$37816 ( \45586 , \45585_nG19222 );
_HMUX g17a18 ( \45587_nG17a18 , RIe1ee858_6173 , \45059 , \45402 );
_HMUX g17a19 ( \45588_nG17a19 , RIe1ee858_6173 , \45587_nG17a18 , \44817 );
_HMUX g17a1a ( \45589_nG17a1a , RIe1ee858_6173 , \45062 , \45406 );
_HMUX g17a1b ( \45590_nG17a1b , \45588_nG17a19 , \45589_nG17a1a , \44829 );
buf \U$37817 ( \45591 , \45590_nG17a1b );
_DC g19224_GF_IsGateDCbyConstraint ( \45592_nG19224 , \45591 , \42503 );
buf \U$37818 ( \45593 , \45592_nG19224 );
_HMUX g17a1c ( \45594_nG17a1c , RIe1f1120_6174 , \45068 , \45402 );
_HMUX g17a1d ( \45595_nG17a1d , RIe1f1120_6174 , \45594_nG17a1c , \44817 );
_HMUX g17a1e ( \45596_nG17a1e , RIe1f1120_6174 , \45071 , \45406 );
_HMUX g17a1f ( \45597_nG17a1f , \45595_nG17a1d , \45596_nG17a1e , \44829 );
buf \U$37819 ( \45598 , \45597_nG17a1f );
_DC g19226_GF_IsGateDCbyConstraint ( \45599_nG19226 , \45598 , \42503 );
buf \U$37820 ( \45600 , \45599_nG19226 );
_HMUX g17a20 ( \45601_nG17a20 , RIe1f47f8_6175 , \45077 , \45402 );
_HMUX g17a21 ( \45602_nG17a21 , RIe1f47f8_6175 , \45601_nG17a20 , \44817 );
_HMUX g17a22 ( \45603_nG17a22 , RIe1f47f8_6175 , \45080 , \45406 );
_HMUX g17a23 ( \45604_nG17a23 , \45602_nG17a21 , \45603_nG17a22 , \44829 );
buf \U$37821 ( \45605 , \45604_nG17a23 );
_DC g19228_GF_IsGateDCbyConstraint ( \45606_nG19228 , \45605 , \42503 );
buf \U$37822 ( \45607 , \45606_nG19228 );
_HMUX g17a24 ( \45608_nG17a24 , RIe1f70c0_6176 , \45086 , \45402 );
_HMUX g17a25 ( \45609_nG17a25 , RIe1f70c0_6176 , \45608_nG17a24 , \44817 );
_HMUX g17a26 ( \45610_nG17a26 , RIe1f70c0_6176 , \45089 , \45406 );
_HMUX g17a27 ( \45611_nG17a27 , \45609_nG17a25 , \45610_nG17a26 , \44829 );
buf \U$37823 ( \45612 , \45611_nG17a27 );
_DC g1922c_GF_IsGateDCbyConstraint ( \45613_nG1922c , \45612 , \42503 );
buf \U$37824 ( \45614 , \45613_nG1922c );
_HMUX g17a28 ( \45615_nG17a28 , RIe1fa180_6177 , \45095 , \45402 );
_HMUX g17a29 ( \45616_nG17a29 , RIe1fa180_6177 , \45615_nG17a28 , \44817 );
_HMUX g17a2a ( \45617_nG17a2a , RIe1fa180_6177 , \45098 , \45406 );
_HMUX g17a2b ( \45618_nG17a2b , \45616_nG17a29 , \45617_nG17a2a , \44829 );
buf \U$37825 ( \45619 , \45618_nG17a2b );
_DC g1922e_GF_IsGateDCbyConstraint ( \45620_nG1922e , \45619 , \42503 );
buf \U$37826 ( \45621 , \45620_nG1922e );
_HMUX g17a2c ( \45622_nG17a2c , RIe1fbad0_6178 , \45104 , \45402 );
_HMUX g17a2d ( \45623_nG17a2d , RIe1fbad0_6178 , \45622_nG17a2c , \44817 );
_HMUX g17a2e ( \45624_nG17a2e , RIe1fbad0_6178 , \45107 , \45406 );
_HMUX g17a2f ( \45625_nG17a2f , \45623_nG17a2d , \45624_nG17a2e , \44829 );
buf \U$37827 ( \45626 , \45625_nG17a2f );
_DC g19230_GF_IsGateDCbyConstraint ( \45627_nG19230 , \45626 , \42503 );
buf \U$37828 ( \45628 , \45627_nG19230 );
_HMUX g17a30 ( \45629_nG17a30 , RIe1fd330_6179 , \45113 , \45402 );
_HMUX g17a31 ( \45630_nG17a31 , RIe1fd330_6179 , \45629_nG17a30 , \44817 );
_HMUX g17a32 ( \45631_nG17a32 , RIe1fd330_6179 , \45116 , \45406 );
_HMUX g17a33 ( \45632_nG17a33 , \45630_nG17a31 , \45631_nG17a32 , \44829 );
buf \U$37829 ( \45633 , \45632_nG17a33 );
_DC g19232_GF_IsGateDCbyConstraint ( \45634_nG19232 , \45633 , \42503 );
buf \U$37830 ( \45635 , \45634_nG19232 );
_HMUX g17a34 ( \45636_nG17a34 , RIe1ff568_6180 , \45122 , \45402 );
_HMUX g17a35 ( \45637_nG17a35 , RIe1ff568_6180 , \45636_nG17a34 , \44817 );
_HMUX g17a36 ( \45638_nG17a36 , RIe1ff568_6180 , \45125 , \45406 );
_HMUX g17a37 ( \45639_nG17a37 , \45637_nG17a35 , \45638_nG17a36 , \44829 );
buf \U$37831 ( \45640 , \45639_nG17a37 );
_DC g19234_GF_IsGateDCbyConstraint ( \45641_nG19234 , \45640 , \42503 );
buf \U$37832 ( \45642 , \45641_nG19234 );
_HMUX g17a38 ( \45643_nG17a38 , RIe2012f0_6181 , \45131 , \45402 );
_HMUX g17a39 ( \45644_nG17a39 , RIe2012f0_6181 , \45643_nG17a38 , \44817 );
_HMUX g17a3a ( \45645_nG17a3a , RIe2012f0_6181 , \45134 , \45406 );
_HMUX g17a3b ( \45646_nG17a3b , \45644_nG17a39 , \45645_nG17a3a , \44829 );
buf \U$37833 ( \45647 , \45646_nG17a3b );
_DC g19236_GF_IsGateDCbyConstraint ( \45648_nG19236 , \45647 , \42503 );
buf \U$37834 ( \45649 , \45648_nG19236 );
_HMUX g17a3c ( \45650_nG17a3c , RIe203000_6182 , \45140 , \45402 );
_HMUX g17a3d ( \45651_nG17a3d , RIe203000_6182 , \45650_nG17a3c , \44817 );
_HMUX g17a3e ( \45652_nG17a3e , RIe203000_6182 , \45143 , \45406 );
_HMUX g17a3f ( \45653_nG17a3f , \45651_nG17a3d , \45652_nG17a3e , \44829 );
buf \U$37835 ( \45654 , \45653_nG17a3f );
_DC g19238_GF_IsGateDCbyConstraint ( \45655_nG19238 , \45654 , \42503 );
buf \U$37836 ( \45656 , \45655_nG19238 );
_HMUX g17a40 ( \45657_nG17a40 , RIe203f00_6183 , \45149 , \45402 );
_HMUX g17a41 ( \45658_nG17a41 , RIe203f00_6183 , \45657_nG17a40 , \44817 );
_HMUX g17a42 ( \45659_nG17a42 , RIe203f00_6183 , \45152 , \45406 );
_HMUX g17a43 ( \45660_nG17a43 , \45658_nG17a41 , \45659_nG17a42 , \44829 );
buf \U$37837 ( \45661 , \45660_nG17a43 );
_DC g1923a_GF_IsGateDCbyConstraint ( \45662_nG1923a , \45661 , \42503 );
buf \U$37838 ( \45663 , \45662_nG1923a );
_HMUX g17a44 ( \45664_nG17a44 , RIe2053a0_6184 , \45158 , \45402 );
_HMUX g17a45 ( \45665_nG17a45 , RIe2053a0_6184 , \45664_nG17a44 , \44817 );
_HMUX g17a46 ( \45666_nG17a46 , RIe2053a0_6184 , \45161 , \45406 );
_HMUX g17a47 ( \45667_nG17a47 , \45665_nG17a45 , \45666_nG17a46 , \44829 );
buf \U$37839 ( \45668 , \45667_nG17a47 );
_DC g1923c_GF_IsGateDCbyConstraint ( \45669_nG1923c , \45668 , \42503 );
buf \U$37840 ( \45670 , \45669_nG1923c );
_HMUX g17a48 ( \45671_nG17a48 , RIe2066d8_6185 , \45167 , \45402 );
_HMUX g17a49 ( \45672_nG17a49 , RIe2066d8_6185 , \45671_nG17a48 , \44817 );
_HMUX g17a4a ( \45673_nG17a4a , RIe2066d8_6185 , \45170 , \45406 );
_HMUX g17a4b ( \45674_nG17a4b , \45672_nG17a49 , \45673_nG17a4a , \44829 );
buf \U$37841 ( \45675 , \45674_nG17a4b );
_DC g1923e_GF_IsGateDCbyConstraint ( \45676_nG1923e , \45675 , \42503 );
buf \U$37842 ( \45677 , \45676_nG1923e );
_HMUX g17a4c ( \45678_nG17a4c , RIe207920_6186 , \45176 , \45402 );
_HMUX g17a4d ( \45679_nG17a4d , RIe207920_6186 , \45678_nG17a4c , \44817 );
_HMUX g17a4e ( \45680_nG17a4e , RIe207920_6186 , \45179 , \45406 );
_HMUX g17a4f ( \45681_nG17a4f , \45679_nG17a4d , \45680_nG17a4e , \44829 );
buf \U$37843 ( \45682 , \45681_nG17a4f );
_DC g19242_GF_IsGateDCbyConstraint ( \45683_nG19242 , \45682 , \42503 );
buf \U$37844 ( \45684 , \45683_nG19242 );
_HMUX g17a50 ( \45685_nG17a50 , RIe208be0_6187 , \45185 , \45402 );
_HMUX g17a51 ( \45686_nG17a51 , RIe208be0_6187 , \45685_nG17a50 , \44817 );
_HMUX g17a52 ( \45687_nG17a52 , RIe208be0_6187 , \45188 , \45406 );
_HMUX g17a53 ( \45688_nG17a53 , \45686_nG17a51 , \45687_nG17a52 , \44829 );
buf \U$37845 ( \45689 , \45688_nG17a53 );
_DC g19244_GF_IsGateDCbyConstraint ( \45690_nG19244 , \45689 , \42503 );
buf \U$37846 ( \45691 , \45690_nG19244 );
_HMUX g17a54 ( \45692_nG17a54 , RIe209d38_6188 , \45194 , \45402 );
_HMUX g17a55 ( \45693_nG17a55 , RIe209d38_6188 , \45692_nG17a54 , \44817 );
_HMUX g17a56 ( \45694_nG17a56 , RIe209d38_6188 , \45197 , \45406 );
_HMUX g17a57 ( \45695_nG17a57 , \45693_nG17a55 , \45694_nG17a56 , \44829 );
buf \U$37847 ( \45696 , \45695_nG17a57 );
_DC g19246_GF_IsGateDCbyConstraint ( \45697_nG19246 , \45696 , \42503 );
buf \U$37848 ( \45698 , \45697_nG19246 );
_HMUX g17a58 ( \45699_nG17a58 , RIe20b958_6189 , \45203 , \45402 );
_HMUX g17a59 ( \45700_nG17a59 , RIe20b958_6189 , \45699_nG17a58 , \44817 );
_HMUX g17a5a ( \45701_nG17a5a , RIe20b958_6189 , \45206 , \45406 );
_HMUX g17a5b ( \45702_nG17a5b , \45700_nG17a59 , \45701_nG17a5a , \44829 );
buf \U$37849 ( \45703 , \45702_nG17a5b );
_DC g19248_GF_IsGateDCbyConstraint ( \45704_nG19248 , \45703 , \42503 );
buf \U$37850 ( \45705 , \45704_nG19248 );
_HMUX g17a5c ( \45706_nG17a5c , RIe20cf60_6190 , \45212 , \45402 );
_HMUX g17a5d ( \45707_nG17a5d , RIe20cf60_6190 , \45706_nG17a5c , \44817 );
_HMUX g17a5e ( \45708_nG17a5e , RIe20cf60_6190 , \45215 , \45406 );
_HMUX g17a5f ( \45709_nG17a5f , \45707_nG17a5d , \45708_nG17a5e , \44829 );
buf \U$37851 ( \45710 , \45709_nG17a5f );
_DC g1924a_GF_IsGateDCbyConstraint ( \45711_nG1924a , \45710 , \42503 );
buf \U$37852 ( \45712 , \45711_nG1924a );
_HMUX g17a60 ( \45713_nG17a60 , RIe20e4f0_6191 , \45221 , \45402 );
_HMUX g17a61 ( \45714_nG17a61 , RIe20e4f0_6191 , \45713_nG17a60 , \44817 );
_HMUX g17a62 ( \45715_nG17a62 , RIe20e4f0_6191 , \45224 , \45406 );
_HMUX g17a63 ( \45716_nG17a63 , \45714_nG17a61 , \45715_nG17a62 , \44829 );
buf \U$37853 ( \45717 , \45716_nG17a63 );
_DC g1924c_GF_IsGateDCbyConstraint ( \45718_nG1924c , \45717 , \42503 );
buf \U$37854 ( \45719 , \45718_nG1924c );
_HMUX g17a64 ( \45720_nG17a64 , RIe20f5d0_6192 , \45230 , \45402 );
_HMUX g17a65 ( \45721_nG17a65 , RIe20f5d0_6192 , \45720_nG17a64 , \44817 );
_HMUX g17a66 ( \45722_nG17a66 , RIe20f5d0_6192 , \45233 , \45406 );
_HMUX g17a67 ( \45723_nG17a67 , \45721_nG17a65 , \45722_nG17a66 , \44829 );
buf \U$37855 ( \45724 , \45723_nG17a67 );
_DC g1924e_GF_IsGateDCbyConstraint ( \45725_nG1924e , \45724 , \42503 );
buf \U$37856 ( \45726 , \45725_nG1924e );
_HMUX g17a68 ( \45727_nG17a68 , RIe211178_6193 , \45239 , \45402 );
_HMUX g17a69 ( \45728_nG17a69 , RIe211178_6193 , \45727_nG17a68 , \44817 );
_HMUX g17a6a ( \45729_nG17a6a , RIe211178_6193 , \45242 , \45406 );
_HMUX g17a6b ( \45730_nG17a6b , \45728_nG17a69 , \45729_nG17a6a , \44829 );
buf \U$37857 ( \45731 , \45730_nG17a6b );
_DC g19250_GF_IsGateDCbyConstraint ( \45732_nG19250 , \45731 , \42503 );
buf \U$37858 ( \45733 , \45732_nG19250 );
_HMUX g17a6c ( \45734_nG17a6c , RIe212c30_6194 , \45248 , \45402 );
_HMUX g17a6d ( \45735_nG17a6d , RIe212c30_6194 , \45734_nG17a6c , \44817 );
_HMUX g17a6e ( \45736_nG17a6e , RIe212c30_6194 , \45251 , \45406 );
_HMUX g17a6f ( \45737_nG17a6f , \45735_nG17a6d , \45736_nG17a6e , \44829 );
buf \U$37859 ( \45738 , \45737_nG17a6f );
_DC g19252_GF_IsGateDCbyConstraint ( \45739_nG19252 , \45738 , \42503 );
buf \U$37860 ( \45740 , \45739_nG19252 );
_HMUX g17a70 ( \45741_nG17a70 , RIe214148_6195 , \45257 , \45402 );
_HMUX g17a71 ( \45742_nG17a71 , RIe214148_6195 , \45741_nG17a70 , \44817 );
_HMUX g17a72 ( \45743_nG17a72 , RIe214148_6195 , \45260 , \45406 );
_HMUX g17a73 ( \45744_nG17a73 , \45742_nG17a71 , \45743_nG17a72 , \44829 );
buf \U$37861 ( \45745 , \45744_nG17a73 );
_DC g19254_GF_IsGateDCbyConstraint ( \45746_nG19254 , \45745 , \42503 );
buf \U$37862 ( \45747 , \45746_nG19254 );
_HMUX g17a74 ( \45748_nG17a74 , RIe215c00_6196 , \45266 , \45402 );
_HMUX g17a75 ( \45749_nG17a75 , RIe215c00_6196 , \45748_nG17a74 , \44817 );
_HMUX g17a76 ( \45750_nG17a76 , RIe215c00_6196 , \45269 , \45406 );
_HMUX g17a77 ( \45751_nG17a77 , \45749_nG17a75 , \45750_nG17a76 , \44829 );
buf \U$37863 ( \45752 , \45751_nG17a77 );
_DC g19258_GF_IsGateDCbyConstraint ( \45753_nG19258 , \45752 , \42503 );
buf \U$37864 ( \45754 , \45753_nG19258 );
_HMUX g17a78 ( \45755_nG17a78 , RIe217460_6197 , \45275 , \45402 );
_HMUX g17a79 ( \45756_nG17a79 , RIe217460_6197 , \45755_nG17a78 , \44817 );
_HMUX g17a7a ( \45757_nG17a7a , RIe217460_6197 , \45278 , \45406 );
_HMUX g17a7b ( \45758_nG17a7b , \45756_nG17a79 , \45757_nG17a7a , \44829 );
buf \U$37865 ( \45759 , \45758_nG17a7b );
_DC g1925a_GF_IsGateDCbyConstraint ( \45760_nG1925a , \45759 , \42503 );
buf \U$37866 ( \45761 , \45760_nG1925a );
_HMUX g17a7c ( \45762_nG17a7c , RIe218798_6198 , \45284 , \45402 );
_HMUX g17a7d ( \45763_nG17a7d , RIe218798_6198 , \45762_nG17a7c , \44817 );
_HMUX g17a7e ( \45764_nG17a7e , RIe218798_6198 , \45287 , \45406 );
_HMUX g17a7f ( \45765_nG17a7f , \45763_nG17a7d , \45764_nG17a7e , \44829 );
buf \U$37867 ( \45766 , \45765_nG17a7f );
_DC g1925c_GF_IsGateDCbyConstraint ( \45767_nG1925c , \45766 , \42503 );
buf \U$37868 ( \45768 , \45767_nG1925c );
_HMUX g17a80 ( \45769_nG17a80 , RIe2199e0_6199 , \45293 , \45402 );
_HMUX g17a81 ( \45770_nG17a81 , RIe2199e0_6199 , \45769_nG17a80 , \44817 );
_HMUX g17a82 ( \45771_nG17a82 , RIe2199e0_6199 , \45296 , \45406 );
_HMUX g17a83 ( \45772_nG17a83 , \45770_nG17a81 , \45771_nG17a82 , \44829 );
buf \U$37869 ( \45773 , \45772_nG17a83 );
_DC g1925e_GF_IsGateDCbyConstraint ( \45774_nG1925e , \45773 , \42503 );
buf \U$37870 ( \45775 , \45774_nG1925e );
_HMUX g17a84 ( \45776_nG17a84 , RIe14e868_6200 , \45302 , \45402 );
_HMUX g17a85 ( \45777_nG17a85 , RIe14e868_6200 , \45776_nG17a84 , \44817 );
_HMUX g17a86 ( \45778_nG17a86 , RIe14e868_6200 , \45305 , \45406 );
_HMUX g17a87 ( \45779_nG17a87 , \45777_nG17a85 , \45778_nG17a86 , \44829 );
buf \U$37871 ( \45780 , \45779_nG17a87 );
_DC g19260_GF_IsGateDCbyConstraint ( \45781_nG19260 , \45780 , \42503 );
buf \U$37872 ( \45782 , \45781_nG19260 );
_HMUX g17a88 ( \45783_nG17a88 , RIe151130_6201 , \45311 , \45402 );
_HMUX g17a89 ( \45784_nG17a89 , RIe151130_6201 , \45783_nG17a88 , \44817 );
_HMUX g17a8a ( \45785_nG17a8a , RIe151130_6201 , \45314 , \45406 );
_HMUX g17a8b ( \45786_nG17a8b , \45784_nG17a89 , \45785_nG17a8a , \44829 );
buf \U$37873 ( \45787 , \45786_nG17a8b );
_DC g19262_GF_IsGateDCbyConstraint ( \45788_nG19262 , \45787 , \42503 );
buf \U$37874 ( \45789 , \45788_nG19262 );
_HMUX g17a8c ( \45790_nG17a8c , RIe153020_6202 , \45320 , \45402 );
_HMUX g17a8d ( \45791_nG17a8d , RIe153020_6202 , \45790_nG17a8c , \44817 );
_HMUX g17a8e ( \45792_nG17a8e , RIe153020_6202 , \45323 , \45406 );
_HMUX g17a8f ( \45793_nG17a8f , \45791_nG17a8d , \45792_nG17a8e , \44829 );
buf \U$37875 ( \45794 , \45793_nG17a8f );
_DC g19264_GF_IsGateDCbyConstraint ( \45795_nG19264 , \45794 , \42503 );
buf \U$37876 ( \45796 , \45795_nG19264 );
_HMUX g17a90 ( \45797_nG17a90 , RIe154ad8_6203 , \45329 , \45402 );
_HMUX g17a91 ( \45798_nG17a91 , RIe154ad8_6203 , \45797_nG17a90 , \44817 );
_HMUX g17a92 ( \45799_nG17a92 , RIe154ad8_6203 , \45332 , \45406 );
_HMUX g17a93 ( \45800_nG17a93 , \45798_nG17a91 , \45799_nG17a92 , \44829 );
buf \U$37877 ( \45801 , \45800_nG17a93 );
_DC g19266_GF_IsGateDCbyConstraint ( \45802_nG19266 , \45801 , \42503 );
buf \U$37878 ( \45803 , \45802_nG19266 );
_HMUX g17a94 ( \45804_nG17a94 , RIe156518_6204 , \45338 , \45402 );
_HMUX g17a95 ( \45805_nG17a95 , RIe156518_6204 , \45804_nG17a94 , \44817 );
_HMUX g17a96 ( \45806_nG17a96 , RIe156518_6204 , \45341 , \45406 );
_HMUX g17a97 ( \45807_nG17a97 , \45805_nG17a95 , \45806_nG17a96 , \44829 );
buf \U$37879 ( \45808 , \45807_nG17a97 );
_DC g19268_GF_IsGateDCbyConstraint ( \45809_nG19268 , \45808 , \42503 );
buf \U$37880 ( \45810 , \45809_nG19268 );
_HMUX g17a98 ( \45811_nG17a98 , RIe158228_6205 , \45347 , \45402 );
_HMUX g17a99 ( \45812_nG17a99 , RIe158228_6205 , \45811_nG17a98 , \44817 );
_HMUX g17a9a ( \45813_nG17a9a , RIe158228_6205 , \45350 , \45406 );
_HMUX g17a9b ( \45814_nG17a9b , \45812_nG17a99 , \45813_nG17a9a , \44829 );
buf \U$37881 ( \45815 , \45814_nG17a9b );
_DC g1926a_GF_IsGateDCbyConstraint ( \45816_nG1926a , \45815 , \42503 );
buf \U$37882 ( \45817 , \45816_nG1926a );
_HMUX g17a9c ( \45818_nG17a9c , RIe15a280_6206 , \45356 , \45402 );
_HMUX g17a9d ( \45819_nG17a9d , RIe15a280_6206 , \45818_nG17a9c , \44817 );
_HMUX g17a9e ( \45820_nG17a9e , RIe15a280_6206 , \45359 , \45406 );
_HMUX g17a9f ( \45821_nG17a9f , \45819_nG17a9d , \45820_nG17a9e , \44829 );
buf \U$37883 ( \45822 , \45821_nG17a9f );
_DC g1926e_GF_IsGateDCbyConstraint ( \45823_nG1926e , \45822 , \42503 );
buf \U$37884 ( \45824 , \45823_nG1926e );
_HMUX g17aa0 ( \45825_nG17aa0 , RIe15c3c8_6207 , \45365 , \45402 );
_HMUX g17aa1 ( \45826_nG17aa1 , RIe15c3c8_6207 , \45825_nG17aa0 , \44817 );
_HMUX g17aa2 ( \45827_nG17aa2 , RIe15c3c8_6207 , \45368 , \45406 );
_HMUX g17aa3 ( \45828_nG17aa3 , \45826_nG17aa1 , \45827_nG17aa2 , \44829 );
buf \U$37885 ( \45829 , \45828_nG17aa3 );
_DC g19270_GF_IsGateDCbyConstraint ( \45830_nG19270 , \45829 , \42503 );
buf \U$37886 ( \45831 , \45830_nG19270 );
_HMUX g17aa4 ( \45832_nG17aa4 , RIe15ef60_6208 , \45374 , \45402 );
_HMUX g17aa5 ( \45833_nG17aa5 , RIe15ef60_6208 , \45832_nG17aa4 , \44817 );
_HMUX g17aa6 ( \45834_nG17aa6 , RIe15ef60_6208 , \45377 , \45406 );
_HMUX g17aa7 ( \45835_nG17aa7 , \45833_nG17aa5 , \45834_nG17aa6 , \44829 );
buf \U$37887 ( \45836 , \45835_nG17aa7 );
_DC g19272_GF_IsGateDCbyConstraint ( \45837_nG19272 , \45836 , \42503 );
buf \U$37888 ( \45838 , \45837_nG19272 );
_HMUX g17aa8 ( \45839_nG17aa8 , RIe1616c0_6209 , \45383 , \45402 );
_HMUX g17aa9 ( \45840_nG17aa9 , RIe1616c0_6209 , \45839_nG17aa8 , \44817 );
_HMUX g17aaa ( \45841_nG17aaa , RIe1616c0_6209 , \45386 , \45406 );
_HMUX g17aab ( \45842_nG17aab , \45840_nG17aa9 , \45841_nG17aaa , \44829 );
buf \U$37889 ( \45843 , \45842_nG17aab );
_DC g19274_GF_IsGateDCbyConstraint ( \45844_nG19274 , \45843 , \42503 );
buf \U$37890 ( \45845 , \45844_nG19274 );
_HMUX g17aac ( \45846_nG17aac , RIe164168_6210 , \45392 , \45402 );
_HMUX g17aad ( \45847_nG17aad , RIe164168_6210 , \45846_nG17aac , \44817 );
_HMUX g17aae ( \45848_nG17aae , RIe164168_6210 , \45395 , \45406 );
_HMUX g17aaf ( \45849_nG17aaf , \45847_nG17aad , \45848_nG17aae , \44829 );
buf \U$37891 ( \45850 , \45849_nG17aaf );
_DC g19276_GF_IsGateDCbyConstraint ( \45851_nG19276 , \45850 , \42503 );
buf \U$37892 ( \45852 , \45851_nG19276 );
nor \U$37893 ( \45853 , \44808 , \45401 );
_HMUX g178ad ( \45854_nG178ad , RIe166c10_6211 , \44807 , \45853 );
_HMUX g178ae ( \45855_nG178ae , RIe166c10_6211 , \45854_nG178ad , \44817 );
nor \U$37894 ( \45856 , \44820 , \45405 );
_HMUX g178b1 ( \45857_nG178b1 , RIe166c10_6211 , \44819 , \45856 );
_HMUX g178b2 ( \45858_nG178b2 , \45855_nG178ae , \45857_nG178b1 , \44829 );
buf \U$37895 ( \45859 , \45858_nG178b2 );
_DC g1917e_GF_IsGateDCbyConstraint ( \45860_nG1917e , \45859 , \42503 );
buf \U$37896 ( \45861 , \45860_nG1917e );
_HMUX g178b3 ( \45862_nG178b3 , RIe39a100_6212 , \44834 , \45853 );
_HMUX g178b4 ( \45863_nG178b4 , RIe39a100_6212 , \45862_nG178b3 , \44817 );
_HMUX g178b5 ( \45864_nG178b5 , RIe39a100_6212 , \44837 , \45856 );
_HMUX g178b6 ( \45865_nG178b6 , \45863_nG178b4 , \45864_nG178b5 , \44829 );
buf \U$37897 ( \45866 , \45865_nG178b6 );
_DC g19194_GF_IsGateDCbyConstraint ( \45867_nG19194 , \45866 , \42503 );
buf \U$37898 ( \45868 , \45867_nG19194 );
_HMUX g178b7 ( \45869_nG178b7 , RIe3984e0_6213 , \44843 , \45853 );
_HMUX g178b8 ( \45870_nG178b8 , RIe3984e0_6213 , \45869_nG178b7 , \44817 );
_HMUX g178b9 ( \45871_nG178b9 , RIe3984e0_6213 , \44846 , \45856 );
_HMUX g178ba ( \45872_nG178ba , \45870_nG178b8 , \45871_nG178b9 , \44829 );
buf \U$37899 ( \45873 , \45872_nG178ba );
_DC g191aa_GF_IsGateDCbyConstraint ( \45874_nG191aa , \45873 , \42503 );
buf \U$37900 ( \45875 , \45874_nG191aa );
_HMUX g178bb ( \45876_nG178bb , RIe3967d0_6214 , \44852 , \45853 );
_HMUX g178bc ( \45877_nG178bc , RIe3967d0_6214 , \45876_nG178bb , \44817 );
_HMUX g178bd ( \45878_nG178bd , RIe3967d0_6214 , \44855 , \45856 );
_HMUX g178be ( \45879_nG178be , \45877_nG178bc , \45878_nG178bd , \44829 );
buf \U$37901 ( \45880 , \45879_nG178be );
_DC g191c0_GF_IsGateDCbyConstraint ( \45881_nG191c0 , \45880 , \42503 );
buf \U$37902 ( \45882 , \45881_nG191c0 );
_HMUX g178bf ( \45883_nG178bf , RIe3941d8_6215 , \44861 , \45853 );
_HMUX g178c0 ( \45884_nG178c0 , RIe3941d8_6215 , \45883_nG178bf , \44817 );
_HMUX g178c1 ( \45885_nG178c1 , RIe3941d8_6215 , \44864 , \45856 );
_HMUX g178c2 ( \45886_nG178c2 , \45884_nG178c0 , \45885_nG178c1 , \44829 );
buf \U$37903 ( \45887 , \45886_nG178c2 );
_DC g191d6_GF_IsGateDCbyConstraint ( \45888_nG191d6 , \45887 , \42503 );
buf \U$37904 ( \45889 , \45888_nG191d6 );
_HMUX g178c3 ( \45890_nG178c3 , RIe391c58_6216 , \44870 , \45853 );
_HMUX g178c4 ( \45891_nG178c4 , RIe391c58_6216 , \45890_nG178c3 , \44817 );
_HMUX g178c5 ( \45892_nG178c5 , RIe391c58_6216 , \44873 , \45856 );
_HMUX g178c6 ( \45893_nG178c6 , \45891_nG178c4 , \45892_nG178c5 , \44829 );
buf \U$37905 ( \45894 , \45893_nG178c6 );
_DC g191ec_GF_IsGateDCbyConstraint ( \45895_nG191ec , \45894 , \42503 );
buf \U$37906 ( \45896 , \45895_nG191ec );
_HMUX g178c7 ( \45897_nG178c7 , RIe38f5e8_6217 , \44879 , \45853 );
_HMUX g178c8 ( \45898_nG178c8 , RIe38f5e8_6217 , \45897_nG178c7 , \44817 );
_HMUX g178c9 ( \45899_nG178c9 , RIe38f5e8_6217 , \44882 , \45856 );
_HMUX g178ca ( \45900_nG178ca , \45898_nG178c8 , \45899_nG178c9 , \44829 );
buf \U$37907 ( \45901 , \45900_nG178ca );
_DC g191f8_GF_IsGateDCbyConstraint ( \45902_nG191f8 , \45901 , \42503 );
buf \U$37908 ( \45903 , \45902_nG191f8 );
_HMUX g178cb ( \45904_nG178cb , RIe38d428_6218 , \44888 , \45853 );
_HMUX g178cc ( \45905_nG178cc , RIe38d428_6218 , \45904_nG178cb , \44817 );
_HMUX g178cd ( \45906_nG178cd , RIe38d428_6218 , \44891 , \45856 );
_HMUX g178ce ( \45907_nG178ce , \45905_nG178cc , \45906_nG178cd , \44829 );
buf \U$37909 ( \45908 , \45907_nG178ce );
_DC g191fa_GF_IsGateDCbyConstraint ( \45909_nG191fa , \45908 , \42503 );
buf \U$37910 ( \45910 , \45909_nG191fa );
_HMUX g178cf ( \45911_nG178cf , RIe38ae30_6219 , \44897 , \45853 );
_HMUX g178d0 ( \45912_nG178d0 , RIe38ae30_6219 , \45911_nG178cf , \44817 );
_HMUX g178d1 ( \45913_nG178d1 , RIe38ae30_6219 , \44900 , \45856 );
_HMUX g178d2 ( \45914_nG178d2 , \45912_nG178d0 , \45913_nG178d1 , \44829 );
buf \U$37911 ( \45915 , \45914_nG178d2 );
_DC g191fc_GF_IsGateDCbyConstraint ( \45916_nG191fc , \45915 , \42503 );
buf \U$37912 ( \45917 , \45916_nG191fc );
_HMUX g178d3 ( \45918_nG178d3 , RIe389030_6220 , \44906 , \45853 );
_HMUX g178d4 ( \45919_nG178d4 , RIe389030_6220 , \45918_nG178d3 , \44817 );
_HMUX g178d5 ( \45920_nG178d5 , RIe389030_6220 , \44909 , \45856 );
_HMUX g178d6 ( \45921_nG178d6 , \45919_nG178d4 , \45920_nG178d5 , \44829 );
buf \U$37913 ( \45922 , \45921_nG178d6 );
_DC g19180_GF_IsGateDCbyConstraint ( \45923_nG19180 , \45922 , \42503 );
buf \U$37914 ( \45924 , \45923_nG19180 );
_HMUX g178d7 ( \45925_nG178d7 , RIe386fd8_6221 , \44915 , \45853 );
_HMUX g178d8 ( \45926_nG178d8 , RIe386fd8_6221 , \45925_nG178d7 , \44817 );
_HMUX g178d9 ( \45927_nG178d9 , RIe386fd8_6221 , \44918 , \45856 );
_HMUX g178da ( \45928_nG178da , \45926_nG178d8 , \45927_nG178d9 , \44829 );
buf \U$37915 ( \45929 , \45928_nG178da );
_DC g19182_GF_IsGateDCbyConstraint ( \45930_nG19182 , \45929 , \42503 );
buf \U$37916 ( \45931 , \45930_nG19182 );
_HMUX g178db ( \45932_nG178db , RIe384ff8_6222 , \44924 , \45853 );
_HMUX g178dc ( \45933_nG178dc , RIe384ff8_6222 , \45932_nG178db , \44817 );
_HMUX g178dd ( \45934_nG178dd , RIe384ff8_6222 , \44927 , \45856 );
_HMUX g178de ( \45935_nG178de , \45933_nG178dc , \45934_nG178dd , \44829 );
buf \U$37917 ( \45936 , \45935_nG178de );
_DC g19184_GF_IsGateDCbyConstraint ( \45937_nG19184 , \45936 , \42503 );
buf \U$37918 ( \45938 , \45937_nG19184 );
_HMUX g178df ( \45939_nG178df , RIe3832e8_6223 , \44933 , \45853 );
_HMUX g178e0 ( \45940_nG178e0 , RIe3832e8_6223 , \45939_nG178df , \44817 );
_HMUX g178e1 ( \45941_nG178e1 , RIe3832e8_6223 , \44936 , \45856 );
_HMUX g178e2 ( \45942_nG178e2 , \45940_nG178e0 , \45941_nG178e1 , \44829 );
buf \U$37919 ( \45943 , \45942_nG178e2 );
_DC g19186_GF_IsGateDCbyConstraint ( \45944_nG19186 , \45943 , \42503 );
buf \U$37920 ( \45945 , \45944_nG19186 );
_HMUX g178e3 ( \45946_nG178e3 , RIe381218_6224 , \44942 , \45853 );
_HMUX g178e4 ( \45947_nG178e4 , RIe381218_6224 , \45946_nG178e3 , \44817 );
_HMUX g178e5 ( \45948_nG178e5 , RIe381218_6224 , \44945 , \45856 );
_HMUX g178e6 ( \45949_nG178e6 , \45947_nG178e4 , \45948_nG178e5 , \44829 );
buf \U$37921 ( \45950 , \45949_nG178e6 );
_DC g19188_GF_IsGateDCbyConstraint ( \45951_nG19188 , \45950 , \42503 );
buf \U$37922 ( \45952 , \45951_nG19188 );
_HMUX g178e7 ( \45953_nG178e7 , RIe37f148_6225 , \44951 , \45853 );
_HMUX g178e8 ( \45954_nG178e8 , RIe37f148_6225 , \45953_nG178e7 , \44817 );
_HMUX g178e9 ( \45955_nG178e9 , RIe37f148_6225 , \44954 , \45856 );
_HMUX g178ea ( \45956_nG178ea , \45954_nG178e8 , \45955_nG178e9 , \44829 );
buf \U$37923 ( \45957 , \45956_nG178ea );
_DC g1918a_GF_IsGateDCbyConstraint ( \45958_nG1918a , \45957 , \42503 );
buf \U$37924 ( \45959 , \45958_nG1918a );
_HMUX g178eb ( \45960_nG178eb , RIe37ce20_6226 , \44960 , \45853 );
_HMUX g178ec ( \45961_nG178ec , RIe37ce20_6226 , \45960_nG178eb , \44817 );
_HMUX g178ed ( \45962_nG178ed , RIe37ce20_6226 , \44963 , \45856 );
_HMUX g178ee ( \45963_nG178ee , \45961_nG178ec , \45962_nG178ed , \44829 );
buf \U$37925 ( \45964 , \45963_nG178ee );
_DC g1918c_GF_IsGateDCbyConstraint ( \45965_nG1918c , \45964 , \42503 );
buf \U$37926 ( \45966 , \45965_nG1918c );
_HMUX g178ef ( \45967_nG178ef , RIe37aeb8_6227 , \44969 , \45853 );
_HMUX g178f0 ( \45968_nG178f0 , RIe37aeb8_6227 , \45967_nG178ef , \44817 );
_HMUX g178f1 ( \45969_nG178f1 , RIe37aeb8_6227 , \44972 , \45856 );
_HMUX g178f2 ( \45970_nG178f2 , \45968_nG178f0 , \45969_nG178f1 , \44829 );
buf \U$37927 ( \45971 , \45970_nG178f2 );
_DC g1918e_GF_IsGateDCbyConstraint ( \45972_nG1918e , \45971 , \42503 );
buf \U$37928 ( \45973 , \45972_nG1918e );
_HMUX g178f3 ( \45974_nG178f3 , RIe378668_6228 , \44978 , \45853 );
_HMUX g178f4 ( \45975_nG178f4 , RIe378668_6228 , \45974_nG178f3 , \44817 );
_HMUX g178f5 ( \45976_nG178f5 , RIe378668_6228 , \44981 , \45856 );
_HMUX g178f6 ( \45977_nG178f6 , \45975_nG178f4 , \45976_nG178f5 , \44829 );
buf \U$37929 ( \45978 , \45977_nG178f6 );
_DC g19190_GF_IsGateDCbyConstraint ( \45979_nG19190 , \45978 , \42503 );
buf \U$37930 ( \45980 , \45979_nG19190 );
_HMUX g178f7 ( \45981_nG178f7 , RIe3755a8_6229 , \44987 , \45853 );
_HMUX g178f8 ( \45982_nG178f8 , RIe3755a8_6229 , \45981_nG178f7 , \44817 );
_HMUX g178f9 ( \45983_nG178f9 , RIe3755a8_6229 , \44990 , \45856 );
_HMUX g178fa ( \45984_nG178fa , \45982_nG178f8 , \45983_nG178f9 , \44829 );
buf \U$37931 ( \45985 , \45984_nG178fa );
_DC g19192_GF_IsGateDCbyConstraint ( \45986_nG19192 , \45985 , \42503 );
buf \U$37932 ( \45987 , \45986_nG19192 );
_HMUX g178fb ( \45988_nG178fb , RIe372c68_6230 , \44996 , \45853 );
_HMUX g178fc ( \45989_nG178fc , RIe372c68_6230 , \45988_nG178fb , \44817 );
_HMUX g178fd ( \45990_nG178fd , RIe372c68_6230 , \44999 , \45856 );
_HMUX g178fe ( \45991_nG178fe , \45989_nG178fc , \45990_nG178fd , \44829 );
buf \U$37933 ( \45992 , \45991_nG178fe );
_DC g19196_GF_IsGateDCbyConstraint ( \45993_nG19196 , \45992 , \42503 );
buf \U$37934 ( \45994 , \45993_nG19196 );
_HMUX g178ff ( \45995_nG178ff , RIe2703f8_6231 , \45005 , \45853 );
_HMUX g17900 ( \45996_nG17900 , RIe2703f8_6231 , \45995_nG178ff , \44817 );
_HMUX g17901 ( \45997_nG17901 , RIe2703f8_6231 , \45008 , \45856 );
_HMUX g17902 ( \45998_nG17902 , \45996_nG17900 , \45997_nG17901 , \44829 );
buf \U$37935 ( \45999 , \45998_nG17902 );
_DC g19198_GF_IsGateDCbyConstraint ( \46000_nG19198 , \45999 , \42503 );
buf \U$37936 ( \46001 , \46000_nG19198 );
_HMUX g17903 ( \46002_nG17903 , RIe26d4a0_6232 , \45014 , \45853 );
_HMUX g17904 ( \46003_nG17904 , RIe26d4a0_6232 , \46002_nG17903 , \44817 );
_HMUX g17905 ( \46004_nG17905 , RIe26d4a0_6232 , \45017 , \45856 );
_HMUX g17906 ( \46005_nG17906 , \46003_nG17904 , \46004_nG17905 , \44829 );
buf \U$37937 ( \46006 , \46005_nG17906 );
_DC g1919a_GF_IsGateDCbyConstraint ( \46007_nG1919a , \46006 , \42503 );
buf \U$37938 ( \46008 , \46007_nG1919a );
_HMUX g17907 ( \46009_nG17907 , RIe26aae8_6233 , \45023 , \45853 );
_HMUX g17908 ( \46010_nG17908 , RIe26aae8_6233 , \46009_nG17907 , \44817 );
_HMUX g17909 ( \46011_nG17909 , RIe26aae8_6233 , \45026 , \45856 );
_HMUX g1790a ( \46012_nG1790a , \46010_nG17908 , \46011_nG17909 , \44829 );
buf \U$37939 ( \46013 , \46012_nG1790a );
_DC g1919c_GF_IsGateDCbyConstraint ( \46014_nG1919c , \46013 , \42503 );
buf \U$37940 ( \46015 , \46014_nG1919c );
_HMUX g1790b ( \46016_nG1790b , RIe2686d0_6234 , \45032 , \45853 );
_HMUX g1790c ( \46017_nG1790c , RIe2686d0_6234 , \46016_nG1790b , \44817 );
_HMUX g1790d ( \46018_nG1790d , RIe2686d0_6234 , \45035 , \45856 );
_HMUX g1790e ( \46019_nG1790e , \46017_nG1790c , \46018_nG1790d , \44829 );
buf \U$37941 ( \46020 , \46019_nG1790e );
_DC g1919e_GF_IsGateDCbyConstraint ( \46021_nG1919e , \46020 , \42503 );
buf \U$37942 ( \46022 , \46021_nG1919e );
_HMUX g1790f ( \46023_nG1790f , RIe265ca0_6235 , \45041 , \45853 );
_HMUX g17910 ( \46024_nG17910 , RIe265ca0_6235 , \46023_nG1790f , \44817 );
_HMUX g17911 ( \46025_nG17911 , RIe265ca0_6235 , \45044 , \45856 );
_HMUX g17912 ( \46026_nG17912 , \46024_nG17910 , \46025_nG17911 , \44829 );
buf \U$37943 ( \46027 , \46026_nG17912 );
_DC g191a0_GF_IsGateDCbyConstraint ( \46028_nG191a0 , \46027 , \42503 );
buf \U$37944 ( \46029 , \46028_nG191a0 );
_HMUX g17913 ( \46030_nG17913 , RIe264170_6236 , \45050 , \45853 );
_HMUX g17914 ( \46031_nG17914 , RIe264170_6236 , \46030_nG17913 , \44817 );
_HMUX g17915 ( \46032_nG17915 , RIe264170_6236 , \45053 , \45856 );
_HMUX g17916 ( \46033_nG17916 , \46031_nG17914 , \46032_nG17915 , \44829 );
buf \U$37945 ( \46034 , \46033_nG17916 );
_DC g191a2_GF_IsGateDCbyConstraint ( \46035_nG191a2 , \46034 , \42503 );
buf \U$37946 ( \46036 , \46035_nG191a2 );
_HMUX g17917 ( \46037_nG17917 , RIe2616c8_6237 , \45059 , \45853 );
_HMUX g17918 ( \46038_nG17918 , RIe2616c8_6237 , \46037_nG17917 , \44817 );
_HMUX g17919 ( \46039_nG17919 , RIe2616c8_6237 , \45062 , \45856 );
_HMUX g1791a ( \46040_nG1791a , \46038_nG17918 , \46039_nG17919 , \44829 );
buf \U$37947 ( \46041 , \46040_nG1791a );
_DC g191a4_GF_IsGateDCbyConstraint ( \46042_nG191a4 , \46041 , \42503 );
buf \U$37948 ( \46043 , \46042_nG191a4 );
_HMUX g1791b ( \46044_nG1791b , RIe25f238_6238 , \45068 , \45853 );
_HMUX g1791c ( \46045_nG1791c , RIe25f238_6238 , \46044_nG1791b , \44817 );
_HMUX g1791d ( \46046_nG1791d , RIe25f238_6238 , \45071 , \45856 );
_HMUX g1791e ( \46047_nG1791e , \46045_nG1791c , \46046_nG1791d , \44829 );
buf \U$37949 ( \46048 , \46047_nG1791e );
_DC g191a6_GF_IsGateDCbyConstraint ( \46049_nG191a6 , \46048 , \42503 );
buf \U$37950 ( \46050 , \46049_nG191a6 );
_HMUX g1791f ( \46051_nG1791f , RIe25c6a0_6239 , \45077 , \45853 );
_HMUX g17920 ( \46052_nG17920 , RIe25c6a0_6239 , \46051_nG1791f , \44817 );
_HMUX g17921 ( \46053_nG17921 , RIe25c6a0_6239 , \45080 , \45856 );
_HMUX g17922 ( \46054_nG17922 , \46052_nG17920 , \46053_nG17921 , \44829 );
buf \U$37951 ( \46055 , \46054_nG17922 );
_DC g191a8_GF_IsGateDCbyConstraint ( \46056_nG191a8 , \46055 , \42503 );
buf \U$37952 ( \46057 , \46056_nG191a8 );
_HMUX g17923 ( \46058_nG17923 , RIe259ec8_6240 , \45086 , \45853 );
_HMUX g17924 ( \46059_nG17924 , RIe259ec8_6240 , \46058_nG17923 , \44817 );
_HMUX g17925 ( \46060_nG17925 , RIe259ec8_6240 , \45089 , \45856 );
_HMUX g17926 ( \46061_nG17926 , \46059_nG17924 , \46060_nG17925 , \44829 );
buf \U$37953 ( \46062 , \46061_nG17926 );
_DC g191ac_GF_IsGateDCbyConstraint ( \46063_nG191ac , \46062 , \42503 );
buf \U$37954 ( \46064 , \46063_nG191ac );
_HMUX g17927 ( \46065_nG17927 , RIe257240_6241 , \45095 , \45853 );
_HMUX g17928 ( \46066_nG17928 , RIe257240_6241 , \46065_nG17927 , \44817 );
_HMUX g17929 ( \46067_nG17929 , RIe257240_6241 , \45098 , \45856 );
_HMUX g1792a ( \46068_nG1792a , \46066_nG17928 , \46067_nG17929 , \44829 );
buf \U$37955 ( \46069 , \46068_nG1792a );
_DC g191ae_GF_IsGateDCbyConstraint ( \46070_nG191ae , \46069 , \42503 );
buf \U$37956 ( \46071 , \46070_nG191ae );
_HMUX g1792b ( \46072_nG1792b , RIe254018_6242 , \45104 , \45853 );
_HMUX g1792c ( \46073_nG1792c , RIe254018_6242 , \46072_nG1792b , \44817 );
_HMUX g1792d ( \46074_nG1792d , RIe254018_6242 , \45107 , \45856 );
_HMUX g1792e ( \46075_nG1792e , \46073_nG1792c , \46074_nG1792d , \44829 );
buf \U$37957 ( \46076 , \46075_nG1792e );
_DC g191b0_GF_IsGateDCbyConstraint ( \46077_nG191b0 , \46076 , \42503 );
buf \U$37958 ( \46078 , \46077_nG191b0 );
_HMUX g1792f ( \46079_nG1792f , RIe251408_6243 , \45113 , \45853 );
_HMUX g17930 ( \46080_nG17930 , RIe251408_6243 , \46079_nG1792f , \44817 );
_HMUX g17931 ( \46081_nG17931 , RIe251408_6243 , \45116 , \45856 );
_HMUX g17932 ( \46082_nG17932 , \46080_nG17930 , \46081_nG17931 , \44829 );
buf \U$37959 ( \46083 , \46082_nG17932 );
_DC g191b2_GF_IsGateDCbyConstraint ( \46084_nG191b2 , \46083 , \42503 );
buf \U$37960 ( \46085 , \46084_nG191b2 );
_HMUX g17933 ( \46086_nG17933 , RIe24e8e8_6244 , \45122 , \45853 );
_HMUX g17934 ( \46087_nG17934 , RIe24e8e8_6244 , \46086_nG17933 , \44817 );
_HMUX g17935 ( \46088_nG17935 , RIe24e8e8_6244 , \45125 , \45856 );
_HMUX g17936 ( \46089_nG17936 , \46087_nG17934 , \46088_nG17935 , \44829 );
buf \U$37961 ( \46090 , \46089_nG17936 );
_DC g191b4_GF_IsGateDCbyConstraint ( \46091_nG191b4 , \46090 , \42503 );
buf \U$37962 ( \46092 , \46091_nG191b4 );
_HMUX g17937 ( \46093_nG17937 , RIe24c110_6245 , \45131 , \45853 );
_HMUX g17938 ( \46094_nG17938 , RIe24c110_6245 , \46093_nG17937 , \44817 );
_HMUX g17939 ( \46095_nG17939 , RIe24c110_6245 , \45134 , \45856 );
_HMUX g1793a ( \46096_nG1793a , \46094_nG17938 , \46095_nG17939 , \44829 );
buf \U$37963 ( \46097 , \46096_nG1793a );
_DC g191b6_GF_IsGateDCbyConstraint ( \46098_nG191b6 , \46097 , \42503 );
buf \U$37964 ( \46099 , \46098_nG191b6 );
_HMUX g1793b ( \46100_nG1793b , RIe248d08_6246 , \45140 , \45853 );
_HMUX g1793c ( \46101_nG1793c , RIe248d08_6246 , \46100_nG1793b , \44817 );
_HMUX g1793d ( \46102_nG1793d , RIe248d08_6246 , \45143 , \45856 );
_HMUX g1793e ( \46103_nG1793e , \46101_nG1793c , \46102_nG1793d , \44829 );
buf \U$37965 ( \46104 , \46103_nG1793e );
_DC g191b8_GF_IsGateDCbyConstraint ( \46105_nG191b8 , \46104 , \42503 );
buf \U$37966 ( \46106 , \46105_nG191b8 );
_HMUX g1793f ( \46107_nG1793f , RIe246170_6247 , \45149 , \45853 );
_HMUX g17940 ( \46108_nG17940 , RIe246170_6247 , \46107_nG1793f , \44817 );
_HMUX g17941 ( \46109_nG17941 , RIe246170_6247 , \45152 , \45856 );
_HMUX g17942 ( \46110_nG17942 , \46108_nG17940 , \46109_nG17941 , \44829 );
buf \U$37967 ( \46111 , \46110_nG17942 );
_DC g191ba_GF_IsGateDCbyConstraint ( \46112_nG191ba , \46111 , \42503 );
buf \U$37968 ( \46113 , \46112_nG191ba );
_HMUX g17943 ( \46114_nG17943 , RIe2435d8_6248 , \45158 , \45853 );
_HMUX g17944 ( \46115_nG17944 , RIe2435d8_6248 , \46114_nG17943 , \44817 );
_HMUX g17945 ( \46116_nG17945 , RIe2435d8_6248 , \45161 , \45856 );
_HMUX g17946 ( \46117_nG17946 , \46115_nG17944 , \46116_nG17945 , \44829 );
buf \U$37969 ( \46118 , \46117_nG17946 );
_DC g191bc_GF_IsGateDCbyConstraint ( \46119_nG191bc , \46118 , \42503 );
buf \U$37970 ( \46120 , \46119_nG191bc );
_HMUX g17947 ( \46121_nG17947 , RIe2418c8_6249 , \45167 , \45853 );
_HMUX g17948 ( \46122_nG17948 , RIe2418c8_6249 , \46121_nG17947 , \44817 );
_HMUX g17949 ( \46123_nG17949 , RIe2418c8_6249 , \45170 , \45856 );
_HMUX g1794a ( \46124_nG1794a , \46122_nG17948 , \46123_nG17949 , \44829 );
buf \U$37971 ( \46125 , \46124_nG1794a );
_DC g191be_GF_IsGateDCbyConstraint ( \46126_nG191be , \46125 , \42503 );
buf \U$37972 ( \46127 , \46126_nG191be );
_HMUX g1794b ( \46128_nG1794b , RIe23fb40_6250 , \45176 , \45853 );
_HMUX g1794c ( \46129_nG1794c , RIe23fb40_6250 , \46128_nG1794b , \44817 );
_HMUX g1794d ( \46130_nG1794d , RIe23fb40_6250 , \45179 , \45856 );
_HMUX g1794e ( \46131_nG1794e , \46129_nG1794c , \46130_nG1794d , \44829 );
buf \U$37973 ( \46132 , \46131_nG1794e );
_DC g191c2_GF_IsGateDCbyConstraint ( \46133_nG191c2 , \46132 , \42503 );
buf \U$37974 ( \46134 , \46133_nG191c2 );
_HMUX g1794f ( \46135_nG1794f , RIe23dcc8_6251 , \45185 , \45853 );
_HMUX g17950 ( \46136_nG17950 , RIe23dcc8_6251 , \46135_nG1794f , \44817 );
_HMUX g17951 ( \46137_nG17951 , RIe23dcc8_6251 , \45188 , \45856 );
_HMUX g17952 ( \46138_nG17952 , \46136_nG17950 , \46137_nG17951 , \44829 );
buf \U$37975 ( \46139 , \46138_nG17952 );
_DC g191c4_GF_IsGateDCbyConstraint ( \46140_nG191c4 , \46139 , \42503 );
buf \U$37976 ( \46141 , \46140_nG191c4 );
_HMUX g17953 ( \46142_nG17953 , RIe23ba18_6252 , \45194 , \45853 );
_HMUX g17954 ( \46143_nG17954 , RIe23ba18_6252 , \46142_nG17953 , \44817 );
_HMUX g17955 ( \46144_nG17955 , RIe23ba18_6252 , \45197 , \45856 );
_HMUX g17956 ( \46145_nG17956 , \46143_nG17954 , \46144_nG17955 , \44829 );
buf \U$37977 ( \46146 , \46145_nG17956 );
_DC g191c6_GF_IsGateDCbyConstraint ( \46147_nG191c6 , \46146 , \42503 );
buf \U$37978 ( \46148 , \46147_nG191c6 );
_HMUX g17957 ( \46149_nG17957 , RIe239948_6253 , \45203 , \45853 );
_HMUX g17958 ( \46150_nG17958 , RIe239948_6253 , \46149_nG17957 , \44817 );
_HMUX g17959 ( \46151_nG17959 , RIe239948_6253 , \45206 , \45856 );
_HMUX g1795a ( \46152_nG1795a , \46150_nG17958 , \46151_nG17959 , \44829 );
buf \U$37979 ( \46153 , \46152_nG1795a );
_DC g191c8_GF_IsGateDCbyConstraint ( \46154_nG191c8 , \46153 , \42503 );
buf \U$37980 ( \46155 , \46154_nG191c8 );
_HMUX g1795b ( \46156_nG1795b , RIe2381d8_6254 , \45212 , \45853 );
_HMUX g1795c ( \46157_nG1795c , RIe2381d8_6254 , \46156_nG1795b , \44817 );
_HMUX g1795d ( \46158_nG1795d , RIe2381d8_6254 , \45215 , \45856 );
_HMUX g1795e ( \46159_nG1795e , \46157_nG1795c , \46158_nG1795d , \44829 );
buf \U$37981 ( \46160 , \46159_nG1795e );
_DC g191ca_GF_IsGateDCbyConstraint ( \46161_nG191ca , \46160 , \42503 );
buf \U$37982 ( \46162 , \46161_nG191ca );
_HMUX g1795f ( \46163_nG1795f , RIe236720_6255 , \45221 , \45853 );
_HMUX g17960 ( \46164_nG17960 , RIe236720_6255 , \46163_nG1795f , \44817 );
_HMUX g17961 ( \46165_nG17961 , RIe236720_6255 , \45224 , \45856 );
_HMUX g17962 ( \46166_nG17962 , \46164_nG17960 , \46165_nG17961 , \44829 );
buf \U$37983 ( \46167 , \46166_nG17962 );
_DC g191cc_GF_IsGateDCbyConstraint ( \46168_nG191cc , \46167 , \42503 );
buf \U$37984 ( \46169 , \46168_nG191cc );
_HMUX g17963 ( \46170_nG17963 , RIe2346c8_6256 , \45230 , \45853 );
_HMUX g17964 ( \46171_nG17964 , RIe2346c8_6256 , \46170_nG17963 , \44817 );
_HMUX g17965 ( \46172_nG17965 , RIe2346c8_6256 , \45233 , \45856 );
_HMUX g17966 ( \46173_nG17966 , \46171_nG17964 , \46172_nG17965 , \44829 );
buf \U$37985 ( \46174 , \46173_nG17966 );
_DC g191ce_GF_IsGateDCbyConstraint ( \46175_nG191ce , \46174 , \42503 );
buf \U$37986 ( \46176 , \46175_nG191ce );
_HMUX g17967 ( \46177_nG17967 , RIe232a30_6257 , \45239 , \45853 );
_HMUX g17968 ( \46178_nG17968 , RIe232a30_6257 , \46177_nG17967 , \44817 );
_HMUX g17969 ( \46179_nG17969 , RIe232a30_6257 , \45242 , \45856 );
_HMUX g1796a ( \46180_nG1796a , \46178_nG17968 , \46179_nG17969 , \44829 );
buf \U$37987 ( \46181 , \46180_nG1796a );
_DC g191d0_GF_IsGateDCbyConstraint ( \46182_nG191d0 , \46181 , \42503 );
buf \U$37988 ( \46183 , \46182_nG191d0 );
_HMUX g1796b ( \46184_nG1796b , RIe230bb8_6258 , \45248 , \45853 );
_HMUX g1796c ( \46185_nG1796c , RIe230bb8_6258 , \46184_nG1796b , \44817 );
_HMUX g1796d ( \46186_nG1796d , RIe230bb8_6258 , \45251 , \45856 );
_HMUX g1796e ( \46187_nG1796e , \46185_nG1796c , \46186_nG1796d , \44829 );
buf \U$37989 ( \46188 , \46187_nG1796e );
_DC g191d2_GF_IsGateDCbyConstraint ( \46189_nG191d2 , \46188 , \42503 );
buf \U$37990 ( \46190 , \46189_nG191d2 );
_HMUX g1796f ( \46191_nG1796f , RIe465cb0_6259 , \45257 , \45853 );
_HMUX g17970 ( \46192_nG17970 , RIe465cb0_6259 , \46191_nG1796f , \44817 );
_HMUX g17971 ( \46193_nG17971 , RIe465cb0_6259 , \45260 , \45856 );
_HMUX g17972 ( \46194_nG17972 , \46192_nG17970 , \46193_nG17971 , \44829 );
buf \U$37991 ( \46195 , \46194_nG17972 );
_DC g191d4_GF_IsGateDCbyConstraint ( \46196_nG191d4 , \46195 , \42503 );
buf \U$37992 ( \46197 , \46196_nG191d4 );
_HMUX g17973 ( \46198_nG17973 , RIe4664a8_6260 , \45266 , \45853 );
_HMUX g17974 ( \46199_nG17974 , RIe4664a8_6260 , \46198_nG17973 , \44817 );
_HMUX g17975 ( \46200_nG17975 , RIe4664a8_6260 , \45269 , \45856 );
_HMUX g17976 ( \46201_nG17976 , \46199_nG17974 , \46200_nG17975 , \44829 );
buf \U$37993 ( \46202 , \46201_nG17976 );
_DC g191d8_GF_IsGateDCbyConstraint ( \46203_nG191d8 , \46202 , \42503 );
buf \U$37994 ( \46204 , \46203_nG191d8 );
_HMUX g17977 ( \46205_nG17977 , RIe466ca0_6261 , \45275 , \45853 );
_HMUX g17978 ( \46206_nG17978 , RIe466ca0_6261 , \46205_nG17977 , \44817 );
_HMUX g17979 ( \46207_nG17979 , RIe466ca0_6261 , \45278 , \45856 );
_HMUX g1797a ( \46208_nG1797a , \46206_nG17978 , \46207_nG17979 , \44829 );
buf \U$37995 ( \46209 , \46208_nG1797a );
_DC g191da_GF_IsGateDCbyConstraint ( \46210_nG191da , \46209 , \42503 );
buf \U$37996 ( \46211 , \46210_nG191da );
_HMUX g1797b ( \46212_nG1797b , RIe467498_6262 , \45284 , \45853 );
_HMUX g1797c ( \46213_nG1797c , RIe467498_6262 , \46212_nG1797b , \44817 );
_HMUX g1797d ( \46214_nG1797d , RIe467498_6262 , \45287 , \45856 );
_HMUX g1797e ( \46215_nG1797e , \46213_nG1797c , \46214_nG1797d , \44829 );
buf \U$37997 ( \46216 , \46215_nG1797e );
_DC g191dc_GF_IsGateDCbyConstraint ( \46217_nG191dc , \46216 , \42503 );
buf \U$37998 ( \46218 , \46217_nG191dc );
_HMUX g1797f ( \46219_nG1797f , RIe467c90_6263 , \45293 , \45853 );
_HMUX g17980 ( \46220_nG17980 , RIe467c90_6263 , \46219_nG1797f , \44817 );
_HMUX g17981 ( \46221_nG17981 , RIe467c90_6263 , \45296 , \45856 );
_HMUX g17982 ( \46222_nG17982 , \46220_nG17980 , \46221_nG17981 , \44829 );
buf \U$37999 ( \46223 , \46222_nG17982 );
_DC g191de_GF_IsGateDCbyConstraint ( \46224_nG191de , \46223 , \42503 );
buf \U$38000 ( \46225 , \46224_nG191de );
_HMUX g17983 ( \46226_nG17983 , RIe468488_6264 , \45302 , \45853 );
_HMUX g17984 ( \46227_nG17984 , RIe468488_6264 , \46226_nG17983 , \44817 );
_HMUX g17985 ( \46228_nG17985 , RIe468488_6264 , \45305 , \45856 );
_HMUX g17986 ( \46229_nG17986 , \46227_nG17984 , \46228_nG17985 , \44829 );
buf \U$38001 ( \46230 , \46229_nG17986 );
_DC g191e0_GF_IsGateDCbyConstraint ( \46231_nG191e0 , \46230 , \42503 );
buf \U$38002 ( \46232 , \46231_nG191e0 );
_HMUX g17987 ( \46233_nG17987 , RIe468c80_6265 , \45311 , \45853 );
_HMUX g17988 ( \46234_nG17988 , RIe468c80_6265 , \46233_nG17987 , \44817 );
_HMUX g17989 ( \46235_nG17989 , RIe468c80_6265 , \45314 , \45856 );
_HMUX g1798a ( \46236_nG1798a , \46234_nG17988 , \46235_nG17989 , \44829 );
buf \U$38003 ( \46237 , \46236_nG1798a );
_DC g191e2_GF_IsGateDCbyConstraint ( \46238_nG191e2 , \46237 , \42503 );
buf \U$38004 ( \46239 , \46238_nG191e2 );
_HMUX g1798b ( \46240_nG1798b , RIe469478_6266 , \45320 , \45853 );
_HMUX g1798c ( \46241_nG1798c , RIe469478_6266 , \46240_nG1798b , \44817 );
_HMUX g1798d ( \46242_nG1798d , RIe469478_6266 , \45323 , \45856 );
_HMUX g1798e ( \46243_nG1798e , \46241_nG1798c , \46242_nG1798d , \44829 );
buf \U$38005 ( \46244 , \46243_nG1798e );
_DC g191e4_GF_IsGateDCbyConstraint ( \46245_nG191e4 , \46244 , \42503 );
buf \U$38006 ( \46246 , \46245_nG191e4 );
_HMUX g1798f ( \46247_nG1798f , RIe469c70_6267 , \45329 , \45853 );
_HMUX g17990 ( \46248_nG17990 , RIe469c70_6267 , \46247_nG1798f , \44817 );
_HMUX g17991 ( \46249_nG17991 , RIe469c70_6267 , \45332 , \45856 );
_HMUX g17992 ( \46250_nG17992 , \46248_nG17990 , \46249_nG17991 , \44829 );
buf \U$38007 ( \46251 , \46250_nG17992 );
_DC g191e6_GF_IsGateDCbyConstraint ( \46252_nG191e6 , \46251 , \42503 );
buf \U$38008 ( \46253 , \46252_nG191e6 );
_HMUX g17993 ( \46254_nG17993 , RIe46a468_6268 , \45338 , \45853 );
_HMUX g17994 ( \46255_nG17994 , RIe46a468_6268 , \46254_nG17993 , \44817 );
_HMUX g17995 ( \46256_nG17995 , RIe46a468_6268 , \45341 , \45856 );
_HMUX g17996 ( \46257_nG17996 , \46255_nG17994 , \46256_nG17995 , \44829 );
buf \U$38009 ( \46258 , \46257_nG17996 );
_DC g191e8_GF_IsGateDCbyConstraint ( \46259_nG191e8 , \46258 , \42503 );
buf \U$38010 ( \46260 , \46259_nG191e8 );
_HMUX g17997 ( \46261_nG17997 , RIe46ac60_6269 , \45347 , \45853 );
_HMUX g17998 ( \46262_nG17998 , RIe46ac60_6269 , \46261_nG17997 , \44817 );
_HMUX g17999 ( \46263_nG17999 , RIe46ac60_6269 , \45350 , \45856 );
_HMUX g1799a ( \46264_nG1799a , \46262_nG17998 , \46263_nG17999 , \44829 );
buf \U$38011 ( \46265 , \46264_nG1799a );
_DC g191ea_GF_IsGateDCbyConstraint ( \46266_nG191ea , \46265 , \42503 );
buf \U$38012 ( \46267 , \46266_nG191ea );
_HMUX g1799b ( \46268_nG1799b , RIe46b458_6270 , \45356 , \45853 );
_HMUX g1799c ( \46269_nG1799c , RIe46b458_6270 , \46268_nG1799b , \44817 );
_HMUX g1799d ( \46270_nG1799d , RIe46b458_6270 , \45359 , \45856 );
_HMUX g1799e ( \46271_nG1799e , \46269_nG1799c , \46270_nG1799d , \44829 );
buf \U$38013 ( \46272 , \46271_nG1799e );
_DC g191ee_GF_IsGateDCbyConstraint ( \46273_nG191ee , \46272 , \42503 );
buf \U$38014 ( \46274 , \46273_nG191ee );
_HMUX g1799f ( \46275_nG1799f , RIe46bc50_6271 , \45365 , \45853 );
_HMUX g179a0 ( \46276_nG179a0 , RIe46bc50_6271 , \46275_nG1799f , \44817 );
_HMUX g179a1 ( \46277_nG179a1 , RIe46bc50_6271 , \45368 , \45856 );
_HMUX g179a2 ( \46278_nG179a2 , \46276_nG179a0 , \46277_nG179a1 , \44829 );
buf \U$38015 ( \46279 , \46278_nG179a2 );
_DC g191f0_GF_IsGateDCbyConstraint ( \46280_nG191f0 , \46279 , \42503 );
buf \U$38016 ( \46281 , \46280_nG191f0 );
_HMUX g179a3 ( \46282_nG179a3 , RIe46c448_6272 , \45374 , \45853 );
_HMUX g179a4 ( \46283_nG179a4 , RIe46c448_6272 , \46282_nG179a3 , \44817 );
_HMUX g179a5 ( \46284_nG179a5 , RIe46c448_6272 , \45377 , \45856 );
_HMUX g179a6 ( \46285_nG179a6 , \46283_nG179a4 , \46284_nG179a5 , \44829 );
buf \U$38017 ( \46286 , \46285_nG179a6 );
_DC g191f2_GF_IsGateDCbyConstraint ( \46287_nG191f2 , \46286 , \42503 );
buf \U$38018 ( \46288 , \46287_nG191f2 );
_HMUX g179a7 ( \46289_nG179a7 , RIe46cc40_6273 , \45383 , \45853 );
_HMUX g179a8 ( \46290_nG179a8 , RIe46cc40_6273 , \46289_nG179a7 , \44817 );
_HMUX g179a9 ( \46291_nG179a9 , RIe46cc40_6273 , \45386 , \45856 );
_HMUX g179aa ( \46292_nG179aa , \46290_nG179a8 , \46291_nG179a9 , \44829 );
buf \U$38019 ( \46293 , \46292_nG179aa );
_DC g191f4_GF_IsGateDCbyConstraint ( \46294_nG191f4 , \46293 , \42503 );
buf \U$38020 ( \46295 , \46294_nG191f4 );
_HMUX g179ab ( \46296_nG179ab , RIe46d438_6274 , \45392 , \45853 );
_HMUX g179ac ( \46297_nG179ac , RIe46d438_6274 , \46296_nG179ab , \44817 );
_HMUX g179ad ( \46298_nG179ad , RIe46d438_6274 , \45395 , \45856 );
_HMUX g179ae ( \46299_nG179ae , \46297_nG179ac , \46298_nG179ad , \44829 );
buf \U$38021 ( \46300 , \46299_nG179ae );
_DC g191f6_GF_IsGateDCbyConstraint ( \46301_nG191f6 , \46300 , \42503 );
buf \U$38022 ( \46302 , \46301_nG191f6 );
and \U$38023 ( \46303 , \44808 , \44809 );
_HMUX g1772b ( \46304_nG1772b , RIe46dc30_6275 , \44807 , \46303 );
_HMUX g1772c ( \46305_nG1772c , RIe46dc30_6275 , \46304_nG1772b , \44817 );
and \U$38024 ( \46306 , \44820 , \44821 );
_HMUX g17731 ( \46307_nG17731 , RIe46dc30_6275 , \44819 , \46306 );
_HMUX g17732 ( \46308_nG17732 , \46305_nG1772c , \46307_nG17731 , \44829 );
buf \U$38025 ( \46309 , \46308_nG17732 );
_DC g190fe_GF_IsGateDCbyConstraint ( \46310_nG190fe , \46309 , \42503 );
buf \U$38026 ( \46311 , \46310_nG190fe );
_HMUX g17734 ( \46312_nG17734 , RIe46e428_6276 , \44834 , \46303 );
_HMUX g17735 ( \46313_nG17735 , RIe46e428_6276 , \46312_nG17734 , \44817 );
_HMUX g17737 ( \46314_nG17737 , RIe46e428_6276 , \44837 , \46306 );
_HMUX g17738 ( \46315_nG17738 , \46313_nG17735 , \46314_nG17737 , \44829 );
buf \U$38027 ( \46316 , \46315_nG17738 );
_DC g19114_GF_IsGateDCbyConstraint ( \46317_nG19114 , \46316 , \42503 );
buf \U$38028 ( \46318 , \46317_nG19114 );
_HMUX g1773a ( \46319_nG1773a , RIe46ec20_6277 , \44843 , \46303 );
_HMUX g1773b ( \46320_nG1773b , RIe46ec20_6277 , \46319_nG1773a , \44817 );
_HMUX g1773d ( \46321_nG1773d , RIe46ec20_6277 , \44846 , \46306 );
_HMUX g1773e ( \46322_nG1773e , \46320_nG1773b , \46321_nG1773d , \44829 );
buf \U$38029 ( \46323 , \46322_nG1773e );
_DC g1912a_GF_IsGateDCbyConstraint ( \46324_nG1912a , \46323 , \42503 );
buf \U$38030 ( \46325 , \46324_nG1912a );
_HMUX g17740 ( \46326_nG17740 , RIe46f418_6278 , \44852 , \46303 );
_HMUX g17741 ( \46327_nG17741 , RIe46f418_6278 , \46326_nG17740 , \44817 );
_HMUX g17743 ( \46328_nG17743 , RIe46f418_6278 , \44855 , \46306 );
_HMUX g17744 ( \46329_nG17744 , \46327_nG17741 , \46328_nG17743 , \44829 );
buf \U$38031 ( \46330 , \46329_nG17744 );
_DC g19140_GF_IsGateDCbyConstraint ( \46331_nG19140 , \46330 , \42503 );
buf \U$38032 ( \46332 , \46331_nG19140 );
_HMUX g17746 ( \46333_nG17746 , RIe46fc10_6279 , \44861 , \46303 );
_HMUX g17747 ( \46334_nG17747 , RIe46fc10_6279 , \46333_nG17746 , \44817 );
_HMUX g17749 ( \46335_nG17749 , RIe46fc10_6279 , \44864 , \46306 );
_HMUX g1774a ( \46336_nG1774a , \46334_nG17747 , \46335_nG17749 , \44829 );
buf \U$38033 ( \46337 , \46336_nG1774a );
_DC g19156_GF_IsGateDCbyConstraint ( \46338_nG19156 , \46337 , \42503 );
buf \U$38034 ( \46339 , \46338_nG19156 );
_HMUX g1774c ( \46340_nG1774c , RIe470408_6280 , \44870 , \46303 );
_HMUX g1774d ( \46341_nG1774d , RIe470408_6280 , \46340_nG1774c , \44817 );
_HMUX g1774f ( \46342_nG1774f , RIe470408_6280 , \44873 , \46306 );
_HMUX g17750 ( \46343_nG17750 , \46341_nG1774d , \46342_nG1774f , \44829 );
buf \U$38035 ( \46344 , \46343_nG17750 );
_DC g1916c_GF_IsGateDCbyConstraint ( \46345_nG1916c , \46344 , \42503 );
buf \U$38036 ( \46346 , \46345_nG1916c );
_HMUX g17752 ( \46347_nG17752 , RIe470c00_6281 , \44879 , \46303 );
_HMUX g17753 ( \46348_nG17753 , RIe470c00_6281 , \46347_nG17752 , \44817 );
_HMUX g17755 ( \46349_nG17755 , RIe470c00_6281 , \44882 , \46306 );
_HMUX g17756 ( \46350_nG17756 , \46348_nG17753 , \46349_nG17755 , \44829 );
buf \U$38037 ( \46351 , \46350_nG17756 );
_DC g19178_GF_IsGateDCbyConstraint ( \46352_nG19178 , \46351 , \42503 );
buf \U$38038 ( \46353 , \46352_nG19178 );
_HMUX g17758 ( \46354_nG17758 , RIe4713f8_6282 , \44888 , \46303 );
_HMUX g17759 ( \46355_nG17759 , RIe4713f8_6282 , \46354_nG17758 , \44817 );
_HMUX g1775b ( \46356_nG1775b , RIe4713f8_6282 , \44891 , \46306 );
_HMUX g1775c ( \46357_nG1775c , \46355_nG17759 , \46356_nG1775b , \44829 );
buf \U$38039 ( \46358 , \46357_nG1775c );
_DC g1917a_GF_IsGateDCbyConstraint ( \46359_nG1917a , \46358 , \42503 );
buf \U$38040 ( \46360 , \46359_nG1917a );
_HMUX g1775e ( \46361_nG1775e , RIe471bf0_6283 , \44897 , \46303 );
_HMUX g1775f ( \46362_nG1775f , RIe471bf0_6283 , \46361_nG1775e , \44817 );
_HMUX g17761 ( \46363_nG17761 , RIe471bf0_6283 , \44900 , \46306 );
_HMUX g17762 ( \46364_nG17762 , \46362_nG1775f , \46363_nG17761 , \44829 );
buf \U$38041 ( \46365 , \46364_nG17762 );
_DC g1917c_GF_IsGateDCbyConstraint ( \46366_nG1917c , \46365 , \42503 );
buf \U$38042 ( \46367 , \46366_nG1917c );
_HMUX g17764 ( \46368_nG17764 , RIe4723e8_6284 , \44906 , \46303 );
_HMUX g17765 ( \46369_nG17765 , RIe4723e8_6284 , \46368_nG17764 , \44817 );
_HMUX g17767 ( \46370_nG17767 , RIe4723e8_6284 , \44909 , \46306 );
_HMUX g17768 ( \46371_nG17768 , \46369_nG17765 , \46370_nG17767 , \44829 );
buf \U$38043 ( \46372 , \46371_nG17768 );
_DC g19100_GF_IsGateDCbyConstraint ( \46373_nG19100 , \46372 , \42503 );
buf \U$38044 ( \46374 , \46373_nG19100 );
_HMUX g1776a ( \46375_nG1776a , RIe472bf8_6285 , \44915 , \46303 );
_HMUX g1776b ( \46376_nG1776b , RIe472bf8_6285 , \46375_nG1776a , \44817 );
_HMUX g1776d ( \46377_nG1776d , RIe472bf8_6285 , \44918 , \46306 );
_HMUX g1776e ( \46378_nG1776e , \46376_nG1776b , \46377_nG1776d , \44829 );
buf \U$38045 ( \46379 , \46378_nG1776e );
_DC g19102_GF_IsGateDCbyConstraint ( \46380_nG19102 , \46379 , \42503 );
buf \U$38046 ( \46381 , \46380_nG19102 );
_HMUX g17770 ( \46382_nG17770 , RIe4733f0_6286 , \44924 , \46303 );
_HMUX g17771 ( \46383_nG17771 , RIe4733f0_6286 , \46382_nG17770 , \44817 );
_HMUX g17773 ( \46384_nG17773 , RIe4733f0_6286 , \44927 , \46306 );
_HMUX g17774 ( \46385_nG17774 , \46383_nG17771 , \46384_nG17773 , \44829 );
buf \U$38047 ( \46386 , \46385_nG17774 );
_DC g19104_GF_IsGateDCbyConstraint ( \46387_nG19104 , \46386 , \42503 );
buf \U$38048 ( \46388 , \46387_nG19104 );
_HMUX g17776 ( \46389_nG17776 , RIe473be8_6287 , \44933 , \46303 );
_HMUX g17777 ( \46390_nG17777 , RIe473be8_6287 , \46389_nG17776 , \44817 );
_HMUX g17779 ( \46391_nG17779 , RIe473be8_6287 , \44936 , \46306 );
_HMUX g1777a ( \46392_nG1777a , \46390_nG17777 , \46391_nG17779 , \44829 );
buf \U$38049 ( \46393 , \46392_nG1777a );
_DC g19106_GF_IsGateDCbyConstraint ( \46394_nG19106 , \46393 , \42503 );
buf \U$38050 ( \46395 , \46394_nG19106 );
_HMUX g1777c ( \46396_nG1777c , RIe4743e0_6288 , \44942 , \46303 );
_HMUX g1777d ( \46397_nG1777d , RIe4743e0_6288 , \46396_nG1777c , \44817 );
_HMUX g1777f ( \46398_nG1777f , RIe4743e0_6288 , \44945 , \46306 );
_HMUX g17780 ( \46399_nG17780 , \46397_nG1777d , \46398_nG1777f , \44829 );
buf \U$38051 ( \46400 , \46399_nG17780 );
_DC g19108_GF_IsGateDCbyConstraint ( \46401_nG19108 , \46400 , \42503 );
buf \U$38052 ( \46402 , \46401_nG19108 );
_HMUX g17782 ( \46403_nG17782 , RIe474bd8_6289 , \44951 , \46303 );
_HMUX g17783 ( \46404_nG17783 , RIe474bd8_6289 , \46403_nG17782 , \44817 );
_HMUX g17785 ( \46405_nG17785 , RIe474bd8_6289 , \44954 , \46306 );
_HMUX g17786 ( \46406_nG17786 , \46404_nG17783 , \46405_nG17785 , \44829 );
buf \U$38053 ( \46407 , \46406_nG17786 );
_DC g1910a_GF_IsGateDCbyConstraint ( \46408_nG1910a , \46407 , \42503 );
buf \U$38054 ( \46409 , \46408_nG1910a );
_HMUX g17788 ( \46410_nG17788 , RIe4753d0_6290 , \44960 , \46303 );
_HMUX g17789 ( \46411_nG17789 , RIe4753d0_6290 , \46410_nG17788 , \44817 );
_HMUX g1778b ( \46412_nG1778b , RIe4753d0_6290 , \44963 , \46306 );
_HMUX g1778c ( \46413_nG1778c , \46411_nG17789 , \46412_nG1778b , \44829 );
buf \U$38055 ( \46414 , \46413_nG1778c );
_DC g1910c_GF_IsGateDCbyConstraint ( \46415_nG1910c , \46414 , \42503 );
buf \U$38056 ( \46416 , \46415_nG1910c );
_HMUX g1778e ( \46417_nG1778e , RIe475bc8_6291 , \44969 , \46303 );
_HMUX g1778f ( \46418_nG1778f , RIe475bc8_6291 , \46417_nG1778e , \44817 );
_HMUX g17791 ( \46419_nG17791 , RIe475bc8_6291 , \44972 , \46306 );
_HMUX g17792 ( \46420_nG17792 , \46418_nG1778f , \46419_nG17791 , \44829 );
buf \U$38057 ( \46421 , \46420_nG17792 );
_DC g1910e_GF_IsGateDCbyConstraint ( \46422_nG1910e , \46421 , \42503 );
buf \U$38058 ( \46423 , \46422_nG1910e );
_HMUX g17794 ( \46424_nG17794 , RIe4763c0_6292 , \44978 , \46303 );
_HMUX g17795 ( \46425_nG17795 , RIe4763c0_6292 , \46424_nG17794 , \44817 );
_HMUX g17797 ( \46426_nG17797 , RIe4763c0_6292 , \44981 , \46306 );
_HMUX g17798 ( \46427_nG17798 , \46425_nG17795 , \46426_nG17797 , \44829 );
buf \U$38059 ( \46428 , \46427_nG17798 );
_DC g19110_GF_IsGateDCbyConstraint ( \46429_nG19110 , \46428 , \42503 );
buf \U$38060 ( \46430 , \46429_nG19110 );
_HMUX g1779a ( \46431_nG1779a , RIe476bb8_6293 , \44987 , \46303 );
_HMUX g1779b ( \46432_nG1779b , RIe476bb8_6293 , \46431_nG1779a , \44817 );
_HMUX g1779d ( \46433_nG1779d , RIe476bb8_6293 , \44990 , \46306 );
_HMUX g1779e ( \46434_nG1779e , \46432_nG1779b , \46433_nG1779d , \44829 );
buf \U$38061 ( \46435 , \46434_nG1779e );
_DC g19112_GF_IsGateDCbyConstraint ( \46436_nG19112 , \46435 , \42503 );
buf \U$38062 ( \46437 , \46436_nG19112 );
_HMUX g177a0 ( \46438_nG177a0 , RIe4773b0_6294 , \44996 , \46303 );
_HMUX g177a1 ( \46439_nG177a1 , RIe4773b0_6294 , \46438_nG177a0 , \44817 );
_HMUX g177a3 ( \46440_nG177a3 , RIe4773b0_6294 , \44999 , \46306 );
_HMUX g177a4 ( \46441_nG177a4 , \46439_nG177a1 , \46440_nG177a3 , \44829 );
buf \U$38063 ( \46442 , \46441_nG177a4 );
_DC g19116_GF_IsGateDCbyConstraint ( \46443_nG19116 , \46442 , \42503 );
buf \U$38064 ( \46444 , \46443_nG19116 );
_HMUX g177a6 ( \46445_nG177a6 , RIe477ba8_6295 , \45005 , \46303 );
_HMUX g177a7 ( \46446_nG177a7 , RIe477ba8_6295 , \46445_nG177a6 , \44817 );
_HMUX g177a9 ( \46447_nG177a9 , RIe477ba8_6295 , \45008 , \46306 );
_HMUX g177aa ( \46448_nG177aa , \46446_nG177a7 , \46447_nG177a9 , \44829 );
buf \U$38065 ( \46449 , \46448_nG177aa );
_DC g19118_GF_IsGateDCbyConstraint ( \46450_nG19118 , \46449 , \42503 );
buf \U$38066 ( \46451 , \46450_nG19118 );
_HMUX g177ac ( \46452_nG177ac , RIe4783a0_6296 , \45014 , \46303 );
_HMUX g177ad ( \46453_nG177ad , RIe4783a0_6296 , \46452_nG177ac , \44817 );
_HMUX g177af ( \46454_nG177af , RIe4783a0_6296 , \45017 , \46306 );
_HMUX g177b0 ( \46455_nG177b0 , \46453_nG177ad , \46454_nG177af , \44829 );
buf \U$38067 ( \46456 , \46455_nG177b0 );
_DC g1911a_GF_IsGateDCbyConstraint ( \46457_nG1911a , \46456 , \42503 );
buf \U$38068 ( \46458 , \46457_nG1911a );
_HMUX g177b2 ( \46459_nG177b2 , RIe478b98_6297 , \45023 , \46303 );
_HMUX g177b3 ( \46460_nG177b3 , RIe478b98_6297 , \46459_nG177b2 , \44817 );
_HMUX g177b5 ( \46461_nG177b5 , RIe478b98_6297 , \45026 , \46306 );
_HMUX g177b6 ( \46462_nG177b6 , \46460_nG177b3 , \46461_nG177b5 , \44829 );
buf \U$38069 ( \46463 , \46462_nG177b6 );
_DC g1911c_GF_IsGateDCbyConstraint ( \46464_nG1911c , \46463 , \42503 );
buf \U$38070 ( \46465 , \46464_nG1911c );
_HMUX g177b8 ( \46466_nG177b8 , RIe479390_6298 , \45032 , \46303 );
_HMUX g177b9 ( \46467_nG177b9 , RIe479390_6298 , \46466_nG177b8 , \44817 );
_HMUX g177bb ( \46468_nG177bb , RIe479390_6298 , \45035 , \46306 );
_HMUX g177bc ( \46469_nG177bc , \46467_nG177b9 , \46468_nG177bb , \44829 );
buf \U$38071 ( \46470 , \46469_nG177bc );
_DC g1911e_GF_IsGateDCbyConstraint ( \46471_nG1911e , \46470 , \42503 );
buf \U$38072 ( \46472 , \46471_nG1911e );
_HMUX g177be ( \46473_nG177be , RIe479b88_6299 , \45041 , \46303 );
_HMUX g177bf ( \46474_nG177bf , RIe479b88_6299 , \46473_nG177be , \44817 );
_HMUX g177c1 ( \46475_nG177c1 , RIe479b88_6299 , \45044 , \46306 );
_HMUX g177c2 ( \46476_nG177c2 , \46474_nG177bf , \46475_nG177c1 , \44829 );
buf \U$38073 ( \46477 , \46476_nG177c2 );
_DC g19120_GF_IsGateDCbyConstraint ( \46478_nG19120 , \46477 , \42503 );
buf \U$38074 ( \46479 , \46478_nG19120 );
_HMUX g177c4 ( \46480_nG177c4 , RIe47a380_6300 , \45050 , \46303 );
_HMUX g177c5 ( \46481_nG177c5 , RIe47a380_6300 , \46480_nG177c4 , \44817 );
_HMUX g177c7 ( \46482_nG177c7 , RIe47a380_6300 , \45053 , \46306 );
_HMUX g177c8 ( \46483_nG177c8 , \46481_nG177c5 , \46482_nG177c7 , \44829 );
buf \U$38075 ( \46484 , \46483_nG177c8 );
_DC g19122_GF_IsGateDCbyConstraint ( \46485_nG19122 , \46484 , \42503 );
buf \U$38076 ( \46486 , \46485_nG19122 );
_HMUX g177ca ( \46487_nG177ca , RIe47ab78_6301 , \45059 , \46303 );
_HMUX g177cb ( \46488_nG177cb , RIe47ab78_6301 , \46487_nG177ca , \44817 );
_HMUX g177cd ( \46489_nG177cd , RIe47ab78_6301 , \45062 , \46306 );
_HMUX g177ce ( \46490_nG177ce , \46488_nG177cb , \46489_nG177cd , \44829 );
buf \U$38077 ( \46491 , \46490_nG177ce );
_DC g19124_GF_IsGateDCbyConstraint ( \46492_nG19124 , \46491 , \42503 );
buf \U$38078 ( \46493 , \46492_nG19124 );
_HMUX g177d0 ( \46494_nG177d0 , RIe47b370_6302 , \45068 , \46303 );
_HMUX g177d1 ( \46495_nG177d1 , RIe47b370_6302 , \46494_nG177d0 , \44817 );
_HMUX g177d3 ( \46496_nG177d3 , RIe47b370_6302 , \45071 , \46306 );
_HMUX g177d4 ( \46497_nG177d4 , \46495_nG177d1 , \46496_nG177d3 , \44829 );
buf \U$38079 ( \46498 , \46497_nG177d4 );
_DC g19126_GF_IsGateDCbyConstraint ( \46499_nG19126 , \46498 , \42503 );
buf \U$38080 ( \46500 , \46499_nG19126 );
_HMUX g177d6 ( \46501_nG177d6 , RIe47bb68_6303 , \45077 , \46303 );
_HMUX g177d7 ( \46502_nG177d7 , RIe47bb68_6303 , \46501_nG177d6 , \44817 );
_HMUX g177d9 ( \46503_nG177d9 , RIe47bb68_6303 , \45080 , \46306 );
_HMUX g177da ( \46504_nG177da , \46502_nG177d7 , \46503_nG177d9 , \44829 );
buf \U$38081 ( \46505 , \46504_nG177da );
_DC g19128_GF_IsGateDCbyConstraint ( \46506_nG19128 , \46505 , \42503 );
buf \U$38082 ( \46507 , \46506_nG19128 );
_HMUX g177dc ( \46508_nG177dc , RIe47c360_6304 , \45086 , \46303 );
_HMUX g177dd ( \46509_nG177dd , RIe47c360_6304 , \46508_nG177dc , \44817 );
_HMUX g177df ( \46510_nG177df , RIe47c360_6304 , \45089 , \46306 );
_HMUX g177e0 ( \46511_nG177e0 , \46509_nG177dd , \46510_nG177df , \44829 );
buf \U$38083 ( \46512 , \46511_nG177e0 );
_DC g1912c_GF_IsGateDCbyConstraint ( \46513_nG1912c , \46512 , \42503 );
buf \U$38084 ( \46514 , \46513_nG1912c );
_HMUX g177e2 ( \46515_nG177e2 , RIe47cb58_6305 , \45095 , \46303 );
_HMUX g177e3 ( \46516_nG177e3 , RIe47cb58_6305 , \46515_nG177e2 , \44817 );
_HMUX g177e5 ( \46517_nG177e5 , RIe47cb58_6305 , \45098 , \46306 );
_HMUX g177e6 ( \46518_nG177e6 , \46516_nG177e3 , \46517_nG177e5 , \44829 );
buf \U$38085 ( \46519 , \46518_nG177e6 );
_DC g1912e_GF_IsGateDCbyConstraint ( \46520_nG1912e , \46519 , \42503 );
buf \U$38086 ( \46521 , \46520_nG1912e );
_HMUX g177e8 ( \46522_nG177e8 , RIe47d350_6306 , \45104 , \46303 );
_HMUX g177e9 ( \46523_nG177e9 , RIe47d350_6306 , \46522_nG177e8 , \44817 );
_HMUX g177eb ( \46524_nG177eb , RIe47d350_6306 , \45107 , \46306 );
_HMUX g177ec ( \46525_nG177ec , \46523_nG177e9 , \46524_nG177eb , \44829 );
buf \U$38087 ( \46526 , \46525_nG177ec );
_DC g19130_GF_IsGateDCbyConstraint ( \46527_nG19130 , \46526 , \42503 );
buf \U$38088 ( \46528 , \46527_nG19130 );
_HMUX g177ee ( \46529_nG177ee , RIe47db48_6307 , \45113 , \46303 );
_HMUX g177ef ( \46530_nG177ef , RIe47db48_6307 , \46529_nG177ee , \44817 );
_HMUX g177f1 ( \46531_nG177f1 , RIe47db48_6307 , \45116 , \46306 );
_HMUX g177f2 ( \46532_nG177f2 , \46530_nG177ef , \46531_nG177f1 , \44829 );
buf \U$38089 ( \46533 , \46532_nG177f2 );
_DC g19132_GF_IsGateDCbyConstraint ( \46534_nG19132 , \46533 , \42503 );
buf \U$38090 ( \46535 , \46534_nG19132 );
_HMUX g177f4 ( \46536_nG177f4 , RIe47e340_6308 , \45122 , \46303 );
_HMUX g177f5 ( \46537_nG177f5 , RIe47e340_6308 , \46536_nG177f4 , \44817 );
_HMUX g177f7 ( \46538_nG177f7 , RIe47e340_6308 , \45125 , \46306 );
_HMUX g177f8 ( \46539_nG177f8 , \46537_nG177f5 , \46538_nG177f7 , \44829 );
buf \U$38091 ( \46540 , \46539_nG177f8 );
_DC g19134_GF_IsGateDCbyConstraint ( \46541_nG19134 , \46540 , \42503 );
buf \U$38092 ( \46542 , \46541_nG19134 );
_HMUX g177fa ( \46543_nG177fa , RIe47eb38_6309 , \45131 , \46303 );
_HMUX g177fb ( \46544_nG177fb , RIe47eb38_6309 , \46543_nG177fa , \44817 );
_HMUX g177fd ( \46545_nG177fd , RIe47eb38_6309 , \45134 , \46306 );
_HMUX g177fe ( \46546_nG177fe , \46544_nG177fb , \46545_nG177fd , \44829 );
buf \U$38093 ( \46547 , \46546_nG177fe );
_DC g19136_GF_IsGateDCbyConstraint ( \46548_nG19136 , \46547 , \42503 );
buf \U$38094 ( \46549 , \46548_nG19136 );
_HMUX g17800 ( \46550_nG17800 , RIe47f330_6310 , \45140 , \46303 );
_HMUX g17801 ( \46551_nG17801 , RIe47f330_6310 , \46550_nG17800 , \44817 );
_HMUX g17803 ( \46552_nG17803 , RIe47f330_6310 , \45143 , \46306 );
_HMUX g17804 ( \46553_nG17804 , \46551_nG17801 , \46552_nG17803 , \44829 );
buf \U$38095 ( \46554 , \46553_nG17804 );
_DC g19138_GF_IsGateDCbyConstraint ( \46555_nG19138 , \46554 , \42503 );
buf \U$38096 ( \46556 , \46555_nG19138 );
_HMUX g17806 ( \46557_nG17806 , RIe47fb28_6311 , \45149 , \46303 );
_HMUX g17807 ( \46558_nG17807 , RIe47fb28_6311 , \46557_nG17806 , \44817 );
_HMUX g17809 ( \46559_nG17809 , RIe47fb28_6311 , \45152 , \46306 );
_HMUX g1780a ( \46560_nG1780a , \46558_nG17807 , \46559_nG17809 , \44829 );
buf \U$38097 ( \46561 , \46560_nG1780a );
_DC g1913a_GF_IsGateDCbyConstraint ( \46562_nG1913a , \46561 , \42503 );
buf \U$38098 ( \46563 , \46562_nG1913a );
_HMUX g1780c ( \46564_nG1780c , RIe480320_6312 , \45158 , \46303 );
_HMUX g1780d ( \46565_nG1780d , RIe480320_6312 , \46564_nG1780c , \44817 );
_HMUX g1780f ( \46566_nG1780f , RIe480320_6312 , \45161 , \46306 );
_HMUX g17810 ( \46567_nG17810 , \46565_nG1780d , \46566_nG1780f , \44829 );
buf \U$38099 ( \46568 , \46567_nG17810 );
_DC g1913c_GF_IsGateDCbyConstraint ( \46569_nG1913c , \46568 , \42503 );
buf \U$38100 ( \46570 , \46569_nG1913c );
_HMUX g17812 ( \46571_nG17812 , RIe480b18_6313 , \45167 , \46303 );
_HMUX g17813 ( \46572_nG17813 , RIe480b18_6313 , \46571_nG17812 , \44817 );
_HMUX g17815 ( \46573_nG17815 , RIe480b18_6313 , \45170 , \46306 );
_HMUX g17816 ( \46574_nG17816 , \46572_nG17813 , \46573_nG17815 , \44829 );
buf \U$38101 ( \46575 , \46574_nG17816 );
_DC g1913e_GF_IsGateDCbyConstraint ( \46576_nG1913e , \46575 , \42503 );
buf \U$38102 ( \46577 , \46576_nG1913e );
_HMUX g17818 ( \46578_nG17818 , RIe481310_6314 , \45176 , \46303 );
_HMUX g17819 ( \46579_nG17819 , RIe481310_6314 , \46578_nG17818 , \44817 );
_HMUX g1781b ( \46580_nG1781b , RIe481310_6314 , \45179 , \46306 );
_HMUX g1781c ( \46581_nG1781c , \46579_nG17819 , \46580_nG1781b , \44829 );
buf \U$38103 ( \46582 , \46581_nG1781c );
_DC g19142_GF_IsGateDCbyConstraint ( \46583_nG19142 , \46582 , \42503 );
buf \U$38104 ( \46584 , \46583_nG19142 );
_HMUX g1781e ( \46585_nG1781e , RIe481b08_6315 , \45185 , \46303 );
_HMUX g1781f ( \46586_nG1781f , RIe481b08_6315 , \46585_nG1781e , \44817 );
_HMUX g17821 ( \46587_nG17821 , RIe481b08_6315 , \45188 , \46306 );
_HMUX g17822 ( \46588_nG17822 , \46586_nG1781f , \46587_nG17821 , \44829 );
buf \U$38105 ( \46589 , \46588_nG17822 );
_DC g19144_GF_IsGateDCbyConstraint ( \46590_nG19144 , \46589 , \42503 );
buf \U$38106 ( \46591 , \46590_nG19144 );
_HMUX g17824 ( \46592_nG17824 , RIe482300_6316 , \45194 , \46303 );
_HMUX g17825 ( \46593_nG17825 , RIe482300_6316 , \46592_nG17824 , \44817 );
_HMUX g17827 ( \46594_nG17827 , RIe482300_6316 , \45197 , \46306 );
_HMUX g17828 ( \46595_nG17828 , \46593_nG17825 , \46594_nG17827 , \44829 );
buf \U$38107 ( \46596 , \46595_nG17828 );
_DC g19146_GF_IsGateDCbyConstraint ( \46597_nG19146 , \46596 , \42503 );
buf \U$38108 ( \46598 , \46597_nG19146 );
_HMUX g1782a ( \46599_nG1782a , RIe482af8_6317 , \45203 , \46303 );
_HMUX g1782b ( \46600_nG1782b , RIe482af8_6317 , \46599_nG1782a , \44817 );
_HMUX g1782d ( \46601_nG1782d , RIe482af8_6317 , \45206 , \46306 );
_HMUX g1782e ( \46602_nG1782e , \46600_nG1782b , \46601_nG1782d , \44829 );
buf \U$38109 ( \46603 , \46602_nG1782e );
_DC g19148_GF_IsGateDCbyConstraint ( \46604_nG19148 , \46603 , \42503 );
buf \U$38110 ( \46605 , \46604_nG19148 );
_HMUX g17830 ( \46606_nG17830 , RIe4832f0_6318 , \45212 , \46303 );
_HMUX g17831 ( \46607_nG17831 , RIe4832f0_6318 , \46606_nG17830 , \44817 );
_HMUX g17833 ( \46608_nG17833 , RIe4832f0_6318 , \45215 , \46306 );
_HMUX g17834 ( \46609_nG17834 , \46607_nG17831 , \46608_nG17833 , \44829 );
buf \U$38111 ( \46610 , \46609_nG17834 );
_DC g1914a_GF_IsGateDCbyConstraint ( \46611_nG1914a , \46610 , \42503 );
buf \U$38112 ( \46612 , \46611_nG1914a );
_HMUX g17836 ( \46613_nG17836 , RIe483ae8_6319 , \45221 , \46303 );
_HMUX g17837 ( \46614_nG17837 , RIe483ae8_6319 , \46613_nG17836 , \44817 );
_HMUX g17839 ( \46615_nG17839 , RIe483ae8_6319 , \45224 , \46306 );
_HMUX g1783a ( \46616_nG1783a , \46614_nG17837 , \46615_nG17839 , \44829 );
buf \U$38113 ( \46617 , \46616_nG1783a );
_DC g1914c_GF_IsGateDCbyConstraint ( \46618_nG1914c , \46617 , \42503 );
buf \U$38114 ( \46619 , \46618_nG1914c );
_HMUX g1783c ( \46620_nG1783c , RIe4842e0_6320 , \45230 , \46303 );
_HMUX g1783d ( \46621_nG1783d , RIe4842e0_6320 , \46620_nG1783c , \44817 );
_HMUX g1783f ( \46622_nG1783f , RIe4842e0_6320 , \45233 , \46306 );
_HMUX g17840 ( \46623_nG17840 , \46621_nG1783d , \46622_nG1783f , \44829 );
buf \U$38115 ( \46624 , \46623_nG17840 );
_DC g1914e_GF_IsGateDCbyConstraint ( \46625_nG1914e , \46624 , \42503 );
buf \U$38116 ( \46626 , \46625_nG1914e );
_HMUX g17842 ( \46627_nG17842 , RIe484ad8_6321 , \45239 , \46303 );
_HMUX g17843 ( \46628_nG17843 , RIe484ad8_6321 , \46627_nG17842 , \44817 );
_HMUX g17845 ( \46629_nG17845 , RIe484ad8_6321 , \45242 , \46306 );
_HMUX g17846 ( \46630_nG17846 , \46628_nG17843 , \46629_nG17845 , \44829 );
buf \U$38117 ( \46631 , \46630_nG17846 );
_DC g19150_GF_IsGateDCbyConstraint ( \46632_nG19150 , \46631 , \42503 );
buf \U$38118 ( \46633 , \46632_nG19150 );
_HMUX g17848 ( \46634_nG17848 , RIe4852d0_6322 , \45248 , \46303 );
_HMUX g17849 ( \46635_nG17849 , RIe4852d0_6322 , \46634_nG17848 , \44817 );
_HMUX g1784b ( \46636_nG1784b , RIe4852d0_6322 , \45251 , \46306 );
_HMUX g1784c ( \46637_nG1784c , \46635_nG17849 , \46636_nG1784b , \44829 );
buf \U$38119 ( \46638 , \46637_nG1784c );
_DC g19152_GF_IsGateDCbyConstraint ( \46639_nG19152 , \46638 , \42503 );
buf \U$38120 ( \46640 , \46639_nG19152 );
_HMUX g1784e ( \46641_nG1784e , RIe485ac8_6323 , \45257 , \46303 );
_HMUX g1784f ( \46642_nG1784f , RIe485ac8_6323 , \46641_nG1784e , \44817 );
_HMUX g17851 ( \46643_nG17851 , RIe485ac8_6323 , \45260 , \46306 );
_HMUX g17852 ( \46644_nG17852 , \46642_nG1784f , \46643_nG17851 , \44829 );
buf \U$38121 ( \46645 , \46644_nG17852 );
_DC g19154_GF_IsGateDCbyConstraint ( \46646_nG19154 , \46645 , \42503 );
buf \U$38122 ( \46647 , \46646_nG19154 );
_HMUX g17854 ( \46648_nG17854 , RIe4862c0_6324 , \45266 , \46303 );
_HMUX g17855 ( \46649_nG17855 , RIe4862c0_6324 , \46648_nG17854 , \44817 );
_HMUX g17857 ( \46650_nG17857 , RIe4862c0_6324 , \45269 , \46306 );
_HMUX g17858 ( \46651_nG17858 , \46649_nG17855 , \46650_nG17857 , \44829 );
buf \U$38123 ( \46652 , \46651_nG17858 );
_DC g19158_GF_IsGateDCbyConstraint ( \46653_nG19158 , \46652 , \42503 );
buf \U$38124 ( \46654 , \46653_nG19158 );
_HMUX g1785a ( \46655_nG1785a , RIe486ab8_6325 , \45275 , \46303 );
_HMUX g1785b ( \46656_nG1785b , RIe486ab8_6325 , \46655_nG1785a , \44817 );
_HMUX g1785d ( \46657_nG1785d , RIe486ab8_6325 , \45278 , \46306 );
_HMUX g1785e ( \46658_nG1785e , \46656_nG1785b , \46657_nG1785d , \44829 );
buf \U$38125 ( \46659 , \46658_nG1785e );
_DC g1915a_GF_IsGateDCbyConstraint ( \46660_nG1915a , \46659 , \42503 );
buf \U$38126 ( \46661 , \46660_nG1915a );
_HMUX g17860 ( \46662_nG17860 , RIe4872b0_6326 , \45284 , \46303 );
_HMUX g17861 ( \46663_nG17861 , RIe4872b0_6326 , \46662_nG17860 , \44817 );
_HMUX g17863 ( \46664_nG17863 , RIe4872b0_6326 , \45287 , \46306 );
_HMUX g17864 ( \46665_nG17864 , \46663_nG17861 , \46664_nG17863 , \44829 );
buf \U$38127 ( \46666 , \46665_nG17864 );
_DC g1915c_GF_IsGateDCbyConstraint ( \46667_nG1915c , \46666 , \42503 );
buf \U$38128 ( \46668 , \46667_nG1915c );
_HMUX g17866 ( \46669_nG17866 , RIe487aa8_6327 , \45293 , \46303 );
_HMUX g17867 ( \46670_nG17867 , RIe487aa8_6327 , \46669_nG17866 , \44817 );
_HMUX g17869 ( \46671_nG17869 , RIe487aa8_6327 , \45296 , \46306 );
_HMUX g1786a ( \46672_nG1786a , \46670_nG17867 , \46671_nG17869 , \44829 );
buf \U$38129 ( \46673 , \46672_nG1786a );
_DC g1915e_GF_IsGateDCbyConstraint ( \46674_nG1915e , \46673 , \42503 );
buf \U$38130 ( \46675 , \46674_nG1915e );
_HMUX g1786c ( \46676_nG1786c , RIe4882a0_6328 , \45302 , \46303 );
_HMUX g1786d ( \46677_nG1786d , RIe4882a0_6328 , \46676_nG1786c , \44817 );
_HMUX g1786f ( \46678_nG1786f , RIe4882a0_6328 , \45305 , \46306 );
_HMUX g17870 ( \46679_nG17870 , \46677_nG1786d , \46678_nG1786f , \44829 );
buf \U$38131 ( \46680 , \46679_nG17870 );
_DC g19160_GF_IsGateDCbyConstraint ( \46681_nG19160 , \46680 , \42503 );
buf \U$38132 ( \46682 , \46681_nG19160 );
_HMUX g17872 ( \46683_nG17872 , RIe488a98_6329 , \45311 , \46303 );
_HMUX g17873 ( \46684_nG17873 , RIe488a98_6329 , \46683_nG17872 , \44817 );
_HMUX g17875 ( \46685_nG17875 , RIe488a98_6329 , \45314 , \46306 );
_HMUX g17876 ( \46686_nG17876 , \46684_nG17873 , \46685_nG17875 , \44829 );
buf \U$38133 ( \46687 , \46686_nG17876 );
_DC g19162_GF_IsGateDCbyConstraint ( \46688_nG19162 , \46687 , \42503 );
buf \U$38134 ( \46689 , \46688_nG19162 );
_HMUX g17878 ( \46690_nG17878 , RIe489290_6330 , \45320 , \46303 );
_HMUX g17879 ( \46691_nG17879 , RIe489290_6330 , \46690_nG17878 , \44817 );
_HMUX g1787b ( \46692_nG1787b , RIe489290_6330 , \45323 , \46306 );
_HMUX g1787c ( \46693_nG1787c , \46691_nG17879 , \46692_nG1787b , \44829 );
buf \U$38135 ( \46694 , \46693_nG1787c );
_DC g19164_GF_IsGateDCbyConstraint ( \46695_nG19164 , \46694 , \42503 );
buf \U$38136 ( \46696 , \46695_nG19164 );
_HMUX g1787e ( \46697_nG1787e , RIe489a88_6331 , \45329 , \46303 );
_HMUX g1787f ( \46698_nG1787f , RIe489a88_6331 , \46697_nG1787e , \44817 );
_HMUX g17881 ( \46699_nG17881 , RIe489a88_6331 , \45332 , \46306 );
_HMUX g17882 ( \46700_nG17882 , \46698_nG1787f , \46699_nG17881 , \44829 );
buf \U$38137 ( \46701 , \46700_nG17882 );
_DC g19166_GF_IsGateDCbyConstraint ( \46702_nG19166 , \46701 , \42503 );
buf \U$38138 ( \46703 , \46702_nG19166 );
_HMUX g17884 ( \46704_nG17884 , RIe48a280_6332 , \45338 , \46303 );
_HMUX g17885 ( \46705_nG17885 , RIe48a280_6332 , \46704_nG17884 , \44817 );
_HMUX g17887 ( \46706_nG17887 , RIe48a280_6332 , \45341 , \46306 );
_HMUX g17888 ( \46707_nG17888 , \46705_nG17885 , \46706_nG17887 , \44829 );
buf \U$38139 ( \46708 , \46707_nG17888 );
_DC g19168_GF_IsGateDCbyConstraint ( \46709_nG19168 , \46708 , \42503 );
buf \U$38140 ( \46710 , \46709_nG19168 );
_HMUX g1788a ( \46711_nG1788a , RIe48aa78_6333 , \45347 , \46303 );
_HMUX g1788b ( \46712_nG1788b , RIe48aa78_6333 , \46711_nG1788a , \44817 );
_HMUX g1788d ( \46713_nG1788d , RIe48aa78_6333 , \45350 , \46306 );
_HMUX g1788e ( \46714_nG1788e , \46712_nG1788b , \46713_nG1788d , \44829 );
buf \U$38141 ( \46715 , \46714_nG1788e );
_DC g1916a_GF_IsGateDCbyConstraint ( \46716_nG1916a , \46715 , \42503 );
buf \U$38142 ( \46717 , \46716_nG1916a );
_HMUX g17890 ( \46718_nG17890 , RIe48b270_6334 , \45356 , \46303 );
_HMUX g17891 ( \46719_nG17891 , RIe48b270_6334 , \46718_nG17890 , \44817 );
_HMUX g17893 ( \46720_nG17893 , RIe48b270_6334 , \45359 , \46306 );
_HMUX g17894 ( \46721_nG17894 , \46719_nG17891 , \46720_nG17893 , \44829 );
buf \U$38143 ( \46722 , \46721_nG17894 );
_DC g1916e_GF_IsGateDCbyConstraint ( \46723_nG1916e , \46722 , \42503 );
buf \U$38144 ( \46724 , \46723_nG1916e );
_HMUX g17896 ( \46725_nG17896 , RIe48ba68_6335 , \45365 , \46303 );
_HMUX g17897 ( \46726_nG17897 , RIe48ba68_6335 , \46725_nG17896 , \44817 );
_HMUX g17899 ( \46727_nG17899 , RIe48ba68_6335 , \45368 , \46306 );
_HMUX g1789a ( \46728_nG1789a , \46726_nG17897 , \46727_nG17899 , \44829 );
buf \U$38145 ( \46729 , \46728_nG1789a );
_DC g19170_GF_IsGateDCbyConstraint ( \46730_nG19170 , \46729 , \42503 );
buf \U$38146 ( \46731 , \46730_nG19170 );
_HMUX g1789c ( \46732_nG1789c , RIe48c260_6336 , \45374 , \46303 );
_HMUX g1789d ( \46733_nG1789d , RIe48c260_6336 , \46732_nG1789c , \44817 );
_HMUX g1789f ( \46734_nG1789f , RIe48c260_6336 , \45377 , \46306 );
_HMUX g178a0 ( \46735_nG178a0 , \46733_nG1789d , \46734_nG1789f , \44829 );
buf \U$38147 ( \46736 , \46735_nG178a0 );
_DC g19172_GF_IsGateDCbyConstraint ( \46737_nG19172 , \46736 , \42503 );
buf \U$38148 ( \46738 , \46737_nG19172 );
_HMUX g178a2 ( \46739_nG178a2 , RIe48ca58_6337 , \45383 , \46303 );
_HMUX g178a3 ( \46740_nG178a3 , RIe48ca58_6337 , \46739_nG178a2 , \44817 );
_HMUX g178a5 ( \46741_nG178a5 , RIe48ca58_6337 , \45386 , \46306 );
_HMUX g178a6 ( \46742_nG178a6 , \46740_nG178a3 , \46741_nG178a5 , \44829 );
buf \U$38149 ( \46743 , \46742_nG178a6 );
_DC g19174_GF_IsGateDCbyConstraint ( \46744_nG19174 , \46743 , \42503 );
buf \U$38150 ( \46745 , \46744_nG19174 );
_HMUX g178a8 ( \46746_nG178a8 , RIe48d250_6338 , \45392 , \46303 );
_HMUX g178a9 ( \46747_nG178a9 , RIe48d250_6338 , \46746_nG178a8 , \44817 );
_HMUX g178ab ( \46748_nG178ab , RIe48d250_6338 , \45395 , \46306 );
_HMUX g178ac ( \46749_nG178ac , \46747_nG178a9 , \46748_nG178ab , \44829 );
buf \U$38151 ( \46750 , \46749_nG178ac );
_DC g19176_GF_IsGateDCbyConstraint ( \46751_nG19176 , \46750 , \42503 );
buf \U$38152 ( \46752 , \46751_nG19176 );
buf \U$38153 ( \46753 , RIb86fc68_77);
_HMUX g176fd ( \46754_nG176fd , RIe3cd190_6051 , \46753 , \44810 );
not \U$38154 ( \46755 , \44817 );
or \U$38155 ( \46756 , \44829 , \46755 );
_HMUX g176fe ( \46757_nG176fe , \46754_nG176fd , RIe3cd190_6051 , \46756 );
buf \U$38156 ( \46758 , \46757_nG176fe );
_DC g190e6_GF_IsGateDCbyConstraint ( \46759_nG190e6 , \46758 , \42503 );
buf \U$38157 ( \46760 , \46759_nG190e6 );
buf \U$38158 ( \46761 , RIb86fce0_76);
_HMUX g176ff ( \46762_nG176ff , RIe3cc3f8_6052 , \46761 , \44810 );
_HMUX g17700 ( \46763_nG17700 , \46762_nG176ff , RIe3cc3f8_6052 , \46756 );
buf \U$38159 ( \46764 , \46763_nG17700 );
_DC g190e8_GF_IsGateDCbyConstraint ( \46765_nG190e8 , \46764 , \42503 );
buf \U$38160 ( \46766 , \46765_nG190e8 );
buf \U$38161 ( \46767 , RIb86fd58_75);
_HMUX g17701 ( \46768_nG17701 , RIe3cb750_6053 , \46767 , \44810 );
_HMUX g17702 ( \46769_nG17702 , \46768_nG17701 , RIe3cb750_6053 , \46756 );
buf \U$38162 ( \46770 , \46769_nG17702 );
_DC g190ea_GF_IsGateDCbyConstraint ( \46771_nG190ea , \46770 , \42503 );
buf \U$38163 ( \46772 , \46771_nG190ea );
buf \U$38164 ( \46773 , RIb87e8a8_74);
_HMUX g17703 ( \46774_nG17703 , RIe3ca9b8_6054 , \46773 , \44810 );
_HMUX g17704 ( \46775_nG17704 , \46774_nG17703 , RIe3ca9b8_6054 , \46756 );
buf \U$38165 ( \46776 , \46775_nG17704 );
_DC g190ec_GF_IsGateDCbyConstraint ( \46777_nG190ec , \46776 , \42503 );
buf \U$38166 ( \46778 , \46777_nG190ec );
buf \U$38167 ( \46779 , RIb87e920_73);
_HMUX g17705 ( \46780_nG17705 , RIe3c9e00_6055 , \46779 , \44810 );
_HMUX g17706 ( \46781_nG17706 , \46780_nG17705 , RIe3c9e00_6055 , \46756 );
buf \U$38168 ( \46782 , \46781_nG17706 );
_DC g190ee_GF_IsGateDCbyConstraint ( \46783_nG190ee , \46782 , \42503 );
buf \U$38169 ( \46784 , \46783_nG190ee );
buf \U$38170 ( \46785 , RIb87e998_72);
_HMUX g17707 ( \46786_nG17707 , RIe3c9248_6056 , \46785 , \44810 );
_HMUX g17708 ( \46787_nG17708 , \46786_nG17707 , RIe3c9248_6056 , \46756 );
buf \U$38171 ( \46788 , \46787_nG17708 );
_DC g190f0_GF_IsGateDCbyConstraint ( \46789_nG190f0 , \46788 , \42503 );
buf \U$38172 ( \46790 , \46789_nG190f0 );
buf \U$38173 ( \46791 , RIb87ea10_71);
_HMUX g17709 ( \46792_nG17709 , RIe3c8708_6057 , \46791 , \44810 );
_HMUX g1770a ( \46793_nG1770a , \46792_nG17709 , RIe3c8708_6057 , \46756 );
buf \U$38174 ( \46794 , \46793_nG1770a );
_DC g190f2_GF_IsGateDCbyConstraint ( \46795_nG190f2 , \46794 , \42503 );
buf \U$38175 ( \46796 , \46795_nG190f2 );
buf \U$38176 ( \46797 , RIb87ea88_70);
_HMUX g1770b ( \46798_nG1770b , RIe3c7bc8_6058 , \46797 , \44810 );
_HMUX g1770c ( \46799_nG1770c , \46798_nG1770b , RIe3c7bc8_6058 , \46756 );
buf \U$38177 ( \46800 , \46799_nG1770c );
_DC g190f4_GF_IsGateDCbyConstraint ( \46801_nG190f4 , \46800 , \42503 );
buf \U$38178 ( \46802 , \46801_nG190f4 );
_HMUX g176ec ( \46803_nG176ec , RIe3c7100_6059 , \46753 , \45402 );
_HMUX g176ed ( \46804_nG176ed , \46803_nG176ec , RIe3c7100_6059 , \46756 );
buf \U$38179 ( \46805 , \46804_nG176ed );
_DC g190d6_GF_IsGateDCbyConstraint ( \46806_nG190d6 , \46805 , \42503 );
buf \U$38180 ( \46807 , \46806_nG190d6 );
_HMUX g176ee ( \46808_nG176ee , RIe3c6638_6060 , \46761 , \45402 );
_HMUX g176ef ( \46809_nG176ef , \46808_nG176ee , RIe3c6638_6060 , \46756 );
buf \U$38181 ( \46810 , \46809_nG176ef );
_DC g190d8_GF_IsGateDCbyConstraint ( \46811_nG190d8 , \46810 , \42503 );
buf \U$38182 ( \46812 , \46811_nG190d8 );
_HMUX g176f0 ( \46813_nG176f0 , RIe3c5af8_6061 , \46767 , \45402 );
_HMUX g176f1 ( \46814_nG176f1 , \46813_nG176f0 , RIe3c5af8_6061 , \46756 );
buf \U$38183 ( \46815 , \46814_nG176f1 );
_DC g190da_GF_IsGateDCbyConstraint ( \46816_nG190da , \46815 , \42503 );
buf \U$38184 ( \46817 , \46816_nG190da );
_HMUX g176f2 ( \46818_nG176f2 , RIe3c4ec8_6062 , \46773 , \45402 );
_HMUX g176f3 ( \46819_nG176f3 , \46818_nG176f2 , RIe3c4ec8_6062 , \46756 );
buf \U$38185 ( \46820 , \46819_nG176f3 );
_DC g190dc_GF_IsGateDCbyConstraint ( \46821_nG190dc , \46820 , \42503 );
buf \U$38186 ( \46822 , \46821_nG190dc );
_HMUX g176f4 ( \46823_nG176f4 , RIe3c4130_6063 , \46779 , \45402 );
_HMUX g176f5 ( \46824_nG176f5 , \46823_nG176f4 , RIe3c4130_6063 , \46756 );
buf \U$38187 ( \46825 , \46824_nG176f5 );
_DC g190de_GF_IsGateDCbyConstraint ( \46826_nG190de , \46825 , \42503 );
buf \U$38188 ( \46827 , \46826_nG190de );
_HMUX g176f6 ( \46828_nG176f6 , RIe3c31b8_6064 , \46785 , \45402 );
_HMUX g176f7 ( \46829_nG176f7 , \46828_nG176f6 , RIe3c31b8_6064 , \46756 );
buf \U$38189 ( \46830 , \46829_nG176f7 );
_DC g190e0_GF_IsGateDCbyConstraint ( \46831_nG190e0 , \46830 , \42503 );
buf \U$38190 ( \46832 , \46831_nG190e0 );
_HMUX g176f8 ( \46833_nG176f8 , RIe3c1bb0_6065 , \46791 , \45402 );
_HMUX g176f9 ( \46834_nG176f9 , \46833_nG176f8 , RIe3c1bb0_6065 , \46756 );
buf \U$38191 ( \46835 , \46834_nG176f9 );
_DC g190e2_GF_IsGateDCbyConstraint ( \46836_nG190e2 , \46835 , \42503 );
buf \U$38192 ( \46837 , \46836_nG190e2 );
_HMUX g176fa ( \46838_nG176fa , RIe3c0a58_6066 , \46797 , \45402 );
_HMUX g176fb ( \46839_nG176fb , \46838_nG176fa , RIe3c0a58_6066 , \46756 );
buf \U$38193 ( \46840 , \46839_nG176fb );
_DC g190e4_GF_IsGateDCbyConstraint ( \46841_nG190e4 , \46840 , \42503 );
buf \U$38194 ( \46842 , \46841_nG190e4 );
_HMUX g176db ( \46843_nG176db , RIe3bf900_6067 , \46753 , \45853 );
_HMUX g176dc ( \46844_nG176dc , \46843_nG176db , RIe3bf900_6067 , \46756 );
buf \U$38195 ( \46845 , \46844_nG176dc );
_DC g190c6_GF_IsGateDCbyConstraint ( \46846_nG190c6 , \46845 , \42503 );
buf \U$38196 ( \46847 , \46846_nG190c6 );
_HMUX g176dd ( \46848_nG176dd , RIe3be2f8_6068 , \46761 , \45853 );
_HMUX g176de ( \46849_nG176de , \46848_nG176dd , RIe3be2f8_6068 , \46756 );
buf \U$38197 ( \46850 , \46849_nG176de );
_DC g190c8_GF_IsGateDCbyConstraint ( \46851_nG190c8 , \46850 , \42503 );
buf \U$38198 ( \46852 , \46851_nG190c8 );
_HMUX g176df ( \46853_nG176df , RIe3bd1a0_6069 , \46767 , \45853 );
_HMUX g176e0 ( \46854_nG176e0 , \46853_nG176df , RIe3bd1a0_6069 , \46756 );
buf \U$38199 ( \46855 , \46854_nG176e0 );
_DC g190ca_GF_IsGateDCbyConstraint ( \46856_nG190ca , \46855 , \42503 );
buf \U$38200 ( \46857 , \46856_nG190ca );
_HMUX g176e1 ( \46858_nG176e1 , RIe3bbb98_6070 , \46773 , \45853 );
_HMUX g176e2 ( \46859_nG176e2 , \46858_nG176e1 , RIe3bbb98_6070 , \46756 );
buf \U$38201 ( \46860 , \46859_nG176e2 );
_DC g190cc_GF_IsGateDCbyConstraint ( \46861_nG190cc , \46860 , \42503 );
buf \U$38202 ( \46862 , \46861_nG190cc );
_HMUX g176e3 ( \46863_nG176e3 , RIe3baa40_6071 , \46779 , \45853 );
_HMUX g176e4 ( \46864_nG176e4 , \46863_nG176e3 , RIe3baa40_6071 , \46756 );
buf \U$38203 ( \46865 , \46864_nG176e4 );
_DC g190ce_GF_IsGateDCbyConstraint ( \46866_nG190ce , \46865 , \42503 );
buf \U$38204 ( \46867 , \46866_nG190ce );
_HMUX g176e5 ( \46868_nG176e5 , RIe3b9438_6072 , \46785 , \45853 );
_HMUX g176e6 ( \46869_nG176e6 , \46868_nG176e5 , RIe3b9438_6072 , \46756 );
buf \U$38205 ( \46870 , \46869_nG176e6 );
_DC g190d0_GF_IsGateDCbyConstraint ( \46871_nG190d0 , \46870 , \42503 );
buf \U$38206 ( \46872 , \46871_nG190d0 );
_HMUX g176e7 ( \46873_nG176e7 , RIe3b82e0_6073 , \46791 , \45853 );
_HMUX g176e8 ( \46874_nG176e8 , \46873_nG176e7 , RIe3b82e0_6073 , \46756 );
buf \U$38207 ( \46875 , \46874_nG176e8 );
_DC g190d2_GF_IsGateDCbyConstraint ( \46876_nG190d2 , \46875 , \42503 );
buf \U$38208 ( \46877 , \46876_nG190d2 );
_HMUX g176e9 ( \46878_nG176e9 , RIe3b7188_6074 , \46797 , \45853 );
_HMUX g176ea ( \46879_nG176ea , \46878_nG176e9 , RIe3b7188_6074 , \46756 );
buf \U$38209 ( \46880 , \46879_nG176ea );
_DC g190d4_GF_IsGateDCbyConstraint ( \46881_nG190d4 , \46880 , \42503 );
buf \U$38210 ( \46882 , \46881_nG190d4 );
_HMUX g176ba ( \46883_nG176ba , RIe3b5b80_6075 , \46753 , \46303 );
_HMUX g176c3 ( \46884_nG176c3 , \46883_nG176ba , RIe3b5b80_6075 , \46756 );
buf \U$38211 ( \46885 , \46884_nG176c3 );
_DC g192fe_GF_IsGateDCbyConstraint ( \46886_nG192fe , \46885 , \42503 );
buf \U$38212 ( \46887 , \46886_nG192fe );
_HMUX g176c5 ( \46888_nG176c5 , RIe3b4a28_6076 , \46761 , \46303 );
_HMUX g176c6 ( \46889_nG176c6 , \46888_nG176c5 , RIe3b4a28_6076 , \46756 );
buf \U$38213 ( \46890 , \46889_nG176c6 );
_DC g19300_GF_IsGateDCbyConstraint ( \46891_nG19300 , \46890 , \42503 );
buf \U$38214 ( \46892 , \46891_nG19300 );
_HMUX g176c8 ( \46893_nG176c8 , RIe3b3420_6077 , \46767 , \46303 );
_HMUX g176c9 ( \46894_nG176c9 , \46893_nG176c8 , RIe3b3420_6077 , \46756 );
buf \U$38215 ( \46895 , \46894_nG176c9 );
_DC g19302_GF_IsGateDCbyConstraint ( \46896_nG19302 , \46895 , \42503 );
buf \U$38216 ( \46897 , \46896_nG19302 );
_HMUX g176cb ( \46898_nG176cb , RIe3b22c8_6078 , \46773 , \46303 );
_HMUX g176cc ( \46899_nG176cc , \46898_nG176cb , RIe3b22c8_6078 , \46756 );
buf \U$38217 ( \46900 , \46899_nG176cc );
_DC g19304_GF_IsGateDCbyConstraint ( \46901_nG19304 , \46900 , \42503 );
buf \U$38218 ( \46902 , \46901_nG19304 );
_HMUX g176ce ( \46903_nG176ce , RIe3b0cc0_6079 , \46779 , \46303 );
_HMUX g176cf ( \46904_nG176cf , \46903_nG176ce , RIe3b0cc0_6079 , \46756 );
buf \U$38219 ( \46905 , \46904_nG176cf );
_DC g19306_GF_IsGateDCbyConstraint ( \46906_nG19306 , \46905 , \42503 );
buf \U$38220 ( \46907 , \46906_nG19306 );
_HMUX g176d1 ( \46908_nG176d1 , RIe3afb68_6080 , \46785 , \46303 );
_HMUX g176d2 ( \46909_nG176d2 , \46908_nG176d1 , RIe3afb68_6080 , \46756 );
buf \U$38221 ( \46910 , \46909_nG176d2 );
_DC g19308_GF_IsGateDCbyConstraint ( \46911_nG19308 , \46910 , \42503 );
buf \U$38222 ( \46912 , \46911_nG19308 );
_HMUX g176d4 ( \46913_nG176d4 , RIe3aea10_6081 , \46791 , \46303 );
_HMUX g176d5 ( \46914_nG176d5 , \46913_nG176d4 , RIe3aea10_6081 , \46756 );
buf \U$38223 ( \46915 , \46914_nG176d5 );
_DC g1930a_GF_IsGateDCbyConstraint ( \46916_nG1930a , \46915 , \42503 );
buf \U$38224 ( \46917 , \46916_nG1930a );
_HMUX g176d7 ( \46918_nG176d7 , RIe3ad408_6082 , \46797 , \46303 );
_HMUX g176d8 ( \46919_nG176d8 , \46918_nG176d7 , RIe3ad408_6082 , \46756 );
buf \U$38225 ( \46920 , \46919_nG176d8 );
_DC g1930c_GF_IsGateDCbyConstraint ( \46921_nG1930c , \46920 , \42503 );
buf \U$38226 ( \46922 , \46921_nG1930c );
buf \U$38227 ( \46923 , RIb7b9680_245);
buf \U$38228 ( \46924 , RIb79b3b0_273);
and \U$38229 ( \46925 , \44825 , \46924 );
_HMUX g175af ( \46926_nG175af , RIe51b690_6365 , \46923 , \46925 );
buf \U$38230 ( \46927 , \46926_nG175af );
_DC g1930d_GF_IsGateDCbyConstraint ( \46928_nG1930d , \46927 , \42503 );
buf \U$38231 ( \46929 , \46928_nG1930d );
buf \U$38232 ( \46930 , RIb7b96f8_244);
_HMUX g1761c ( \46931_nG1761c , RIe500d68_6388 , \46930 , \46925 );
buf \U$38233 ( \46932 , \46931_nG1761c );
_DC g190aa_GF_IsGateDCbyConstraint ( \46933_nG190aa , \46932 , \42503 );
buf \U$38234 ( \46934 , \46933_nG190aa );
buf \U$38235 ( \46935 , RIb7c20c8_243);
_HMUX g1761e ( \46936_nG1761e , RIe501998_6387 , \46935 , \46925 );
buf \U$38236 ( \46937 , \46936_nG1761e );
_DC g190ac_GF_IsGateDCbyConstraint ( \46938_nG190ac , \46937 , \42503 );
buf \U$38237 ( \46939 , \46938_nG190ac );
buf \U$38238 ( \46940 , RIb7c5728_242);
_HMUX g17620 ( \46941_nG17620 , RIe5026b8_6386 , \46940 , \46925 );
buf \U$38239 ( \46942 , \46941_nG17620 );
_DC g190ae_GF_IsGateDCbyConstraint ( \46943_nG190ae , \46942 , \42503 );
buf \U$38240 ( \46944 , \46943_nG190ae );
buf \U$38241 ( \46945 , RIb7c57a0_241);
_HMUX g17622 ( \46946_nG17622 , RIe5032e8_6385 , \46945 , \46925 );
buf \U$38242 ( \46947 , \46946_nG17622 );
_DC g190b0_GF_IsGateDCbyConstraint ( \46948_nG190b0 , \46947 , \42503 );
buf \U$38243 ( \46949 , \46948_nG190b0 );
buf \U$38244 ( \46950 , RIb7c5818_240);
_HMUX g17624 ( \46951_nG17624 , RIe503f90_6384 , \46950 , \46925 );
buf \U$38245 ( \46952 , \46951_nG17624 );
_DC g190b2_GF_IsGateDCbyConstraint ( \46953_nG190b2 , \46952 , \42503 );
buf \U$38246 ( \46954 , \46953_nG190b2 );
buf \U$38247 ( \46955 , RIb7c5890_239);
_HMUX g17626 ( \46956_nG17626 , RIe504d28_6383 , \46955 , \46925 );
buf \U$38248 ( \46957 , \46956_nG17626 );
_DC g190b4_GF_IsGateDCbyConstraint ( \46958_nG190b4 , \46957 , \42503 );
buf \U$38249 ( \46959 , \46958_nG190b4 );
buf \U$38250 ( \46960 , RIb7c5908_238);
_HMUX g17628 ( \46961_nG17628 , RIe505958_6382 , \46960 , \46925 );
buf \U$38251 ( \46962 , \46961_nG17628 );
_DC g190b6_GF_IsGateDCbyConstraint ( \46963_nG190b6 , \46962 , \42503 );
buf \U$38252 ( \46964 , \46963_nG190b6 );
buf \U$38253 ( \46965 , RIb7a09f0_266);
_HMUX g1761a ( \46966_nG1761a , RIe50ef58_6371 , \46965 , \46925 );
buf \U$38254 ( \46967 , \46966_nG1761a );
_DC g190a8_GF_IsGateDCbyConstraint ( \46968_nG190a8 , \46967 , \42503 );
buf \U$38255 ( \46969 , \46968_nG190a8 );
buf \U$38256 ( \46970 , RIb7a0a68_265);
_HMUX g17612 ( \46971_nG17612 , RIe50ac50_6376 , \46970 , \46925 );
buf \U$38257 ( \46972 , \46971_nG17612 );
_DC g190a0_GF_IsGateDCbyConstraint ( \46973_nG190a0 , \46972 , \42503 );
buf \U$38258 ( \46974 , \46973_nG190a0 );
buf \U$38259 ( \46975 , RIb7a0ae0_264);
_HMUX g17614 ( \46976_nG17614 , RIe50b880_6375 , \46975 , \46925 );
buf \U$38260 ( \46977 , \46976_nG17614 );
_DC g190a2_GF_IsGateDCbyConstraint ( \46978_nG190a2 , \46977 , \42503 );
buf \U$38261 ( \46979 , \46978_nG190a2 );
buf \U$38262 ( \46980 , RIb7a0b58_263);
_HMUX g17616 ( \46981_nG17616 , RIe50c690_6374 , \46980 , \46925 );
buf \U$38263 ( \46982 , \46981_nG17616 );
_DC g190a4_GF_IsGateDCbyConstraint ( \46983_nG190a4 , \46982 , \42503 );
buf \U$38264 ( \46984 , \46983_nG190a4 );
buf \U$38265 ( \46985 , RIb7a0bd0_262);
_HMUX g17618 ( \46986_nG17618 , RIe50d428_6373 , \46985 , \46925 );
buf \U$38266 ( \46987 , \46986_nG17618 );
_DC g190a6_GF_IsGateDCbyConstraint ( \46988_nG190a6 , \46987 , \42503 );
buf \U$38267 ( \46989 , \46988_nG190a6 );
buf \U$38268 ( \46990 , RIe523688_6352);
not \U$38269 ( \46991 , \46990 );
buf \U$38270 ( \46992 , \46991 );
nor \U$38272 ( \46993 , RIe523688_6352, RIe524060_6351, RIe524948_6350);
_HMUX g17482 ( \46994_nG17482 , \46992 , 1'b0 , \46993 );
and \U$38273 ( \46995 , RIe5319e0_6884, RIe549ef0_6842, RIe549770_6843, RIe548ff0_6844, \7063 );
buf \U$38274 ( \46996 , \46995 );
buf \U$38275 ( \46997 , RIb79b4a0_271);
and \U$38276 ( \46998 , \46996 , \46997 );
_HMUX g17483 ( \46999_nG17483 , RIe523688_6352 , \46994_nG17482 , \46998 );
buf \U$38277 ( \47000 , RIe523688_6352);
not \U$38278 ( \47001 , \47000 );
buf \U$38279 ( \47002 , \47001 );
not \U$38280 ( \47003 , RIe524948_6350);
nor \U$38281 ( \47004 , RIe523688_6352, RIe524060_6351, \47003 );
_HMUX g17489 ( \47005_nG17489 , \47002 , RIe523688_6352 , \47004 );
and \U$38282 ( \47006 , \44827 , \44825 );
_HMUX g1748d ( \47007_nG1748d , \46999_nG17483 , \47005_nG17489 , \47006 );
and \U$38283 ( \47008 , \47006 , \46997 );
and \U$38284 ( \47009 , \47008 , \46996 );
_HMUX g17490 ( \47010_nG17490 , \47007_nG1748d , RIe523688_6352 , \47009 );
not \U$38285 ( \47011 , RIe5117a8_6369);
and \U$38286 ( \47012 , RIe5117a8_6369, \46923 );
or \U$38287 ( \47013 , \47011 , \47012 );
and \U$38288 ( \47014 , \47013 , \44827 );
and \U$38289 ( \47015 , \47014 , \44825 );
_HMUX g17497 ( \47016_nG17497 , \47010_nG17490 , RIe51c158_6364 , \47015 );
buf \U$38291 ( \47017 , RIb79b338_274);
and \U$38292 ( \47018 , \46996 , \47017 );
_HMUX g17498 ( \47019_nG17498 , \47016_nG17497 , 1'b0 , \47018 );
buf \U$38293 ( \47020 , \47019_nG17498 );
buf \U$38294 ( \47021 , RIe524060_6351);
xnor \U$38295 ( \47022 , \47021 , \46990 );
buf \U$38296 ( \47023 , \47022 );
_HMUX g1749c ( \47024_nG1749c , \47023 , 1'b0 , \46993 );
_HMUX g1749d ( \47025_nG1749d , RIe524060_6351 , \47024_nG1749c , \46998 );
buf \U$38298 ( \47026 , RIe524060_6351);
xor \U$38299 ( \47027 , \47026 , \47000 );
buf \U$38300 ( \47028 , \47027 );
_HMUX g174a1 ( \47029_nG174a1 , \47028 , RIe524060_6351 , \47004 );
_HMUX g174a2 ( \47030_nG174a2 , \47025_nG1749d , \47029_nG174a1 , \47006 );
_HMUX g174a3 ( \47031_nG174a3 , \47030_nG174a2 , RIe524060_6351 , \47009 );
_HMUX g174a4 ( \47032_nG174a4 , \47031_nG174a3 , RIe51cc20_6363 , \47015 );
_HMUX g174a5 ( \47033_nG174a5 , \47032_nG174a4 , 1'b0 , \47018 );
buf \U$38302 ( \47034 , \47033_nG174a5 );
buf \U$38303 ( \47035 , RIe524948_6350);
or \U$38304 ( \47036 , \47021 , \46990 );
xnor \U$38305 ( \47037 , \47035 , \47036 );
buf \U$38306 ( \47038 , \47037 );
_HMUX g174aa ( \47039_nG174aa , \47038 , 1'b0 , \46993 );
_HMUX g174ab ( \47040_nG174ab , RIe524948_6350 , \47039_nG174aa , \46998 );
buf \U$38308 ( \47041 , RIe524948_6350);
and \U$38309 ( \47042 , \47026 , \47000 );
xor \U$38310 ( \47043 , \47041 , \47042 );
buf \U$38311 ( \47044 , \47043 );
_HMUX g174b0 ( \47045_nG174b0 , \47044 , RIe524948_6350 , \47004 );
_HMUX g174b1 ( \47046_nG174b1 , \47040_nG174ab , \47045_nG174b0 , \47006 );
_HMUX g174b2 ( \47047_nG174b2 , \47046_nG174b1 , RIe524948_6350 , \47009 );
_HMUX g174b3 ( \47048_nG174b3 , \47047_nG174b2 , RIe51d5f8_6362 , \47015 );
_HMUX g174b4 ( \47049_nG174b4 , \47048_nG174b3 , 1'b0 , \47018 );
buf \U$38313 ( \47050 , \47049_nG174b4 );
or \U$38314 ( \47051 , \47020 , \47034 , \47050 );
buf \U$38315 ( \47052 , \47051 );
buf \U$38316 ( \47053 , RIe5267c0_6347);
buf \U$38317 ( \47054 , RIe525d70_6348);
buf \U$38318 ( \47055 , RIe525410_6349);
and \U$38319 ( \47056 , \47054 , \47055 );
xor \U$38320 ( \47057 , \47053 , \47056 );
buf \U$38321 ( \47058 , \47057 );
not \U$38322 ( \47059 , RIe5267c0_6347);
nor \U$38323 ( \47060 , RIe525410_6349, RIe525d70_6348, \47059 );
not \U$38324 ( \47061 , \47060 );
and \U$38325 ( \47062 , \46998 , \47061 );
_HMUX g17479 ( \47063_nG17479 , RIe5267c0_6347 , \47058 , \47062 );
_HMUX g1747a ( \47064_nG1747a , \47063_nG17479 , 1'b0 , \47018 );
buf \U$38327 ( \47065 , \47064_nG1747a );
not \U$38328 ( \47066 , \47065 );
buf \U$38329 ( \47067 , RIe51f290_6359);
buf \U$38330 ( \47068 , RIe51e840_6360);
buf \U$38331 ( \47069 , RIe51dee0_6361);
and \U$38332 ( \47070 , \47068 , \47069 );
xor \U$38333 ( \47071 , \47067 , \47070 );
buf \U$38334 ( \47072 , \47071 );
buf \U$38335 ( \47073 , RIb839848_152);
and \U$38336 ( \47074 , \44813 , \47073 );
not \U$38337 ( \47075 , RIe51e840_6360);
and \U$38338 ( \47076 , RIe51dee0_6361, \47075 , RIe51f290_6359);
not \U$38339 ( \47077 , \47076 );
and \U$38340 ( \47078 , \47074 , \47077 );
_HMUX g17537 ( \47079_nG17537 , RIe51f290_6359 , \47072 , \47078 );
buf \U$38341 ( \47080 , RIe51f290_6359);
buf \U$38342 ( \47081 , RIe51e840_6360);
xor \U$38343 ( \47082 , \47080 , \47081 );
buf \U$38344 ( \47083 , \47082 );
not \U$38345 ( \47084 , RIe51dee0_6361);
and \U$38346 ( \47085 , \47084 , \47075 , RIe51f290_6359);
or \U$38347 ( \47086 , \47085 , \47076 );
_HMUX g1753b ( \47087_nG1753b , \47083 , RIe51f290_6359 , \47086 );
buf \U$38348 ( \47088 , RIb839668_156);
and \U$38349 ( \47089 , \44813 , \47088 );
_HMUX g1753c ( \47090_nG1753c , \47079_nG17537 , \47087_nG1753b , \47089 );
buf \U$38351 ( \47091 , RIb8396e0_155);
and \U$38352 ( \47092 , \44813 , \47091 );
_HMUX g1753d ( \47093_nG1753d , \47090_nG1753c , 1'b0 , \47092 );
and \U$38354 ( \47094 , \47092 , \47088 );
_HMUX g1753e ( \47095_nG1753e , \47093_nG1753d , 1'b0 , \47094 );
buf \U$38355 ( \47096 , \47095_nG1753e );
and \U$38356 ( \47097 , \47066 , \47096 );
xor \U$38357 ( \47098 , \47054 , \47055 );
buf \U$38358 ( \47099 , \47098 );
_HMUX g17473 ( \47100_nG17473 , RIe525d70_6348 , \47099 , \47062 );
_HMUX g17474 ( \47101_nG17474 , \47100_nG17473 , 1'b0 , \47018 );
buf \U$38360 ( \47102 , \47101_nG17474 );
not \U$38361 ( \47103 , \47102 );
xor \U$38362 ( \47104 , \47068 , \47069 );
buf \U$38363 ( \47105 , \47104 );
_HMUX g17528 ( \47106_nG17528 , RIe51e840_6360 , \47105 , \47078 );
not \U$38364 ( \47107 , \47081 );
buf \U$38365 ( \47108 , \47107 );
_HMUX g1752f ( \47109_nG1752f , \47108 , RIe51e840_6360 , \47086 );
_HMUX g17530 ( \47110_nG17530 , \47106_nG17528 , \47109_nG1752f , \47089 );
_HMUX g17531 ( \47111_nG17531 , \47110_nG17530 , 1'b0 , \47092 );
_HMUX g17532 ( \47112_nG17532 , \47111_nG17531 , 1'b1 , \47094 );
buf \U$38368 ( \47113 , \47112_nG17532 );
and \U$38369 ( \47114 , \47103 , \47113 );
not \U$38370 ( \47115 , \47055 );
buf \U$38371 ( \47116 , \47115 );
_HMUX g1746c ( \47117_nG1746c , RIe525410_6349 , \47116 , \47062 );
_HMUX g1746f ( \47118_nG1746f , \47117_nG1746c , 1'b0 , \47018 );
buf \U$38373 ( \47119 , \47118_nG1746f );
not \U$38374 ( \47120 , \47119 );
not \U$38375 ( \47121 , \47069 );
buf \U$38376 ( \47122 , \47121 );
_HMUX g17518 ( \47123_nG17518 , RIe51dee0_6361 , \47122 , \47078 );
buf \U$38377 ( \47124 , RIe51dee0_6361);
buf g1751c( \47125_nG1751c , \47124 );
_HMUX g1751f ( \47126_nG1751f , \47123_nG17518 , \47125_nG1751c , \47089 );
_HMUX g17522 ( \47127_nG17522 , \47126_nG1751f , 1'b1 , \47092 );
_HMUX g17524 ( \47128_nG17524 , \47127_nG17522 , 1'b0 , \47094 );
buf \U$38382 ( \47129 , \47128_nG17524 );
and \U$38383 ( \47130 , \47120 , \47129 );
xnor \U$38384 ( \47131 , \47113 , \47102 );
and \U$38385 ( \47132 , \47130 , \47131 );
or \U$38386 ( \47133 , \47114 , \47132 );
xnor \U$38387 ( \47134 , \47096 , \47065 );
and \U$38388 ( \47135 , \47133 , \47134 );
or \U$38389 ( \47136 , \47097 , \47135 );
buf \U$38390 ( \47137 , \47136 );
and \U$38391 ( \47138 , \47052 , \47137 );
not \U$38393 ( \47139 , \46926_nG175af );
or \U$38394 ( \47140 , \47139 , \47011 );
and \U$38395 ( \47141 , \47052 , \47140 );
_HMUX g175b3 ( \47142_nG175b3 , \47138 , 1'b1 , \47141 );
buf \U$38396 ( \47143 , \47142_nG175b3 );
_DC g190c4_GF_IsGateDCbyConstraint ( \47144_nG190c4 , \47143 , \42503 );
buf \U$38397 ( \47145 , \47144_nG190c4 );
buf \U$38398 ( \47146 , \47019_nG17498 );
_DC g19311_GF_IsGateDCbyConstraint ( \47147_nG19311 , \47146 , \42503 );
buf \U$38399 ( \47148 , \47147_nG19311 );
buf \U$38400 ( \47149 , \47033_nG174a5 );
_DC g19312_GF_IsGateDCbyConstraint ( \47150_nG19312 , \47149 , \42503 );
buf \U$38401 ( \47151 , \47150_nG19312 );
buf \U$38402 ( \47152 , \47049_nG174b4 );
_DC g19313_GF_IsGateDCbyConstraint ( \47153_nG19313 , \47152 , \42503 );
buf \U$38403 ( \47154 , \47153_nG19313 );
buf \U$38404 ( \47155 , RIb87eb00_69);
buf \U$38405 ( \47156 , RIe667bb0_6885);
buf \U$38406 ( \47157 , RIe667f70_6886);
nor \U$38407 ( \47158 , \47156 , \47157 );
_HMUX g1735d ( \47159_nG1735d , RIe1e2210_5688 , \47155 , \47158 );
not \U$38408 ( \47160 , RIea90778_6887);
and \U$38409 ( \47161 , \47160 , RIe546890_6849, RIe546098_6850, RIe545dc8_6851, \42389 );
buf \U$38410 ( \47162 , \47161 );
buf \U$38411 ( \47163 , \47162 );
buf \U$38412 ( \47164 , \42587 );
buf \U$38413 ( \47165 , \47164 );
and \U$38414 ( \47166 , \47163 , \47165 );
_HMUX g1735e ( \47167_nG1735e , RIe1e2210_5688 , \47159_nG1735d , \47166 );
buf \U$38415 ( \47168 , RIb7c5980_237);
buf \U$38416 ( \47169 , RIeab7058_6894);
buf \U$38417 ( \47170 , RIea91768_6889);
nor \U$38418 ( \47171 , \47169 , \47170 );
_HMUX g17360 ( \47172_nG17360 , RIe1e2210_5688 , \47168 , \47171 );
and \U$38419 ( \47173 , \44707 , \42169_nGbbec , \42218_nGbc1c , \42267_nGbc4c , \42316 );
buf \U$38420 ( \47174 , \47173 );
buf \U$38421 ( \47175 , \47174 );
buf \U$38422 ( \47176 , RIb79b518_270);
buf \U$38423 ( \47177 , \47176 );
and \U$38424 ( \47178 , \47175 , \47177 );
_HMUX g17361 ( \47179_nG17361 , \47167_nG1735e , \47172_nG17360 , \47178 );
buf \U$38425 ( \47180 , \47179_nG17361 );
_DC g19001_GF_IsGateDCbyConstraint ( \47181_nG19001 , \47180 , \42503 );
buf \U$38426 ( \47182 , \47181_nG19001 );
buf \U$38427 ( \47183 , RIb87eb78_68);
_HMUX g17362 ( \47184_nG17362 , RIe1e10b8_5689 , \47183 , \47158 );
_HMUX g17363 ( \47185_nG17363 , RIe1e10b8_5689 , \47184_nG17362 , \47166 );
buf \U$38428 ( \47186 , RIb7c59f8_236);
_HMUX g17364 ( \47187_nG17364 , RIe1e10b8_5689 , \47186 , \47171 );
_HMUX g17365 ( \47188_nG17365 , \47185_nG17363 , \47187_nG17364 , \47178 );
buf \U$38429 ( \47189 , \47188_nG17365 );
_DC g19017_GF_IsGateDCbyConstraint ( \47190_nG19017 , \47189 , \42503 );
buf \U$38430 ( \47191 , \47190_nG19017 );
buf \U$38431 ( \47192 , RIb87ebf0_67);
_HMUX g17366 ( \47193_nG17366 , RIe1dfab0_5690 , \47192 , \47158 );
_HMUX g17367 ( \47194_nG17367 , RIe1dfab0_5690 , \47193_nG17366 , \47166 );
buf \U$38432 ( \47195 , RIb7c5a70_235);
_HMUX g17368 ( \47196_nG17368 , RIe1dfab0_5690 , \47195 , \47171 );
_HMUX g17369 ( \47197_nG17369 , \47194_nG17367 , \47196_nG17368 , \47178 );
buf \U$38433 ( \47198 , \47197_nG17369 );
_DC g1902d_GF_IsGateDCbyConstraint ( \47199_nG1902d , \47198 , \42503 );
buf \U$38434 ( \47200 , \47199_nG1902d );
buf \U$38435 ( \47201 , RIb882ca0_66);
_HMUX g1736a ( \47202_nG1736a , RIe1de958_5691 , \47201 , \47158 );
_HMUX g1736b ( \47203_nG1736b , RIe1de958_5691 , \47202_nG1736a , \47166 );
buf \U$38436 ( \47204 , RIb7cade0_234);
_HMUX g1736c ( \47205_nG1736c , RIe1de958_5691 , \47204 , \47171 );
_HMUX g1736d ( \47206_nG1736d , \47203_nG1736b , \47205_nG1736c , \47178 );
buf \U$38437 ( \47207 , \47206_nG1736d );
_DC g19043_GF_IsGateDCbyConstraint ( \47208_nG19043 , \47207 , \42503 );
buf \U$38438 ( \47209 , \47208_nG19043 );
buf \U$38439 ( \47210 , RIb885310_65);
_HMUX g1736e ( \47211_nG1736e , RIe1dd350_5692 , \47210 , \47158 );
_HMUX g1736f ( \47212_nG1736f , RIe1dd350_5692 , \47211_nG1736e , \47166 );
buf \U$38440 ( \47213 , RIb7cae58_233);
_HMUX g17370 ( \47214_nG17370 , RIe1dd350_5692 , \47213 , \47171 );
_HMUX g17371 ( \47215_nG17371 , \47212_nG1736f , \47214_nG17370 , \47178 );
buf \U$38441 ( \47216 , \47215_nG17371 );
_DC g19059_GF_IsGateDCbyConstraint ( \47217_nG19059 , \47216 , \42503 );
buf \U$38442 ( \47218 , \47217_nG19059 );
buf \U$38443 ( \47219 , RIb885388_64);
_HMUX g17372 ( \47220_nG17372 , RIe1dc1f8_5693 , \47219 , \47158 );
_HMUX g17373 ( \47221_nG17373 , RIe1dc1f8_5693 , \47220_nG17372 , \47166 );
buf \U$38444 ( \47222 , RIb7caed0_232);
_HMUX g17374 ( \47223_nG17374 , RIe1dc1f8_5693 , \47222 , \47171 );
_HMUX g17375 ( \47224_nG17375 , \47221_nG17373 , \47223_nG17374 , \47178 );
buf \U$38445 ( \47225 , \47224_nG17375 );
_DC g1906f_GF_IsGateDCbyConstraint ( \47226_nG1906f , \47225 , \42503 );
buf \U$38446 ( \47227 , \47226_nG1906f );
buf \U$38447 ( \47228 , RIb885400_63);
_HMUX g17376 ( \47229_nG17376 , RIe1dabf0_5694 , \47228 , \47158 );
_HMUX g17377 ( \47230_nG17377 , RIe1dabf0_5694 , \47229_nG17376 , \47166 );
buf \U$38448 ( \47231 , RIb7caf48_231);
_HMUX g17378 ( \47232_nG17378 , RIe1dabf0_5694 , \47231 , \47171 );
_HMUX g17379 ( \47233_nG17379 , \47230_nG17377 , \47232_nG17378 , \47178 );
buf \U$38449 ( \47234 , \47233_nG17379 );
_DC g1907b_GF_IsGateDCbyConstraint ( \47235_nG1907b , \47234 , \42503 );
buf \U$38450 ( \47236 , \47235_nG1907b );
buf \U$38451 ( \47237 , RIb885478_62);
_HMUX g1737a ( \47238_nG1737a , RIe1d9a98_5695 , \47237 , \47158 );
_HMUX g1737b ( \47239_nG1737b , RIe1d9a98_5695 , \47238_nG1737a , \47166 );
buf \U$38452 ( \47240 , RIb7cafc0_230);
_HMUX g1737c ( \47241_nG1737c , RIe1d9a98_5695 , \47240 , \47171 );
_HMUX g1737d ( \47242_nG1737d , \47239_nG1737b , \47241_nG1737c , \47178 );
buf \U$38453 ( \47243 , \47242_nG1737d );
_DC g1907d_GF_IsGateDCbyConstraint ( \47244_nG1907d , \47243 , \42503 );
buf \U$38454 ( \47245 , \47244_nG1907d );
buf \U$38455 ( \47246 , RIb8854f0_61);
_HMUX g1737e ( \47247_nG1737e , RIe1d8940_5696 , \47246 , \47158 );
_HMUX g1737f ( \47248_nG1737f , RIe1d8940_5696 , \47247_nG1737e , \47166 );
buf \U$38456 ( \47249 , RIb7cb038_229);
_HMUX g17380 ( \47250_nG17380 , RIe1d8940_5696 , \47249 , \47171 );
_HMUX g17381 ( \47251_nG17381 , \47248_nG1737f , \47250_nG17380 , \47178 );
buf \U$38457 ( \47252 , \47251_nG17381 );
_DC g1907f_GF_IsGateDCbyConstraint ( \47253_nG1907f , \47252 , \42503 );
buf \U$38458 ( \47254 , \47253_nG1907f );
buf \U$38459 ( \47255 , RIb885568_60);
_HMUX g17382 ( \47256_nG17382 , RIe1d7338_5697 , \47255 , \47158 );
_HMUX g17383 ( \47257_nG17383 , RIe1d7338_5697 , \47256_nG17382 , \47166 );
buf \U$38460 ( \47258 , RIb7cb0b0_228);
_HMUX g17384 ( \47259_nG17384 , RIe1d7338_5697 , \47258 , \47171 );
_HMUX g17385 ( \47260_nG17385 , \47257_nG17383 , \47259_nG17384 , \47178 );
buf \U$38461 ( \47261 , \47260_nG17385 );
_DC g19003_GF_IsGateDCbyConstraint ( \47262_nG19003 , \47261 , \42503 );
buf \U$38462 ( \47263 , \47262_nG19003 );
buf \U$38463 ( \47264 , RIb8855e0_59);
_HMUX g17386 ( \47265_nG17386 , RIe1d61e0_5698 , \47264 , \47158 );
_HMUX g17387 ( \47266_nG17387 , RIe1d61e0_5698 , \47265_nG17386 , \47166 );
buf \U$38464 ( \47267 , RIb7cb128_227);
_HMUX g17388 ( \47268_nG17388 , RIe1d61e0_5698 , \47267 , \47171 );
_HMUX g17389 ( \47269_nG17389 , \47266_nG17387 , \47268_nG17388 , \47178 );
buf \U$38465 ( \47270 , \47269_nG17389 );
_DC g19005_GF_IsGateDCbyConstraint ( \47271_nG19005 , \47270 , \42503 );
buf \U$38466 ( \47272 , \47271_nG19005 );
buf \U$38467 ( \47273 , RIb885658_58);
_HMUX g1738a ( \47274_nG1738a , RIe1d4bd8_5699 , \47273 , \47158 );
_HMUX g1738b ( \47275_nG1738b , RIe1d4bd8_5699 , \47274_nG1738a , \47166 );
buf \U$38468 ( \47276 , RIb7d00d8_226);
_HMUX g1738c ( \47277_nG1738c , RIe1d4bd8_5699 , \47276 , \47171 );
_HMUX g1738d ( \47278_nG1738d , \47275_nG1738b , \47277_nG1738c , \47178 );
buf \U$38469 ( \47279 , \47278_nG1738d );
_DC g19007_GF_IsGateDCbyConstraint ( \47280_nG19007 , \47279 , \42503 );
buf \U$38470 ( \47281 , \47280_nG19007 );
buf \U$38471 ( \47282 , RIb8856d0_57);
_HMUX g1738e ( \47283_nG1738e , RIe1d3a80_5700 , \47282 , \47158 );
_HMUX g1738f ( \47284_nG1738f , RIe1d3a80_5700 , \47283_nG1738e , \47166 );
buf \U$38472 ( \47285 , RIb8263d8_225);
_HMUX g17390 ( \47286_nG17390 , RIe1d3a80_5700 , \47285 , \47171 );
_HMUX g17391 ( \47287_nG17391 , \47284_nG1738f , \47286_nG17390 , \47178 );
buf \U$38473 ( \47288 , \47287_nG17391 );
_DC g19009_GF_IsGateDCbyConstraint ( \47289_nG19009 , \47288 , \42503 );
buf \U$38474 ( \47290 , \47289_nG19009 );
buf \U$38475 ( \47291 , RIb885748_56);
_HMUX g17392 ( \47292_nG17392 , RIe1d2478_5701 , \47291 , \47158 );
_HMUX g17393 ( \47293_nG17393 , RIe1d2478_5701 , \47292_nG17392 , \47166 );
buf \U$38476 ( \47294 , RIb826e28_224);
_HMUX g17394 ( \47295_nG17394 , RIe1d2478_5701 , \47294 , \47171 );
_HMUX g17395 ( \47296_nG17395 , \47293_nG17393 , \47295_nG17394 , \47178 );
buf \U$38477 ( \47297 , \47296_nG17395 );
_DC g1900b_GF_IsGateDCbyConstraint ( \47298_nG1900b , \47297 , \42503 );
buf \U$38478 ( \47299 , \47298_nG1900b );
buf \U$38479 ( \47300 , RIb8857c0_55);
_HMUX g17396 ( \47301_nG17396 , RIe099530_5702 , \47300 , \47158 );
_HMUX g17397 ( \47302_nG17397 , RIe099530_5702 , \47301_nG17396 , \47166 );
buf \U$38480 ( \47303 , RIb826ea0_223);
_HMUX g17398 ( \47304_nG17398 , RIe099530_5702 , \47303 , \47171 );
_HMUX g17399 ( \47305_nG17399 , \47302_nG17397 , \47304_nG17398 , \47178 );
buf \U$38481 ( \47306 , \47305_nG17399 );
_DC g1900d_GF_IsGateDCbyConstraint ( \47307_nG1900d , \47306 , \42503 );
buf \U$38482 ( \47308 , \47307_nG1900d );
buf \U$38483 ( \47309 , RIb885838_54);
_HMUX g1739a ( \47310_nG1739a , RIe09d298_5703 , \47309 , \47158 );
_HMUX g1739b ( \47311_nG1739b , RIe09d298_5703 , \47310_nG1739a , \47166 );
buf \U$38484 ( \47312 , RIb826f18_222);
_HMUX g1739c ( \47313_nG1739c , RIe09d298_5703 , \47312 , \47171 );
_HMUX g1739d ( \47314_nG1739d , \47311_nG1739b , \47313_nG1739c , \47178 );
buf \U$38485 ( \47315 , \47314_nG1739d );
_DC g1900f_GF_IsGateDCbyConstraint ( \47316_nG1900f , \47315 , \42503 );
buf \U$38486 ( \47317 , \47316_nG1900f );
buf \U$38487 ( \47318 , RIb8858b0_53);
_HMUX g1739e ( \47319_nG1739e , RIe0a2338_5704 , \47318 , \47158 );
_HMUX g1739f ( \47320_nG1739f , RIe0a2338_5704 , \47319_nG1739e , \47166 );
buf \U$38488 ( \47321 , RIb826f90_221);
_HMUX g173a0 ( \47322_nG173a0 , RIe0a2338_5704 , \47321 , \47171 );
_HMUX g173a1 ( \47323_nG173a1 , \47320_nG1739f , \47322_nG173a0 , \47178 );
buf \U$38489 ( \47324 , \47323_nG173a1 );
_DC g19011_GF_IsGateDCbyConstraint ( \47325_nG19011 , \47324 , \42503 );
buf \U$38490 ( \47326 , \47325_nG19011 );
buf \U$38491 ( \47327 , RIb885928_52);
_HMUX g173a2 ( \47328_nG173a2 , RIe0a6fa0_5705 , \47327 , \47158 );
_HMUX g173a3 ( \47329_nG173a3 , RIe0a6fa0_5705 , \47328_nG173a2 , \47166 );
buf \U$38492 ( \47330 , RIb8293a8_220);
_HMUX g173a4 ( \47331_nG173a4 , RIe0a6fa0_5705 , \47330 , \47171 );
_HMUX g173a5 ( \47332_nG173a5 , \47329_nG173a3 , \47331_nG173a4 , \47178 );
buf \U$38493 ( \47333 , \47332_nG173a5 );
_DC g19013_GF_IsGateDCbyConstraint ( \47334_nG19013 , \47333 , \42503 );
buf \U$38494 ( \47335 , \47334_nG19013 );
buf \U$38495 ( \47336 , RIb8859a0_51);
_HMUX g173a6 ( \47337_nG173a6 , RIe0ac310_5706 , \47336 , \47158 );
_HMUX g173a7 ( \47338_nG173a7 , RIe0ac310_5706 , \47337_nG173a6 , \47166 );
buf \U$38496 ( \47339 , RIb829420_219);
_HMUX g173a8 ( \47340_nG173a8 , RIe0ac310_5706 , \47339 , \47171 );
_HMUX g173a9 ( \47341_nG173a9 , \47338_nG173a7 , \47340_nG173a8 , \47178 );
buf \U$38497 ( \47342 , \47341_nG173a9 );
_DC g19015_GF_IsGateDCbyConstraint ( \47343_nG19015 , \47342 , \42503 );
buf \U$38498 ( \47344 , \47343_nG19015 );
buf \U$38499 ( \47345 , RIb885a18_50);
_HMUX g173aa ( \47346_nG173aa , RIe0b16f8_5707 , \47345 , \47158 );
_HMUX g173ab ( \47347_nG173ab , RIe0b16f8_5707 , \47346_nG173aa , \47166 );
buf \U$38500 ( \47348 , RIb829498_218);
_HMUX g173ac ( \47349_nG173ac , RIe0b16f8_5707 , \47348 , \47171 );
_HMUX g173ad ( \47350_nG173ad , \47347_nG173ab , \47349_nG173ac , \47178 );
buf \U$38501 ( \47351 , \47350_nG173ad );
_DC g19019_GF_IsGateDCbyConstraint ( \47352_nG19019 , \47351 , \42503 );
buf \U$38502 ( \47353 , \47352_nG19019 );
buf \U$38503 ( \47354 , RIb885a90_49);
_HMUX g173ae ( \47355_nG173ae , RIe0b9240_5708 , \47354 , \47158 );
_HMUX g173af ( \47356_nG173af , RIe0b9240_5708 , \47355_nG173ae , \47166 );
buf \U$38504 ( \47357 , RIb829510_217);
_HMUX g173b0 ( \47358_nG173b0 , RIe0b9240_5708 , \47357 , \47171 );
_HMUX g173b1 ( \47359_nG173b1 , \47356_nG173af , \47358_nG173b0 , \47178 );
buf \U$38505 ( \47360 , \47359_nG173b1 );
_DC g1901b_GF_IsGateDCbyConstraint ( \47361_nG1901b , \47360 , \42503 );
buf \U$38506 ( \47362 , \47361_nG1901b );
buf \U$38507 ( \47363 , RIb885b08_48);
_HMUX g173b2 ( \47364_nG173b2 , RIe0bf438_5709 , \47363 , \47158 );
_HMUX g173b3 ( \47365_nG173b3 , RIe0bf438_5709 , \47364_nG173b2 , \47166 );
buf \U$38508 ( \47366 , RIb829588_216);
_HMUX g173b4 ( \47367_nG173b4 , RIe0bf438_5709 , \47366 , \47171 );
_HMUX g173b5 ( \47368_nG173b5 , \47365_nG173b3 , \47367_nG173b4 , \47178 );
buf \U$38509 ( \47369 , \47368_nG173b5 );
_DC g1901d_GF_IsGateDCbyConstraint ( \47370_nG1901d , \47369 , \42503 );
buf \U$38510 ( \47371 , \47370_nG1901d );
buf \U$38511 ( \47372 , RIb885b80_47);
_HMUX g173b6 ( \47373_nG173b6 , RIe0c4730_5710 , \47372 , \47158 );
_HMUX g173b7 ( \47374_nG173b7 , RIe0c4730_5710 , \47373_nG173b6 , \47166 );
buf \U$38512 ( \47375 , RIb829600_215);
_HMUX g173b8 ( \47376_nG173b8 , RIe0c4730_5710 , \47375 , \47171 );
_HMUX g173b9 ( \47377_nG173b9 , \47374_nG173b7 , \47376_nG173b8 , \47178 );
buf \U$38513 ( \47378 , \47377_nG173b9 );
_DC g1901f_GF_IsGateDCbyConstraint ( \47379_nG1901f , \47378 , \42503 );
buf \U$38514 ( \47380 , \47379_nG1901f );
buf \U$38515 ( \47381 , RIb885bf8_46);
_HMUX g173ba ( \47382_nG173ba , RIe0cb0a8_5711 , \47381 , \47158 );
_HMUX g173bb ( \47383_nG173bb , RIe0cb0a8_5711 , \47382_nG173ba , \47166 );
buf \U$38516 ( \47384 , RIb829678_214);
_HMUX g173bc ( \47385_nG173bc , RIe0cb0a8_5711 , \47384 , \47171 );
_HMUX g173bd ( \47386_nG173bd , \47383_nG173bb , \47385_nG173bc , \47178 );
buf \U$38517 ( \47387 , \47386_nG173bd );
_DC g19021_GF_IsGateDCbyConstraint ( \47388_nG19021 , \47387 , \42503 );
buf \U$38518 ( \47389 , \47388_nG19021 );
buf \U$38519 ( \47390 , RIb885c70_45);
_HMUX g173be ( \47391_nG173be , RIe0d0df0_5712 , \47390 , \47158 );
_HMUX g173bf ( \47392_nG173bf , RIe0d0df0_5712 , \47391_nG173be , \47166 );
buf \U$38520 ( \47393 , RIb8296f0_213);
_HMUX g173c0 ( \47394_nG173c0 , RIe0d0df0_5712 , \47393 , \47171 );
_HMUX g173c1 ( \47395_nG173c1 , \47392_nG173bf , \47394_nG173c0 , \47178 );
buf \U$38521 ( \47396 , \47395_nG173c1 );
_DC g19023_GF_IsGateDCbyConstraint ( \47397_nG19023 , \47396 , \42503 );
buf \U$38522 ( \47398 , \47397_nG19023 );
buf \U$38523 ( \47399 , RIb885ce8_44);
_HMUX g173c2 ( \47400_nG173c2 , RIe0d8aa0_5713 , \47399 , \47158 );
_HMUX g173c3 ( \47401_nG173c3 , RIe0d8aa0_5713 , \47400_nG173c2 , \47166 );
buf \U$38524 ( \47402 , RIb82dae8_212);
_HMUX g173c4 ( \47403_nG173c4 , RIe0d8aa0_5713 , \47402 , \47171 );
_HMUX g173c5 ( \47404_nG173c5 , \47401_nG173c3 , \47403_nG173c4 , \47178 );
buf \U$38525 ( \47405 , \47404_nG173c5 );
_DC g19025_GF_IsGateDCbyConstraint ( \47406_nG19025 , \47405 , \42503 );
buf \U$38526 ( \47407 , \47406_nG19025 );
buf \U$38527 ( \47408 , RIb885d60_43);
_HMUX g173c6 ( \47409_nG173c6 , RIe0de608_5714 , \47408 , \47158 );
_HMUX g173c7 ( \47410_nG173c7 , RIe0de608_5714 , \47409_nG173c6 , \47166 );
buf \U$38528 ( \47411 , RIb82db60_211);
_HMUX g173c8 ( \47412_nG173c8 , RIe0de608_5714 , \47411 , \47171 );
_HMUX g173c9 ( \47413_nG173c9 , \47410_nG173c7 , \47412_nG173c8 , \47178 );
buf \U$38529 ( \47414 , \47413_nG173c9 );
_DC g19027_GF_IsGateDCbyConstraint ( \47415_nG19027 , \47414 , \42503 );
buf \U$38530 ( \47416 , \47415_nG19027 );
buf \U$38531 ( \47417 , RIb885dd8_42);
_HMUX g173ca ( \47418_nG173ca , RIe0e5ca0_5715 , \47417 , \47158 );
_HMUX g173cb ( \47419_nG173cb , RIe0e5ca0_5715 , \47418_nG173ca , \47166 );
buf \U$38532 ( \47420 , RIb82dbd8_210);
_HMUX g173cc ( \47421_nG173cc , RIe0e5ca0_5715 , \47420 , \47171 );
_HMUX g173cd ( \47422_nG173cd , \47419_nG173cb , \47421_nG173cc , \47178 );
buf \U$38533 ( \47423 , \47422_nG173cd );
_DC g19029_GF_IsGateDCbyConstraint ( \47424_nG19029 , \47423 , \42503 );
buf \U$38534 ( \47425 , \47424_nG19029 );
buf \U$38535 ( \47426 , RIb885e50_41);
_HMUX g173ce ( \47427_nG173ce , RIe0eb358_5716 , \47426 , \47158 );
_HMUX g173cf ( \47428_nG173cf , RIe0eb358_5716 , \47427_nG173ce , \47166 );
buf \U$38536 ( \47429 , RIb82dc50_209);
_HMUX g173d0 ( \47430_nG173d0 , RIe0eb358_5716 , \47429 , \47171 );
_HMUX g173d1 ( \47431_nG173d1 , \47428_nG173cf , \47430_nG173d0 , \47178 );
buf \U$38537 ( \47432 , \47431_nG173d1 );
_DC g1902b_GF_IsGateDCbyConstraint ( \47433_nG1902b , \47432 , \42503 );
buf \U$38538 ( \47434 , \47433_nG1902b );
buf \U$38539 ( \47435 , RIb885ec8_40);
_HMUX g173d2 ( \47436_nG173d2 , RIe0ef138_5717 , \47435 , \47158 );
_HMUX g173d3 ( \47437_nG173d3 , RIe0ef138_5717 , \47436_nG173d2 , \47166 );
buf \U$38540 ( \47438 , RIb82dcc8_208);
_HMUX g173d4 ( \47439_nG173d4 , RIe0ef138_5717 , \47438 , \47171 );
_HMUX g173d5 ( \47440_nG173d5 , \47437_nG173d3 , \47439_nG173d4 , \47178 );
buf \U$38541 ( \47441 , \47440_nG173d5 );
_DC g1902f_GF_IsGateDCbyConstraint ( \47442_nG1902f , \47441 , \42503 );
buf \U$38542 ( \47443 , \47442_nG1902f );
buf \U$38543 ( \47444 , RIb885f40_39);
_HMUX g173d6 ( \47445_nG173d6 , RIe0f3bc0_5718 , \47444 , \47158 );
_HMUX g173d7 ( \47446_nG173d7 , RIe0f3bc0_5718 , \47445_nG173d6 , \47166 );
buf \U$38544 ( \47447 , RIb82dd40_207);
_HMUX g173d8 ( \47448_nG173d8 , RIe0f3bc0_5718 , \47447 , \47171 );
_HMUX g173d9 ( \47449_nG173d9 , \47446_nG173d7 , \47448_nG173d8 , \47178 );
buf \U$38545 ( \47450 , \47449_nG173d9 );
_DC g19031_GF_IsGateDCbyConstraint ( \47451_nG19031 , \47450 , \42503 );
buf \U$38546 ( \47452 , \47451_nG19031 );
buf \U$38547 ( \47453 , RIb885fb8_38);
_HMUX g173da ( \47454_nG173da , RIe0f8300_5719 , \47453 , \47158 );
_HMUX g173db ( \47455_nG173db , RIe0f8300_5719 , \47454_nG173da , \47166 );
buf \U$38548 ( \47456 , RIb82ddb8_206);
_HMUX g173dc ( \47457_nG173dc , RIe0f8300_5719 , \47456 , \47171 );
_HMUX g173dd ( \47458_nG173dd , \47455_nG173db , \47457_nG173dc , \47178 );
buf \U$38549 ( \47459 , \47458_nG173dd );
_DC g19033_GF_IsGateDCbyConstraint ( \47460_nG19033 , \47459 , \42503 );
buf \U$38550 ( \47461 , \47460_nG19033 );
buf \U$38551 ( \47462 , RIb886030_37);
_HMUX g173de ( \47463_nG173de , RIe0ff380_5720 , \47462 , \47158 );
_HMUX g173df ( \47464_nG173df , RIe0ff380_5720 , \47463_nG173de , \47166 );
buf \U$38552 ( \47465 , RIb82de30_205);
_HMUX g173e0 ( \47466_nG173e0 , RIe0ff380_5720 , \47465 , \47171 );
_HMUX g173e1 ( \47467_nG173e1 , \47464_nG173df , \47466_nG173e0 , \47178 );
buf \U$38553 ( \47468 , \47467_nG173e1 );
_DC g19035_GF_IsGateDCbyConstraint ( \47469_nG19035 , \47468 , \42503 );
buf \U$38554 ( \47470 , \47469_nG19035 );
buf \U$38555 ( \47471 , RIb8860a8_36);
_HMUX g173e2 ( \47472_nG173e2 , RIe103430_5721 , \47471 , \47158 );
_HMUX g173e3 ( \47473_nG173e3 , RIe103430_5721 , \47472_nG173e2 , \47166 );
buf \U$38556 ( \47474 , RIb832228_204);
_HMUX g173e4 ( \47475_nG173e4 , RIe103430_5721 , \47474 , \47171 );
_HMUX g173e5 ( \47476_nG173e5 , \47473_nG173e3 , \47475_nG173e4 , \47178 );
buf \U$38557 ( \47477 , \47476_nG173e5 );
_DC g19037_GF_IsGateDCbyConstraint ( \47478_nG19037 , \47477 , \42503 );
buf \U$38558 ( \47479 , \47478_nG19037 );
buf \U$38559 ( \47480 , RIb886120_35);
_HMUX g173e6 ( \47481_nG173e6 , RIdfce868_5722 , \47480 , \47158 );
_HMUX g173e7 ( \47482_nG173e7 , RIdfce868_5722 , \47481_nG173e6 , \47166 );
buf \U$38560 ( \47483 , RIb8322a0_203);
_HMUX g173e8 ( \47484_nG173e8 , RIdfce868_5722 , \47483 , \47171 );
_HMUX g173e9 ( \47485_nG173e9 , \47482_nG173e7 , \47484_nG173e8 , \47178 );
buf \U$38561 ( \47486 , \47485_nG173e9 );
_DC g19039_GF_IsGateDCbyConstraint ( \47487_nG19039 , \47486 , \42503 );
buf \U$38562 ( \47488 , \47487_nG19039 );
buf \U$38563 ( \47489 , RIb886198_34);
_HMUX g173ea ( \47490_nG173ea , RIdfc9fc0_5723 , \47489 , \47158 );
_HMUX g173eb ( \47491_nG173eb , RIdfc9fc0_5723 , \47490_nG173ea , \47166 );
buf \U$38564 ( \47492 , RIb832318_202);
_HMUX g173ec ( \47493_nG173ec , RIdfc9fc0_5723 , \47492 , \47171 );
_HMUX g173ed ( \47494_nG173ed , \47491_nG173eb , \47493_nG173ec , \47178 );
buf \U$38565 ( \47495 , \47494_nG173ed );
_DC g1903b_GF_IsGateDCbyConstraint ( \47496_nG1903b , \47495 , \42503 );
buf \U$38566 ( \47497 , \47496_nG1903b );
buf \U$38567 ( \47498 , RIb886210_33);
_HMUX g173ee ( \47499_nG173ee , RIdfc6000_5724 , \47498 , \47158 );
_HMUX g173ef ( \47500_nG173ef , RIdfc6000_5724 , \47499_nG173ee , \47166 );
buf \U$38568 ( \47501 , RIb832390_201);
_HMUX g173f0 ( \47502_nG173f0 , RIdfc6000_5724 , \47501 , \47171 );
_HMUX g173f1 ( \47503_nG173f1 , \47500_nG173ef , \47502_nG173f0 , \47178 );
buf \U$38569 ( \47504 , \47503_nG173f1 );
_DC g1903d_GF_IsGateDCbyConstraint ( \47505_nG1903d , \47504 , \42503 );
buf \U$38570 ( \47506 , \47505_nG1903d );
buf \U$38571 ( \47507 , RIb886288_32);
_HMUX g173f2 ( \47508_nG173f2 , RIdfc1410_5725 , \47507 , \47158 );
_HMUX g173f3 ( \47509_nG173f3 , RIdfc1410_5725 , \47508_nG173f2 , \47166 );
buf \U$38572 ( \47510 , RIb832408_200);
_HMUX g173f4 ( \47511_nG173f4 , RIdfc1410_5725 , \47510 , \47171 );
_HMUX g173f5 ( \47512_nG173f5 , \47509_nG173f3 , \47511_nG173f4 , \47178 );
buf \U$38573 ( \47513 , \47512_nG173f5 );
_DC g1903f_GF_IsGateDCbyConstraint ( \47514_nG1903f , \47513 , \42503 );
buf \U$38574 ( \47515 , \47514_nG1903f );
buf \U$38575 ( \47516 , RIb886300_31);
_HMUX g173f6 ( \47517_nG173f6 , RIdfbcc58_5726 , \47516 , \47158 );
_HMUX g173f7 ( \47518_nG173f7 , RIdfbcc58_5726 , \47517_nG173f6 , \47166 );
buf \U$38576 ( \47519 , RIb832480_199);
_HMUX g173f8 ( \47520_nG173f8 , RIdfbcc58_5726 , \47519 , \47171 );
_HMUX g173f9 ( \47521_nG173f9 , \47518_nG173f7 , \47520_nG173f8 , \47178 );
buf \U$38577 ( \47522 , \47521_nG173f9 );
_DC g19041_GF_IsGateDCbyConstraint ( \47523_nG19041 , \47522 , \42503 );
buf \U$38578 ( \47524 , \47523_nG19041 );
buf \U$38579 ( \47525 , RIb886378_30);
_HMUX g173fa ( \47526_nG173fa , RIe082f10_5727 , \47525 , \47158 );
_HMUX g173fb ( \47527_nG173fb , RIe082f10_5727 , \47526_nG173fa , \47166 );
buf \U$38580 ( \47528 , RIb8324f8_198);
_HMUX g173fc ( \47529_nG173fc , RIe082f10_5727 , \47528 , \47171 );
_HMUX g173fd ( \47530_nG173fd , \47527_nG173fb , \47529_nG173fc , \47178 );
buf \U$38581 ( \47531 , \47530_nG173fd );
_DC g19045_GF_IsGateDCbyConstraint ( \47532_nG19045 , \47531 , \42503 );
buf \U$38582 ( \47533 , \47532_nG19045 );
buf \U$38583 ( \47534 , RIb8863f0_29);
_HMUX g173fe ( \47535_nG173fe , RIe0800a8_5728 , \47534 , \47158 );
_HMUX g173ff ( \47536_nG173ff , RIe0800a8_5728 , \47535_nG173fe , \47166 );
buf \U$38584 ( \47537 , RIb832570_197);
_HMUX g17400 ( \47538_nG17400 , RIe0800a8_5728 , \47537 , \47171 );
_HMUX g17401 ( \47539_nG17401 , \47536_nG173ff , \47538_nG17400 , \47178 );
buf \U$38585 ( \47540 , \47539_nG17401 );
_DC g19047_GF_IsGateDCbyConstraint ( \47541_nG19047 , \47540 , \42503 );
buf \U$38586 ( \47542 , \47541_nG19047 );
buf \U$38587 ( \47543 , RIb886468_28);
_HMUX g17402 ( \47544_nG17402 , RIe07bd28_5729 , \47543 , \47158 );
_HMUX g17403 ( \47545_nG17403 , RIe07bd28_5729 , \47544_nG17402 , \47166 );
buf \U$38588 ( \47546 , RIb8383a8_196);
_HMUX g17404 ( \47547_nG17404 , RIe07bd28_5729 , \47546 , \47171 );
_HMUX g17405 ( \47548_nG17405 , \47545_nG17403 , \47547_nG17404 , \47178 );
buf \U$38589 ( \47549 , \47548_nG17405 );
_DC g19049_GF_IsGateDCbyConstraint ( \47550_nG19049 , \47549 , \42503 );
buf \U$38590 ( \47551 , \47550_nG19049 );
buf \U$38591 ( \47552 , RIb8864e0_27);
_HMUX g17406 ( \47553_nG17406 , RIe078ec0_5730 , \47552 , \47158 );
_HMUX g17407 ( \47554_nG17407 , RIe078ec0_5730 , \47553_nG17406 , \47166 );
buf \U$38592 ( \47555 , RIb838420_195);
_HMUX g17408 ( \47556_nG17408 , RIe078ec0_5730 , \47555 , \47171 );
_HMUX g17409 ( \47557_nG17409 , \47554_nG17407 , \47556_nG17408 , \47178 );
buf \U$38593 ( \47558 , \47557_nG17409 );
_DC g1904b_GF_IsGateDCbyConstraint ( \47559_nG1904b , \47558 , \42503 );
buf \U$38594 ( \47560 , \47559_nG1904b );
buf \U$38595 ( \47561 , RIb886558_26);
_HMUX g1740a ( \47562_nG1740a , RIe075ab8_5731 , \47561 , \47158 );
_HMUX g1740b ( \47563_nG1740b , RIe075ab8_5731 , \47562_nG1740a , \47166 );
buf \U$38596 ( \47564 , RIb838498_194);
_HMUX g1740c ( \47565_nG1740c , RIe075ab8_5731 , \47564 , \47171 );
_HMUX g1740d ( \47566_nG1740d , \47563_nG1740b , \47565_nG1740c , \47178 );
buf \U$38597 ( \47567 , \47566_nG1740d );
_DC g1904d_GF_IsGateDCbyConstraint ( \47568_nG1904d , \47567 , \42503 );
buf \U$38598 ( \47569 , \47568_nG1904d );
buf \U$38599 ( \47570 , RIb8865d0_25);
_HMUX g1740e ( \47571_nG1740e , RIe071f18_5732 , \47570 , \47158 );
_HMUX g1740f ( \47572_nG1740f , RIe071f18_5732 , \47571_nG1740e , \47166 );
buf \U$38600 ( \47573 , RIb838510_193);
_HMUX g17410 ( \47574_nG17410 , RIe071f18_5732 , \47573 , \47171 );
_HMUX g17411 ( \47575_nG17411 , \47572_nG1740f , \47574_nG17410 , \47178 );
buf \U$38601 ( \47576 , \47575_nG17411 );
_DC g1904f_GF_IsGateDCbyConstraint ( \47577_nG1904f , \47576 , \42503 );
buf \U$38602 ( \47578 , \47577_nG1904f );
buf \U$38603 ( \47579 , RIb886648_24);
_HMUX g17412 ( \47580_nG17412 , RIe06f308_5733 , \47579 , \47158 );
_HMUX g17413 ( \47581_nG17413 , RIe06f308_5733 , \47580_nG17412 , \47166 );
buf \U$38604 ( \47582 , RIb838588_192);
_HMUX g17414 ( \47583_nG17414 , RIe06f308_5733 , \47582 , \47171 );
_HMUX g17415 ( \47584_nG17415 , \47581_nG17413 , \47583_nG17414 , \47178 );
buf \U$38605 ( \47585 , \47584_nG17415 );
_DC g19051_GF_IsGateDCbyConstraint ( \47586_nG19051 , \47585 , \42503 );
buf \U$38606 ( \47587 , \47586_nG19051 );
buf \U$38607 ( \47588 , RIb8866c0_23);
_HMUX g17416 ( \47589_nG17416 , RIe06b0f0_5734 , \47588 , \47158 );
_HMUX g17417 ( \47590_nG17417 , RIe06b0f0_5734 , \47589_nG17416 , \47166 );
buf \U$38608 ( \47591 , RIb838600_191);
_HMUX g17418 ( \47592_nG17418 , RIe06b0f0_5734 , \47591 , \47171 );
_HMUX g17419 ( \47593_nG17419 , \47590_nG17417 , \47592_nG17418 , \47178 );
buf \U$38609 ( \47594 , \47593_nG17419 );
_DC g19053_GF_IsGateDCbyConstraint ( \47595_nG19053 , \47594 , \42503 );
buf \U$38610 ( \47596 , \47595_nG19053 );
buf \U$38611 ( \47597 , RIb886738_22);
_HMUX g1741a ( \47598_nG1741a , RIe067928_5735 , \47597 , \47158 );
_HMUX g1741b ( \47599_nG1741b , RIe067928_5735 , \47598_nG1741a , \47166 );
buf \U$38612 ( \47600 , RIb838678_190);
_HMUX g1741c ( \47601_nG1741c , RIe067928_5735 , \47600 , \47171 );
_HMUX g1741d ( \47602_nG1741d , \47599_nG1741b , \47601_nG1741c , \47178 );
buf \U$38613 ( \47603 , \47602_nG1741d );
_DC g19055_GF_IsGateDCbyConstraint ( \47604_nG19055 , \47603 , \42503 );
buf \U$38614 ( \47605 , \47604_nG19055 );
buf \U$38615 ( \47606 , RIb8867b0_21);
_HMUX g1741e ( \47607_nG1741e , RIe0608a8_5736 , \47606 , \47158 );
_HMUX g1741f ( \47608_nG1741f , RIe0608a8_5736 , \47607_nG1741e , \47166 );
buf \U$38616 ( \47609 , RIb8386f0_189);
_HMUX g17420 ( \47610_nG17420 , RIe0608a8_5736 , \47609 , \47171 );
_HMUX g17421 ( \47611_nG17421 , \47608_nG1741f , \47610_nG17420 , \47178 );
buf \U$38617 ( \47612 , \47611_nG17421 );
_DC g19057_GF_IsGateDCbyConstraint ( \47613_nG19057 , \47612 , \42503 );
buf \U$38618 ( \47614 , \47613_nG19057 );
buf \U$38619 ( \47615 , RIb886828_20);
_HMUX g17422 ( \47616_nG17422 , RIe05a2f0_5737 , \47615 , \47158 );
_HMUX g17423 ( \47617_nG17423 , RIe05a2f0_5737 , \47616_nG17422 , \47166 );
buf \U$38620 ( \47618 , RIb838768_188);
_HMUX g17424 ( \47619_nG17424 , RIe05a2f0_5737 , \47618 , \47171 );
_HMUX g17425 ( \47620_nG17425 , \47617_nG17423 , \47619_nG17424 , \47178 );
buf \U$38621 ( \47621 , \47620_nG17425 );
_DC g1905b_GF_IsGateDCbyConstraint ( \47622_nG1905b , \47621 , \42503 );
buf \U$38622 ( \47623 , \47622_nG1905b );
buf \U$38623 ( \47624 , RIb8868a0_19);
_HMUX g17426 ( \47625_nG17426 , RIe0541e8_5738 , \47624 , \47158 );
_HMUX g17427 ( \47626_nG17427 , RIe0541e8_5738 , \47625_nG17426 , \47166 );
buf \U$38624 ( \47627 , RIb8387e0_187);
_HMUX g17428 ( \47628_nG17428 , RIe0541e8_5738 , \47627 , \47171 );
_HMUX g17429 ( \47629_nG17429 , \47626_nG17427 , \47628_nG17428 , \47178 );
buf \U$38625 ( \47630 , \47629_nG17429 );
_DC g1905d_GF_IsGateDCbyConstraint ( \47631_nG1905d , \47630 , \42503 );
buf \U$38626 ( \47632 , \47631_nG1905d );
buf \U$38627 ( \47633 , RIb886918_18);
_HMUX g1742a ( \47634_nG1742a , RIe04bb60_5739 , \47633 , \47158 );
_HMUX g1742b ( \47635_nG1742b , RIe04bb60_5739 , \47634_nG1742a , \47166 );
buf \U$38628 ( \47636 , RIb838858_186);
_HMUX g1742c ( \47637_nG1742c , RIe04bb60_5739 , \47636 , \47171 );
_HMUX g1742d ( \47638_nG1742d , \47635_nG1742b , \47637_nG1742c , \47178 );
buf \U$38629 ( \47639 , \47638_nG1742d );
_DC g1905f_GF_IsGateDCbyConstraint ( \47640_nG1905f , \47639 , \42503 );
buf \U$38630 ( \47641 , \47640_nG1905f );
buf \U$38631 ( \47642 , RIb886990_17);
_HMUX g1742e ( \47643_nG1742e , RIe045a58_5740 , \47642 , \47158 );
_HMUX g1742f ( \47644_nG1742f , RIe045a58_5740 , \47643_nG1742e , \47166 );
buf \U$38632 ( \47645 , RIb8388d0_185);
_HMUX g17430 ( \47646_nG17430 , RIe045a58_5740 , \47645 , \47171 );
_HMUX g17431 ( \47647_nG17431 , \47644_nG1742f , \47646_nG17430 , \47178 );
buf \U$38633 ( \47648 , \47647_nG17431 );
_DC g19061_GF_IsGateDCbyConstraint ( \47649_nG19061 , \47648 , \42503 );
buf \U$38634 ( \47650 , \47649_nG19061 );
buf \U$38635 ( \47651 , RIb886a08_16);
_HMUX g17432 ( \47652_nG17432 , RIe03d3d0_5741 , \47651 , \47158 );
_HMUX g17433 ( \47653_nG17433 , RIe03d3d0_5741 , \47652_nG17432 , \47166 );
buf \U$38636 ( \47654 , RIb838948_184);
_HMUX g17434 ( \47655_nG17434 , RIe03d3d0_5741 , \47654 , \47171 );
_HMUX g17435 ( \47656_nG17435 , \47653_nG17433 , \47655_nG17434 , \47178 );
buf \U$38637 ( \47657 , \47656_nG17435 );
_DC g19063_GF_IsGateDCbyConstraint ( \47658_nG19063 , \47657 , \42503 );
buf \U$38638 ( \47659 , \47658_nG19063 );
buf \U$38639 ( \47660 , RIb886a80_15);
_HMUX g17436 ( \47661_nG17436 , RIde1d908_5742 , \47660 , \47158 );
_HMUX g17437 ( \47662_nG17437 , RIde1d908_5742 , \47661_nG17436 , \47166 );
buf \U$38640 ( \47663 , RIb8389c0_183);
_HMUX g17438 ( \47664_nG17438 , RIde1d908_5742 , \47663 , \47171 );
_HMUX g17439 ( \47665_nG17439 , \47662_nG17437 , \47664_nG17438 , \47178 );
buf \U$38641 ( \47666 , \47665_nG17439 );
_DC g19065_GF_IsGateDCbyConstraint ( \47667_nG19065 , \47666 , \42503 );
buf \U$38642 ( \47668 , \47667_nG19065 );
buf \U$38643 ( \47669 , RIb886af8_14);
_HMUX g1743a ( \47670_nG1743a , RIde4a200_5743 , \47669 , \47158 );
_HMUX g1743b ( \47671_nG1743b , RIde4a200_5743 , \47670_nG1743a , \47166 );
buf \U$38644 ( \47672 , RIb838a38_182);
_HMUX g1743c ( \47673_nG1743c , RIde4a200_5743 , \47672 , \47171 );
_HMUX g1743d ( \47674_nG1743d , \47671_nG1743b , \47673_nG1743c , \47178 );
buf \U$38645 ( \47675 , \47674_nG1743d );
_DC g19067_GF_IsGateDCbyConstraint ( \47676_nG19067 , \47675 , \42503 );
buf \U$38646 ( \47677 , \47676_nG19067 );
buf \U$38647 ( \47678 , RIb886b70_13);
_HMUX g1743e ( \47679_nG1743e , RIde62e18_5744 , \47678 , \47158 );
_HMUX g1743f ( \47680_nG1743f , RIde62e18_5744 , \47679_nG1743e , \47166 );
buf \U$38648 ( \47681 , RIb838ab0_181);
_HMUX g17440 ( \47682_nG17440 , RIde62e18_5744 , \47681 , \47171 );
_HMUX g17441 ( \47683_nG17441 , \47680_nG1743f , \47682_nG17440 , \47178 );
buf \U$38649 ( \47684 , \47683_nG17441 );
_DC g19069_GF_IsGateDCbyConstraint ( \47685_nG19069 , \47684 , \42503 );
buf \U$38650 ( \47686 , \47685_nG19069 );
buf \U$38651 ( \47687 , RIb886be8_12);
_HMUX g17442 ( \47688_nG17442 , RIdc30d68_5745 , \47687 , \47158 );
_HMUX g17443 ( \47689_nG17443 , RIdc30d68_5745 , \47688_nG17442 , \47166 );
buf \U$38652 ( \47690 , RIb838b28_180);
_HMUX g17444 ( \47691_nG17444 , RIdc30d68_5745 , \47690 , \47171 );
_HMUX g17445 ( \47692_nG17445 , \47689_nG17443 , \47691_nG17444 , \47178 );
buf \U$38653 ( \47693 , \47692_nG17445 );
_DC g1906b_GF_IsGateDCbyConstraint ( \47694_nG1906b , \47693 , \42503 );
buf \U$38654 ( \47695 , \47694_nG1906b );
buf \U$38655 ( \47696 , RIb886c60_11);
_HMUX g17446 ( \47697_nG17446 , RIdde3e10_5746 , \47696 , \47158 );
_HMUX g17447 ( \47698_nG17447 , RIdde3e10_5746 , \47697_nG17446 , \47166 );
buf \U$38656 ( \47699 , RIb838ba0_179);
_HMUX g17448 ( \47700_nG17448 , RIdde3e10_5746 , \47699 , \47171 );
_HMUX g17449 ( \47701_nG17449 , \47698_nG17447 , \47700_nG17448 , \47178 );
buf \U$38657 ( \47702 , \47701_nG17449 );
_DC g1906d_GF_IsGateDCbyConstraint ( \47703_nG1906d , \47702 , \42503 );
buf \U$38658 ( \47704 , \47703_nG1906d );
buf \U$38659 ( \47705 , RIb886cd8_10);
_HMUX g1744a ( \47706_nG1744a , RIddce948_5747 , \47705 , \47158 );
_HMUX g1744b ( \47707_nG1744b , RIddce948_5747 , \47706_nG1744a , \47166 );
buf \U$38660 ( \47708 , RIb838c18_178);
_HMUX g1744c ( \47709_nG1744c , RIddce948_5747 , \47708 , \47171 );
_HMUX g1744d ( \47710_nG1744d , \47707_nG1744b , \47709_nG1744c , \47178 );
buf \U$38661 ( \47711 , \47710_nG1744d );
_DC g19071_GF_IsGateDCbyConstraint ( \47712_nG19071 , \47711 , \42503 );
buf \U$38662 ( \47713 , \47712_nG19071 );
buf \U$38663 ( \47714 , RIb886d50_9);
_HMUX g1744e ( \47715_nG1744e , RIdb96b50_5748 , \47714 , \47158 );
_HMUX g1744f ( \47716_nG1744f , RIdb96b50_5748 , \47715_nG1744e , \47166 );
buf \U$38664 ( \47717 , RIb838c90_177);
_HMUX g17450 ( \47718_nG17450 , RIdb96b50_5748 , \47717 , \47171 );
_HMUX g17451 ( \47719_nG17451 , \47716_nG1744f , \47718_nG17450 , \47178 );
buf \U$38665 ( \47720 , \47719_nG17451 );
_DC g19073_GF_IsGateDCbyConstraint ( \47721_nG19073 , \47720 , \42503 );
buf \U$38666 ( \47722 , \47721_nG19073 );
buf \U$38667 ( \47723 , RIb886dc8_8);
_HMUX g17452 ( \47724_nG17452 , RIda0b300_5749 , \47723 , \47158 );
_HMUX g17453 ( \47725_nG17453 , RIda0b300_5749 , \47724_nG17452 , \47166 );
buf \U$38668 ( \47726 , RIb838d08_176);
_HMUX g17454 ( \47727_nG17454 , RIda0b300_5749 , \47726 , \47171 );
_HMUX g17455 ( \47728_nG17455 , \47725_nG17453 , \47727_nG17454 , \47178 );
buf \U$38669 ( \47729 , \47728_nG17455 );
_DC g19075_GF_IsGateDCbyConstraint ( \47730_nG19075 , \47729 , \42503 );
buf \U$38670 ( \47731 , \47730_nG19075 );
buf \U$38671 ( \47732 , RIb886e40_7);
_HMUX g17456 ( \47733_nG17456 , RIdc00960_5750 , \47732 , \47158 );
_HMUX g17457 ( \47734_nG17457 , RIdc00960_5750 , \47733_nG17456 , \47166 );
buf \U$38672 ( \47735 , RIb838d80_175);
_HMUX g17458 ( \47736_nG17458 , RIdc00960_5750 , \47735 , \47171 );
_HMUX g17459 ( \47737_nG17459 , \47734_nG17457 , \47736_nG17458 , \47178 );
buf \U$38673 ( \47738 , \47737_nG17459 );
_DC g19077_GF_IsGateDCbyConstraint ( \47739_nG19077 , \47738 , \42503 );
buf \U$38674 ( \47740 , \47739_nG19077 );
buf \U$38675 ( \47741 , RIb886eb8_6);
_HMUX g1745a ( \47742_nG1745a , RIdb708e8_5751 , \47741 , \47158 );
_HMUX g1745b ( \47743_nG1745b , RIdb708e8_5751 , \47742_nG1745a , \47166 );
buf \U$38676 ( \47744 , RIb838df8_174);
_HMUX g1745c ( \47745_nG1745c , RIdb708e8_5751 , \47744 , \47171 );
_HMUX g1745d ( \47746_nG1745d , \47743_nG1745b , \47745_nG1745c , \47178 );
buf \U$38677 ( \47747 , \47746_nG1745d );
_DC g19079_GF_IsGateDCbyConstraint ( \47748_nG19079 , \47747 , \42503 );
buf \U$38678 ( \47749 , \47748_nG19079 );
not \U$38679 ( \47750 , \47157 );
and \U$38680 ( \47751 , \47156 , \47750 );
_HMUX g1725c ( \47752_nG1725c , RIdc692d0_5752 , \47155 , \47751 );
_HMUX g1725d ( \47753_nG1725d , RIdc692d0_5752 , \47752_nG1725c , \47166 );
not \U$38681 ( \47754 , \47170 );
and \U$38682 ( \47755 , \47169 , \47754 );
_HMUX g1725f ( \47756_nG1725f , RIdc692d0_5752 , \47168 , \47755 );
_HMUX g17260 ( \47757_nG17260 , \47753_nG1725d , \47756_nG1725f , \47178 );
buf \U$38683 ( \47758 , \47757_nG17260 );
_DC g18f81_GF_IsGateDCbyConstraint ( \47759_nG18f81 , \47758 , \42503 );
buf \U$38684 ( \47760 , \47759_nG18f81 );
_HMUX g17261 ( \47761_nG17261 , RIdf7e930_5753 , \47183 , \47751 );
_HMUX g17262 ( \47762_nG17262 , RIdf7e930_5753 , \47761_nG17261 , \47166 );
_HMUX g17263 ( \47763_nG17263 , RIdf7e930_5753 , \47186 , \47755 );
_HMUX g17264 ( \47764_nG17264 , \47762_nG17262 , \47763_nG17263 , \47178 );
buf \U$38685 ( \47765 , \47764_nG17264 );
_DC g18f97_GF_IsGateDCbyConstraint ( \47766_nG18f97 , \47765 , \42503 );
buf \U$38686 ( \47767 , \47766_nG18f97 );
_HMUX g17265 ( \47768_nG17265 , RIdf8d6d8_5754 , \47192 , \47751 );
_HMUX g17266 ( \47769_nG17266 , RIdf8d6d8_5754 , \47768_nG17265 , \47166 );
_HMUX g17267 ( \47770_nG17267 , RIdf8d6d8_5754 , \47195 , \47755 );
_HMUX g17268 ( \47771_nG17268 , \47769_nG17266 , \47770_nG17267 , \47178 );
buf \U$38687 ( \47772 , \47771_nG17268 );
_DC g18fad_GF_IsGateDCbyConstraint ( \47773_nG18fad , \47772 , \42503 );
buf \U$38688 ( \47774 , \47773_nG18fad );
_HMUX g17269 ( \47775_nG17269 , RIdf9f978_5755 , \47201 , \47751 );
_HMUX g1726a ( \47776_nG1726a , RIdf9f978_5755 , \47775_nG17269 , \47166 );
_HMUX g1726b ( \47777_nG1726b , RIdf9f978_5755 , \47204 , \47755 );
_HMUX g1726c ( \47778_nG1726c , \47776_nG1726a , \47777_nG1726b , \47178 );
buf \U$38689 ( \47779 , \47778_nG1726c );
_DC g18fc3_GF_IsGateDCbyConstraint ( \47780_nG18fc3 , \47779 , \42503 );
buf \U$38690 ( \47781 , \47780_nG18fc3 );
_HMUX g1726d ( \47782_nG1726d , RIdfa6f20_5756 , \47210 , \47751 );
_HMUX g1726e ( \47783_nG1726e , RIdfa6f20_5756 , \47782_nG1726d , \47166 );
_HMUX g1726f ( \47784_nG1726f , RIdfa6f20_5756 , \47213 , \47755 );
_HMUX g17270 ( \47785_nG17270 , \47783_nG1726e , \47784_nG1726f , \47178 );
buf \U$38691 ( \47786 , \47785_nG17270 );
_DC g18fd9_GF_IsGateDCbyConstraint ( \47787_nG18fd9 , \47786 , \42503 );
buf \U$38692 ( \47788 , \47787_nG18fd9 );
_HMUX g17271 ( \47789_nG17271 , RIdfaf968_5757 , \47219 , \47751 );
_HMUX g17272 ( \47790_nG17272 , RIdfaf968_5757 , \47789_nG17271 , \47166 );
_HMUX g17273 ( \47791_nG17273 , RIdfaf968_5757 , \47222 , \47755 );
_HMUX g17274 ( \47792_nG17274 , \47790_nG17272 , \47791_nG17273 , \47178 );
buf \U$38693 ( \47793 , \47792_nG17274 );
_DC g18fef_GF_IsGateDCbyConstraint ( \47794_nG18fef , \47793 , \42503 );
buf \U$38694 ( \47795 , \47794_nG18fef );
_HMUX g17275 ( \47796_nG17275 , RIdfb74b0_5758 , \47228 , \47751 );
_HMUX g17276 ( \47797_nG17276 , RIdfb74b0_5758 , \47796_nG17275 , \47166 );
_HMUX g17277 ( \47798_nG17277 , RIdfb74b0_5758 , \47231 , \47755 );
_HMUX g17278 ( \47799_nG17278 , \47797_nG17276 , \47798_nG17277 , \47178 );
buf \U$38695 ( \47800 , \47799_nG17278 );
_DC g18ffb_GF_IsGateDCbyConstraint ( \47801_nG18ffb , \47800 , \42503 );
buf \U$38696 ( \47802 , \47801_nG18ffb );
_HMUX g17279 ( \47803_nG17279 , RIddf5a98_5759 , \47237 , \47751 );
_HMUX g1727a ( \47804_nG1727a , RIddf5a98_5759 , \47803_nG17279 , \47166 );
_HMUX g1727b ( \47805_nG1727b , RIddf5a98_5759 , \47240 , \47755 );
_HMUX g1727c ( \47806_nG1727c , \47804_nG1727a , \47805_nG1727b , \47178 );
buf \U$38697 ( \47807 , \47806_nG1727c );
_DC g18ffd_GF_IsGateDCbyConstraint ( \47808_nG18ffd , \47807 , \42503 );
buf \U$38698 ( \47809 , \47808_nG18ffd );
_HMUX g1727d ( \47810_nG1727d , RIde028d8_5760 , \47246 , \47751 );
_HMUX g1727e ( \47811_nG1727e , RIde028d8_5760 , \47810_nG1727d , \47166 );
_HMUX g1727f ( \47812_nG1727f , RIde028d8_5760 , \47249 , \47755 );
_HMUX g17280 ( \47813_nG17280 , \47811_nG1727e , \47812_nG1727f , \47178 );
buf \U$38699 ( \47814 , \47813_nG17280 );
_DC g18fff_GF_IsGateDCbyConstraint ( \47815_nG18fff , \47814 , \42503 );
buf \U$38700 ( \47816 , \47815_nG18fff );
_HMUX g17281 ( \47817_nG17281 , RIe036620_5761 , \47255 , \47751 );
_HMUX g17282 ( \47818_nG17282 , RIe036620_5761 , \47817_nG17281 , \47166 );
_HMUX g17283 ( \47819_nG17283 , RIe036620_5761 , \47258 , \47755 );
_HMUX g17284 ( \47820_nG17284 , \47818_nG17282 , \47819_nG17283 , \47178 );
buf \U$38701 ( \47821 , \47820_nG17284 );
_DC g18f83_GF_IsGateDCbyConstraint ( \47822_nG18f83 , \47821 , \42503 );
buf \U$38702 ( \47823 , \47822_nG18f83 );
_HMUX g17285 ( \47824_nG17285 , RIe027530_5762 , \47264 , \47751 );
_HMUX g17286 ( \47825_nG17286 , RIe027530_5762 , \47824_nG17285 , \47166 );
_HMUX g17287 ( \47826_nG17287 , RIe027530_5762 , \47267 , \47755 );
_HMUX g17288 ( \47827_nG17288 , \47825_nG17286 , \47826_nG17287 , \47178 );
buf \U$38703 ( \47828 , \47827_nG17288 );
_DC g18f85_GF_IsGateDCbyConstraint ( \47829_nG18f85 , \47828 , \42503 );
buf \U$38704 ( \47830 , \47829_nG18f85 );
_HMUX g17289 ( \47831_nG17289 , RIe01deb8_5763 , \47273 , \47751 );
_HMUX g1728a ( \47832_nG1728a , RIe01deb8_5763 , \47831_nG17289 , \47166 );
_HMUX g1728b ( \47833_nG1728b , RIe01deb8_5763 , \47276 , \47755 );
_HMUX g1728c ( \47834_nG1728c , \47832_nG1728a , \47833_nG1728b , \47178 );
buf \U$38705 ( \47835 , \47834_nG1728c );
_DC g18f87_GF_IsGateDCbyConstraint ( \47836_nG18f87 , \47835 , \42503 );
buf \U$38706 ( \47837 , \47836_nG18f87 );
_HMUX g1728d ( \47838_nG1728d , RIe00b3a8_5764 , \47282 , \47751 );
_HMUX g1728e ( \47839_nG1728e , RIe00b3a8_5764 , \47838_nG1728d , \47166 );
_HMUX g1728f ( \47840_nG1728f , RIe00b3a8_5764 , \47285 , \47755 );
_HMUX g17290 ( \47841_nG17290 , \47839_nG1728e , \47840_nG1728f , \47178 );
buf \U$38707 ( \47842 , \47841_nG17290 );
_DC g18f89_GF_IsGateDCbyConstraint ( \47843_nG18f89 , \47842 , \42503 );
buf \U$38708 ( \47844 , \47843_nG18f89 );
_HMUX g17291 ( \47845_nG17291 , RIdffd938_5765 , \47291 , \47751 );
_HMUX g17292 ( \47846_nG17292 , RIdffd938_5765 , \47845_nG17291 , \47166 );
_HMUX g17293 ( \47847_nG17293 , RIdffd938_5765 , \47294 , \47755 );
_HMUX g17294 ( \47848_nG17294 , \47846_nG17292 , \47847_nG17293 , \47178 );
buf \U$38709 ( \47849 , \47848_nG17294 );
_DC g18f8b_GF_IsGateDCbyConstraint ( \47850_nG18f8b , \47849 , \42503 );
buf \U$38710 ( \47851 , \47850_nG18f8b );
_HMUX g17295 ( \47852_nG17295 , RIdfefb08_5766 , \47300 , \47751 );
_HMUX g17296 ( \47853_nG17296 , RIdfefb08_5766 , \47852_nG17295 , \47166 );
_HMUX g17297 ( \47854_nG17297 , RIdfefb08_5766 , \47303 , \47755 );
_HMUX g17298 ( \47855_nG17298 , \47853_nG17296 , \47854_nG17297 , \47178 );
buf \U$38711 ( \47856 , \47855_nG17298 );
_DC g18f8d_GF_IsGateDCbyConstraint ( \47857_nG18f8d , \47856 , \42503 );
buf \U$38712 ( \47858 , \47857_nG18f8d );
_HMUX g17299 ( \47859_nG17299 , RIdfe0838_5767 , \47309 , \47751 );
_HMUX g1729a ( \47860_nG1729a , RIdfe0838_5767 , \47859_nG17299 , \47166 );
_HMUX g1729b ( \47861_nG1729b , RIdfe0838_5767 , \47312 , \47755 );
_HMUX g1729c ( \47862_nG1729c , \47860_nG1729a , \47861_nG1729b , \47178 );
buf \U$38713 ( \47863 , \47862_nG1729c );
_DC g18f8f_GF_IsGateDCbyConstraint ( \47864_nG18f8f , \47863 , \42503 );
buf \U$38714 ( \47865 , \47864_nG18f8f );
_HMUX g1729d ( \47866_nG1729d , RIdfd6680_5768 , \47318 , \47751 );
_HMUX g1729e ( \47867_nG1729e , RIdfd6680_5768 , \47866_nG1729d , \47166 );
_HMUX g1729f ( \47868_nG1729f , RIdfd6680_5768 , \47321 , \47755 );
_HMUX g172a0 ( \47869_nG172a0 , \47867_nG1729e , \47868_nG1729f , \47178 );
buf \U$38715 ( \47870 , \47869_nG172a0 );
_DC g18f91_GF_IsGateDCbyConstraint ( \47871_nG18f91 , \47870 , \42503 );
buf \U$38716 ( \47872 , \47871_nG18f91 );
_HMUX g172a1 ( \47873_nG172a1 , RIe1084d0_5769 , \47327 , \47751 );
_HMUX g172a2 ( \47874_nG172a2 , RIe1084d0_5769 , \47873_nG172a1 , \47166 );
_HMUX g172a3 ( \47875_nG172a3 , RIe1084d0_5769 , \47330 , \47755 );
_HMUX g172a4 ( \47876_nG172a4 , \47874_nG172a2 , \47875_nG172a3 , \47178 );
buf \U$38717 ( \47877 , \47876_nG172a4 );
_DC g18f93_GF_IsGateDCbyConstraint ( \47878_nG18f93 , \47877 , \42503 );
buf \U$38718 ( \47879 , \47878_nG18f93 );
_HMUX g172a5 ( \47880_nG172a5 , RIe10ad98_5770 , \47336 , \47751 );
_HMUX g172a6 ( \47881_nG172a6 , RIe10ad98_5770 , \47880_nG172a5 , \47166 );
_HMUX g172a7 ( \47882_nG172a7 , RIe10ad98_5770 , \47339 , \47755 );
_HMUX g172a8 ( \47883_nG172a8 , \47881_nG172a6 , \47882_nG172a7 , \47178 );
buf \U$38719 ( \47884 , \47883_nG172a8 );
_DC g18f95_GF_IsGateDCbyConstraint ( \47885_nG18f95 , \47884 , \42503 );
buf \U$38720 ( \47886 , \47885_nG18f95 );
_HMUX g172a9 ( \47887_nG172a9 , RIe10e470_5771 , \47345 , \47751 );
_HMUX g172aa ( \47888_nG172aa , RIe10e470_5771 , \47887_nG172a9 , \47166 );
_HMUX g172ab ( \47889_nG172ab , RIe10e470_5771 , \47348 , \47755 );
_HMUX g172ac ( \47890_nG172ac , \47888_nG172aa , \47889_nG172ab , \47178 );
buf \U$38721 ( \47891 , \47890_nG172ac );
_DC g18f99_GF_IsGateDCbyConstraint ( \47892_nG18f99 , \47891 , \42503 );
buf \U$38722 ( \47893 , \47892_nG18f99 );
_HMUX g172ad ( \47894_nG172ad , RIe110d38_5772 , \47354 , \47751 );
_HMUX g172ae ( \47895_nG172ae , RIe110d38_5772 , \47894_nG172ad , \47166 );
_HMUX g172af ( \47896_nG172af , RIe110d38_5772 , \47357 , \47755 );
_HMUX g172b0 ( \47897_nG172b0 , \47895_nG172ae , \47896_nG172af , \47178 );
buf \U$38723 ( \47898 , \47897_nG172b0 );
_DC g18f9b_GF_IsGateDCbyConstraint ( \47899_nG18f9b , \47898 , \42503 );
buf \U$38724 ( \47900 , \47899_nG18f9b );
_HMUX g172b1 ( \47901_nG172b1 , RIe113ab0_5773 , \47363 , \47751 );
_HMUX g172b2 ( \47902_nG172b2 , RIe113ab0_5773 , \47901_nG172b1 , \47166 );
_HMUX g172b3 ( \47903_nG172b3 , RIe113ab0_5773 , \47366 , \47755 );
_HMUX g172b4 ( \47904_nG172b4 , \47902_nG172b2 , \47903_nG172b3 , \47178 );
buf \U$38725 ( \47905 , \47904_nG172b4 );
_DC g18f9d_GF_IsGateDCbyConstraint ( \47906_nG18f9d , \47905 , \42503 );
buf \U$38726 ( \47907 , \47906_nG18f9d );
_HMUX g172b5 ( \47908_nG172b5 , RIe116cd8_5774 , \47372 , \47751 );
_HMUX g172b6 ( \47909_nG172b6 , RIe116cd8_5774 , \47908_nG172b5 , \47166 );
_HMUX g172b7 ( \47910_nG172b7 , RIe116cd8_5774 , \47375 , \47755 );
_HMUX g172b8 ( \47911_nG172b8 , \47909_nG172b6 , \47910_nG172b7 , \47178 );
buf \U$38727 ( \47912 , \47911_nG172b8 );
_DC g18f9f_GF_IsGateDCbyConstraint ( \47913_nG18f9f , \47912 , \42503 );
buf \U$38728 ( \47914 , \47913_nG18f9f );
_HMUX g172b9 ( \47915_nG172b9 , RIe119a50_5775 , \47381 , \47751 );
_HMUX g172ba ( \47916_nG172ba , RIe119a50_5775 , \47915_nG172b9 , \47166 );
_HMUX g172bb ( \47917_nG172bb , RIe119a50_5775 , \47384 , \47755 );
_HMUX g172bc ( \47918_nG172bc , \47916_nG172ba , \47917_nG172bb , \47178 );
buf \U$38729 ( \47919 , \47918_nG172bc );
_DC g18fa1_GF_IsGateDCbyConstraint ( \47920_nG18fa1 , \47919 , \42503 );
buf \U$38730 ( \47921 , \47920_nG18fa1 );
_HMUX g172bd ( \47922_nG172bd , RIe11cc78_5776 , \47390 , \47751 );
_HMUX g172be ( \47923_nG172be , RIe11cc78_5776 , \47922_nG172bd , \47166 );
_HMUX g172bf ( \47924_nG172bf , RIe11cc78_5776 , \47393 , \47755 );
_HMUX g172c0 ( \47925_nG172c0 , \47923_nG172be , \47924_nG172bf , \47178 );
buf \U$38731 ( \47926 , \47925_nG172c0 );
_DC g18fa3_GF_IsGateDCbyConstraint ( \47927_nG18fa3 , \47926 , \42503 );
buf \U$38732 ( \47928 , \47927_nG18fa3 );
_HMUX g172c1 ( \47929_nG172c1 , RIe11f9f0_5777 , \47399 , \47751 );
_HMUX g172c2 ( \47930_nG172c2 , RIe11f9f0_5777 , \47929_nG172c1 , \47166 );
_HMUX g172c3 ( \47931_nG172c3 , RIe11f9f0_5777 , \47402 , \47755 );
_HMUX g172c4 ( \47932_nG172c4 , \47930_nG172c2 , \47931_nG172c3 , \47178 );
buf \U$38733 ( \47933 , \47932_nG172c4 );
_DC g18fa5_GF_IsGateDCbyConstraint ( \47934_nG18fa5 , \47933 , \42503 );
buf \U$38734 ( \47935 , \47934_nG18fa5 );
_HMUX g172c5 ( \47936_nG172c5 , RIe122c18_5778 , \47408 , \47751 );
_HMUX g172c6 ( \47937_nG172c6 , RIe122c18_5778 , \47936_nG172c5 , \47166 );
_HMUX g172c7 ( \47938_nG172c7 , RIe122c18_5778 , \47411 , \47755 );
_HMUX g172c8 ( \47939_nG172c8 , \47937_nG172c6 , \47938_nG172c7 , \47178 );
buf \U$38735 ( \47940 , \47939_nG172c8 );
_DC g18fa7_GF_IsGateDCbyConstraint ( \47941_nG18fa7 , \47940 , \42503 );
buf \U$38736 ( \47942 , \47941_nG18fa7 );
_HMUX g172c9 ( \47943_nG172c9 , RIe125990_5779 , \47417 , \47751 );
_HMUX g172ca ( \47944_nG172ca , RIe125990_5779 , \47943_nG172c9 , \47166 );
_HMUX g172cb ( \47945_nG172cb , RIe125990_5779 , \47420 , \47755 );
_HMUX g172cc ( \47946_nG172cc , \47944_nG172ca , \47945_nG172cb , \47178 );
buf \U$38737 ( \47947 , \47946_nG172cc );
_DC g18fa9_GF_IsGateDCbyConstraint ( \47948_nG18fa9 , \47947 , \42503 );
buf \U$38738 ( \47949 , \47948_nG18fa9 );
_HMUX g172cd ( \47950_nG172cd , RIe128258_5780 , \47426 , \47751 );
_HMUX g172ce ( \47951_nG172ce , RIe128258_5780 , \47950_nG172cd , \47166 );
_HMUX g172cf ( \47952_nG172cf , RIe128258_5780 , \47429 , \47755 );
_HMUX g172d0 ( \47953_nG172d0 , \47951_nG172ce , \47952_nG172cf , \47178 );
buf \U$38739 ( \47954 , \47953_nG172d0 );
_DC g18fab_GF_IsGateDCbyConstraint ( \47955_nG18fab , \47954 , \42503 );
buf \U$38740 ( \47956 , \47955_nG18fab );
_HMUX g172d1 ( \47957_nG172d1 , RIe12b930_5781 , \47435 , \47751 );
_HMUX g172d2 ( \47958_nG172d2 , RIe12b930_5781 , \47957_nG172d1 , \47166 );
_HMUX g172d3 ( \47959_nG172d3 , RIe12b930_5781 , \47438 , \47755 );
_HMUX g172d4 ( \47960_nG172d4 , \47958_nG172d2 , \47959_nG172d3 , \47178 );
buf \U$38741 ( \47961 , \47960_nG172d4 );
_DC g18faf_GF_IsGateDCbyConstraint ( \47962_nG18faf , \47961 , \42503 );
buf \U$38742 ( \47963 , \47962_nG18faf );
_HMUX g172d5 ( \47964_nG172d5 , RIe12e1f8_5782 , \47444 , \47751 );
_HMUX g172d6 ( \47965_nG172d6 , RIe12e1f8_5782 , \47964_nG172d5 , \47166 );
_HMUX g172d7 ( \47966_nG172d7 , RIe12e1f8_5782 , \47447 , \47755 );
_HMUX g172d8 ( \47967_nG172d8 , \47965_nG172d6 , \47966_nG172d7 , \47178 );
buf \U$38743 ( \47968 , \47967_nG172d8 );
_DC g18fb1_GF_IsGateDCbyConstraint ( \47969_nG18fb1 , \47968 , \42503 );
buf \U$38744 ( \47970 , \47969_nG18fb1 );
_HMUX g172d9 ( \47971_nG172d9 , RIe1308e0_5783 , \47453 , \47751 );
_HMUX g172da ( \47972_nG172da , RIe1308e0_5783 , \47971_nG172d9 , \47166 );
_HMUX g172db ( \47973_nG172db , RIe1308e0_5783 , \47456 , \47755 );
_HMUX g172dc ( \47974_nG172dc , \47972_nG172da , \47973_nG172db , \47178 );
buf \U$38745 ( \47975 , \47974_nG172dc );
_DC g18fb3_GF_IsGateDCbyConstraint ( \47976_nG18fb3 , \47975 , \42503 );
buf \U$38746 ( \47977 , \47976_nG18fb3 );
_HMUX g172dd ( \47978_nG172dd , RIe132398_5784 , \47462 , \47751 );
_HMUX g172de ( \47979_nG172de , RIe132398_5784 , \47978_nG172dd , \47166 );
_HMUX g172df ( \47980_nG172df , RIe132398_5784 , \47465 , \47755 );
_HMUX g172e0 ( \47981_nG172e0 , \47979_nG172de , \47980_nG172df , \47178 );
buf \U$38747 ( \47982 , \47981_nG172e0 );
_DC g18fb5_GF_IsGateDCbyConstraint ( \47983_nG18fb5 , \47982 , \42503 );
buf \U$38748 ( \47984 , \47983_nG18fb5 );
_HMUX g172e1 ( \47985_nG172e1 , RIe134300_5785 , \47471 , \47751 );
_HMUX g172e2 ( \47986_nG172e2 , RIe134300_5785 , \47985_nG172e1 , \47166 );
_HMUX g172e3 ( \47987_nG172e3 , RIe134300_5785 , \47474 , \47755 );
_HMUX g172e4 ( \47988_nG172e4 , \47986_nG172e2 , \47987_nG172e3 , \47178 );
buf \U$38749 ( \47989 , \47988_nG172e4 );
_DC g18fb7_GF_IsGateDCbyConstraint ( \47990_nG18fb7 , \47989 , \42503 );
buf \U$38750 ( \47991 , \47990_nG18fb7 );
_HMUX g172e5 ( \47992_nG172e5 , RIe135ae8_5786 , \47480 , \47751 );
_HMUX g172e6 ( \47993_nG172e6 , RIe135ae8_5786 , \47992_nG172e5 , \47166 );
_HMUX g172e7 ( \47994_nG172e7 , RIe135ae8_5786 , \47483 , \47755 );
_HMUX g172e8 ( \47995_nG172e8 , \47993_nG172e6 , \47994_nG172e7 , \47178 );
buf \U$38751 ( \47996 , \47995_nG172e8 );
_DC g18fb9_GF_IsGateDCbyConstraint ( \47997_nG18fb9 , \47996 , \42503 );
buf \U$38752 ( \47998 , \47997_nG18fb9 );
_HMUX g172e9 ( \47999_nG172e9 , RIe137258_5787 , \47489 , \47751 );
_HMUX g172ea ( \48000_nG172ea , RIe137258_5787 , \47999_nG172e9 , \47166 );
_HMUX g172eb ( \48001_nG172eb , RIe137258_5787 , \47492 , \47755 );
_HMUX g172ec ( \48002_nG172ec , \48000_nG172ea , \48001_nG172eb , \47178 );
buf \U$38753 ( \48003 , \48002_nG172ec );
_DC g18fbb_GF_IsGateDCbyConstraint ( \48004_nG18fbb , \48003 , \42503 );
buf \U$38754 ( \48005 , \48004_nG18fbb );
_HMUX g172ed ( \48006_nG172ed , RIe138608_5788 , \47498 , \47751 );
_HMUX g172ee ( \48007_nG172ee , RIe138608_5788 , \48006_nG172ed , \47166 );
_HMUX g172ef ( \48008_nG172ef , RIe138608_5788 , \47501 , \47755 );
_HMUX g172f0 ( \48009_nG172f0 , \48007_nG172ee , \48008_nG172ef , \47178 );
buf \U$38755 ( \48010 , \48009_nG172f0 );
_DC g18fbd_GF_IsGateDCbyConstraint ( \48011_nG18fbd , \48010 , \42503 );
buf \U$38756 ( \48012 , \48011_nG18fbd );
_HMUX g172f1 ( \48013_nG172f1 , RIe139850_5789 , \47507 , \47751 );
_HMUX g172f2 ( \48014_nG172f2 , RIe139850_5789 , \48013_nG172f1 , \47166 );
_HMUX g172f3 ( \48015_nG172f3 , RIe139850_5789 , \47510 , \47755 );
_HMUX g172f4 ( \48016_nG172f4 , \48014_nG172f2 , \48015_nG172f3 , \47178 );
buf \U$38757 ( \48017 , \48016_nG172f4 );
_DC g18fbf_GF_IsGateDCbyConstraint ( \48018_nG18fbf , \48017 , \42503 );
buf \U$38758 ( \48019 , \48018_nG18fbf );
_HMUX g172f5 ( \48020_nG172f5 , RIe13ab88_5790 , \47516 , \47751 );
_HMUX g172f6 ( \48021_nG172f6 , RIe13ab88_5790 , \48020_nG172f5 , \47166 );
_HMUX g172f7 ( \48022_nG172f7 , RIe13ab88_5790 , \47519 , \47755 );
_HMUX g172f8 ( \48023_nG172f8 , \48021_nG172f6 , \48022_nG172f7 , \47178 );
buf \U$38759 ( \48024 , \48023_nG172f8 );
_DC g18fc1_GF_IsGateDCbyConstraint ( \48025_nG18fc1 , \48024 , \42503 );
buf \U$38760 ( \48026 , \48025_nG18fc1 );
_HMUX g172f9 ( \48027_nG172f9 , RIe13c028_5791 , \47525 , \47751 );
_HMUX g172fa ( \48028_nG172fa , RIe13c028_5791 , \48027_nG172f9 , \47166 );
_HMUX g172fb ( \48029_nG172fb , RIe13c028_5791 , \47528 , \47755 );
_HMUX g172fc ( \48030_nG172fc , \48028_nG172fa , \48029_nG172fb , \47178 );
buf \U$38761 ( \48031 , \48030_nG172fc );
_DC g18fc5_GF_IsGateDCbyConstraint ( \48032_nG18fc5 , \48031 , \42503 );
buf \U$38762 ( \48033 , \48032_nG18fc5 );
_HMUX g172fd ( \48034_nG172fd , RIe13d5b8_5792 , \47534 , \47751 );
_HMUX g172fe ( \48035_nG172fe , RIe13d5b8_5792 , \48034_nG172fd , \47166 );
_HMUX g172ff ( \48036_nG172ff , RIe13d5b8_5792 , \47537 , \47755 );
_HMUX g17300 ( \48037_nG17300 , \48035_nG172fe , \48036_nG172ff , \47178 );
buf \U$38763 ( \48038 , \48037_nG17300 );
_DC g18fc7_GF_IsGateDCbyConstraint ( \48039_nG18fc7 , \48038 , \42503 );
buf \U$38764 ( \48040 , \48039_nG18fc7 );
_HMUX g17301 ( \48041_nG17301 , RIe13ead0_5793 , \47543 , \47751 );
_HMUX g17302 ( \48042_nG17302 , RIe13ead0_5793 , \48041_nG17301 , \47166 );
_HMUX g17303 ( \48043_nG17303 , RIe13ead0_5793 , \47546 , \47755 );
_HMUX g17304 ( \48044_nG17304 , \48042_nG17302 , \48043_nG17303 , \47178 );
buf \U$38765 ( \48045 , \48044_nG17304 );
_DC g18fc9_GF_IsGateDCbyConstraint ( \48046_nG18fc9 , \48045 , \42503 );
buf \U$38766 ( \48047 , \48046_nG18fc9 );
_HMUX g17305 ( \48048_nG17305 , RIe13fef8_5794 , \47552 , \47751 );
_HMUX g17306 ( \48049_nG17306 , RIe13fef8_5794 , \48048_nG17305 , \47166 );
_HMUX g17307 ( \48050_nG17307 , RIe13fef8_5794 , \47555 , \47755 );
_HMUX g17308 ( \48051_nG17308 , \48049_nG17306 , \48050_nG17307 , \47178 );
buf \U$38767 ( \48052 , \48051_nG17308 );
_DC g18fcb_GF_IsGateDCbyConstraint ( \48053_nG18fcb , \48052 , \42503 );
buf \U$38768 ( \48054 , \48053_nG18fcb );
_HMUX g17309 ( \48055_nG17309 , RIe141230_5795 , \47561 , \47751 );
_HMUX g1730a ( \48056_nG1730a , RIe141230_5795 , \48055_nG17309 , \47166 );
_HMUX g1730b ( \48057_nG1730b , RIe141230_5795 , \47564 , \47755 );
_HMUX g1730c ( \48058_nG1730c , \48056_nG1730a , \48057_nG1730b , \47178 );
buf \U$38769 ( \48059 , \48058_nG1730c );
_DC g18fcd_GF_IsGateDCbyConstraint ( \48060_nG18fcd , \48059 , \42503 );
buf \U$38770 ( \48061 , \48060_nG18fcd );
_HMUX g1730d ( \48062_nG1730d , RIe142568_5796 , \47570 , \47751 );
_HMUX g1730e ( \48063_nG1730e , RIe142568_5796 , \48062_nG1730d , \47166 );
_HMUX g1730f ( \48064_nG1730f , RIe142568_5796 , \47573 , \47755 );
_HMUX g17310 ( \48065_nG17310 , \48063_nG1730e , \48064_nG1730f , \47178 );
buf \U$38771 ( \48066 , \48065_nG17310 );
_DC g18fcf_GF_IsGateDCbyConstraint ( \48067_nG18fcf , \48066 , \42503 );
buf \U$38772 ( \48068 , \48067_nG18fcf );
_HMUX g17311 ( \48069_nG17311 , RIe1434e0_5797 , \47579 , \47751 );
_HMUX g17312 ( \48070_nG17312 , RIe1434e0_5797 , \48069_nG17311 , \47166 );
_HMUX g17313 ( \48071_nG17313 , RIe1434e0_5797 , \47582 , \47755 );
_HMUX g17314 ( \48072_nG17314 , \48070_nG17312 , \48071_nG17313 , \47178 );
buf \U$38773 ( \48073 , \48072_nG17314 );
_DC g18fd1_GF_IsGateDCbyConstraint ( \48074_nG18fd1 , \48073 , \42503 );
buf \U$38774 ( \48075 , \48074_nG18fd1 );
_HMUX g17315 ( \48076_nG17315 , RIe144638_5798 , \47588 , \47751 );
_HMUX g17316 ( \48077_nG17316 , RIe144638_5798 , \48076_nG17315 , \47166 );
_HMUX g17317 ( \48078_nG17317 , RIe144638_5798 , \47591 , \47755 );
_HMUX g17318 ( \48079_nG17318 , \48077_nG17316 , \48078_nG17317 , \47178 );
buf \U$38775 ( \48080 , \48079_nG17318 );
_DC g18fd3_GF_IsGateDCbyConstraint ( \48081_nG18fd3 , \48080 , \42503 );
buf \U$38776 ( \48082 , \48081_nG18fd3 );
_HMUX g17319 ( \48083_nG17319 , RIe145880_5799 , \47597 , \47751 );
_HMUX g1731a ( \48084_nG1731a , RIe145880_5799 , \48083_nG17319 , \47166 );
_HMUX g1731b ( \48085_nG1731b , RIe145880_5799 , \47600 , \47755 );
_HMUX g1731c ( \48086_nG1731c , \48084_nG1731a , \48085_nG1731b , \47178 );
buf \U$38777 ( \48087 , \48086_nG1731c );
_DC g18fd5_GF_IsGateDCbyConstraint ( \48088_nG18fd5 , \48087 , \42503 );
buf \U$38778 ( \48089 , \48088_nG18fd5 );
_HMUX g1731d ( \48090_nG1731d , RIe146ac8_5800 , \47606 , \47751 );
_HMUX g1731e ( \48091_nG1731e , RIe146ac8_5800 , \48090_nG1731d , \47166 );
_HMUX g1731f ( \48092_nG1731f , RIe146ac8_5800 , \47609 , \47755 );
_HMUX g17320 ( \48093_nG17320 , \48091_nG1731e , \48092_nG1731f , \47178 );
buf \U$38779 ( \48094 , \48093_nG17320 );
_DC g18fd7_GF_IsGateDCbyConstraint ( \48095_nG18fd7 , \48094 , \42503 );
buf \U$38780 ( \48096 , \48095_nG18fd7 );
_HMUX g17321 ( \48097_nG17321 , RIe1486e8_5801 , \47615 , \47751 );
_HMUX g17322 ( \48098_nG17322 , RIe1486e8_5801 , \48097_nG17321 , \47166 );
_HMUX g17323 ( \48099_nG17323 , RIe1486e8_5801 , \47618 , \47755 );
_HMUX g17324 ( \48100_nG17324 , \48098_nG17322 , \48099_nG17323 , \47178 );
buf \U$38781 ( \48101 , \48100_nG17324 );
_DC g18fdb_GF_IsGateDCbyConstraint ( \48102_nG18fdb , \48101 , \42503 );
buf \U$38782 ( \48103 , \48102_nG18fdb );
_HMUX g17325 ( \48104_nG17325 , RIe149f48_5802 , \47624 , \47751 );
_HMUX g17326 ( \48105_nG17326 , RIe149f48_5802 , \48104_nG17325 , \47166 );
_HMUX g17327 ( \48106_nG17327 , RIe149f48_5802 , \47627 , \47755 );
_HMUX g17328 ( \48107_nG17328 , \48105_nG17326 , \48106_nG17327 , \47178 );
buf \U$38783 ( \48108 , \48107_nG17328 );
_DC g18fdd_GF_IsGateDCbyConstraint ( \48109_nG18fdd , \48108 , \42503 );
buf \U$38784 ( \48110 , \48109_nG18fdd );
_HMUX g17329 ( \48111_nG17329 , RIe14b550_5803 , \47633 , \47751 );
_HMUX g1732a ( \48112_nG1732a , RIe14b550_5803 , \48111_nG17329 , \47166 );
_HMUX g1732b ( \48113_nG1732b , RIe14b550_5803 , \47636 , \47755 );
_HMUX g1732c ( \48114_nG1732c , \48112_nG1732a , \48113_nG1732b , \47178 );
buf \U$38785 ( \48115 , \48114_nG1732c );
_DC g18fdf_GF_IsGateDCbyConstraint ( \48116_nG18fdf , \48115 , \42503 );
buf \U$38786 ( \48117 , \48116_nG18fdf );
_HMUX g1732d ( \48118_nG1732d , RIe14c978_5804 , \47642 , \47751 );
_HMUX g1732e ( \48119_nG1732e , RIe14c978_5804 , \48118_nG1732d , \47166 );
_HMUX g1732f ( \48120_nG1732f , RIe14c978_5804 , \47645 , \47755 );
_HMUX g17330 ( \48121_nG17330 , \48119_nG1732e , \48120_nG1732f , \47178 );
buf \U$38787 ( \48122 , \48121_nG17330 );
_DC g18fe1_GF_IsGateDCbyConstraint ( \48123_nG18fe1 , \48122 , \42503 );
buf \U$38788 ( \48124 , \48123_nG18fe1 );
_HMUX g17331 ( \48125_nG17331 , RIe14e430_5805 , \47651 , \47751 );
_HMUX g17332 ( \48126_nG17332 , RIe14e430_5805 , \48125_nG17331 , \47166 );
_HMUX g17333 ( \48127_nG17333 , RIe14e430_5805 , \47654 , \47755 );
_HMUX g17334 ( \48128_nG17334 , \48126_nG17332 , \48127_nG17333 , \47178 );
buf \U$38789 ( \48129 , \48128_nG17334 );
_DC g18fe3_GF_IsGateDCbyConstraint ( \48130_nG18fe3 , \48129 , \42503 );
buf \U$38790 ( \48131 , \48130_nG18fe3 );
_HMUX g17335 ( \48132_nG17335 , RIe0865e8_5806 , \47660 , \47751 );
_HMUX g17336 ( \48133_nG17336 , RIe0865e8_5806 , \48132_nG17335 , \47166 );
_HMUX g17337 ( \48134_nG17337 , RIe0865e8_5806 , \47663 , \47755 );
_HMUX g17338 ( \48135_nG17338 , \48133_nG17336 , \48134_nG17337 , \47178 );
buf \U$38791 ( \48136 , \48135_nG17338 );
_DC g18fe5_GF_IsGateDCbyConstraint ( \48137_nG18fe5 , \48136 , \42503 );
buf \U$38792 ( \48138 , \48137_nG18fe5 );
_HMUX g17339 ( \48139_nG17339 , RIe087f38_5807 , \47669 , \47751 );
_HMUX g1733a ( \48140_nG1733a , RIe087f38_5807 , \48139_nG17339 , \47166 );
_HMUX g1733b ( \48141_nG1733b , RIe087f38_5807 , \47672 , \47755 );
_HMUX g1733c ( \48142_nG1733c , \48140_nG1733a , \48141_nG1733b , \47178 );
buf \U$38793 ( \48143 , \48142_nG1733c );
_DC g18fe7_GF_IsGateDCbyConstraint ( \48144_nG18fe7 , \48143 , \42503 );
buf \U$38794 ( \48145 , \48144_nG18fe7 );
_HMUX g1733d ( \48146_nG1733d , RIe089db0_5808 , \47678 , \47751 );
_HMUX g1733e ( \48147_nG1733e , RIe089db0_5808 , \48146_nG1733d , \47166 );
_HMUX g1733f ( \48148_nG1733f , RIe089db0_5808 , \47681 , \47755 );
_HMUX g17340 ( \48149_nG17340 , \48147_nG1733e , \48148_nG1733f , \47178 );
buf \U$38795 ( \48150 , \48149_nG17340 );
_DC g18fe9_GF_IsGateDCbyConstraint ( \48151_nG18fe9 , \48150 , \42503 );
buf \U$38796 ( \48152 , \48151_nG18fe9 );
_HMUX g17341 ( \48153_nG17341 , RIe08b7f0_5809 , \47687 , \47751 );
_HMUX g17342 ( \48154_nG17342 , RIe08b7f0_5809 , \48153_nG17341 , \47166 );
_HMUX g17343 ( \48155_nG17343 , RIe08b7f0_5809 , \47690 , \47755 );
_HMUX g17344 ( \48156_nG17344 , \48154_nG17342 , \48155_nG17343 , \47178 );
buf \U$38797 ( \48157 , \48156_nG17344 );
_DC g18feb_GF_IsGateDCbyConstraint ( \48158_nG18feb , \48157 , \42503 );
buf \U$38798 ( \48159 , \48158_nG18feb );
_HMUX g17345 ( \48160_nG17345 , RIe08d578_5810 , \47696 , \47751 );
_HMUX g17346 ( \48161_nG17346 , RIe08d578_5810 , \48160_nG17345 , \47166 );
_HMUX g17347 ( \48162_nG17347 , RIe08d578_5810 , \47699 , \47755 );
_HMUX g17348 ( \48163_nG17348 , \48161_nG17346 , \48162_nG17347 , \47178 );
buf \U$38799 ( \48164 , \48163_nG17348 );
_DC g18fed_GF_IsGateDCbyConstraint ( \48165_nG18fed , \48164 , \42503 );
buf \U$38800 ( \48166 , \48165_nG18fed );
_HMUX g17349 ( \48167_nG17349 , RIe08f120_5811 , \47705 , \47751 );
_HMUX g1734a ( \48168_nG1734a , RIe08f120_5811 , \48167_nG17349 , \47166 );
_HMUX g1734b ( \48169_nG1734b , RIe08f120_5811 , \47708 , \47755 );
_HMUX g1734c ( \48170_nG1734c , \48168_nG1734a , \48169_nG1734b , \47178 );
buf \U$38801 ( \48171 , \48170_nG1734c );
_DC g18ff1_GF_IsGateDCbyConstraint ( \48172_nG18ff1 , \48171 , \42503 );
buf \U$38802 ( \48173 , \48172_nG18ff1 );
_HMUX g1734d ( \48174_nG1734d , RIe091100_5812 , \47714 , \47751 );
_HMUX g1734e ( \48175_nG1734e , RIe091100_5812 , \48174_nG1734d , \47166 );
_HMUX g1734f ( \48176_nG1734f , RIe091100_5812 , \47717 , \47755 );
_HMUX g17350 ( \48177_nG17350 , \48175_nG1734e , \48176_nG1734f , \47178 );
buf \U$38803 ( \48178 , \48177_nG17350 );
_DC g18ff3_GF_IsGateDCbyConstraint ( \48179_nG18ff3 , \48178 , \42503 );
buf \U$38804 ( \48180 , \48179_nG18ff3 );
_HMUX g17351 ( \48181_nG17351 , RIe093248_5813 , \47723 , \47751 );
_HMUX g17352 ( \48182_nG17352 , RIe093248_5813 , \48181_nG17351 , \47166 );
_HMUX g17353 ( \48183_nG17353 , RIe093248_5813 , \47726 , \47755 );
_HMUX g17354 ( \48184_nG17354 , \48182_nG17352 , \48183_nG17353 , \47178 );
buf \U$38805 ( \48185 , \48184_nG17354 );
_DC g18ff5_GF_IsGateDCbyConstraint ( \48186_nG18ff5 , \48185 , \42503 );
buf \U$38806 ( \48187 , \48186_nG18ff5 );
_HMUX g17355 ( \48188_nG17355 , RIe0950c0_5814 , \47732 , \47751 );
_HMUX g17356 ( \48189_nG17356 , RIe0950c0_5814 , \48188_nG17355 , \47166 );
_HMUX g17357 ( \48190_nG17357 , RIe0950c0_5814 , \47735 , \47755 );
_HMUX g17358 ( \48191_nG17358 , \48189_nG17356 , \48190_nG17357 , \47178 );
buf \U$38807 ( \48192 , \48191_nG17358 );
_DC g18ff7_GF_IsGateDCbyConstraint ( \48193_nG18ff7 , \48192 , \42503 );
buf \U$38808 ( \48194 , \48193_nG18ff7 );
_HMUX g17359 ( \48195_nG17359 , RIe096998_5815 , \47741 , \47751 );
_HMUX g1735a ( \48196_nG1735a , RIe096998_5815 , \48195_nG17359 , \47166 );
_HMUX g1735b ( \48197_nG1735b , RIe096998_5815 , \47744 , \47755 );
_HMUX g1735c ( \48198_nG1735c , \48196_nG1735a , \48197_nG1735b , \47178 );
buf \U$38809 ( \48199 , \48198_nG1735c );
_DC g18ff9_GF_IsGateDCbyConstraint ( \48200_nG18ff9 , \48199 , \42503 );
buf \U$38810 ( \48201 , \48200_nG18ff9 );
nor \U$38811 ( \48202 , \47156 , \47750 );
_HMUX g1715a ( \48203_nG1715a , RIe0986a8_5816 , \47155 , \48202 );
_HMUX g1715b ( \48204_nG1715b , RIe0986a8_5816 , \48203_nG1715a , \47166 );
nor \U$38812 ( \48205 , \47169 , \47754 );
_HMUX g1715e ( \48206_nG1715e , RIe0986a8_5816 , \47168 , \48205 );
_HMUX g1715f ( \48207_nG1715f , \48204_nG1715b , \48206_nG1715e , \47178 );
buf \U$38813 ( \48208 , \48207_nG1715f );
_DC g18f01_GF_IsGateDCbyConstraint ( \48209_nG18f01 , \48208 , \42503 );
buf \U$38814 ( \48210 , \48209_nG18f01 );
_HMUX g17160 ( \48211_nG17160 , RIe1cfd18_5817 , \47183 , \48202 );
_HMUX g17161 ( \48212_nG17161 , RIe1cfd18_5817 , \48211_nG17160 , \47166 );
_HMUX g17162 ( \48213_nG17162 , RIe1cfd18_5817 , \47186 , \48205 );
_HMUX g17163 ( \48214_nG17163 , \48212_nG17161 , \48213_nG17162 , \47178 );
buf \U$38815 ( \48215 , \48214_nG17163 );
_DC g18f17_GF_IsGateDCbyConstraint ( \48216_nG18f17 , \48215 , \42503 );
buf \U$38816 ( \48217 , \48216_nG18f17 );
_HMUX g17164 ( \48218_nG17164 , RIe1ce080_5818 , \47192 , \48202 );
_HMUX g17165 ( \48219_nG17165 , RIe1ce080_5818 , \48218_nG17164 , \47166 );
_HMUX g17166 ( \48220_nG17166 , RIe1ce080_5818 , \47195 , \48205 );
_HMUX g17167 ( \48221_nG17167 , \48219_nG17165 , \48220_nG17166 , \47178 );
buf \U$38817 ( \48222 , \48221_nG17167 );
_DC g18f2d_GF_IsGateDCbyConstraint ( \48223_nG18f2d , \48222 , \42503 );
buf \U$38818 ( \48224 , \48223_nG18f2d );
_HMUX g17168 ( \48225_nG17168 , RIe1cc550_5819 , \47201 , \48202 );
_HMUX g17169 ( \48226_nG17169 , RIe1cc550_5819 , \48225_nG17168 , \47166 );
_HMUX g1716a ( \48227_nG1716a , RIe1cc550_5819 , \47204 , \48205 );
_HMUX g1716b ( \48228_nG1716b , \48226_nG17169 , \48227_nG1716a , \47178 );
buf \U$38819 ( \48229 , \48228_nG1716b );
_DC g18f43_GF_IsGateDCbyConstraint ( \48230_nG18f43 , \48229 , \42503 );
buf \U$38820 ( \48231 , \48230_nG18f43 );
_HMUX g1716c ( \48232_nG1716c , RIe1ca048_5820 , \47210 , \48202 );
_HMUX g1716d ( \48233_nG1716d , RIe1ca048_5820 , \48232_nG1716c , \47166 );
_HMUX g1716e ( \48234_nG1716e , RIe1ca048_5820 , \47213 , \48205 );
_HMUX g1716f ( \48235_nG1716f , \48233_nG1716d , \48234_nG1716e , \47178 );
buf \U$38821 ( \48236 , \48235_nG1716f );
_DC g18f59_GF_IsGateDCbyConstraint ( \48237_nG18f59 , \48236 , \42503 );
buf \U$38822 ( \48238 , \48237_nG18f59 );
_HMUX g17170 ( \48239_nG17170 , RIe1c78e8_5821 , \47219 , \48202 );
_HMUX g17171 ( \48240_nG17171 , RIe1c78e8_5821 , \48239_nG17170 , \47166 );
_HMUX g17172 ( \48241_nG17172 , RIe1c78e8_5821 , \47222 , \48205 );
_HMUX g17173 ( \48242_nG17173 , \48240_nG17171 , \48241_nG17172 , \47178 );
buf \U$38823 ( \48243 , \48242_nG17173 );
_DC g18f6f_GF_IsGateDCbyConstraint ( \48244_nG18f6f , \48243 , \42503 );
buf \U$38824 ( \48245 , \48244_nG18f6f );
_HMUX g17174 ( \48246_nG17174 , RIe1c4f30_5822 , \47228 , \48202 );
_HMUX g17175 ( \48247_nG17175 , RIe1c4f30_5822 , \48246_nG17174 , \47166 );
_HMUX g17176 ( \48248_nG17176 , RIe1c4f30_5822 , \47231 , \48205 );
_HMUX g17177 ( \48249_nG17177 , \48247_nG17175 , \48248_nG17176 , \47178 );
buf \U$38825 ( \48250 , \48249_nG17177 );
_DC g18f7b_GF_IsGateDCbyConstraint ( \48251_nG18f7b , \48250 , \42503 );
buf \U$38826 ( \48252 , \48251_nG18f7b );
_HMUX g17178 ( \48253_nG17178 , RIe1c26e0_5823 , \47237 , \48202 );
_HMUX g17179 ( \48254_nG17179 , RIe1c26e0_5823 , \48253_nG17178 , \47166 );
_HMUX g1717a ( \48255_nG1717a , RIe1c26e0_5823 , \47240 , \48205 );
_HMUX g1717b ( \48256_nG1717b , \48254_nG17179 , \48255_nG1717a , \47178 );
buf \U$38827 ( \48257 , \48256_nG1717b );
_DC g18f7d_GF_IsGateDCbyConstraint ( \48258_nG18f7d , \48257 , \42503 );
buf \U$38828 ( \48259 , \48258_nG18f7d );
_HMUX g1717c ( \48260_nG1717c , RIe1c0b38_5824 , \47246 , \48202 );
_HMUX g1717d ( \48261_nG1717d , RIe1c0b38_5824 , \48260_nG1717c , \47166 );
_HMUX g1717e ( \48262_nG1717e , RIe1c0b38_5824 , \47249 , \48205 );
_HMUX g1717f ( \48263_nG1717f , \48261_nG1717d , \48262_nG1717e , \47178 );
buf \U$38829 ( \48264 , \48263_nG1717f );
_DC g18f7f_GF_IsGateDCbyConstraint ( \48265_nG18f7f , \48264 , \42503 );
buf \U$38830 ( \48266 , \48265_nG18f7f );
_HMUX g17180 ( \48267_nG17180 , RIe1be9f0_5825 , \47255 , \48202 );
_HMUX g17181 ( \48268_nG17181 , RIe1be9f0_5825 , \48267_nG17180 , \47166 );
_HMUX g17182 ( \48269_nG17182 , RIe1be9f0_5825 , \47258 , \48205 );
_HMUX g17183 ( \48270_nG17183 , \48268_nG17181 , \48269_nG17182 , \47178 );
buf \U$38831 ( \48271 , \48270_nG17183 );
_DC g18f03_GF_IsGateDCbyConstraint ( \48272_nG18f03 , \48271 , \42503 );
buf \U$38832 ( \48273 , \48272_nG18f03 );
_HMUX g17184 ( \48274_nG17184 , RIe1bcce0_5826 , \47264 , \48202 );
_HMUX g17185 ( \48275_nG17185 , RIe1bcce0_5826 , \48274_nG17184 , \47166 );
_HMUX g17186 ( \48276_nG17186 , RIe1bcce0_5826 , \47267 , \48205 );
_HMUX g17187 ( \48277_nG17187 , \48275_nG17185 , \48276_nG17186 , \47178 );
buf \U$38833 ( \48278 , \48277_nG17187 );
_DC g18f05_GF_IsGateDCbyConstraint ( \48279_nG18f05 , \48278 , \42503 );
buf \U$38834 ( \48280 , \48279_nG18f05 );
_HMUX g17188 ( \48281_nG17188 , RIe1baf58_5827 , \47273 , \48202 );
_HMUX g17189 ( \48282_nG17189 , RIe1baf58_5827 , \48281_nG17188 , \47166 );
_HMUX g1718a ( \48283_nG1718a , RIe1baf58_5827 , \47276 , \48205 );
_HMUX g1718b ( \48284_nG1718b , \48282_nG17189 , \48283_nG1718a , \47178 );
buf \U$38835 ( \48285 , \48284_nG1718b );
_DC g18f07_GF_IsGateDCbyConstraint ( \48286_nG18f07 , \48285 , \42503 );
buf \U$38836 ( \48287 , \48286_nG18f07 );
_HMUX g1718c ( \48288_nG1718c , RIe1b9158_5828 , \47282 , \48202 );
_HMUX g1718d ( \48289_nG1718d , RIe1b9158_5828 , \48288_nG1718c , \47166 );
_HMUX g1718e ( \48290_nG1718e , RIe1b9158_5828 , \47285 , \48205 );
_HMUX g1718f ( \48291_nG1718f , \48289_nG1718d , \48290_nG1718e , \47178 );
buf \U$38837 ( \48292 , \48291_nG1718f );
_DC g18f09_GF_IsGateDCbyConstraint ( \48293_nG18f09 , \48292 , \42503 );
buf \U$38838 ( \48294 , \48293_nG18f09 );
_HMUX g17190 ( \48295_nG17190 , RIe1b6908_5829 , \47291 , \48202 );
_HMUX g17191 ( \48296_nG17191 , RIe1b6908_5829 , \48295_nG17190 , \47166 );
_HMUX g17192 ( \48297_nG17192 , RIe1b6908_5829 , \47294 , \48205 );
_HMUX g17193 ( \48298_nG17193 , \48296_nG17191 , \48297_nG17192 , \47178 );
buf \U$38839 ( \48299 , \48298_nG17193 );
_DC g18f0b_GF_IsGateDCbyConstraint ( \48300_nG18f0b , \48299 , \42503 );
buf \U$38840 ( \48301 , \48300_nG18f0b );
_HMUX g17194 ( \48302_nG17194 , RIe1b3b90_5830 , \47300 , \48202 );
_HMUX g17195 ( \48303_nG17195 , RIe1b3b90_5830 , \48302_nG17194 , \47166 );
_HMUX g17196 ( \48304_nG17196 , RIe1b3b90_5830 , \47303 , \48205 );
_HMUX g17197 ( \48305_nG17197 , \48303_nG17195 , \48304_nG17196 , \47178 );
buf \U$38841 ( \48306 , \48305_nG17197 );
_DC g18f0d_GF_IsGateDCbyConstraint ( \48307_nG18f0d , \48306 , \42503 );
buf \U$38842 ( \48308 , \48307_nG18f0d );
_HMUX g17198 ( \48309_nG17198 , RIe1b1d18_5831 , \47309 , \48202 );
_HMUX g17199 ( \48310_nG17199 , RIe1b1d18_5831 , \48309_nG17198 , \47166 );
_HMUX g1719a ( \48311_nG1719a , RIe1b1d18_5831 , \47312 , \48205 );
_HMUX g1719b ( \48312_nG1719b , \48310_nG17199 , \48311_nG1719a , \47178 );
buf \U$38843 ( \48313 , \48312_nG1719b );
_DC g18f0f_GF_IsGateDCbyConstraint ( \48314_nG18f0f , \48313 , \42503 );
buf \U$38844 ( \48315 , \48314_nG18f0f );
_HMUX g1719c ( \48316_nG1719c , RIe1aff90_5832 , \47318 , \48202 );
_HMUX g1719d ( \48317_nG1719d , RIe1aff90_5832 , \48316_nG1719c , \47166 );
_HMUX g1719e ( \48318_nG1719e , RIe1aff90_5832 , \47321 , \48205 );
_HMUX g1719f ( \48319_nG1719f , \48317_nG1719d , \48318_nG1719e , \47178 );
buf \U$38845 ( \48320 , \48319_nG1719f );
_DC g18f11_GF_IsGateDCbyConstraint ( \48321_nG18f11 , \48320 , \42503 );
buf \U$38846 ( \48322 , \48321_nG18f11 );
_HMUX g171a0 ( \48323_nG171a0 , RIe1ae2f8_5833 , \47327 , \48202 );
_HMUX g171a1 ( \48324_nG171a1 , RIe1ae2f8_5833 , \48323_nG171a0 , \47166 );
_HMUX g171a2 ( \48325_nG171a2 , RIe1ae2f8_5833 , \47330 , \48205 );
_HMUX g171a3 ( \48326_nG171a3 , \48324_nG171a1 , \48325_nG171a2 , \47178 );
buf \U$38847 ( \48327 , \48326_nG171a3 );
_DC g18f13_GF_IsGateDCbyConstraint ( \48328_nG18f13 , \48327 , \42503 );
buf \U$38848 ( \48329 , \48328_nG18f13 );
_HMUX g171a4 ( \48330_nG171a4 , RIe1ab940_5834 , \47336 , \48202 );
_HMUX g171a5 ( \48331_nG171a5 , RIe1ab940_5834 , \48330_nG171a4 , \47166 );
_HMUX g171a6 ( \48332_nG171a6 , RIe1ab940_5834 , \47339 , \48205 );
_HMUX g171a7 ( \48333_nG171a7 , \48331_nG171a5 , \48332_nG171a6 , \47178 );
buf \U$38849 ( \48334 , \48333_nG171a7 );
_DC g18f15_GF_IsGateDCbyConstraint ( \48335_nG18f15 , \48334 , \42503 );
buf \U$38850 ( \48336 , \48335_nG18f15 );
_HMUX g171a8 ( \48337_nG171a8 , RIe1a8628_5835 , \47345 , \48202 );
_HMUX g171a9 ( \48338_nG171a9 , RIe1a8628_5835 , \48337_nG171a8 , \47166 );
_HMUX g171aa ( \48339_nG171aa , RIe1a8628_5835 , \47348 , \48205 );
_HMUX g171ab ( \48340_nG171ab , \48338_nG171a9 , \48339_nG171aa , \47178 );
buf \U$38851 ( \48341 , \48340_nG171ab );
_DC g18f19_GF_IsGateDCbyConstraint ( \48342_nG18f19 , \48341 , \42503 );
buf \U$38852 ( \48343 , \48342_nG18f19 );
_HMUX g171ac ( \48344_nG171ac , RIe1a6030_5836 , \47354 , \48202 );
_HMUX g171ad ( \48345_nG171ad , RIe1a6030_5836 , \48344_nG171ac , \47166 );
_HMUX g171ae ( \48346_nG171ae , RIe1a6030_5836 , \47357 , \48205 );
_HMUX g171af ( \48347_nG171af , \48345_nG171ad , \48346_nG171ae , \47178 );
buf \U$38853 ( \48348 , \48347_nG171af );
_DC g18f1b_GF_IsGateDCbyConstraint ( \48349_nG18f1b , \48348 , \42503 );
buf \U$38854 ( \48350 , \48349_nG18f1b );
_HMUX g171b0 ( \48351_nG171b0 , RIe1a2d90_5837 , \47363 , \48202 );
_HMUX g171b1 ( \48352_nG171b1 , RIe1a2d90_5837 , \48351_nG171b0 , \47166 );
_HMUX g171b2 ( \48353_nG171b2 , RIe1a2d90_5837 , \47366 , \48205 );
_HMUX g171b3 ( \48354_nG171b3 , \48352_nG171b1 , \48353_nG171b2 , \47178 );
buf \U$38855 ( \48355 , \48354_nG171b3 );
_DC g18f1d_GF_IsGateDCbyConstraint ( \48356_nG18f1d , \48355 , \42503 );
buf \U$38856 ( \48357 , \48356_nG18f1d );
_HMUX g171b4 ( \48358_nG171b4 , RIe1a0540_5838 , \47372 , \48202 );
_HMUX g171b5 ( \48359_nG171b5 , RIe1a0540_5838 , \48358_nG171b4 , \47166 );
_HMUX g171b6 ( \48360_nG171b6 , RIe1a0540_5838 , \47375 , \48205 );
_HMUX g171b7 ( \48361_nG171b7 , \48359_nG171b5 , \48360_nG171b6 , \47178 );
buf \U$38857 ( \48362 , \48361_nG171b7 );
_DC g18f1f_GF_IsGateDCbyConstraint ( \48363_nG18f1f , \48362 , \42503 );
buf \U$38858 ( \48364 , \48363_nG18f1f );
_HMUX g171b8 ( \48365_nG171b8 , RIe19da20_5839 , \47381 , \48202 );
_HMUX g171b9 ( \48366_nG171b9 , RIe19da20_5839 , \48365_nG171b8 , \47166 );
_HMUX g171ba ( \48367_nG171ba , RIe19da20_5839 , \47384 , \48205 );
_HMUX g171bb ( \48368_nG171bb , \48366_nG171b9 , \48367_nG171ba , \47178 );
buf \U$38859 ( \48369 , \48368_nG171bb );
_DC g18f21_GF_IsGateDCbyConstraint ( \48370_nG18f21 , \48369 , \42503 );
buf \U$38860 ( \48371 , \48370_nG18f21 );
_HMUX g171bc ( \48372_nG171bc , RIe19a870_5840 , \47390 , \48202 );
_HMUX g171bd ( \48373_nG171bd , RIe19a870_5840 , \48372_nG171bc , \47166 );
_HMUX g171be ( \48374_nG171be , RIe19a870_5840 , \47393 , \48205 );
_HMUX g171bf ( \48375_nG171bf , \48373_nG171bd , \48374_nG171be , \47178 );
buf \U$38861 ( \48376 , \48375_nG171bf );
_DC g18f23_GF_IsGateDCbyConstraint ( \48377_nG18f23 , \48376 , \42503 );
buf \U$38862 ( \48378 , \48377_nG18f23 );
_HMUX g171c0 ( \48379_nG171c0 , RIe197cd8_5841 , \47399 , \48202 );
_HMUX g171c1 ( \48380_nG171c1 , RIe197cd8_5841 , \48379_nG171c0 , \47166 );
_HMUX g171c2 ( \48381_nG171c2 , RIe197cd8_5841 , \47402 , \48205 );
_HMUX g171c3 ( \48382_nG171c3 , \48380_nG171c1 , \48381_nG171c2 , \47178 );
buf \U$38863 ( \48383 , \48382_nG171c3 );
_DC g18f25_GF_IsGateDCbyConstraint ( \48384_nG18f25 , \48383 , \42503 );
buf \U$38864 ( \48385 , \48384_nG18f25 );
_HMUX g171c4 ( \48386_nG171c4 , RIe195410_5842 , \47408 , \48202 );
_HMUX g171c5 ( \48387_nG171c5 , RIe195410_5842 , \48386_nG171c4 , \47166 );
_HMUX g171c6 ( \48388_nG171c6 , RIe195410_5842 , \47411 , \48205 );
_HMUX g171c7 ( \48389_nG171c7 , \48387_nG171c5 , \48388_nG171c6 , \47178 );
buf \U$38865 ( \48390 , \48389_nG171c7 );
_DC g18f27_GF_IsGateDCbyConstraint ( \48391_nG18f27 , \48390 , \42503 );
buf \U$38866 ( \48392 , \48391_nG18f27 );
_HMUX g171c8 ( \48393_nG171c8 , RIe192e90_5843 , \47417 , \48202 );
_HMUX g171c9 ( \48394_nG171c9 , RIe192e90_5843 , \48393_nG171c8 , \47166 );
_HMUX g171ca ( \48395_nG171ca , RIe192e90_5843 , \47420 , \48205 );
_HMUX g171cb ( \48396_nG171cb , \48394_nG171c9 , \48395_nG171ca , \47178 );
buf \U$38867 ( \48397 , \48396_nG171cb );
_DC g18f29_GF_IsGateDCbyConstraint ( \48398_nG18f29 , \48397 , \42503 );
buf \U$38868 ( \48399 , \48398_nG18f29 );
_HMUX g171cc ( \48400_nG171cc , RIe190460_5844 , \47426 , \48202 );
_HMUX g171cd ( \48401_nG171cd , RIe190460_5844 , \48400_nG171cc , \47166 );
_HMUX g171ce ( \48402_nG171ce , RIe190460_5844 , \47429 , \48205 );
_HMUX g171cf ( \48403_nG171cf , \48401_nG171cd , \48402_nG171ce , \47178 );
buf \U$38869 ( \48404 , \48403_nG171cf );
_DC g18f2b_GF_IsGateDCbyConstraint ( \48405_nG18f2b , \48404 , \42503 );
buf \U$38870 ( \48406 , \48405_nG18f2b );
_HMUX g171d0 ( \48407_nG171d0 , RIe18e0c0_5845 , \47435 , \48202 );
_HMUX g171d1 ( \48408_nG171d1 , RIe18e0c0_5845 , \48407_nG171d0 , \47166 );
_HMUX g171d2 ( \48409_nG171d2 , RIe18e0c0_5845 , \47438 , \48205 );
_HMUX g171d3 ( \48410_nG171d3 , \48408_nG171d1 , \48409_nG171d2 , \47178 );
buf \U$38871 ( \48411 , \48410_nG171d3 );
_DC g18f2f_GF_IsGateDCbyConstraint ( \48412_nG18f2f , \48411 , \42503 );
buf \U$38872 ( \48413 , \48412_nG18f2f );
_HMUX g171d4 ( \48414_nG171d4 , RIe18bc30_5846 , \47444 , \48202 );
_HMUX g171d5 ( \48415_nG171d5 , RIe18bc30_5846 , \48414_nG171d4 , \47166 );
_HMUX g171d6 ( \48416_nG171d6 , RIe18bc30_5846 , \47447 , \48205 );
_HMUX g171d7 ( \48417_nG171d7 , \48415_nG171d5 , \48416_nG171d6 , \47178 );
buf \U$38873 ( \48418 , \48417_nG171d7 );
_DC g18f31_GF_IsGateDCbyConstraint ( \48419_nG18f31 , \48418 , \42503 );
buf \U$38874 ( \48420 , \48419_nG18f31 );
_HMUX g171d8 ( \48421_nG171d8 , RIe189098_5847 , \47453 , \48202 );
_HMUX g171d9 ( \48422_nG171d9 , RIe189098_5847 , \48421_nG171d8 , \47166 );
_HMUX g171da ( \48423_nG171da , RIe189098_5847 , \47456 , \48205 );
_HMUX g171db ( \48424_nG171db , \48422_nG171d9 , \48423_nG171da , \47178 );
buf \U$38875 ( \48425 , \48424_nG171db );
_DC g18f33_GF_IsGateDCbyConstraint ( \48426_nG18f33 , \48425 , \42503 );
buf \U$38876 ( \48427 , \48426_nG18f33 );
_HMUX g171dc ( \48428_nG171dc , RIe186c08_5848 , \47462 , \48202 );
_HMUX g171dd ( \48429_nG171dd , RIe186c08_5848 , \48428_nG171dc , \47166 );
_HMUX g171de ( \48430_nG171de , RIe186c08_5848 , \47465 , \48205 );
_HMUX g171df ( \48431_nG171df , \48429_nG171dd , \48430_nG171de , \47178 );
buf \U$38877 ( \48432 , \48431_nG171df );
_DC g18f35_GF_IsGateDCbyConstraint ( \48433_nG18f35 , \48432 , \42503 );
buf \U$38878 ( \48434 , \48433_nG18f35 );
_HMUX g171e0 ( \48435_nG171e0 , RIe1839e0_5849 , \47471 , \48202 );
_HMUX g171e1 ( \48436_nG171e1 , RIe1839e0_5849 , \48435_nG171e0 , \47166 );
_HMUX g171e2 ( \48437_nG171e2 , RIe1839e0_5849 , \47474 , \48205 );
_HMUX g171e3 ( \48438_nG171e3 , \48436_nG171e1 , \48437_nG171e2 , \47178 );
buf \U$38879 ( \48439 , \48438_nG171e3 );
_DC g18f37_GF_IsGateDCbyConstraint ( \48440_nG18f37 , \48439 , \42503 );
buf \U$38880 ( \48441 , \48440_nG18f37 );
_HMUX g171e4 ( \48442_nG171e4 , RIe1817a8_5850 , \47480 , \48202 );
_HMUX g171e5 ( \48443_nG171e5 , RIe1817a8_5850 , \48442_nG171e4 , \47166 );
_HMUX g171e6 ( \48444_nG171e6 , RIe1817a8_5850 , \47483 , \48205 );
_HMUX g171e7 ( \48445_nG171e7 , \48443_nG171e5 , \48444_nG171e6 , \47178 );
buf \U$38881 ( \48446 , \48445_nG171e7 );
_DC g18f39_GF_IsGateDCbyConstraint ( \48447_nG18f39 , \48446 , \42503 );
buf \U$38882 ( \48448 , \48447_nG18f39 );
_HMUX g171e8 ( \48449_nG171e8 , RIe17fb88_5851 , \47489 , \48202 );
_HMUX g171e9 ( \48450_nG171e9 , RIe17fb88_5851 , \48449_nG171e8 , \47166 );
_HMUX g171ea ( \48451_nG171ea , RIe17fb88_5851 , \47492 , \48205 );
_HMUX g171eb ( \48452_nG171eb , \48450_nG171e9 , \48451_nG171ea , \47178 );
buf \U$38883 ( \48453 , \48452_nG171eb );
_DC g18f3b_GF_IsGateDCbyConstraint ( \48454_nG18f3b , \48453 , \42503 );
buf \U$38884 ( \48455 , \48454_nG18f3b );
_HMUX g171ec ( \48456_nG171ec , RIe17def0_5852 , \47498 , \48202 );
_HMUX g171ed ( \48457_nG171ed , RIe17def0_5852 , \48456_nG171ec , \47166 );
_HMUX g171ee ( \48458_nG171ee , RIe17def0_5852 , \47501 , \48205 );
_HMUX g171ef ( \48459_nG171ef , \48457_nG171ed , \48458_nG171ee , \47178 );
buf \U$38885 ( \48460 , \48459_nG171ef );
_DC g18f3d_GF_IsGateDCbyConstraint ( \48461_nG18f3d , \48460 , \42503 );
buf \U$38886 ( \48462 , \48461_nG18f3d );
_HMUX g171f0 ( \48463_nG171f0 , RIe17c3c0_5853 , \47507 , \48202 );
_HMUX g171f1 ( \48464_nG171f1 , RIe17c3c0_5853 , \48463_nG171f0 , \47166 );
_HMUX g171f2 ( \48465_nG171f2 , RIe17c3c0_5853 , \47510 , \48205 );
_HMUX g171f3 ( \48466_nG171f3 , \48464_nG171f1 , \48465_nG171f2 , \47178 );
buf \U$38887 ( \48467 , \48466_nG171f3 );
_DC g18f3f_GF_IsGateDCbyConstraint ( \48468_nG18f3f , \48467 , \42503 );
buf \U$38888 ( \48469 , \48468_nG18f3f );
_HMUX g171f4 ( \48470_nG171f4 , RIe17a458_5854 , \47516 , \48202 );
_HMUX g171f5 ( \48471_nG171f5 , RIe17a458_5854 , \48470_nG171f4 , \47166 );
_HMUX g171f6 ( \48472_nG171f6 , RIe17a458_5854 , \47519 , \48205 );
_HMUX g171f7 ( \48473_nG171f7 , \48471_nG171f5 , \48472_nG171f6 , \47178 );
buf \U$38889 ( \48474 , \48473_nG171f7 );
_DC g18f41_GF_IsGateDCbyConstraint ( \48475_nG18f41 , \48474 , \42503 );
buf \U$38890 ( \48476 , \48475_nG18f41 );
_HMUX g171f8 ( \48477_nG171f8 , RIe1781a8_5855 , \47525 , \48202 );
_HMUX g171f9 ( \48478_nG171f9 , RIe1781a8_5855 , \48477_nG171f8 , \47166 );
_HMUX g171fa ( \48479_nG171fa , RIe1781a8_5855 , \47528 , \48205 );
_HMUX g171fb ( \48480_nG171fb , \48478_nG171f9 , \48479_nG171fa , \47178 );
buf \U$38891 ( \48481 , \48480_nG171fb );
_DC g18f45_GF_IsGateDCbyConstraint ( \48482_nG18f45 , \48481 , \42503 );
buf \U$38892 ( \48483 , \48482_nG18f45 );
_HMUX g171fc ( \48484_nG171fc , RIe176240_5856 , \47534 , \48202 );
_HMUX g171fd ( \48485_nG171fd , RIe176240_5856 , \48484_nG171fc , \47166 );
_HMUX g171fe ( \48486_nG171fe , RIe176240_5856 , \47537 , \48205 );
_HMUX g171ff ( \48487_nG171ff , \48485_nG171fd , \48486_nG171fe , \47178 );
buf \U$38893 ( \48488 , \48487_nG171ff );
_DC g18f47_GF_IsGateDCbyConstraint ( \48489_nG18f47 , \48488 , \42503 );
buf \U$38894 ( \48490 , \48489_nG18f47 );
_HMUX g17200 ( \48491_nG17200 , RIe174530_5857 , \47543 , \48202 );
_HMUX g17201 ( \48492_nG17201 , RIe174530_5857 , \48491_nG17200 , \47166 );
_HMUX g17202 ( \48493_nG17202 , RIe174530_5857 , \47546 , \48205 );
_HMUX g17203 ( \48494_nG17203 , \48492_nG17201 , \48493_nG17202 , \47178 );
buf \U$38895 ( \48495 , \48494_nG17203 );
_DC g18f49_GF_IsGateDCbyConstraint ( \48496_nG18f49 , \48495 , \42503 );
buf \U$38896 ( \48497 , \48496_nG18f49 );
_HMUX g17204 ( \48498_nG17204 , RIe172988_5858 , \47552 , \48202 );
_HMUX g17205 ( \48499_nG17205 , RIe172988_5858 , \48498_nG17204 , \47166 );
_HMUX g17206 ( \48500_nG17206 , RIe172988_5858 , \47555 , \48205 );
_HMUX g17207 ( \48501_nG17207 , \48499_nG17205 , \48500_nG17206 , \47178 );
buf \U$38897 ( \48502 , \48501_nG17207 );
_DC g18f4b_GF_IsGateDCbyConstraint ( \48503_nG18f4b , \48502 , \42503 );
buf \U$38898 ( \48504 , \48503_nG18f4b );
_HMUX g17208 ( \48505_nG17208 , RIe16fc70_5859 , \47561 , \48202 );
_HMUX g17209 ( \48506_nG17209 , RIe16fc70_5859 , \48505_nG17208 , \47166 );
_HMUX g1720a ( \48507_nG1720a , RIe16fc70_5859 , \47564 , \48205 );
_HMUX g1720b ( \48508_nG1720b , \48506_nG17209 , \48507_nG1720a , \47178 );
buf \U$38899 ( \48509 , \48508_nG1720b );
_DC g18f4d_GF_IsGateDCbyConstraint ( \48510_nG18f4d , \48509 , \42503 );
buf \U$38900 ( \48511 , \48510_nG18f4d );
_HMUX g1720c ( \48512_nG1720c , RIe16e140_5860 , \47570 , \48202 );
_HMUX g1720d ( \48513_nG1720d , RIe16e140_5860 , \48512_nG1720c , \47166 );
_HMUX g1720e ( \48514_nG1720e , RIe16e140_5860 , \47573 , \48205 );
_HMUX g1720f ( \48515_nG1720f , \48513_nG1720d , \48514_nG1720e , \47178 );
buf \U$38901 ( \48516 , \48515_nG1720f );
_DC g18f4f_GF_IsGateDCbyConstraint ( \48517_nG18f4f , \48516 , \42503 );
buf \U$38902 ( \48518 , \48517_nG18f4f );
_HMUX g17210 ( \48519_nG17210 , RIe16c1d8_5861 , \47579 , \48202 );
_HMUX g17211 ( \48520_nG17211 , RIe16c1d8_5861 , \48519_nG17210 , \47166 );
_HMUX g17212 ( \48521_nG17212 , RIe16c1d8_5861 , \47582 , \48205 );
_HMUX g17213 ( \48522_nG17213 , \48520_nG17211 , \48521_nG17212 , \47178 );
buf \U$38903 ( \48523 , \48522_nG17213 );
_DC g18f51_GF_IsGateDCbyConstraint ( \48524_nG18f51 , \48523 , \42503 );
buf \U$38904 ( \48525 , \48524_nG18f51 );
_HMUX g17214 ( \48526_nG17214 , RIe16a5b8_5862 , \47588 , \48202 );
_HMUX g17215 ( \48527_nG17215 , RIe16a5b8_5862 , \48526_nG17214 , \47166 );
_HMUX g17216 ( \48528_nG17216 , RIe16a5b8_5862 , \47591 , \48205 );
_HMUX g17217 ( \48529_nG17217 , \48527_nG17215 , \48528_nG17216 , \47178 );
buf \U$38905 ( \48530 , \48529_nG17217 );
_DC g18f53_GF_IsGateDCbyConstraint ( \48531_nG18f53 , \48530 , \42503 );
buf \U$38906 ( \48532 , \48531_nG18f53 );
_HMUX g17218 ( \48533_nG17218 , RIe168a88_5863 , \47597 , \48202 );
_HMUX g17219 ( \48534_nG17219 , RIe168a88_5863 , \48533_nG17218 , \47166 );
_HMUX g1721a ( \48535_nG1721a , RIe168a88_5863 , \47600 , \48205 );
_HMUX g1721b ( \48536_nG1721b , \48534_nG17219 , \48535_nG1721a , \47178 );
buf \U$38907 ( \48537 , \48536_nG1721b );
_DC g18f55_GF_IsGateDCbyConstraint ( \48538_nG18f55 , \48537 , \42503 );
buf \U$38908 ( \48539 , \48538_nG18f55 );
_HMUX g1721c ( \48540_nG1721c , RIe167138_5864 , \47606 , \48202 );
_HMUX g1721d ( \48541_nG1721d , RIe167138_5864 , \48540_nG1721c , \47166 );
_HMUX g1721e ( \48542_nG1721e , RIe167138_5864 , \47609 , \48205 );
_HMUX g1721f ( \48543_nG1721f , \48541_nG1721d , \48542_nG1721e , \47178 );
buf \U$38909 ( \48544 , \48543_nG1721f );
_DC g18f57_GF_IsGateDCbyConstraint ( \48545_nG18f57 , \48544 , \42503 );
buf \U$38910 ( \48546 , \48545_nG18f57 );
_HMUX g17220 ( \48547_nG17220 , RIe39c680_5865 , \47615 , \48202 );
_HMUX g17221 ( \48548_nG17221 , RIe39c680_5865 , \48547_nG17220 , \47166 );
_HMUX g17222 ( \48549_nG17222 , RIe39c680_5865 , \47618 , \48205 );
_HMUX g17223 ( \48550_nG17223 , \48548_nG17221 , \48549_nG17222 , \47178 );
buf \U$38911 ( \48551 , \48550_nG17223 );
_DC g18f5b_GF_IsGateDCbyConstraint ( \48552_nG18f5b , \48551 , \42503 );
buf \U$38912 ( \48553 , \48552_nG18f5b );
_HMUX g17224 ( \48554_nG17224 , RIe39ce78_5866 , \47624 , \48202 );
_HMUX g17225 ( \48555_nG17225 , RIe39ce78_5866 , \48554_nG17224 , \47166 );
_HMUX g17226 ( \48556_nG17226 , RIe39ce78_5866 , \47627 , \48205 );
_HMUX g17227 ( \48557_nG17227 , \48555_nG17225 , \48556_nG17226 , \47178 );
buf \U$38913 ( \48558 , \48557_nG17227 );
_DC g18f5d_GF_IsGateDCbyConstraint ( \48559_nG18f5d , \48558 , \42503 );
buf \U$38914 ( \48560 , \48559_nG18f5d );
_HMUX g17228 ( \48561_nG17228 , RIe39d670_5867 , \47633 , \48202 );
_HMUX g17229 ( \48562_nG17229 , RIe39d670_5867 , \48561_nG17228 , \47166 );
_HMUX g1722a ( \48563_nG1722a , RIe39d670_5867 , \47636 , \48205 );
_HMUX g1722b ( \48564_nG1722b , \48562_nG17229 , \48563_nG1722a , \47178 );
buf \U$38915 ( \48565 , \48564_nG1722b );
_DC g18f5f_GF_IsGateDCbyConstraint ( \48566_nG18f5f , \48565 , \42503 );
buf \U$38916 ( \48567 , \48566_nG18f5f );
_HMUX g1722c ( \48568_nG1722c , RIe39de68_5868 , \47642 , \48202 );
_HMUX g1722d ( \48569_nG1722d , RIe39de68_5868 , \48568_nG1722c , \47166 );
_HMUX g1722e ( \48570_nG1722e , RIe39de68_5868 , \47645 , \48205 );
_HMUX g1722f ( \48571_nG1722f , \48569_nG1722d , \48570_nG1722e , \47178 );
buf \U$38917 ( \48572 , \48571_nG1722f );
_DC g18f61_GF_IsGateDCbyConstraint ( \48573_nG18f61 , \48572 , \42503 );
buf \U$38918 ( \48574 , \48573_nG18f61 );
_HMUX g17230 ( \48575_nG17230 , RIe39e660_5869 , \47651 , \48202 );
_HMUX g17231 ( \48576_nG17231 , RIe39e660_5869 , \48575_nG17230 , \47166 );
_HMUX g17232 ( \48577_nG17232 , RIe39e660_5869 , \47654 , \48205 );
_HMUX g17233 ( \48578_nG17233 , \48576_nG17231 , \48577_nG17232 , \47178 );
buf \U$38919 ( \48579 , \48578_nG17233 );
_DC g18f63_GF_IsGateDCbyConstraint ( \48580_nG18f63 , \48579 , \42503 );
buf \U$38920 ( \48581 , \48580_nG18f63 );
_HMUX g17234 ( \48582_nG17234 , RIe39ee58_5870 , \47660 , \48202 );
_HMUX g17235 ( \48583_nG17235 , RIe39ee58_5870 , \48582_nG17234 , \47166 );
_HMUX g17236 ( \48584_nG17236 , RIe39ee58_5870 , \47663 , \48205 );
_HMUX g17237 ( \48585_nG17237 , \48583_nG17235 , \48584_nG17236 , \47178 );
buf \U$38921 ( \48586 , \48585_nG17237 );
_DC g18f65_GF_IsGateDCbyConstraint ( \48587_nG18f65 , \48586 , \42503 );
buf \U$38922 ( \48588 , \48587_nG18f65 );
_HMUX g17238 ( \48589_nG17238 , RIe39f650_5871 , \47669 , \48202 );
_HMUX g17239 ( \48590_nG17239 , RIe39f650_5871 , \48589_nG17238 , \47166 );
_HMUX g1723a ( \48591_nG1723a , RIe39f650_5871 , \47672 , \48205 );
_HMUX g1723b ( \48592_nG1723b , \48590_nG17239 , \48591_nG1723a , \47178 );
buf \U$38923 ( \48593 , \48592_nG1723b );
_DC g18f67_GF_IsGateDCbyConstraint ( \48594_nG18f67 , \48593 , \42503 );
buf \U$38924 ( \48595 , \48594_nG18f67 );
_HMUX g1723c ( \48596_nG1723c , RIe39fe48_5872 , \47678 , \48202 );
_HMUX g1723d ( \48597_nG1723d , RIe39fe48_5872 , \48596_nG1723c , \47166 );
_HMUX g1723e ( \48598_nG1723e , RIe39fe48_5872 , \47681 , \48205 );
_HMUX g1723f ( \48599_nG1723f , \48597_nG1723d , \48598_nG1723e , \47178 );
buf \U$38925 ( \48600 , \48599_nG1723f );
_DC g18f69_GF_IsGateDCbyConstraint ( \48601_nG18f69 , \48600 , \42503 );
buf \U$38926 ( \48602 , \48601_nG18f69 );
_HMUX g17240 ( \48603_nG17240 , RIe3a0640_5873 , \47687 , \48202 );
_HMUX g17241 ( \48604_nG17241 , RIe3a0640_5873 , \48603_nG17240 , \47166 );
_HMUX g17242 ( \48605_nG17242 , RIe3a0640_5873 , \47690 , \48205 );
_HMUX g17243 ( \48606_nG17243 , \48604_nG17241 , \48605_nG17242 , \47178 );
buf \U$38927 ( \48607 , \48606_nG17243 );
_DC g18f6b_GF_IsGateDCbyConstraint ( \48608_nG18f6b , \48607 , \42503 );
buf \U$38928 ( \48609 , \48608_nG18f6b );
_HMUX g17244 ( \48610_nG17244 , RIe3a0e38_5874 , \47696 , \48202 );
_HMUX g17245 ( \48611_nG17245 , RIe3a0e38_5874 , \48610_nG17244 , \47166 );
_HMUX g17246 ( \48612_nG17246 , RIe3a0e38_5874 , \47699 , \48205 );
_HMUX g17247 ( \48613_nG17247 , \48611_nG17245 , \48612_nG17246 , \47178 );
buf \U$38929 ( \48614 , \48613_nG17247 );
_DC g18f6d_GF_IsGateDCbyConstraint ( \48615_nG18f6d , \48614 , \42503 );
buf \U$38930 ( \48616 , \48615_nG18f6d );
_HMUX g17248 ( \48617_nG17248 , RIe3a1630_5875 , \47705 , \48202 );
_HMUX g17249 ( \48618_nG17249 , RIe3a1630_5875 , \48617_nG17248 , \47166 );
_HMUX g1724a ( \48619_nG1724a , RIe3a1630_5875 , \47708 , \48205 );
_HMUX g1724b ( \48620_nG1724b , \48618_nG17249 , \48619_nG1724a , \47178 );
buf \U$38931 ( \48621 , \48620_nG1724b );
_DC g18f71_GF_IsGateDCbyConstraint ( \48622_nG18f71 , \48621 , \42503 );
buf \U$38932 ( \48623 , \48622_nG18f71 );
_HMUX g1724c ( \48624_nG1724c , RIe3a1e28_5876 , \47714 , \48202 );
_HMUX g1724d ( \48625_nG1724d , RIe3a1e28_5876 , \48624_nG1724c , \47166 );
_HMUX g1724e ( \48626_nG1724e , RIe3a1e28_5876 , \47717 , \48205 );
_HMUX g1724f ( \48627_nG1724f , \48625_nG1724d , \48626_nG1724e , \47178 );
buf \U$38933 ( \48628 , \48627_nG1724f );
_DC g18f73_GF_IsGateDCbyConstraint ( \48629_nG18f73 , \48628 , \42503 );
buf \U$38934 ( \48630 , \48629_nG18f73 );
_HMUX g17250 ( \48631_nG17250 , RIe3a2620_5877 , \47723 , \48202 );
_HMUX g17251 ( \48632_nG17251 , RIe3a2620_5877 , \48631_nG17250 , \47166 );
_HMUX g17252 ( \48633_nG17252 , RIe3a2620_5877 , \47726 , \48205 );
_HMUX g17253 ( \48634_nG17253 , \48632_nG17251 , \48633_nG17252 , \47178 );
buf \U$38935 ( \48635 , \48634_nG17253 );
_DC g18f75_GF_IsGateDCbyConstraint ( \48636_nG18f75 , \48635 , \42503 );
buf \U$38936 ( \48637 , \48636_nG18f75 );
_HMUX g17254 ( \48638_nG17254 , RIe3a2e18_5878 , \47732 , \48202 );
_HMUX g17255 ( \48639_nG17255 , RIe3a2e18_5878 , \48638_nG17254 , \47166 );
_HMUX g17256 ( \48640_nG17256 , RIe3a2e18_5878 , \47735 , \48205 );
_HMUX g17257 ( \48641_nG17257 , \48639_nG17255 , \48640_nG17256 , \47178 );
buf \U$38937 ( \48642 , \48641_nG17257 );
_DC g18f77_GF_IsGateDCbyConstraint ( \48643_nG18f77 , \48642 , \42503 );
buf \U$38938 ( \48644 , \48643_nG18f77 );
_HMUX g17258 ( \48645_nG17258 , RIe3a3610_5879 , \47741 , \48202 );
_HMUX g17259 ( \48646_nG17259 , RIe3a3610_5879 , \48645_nG17258 , \47166 );
_HMUX g1725a ( \48647_nG1725a , RIe3a3610_5879 , \47744 , \48205 );
_HMUX g1725b ( \48648_nG1725b , \48646_nG17259 , \48647_nG1725a , \47178 );
buf \U$38939 ( \48649 , \48648_nG1725b );
_DC g18f79_GF_IsGateDCbyConstraint ( \48650_nG18f79 , \48649 , \42503 );
buf \U$38940 ( \48651 , \48650_nG18f79 );
and \U$38941 ( \48652 , \47156 , \47157 );
_HMUX g16fd8 ( \48653_nG16fd8 , RIe3a3e08_5880 , \47155 , \48652 );
_HMUX g16fd9 ( \48654_nG16fd9 , RIe3a3e08_5880 , \48653_nG16fd8 , \47166 );
and \U$38942 ( \48655 , \47169 , \47170 );
_HMUX g16fde ( \48656_nG16fde , RIe3a3e08_5880 , \47168 , \48655 );
_HMUX g16fdf ( \48657_nG16fdf , \48654_nG16fd9 , \48656_nG16fde , \47178 );
buf \U$38943 ( \48658 , \48657_nG16fdf );
_DC g18e81_GF_IsGateDCbyConstraint ( \48659_nG18e81 , \48658 , \42503 );
buf \U$38944 ( \48660 , \48659_nG18e81 );
_HMUX g16fe1 ( \48661_nG16fe1 , RIe3a4600_5881 , \47183 , \48652 );
_HMUX g16fe2 ( \48662_nG16fe2 , RIe3a4600_5881 , \48661_nG16fe1 , \47166 );
_HMUX g16fe4 ( \48663_nG16fe4 , RIe3a4600_5881 , \47186 , \48655 );
_HMUX g16fe5 ( \48664_nG16fe5 , \48662_nG16fe2 , \48663_nG16fe4 , \47178 );
buf \U$38945 ( \48665 , \48664_nG16fe5 );
_DC g18e97_GF_IsGateDCbyConstraint ( \48666_nG18e97 , \48665 , \42503 );
buf \U$38946 ( \48667 , \48666_nG18e97 );
_HMUX g16fe7 ( \48668_nG16fe7 , RIe3a4df8_5882 , \47192 , \48652 );
_HMUX g16fe8 ( \48669_nG16fe8 , RIe3a4df8_5882 , \48668_nG16fe7 , \47166 );
_HMUX g16fea ( \48670_nG16fea , RIe3a4df8_5882 , \47195 , \48655 );
_HMUX g16feb ( \48671_nG16feb , \48669_nG16fe8 , \48670_nG16fea , \47178 );
buf \U$38947 ( \48672 , \48671_nG16feb );
_DC g18ead_GF_IsGateDCbyConstraint ( \48673_nG18ead , \48672 , \42503 );
buf \U$38948 ( \48674 , \48673_nG18ead );
_HMUX g16fed ( \48675_nG16fed , RIe3a55f0_5883 , \47201 , \48652 );
_HMUX g16fee ( \48676_nG16fee , RIe3a55f0_5883 , \48675_nG16fed , \47166 );
_HMUX g16ff0 ( \48677_nG16ff0 , RIe3a55f0_5883 , \47204 , \48655 );
_HMUX g16ff1 ( \48678_nG16ff1 , \48676_nG16fee , \48677_nG16ff0 , \47178 );
buf \U$38949 ( \48679 , \48678_nG16ff1 );
_DC g18ec3_GF_IsGateDCbyConstraint ( \48680_nG18ec3 , \48679 , \42503 );
buf \U$38950 ( \48681 , \48680_nG18ec3 );
_HMUX g16ff3 ( \48682_nG16ff3 , RIe3a5de8_5884 , \47210 , \48652 );
_HMUX g16ff4 ( \48683_nG16ff4 , RIe3a5de8_5884 , \48682_nG16ff3 , \47166 );
_HMUX g16ff6 ( \48684_nG16ff6 , RIe3a5de8_5884 , \47213 , \48655 );
_HMUX g16ff7 ( \48685_nG16ff7 , \48683_nG16ff4 , \48684_nG16ff6 , \47178 );
buf \U$38951 ( \48686 , \48685_nG16ff7 );
_DC g18ed9_GF_IsGateDCbyConstraint ( \48687_nG18ed9 , \48686 , \42503 );
buf \U$38952 ( \48688 , \48687_nG18ed9 );
_HMUX g16ff9 ( \48689_nG16ff9 , RIe3a65e0_5885 , \47219 , \48652 );
_HMUX g16ffa ( \48690_nG16ffa , RIe3a65e0_5885 , \48689_nG16ff9 , \47166 );
_HMUX g16ffc ( \48691_nG16ffc , RIe3a65e0_5885 , \47222 , \48655 );
_HMUX g16ffd ( \48692_nG16ffd , \48690_nG16ffa , \48691_nG16ffc , \47178 );
buf \U$38953 ( \48693 , \48692_nG16ffd );
_DC g18eef_GF_IsGateDCbyConstraint ( \48694_nG18eef , \48693 , \42503 );
buf \U$38954 ( \48695 , \48694_nG18eef );
_HMUX g16fff ( \48696_nG16fff , RIe3a6dd8_5886 , \47228 , \48652 );
_HMUX g17000 ( \48697_nG17000 , RIe3a6dd8_5886 , \48696_nG16fff , \47166 );
_HMUX g17002 ( \48698_nG17002 , RIe3a6dd8_5886 , \47231 , \48655 );
_HMUX g17003 ( \48699_nG17003 , \48697_nG17000 , \48698_nG17002 , \47178 );
buf \U$38955 ( \48700 , \48699_nG17003 );
_DC g18efb_GF_IsGateDCbyConstraint ( \48701_nG18efb , \48700 , \42503 );
buf \U$38956 ( \48702 , \48701_nG18efb );
_HMUX g17005 ( \48703_nG17005 , RIe3a75d0_5887 , \47237 , \48652 );
_HMUX g17006 ( \48704_nG17006 , RIe3a75d0_5887 , \48703_nG17005 , \47166 );
_HMUX g17008 ( \48705_nG17008 , RIe3a75d0_5887 , \47240 , \48655 );
_HMUX g17009 ( \48706_nG17009 , \48704_nG17006 , \48705_nG17008 , \47178 );
buf \U$38957 ( \48707 , \48706_nG17009 );
_DC g18efd_GF_IsGateDCbyConstraint ( \48708_nG18efd , \48707 , \42503 );
buf \U$38958 ( \48709 , \48708_nG18efd );
_HMUX g1700b ( \48710_nG1700b , RIe3a7dc8_5888 , \47246 , \48652 );
_HMUX g1700c ( \48711_nG1700c , RIe3a7dc8_5888 , \48710_nG1700b , \47166 );
_HMUX g1700e ( \48712_nG1700e , RIe3a7dc8_5888 , \47249 , \48655 );
_HMUX g1700f ( \48713_nG1700f , \48711_nG1700c , \48712_nG1700e , \47178 );
buf \U$38959 ( \48714 , \48713_nG1700f );
_DC g18eff_GF_IsGateDCbyConstraint ( \48715_nG18eff , \48714 , \42503 );
buf \U$38960 ( \48716 , \48715_nG18eff );
_HMUX g17011 ( \48717_nG17011 , RIe3a85c0_5889 , \47255 , \48652 );
_HMUX g17012 ( \48718_nG17012 , RIe3a85c0_5889 , \48717_nG17011 , \47166 );
_HMUX g17014 ( \48719_nG17014 , RIe3a85c0_5889 , \47258 , \48655 );
_HMUX g17015 ( \48720_nG17015 , \48718_nG17012 , \48719_nG17014 , \47178 );
buf \U$38961 ( \48721 , \48720_nG17015 );
_DC g18e83_GF_IsGateDCbyConstraint ( \48722_nG18e83 , \48721 , \42503 );
buf \U$38962 ( \48723 , \48722_nG18e83 );
_HMUX g17017 ( \48724_nG17017 , RIe3a8db8_5890 , \47264 , \48652 );
_HMUX g17018 ( \48725_nG17018 , RIe3a8db8_5890 , \48724_nG17017 , \47166 );
_HMUX g1701a ( \48726_nG1701a , RIe3a8db8_5890 , \47267 , \48655 );
_HMUX g1701b ( \48727_nG1701b , \48725_nG17018 , \48726_nG1701a , \47178 );
buf \U$38963 ( \48728 , \48727_nG1701b );
_DC g18e85_GF_IsGateDCbyConstraint ( \48729_nG18e85 , \48728 , \42503 );
buf \U$38964 ( \48730 , \48729_nG18e85 );
_HMUX g1701d ( \48731_nG1701d , RIe3a95b0_5891 , \47273 , \48652 );
_HMUX g1701e ( \48732_nG1701e , RIe3a95b0_5891 , \48731_nG1701d , \47166 );
_HMUX g17020 ( \48733_nG17020 , RIe3a95b0_5891 , \47276 , \48655 );
_HMUX g17021 ( \48734_nG17021 , \48732_nG1701e , \48733_nG17020 , \47178 );
buf \U$38965 ( \48735 , \48734_nG17021 );
_DC g18e87_GF_IsGateDCbyConstraint ( \48736_nG18e87 , \48735 , \42503 );
buf \U$38966 ( \48737 , \48736_nG18e87 );
_HMUX g17023 ( \48738_nG17023 , RIe3a9da8_5892 , \47282 , \48652 );
_HMUX g17024 ( \48739_nG17024 , RIe3a9da8_5892 , \48738_nG17023 , \47166 );
_HMUX g17026 ( \48740_nG17026 , RIe3a9da8_5892 , \47285 , \48655 );
_HMUX g17027 ( \48741_nG17027 , \48739_nG17024 , \48740_nG17026 , \47178 );
buf \U$38967 ( \48742 , \48741_nG17027 );
_DC g18e89_GF_IsGateDCbyConstraint ( \48743_nG18e89 , \48742 , \42503 );
buf \U$38968 ( \48744 , \48743_nG18e89 );
_HMUX g17029 ( \48745_nG17029 , RIe3aa5a0_5893 , \47291 , \48652 );
_HMUX g1702a ( \48746_nG1702a , RIe3aa5a0_5893 , \48745_nG17029 , \47166 );
_HMUX g1702c ( \48747_nG1702c , RIe3aa5a0_5893 , \47294 , \48655 );
_HMUX g1702d ( \48748_nG1702d , \48746_nG1702a , \48747_nG1702c , \47178 );
buf \U$38969 ( \48749 , \48748_nG1702d );
_DC g18e8b_GF_IsGateDCbyConstraint ( \48750_nG18e8b , \48749 , \42503 );
buf \U$38970 ( \48751 , \48750_nG18e8b );
_HMUX g1702f ( \48752_nG1702f , RIe3aad98_5894 , \47300 , \48652 );
_HMUX g17030 ( \48753_nG17030 , RIe3aad98_5894 , \48752_nG1702f , \47166 );
_HMUX g17032 ( \48754_nG17032 , RIe3aad98_5894 , \47303 , \48655 );
_HMUX g17033 ( \48755_nG17033 , \48753_nG17030 , \48754_nG17032 , \47178 );
buf \U$38971 ( \48756 , \48755_nG17033 );
_DC g18e8d_GF_IsGateDCbyConstraint ( \48757_nG18e8d , \48756 , \42503 );
buf \U$38972 ( \48758 , \48757_nG18e8d );
_HMUX g17035 ( \48759_nG17035 , RIe3ab590_5895 , \47309 , \48652 );
_HMUX g17036 ( \48760_nG17036 , RIe3ab590_5895 , \48759_nG17035 , \47166 );
_HMUX g17038 ( \48761_nG17038 , RIe3ab590_5895 , \47312 , \48655 );
_HMUX g17039 ( \48762_nG17039 , \48760_nG17036 , \48761_nG17038 , \47178 );
buf \U$38973 ( \48763 , \48762_nG17039 );
_DC g18e8f_GF_IsGateDCbyConstraint ( \48764_nG18e8f , \48763 , \42503 );
buf \U$38974 ( \48765 , \48764_nG18e8f );
_HMUX g1703b ( \48766_nG1703b , RIe3abd88_5896 , \47318 , \48652 );
_HMUX g1703c ( \48767_nG1703c , RIe3abd88_5896 , \48766_nG1703b , \47166 );
_HMUX g1703e ( \48768_nG1703e , RIe3abd88_5896 , \47321 , \48655 );
_HMUX g1703f ( \48769_nG1703f , \48767_nG1703c , \48768_nG1703e , \47178 );
buf \U$38975 ( \48770 , \48769_nG1703f );
_DC g18e91_GF_IsGateDCbyConstraint ( \48771_nG18e91 , \48770 , \42503 );
buf \U$38976 ( \48772 , \48771_nG18e91 );
_HMUX g17041 ( \48773_nG17041 , RIe3ac580_5897 , \47327 , \48652 );
_HMUX g17042 ( \48774_nG17042 , RIe3ac580_5897 , \48773_nG17041 , \47166 );
_HMUX g17044 ( \48775_nG17044 , RIe3ac580_5897 , \47330 , \48655 );
_HMUX g17045 ( \48776_nG17045 , \48774_nG17042 , \48775_nG17044 , \47178 );
buf \U$38977 ( \48777 , \48776_nG17045 );
_DC g18e93_GF_IsGateDCbyConstraint ( \48778_nG18e93 , \48777 , \42503 );
buf \U$38978 ( \48779 , \48778_nG18e93 );
_HMUX g17047 ( \48780_nG17047 , RIe3acd78_5898 , \47336 , \48652 );
_HMUX g17048 ( \48781_nG17048 , RIe3acd78_5898 , \48780_nG17047 , \47166 );
_HMUX g1704a ( \48782_nG1704a , RIe3acd78_5898 , \47339 , \48655 );
_HMUX g1704b ( \48783_nG1704b , \48781_nG17048 , \48782_nG1704a , \47178 );
buf \U$38979 ( \48784 , \48783_nG1704b );
_DC g18e95_GF_IsGateDCbyConstraint ( \48785_nG18e95 , \48784 , \42503 );
buf \U$38980 ( \48786 , \48785_nG18e95 );
_HMUX g1704d ( \48787_nG1704d , RIe3ad570_5899 , \47345 , \48652 );
_HMUX g1704e ( \48788_nG1704e , RIe3ad570_5899 , \48787_nG1704d , \47166 );
_HMUX g17050 ( \48789_nG17050 , RIe3ad570_5899 , \47348 , \48655 );
_HMUX g17051 ( \48790_nG17051 , \48788_nG1704e , \48789_nG17050 , \47178 );
buf \U$38981 ( \48791 , \48790_nG17051 );
_DC g18e99_GF_IsGateDCbyConstraint ( \48792_nG18e99 , \48791 , \42503 );
buf \U$38982 ( \48793 , \48792_nG18e99 );
_HMUX g17053 ( \48794_nG17053 , RIe3add68_5900 , \47354 , \48652 );
_HMUX g17054 ( \48795_nG17054 , RIe3add68_5900 , \48794_nG17053 , \47166 );
_HMUX g17056 ( \48796_nG17056 , RIe3add68_5900 , \47357 , \48655 );
_HMUX g17057 ( \48797_nG17057 , \48795_nG17054 , \48796_nG17056 , \47178 );
buf \U$38983 ( \48798 , \48797_nG17057 );
_DC g18e9b_GF_IsGateDCbyConstraint ( \48799_nG18e9b , \48798 , \42503 );
buf \U$38984 ( \48800 , \48799_nG18e9b );
_HMUX g17059 ( \48801_nG17059 , RIe3ae560_5901 , \47363 , \48652 );
_HMUX g1705a ( \48802_nG1705a , RIe3ae560_5901 , \48801_nG17059 , \47166 );
_HMUX g1705c ( \48803_nG1705c , RIe3ae560_5901 , \47366 , \48655 );
_HMUX g1705d ( \48804_nG1705d , \48802_nG1705a , \48803_nG1705c , \47178 );
buf \U$38985 ( \48805 , \48804_nG1705d );
_DC g18e9d_GF_IsGateDCbyConstraint ( \48806_nG18e9d , \48805 , \42503 );
buf \U$38986 ( \48807 , \48806_nG18e9d );
_HMUX g1705f ( \48808_nG1705f , RIe3aed58_5902 , \47372 , \48652 );
_HMUX g17060 ( \48809_nG17060 , RIe3aed58_5902 , \48808_nG1705f , \47166 );
_HMUX g17062 ( \48810_nG17062 , RIe3aed58_5902 , \47375 , \48655 );
_HMUX g17063 ( \48811_nG17063 , \48809_nG17060 , \48810_nG17062 , \47178 );
buf \U$38987 ( \48812 , \48811_nG17063 );
_DC g18e9f_GF_IsGateDCbyConstraint ( \48813_nG18e9f , \48812 , \42503 );
buf \U$38988 ( \48814 , \48813_nG18e9f );
_HMUX g17065 ( \48815_nG17065 , RIe3af550_5903 , \47381 , \48652 );
_HMUX g17066 ( \48816_nG17066 , RIe3af550_5903 , \48815_nG17065 , \47166 );
_HMUX g17068 ( \48817_nG17068 , RIe3af550_5903 , \47384 , \48655 );
_HMUX g17069 ( \48818_nG17069 , \48816_nG17066 , \48817_nG17068 , \47178 );
buf \U$38989 ( \48819 , \48818_nG17069 );
_DC g18ea1_GF_IsGateDCbyConstraint ( \48820_nG18ea1 , \48819 , \42503 );
buf \U$38990 ( \48821 , \48820_nG18ea1 );
_HMUX g1706b ( \48822_nG1706b , RIe3afd48_5904 , \47390 , \48652 );
_HMUX g1706c ( \48823_nG1706c , RIe3afd48_5904 , \48822_nG1706b , \47166 );
_HMUX g1706e ( \48824_nG1706e , RIe3afd48_5904 , \47393 , \48655 );
_HMUX g1706f ( \48825_nG1706f , \48823_nG1706c , \48824_nG1706e , \47178 );
buf \U$38991 ( \48826 , \48825_nG1706f );
_DC g18ea3_GF_IsGateDCbyConstraint ( \48827_nG18ea3 , \48826 , \42503 );
buf \U$38992 ( \48828 , \48827_nG18ea3 );
_HMUX g17071 ( \48829_nG17071 , RIe3b0540_5905 , \47399 , \48652 );
_HMUX g17072 ( \48830_nG17072 , RIe3b0540_5905 , \48829_nG17071 , \47166 );
_HMUX g17074 ( \48831_nG17074 , RIe3b0540_5905 , \47402 , \48655 );
_HMUX g17075 ( \48832_nG17075 , \48830_nG17072 , \48831_nG17074 , \47178 );
buf \U$38993 ( \48833 , \48832_nG17075 );
_DC g18ea5_GF_IsGateDCbyConstraint ( \48834_nG18ea5 , \48833 , \42503 );
buf \U$38994 ( \48835 , \48834_nG18ea5 );
_HMUX g17077 ( \48836_nG17077 , RIe3b0d38_5906 , \47408 , \48652 );
_HMUX g17078 ( \48837_nG17078 , RIe3b0d38_5906 , \48836_nG17077 , \47166 );
_HMUX g1707a ( \48838_nG1707a , RIe3b0d38_5906 , \47411 , \48655 );
_HMUX g1707b ( \48839_nG1707b , \48837_nG17078 , \48838_nG1707a , \47178 );
buf \U$38995 ( \48840 , \48839_nG1707b );
_DC g18ea7_GF_IsGateDCbyConstraint ( \48841_nG18ea7 , \48840 , \42503 );
buf \U$38996 ( \48842 , \48841_nG18ea7 );
_HMUX g1707d ( \48843_nG1707d , RIe3b1530_5907 , \47417 , \48652 );
_HMUX g1707e ( \48844_nG1707e , RIe3b1530_5907 , \48843_nG1707d , \47166 );
_HMUX g17080 ( \48845_nG17080 , RIe3b1530_5907 , \47420 , \48655 );
_HMUX g17081 ( \48846_nG17081 , \48844_nG1707e , \48845_nG17080 , \47178 );
buf \U$38997 ( \48847 , \48846_nG17081 );
_DC g18ea9_GF_IsGateDCbyConstraint ( \48848_nG18ea9 , \48847 , \42503 );
buf \U$38998 ( \48849 , \48848_nG18ea9 );
_HMUX g17083 ( \48850_nG17083 , RIe3b1d28_5908 , \47426 , \48652 );
_HMUX g17084 ( \48851_nG17084 , RIe3b1d28_5908 , \48850_nG17083 , \47166 );
_HMUX g17086 ( \48852_nG17086 , RIe3b1d28_5908 , \47429 , \48655 );
_HMUX g17087 ( \48853_nG17087 , \48851_nG17084 , \48852_nG17086 , \47178 );
buf \U$38999 ( \48854 , \48853_nG17087 );
_DC g18eab_GF_IsGateDCbyConstraint ( \48855_nG18eab , \48854 , \42503 );
buf \U$39000 ( \48856 , \48855_nG18eab );
_HMUX g17089 ( \48857_nG17089 , RIe3b2520_5909 , \47435 , \48652 );
_HMUX g1708a ( \48858_nG1708a , RIe3b2520_5909 , \48857_nG17089 , \47166 );
_HMUX g1708c ( \48859_nG1708c , RIe3b2520_5909 , \47438 , \48655 );
_HMUX g1708d ( \48860_nG1708d , \48858_nG1708a , \48859_nG1708c , \47178 );
buf \U$39001 ( \48861 , \48860_nG1708d );
_DC g18eaf_GF_IsGateDCbyConstraint ( \48862_nG18eaf , \48861 , \42503 );
buf \U$39002 ( \48863 , \48862_nG18eaf );
_HMUX g1708f ( \48864_nG1708f , RIe3b2d18_5910 , \47444 , \48652 );
_HMUX g17090 ( \48865_nG17090 , RIe3b2d18_5910 , \48864_nG1708f , \47166 );
_HMUX g17092 ( \48866_nG17092 , RIe3b2d18_5910 , \47447 , \48655 );
_HMUX g17093 ( \48867_nG17093 , \48865_nG17090 , \48866_nG17092 , \47178 );
buf \U$39003 ( \48868 , \48867_nG17093 );
_DC g18eb1_GF_IsGateDCbyConstraint ( \48869_nG18eb1 , \48868 , \42503 );
buf \U$39004 ( \48870 , \48869_nG18eb1 );
_HMUX g17095 ( \48871_nG17095 , RIe3b3510_5911 , \47453 , \48652 );
_HMUX g17096 ( \48872_nG17096 , RIe3b3510_5911 , \48871_nG17095 , \47166 );
_HMUX g17098 ( \48873_nG17098 , RIe3b3510_5911 , \47456 , \48655 );
_HMUX g17099 ( \48874_nG17099 , \48872_nG17096 , \48873_nG17098 , \47178 );
buf \U$39005 ( \48875 , \48874_nG17099 );
_DC g18eb3_GF_IsGateDCbyConstraint ( \48876_nG18eb3 , \48875 , \42503 );
buf \U$39006 ( \48877 , \48876_nG18eb3 );
_HMUX g1709b ( \48878_nG1709b , RIe3b3d08_5912 , \47462 , \48652 );
_HMUX g1709c ( \48879_nG1709c , RIe3b3d08_5912 , \48878_nG1709b , \47166 );
_HMUX g1709e ( \48880_nG1709e , RIe3b3d08_5912 , \47465 , \48655 );
_HMUX g1709f ( \48881_nG1709f , \48879_nG1709c , \48880_nG1709e , \47178 );
buf \U$39007 ( \48882 , \48881_nG1709f );
_DC g18eb5_GF_IsGateDCbyConstraint ( \48883_nG18eb5 , \48882 , \42503 );
buf \U$39008 ( \48884 , \48883_nG18eb5 );
_HMUX g170a1 ( \48885_nG170a1 , RIe3b4500_5913 , \47471 , \48652 );
_HMUX g170a2 ( \48886_nG170a2 , RIe3b4500_5913 , \48885_nG170a1 , \47166 );
_HMUX g170a4 ( \48887_nG170a4 , RIe3b4500_5913 , \47474 , \48655 );
_HMUX g170a5 ( \48888_nG170a5 , \48886_nG170a2 , \48887_nG170a4 , \47178 );
buf \U$39009 ( \48889 , \48888_nG170a5 );
_DC g18eb7_GF_IsGateDCbyConstraint ( \48890_nG18eb7 , \48889 , \42503 );
buf \U$39010 ( \48891 , \48890_nG18eb7 );
_HMUX g170a7 ( \48892_nG170a7 , RIe3b4cf8_5914 , \47480 , \48652 );
_HMUX g170a8 ( \48893_nG170a8 , RIe3b4cf8_5914 , \48892_nG170a7 , \47166 );
_HMUX g170aa ( \48894_nG170aa , RIe3b4cf8_5914 , \47483 , \48655 );
_HMUX g170ab ( \48895_nG170ab , \48893_nG170a8 , \48894_nG170aa , \47178 );
buf \U$39011 ( \48896 , \48895_nG170ab );
_DC g18eb9_GF_IsGateDCbyConstraint ( \48897_nG18eb9 , \48896 , \42503 );
buf \U$39012 ( \48898 , \48897_nG18eb9 );
_HMUX g170ad ( \48899_nG170ad , RIe3b54f0_5915 , \47489 , \48652 );
_HMUX g170ae ( \48900_nG170ae , RIe3b54f0_5915 , \48899_nG170ad , \47166 );
_HMUX g170b0 ( \48901_nG170b0 , RIe3b54f0_5915 , \47492 , \48655 );
_HMUX g170b1 ( \48902_nG170b1 , \48900_nG170ae , \48901_nG170b0 , \47178 );
buf \U$39013 ( \48903 , \48902_nG170b1 );
_DC g18ebb_GF_IsGateDCbyConstraint ( \48904_nG18ebb , \48903 , \42503 );
buf \U$39014 ( \48905 , \48904_nG18ebb );
_HMUX g170b3 ( \48906_nG170b3 , RIe3b5ce8_5916 , \47498 , \48652 );
_HMUX g170b4 ( \48907_nG170b4 , RIe3b5ce8_5916 , \48906_nG170b3 , \47166 );
_HMUX g170b6 ( \48908_nG170b6 , RIe3b5ce8_5916 , \47501 , \48655 );
_HMUX g170b7 ( \48909_nG170b7 , \48907_nG170b4 , \48908_nG170b6 , \47178 );
buf \U$39015 ( \48910 , \48909_nG170b7 );
_DC g18ebd_GF_IsGateDCbyConstraint ( \48911_nG18ebd , \48910 , \42503 );
buf \U$39016 ( \48912 , \48911_nG18ebd );
_HMUX g170b9 ( \48913_nG170b9 , RIe3b64e0_5917 , \47507 , \48652 );
_HMUX g170ba ( \48914_nG170ba , RIe3b64e0_5917 , \48913_nG170b9 , \47166 );
_HMUX g170bc ( \48915_nG170bc , RIe3b64e0_5917 , \47510 , \48655 );
_HMUX g170bd ( \48916_nG170bd , \48914_nG170ba , \48915_nG170bc , \47178 );
buf \U$39017 ( \48917 , \48916_nG170bd );
_DC g18ebf_GF_IsGateDCbyConstraint ( \48918_nG18ebf , \48917 , \42503 );
buf \U$39018 ( \48919 , \48918_nG18ebf );
_HMUX g170bf ( \48920_nG170bf , RIe3b6cd8_5918 , \47516 , \48652 );
_HMUX g170c0 ( \48921_nG170c0 , RIe3b6cd8_5918 , \48920_nG170bf , \47166 );
_HMUX g170c2 ( \48922_nG170c2 , RIe3b6cd8_5918 , \47519 , \48655 );
_HMUX g170c3 ( \48923_nG170c3 , \48921_nG170c0 , \48922_nG170c2 , \47178 );
buf \U$39019 ( \48924 , \48923_nG170c3 );
_DC g18ec1_GF_IsGateDCbyConstraint ( \48925_nG18ec1 , \48924 , \42503 );
buf \U$39020 ( \48926 , \48925_nG18ec1 );
_HMUX g170c5 ( \48927_nG170c5 , RIe3b74d0_5919 , \47525 , \48652 );
_HMUX g170c6 ( \48928_nG170c6 , RIe3b74d0_5919 , \48927_nG170c5 , \47166 );
_HMUX g170c8 ( \48929_nG170c8 , RIe3b74d0_5919 , \47528 , \48655 );
_HMUX g170c9 ( \48930_nG170c9 , \48928_nG170c6 , \48929_nG170c8 , \47178 );
buf \U$39021 ( \48931 , \48930_nG170c9 );
_DC g18ec5_GF_IsGateDCbyConstraint ( \48932_nG18ec5 , \48931 , \42503 );
buf \U$39022 ( \48933 , \48932_nG18ec5 );
_HMUX g170cb ( \48934_nG170cb , RIe3b7cc8_5920 , \47534 , \48652 );
_HMUX g170cc ( \48935_nG170cc , RIe3b7cc8_5920 , \48934_nG170cb , \47166 );
_HMUX g170ce ( \48936_nG170ce , RIe3b7cc8_5920 , \47537 , \48655 );
_HMUX g170cf ( \48937_nG170cf , \48935_nG170cc , \48936_nG170ce , \47178 );
buf \U$39023 ( \48938 , \48937_nG170cf );
_DC g18ec7_GF_IsGateDCbyConstraint ( \48939_nG18ec7 , \48938 , \42503 );
buf \U$39024 ( \48940 , \48939_nG18ec7 );
_HMUX g170d1 ( \48941_nG170d1 , RIe3b84c0_5921 , \47543 , \48652 );
_HMUX g170d2 ( \48942_nG170d2 , RIe3b84c0_5921 , \48941_nG170d1 , \47166 );
_HMUX g170d4 ( \48943_nG170d4 , RIe3b84c0_5921 , \47546 , \48655 );
_HMUX g170d5 ( \48944_nG170d5 , \48942_nG170d2 , \48943_nG170d4 , \47178 );
buf \U$39025 ( \48945 , \48944_nG170d5 );
_DC g18ec9_GF_IsGateDCbyConstraint ( \48946_nG18ec9 , \48945 , \42503 );
buf \U$39026 ( \48947 , \48946_nG18ec9 );
_HMUX g170d7 ( \48948_nG170d7 , RIe3b8cb8_5922 , \47552 , \48652 );
_HMUX g170d8 ( \48949_nG170d8 , RIe3b8cb8_5922 , \48948_nG170d7 , \47166 );
_HMUX g170da ( \48950_nG170da , RIe3b8cb8_5922 , \47555 , \48655 );
_HMUX g170db ( \48951_nG170db , \48949_nG170d8 , \48950_nG170da , \47178 );
buf \U$39027 ( \48952 , \48951_nG170db );
_DC g18ecb_GF_IsGateDCbyConstraint ( \48953_nG18ecb , \48952 , \42503 );
buf \U$39028 ( \48954 , \48953_nG18ecb );
_HMUX g170dd ( \48955_nG170dd , RIe3b94b0_5923 , \47561 , \48652 );
_HMUX g170de ( \48956_nG170de , RIe3b94b0_5923 , \48955_nG170dd , \47166 );
_HMUX g170e0 ( \48957_nG170e0 , RIe3b94b0_5923 , \47564 , \48655 );
_HMUX g170e1 ( \48958_nG170e1 , \48956_nG170de , \48957_nG170e0 , \47178 );
buf \U$39029 ( \48959 , \48958_nG170e1 );
_DC g18ecd_GF_IsGateDCbyConstraint ( \48960_nG18ecd , \48959 , \42503 );
buf \U$39030 ( \48961 , \48960_nG18ecd );
_HMUX g170e3 ( \48962_nG170e3 , RIe3b9ca8_5924 , \47570 , \48652 );
_HMUX g170e4 ( \48963_nG170e4 , RIe3b9ca8_5924 , \48962_nG170e3 , \47166 );
_HMUX g170e6 ( \48964_nG170e6 , RIe3b9ca8_5924 , \47573 , \48655 );
_HMUX g170e7 ( \48965_nG170e7 , \48963_nG170e4 , \48964_nG170e6 , \47178 );
buf \U$39031 ( \48966 , \48965_nG170e7 );
_DC g18ecf_GF_IsGateDCbyConstraint ( \48967_nG18ecf , \48966 , \42503 );
buf \U$39032 ( \48968 , \48967_nG18ecf );
_HMUX g170e9 ( \48969_nG170e9 , RIe3ba4a0_5925 , \47579 , \48652 );
_HMUX g170ea ( \48970_nG170ea , RIe3ba4a0_5925 , \48969_nG170e9 , \47166 );
_HMUX g170ec ( \48971_nG170ec , RIe3ba4a0_5925 , \47582 , \48655 );
_HMUX g170ed ( \48972_nG170ed , \48970_nG170ea , \48971_nG170ec , \47178 );
buf \U$39033 ( \48973 , \48972_nG170ed );
_DC g18ed1_GF_IsGateDCbyConstraint ( \48974_nG18ed1 , \48973 , \42503 );
buf \U$39034 ( \48975 , \48974_nG18ed1 );
_HMUX g170ef ( \48976_nG170ef , RIe3bac98_5926 , \47588 , \48652 );
_HMUX g170f0 ( \48977_nG170f0 , RIe3bac98_5926 , \48976_nG170ef , \47166 );
_HMUX g170f2 ( \48978_nG170f2 , RIe3bac98_5926 , \47591 , \48655 );
_HMUX g170f3 ( \48979_nG170f3 , \48977_nG170f0 , \48978_nG170f2 , \47178 );
buf \U$39035 ( \48980 , \48979_nG170f3 );
_DC g18ed3_GF_IsGateDCbyConstraint ( \48981_nG18ed3 , \48980 , \42503 );
buf \U$39036 ( \48982 , \48981_nG18ed3 );
_HMUX g170f5 ( \48983_nG170f5 , RIe3bb490_5927 , \47597 , \48652 );
_HMUX g170f6 ( \48984_nG170f6 , RIe3bb490_5927 , \48983_nG170f5 , \47166 );
_HMUX g170f8 ( \48985_nG170f8 , RIe3bb490_5927 , \47600 , \48655 );
_HMUX g170f9 ( \48986_nG170f9 , \48984_nG170f6 , \48985_nG170f8 , \47178 );
buf \U$39037 ( \48987 , \48986_nG170f9 );
_DC g18ed5_GF_IsGateDCbyConstraint ( \48988_nG18ed5 , \48987 , \42503 );
buf \U$39038 ( \48989 , \48988_nG18ed5 );
_HMUX g170fb ( \48990_nG170fb , RIe3bbc88_5928 , \47606 , \48652 );
_HMUX g170fc ( \48991_nG170fc , RIe3bbc88_5928 , \48990_nG170fb , \47166 );
_HMUX g170fe ( \48992_nG170fe , RIe3bbc88_5928 , \47609 , \48655 );
_HMUX g170ff ( \48993_nG170ff , \48991_nG170fc , \48992_nG170fe , \47178 );
buf \U$39039 ( \48994 , \48993_nG170ff );
_DC g18ed7_GF_IsGateDCbyConstraint ( \48995_nG18ed7 , \48994 , \42503 );
buf \U$39040 ( \48996 , \48995_nG18ed7 );
_HMUX g17101 ( \48997_nG17101 , RIe3bc480_5929 , \47615 , \48652 );
_HMUX g17102 ( \48998_nG17102 , RIe3bc480_5929 , \48997_nG17101 , \47166 );
_HMUX g17104 ( \48999_nG17104 , RIe3bc480_5929 , \47618 , \48655 );
_HMUX g17105 ( \49000_nG17105 , \48998_nG17102 , \48999_nG17104 , \47178 );
buf \U$39041 ( \49001 , \49000_nG17105 );
_DC g18edb_GF_IsGateDCbyConstraint ( \49002_nG18edb , \49001 , \42503 );
buf \U$39042 ( \49003 , \49002_nG18edb );
_HMUX g17107 ( \49004_nG17107 , RIe3bcc78_5930 , \47624 , \48652 );
_HMUX g17108 ( \49005_nG17108 , RIe3bcc78_5930 , \49004_nG17107 , \47166 );
_HMUX g1710a ( \49006_nG1710a , RIe3bcc78_5930 , \47627 , \48655 );
_HMUX g1710b ( \49007_nG1710b , \49005_nG17108 , \49006_nG1710a , \47178 );
buf \U$39043 ( \49008 , \49007_nG1710b );
_DC g18edd_GF_IsGateDCbyConstraint ( \49009_nG18edd , \49008 , \42503 );
buf \U$39044 ( \49010 , \49009_nG18edd );
_HMUX g1710d ( \49011_nG1710d , RIe3bd470_5931 , \47633 , \48652 );
_HMUX g1710e ( \49012_nG1710e , RIe3bd470_5931 , \49011_nG1710d , \47166 );
_HMUX g17110 ( \49013_nG17110 , RIe3bd470_5931 , \47636 , \48655 );
_HMUX g17111 ( \49014_nG17111 , \49012_nG1710e , \49013_nG17110 , \47178 );
buf \U$39045 ( \49015 , \49014_nG17111 );
_DC g18edf_GF_IsGateDCbyConstraint ( \49016_nG18edf , \49015 , \42503 );
buf \U$39046 ( \49017 , \49016_nG18edf );
_HMUX g17113 ( \49018_nG17113 , RIe3bdc68_5932 , \47642 , \48652 );
_HMUX g17114 ( \49019_nG17114 , RIe3bdc68_5932 , \49018_nG17113 , \47166 );
_HMUX g17116 ( \49020_nG17116 , RIe3bdc68_5932 , \47645 , \48655 );
_HMUX g17117 ( \49021_nG17117 , \49019_nG17114 , \49020_nG17116 , \47178 );
buf \U$39047 ( \49022 , \49021_nG17117 );
_DC g18ee1_GF_IsGateDCbyConstraint ( \49023_nG18ee1 , \49022 , \42503 );
buf \U$39048 ( \49024 , \49023_nG18ee1 );
_HMUX g17119 ( \49025_nG17119 , RIe3be460_5933 , \47651 , \48652 );
_HMUX g1711a ( \49026_nG1711a , RIe3be460_5933 , \49025_nG17119 , \47166 );
_HMUX g1711c ( \49027_nG1711c , RIe3be460_5933 , \47654 , \48655 );
_HMUX g1711d ( \49028_nG1711d , \49026_nG1711a , \49027_nG1711c , \47178 );
buf \U$39049 ( \49029 , \49028_nG1711d );
_DC g18ee3_GF_IsGateDCbyConstraint ( \49030_nG18ee3 , \49029 , \42503 );
buf \U$39050 ( \49031 , \49030_nG18ee3 );
_HMUX g1711f ( \49032_nG1711f , RIe3bec58_5934 , \47660 , \48652 );
_HMUX g17120 ( \49033_nG17120 , RIe3bec58_5934 , \49032_nG1711f , \47166 );
_HMUX g17122 ( \49034_nG17122 , RIe3bec58_5934 , \47663 , \48655 );
_HMUX g17123 ( \49035_nG17123 , \49033_nG17120 , \49034_nG17122 , \47178 );
buf \U$39051 ( \49036 , \49035_nG17123 );
_DC g18ee5_GF_IsGateDCbyConstraint ( \49037_nG18ee5 , \49036 , \42503 );
buf \U$39052 ( \49038 , \49037_nG18ee5 );
_HMUX g17125 ( \49039_nG17125 , RIe3bf450_5935 , \47669 , \48652 );
_HMUX g17126 ( \49040_nG17126 , RIe3bf450_5935 , \49039_nG17125 , \47166 );
_HMUX g17128 ( \49041_nG17128 , RIe3bf450_5935 , \47672 , \48655 );
_HMUX g17129 ( \49042_nG17129 , \49040_nG17126 , \49041_nG17128 , \47178 );
buf \U$39053 ( \49043 , \49042_nG17129 );
_DC g18ee7_GF_IsGateDCbyConstraint ( \49044_nG18ee7 , \49043 , \42503 );
buf \U$39054 ( \49045 , \49044_nG18ee7 );
_HMUX g1712b ( \49046_nG1712b , RIe3bfc48_5936 , \47678 , \48652 );
_HMUX g1712c ( \49047_nG1712c , RIe3bfc48_5936 , \49046_nG1712b , \47166 );
_HMUX g1712e ( \49048_nG1712e , RIe3bfc48_5936 , \47681 , \48655 );
_HMUX g1712f ( \49049_nG1712f , \49047_nG1712c , \49048_nG1712e , \47178 );
buf \U$39055 ( \49050 , \49049_nG1712f );
_DC g18ee9_GF_IsGateDCbyConstraint ( \49051_nG18ee9 , \49050 , \42503 );
buf \U$39056 ( \49052 , \49051_nG18ee9 );
_HMUX g17131 ( \49053_nG17131 , RIe3c0440_5937 , \47687 , \48652 );
_HMUX g17132 ( \49054_nG17132 , RIe3c0440_5937 , \49053_nG17131 , \47166 );
_HMUX g17134 ( \49055_nG17134 , RIe3c0440_5937 , \47690 , \48655 );
_HMUX g17135 ( \49056_nG17135 , \49054_nG17132 , \49055_nG17134 , \47178 );
buf \U$39057 ( \49057 , \49056_nG17135 );
_DC g18eeb_GF_IsGateDCbyConstraint ( \49058_nG18eeb , \49057 , \42503 );
buf \U$39058 ( \49059 , \49058_nG18eeb );
_HMUX g17137 ( \49060_nG17137 , RIe3c0c38_5938 , \47696 , \48652 );
_HMUX g17138 ( \49061_nG17138 , RIe3c0c38_5938 , \49060_nG17137 , \47166 );
_HMUX g1713a ( \49062_nG1713a , RIe3c0c38_5938 , \47699 , \48655 );
_HMUX g1713b ( \49063_nG1713b , \49061_nG17138 , \49062_nG1713a , \47178 );
buf \U$39059 ( \49064 , \49063_nG1713b );
_DC g18eed_GF_IsGateDCbyConstraint ( \49065_nG18eed , \49064 , \42503 );
buf \U$39060 ( \49066 , \49065_nG18eed );
_HMUX g1713d ( \49067_nG1713d , RIe3c1430_5939 , \47705 , \48652 );
_HMUX g1713e ( \49068_nG1713e , RIe3c1430_5939 , \49067_nG1713d , \47166 );
_HMUX g17140 ( \49069_nG17140 , RIe3c1430_5939 , \47708 , \48655 );
_HMUX g17141 ( \49070_nG17141 , \49068_nG1713e , \49069_nG17140 , \47178 );
buf \U$39061 ( \49071 , \49070_nG17141 );
_DC g18ef1_GF_IsGateDCbyConstraint ( \49072_nG18ef1 , \49071 , \42503 );
buf \U$39062 ( \49073 , \49072_nG18ef1 );
_HMUX g17143 ( \49074_nG17143 , RIe3c1c28_5940 , \47714 , \48652 );
_HMUX g17144 ( \49075_nG17144 , RIe3c1c28_5940 , \49074_nG17143 , \47166 );
_HMUX g17146 ( \49076_nG17146 , RIe3c1c28_5940 , \47717 , \48655 );
_HMUX g17147 ( \49077_nG17147 , \49075_nG17144 , \49076_nG17146 , \47178 );
buf \U$39063 ( \49078 , \49077_nG17147 );
_DC g18ef3_GF_IsGateDCbyConstraint ( \49079_nG18ef3 , \49078 , \42503 );
buf \U$39064 ( \49080 , \49079_nG18ef3 );
_HMUX g17149 ( \49081_nG17149 , RIe3c2420_5941 , \47723 , \48652 );
_HMUX g1714a ( \49082_nG1714a , RIe3c2420_5941 , \49081_nG17149 , \47166 );
_HMUX g1714c ( \49083_nG1714c , RIe3c2420_5941 , \47726 , \48655 );
_HMUX g1714d ( \49084_nG1714d , \49082_nG1714a , \49083_nG1714c , \47178 );
buf \U$39065 ( \49085 , \49084_nG1714d );
_DC g18ef5_GF_IsGateDCbyConstraint ( \49086_nG18ef5 , \49085 , \42503 );
buf \U$39066 ( \49087 , \49086_nG18ef5 );
_HMUX g1714f ( \49088_nG1714f , RIe3c2c18_5942 , \47732 , \48652 );
_HMUX g17150 ( \49089_nG17150 , RIe3c2c18_5942 , \49088_nG1714f , \47166 );
_HMUX g17152 ( \49090_nG17152 , RIe3c2c18_5942 , \47735 , \48655 );
_HMUX g17153 ( \49091_nG17153 , \49089_nG17150 , \49090_nG17152 , \47178 );
buf \U$39067 ( \49092 , \49091_nG17153 );
_DC g18ef7_GF_IsGateDCbyConstraint ( \49093_nG18ef7 , \49092 , \42503 );
buf \U$39068 ( \49094 , \49093_nG18ef7 );
_HMUX g17155 ( \49095_nG17155 , RIe3c3410_5943 , \47741 , \48652 );
_HMUX g17156 ( \49096_nG17156 , RIe3c3410_5943 , \49095_nG17155 , \47166 );
_HMUX g17158 ( \49097_nG17158 , RIe3c3410_5943 , \47744 , \48655 );
_HMUX g17159 ( \49098_nG17159 , \49096_nG17156 , \49097_nG17158 , \47178 );
buf \U$39069 ( \49099 , \49098_nG17159 );
_DC g18ef9_GF_IsGateDCbyConstraint ( \49100_nG18ef9 , \49099 , \42503 );
buf \U$39070 ( \49101 , \49100_nG18ef9 );
buf \U$39071 ( \49102 , RIb86fc68_77);
_HMUX g16faa ( \49103_nG16faa , RIe202f10_5656 , \49102 , \47158 );
not \U$39072 ( \49104 , \47166 );
or \U$39073 ( \49105 , \47178 , \49104 );
_HMUX g16fab ( \49106_nG16fab , \49103_nG16faa , RIe202f10_5656 , \49105 );
buf \U$39074 ( \49107 , \49106_nG16fab );
_DC g18e69_GF_IsGateDCbyConstraint ( \49108_nG18e69 , \49107 , \42503 );
buf \U$39075 ( \49109 , \49108_nG18e69 );
buf \U$39076 ( \49110 , RIb86fce0_76);
_HMUX g16fac ( \49111_nG16fac , RIe202448_5657 , \49110 , \47158 );
_HMUX g16fad ( \49112_nG16fad , \49111_nG16fac , RIe202448_5657 , \49105 );
buf \U$39077 ( \49113 , \49112_nG16fad );
_DC g18e6b_GF_IsGateDCbyConstraint ( \49114_nG18e6b , \49113 , \42503 );
buf \U$39078 ( \49115 , \49114_nG18e6b );
buf \U$39079 ( \49116 , RIb86fd58_75);
_HMUX g16fae ( \49117_nG16fae , RIe201980_5658 , \49116 , \47158 );
_HMUX g16faf ( \49118_nG16faf , \49117_nG16fae , RIe201980_5658 , \49105 );
buf \U$39080 ( \49119 , \49118_nG16faf );
_DC g18e6d_GF_IsGateDCbyConstraint ( \49120_nG18e6d , \49119 , \42503 );
buf \U$39081 ( \49121 , \49120_nG18e6d );
buf \U$39082 ( \49122 , RIb87e8a8_74);
_HMUX g16fb0 ( \49123_nG16fb0 , RIe200e40_5659 , \49122 , \47158 );
_HMUX g16fb1 ( \49124_nG16fb1 , \49123_nG16fb0 , RIe200e40_5659 , \49105 );
buf \U$39083 ( \49125 , \49124_nG16fb1 );
_DC g18e6f_GF_IsGateDCbyConstraint ( \49126_nG18e6f , \49125 , \42503 );
buf \U$39084 ( \49127 , \49126_nG18e6f );
buf \U$39085 ( \49128 , RIb87e920_73);
_HMUX g16fb2 ( \49129_nG16fb2 , RIe2000a8_5660 , \49128 , \47158 );
_HMUX g16fb3 ( \49130_nG16fb3 , \49129_nG16fb2 , RIe2000a8_5660 , \49105 );
buf \U$39086 ( \49131 , \49130_nG16fb3 );
_DC g18e71_GF_IsGateDCbyConstraint ( \49132_nG18e71 , \49131 , \42503 );
buf \U$39087 ( \49133 , \49132_nG18e71 );
buf \U$39088 ( \49134 , RIb87e998_72);
_HMUX g16fb4 ( \49135_nG16fb4 , RIe1ff310_5661 , \49134 , \47158 );
_HMUX g16fb5 ( \49136_nG16fb5 , \49135_nG16fb4 , RIe1ff310_5661 , \49105 );
buf \U$39089 ( \49137 , \49136_nG16fb5 );
_DC g18e73_GF_IsGateDCbyConstraint ( \49138_nG18e73 , \49137 , \42503 );
buf \U$39090 ( \49139 , \49138_nG18e73 );
buf \U$39091 ( \49140 , RIb87ea10_71);
_HMUX g16fb6 ( \49141_nG16fb6 , RIe1fe668_5662 , \49140 , \47158 );
_HMUX g16fb7 ( \49142_nG16fb7 , \49141_nG16fb6 , RIe1fe668_5662 , \49105 );
buf \U$39092 ( \49143 , \49142_nG16fb7 );
_DC g18e75_GF_IsGateDCbyConstraint ( \49144_nG18e75 , \49143 , \42503 );
buf \U$39093 ( \49145 , \49144_nG18e75 );
buf \U$39094 ( \49146 , RIb87ea88_70);
_HMUX g16fb8 ( \49147_nG16fb8 , RIe1fd9c0_5663 , \49146 , \47158 );
_HMUX g16fb9 ( \49148_nG16fb9 , \49147_nG16fb8 , RIe1fd9c0_5663 , \49105 );
buf \U$39095 ( \49149 , \49148_nG16fb9 );
_DC g18e77_GF_IsGateDCbyConstraint ( \49150_nG18e77 , \49149 , \42503 );
buf \U$39096 ( \49151 , \49150_nG18e77 );
_HMUX g16f99 ( \49152_nG16f99 , RIe1fce80_5664 , \49102 , \47751 );
_HMUX g16f9a ( \49153_nG16f9a , \49152_nG16f99 , RIe1fce80_5664 , \49105 );
buf \U$39097 ( \49154 , \49153_nG16f9a );
_DC g18e59_GF_IsGateDCbyConstraint ( \49155_nG18e59 , \49154 , \42503 );
buf \U$39098 ( \49156 , \49155_nG18e59 );
_HMUX g16f9b ( \49157_nG16f9b , RIe1fc340_5665 , \49110 , \47751 );
_HMUX g16f9c ( \49158_nG16f9c , \49157_nG16f9b , RIe1fc340_5665 , \49105 );
buf \U$39099 ( \49159 , \49158_nG16f9c );
_DC g18e5b_GF_IsGateDCbyConstraint ( \49160_nG18e5b , \49159 , \42503 );
buf \U$39100 ( \49161 , \49160_nG18e5b );
_HMUX g16f9d ( \49162_nG16f9d , RIe1fb878_5666 , \49116 , \47751 );
_HMUX g16f9e ( \49163_nG16f9e , \49162_nG16f9d , RIe1fb878_5666 , \49105 );
buf \U$39101 ( \49164 , \49163_nG16f9e );
_DC g18e5d_GF_IsGateDCbyConstraint ( \49165_nG18e5d , \49164 , \42503 );
buf \U$39102 ( \49166 , \49165_nG18e5d );
_HMUX g16f9f ( \49167_nG16f9f , RIe1facc0_5667 , \49122 , \47751 );
_HMUX g16fa0 ( \49168_nG16fa0 , \49167_nG16f9f , RIe1facc0_5667 , \49105 );
buf \U$39103 ( \49169 , \49168_nG16fa0 );
_DC g18e5f_GF_IsGateDCbyConstraint ( \49170_nG18e5f , \49169 , \42503 );
buf \U$39104 ( \49171 , \49170_nG18e5f );
_HMUX g16fa1 ( \49172_nG16fa1 , RIe1fa090_5668 , \49128 , \47751 );
_HMUX g16fa2 ( \49173_nG16fa2 , \49172_nG16fa1 , RIe1fa090_5668 , \49105 );
buf \U$39105 ( \49174 , \49173_nG16fa2 );
_DC g18e61_GF_IsGateDCbyConstraint ( \49175_nG18e61 , \49174 , \42503 );
buf \U$39106 ( \49176 , \49175_nG18e61 );
_HMUX g16fa3 ( \49177_nG16fa3 , RIe1f9118_5669 , \49134 , \47751 );
_HMUX g16fa4 ( \49178_nG16fa4 , \49177_nG16fa3 , RIe1f9118_5669 , \49105 );
buf \U$39107 ( \49179 , \49178_nG16fa4 );
_DC g18e63_GF_IsGateDCbyConstraint ( \49180_nG18e63 , \49179 , \42503 );
buf \U$39108 ( \49181 , \49180_nG18e63 );
_HMUX g16fa5 ( \49182_nG16fa5 , RIe1f7fc0_5670 , \49140 , \47751 );
_HMUX g16fa6 ( \49183_nG16fa6 , \49182_nG16fa5 , RIe1f7fc0_5670 , \49105 );
buf \U$39109 ( \49184 , \49183_nG16fa6 );
_DC g18e65_GF_IsGateDCbyConstraint ( \49185_nG18e65 , \49184 , \42503 );
buf \U$39110 ( \49186 , \49185_nG18e65 );
_HMUX g16fa7 ( \49187_nG16fa7 , RIe1f69b8_5671 , \49146 , \47751 );
_HMUX g16fa8 ( \49188_nG16fa8 , \49187_nG16fa7 , RIe1f69b8_5671 , \49105 );
buf \U$39111 ( \49189 , \49188_nG16fa8 );
_DC g18e67_GF_IsGateDCbyConstraint ( \49190_nG18e67 , \49189 , \42503 );
buf \U$39112 ( \49191 , \49190_nG18e67 );
_HMUX g16f88 ( \49192_nG16f88 , RIe1f5860_5672 , \49102 , \48202 );
_HMUX g16f89 ( \49193_nG16f89 , \49192_nG16f88 , RIe1f5860_5672 , \49105 );
buf \U$39113 ( \49194 , \49193_nG16f89 );
_DC g18e49_GF_IsGateDCbyConstraint ( \49195_nG18e49 , \49194 , \42503 );
buf \U$39114 ( \49196 , \49195_nG18e49 );
_HMUX g16f8a ( \49197_nG16f8a , RIe1f4258_5673 , \49110 , \48202 );
_HMUX g16f8b ( \49198_nG16f8b , \49197_nG16f8a , RIe1f4258_5673 , \49105 );
buf \U$39115 ( \49199 , \49198_nG16f8b );
_DC g18e4b_GF_IsGateDCbyConstraint ( \49200_nG18e4b , \49199 , \42503 );
buf \U$39116 ( \49201 , \49200_nG18e4b );
_HMUX g16f8c ( \49202_nG16f8c , RIe1f3100_5674 , \49116 , \48202 );
_HMUX g16f8d ( \49203_nG16f8d , \49202_nG16f8c , RIe1f3100_5674 , \49105 );
buf \U$39117 ( \49204 , \49203_nG16f8d );
_DC g18e4d_GF_IsGateDCbyConstraint ( \49205_nG18e4d , \49204 , \42503 );
buf \U$39118 ( \49206 , \49205_nG18e4d );
_HMUX g16f8e ( \49207_nG16f8e , RIe1f1fa8_5675 , \49122 , \48202 );
_HMUX g16f8f ( \49208_nG16f8f , \49207_nG16f8e , RIe1f1fa8_5675 , \49105 );
buf \U$39119 ( \49209 , \49208_nG16f8f );
_DC g18e4f_GF_IsGateDCbyConstraint ( \49210_nG18e4f , \49209 , \42503 );
buf \U$39120 ( \49211 , \49210_nG18e4f );
_HMUX g16f90 ( \49212_nG16f90 , RIe1f09a0_5676 , \49128 , \48202 );
_HMUX g16f91 ( \49213_nG16f91 , \49212_nG16f90 , RIe1f09a0_5676 , \49105 );
buf \U$39121 ( \49214 , \49213_nG16f91 );
_DC g18e51_GF_IsGateDCbyConstraint ( \49215_nG18e51 , \49214 , \42503 );
buf \U$39122 ( \49216 , \49215_nG18e51 );
_HMUX g16f92 ( \49217_nG16f92 , RIe1ef848_5677 , \49134 , \48202 );
_HMUX g16f93 ( \49218_nG16f93 , \49217_nG16f92 , RIe1ef848_5677 , \49105 );
buf \U$39123 ( \49219 , \49218_nG16f93 );
_DC g18e53_GF_IsGateDCbyConstraint ( \49220_nG18e53 , \49219 , \42503 );
buf \U$39124 ( \49221 , \49220_nG18e53 );
_HMUX g16f94 ( \49222_nG16f94 , RIe1ee240_5678 , \49140 , \48202 );
_HMUX g16f95 ( \49223_nG16f95 , \49222_nG16f94 , RIe1ee240_5678 , \49105 );
buf \U$39125 ( \49224 , \49223_nG16f95 );
_DC g18e55_GF_IsGateDCbyConstraint ( \49225_nG18e55 , \49224 , \42503 );
buf \U$39126 ( \49226 , \49225_nG18e55 );
_HMUX g16f96 ( \49227_nG16f96 , RIe1ed0e8_5679 , \49146 , \48202 );
_HMUX g16f97 ( \49228_nG16f97 , \49227_nG16f96 , RIe1ed0e8_5679 , \49105 );
buf \U$39127 ( \49229 , \49228_nG16f97 );
_DC g18e57_GF_IsGateDCbyConstraint ( \49230_nG18e57 , \49229 , \42503 );
buf \U$39128 ( \49231 , \49230_nG18e57 );
_HMUX g16f67 ( \49232_nG16f67 , RIe1ebae0_5680 , \49102 , \48652 );
_HMUX g16f70 ( \49233_nG16f70 , \49232_nG16f67 , RIe1ebae0_5680 , \49105 );
buf \U$39129 ( \49234 , \49233_nG16f70 );
_DC g19081_GF_IsGateDCbyConstraint ( \49235_nG19081 , \49234 , \42503 );
buf \U$39130 ( \49236 , \49235_nG19081 );
_HMUX g16f72 ( \49237_nG16f72 , RIe1ea988_5681 , \49110 , \48652 );
_HMUX g16f73 ( \49238_nG16f73 , \49237_nG16f72 , RIe1ea988_5681 , \49105 );
buf \U$39131 ( \49239 , \49238_nG16f73 );
_DC g19083_GF_IsGateDCbyConstraint ( \49240_nG19083 , \49239 , \42503 );
buf \U$39132 ( \49241 , \49240_nG19083 );
_HMUX g16f75 ( \49242_nG16f75 , RIe1e9830_5682 , \49116 , \48652 );
_HMUX g16f76 ( \49243_nG16f76 , \49242_nG16f75 , RIe1e9830_5682 , \49105 );
buf \U$39133 ( \49244 , \49243_nG16f76 );
_DC g19085_GF_IsGateDCbyConstraint ( \49245_nG19085 , \49244 , \42503 );
buf \U$39134 ( \49246 , \49245_nG19085 );
_HMUX g16f78 ( \49247_nG16f78 , RIe1e8228_5683 , \49122 , \48652 );
_HMUX g16f79 ( \49248_nG16f79 , \49247_nG16f78 , RIe1e8228_5683 , \49105 );
buf \U$39135 ( \49249 , \49248_nG16f79 );
_DC g19087_GF_IsGateDCbyConstraint ( \49250_nG19087 , \49249 , \42503 );
buf \U$39136 ( \49251 , \49250_nG19087 );
_HMUX g16f7b ( \49252_nG16f7b , RIe1e70d0_5684 , \49128 , \48652 );
_HMUX g16f7c ( \49253_nG16f7c , \49252_nG16f7b , RIe1e70d0_5684 , \49105 );
buf \U$39137 ( \49254 , \49253_nG16f7c );
_DC g19089_GF_IsGateDCbyConstraint ( \49255_nG19089 , \49254 , \42503 );
buf \U$39138 ( \49256 , \49255_nG19089 );
_HMUX g16f7e ( \49257_nG16f7e , RIe1e5ac8_5685 , \49134 , \48652 );
_HMUX g16f7f ( \49258_nG16f7f , \49257_nG16f7e , RIe1e5ac8_5685 , \49105 );
buf \U$39139 ( \49259 , \49258_nG16f7f );
_DC g1908b_GF_IsGateDCbyConstraint ( \49260_nG1908b , \49259 , \42503 );
buf \U$39140 ( \49261 , \49260_nG1908b );
_HMUX g16f81 ( \49262_nG16f81 , RIe1e4970_5686 , \49140 , \48652 );
_HMUX g16f82 ( \49263_nG16f82 , \49262_nG16f81 , RIe1e4970_5686 , \49105 );
buf \U$39141 ( \49264 , \49263_nG16f82 );
_DC g1908d_GF_IsGateDCbyConstraint ( \49265_nG1908d , \49264 , \42503 );
buf \U$39142 ( \49266 , \49265_nG1908d );
_HMUX g16f84 ( \49267_nG16f84 , RIe1e3368_5687 , \49146 , \48652 );
_HMUX g16f85 ( \49268_nG16f85 , \49267_nG16f84 , RIe1e3368_5687 , \49105 );
buf \U$39143 ( \49269 , \49268_nG16f85 );
_DC g1908f_GF_IsGateDCbyConstraint ( \49270_nG1908f , \49269 , \42503 );
buf \U$39144 ( \49271 , \49270_nG1908f );
buf \U$39145 ( \49272 , RIb7b9680_245);
buf \U$39146 ( \49273 , RIb79b3b0_273);
and \U$39147 ( \49274 , \47174 , \49273 );
_HMUX g16e5c ( \49275_nG16e5c , RIe4520c0_5970 , \49272 , \49274 );
buf \U$39148 ( \49276 , \49275_nG16e5c );
_DC g19090_GF_IsGateDCbyConstraint ( \49277_nG19090 , \49276 , \42503 );
buf \U$39149 ( \49278 , \49277_nG19090 );
buf \U$39150 ( \49279 , RIb7b96f8_244);
_HMUX g16ec9 ( \49280_nG16ec9 , RIe438440_5990 , \49279 , \49274 );
buf \U$39151 ( \49281 , \49280_nG16ec9 );
_DC g18e2d_GF_IsGateDCbyConstraint ( \49282_nG18e2d , \49281 , \42503 );
buf \U$39152 ( \49283 , \49282_nG18e2d );
buf \U$39153 ( \49284 , RIb7c20c8_243);
_HMUX g16ecb ( \49285_nG16ecb , RIe4390e8_5989 , \49284 , \49274 );
buf \U$39154 ( \49286 , \49285_nG16ecb );
_DC g18e2f_GF_IsGateDCbyConstraint ( \49287_nG18e2f , \49286 , \42503 );
buf \U$39155 ( \49288 , \49287_nG18e2f );
buf \U$39156 ( \49289 , RIb7c5728_242);
_HMUX g16ecd ( \49290_nG16ecd , RIe439f70_5988 , \49289 , \49274 );
buf \U$39157 ( \49291 , \49290_nG16ecd );
_DC g18e31_GF_IsGateDCbyConstraint ( \49292_nG18e31 , \49291 , \42503 );
buf \U$39158 ( \49293 , \49292_nG18e31 );
buf \U$39159 ( \49294 , RIb7c57a0_241);
_HMUX g16ecf ( \49295_nG16ecf , RIe43ad80_5987 , \49294 , \49274 );
buf \U$39160 ( \49296 , \49295_nG16ecf );
_DC g18e33_GF_IsGateDCbyConstraint ( \49297_nG18e33 , \49296 , \42503 );
buf \U$39161 ( \49298 , \49297_nG18e33 );
buf \U$39162 ( \49299 , RIb7c5818_240);
_HMUX g16ed1 ( \49300_nG16ed1 , RIe43ba28_5986 , \49299 , \49274 );
buf \U$39163 ( \49301 , \49300_nG16ed1 );
_DC g18e35_GF_IsGateDCbyConstraint ( \49302_nG18e35 , \49301 , \42503 );
buf \U$39164 ( \49303 , \49302_nG18e35 );
buf \U$39165 ( \49304 , RIb7c5890_239);
_HMUX g16ed3 ( \49305_nG16ed3 , RIe43c7c0_5985 , \49304 , \49274 );
buf \U$39166 ( \49306 , \49305_nG16ed3 );
_DC g18e37_GF_IsGateDCbyConstraint ( \49307_nG18e37 , \49306 , \42503 );
buf \U$39167 ( \49308 , \49307_nG18e37 );
buf \U$39168 ( \49309 , RIb7c5908_238);
_HMUX g16ed5 ( \49310_nG16ed5 , RIe43d5d0_5984 , \49309 , \49274 );
buf \U$39169 ( \49311 , \49310_nG16ed5 );
_DC g18e39_GF_IsGateDCbyConstraint ( \49312_nG18e39 , \49311 , \42503 );
buf \U$39170 ( \49313 , \49312_nG18e39 );
buf \U$39171 ( \49314 , RIb7a09f0_266);
_HMUX g16ec7 ( \49315_nG16ec7 , RIe445e38_5974 , \49314 , \49274 );
buf \U$39172 ( \49316 , \49315_nG16ec7 );
_DC g18e2b_GF_IsGateDCbyConstraint ( \49317_nG18e2b , \49316 , \42503 );
buf \U$39173 ( \49318 , \49317_nG18e2b );
buf \U$39174 ( \49319 , RIb7a0a68_265);
_HMUX g16ebf ( \49320_nG16ebf , RIe441c98_5979 , \49319 , \49274 );
buf \U$39175 ( \49321 , \49320_nG16ebf );
_DC g18e23_GF_IsGateDCbyConstraint ( \49322_nG18e23 , \49321 , \42503 );
buf \U$39176 ( \49323 , \49322_nG18e23 );
buf \U$39177 ( \49324 , RIb7a0ae0_264);
_HMUX g16ec1 ( \49325_nG16ec1 , RIe4429b8_5978 , \49324 , \49274 );
buf \U$39178 ( \49326 , \49325_nG16ec1 );
_DC g18e25_GF_IsGateDCbyConstraint ( \49327_nG18e25 , \49326 , \42503 );
buf \U$39179 ( \49328 , \49327_nG18e25 );
buf \U$39180 ( \49329 , RIb7a0b58_263);
_HMUX g16ec3 ( \49330_nG16ec3 , RIe443750_5977 , \49329 , \49274 );
buf \U$39181 ( \49331 , \49330_nG16ec3 );
_DC g18e27_GF_IsGateDCbyConstraint ( \49332_nG18e27 , \49331 , \42503 );
buf \U$39182 ( \49333 , \49332_nG18e27 );
buf \U$39183 ( \49334 , RIb7a0bd0_262);
_HMUX g16ec5 ( \49335_nG16ec5 , RIe437630_5991 , \49334 , \49274 );
buf \U$39184 ( \49336 , \49335_nG16ec5 );
_DC g18e29_GF_IsGateDCbyConstraint ( \49337_nG18e29 , \49336 , \42503 );
buf \U$39185 ( \49338 , \49337_nG18e29 );
buf \U$39186 ( \49339 , RIe45a478_5957);
not \U$39187 ( \49340 , \49339 );
buf \U$39188 ( \49341 , \49340 );
nor \U$39190 ( \49342 , RIe45a478_5957, RIe45aec8_5956, RIe45b8a0_5955);
_HMUX g16d2f ( \49343_nG16d2f , \49341 , 1'b0 , \49342 );
and \U$39191 ( \49344 , \40007 , RIe549ef0_6842, RIe549770_6843, RIe548ff0_6844, \7063 );
buf \U$39192 ( \49345 , \49344 );
buf \U$39193 ( \49346 , RIb79b4a0_271);
and \U$39194 ( \49347 , \49345 , \49346 );
_HMUX g16d30 ( \49348_nG16d30 , RIe45a478_5957 , \49343_nG16d2f , \49347 );
buf \U$39195 ( \49349 , RIe45a478_5957);
not \U$39196 ( \49350 , \49349 );
buf \U$39197 ( \49351 , \49350 );
not \U$39198 ( \49352 , RIe45b8a0_5955);
nor \U$39199 ( \49353 , RIe45a478_5957, RIe45aec8_5956, \49352 );
_HMUX g16d36 ( \49354_nG16d36 , \49351 , RIe45a478_5957 , \49353 );
and \U$39200 ( \49355 , \47176 , \47174 );
_HMUX g16d3a ( \49356_nG16d3a , \49348_nG16d30 , \49354_nG16d36 , \49355 );
and \U$39201 ( \49357 , \49355 , \49346 );
and \U$39202 ( \49358 , \49357 , \49345 );
_HMUX g16d3d ( \49359_nG16d3d , \49356_nG16d3a , RIe45a478_5957 , \49358 );
not \U$39203 ( \49360 , RIe444fb0_5975);
and \U$39204 ( \49361 , RIe444fb0_5975, \49272 );
or \U$39205 ( \49362 , \49360 , \49361 );
and \U$39206 ( \49363 , \49362 , \47176 );
and \U$39207 ( \49364 , \49363 , \47174 );
_HMUX g16d44 ( \49365_nG16d44 , \49359_nG16d3d , RIe452b88_5969 , \49364 );
buf \U$39209 ( \49366 , RIb79b338_274);
and \U$39210 ( \49367 , \49345 , \49366 );
_HMUX g16d45 ( \49368_nG16d45 , \49365_nG16d44 , 1'b0 , \49367 );
buf \U$39211 ( \49369 , \49368_nG16d45 );
buf \U$39212 ( \49370 , RIe45aec8_5956);
xnor \U$39213 ( \49371 , \49370 , \49339 );
buf \U$39214 ( \49372 , \49371 );
_HMUX g16d49 ( \49373_nG16d49 , \49372 , 1'b0 , \49342 );
_HMUX g16d4a ( \49374_nG16d4a , RIe45aec8_5956 , \49373_nG16d49 , \49347 );
buf \U$39216 ( \49375 , RIe45aec8_5956);
xor \U$39217 ( \49376 , \49375 , \49349 );
buf \U$39218 ( \49377 , \49376 );
_HMUX g16d4e ( \49378_nG16d4e , \49377 , RIe45aec8_5956 , \49353 );
_HMUX g16d4f ( \49379_nG16d4f , \49374_nG16d4a , \49378_nG16d4e , \49355 );
_HMUX g16d50 ( \49380_nG16d50 , \49379_nG16d4f , RIe45aec8_5956 , \49358 );
_HMUX g16d51 ( \49381_nG16d51 , \49380_nG16d50 , RIe4534e8_5968 , \49364 );
_HMUX g16d52 ( \49382_nG16d52 , \49381_nG16d51 , 1'b0 , \49367 );
buf \U$39219 ( \49383 , \49382_nG16d52 );
buf \U$39220 ( \49384 , RIe45b8a0_5955);
or \U$39221 ( \49385 , \49370 , \49339 );
xnor \U$39222 ( \49386 , \49384 , \49385 );
buf \U$39223 ( \49387 , \49386 );
_HMUX g16d57 ( \49388_nG16d57 , \49387 , 1'b0 , \49342 );
_HMUX g16d58 ( \49389_nG16d58 , RIe45b8a0_5955 , \49388_nG16d57 , \49347 );
buf \U$39225 ( \49390 , RIe45b8a0_5955);
and \U$39226 ( \49391 , \49375 , \49349 );
xor \U$39227 ( \49392 , \49390 , \49391 );
buf \U$39228 ( \49393 , \49392 );
_HMUX g16d5d ( \49394_nG16d5d , \49393 , RIe45b8a0_5955 , \49353 );
_HMUX g16d5e ( \49395_nG16d5e , \49389_nG16d58 , \49394_nG16d5d , \49355 );
_HMUX g16d5f ( \49396_nG16d5f , \49395_nG16d5e , RIe45b8a0_5955 , \49358 );
_HMUX g16d60 ( \49397_nG16d60 , \49396_nG16d5f , RIe453fb0_5967 , \49364 );
_HMUX g16d61 ( \49398_nG16d61 , \49397_nG16d60 , 1'b0 , \49367 );
buf \U$39230 ( \49399 , \49398_nG16d61 );
or \U$39231 ( \49400 , \49369 , \49383 , \49399 );
buf \U$39232 ( \49401 , \49400 );
buf \U$39233 ( \49402 , RIe45d880_5952);
buf \U$39234 ( \49403 , RIe45cdb8_5953);
buf \U$39235 ( \49404 , RIe45c278_5954);
and \U$39236 ( \49405 , \49403 , \49404 );
xor \U$39237 ( \49406 , \49402 , \49405 );
buf \U$39238 ( \49407 , \49406 );
not \U$39239 ( \49408 , RIe45d880_5952);
nor \U$39240 ( \49409 , RIe45c278_5954, RIe45cdb8_5953, \49408 );
not \U$39241 ( \49410 , \49409 );
and \U$39242 ( \49411 , \49347 , \49410 );
_HMUX g16d26 ( \49412_nG16d26 , RIe45d880_5952 , \49407 , \49411 );
_HMUX g16d27 ( \49413_nG16d27 , \49412_nG16d26 , 1'b0 , \49367 );
buf \U$39244 ( \49414 , \49413_nG16d27 );
not \U$39245 ( \49415 , \49414 );
buf \U$39246 ( \49416 , RIe455e28_5964);
buf \U$39247 ( \49417 , RIe4554c8_5965);
buf \U$39248 ( \49418 , RIe454988_5966);
and \U$39249 ( \49419 , \49417 , \49418 );
xor \U$39250 ( \49420 , \49416 , \49419 );
buf \U$39251 ( \49421 , \49420 );
buf \U$39252 ( \49422 , RIb839848_152);
and \U$39253 ( \49423 , \47162 , \49422 );
not \U$39254 ( \49424 , RIe4554c8_5965);
and \U$39255 ( \49425 , RIe454988_5966, \49424 , RIe455e28_5964);
not \U$39256 ( \49426 , \49425 );
and \U$39257 ( \49427 , \49423 , \49426 );
_HMUX g16de4 ( \49428_nG16de4 , RIe455e28_5964 , \49421 , \49427 );
buf \U$39258 ( \49429 , RIe455e28_5964);
buf \U$39259 ( \49430 , RIe4554c8_5965);
xor \U$39260 ( \49431 , \49429 , \49430 );
buf \U$39261 ( \49432 , \49431 );
not \U$39262 ( \49433 , RIe454988_5966);
and \U$39263 ( \49434 , \49433 , \49424 , RIe455e28_5964);
or \U$39264 ( \49435 , \49434 , \49425 );
_HMUX g16de8 ( \49436_nG16de8 , \49432 , RIe455e28_5964 , \49435 );
buf \U$39265 ( \49437 , RIb839668_156);
and \U$39266 ( \49438 , \47162 , \49437 );
_HMUX g16de9 ( \49439_nG16de9 , \49428_nG16de4 , \49436_nG16de8 , \49438 );
buf \U$39268 ( \49440 , RIb8396e0_155);
and \U$39269 ( \49441 , \47162 , \49440 );
_HMUX g16dea ( \49442_nG16dea , \49439_nG16de9 , 1'b0 , \49441 );
and \U$39271 ( \49443 , \49441 , \49437 );
_HMUX g16deb ( \49444_nG16deb , \49442_nG16dea , 1'b0 , \49443 );
buf \U$39272 ( \49445 , \49444_nG16deb );
and \U$39273 ( \49446 , \49415 , \49445 );
xor \U$39274 ( \49447 , \49403 , \49404 );
buf \U$39275 ( \49448 , \49447 );
_HMUX g16d20 ( \49449_nG16d20 , RIe45cdb8_5953 , \49448 , \49411 );
_HMUX g16d21 ( \49450_nG16d21 , \49449_nG16d20 , 1'b0 , \49367 );
buf \U$39277 ( \49451 , \49450_nG16d21 );
not \U$39278 ( \49452 , \49451 );
xor \U$39279 ( \49453 , \49417 , \49418 );
buf \U$39280 ( \49454 , \49453 );
_HMUX g16dd5 ( \49455_nG16dd5 , RIe4554c8_5965 , \49454 , \49427 );
not \U$39281 ( \49456 , \49430 );
buf \U$39282 ( \49457 , \49456 );
_HMUX g16ddc ( \49458_nG16ddc , \49457 , RIe4554c8_5965 , \49435 );
_HMUX g16ddd ( \49459_nG16ddd , \49455_nG16dd5 , \49458_nG16ddc , \49438 );
_HMUX g16dde ( \49460_nG16dde , \49459_nG16ddd , 1'b0 , \49441 );
_HMUX g16ddf ( \49461_nG16ddf , \49460_nG16dde , 1'b1 , \49443 );
buf \U$39285 ( \49462 , \49461_nG16ddf );
and \U$39286 ( \49463 , \49452 , \49462 );
not \U$39287 ( \49464 , \49404 );
buf \U$39288 ( \49465 , \49464 );
_HMUX g16d19 ( \49466_nG16d19 , RIe45c278_5954 , \49465 , \49411 );
_HMUX g16d1c ( \49467_nG16d1c , \49466_nG16d19 , 1'b0 , \49367 );
buf \U$39290 ( \49468 , \49467_nG16d1c );
not \U$39291 ( \49469 , \49468 );
not \U$39292 ( \49470 , \49418 );
buf \U$39293 ( \49471 , \49470 );
_HMUX g16dc5 ( \49472_nG16dc5 , RIe454988_5966 , \49471 , \49427 );
buf \U$39294 ( \49473 , RIe454988_5966);
buf g16dc9( \49474_nG16dc9 , \49473 );
_HMUX g16dcc ( \49475_nG16dcc , \49472_nG16dc5 , \49474_nG16dc9 , \49438 );
_HMUX g16dcf ( \49476_nG16dcf , \49475_nG16dcc , 1'b1 , \49441 );
_HMUX g16dd1 ( \49477_nG16dd1 , \49476_nG16dcf , 1'b0 , \49443 );
buf \U$39299 ( \49478 , \49477_nG16dd1 );
and \U$39300 ( \49479 , \49469 , \49478 );
xnor \U$39301 ( \49480 , \49462 , \49451 );
and \U$39302 ( \49481 , \49479 , \49480 );
or \U$39303 ( \49482 , \49463 , \49481 );
xnor \U$39304 ( \49483 , \49445 , \49414 );
and \U$39305 ( \49484 , \49482 , \49483 );
or \U$39306 ( \49485 , \49446 , \49484 );
buf \U$39307 ( \49486 , \49485 );
and \U$39308 ( \49487 , \49401 , \49486 );
not \U$39310 ( \49488 , \49275_nG16e5c );
or \U$39311 ( \49489 , \49488 , \49360 );
and \U$39312 ( \49490 , \49401 , \49489 );
_HMUX g16e60 ( \49491_nG16e60 , \49487 , 1'b1 , \49490 );
buf \U$39313 ( \49492 , \49491_nG16e60 );
_DC g18e47_GF_IsGateDCbyConstraint ( \49493_nG18e47 , \49492 , \42503 );
buf \U$39314 ( \49494 , \49493_nG18e47 );
buf \U$39315 ( \49495 , \49368_nG16d45 );
_DC g19094_GF_IsGateDCbyConstraint ( \49496_nG19094 , \49495 , \42503 );
buf \U$39316 ( \49497 , \49496_nG19094 );
buf \U$39317 ( \49498 , \49382_nG16d52 );
_DC g19095_GF_IsGateDCbyConstraint ( \49499_nG19095 , \49498 , \42503 );
buf \U$39318 ( \49500 , \49499_nG19095 );
buf \U$39319 ( \49501 , \49398_nG16d61 );
_DC g19096_GF_IsGateDCbyConstraint ( \49502_nG19096 , \49501 , \42503 );
buf \U$39320 ( \49503 , \49502_nG19096 );
buf \U$39321 ( \49504 , RIb87eb00_69);
buf \U$39322 ( \49505 , RIe667bb0_6885);
buf \U$39323 ( \49506 , RIe667f70_6886);
nor \U$39324 ( \49507 , \49505 , \49506 );
_HMUX g16c0a ( \49508_nG16c0a , RIe116b70_5293 , \49504 , \49507 );
and \U$39325 ( \49509 , RIea90778_6887, \42387 , RIe546098_6850, RIe545dc8_6851, \42389 );
buf \U$39326 ( \49510 , \49509 );
buf \U$39327 ( \49511 , \49510 );
buf \U$39328 ( \49512 , \42587 );
buf \U$39329 ( \49513 , \49512 );
and \U$39330 ( \49514 , \49511 , \49513 );
_HMUX g16c0b ( \49515_nG16c0b , RIe116b70_5293 , \49508_nG16c0a , \49514 );
buf \U$39331 ( \49516 , RIb7c5980_237);
buf \U$39332 ( \49517 , RIeab7058_6894);
buf \U$39333 ( \49518 , RIea91768_6889);
nor \U$39334 ( \49519 , \49517 , \49518 );
_HMUX g16c0d ( \49520_nG16c0d , RIe116b70_5293 , \49516 , \49519 );
and \U$39335 ( \49521 , \42121_nGbbbc , \42170 , \42218_nGbc1c , \42267_nGbc4c , \42316 );
buf \U$39336 ( \49522 , \49521 );
buf \U$39337 ( \49523 , \49522 );
buf \U$39338 ( \49524 , RIb79b518_270);
buf \U$39339 ( \49525 , \49524 );
and \U$39340 ( \49526 , \49523 , \49525 );
_HMUX g16c0e ( \49527_nG16c0e , \49515_nG16c0b , \49520_nG16c0d , \49526 );
buf \U$39341 ( \49528 , \49527_nG16c0e );
_DC g18d84_GF_IsGateDCbyConstraint ( \49529_nG18d84 , \49528 , \42503 );
buf \U$39342 ( \49530 , \49529_nG18d84 );
buf \U$39343 ( \49531 , RIb87eb78_68);
_HMUX g16c0f ( \49532_nG16c0f , RIe115a18_5294 , \49531 , \49507 );
_HMUX g16c10 ( \49533_nG16c10 , RIe115a18_5294 , \49532_nG16c0f , \49514 );
buf \U$39344 ( \49534 , RIb7c59f8_236);
_HMUX g16c11 ( \49535_nG16c11 , RIe115a18_5294 , \49534 , \49519 );
_HMUX g16c12 ( \49536_nG16c12 , \49533_nG16c10 , \49535_nG16c11 , \49526 );
buf \U$39345 ( \49537 , \49536_nG16c12 );
_DC g18d9a_GF_IsGateDCbyConstraint ( \49538_nG18d9a , \49537 , \42503 );
buf \U$39346 ( \49539 , \49538_nG18d9a );
buf \U$39347 ( \49540 , RIb87ebf0_67);
_HMUX g16c13 ( \49541_nG16c13 , RIe114410_5295 , \49540 , \49507 );
_HMUX g16c14 ( \49542_nG16c14 , RIe114410_5295 , \49541_nG16c13 , \49514 );
buf \U$39348 ( \49543 , RIb7c5a70_235);
_HMUX g16c15 ( \49544_nG16c15 , RIe114410_5295 , \49543 , \49519 );
_HMUX g16c16 ( \49545_nG16c16 , \49542_nG16c14 , \49544_nG16c15 , \49526 );
buf \U$39349 ( \49546 , \49545_nG16c16 );
_DC g18db0_GF_IsGateDCbyConstraint ( \49547_nG18db0 , \49546 , \42503 );
buf \U$39350 ( \49548 , \49547_nG18db0 );
buf \U$39351 ( \49549 , RIb882ca0_66);
_HMUX g16c17 ( \49550_nG16c17 , RIe1132b8_5296 , \49549 , \49507 );
_HMUX g16c18 ( \49551_nG16c18 , RIe1132b8_5296 , \49550_nG16c17 , \49514 );
buf \U$39352 ( \49552 , RIb7cade0_234);
_HMUX g16c19 ( \49553_nG16c19 , RIe1132b8_5296 , \49552 , \49519 );
_HMUX g16c1a ( \49554_nG16c1a , \49551_nG16c18 , \49553_nG16c19 , \49526 );
buf \U$39353 ( \49555 , \49554_nG16c1a );
_DC g18dc6_GF_IsGateDCbyConstraint ( \49556_nG18dc6 , \49555 , \42503 );
buf \U$39354 ( \49557 , \49556_nG18dc6 );
buf \U$39355 ( \49558 , RIb885310_65);
_HMUX g16c1b ( \49559_nG16c1b , RIe111cb0_5297 , \49558 , \49507 );
_HMUX g16c1c ( \49560_nG16c1c , RIe111cb0_5297 , \49559_nG16c1b , \49514 );
buf \U$39356 ( \49561 , RIb7cae58_233);
_HMUX g16c1d ( \49562_nG16c1d , RIe111cb0_5297 , \49561 , \49519 );
_HMUX g16c1e ( \49563_nG16c1e , \49560_nG16c1c , \49562_nG16c1d , \49526 );
buf \U$39357 ( \49564 , \49563_nG16c1e );
_DC g18ddc_GF_IsGateDCbyConstraint ( \49565_nG18ddc , \49564 , \42503 );
buf \U$39358 ( \49566 , \49565_nG18ddc );
buf \U$39359 ( \49567 , RIb885388_64);
_HMUX g16c1f ( \49568_nG16c1f , RIe110b58_5298 , \49567 , \49507 );
_HMUX g16c20 ( \49569_nG16c20 , RIe110b58_5298 , \49568_nG16c1f , \49514 );
buf \U$39360 ( \49570 , RIb7caed0_232);
_HMUX g16c21 ( \49571_nG16c21 , RIe110b58_5298 , \49570 , \49519 );
_HMUX g16c22 ( \49572_nG16c22 , \49569_nG16c20 , \49571_nG16c21 , \49526 );
buf \U$39361 ( \49573 , \49572_nG16c22 );
_DC g18df2_GF_IsGateDCbyConstraint ( \49574_nG18df2 , \49573 , \42503 );
buf \U$39362 ( \49575 , \49574_nG18df2 );
buf \U$39363 ( \49576 , RIb885400_63);
_HMUX g16c23 ( \49577_nG16c23 , RIe10f550_5299 , \49576 , \49507 );
_HMUX g16c24 ( \49578_nG16c24 , RIe10f550_5299 , \49577_nG16c23 , \49514 );
buf \U$39364 ( \49579 , RIb7caf48_231);
_HMUX g16c25 ( \49580_nG16c25 , RIe10f550_5299 , \49579 , \49519 );
_HMUX g16c26 ( \49581_nG16c26 , \49578_nG16c24 , \49580_nG16c25 , \49526 );
buf \U$39365 ( \49582 , \49581_nG16c26 );
_DC g18dfe_GF_IsGateDCbyConstraint ( \49583_nG18dfe , \49582 , \42503 );
buf \U$39366 ( \49584 , \49583_nG18dfe );
buf \U$39367 ( \49585 , RIb885478_62);
_HMUX g16c27 ( \49586_nG16c27 , RIe10e3f8_5300 , \49585 , \49507 );
_HMUX g16c28 ( \49587_nG16c28 , RIe10e3f8_5300 , \49586_nG16c27 , \49514 );
buf \U$39368 ( \49588 , RIb7cafc0_230);
_HMUX g16c29 ( \49589_nG16c29 , RIe10e3f8_5300 , \49588 , \49519 );
_HMUX g16c2a ( \49590_nG16c2a , \49587_nG16c28 , \49589_nG16c29 , \49526 );
buf \U$39369 ( \49591 , \49590_nG16c2a );
_DC g18e00_GF_IsGateDCbyConstraint ( \49592_nG18e00 , \49591 , \42503 );
buf \U$39370 ( \49593 , \49592_nG18e00 );
buf \U$39371 ( \49594 , RIb8854f0_61);
_HMUX g16c2b ( \49595_nG16c2b , RIe10d2a0_5301 , \49594 , \49507 );
_HMUX g16c2c ( \49596_nG16c2c , RIe10d2a0_5301 , \49595_nG16c2b , \49514 );
buf \U$39372 ( \49597 , RIb7cb038_229);
_HMUX g16c2d ( \49598_nG16c2d , RIe10d2a0_5301 , \49597 , \49519 );
_HMUX g16c2e ( \49599_nG16c2e , \49596_nG16c2c , \49598_nG16c2d , \49526 );
buf \U$39373 ( \49600 , \49599_nG16c2e );
_DC g18e02_GF_IsGateDCbyConstraint ( \49601_nG18e02 , \49600 , \42503 );
buf \U$39374 ( \49602 , \49601_nG18e02 );
buf \U$39375 ( \49603 , RIb885568_60);
_HMUX g16c2f ( \49604_nG16c2f , RIe10bc98_5302 , \49603 , \49507 );
_HMUX g16c30 ( \49605_nG16c30 , RIe10bc98_5302 , \49604_nG16c2f , \49514 );
buf \U$39376 ( \49606 , RIb7cb0b0_228);
_HMUX g16c31 ( \49607_nG16c31 , RIe10bc98_5302 , \49606 , \49519 );
_HMUX g16c32 ( \49608_nG16c32 , \49605_nG16c30 , \49607_nG16c31 , \49526 );
buf \U$39377 ( \49609 , \49608_nG16c32 );
_DC g18d86_GF_IsGateDCbyConstraint ( \49610_nG18d86 , \49609 , \42503 );
buf \U$39378 ( \49611 , \49610_nG18d86 );
buf \U$39379 ( \49612 , RIb8855e0_59);
_HMUX g16c33 ( \49613_nG16c33 , RIe10ab40_5303 , \49612 , \49507 );
_HMUX g16c34 ( \49614_nG16c34 , RIe10ab40_5303 , \49613_nG16c33 , \49514 );
buf \U$39380 ( \49615 , RIb7cb128_227);
_HMUX g16c35 ( \49616_nG16c35 , RIe10ab40_5303 , \49615 , \49519 );
_HMUX g16c36 ( \49617_nG16c36 , \49614_nG16c34 , \49616_nG16c35 , \49526 );
buf \U$39381 ( \49618 , \49617_nG16c36 );
_DC g18d88_GF_IsGateDCbyConstraint ( \49619_nG18d88 , \49618 , \42503 );
buf \U$39382 ( \49620 , \49619_nG18d88 );
buf \U$39383 ( \49621 , RIb885658_58);
_HMUX g16c37 ( \49622_nG16c37 , RIe109538_5304 , \49621 , \49507 );
_HMUX g16c38 ( \49623_nG16c38 , RIe109538_5304 , \49622_nG16c37 , \49514 );
buf \U$39384 ( \49624 , RIb7d00d8_226);
_HMUX g16c39 ( \49625_nG16c39 , RIe109538_5304 , \49624 , \49519 );
_HMUX g16c3a ( \49626_nG16c3a , \49623_nG16c38 , \49625_nG16c39 , \49526 );
buf \U$39385 ( \49627 , \49626_nG16c3a );
_DC g18d8a_GF_IsGateDCbyConstraint ( \49628_nG18d8a , \49627 , \42503 );
buf \U$39386 ( \49629 , \49628_nG18d8a );
buf \U$39387 ( \49630 , RIb8856d0_57);
_HMUX g16c3b ( \49631_nG16c3b , RIe1083e0_5305 , \49630 , \49507 );
_HMUX g16c3c ( \49632_nG16c3c , RIe1083e0_5305 , \49631_nG16c3b , \49514 );
buf \U$39388 ( \49633 , RIb8263d8_225);
_HMUX g16c3d ( \49634_nG16c3d , RIe1083e0_5305 , \49633 , \49519 );
_HMUX g16c3e ( \49635_nG16c3e , \49632_nG16c3c , \49634_nG16c3d , \49526 );
buf \U$39389 ( \49636 , \49635_nG16c3e );
_DC g18d8c_GF_IsGateDCbyConstraint ( \49637_nG18d8c , \49636 , \42503 );
buf \U$39390 ( \49638 , \49637_nG18d8c );
buf \U$39391 ( \49639 , RIb885748_56);
_HMUX g16c3f ( \49640_nG16c3f , RIe106dd8_5306 , \49639 , \49507 );
_HMUX g16c40 ( \49641_nG16c40 , RIe106dd8_5306 , \49640_nG16c3f , \49514 );
buf \U$39392 ( \49642 , RIb826e28_224);
_HMUX g16c41 ( \49643_nG16c41 , RIe106dd8_5306 , \49642 , \49519 );
_HMUX g16c42 ( \49644_nG16c42 , \49641_nG16c40 , \49643_nG16c41 , \49526 );
buf \U$39393 ( \49645 , \49644_nG16c42 );
_DC g18d8e_GF_IsGateDCbyConstraint ( \49646_nG18d8e , \49645 , \42503 );
buf \U$39394 ( \49647 , \49646_nG18d8e );
buf \U$39395 ( \49648 , RIb8857c0_55);
_HMUX g16c43 ( \49649_nG16c43 , RIdfd3728_5307 , \49648 , \49507 );
_HMUX g16c44 ( \49650_nG16c44 , RIdfd3728_5307 , \49649_nG16c43 , \49514 );
buf \U$39396 ( \49651 , RIb826ea0_223);
_HMUX g16c45 ( \49652_nG16c45 , RIdfd3728_5307 , \49651 , \49519 );
_HMUX g16c46 ( \49653_nG16c46 , \49650_nG16c44 , \49652_nG16c45 , \49526 );
buf \U$39397 ( \49654 , \49653_nG16c46 );
_DC g18d90_GF_IsGateDCbyConstraint ( \49655_nG18d90 , \49654 , \42503 );
buf \U$39398 ( \49656 , \49655_nG18d90 );
buf \U$39399 ( \49657 , RIb885838_54);
_HMUX g16c47 ( \49658_nG16c47 , RIdfd71c0_5308 , \49657 , \49507 );
_HMUX g16c48 ( \49659_nG16c48 , RIdfd71c0_5308 , \49658_nG16c47 , \49514 );
buf \U$39400 ( \49660 , RIb826f18_222);
_HMUX g16c49 ( \49661_nG16c49 , RIdfd71c0_5308 , \49660 , \49519 );
_HMUX g16c4a ( \49662_nG16c4a , \49659_nG16c48 , \49661_nG16c49 , \49526 );
buf \U$39401 ( \49663 , \49662_nG16c4a );
_DC g18d92_GF_IsGateDCbyConstraint ( \49664_nG18d92 , \49663 , \42503 );
buf \U$39402 ( \49665 , \49664_nG18d92 );
buf \U$39403 ( \49666 , RIb8858b0_53);
_HMUX g16c4b ( \49667_nG16c4b , RIdfdc8f0_5309 , \49666 , \49507 );
_HMUX g16c4c ( \49668_nG16c4c , RIdfdc8f0_5309 , \49667_nG16c4b , \49514 );
buf \U$39404 ( \49669 , RIb826f90_221);
_HMUX g16c4d ( \49670_nG16c4d , RIdfdc8f0_5309 , \49669 , \49519 );
_HMUX g16c4e ( \49671_nG16c4e , \49668_nG16c4c , \49670_nG16c4d , \49526 );
buf \U$39405 ( \49672 , \49671_nG16c4e );
_DC g18d94_GF_IsGateDCbyConstraint ( \49673_nG18d94 , \49672 , \42503 );
buf \U$39406 ( \49674 , \49673_nG18d94 );
buf \U$39407 ( \49675 , RIb885928_52);
_HMUX g16c4f ( \49676_nG16c4f , RIdfe0b80_5310 , \49675 , \49507 );
_HMUX g16c50 ( \49677_nG16c50 , RIdfe0b80_5310 , \49676_nG16c4f , \49514 );
buf \U$39408 ( \49678 , RIb8293a8_220);
_HMUX g16c51 ( \49679_nG16c51 , RIdfe0b80_5310 , \49678 , \49519 );
_HMUX g16c52 ( \49680_nG16c52 , \49677_nG16c50 , \49679_nG16c51 , \49526 );
buf \U$39409 ( \49681 , \49680_nG16c52 );
_DC g18d96_GF_IsGateDCbyConstraint ( \49682_nG18d96 , \49681 , \42503 );
buf \U$39410 ( \49683 , \49682_nG18d96 );
buf \U$39411 ( \49684 , RIb8859a0_51);
_HMUX g16c53 ( \49685_nG16c53 , RIdfe6760_5311 , \49684 , \49507 );
_HMUX g16c54 ( \49686_nG16c54 , RIdfe6760_5311 , \49685_nG16c53 , \49514 );
buf \U$39412 ( \49687 , RIb829420_219);
_HMUX g16c55 ( \49688_nG16c55 , RIdfe6760_5311 , \49687 , \49519 );
_HMUX g16c56 ( \49689_nG16c56 , \49686_nG16c54 , \49688_nG16c55 , \49526 );
buf \U$39413 ( \49690 , \49689_nG16c56 );
_DC g18d98_GF_IsGateDCbyConstraint ( \49691_nG18d98 , \49690 , \42503 );
buf \U$39414 ( \49692 , \49691_nG18d98 );
buf \U$39415 ( \49693 , RIb885a18_50);
_HMUX g16c57 ( \49694_nG16c57 , RIdfeb788_5312 , \49693 , \49507 );
_HMUX g16c58 ( \49695_nG16c58 , RIdfeb788_5312 , \49694_nG16c57 , \49514 );
buf \U$39416 ( \49696 , RIb829498_218);
_HMUX g16c59 ( \49697_nG16c59 , RIdfeb788_5312 , \49696 , \49519 );
_HMUX g16c5a ( \49698_nG16c5a , \49695_nG16c58 , \49697_nG16c59 , \49526 );
buf \U$39417 ( \49699 , \49698_nG16c5a );
_DC g18d9c_GF_IsGateDCbyConstraint ( \49700_nG18d9c , \49699 , \42503 );
buf \U$39418 ( \49701 , \49700_nG18d9c );
buf \U$39419 ( \49702 , RIb885a90_49);
_HMUX g16c5b ( \49703_nG16c5b , RIdff1f98_5313 , \49702 , \49507 );
_HMUX g16c5c ( \49704_nG16c5c , RIdff1f98_5313 , \49703_nG16c5b , \49514 );
buf \U$39420 ( \49705 , RIb829510_217);
_HMUX g16c5d ( \49706_nG16c5d , RIdff1f98_5313 , \49705 , \49519 );
_HMUX g16c5e ( \49707_nG16c5e , \49704_nG16c5c , \49706_nG16c5d , \49526 );
buf \U$39421 ( \49708 , \49707_nG16c5e );
_DC g18d9e_GF_IsGateDCbyConstraint ( \49709_nG18d9e , \49708 , \42503 );
buf \U$39422 ( \49710 , \49709_nG18d9e );
buf \U$39423 ( \49711 , RIb885b08_48);
_HMUX g16c5f ( \49712_nG16c5f , RIdff7f38_5314 , \49711 , \49507 );
_HMUX g16c60 ( \49713_nG16c60 , RIdff7f38_5314 , \49712_nG16c5f , \49514 );
buf \U$39424 ( \49714 , RIb829588_216);
_HMUX g16c61 ( \49715_nG16c61 , RIdff7f38_5314 , \49714 , \49519 );
_HMUX g16c62 ( \49716_nG16c62 , \49713_nG16c60 , \49715_nG16c61 , \49526 );
buf \U$39425 ( \49717 , \49716_nG16c62 );
_DC g18da0_GF_IsGateDCbyConstraint ( \49718_nG18da0 , \49717 , \42503 );
buf \U$39426 ( \49719 , \49718_nG18da0 );
buf \U$39427 ( \49720 , RIb885b80_47);
_HMUX g16c63 ( \49721_nG16c63 , RIdffe400_5315 , \49720 , \49507 );
_HMUX g16c64 ( \49722_nG16c64 , RIdffe400_5315 , \49721_nG16c63 , \49514 );
buf \U$39428 ( \49723 , RIb829600_215);
_HMUX g16c65 ( \49724_nG16c65 , RIdffe400_5315 , \49723 , \49519 );
_HMUX g16c66 ( \49725_nG16c66 , \49722_nG16c64 , \49724_nG16c65 , \49526 );
buf \U$39429 ( \49726 , \49725_nG16c66 );
_DC g18da2_GF_IsGateDCbyConstraint ( \49727_nG18da2 , \49726 , \42503 );
buf \U$39430 ( \49728 , \49727_nG18da2 );
buf \U$39431 ( \49729 , RIb885bf8_46);
_HMUX g16c67 ( \49730_nG16c67 , RIe005750_5316 , \49729 , \49507 );
_HMUX g16c68 ( \49731_nG16c68 , RIe005750_5316 , \49730_nG16c67 , \49514 );
buf \U$39432 ( \49732 , RIb829678_214);
_HMUX g16c69 ( \49733_nG16c69 , RIe005750_5316 , \49732 , \49519 );
_HMUX g16c6a ( \49734_nG16c6a , \49731_nG16c68 , \49733_nG16c69 , \49526 );
buf \U$39433 ( \49735 , \49734_nG16c6a );
_DC g18da4_GF_IsGateDCbyConstraint ( \49736_nG18da4 , \49735 , \42503 );
buf \U$39434 ( \49737 , \49736_nG18da4 );
buf \U$39435 ( \49738 , RIb885c70_45);
_HMUX g16c6b ( \49739_nG16c6b , RIe00b420_5317 , \49738 , \49507 );
_HMUX g16c6c ( \49740_nG16c6c , RIe00b420_5317 , \49739_nG16c6b , \49514 );
buf \U$39436 ( \49741 , RIb8296f0_213);
_HMUX g16c6d ( \49742_nG16c6d , RIe00b420_5317 , \49741 , \49519 );
_HMUX g16c6e ( \49743_nG16c6e , \49740_nG16c6c , \49742_nG16c6d , \49526 );
buf \U$39437 ( \49744 , \49743_nG16c6e );
_DC g18da6_GF_IsGateDCbyConstraint ( \49745_nG18da6 , \49744 , \42503 );
buf \U$39438 ( \49746 , \49745_nG18da6 );
buf \U$39439 ( \49747 , RIb885ce8_44);
_HMUX g16c6f ( \49748_nG16c6f , RIe0132b0_5318 , \49747 , \49507 );
_HMUX g16c70 ( \49749_nG16c70 , RIe0132b0_5318 , \49748_nG16c6f , \49514 );
buf \U$39440 ( \49750 , RIb82dae8_212);
_HMUX g16c71 ( \49751_nG16c71 , RIe0132b0_5318 , \49750 , \49519 );
_HMUX g16c72 ( \49752_nG16c72 , \49749_nG16c70 , \49751_nG16c71 , \49526 );
buf \U$39441 ( \49753 , \49752_nG16c72 );
_DC g18da8_GF_IsGateDCbyConstraint ( \49754_nG18da8 , \49753 , \42503 );
buf \U$39442 ( \49755 , \49754_nG18da8 );
buf \U$39443 ( \49756 , RIb885d60_43);
_HMUX g16c73 ( \49757_nG16c73 , RIe0193b8_5319 , \49756 , \49507 );
_HMUX g16c74 ( \49758_nG16c74 , RIe0193b8_5319 , \49757_nG16c73 , \49514 );
buf \U$39444 ( \49759 , RIb82db60_211);
_HMUX g16c75 ( \49760_nG16c75 , RIe0193b8_5319 , \49759 , \49519 );
_HMUX g16c76 ( \49761_nG16c76 , \49758_nG16c74 , \49760_nG16c75 , \49526 );
buf \U$39445 ( \49762 , \49761_nG16c76 );
_DC g18daa_GF_IsGateDCbyConstraint ( \49763_nG18daa , \49762 , \42503 );
buf \U$39446 ( \49764 , \49763_nG18daa );
buf \U$39447 ( \49765 , RIb885dd8_42);
_HMUX g16c77 ( \49766_nG16c77 , RIe0202d0_5320 , \49765 , \49507 );
_HMUX g16c78 ( \49767_nG16c78 , RIe0202d0_5320 , \49766_nG16c77 , \49514 );
buf \U$39448 ( \49768 , RIb82dbd8_210);
_HMUX g16c79 ( \49769_nG16c79 , RIe0202d0_5320 , \49768 , \49519 );
_HMUX g16c7a ( \49770_nG16c7a , \49767_nG16c78 , \49769_nG16c79 , \49526 );
buf \U$39449 ( \49771 , \49770_nG16c7a );
_DC g18dac_GF_IsGateDCbyConstraint ( \49772_nG18dac , \49771 , \42503 );
buf \U$39450 ( \49773 , \49772_nG18dac );
buf \U$39451 ( \49774 , RIb885e50_41);
_HMUX g16c7b ( \49775_nG16c7b , RIe023de0_5321 , \49774 , \49507 );
_HMUX g16c7c ( \49776_nG16c7c , RIe023de0_5321 , \49775_nG16c7b , \49514 );
buf \U$39452 ( \49777 , RIb82dc50_209);
_HMUX g16c7d ( \49778_nG16c7d , RIe023de0_5321 , \49777 , \49519 );
_HMUX g16c7e ( \49779_nG16c7e , \49776_nG16c7c , \49778_nG16c7d , \49526 );
buf \U$39453 ( \49780 , \49779_nG16c7e );
_DC g18dae_GF_IsGateDCbyConstraint ( \49781_nG18dae , \49780 , \42503 );
buf \U$39454 ( \49782 , \49781_nG18dae );
buf \U$39455 ( \49783 , RIb885ec8_40);
_HMUX g16c7f ( \49784_nG16c7f , RIe027878_5322 , \49783 , \49507 );
_HMUX g16c80 ( \49785_nG16c80 , RIe027878_5322 , \49784_nG16c7f , \49514 );
buf \U$39456 ( \49786 , RIb82dcc8_208);
_HMUX g16c81 ( \49787_nG16c81 , RIe027878_5322 , \49786 , \49519 );
_HMUX g16c82 ( \49788_nG16c82 , \49785_nG16c80 , \49787_nG16c81 , \49526 );
buf \U$39457 ( \49789 , \49788_nG16c82 );
_DC g18db2_GF_IsGateDCbyConstraint ( \49790_nG18db2 , \49789 , \42503 );
buf \U$39458 ( \49791 , \49790_nG18db2 );
buf \U$39459 ( \49792 , RIb885f40_39);
_HMUX g16c83 ( \49793_nG16c83 , RIe02ccd8_5323 , \49792 , \49507 );
_HMUX g16c84 ( \49794_nG16c84 , RIe02ccd8_5323 , \49793_nG16c83 , \49514 );
buf \U$39460 ( \49795 , RIb82dd40_207);
_HMUX g16c85 ( \49796_nG16c85 , RIe02ccd8_5323 , \49795 , \49519 );
_HMUX g16c86 ( \49797_nG16c86 , \49794_nG16c84 , \49796_nG16c85 , \49526 );
buf \U$39461 ( \49798 , \49797_nG16c86 );
_DC g18db4_GF_IsGateDCbyConstraint ( \49799_nG18db4 , \49798 , \42503 );
buf \U$39462 ( \49800 , \49799_nG18db4 );
buf \U$39463 ( \49801 , RIb885fb8_38);
_HMUX g16c87 ( \49802_nG16c87 , RIe0322a0_5324 , \49801 , \49507 );
_HMUX g16c88 ( \49803_nG16c88 , RIe0322a0_5324 , \49802_nG16c87 , \49514 );
buf \U$39464 ( \49804 , RIb82ddb8_206);
_HMUX g16c89 ( \49805_nG16c89 , RIe0322a0_5324 , \49804 , \49519 );
_HMUX g16c8a ( \49806_nG16c8a , \49803_nG16c88 , \49805_nG16c89 , \49526 );
buf \U$39465 ( \49807 , \49806_nG16c8a );
_DC g18db6_GF_IsGateDCbyConstraint ( \49808_nG18db6 , \49807 , \42503 );
buf \U$39466 ( \49809 , \49808_nG18db6 );
buf \U$39467 ( \49810 , RIb886030_37);
_HMUX g16c8b ( \49811_nG16c8b , RIe038768_5325 , \49810 , \49507 );
_HMUX g16c8c ( \49812_nG16c8c , RIe038768_5325 , \49811_nG16c8b , \49514 );
buf \U$39468 ( \49813 , RIb82de30_205);
_HMUX g16c8d ( \49814_nG16c8d , RIe038768_5325 , \49813 , \49519 );
_HMUX g16c8e ( \49815_nG16c8e , \49812_nG16c8c , \49814_nG16c8d , \49526 );
buf \U$39469 ( \49816 , \49815_nG16c8e );
_DC g18db8_GF_IsGateDCbyConstraint ( \49817_nG18db8 , \49816 , \42503 );
buf \U$39470 ( \49818 , \49817_nG18db8 );
buf \U$39471 ( \49819 , RIb8860a8_36);
_HMUX g16c8f ( \49820_nG16c8f , RIe03c728_5326 , \49819 , \49507 );
_HMUX g16c90 ( \49821_nG16c90 , RIe03c728_5326 , \49820_nG16c8f , \49514 );
buf \U$39472 ( \49822 , RIb832228_204);
_HMUX g16c91 ( \49823_nG16c91 , RIe03c728_5326 , \49822 , \49519 );
_HMUX g16c92 ( \49824_nG16c92 , \49821_nG16c90 , \49823_nG16c91 , \49526 );
buf \U$39473 ( \49825 , \49824_nG16c92 );
_DC g18dba_GF_IsGateDCbyConstraint ( \49826_nG18dba , \49825 , \42503 );
buf \U$39474 ( \49827 , \49826_nG18dba );
buf \U$39475 ( \49828 , RIb886120_35);
_HMUX g16c93 ( \49829_nG16c93 , RIde01258_5327 , \49828 , \49507 );
_HMUX g16c94 ( \49830_nG16c94 , RIde01258_5327 , \49829_nG16c93 , \49514 );
buf \U$39476 ( \49831 , RIb8322a0_203);
_HMUX g16c95 ( \49832_nG16c95 , RIde01258_5327 , \49831 , \49519 );
_HMUX g16c96 ( \49833_nG16c96 , \49830_nG16c94 , \49832_nG16c95 , \49526 );
buf \U$39477 ( \49834 , \49833_nG16c96 );
_DC g18dbc_GF_IsGateDCbyConstraint ( \49835_nG18dbc , \49834 , \42503 );
buf \U$39478 ( \49836 , \49835_nG18dbc );
buf \U$39479 ( \49837 , RIb886198_34);
_HMUX g16c97 ( \49838_nG16c97 , RIddfd748_5328 , \49837 , \49507 );
_HMUX g16c98 ( \49839_nG16c98 , RIddfd748_5328 , \49838_nG16c97 , \49514 );
buf \U$39480 ( \49840 , RIb832318_202);
_HMUX g16c99 ( \49841_nG16c99 , RIddfd748_5328 , \49840 , \49519 );
_HMUX g16c9a ( \49842_nG16c9a , \49839_nG16c98 , \49841_nG16c99 , \49526 );
buf \U$39481 ( \49843 , \49842_nG16c9a );
_DC g18dbe_GF_IsGateDCbyConstraint ( \49844_nG18dbe , \49843 , \42503 );
buf \U$39482 ( \49845 , \49844_nG18dbe );
buf \U$39483 ( \49846 , RIb886210_33);
_HMUX g16c9b ( \49847_nG16c9b , RIddf9788_5329 , \49846 , \49507 );
_HMUX g16c9c ( \49848_nG16c9c , RIddf9788_5329 , \49847_nG16c9b , \49514 );
buf \U$39484 ( \49849 , RIb832390_201);
_HMUX g16c9d ( \49850_nG16c9d , RIddf9788_5329 , \49849 , \49519 );
_HMUX g16c9e ( \49851_nG16c9e , \49848_nG16c9c , \49850_nG16c9d , \49526 );
buf \U$39485 ( \49852 , \49851_nG16c9e );
_DC g18dc0_GF_IsGateDCbyConstraint ( \49853_nG18dc0 , \49852 , \42503 );
buf \U$39486 ( \49854 , \49853_nG18dc0 );
buf \U$39487 ( \49855 , RIb886288_32);
_HMUX g16c9f ( \49856_nG16c9f , RIddf3d88_5330 , \49855 , \49507 );
_HMUX g16ca0 ( \49857_nG16ca0 , RIddf3d88_5330 , \49856_nG16c9f , \49514 );
buf \U$39488 ( \49858 , RIb832408_200);
_HMUX g16ca1 ( \49859_nG16ca1 , RIddf3d88_5330 , \49858 , \49519 );
_HMUX g16ca2 ( \49860_nG16ca2 , \49857_nG16ca0 , \49859_nG16ca1 , \49526 );
buf \U$39489 ( \49861 , \49860_nG16ca2 );
_DC g18dc2_GF_IsGateDCbyConstraint ( \49862_nG18dc2 , \49861 , \42503 );
buf \U$39490 ( \49863 , \49862_nG18dc2 );
buf \U$39491 ( \49864 , RIb886300_31);
_HMUX g16ca3 ( \49865_nG16ca3 , RIdfba228_5331 , \49864 , \49507 );
_HMUX g16ca4 ( \49866_nG16ca4 , RIdfba228_5331 , \49865_nG16ca3 , \49514 );
buf \U$39492 ( \49867 , RIb832480_199);
_HMUX g16ca5 ( \49868_nG16ca5 , RIdfba228_5331 , \49867 , \49519 );
_HMUX g16ca6 ( \49869_nG16ca6 , \49866_nG16ca4 , \49868_nG16ca5 , \49526 );
buf \U$39493 ( \49870 , \49869_nG16ca6 );
_DC g18dc4_GF_IsGateDCbyConstraint ( \49871_nG18dc4 , \49870 , \42503 );
buf \U$39494 ( \49872 , \49871_nG18dc4 );
buf \U$39495 ( \49873 , RIb886378_30);
_HMUX g16ca7 ( \49874_nG16ca7 , RIdfb5e30_5332 , \49873 , \49507 );
_HMUX g16ca8 ( \49875_nG16ca8 , RIdfb5e30_5332 , \49874_nG16ca7 , \49514 );
buf \U$39496 ( \49876 , RIb8324f8_198);
_HMUX g16ca9 ( \49877_nG16ca9 , RIdfb5e30_5332 , \49876 , \49519 );
_HMUX g16caa ( \49878_nG16caa , \49875_nG16ca8 , \49877_nG16ca9 , \49526 );
buf \U$39497 ( \49879 , \49878_nG16caa );
_DC g18dc8_GF_IsGateDCbyConstraint ( \49880_nG18dc8 , \49879 , \42503 );
buf \U$39498 ( \49881 , \49880_nG18dc8 );
buf \U$39499 ( \49882 , RIb8863f0_29);
_HMUX g16cab ( \49883_nG16cab , RIdfb2aa0_5333 , \49882 , \49507 );
_HMUX g16cac ( \49884_nG16cac , RIdfb2aa0_5333 , \49883_nG16cab , \49514 );
buf \U$39500 ( \49885 , RIb832570_197);
_HMUX g16cad ( \49886_nG16cad , RIdfb2aa0_5333 , \49885 , \49519 );
_HMUX g16cae ( \49887_nG16cae , \49884_nG16cac , \49886_nG16cad , \49526 );
buf \U$39501 ( \49888 , \49887_nG16cae );
_DC g18dca_GF_IsGateDCbyConstraint ( \49889_nG18dca , \49888 , \42503 );
buf \U$39502 ( \49890 , \49889_nG18dca );
buf \U$39503 ( \49891 , RIb886468_28);
_HMUX g16caf ( \49892_nG16caf , RIdfaec48_5334 , \49891 , \49507 );
_HMUX g16cb0 ( \49893_nG16cb0 , RIdfaec48_5334 , \49892_nG16caf , \49514 );
buf \U$39504 ( \49894 , RIb8383a8_196);
_HMUX g16cb1 ( \49895_nG16cb1 , RIdfaec48_5334 , \49894 , \49519 );
_HMUX g16cb2 ( \49896_nG16cb2 , \49893_nG16cb0 , \49895_nG16cb1 , \49526 );
buf \U$39505 ( \49897 , \49896_nG16cb2 );
_DC g18dcc_GF_IsGateDCbyConstraint ( \49898_nG18dcc , \49897 , \42503 );
buf \U$39506 ( \49899 , \49898_nG18dcc );
buf \U$39507 ( \49900 , RIb8864e0_27);
_HMUX g16cb3 ( \49901_nG16cb3 , RIdfabf48_5335 , \49900 , \49507 );
_HMUX g16cb4 ( \49902_nG16cb4 , RIdfabf48_5335 , \49901_nG16cb3 , \49514 );
buf \U$39508 ( \49903 , RIb838420_195);
_HMUX g16cb5 ( \49904_nG16cb5 , RIdfabf48_5335 , \49903 , \49519 );
_HMUX g16cb6 ( \49905_nG16cb6 , \49902_nG16cb4 , \49904_nG16cb5 , \49526 );
buf \U$39509 ( \49906 , \49905_nG16cb6 );
_DC g18dce_GF_IsGateDCbyConstraint ( \49907_nG18dce , \49906 , \42503 );
buf \U$39510 ( \49908 , \49907_nG18dce );
buf \U$39511 ( \49909 , RIb886558_26);
_HMUX g16cb7 ( \49910_nG16cb7 , RIdfa97e8_5336 , \49909 , \49507 );
_HMUX g16cb8 ( \49911_nG16cb8 , RIdfa97e8_5336 , \49910_nG16cb7 , \49514 );
buf \U$39512 ( \49912 , RIb838498_194);
_HMUX g16cb9 ( \49913_nG16cb9 , RIdfa97e8_5336 , \49912 , \49519 );
_HMUX g16cba ( \49914_nG16cba , \49911_nG16cb8 , \49913_nG16cb9 , \49526 );
buf \U$39513 ( \49915 , \49914_nG16cba );
_DC g18dd0_GF_IsGateDCbyConstraint ( \49916_nG18dd0 , \49915 , \42503 );
buf \U$39514 ( \49917 , \49916_nG18dd0 );
buf \U$39515 ( \49918 , RIb8865d0_25);
_HMUX g16cbb ( \49919_nG16cbb , RIdfa5e40_5337 , \49918 , \49507 );
_HMUX g16cbc ( \49920_nG16cbc , RIdfa5e40_5337 , \49919_nG16cbb , \49514 );
buf \U$39516 ( \49921 , RIb838510_193);
_HMUX g16cbd ( \49922_nG16cbd , RIdfa5e40_5337 , \49921 , \49519 );
_HMUX g16cbe ( \49923_nG16cbe , \49920_nG16cbc , \49922_nG16cbd , \49526 );
buf \U$39517 ( \49924 , \49923_nG16cbe );
_DC g18dd2_GF_IsGateDCbyConstraint ( \49925_nG18dd2 , \49924 , \42503 );
buf \U$39518 ( \49926 , \49925_nG18dd2 );
buf \U$39519 ( \49927 , RIb886648_24);
_HMUX g16cbf ( \49928_nG16cbf , RIdfa2f60_5338 , \49927 , \49507 );
_HMUX g16cc0 ( \49929_nG16cc0 , RIdfa2f60_5338 , \49928_nG16cbf , \49514 );
buf \U$39520 ( \49930 , RIb838588_192);
_HMUX g16cc1 ( \49931_nG16cc1 , RIdfa2f60_5338 , \49930 , \49519 );
_HMUX g16cc2 ( \49932_nG16cc2 , \49929_nG16cc0 , \49931_nG16cc1 , \49526 );
buf \U$39521 ( \49933 , \49932_nG16cc2 );
_DC g18dd4_GF_IsGateDCbyConstraint ( \49934_nG18dd4 , \49933 , \42503 );
buf \U$39522 ( \49935 , \49934_nG18dd4 );
buf \U$39523 ( \49936 , RIb8866c0_23);
_HMUX g16cc3 ( \49937_nG16cc3 , RIdf9e4d8_5339 , \49936 , \49507 );
_HMUX g16cc4 ( \49938_nG16cc4 , RIdf9e4d8_5339 , \49937_nG16cc3 , \49514 );
buf \U$39524 ( \49939 , RIb838600_191);
_HMUX g16cc5 ( \49940_nG16cc5 , RIdf9e4d8_5339 , \49939 , \49519 );
_HMUX g16cc6 ( \49941_nG16cc6 , \49938_nG16cc4 , \49940_nG16cc5 , \49526 );
buf \U$39525 ( \49942 , \49941_nG16cc6 );
_DC g18dd6_GF_IsGateDCbyConstraint ( \49943_nG18dd6 , \49942 , \42503 );
buf \U$39526 ( \49944 , \49943_nG18dd6 );
buf \U$39527 ( \49945 , RIb886738_22);
_HMUX g16cc7 ( \49946_nG16cc7 , RIdf99618_5340 , \49945 , \49507 );
_HMUX g16cc8 ( \49947_nG16cc8 , RIdf99618_5340 , \49946_nG16cc7 , \49514 );
buf \U$39528 ( \49948 , RIb838678_190);
_HMUX g16cc9 ( \49949_nG16cc9 , RIdf99618_5340 , \49948 , \49519 );
_HMUX g16cca ( \49950_nG16cca , \49947_nG16cc8 , \49949_nG16cc9 , \49526 );
buf \U$39529 ( \49951 , \49950_nG16cca );
_DC g18dd8_GF_IsGateDCbyConstraint ( \49952_nG18dd8 , \49951 , \42503 );
buf \U$39530 ( \49953 , \49952_nG18dd8 );
buf \U$39531 ( \49954 , RIb8867b0_21);
_HMUX g16ccb ( \49955_nG16ccb , RIdf90f90_5341 , \49954 , \49507 );
_HMUX g16ccc ( \49956_nG16ccc , RIdf90f90_5341 , \49955_nG16ccb , \49514 );
buf \U$39532 ( \49957 , RIb8386f0_189);
_HMUX g16ccd ( \49958_nG16ccd , RIdf90f90_5341 , \49957 , \49519 );
_HMUX g16cce ( \49959_nG16cce , \49956_nG16ccc , \49958_nG16ccd , \49526 );
buf \U$39533 ( \49960 , \49959_nG16cce );
_DC g18dda_GF_IsGateDCbyConstraint ( \49961_nG18dda , \49960 , \42503 );
buf \U$39534 ( \49962 , \49961_nG18dda );
buf \U$39535 ( \49963 , RIb886828_20);
_HMUX g16ccf ( \49964_nG16ccf , RIdf8ae88_5342 , \49963 , \49507 );
_HMUX g16cd0 ( \49965_nG16cd0 , RIdf8ae88_5342 , \49964_nG16ccf , \49514 );
buf \U$39536 ( \49966 , RIb838768_188);
_HMUX g16cd1 ( \49967_nG16cd1 , RIdf8ae88_5342 , \49966 , \49519 );
_HMUX g16cd2 ( \49968_nG16cd2 , \49965_nG16cd0 , \49967_nG16cd1 , \49526 );
buf \U$39537 ( \49969 , \49968_nG16cd2 );
_DC g18dde_GF_IsGateDCbyConstraint ( \49970_nG18dde , \49969 , \42503 );
buf \U$39538 ( \49971 , \49970_nG18dde );
buf \U$39539 ( \49972 , RIb8868a0_19);
_HMUX g16cd3 ( \49973_nG16cd3 , RIdf848d0_5343 , \49972 , \49507 );
_HMUX g16cd4 ( \49974_nG16cd4 , RIdf848d0_5343 , \49973_nG16cd3 , \49514 );
buf \U$39540 ( \49975 , RIb8387e0_187);
_HMUX g16cd5 ( \49976_nG16cd5 , RIdf848d0_5343 , \49975 , \49519 );
_HMUX g16cd6 ( \49977_nG16cd6 , \49974_nG16cd4 , \49976_nG16cd5 , \49526 );
buf \U$39541 ( \49978 , \49977_nG16cd6 );
_DC g18de0_GF_IsGateDCbyConstraint ( \49979_nG18de0 , \49978 , \42503 );
buf \U$39542 ( \49980 , \49979_nG18de0 );
buf \U$39543 ( \49981 , RIb886918_18);
_HMUX g16cd7 ( \49982_nG16cd7 , RIdf7c248_5344 , \49981 , \49507 );
_HMUX g16cd8 ( \49983_nG16cd8 , RIdf7c248_5344 , \49982_nG16cd7 , \49514 );
buf \U$39544 ( \49984 , RIb838858_186);
_HMUX g16cd9 ( \49985_nG16cd9 , RIdf7c248_5344 , \49984 , \49519 );
_HMUX g16cda ( \49986_nG16cda , \49983_nG16cd8 , \49985_nG16cd9 , \49526 );
buf \U$39545 ( \49987 , \49986_nG16cda );
_DC g18de2_GF_IsGateDCbyConstraint ( \49988_nG18de2 , \49987 , \42503 );
buf \U$39546 ( \49989 , \49988_nG18de2 );
buf \U$39547 ( \49990 , RIb886990_17);
_HMUX g16cdb ( \49991_nG16cdb , RIdf76140_5345 , \49990 , \49507 );
_HMUX g16cdc ( \49992_nG16cdc , RIdf76140_5345 , \49991_nG16cdb , \49514 );
buf \U$39548 ( \49993 , RIb8388d0_185);
_HMUX g16cdd ( \49994_nG16cdd , RIdf76140_5345 , \49993 , \49519 );
_HMUX g16cde ( \49995_nG16cde , \49992_nG16cdc , \49994_nG16cdd , \49526 );
buf \U$39549 ( \49996 , \49995_nG16cde );
_DC g18de4_GF_IsGateDCbyConstraint ( \49997_nG18de4 , \49996 , \42503 );
buf \U$39550 ( \49998 , \49997_nG18de4 );
buf \U$39551 ( \49999 , RIb886a08_16);
_HMUX g16cdf ( \50000_nG16cdf , RIdc56298_5346 , \49999 , \49507 );
_HMUX g16ce0 ( \50001_nG16ce0 , RIdc56298_5346 , \50000_nG16cdf , \49514 );
buf \U$39552 ( \50002 , RIb838948_184);
_HMUX g16ce1 ( \50003_nG16ce1 , RIdc56298_5346 , \50002 , \49519 );
_HMUX g16ce2 ( \50004_nG16ce2 , \50001_nG16ce0 , \50003_nG16ce1 , \49526 );
buf \U$39553 ( \50005 , \50004_nG16ce2 );
_DC g18de6_GF_IsGateDCbyConstraint ( \50006_nG18de6 , \50005 , \42503 );
buf \U$39554 ( \50007 , \50006_nG18de6 );
buf \U$39555 ( \50008 , RIb886a80_15);
_HMUX g16ce3 ( \50009_nG16ce3 , RIdd75f50_5347 , \50008 , \49507 );
_HMUX g16ce4 ( \50010_nG16ce4 , RIdd75f50_5347 , \50009_nG16ce3 , \49514 );
buf \U$39556 ( \50011 , RIb8389c0_183);
_HMUX g16ce5 ( \50012_nG16ce5 , RIdd75f50_5347 , \50011 , \49519 );
_HMUX g16ce6 ( \50013_nG16ce6 , \50010_nG16ce4 , \50012_nG16ce5 , \49526 );
buf \U$39557 ( \50014 , \50013_nG16ce6 );
_DC g18de8_GF_IsGateDCbyConstraint ( \50015_nG18de8 , \50014 , \42503 );
buf \U$39558 ( \50016 , \50015_nG18de8 );
buf \U$39559 ( \50017 , RIb886af8_14);
_HMUX g16ce7 ( \50018_nG16ce7 , RIdd9d6b8_5348 , \50017 , \49507 );
_HMUX g16ce8 ( \50019_nG16ce8 , RIdd9d6b8_5348 , \50018_nG16ce7 , \49514 );
buf \U$39560 ( \50020 , RIb838a38_182);
_HMUX g16ce9 ( \50021_nG16ce9 , RIdd9d6b8_5348 , \50020 , \49519 );
_HMUX g16cea ( \50022_nG16cea , \50019_nG16ce8 , \50021_nG16ce9 , \49526 );
buf \U$39561 ( \50023 , \50022_nG16cea );
_DC g18dea_GF_IsGateDCbyConstraint ( \50024_nG18dea , \50023 , \42503 );
buf \U$39562 ( \50025 , \50024_nG18dea );
buf \U$39563 ( \50026 , RIb886b70_13);
_HMUX g16ceb ( \50027_nG16ceb , RIdb67180_5349 , \50026 , \49507 );
_HMUX g16cec ( \50028_nG16cec , RIdb67180_5349 , \50027_nG16ceb , \49514 );
buf \U$39564 ( \50029 , RIb838ab0_181);
_HMUX g16ced ( \50030_nG16ced , RIdb67180_5349 , \50029 , \49519 );
_HMUX g16cee ( \50031_nG16cee , \50028_nG16cec , \50030_nG16ced , \49526 );
buf \U$39565 ( \50032 , \50031_nG16cee );
_DC g18dec_GF_IsGateDCbyConstraint ( \50033_nG18dec , \50032 , \42503 );
buf \U$39566 ( \50034 , \50033_nG18dec );
buf \U$39567 ( \50035 , RIb886be8_12);
_HMUX g16cef ( \50036_nG16cef , RIdc198c0_5350 , \50035 , \49507 );
_HMUX g16cf0 ( \50037_nG16cf0 , RIdc198c0_5350 , \50036_nG16cef , \49514 );
buf \U$39568 ( \50038 , RIb838b28_180);
_HMUX g16cf1 ( \50039_nG16cf1 , RIdc198c0_5350 , \50038 , \49519 );
_HMUX g16cf2 ( \50040_nG16cf2 , \50037_nG16cf0 , \50039_nG16cf1 , \49526 );
buf \U$39569 ( \50041 , \50040_nG16cf2 );
_DC g18dee_GF_IsGateDCbyConstraint ( \50042_nG18dee , \50041 , \42503 );
buf \U$39570 ( \50043 , \50042_nG18dee );
buf \U$39571 ( \50044 , RIb886c60_11);
_HMUX g16cf3 ( \50045_nG16cf3 , RIdc008e8_5351 , \50044 , \49507 );
_HMUX g16cf4 ( \50046_nG16cf4 , RIdc008e8_5351 , \50045_nG16cf3 , \49514 );
buf \U$39572 ( \50047 , RIb838ba0_179);
_HMUX g16cf5 ( \50048_nG16cf5 , RIdc008e8_5351 , \50047 , \49519 );
_HMUX g16cf6 ( \50049_nG16cf6 , \50046_nG16cf4 , \50048_nG16cf5 , \49526 );
buf \U$39573 ( \50050 , \50049_nG16cf6 );
_DC g18df0_GF_IsGateDCbyConstraint ( \50051_nG18df0 , \50050 , \42503 );
buf \U$39574 ( \50052 , \50051_nG18df0 );
buf \U$39575 ( \50053 , RIb886cd8_10);
_HMUX g16cf7 ( \50054_nG16cf7 , RIdacdc88_5352 , \50053 , \49507 );
_HMUX g16cf8 ( \50055_nG16cf8 , RIdacdc88_5352 , \50054_nG16cf7 , \49514 );
buf \U$39576 ( \50056 , RIb838c18_178);
_HMUX g16cf9 ( \50057_nG16cf9 , RIdacdc88_5352 , \50056 , \49519 );
_HMUX g16cfa ( \50058_nG16cfa , \50055_nG16cf8 , \50057_nG16cf9 , \49526 );
buf \U$39577 ( \50059 , \50058_nG16cfa );
_DC g18df4_GF_IsGateDCbyConstraint ( \50060_nG18df4 , \50059 , \42503 );
buf \U$39578 ( \50061 , \50060_nG18df4 );
buf \U$39579 ( \50062 , RIb886d50_9);
_HMUX g16cfb ( \50063_nG16cfb , RId8fd180_5353 , \50062 , \49507 );
_HMUX g16cfc ( \50064_nG16cfc , RId8fd180_5353 , \50063_nG16cfb , \49514 );
buf \U$39580 ( \50065 , RIb838c90_177);
_HMUX g16cfd ( \50066_nG16cfd , RId8fd180_5353 , \50065 , \49519 );
_HMUX g16cfe ( \50067_nG16cfe , \50064_nG16cfc , \50066_nG16cfd , \49526 );
buf \U$39581 ( \50068 , \50067_nG16cfe );
_DC g18df6_GF_IsGateDCbyConstraint ( \50069_nG18df6 , \50068 , \42503 );
buf \U$39582 ( \50070 , \50069_nG18df6 );
buf \U$39583 ( \50071 , RIb886dc8_8);
_HMUX g16cff ( \50072_nG16cff , RIdb353b0_5354 , \50071 , \49507 );
_HMUX g16d00 ( \50073_nG16d00 , RIdb353b0_5354 , \50072_nG16cff , \49514 );
buf \U$39584 ( \50074 , RIb838d08_176);
_HMUX g16d01 ( \50075_nG16d01 , RIdb353b0_5354 , \50074 , \49519 );
_HMUX g16d02 ( \50076_nG16d02 , \50073_nG16d00 , \50075_nG16d01 , \49526 );
buf \U$39585 ( \50077 , \50076_nG16d02 );
_DC g18df8_GF_IsGateDCbyConstraint ( \50078_nG18df8 , \50077 , \42503 );
buf \U$39586 ( \50079 , \50078_nG18df8 );
buf \U$39587 ( \50080 , RIb886e40_7);
_HMUX g16d03 ( \50081_nG16d03 , RIdbdbca0_5355 , \50080 , \49507 );
_HMUX g16d04 ( \50082_nG16d04 , RIdbdbca0_5355 , \50081_nG16d03 , \49514 );
buf \U$39588 ( \50083 , RIb838d80_175);
_HMUX g16d05 ( \50084_nG16d05 , RIdbdbca0_5355 , \50083 , \49519 );
_HMUX g16d06 ( \50085_nG16d06 , \50082_nG16d04 , \50084_nG16d05 , \49526 );
buf \U$39589 ( \50086 , \50085_nG16d06 );
_DC g18dfa_GF_IsGateDCbyConstraint ( \50087_nG18dfa , \50086 , \42503 );
buf \U$39590 ( \50088 , \50087_nG18dfa );
buf \U$39591 ( \50089 , RIb886eb8_6);
_HMUX g16d07 ( \50090_nG16d07 , RIdb8b8b8_5356 , \50089 , \49507 );
_HMUX g16d08 ( \50091_nG16d08 , RIdb8b8b8_5356 , \50090_nG16d07 , \49514 );
buf \U$39592 ( \50092 , RIb838df8_174);
_HMUX g16d09 ( \50093_nG16d09 , RIdb8b8b8_5356 , \50092 , \49519 );
_HMUX g16d0a ( \50094_nG16d0a , \50091_nG16d08 , \50093_nG16d09 , \49526 );
buf \U$39593 ( \50095 , \50094_nG16d0a );
_DC g18dfc_GF_IsGateDCbyConstraint ( \50096_nG18dfc , \50095 , \42503 );
buf \U$39594 ( \50097 , \50096_nG18dfc );
not \U$39595 ( \50098 , \49506 );
and \U$39596 ( \50099 , \49505 , \50098 );
_HMUX g16b09 ( \50100_nG16b09 , RIddb1a28_5357 , \49504 , \50099 );
_HMUX g16b0a ( \50101_nG16b0a , RIddb1a28_5357 , \50100_nG16b09 , \49514 );
not \U$39597 ( \50102 , \49518 );
and \U$39598 ( \50103 , \49517 , \50102 );
_HMUX g16b0c ( \50104_nG16b0c , RIddb1a28_5357 , \49516 , \50103 );
_HMUX g16b0d ( \50105_nG16b0d , \50101_nG16b0a , \50104_nG16b0c , \49526 );
buf \U$39599 ( \50106 , \50105_nG16b0d );
_DC g18d04_GF_IsGateDCbyConstraint ( \50107_nG18d04 , \50106 , \42503 );
buf \U$39600 ( \50108 , \50107_nG18d04 );
_HMUX g16b0e ( \50109_nG16b0e , RIddc60e0_5358 , \49531 , \50099 );
_HMUX g16b0f ( \50110_nG16b0f , RIddc60e0_5358 , \50109_nG16b0e , \49514 );
_HMUX g16b10 ( \50111_nG16b10 , RIddc60e0_5358 , \49534 , \50103 );
_HMUX g16b11 ( \50112_nG16b11 , \50110_nG16b0f , \50111_nG16b10 , \49526 );
buf \U$39601 ( \50113 , \50112_nG16b11 );
_DC g18d1a_GF_IsGateDCbyConstraint ( \50114_nG18d1a , \50113 , \42503 );
buf \U$39602 ( \50115 , \50114_nG18d1a );
_HMUX g16b12 ( \50116_nG16b12 , RIddd3cb8_5359 , \49540 , \50099 );
_HMUX g16b13 ( \50117_nG16b13 , RIddd3cb8_5359 , \50116_nG16b12 , \49514 );
_HMUX g16b14 ( \50118_nG16b14 , RIddd3cb8_5359 , \49543 , \50103 );
_HMUX g16b15 ( \50119_nG16b15 , \50117_nG16b13 , \50118_nG16b14 , \49526 );
buf \U$39603 ( \50120 , \50119_nG16b15 );
_DC g18d30_GF_IsGateDCbyConstraint ( \50121_nG18d30 , \50120 , \42503 );
buf \U$39604 ( \50122 , \50121_nG18d30 );
_HMUX g16b16 ( \50123_nG16b16 , RIdddeaa0_5360 , \49549 , \50099 );
_HMUX g16b17 ( \50124_nG16b17 , RIdddeaa0_5360 , \50123_nG16b16 , \49514 );
_HMUX g16b18 ( \50125_nG16b18 , RIdddeaa0_5360 , \49552 , \50103 );
_HMUX g16b19 ( \50126_nG16b19 , \50124_nG16b17 , \50125_nG16b18 , \49526 );
buf \U$39605 ( \50127 , \50126_nG16b19 );
_DC g18d46_GF_IsGateDCbyConstraint ( \50128_nG18d46 , \50127 , \42503 );
buf \U$39606 ( \50129 , \50128_nG18d46 );
_HMUX g16b1a ( \50130_nG16b1a , RIdde50d0_5361 , \49558 , \50099 );
_HMUX g16b1b ( \50131_nG16b1b , RIdde50d0_5361 , \50130_nG16b1a , \49514 );
_HMUX g16b1c ( \50132_nG16b1c , RIdde50d0_5361 , \49561 , \50103 );
_HMUX g16b1d ( \50133_nG16b1d , \50131_nG16b1b , \50132_nG16b1c , \49526 );
buf \U$39607 ( \50134 , \50133_nG16b1d );
_DC g18d5c_GF_IsGateDCbyConstraint ( \50135_nG18d5c , \50134 , \42503 );
buf \U$39608 ( \50136 , \50135_nG18d5c );
_HMUX g16b1e ( \50137_nG16b1e , RIddeee50_5362 , \49567 , \50099 );
_HMUX g16b1f ( \50138_nG16b1f , RIddeee50_5362 , \50137_nG16b1e , \49514 );
_HMUX g16b20 ( \50139_nG16b20 , RIddeee50_5362 , \49570 , \50103 );
_HMUX g16b21 ( \50140_nG16b21 , \50138_nG16b1f , \50139_nG16b20 , \49526 );
buf \U$39609 ( \50141 , \50140_nG16b21 );
_DC g18d72_GF_IsGateDCbyConstraint ( \50142_nG18d72 , \50141 , \42503 );
buf \U$39610 ( \50143 , \50142_nG18d72 );
_HMUX g16b22 ( \50144_nG16b22 , RIdc2bb60_5363 , \49576 , \50099 );
_HMUX g16b23 ( \50145_nG16b23 , RIdc2bb60_5363 , \50144_nG16b22 , \49514 );
_HMUX g16b24 ( \50146_nG16b24 , RIdc2bb60_5363 , \49579 , \50103 );
_HMUX g16b25 ( \50147_nG16b25 , \50145_nG16b23 , \50146_nG16b24 , \49526 );
buf \U$39611 ( \50148 , \50147_nG16b25 );
_DC g18d7e_GF_IsGateDCbyConstraint ( \50149_nG18d7e , \50148 , \42503 );
buf \U$39612 ( \50150 , \50149_nG18d7e );
_HMUX g16b26 ( \50151_nG16b26 , RIdc34788_5364 , \49585 , \50099 );
_HMUX g16b27 ( \50152_nG16b27 , RIdc34788_5364 , \50151_nG16b26 , \49514 );
_HMUX g16b28 ( \50153_nG16b28 , RIdc34788_5364 , \49588 , \50103 );
_HMUX g16b29 ( \50154_nG16b29 , \50152_nG16b27 , \50153_nG16b28 , \49526 );
buf \U$39613 ( \50155 , \50154_nG16b29 );
_DC g18d80_GF_IsGateDCbyConstraint ( \50156_nG18d80 , \50155 , \42503 );
buf \U$39614 ( \50157 , \50156_nG18d80 );
_HMUX g16b2a ( \50158_nG16b2a , RIde6e7b8_5365 , \49594 , \50099 );
_HMUX g16b2b ( \50159_nG16b2b , RIde6e7b8_5365 , \50158_nG16b2a , \49514 );
_HMUX g16b2c ( \50160_nG16b2c , RIde6e7b8_5365 , \49597 , \50103 );
_HMUX g16b2d ( \50161_nG16b2d , \50159_nG16b2b , \50160_nG16b2c , \49526 );
buf \U$39615 ( \50162 , \50161_nG16b2d );
_DC g18d82_GF_IsGateDCbyConstraint ( \50163_nG18d82 , \50162 , \42503 );
buf \U$39616 ( \50164 , \50163_nG18d82 );
_HMUX g16b2e ( \50165_nG16b2e , RIde62ad0_5366 , \49603 , \50099 );
_HMUX g16b2f ( \50166_nG16b2f , RIde62ad0_5366 , \50165_nG16b2e , \49514 );
_HMUX g16b30 ( \50167_nG16b30 , RIde62ad0_5366 , \49606 , \50103 );
_HMUX g16b31 ( \50168_nG16b31 , \50166_nG16b2f , \50167_nG16b30 , \49526 );
buf \U$39617 ( \50169 , \50168_nG16b31 );
_DC g18d06_GF_IsGateDCbyConstraint ( \50170_nG18d06 , \50169 , \42503 );
buf \U$39618 ( \50171 , \50170_nG18d06 );
_HMUX g16b32 ( \50172_nG16b32 , RIde55510_5367 , \49612 , \50099 );
_HMUX g16b33 ( \50173_nG16b33 , RIde55510_5367 , \50172_nG16b32 , \49514 );
_HMUX g16b34 ( \50174_nG16b34 , RIde55510_5367 , \49615 , \50103 );
_HMUX g16b35 ( \50175_nG16b35 , \50173_nG16b33 , \50174_nG16b34 , \49526 );
buf \U$39619 ( \50176 , \50175_nG16b35 );
_DC g18d08_GF_IsGateDCbyConstraint ( \50177_nG18d08 , \50176 , \42503 );
buf \U$39620 ( \50178 , \50177_nG18d08 );
_HMUX g16b36 ( \50179_nG16b36 , RIde4a188_5368 , \49621 , \50099 );
_HMUX g16b37 ( \50180_nG16b37 , RIde4a188_5368 , \50179_nG16b36 , \49514 );
_HMUX g16b38 ( \50181_nG16b38 , RIde4a188_5368 , \49624 , \50103 );
_HMUX g16b39 ( \50182_nG16b39 , \50180_nG16b37 , \50181_nG16b38 , \49526 );
buf \U$39621 ( \50183 , \50182_nG16b39 );
_DC g18d0a_GF_IsGateDCbyConstraint ( \50184_nG18d0a , \50183 , \42503 );
buf \U$39622 ( \50185 , \50184_nG18d0a );
_HMUX g16b3a ( \50186_nG16b3a , RIde36d90_5369 , \49630 , \50099 );
_HMUX g16b3b ( \50187_nG16b3b , RIde36d90_5369 , \50186_nG16b3a , \49514 );
_HMUX g16b3c ( \50188_nG16b3c , RIde36d90_5369 , \49633 , \50103 );
_HMUX g16b3d ( \50189_nG16b3d , \50187_nG16b3b , \50188_nG16b3c , \49526 );
buf \U$39623 ( \50190 , \50189_nG16b3d );
_DC g18d0c_GF_IsGateDCbyConstraint ( \50191_nG18d0c , \50190 , \42503 );
buf \U$39624 ( \50192 , \50191_nG18d0c );
_HMUX g16b3e ( \50193_nG16b3e , RIde29c80_5370 , \49639 , \50099 );
_HMUX g16b3f ( \50194_nG16b3f , RIde29c80_5370 , \50193_nG16b3e , \49514 );
_HMUX g16b40 ( \50195_nG16b40 , RIde29c80_5370 , \49642 , \50103 );
_HMUX g16b41 ( \50196_nG16b41 , \50194_nG16b3f , \50195_nG16b40 , \49526 );
buf \U$39625 ( \50197 , \50196_nG16b41 );
_DC g18d0e_GF_IsGateDCbyConstraint ( \50198_nG18d0e , \50197 , \42503 );
buf \U$39626 ( \50199 , \50198_nG18d0e );
_HMUX g16b42 ( \50200_nG16b42 , RIde1c210_5371 , \49648 , \50099 );
_HMUX g16b43 ( \50201_nG16b43 , RIde1c210_5371 , \50200_nG16b42 , \49514 );
_HMUX g16b44 ( \50202_nG16b44 , RIde1c210_5371 , \49651 , \50103 );
_HMUX g16b45 ( \50203_nG16b45 , \50201_nG16b43 , \50202_nG16b44 , \49526 );
buf \U$39627 ( \50204 , \50203_nG16b45 );
_DC g18d10_GF_IsGateDCbyConstraint ( \50205_nG18d10 , \50204 , \42503 );
buf \U$39628 ( \50206 , \50205_nG18d10 );
_HMUX g16b46 ( \50207_nG16b46 , RIde0cb08_5372 , \49657 , \50099 );
_HMUX g16b47 ( \50208_nG16b47 , RIde0cb08_5372 , \50207_nG16b46 , \49514 );
_HMUX g16b48 ( \50209_nG16b48 , RIde0cb08_5372 , \49660 , \50103 );
_HMUX g16b49 ( \50210_nG16b49 , \50208_nG16b47 , \50209_nG16b48 , \49526 );
buf \U$39629 ( \50211 , \50210_nG16b49 );
_DC g18d12_GF_IsGateDCbyConstraint ( \50212_nG18d12 , \50211 , \42503 );
buf \U$39630 ( \50213 , \50212_nG18d12 );
_HMUX g16b4a ( \50214_nG16b4a , RIe03d4c0_5373 , \49666 , \50099 );
_HMUX g16b4b ( \50215_nG16b4b , RIe03d4c0_5373 , \50214_nG16b4a , \49514 );
_HMUX g16b4c ( \50216_nG16b4c , RIe03d4c0_5373 , \49669 , \50103 );
_HMUX g16b4d ( \50217_nG16b4d , \50215_nG16b4b , \50216_nG16b4c , \49526 );
buf \U$39631 ( \50218 , \50217_nG16b4d );
_DC g18d14_GF_IsGateDCbyConstraint ( \50219_nG18d14 , \50218 , \42503 );
buf \U$39632 ( \50220 , \50219_nG18d14 );
_HMUX g16b4e ( \50221_nG16b4e , RIe040b98_5374 , \49675 , \50099 );
_HMUX g16b4f ( \50222_nG16b4f , RIe040b98_5374 , \50221_nG16b4e , \49514 );
_HMUX g16b50 ( \50223_nG16b50 , RIe040b98_5374 , \49678 , \50103 );
_HMUX g16b51 ( \50224_nG16b51 , \50222_nG16b4f , \50223_nG16b50 , \49526 );
buf \U$39633 ( \50225 , \50224_nG16b51 );
_DC g18d16_GF_IsGateDCbyConstraint ( \50226_nG18d16 , \50225 , \42503 );
buf \U$39634 ( \50227 , \50226_nG18d16 );
_HMUX g16b52 ( \50228_nG16b52 , RIe043460_5375 , \49684 , \50099 );
_HMUX g16b53 ( \50229_nG16b53 , RIe043460_5375 , \50228_nG16b52 , \49514 );
_HMUX g16b54 ( \50230_nG16b54 , RIe043460_5375 , \49687 , \50103 );
_HMUX g16b55 ( \50231_nG16b55 , \50229_nG16b53 , \50230_nG16b54 , \49526 );
buf \U$39635 ( \50232 , \50231_nG16b55 );
_DC g18d18_GF_IsGateDCbyConstraint ( \50233_nG18d18 , \50232 , \42503 );
buf \U$39636 ( \50234 , \50233_nG18d18 );
_HMUX g16b56 ( \50235_nG16b56 , RIe046b38_5376 , \49693 , \50099 );
_HMUX g16b57 ( \50236_nG16b57 , RIe046b38_5376 , \50235_nG16b56 , \49514 );
_HMUX g16b58 ( \50237_nG16b58 , RIe046b38_5376 , \49696 , \50103 );
_HMUX g16b59 ( \50238_nG16b59 , \50236_nG16b57 , \50237_nG16b58 , \49526 );
buf \U$39637 ( \50239 , \50238_nG16b59 );
_DC g18d1c_GF_IsGateDCbyConstraint ( \50240_nG18d1c , \50239 , \42503 );
buf \U$39638 ( \50241 , \50240_nG18d1c );
_HMUX g16b5a ( \50242_nG16b5a , RIe049400_5377 , \49702 , \50099 );
_HMUX g16b5b ( \50243_nG16b5b , RIe049400_5377 , \50242_nG16b5a , \49514 );
_HMUX g16b5c ( \50244_nG16b5c , RIe049400_5377 , \49705 , \50103 );
_HMUX g16b5d ( \50245_nG16b5d , \50243_nG16b5b , \50244_nG16b5c , \49526 );
buf \U$39639 ( \50246 , \50245_nG16b5d );
_DC g18d1e_GF_IsGateDCbyConstraint ( \50247_nG18d1e , \50246 , \42503 );
buf \U$39640 ( \50248 , \50247_nG18d1e );
_HMUX g16b5e ( \50249_nG16b5e , RIe04c178_5378 , \49711 , \50099 );
_HMUX g16b5f ( \50250_nG16b5f , RIe04c178_5378 , \50249_nG16b5e , \49514 );
_HMUX g16b60 ( \50251_nG16b60 , RIe04c178_5378 , \49714 , \50103 );
_HMUX g16b61 ( \50252_nG16b61 , \50250_nG16b5f , \50251_nG16b60 , \49526 );
buf \U$39641 ( \50253 , \50252_nG16b61 );
_DC g18d20_GF_IsGateDCbyConstraint ( \50254_nG18d20 , \50253 , \42503 );
buf \U$39642 ( \50255 , \50254_nG18d20 );
_HMUX g16b62 ( \50256_nG16b62 , RIe04f3a0_5379 , \49720 , \50099 );
_HMUX g16b63 ( \50257_nG16b63 , RIe04f3a0_5379 , \50256_nG16b62 , \49514 );
_HMUX g16b64 ( \50258_nG16b64 , RIe04f3a0_5379 , \49723 , \50103 );
_HMUX g16b65 ( \50259_nG16b65 , \50257_nG16b63 , \50258_nG16b64 , \49526 );
buf \U$39643 ( \50260 , \50259_nG16b65 );
_DC g18d22_GF_IsGateDCbyConstraint ( \50261_nG18d22 , \50260 , \42503 );
buf \U$39644 ( \50262 , \50261_nG18d22 );
_HMUX g16b66 ( \50263_nG16b66 , RIe052118_5380 , \49729 , \50099 );
_HMUX g16b67 ( \50264_nG16b67 , RIe052118_5380 , \50263_nG16b66 , \49514 );
_HMUX g16b68 ( \50265_nG16b68 , RIe052118_5380 , \49732 , \50103 );
_HMUX g16b69 ( \50266_nG16b69 , \50264_nG16b67 , \50265_nG16b68 , \49526 );
buf \U$39645 ( \50267 , \50266_nG16b69 );
_DC g18d24_GF_IsGateDCbyConstraint ( \50268_nG18d24 , \50267 , \42503 );
buf \U$39646 ( \50269 , \50268_nG18d24 );
_HMUX g16b6a ( \50270_nG16b6a , RIe055340_5381 , \49738 , \50099 );
_HMUX g16b6b ( \50271_nG16b6b , RIe055340_5381 , \50270_nG16b6a , \49514 );
_HMUX g16b6c ( \50272_nG16b6c , RIe055340_5381 , \49741 , \50103 );
_HMUX g16b6d ( \50273_nG16b6d , \50271_nG16b6b , \50272_nG16b6c , \49526 );
buf \U$39647 ( \50274 , \50273_nG16b6d );
_DC g18d26_GF_IsGateDCbyConstraint ( \50275_nG18d26 , \50274 , \42503 );
buf \U$39648 ( \50276 , \50275_nG18d26 );
_HMUX g16b6e ( \50277_nG16b6e , RIe0580b8_5382 , \49747 , \50099 );
_HMUX g16b6f ( \50278_nG16b6f , RIe0580b8_5382 , \50277_nG16b6e , \49514 );
_HMUX g16b70 ( \50279_nG16b70 , RIe0580b8_5382 , \49750 , \50103 );
_HMUX g16b71 ( \50280_nG16b71 , \50278_nG16b6f , \50279_nG16b70 , \49526 );
buf \U$39649 ( \50281 , \50280_nG16b71 );
_DC g18d28_GF_IsGateDCbyConstraint ( \50282_nG18d28 , \50281 , \42503 );
buf \U$39650 ( \50283 , \50282_nG18d28 );
_HMUX g16b72 ( \50284_nG16b72 , RIe05b2e0_5383 , \49756 , \50099 );
_HMUX g16b73 ( \50285_nG16b73 , RIe05b2e0_5383 , \50284_nG16b72 , \49514 );
_HMUX g16b74 ( \50286_nG16b74 , RIe05b2e0_5383 , \49759 , \50103 );
_HMUX g16b75 ( \50287_nG16b75 , \50285_nG16b73 , \50286_nG16b74 , \49526 );
buf \U$39651 ( \50288 , \50287_nG16b75 );
_DC g18d2a_GF_IsGateDCbyConstraint ( \50289_nG18d2a , \50288 , \42503 );
buf \U$39652 ( \50290 , \50289_nG18d2a );
_HMUX g16b76 ( \50291_nG16b76 , RIe05e058_5384 , \49765 , \50099 );
_HMUX g16b77 ( \50292_nG16b77 , RIe05e058_5384 , \50291_nG16b76 , \49514 );
_HMUX g16b78 ( \50293_nG16b78 , RIe05e058_5384 , \49768 , \50103 );
_HMUX g16b79 ( \50294_nG16b79 , \50292_nG16b77 , \50293_nG16b78 , \49526 );
buf \U$39653 ( \50295 , \50294_nG16b79 );
_DC g18d2c_GF_IsGateDCbyConstraint ( \50296_nG18d2c , \50295 , \42503 );
buf \U$39654 ( \50297 , \50296_nG18d2c );
_HMUX g16b7a ( \50298_nG16b7a , RIe060920_5385 , \49774 , \50099 );
_HMUX g16b7b ( \50299_nG16b7b , RIe060920_5385 , \50298_nG16b7a , \49514 );
_HMUX g16b7c ( \50300_nG16b7c , RIe060920_5385 , \49777 , \50103 );
_HMUX g16b7d ( \50301_nG16b7d , \50299_nG16b7b , \50300_nG16b7c , \49526 );
buf \U$39655 ( \50302 , \50301_nG16b7d );
_DC g18d2e_GF_IsGateDCbyConstraint ( \50303_nG18d2e , \50302 , \42503 );
buf \U$39656 ( \50304 , \50303_nG18d2e );
_HMUX g16b7e ( \50305_nG16b7e , RIe063ff8_5386 , \49783 , \50099 );
_HMUX g16b7f ( \50306_nG16b7f , RIe063ff8_5386 , \50305_nG16b7e , \49514 );
_HMUX g16b80 ( \50307_nG16b80 , RIe063ff8_5386 , \49786 , \50103 );
_HMUX g16b81 ( \50308_nG16b81 , \50306_nG16b7f , \50307_nG16b80 , \49526 );
buf \U$39657 ( \50309 , \50308_nG16b81 );
_DC g18d32_GF_IsGateDCbyConstraint ( \50310_nG18d32 , \50309 , \42503 );
buf \U$39658 ( \50311 , \50310_nG18d32 );
_HMUX g16b82 ( \50312_nG16b82 , RIe0662a8_5387 , \49792 , \50099 );
_HMUX g16b83 ( \50313_nG16b83 , RIe0662a8_5387 , \50312_nG16b82 , \49514 );
_HMUX g16b84 ( \50314_nG16b84 , RIe0662a8_5387 , \49795 , \50103 );
_HMUX g16b85 ( \50315_nG16b85 , \50313_nG16b83 , \50314_nG16b84 , \49526 );
buf \U$39659 ( \50316 , \50315_nG16b85 );
_DC g18d34_GF_IsGateDCbyConstraint ( \50317_nG18d34 , \50316 , \42503 );
buf \U$39660 ( \50318 , \50317_nG18d34 );
_HMUX g16b86 ( \50319_nG16b86 , RIe068288_5388 , \49801 , \50099 );
_HMUX g16b87 ( \50320_nG16b87 , RIe068288_5388 , \50319_nG16b86 , \49514 );
_HMUX g16b88 ( \50321_nG16b88 , RIe068288_5388 , \49804 , \50103 );
_HMUX g16b89 ( \50322_nG16b89 , \50320_nG16b87 , \50321_nG16b88 , \49526 );
buf \U$39661 ( \50323 , \50322_nG16b89 );
_DC g18d36_GF_IsGateDCbyConstraint ( \50324_nG18d36 , \50323 , \42503 );
buf \U$39662 ( \50325 , \50324_nG18d36 );
_HMUX g16b8a ( \50326_nG16b8a , RIe069a70_5389 , \49810 , \50099 );
_HMUX g16b8b ( \50327_nG16b8b , RIe069a70_5389 , \50326_nG16b8a , \49514 );
_HMUX g16b8c ( \50328_nG16b8c , RIe069a70_5389 , \49813 , \50103 );
_HMUX g16b8d ( \50329_nG16b8d , \50327_nG16b8b , \50328_nG16b8c , \49526 );
buf \U$39663 ( \50330 , \50329_nG16b8d );
_DC g18d38_GF_IsGateDCbyConstraint ( \50331_nG18d38 , \50330 , \42503 );
buf \U$39664 ( \50332 , \50331_nG18d38 );
_HMUX g16b8e ( \50333_nG16b8e , RIe06b870_5390 , \49819 , \50099 );
_HMUX g16b8f ( \50334_nG16b8f , RIe06b870_5390 , \50333_nG16b8e , \49514 );
_HMUX g16b90 ( \50335_nG16b90 , RIe06b870_5390 , \49822 , \50103 );
_HMUX g16b91 ( \50336_nG16b91 , \50334_nG16b8f , \50335_nG16b90 , \49526 );
buf \U$39665 ( \50337 , \50336_nG16b91 );
_DC g18d3a_GF_IsGateDCbyConstraint ( \50338_nG18d3a , \50337 , \42503 );
buf \U$39666 ( \50339 , \50338_nG18d3a );
_HMUX g16b92 ( \50340_nG16b92 , RIe06cf68_5391 , \49828 , \50099 );
_HMUX g16b93 ( \50341_nG16b93 , RIe06cf68_5391 , \50340_nG16b92 , \49514 );
_HMUX g16b94 ( \50342_nG16b94 , RIe06cf68_5391 , \49831 , \50103 );
_HMUX g16b95 ( \50343_nG16b95 , \50341_nG16b93 , \50342_nG16b94 , \49526 );
buf \U$39667 ( \50344 , \50343_nG16b95 );
_DC g18d3c_GF_IsGateDCbyConstraint ( \50345_nG18d3c , \50344 , \42503 );
buf \U$39668 ( \50346 , \50345_nG18d3c );
_HMUX g16b96 ( \50347_nG16b96 , RIe06e6d8_5392 , \49837 , \50099 );
_HMUX g16b97 ( \50348_nG16b97 , RIe06e6d8_5392 , \50347_nG16b96 , \49514 );
_HMUX g16b98 ( \50349_nG16b98 , RIe06e6d8_5392 , \49840 , \50103 );
_HMUX g16b99 ( \50350_nG16b99 , \50348_nG16b97 , \50349_nG16b98 , \49526 );
buf \U$39669 ( \50351 , \50350_nG16b99 );
_DC g18d3e_GF_IsGateDCbyConstraint ( \50352_nG18d3e , \50351 , \42503 );
buf \U$39670 ( \50353 , \50352_nG18d3e );
_HMUX g16b9a ( \50354_nG16b9a , RIe06fa10_5393 , \49846 , \50099 );
_HMUX g16b9b ( \50355_nG16b9b , RIe06fa10_5393 , \50354_nG16b9a , \49514 );
_HMUX g16b9c ( \50356_nG16b9c , RIe06fa10_5393 , \49849 , \50103 );
_HMUX g16b9d ( \50357_nG16b9d , \50355_nG16b9b , \50356_nG16b9c , \49526 );
buf \U$39671 ( \50358 , \50357_nG16b9d );
_DC g18d40_GF_IsGateDCbyConstraint ( \50359_nG18d40 , \50358 , \42503 );
buf \U$39672 ( \50360 , \50359_nG18d40 );
_HMUX g16b9e ( \50361_nG16b9e , RIe070eb0_5394 , \49855 , \50099 );
_HMUX g16b9f ( \50362_nG16b9f , RIe070eb0_5394 , \50361_nG16b9e , \49514 );
_HMUX g16ba0 ( \50363_nG16ba0 , RIe070eb0_5394 , \49858 , \50103 );
_HMUX g16ba1 ( \50364_nG16ba1 , \50362_nG16b9f , \50363_nG16ba0 , \49526 );
buf \U$39673 ( \50365 , \50364_nG16ba1 );
_DC g18d42_GF_IsGateDCbyConstraint ( \50366_nG18d42 , \50365 , \42503 );
buf \U$39674 ( \50367 , \50366_nG18d42 );
_HMUX g16ba2 ( \50368_nG16ba2 , RIe0721e8_5395 , \49864 , \50099 );
_HMUX g16ba3 ( \50369_nG16ba3 , RIe0721e8_5395 , \50368_nG16ba2 , \49514 );
_HMUX g16ba4 ( \50370_nG16ba4 , RIe0721e8_5395 , \49867 , \50103 );
_HMUX g16ba5 ( \50371_nG16ba5 , \50369_nG16ba3 , \50370_nG16ba4 , \49526 );
buf \U$39675 ( \50372 , \50371_nG16ba5 );
_DC g18d44_GF_IsGateDCbyConstraint ( \50373_nG18d44 , \50372 , \42503 );
buf \U$39676 ( \50374 , \50373_nG18d44 );
_HMUX g16ba6 ( \50375_nG16ba6 , RIe073808_5396 , \49873 , \50099 );
_HMUX g16ba7 ( \50376_nG16ba7 , RIe073808_5396 , \50375_nG16ba6 , \49514 );
_HMUX g16ba8 ( \50377_nG16ba8 , RIe073808_5396 , \49876 , \50103 );
_HMUX g16ba9 ( \50378_nG16ba9 , \50376_nG16ba7 , \50377_nG16ba8 , \49526 );
buf \U$39677 ( \50379 , \50378_nG16ba9 );
_DC g18d48_GF_IsGateDCbyConstraint ( \50380_nG18d48 , \50379 , \42503 );
buf \U$39678 ( \50381 , \50380_nG18d48 );
_HMUX g16baa ( \50382_nG16baa , RIe074960_5397 , \49882 , \50099 );
_HMUX g16bab ( \50383_nG16bab , RIe074960_5397 , \50382_nG16baa , \49514 );
_HMUX g16bac ( \50384_nG16bac , RIe074960_5397 , \49885 , \50103 );
_HMUX g16bad ( \50385_nG16bad , \50383_nG16bab , \50384_nG16bac , \49526 );
buf \U$39679 ( \50386 , \50385_nG16bad );
_DC g18d4a_GF_IsGateDCbyConstraint ( \50387_nG18d4a , \50386 , \42503 );
buf \U$39680 ( \50388 , \50387_nG18d4a );
_HMUX g16bae ( \50389_nG16bae , RIe0762b0_5398 , \49891 , \50099 );
_HMUX g16baf ( \50390_nG16baf , RIe0762b0_5398 , \50389_nG16bae , \49514 );
_HMUX g16bb0 ( \50391_nG16bb0 , RIe0762b0_5398 , \49894 , \50103 );
_HMUX g16bb1 ( \50392_nG16bb1 , \50390_nG16baf , \50391_nG16bb0 , \49526 );
buf \U$39681 ( \50393 , \50392_nG16bb1 );
_DC g18d4c_GF_IsGateDCbyConstraint ( \50394_nG18d4c , \50393 , \42503 );
buf \U$39682 ( \50395 , \50394_nG18d4c );
_HMUX g16bb2 ( \50396_nG16bb2 , RIe0779a8_5399 , \49900 , \50099 );
_HMUX g16bb3 ( \50397_nG16bb3 , RIe0779a8_5399 , \50396_nG16bb2 , \49514 );
_HMUX g16bb4 ( \50398_nG16bb4 , RIe0779a8_5399 , \49903 , \50103 );
_HMUX g16bb5 ( \50399_nG16bb5 , \50397_nG16bb3 , \50398_nG16bb4 , \49526 );
buf \U$39683 ( \50400 , \50399_nG16bb5 );
_DC g18d4e_GF_IsGateDCbyConstraint ( \50401_nG18d4e , \50400 , \42503 );
buf \U$39684 ( \50402 , \50401_nG18d4e );
_HMUX g16bb6 ( \50403_nG16bb6 , RIe079118_5400 , \49909 , \50099 );
_HMUX g16bb7 ( \50404_nG16bb7 , RIe079118_5400 , \50403_nG16bb6 , \49514 );
_HMUX g16bb8 ( \50405_nG16bb8 , RIe079118_5400 , \49912 , \50103 );
_HMUX g16bb9 ( \50406_nG16bb9 , \50404_nG16bb7 , \50405_nG16bb8 , \49526 );
buf \U$39685 ( \50407 , \50406_nG16bb9 );
_DC g18d50_GF_IsGateDCbyConstraint ( \50408_nG18d50 , \50407 , \42503 );
buf \U$39686 ( \50409 , \50408_nG18d50 );
_HMUX g16bba ( \50410_nG16bba , RIe07a798_5401 , \49918 , \50099 );
_HMUX g16bbb ( \50411_nG16bbb , RIe07a798_5401 , \50410_nG16bba , \49514 );
_HMUX g16bbc ( \50412_nG16bbc , RIe07a798_5401 , \49921 , \50103 );
_HMUX g16bbd ( \50413_nG16bbd , \50411_nG16bbb , \50412_nG16bbc , \49526 );
buf \U$39687 ( \50414 , \50413_nG16bbd );
_DC g18d52_GF_IsGateDCbyConstraint ( \50415_nG18d52 , \50414 , \42503 );
buf \U$39688 ( \50416 , \50415_nG18d52 );
_HMUX g16bbe ( \50417_nG16bbe , RIe07bcb0_5402 , \49927 , \50099 );
_HMUX g16bbf ( \50418_nG16bbf , RIe07bcb0_5402 , \50417_nG16bbe , \49514 );
_HMUX g16bc0 ( \50419_nG16bc0 , RIe07bcb0_5402 , \49930 , \50103 );
_HMUX g16bc1 ( \50420_nG16bc1 , \50418_nG16bbf , \50419_nG16bc0 , \49526 );
buf \U$39689 ( \50421 , \50420_nG16bc1 );
_DC g18d54_GF_IsGateDCbyConstraint ( \50422_nG18d54 , \50421 , \42503 );
buf \U$39690 ( \50423 , \50422_nG18d54 );
_HMUX g16bc2 ( \50424_nG16bc2 , RIe07d768_5403 , \49936 , \50099 );
_HMUX g16bc3 ( \50425_nG16bc3 , RIe07d768_5403 , \50424_nG16bc2 , \49514 );
_HMUX g16bc4 ( \50426_nG16bc4 , RIe07d768_5403 , \49939 , \50103 );
_HMUX g16bc5 ( \50427_nG16bc5 , \50425_nG16bc3 , \50426_nG16bc4 , \49526 );
buf \U$39691 ( \50428 , \50427_nG16bc5 );
_DC g18d56_GF_IsGateDCbyConstraint ( \50429_nG18d56 , \50428 , \42503 );
buf \U$39692 ( \50430 , \50429_nG18d56 );
_HMUX g16bc6 ( \50431_nG16bc6 , RIe07f220_5404 , \49945 , \50099 );
_HMUX g16bc7 ( \50432_nG16bc7 , RIe07f220_5404 , \50431_nG16bc6 , \49514 );
_HMUX g16bc8 ( \50433_nG16bc8 , RIe07f220_5404 , \49948 , \50103 );
_HMUX g16bc9 ( \50434_nG16bc9 , \50432_nG16bc7 , \50433_nG16bc8 , \49526 );
buf \U$39693 ( \50435 , \50434_nG16bc9 );
_DC g18d58_GF_IsGateDCbyConstraint ( \50436_nG18d58 , \50435 , \42503 );
buf \U$39694 ( \50437 , \50436_nG18d58 );
_HMUX g16bca ( \50438_nG16bca , RIe080cd8_5405 , \49954 , \50099 );
_HMUX g16bcb ( \50439_nG16bcb , RIe080cd8_5405 , \50438_nG16bca , \49514 );
_HMUX g16bcc ( \50440_nG16bcc , RIe080cd8_5405 , \49957 , \50103 );
_HMUX g16bcd ( \50441_nG16bcd , \50439_nG16bcb , \50440_nG16bcc , \49526 );
buf \U$39695 ( \50442 , \50441_nG16bcd );
_DC g18d5a_GF_IsGateDCbyConstraint ( \50443_nG18d5a , \50442 , \42503 );
buf \U$39696 ( \50444 , \50443_nG18d5a );
_HMUX g16bce ( \50445_nG16bce , RIe082088_5406 , \49963 , \50099 );
_HMUX g16bcf ( \50446_nG16bcf , RIe082088_5406 , \50445_nG16bce , \49514 );
_HMUX g16bd0 ( \50447_nG16bd0 , RIe082088_5406 , \49966 , \50103 );
_HMUX g16bd1 ( \50448_nG16bd1 , \50446_nG16bcf , \50447_nG16bd0 , \49526 );
buf \U$39697 ( \50449 , \50448_nG16bd1 );
_DC g18d5e_GF_IsGateDCbyConstraint ( \50450_nG18d5e , \50449 , \42503 );
buf \U$39698 ( \50451 , \50450_nG18d5e );
_HMUX g16bd2 ( \50452_nG16bd2 , RIe083078_5407 , \49972 , \50099 );
_HMUX g16bd3 ( \50453_nG16bd3 , RIe083078_5407 , \50452_nG16bd2 , \49514 );
_HMUX g16bd4 ( \50454_nG16bd4 , RIe083078_5407 , \49975 , \50103 );
_HMUX g16bd5 ( \50455_nG16bd5 , \50453_nG16bd3 , \50454_nG16bd4 , \49526 );
buf \U$39699 ( \50456 , \50455_nG16bd5 );
_DC g18d60_GF_IsGateDCbyConstraint ( \50457_nG18d60 , \50456 , \42503 );
buf \U$39700 ( \50458 , \50457_nG18d60 );
_HMUX g16bd6 ( \50459_nG16bd6 , RIe0843b0_5408 , \49981 , \50099 );
_HMUX g16bd7 ( \50460_nG16bd7 , RIe0843b0_5408 , \50459_nG16bd6 , \49514 );
_HMUX g16bd8 ( \50461_nG16bd8 , RIe0843b0_5408 , \49984 , \50103 );
_HMUX g16bd9 ( \50462_nG16bd9 , \50460_nG16bd7 , \50461_nG16bd8 , \49526 );
buf \U$39701 ( \50463 , \50462_nG16bd9 );
_DC g18d62_GF_IsGateDCbyConstraint ( \50464_nG18d62 , \50463 , \42503 );
buf \U$39702 ( \50465 , \50464_nG18d62 );
_HMUX g16bda ( \50466_nG16bda , RIdfbbbf0_5409 , \49990 , \50099 );
_HMUX g16bdb ( \50467_nG16bdb , RIdfbbbf0_5409 , \50466_nG16bda , \49514 );
_HMUX g16bdc ( \50468_nG16bdc , RIdfbbbf0_5409 , \49993 , \50103 );
_HMUX g16bdd ( \50469_nG16bdd , \50467_nG16bdb , \50468_nG16bdc , \49526 );
buf \U$39703 ( \50470 , \50469_nG16bdd );
_DC g18d64_GF_IsGateDCbyConstraint ( \50471_nG18d64 , \50470 , \42503 );
buf \U$39704 ( \50472 , \50471_nG18d64 );
_HMUX g16bde ( \50473_nG16bde , RIdfbd5b8_5410 , \49999 , \50099 );
_HMUX g16bdf ( \50474_nG16bdf , RIdfbd5b8_5410 , \50473_nG16bde , \49514 );
_HMUX g16be0 ( \50475_nG16be0 , RIdfbd5b8_5410 , \50002 , \50103 );
_HMUX g16be1 ( \50476_nG16be1 , \50474_nG16bdf , \50475_nG16be0 , \49526 );
buf \U$39705 ( \50477 , \50476_nG16be1 );
_DC g18d66_GF_IsGateDCbyConstraint ( \50478_nG18d66 , \50477 , \42503 );
buf \U$39706 ( \50479 , \50478_nG18d66 );
_HMUX g16be2 ( \50480_nG16be2 , RIdfbf3b8_5411 , \50008 , \50099 );
_HMUX g16be3 ( \50481_nG16be3 , RIdfbf3b8_5411 , \50480_nG16be2 , \49514 );
_HMUX g16be4 ( \50482_nG16be4 , RIdfbf3b8_5411 , \50011 , \50103 );
_HMUX g16be5 ( \50483_nG16be5 , \50481_nG16be3 , \50482_nG16be4 , \49526 );
buf \U$39707 ( \50484 , \50483_nG16be5 );
_DC g18d68_GF_IsGateDCbyConstraint ( \50485_nG18d68 , \50484 , \42503 );
buf \U$39708 ( \50486 , \50485_nG18d68 );
_HMUX g16be6 ( \50487_nG16be6 , RIdfc15f0_5412 , \50017 , \50099 );
_HMUX g16be7 ( \50488_nG16be7 , RIdfc15f0_5412 , \50487_nG16be6 , \49514 );
_HMUX g16be8 ( \50489_nG16be8 , RIdfc15f0_5412 , \50020 , \50103 );
_HMUX g16be9 ( \50490_nG16be9 , \50488_nG16be7 , \50489_nG16be8 , \49526 );
buf \U$39709 ( \50491 , \50490_nG16be9 );
_DC g18d6a_GF_IsGateDCbyConstraint ( \50492_nG18d6a , \50491 , \42503 );
buf \U$39710 ( \50493 , \50492_nG18d6a );
_HMUX g16bea ( \50494_nG16bea , RIdfc30a8_5413 , \50026 , \50099 );
_HMUX g16beb ( \50495_nG16beb , RIdfc30a8_5413 , \50494_nG16bea , \49514 );
_HMUX g16bec ( \50496_nG16bec , RIdfc30a8_5413 , \50029 , \50103 );
_HMUX g16bed ( \50497_nG16bed , \50495_nG16beb , \50496_nG16bec , \49526 );
buf \U$39711 ( \50498 , \50497_nG16bed );
_DC g18d6c_GF_IsGateDCbyConstraint ( \50499_nG18d6c , \50498 , \42503 );
buf \U$39712 ( \50500 , \50499_nG18d6c );
_HMUX g16bee ( \50501_nG16bee , RIdfc4f20_5414 , \50035 , \50099 );
_HMUX g16bef ( \50502_nG16bef , RIdfc4f20_5414 , \50501_nG16bee , \49514 );
_HMUX g16bf0 ( \50503_nG16bf0 , RIdfc4f20_5414 , \50038 , \50103 );
_HMUX g16bf1 ( \50504_nG16bf1 , \50502_nG16bef , \50503_nG16bf0 , \49526 );
buf \U$39713 ( \50505 , \50504_nG16bf1 );
_DC g18d6e_GF_IsGateDCbyConstraint ( \50506_nG18d6e , \50505 , \42503 );
buf \U$39714 ( \50507 , \50506_nG18d6e );
_HMUX g16bf2 ( \50508_nG16bf2 , RIdfc6f00_5415 , \50044 , \50099 );
_HMUX g16bf3 ( \50509_nG16bf3 , RIdfc6f00_5415 , \50508_nG16bf2 , \49514 );
_HMUX g16bf4 ( \50510_nG16bf4 , RIdfc6f00_5415 , \50047 , \50103 );
_HMUX g16bf5 ( \50511_nG16bf5 , \50509_nG16bf3 , \50510_nG16bf4 , \49526 );
buf \U$39715 ( \50512 , \50511_nG16bf5 );
_DC g18d70_GF_IsGateDCbyConstraint ( \50513_nG18d70 , \50512 , \42503 );
buf \U$39716 ( \50514 , \50513_nG18d70 );
_HMUX g16bf6 ( \50515_nG16bf6 , RIdfc85f8_5416 , \50053 , \50099 );
_HMUX g16bf7 ( \50516_nG16bf7 , RIdfc85f8_5416 , \50515_nG16bf6 , \49514 );
_HMUX g16bf8 ( \50517_nG16bf8 , RIdfc85f8_5416 , \50056 , \50103 );
_HMUX g16bf9 ( \50518_nG16bf9 , \50516_nG16bf7 , \50517_nG16bf8 , \49526 );
buf \U$39717 ( \50519 , \50518_nG16bf9 );
_DC g18d74_GF_IsGateDCbyConstraint ( \50520_nG18d74 , \50519 , \42503 );
buf \U$39718 ( \50521 , \50520_nG18d74 );
_HMUX g16bfa ( \50522_nG16bfa , RIdfca3f8_5417 , \50062 , \50099 );
_HMUX g16bfb ( \50523_nG16bfb , RIdfca3f8_5417 , \50522_nG16bfa , \49514 );
_HMUX g16bfc ( \50524_nG16bfc , RIdfca3f8_5417 , \50065 , \50103 );
_HMUX g16bfd ( \50525_nG16bfd , \50523_nG16bfb , \50524_nG16bfc , \49526 );
buf \U$39719 ( \50526 , \50525_nG16bfd );
_DC g18d76_GF_IsGateDCbyConstraint ( \50527_nG18d76 , \50526 , \42503 );
buf \U$39720 ( \50528 , \50527_nG18d76 );
_HMUX g16bfe ( \50529_nG16bfe , RIdfcc720_5418 , \50071 , \50099 );
_HMUX g16bff ( \50530_nG16bff , RIdfcc720_5418 , \50529_nG16bfe , \49514 );
_HMUX g16c00 ( \50531_nG16c00 , RIdfcc720_5418 , \50074 , \50103 );
_HMUX g16c01 ( \50532_nG16c01 , \50530_nG16bff , \50531_nG16c00 , \49526 );
buf \U$39721 ( \50533 , \50532_nG16c01 );
_DC g18d78_GF_IsGateDCbyConstraint ( \50534_nG18d78 , \50533 , \42503 );
buf \U$39722 ( \50535 , \50534_nG18d78 );
_HMUX g16c02 ( \50536_nG16c02 , RIdfce8e0_5419 , \50080 , \50099 );
_HMUX g16c03 ( \50537_nG16c03 , RIdfce8e0_5419 , \50536_nG16c02 , \49514 );
_HMUX g16c04 ( \50538_nG16c04 , RIdfce8e0_5419 , \50083 , \50103 );
_HMUX g16c05 ( \50539_nG16c05 , \50537_nG16c03 , \50538_nG16c04 , \49526 );
buf \U$39723 ( \50540 , \50539_nG16c05 );
_DC g18d7a_GF_IsGateDCbyConstraint ( \50541_nG18d7a , \50540 , \42503 );
buf \U$39724 ( \50542 , \50541_nG18d7a );
_HMUX g16c06 ( \50543_nG16c06 , RIe106478_5420 , \50089 , \50099 );
_HMUX g16c07 ( \50544_nG16c07 , RIe106478_5420 , \50543_nG16c06 , \49514 );
_HMUX g16c08 ( \50545_nG16c08 , RIe106478_5420 , \50092 , \50103 );
_HMUX g16c09 ( \50546_nG16c09 , \50544_nG16c07 , \50545_nG16c08 , \49526 );
buf \U$39725 ( \50547 , \50546_nG16c09 );
_DC g18d7c_GF_IsGateDCbyConstraint ( \50548_nG18d7c , \50547 , \42503 );
buf \U$39726 ( \50549 , \50548_nG18d7c );
nor \U$39727 ( \50550 , \49505 , \50098 );
_HMUX g16a07 ( \50551_nG16a07 , RIe104948_5421 , \49504 , \50550 );
_HMUX g16a08 ( \50552_nG16a08 , RIe104948_5421 , \50551_nG16a07 , \49514 );
nor \U$39728 ( \50553 , \49517 , \50102 );
_HMUX g16a0b ( \50554_nG16a0b , RIe104948_5421 , \49516 , \50553 );
_HMUX g16a0c ( \50555_nG16a0c , \50552_nG16a08 , \50554_nG16a0b , \49526 );
buf \U$39729 ( \50556 , \50555_nG16a0c );
_DC g18c84_GF_IsGateDCbyConstraint ( \50557_nG18c84 , \50556 , \42503 );
buf \U$39730 ( \50558 , \50557_nG18c84 );
_HMUX g16a0d ( \50559_nG16a0d , RIe102b48_5422 , \49531 , \50550 );
_HMUX g16a0e ( \50560_nG16a0e , RIe102b48_5422 , \50559_nG16a0d , \49514 );
_HMUX g16a0f ( \50561_nG16a0f , RIe102b48_5422 , \49534 , \50553 );
_HMUX g16a10 ( \50562_nG16a10 , \50560_nG16a0e , \50561_nG16a0f , \49526 );
buf \U$39731 ( \50563 , \50562_nG16a10 );
_DC g18c9a_GF_IsGateDCbyConstraint ( \50564_nG18c9a , \50563 , \42503 );
buf \U$39732 ( \50565 , \50564_nG18c9a );
_HMUX g16a11 ( \50566_nG16a11 , RIe100f28_5423 , \49540 , \50550 );
_HMUX g16a12 ( \50567_nG16a12 , RIe100f28_5423 , \50566_nG16a11 , \49514 );
_HMUX g16a13 ( \50568_nG16a13 , RIe100f28_5423 , \49543 , \50553 );
_HMUX g16a14 ( \50569_nG16a14 , \50567_nG16a12 , \50568_nG16a13 , \49526 );
buf \U$39733 ( \50570 , \50569_nG16a14 );
_DC g18cb0_GF_IsGateDCbyConstraint ( \50571_nG18cb0 , \50570 , \42503 );
buf \U$39734 ( \50572 , \50571_nG18cb0 );
_HMUX g16a15 ( \50573_nG16a15 , RIe0fea20_5424 , \49549 , \50550 );
_HMUX g16a16 ( \50574_nG16a16 , RIe0fea20_5424 , \50573_nG16a15 , \49514 );
_HMUX g16a17 ( \50575_nG16a17 , RIe0fea20_5424 , \49552 , \50553 );
_HMUX g16a18 ( \50576_nG16a18 , \50574_nG16a16 , \50575_nG16a17 , \49526 );
buf \U$39735 ( \50577 , \50576_nG16a18 );
_DC g18cc6_GF_IsGateDCbyConstraint ( \50578_nG18cc6 , \50577 , \42503 );
buf \U$39736 ( \50579 , \50578_nG18cc6 );
_HMUX g16a19 ( \50580_nG16a19 , RIe0fcd10_5425 , \49558 , \50550 );
_HMUX g16a1a ( \50581_nG16a1a , RIe0fcd10_5425 , \50580_nG16a19 , \49514 );
_HMUX g16a1b ( \50582_nG16a1b , RIe0fcd10_5425 , \49561 , \50553 );
_HMUX g16a1c ( \50583_nG16a1c , \50581_nG16a1a , \50582_nG16a1b , \49526 );
buf \U$39737 ( \50584 , \50583_nG16a1c );
_DC g18cdc_GF_IsGateDCbyConstraint ( \50585_nG18cdc , \50584 , \42503 );
buf \U$39738 ( \50586 , \50585_nG18cdc );
_HMUX g16a1d ( \50587_nG16a1d , RIe0fa3d0_5426 , \49567 , \50550 );
_HMUX g16a1e ( \50588_nG16a1e , RIe0fa3d0_5426 , \50587_nG16a1d , \49514 );
_HMUX g16a1f ( \50589_nG16a1f , RIe0fa3d0_5426 , \49570 , \50553 );
_HMUX g16a20 ( \50590_nG16a20 , \50588_nG16a1e , \50589_nG16a1f , \49526 );
buf \U$39739 ( \50591 , \50590_nG16a20 );
_DC g18cf2_GF_IsGateDCbyConstraint ( \50592_nG18cf2 , \50591 , \42503 );
buf \U$39740 ( \50593 , \50592_nG18cf2 );
_HMUX g16a21 ( \50594_nG16a21 , RIe0f7838_5427 , \49576 , \50550 );
_HMUX g16a22 ( \50595_nG16a22 , RIe0f7838_5427 , \50594_nG16a21 , \49514 );
_HMUX g16a23 ( \50596_nG16a23 , RIe0f7838_5427 , \49579 , \50553 );
_HMUX g16a24 ( \50597_nG16a24 , \50595_nG16a22 , \50596_nG16a23 , \49526 );
buf \U$39741 ( \50598 , \50597_nG16a24 );
_DC g18cfe_GF_IsGateDCbyConstraint ( \50599_nG18cfe , \50598 , \42503 );
buf \U$39742 ( \50600 , \50599_nG18cfe );
_HMUX g16a25 ( \50601_nG16a25 , RIe0f5a38_5428 , \49585 , \50550 );
_HMUX g16a26 ( \50602_nG16a26 , RIe0f5a38_5428 , \50601_nG16a25 , \49514 );
_HMUX g16a27 ( \50603_nG16a27 , RIe0f5a38_5428 , \49588 , \50553 );
_HMUX g16a28 ( \50604_nG16a28 , \50602_nG16a26 , \50603_nG16a27 , \49526 );
buf \U$39743 ( \50605 , \50604_nG16a28 );
_DC g18d00_GF_IsGateDCbyConstraint ( \50606_nG18d00 , \50605 , \42503 );
buf \U$39744 ( \50607 , \50606_nG18d00 );
_HMUX g16a29 ( \50608_nG16a29 , RIe0f3968_5429 , \49594 , \50550 );
_HMUX g16a2a ( \50609_nG16a2a , RIe0f3968_5429 , \50608_nG16a29 , \49514 );
_HMUX g16a2b ( \50610_nG16a2b , RIe0f3968_5429 , \49597 , \50553 );
_HMUX g16a2c ( \50611_nG16a2c , \50609_nG16a2a , \50610_nG16a2b , \49526 );
buf \U$39745 ( \50612 , \50611_nG16a2c );
_DC g18d02_GF_IsGateDCbyConstraint ( \50613_nG18d02 , \50612 , \42503 );
buf \U$39746 ( \50614 , \50613_nG18d02 );
_HMUX g16a2d ( \50615_nG16a2d , RIe0f1b68_5430 , \49603 , \50550 );
_HMUX g16a2e ( \50616_nG16a2e , RIe0f1b68_5430 , \50615_nG16a2d , \49514 );
_HMUX g16a2f ( \50617_nG16a2f , RIe0f1b68_5430 , \49606 , \50553 );
_HMUX g16a30 ( \50618_nG16a30 , \50616_nG16a2e , \50617_nG16a2f , \49526 );
buf \U$39747 ( \50619 , \50618_nG16a30 );
_DC g18c86_GF_IsGateDCbyConstraint ( \50620_nG18c86 , \50619 , \42503 );
buf \U$39748 ( \50621 , \50620_nG18c86 );
_HMUX g16a31 ( \50622_nG16a31 , RIe0f0290_5431 , \49612 , \50550 );
_HMUX g16a32 ( \50623_nG16a32 , RIe0f0290_5431 , \50622_nG16a31 , \49514 );
_HMUX g16a33 ( \50624_nG16a33 , RIe0f0290_5431 , \49615 , \50553 );
_HMUX g16a34 ( \50625_nG16a34 , \50623_nG16a32 , \50624_nG16a33 , \49526 );
buf \U$39749 ( \50626 , \50625_nG16a34 );
_DC g18c88_GF_IsGateDCbyConstraint ( \50627_nG18c88 , \50626 , \42503 );
buf \U$39750 ( \50628 , \50627_nG18c88 );
_HMUX g16a35 ( \50629_nG16a35 , RIe0ee508_5432 , \49621 , \50550 );
_HMUX g16a36 ( \50630_nG16a36 , RIe0ee508_5432 , \50629_nG16a35 , \49514 );
_HMUX g16a37 ( \50631_nG16a37 , RIe0ee508_5432 , \49624 , \50553 );
_HMUX g16a38 ( \50632_nG16a38 , \50630_nG16a36 , \50631_nG16a37 , \49526 );
buf \U$39751 ( \50633 , \50632_nG16a38 );
_DC g18c8a_GF_IsGateDCbyConstraint ( \50634_nG18c8a , \50633 , \42503 );
buf \U$39752 ( \50635 , \50634_nG18c8a );
_HMUX g16a39 ( \50636_nG16a39 , RIe0ec690_5433 , \49630 , \50550 );
_HMUX g16a3a ( \50637_nG16a3a , RIe0ec690_5433 , \50636_nG16a39 , \49514 );
_HMUX g16a3b ( \50638_nG16a3b , RIe0ec690_5433 , \49633 , \50553 );
_HMUX g16a3c ( \50639_nG16a3c , \50637_nG16a3a , \50638_nG16a3b , \49526 );
buf \U$39753 ( \50640 , \50639_nG16a3c );
_DC g18c8c_GF_IsGateDCbyConstraint ( \50641_nG18c8c , \50640 , \42503 );
buf \U$39754 ( \50642 , \50641_nG18c8c );
_HMUX g16a3d ( \50643_nG16a3d , RIe0eaea8_5434 , \49639 , \50550 );
_HMUX g16a3e ( \50644_nG16a3e , RIe0eaea8_5434 , \50643_nG16a3d , \49514 );
_HMUX g16a3f ( \50645_nG16a3f , RIe0eaea8_5434 , \49642 , \50553 );
_HMUX g16a40 ( \50646_nG16a40 , \50644_nG16a3e , \50645_nG16a3f , \49526 );
buf \U$39755 ( \50647 , \50646_nG16a40 );
_DC g18c8e_GF_IsGateDCbyConstraint ( \50648_nG18c8e , \50647 , \42503 );
buf \U$39756 ( \50649 , \50648_nG18c8e );
_HMUX g16a41 ( \50650_nG16a41 , RIe0e8658_5435 , \49648 , \50550 );
_HMUX g16a42 ( \50651_nG16a42 , RIe0e8658_5435 , \50650_nG16a41 , \49514 );
_HMUX g16a43 ( \50652_nG16a43 , RIe0e8658_5435 , \49651 , \50553 );
_HMUX g16a44 ( \50653_nG16a44 , \50651_nG16a42 , \50652_nG16a43 , \49526 );
buf \U$39757 ( \50654 , \50653_nG16a44 );
_DC g18c90_GF_IsGateDCbyConstraint ( \50655_nG18c90 , \50654 , \42503 );
buf \U$39758 ( \50656 , \50655_nG18c90 );
_HMUX g16a45 ( \50657_nG16a45 , RIe0e54a8_5436 , \49657 , \50550 );
_HMUX g16a46 ( \50658_nG16a46 , RIe0e54a8_5436 , \50657_nG16a45 , \49514 );
_HMUX g16a47 ( \50659_nG16a47 , RIe0e54a8_5436 , \49660 , \50553 );
_HMUX g16a48 ( \50660_nG16a48 , \50658_nG16a46 , \50659_nG16a47 , \49526 );
buf \U$39759 ( \50661 , \50660_nG16a48 );
_DC g18c92_GF_IsGateDCbyConstraint ( \50662_nG18c92 , \50661 , \42503 );
buf \U$39760 ( \50663 , \50662_nG18c92 );
_HMUX g16a49 ( \50664_nG16a49 , RIe0e2988_5437 , \49666 , \50550 );
_HMUX g16a4a ( \50665_nG16a4a , RIe0e2988_5437 , \50664_nG16a49 , \49514 );
_HMUX g16a4b ( \50666_nG16a4b , RIe0e2988_5437 , \49669 , \50553 );
_HMUX g16a4c ( \50667_nG16a4c , \50665_nG16a4a , \50666_nG16a4b , \49526 );
buf \U$39761 ( \50668 , \50667_nG16a4c );
_DC g18c94_GF_IsGateDCbyConstraint ( \50669_nG18c94 , \50668 , \42503 );
buf \U$39762 ( \50670 , \50669_nG18c94 );
_HMUX g16a4d ( \50671_nG16a4d , RIe0e0228_5438 , \49675 , \50550 );
_HMUX g16a4e ( \50672_nG16a4e , RIe0e0228_5438 , \50671_nG16a4d , \49514 );
_HMUX g16a4f ( \50673_nG16a4f , RIe0e0228_5438 , \49678 , \50553 );
_HMUX g16a50 ( \50674_nG16a50 , \50672_nG16a4e , \50673_nG16a4f , \49526 );
buf \U$39763 ( \50675 , \50674_nG16a50 );
_DC g18c96_GF_IsGateDCbyConstraint ( \50676_nG18c96 , \50675 , \42503 );
buf \U$39764 ( \50677 , \50676_nG18c96 );
_HMUX g16a51 ( \50678_nG16a51 , RIe0dd7f8_5439 , \49684 , \50550 );
_HMUX g16a52 ( \50679_nG16a52 , RIe0dd7f8_5439 , \50678_nG16a51 , \49514 );
_HMUX g16a53 ( \50680_nG16a53 , RIe0dd7f8_5439 , \49687 , \50553 );
_HMUX g16a54 ( \50681_nG16a54 , \50679_nG16a52 , \50680_nG16a53 , \49526 );
buf \U$39765 ( \50682 , \50681_nG16a54 );
_DC g18c98_GF_IsGateDCbyConstraint ( \50683_nG18c98 , \50682 , \42503 );
buf \U$39766 ( \50684 , \50683_nG18c98 );
_HMUX g16a55 ( \50685_nG16a55 , RIe0da828_5440 , \49693 , \50550 );
_HMUX g16a56 ( \50686_nG16a56 , RIe0da828_5440 , \50685_nG16a55 , \49514 );
_HMUX g16a57 ( \50687_nG16a57 , RIe0da828_5440 , \49696 , \50553 );
_HMUX g16a58 ( \50688_nG16a58 , \50686_nG16a56 , \50687_nG16a57 , \49526 );
buf \U$39767 ( \50689 , \50688_nG16a58 );
_DC g18c9c_GF_IsGateDCbyConstraint ( \50690_nG18c9c , \50689 , \42503 );
buf \U$39768 ( \50691 , \50690_nG18c9c );
_HMUX g16a59 ( \50692_nG16a59 , RIe0d7f60_5441 , \49702 , \50550 );
_HMUX g16a5a ( \50693_nG16a5a , RIe0d7f60_5441 , \50692_nG16a59 , \49514 );
_HMUX g16a5b ( \50694_nG16a5b , RIe0d7f60_5441 , \49705 , \50553 );
_HMUX g16a5c ( \50695_nG16a5c , \50693_nG16a5a , \50694_nG16a5b , \49526 );
buf \U$39769 ( \50696 , \50695_nG16a5c );
_DC g18c9e_GF_IsGateDCbyConstraint ( \50697_nG18c9e , \50696 , \42503 );
buf \U$39770 ( \50698 , \50697_nG18c9e );
_HMUX g16a5d ( \50699_nG16a5d , RIe0d4f18_5442 , \49711 , \50550 );
_HMUX g16a5e ( \50700_nG16a5e , RIe0d4f18_5442 , \50699_nG16a5d , \49514 );
_HMUX g16a5f ( \50701_nG16a5f , RIe0d4f18_5442 , \49714 , \50553 );
_HMUX g16a60 ( \50702_nG16a60 , \50700_nG16a5e , \50701_nG16a5f , \49526 );
buf \U$39771 ( \50703 , \50702_nG16a60 );
_DC g18ca0_GF_IsGateDCbyConstraint ( \50704_nG18ca0 , \50703 , \42503 );
buf \U$39772 ( \50705 , \50704_nG18ca0 );
_HMUX g16a61 ( \50706_nG16a61 , RIe0d3280_5443 , \49720 , \50550 );
_HMUX g16a62 ( \50707_nG16a62 , RIe0d3280_5443 , \50706_nG16a61 , \49514 );
_HMUX g16a63 ( \50708_nG16a63 , RIe0d3280_5443 , \49723 , \50553 );
_HMUX g16a64 ( \50709_nG16a64 , \50707_nG16a62 , \50708_nG16a63 , \49526 );
buf \U$39773 ( \50710 , \50709_nG16a64 );
_DC g18ca2_GF_IsGateDCbyConstraint ( \50711_nG18ca2 , \50710 , \42503 );
buf \U$39774 ( \50712 , \50711_nG18ca2 );
_HMUX g16a65 ( \50713_nG16a65 , RIe0d02b0_5444 , \49729 , \50550 );
_HMUX g16a66 ( \50714_nG16a66 , RIe0d02b0_5444 , \50713_nG16a65 , \49514 );
_HMUX g16a67 ( \50715_nG16a67 , RIe0d02b0_5444 , \49732 , \50553 );
_HMUX g16a68 ( \50716_nG16a68 , \50714_nG16a66 , \50715_nG16a67 , \49526 );
buf \U$39775 ( \50717 , \50716_nG16a68 );
_DC g18ca4_GF_IsGateDCbyConstraint ( \50718_nG18ca4 , \50717 , \42503 );
buf \U$39776 ( \50719 , \50718_nG18ca4 );
_HMUX g16a69 ( \50720_nG16a69 , RIe0cdad8_5445 , \49738 , \50550 );
_HMUX g16a6a ( \50721_nG16a6a , RIe0cdad8_5445 , \50720_nG16a69 , \49514 );
_HMUX g16a6b ( \50722_nG16a6b , RIe0cdad8_5445 , \49741 , \50553 );
_HMUX g16a6c ( \50723_nG16a6c , \50721_nG16a6a , \50722_nG16a6b , \49526 );
buf \U$39777 ( \50724 , \50723_nG16a6c );
_DC g18ca6_GF_IsGateDCbyConstraint ( \50725_nG18ca6 , \50724 , \42503 );
buf \U$39778 ( \50726 , \50725_nG18ca6 );
_HMUX g16a6d ( \50727_nG16a6d , RIe0cae50_5446 , \49747 , \50550 );
_HMUX g16a6e ( \50728_nG16a6e , RIe0cae50_5446 , \50727_nG16a6d , \49514 );
_HMUX g16a6f ( \50729_nG16a6f , RIe0cae50_5446 , \49750 , \50553 );
_HMUX g16a70 ( \50730_nG16a70 , \50728_nG16a6e , \50729_nG16a6f , \49526 );
buf \U$39779 ( \50731 , \50730_nG16a70 );
_DC g18ca8_GF_IsGateDCbyConstraint ( \50732_nG18ca8 , \50731 , \42503 );
buf \U$39780 ( \50733 , \50732_nG18ca8 );
_HMUX g16a71 ( \50734_nG16a71 , RIe0c8150_5447 , \49756 , \50550 );
_HMUX g16a72 ( \50735_nG16a72 , RIe0c8150_5447 , \50734_nG16a71 , \49514 );
_HMUX g16a73 ( \50736_nG16a73 , RIe0c8150_5447 , \49759 , \50553 );
_HMUX g16a74 ( \50737_nG16a74 , \50735_nG16a72 , \50736_nG16a73 , \49526 );
buf \U$39781 ( \50738 , \50737_nG16a74 );
_DC g18caa_GF_IsGateDCbyConstraint ( \50739_nG18caa , \50738 , \42503 );
buf \U$39782 ( \50740 , \50739_nG18caa );
_HMUX g16a75 ( \50741_nG16a75 , RIe0c5d38_5448 , \49765 , \50550 );
_HMUX g16a76 ( \50742_nG16a76 , RIe0c5d38_5448 , \50741_nG16a75 , \49514 );
_HMUX g16a77 ( \50743_nG16a77 , RIe0c5d38_5448 , \49768 , \50553 );
_HMUX g16a78 ( \50744_nG16a78 , \50742_nG16a76 , \50743_nG16a77 , \49526 );
buf \U$39783 ( \50745 , \50744_nG16a78 );
_DC g18cac_GF_IsGateDCbyConstraint ( \50746_nG18cac , \50745 , \42503 );
buf \U$39784 ( \50747 , \50746_nG18cac );
_HMUX g16a79 ( \50748_nG16a79 , RIe0c3290_5449 , \49774 , \50550 );
_HMUX g16a7a ( \50749_nG16a7a , RIe0c3290_5449 , \50748_nG16a79 , \49514 );
_HMUX g16a7b ( \50750_nG16a7b , RIe0c3290_5449 , \49777 , \50553 );
_HMUX g16a7c ( \50751_nG16a7c , \50749_nG16a7a , \50750_nG16a7b , \49526 );
buf \U$39785 ( \50752 , \50751_nG16a7c );
_DC g18cae_GF_IsGateDCbyConstraint ( \50753_nG18cae , \50752 , \42503 );
buf \U$39786 ( \50754 , \50753_nG18cae );
_HMUX g16a7d ( \50755_nG16a7d , RIe0c0d88_5450 , \49783 , \50550 );
_HMUX g16a7e ( \50756_nG16a7e , RIe0c0d88_5450 , \50755_nG16a7d , \49514 );
_HMUX g16a7f ( \50757_nG16a7f , RIe0c0d88_5450 , \49786 , \50553 );
_HMUX g16a80 ( \50758_nG16a80 , \50756_nG16a7e , \50757_nG16a7f , \49526 );
buf \U$39787 ( \50759 , \50758_nG16a80 );
_DC g18cb2_GF_IsGateDCbyConstraint ( \50760_nG18cb2 , \50759 , \42503 );
buf \U$39788 ( \50761 , \50760_nG18cb2 );
_HMUX g16a81 ( \50762_nG16a81 , RIe0be628_5451 , \49792 , \50550 );
_HMUX g16a82 ( \50763_nG16a82 , RIe0be628_5451 , \50762_nG16a81 , \49514 );
_HMUX g16a83 ( \50764_nG16a83 , RIe0be628_5451 , \49795 , \50553 );
_HMUX g16a84 ( \50765_nG16a84 , \50763_nG16a82 , \50764_nG16a83 , \49526 );
buf \U$39789 ( \50766 , \50765_nG16a84 );
_DC g18cb4_GF_IsGateDCbyConstraint ( \50767_nG18cb4 , \50766 , \42503 );
buf \U$39790 ( \50768 , \50767_nG18cb4 );
_HMUX g16a85 ( \50769_nG16a85 , RIe0bbdd8_5452 , \49801 , \50550 );
_HMUX g16a86 ( \50770_nG16a86 , RIe0bbdd8_5452 , \50769_nG16a85 , \49514 );
_HMUX g16a87 ( \50771_nG16a87 , RIe0bbdd8_5452 , \49804 , \50553 );
_HMUX g16a88 ( \50772_nG16a88 , \50770_nG16a86 , \50771_nG16a87 , \49526 );
buf \U$39791 ( \50773 , \50772_nG16a88 );
_DC g18cb6_GF_IsGateDCbyConstraint ( \50774_nG18cb6 , \50773 , \42503 );
buf \U$39792 ( \50775 , \50774_nG18cb6 );
_HMUX g16a89 ( \50776_nG16a89 , RIe0b91c8_5453 , \49810 , \50550 );
_HMUX g16a8a ( \50777_nG16a8a , RIe0b91c8_5453 , \50776_nG16a89 , \49514 );
_HMUX g16a8b ( \50778_nG16a8b , RIe0b91c8_5453 , \49813 , \50553 );
_HMUX g16a8c ( \50779_nG16a8c , \50777_nG16a8a , \50778_nG16a8b , \49526 );
buf \U$39793 ( \50780 , \50779_nG16a8c );
_DC g18cb8_GF_IsGateDCbyConstraint ( \50781_nG18cb8 , \50780 , \42503 );
buf \U$39794 ( \50782 , \50781_nG18cb8 );
_HMUX g16a8d ( \50783_nG16a8d , RIe0b5f28_5454 , \49819 , \50550 );
_HMUX g16a8e ( \50784_nG16a8e , RIe0b5f28_5454 , \50783_nG16a8d , \49514 );
_HMUX g16a8f ( \50785_nG16a8f , RIe0b5f28_5454 , \49822 , \50553 );
_HMUX g16a90 ( \50786_nG16a90 , \50784_nG16a8e , \50785_nG16a8f , \49526 );
buf \U$39795 ( \50787 , \50786_nG16a90 );
_DC g18cba_GF_IsGateDCbyConstraint ( \50788_nG18cba , \50787 , \42503 );
buf \U$39796 ( \50789 , \50788_nG18cba );
_HMUX g16a91 ( \50790_nG16a91 , RIe0b3318_5455 , \49828 , \50550 );
_HMUX g16a92 ( \50791_nG16a92 , RIe0b3318_5455 , \50790_nG16a91 , \49514 );
_HMUX g16a93 ( \50792_nG16a93 , RIe0b3318_5455 , \49831 , \50553 );
_HMUX g16a94 ( \50793_nG16a94 , \50791_nG16a92 , \50792_nG16a93 , \49526 );
buf \U$39797 ( \50794 , \50793_nG16a94 );
_DC g18cbc_GF_IsGateDCbyConstraint ( \50795_nG18cbc , \50794 , \42503 );
buf \U$39798 ( \50796 , \50795_nG18cbc );
_HMUX g16a95 ( \50797_nG16a95 , RIe0b02d0_5456 , \49837 , \50550 );
_HMUX g16a96 ( \50798_nG16a96 , RIe0b02d0_5456 , \50797_nG16a95 , \49514 );
_HMUX g16a97 ( \50799_nG16a97 , RIe0b02d0_5456 , \49840 , \50553 );
_HMUX g16a98 ( \50800_nG16a98 , \50798_nG16a96 , \50799_nG16a97 , \49526 );
buf \U$39799 ( \50801 , \50800_nG16a98 );
_DC g18cbe_GF_IsGateDCbyConstraint ( \50802_nG18cbe , \50801 , \42503 );
buf \U$39800 ( \50803 , \50802_nG18cbe );
_HMUX g16a99 ( \50804_nG16a99 , RIe0adeb8_5457 , \49846 , \50550 );
_HMUX g16a9a ( \50805_nG16a9a , RIe0adeb8_5457 , \50804_nG16a99 , \49514 );
_HMUX g16a9b ( \50806_nG16a9b , RIe0adeb8_5457 , \49849 , \50553 );
_HMUX g16a9c ( \50807_nG16a9c , \50805_nG16a9a , \50806_nG16a9b , \49526 );
buf \U$39801 ( \50808 , \50807_nG16a9c );
_DC g18cc0_GF_IsGateDCbyConstraint ( \50809_nG18cc0 , \50808 , \42503 );
buf \U$39802 ( \50810 , \50809_nG18cc0 );
_HMUX g16a9d ( \50811_nG16a9d , RIe0ac0b8_5458 , \49855 , \50550 );
_HMUX g16a9e ( \50812_nG16a9e , RIe0ac0b8_5458 , \50811_nG16a9d , \49514 );
_HMUX g16a9f ( \50813_nG16a9f , RIe0ac0b8_5458 , \49858 , \50553 );
_HMUX g16aa0 ( \50814_nG16aa0 , \50812_nG16a9e , \50813_nG16a9f , \49526 );
buf \U$39803 ( \50815 , \50814_nG16aa0 );
_DC g18cc2_GF_IsGateDCbyConstraint ( \50816_nG18cc2 , \50815 , \42503 );
buf \U$39804 ( \50817 , \50816_nG18cc2 );
_HMUX g16aa1 ( \50818_nG16aa1 , RIe0aa330_5459 , \49864 , \50550 );
_HMUX g16aa2 ( \50819_nG16aa2 , RIe0aa330_5459 , \50818_nG16aa1 , \49514 );
_HMUX g16aa3 ( \50820_nG16aa3 , RIe0aa330_5459 , \49867 , \50553 );
_HMUX g16aa4 ( \50821_nG16aa4 , \50819_nG16aa2 , \50820_nG16aa3 , \49526 );
buf \U$39805 ( \50822 , \50821_nG16aa4 );
_DC g18cc4_GF_IsGateDCbyConstraint ( \50823_nG18cc4 , \50822 , \42503 );
buf \U$39806 ( \50824 , \50823_nG18cc4 );
_HMUX g16aa5 ( \50825_nG16aa5 , RIe0a83c8_5460 , \49873 , \50550 );
_HMUX g16aa6 ( \50826_nG16aa6 , RIe0a83c8_5460 , \50825_nG16aa5 , \49514 );
_HMUX g16aa7 ( \50827_nG16aa7 , RIe0a83c8_5460 , \49876 , \50553 );
_HMUX g16aa8 ( \50828_nG16aa8 , \50826_nG16aa6 , \50827_nG16aa7 , \49526 );
buf \U$39807 ( \50829 , \50828_nG16aa8 );
_DC g18cc8_GF_IsGateDCbyConstraint ( \50830_nG18cc8 , \50829 , \42503 );
buf \U$39808 ( \50831 , \50830_nG18cc8 );
_HMUX g16aa9 ( \50832_nG16aa9 , RIe0a6a00_5461 , \49882 , \50550 );
_HMUX g16aaa ( \50833_nG16aaa , RIe0a6a00_5461 , \50832_nG16aa9 , \49514 );
_HMUX g16aab ( \50834_nG16aab , RIe0a6a00_5461 , \49885 , \50553 );
_HMUX g16aac ( \50835_nG16aac , \50833_nG16aaa , \50834_nG16aab , \49526 );
buf \U$39809 ( \50836 , \50835_nG16aac );
_DC g18cca_GF_IsGateDCbyConstraint ( \50837_nG18cca , \50836 , \42503 );
buf \U$39810 ( \50838 , \50837_nG18cca );
_HMUX g16aad ( \50839_nG16aad , RIe0a40c0_5462 , \49891 , \50550 );
_HMUX g16aae ( \50840_nG16aae , RIe0a40c0_5462 , \50839_nG16aad , \49514 );
_HMUX g16aaf ( \50841_nG16aaf , RIe0a40c0_5462 , \49894 , \50553 );
_HMUX g16ab0 ( \50842_nG16ab0 , \50840_nG16aae , \50841_nG16aaf , \49526 );
buf \U$39811 ( \50843 , \50842_nG16ab0 );
_DC g18ccc_GF_IsGateDCbyConstraint ( \50844_nG18ccc , \50843 , \42503 );
buf \U$39812 ( \50845 , \50844_nG18ccc );
_HMUX g16ab1 ( \50846_nG16ab1 , RIe0a2158_5463 , \49900 , \50550 );
_HMUX g16ab2 ( \50847_nG16ab2 , RIe0a2158_5463 , \50846_nG16ab1 , \49514 );
_HMUX g16ab3 ( \50848_nG16ab3 , RIe0a2158_5463 , \49903 , \50553 );
_HMUX g16ab4 ( \50849_nG16ab4 , \50847_nG16ab2 , \50848_nG16ab3 , \49526 );
buf \U$39813 ( \50850 , \50849_nG16ab4 );
_DC g18cce_GF_IsGateDCbyConstraint ( \50851_nG18cce , \50850 , \42503 );
buf \U$39814 ( \50852 , \50851_nG18cce );
_HMUX g16ab5 ( \50853_nG16ab5 , RIe0a0010_5464 , \49909 , \50550 );
_HMUX g16ab6 ( \50854_nG16ab6 , RIe0a0010_5464 , \50853_nG16ab5 , \49514 );
_HMUX g16ab7 ( \50855_nG16ab7 , RIe0a0010_5464 , \49912 , \50553 );
_HMUX g16ab8 ( \50856_nG16ab8 , \50854_nG16ab6 , \50855_nG16ab7 , \49526 );
buf \U$39815 ( \50857 , \50856_nG16ab8 );
_DC g18cd0_GF_IsGateDCbyConstraint ( \50858_nG18cd0 , \50857 , \42503 );
buf \U$39816 ( \50859 , \50858_nG18cd0 );
_HMUX g16ab9 ( \50860_nG16ab9 , RIe09e378_5465 , \49918 , \50550 );
_HMUX g16aba ( \50861_nG16aba , RIe09e378_5465 , \50860_nG16ab9 , \49514 );
_HMUX g16abb ( \50862_nG16abb , RIe09e378_5465 , \49921 , \50553 );
_HMUX g16abc ( \50863_nG16abc , \50861_nG16aba , \50862_nG16abb , \49526 );
buf \U$39817 ( \50864 , \50863_nG16abc );
_DC g18cd2_GF_IsGateDCbyConstraint ( \50865_nG18cd2 , \50864 , \42503 );
buf \U$39818 ( \50866 , \50865_nG18cd2 );
_HMUX g16abd ( \50867_nG16abd , RIe09c668_5466 , \49927 , \50550 );
_HMUX g16abe ( \50868_nG16abe , RIe09c668_5466 , \50867_nG16abd , \49514 );
_HMUX g16abf ( \50869_nG16abf , RIe09c668_5466 , \49930 , \50553 );
_HMUX g16ac0 ( \50870_nG16ac0 , \50868_nG16abe , \50869_nG16abf , \49526 );
buf \U$39819 ( \50871 , \50870_nG16ac0 );
_DC g18cd4_GF_IsGateDCbyConstraint ( \50872_nG18cd4 , \50871 , \42503 );
buf \U$39820 ( \50873 , \50872_nG18cd4 );
_HMUX g16ac1 ( \50874_nG16ac1 , RIe09a8e0_5467 , \49936 , \50550 );
_HMUX g16ac2 ( \50875_nG16ac2 , RIe09a8e0_5467 , \50874_nG16ac1 , \49514 );
_HMUX g16ac3 ( \50876_nG16ac3 , RIe09a8e0_5467 , \49939 , \50553 );
_HMUX g16ac4 ( \50877_nG16ac4 , \50875_nG16ac2 , \50876_nG16ac3 , \49526 );
buf \U$39821 ( \50878 , \50877_nG16ac4 );
_DC g18cd6_GF_IsGateDCbyConstraint ( \50879_nG18cd6 , \50878 , \42503 );
buf \U$39822 ( \50880 , \50879_nG18cd6 );
_HMUX g16ac5 ( \50881_nG16ac5 , RIe099080_5468 , \49945 , \50550 );
_HMUX g16ac6 ( \50882_nG16ac6 , RIe099080_5468 , \50881_nG16ac5 , \49514 );
_HMUX g16ac7 ( \50883_nG16ac7 , RIe099080_5468 , \49948 , \50553 );
_HMUX g16ac8 ( \50884_nG16ac8 , \50882_nG16ac6 , \50883_nG16ac7 , \49526 );
buf \U$39823 ( \50885 , \50884_nG16ac8 );
_DC g18cd8_GF_IsGateDCbyConstraint ( \50886_nG18cd8 , \50885 , \42503 );
buf \U$39824 ( \50887 , \50886_nG18cd8 );
_HMUX g16ac9 ( \50888_nG16ac9 , RIe1d1cf8_5469 , \49954 , \50550 );
_HMUX g16aca ( \50889_nG16aca , RIe1d1cf8_5469 , \50888_nG16ac9 , \49514 );
_HMUX g16acb ( \50890_nG16acb , RIe1d1cf8_5469 , \49957 , \50553 );
_HMUX g16acc ( \50891_nG16acc , \50889_nG16aca , \50890_nG16acb , \49526 );
buf \U$39825 ( \50892 , \50891_nG16acc );
_DC g18cda_GF_IsGateDCbyConstraint ( \50893_nG18cda , \50892 , \42503 );
buf \U$39826 ( \50894 , \50893_nG18cda );
_HMUX g16acd ( \50895_nG16acd , RIe1d24f0_5470 , \49963 , \50550 );
_HMUX g16ace ( \50896_nG16ace , RIe1d24f0_5470 , \50895_nG16acd , \49514 );
_HMUX g16acf ( \50897_nG16acf , RIe1d24f0_5470 , \49966 , \50553 );
_HMUX g16ad0 ( \50898_nG16ad0 , \50896_nG16ace , \50897_nG16acf , \49526 );
buf \U$39827 ( \50899 , \50898_nG16ad0 );
_DC g18cde_GF_IsGateDCbyConstraint ( \50900_nG18cde , \50899 , \42503 );
buf \U$39828 ( \50901 , \50900_nG18cde );
_HMUX g16ad1 ( \50902_nG16ad1 , RIe1d2ce8_5471 , \49972 , \50550 );
_HMUX g16ad2 ( \50903_nG16ad2 , RIe1d2ce8_5471 , \50902_nG16ad1 , \49514 );
_HMUX g16ad3 ( \50904_nG16ad3 , RIe1d2ce8_5471 , \49975 , \50553 );
_HMUX g16ad4 ( \50905_nG16ad4 , \50903_nG16ad2 , \50904_nG16ad3 , \49526 );
buf \U$39829 ( \50906 , \50905_nG16ad4 );
_DC g18ce0_GF_IsGateDCbyConstraint ( \50907_nG18ce0 , \50906 , \42503 );
buf \U$39830 ( \50908 , \50907_nG18ce0 );
_HMUX g16ad5 ( \50909_nG16ad5 , RIe1d34e0_5472 , \49981 , \50550 );
_HMUX g16ad6 ( \50910_nG16ad6 , RIe1d34e0_5472 , \50909_nG16ad5 , \49514 );
_HMUX g16ad7 ( \50911_nG16ad7 , RIe1d34e0_5472 , \49984 , \50553 );
_HMUX g16ad8 ( \50912_nG16ad8 , \50910_nG16ad6 , \50911_nG16ad7 , \49526 );
buf \U$39831 ( \50913 , \50912_nG16ad8 );
_DC g18ce2_GF_IsGateDCbyConstraint ( \50914_nG18ce2 , \50913 , \42503 );
buf \U$39832 ( \50915 , \50914_nG18ce2 );
_HMUX g16ad9 ( \50916_nG16ad9 , RIe1d3cd8_5473 , \49990 , \50550 );
_HMUX g16ada ( \50917_nG16ada , RIe1d3cd8_5473 , \50916_nG16ad9 , \49514 );
_HMUX g16adb ( \50918_nG16adb , RIe1d3cd8_5473 , \49993 , \50553 );
_HMUX g16adc ( \50919_nG16adc , \50917_nG16ada , \50918_nG16adb , \49526 );
buf \U$39833 ( \50920 , \50919_nG16adc );
_DC g18ce4_GF_IsGateDCbyConstraint ( \50921_nG18ce4 , \50920 , \42503 );
buf \U$39834 ( \50922 , \50921_nG18ce4 );
_HMUX g16add ( \50923_nG16add , RIe1d44d0_5474 , \49999 , \50550 );
_HMUX g16ade ( \50924_nG16ade , RIe1d44d0_5474 , \50923_nG16add , \49514 );
_HMUX g16adf ( \50925_nG16adf , RIe1d44d0_5474 , \50002 , \50553 );
_HMUX g16ae0 ( \50926_nG16ae0 , \50924_nG16ade , \50925_nG16adf , \49526 );
buf \U$39835 ( \50927 , \50926_nG16ae0 );
_DC g18ce6_GF_IsGateDCbyConstraint ( \50928_nG18ce6 , \50927 , \42503 );
buf \U$39836 ( \50929 , \50928_nG18ce6 );
_HMUX g16ae1 ( \50930_nG16ae1 , RIe1d4cc8_5475 , \50008 , \50550 );
_HMUX g16ae2 ( \50931_nG16ae2 , RIe1d4cc8_5475 , \50930_nG16ae1 , \49514 );
_HMUX g16ae3 ( \50932_nG16ae3 , RIe1d4cc8_5475 , \50011 , \50553 );
_HMUX g16ae4 ( \50933_nG16ae4 , \50931_nG16ae2 , \50932_nG16ae3 , \49526 );
buf \U$39837 ( \50934 , \50933_nG16ae4 );
_DC g18ce8_GF_IsGateDCbyConstraint ( \50935_nG18ce8 , \50934 , \42503 );
buf \U$39838 ( \50936 , \50935_nG18ce8 );
_HMUX g16ae5 ( \50937_nG16ae5 , RIe1d54c0_5476 , \50017 , \50550 );
_HMUX g16ae6 ( \50938_nG16ae6 , RIe1d54c0_5476 , \50937_nG16ae5 , \49514 );
_HMUX g16ae7 ( \50939_nG16ae7 , RIe1d54c0_5476 , \50020 , \50553 );
_HMUX g16ae8 ( \50940_nG16ae8 , \50938_nG16ae6 , \50939_nG16ae7 , \49526 );
buf \U$39839 ( \50941 , \50940_nG16ae8 );
_DC g18cea_GF_IsGateDCbyConstraint ( \50942_nG18cea , \50941 , \42503 );
buf \U$39840 ( \50943 , \50942_nG18cea );
_HMUX g16ae9 ( \50944_nG16ae9 , RIe1d5cb8_5477 , \50026 , \50550 );
_HMUX g16aea ( \50945_nG16aea , RIe1d5cb8_5477 , \50944_nG16ae9 , \49514 );
_HMUX g16aeb ( \50946_nG16aeb , RIe1d5cb8_5477 , \50029 , \50553 );
_HMUX g16aec ( \50947_nG16aec , \50945_nG16aea , \50946_nG16aeb , \49526 );
buf \U$39841 ( \50948 , \50947_nG16aec );
_DC g18cec_GF_IsGateDCbyConstraint ( \50949_nG18cec , \50948 , \42503 );
buf \U$39842 ( \50950 , \50949_nG18cec );
_HMUX g16aed ( \50951_nG16aed , RIe1d64b0_5478 , \50035 , \50550 );
_HMUX g16aee ( \50952_nG16aee , RIe1d64b0_5478 , \50951_nG16aed , \49514 );
_HMUX g16aef ( \50953_nG16aef , RIe1d64b0_5478 , \50038 , \50553 );
_HMUX g16af0 ( \50954_nG16af0 , \50952_nG16aee , \50953_nG16aef , \49526 );
buf \U$39843 ( \50955 , \50954_nG16af0 );
_DC g18cee_GF_IsGateDCbyConstraint ( \50956_nG18cee , \50955 , \42503 );
buf \U$39844 ( \50957 , \50956_nG18cee );
_HMUX g16af1 ( \50958_nG16af1 , RIe1d6ca8_5479 , \50044 , \50550 );
_HMUX g16af2 ( \50959_nG16af2 , RIe1d6ca8_5479 , \50958_nG16af1 , \49514 );
_HMUX g16af3 ( \50960_nG16af3 , RIe1d6ca8_5479 , \50047 , \50553 );
_HMUX g16af4 ( \50961_nG16af4 , \50959_nG16af2 , \50960_nG16af3 , \49526 );
buf \U$39845 ( \50962 , \50961_nG16af4 );
_DC g18cf0_GF_IsGateDCbyConstraint ( \50963_nG18cf0 , \50962 , \42503 );
buf \U$39846 ( \50964 , \50963_nG18cf0 );
_HMUX g16af5 ( \50965_nG16af5 , RIe1d74a0_5480 , \50053 , \50550 );
_HMUX g16af6 ( \50966_nG16af6 , RIe1d74a0_5480 , \50965_nG16af5 , \49514 );
_HMUX g16af7 ( \50967_nG16af7 , RIe1d74a0_5480 , \50056 , \50553 );
_HMUX g16af8 ( \50968_nG16af8 , \50966_nG16af6 , \50967_nG16af7 , \49526 );
buf \U$39847 ( \50969 , \50968_nG16af8 );
_DC g18cf4_GF_IsGateDCbyConstraint ( \50970_nG18cf4 , \50969 , \42503 );
buf \U$39848 ( \50971 , \50970_nG18cf4 );
_HMUX g16af9 ( \50972_nG16af9 , RIe1d7c98_5481 , \50062 , \50550 );
_HMUX g16afa ( \50973_nG16afa , RIe1d7c98_5481 , \50972_nG16af9 , \49514 );
_HMUX g16afb ( \50974_nG16afb , RIe1d7c98_5481 , \50065 , \50553 );
_HMUX g16afc ( \50975_nG16afc , \50973_nG16afa , \50974_nG16afb , \49526 );
buf \U$39849 ( \50976 , \50975_nG16afc );
_DC g18cf6_GF_IsGateDCbyConstraint ( \50977_nG18cf6 , \50976 , \42503 );
buf \U$39850 ( \50978 , \50977_nG18cf6 );
_HMUX g16afd ( \50979_nG16afd , RIe1d8490_5482 , \50071 , \50550 );
_HMUX g16afe ( \50980_nG16afe , RIe1d8490_5482 , \50979_nG16afd , \49514 );
_HMUX g16aff ( \50981_nG16aff , RIe1d8490_5482 , \50074 , \50553 );
_HMUX g16b00 ( \50982_nG16b00 , \50980_nG16afe , \50981_nG16aff , \49526 );
buf \U$39851 ( \50983 , \50982_nG16b00 );
_DC g18cf8_GF_IsGateDCbyConstraint ( \50984_nG18cf8 , \50983 , \42503 );
buf \U$39852 ( \50985 , \50984_nG18cf8 );
_HMUX g16b01 ( \50986_nG16b01 , RIe1d8c88_5483 , \50080 , \50550 );
_HMUX g16b02 ( \50987_nG16b02 , RIe1d8c88_5483 , \50986_nG16b01 , \49514 );
_HMUX g16b03 ( \50988_nG16b03 , RIe1d8c88_5483 , \50083 , \50553 );
_HMUX g16b04 ( \50989_nG16b04 , \50987_nG16b02 , \50988_nG16b03 , \49526 );
buf \U$39853 ( \50990 , \50989_nG16b04 );
_DC g18cfa_GF_IsGateDCbyConstraint ( \50991_nG18cfa , \50990 , \42503 );
buf \U$39854 ( \50992 , \50991_nG18cfa );
_HMUX g16b05 ( \50993_nG16b05 , RIe1d9480_5484 , \50089 , \50550 );
_HMUX g16b06 ( \50994_nG16b06 , RIe1d9480_5484 , \50993_nG16b05 , \49514 );
_HMUX g16b07 ( \50995_nG16b07 , RIe1d9480_5484 , \50092 , \50553 );
_HMUX g16b08 ( \50996_nG16b08 , \50994_nG16b06 , \50995_nG16b07 , \49526 );
buf \U$39855 ( \50997 , \50996_nG16b08 );
_DC g18cfc_GF_IsGateDCbyConstraint ( \50998_nG18cfc , \50997 , \42503 );
buf \U$39856 ( \50999 , \50998_nG18cfc );
and \U$39857 ( \51000 , \49505 , \49506 );
_HMUX g16885 ( \51001_nG16885 , RIe1d9c78_5485 , \49504 , \51000 );
_HMUX g16886 ( \51002_nG16886 , RIe1d9c78_5485 , \51001_nG16885 , \49514 );
and \U$39858 ( \51003 , \49517 , \49518 );
_HMUX g1688b ( \51004_nG1688b , RIe1d9c78_5485 , \49516 , \51003 );
_HMUX g1688c ( \51005_nG1688c , \51002_nG16886 , \51004_nG1688b , \49526 );
buf \U$39859 ( \51006 , \51005_nG1688c );
_DC g18c04_GF_IsGateDCbyConstraint ( \51007_nG18c04 , \51006 , \42503 );
buf \U$39860 ( \51008 , \51007_nG18c04 );
_HMUX g1688e ( \51009_nG1688e , RIe1da470_5486 , \49531 , \51000 );
_HMUX g1688f ( \51010_nG1688f , RIe1da470_5486 , \51009_nG1688e , \49514 );
_HMUX g16891 ( \51011_nG16891 , RIe1da470_5486 , \49534 , \51003 );
_HMUX g16892 ( \51012_nG16892 , \51010_nG1688f , \51011_nG16891 , \49526 );
buf \U$39861 ( \51013 , \51012_nG16892 );
_DC g18c1a_GF_IsGateDCbyConstraint ( \51014_nG18c1a , \51013 , \42503 );
buf \U$39862 ( \51015 , \51014_nG18c1a );
_HMUX g16894 ( \51016_nG16894 , RIe1dac68_5487 , \49540 , \51000 );
_HMUX g16895 ( \51017_nG16895 , RIe1dac68_5487 , \51016_nG16894 , \49514 );
_HMUX g16897 ( \51018_nG16897 , RIe1dac68_5487 , \49543 , \51003 );
_HMUX g16898 ( \51019_nG16898 , \51017_nG16895 , \51018_nG16897 , \49526 );
buf \U$39863 ( \51020 , \51019_nG16898 );
_DC g18c30_GF_IsGateDCbyConstraint ( \51021_nG18c30 , \51020 , \42503 );
buf \U$39864 ( \51022 , \51021_nG18c30 );
_HMUX g1689a ( \51023_nG1689a , RIe1db460_5488 , \49549 , \51000 );
_HMUX g1689b ( \51024_nG1689b , RIe1db460_5488 , \51023_nG1689a , \49514 );
_HMUX g1689d ( \51025_nG1689d , RIe1db460_5488 , \49552 , \51003 );
_HMUX g1689e ( \51026_nG1689e , \51024_nG1689b , \51025_nG1689d , \49526 );
buf \U$39865 ( \51027 , \51026_nG1689e );
_DC g18c46_GF_IsGateDCbyConstraint ( \51028_nG18c46 , \51027 , \42503 );
buf \U$39866 ( \51029 , \51028_nG18c46 );
_HMUX g168a0 ( \51030_nG168a0 , RIe1dbc58_5489 , \49558 , \51000 );
_HMUX g168a1 ( \51031_nG168a1 , RIe1dbc58_5489 , \51030_nG168a0 , \49514 );
_HMUX g168a3 ( \51032_nG168a3 , RIe1dbc58_5489 , \49561 , \51003 );
_HMUX g168a4 ( \51033_nG168a4 , \51031_nG168a1 , \51032_nG168a3 , \49526 );
buf \U$39867 ( \51034 , \51033_nG168a4 );
_DC g18c5c_GF_IsGateDCbyConstraint ( \51035_nG18c5c , \51034 , \42503 );
buf \U$39868 ( \51036 , \51035_nG18c5c );
_HMUX g168a6 ( \51037_nG168a6 , RIe1dc450_5490 , \49567 , \51000 );
_HMUX g168a7 ( \51038_nG168a7 , RIe1dc450_5490 , \51037_nG168a6 , \49514 );
_HMUX g168a9 ( \51039_nG168a9 , RIe1dc450_5490 , \49570 , \51003 );
_HMUX g168aa ( \51040_nG168aa , \51038_nG168a7 , \51039_nG168a9 , \49526 );
buf \U$39869 ( \51041 , \51040_nG168aa );
_DC g18c72_GF_IsGateDCbyConstraint ( \51042_nG18c72 , \51041 , \42503 );
buf \U$39870 ( \51043 , \51042_nG18c72 );
_HMUX g168ac ( \51044_nG168ac , RIe1dcc48_5491 , \49576 , \51000 );
_HMUX g168ad ( \51045_nG168ad , RIe1dcc48_5491 , \51044_nG168ac , \49514 );
_HMUX g168af ( \51046_nG168af , RIe1dcc48_5491 , \49579 , \51003 );
_HMUX g168b0 ( \51047_nG168b0 , \51045_nG168ad , \51046_nG168af , \49526 );
buf \U$39871 ( \51048 , \51047_nG168b0 );
_DC g18c7e_GF_IsGateDCbyConstraint ( \51049_nG18c7e , \51048 , \42503 );
buf \U$39872 ( \51050 , \51049_nG18c7e );
_HMUX g168b2 ( \51051_nG168b2 , RIe1dd440_5492 , \49585 , \51000 );
_HMUX g168b3 ( \51052_nG168b3 , RIe1dd440_5492 , \51051_nG168b2 , \49514 );
_HMUX g168b5 ( \51053_nG168b5 , RIe1dd440_5492 , \49588 , \51003 );
_HMUX g168b6 ( \51054_nG168b6 , \51052_nG168b3 , \51053_nG168b5 , \49526 );
buf \U$39873 ( \51055 , \51054_nG168b6 );
_DC g18c80_GF_IsGateDCbyConstraint ( \51056_nG18c80 , \51055 , \42503 );
buf \U$39874 ( \51057 , \51056_nG18c80 );
_HMUX g168b8 ( \51058_nG168b8 , RIe1ddc38_5493 , \49594 , \51000 );
_HMUX g168b9 ( \51059_nG168b9 , RIe1ddc38_5493 , \51058_nG168b8 , \49514 );
_HMUX g168bb ( \51060_nG168bb , RIe1ddc38_5493 , \49597 , \51003 );
_HMUX g168bc ( \51061_nG168bc , \51059_nG168b9 , \51060_nG168bb , \49526 );
buf \U$39875 ( \51062 , \51061_nG168bc );
_DC g18c82_GF_IsGateDCbyConstraint ( \51063_nG18c82 , \51062 , \42503 );
buf \U$39876 ( \51064 , \51063_nG18c82 );
_HMUX g168be ( \51065_nG168be , RIe1de430_5494 , \49603 , \51000 );
_HMUX g168bf ( \51066_nG168bf , RIe1de430_5494 , \51065_nG168be , \49514 );
_HMUX g168c1 ( \51067_nG168c1 , RIe1de430_5494 , \49606 , \51003 );
_HMUX g168c2 ( \51068_nG168c2 , \51066_nG168bf , \51067_nG168c1 , \49526 );
buf \U$39877 ( \51069 , \51068_nG168c2 );
_DC g18c06_GF_IsGateDCbyConstraint ( \51070_nG18c06 , \51069 , \42503 );
buf \U$39878 ( \51071 , \51070_nG18c06 );
_HMUX g168c4 ( \51072_nG168c4 , RIe1dec28_5495 , \49612 , \51000 );
_HMUX g168c5 ( \51073_nG168c5 , RIe1dec28_5495 , \51072_nG168c4 , \49514 );
_HMUX g168c7 ( \51074_nG168c7 , RIe1dec28_5495 , \49615 , \51003 );
_HMUX g168c8 ( \51075_nG168c8 , \51073_nG168c5 , \51074_nG168c7 , \49526 );
buf \U$39879 ( \51076 , \51075_nG168c8 );
_DC g18c08_GF_IsGateDCbyConstraint ( \51077_nG18c08 , \51076 , \42503 );
buf \U$39880 ( \51078 , \51077_nG18c08 );
_HMUX g168ca ( \51079_nG168ca , RIe1df420_5496 , \49621 , \51000 );
_HMUX g168cb ( \51080_nG168cb , RIe1df420_5496 , \51079_nG168ca , \49514 );
_HMUX g168cd ( \51081_nG168cd , RIe1df420_5496 , \49624 , \51003 );
_HMUX g168ce ( \51082_nG168ce , \51080_nG168cb , \51081_nG168cd , \49526 );
buf \U$39881 ( \51083 , \51082_nG168ce );
_DC g18c0a_GF_IsGateDCbyConstraint ( \51084_nG18c0a , \51083 , \42503 );
buf \U$39882 ( \51085 , \51084_nG18c0a );
_HMUX g168d0 ( \51086_nG168d0 , RIe1dfc18_5497 , \49630 , \51000 );
_HMUX g168d1 ( \51087_nG168d1 , RIe1dfc18_5497 , \51086_nG168d0 , \49514 );
_HMUX g168d3 ( \51088_nG168d3 , RIe1dfc18_5497 , \49633 , \51003 );
_HMUX g168d4 ( \51089_nG168d4 , \51087_nG168d1 , \51088_nG168d3 , \49526 );
buf \U$39883 ( \51090 , \51089_nG168d4 );
_DC g18c0c_GF_IsGateDCbyConstraint ( \51091_nG18c0c , \51090 , \42503 );
buf \U$39884 ( \51092 , \51091_nG18c0c );
_HMUX g168d6 ( \51093_nG168d6 , RIe1e0410_5498 , \49639 , \51000 );
_HMUX g168d7 ( \51094_nG168d7 , RIe1e0410_5498 , \51093_nG168d6 , \49514 );
_HMUX g168d9 ( \51095_nG168d9 , RIe1e0410_5498 , \49642 , \51003 );
_HMUX g168da ( \51096_nG168da , \51094_nG168d7 , \51095_nG168d9 , \49526 );
buf \U$39885 ( \51097 , \51096_nG168da );
_DC g18c0e_GF_IsGateDCbyConstraint ( \51098_nG18c0e , \51097 , \42503 );
buf \U$39886 ( \51099 , \51098_nG18c0e );
_HMUX g168dc ( \51100_nG168dc , RIe1e0c08_5499 , \49648 , \51000 );
_HMUX g168dd ( \51101_nG168dd , RIe1e0c08_5499 , \51100_nG168dc , \49514 );
_HMUX g168df ( \51102_nG168df , RIe1e0c08_5499 , \49651 , \51003 );
_HMUX g168e0 ( \51103_nG168e0 , \51101_nG168dd , \51102_nG168df , \49526 );
buf \U$39887 ( \51104 , \51103_nG168e0 );
_DC g18c10_GF_IsGateDCbyConstraint ( \51105_nG18c10 , \51104 , \42503 );
buf \U$39888 ( \51106 , \51105_nG18c10 );
_HMUX g168e2 ( \51107_nG168e2 , RIe1e1400_5500 , \49657 , \51000 );
_HMUX g168e3 ( \51108_nG168e3 , RIe1e1400_5500 , \51107_nG168e2 , \49514 );
_HMUX g168e5 ( \51109_nG168e5 , RIe1e1400_5500 , \49660 , \51003 );
_HMUX g168e6 ( \51110_nG168e6 , \51108_nG168e3 , \51109_nG168e5 , \49526 );
buf \U$39889 ( \51111 , \51110_nG168e6 );
_DC g18c12_GF_IsGateDCbyConstraint ( \51112_nG18c12 , \51111 , \42503 );
buf \U$39890 ( \51113 , \51112_nG18c12 );
_HMUX g168e8 ( \51114_nG168e8 , RIe1e1bf8_5501 , \49666 , \51000 );
_HMUX g168e9 ( \51115_nG168e9 , RIe1e1bf8_5501 , \51114_nG168e8 , \49514 );
_HMUX g168eb ( \51116_nG168eb , RIe1e1bf8_5501 , \49669 , \51003 );
_HMUX g168ec ( \51117_nG168ec , \51115_nG168e9 , \51116_nG168eb , \49526 );
buf \U$39891 ( \51118 , \51117_nG168ec );
_DC g18c14_GF_IsGateDCbyConstraint ( \51119_nG18c14 , \51118 , \42503 );
buf \U$39892 ( \51120 , \51119_nG18c14 );
_HMUX g168ee ( \51121_nG168ee , RIe1e23f0_5502 , \49675 , \51000 );
_HMUX g168ef ( \51122_nG168ef , RIe1e23f0_5502 , \51121_nG168ee , \49514 );
_HMUX g168f1 ( \51123_nG168f1 , RIe1e23f0_5502 , \49678 , \51003 );
_HMUX g168f2 ( \51124_nG168f2 , \51122_nG168ef , \51123_nG168f1 , \49526 );
buf \U$39893 ( \51125 , \51124_nG168f2 );
_DC g18c16_GF_IsGateDCbyConstraint ( \51126_nG18c16 , \51125 , \42503 );
buf \U$39894 ( \51127 , \51126_nG18c16 );
_HMUX g168f4 ( \51128_nG168f4 , RIe1e2be8_5503 , \49684 , \51000 );
_HMUX g168f5 ( \51129_nG168f5 , RIe1e2be8_5503 , \51128_nG168f4 , \49514 );
_HMUX g168f7 ( \51130_nG168f7 , RIe1e2be8_5503 , \49687 , \51003 );
_HMUX g168f8 ( \51131_nG168f8 , \51129_nG168f5 , \51130_nG168f7 , \49526 );
buf \U$39895 ( \51132 , \51131_nG168f8 );
_DC g18c18_GF_IsGateDCbyConstraint ( \51133_nG18c18 , \51132 , \42503 );
buf \U$39896 ( \51134 , \51133_nG18c18 );
_HMUX g168fa ( \51135_nG168fa , RIe1e33e0_5504 , \49693 , \51000 );
_HMUX g168fb ( \51136_nG168fb , RIe1e33e0_5504 , \51135_nG168fa , \49514 );
_HMUX g168fd ( \51137_nG168fd , RIe1e33e0_5504 , \49696 , \51003 );
_HMUX g168fe ( \51138_nG168fe , \51136_nG168fb , \51137_nG168fd , \49526 );
buf \U$39897 ( \51139 , \51138_nG168fe );
_DC g18c1c_GF_IsGateDCbyConstraint ( \51140_nG18c1c , \51139 , \42503 );
buf \U$39898 ( \51141 , \51140_nG18c1c );
_HMUX g16900 ( \51142_nG16900 , RIe1e3bd8_5505 , \49702 , \51000 );
_HMUX g16901 ( \51143_nG16901 , RIe1e3bd8_5505 , \51142_nG16900 , \49514 );
_HMUX g16903 ( \51144_nG16903 , RIe1e3bd8_5505 , \49705 , \51003 );
_HMUX g16904 ( \51145_nG16904 , \51143_nG16901 , \51144_nG16903 , \49526 );
buf \U$39899 ( \51146 , \51145_nG16904 );
_DC g18c1e_GF_IsGateDCbyConstraint ( \51147_nG18c1e , \51146 , \42503 );
buf \U$39900 ( \51148 , \51147_nG18c1e );
_HMUX g16906 ( \51149_nG16906 , RIe1e43d0_5506 , \49711 , \51000 );
_HMUX g16907 ( \51150_nG16907 , RIe1e43d0_5506 , \51149_nG16906 , \49514 );
_HMUX g16909 ( \51151_nG16909 , RIe1e43d0_5506 , \49714 , \51003 );
_HMUX g1690a ( \51152_nG1690a , \51150_nG16907 , \51151_nG16909 , \49526 );
buf \U$39901 ( \51153 , \51152_nG1690a );
_DC g18c20_GF_IsGateDCbyConstraint ( \51154_nG18c20 , \51153 , \42503 );
buf \U$39902 ( \51155 , \51154_nG18c20 );
_HMUX g1690c ( \51156_nG1690c , RIe1e4bc8_5507 , \49720 , \51000 );
_HMUX g1690d ( \51157_nG1690d , RIe1e4bc8_5507 , \51156_nG1690c , \49514 );
_HMUX g1690f ( \51158_nG1690f , RIe1e4bc8_5507 , \49723 , \51003 );
_HMUX g16910 ( \51159_nG16910 , \51157_nG1690d , \51158_nG1690f , \49526 );
buf \U$39903 ( \51160 , \51159_nG16910 );
_DC g18c22_GF_IsGateDCbyConstraint ( \51161_nG18c22 , \51160 , \42503 );
buf \U$39904 ( \51162 , \51161_nG18c22 );
_HMUX g16912 ( \51163_nG16912 , RIe1e53c0_5508 , \49729 , \51000 );
_HMUX g16913 ( \51164_nG16913 , RIe1e53c0_5508 , \51163_nG16912 , \49514 );
_HMUX g16915 ( \51165_nG16915 , RIe1e53c0_5508 , \49732 , \51003 );
_HMUX g16916 ( \51166_nG16916 , \51164_nG16913 , \51165_nG16915 , \49526 );
buf \U$39905 ( \51167 , \51166_nG16916 );
_DC g18c24_GF_IsGateDCbyConstraint ( \51168_nG18c24 , \51167 , \42503 );
buf \U$39906 ( \51169 , \51168_nG18c24 );
_HMUX g16918 ( \51170_nG16918 , RIe1e5bb8_5509 , \49738 , \51000 );
_HMUX g16919 ( \51171_nG16919 , RIe1e5bb8_5509 , \51170_nG16918 , \49514 );
_HMUX g1691b ( \51172_nG1691b , RIe1e5bb8_5509 , \49741 , \51003 );
_HMUX g1691c ( \51173_nG1691c , \51171_nG16919 , \51172_nG1691b , \49526 );
buf \U$39907 ( \51174 , \51173_nG1691c );
_DC g18c26_GF_IsGateDCbyConstraint ( \51175_nG18c26 , \51174 , \42503 );
buf \U$39908 ( \51176 , \51175_nG18c26 );
_HMUX g1691e ( \51177_nG1691e , RIe1e63b0_5510 , \49747 , \51000 );
_HMUX g1691f ( \51178_nG1691f , RIe1e63b0_5510 , \51177_nG1691e , \49514 );
_HMUX g16921 ( \51179_nG16921 , RIe1e63b0_5510 , \49750 , \51003 );
_HMUX g16922 ( \51180_nG16922 , \51178_nG1691f , \51179_nG16921 , \49526 );
buf \U$39909 ( \51181 , \51180_nG16922 );
_DC g18c28_GF_IsGateDCbyConstraint ( \51182_nG18c28 , \51181 , \42503 );
buf \U$39910 ( \51183 , \51182_nG18c28 );
_HMUX g16924 ( \51184_nG16924 , RIe1e6ba8_5511 , \49756 , \51000 );
_HMUX g16925 ( \51185_nG16925 , RIe1e6ba8_5511 , \51184_nG16924 , \49514 );
_HMUX g16927 ( \51186_nG16927 , RIe1e6ba8_5511 , \49759 , \51003 );
_HMUX g16928 ( \51187_nG16928 , \51185_nG16925 , \51186_nG16927 , \49526 );
buf \U$39911 ( \51188 , \51187_nG16928 );
_DC g18c2a_GF_IsGateDCbyConstraint ( \51189_nG18c2a , \51188 , \42503 );
buf \U$39912 ( \51190 , \51189_nG18c2a );
_HMUX g1692a ( \51191_nG1692a , RIe1e73a0_5512 , \49765 , \51000 );
_HMUX g1692b ( \51192_nG1692b , RIe1e73a0_5512 , \51191_nG1692a , \49514 );
_HMUX g1692d ( \51193_nG1692d , RIe1e73a0_5512 , \49768 , \51003 );
_HMUX g1692e ( \51194_nG1692e , \51192_nG1692b , \51193_nG1692d , \49526 );
buf \U$39913 ( \51195 , \51194_nG1692e );
_DC g18c2c_GF_IsGateDCbyConstraint ( \51196_nG18c2c , \51195 , \42503 );
buf \U$39914 ( \51197 , \51196_nG18c2c );
_HMUX g16930 ( \51198_nG16930 , RIe1e7b98_5513 , \49774 , \51000 );
_HMUX g16931 ( \51199_nG16931 , RIe1e7b98_5513 , \51198_nG16930 , \49514 );
_HMUX g16933 ( \51200_nG16933 , RIe1e7b98_5513 , \49777 , \51003 );
_HMUX g16934 ( \51201_nG16934 , \51199_nG16931 , \51200_nG16933 , \49526 );
buf \U$39915 ( \51202 , \51201_nG16934 );
_DC g18c2e_GF_IsGateDCbyConstraint ( \51203_nG18c2e , \51202 , \42503 );
buf \U$39916 ( \51204 , \51203_nG18c2e );
_HMUX g16936 ( \51205_nG16936 , RIe1e8390_5514 , \49783 , \51000 );
_HMUX g16937 ( \51206_nG16937 , RIe1e8390_5514 , \51205_nG16936 , \49514 );
_HMUX g16939 ( \51207_nG16939 , RIe1e8390_5514 , \49786 , \51003 );
_HMUX g1693a ( \51208_nG1693a , \51206_nG16937 , \51207_nG16939 , \49526 );
buf \U$39917 ( \51209 , \51208_nG1693a );
_DC g18c32_GF_IsGateDCbyConstraint ( \51210_nG18c32 , \51209 , \42503 );
buf \U$39918 ( \51211 , \51210_nG18c32 );
_HMUX g1693c ( \51212_nG1693c , RIe1e8b88_5515 , \49792 , \51000 );
_HMUX g1693d ( \51213_nG1693d , RIe1e8b88_5515 , \51212_nG1693c , \49514 );
_HMUX g1693f ( \51214_nG1693f , RIe1e8b88_5515 , \49795 , \51003 );
_HMUX g16940 ( \51215_nG16940 , \51213_nG1693d , \51214_nG1693f , \49526 );
buf \U$39919 ( \51216 , \51215_nG16940 );
_DC g18c34_GF_IsGateDCbyConstraint ( \51217_nG18c34 , \51216 , \42503 );
buf \U$39920 ( \51218 , \51217_nG18c34 );
_HMUX g16942 ( \51219_nG16942 , RIe1e9380_5516 , \49801 , \51000 );
_HMUX g16943 ( \51220_nG16943 , RIe1e9380_5516 , \51219_nG16942 , \49514 );
_HMUX g16945 ( \51221_nG16945 , RIe1e9380_5516 , \49804 , \51003 );
_HMUX g16946 ( \51222_nG16946 , \51220_nG16943 , \51221_nG16945 , \49526 );
buf \U$39921 ( \51223 , \51222_nG16946 );
_DC g18c36_GF_IsGateDCbyConstraint ( \51224_nG18c36 , \51223 , \42503 );
buf \U$39922 ( \51225 , \51224_nG18c36 );
_HMUX g16948 ( \51226_nG16948 , RIe1e9b78_5517 , \49810 , \51000 );
_HMUX g16949 ( \51227_nG16949 , RIe1e9b78_5517 , \51226_nG16948 , \49514 );
_HMUX g1694b ( \51228_nG1694b , RIe1e9b78_5517 , \49813 , \51003 );
_HMUX g1694c ( \51229_nG1694c , \51227_nG16949 , \51228_nG1694b , \49526 );
buf \U$39923 ( \51230 , \51229_nG1694c );
_DC g18c38_GF_IsGateDCbyConstraint ( \51231_nG18c38 , \51230 , \42503 );
buf \U$39924 ( \51232 , \51231_nG18c38 );
_HMUX g1694e ( \51233_nG1694e , RIe1ea370_5518 , \49819 , \51000 );
_HMUX g1694f ( \51234_nG1694f , RIe1ea370_5518 , \51233_nG1694e , \49514 );
_HMUX g16951 ( \51235_nG16951 , RIe1ea370_5518 , \49822 , \51003 );
_HMUX g16952 ( \51236_nG16952 , \51234_nG1694f , \51235_nG16951 , \49526 );
buf \U$39925 ( \51237 , \51236_nG16952 );
_DC g18c3a_GF_IsGateDCbyConstraint ( \51238_nG18c3a , \51237 , \42503 );
buf \U$39926 ( \51239 , \51238_nG18c3a );
_HMUX g16954 ( \51240_nG16954 , RIe1eab68_5519 , \49828 , \51000 );
_HMUX g16955 ( \51241_nG16955 , RIe1eab68_5519 , \51240_nG16954 , \49514 );
_HMUX g16957 ( \51242_nG16957 , RIe1eab68_5519 , \49831 , \51003 );
_HMUX g16958 ( \51243_nG16958 , \51241_nG16955 , \51242_nG16957 , \49526 );
buf \U$39927 ( \51244 , \51243_nG16958 );
_DC g18c3c_GF_IsGateDCbyConstraint ( \51245_nG18c3c , \51244 , \42503 );
buf \U$39928 ( \51246 , \51245_nG18c3c );
_HMUX g1695a ( \51247_nG1695a , RIe1eb360_5520 , \49837 , \51000 );
_HMUX g1695b ( \51248_nG1695b , RIe1eb360_5520 , \51247_nG1695a , \49514 );
_HMUX g1695d ( \51249_nG1695d , RIe1eb360_5520 , \49840 , \51003 );
_HMUX g1695e ( \51250_nG1695e , \51248_nG1695b , \51249_nG1695d , \49526 );
buf \U$39929 ( \51251 , \51250_nG1695e );
_DC g18c3e_GF_IsGateDCbyConstraint ( \51252_nG18c3e , \51251 , \42503 );
buf \U$39930 ( \51253 , \51252_nG18c3e );
_HMUX g16960 ( \51254_nG16960 , RIe1ebb58_5521 , \49846 , \51000 );
_HMUX g16961 ( \51255_nG16961 , RIe1ebb58_5521 , \51254_nG16960 , \49514 );
_HMUX g16963 ( \51256_nG16963 , RIe1ebb58_5521 , \49849 , \51003 );
_HMUX g16964 ( \51257_nG16964 , \51255_nG16961 , \51256_nG16963 , \49526 );
buf \U$39931 ( \51258 , \51257_nG16964 );
_DC g18c40_GF_IsGateDCbyConstraint ( \51259_nG18c40 , \51258 , \42503 );
buf \U$39932 ( \51260 , \51259_nG18c40 );
_HMUX g16966 ( \51261_nG16966 , RIe1ec350_5522 , \49855 , \51000 );
_HMUX g16967 ( \51262_nG16967 , RIe1ec350_5522 , \51261_nG16966 , \49514 );
_HMUX g16969 ( \51263_nG16969 , RIe1ec350_5522 , \49858 , \51003 );
_HMUX g1696a ( \51264_nG1696a , \51262_nG16967 , \51263_nG16969 , \49526 );
buf \U$39933 ( \51265 , \51264_nG1696a );
_DC g18c42_GF_IsGateDCbyConstraint ( \51266_nG18c42 , \51265 , \42503 );
buf \U$39934 ( \51267 , \51266_nG18c42 );
_HMUX g1696c ( \51268_nG1696c , RIe1ecb48_5523 , \49864 , \51000 );
_HMUX g1696d ( \51269_nG1696d , RIe1ecb48_5523 , \51268_nG1696c , \49514 );
_HMUX g1696f ( \51270_nG1696f , RIe1ecb48_5523 , \49867 , \51003 );
_HMUX g16970 ( \51271_nG16970 , \51269_nG1696d , \51270_nG1696f , \49526 );
buf \U$39935 ( \51272 , \51271_nG16970 );
_DC g18c44_GF_IsGateDCbyConstraint ( \51273_nG18c44 , \51272 , \42503 );
buf \U$39936 ( \51274 , \51273_nG18c44 );
_HMUX g16972 ( \51275_nG16972 , RIe1ed340_5524 , \49873 , \51000 );
_HMUX g16973 ( \51276_nG16973 , RIe1ed340_5524 , \51275_nG16972 , \49514 );
_HMUX g16975 ( \51277_nG16975 , RIe1ed340_5524 , \49876 , \51003 );
_HMUX g16976 ( \51278_nG16976 , \51276_nG16973 , \51277_nG16975 , \49526 );
buf \U$39937 ( \51279 , \51278_nG16976 );
_DC g18c48_GF_IsGateDCbyConstraint ( \51280_nG18c48 , \51279 , \42503 );
buf \U$39938 ( \51281 , \51280_nG18c48 );
_HMUX g16978 ( \51282_nG16978 , RIe1edb38_5525 , \49882 , \51000 );
_HMUX g16979 ( \51283_nG16979 , RIe1edb38_5525 , \51282_nG16978 , \49514 );
_HMUX g1697b ( \51284_nG1697b , RIe1edb38_5525 , \49885 , \51003 );
_HMUX g1697c ( \51285_nG1697c , \51283_nG16979 , \51284_nG1697b , \49526 );
buf \U$39939 ( \51286 , \51285_nG1697c );
_DC g18c4a_GF_IsGateDCbyConstraint ( \51287_nG18c4a , \51286 , \42503 );
buf \U$39940 ( \51288 , \51287_nG18c4a );
_HMUX g1697e ( \51289_nG1697e , RIe1ee330_5526 , \49891 , \51000 );
_HMUX g1697f ( \51290_nG1697f , RIe1ee330_5526 , \51289_nG1697e , \49514 );
_HMUX g16981 ( \51291_nG16981 , RIe1ee330_5526 , \49894 , \51003 );
_HMUX g16982 ( \51292_nG16982 , \51290_nG1697f , \51291_nG16981 , \49526 );
buf \U$39941 ( \51293 , \51292_nG16982 );
_DC g18c4c_GF_IsGateDCbyConstraint ( \51294_nG18c4c , \51293 , \42503 );
buf \U$39942 ( \51295 , \51294_nG18c4c );
_HMUX g16984 ( \51296_nG16984 , RIe1eeb28_5527 , \49900 , \51000 );
_HMUX g16985 ( \51297_nG16985 , RIe1eeb28_5527 , \51296_nG16984 , \49514 );
_HMUX g16987 ( \51298_nG16987 , RIe1eeb28_5527 , \49903 , \51003 );
_HMUX g16988 ( \51299_nG16988 , \51297_nG16985 , \51298_nG16987 , \49526 );
buf \U$39943 ( \51300 , \51299_nG16988 );
_DC g18c4e_GF_IsGateDCbyConstraint ( \51301_nG18c4e , \51300 , \42503 );
buf \U$39944 ( \51302 , \51301_nG18c4e );
_HMUX g1698a ( \51303_nG1698a , RIe1ef320_5528 , \49909 , \51000 );
_HMUX g1698b ( \51304_nG1698b , RIe1ef320_5528 , \51303_nG1698a , \49514 );
_HMUX g1698d ( \51305_nG1698d , RIe1ef320_5528 , \49912 , \51003 );
_HMUX g1698e ( \51306_nG1698e , \51304_nG1698b , \51305_nG1698d , \49526 );
buf \U$39945 ( \51307 , \51306_nG1698e );
_DC g18c50_GF_IsGateDCbyConstraint ( \51308_nG18c50 , \51307 , \42503 );
buf \U$39946 ( \51309 , \51308_nG18c50 );
_HMUX g16990 ( \51310_nG16990 , RIe1efb18_5529 , \49918 , \51000 );
_HMUX g16991 ( \51311_nG16991 , RIe1efb18_5529 , \51310_nG16990 , \49514 );
_HMUX g16993 ( \51312_nG16993 , RIe1efb18_5529 , \49921 , \51003 );
_HMUX g16994 ( \51313_nG16994 , \51311_nG16991 , \51312_nG16993 , \49526 );
buf \U$39947 ( \51314 , \51313_nG16994 );
_DC g18c52_GF_IsGateDCbyConstraint ( \51315_nG18c52 , \51314 , \42503 );
buf \U$39948 ( \51316 , \51315_nG18c52 );
_HMUX g16996 ( \51317_nG16996 , RIe1f0310_5530 , \49927 , \51000 );
_HMUX g16997 ( \51318_nG16997 , RIe1f0310_5530 , \51317_nG16996 , \49514 );
_HMUX g16999 ( \51319_nG16999 , RIe1f0310_5530 , \49930 , \51003 );
_HMUX g1699a ( \51320_nG1699a , \51318_nG16997 , \51319_nG16999 , \49526 );
buf \U$39949 ( \51321 , \51320_nG1699a );
_DC g18c54_GF_IsGateDCbyConstraint ( \51322_nG18c54 , \51321 , \42503 );
buf \U$39950 ( \51323 , \51322_nG18c54 );
_HMUX g1699c ( \51324_nG1699c , RIe1f0b08_5531 , \49936 , \51000 );
_HMUX g1699d ( \51325_nG1699d , RIe1f0b08_5531 , \51324_nG1699c , \49514 );
_HMUX g1699f ( \51326_nG1699f , RIe1f0b08_5531 , \49939 , \51003 );
_HMUX g169a0 ( \51327_nG169a0 , \51325_nG1699d , \51326_nG1699f , \49526 );
buf \U$39951 ( \51328 , \51327_nG169a0 );
_DC g18c56_GF_IsGateDCbyConstraint ( \51329_nG18c56 , \51328 , \42503 );
buf \U$39952 ( \51330 , \51329_nG18c56 );
_HMUX g169a2 ( \51331_nG169a2 , RIe1f1300_5532 , \49945 , \51000 );
_HMUX g169a3 ( \51332_nG169a3 , RIe1f1300_5532 , \51331_nG169a2 , \49514 );
_HMUX g169a5 ( \51333_nG169a5 , RIe1f1300_5532 , \49948 , \51003 );
_HMUX g169a6 ( \51334_nG169a6 , \51332_nG169a3 , \51333_nG169a5 , \49526 );
buf \U$39953 ( \51335 , \51334_nG169a6 );
_DC g18c58_GF_IsGateDCbyConstraint ( \51336_nG18c58 , \51335 , \42503 );
buf \U$39954 ( \51337 , \51336_nG18c58 );
_HMUX g169a8 ( \51338_nG169a8 , RIe1f1af8_5533 , \49954 , \51000 );
_HMUX g169a9 ( \51339_nG169a9 , RIe1f1af8_5533 , \51338_nG169a8 , \49514 );
_HMUX g169ab ( \51340_nG169ab , RIe1f1af8_5533 , \49957 , \51003 );
_HMUX g169ac ( \51341_nG169ac , \51339_nG169a9 , \51340_nG169ab , \49526 );
buf \U$39955 ( \51342 , \51341_nG169ac );
_DC g18c5a_GF_IsGateDCbyConstraint ( \51343_nG18c5a , \51342 , \42503 );
buf \U$39956 ( \51344 , \51343_nG18c5a );
_HMUX g169ae ( \51345_nG169ae , RIe1f22f0_5534 , \49963 , \51000 );
_HMUX g169af ( \51346_nG169af , RIe1f22f0_5534 , \51345_nG169ae , \49514 );
_HMUX g169b1 ( \51347_nG169b1 , RIe1f22f0_5534 , \49966 , \51003 );
_HMUX g169b2 ( \51348_nG169b2 , \51346_nG169af , \51347_nG169b1 , \49526 );
buf \U$39957 ( \51349 , \51348_nG169b2 );
_DC g18c5e_GF_IsGateDCbyConstraint ( \51350_nG18c5e , \51349 , \42503 );
buf \U$39958 ( \51351 , \51350_nG18c5e );
_HMUX g169b4 ( \51352_nG169b4 , RIe1f2ae8_5535 , \49972 , \51000 );
_HMUX g169b5 ( \51353_nG169b5 , RIe1f2ae8_5535 , \51352_nG169b4 , \49514 );
_HMUX g169b7 ( \51354_nG169b7 , RIe1f2ae8_5535 , \49975 , \51003 );
_HMUX g169b8 ( \51355_nG169b8 , \51353_nG169b5 , \51354_nG169b7 , \49526 );
buf \U$39959 ( \51356 , \51355_nG169b8 );
_DC g18c60_GF_IsGateDCbyConstraint ( \51357_nG18c60 , \51356 , \42503 );
buf \U$39960 ( \51358 , \51357_nG18c60 );
_HMUX g169ba ( \51359_nG169ba , RIe1f32e0_5536 , \49981 , \51000 );
_HMUX g169bb ( \51360_nG169bb , RIe1f32e0_5536 , \51359_nG169ba , \49514 );
_HMUX g169bd ( \51361_nG169bd , RIe1f32e0_5536 , \49984 , \51003 );
_HMUX g169be ( \51362_nG169be , \51360_nG169bb , \51361_nG169bd , \49526 );
buf \U$39961 ( \51363 , \51362_nG169be );
_DC g18c62_GF_IsGateDCbyConstraint ( \51364_nG18c62 , \51363 , \42503 );
buf \U$39962 ( \51365 , \51364_nG18c62 );
_HMUX g169c0 ( \51366_nG169c0 , RIe1f3ad8_5537 , \49990 , \51000 );
_HMUX g169c1 ( \51367_nG169c1 , RIe1f3ad8_5537 , \51366_nG169c0 , \49514 );
_HMUX g169c3 ( \51368_nG169c3 , RIe1f3ad8_5537 , \49993 , \51003 );
_HMUX g169c4 ( \51369_nG169c4 , \51367_nG169c1 , \51368_nG169c3 , \49526 );
buf \U$39963 ( \51370 , \51369_nG169c4 );
_DC g18c64_GF_IsGateDCbyConstraint ( \51371_nG18c64 , \51370 , \42503 );
buf \U$39964 ( \51372 , \51371_nG18c64 );
_HMUX g169c6 ( \51373_nG169c6 , RIe1f42d0_5538 , \49999 , \51000 );
_HMUX g169c7 ( \51374_nG169c7 , RIe1f42d0_5538 , \51373_nG169c6 , \49514 );
_HMUX g169c9 ( \51375_nG169c9 , RIe1f42d0_5538 , \50002 , \51003 );
_HMUX g169ca ( \51376_nG169ca , \51374_nG169c7 , \51375_nG169c9 , \49526 );
buf \U$39965 ( \51377 , \51376_nG169ca );
_DC g18c66_GF_IsGateDCbyConstraint ( \51378_nG18c66 , \51377 , \42503 );
buf \U$39966 ( \51379 , \51378_nG18c66 );
_HMUX g169cc ( \51380_nG169cc , RIe1f4ac8_5539 , \50008 , \51000 );
_HMUX g169cd ( \51381_nG169cd , RIe1f4ac8_5539 , \51380_nG169cc , \49514 );
_HMUX g169cf ( \51382_nG169cf , RIe1f4ac8_5539 , \50011 , \51003 );
_HMUX g169d0 ( \51383_nG169d0 , \51381_nG169cd , \51382_nG169cf , \49526 );
buf \U$39967 ( \51384 , \51383_nG169d0 );
_DC g18c68_GF_IsGateDCbyConstraint ( \51385_nG18c68 , \51384 , \42503 );
buf \U$39968 ( \51386 , \51385_nG18c68 );
_HMUX g169d2 ( \51387_nG169d2 , RIe1f52c0_5540 , \50017 , \51000 );
_HMUX g169d3 ( \51388_nG169d3 , RIe1f52c0_5540 , \51387_nG169d2 , \49514 );
_HMUX g169d5 ( \51389_nG169d5 , RIe1f52c0_5540 , \50020 , \51003 );
_HMUX g169d6 ( \51390_nG169d6 , \51388_nG169d3 , \51389_nG169d5 , \49526 );
buf \U$39969 ( \51391 , \51390_nG169d6 );
_DC g18c6a_GF_IsGateDCbyConstraint ( \51392_nG18c6a , \51391 , \42503 );
buf \U$39970 ( \51393 , \51392_nG18c6a );
_HMUX g169d8 ( \51394_nG169d8 , RIe1f5ab8_5541 , \50026 , \51000 );
_HMUX g169d9 ( \51395_nG169d9 , RIe1f5ab8_5541 , \51394_nG169d8 , \49514 );
_HMUX g169db ( \51396_nG169db , RIe1f5ab8_5541 , \50029 , \51003 );
_HMUX g169dc ( \51397_nG169dc , \51395_nG169d9 , \51396_nG169db , \49526 );
buf \U$39971 ( \51398 , \51397_nG169dc );
_DC g18c6c_GF_IsGateDCbyConstraint ( \51399_nG18c6c , \51398 , \42503 );
buf \U$39972 ( \51400 , \51399_nG18c6c );
_HMUX g169de ( \51401_nG169de , RIe1f62b0_5542 , \50035 , \51000 );
_HMUX g169df ( \51402_nG169df , RIe1f62b0_5542 , \51401_nG169de , \49514 );
_HMUX g169e1 ( \51403_nG169e1 , RIe1f62b0_5542 , \50038 , \51003 );
_HMUX g169e2 ( \51404_nG169e2 , \51402_nG169df , \51403_nG169e1 , \49526 );
buf \U$39973 ( \51405 , \51404_nG169e2 );
_DC g18c6e_GF_IsGateDCbyConstraint ( \51406_nG18c6e , \51405 , \42503 );
buf \U$39974 ( \51407 , \51406_nG18c6e );
_HMUX g169e4 ( \51408_nG169e4 , RIe1f6aa8_5543 , \50044 , \51000 );
_HMUX g169e5 ( \51409_nG169e5 , RIe1f6aa8_5543 , \51408_nG169e4 , \49514 );
_HMUX g169e7 ( \51410_nG169e7 , RIe1f6aa8_5543 , \50047 , \51003 );
_HMUX g169e8 ( \51411_nG169e8 , \51409_nG169e5 , \51410_nG169e7 , \49526 );
buf \U$39975 ( \51412 , \51411_nG169e8 );
_DC g18c70_GF_IsGateDCbyConstraint ( \51413_nG18c70 , \51412 , \42503 );
buf \U$39976 ( \51414 , \51413_nG18c70 );
_HMUX g169ea ( \51415_nG169ea , RIe1f72a0_5544 , \50053 , \51000 );
_HMUX g169eb ( \51416_nG169eb , RIe1f72a0_5544 , \51415_nG169ea , \49514 );
_HMUX g169ed ( \51417_nG169ed , RIe1f72a0_5544 , \50056 , \51003 );
_HMUX g169ee ( \51418_nG169ee , \51416_nG169eb , \51417_nG169ed , \49526 );
buf \U$39977 ( \51419 , \51418_nG169ee );
_DC g18c74_GF_IsGateDCbyConstraint ( \51420_nG18c74 , \51419 , \42503 );
buf \U$39978 ( \51421 , \51420_nG18c74 );
_HMUX g169f0 ( \51422_nG169f0 , RIe1f7a98_5545 , \50062 , \51000 );
_HMUX g169f1 ( \51423_nG169f1 , RIe1f7a98_5545 , \51422_nG169f0 , \49514 );
_HMUX g169f3 ( \51424_nG169f3 , RIe1f7a98_5545 , \50065 , \51003 );
_HMUX g169f4 ( \51425_nG169f4 , \51423_nG169f1 , \51424_nG169f3 , \49526 );
buf \U$39979 ( \51426 , \51425_nG169f4 );
_DC g18c76_GF_IsGateDCbyConstraint ( \51427_nG18c76 , \51426 , \42503 );
buf \U$39980 ( \51428 , \51427_nG18c76 );
_HMUX g169f6 ( \51429_nG169f6 , RIe1f8290_5546 , \50071 , \51000 );
_HMUX g169f7 ( \51430_nG169f7 , RIe1f8290_5546 , \51429_nG169f6 , \49514 );
_HMUX g169f9 ( \51431_nG169f9 , RIe1f8290_5546 , \50074 , \51003 );
_HMUX g169fa ( \51432_nG169fa , \51430_nG169f7 , \51431_nG169f9 , \49526 );
buf \U$39981 ( \51433 , \51432_nG169fa );
_DC g18c78_GF_IsGateDCbyConstraint ( \51434_nG18c78 , \51433 , \42503 );
buf \U$39982 ( \51435 , \51434_nG18c78 );
_HMUX g169fc ( \51436_nG169fc , RIe1f8a88_5547 , \50080 , \51000 );
_HMUX g169fd ( \51437_nG169fd , RIe1f8a88_5547 , \51436_nG169fc , \49514 );
_HMUX g169ff ( \51438_nG169ff , RIe1f8a88_5547 , \50083 , \51003 );
_HMUX g16a00 ( \51439_nG16a00 , \51437_nG169fd , \51438_nG169ff , \49526 );
buf \U$39983 ( \51440 , \51439_nG16a00 );
_DC g18c7a_GF_IsGateDCbyConstraint ( \51441_nG18c7a , \51440 , \42503 );
buf \U$39984 ( \51442 , \51441_nG18c7a );
_HMUX g16a02 ( \51443_nG16a02 , RIe1f9280_5548 , \50089 , \51000 );
_HMUX g16a03 ( \51444_nG16a03 , RIe1f9280_5548 , \51443_nG16a02 , \49514 );
_HMUX g16a05 ( \51445_nG16a05 , RIe1f9280_5548 , \50092 , \51003 );
_HMUX g16a06 ( \51446_nG16a06 , \51444_nG16a03 , \51445_nG16a05 , \49526 );
buf \U$39985 ( \51447 , \51446_nG16a06 );
_DC g18c7c_GF_IsGateDCbyConstraint ( \51448_nG18c7c , \51447 , \42503 );
buf \U$39986 ( \51449 , \51448_nG18c7c );
buf \U$39987 ( \51450 , RIb86fc68_77);
_HMUX g16857 ( \51451_nG16857 , RIe137870_5261 , \51450 , \49507 );
not \U$39988 ( \51452 , \49514 );
or \U$39989 ( \51453 , \49526 , \51452 );
_HMUX g16858 ( \51454_nG16858 , \51451_nG16857 , RIe137870_5261 , \51453 );
buf \U$39990 ( \51455 , \51454_nG16858 );
_DC g18bec_GF_IsGateDCbyConstraint ( \51456_nG18bec , \51455 , \42503 );
buf \U$39991 ( \51457 , \51456_nG18bec );
buf \U$39992 ( \51458 , RIb86fce0_76);
_HMUX g16859 ( \51459_nG16859 , RIe136da8_5262 , \51458 , \49507 );
_HMUX g1685a ( \51460_nG1685a , \51459_nG16859 , RIe136da8_5262 , \51453 );
buf \U$39993 ( \51461 , \51460_nG1685a );
_DC g18bee_GF_IsGateDCbyConstraint ( \51462_nG18bee , \51461 , \42503 );
buf \U$39994 ( \51463 , \51462_nG18bee );
buf \U$39995 ( \51464 , RIb86fd58_75);
_HMUX g1685b ( \51465_nG1685b , RIe136358_5263 , \51464 , \49507 );
_HMUX g1685c ( \51466_nG1685c , \51465_nG1685b , RIe136358_5263 , \51453 );
buf \U$39996 ( \51467 , \51466_nG1685c );
_DC g18bf0_GF_IsGateDCbyConstraint ( \51468_nG18bf0 , \51467 , \42503 );
buf \U$39997 ( \51469 , \51468_nG18bf0 );
buf \U$39998 ( \51470 , RIb87e8a8_74);
_HMUX g1685d ( \51471_nG1685d , RIe135890_5264 , \51470 , \49507 );
_HMUX g1685e ( \51472_nG1685e , \51471_nG1685d , RIe135890_5264 , \51453 );
buf \U$39999 ( \51473 , \51472_nG1685e );
_DC g18bf2_GF_IsGateDCbyConstraint ( \51474_nG18bf2 , \51473 , \42503 );
buf \U$40000 ( \51475 , \51474_nG18bf2 );
buf \U$40001 ( \51476 , RIb87e920_73);
_HMUX g1685f ( \51477_nG1685f , RIe134d50_5265 , \51476 , \49507 );
_HMUX g16860 ( \51478_nG16860 , \51477_nG1685f , RIe134d50_5265 , \51453 );
buf \U$40002 ( \51479 , \51478_nG16860 );
_DC g18bf4_GF_IsGateDCbyConstraint ( \51480_nG18bf4 , \51479 , \42503 );
buf \U$40003 ( \51481 , \51480_nG18bf4 );
buf \U$40004 ( \51482 , RIb87e998_72);
_HMUX g16861 ( \51483_nG16861 , RIe134288_5266 , \51482 , \49507 );
_HMUX g16862 ( \51484_nG16862 , \51483_nG16861 , RIe134288_5266 , \51453 );
buf \U$40005 ( \51485 , \51484_nG16862 );
_DC g18bf6_GF_IsGateDCbyConstraint ( \51486_nG18bf6 , \51485 , \42503 );
buf \U$40006 ( \51487 , \51486_nG18bf6 );
buf \U$40007 ( \51488 , RIb87ea10_71);
_HMUX g16863 ( \51489_nG16863 , RIe1337c0_5267 , \51488 , \49507 );
_HMUX g16864 ( \51490_nG16864 , \51489_nG16863 , RIe1337c0_5267 , \51453 );
buf \U$40008 ( \51491 , \51490_nG16864 );
_DC g18bf8_GF_IsGateDCbyConstraint ( \51492_nG18bf8 , \51491 , \42503 );
buf \U$40009 ( \51493 , \51492_nG18bf8 );
buf \U$40010 ( \51494 , RIb87ea88_70);
_HMUX g16865 ( \51495_nG16865 , RIe132c08_5268 , \51494 , \49507 );
_HMUX g16866 ( \51496_nG16866 , \51495_nG16865 , RIe132c08_5268 , \51453 );
buf \U$40011 ( \51497 , \51496_nG16866 );
_DC g18bfa_GF_IsGateDCbyConstraint ( \51498_nG18bfa , \51497 , \42503 );
buf \U$40012 ( \51499 , \51498_nG18bfa );
_HMUX g16846 ( \51500_nG16846 , RIe131fd8_5269 , \51450 , \50099 );
_HMUX g16847 ( \51501_nG16847 , \51500_nG16846 , RIe131fd8_5269 , \51453 );
buf \U$40013 ( \51502 , \51501_nG16847 );
_DC g18bdc_GF_IsGateDCbyConstraint ( \51503_nG18bdc , \51502 , \42503 );
buf \U$40014 ( \51504 , \51503_nG18bdc );
_HMUX g16848 ( \51505_nG16848 , RIe1313a8_5270 , \51458 , \50099 );
_HMUX g16849 ( \51506_nG16849 , \51505_nG16848 , RIe1313a8_5270 , \51453 );
buf \U$40015 ( \51507 , \51506_nG16849 );
_DC g18bde_GF_IsGateDCbyConstraint ( \51508_nG18bde , \51507 , \42503 );
buf \U$40016 ( \51509 , \51508_nG18bde );
_HMUX g1684a ( \51510_nG1684a , RIe1307f0_5271 , \51464 , \50099 );
_HMUX g1684b ( \51511_nG1684b , \51510_nG1684a , RIe1307f0_5271 , \51453 );
buf \U$40017 ( \51512 , \51511_nG1684b );
_DC g18be0_GF_IsGateDCbyConstraint ( \51513_nG18be0 , \51512 , \42503 );
buf \U$40018 ( \51514 , \51513_nG18be0 );
_HMUX g1684c ( \51515_nG1684c , RIe12fbc0_5272 , \51470 , \50099 );
_HMUX g1684d ( \51516_nG1684d , \51515_nG1684c , RIe12fbc0_5272 , \51453 );
buf \U$40019 ( \51517 , \51516_nG1684d );
_DC g18be2_GF_IsGateDCbyConstraint ( \51518_nG18be2 , \51517 , \42503 );
buf \U$40020 ( \51519 , \51518_nG18be2 );
_HMUX g1684e ( \51520_nG1684e , RIe12f080_5273 , \51476 , \50099 );
_HMUX g1684f ( \51521_nG1684f , \51520_nG1684e , RIe12f080_5273 , \51453 );
buf \U$40021 ( \51522 , \51521_nG1684f );
_DC g18be4_GF_IsGateDCbyConstraint ( \51523_nG18be4 , \51522 , \42503 );
buf \U$40022 ( \51524 , \51523_nG18be4 );
_HMUX g16850 ( \51525_nG16850 , RIe12da78_5274 , \51482 , \50099 );
_HMUX g16851 ( \51526_nG16851 , \51525_nG16850 , RIe12da78_5274 , \51453 );
buf \U$40023 ( \51527 , \51526_nG16851 );
_DC g18be6_GF_IsGateDCbyConstraint ( \51528_nG18be6 , \51527 , \42503 );
buf \U$40024 ( \51529 , \51528_nG18be6 );
_HMUX g16852 ( \51530_nG16852 , RIe12c920_5275 , \51488 , \50099 );
_HMUX g16853 ( \51531_nG16853 , \51530_nG16852 , RIe12c920_5275 , \51453 );
buf \U$40025 ( \51532 , \51531_nG16853 );
_DC g18be8_GF_IsGateDCbyConstraint ( \51533_nG18be8 , \51532 , \42503 );
buf \U$40026 ( \51534 , \51533_nG18be8 );
_HMUX g16854 ( \51535_nG16854 , RIe12b318_5276 , \51494 , \50099 );
_HMUX g16855 ( \51536_nG16855 , \51535_nG16854 , RIe12b318_5276 , \51453 );
buf \U$40027 ( \51537 , \51536_nG16855 );
_DC g18bea_GF_IsGateDCbyConstraint ( \51538_nG18bea , \51537 , \42503 );
buf \U$40028 ( \51539 , \51538_nG18bea );
_HMUX g16835 ( \51540_nG16835 , RIe12a1c0_5277 , \51450 , \50550 );
_HMUX g16836 ( \51541_nG16836 , \51540_nG16835 , RIe12a1c0_5277 , \51453 );
buf \U$40029 ( \51542 , \51541_nG16836 );
_DC g18bcc_GF_IsGateDCbyConstraint ( \51543_nG18bcc , \51542 , \42503 );
buf \U$40030 ( \51544 , \51543_nG18bcc );
_HMUX g16837 ( \51545_nG16837 , RIe128bb8_5278 , \51458 , \50550 );
_HMUX g16838 ( \51546_nG16838 , \51545_nG16837 , RIe128bb8_5278 , \51453 );
buf \U$40031 ( \51547 , \51546_nG16838 );
_DC g18bce_GF_IsGateDCbyConstraint ( \51548_nG18bce , \51547 , \42503 );
buf \U$40032 ( \51549 , \51548_nG18bce );
_HMUX g16839 ( \51550_nG16839 , RIe127a60_5279 , \51464 , \50550 );
_HMUX g1683a ( \51551_nG1683a , \51550_nG16839 , RIe127a60_5279 , \51453 );
buf \U$40033 ( \51552 , \51551_nG1683a );
_DC g18bd0_GF_IsGateDCbyConstraint ( \51553_nG18bd0 , \51552 , \42503 );
buf \U$40034 ( \51554 , \51553_nG18bd0 );
_HMUX g1683b ( \51555_nG1683b , RIe126908_5280 , \51470 , \50550 );
_HMUX g1683c ( \51556_nG1683c , \51555_nG1683b , RIe126908_5280 , \51453 );
buf \U$40035 ( \51557 , \51556_nG1683c );
_DC g18bd2_GF_IsGateDCbyConstraint ( \51558_nG18bd2 , \51557 , \42503 );
buf \U$40036 ( \51559 , \51558_nG18bd2 );
_HMUX g1683d ( \51560_nG1683d , RIe125300_5281 , \51476 , \50550 );
_HMUX g1683e ( \51561_nG1683e , \51560_nG1683d , RIe125300_5281 , \51453 );
buf \U$40037 ( \51562 , \51561_nG1683e );
_DC g18bd4_GF_IsGateDCbyConstraint ( \51563_nG18bd4 , \51562 , \42503 );
buf \U$40038 ( \51564 , \51563_nG18bd4 );
_HMUX g1683f ( \51565_nG1683f , RIe1241a8_5282 , \51482 , \50550 );
_HMUX g16840 ( \51566_nG16840 , \51565_nG1683f , RIe1241a8_5282 , \51453 );
buf \U$40039 ( \51567 , \51566_nG16840 );
_DC g18bd6_GF_IsGateDCbyConstraint ( \51568_nG18bd6 , \51567 , \42503 );
buf \U$40040 ( \51569 , \51568_nG18bd6 );
_HMUX g16841 ( \51570_nG16841 , RIe122ba0_5283 , \51488 , \50550 );
_HMUX g16842 ( \51571_nG16842 , \51570_nG16841 , RIe122ba0_5283 , \51453 );
buf \U$40041 ( \51572 , \51571_nG16842 );
_DC g18bd8_GF_IsGateDCbyConstraint ( \51573_nG18bd8 , \51572 , \42503 );
buf \U$40042 ( \51574 , \51573_nG18bd8 );
_HMUX g16843 ( \51575_nG16843 , RIe121a48_5284 , \51494 , \50550 );
_HMUX g16844 ( \51576_nG16844 , \51575_nG16843 , RIe121a48_5284 , \51453 );
buf \U$40043 ( \51577 , \51576_nG16844 );
_DC g18bda_GF_IsGateDCbyConstraint ( \51578_nG18bda , \51577 , \42503 );
buf \U$40044 ( \51579 , \51578_nG18bda );
_HMUX g16814 ( \51580_nG16814 , RIe120440_5285 , \51450 , \51000 );
_HMUX g1681d ( \51581_nG1681d , \51580_nG16814 , RIe120440_5285 , \51453 );
buf \U$40045 ( \51582 , \51581_nG1681d );
_DC g18e04_GF_IsGateDCbyConstraint ( \51583_nG18e04 , \51582 , \42503 );
buf \U$40046 ( \51584 , \51583_nG18e04 );
_HMUX g1681f ( \51585_nG1681f , RIe11f2e8_5286 , \51458 , \51000 );
_HMUX g16820 ( \51586_nG16820 , \51585_nG1681f , RIe11f2e8_5286 , \51453 );
buf \U$40047 ( \51587 , \51586_nG16820 );
_DC g18e06_GF_IsGateDCbyConstraint ( \51588_nG18e06 , \51587 , \42503 );
buf \U$40048 ( \51589 , \51588_nG18e06 );
_HMUX g16822 ( \51590_nG16822 , RIe11e190_5287 , \51464 , \51000 );
_HMUX g16823 ( \51591_nG16823 , \51590_nG16822 , RIe11e190_5287 , \51453 );
buf \U$40049 ( \51592 , \51591_nG16823 );
_DC g18e08_GF_IsGateDCbyConstraint ( \51593_nG18e08 , \51592 , \42503 );
buf \U$40050 ( \51594 , \51593_nG18e08 );
_HMUX g16825 ( \51595_nG16825 , RIe11cb88_5288 , \51470 , \51000 );
_HMUX g16826 ( \51596_nG16826 , \51595_nG16825 , RIe11cb88_5288 , \51453 );
buf \U$40051 ( \51597 , \51596_nG16826 );
_DC g18e0a_GF_IsGateDCbyConstraint ( \51598_nG18e0a , \51597 , \42503 );
buf \U$40052 ( \51599 , \51598_nG18e0a );
_HMUX g16828 ( \51600_nG16828 , RIe11ba30_5289 , \51476 , \51000 );
_HMUX g16829 ( \51601_nG16829 , \51600_nG16828 , RIe11ba30_5289 , \51453 );
buf \U$40053 ( \51602 , \51601_nG16829 );
_DC g18e0c_GF_IsGateDCbyConstraint ( \51603_nG18e0c , \51602 , \42503 );
buf \U$40054 ( \51604 , \51603_nG18e0c );
_HMUX g1682b ( \51605_nG1682b , RIe11a428_5290 , \51482 , \51000 );
_HMUX g1682c ( \51606_nG1682c , \51605_nG1682b , RIe11a428_5290 , \51453 );
buf \U$40055 ( \51607 , \51606_nG1682c );
_DC g18e0e_GF_IsGateDCbyConstraint ( \51608_nG18e0e , \51607 , \42503 );
buf \U$40056 ( \51609 , \51608_nG18e0e );
_HMUX g1682e ( \51610_nG1682e , RIe1192d0_5291 , \51488 , \51000 );
_HMUX g1682f ( \51611_nG1682f , \51610_nG1682e , RIe1192d0_5291 , \51453 );
buf \U$40057 ( \51612 , \51611_nG1682f );
_DC g18e10_GF_IsGateDCbyConstraint ( \51613_nG18e10 , \51612 , \42503 );
buf \U$40058 ( \51614 , \51613_nG18e10 );
_HMUX g16831 ( \51615_nG16831 , RIe117cc8_5292 , \51494 , \51000 );
_HMUX g16832 ( \51616_nG16832 , \51615_nG16831 , RIe117cc8_5292 , \51453 );
buf \U$40059 ( \51617 , \51616_nG16832 );
_DC g18e12_GF_IsGateDCbyConstraint ( \51618_nG18e12 , \51617 , \42503 );
buf \U$40060 ( \51619 , \51618_nG18e12 );
buf \U$40061 ( \51620 , RIb7b9680_245);
buf \U$40062 ( \51621 , RIb79b3b0_273);
and \U$40063 ( \51622 , \49522 , \51621 );
_HMUX g16709 ( \51623_nG16709 , RIe38a110_5575 , \51620 , \51622 );
buf \U$40064 ( \51624 , \51623_nG16709 );
_DC g18e13_GF_IsGateDCbyConstraint ( \51625_nG18e13 , \51624 , \42503 );
buf \U$40065 ( \51626 , \51625_nG18e13 );
buf \U$40066 ( \51627 , RIb7b96f8_244);
_HMUX g16776 ( \51628_nG16776 , RIe378410_5590 , \51627 , \51622 );
buf \U$40067 ( \51629 , \51628_nG16776 );
_DC g18bb0_GF_IsGateDCbyConstraint ( \51630_nG18bb0 , \51629 , \42503 );
buf \U$40068 ( \51631 , \51630_nG18bb0 );
buf \U$40069 ( \51632 , RIb7c20c8_243);
_HMUX g16778 ( \51633_nG16778 , RIe379220_5589 , \51632 , \51622 );
buf \U$40070 ( \51634 , \51633_nG16778 );
_DC g18bb2_GF_IsGateDCbyConstraint ( \51635_nG18bb2 , \51634 , \42503 );
buf \U$40071 ( \51636 , \51635_nG18bb2 );
buf \U$40072 ( \51637 , RIb7c5728_242);
_HMUX g1677a ( \51638_nG1677a , RIe379e50_5588 , \51637 , \51622 );
buf \U$40073 ( \51639 , \51638_nG1677a );
_DC g18bb4_GF_IsGateDCbyConstraint ( \51640_nG18bb4 , \51639 , \42503 );
buf \U$40074 ( \51641 , \51640_nG18bb4 );
buf \U$40075 ( \51642 , RIb7c57a0_241);
_HMUX g1677c ( \51643_nG1677c , RIe26f4f8_5601 , \51642 , \51622 );
buf \U$40076 ( \51644 , \51643_nG1677c );
_DC g18bb6_GF_IsGateDCbyConstraint ( \51645_nG18bb6 , \51644 , \42503 );
buf \U$40077 ( \51646 , \51645_nG18bb6 );
buf \U$40078 ( \51647 , RIb7c5818_240);
_HMUX g1677e ( \51648_nG1677e , RIe270290_5600 , \51647 , \51622 );
buf \U$40079 ( \51649 , \51648_nG1677e );
_DC g18bb8_GF_IsGateDCbyConstraint ( \51650_nG18bb8 , \51649 , \42503 );
buf \U$40080 ( \51651 , \51650_nG18bb8 );
buf \U$40081 ( \51652 , RIb7c5890_239);
_HMUX g16780 ( \51653_nG16780 , RIe270ec0_5599 , \51652 , \51622 );
buf \U$40082 ( \51654 , \51653_nG16780 );
_DC g18bba_GF_IsGateDCbyConstraint ( \51655_nG18bba , \51654 , \42503 );
buf \U$40083 ( \51656 , \51655_nG18bba );
buf \U$40084 ( \51657 , RIb7c5908_238);
_HMUX g16782 ( \51658_nG16782 , RIe271be0_5598 , \51657 , \51622 );
buf \U$40085 ( \51659 , \51658_nG16782 );
_DC g18bbc_GF_IsGateDCbyConstraint ( \51660_nG18bbc , \51659 , \42503 );
buf \U$40086 ( \51661 , \51660_nG18bbc );
buf \U$40087 ( \51662 , RIb7a09f0_266);
_HMUX g16774 ( \51663_nG16774 , RIe37b908_5586 , \51662 , \51622 );
buf \U$40088 ( \51664 , \51663_nG16774 );
_DC g18bae_GF_IsGateDCbyConstraint ( \51665_nG18bae , \51664 , \42503 );
buf \U$40089 ( \51666 , \51665_nG18bae );
buf \U$40090 ( \51667 , RIb7a0a68_265);
_HMUX g1676c ( \51668_nG1676c , RIe375008_5594 , \51667 , \51622 );
buf \U$40091 ( \51669 , \51668_nG1676c );
_DC g18ba6_GF_IsGateDCbyConstraint ( \51670_nG18ba6 , \51669 , \42503 );
buf \U$40092 ( \51671 , \51670_nG18ba6 );
buf \U$40093 ( \51672 , RIb7a0ae0_264);
_HMUX g1676e ( \51673_nG1676e , RIe375da0_5593 , \51672 , \51622 );
buf \U$40094 ( \51674 , \51673_nG1676e );
_DC g18ba8_GF_IsGateDCbyConstraint ( \51675_nG18ba8 , \51674 , \42503 );
buf \U$40095 ( \51676 , \51675_nG18ba8 );
buf \U$40096 ( \51677 , RIb7a0b58_263);
_HMUX g16770 ( \51678_nG16770 , RIe376a48_5592 , \51677 , \51622 );
buf \U$40097 ( \51679 , \51678_nG16770 );
_DC g18baa_GF_IsGateDCbyConstraint ( \51680_nG18baa , \51679 , \42503 );
buf \U$40098 ( \51681 , \51680_nG18baa );
buf \U$40099 ( \51682 , RIb7a0bd0_262);
_HMUX g16772 ( \51683_nG16772 , RIe377768_5591 , \51682 , \51622 );
buf \U$40100 ( \51684 , \51683_nG16772 );
_DC g18bac_GF_IsGateDCbyConstraint ( \51685_nG18bac , \51684 , \42503 );
buf \U$40101 ( \51686 , \51685_nG18bac );
buf \U$40102 ( \51687 , RIe3921f8_5562);
not \U$40103 ( \51688 , \51687 );
buf \U$40104 ( \51689 , \51688 );
nor \U$40106 ( \51690 , RIe3921f8_5562, RIe392b58_5561, RIe3934b8_5560);
_HMUX g165dc ( \51691_nG165dc , \51689 , 1'b0 , \51690 );
and \U$40107 ( \51692 , RIe5319e0_6884, \7061 , RIe549770_6843, RIe548ff0_6844, \7063 );
buf \U$40108 ( \51693 , \51692 );
buf \U$40109 ( \51694 , RIb79b4a0_271);
and \U$40110 ( \51695 , \51693 , \51694 );
_HMUX g165dd ( \51696_nG165dd , RIe3921f8_5562 , \51691_nG165dc , \51695 );
buf \U$40111 ( \51697 , RIe3921f8_5562);
not \U$40112 ( \51698 , \51697 );
buf \U$40113 ( \51699 , \51698 );
not \U$40114 ( \51700 , RIe3934b8_5560);
nor \U$40115 ( \51701 , RIe3921f8_5562, RIe392b58_5561, \51700 );
_HMUX g165e3 ( \51702_nG165e3 , \51699 , RIe3921f8_5562 , \51701 );
and \U$40116 ( \51703 , \49524 , \49522 );
_HMUX g165e7 ( \51704_nG165e7 , \51696_nG165dd , \51702_nG165e3 , \51703 );
and \U$40117 ( \51705 , \51703 , \51694 );
and \U$40118 ( \51706 , \51705 , \51693 );
_HMUX g165ea ( \51707_nG165ea , \51704_nG165e7 , RIe3921f8_5562 , \51706 );
not \U$40119 ( \51708 , RIe37f9b8_5584);
and \U$40120 ( \51709 , RIe37f9b8_5584, \51620 );
or \U$40121 ( \51710 , \51708 , \51709 );
and \U$40122 ( \51711 , \51710 , \49524 );
and \U$40123 ( \51712 , \51711 , \49522 );
_HMUX g165f1 ( \51713_nG165f1 , \51707_nG165ea , RIe38a908_5574 , \51712 );
buf \U$40125 ( \51714 , RIb79b338_274);
and \U$40126 ( \51715 , \51693 , \51714 );
_HMUX g165f2 ( \51716_nG165f2 , \51713_nG165f1 , 1'b0 , \51715 );
buf \U$40127 ( \51717 , \51716_nG165f2 );
buf \U$40128 ( \51718 , RIe392b58_5561);
xnor \U$40129 ( \51719 , \51718 , \51687 );
buf \U$40130 ( \51720 , \51719 );
_HMUX g165f6 ( \51721_nG165f6 , \51720 , 1'b0 , \51690 );
_HMUX g165f7 ( \51722_nG165f7 , RIe392b58_5561 , \51721_nG165f6 , \51695 );
buf \U$40132 ( \51723 , RIe392b58_5561);
xor \U$40133 ( \51724 , \51723 , \51697 );
buf \U$40134 ( \51725 , \51724 );
_HMUX g165fb ( \51726_nG165fb , \51725 , RIe392b58_5561 , \51701 );
_HMUX g165fc ( \51727_nG165fc , \51722_nG165f7 , \51726_nG165fb , \51703 );
_HMUX g165fd ( \51728_nG165fd , \51727_nG165fc , RIe392b58_5561 , \51706 );
_HMUX g165fe ( \51729_nG165fe , \51728_nG165fd , RIe38b1f0_5573 , \51712 );
_HMUX g165ff ( \51730_nG165ff , \51729_nG165fe , 1'b0 , \51715 );
buf \U$40136 ( \51731 , \51730_nG165ff );
buf \U$40137 ( \51732 , RIe3934b8_5560);
or \U$40138 ( \51733 , \51718 , \51687 );
xnor \U$40139 ( \51734 , \51732 , \51733 );
buf \U$40140 ( \51735 , \51734 );
_HMUX g16604 ( \51736_nG16604 , \51735 , 1'b0 , \51690 );
_HMUX g16605 ( \51737_nG16605 , RIe3934b8_5560 , \51736_nG16604 , \51695 );
buf \U$40142 ( \51738 , RIe3934b8_5560);
and \U$40143 ( \51739 , \51723 , \51697 );
xor \U$40144 ( \51740 , \51738 , \51739 );
buf \U$40145 ( \51741 , \51740 );
_HMUX g1660a ( \51742_nG1660a , \51741 , RIe3934b8_5560 , \51701 );
_HMUX g1660b ( \51743_nG1660b , \51737_nG16605 , \51742_nG1660a , \51703 );
_HMUX g1660c ( \51744_nG1660c , \51743_nG1660b , RIe3934b8_5560 , \51706 );
_HMUX g1660d ( \51745_nG1660d , \51744_nG1660c , RIe38b9e8_5572 , \51712 );
_HMUX g1660e ( \51746_nG1660e , \51745_nG1660d , 1'b0 , \51715 );
buf \U$40147 ( \51747 , \51746_nG1660e );
or \U$40148 ( \51748 , \51717 , \51731 , \51747 );
buf \U$40149 ( \51749 , \51748 );
buf \U$40150 ( \51750 , RIe3951c8_5557);
buf \U$40151 ( \51751 , RIe394868_5558);
buf \U$40152 ( \51752 , RIe393e90_5559);
and \U$40153 ( \51753 , \51751 , \51752 );
xor \U$40154 ( \51754 , \51750 , \51753 );
buf \U$40155 ( \51755 , \51754 );
not \U$40156 ( \51756 , RIe3951c8_5557);
nor \U$40157 ( \51757 , RIe393e90_5559, RIe394868_5558, \51756 );
not \U$40158 ( \51758 , \51757 );
and \U$40159 ( \51759 , \51695 , \51758 );
_HMUX g165d3 ( \51760_nG165d3 , RIe3951c8_5557 , \51755 , \51759 );
_HMUX g165d4 ( \51761_nG165d4 , \51760_nG165d3 , 1'b0 , \51715 );
buf \U$40161 ( \51762 , \51761_nG165d4 );
not \U$40162 ( \51763 , \51762 );
buf \U$40163 ( \51764 , RIe38da40_5569);
buf \U$40164 ( \51765 , RIe38cf78_5570);
buf \U$40165 ( \51766 , RIe38c4b0_5571);
and \U$40166 ( \51767 , \51765 , \51766 );
xor \U$40167 ( \51768 , \51764 , \51767 );
buf \U$40168 ( \51769 , \51768 );
buf \U$40169 ( \51770 , RIb839848_152);
and \U$40170 ( \51771 , \49510 , \51770 );
not \U$40171 ( \51772 , RIe38cf78_5570);
and \U$40172 ( \51773 , RIe38c4b0_5571, \51772 , RIe38da40_5569);
not \U$40173 ( \51774 , \51773 );
and \U$40174 ( \51775 , \51771 , \51774 );
_HMUX g16691 ( \51776_nG16691 , RIe38da40_5569 , \51769 , \51775 );
buf \U$40175 ( \51777 , RIe38da40_5569);
buf \U$40176 ( \51778 , RIe38cf78_5570);
xor \U$40177 ( \51779 , \51777 , \51778 );
buf \U$40178 ( \51780 , \51779 );
not \U$40179 ( \51781 , RIe38c4b0_5571);
and \U$40180 ( \51782 , \51781 , \51772 , RIe38da40_5569);
or \U$40181 ( \51783 , \51782 , \51773 );
_HMUX g16695 ( \51784_nG16695 , \51780 , RIe38da40_5569 , \51783 );
buf \U$40182 ( \51785 , RIb839668_156);
and \U$40183 ( \51786 , \49510 , \51785 );
_HMUX g16696 ( \51787_nG16696 , \51776_nG16691 , \51784_nG16695 , \51786 );
buf \U$40185 ( \51788 , RIb8396e0_155);
and \U$40186 ( \51789 , \49510 , \51788 );
_HMUX g16697 ( \51790_nG16697 , \51787_nG16696 , 1'b0 , \51789 );
and \U$40188 ( \51791 , \51789 , \51785 );
_HMUX g16698 ( \51792_nG16698 , \51790_nG16697 , 1'b0 , \51791 );
buf \U$40189 ( \51793 , \51792_nG16698 );
and \U$40190 ( \51794 , \51763 , \51793 );
xor \U$40191 ( \51795 , \51751 , \51752 );
buf \U$40192 ( \51796 , \51795 );
_HMUX g165cd ( \51797_nG165cd , RIe394868_5558 , \51796 , \51759 );
_HMUX g165ce ( \51798_nG165ce , \51797_nG165cd , 1'b0 , \51715 );
buf \U$40194 ( \51799 , \51798_nG165ce );
not \U$40195 ( \51800 , \51799 );
xor \U$40196 ( \51801 , \51765 , \51766 );
buf \U$40197 ( \51802 , \51801 );
_HMUX g16682 ( \51803_nG16682 , RIe38cf78_5570 , \51802 , \51775 );
not \U$40198 ( \51804 , \51778 );
buf \U$40199 ( \51805 , \51804 );
_HMUX g16689 ( \51806_nG16689 , \51805 , RIe38cf78_5570 , \51783 );
_HMUX g1668a ( \51807_nG1668a , \51803_nG16682 , \51806_nG16689 , \51786 );
_HMUX g1668b ( \51808_nG1668b , \51807_nG1668a , 1'b0 , \51789 );
_HMUX g1668c ( \51809_nG1668c , \51808_nG1668b , 1'b1 , \51791 );
buf \U$40202 ( \51810 , \51809_nG1668c );
and \U$40203 ( \51811 , \51800 , \51810 );
not \U$40204 ( \51812 , \51752 );
buf \U$40205 ( \51813 , \51812 );
_HMUX g165c6 ( \51814_nG165c6 , RIe393e90_5559 , \51813 , \51759 );
_HMUX g165c9 ( \51815_nG165c9 , \51814_nG165c6 , 1'b0 , \51715 );
buf \U$40207 ( \51816 , \51815_nG165c9 );
not \U$40208 ( \51817 , \51816 );
not \U$40209 ( \51818 , \51766 );
buf \U$40210 ( \51819 , \51818 );
_HMUX g16672 ( \51820_nG16672 , RIe38c4b0_5571 , \51819 , \51775 );
buf \U$40211 ( \51821 , RIe38c4b0_5571);
buf g16676( \51822_nG16676 , \51821 );
_HMUX g16679 ( \51823_nG16679 , \51820_nG16672 , \51822_nG16676 , \51786 );
_HMUX g1667c ( \51824_nG1667c , \51823_nG16679 , 1'b1 , \51789 );
_HMUX g1667e ( \51825_nG1667e , \51824_nG1667c , 1'b0 , \51791 );
buf \U$40216 ( \51826 , \51825_nG1667e );
and \U$40217 ( \51827 , \51817 , \51826 );
xnor \U$40218 ( \51828 , \51810 , \51799 );
and \U$40219 ( \51829 , \51827 , \51828 );
or \U$40220 ( \51830 , \51811 , \51829 );
xnor \U$40221 ( \51831 , \51793 , \51762 );
and \U$40222 ( \51832 , \51830 , \51831 );
or \U$40223 ( \51833 , \51794 , \51832 );
buf \U$40224 ( \51834 , \51833 );
and \U$40225 ( \51835 , \51749 , \51834 );
not \U$40227 ( \51836 , \51623_nG16709 );
or \U$40228 ( \51837 , \51836 , \51708 );
and \U$40229 ( \51838 , \51749 , \51837 );
_HMUX g1670d ( \51839_nG1670d , \51835 , 1'b1 , \51838 );
buf \U$40230 ( \51840 , \51839_nG1670d );
_DC g18bca_GF_IsGateDCbyConstraint ( \51841_nG18bca , \51840 , \42503 );
buf \U$40231 ( \51842 , \51841_nG18bca );
buf \U$40232 ( \51843 , \51716_nG165f2 );
_DC g18e17_GF_IsGateDCbyConstraint ( \51844_nG18e17 , \51843 , \42503 );
buf \U$40233 ( \51845 , \51844_nG18e17 );
buf \U$40234 ( \51846 , \51730_nG165ff );
_DC g18e18_GF_IsGateDCbyConstraint ( \51847_nG18e18 , \51846 , \42503 );
buf \U$40235 ( \51848 , \51847_nG18e18 );
buf \U$40236 ( \51849 , \51746_nG1660e );
_DC g18e19_GF_IsGateDCbyConstraint ( \51850_nG18e19 , \51849 , \42503 );
buf \U$40237 ( \51851 , \51850_nG18e19 );
buf \U$40238 ( \51852 , RIb87eb00_69);
buf \U$40239 ( \51853 , RIe667bb0_6885);
buf \U$40240 ( \51854 , RIe667f70_6886);
nor \U$40241 ( \51855 , \51853 , \51854 );
_HMUX g164b7 ( \51856_nG164b7 , RIe04cad8_4898 , \51852 , \51855 );
and \U$40242 ( \51857 , \47160 , \42387 , RIe546098_6850, RIe545dc8_6851, \42389 );
buf \U$40243 ( \51858 , \51857 );
buf \U$40244 ( \51859 , \51858 );
buf \U$40245 ( \51860 , \42587 );
buf \U$40246 ( \51861 , \51860 );
and \U$40247 ( \51862 , \51859 , \51861 );
_HMUX g164b8 ( \51863_nG164b8 , RIe04cad8_4898 , \51856_nG164b7 , \51862 );
buf \U$40248 ( \51864 , RIb7c5980_237);
buf \U$40249 ( \51865 , RIeab7058_6894);
buf \U$40250 ( \51866 , RIea91768_6889);
nor \U$40251 ( \51867 , \51865 , \51866 );
_HMUX g164ba ( \51868_nG164ba , RIe04cad8_4898 , \51864 , \51867 );
and \U$40252 ( \51869 , \44707 , \42170 , \42218_nGbc1c , \42267_nGbc4c , \42316 );
buf \U$40253 ( \51870 , \51869 );
buf \U$40254 ( \51871 , \51870 );
buf \U$40255 ( \51872 , RIb79b518_270);
buf \U$40256 ( \51873 , \51872 );
and \U$40257 ( \51874 , \51871 , \51873 );
_HMUX g164bb ( \51875_nG164bb , \51863_nG164b8 , \51868_nG164ba , \51874 );
buf \U$40258 ( \51876 , \51875_nG164bb );
_DC g18b07_GF_IsGateDCbyConstraint ( \51877_nG18b07 , \51876 , \42503 );
buf \U$40259 ( \51878 , \51877_nG18b07 );
buf \U$40260 ( \51879 , RIb87eb78_68);
_HMUX g164bc ( \51880_nG164bc , RIe04b980_4899 , \51879 , \51855 );
_HMUX g164bd ( \51881_nG164bd , RIe04b980_4899 , \51880_nG164bc , \51862 );
buf \U$40261 ( \51882 , RIb7c59f8_236);
_HMUX g164be ( \51883_nG164be , RIe04b980_4899 , \51882 , \51867 );
_HMUX g164bf ( \51884_nG164bf , \51881_nG164bd , \51883_nG164be , \51874 );
buf \U$40262 ( \51885 , \51884_nG164bf );
_DC g18b1d_GF_IsGateDCbyConstraint ( \51886_nG18b1d , \51885 , \42503 );
buf \U$40263 ( \51887 , \51886_nG18b1d );
buf \U$40264 ( \51888 , RIb87ebf0_67);
_HMUX g164c0 ( \51889_nG164c0 , RIe04a378_4900 , \51888 , \51855 );
_HMUX g164c1 ( \51890_nG164c1 , RIe04a378_4900 , \51889_nG164c0 , \51862 );
buf \U$40265 ( \51891 , RIb7c5a70_235);
_HMUX g164c2 ( \51892_nG164c2 , RIe04a378_4900 , \51891 , \51867 );
_HMUX g164c3 ( \51893_nG164c3 , \51890_nG164c1 , \51892_nG164c2 , \51874 );
buf \U$40266 ( \51894 , \51893_nG164c3 );
_DC g18b33_GF_IsGateDCbyConstraint ( \51895_nG18b33 , \51894 , \42503 );
buf \U$40267 ( \51896 , \51895_nG18b33 );
buf \U$40268 ( \51897 , RIb882ca0_66);
_HMUX g164c4 ( \51898_nG164c4 , RIe049220_4901 , \51897 , \51855 );
_HMUX g164c5 ( \51899_nG164c5 , RIe049220_4901 , \51898_nG164c4 , \51862 );
buf \U$40269 ( \51900 , RIb7cade0_234);
_HMUX g164c6 ( \51901_nG164c6 , RIe049220_4901 , \51900 , \51867 );
_HMUX g164c7 ( \51902_nG164c7 , \51899_nG164c5 , \51901_nG164c6 , \51874 );
buf \U$40270 ( \51903 , \51902_nG164c7 );
_DC g18b49_GF_IsGateDCbyConstraint ( \51904_nG18b49 , \51903 , \42503 );
buf \U$40271 ( \51905 , \51904_nG18b49 );
buf \U$40272 ( \51906 , RIb885310_65);
_HMUX g164c8 ( \51907_nG164c8 , RIe047c18_4902 , \51906 , \51855 );
_HMUX g164c9 ( \51908_nG164c9 , RIe047c18_4902 , \51907_nG164c8 , \51862 );
buf \U$40273 ( \51909 , RIb7cae58_233);
_HMUX g164ca ( \51910_nG164ca , RIe047c18_4902 , \51909 , \51867 );
_HMUX g164cb ( \51911_nG164cb , \51908_nG164c9 , \51910_nG164ca , \51874 );
buf \U$40274 ( \51912 , \51911_nG164cb );
_DC g18b5f_GF_IsGateDCbyConstraint ( \51913_nG18b5f , \51912 , \42503 );
buf \U$40275 ( \51914 , \51913_nG18b5f );
buf \U$40276 ( \51915 , RIb885388_64);
_HMUX g164cc ( \51916_nG164cc , RIe046ac0_4903 , \51915 , \51855 );
_HMUX g164cd ( \51917_nG164cd , RIe046ac0_4903 , \51916_nG164cc , \51862 );
buf \U$40277 ( \51918 , RIb7caed0_232);
_HMUX g164ce ( \51919_nG164ce , RIe046ac0_4903 , \51918 , \51867 );
_HMUX g164cf ( \51920_nG164cf , \51917_nG164cd , \51919_nG164ce , \51874 );
buf \U$40278 ( \51921 , \51920_nG164cf );
_DC g18b75_GF_IsGateDCbyConstraint ( \51922_nG18b75 , \51921 , \42503 );
buf \U$40279 ( \51923 , \51922_nG18b75 );
buf \U$40280 ( \51924 , RIb885400_63);
_HMUX g164d0 ( \51925_nG164d0 , RIe045968_4904 , \51924 , \51855 );
_HMUX g164d1 ( \51926_nG164d1 , RIe045968_4904 , \51925_nG164d0 , \51862 );
buf \U$40281 ( \51927 , RIb7caf48_231);
_HMUX g164d2 ( \51928_nG164d2 , RIe045968_4904 , \51927 , \51867 );
_HMUX g164d3 ( \51929_nG164d3 , \51926_nG164d1 , \51928_nG164d2 , \51874 );
buf \U$40282 ( \51930 , \51929_nG164d3 );
_DC g18b81_GF_IsGateDCbyConstraint ( \51931_nG18b81 , \51930 , \42503 );
buf \U$40283 ( \51932 , \51931_nG18b81 );
buf \U$40284 ( \51933 , RIb885478_62);
_HMUX g164d4 ( \51934_nG164d4 , RIe044360_4905 , \51933 , \51855 );
_HMUX g164d5 ( \51935_nG164d5 , RIe044360_4905 , \51934_nG164d4 , \51862 );
buf \U$40285 ( \51936 , RIb7cafc0_230);
_HMUX g164d6 ( \51937_nG164d6 , RIe044360_4905 , \51936 , \51867 );
_HMUX g164d7 ( \51938_nG164d7 , \51935_nG164d5 , \51937_nG164d6 , \51874 );
buf \U$40286 ( \51939 , \51938_nG164d7 );
_DC g18b83_GF_IsGateDCbyConstraint ( \51940_nG18b83 , \51939 , \42503 );
buf \U$40287 ( \51941 , \51940_nG18b83 );
buf \U$40288 ( \51942 , RIb8854f0_61);
_HMUX g164d8 ( \51943_nG164d8 , RIe043208_4906 , \51942 , \51855 );
_HMUX g164d9 ( \51944_nG164d9 , RIe043208_4906 , \51943_nG164d8 , \51862 );
buf \U$40289 ( \51945 , RIb7cb038_229);
_HMUX g164da ( \51946_nG164da , RIe043208_4906 , \51945 , \51867 );
_HMUX g164db ( \51947_nG164db , \51944_nG164d9 , \51946_nG164da , \51874 );
buf \U$40290 ( \51948 , \51947_nG164db );
_DC g18b85_GF_IsGateDCbyConstraint ( \51949_nG18b85 , \51948 , \42503 );
buf \U$40291 ( \51950 , \51949_nG18b85 );
buf \U$40292 ( \51951 , RIb885568_60);
_HMUX g164dc ( \51952_nG164dc , RIe041c00_4907 , \51951 , \51855 );
_HMUX g164dd ( \51953_nG164dd , RIe041c00_4907 , \51952_nG164dc , \51862 );
buf \U$40293 ( \51954 , RIb7cb0b0_228);
_HMUX g164de ( \51955_nG164de , RIe041c00_4907 , \51954 , \51867 );
_HMUX g164df ( \51956_nG164df , \51953_nG164dd , \51955_nG164de , \51874 );
buf \U$40294 ( \51957 , \51956_nG164df );
_DC g18b09_GF_IsGateDCbyConstraint ( \51958_nG18b09 , \51957 , \42503 );
buf \U$40295 ( \51959 , \51958_nG18b09 );
buf \U$40296 ( \51960 , RIb8855e0_59);
_HMUX g164e0 ( \51961_nG164e0 , RIe040aa8_4908 , \51960 , \51855 );
_HMUX g164e1 ( \51962_nG164e1 , RIe040aa8_4908 , \51961_nG164e0 , \51862 );
buf \U$40297 ( \51963 , RIb7cb128_227);
_HMUX g164e2 ( \51964_nG164e2 , RIe040aa8_4908 , \51963 , \51867 );
_HMUX g164e3 ( \51965_nG164e3 , \51962_nG164e1 , \51964_nG164e2 , \51874 );
buf \U$40298 ( \51966 , \51965_nG164e3 );
_DC g18b0b_GF_IsGateDCbyConstraint ( \51967_nG18b0b , \51966 , \42503 );
buf \U$40299 ( \51968 , \51967_nG18b0b );
buf \U$40300 ( \51969 , RIb885658_58);
_HMUX g164e4 ( \51970_nG164e4 , RIe03f4a0_4909 , \51969 , \51855 );
_HMUX g164e5 ( \51971_nG164e5 , RIe03f4a0_4909 , \51970_nG164e4 , \51862 );
buf \U$40301 ( \51972 , RIb7d00d8_226);
_HMUX g164e6 ( \51973_nG164e6 , RIe03f4a0_4909 , \51972 , \51867 );
_HMUX g164e7 ( \51974_nG164e7 , \51971_nG164e5 , \51973_nG164e6 , \51874 );
buf \U$40302 ( \51975 , \51974_nG164e7 );
_DC g18b0d_GF_IsGateDCbyConstraint ( \51976_nG18b0d , \51975 , \42503 );
buf \U$40303 ( \51977 , \51976_nG18b0d );
buf \U$40304 ( \51978 , RIb8856d0_57);
_HMUX g164e8 ( \51979_nG164e8 , RIe03e348_4910 , \51978 , \51855 );
_HMUX g164e9 ( \51980_nG164e9 , RIe03e348_4910 , \51979_nG164e8 , \51862 );
buf \U$40305 ( \51981 , RIb8263d8_225);
_HMUX g164ea ( \51982_nG164ea , RIe03e348_4910 , \51981 , \51867 );
_HMUX g164eb ( \51983_nG164eb , \51980_nG164e9 , \51982_nG164ea , \51874 );
buf \U$40306 ( \51984 , \51983_nG164eb );
_DC g18b0f_GF_IsGateDCbyConstraint ( \51985_nG18b0f , \51984 , \42503 );
buf \U$40307 ( \51986 , \51985_nG18b0f );
buf \U$40308 ( \51987 , RIb885748_56);
_HMUX g164ec ( \51988_nG164ec , RIe03d1f0_4911 , \51987 , \51855 );
_HMUX g164ed ( \51989_nG164ed , RIe03d1f0_4911 , \51988_nG164ec , \51862 );
buf \U$40309 ( \51990 , RIb826e28_224);
_HMUX g164ee ( \51991_nG164ee , RIe03d1f0_4911 , \51990 , \51867 );
_HMUX g164ef ( \51992_nG164ef , \51989_nG164ed , \51991_nG164ee , \51874 );
buf \U$40310 ( \51993 , \51992_nG164ef );
_DC g18b11_GF_IsGateDCbyConstraint ( \51994_nG18b11 , \51993 , \42503 );
buf \U$40311 ( \51995 , \51994_nG18b11 );
buf \U$40312 ( \51996 , RIb8857c0_55);
_HMUX g164f0 ( \51997_nG164f0 , RIde08bc0_4912 , \51996 , \51855 );
_HMUX g164f1 ( \51998_nG164f1 , RIde08bc0_4912 , \51997_nG164f0 , \51862 );
buf \U$40313 ( \51999 , RIb826ea0_223);
_HMUX g164f2 ( \52000_nG164f2 , RIde08bc0_4912 , \51999 , \51867 );
_HMUX g164f3 ( \52001_nG164f3 , \51998_nG164f1 , \52000_nG164f2 , \51874 );
buf \U$40314 ( \52002 , \52001_nG164f3 );
_DC g18b13_GF_IsGateDCbyConstraint ( \52003_nG18b13 , \52002 , \42503 );
buf \U$40315 ( \52004 , \52003_nG18b13 );
buf \U$40316 ( \52005 , RIb885838_54);
_HMUX g164f4 ( \52006_nG164f4 , RIde0d030_4913 , \52005 , \51855 );
_HMUX g164f5 ( \52007_nG164f5 , RIde0d030_4913 , \52006_nG164f4 , \51862 );
buf \U$40317 ( \52008 , RIb826f18_222);
_HMUX g164f6 ( \52009_nG164f6 , RIde0d030_4913 , \52008 , \51867 );
_HMUX g164f7 ( \52010_nG164f7 , \52007_nG164f5 , \52009_nG164f6 , \51874 );
buf \U$40318 ( \52011 , \52010_nG164f7 );
_DC g18b15_GF_IsGateDCbyConstraint ( \52012_nG18b15 , \52011 , \42503 );
buf \U$40319 ( \52013 , \52012_nG18b15 );
buf \U$40320 ( \52014 , RIb8858b0_53);
_HMUX g164f8 ( \52015_nG164f8 , RIde131b0_4914 , \52014 , \51855 );
_HMUX g164f9 ( \52016_nG164f9 , RIde131b0_4914 , \52015_nG164f8 , \51862 );
buf \U$40321 ( \52017 , RIb826f90_221);
_HMUX g164fa ( \52018_nG164fa , RIde131b0_4914 , \52017 , \51867 );
_HMUX g164fb ( \52019_nG164fb , \52016_nG164f9 , \52018_nG164fa , \51874 );
buf \U$40322 ( \52020 , \52019_nG164fb );
_DC g18b17_GF_IsGateDCbyConstraint ( \52021_nG18b17 , \52020 , \42503 );
buf \U$40323 ( \52022 , \52021_nG18b17 );
buf \U$40324 ( \52023 , RIb885928_52);
_HMUX g164fc ( \52024_nG164fc , RIde17968_4915 , \52023 , \51855 );
_HMUX g164fd ( \52025_nG164fd , RIde17968_4915 , \52024_nG164fc , \51862 );
buf \U$40325 ( \52026 , RIb8293a8_220);
_HMUX g164fe ( \52027_nG164fe , RIde17968_4915 , \52026 , \51867 );
_HMUX g164ff ( \52028_nG164ff , \52025_nG164fd , \52027_nG164fe , \51874 );
buf \U$40326 ( \52029 , \52028_nG164ff );
_DC g18b19_GF_IsGateDCbyConstraint ( \52030_nG18b19 , \52029 , \42503 );
buf \U$40327 ( \52031 , \52030_nG18b19 );
buf \U$40328 ( \52032 , RIb8859a0_51);
_HMUX g16500 ( \52033_nG16500 , RIde1f528_4916 , \52032 , \51855 );
_HMUX g16501 ( \52034_nG16501 , RIde1f528_4916 , \52033_nG16500 , \51862 );
buf \U$40329 ( \52035 , RIb829420_219);
_HMUX g16502 ( \52036_nG16502 , RIde1f528_4916 , \52035 , \51867 );
_HMUX g16503 ( \52037_nG16503 , \52034_nG16501 , \52036_nG16502 , \51874 );
buf \U$40330 ( \52038 , \52037_nG16503 );
_DC g18b1b_GF_IsGateDCbyConstraint ( \52039_nG18b1b , \52038 , \42503 );
buf \U$40331 ( \52040 , \52039_nG18b1b );
buf \U$40332 ( \52041 , RIb885a18_50);
_HMUX g16504 ( \52042_nG16504 , RIde24e38_4917 , \52041 , \51855 );
_HMUX g16505 ( \52043_nG16505 , RIde24e38_4917 , \52042_nG16504 , \51862 );
buf \U$40333 ( \52044 , RIb829498_218);
_HMUX g16506 ( \52045_nG16506 , RIde24e38_4917 , \52044 , \51867 );
_HMUX g16507 ( \52046_nG16507 , \52043_nG16505 , \52045_nG16506 , \51874 );
buf \U$40334 ( \52047 , \52046_nG16507 );
_DC g18b1f_GF_IsGateDCbyConstraint ( \52048_nG18b1f , \52047 , \42503 );
buf \U$40335 ( \52049 , \52048_nG18b1f );
buf \U$40336 ( \52050 , RIb885a90_49);
_HMUX g16508 ( \52051_nG16508 , RIde29ed8_4918 , \52050 , \51855 );
_HMUX g16509 ( \52052_nG16509 , RIde29ed8_4918 , \52051_nG16508 , \51862 );
buf \U$40337 ( \52053 , RIb829510_217);
_HMUX g1650a ( \52054_nG1650a , RIde29ed8_4918 , \52053 , \51867 );
_HMUX g1650b ( \52055_nG1650b , \52052_nG16509 , \52054_nG1650a , \51874 );
buf \U$40338 ( \52056 , \52055_nG1650b );
_DC g18b21_GF_IsGateDCbyConstraint ( \52057_nG18b21 , \52056 , \42503 );
buf \U$40339 ( \52058 , \52057_nG18b21 );
buf \U$40340 ( \52059 , RIb885b08_48);
_HMUX g1650c ( \52060_nG1650c , RIde31390_4919 , \52059 , \51855 );
_HMUX g1650d ( \52061_nG1650d , RIde31390_4919 , \52060_nG1650c , \51862 );
buf \U$40341 ( \52062 , RIb829588_216);
_HMUX g1650e ( \52063_nG1650e , RIde31390_4919 , \52062 , \51867 );
_HMUX g1650f ( \52064_nG1650f , \52061_nG1650d , \52063_nG1650e , \51874 );
buf \U$40342 ( \52065 , \52064_nG1650f );
_DC g18b23_GF_IsGateDCbyConstraint ( \52066_nG18b23 , \52065 , \42503 );
buf \U$40343 ( \52067 , \52066_nG18b23 );
buf \U$40344 ( \52068 , RIb885b80_47);
_HMUX g16510 ( \52069_nG16510 , RIde36e08_4920 , \52068 , \51855 );
_HMUX g16511 ( \52070_nG16511 , RIde36e08_4920 , \52069_nG16510 , \51862 );
buf \U$40345 ( \52071 , RIb829600_215);
_HMUX g16512 ( \52072_nG16512 , RIde36e08_4920 , \52071 , \51867 );
_HMUX g16513 ( \52073_nG16513 , \52070_nG16511 , \52072_nG16512 , \51874 );
buf \U$40346 ( \52074 , \52073_nG16513 );
_DC g18b25_GF_IsGateDCbyConstraint ( \52075_nG18b25 , \52074 , \42503 );
buf \U$40347 ( \52076 , \52075_nG18b25 );
buf \U$40348 ( \52077 , RIb885bf8_46);
_HMUX g16514 ( \52078_nG16514 , RIde3efe0_4921 , \52077 , \51855 );
_HMUX g16515 ( \52079_nG16515 , RIde3efe0_4921 , \52078_nG16514 , \51862 );
buf \U$40349 ( \52080 , RIb829678_214);
_HMUX g16516 ( \52081_nG16516 , RIde3efe0_4921 , \52080 , \51867 );
_HMUX g16517 ( \52082_nG16517 , \52079_nG16515 , \52081_nG16516 , \51874 );
buf \U$40350 ( \52083 , \52082_nG16517 );
_DC g18b27_GF_IsGateDCbyConstraint ( \52084_nG18b27 , \52083 , \42503 );
buf \U$40351 ( \52085 , \52084_nG18b27 );
buf \U$40352 ( \52086 , RIb885c70_45);
_HMUX g16518 ( \52087_nG16518 , RIde45070_4922 , \52086 , \51855 );
_HMUX g16519 ( \52088_nG16519 , RIde45070_4922 , \52087_nG16518 , \51862 );
buf \U$40353 ( \52089 , RIb8296f0_213);
_HMUX g1651a ( \52090_nG1651a , RIde45070_4922 , \52089 , \51867 );
_HMUX g1651b ( \52091_nG1651b , \52088_nG16519 , \52090_nG1651a , \51874 );
buf \U$40354 ( \52092 , \52091_nG1651b );
_DC g18b29_GF_IsGateDCbyConstraint ( \52093_nG18b29 , \52092 , \42503 );
buf \U$40355 ( \52094 , \52093_nG18b29 );
buf \U$40356 ( \52095 , RIb885ce8_44);
_HMUX g1651c ( \52096_nG1651c , RIde4c9d8_4923 , \52095 , \51855 );
_HMUX g1651d ( \52097_nG1651d , RIde4c9d8_4923 , \52096_nG1651c , \51862 );
buf \U$40357 ( \52098 , RIb82dae8_212);
_HMUX g1651e ( \52099_nG1651e , RIde4c9d8_4923 , \52098 , \51867 );
_HMUX g1651f ( \52100_nG1651f , \52097_nG1651d , \52099_nG1651e , \51874 );
buf \U$40358 ( \52101 , \52100_nG1651f );
_DC g18b2b_GF_IsGateDCbyConstraint ( \52102_nG18b2b , \52101 , \42503 );
buf \U$40359 ( \52103 , \52102_nG18b2b );
buf \U$40360 ( \52104 , RIb885d60_43);
_HMUX g16520 ( \52105_nG16520 , RIde51b68_4924 , \52104 , \51855 );
_HMUX g16521 ( \52106_nG16521 , RIde51b68_4924 , \52105_nG16520 , \51862 );
buf \U$40361 ( \52107 , RIb82db60_211);
_HMUX g16522 ( \52108_nG16522 , RIde51b68_4924 , \52107 , \51867 );
_HMUX g16523 ( \52109_nG16523 , \52106_nG16521 , \52108_nG16522 , \51874 );
buf \U$40362 ( \52110 , \52109_nG16523 );
_DC g18b2d_GF_IsGateDCbyConstraint ( \52111_nG18b2d , \52110 , \42503 );
buf \U$40363 ( \52112 , \52111_nG18b2d );
buf \U$40364 ( \52113 , RIb885dd8_42);
_HMUX g16524 ( \52114_nG16524 , RIde553a8_4925 , \52113 , \51855 );
_HMUX g16525 ( \52115_nG16525 , RIde553a8_4925 , \52114_nG16524 , \51862 );
buf \U$40365 ( \52116 , RIb82dbd8_210);
_HMUX g16526 ( \52117_nG16526 , RIde553a8_4925 , \52116 , \51867 );
_HMUX g16527 ( \52118_nG16527 , \52115_nG16525 , \52117_nG16526 , \51874 );
buf \U$40366 ( \52119 , \52118_nG16527 );
_DC g18b2f_GF_IsGateDCbyConstraint ( \52120_nG18b2f , \52119 , \42503 );
buf \U$40367 ( \52121 , \52120_nG18b2f );
buf \U$40368 ( \52122 , RIb885e50_41);
_HMUX g16528 ( \52123_nG16528 , RIde59c50_4926 , \52122 , \51855 );
_HMUX g16529 ( \52124_nG16529 , RIde59c50_4926 , \52123_nG16528 , \51862 );
buf \U$40369 ( \52125 , RIb82dc50_209);
_HMUX g1652a ( \52126_nG1652a , RIde59c50_4926 , \52125 , \51867 );
_HMUX g1652b ( \52127_nG1652b , \52124_nG16529 , \52126_nG1652a , \51874 );
buf \U$40370 ( \52128 , \52127_nG1652b );
_DC g18b31_GF_IsGateDCbyConstraint ( \52129_nG18b31 , \52128 , \42503 );
buf \U$40371 ( \52130 , \52129_nG18b31 );
buf \U$40372 ( \52131 , RIb885ec8_40);
_HMUX g1652c ( \52132_nG1652c , RIde5e390_4927 , \52131 , \51855 );
_HMUX g1652d ( \52133_nG1652d , RIde5e390_4927 , \52132_nG1652c , \51862 );
buf \U$40373 ( \52134 , RIb82dcc8_208);
_HMUX g1652e ( \52135_nG1652e , RIde5e390_4927 , \52134 , \51867 );
_HMUX g1652f ( \52136_nG1652f , \52133_nG1652d , \52135_nG1652e , \51874 );
buf \U$40374 ( \52137 , \52136_nG1652f );
_DC g18b35_GF_IsGateDCbyConstraint ( \52138_nG18b35 , \52137 , \42503 );
buf \U$40375 ( \52139 , \52138_nG18b35 );
buf \U$40376 ( \52140 , RIb885f40_39);
_HMUX g16530 ( \52141_nG16530 , RIde65668_4928 , \52140 , \51855 );
_HMUX g16531 ( \52142_nG16531 , RIde65668_4928 , \52141_nG16530 , \51862 );
buf \U$40377 ( \52143 , RIb82dd40_207);
_HMUX g16532 ( \52144_nG16532 , RIde65668_4928 , \52143 , \51867 );
_HMUX g16533 ( \52145_nG16533 , \52142_nG16531 , \52144_nG16532 , \51874 );
buf \U$40378 ( \52146 , \52145_nG16533 );
_DC g18b37_GF_IsGateDCbyConstraint ( \52147_nG18b37 , \52146 , \42503 );
buf \U$40379 ( \52148 , \52147_nG18b37 );
buf \U$40380 ( \52149 , RIb885fb8_38);
_HMUX g16534 ( \52150_nG16534 , RIde6a4b0_4929 , \52149 , \51855 );
_HMUX g16535 ( \52151_nG16535 , RIde6a4b0_4929 , \52150_nG16534 , \51862 );
buf \U$40381 ( \52152 , RIb82ddb8_206);
_HMUX g16536 ( \52153_nG16536 , RIde6a4b0_4929 , \52152 , \51867 );
_HMUX g16537 ( \52154_nG16537 , \52151_nG16535 , \52153_nG16536 , \51874 );
buf \U$40382 ( \52155 , \52154_nG16537 );
_DC g18b39_GF_IsGateDCbyConstraint ( \52156_nG18b39 , \52155 , \42503 );
buf \U$40383 ( \52157 , \52156_nG18b39 );
buf \U$40384 ( \52158 , RIb886030_37);
_HMUX g16538 ( \52159_nG16538 , RIde6f820_4930 , \52158 , \51855 );
_HMUX g16539 ( \52160_nG16539 , RIde6f820_4930 , \52159_nG16538 , \51862 );
buf \U$40385 ( \52161 , RIb82de30_205);
_HMUX g1653a ( \52162_nG1653a , RIde6f820_4930 , \52161 , \51867 );
_HMUX g1653b ( \52163_nG1653b , \52160_nG16539 , \52162_nG1653a , \51874 );
buf \U$40386 ( \52164 , \52163_nG1653b );
_DC g18b3b_GF_IsGateDCbyConstraint ( \52165_nG18b3b , \52164 , \42503 );
buf \U$40387 ( \52166 , \52165_nG18b3b );
buf \U$40388 ( \52167 , RIb8860a8_36);
_HMUX g1653c ( \52168_nG1653c , RIdf73710_4931 , \52167 , \51855 );
_HMUX g1653d ( \52169_nG1653d , RIdf73710_4931 , \52168_nG1653c , \51862 );
buf \U$40389 ( \52170 , RIb832228_204);
_HMUX g1653e ( \52171_nG1653e , RIdf73710_4931 , \52170 , \51867 );
_HMUX g1653f ( \52172_nG1653f , \52169_nG1653d , \52171_nG1653e , \51874 );
buf \U$40390 ( \52173 , \52172_nG1653f );
_DC g18b3d_GF_IsGateDCbyConstraint ( \52174_nG18b3d , \52173 , \42503 );
buf \U$40391 ( \52175 , \52174_nG18b3d );
buf \U$40392 ( \52176 , RIb886120_35);
_HMUX g16540 ( \52177_nG16540 , RIdc38040_4932 , \52176 , \51855 );
_HMUX g16541 ( \52178_nG16541 , RIdc38040_4932 , \52177_nG16540 , \51862 );
buf \U$40393 ( \52179 , RIb8322a0_203);
_HMUX g16542 ( \52180_nG16542 , RIdc38040_4932 , \52179 , \51867 );
_HMUX g16543 ( \52181_nG16543 , \52178_nG16541 , \52180_nG16542 , \51874 );
buf \U$40394 ( \52182 , \52181_nG16543 );
_DC g18b3f_GF_IsGateDCbyConstraint ( \52183_nG18b3f , \52182 , \42503 );
buf \U$40395 ( \52184 , \52183_nG18b3f );
buf \U$40396 ( \52185 , RIb886198_34);
_HMUX g16544 ( \52186_nG16544 , RIdc32b68_4933 , \52185 , \51855 );
_HMUX g16545 ( \52187_nG16545 , RIdc32b68_4933 , \52186_nG16544 , \51862 );
buf \U$40397 ( \52188 , RIb832318_202);
_HMUX g16546 ( \52189_nG16546 , RIdc32b68_4933 , \52188 , \51867 );
_HMUX g16547 ( \52190_nG16547 , \52187_nG16545 , \52189_nG16546 , \51874 );
buf \U$40398 ( \52191 , \52190_nG16547 );
_DC g18b41_GF_IsGateDCbyConstraint ( \52192_nG18b41 , \52191 , \42503 );
buf \U$40399 ( \52193 , \52192_nG18b41 );
buf \U$40400 ( \52194 , RIb886210_33);
_HMUX g16548 ( \52195_nG16548 , RIdc2ee78_4934 , \52194 , \51855 );
_HMUX g16549 ( \52196_nG16549 , RIdc2ee78_4934 , \52195_nG16548 , \51862 );
buf \U$40401 ( \52197 , RIb832390_201);
_HMUX g1654a ( \52198_nG1654a , RIdc2ee78_4934 , \52197 , \51867 );
_HMUX g1654b ( \52199_nG1654b , \52196_nG16549 , \52198_nG1654a , \51874 );
buf \U$40402 ( \52200 , \52199_nG1654b );
_DC g18b43_GF_IsGateDCbyConstraint ( \52201_nG18b43 , \52200 , \42503 );
buf \U$40403 ( \52202 , \52201_nG18b43 );
buf \U$40404 ( \52203 , RIb886288_32);
_HMUX g1654c ( \52204_nG1654c , RIdc29bf8_4935 , \52203 , \51855 );
_HMUX g1654d ( \52205_nG1654d , RIdc29bf8_4935 , \52204_nG1654c , \51862 );
buf \U$40405 ( \52206 , RIb832408_200);
_HMUX g1654e ( \52207_nG1654e , RIdc29bf8_4935 , \52206 , \51867 );
_HMUX g1654f ( \52208_nG1654f , \52205_nG1654d , \52207_nG1654e , \51874 );
buf \U$40406 ( \52209 , \52208_nG1654f );
_DC g18b45_GF_IsGateDCbyConstraint ( \52210_nG18b45 , \52209 , \42503 );
buf \U$40407 ( \52211 , \52210_nG18b45 );
buf \U$40408 ( \52212 , RIb886300_31);
_HMUX g16550 ( \52213_nG16550 , RIddf1628_4936 , \52212 , \51855 );
_HMUX g16551 ( \52214_nG16551 , RIddf1628_4936 , \52213_nG16550 , \51862 );
buf \U$40409 ( \52215 , RIb832480_199);
_HMUX g16552 ( \52216_nG16552 , RIddf1628_4936 , \52215 , \51867 );
_HMUX g16553 ( \52217_nG16553 , \52214_nG16551 , \52216_nG16552 , \51874 );
buf \U$40410 ( \52218 , \52217_nG16553 );
_DC g18b47_GF_IsGateDCbyConstraint ( \52219_nG18b47 , \52218 , \42503 );
buf \U$40411 ( \52220 , \52219_nG18b47 );
buf \U$40412 ( \52221 , RIb886378_30);
_HMUX g16554 ( \52222_nG16554 , RIddee388_4937 , \52221 , \51855 );
_HMUX g16555 ( \52223_nG16555 , RIddee388_4937 , \52222_nG16554 , \51862 );
buf \U$40413 ( \52224 , RIb8324f8_198);
_HMUX g16556 ( \52225_nG16556 , RIddee388_4937 , \52224 , \51867 );
_HMUX g16557 ( \52226_nG16557 , \52223_nG16555 , \52225_nG16556 , \51874 );
buf \U$40414 ( \52227 , \52226_nG16557 );
_DC g18b4b_GF_IsGateDCbyConstraint ( \52228_nG18b4b , \52227 , \42503 );
buf \U$40415 ( \52229 , \52228_nG18b4b );
buf \U$40416 ( \52230 , RIb8863f0_29);
_HMUX g16558 ( \52231_nG16558 , RIddeaa58_4938 , \52230 , \51855 );
_HMUX g16559 ( \52232_nG16559 , RIddeaa58_4938 , \52231_nG16558 , \51862 );
buf \U$40417 ( \52233 , RIb832570_197);
_HMUX g1655a ( \52234_nG1655a , RIddeaa58_4938 , \52233 , \51867 );
_HMUX g1655b ( \52235_nG1655b , \52232_nG16559 , \52234_nG1655a , \51874 );
buf \U$40418 ( \52236 , \52235_nG1655b );
_DC g18b4d_GF_IsGateDCbyConstraint ( \52237_nG18b4d , \52236 , \42503 );
buf \U$40419 ( \52238 , \52237_nG18b4d );
buf \U$40420 ( \52239 , RIb886468_28);
_HMUX g1655c ( \52240_nG1655c , RIdde7a88_4939 , \52239 , \51855 );
_HMUX g1655d ( \52241_nG1655d , RIdde7a88_4939 , \52240_nG1655c , \51862 );
buf \U$40421 ( \52242 , RIb8383a8_196);
_HMUX g1655e ( \52243_nG1655e , RIdde7a88_4939 , \52242 , \51867 );
_HMUX g1655f ( \52244_nG1655f , \52241_nG1655d , \52243_nG1655e , \51874 );
buf \U$40422 ( \52245 , \52244_nG1655f );
_DC g18b4f_GF_IsGateDCbyConstraint ( \52246_nG18b4f , \52245 , \42503 );
buf \U$40423 ( \52247 , \52246_nG18b4f );
buf \U$40424 ( \52248 , RIb8864e0_27);
_HMUX g16560 ( \52249_nG16560 , RIdde35a0_4940 , \52248 , \51855 );
_HMUX g16561 ( \52250_nG16561 , RIdde35a0_4940 , \52249_nG16560 , \51862 );
buf \U$40425 ( \52251 , RIb838420_195);
_HMUX g16562 ( \52252_nG16562 , RIdde35a0_4940 , \52251 , \51867 );
_HMUX g16563 ( \52253_nG16563 , \52250_nG16561 , \52252_nG16562 , \51874 );
buf \U$40426 ( \52254 , \52253_nG16563 );
_DC g18b51_GF_IsGateDCbyConstraint ( \52255_nG18b51 , \52254 , \42503 );
buf \U$40427 ( \52256 , \52255_nG18b51 );
buf \U$40428 ( \52257 , RIb886558_26);
_HMUX g16564 ( \52258_nG16564 , RIdde0cd8_4941 , \52257 , \51855 );
_HMUX g16565 ( \52259_nG16565 , RIdde0cd8_4941 , \52258_nG16564 , \51862 );
buf \U$40429 ( \52260 , RIb838498_194);
_HMUX g16566 ( \52261_nG16566 , RIdde0cd8_4941 , \52260 , \51867 );
_HMUX g16567 ( \52262_nG16567 , \52259_nG16565 , \52261_nG16566 , \51874 );
buf \U$40430 ( \52263 , \52262_nG16567 );
_DC g18b53_GF_IsGateDCbyConstraint ( \52264_nG18b53 , \52263 , \42503 );
buf \U$40431 ( \52265 , \52264_nG18b53 );
buf \U$40432 ( \52266 , RIb8865d0_25);
_HMUX g16568 ( \52267_nG16568 , RIddddf60_4942 , \52266 , \51855 );
_HMUX g16569 ( \52268_nG16569 , RIddddf60_4942 , \52267_nG16568 , \51862 );
buf \U$40433 ( \52269 , RIb838510_193);
_HMUX g1656a ( \52270_nG1656a , RIddddf60_4942 , \52269 , \51867 );
_HMUX g1656b ( \52271_nG1656b , \52268_nG16569 , \52270_nG1656a , \51874 );
buf \U$40434 ( \52272 , \52271_nG1656b );
_DC g18b55_GF_IsGateDCbyConstraint ( \52273_nG18b55 , \52272 , \42503 );
buf \U$40435 ( \52274 , \52273_nG18b55 );
buf \U$40436 ( \52275 , RIb886648_24);
_HMUX g1656c ( \52276_nG1656c , RIdddb710_4943 , \52275 , \51855 );
_HMUX g1656d ( \52277_nG1656d , RIdddb710_4943 , \52276_nG1656c , \51862 );
buf \U$40437 ( \52278 , RIb838588_192);
_HMUX g1656e ( \52279_nG1656e , RIdddb710_4943 , \52278 , \51867 );
_HMUX g1656f ( \52280_nG1656f , \52277_nG1656d , \52279_nG1656e , \51874 );
buf \U$40438 ( \52281 , \52280_nG1656f );
_DC g18b57_GF_IsGateDCbyConstraint ( \52282_nG18b57 , \52281 , \42503 );
buf \U$40439 ( \52283 , \52282_nG18b57 );
buf \U$40440 ( \52284 , RIb8866c0_23);
_HMUX g16570 ( \52285_nG16570 , RIddd5e78_4944 , \52284 , \51855 );
_HMUX g16571 ( \52286_nG16571 , RIddd5e78_4944 , \52285_nG16570 , \51862 );
buf \U$40441 ( \52287 , RIb838600_191);
_HMUX g16572 ( \52288_nG16572 , RIddd5e78_4944 , \52287 , \51867 );
_HMUX g16573 ( \52289_nG16573 , \52286_nG16571 , \52288_nG16572 , \51874 );
buf \U$40442 ( \52290 , \52289_nG16573 );
_DC g18b59_GF_IsGateDCbyConstraint ( \52291_nG18b59 , \52290 , \42503 );
buf \U$40443 ( \52292 , \52291_nG18b59 );
buf \U$40444 ( \52293 , RIb886738_22);
_HMUX g16574 ( \52294_nG16574 , RIddd2278_4945 , \52293 , \51855 );
_HMUX g16575 ( \52295_nG16575 , RIddd2278_4945 , \52294_nG16574 , \51862 );
buf \U$40445 ( \52296 , RIb838678_190);
_HMUX g16576 ( \52297_nG16576 , RIddd2278_4945 , \52296 , \51867 );
_HMUX g16577 ( \52298_nG16577 , \52295_nG16575 , \52297_nG16576 , \51874 );
buf \U$40446 ( \52299 , \52298_nG16577 );
_DC g18b5b_GF_IsGateDCbyConstraint ( \52300_nG18b5b , \52299 , \42503 );
buf \U$40447 ( \52301 , \52300_nG18b5b );
buf \U$40448 ( \52302 , RIb8867b0_21);
_HMUX g16578 ( \52303_nG16578 , RIddcc080_4946 , \52302 , \51855 );
_HMUX g16579 ( \52304_nG16579 , RIddcc080_4946 , \52303_nG16578 , \51862 );
buf \U$40449 ( \52305 , RIb8386f0_189);
_HMUX g1657a ( \52306_nG1657a , RIddcc080_4946 , \52305 , \51867 );
_HMUX g1657b ( \52307_nG1657b , \52304_nG16579 , \52306_nG1657a , \51874 );
buf \U$40450 ( \52308 , \52307_nG1657b );
_DC g18b5d_GF_IsGateDCbyConstraint ( \52309_nG18b5d , \52308 , \42503 );
buf \U$40451 ( \52310 , \52309_nG18b5d );
buf \U$40452 ( \52311 , RIb886828_20);
_HMUX g1657c ( \52312_nG1657c , RIddc39f8_4947 , \52311 , \51855 );
_HMUX g1657d ( \52313_nG1657d , RIddc39f8_4947 , \52312_nG1657c , \51862 );
buf \U$40453 ( \52314 , RIb838768_188);
_HMUX g1657e ( \52315_nG1657e , RIddc39f8_4947 , \52314 , \51867 );
_HMUX g1657f ( \52316_nG1657f , \52313_nG1657d , \52315_nG1657e , \51874 );
buf \U$40454 ( \52317 , \52316_nG1657f );
_DC g18b61_GF_IsGateDCbyConstraint ( \52318_nG18b61 , \52317 , \42503 );
buf \U$40455 ( \52319 , \52318_nG18b61 );
buf \U$40456 ( \52320 , RIb8868a0_19);
_HMUX g16580 ( \52321_nG16580 , RIddbd8f0_4948 , \52320 , \51855 );
_HMUX g16581 ( \52322_nG16581 , RIddbd8f0_4948 , \52321_nG16580 , \51862 );
buf \U$40457 ( \52323 , RIb8387e0_187);
_HMUX g16582 ( \52324_nG16582 , RIddbd8f0_4948 , \52323 , \51867 );
_HMUX g16583 ( \52325_nG16583 , \52322_nG16581 , \52324_nG16582 , \51874 );
buf \U$40458 ( \52326 , \52325_nG16583 );
_DC g18b63_GF_IsGateDCbyConstraint ( \52327_nG18b63 , \52326 , \42503 );
buf \U$40459 ( \52328 , \52327_nG18b63 );
buf \U$40460 ( \52329 , RIb886918_18);
_HMUX g16584 ( \52330_nG16584 , RIddb5268_4949 , \52329 , \51855 );
_HMUX g16585 ( \52331_nG16585 , RIddb5268_4949 , \52330_nG16584 , \51862 );
buf \U$40461 ( \52332 , RIb838858_186);
_HMUX g16586 ( \52333_nG16586 , RIddb5268_4949 , \52332 , \51867 );
_HMUX g16587 ( \52334_nG16587 , \52331_nG16585 , \52333_nG16586 , \51874 );
buf \U$40462 ( \52335 , \52334_nG16587 );
_DC g18b65_GF_IsGateDCbyConstraint ( \52336_nG18b65 , \52335 , \42503 );
buf \U$40463 ( \52337 , \52336_nG18b65 );
buf \U$40464 ( \52338 , RIb886990_17);
_HMUX g16588 ( \52339_nG16588 , RIddaf160_4950 , \52338 , \51855 );
_HMUX g16589 ( \52340_nG16589 , RIddaf160_4950 , \52339_nG16588 , \51862 );
buf \U$40465 ( \52341 , RIb8388d0_185);
_HMUX g1658a ( \52342_nG1658a , RIddaf160_4950 , \52341 , \51867 );
_HMUX g1658b ( \52343_nG1658b , \52340_nG16589 , \52342_nG1658a , \51874 );
buf \U$40466 ( \52344 , \52343_nG1658b );
_DC g18b67_GF_IsGateDCbyConstraint ( \52345_nG18b67 , \52344 , \42503 );
buf \U$40467 ( \52346 , \52345_nG18b67 );
buf \U$40468 ( \52347 , RIb886a08_16);
_HMUX g1658c ( \52348_nG1658c , RIdb7c228_4951 , \52347 , \51855 );
_HMUX g1658d ( \52349_nG1658d , RIdb7c228_4951 , \52348_nG1658c , \51862 );
buf \U$40469 ( \52350 , RIb838948_184);
_HMUX g1658e ( \52351_nG1658e , RIdb7c228_4951 , \52350 , \51867 );
_HMUX g1658f ( \52352_nG1658f , \52349_nG1658d , \52351_nG1658e , \51874 );
buf \U$40470 ( \52353 , \52352_nG1658f );
_DC g18b69_GF_IsGateDCbyConstraint ( \52354_nG18b69 , \52353 , \42503 );
buf \U$40471 ( \52355 , \52354_nG18b69 );
buf \U$40472 ( \52356 , RIb886a80_15);
_HMUX g16590 ( \52357_nG16590 , RIdb96c40_4952 , \52356 , \51855 );
_HMUX g16591 ( \52358_nG16591 , RIdb96c40_4952 , \52357_nG16590 , \51862 );
buf \U$40473 ( \52359 , RIb8389c0_183);
_HMUX g16592 ( \52360_nG16592 , RIdb96c40_4952 , \52359 , \51867 );
_HMUX g16593 ( \52361_nG16593 , \52358_nG16591 , \52360_nG16592 , \51874 );
buf \U$40474 ( \52362 , \52361_nG16593 );
_DC g18b6b_GF_IsGateDCbyConstraint ( \52363_nG18b6b , \52362 , \42503 );
buf \U$40475 ( \52364 , \52363_nG18b6b );
buf \U$40476 ( \52365 , RIb886af8_14);
_HMUX g16594 ( \52366_nG16594 , RIdbbbd38_4953 , \52365 , \51855 );
_HMUX g16595 ( \52367_nG16595 , RIdbbbd38_4953 , \52366_nG16594 , \51862 );
buf \U$40477 ( \52368 , RIb838a38_182);
_HMUX g16596 ( \52369_nG16596 , RIdbbbd38_4953 , \52368 , \51867 );
_HMUX g16597 ( \52370_nG16597 , \52367_nG16595 , \52369_nG16596 , \51874 );
buf \U$40478 ( \52371 , \52370_nG16597 );
_DC g18b6d_GF_IsGateDCbyConstraint ( \52372_nG18b6d , \52371 , \42503 );
buf \U$40479 ( \52373 , \52372_nG18b6d );
buf \U$40480 ( \52374 , RIb886b70_13);
_HMUX g16598 ( \52375_nG16598 , RIdbdcdf8_4954 , \52374 , \51855 );
_HMUX g16599 ( \52376_nG16599 , RIdbdcdf8_4954 , \52375_nG16598 , \51862 );
buf \U$40481 ( \52377 , RIb838ab0_181);
_HMUX g1659a ( \52378_nG1659a , RIdbdcdf8_4954 , \52377 , \51867 );
_HMUX g1659b ( \52379_nG1659b , \52376_nG16599 , \52378_nG1659a , \51874 );
buf \U$40482 ( \52380 , \52379_nG1659b );
_DC g18b6f_GF_IsGateDCbyConstraint ( \52381_nG18b6f , \52380 , \42503 );
buf \U$40483 ( \52382 , \52381_nG18b6f );
buf \U$40484 ( \52383 , RIb886be8_12);
_HMUX g1659c ( \52384_nG1659c , RIdb5db80_4955 , \52383 , \51855 );
_HMUX g1659d ( \52385_nG1659d , RIdb5db80_4955 , \52384_nG1659c , \51862 );
buf \U$40485 ( \52386 , RIb838b28_180);
_HMUX g1659e ( \52387_nG1659e , RIdb5db80_4955 , \52386 , \51867 );
_HMUX g1659f ( \52388_nG1659f , \52385_nG1659d , \52387_nG1659e , \51874 );
buf \U$40486 ( \52389 , \52388_nG1659f );
_DC g18b71_GF_IsGateDCbyConstraint ( \52390_nG18b71 , \52389 , \42503 );
buf \U$40487 ( \52391 , \52390_nG18b71 );
buf \U$40488 ( \52392 , RIb886c60_11);
_HMUX g165a0 ( \52393_nG165a0 , RIdb48190_4956 , \52392 , \51855 );
_HMUX g165a1 ( \52394_nG165a1 , RIdb48190_4956 , \52393_nG165a0 , \51862 );
buf \U$40489 ( \52395 , RIb838ba0_179);
_HMUX g165a2 ( \52396_nG165a2 , RIdb48190_4956 , \52395 , \51867 );
_HMUX g165a3 ( \52397_nG165a3 , \52394_nG165a1 , \52396_nG165a2 , \51874 );
buf \U$40490 ( \52398 , \52397_nG165a3 );
_DC g18b73_GF_IsGateDCbyConstraint ( \52399_nG18b73 , \52398 , \42503 );
buf \U$40491 ( \52400 , \52399_nG18b73 );
buf \U$40492 ( \52401 , RIb886cd8_10);
_HMUX g165a4 ( \52402_nG165a4 , RIdb26ba8_4957 , \52401 , \51855 );
_HMUX g165a5 ( \52403_nG165a5 , RIdb26ba8_4957 , \52402_nG165a4 , \51862 );
buf \U$40493 ( \52404 , RIb838c18_178);
_HMUX g165a6 ( \52405_nG165a6 , RIdb26ba8_4957 , \52404 , \51867 );
_HMUX g165a7 ( \52406_nG165a7 , \52403_nG165a5 , \52405_nG165a6 , \51874 );
buf \U$40494 ( \52407 , \52406_nG165a7 );
_DC g18b77_GF_IsGateDCbyConstraint ( \52408_nG18b77 , \52407 , \42503 );
buf \U$40495 ( \52409 , \52408_nG18b77 );
buf \U$40496 ( \52410 , RIb886d50_9);
_HMUX g165a8 ( \52411_nG165a8 , RId917aa8_4958 , \52410 , \51855 );
_HMUX g165a9 ( \52412_nG165a9 , RId917aa8_4958 , \52411_nG165a8 , \51862 );
buf \U$40497 ( \52413 , RIb838c90_177);
_HMUX g165aa ( \52414_nG165aa , RId917aa8_4958 , \52413 , \51867 );
_HMUX g165ab ( \52415_nG165ab , \52412_nG165a9 , \52414_nG165aa , \51874 );
buf \U$40498 ( \52416 , \52415_nG165ab );
_DC g18b79_GF_IsGateDCbyConstraint ( \52417_nG18b79 , \52416 , \42503 );
buf \U$40499 ( \52418 , \52417_nG18b79 );
buf \U$40500 ( \52419 , RIb886dc8_8);
_HMUX g165ac ( \52420_nG165ac , RId986da8_4959 , \52419 , \51855 );
_HMUX g165ad ( \52421_nG165ad , RId986da8_4959 , \52420_nG165ac , \51862 );
buf \U$40501 ( \52422 , RIb838d08_176);
_HMUX g165ae ( \52423_nG165ae , RId986da8_4959 , \52422 , \51867 );
_HMUX g165af ( \52424_nG165af , \52421_nG165ad , \52423_nG165ae , \51874 );
buf \U$40502 ( \52425 , \52424_nG165af );
_DC g18b7b_GF_IsGateDCbyConstraint ( \52426_nG18b7b , \52425 , \42503 );
buf \U$40503 ( \52427 , \52426_nG18b7b );
buf \U$40504 ( \52428 , RIb886e40_7);
_HMUX g165b0 ( \52429_nG165b0 , RIda7eb60_4960 , \52428 , \51855 );
_HMUX g165b1 ( \52430_nG165b1 , RIda7eb60_4960 , \52429_nG165b0 , \51862 );
buf \U$40505 ( \52431 , RIb838d80_175);
_HMUX g165b2 ( \52432_nG165b2 , RIda7eb60_4960 , \52431 , \51867 );
_HMUX g165b3 ( \52433_nG165b3 , \52430_nG165b1 , \52432_nG165b2 , \51874 );
buf \U$40506 ( \52434 , \52433_nG165b3 );
_DC g18b7d_GF_IsGateDCbyConstraint ( \52435_nG18b7d , \52434 , \42503 );
buf \U$40507 ( \52436 , \52435_nG18b7d );
buf \U$40508 ( \52437 , RIb886eb8_6);
_HMUX g165b4 ( \52438_nG165b4 , RIdaf90e0_4961 , \52437 , \51855 );
_HMUX g165b5 ( \52439_nG165b5 , RIdaf90e0_4961 , \52438_nG165b4 , \51862 );
buf \U$40509 ( \52440 , RIb838df8_174);
_HMUX g165b6 ( \52441_nG165b6 , RIdaf90e0_4961 , \52440 , \51867 );
_HMUX g165b7 ( \52442_nG165b7 , \52439_nG165b5 , \52441_nG165b6 , \51874 );
buf \U$40510 ( \52443 , \52442_nG165b7 );
_DC g18b7f_GF_IsGateDCbyConstraint ( \52444_nG18b7f , \52443 , \42503 );
buf \U$40511 ( \52445 , \52444_nG18b7f );
not \U$40512 ( \52446 , \51854 );
and \U$40513 ( \52447 , \51853 , \52446 );
_HMUX g163b6 ( \52448_nG163b6 , RIdab27a8_4962 , \51852 , \52447 );
_HMUX g163b7 ( \52449_nG163b7 , RIdab27a8_4962 , \52448_nG163b6 , \51862 );
not \U$40514 ( \52450 , \51866 );
and \U$40515 ( \52451 , \51865 , \52450 );
_HMUX g163b9 ( \52452_nG163b9 , RIdab27a8_4962 , \51864 , \52451 );
_HMUX g163ba ( \52453_nG163ba , \52449_nG163b7 , \52452_nG163b9 , \51874 );
buf \U$40516 ( \52454 , \52453_nG163ba );
_DC g18a87_GF_IsGateDCbyConstraint ( \52455_nG18a87 , \52454 , \42503 );
buf \U$40517 ( \52456 , \52455_nG18a87 );
_HMUX g163bb ( \52457_nG163bb , RIdbf1ca8_4963 , \51879 , \52447 );
_HMUX g163bc ( \52458_nG163bc , RIdbf1ca8_4963 , \52457_nG163bb , \51862 );
_HMUX g163bd ( \52459_nG163bd , RIdbf1ca8_4963 , \51882 , \52451 );
_HMUX g163be ( \52460_nG163be , \52458_nG163bc , \52459_nG163bd , \51874 );
buf \U$40518 ( \52461 , \52460_nG163be );
_DC g18a9d_GF_IsGateDCbyConstraint ( \52462_nG18a9d , \52461 , \42503 );
buf \U$40519 ( \52463 , \52462_nG18a9d );
_HMUX g163bf ( \52464_nG163bf , RIdc00a50_4964 , \51888 , \52447 );
_HMUX g163c0 ( \52465_nG163c0 , RIdc00a50_4964 , \52464_nG163bf , \51862 );
_HMUX g163c1 ( \52466_nG163c1 , RIdc00a50_4964 , \51891 , \52451 );
_HMUX g163c2 ( \52467_nG163c2 , \52465_nG163c0 , \52466_nG163c1 , \51874 );
buf \U$40520 ( \52468 , \52467_nG163c2 );
_DC g18ab3_GF_IsGateDCbyConstraint ( \52469_nG18ab3 , \52468 , \42503 );
buf \U$40521 ( \52470 , \52469_nG18ab3 );
_HMUX g163c3 ( \52471_nG163c3 , RIdc0fe88_4965 , \51897 , \52447 );
_HMUX g163c4 ( \52472_nG163c4 , RIdc0fe88_4965 , \52471_nG163c3 , \51862 );
_HMUX g163c5 ( \52473_nG163c5 , RIdc0fe88_4965 , \51900 , \52451 );
_HMUX g163c6 ( \52474_nG163c6 , \52472_nG163c4 , \52473_nG163c5 , \51874 );
buf \U$40522 ( \52475 , \52474_nG163c6 );
_DC g18ac9_GF_IsGateDCbyConstraint ( \52476_nG18ac9 , \52475 , \42503 );
buf \U$40523 ( \52477 , \52476_nG18ac9 );
_HMUX g163c7 ( \52478_nG163c7 , RIdc16080_4966 , \51906 , \52447 );
_HMUX g163c8 ( \52479_nG163c8 , RIdc16080_4966 , \52478_nG163c7 , \51862 );
_HMUX g163c9 ( \52480_nG163c9 , RIdc16080_4966 , \51909 , \52451 );
_HMUX g163ca ( \52481_nG163ca , \52479_nG163c8 , \52480_nG163c9 , \51874 );
buf \U$40524 ( \52482 , \52481_nG163ca );
_DC g18adf_GF_IsGateDCbyConstraint ( \52483_nG18adf , \52482 , \42503 );
buf \U$40525 ( \52484 , \52483_nG18adf );
_HMUX g163cb ( \52485_nG163cb , RIdc1c098_4967 , \51915 , \52447 );
_HMUX g163cc ( \52486_nG163cc , RIdc1c098_4967 , \52485_nG163cb , \51862 );
_HMUX g163cd ( \52487_nG163cd , RIdc1c098_4967 , \51918 , \52451 );
_HMUX g163ce ( \52488_nG163ce , \52486_nG163cc , \52487_nG163cd , \51874 );
buf \U$40526 ( \52489 , \52488_nG163ce );
_DC g18af5_GF_IsGateDCbyConstraint ( \52490_nG18af5 , \52489 , \42503 );
buf \U$40527 ( \52491 , \52490_nG18af5 );
_HMUX g163cf ( \52492_nG163cf , RIdc25080_4968 , \51924 , \52447 );
_HMUX g163d0 ( \52493_nG163d0 , RIdc25080_4968 , \52492_nG163cf , \51862 );
_HMUX g163d1 ( \52494_nG163d1 , RIdc25080_4968 , \51927 , \52451 );
_HMUX g163d2 ( \52495_nG163d2 , \52493_nG163d0 , \52494_nG163d1 , \51874 );
buf \U$40528 ( \52496 , \52495_nG163d2 );
_DC g18b01_GF_IsGateDCbyConstraint ( \52497_nG18b01 , \52496 , \42503 );
buf \U$40529 ( \52498 , \52497_nG18b01 );
_HMUX g163d3 ( \52499_nG163d3 , RIdb67810_4969 , \51933 , \52447 );
_HMUX g163d4 ( \52500_nG163d4 , RIdb67810_4969 , \52499_nG163d3 , \51862 );
_HMUX g163d5 ( \52501_nG163d5 , RIdb67810_4969 , \51936 , \52451 );
_HMUX g163d6 ( \52502_nG163d6 , \52500_nG163d4 , \52501_nG163d5 , \51874 );
buf \U$40530 ( \52503 , \52502_nG163d6 );
_DC g18b03_GF_IsGateDCbyConstraint ( \52504_nG18b03 , \52503 , \42503 );
buf \U$40531 ( \52505 , \52504_nG18b03 );
_HMUX g163d7 ( \52506_nG163d7 , RIdda8518_4970 , \51942 , \52447 );
_HMUX g163d8 ( \52507_nG163d8 , RIdda8518_4970 , \52506_nG163d7 , \51862 );
_HMUX g163d9 ( \52508_nG163d9 , RIdda8518_4970 , \51945 , \52451 );
_HMUX g163da ( \52509_nG163da , \52507_nG163d8 , \52508_nG163d9 , \51874 );
buf \U$40532 ( \52510 , \52509_nG163da );
_DC g18b05_GF_IsGateDCbyConstraint ( \52511_nG18b05 , \52510 , \42503 );
buf \U$40533 ( \52512 , \52511_nG18b05 );
_HMUX g163db ( \52513_nG163db , RIdd9d5c8_4971 , \51951 , \52447 );
_HMUX g163dc ( \52514_nG163dc , RIdd9d5c8_4971 , \52513_nG163db , \51862 );
_HMUX g163dd ( \52515_nG163dd , RIdd9d5c8_4971 , \51954 , \52451 );
_HMUX g163de ( \52516_nG163de , \52514_nG163dc , \52515_nG163dd , \51874 );
buf \U$40534 ( \52517 , \52516_nG163de );
_DC g18a89_GF_IsGateDCbyConstraint ( \52518_nG18a89 , \52517 , \42503 );
buf \U$40535 ( \52519 , \52518_nG18a89 );
_HMUX g163df ( \52520_nG163df , RIdd8f270_4972 , \51960 , \52447 );
_HMUX g163e0 ( \52521_nG163e0 , RIdd8f270_4972 , \52520_nG163df , \51862 );
_HMUX g163e1 ( \52522_nG163e1 , RIdd8f270_4972 , \51963 , \52451 );
_HMUX g163e2 ( \52523_nG163e2 , \52521_nG163e0 , \52522_nG163e1 , \51874 );
buf \U$40536 ( \52524 , \52523_nG163e2 );
_DC g18a8b_GF_IsGateDCbyConstraint ( \52525_nG18a8b , \52524 , \42503 );
buf \U$40537 ( \52526 , \52525_nG18a8b );
_HMUX g163e3 ( \52527_nG163e3 , RIdd82fe8_4973 , \51969 , \52447 );
_HMUX g163e4 ( \52528_nG163e4 , RIdd82fe8_4973 , \52527_nG163e3 , \51862 );
_HMUX g163e5 ( \52529_nG163e5 , RIdd82fe8_4973 , \51972 , \52451 );
_HMUX g163e6 ( \52530_nG163e6 , \52528_nG163e4 , \52529_nG163e5 , \51874 );
buf \U$40538 ( \52531 , \52530_nG163e6 );
_DC g18a8d_GF_IsGateDCbyConstraint ( \52532_nG18a8d , \52531 , \42503 );
buf \U$40539 ( \52533 , \52532_nG18a8d );
_HMUX g163e7 ( \52534_nG163e7 , RIdd74150_4974 , \51978 , \52447 );
_HMUX g163e8 ( \52535_nG163e8 , RIdd74150_4974 , \52534_nG163e7 , \51862 );
_HMUX g163e9 ( \52536_nG163e9 , RIdd74150_4974 , \51981 , \52451 );
_HMUX g163ea ( \52537_nG163ea , \52535_nG163e8 , \52536_nG163e9 , \51874 );
buf \U$40540 ( \52538 , \52537_nG163ea );
_DC g18a8f_GF_IsGateDCbyConstraint ( \52539_nG18a8f , \52538 , \42503 );
buf \U$40541 ( \52540 , \52539_nG18a8f );
_HMUX g163eb ( \52541_nG163eb , RIdc641b8_4975 , \51987 , \52447 );
_HMUX g163ec ( \52542_nG163ec , RIdc641b8_4975 , \52541_nG163eb , \51862 );
_HMUX g163ed ( \52543_nG163ed , RIdc641b8_4975 , \51990 , \52451 );
_HMUX g163ee ( \52544_nG163ee , \52542_nG163ec , \52543_nG163ed , \51874 );
buf \U$40542 ( \52545 , \52544_nG163ee );
_DC g18a91_GF_IsGateDCbyConstraint ( \52546_nG18a91 , \52545 , \42503 );
buf \U$40543 ( \52547 , \52546_nG18a91 );
_HMUX g163ef ( \52548_nG163ef , RIdc54600_4976 , \51996 , \52447 );
_HMUX g163f0 ( \52549_nG163f0 , RIdc54600_4976 , \52548_nG163ef , \51862 );
_HMUX g163f1 ( \52550_nG163f1 , RIdc54600_4976 , \51999 , \52451 );
_HMUX g163f2 ( \52551_nG163f2 , \52549_nG163f0 , \52550_nG163f1 , \51874 );
buf \U$40544 ( \52552 , \52551_nG163f2 );
_DC g18a93_GF_IsGateDCbyConstraint ( \52553_nG18a93 , \52552 , \42503 );
buf \U$40545 ( \52554 , \52553_nG18a93 );
_HMUX g163f3 ( \52555_nG163f3 , RIdc46848_4977 , \52005 , \52447 );
_HMUX g163f4 ( \52556_nG163f4 , RIdc46848_4977 , \52555_nG163f3 , \51862 );
_HMUX g163f5 ( \52557_nG163f5 , RIdc46848_4977 , \52008 , \52451 );
_HMUX g163f6 ( \52558_nG163f6 , \52556_nG163f4 , \52557_nG163f5 , \51874 );
buf \U$40546 ( \52559 , \52558_nG163f6 );
_DC g18a95_GF_IsGateDCbyConstraint ( \52560_nG18a95 , \52559 , \42503 );
buf \U$40547 ( \52561 , \52560_nG18a95 );
_HMUX g163f7 ( \52562_nG163f7 , RIdc3b970_4978 , \52014 , \52447 );
_HMUX g163f8 ( \52563_nG163f8 , RIdc3b970_4978 , \52562_nG163f7 , \51862 );
_HMUX g163f9 ( \52564_nG163f9 , RIdc3b970_4978 , \52017 , \52451 );
_HMUX g163fa ( \52565_nG163fa , \52563_nG163f8 , \52564_nG163f9 , \51874 );
buf \U$40548 ( \52566 , \52565_nG163fa );
_DC g18a97_GF_IsGateDCbyConstraint ( \52567_nG18a97 , \52566 , \42503 );
buf \U$40549 ( \52568 , \52567_nG18a97 );
_HMUX g163fb ( \52569_nG163fb , RIdf77220_4979 , \52023 , \52447 );
_HMUX g163fc ( \52570_nG163fc , RIdf77220_4979 , \52569_nG163fb , \51862 );
_HMUX g163fd ( \52571_nG163fd , RIdf77220_4979 , \52026 , \52451 );
_HMUX g163fe ( \52572_nG163fe , \52570_nG163fc , \52571_nG163fd , \51874 );
buf \U$40550 ( \52573 , \52572_nG163fe );
_DC g18a99_GF_IsGateDCbyConstraint ( \52574_nG18a99 , \52573 , \42503 );
buf \U$40551 ( \52575 , \52574_nG18a99 );
_HMUX g163ff ( \52576_nG163ff , RIdf79f98_4980 , \52032 , \52447 );
_HMUX g16400 ( \52577_nG16400 , RIdf79f98_4980 , \52576_nG163ff , \51862 );
_HMUX g16401 ( \52578_nG16401 , RIdf79f98_4980 , \52035 , \52451 );
_HMUX g16402 ( \52579_nG16402 , \52577_nG16400 , \52578_nG16401 , \51874 );
buf \U$40552 ( \52580 , \52579_nG16402 );
_DC g18a9b_GF_IsGateDCbyConstraint ( \52581_nG18a9b , \52580 , \42503 );
buf \U$40553 ( \52582 , \52581_nG18a9b );
_HMUX g16403 ( \52583_nG16403 , RIdf7c860_4981 , \52041 , \52447 );
_HMUX g16404 ( \52584_nG16404 , RIdf7c860_4981 , \52583_nG16403 , \51862 );
_HMUX g16405 ( \52585_nG16405 , RIdf7c860_4981 , \52044 , \52451 );
_HMUX g16406 ( \52586_nG16406 , \52584_nG16404 , \52585_nG16405 , \51874 );
buf \U$40554 ( \52587 , \52586_nG16406 );
_DC g18a9f_GF_IsGateDCbyConstraint ( \52588_nG18a9f , \52587 , \42503 );
buf \U$40555 ( \52589 , \52588_nG18a9f );
_HMUX g16407 ( \52590_nG16407 , RIdf7ff38_4982 , \52050 , \52447 );
_HMUX g16408 ( \52591_nG16408 , RIdf7ff38_4982 , \52590_nG16407 , \51862 );
_HMUX g16409 ( \52592_nG16409 , RIdf7ff38_4982 , \52053 , \52451 );
_HMUX g1640a ( \52593_nG1640a , \52591_nG16408 , \52592_nG16409 , \51874 );
buf \U$40556 ( \52594 , \52593_nG1640a );
_DC g18aa1_GF_IsGateDCbyConstraint ( \52595_nG18aa1 , \52594 , \42503 );
buf \U$40557 ( \52596 , \52595_nG18aa1 );
_HMUX g1640b ( \52597_nG1640b , RIdf82800_4983 , \52059 , \52447 );
_HMUX g1640c ( \52598_nG1640c , RIdf82800_4983 , \52597_nG1640b , \51862 );
_HMUX g1640d ( \52599_nG1640d , RIdf82800_4983 , \52062 , \52451 );
_HMUX g1640e ( \52600_nG1640e , \52598_nG1640c , \52599_nG1640d , \51874 );
buf \U$40558 ( \52601 , \52600_nG1640e );
_DC g18aa3_GF_IsGateDCbyConstraint ( \52602_nG18aa3 , \52601 , \42503 );
buf \U$40559 ( \52603 , \52602_nG18aa3 );
_HMUX g1640f ( \52604_nG1640f , RIdf85ed8_4984 , \52068 , \52447 );
_HMUX g16410 ( \52605_nG16410 , RIdf85ed8_4984 , \52604_nG1640f , \51862 );
_HMUX g16411 ( \52606_nG16411 , RIdf85ed8_4984 , \52071 , \52451 );
_HMUX g16412 ( \52607_nG16412 , \52605_nG16410 , \52606_nG16411 , \51874 );
buf \U$40560 ( \52608 , \52607_nG16412 );
_DC g18aa5_GF_IsGateDCbyConstraint ( \52609_nG18aa5 , \52608 , \42503 );
buf \U$40561 ( \52610 , \52609_nG18aa5 );
_HMUX g16413 ( \52611_nG16413 , RIdf887a0_4985 , \52077 , \52447 );
_HMUX g16414 ( \52612_nG16414 , RIdf887a0_4985 , \52611_nG16413 , \51862 );
_HMUX g16415 ( \52613_nG16415 , RIdf887a0_4985 , \52080 , \52451 );
_HMUX g16416 ( \52614_nG16416 , \52612_nG16414 , \52613_nG16415 , \51874 );
buf \U$40562 ( \52615 , \52614_nG16416 );
_DC g18aa7_GF_IsGateDCbyConstraint ( \52616_nG18aa7 , \52615 , \42503 );
buf \U$40563 ( \52617 , \52616_nG18aa7 );
_HMUX g16417 ( \52618_nG16417 , RIdf8be78_4986 , \52086 , \52447 );
_HMUX g16418 ( \52619_nG16418 , RIdf8be78_4986 , \52618_nG16417 , \51862 );
_HMUX g16419 ( \52620_nG16419 , RIdf8be78_4986 , \52089 , \52451 );
_HMUX g1641a ( \52621_nG1641a , \52619_nG16418 , \52620_nG16419 , \51874 );
buf \U$40564 ( \52622 , \52621_nG1641a );
_DC g18aa9_GF_IsGateDCbyConstraint ( \52623_nG18aa9 , \52622 , \42503 );
buf \U$40565 ( \52624 , \52623_nG18aa9 );
_HMUX g1641b ( \52625_nG1641b , RIdf8e740_4987 , \52095 , \52447 );
_HMUX g1641c ( \52626_nG1641c , RIdf8e740_4987 , \52625_nG1641b , \51862 );
_HMUX g1641d ( \52627_nG1641d , RIdf8e740_4987 , \52098 , \52451 );
_HMUX g1641e ( \52628_nG1641e , \52626_nG1641c , \52627_nG1641d , \51874 );
buf \U$40566 ( \52629 , \52628_nG1641e );
_DC g18aab_GF_IsGateDCbyConstraint ( \52630_nG18aab , \52629 , \42503 );
buf \U$40567 ( \52631 , \52630_nG18aab );
_HMUX g1641f ( \52632_nG1641f , RIdf91008_4988 , \52104 , \52447 );
_HMUX g16420 ( \52633_nG16420 , RIdf91008_4988 , \52632_nG1641f , \51862 );
_HMUX g16421 ( \52634_nG16421 , RIdf91008_4988 , \52107 , \52451 );
_HMUX g16422 ( \52635_nG16422 , \52633_nG16420 , \52634_nG16421 , \51874 );
buf \U$40568 ( \52636 , \52635_nG16422 );
_DC g18aad_GF_IsGateDCbyConstraint ( \52637_nG18aad , \52636 , \42503 );
buf \U$40569 ( \52638 , \52637_nG18aad );
_HMUX g16423 ( \52639_nG16423 , RIdf946e0_4989 , \52113 , \52447 );
_HMUX g16424 ( \52640_nG16424 , RIdf946e0_4989 , \52639_nG16423 , \51862 );
_HMUX g16425 ( \52641_nG16425 , RIdf946e0_4989 , \52116 , \52451 );
_HMUX g16426 ( \52642_nG16426 , \52640_nG16424 , \52641_nG16425 , \51874 );
buf \U$40570 ( \52643 , \52642_nG16426 );
_DC g18aaf_GF_IsGateDCbyConstraint ( \52644_nG18aaf , \52643 , \42503 );
buf \U$40571 ( \52645 , \52644_nG18aaf );
_HMUX g16427 ( \52646_nG16427 , RIdf96fa8_4990 , \52122 , \52447 );
_HMUX g16428 ( \52647_nG16428 , RIdf96fa8_4990 , \52646_nG16427 , \51862 );
_HMUX g16429 ( \52648_nG16429 , RIdf96fa8_4990 , \52125 , \52451 );
_HMUX g1642a ( \52649_nG1642a , \52647_nG16428 , \52648_nG16429 , \51874 );
buf \U$40572 ( \52650 , \52649_nG1642a );
_DC g18ab1_GF_IsGateDCbyConstraint ( \52651_nG18ab1 , \52650 , \42503 );
buf \U$40573 ( \52652 , \52651_nG18ab1 );
_HMUX g1642b ( \52653_nG1642b , RIdf9a680_4991 , \52131 , \52447 );
_HMUX g1642c ( \52654_nG1642c , RIdf9a680_4991 , \52653_nG1642b , \51862 );
_HMUX g1642d ( \52655_nG1642d , RIdf9a680_4991 , \52134 , \52451 );
_HMUX g1642e ( \52656_nG1642e , \52654_nG1642c , \52655_nG1642d , \51874 );
buf \U$40574 ( \52657 , \52656_nG1642e );
_DC g18ab5_GF_IsGateDCbyConstraint ( \52658_nG18ab5 , \52657 , \42503 );
buf \U$40575 ( \52659 , \52658_nG18ab5 );
_HMUX g1642f ( \52660_nG1642f , RIdf9ccf0_4992 , \52140 , \52447 );
_HMUX g16430 ( \52661_nG16430 , RIdf9ccf0_4992 , \52660_nG1642f , \51862 );
_HMUX g16431 ( \52662_nG16431 , RIdf9ccf0_4992 , \52143 , \52451 );
_HMUX g16432 ( \52663_nG16432 , \52661_nG16430 , \52662_nG16431 , \51874 );
buf \U$40576 ( \52664 , \52663_nG16432 );
_DC g18ab7_GF_IsGateDCbyConstraint ( \52665_nG18ab7 , \52664 , \42503 );
buf \U$40577 ( \52666 , \52665_nG18ab7 );
_HMUX g16433 ( \52667_nG16433 , RIdf9ec58_4993 , \52149 , \52447 );
_HMUX g16434 ( \52668_nG16434 , RIdf9ec58_4993 , \52667_nG16433 , \51862 );
_HMUX g16435 ( \52669_nG16435 , RIdf9ec58_4993 , \52152 , \52451 );
_HMUX g16436 ( \52670_nG16436 , \52668_nG16434 , \52669_nG16435 , \51874 );
buf \U$40578 ( \52671 , \52670_nG16436 );
_DC g18ab9_GF_IsGateDCbyConstraint ( \52672_nG18ab9 , \52671 , \42503 );
buf \U$40579 ( \52673 , \52672_nG18ab9 );
_HMUX g16437 ( \52674_nG16437 , RIdfa04b8_4994 , \52158 , \52447 );
_HMUX g16438 ( \52675_nG16438 , RIdfa04b8_4994 , \52674_nG16437 , \51862 );
_HMUX g16439 ( \52676_nG16439 , RIdfa04b8_4994 , \52161 , \52451 );
_HMUX g1643a ( \52677_nG1643a , \52675_nG16438 , \52676_nG16439 , \51874 );
buf \U$40580 ( \52678 , \52677_nG1643a );
_DC g18abb_GF_IsGateDCbyConstraint ( \52679_nG18abb , \52678 , \42503 );
buf \U$40581 ( \52680 , \52679_nG18abb );
_HMUX g1643b ( \52681_nG1643b , RIdfa1bb0_4995 , \52167 , \52447 );
_HMUX g1643c ( \52682_nG1643c , RIdfa1bb0_4995 , \52681_nG1643b , \51862 );
_HMUX g1643d ( \52683_nG1643d , RIdfa1bb0_4995 , \52170 , \52451 );
_HMUX g1643e ( \52684_nG1643e , \52682_nG1643c , \52683_nG1643d , \51874 );
buf \U$40582 ( \52685 , \52684_nG1643e );
_DC g18abd_GF_IsGateDCbyConstraint ( \52686_nG18abd , \52685 , \42503 );
buf \U$40583 ( \52687 , \52686_nG18abd );
_HMUX g1643f ( \52688_nG1643f , RIdfa3b18_4996 , \52176 , \52447 );
_HMUX g16440 ( \52689_nG16440 , RIdfa3b18_4996 , \52688_nG1643f , \51862 );
_HMUX g16441 ( \52690_nG16441 , RIdfa3b18_4996 , \52179 , \52451 );
_HMUX g16442 ( \52691_nG16442 , \52689_nG16440 , \52690_nG16441 , \51874 );
buf \U$40584 ( \52692 , \52691_nG16442 );
_DC g18abf_GF_IsGateDCbyConstraint ( \52693_nG18abf , \52692 , \42503 );
buf \U$40585 ( \52694 , \52693_nG18abf );
_HMUX g16443 ( \52695_nG16443 , RIdfa4dd8_4997 , \52185 , \52447 );
_HMUX g16444 ( \52696_nG16444 , RIdfa4dd8_4997 , \52695_nG16443 , \51862 );
_HMUX g16445 ( \52697_nG16445 , RIdfa4dd8_4997 , \52188 , \52451 );
_HMUX g16446 ( \52698_nG16446 , \52696_nG16444 , \52697_nG16445 , \51874 );
buf \U$40586 ( \52699 , \52698_nG16446 );
_DC g18ac1_GF_IsGateDCbyConstraint ( \52700_nG18ac1 , \52699 , \42503 );
buf \U$40587 ( \52701 , \52700_nG18ac1 );
_HMUX g16447 ( \52702_nG16447 , RIdfa6110_4998 , \52194 , \52447 );
_HMUX g16448 ( \52703_nG16448 , RIdfa6110_4998 , \52702_nG16447 , \51862 );
_HMUX g16449 ( \52704_nG16449 , RIdfa6110_4998 , \52197 , \52451 );
_HMUX g1644a ( \52705_nG1644a , \52703_nG16448 , \52704_nG16449 , \51874 );
buf \U$40588 ( \52706 , \52705_nG1644a );
_DC g18ac3_GF_IsGateDCbyConstraint ( \52707_nG18ac3 , \52706 , \42503 );
buf \U$40589 ( \52708 , \52707_nG18ac3 );
_HMUX g1644b ( \52709_nG1644b , RIdfa75b0_4999 , \52203 , \52447 );
_HMUX g1644c ( \52710_nG1644c , RIdfa75b0_4999 , \52709_nG1644b , \51862 );
_HMUX g1644d ( \52711_nG1644d , RIdfa75b0_4999 , \52206 , \52451 );
_HMUX g1644e ( \52712_nG1644e , \52710_nG1644c , \52711_nG1644d , \51874 );
buf \U$40590 ( \52713 , \52712_nG1644e );
_DC g18ac5_GF_IsGateDCbyConstraint ( \52714_nG18ac5 , \52713 , \42503 );
buf \U$40591 ( \52715 , \52714_nG18ac5 );
_HMUX g1644f ( \52716_nG1644f , RIdfa88e8_5000 , \52212 , \52447 );
_HMUX g16450 ( \52717_nG16450 , RIdfa88e8_5000 , \52716_nG1644f , \51862 );
_HMUX g16451 ( \52718_nG16451 , RIdfa88e8_5000 , \52215 , \52451 );
_HMUX g16452 ( \52719_nG16452 , \52717_nG16450 , \52718_nG16451 , \51874 );
buf \U$40592 ( \52720 , \52719_nG16452 );
_DC g18ac7_GF_IsGateDCbyConstraint ( \52721_nG18ac7 , \52720 , \42503 );
buf \U$40593 ( \52722 , \52721_nG18ac7 );
_HMUX g16453 ( \52723_nG16453 , RIdfa9d10_5001 , \52221 , \52447 );
_HMUX g16454 ( \52724_nG16454 , RIdfa9d10_5001 , \52723_nG16453 , \51862 );
_HMUX g16455 ( \52725_nG16455 , RIdfa9d10_5001 , \52224 , \52451 );
_HMUX g16456 ( \52726_nG16456 , \52724_nG16454 , \52725_nG16455 , \51874 );
buf \U$40594 ( \52727 , \52726_nG16456 );
_DC g18acb_GF_IsGateDCbyConstraint ( \52728_nG18acb , \52727 , \42503 );
buf \U$40595 ( \52729 , \52728_nG18acb );
_HMUX g16457 ( \52730_nG16457 , RIdfab048_5002 , \52230 , \52447 );
_HMUX g16458 ( \52731_nG16458 , RIdfab048_5002 , \52730_nG16457 , \51862 );
_HMUX g16459 ( \52732_nG16459 , RIdfab048_5002 , \52233 , \52451 );
_HMUX g1645a ( \52733_nG1645a , \52731_nG16458 , \52732_nG16459 , \51874 );
buf \U$40596 ( \52734 , \52733_nG1645a );
_DC g18acd_GF_IsGateDCbyConstraint ( \52735_nG18acd , \52734 , \42503 );
buf \U$40597 ( \52736 , \52735_nG18acd );
_HMUX g1645b ( \52737_nG1645b , RIdfac218_5003 , \52239 , \52447 );
_HMUX g1645c ( \52738_nG1645c , RIdfac218_5003 , \52737_nG1645b , \51862 );
_HMUX g1645d ( \52739_nG1645d , RIdfac218_5003 , \52242 , \52451 );
_HMUX g1645e ( \52740_nG1645e , \52738_nG1645c , \52739_nG1645d , \51874 );
buf \U$40598 ( \52741 , \52740_nG1645e );
_DC g18acf_GF_IsGateDCbyConstraint ( \52742_nG18acf , \52741 , \42503 );
buf \U$40599 ( \52743 , \52742_nG18acf );
_HMUX g1645f ( \52744_nG1645f , RIdfad460_5004 , \52248 , \52447 );
_HMUX g16460 ( \52745_nG16460 , RIdfad460_5004 , \52744_nG1645f , \51862 );
_HMUX g16461 ( \52746_nG16461 , RIdfad460_5004 , \52251 , \52451 );
_HMUX g16462 ( \52747_nG16462 , \52745_nG16460 , \52746_nG16461 , \51874 );
buf \U$40600 ( \52748 , \52747_nG16462 );
_DC g18ad1_GF_IsGateDCbyConstraint ( \52749_nG18ad1 , \52748 , \42503 );
buf \U$40601 ( \52750 , \52749_nG18ad1 );
_HMUX g16463 ( \52751_nG16463 , RIdfaecc0_5005 , \52257 , \52447 );
_HMUX g16464 ( \52752_nG16464 , RIdfaecc0_5005 , \52751_nG16463 , \51862 );
_HMUX g16465 ( \52753_nG16465 , RIdfaecc0_5005 , \52260 , \52451 );
_HMUX g16466 ( \52754_nG16466 , \52752_nG16464 , \52753_nG16465 , \51874 );
buf \U$40602 ( \52755 , \52754_nG16466 );
_DC g18ad3_GF_IsGateDCbyConstraint ( \52756_nG18ad3 , \52755 , \42503 );
buf \U$40603 ( \52757 , \52756_nG18ad3 );
_HMUX g16467 ( \52758_nG16467 , RIdfb0610_5006 , \52266 , \52447 );
_HMUX g16468 ( \52759_nG16468 , RIdfb0610_5006 , \52758_nG16467 , \51862 );
_HMUX g16469 ( \52760_nG16469 , RIdfb0610_5006 , \52269 , \52451 );
_HMUX g1646a ( \52761_nG1646a , \52759_nG16468 , \52760_nG16469 , \51874 );
buf \U$40604 ( \52762 , \52761_nG1646a );
_DC g18ad5_GF_IsGateDCbyConstraint ( \52763_nG18ad5 , \52762 , \42503 );
buf \U$40605 ( \52764 , \52763_nG18ad5 );
_HMUX g1646b ( \52765_nG1646b , RIdfb1c90_5007 , \52275 , \52447 );
_HMUX g1646c ( \52766_nG1646c , RIdfb1c90_5007 , \52765_nG1646b , \51862 );
_HMUX g1646d ( \52767_nG1646d , RIdfb1c90_5007 , \52278 , \52451 );
_HMUX g1646e ( \52768_nG1646e , \52766_nG1646c , \52767_nG1646d , \51874 );
buf \U$40606 ( \52769 , \52768_nG1646e );
_DC g18ad7_GF_IsGateDCbyConstraint ( \52770_nG18ad7 , \52769 , \42503 );
buf \U$40607 ( \52771 , \52770_nG18ad7 );
_HMUX g1646f ( \52772_nG1646f , RIdfb3310_5008 , \52284 , \52447 );
_HMUX g16470 ( \52773_nG16470 , RIdfb3310_5008 , \52772_nG1646f , \51862 );
_HMUX g16471 ( \52774_nG16471 , RIdfb3310_5008 , \52287 , \52451 );
_HMUX g16472 ( \52775_nG16472 , \52773_nG16470 , \52774_nG16471 , \51874 );
buf \U$40608 ( \52776 , \52775_nG16472 );
_DC g18ad9_GF_IsGateDCbyConstraint ( \52777_nG18ad9 , \52776 , \42503 );
buf \U$40609 ( \52778 , \52777_nG18ad9 );
_HMUX g16473 ( \52779_nG16473 , RIdfb4828_5009 , \52293 , \52447 );
_HMUX g16474 ( \52780_nG16474 , RIdfb4828_5009 , \52779_nG16473 , \51862 );
_HMUX g16475 ( \52781_nG16475 , RIdfb4828_5009 , \52296 , \52451 );
_HMUX g16476 ( \52782_nG16476 , \52780_nG16474 , \52781_nG16475 , \51874 );
buf \U$40610 ( \52783 , \52782_nG16476 );
_DC g18adb_GF_IsGateDCbyConstraint ( \52784_nG18adb , \52783 , \42503 );
buf \U$40611 ( \52785 , \52784_nG18adb );
_HMUX g16477 ( \52786_nG16477 , RIdfb5d40_5010 , \52302 , \52447 );
_HMUX g16478 ( \52787_nG16478 , RIdfb5d40_5010 , \52786_nG16477 , \51862 );
_HMUX g16479 ( \52788_nG16479 , RIdfb5d40_5010 , \52305 , \52451 );
_HMUX g1647a ( \52789_nG1647a , \52787_nG16478 , \52788_nG16479 , \51874 );
buf \U$40612 ( \52790 , \52789_nG1647a );
_DC g18add_GF_IsGateDCbyConstraint ( \52791_nG18add , \52790 , \42503 );
buf \U$40613 ( \52792 , \52791_nG18add );
_HMUX g1647b ( \52793_nG1647b , RIdfb77f8_5011 , \52311 , \52447 );
_HMUX g1647c ( \52794_nG1647c , RIdfb77f8_5011 , \52793_nG1647b , \51862 );
_HMUX g1647d ( \52795_nG1647d , RIdfb77f8_5011 , \52314 , \52451 );
_HMUX g1647e ( \52796_nG1647e , \52794_nG1647c , \52795_nG1647d , \51874 );
buf \U$40614 ( \52797 , \52796_nG1647e );
_DC g18ae1_GF_IsGateDCbyConstraint ( \52798_nG18ae1 , \52797 , \42503 );
buf \U$40615 ( \52799 , \52798_nG18ae1 );
_HMUX g1647f ( \52800_nG1647f , RIdfb92b0_5012 , \52320 , \52447 );
_HMUX g16480 ( \52801_nG16480 , RIdfb92b0_5012 , \52800_nG1647f , \51862 );
_HMUX g16481 ( \52802_nG16481 , RIdfb92b0_5012 , \52323 , \52451 );
_HMUX g16482 ( \52803_nG16482 , \52801_nG16480 , \52802_nG16481 , \51874 );
buf \U$40616 ( \52804 , \52803_nG16482 );
_DC g18ae3_GF_IsGateDCbyConstraint ( \52805_nG18ae3 , \52804 , \42503 );
buf \U$40617 ( \52806 , \52805_nG18ae3 );
_HMUX g16483 ( \52807_nG16483 , RIdfba9a8_5013 , \52329 , \52447 );
_HMUX g16484 ( \52808_nG16484 , RIdfba9a8_5013 , \52807_nG16483 , \51862 );
_HMUX g16485 ( \52809_nG16485 , RIdfba9a8_5013 , \52332 , \52451 );
_HMUX g16486 ( \52810_nG16486 , \52808_nG16484 , \52809_nG16485 , \51874 );
buf \U$40618 ( \52811 , \52810_nG16486 );
_DC g18ae5_GF_IsGateDCbyConstraint ( \52812_nG18ae5 , \52811 , \42503 );
buf \U$40619 ( \52813 , \52812_nG18ae5 );
_HMUX g16487 ( \52814_nG16487 , RIddf2ca8_5014 , \52338 , \52447 );
_HMUX g16488 ( \52815_nG16488 , RIddf2ca8_5014 , \52814_nG16487 , \51862 );
_HMUX g16489 ( \52816_nG16489 , RIddf2ca8_5014 , \52341 , \52451 );
_HMUX g1648a ( \52817_nG1648a , \52815_nG16488 , \52816_nG16489 , \51874 );
buf \U$40620 ( \52818 , \52817_nG1648a );
_DC g18ae7_GF_IsGateDCbyConstraint ( \52819_nG18ae7 , \52818 , \42503 );
buf \U$40621 ( \52820 , \52819_nG18ae7 );
_HMUX g1648b ( \52821_nG1648b , RIddf4580_5015 , \52347 , \52447 );
_HMUX g1648c ( \52822_nG1648c , RIddf4580_5015 , \52821_nG1648b , \51862 );
_HMUX g1648d ( \52823_nG1648d , RIddf4580_5015 , \52350 , \52451 );
_HMUX g1648e ( \52824_nG1648e , \52822_nG1648c , \52823_nG1648d , \51874 );
buf \U$40622 ( \52825 , \52824_nG1648e );
_DC g18ae9_GF_IsGateDCbyConstraint ( \52826_nG18ae9 , \52825 , \42503 );
buf \U$40623 ( \52827 , \52826_nG18ae9 );
_HMUX g1648f ( \52828_nG1648f , RIddf6308_5016 , \52356 , \52447 );
_HMUX g16490 ( \52829_nG16490 , RIddf6308_5016 , \52828_nG1648f , \51862 );
_HMUX g16491 ( \52830_nG16491 , RIddf6308_5016 , \52359 , \52451 );
_HMUX g16492 ( \52831_nG16492 , \52829_nG16490 , \52830_nG16491 , \51874 );
buf \U$40624 ( \52832 , \52831_nG16492 );
_DC g18aeb_GF_IsGateDCbyConstraint ( \52833_nG18aeb , \52832 , \42503 );
buf \U$40625 ( \52834 , \52833_nG18aeb );
_HMUX g16493 ( \52835_nG16493 , RIddf8270_5017 , \52365 , \52447 );
_HMUX g16494 ( \52836_nG16494 , RIddf8270_5017 , \52835_nG16493 , \51862 );
_HMUX g16495 ( \52837_nG16495 , RIddf8270_5017 , \52368 , \52451 );
_HMUX g16496 ( \52838_nG16496 , \52836_nG16494 , \52837_nG16495 , \51874 );
buf \U$40626 ( \52839 , \52838_nG16496 );
_DC g18aed_GF_IsGateDCbyConstraint ( \52840_nG18aed , \52839 , \42503 );
buf \U$40627 ( \52841 , \52840_nG18aed );
_HMUX g16497 ( \52842_nG16497 , RIddf9e90_5018 , \52374 , \52447 );
_HMUX g16498 ( \52843_nG16498 , RIddf9e90_5018 , \52842_nG16497 , \51862 );
_HMUX g16499 ( \52844_nG16499 , RIddf9e90_5018 , \52377 , \52451 );
_HMUX g1649a ( \52845_nG1649a , \52843_nG16498 , \52844_nG16499 , \51874 );
buf \U$40628 ( \52846 , \52845_nG1649a );
_DC g18aef_GF_IsGateDCbyConstraint ( \52847_nG18aef , \52846 , \42503 );
buf \U$40629 ( \52848 , \52847_nG18aef );
_HMUX g1649b ( \52849_nG1649b , RIddfbdf8_5019 , \52383 , \52447 );
_HMUX g1649c ( \52850_nG1649c , RIddfbdf8_5019 , \52849_nG1649b , \51862 );
_HMUX g1649d ( \52851_nG1649d , RIddfbdf8_5019 , \52386 , \52451 );
_HMUX g1649e ( \52852_nG1649e , \52850_nG1649c , \52851_nG1649d , \51874 );
buf \U$40630 ( \52853 , \52852_nG1649e );
_DC g18af1_GF_IsGateDCbyConstraint ( \52854_nG18af1 , \52853 , \42503 );
buf \U$40631 ( \52855 , \52854_nG18af1 );
_HMUX g1649f ( \52856_nG1649f , RIddfdb08_5020 , \52392 , \52447 );
_HMUX g164a0 ( \52857_nG164a0 , RIddfdb08_5020 , \52856_nG1649f , \51862 );
_HMUX g164a1 ( \52858_nG164a1 , RIddfdb08_5020 , \52395 , \52451 );
_HMUX g164a2 ( \52859_nG164a2 , \52857_nG164a0 , \52858_nG164a1 , \51874 );
buf \U$40632 ( \52860 , \52859_nG164a2 );
_DC g18af3_GF_IsGateDCbyConstraint ( \52861_nG18af3 , \52860 , \42503 );
buf \U$40633 ( \52862 , \52861_nG18af3 );
_HMUX g164a3 ( \52863_nG164a3 , RIddff548_5021 , \52401 , \52447 );
_HMUX g164a4 ( \52864_nG164a4 , RIddff548_5021 , \52863_nG164a3 , \51862 );
_HMUX g164a5 ( \52865_nG164a5 , RIddff548_5021 , \52404 , \52451 );
_HMUX g164a6 ( \52866_nG164a6 , \52864_nG164a4 , \52865_nG164a5 , \51874 );
buf \U$40634 ( \52867 , \52866_nG164a6 );
_DC g18af7_GF_IsGateDCbyConstraint ( \52868_nG18af7 , \52867 , \42503 );
buf \U$40635 ( \52869 , \52868_nG18af7 );
_HMUX g164a7 ( \52870_nG164a7 , RIde015a0_5022 , \52410 , \52447 );
_HMUX g164a8 ( \52871_nG164a8 , RIde015a0_5022 , \52870_nG164a7 , \51862 );
_HMUX g164a9 ( \52872_nG164a9 , RIde015a0_5022 , \52413 , \52451 );
_HMUX g164aa ( \52873_nG164aa , \52871_nG164a8 , \52872_nG164a9 , \51874 );
buf \U$40636 ( \52874 , \52873_nG164aa );
_DC g18af9_GF_IsGateDCbyConstraint ( \52875_nG18af9 , \52874 , \42503 );
buf \U$40637 ( \52876 , \52875_nG18af9 );
_HMUX g164ab ( \52877_nG164ab , RIde03508_5023 , \52419 , \52447 );
_HMUX g164ac ( \52878_nG164ac , RIde03508_5023 , \52877_nG164ab , \51862 );
_HMUX g164ad ( \52879_nG164ad , RIde03508_5023 , \52422 , \52451 );
_HMUX g164ae ( \52880_nG164ae , \52878_nG164ac , \52879_nG164ad , \51874 );
buf \U$40638 ( \52881 , \52880_nG164ae );
_DC g18afb_GF_IsGateDCbyConstraint ( \52882_nG18afb , \52881 , \42503 );
buf \U$40639 ( \52883 , \52882_nG18afb );
_HMUX g164af ( \52884_nG164af , RIde04fc0_5024 , \52428 , \52447 );
_HMUX g164b0 ( \52885_nG164b0 , RIde04fc0_5024 , \52884_nG164af , \51862 );
_HMUX g164b1 ( \52886_nG164b1 , RIde04fc0_5024 , \52431 , \52451 );
_HMUX g164b2 ( \52887_nG164b2 , \52885_nG164b0 , \52886_nG164b1 , \51874 );
buf \U$40640 ( \52888 , \52887_nG164b2 );
_DC g18afd_GF_IsGateDCbyConstraint ( \52889_nG18afd , \52888 , \42503 );
buf \U$40641 ( \52890 , \52889_nG18afd );
_HMUX g164b3 ( \52891_nG164b3 , RIe03bbe8_5025 , \52437 , \52447 );
_HMUX g164b4 ( \52892_nG164b4 , RIe03bbe8_5025 , \52891_nG164b3 , \51862 );
_HMUX g164b5 ( \52893_nG164b5 , RIe03bbe8_5025 , \52440 , \52451 );
_HMUX g164b6 ( \52894_nG164b6 , \52892_nG164b4 , \52893_nG164b5 , \51874 );
buf \U$40642 ( \52895 , \52894_nG164b6 );
_DC g18aff_GF_IsGateDCbyConstraint ( \52896_nG18aff , \52895 , \42503 );
buf \U$40643 ( \52897 , \52896_nG18aff );
nor \U$40644 ( \52898 , \51853 , \52446 );
_HMUX g162b4 ( \52899_nG162b4 , RIe039cf8_5026 , \51852 , \52898 );
_HMUX g162b5 ( \52900_nG162b5 , RIe039cf8_5026 , \52899_nG162b4 , \51862 );
nor \U$40645 ( \52901 , \51865 , \52450 );
_HMUX g162b8 ( \52902_nG162b8 , RIe039cf8_5026 , \51864 , \52901 );
_HMUX g162b9 ( \52903_nG162b9 , \52900_nG162b5 , \52902_nG162b8 , \51874 );
buf \U$40646 ( \52904 , \52903_nG162b9 );
_DC g18a07_GF_IsGateDCbyConstraint ( \52905_nG18a07 , \52904 , \42503 );
buf \U$40647 ( \52906 , \52905_nG18a07 );
_HMUX g162ba ( \52907_nG162ba , RIe038600_5027 , \51879 , \52898 );
_HMUX g162bb ( \52908_nG162bb , RIe038600_5027 , \52907_nG162ba , \51862 );
_HMUX g162bc ( \52909_nG162bc , RIe038600_5027 , \51882 , \52901 );
_HMUX g162bd ( \52910_nG162bd , \52908_nG162bb , \52909_nG162bc , \51874 );
buf \U$40648 ( \52911 , \52910_nG162bd );
_DC g18a1d_GF_IsGateDCbyConstraint ( \52912_nG18a1d , \52911 , \42503 );
buf \U$40649 ( \52913 , \52912_nG18a1d );
_HMUX g162be ( \52914_nG162be , RIe0363c8_5028 , \51888 , \52898 );
_HMUX g162bf ( \52915_nG162bf , RIe0363c8_5028 , \52914_nG162be , \51862 );
_HMUX g162c0 ( \52916_nG162c0 , RIe0363c8_5028 , \51891 , \52901 );
_HMUX g162c1 ( \52917_nG162c1 , \52915_nG162bf , \52916_nG162c0 , \51874 );
buf \U$40650 ( \52918 , \52917_nG162c1 );
_DC g18a33_GF_IsGateDCbyConstraint ( \52919_nG18a33 , \52918 , \42503 );
buf \U$40651 ( \52920 , \52919_nG18a33 );
_HMUX g162c2 ( \52921_nG162c2 , RIe033b78_5029 , \51897 , \52898 );
_HMUX g162c3 ( \52922_nG162c3 , RIe033b78_5029 , \52921_nG162c2 , \51862 );
_HMUX g162c4 ( \52923_nG162c4 , RIe033b78_5029 , \51900 , \52901 );
_HMUX g162c5 ( \52924_nG162c5 , \52922_nG162c3 , \52923_nG162c4 , \51874 );
buf \U$40652 ( \52925 , \52924_nG162c5 );
_DC g18a49_GF_IsGateDCbyConstraint ( \52926_nG18a49 , \52925 , \42503 );
buf \U$40653 ( \52927 , \52926_nG18a49 );
_HMUX g162c6 ( \52928_nG162c6 , RIe031580_5030 , \51906 , \52898 );
_HMUX g162c7 ( \52929_nG162c7 , RIe031580_5030 , \52928_nG162c6 , \51862 );
_HMUX g162c8 ( \52930_nG162c8 , RIe031580_5030 , \51909 , \52901 );
_HMUX g162c9 ( \52931_nG162c9 , \52929_nG162c7 , \52930_nG162c8 , \51874 );
buf \U$40654 ( \52932 , \52931_nG162c9 );
_DC g18a5f_GF_IsGateDCbyConstraint ( \52933_nG18a5f , \52932 , \42503 );
buf \U$40655 ( \52934 , \52933_nG18a5f );
_HMUX g162ca ( \52935_nG162ca , RIe02ee98_5031 , \51915 , \52898 );
_HMUX g162cb ( \52936_nG162cb , RIe02ee98_5031 , \52935_nG162ca , \51862 );
_HMUX g162cc ( \52937_nG162cc , RIe02ee98_5031 , \51918 , \52901 );
_HMUX g162cd ( \52938_nG162cd , \52936_nG162cb , \52937_nG162cc , \51874 );
buf \U$40656 ( \52939 , \52938_nG162cd );
_DC g18a75_GF_IsGateDCbyConstraint ( \52940_nG18a75 , \52939 , \42503 );
buf \U$40657 ( \52941 , \52940_nG18a75 );
_HMUX g162ce ( \52942_nG162ce , RIe02c4e0_5032 , \51924 , \52898 );
_HMUX g162cf ( \52943_nG162cf , RIe02c4e0_5032 , \52942_nG162ce , \51862 );
_HMUX g162d0 ( \52944_nG162d0 , RIe02c4e0_5032 , \51927 , \52901 );
_HMUX g162d1 ( \52945_nG162d1 , \52943_nG162cf , \52944_nG162d0 , \51874 );
buf \U$40658 ( \52946 , \52945_nG162d1 );
_DC g18a81_GF_IsGateDCbyConstraint ( \52947_nG18a81 , \52946 , \42503 );
buf \U$40659 ( \52948 , \52947_nG18a81 );
_HMUX g162d2 ( \52949_nG162d2 , RIe02a488_5033 , \51933 , \52898 );
_HMUX g162d3 ( \52950_nG162d3 , RIe02a488_5033 , \52949_nG162d2 , \51862 );
_HMUX g162d4 ( \52951_nG162d4 , RIe02a488_5033 , \51936 , \52901 );
_HMUX g162d5 ( \52952_nG162d5 , \52950_nG162d3 , \52951_nG162d4 , \51874 );
buf \U$40660 ( \52953 , \52952_nG162d5 );
_DC g18a83_GF_IsGateDCbyConstraint ( \52954_nG18a83 , \52953 , \42503 );
buf \U$40661 ( \52955 , \52954_nG18a83 );
_HMUX g162d6 ( \52956_nG162d6 , RIe028958_5034 , \51942 , \52898 );
_HMUX g162d7 ( \52957_nG162d7 , RIe028958_5034 , \52956_nG162d6 , \51862 );
_HMUX g162d8 ( \52958_nG162d8 , RIe028958_5034 , \51945 , \52901 );
_HMUX g162d9 ( \52959_nG162d9 , \52957_nG162d7 , \52958_nG162d8 , \51874 );
buf \U$40662 ( \52960 , \52959_nG162d9 );
_DC g18a85_GF_IsGateDCbyConstraint ( \52961_nG18a85 , \52960 , \42503 );
buf \U$40663 ( \52962 , \52961_nG18a85 );
_HMUX g162da ( \52963_nG162da , RIe026b58_5035 , \51951 , \52898 );
_HMUX g162db ( \52964_nG162db , RIe026b58_5035 , \52963_nG162da , \51862 );
_HMUX g162dc ( \52965_nG162dc , RIe026b58_5035 , \51954 , \52901 );
_HMUX g162dd ( \52966_nG162dd , \52964_nG162db , \52965_nG162dc , \51874 );
buf \U$40664 ( \52967 , \52966_nG162dd );
_DC g18a09_GF_IsGateDCbyConstraint ( \52968_nG18a09 , \52967 , \42503 );
buf \U$40665 ( \52969 , \52968_nG18a09 );
_HMUX g162de ( \52970_nG162de , RIe025460_5036 , \51960 , \52898 );
_HMUX g162df ( \52971_nG162df , RIe025460_5036 , \52970_nG162de , \51862 );
_HMUX g162e0 ( \52972_nG162e0 , RIe025460_5036 , \51963 , \52901 );
_HMUX g162e1 ( \52973_nG162e1 , \52971_nG162df , \52972_nG162e0 , \51874 );
buf \U$40666 ( \52974 , \52973_nG162e1 );
_DC g18a0b_GF_IsGateDCbyConstraint ( \52975_nG18a0b , \52974 , \42503 );
buf \U$40667 ( \52976 , \52975_nG18a0b );
_HMUX g162e2 ( \52977_nG162e2 , RIe023b88_5037 , \51969 , \52898 );
_HMUX g162e3 ( \52978_nG162e3 , RIe023b88_5037 , \52977_nG162e2 , \51862 );
_HMUX g162e4 ( \52979_nG162e4 , RIe023b88_5037 , \51972 , \52901 );
_HMUX g162e5 ( \52980_nG162e5 , \52978_nG162e3 , \52979_nG162e4 , \51874 );
buf \U$40668 ( \52981 , \52980_nG162e5 );
_DC g18a0d_GF_IsGateDCbyConstraint ( \52982_nG18a0d , \52981 , \42503 );
buf \U$40669 ( \52983 , \52982_nG18a0d );
_HMUX g162e6 ( \52984_nG162e6 , RIe021fe0_5038 , \51978 , \52898 );
_HMUX g162e7 ( \52985_nG162e7 , RIe021fe0_5038 , \52984_nG162e6 , \51862 );
_HMUX g162e8 ( \52986_nG162e8 , RIe021fe0_5038 , \51981 , \52901 );
_HMUX g162e9 ( \52987_nG162e9 , \52985_nG162e7 , \52986_nG162e8 , \51874 );
buf \U$40670 ( \52988 , \52987_nG162e9 );
_DC g18a0f_GF_IsGateDCbyConstraint ( \52989_nG18a0f , \52988 , \42503 );
buf \U$40671 ( \52990 , \52989_nG18a0f );
_HMUX g162ea ( \52991_nG162ea , RIe020168_5039 , \51987 , \52898 );
_HMUX g162eb ( \52992_nG162eb , RIe020168_5039 , \52991_nG162ea , \51862 );
_HMUX g162ec ( \52993_nG162ec , RIe020168_5039 , \51990 , \52901 );
_HMUX g162ed ( \52994_nG162ed , \52992_nG162eb , \52993_nG162ec , \51874 );
buf \U$40672 ( \52995 , \52994_nG162ed );
_DC g18a11_GF_IsGateDCbyConstraint ( \52996_nG18a11 , \52995 , \42503 );
buf \U$40673 ( \52997 , \52996_nG18a11 );
_HMUX g162ee ( \52998_nG162ee , RIe01dcd8_5040 , \51996 , \52898 );
_HMUX g162ef ( \52999_nG162ef , RIe01dcd8_5040 , \52998_nG162ee , \51862 );
_HMUX g162f0 ( \53000_nG162f0 , RIe01dcd8_5040 , \51999 , \52901 );
_HMUX g162f1 ( \53001_nG162f1 , \52999_nG162ef , \53000_nG162f0 , \51874 );
buf \U$40674 ( \53002 , \53001_nG162f1 );
_DC g18a13_GF_IsGateDCbyConstraint ( \53003_nG18a13 , \53002 , \42503 );
buf \U$40675 ( \53004 , \53003_nG18a13 );
_HMUX g162f2 ( \53005_nG162f2 , RIe01b758_5041 , \52005 , \52898 );
_HMUX g162f3 ( \53006_nG162f3 , RIe01b758_5041 , \53005_nG162f2 , \51862 );
_HMUX g162f4 ( \53007_nG162f4 , RIe01b758_5041 , \52008 , \52901 );
_HMUX g162f5 ( \53008_nG162f5 , \53006_nG162f3 , \53007_nG162f4 , \51874 );
buf \U$40676 ( \53009 , \53008_nG162f5 );
_DC g18a15_GF_IsGateDCbyConstraint ( \53010_nG18a15 , \53009 , \42503 );
buf \U$40677 ( \53011 , \53010_nG18a15 );
_HMUX g162f6 ( \53012_nG162f6 , RIe018440_5042 , \52014 , \52898 );
_HMUX g162f7 ( \53013_nG162f7 , RIe018440_5042 , \53012_nG162f6 , \51862 );
_HMUX g162f8 ( \53014_nG162f8 , RIe018440_5042 , \52017 , \52901 );
_HMUX g162f9 ( \53015_nG162f9 , \53013_nG162f7 , \53014_nG162f8 , \51874 );
buf \U$40678 ( \53016 , \53015_nG162f9 );
_DC g18a17_GF_IsGateDCbyConstraint ( \53017_nG18a17 , \53016 , \42503 );
buf \U$40679 ( \53018 , \53017_nG18a17 );
_HMUX g162fa ( \53019_nG162fa , RIe0157b8_5043 , \52023 , \52898 );
_HMUX g162fb ( \53020_nG162fb , RIe0157b8_5043 , \53019_nG162fa , \51862 );
_HMUX g162fc ( \53021_nG162fc , RIe0157b8_5043 , \52026 , \52901 );
_HMUX g162fd ( \53022_nG162fd , \53020_nG162fb , \53021_nG162fc , \51874 );
buf \U$40680 ( \53023 , \53022_nG162fd );
_DC g18a19_GF_IsGateDCbyConstraint ( \53024_nG18a19 , \53023 , \42503 );
buf \U$40681 ( \53025 , \53024_nG18a19 );
_HMUX g162fe ( \53026_nG162fe , RIe012590_5044 , \52032 , \52898 );
_HMUX g162ff ( \53027_nG162ff , RIe012590_5044 , \53026_nG162fe , \51862 );
_HMUX g16300 ( \53028_nG16300 , RIe012590_5044 , \52035 , \52901 );
_HMUX g16301 ( \53029_nG16301 , \53027_nG162ff , \53028_nG16300 , \51874 );
buf \U$40682 ( \53030 , \53029_nG16301 );
_DC g18a1b_GF_IsGateDCbyConstraint ( \53031_nG18a1b , \53030 , \42503 );
buf \U$40683 ( \53032 , \53031_nG18a1b );
_HMUX g16302 ( \53033_nG16302 , RIe010628_5045 , \52041 , \52898 );
_HMUX g16303 ( \53034_nG16303 , RIe010628_5045 , \53033_nG16302 , \51862 );
_HMUX g16304 ( \53035_nG16304 , RIe010628_5045 , \52044 , \52901 );
_HMUX g16305 ( \53036_nG16305 , \53034_nG16303 , \53035_nG16304 , \51874 );
buf \U$40684 ( \53037 , \53036_nG16305 );
_DC g18a1f_GF_IsGateDCbyConstraint ( \53038_nG18a1f , \53037 , \42503 );
buf \U$40685 ( \53039 , \53038_nG18a1f );
_HMUX g16306 ( \53040_nG16306 , RIe00d298_5046 , \52050 , \52898 );
_HMUX g16307 ( \53041_nG16307 , RIe00d298_5046 , \53040_nG16306 , \51862 );
_HMUX g16308 ( \53042_nG16308 , RIe00d298_5046 , \52053 , \52901 );
_HMUX g16309 ( \53043_nG16309 , \53041_nG16307 , \53042_nG16308 , \51874 );
buf \U$40686 ( \53044 , \53043_nG16309 );
_DC g18a21_GF_IsGateDCbyConstraint ( \53045_nG18a21 , \53044 , \42503 );
buf \U$40687 ( \53046 , \53045_nG18a21 );
_HMUX g1630a ( \53047_nG1630a , RIe00a778_5047 , \52059 , \52898 );
_HMUX g1630b ( \53048_nG1630b , RIe00a778_5047 , \53047_nG1630a , \51862 );
_HMUX g1630c ( \53049_nG1630c , RIe00a778_5047 , \52062 , \52901 );
_HMUX g1630d ( \53050_nG1630d , \53048_nG1630b , \53049_nG1630c , \51874 );
buf \U$40688 ( \53051 , \53050_nG1630d );
_DC g18a23_GF_IsGateDCbyConstraint ( \53052_nG18a23 , \53051 , \42503 );
buf \U$40689 ( \53053 , \53052_nG18a23 );
_HMUX g1630e ( \53054_nG1630e , RIe007e38_5048 , \52068 , \52898 );
_HMUX g1630f ( \53055_nG1630f , RIe007e38_5048 , \53054_nG1630e , \51862 );
_HMUX g16310 ( \53056_nG16310 , RIe007e38_5048 , \52071 , \52901 );
_HMUX g16311 ( \53057_nG16311 , \53055_nG1630f , \53056_nG16310 , \51874 );
buf \U$40690 ( \53058 , \53057_nG16311 );
_DC g18a25_GF_IsGateDCbyConstraint ( \53059_nG18a25 , \53058 , \42503 );
buf \U$40691 ( \53060 , \53059_nG18a25 );
_HMUX g16312 ( \53061_nG16312 , RIe004df0_5049 , \52077 , \52898 );
_HMUX g16313 ( \53062_nG16313 , RIe004df0_5049 , \53061_nG16312 , \51862 );
_HMUX g16314 ( \53063_nG16314 , RIe004df0_5049 , \52080 , \52901 );
_HMUX g16315 ( \53064_nG16315 , \53062_nG16313 , \53063_nG16314 , \51874 );
buf \U$40692 ( \53065 , \53064_nG16315 );
_DC g18a27_GF_IsGateDCbyConstraint ( \53066_nG18a27 , \53065 , \42503 );
buf \U$40693 ( \53067 , \53066_nG18a27 );
_HMUX g16316 ( \53068_nG16316 , RIe0024b0_5050 , \52086 , \52898 );
_HMUX g16317 ( \53069_nG16317 , RIe0024b0_5050 , \53068_nG16316 , \51862 );
_HMUX g16318 ( \53070_nG16318 , RIe0024b0_5050 , \52089 , \52901 );
_HMUX g16319 ( \53071_nG16319 , \53069_nG16317 , \53070_nG16318 , \51874 );
buf \U$40694 ( \53072 , \53071_nG16319 );
_DC g18a29_GF_IsGateDCbyConstraint ( \53073_nG18a29 , \53072 , \42503 );
buf \U$40695 ( \53074 , \53073_nG18a29 );
_HMUX g1631a ( \53075_nG1631a , RIdfff558_5051 , \52095 , \52898 );
_HMUX g1631b ( \53076_nG1631b , RIdfff558_5051 , \53075_nG1631a , \51862 );
_HMUX g1631c ( \53077_nG1631c , RIdfff558_5051 , \52098 , \52901 );
_HMUX g1631d ( \53078_nG1631d , \53076_nG1631b , \53077_nG1631c , \51874 );
buf \U$40696 ( \53079 , \53078_nG1631d );
_DC g18a2b_GF_IsGateDCbyConstraint ( \53080_nG18a2b , \53079 , \42503 );
buf \U$40697 ( \53081 , \53080_nG18a2b );
_HMUX g1631e ( \53082_nG1631e , RIdffcd08_5052 , \52104 , \52898 );
_HMUX g1631f ( \53083_nG1631f , RIdffcd08_5052 , \53082_nG1631e , \51862 );
_HMUX g16320 ( \53084_nG16320 , RIdffcd08_5052 , \52107 , \52901 );
_HMUX g16321 ( \53085_nG16321 , \53083_nG1631f , \53084_nG16320 , \51874 );
buf \U$40698 ( \53086 , \53085_nG16321 );
_DC g18a2d_GF_IsGateDCbyConstraint ( \53087_nG18a2d , \53086 , \42503 );
buf \U$40699 ( \53088 , \53087_nG18a2d );
_HMUX g16322 ( \53089_nG16322 , RIdffa260_5053 , \52113 , \52898 );
_HMUX g16323 ( \53090_nG16323 , RIdffa260_5053 , \53089_nG16322 , \51862 );
_HMUX g16324 ( \53091_nG16324 , RIdffa260_5053 , \52116 , \52901 );
_HMUX g16325 ( \53092_nG16325 , \53090_nG16323 , \53091_nG16324 , \51874 );
buf \U$40700 ( \53093 , \53092_nG16325 );
_DC g18a2f_GF_IsGateDCbyConstraint ( \53094_nG18a2f , \53093 , \42503 );
buf \U$40701 ( \53095 , \53094_nG18a2f );
_HMUX g16326 ( \53096_nG16326 , RIdff7b78_5054 , \52122 , \52898 );
_HMUX g16327 ( \53097_nG16327 , RIdff7b78_5054 , \53096_nG16326 , \51862 );
_HMUX g16328 ( \53098_nG16328 , RIdff7b78_5054 , \52125 , \52901 );
_HMUX g16329 ( \53099_nG16329 , \53097_nG16327 , \53098_nG16328 , \51874 );
buf \U$40702 ( \53100 , \53099_nG16329 );
_DC g18a31_GF_IsGateDCbyConstraint ( \53101_nG18a31 , \53100 , \42503 );
buf \U$40703 ( \53102 , \53101_nG18a31 );
_HMUX g1632a ( \53103_nG1632a , RIdff4f68_5055 , \52131 , \52898 );
_HMUX g1632b ( \53104_nG1632b , RIdff4f68_5055 , \53103_nG1632a , \51862 );
_HMUX g1632c ( \53105_nG1632c , RIdff4f68_5055 , \52134 , \52901 );
_HMUX g1632d ( \53106_nG1632d , \53104_nG1632b , \53105_nG1632c , \51874 );
buf \U$40704 ( \53107 , \53106_nG1632d );
_DC g18a35_GF_IsGateDCbyConstraint ( \53108_nG18a35 , \53107 , \42503 );
buf \U$40705 ( \53109 , \53108_nG18a35 );
_HMUX g1632e ( \53110_nG1632e , RIdff1ea8_5056 , \52140 , \52898 );
_HMUX g1632f ( \53111_nG1632f , RIdff1ea8_5056 , \53110_nG1632e , \51862 );
_HMUX g16330 ( \53112_nG16330 , RIdff1ea8_5056 , \52143 , \52901 );
_HMUX g16331 ( \53113_nG16331 , \53111_nG1632f , \53112_nG16330 , \51874 );
buf \U$40706 ( \53114 , \53113_nG16331 );
_DC g18a37_GF_IsGateDCbyConstraint ( \53115_nG18a37 , \53114 , \42503 );
buf \U$40707 ( \53116 , \53115_nG18a37 );
endmodule

