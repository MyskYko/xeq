//
// Conformal-LEC Version 20.10-d130 (26-Jun-2020)
//
module top(RIbb2f070_13,RIbb2eff8_14,RIbb2ef80_15,RIbb2d798_66,RIbb2f160_11,RIbb2f0e8_12,RIbb2d810_65,RIbb2d6a8_68,RIbb2f250_9,
        RIbb2f1d8_10,RIbb2d720_67,RIbb2d5b8_70,RIbb2f340_7,RIbb2f2c8_8,RIbb2d630_69,RIbb2d4c8_72,RIbb2f430_5,RIbb2f3b8_6,RIbb2d540_71,
        RIbb2d3d8_74,RIbb2f520_3,RIbb2f4a8_4,RIbb2d450_73,RIbb2d2e8_76,RIbb2f610_1,RIbb2f598_2,RIbb2d360_75,RIbb2d270_77,RIbb2d1f8_78,
        RIbb2ef08_16,RIbb2ee90_17,RIbb2d180_79,RIbb2d108_80,RIbb2ee18_18,RIbb2eda0_19,RIbb2d090_81,RIbb2ed28_20,RIbb2ecb0_21,RIbb2d018_82,
        RIbb2cfa0_83,RIbb2cf28_84,RIbb2ec38_22,RIbb2ebc0_23,RIbb2ceb0_85,RIbb2ce38_86,RIbb2eb48_24,RIbb2ead0_25,RIbb2cdc0_87,RIbb2cd48_88,
        RIbb2ea58_26,RIbb2e9e0_27,RIbb2ccd0_89,RIbb2cc58_90,RIbb2e968_28,RIbb2e8f0_29,RIbb2cbe0_91,RIbb2cb68_92,RIbb2e878_30,RIbb2e800_31,
        RIbb2caf0_93,RIbb2ca78_94,RIbb2e788_32,RIbb2e710_33,RIbb2ca00_95,RIbb2c988_96,RIbb2e698_34,RIbb2e620_35,RIbb2c910_97,RIbb2c898_98,
        RIbb2e5a8_36,RIbb2e530_37,RIbb2c820_99,RIbb2e4b8_38,RIbb2e440_39,RIbb2c7a8_100,RIbb2c730_101,RIbb2c6b8_102,RIbb2e3c8_40,RIbb2e350_41,
        RIbb2c640_103,RIbb2c5c8_104,RIbb2e2d8_42,RIbb2e260_43,RIbb2c550_105,RIbb2c4d8_106,RIbb2e1e8_44,RIbb2e170_45,RIbb2c460_107,RIbb2c3e8_108,
        RIbb2e0f8_46,RIbb2e080_47,RIbb2c370_109,RIbb2c2f8_110,RIbb2e008_48,RIbb2df90_49,RIbb2c280_111,RIbb2c208_112,RIbb2df18_50,RIbb2dea0_51,
        RIbb2c190_113,RIbb2c118_114,RIbb2de28_52,RIbb2ddb0_53,RIbb2c0a0_115,RIbb2c028_116,RIbb2dd38_54,RIbb2dcc0_55,RIbb2bfb0_117,RIbb2dc48_56,
        RIbb2dbd0_57,RIbb2bf38_118,RIbb2bec0_119,RIbb2be48_120,RIbb2db58_58,RIbb2dae0_59,RIbb2bdd0_121,RIbb2bd58_122,RIbb2da68_60,RIbb2d9f0_61,
        RIbb2bce0_123,RIbb2bc68_124,RIbb2d978_62,RIbb2d900_63,RIbb2bbf0_125,RIbb2bb78_126,RIbb31500_127,RIbb2d888_64,RIbb31578_128,RIbb31668_130,
        RIbb315f0_129,RIbb31758_132,RIbb316e0_131,RIbb31848_134,RIbb317d0_133,RIbb31938_136,RIbb318c0_135,RIbb31a28_138,RIbb319b0_137,RIbb31b18_140,
        RIbb31aa0_139,RIbb31b90_141,RIbb31c08_142,RIbb31c80_143,RIbb31cf8_144,RIbb31d70_145,RIbb31de8_146,RIbb31e60_147,RIbb31ed8_148,RIbb31f50_149,
        RIbb31fc8_150,RIbb32040_151,RIbb320b8_152,RIbb32130_153,RIbb321a8_154,RIbb32220_155,RIbb32298_156,RIbb32310_157,RIbb32388_158,RIbb32400_159,
        RIbb32478_160,RIbb324f0_161,RIbb32568_162,RIbb325e0_163,RIbb32658_164,RIbb326d0_165,RIbb32748_166,RIbb327c0_167,RIbb32838_168,RIbb328b0_169,
        RIbb32928_170,RIbb329a0_171,RIbb32a18_172,RIbb32a90_173,RIbb32b08_174,RIbb32b80_175,RIbb32bf8_176,RIbb32c70_177,RIbb32ce8_178,RIbb32d60_179,
        RIbb32dd8_180,RIbb32e50_181,RIbb32ec8_182,RIbb32f40_183,RIbb32fb8_184,RIbb33030_185,RIbb330a8_186,RIbb33120_187,RIbb33198_188,RIbb33210_189,
        RIbb33288_190,RIbb33300_191,RIbb33378_192,RIbb333f0_193,RIbb33468_194,RIbb334e0_195,RIbb33558_196,RIbb335d0_197,RIbb33648_198,RIbb336c0_199,
        RIbb33738_200,RIbb337b0_201,RIbb33828_202,RIbb338a0_203,RIbb33918_204,RIbb33990_205,RIbb33a08_206,RIbb33a80_207,RIbb33af8_208,RIbb33b70_209,
        RIbb33be8_210,RIbb33c60_211,RIbb33cd8_212,RIbb33d50_213,RIbb33dc8_214,RIbb33e40_215,RIbb33eb8_216,RIbb33f30_217,RIbb33fa8_218,RIbb34020_219,
        RIbb34098_220,RIbb34110_221,RIbb34188_222,RIbb34200_223,RIbb34278_224,RIbb342f0_225,RIbb34368_226,RIbb343e0_227,RIbb34458_228,RIbb344d0_229,
        RIbb34548_230,RIbb345c0_231,RIbb34638_232,RIbb346b0_233,RIbb34728_234,RIbb347a0_235,RIbb34818_236,RIbb34890_237,RIbb34908_238,RIbb34980_239,
        RIbb349f8_240,RIbb34a70_241,RIbb34ae8_242,RIbb34b60_243,RIbb34bd8_244,RIbb34c50_245,RIbb34cc8_246,RIbb34d40_247,RIbb34db8_248,RIbb34e30_249,
        RIbb34ea8_250,RIbb34f20_251,RIbb34f98_252,RIbb35010_253,RIbb35088_254,RIbb35100_255,RIbb35178_256,R_109_95e4d78,R_10a_95e4e20,R_10c_95e4f70,
        R_10f_95e5168,R_111_95e52b8,R_119_95e57f8,R_11c_95e59f0,R_11d_95e5a98,R_11f_95e5be8,R_122_95e5de0,R_123_95e5e88,R_124_95e5f30,R_125_95e5fd8,
        R_127_95e6128,R_128_95e61d0,R_129_95e6278,R_12b_95e63c8,R_12c_95e6470,R_12e_95e65c0,R_12f_95e6668,R_130_95e6710,R_131_95e67b8,R_135_95e6a58,
        R_136_95e6b00,R_137_95e6ba8,R_138_95e6c50,R_139_95e6cf8,R_13b_95e6e48,R_13d_95e6f98,R_13e_95e7040,R_13f_95e70e8,R_140_95e7190,R_141_95e7238,
        R_143_95e7388,R_144_95e7430,R_145_95e74d8,R_146_95e7580,R_147_95e7628,R_148_95e76d0,R_149_95e7778,R_14a_95e7820,R_14b_95e78c8,R_14c_95e7970,
        R_14d_95e7a18,R_14e_95e7ac0,R_14f_95e7b68,R_150_95e7c10,R_151_95e7cb8,R_152_95e7d60,R_153_95e7e08,R_154_95e7eb0,R_155_95e7f58,R_156_95e8000,
        R_157_95e80a8,R_158_95e8150,R_159_95e81f8,R_15a_95e82a0,R_15b_95e8348,R_15c_95e83f0,R_15d_95e8498,R_15e_95e8540,R_15f_95e85e8,R_160_95e8690,
        R_161_95e8738,R_162_95e87e0,R_163_95e8888,R_164_95e8930,R_165_95e89d8,R_166_95e8a80,R_167_95e8b28,R_168_95e8bd0,R_169_95e8c78,R_16a_95e8d20,
        R_16b_95e8dc8,R_16c_95e8e70,R_16d_95e8f18,R_16e_95e8fc0,R_16f_95e9068,R_170_95e9110,R_171_95e91b8,R_172_95e9260,R_173_95e9308,R_174_95e93b0,
        R_175_95e9458,R_176_95e9500);
input RIbb2f070_13,RIbb2eff8_14,RIbb2ef80_15,RIbb2d798_66,RIbb2f160_11,RIbb2f0e8_12,RIbb2d810_65,RIbb2d6a8_68,RIbb2f250_9,
        RIbb2f1d8_10,RIbb2d720_67,RIbb2d5b8_70,RIbb2f340_7,RIbb2f2c8_8,RIbb2d630_69,RIbb2d4c8_72,RIbb2f430_5,RIbb2f3b8_6,RIbb2d540_71,
        RIbb2d3d8_74,RIbb2f520_3,RIbb2f4a8_4,RIbb2d450_73,RIbb2d2e8_76,RIbb2f610_1,RIbb2f598_2,RIbb2d360_75,RIbb2d270_77,RIbb2d1f8_78,
        RIbb2ef08_16,RIbb2ee90_17,RIbb2d180_79,RIbb2d108_80,RIbb2ee18_18,RIbb2eda0_19,RIbb2d090_81,RIbb2ed28_20,RIbb2ecb0_21,RIbb2d018_82,
        RIbb2cfa0_83,RIbb2cf28_84,RIbb2ec38_22,RIbb2ebc0_23,RIbb2ceb0_85,RIbb2ce38_86,RIbb2eb48_24,RIbb2ead0_25,RIbb2cdc0_87,RIbb2cd48_88,
        RIbb2ea58_26,RIbb2e9e0_27,RIbb2ccd0_89,RIbb2cc58_90,RIbb2e968_28,RIbb2e8f0_29,RIbb2cbe0_91,RIbb2cb68_92,RIbb2e878_30,RIbb2e800_31,
        RIbb2caf0_93,RIbb2ca78_94,RIbb2e788_32,RIbb2e710_33,RIbb2ca00_95,RIbb2c988_96,RIbb2e698_34,RIbb2e620_35,RIbb2c910_97,RIbb2c898_98,
        RIbb2e5a8_36,RIbb2e530_37,RIbb2c820_99,RIbb2e4b8_38,RIbb2e440_39,RIbb2c7a8_100,RIbb2c730_101,RIbb2c6b8_102,RIbb2e3c8_40,RIbb2e350_41,
        RIbb2c640_103,RIbb2c5c8_104,RIbb2e2d8_42,RIbb2e260_43,RIbb2c550_105,RIbb2c4d8_106,RIbb2e1e8_44,RIbb2e170_45,RIbb2c460_107,RIbb2c3e8_108,
        RIbb2e0f8_46,RIbb2e080_47,RIbb2c370_109,RIbb2c2f8_110,RIbb2e008_48,RIbb2df90_49,RIbb2c280_111,RIbb2c208_112,RIbb2df18_50,RIbb2dea0_51,
        RIbb2c190_113,RIbb2c118_114,RIbb2de28_52,RIbb2ddb0_53,RIbb2c0a0_115,RIbb2c028_116,RIbb2dd38_54,RIbb2dcc0_55,RIbb2bfb0_117,RIbb2dc48_56,
        RIbb2dbd0_57,RIbb2bf38_118,RIbb2bec0_119,RIbb2be48_120,RIbb2db58_58,RIbb2dae0_59,RIbb2bdd0_121,RIbb2bd58_122,RIbb2da68_60,RIbb2d9f0_61,
        RIbb2bce0_123,RIbb2bc68_124,RIbb2d978_62,RIbb2d900_63,RIbb2bbf0_125,RIbb2bb78_126,RIbb31500_127,RIbb2d888_64,RIbb31578_128,RIbb31668_130,
        RIbb315f0_129,RIbb31758_132,RIbb316e0_131,RIbb31848_134,RIbb317d0_133,RIbb31938_136,RIbb318c0_135,RIbb31a28_138,RIbb319b0_137,RIbb31b18_140,
        RIbb31aa0_139,RIbb31b90_141,RIbb31c08_142,RIbb31c80_143,RIbb31cf8_144,RIbb31d70_145,RIbb31de8_146,RIbb31e60_147,RIbb31ed8_148,RIbb31f50_149,
        RIbb31fc8_150,RIbb32040_151,RIbb320b8_152,RIbb32130_153,RIbb321a8_154,RIbb32220_155,RIbb32298_156,RIbb32310_157,RIbb32388_158,RIbb32400_159,
        RIbb32478_160,RIbb324f0_161,RIbb32568_162,RIbb325e0_163,RIbb32658_164,RIbb326d0_165,RIbb32748_166,RIbb327c0_167,RIbb32838_168,RIbb328b0_169,
        RIbb32928_170,RIbb329a0_171,RIbb32a18_172,RIbb32a90_173,RIbb32b08_174,RIbb32b80_175,RIbb32bf8_176,RIbb32c70_177,RIbb32ce8_178,RIbb32d60_179,
        RIbb32dd8_180,RIbb32e50_181,RIbb32ec8_182,RIbb32f40_183,RIbb32fb8_184,RIbb33030_185,RIbb330a8_186,RIbb33120_187,RIbb33198_188,RIbb33210_189,
        RIbb33288_190,RIbb33300_191,RIbb33378_192,RIbb333f0_193,RIbb33468_194,RIbb334e0_195,RIbb33558_196,RIbb335d0_197,RIbb33648_198,RIbb336c0_199,
        RIbb33738_200,RIbb337b0_201,RIbb33828_202,RIbb338a0_203,RIbb33918_204,RIbb33990_205,RIbb33a08_206,RIbb33a80_207,RIbb33af8_208,RIbb33b70_209,
        RIbb33be8_210,RIbb33c60_211,RIbb33cd8_212,RIbb33d50_213,RIbb33dc8_214,RIbb33e40_215,RIbb33eb8_216,RIbb33f30_217,RIbb33fa8_218,RIbb34020_219,
        RIbb34098_220,RIbb34110_221,RIbb34188_222,RIbb34200_223,RIbb34278_224,RIbb342f0_225,RIbb34368_226,RIbb343e0_227,RIbb34458_228,RIbb344d0_229,
        RIbb34548_230,RIbb345c0_231,RIbb34638_232,RIbb346b0_233,RIbb34728_234,RIbb347a0_235,RIbb34818_236,RIbb34890_237,RIbb34908_238,RIbb34980_239,
        RIbb349f8_240,RIbb34a70_241,RIbb34ae8_242,RIbb34b60_243,RIbb34bd8_244,RIbb34c50_245,RIbb34cc8_246,RIbb34d40_247,RIbb34db8_248,RIbb34e30_249,
        RIbb34ea8_250,RIbb34f20_251,RIbb34f98_252,RIbb35010_253,RIbb35088_254,RIbb35100_255,RIbb35178_256;
output R_109_95e4d78,R_10a_95e4e20,R_10c_95e4f70,R_10f_95e5168,R_111_95e52b8,R_119_95e57f8,R_11c_95e59f0,R_11d_95e5a98,R_11f_95e5be8,
        R_122_95e5de0,R_123_95e5e88,R_124_95e5f30,R_125_95e5fd8,R_127_95e6128,R_128_95e61d0,R_129_95e6278,R_12b_95e63c8,R_12c_95e6470,R_12e_95e65c0,
        R_12f_95e6668,R_130_95e6710,R_131_95e67b8,R_135_95e6a58,R_136_95e6b00,R_137_95e6ba8,R_138_95e6c50,R_139_95e6cf8,R_13b_95e6e48,R_13d_95e6f98,
        R_13e_95e7040,R_13f_95e70e8,R_140_95e7190,R_141_95e7238,R_143_95e7388,R_144_95e7430,R_145_95e74d8,R_146_95e7580,R_147_95e7628,R_148_95e76d0,
        R_149_95e7778,R_14a_95e7820,R_14b_95e78c8,R_14c_95e7970,R_14d_95e7a18,R_14e_95e7ac0,R_14f_95e7b68,R_150_95e7c10,R_151_95e7cb8,R_152_95e7d60,
        R_153_95e7e08,R_154_95e7eb0,R_155_95e7f58,R_156_95e8000,R_157_95e80a8,R_158_95e8150,R_159_95e81f8,R_15a_95e82a0,R_15b_95e8348,R_15c_95e83f0,
        R_15d_95e8498,R_15e_95e8540,R_15f_95e85e8,R_160_95e8690,R_161_95e8738,R_162_95e87e0,R_163_95e8888,R_164_95e8930,R_165_95e89d8,R_166_95e8a80,
        R_167_95e8b28,R_168_95e8bd0,R_169_95e8c78,R_16a_95e8d20,R_16b_95e8dc8,R_16c_95e8e70,R_16d_95e8f18,R_16e_95e8fc0,R_16f_95e9068,R_170_95e9110,
        R_171_95e91b8,R_172_95e9260,R_173_95e9308,R_174_95e93b0,R_175_95e9458,R_176_95e9500;

wire \342_ZERO , \343_ONE , \344 , \345 , \346 , \347 , \348 , \349 , \350 ,
         \351 , \352 , \353 , \354 , \355 , \356 , \357 , \358 , \359 , \360 ,
         \361 , \362 , \363 , \364 , \365 , \366 , \367 , \368 , \369 , \370 ,
         \371 , \372 , \373 , \374 , \375 , \376 , \377 , \378 , \379 , \380 ,
         \381 , \382 , \383 , \384 , \385 , \386 , \387 , \388 , \389 , \390 ,
         \391 , \392 , \393 , \394 , \395 , \396 , \397 , \398 , \399 , \400 ,
         \401 , \402 , \403 , \404 , \405 , \406 , \407 , \408 , \409 , \410 ,
         \411 , \412 , \413 , \414 , \415 , \416 , \417 , \418 , \419 , \420 ,
         \421 , \422 , \423 , \424 , \425 , \426 , \427 , \428 , \429 , \430 ,
         \431 , \432 , \433 , \434 , \435 , \436 , \437 , \438 , \439 , \440 ,
         \441 , \442 , \443 , \444 , \445 , \446 , \447 , \448 , \449 , \450 ,
         \451 , \452 , \453 , \454 , \455 , \456 , \457 , \458 , \459 , \460 ,
         \461 , \462 , \463 , \464 , \465 , \466 , \467 , \468 , \469 , \470 ,
         \471 , \472 , \473 , \474 , \475 , \476 , \477 , \478 , \479 , \480 ,
         \481 , \482 , \483 , \484 , \485 , \486 , \487 , \488 , \489 , \490 ,
         \491 , \492 , \493 , \494 , \495 , \496 , \497 , \498 , \499 , \500 ,
         \501 , \502 , \503 , \504 , \505 , \506 , \507 , \508 , \509 , \510 ,
         \511 , \512 , \513 , \514 , \515 , \516 , \517 , \518 , \519 , \520 ,
         \521 , \522 , \523 , \524 , \525 , \526 , \527 , \528 , \529 , \530 ,
         \531 , \532 , \533 , \534 , \535 , \536 , \537 , \538 , \539 , \540 ,
         \541 , \542 , \543 , \544 , \545 , \546 , \547 , \548 , \549 , \550 ,
         \551 , \552 , \553 , \554 , \555 , \556 , \557 , \558 , \559 , \560 ,
         \561 , \562 , \563 , \564 , \565 , \566 , \567 , \568 , \569 , \570 ,
         \571 , \572 , \573 , \574 , \575 , \576 , \577 , \578 , \579 , \580 ,
         \581 , \582 , \583 , \584 , \585 , \586 , \587 , \588 , \589 , \590 ,
         \591 , \592 , \593 , \594 , \595 , \596 , \597 , \598 , \599 , \600 ,
         \601 , \602 , \603 , \604 , \605 , \606 , \607 , \608 , \609 , \610 ,
         \611 , \612 , \613 , \614 , \615 , \616 , \617 , \618 , \619 , \620 ,
         \621 , \622 , \623 , \624 , \625 , \626 , \627 , \628 , \629 , \630 ,
         \631 , \632 , \633 , \634 , \635 , \636 , \637 , \638 , \639 , \640 ,
         \641 , \642 , \643 , \644 , \645 , \646 , \647 , \648 , \649 , \650 ,
         \651 , \652 , \653 , \654 , \655 , \656 , \657 , \658 , \659 , \660 ,
         \661 , \662 , \663 , \664 , \665 , \666 , \667 , \668 , \669 , \670 ,
         \671 , \672 , \673 , \674 , \675 , \676 , \677 , \678 , \679 , \680 ,
         \681 , \682 , \683 , \684 , \685 , \686 , \687 , \688 , \689 , \690 ,
         \691 , \692 , \693 , \694 , \695 , \696 , \697 , \698 , \699 , \700 ,
         \701 , \702 , \703 , \704 , \705 , \706 , \707 , \708 , \709 , \710 ,
         \711 , \712 , \713 , \714 , \715 , \716 , \717 , \718 , \719 , \720 ,
         \721 , \722 , \723 , \724 , \725 , \726 , \727 , \728 , \729 , \730 ,
         \731 , \732 , \733 , \734 , \735 , \736 , \737 , \738 , \739 , \740 ,
         \741 , \742 , \743 , \744 , \745 , \746 , \747 , \748 , \749 , \750 ,
         \751 , \752 , \753 , \754 , \755 , \756 , \757 , \758 , \759 , \760 ,
         \761 , \762 , \763 , \764 , \765 , \766 , \767 , \768 , \769 , \770 ,
         \771 , \772 , \773 , \774 , \775 , \776 , \777 , \778 , \779 , \780 ,
         \781 , \782 , \783 , \784 , \785 , \786 , \787 , \788 , \789 , \790 ,
         \791 , \792 , \793 , \794 , \795 , \796 , \797 , \798 , \799 , \800 ,
         \801 , \802 , \803 , \804 , \805 , \806 , \807 , \808 , \809 , \810 ,
         \811 , \812 , \813 , \814 , \815 , \816 , \817 , \818 , \819 , \820 ,
         \821 , \822 , \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 ,
         \831 , \832 , \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 ,
         \841 , \842 , \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 ,
         \851 , \852 , \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 ,
         \861 , \862 , \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 ,
         \871 , \872 , \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 ,
         \881 , \882 , \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 ,
         \891 , \892 , \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 ,
         \901 , \902 , \903 , \904 , \905 , \906 , \907 , \908 , \909 , \910 ,
         \911 , \912 , \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 ,
         \921 , \922 , \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 ,
         \931 , \932 , \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 ,
         \941 , \942 , \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 ,
         \951 , \952 , \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 ,
         \961 , \962 , \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 ,
         \971 , \972 , \973 , \974 , \975 , \976 , \977 , \978 , \979 , \980 ,
         \981 , \982 , \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 ,
         \991 , \992 , \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 ,
         \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 ,
         \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 ,
         \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 ,
         \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 ,
         \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 ,
         \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 ,
         \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 ,
         \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 ,
         \1081 , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 ,
         \1091 , \1092 , \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 ,
         \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 ,
         \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 ,
         \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 ,
         \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 ,
         \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 ,
         \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 ,
         \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 ,
         \1171 , \1172 , \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 ,
         \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 ,
         \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 ,
         \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 ,
         \1211 , \1212 , \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 ,
         \1221 , \1222 , \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 ,
         \1231 , \1232 , \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 ,
         \1241 , \1242 , \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 ,
         \1251 , \1252 , \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 ,
         \1261 , \1262 , \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 ,
         \1271 , \1272 , \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 ,
         \1281 , \1282 , \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 ,
         \1291 , \1292 , \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 ,
         \1301 , \1302 , \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 ,
         \1311 , \1312 , \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 ,
         \1321 , \1322 , \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 ,
         \1331 , \1332 , \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 ,
         \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 ,
         \1351 , \1352 , \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 ,
         \1361 , \1362 , \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 ,
         \1371 , \1372 , \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 ,
         \1381 , \1382 , \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 ,
         \1391 , \1392 , \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 ,
         \1401 , \1402 , \1403 , \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 ,
         \1411 , \1412 , \1413 , \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 ,
         \1421 , \1422 , \1423 , \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 ,
         \1431 , \1432 , \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 ,
         \1441 , \1442 , \1443 , \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 ,
         \1451 , \1452 , \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 ,
         \1461 , \1462 , \1463 , \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 ,
         \1471 , \1472 , \1473 , \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 ,
         \1481 , \1482 , \1483 , \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 ,
         \1491 , \1492 , \1493 , \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 ,
         \1501 , \1502 , \1503 , \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 ,
         \1511 , \1512 , \1513 , \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 ,
         \1521 , \1522 , \1523 , \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 ,
         \1531 , \1532 , \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 ,
         \1541 , \1542 , \1543 , \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 ,
         \1551 , \1552 , \1553 , \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 ,
         \1561 , \1562 , \1563 , \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 ,
         \1571 , \1572 , \1573 , \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 ,
         \1581 , \1582 , \1583 , \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 ,
         \1591 , \1592 , \1593 , \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 ,
         \1601 , \1602 , \1603 , \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 ,
         \1611 , \1612 , \1613 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 ,
         \1621 , \1622 , \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 ,
         \1631 , \1632 , \1633 , \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 ,
         \1641 , \1642 , \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 ,
         \1651 , \1652 , \1653 , \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 ,
         \1661 , \1662 , \1663 , \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 ,
         \1671 , \1672 , \1673 , \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 ,
         \1681 , \1682 , \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 ,
         \1691 , \1692 , \1693 , \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 ,
         \1701 , \1702 , \1703 , \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 ,
         \1711 , \1712 , \1713 , \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 ,
         \1721 , \1722 , \1723 , \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 ,
         \1731 , \1732 , \1733 , \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 ,
         \1741 , \1742 , \1743 , \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 ,
         \1751 , \1752 , \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 ,
         \1761 , \1762 , \1763 , \1764 , \1765 , \1766 , \1767 , \1768 , \1769 , \1770 ,
         \1771 , \1772 , \1773 , \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 ,
         \1781 , \1782 , \1783 , \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 ,
         \1791 , \1792 , \1793 , \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 ,
         \1801 , \1802 , \1803 , \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 ,
         \1811 , \1812 , \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 ,
         \1821 , \1822 , \1823 , \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 ,
         \1831 , \1832 , \1833 , \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 ,
         \1841 , \1842 , \1843 , \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 ,
         \1851 , \1852 , \1853 , \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 ,
         \1861 , \1862 , \1863 , \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 ,
         \1871 , \1872 , \1873 , \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 ,
         \1881 , \1882 , \1883 , \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 ,
         \1891 , \1892 , \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 ,
         \1901 , \1902 , \1903 , \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 ,
         \1911 , \1912 , \1913 , \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 ,
         \1921 , \1922 , \1923 , \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 ,
         \1931 , \1932 , \1933 , \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 ,
         \1941 , \1942 , \1943 , \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 ,
         \1951 , \1952 , \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 ,
         \1961 , \1962 , \1963 , \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 ,
         \1971 , \1972 , \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 ,
         \1981 , \1982 , \1983 , \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 ,
         \1991 , \1992 , \1993 , \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 ,
         \2001 , \2002 , \2003 , \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 ,
         \2011 , \2012 , \2013 , \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 ,
         \2021 , \2022 , \2023 , \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 ,
         \2031 , \2032 , \2033 , \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 ,
         \2041 , \2042 , \2043 , \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 ,
         \2051 , \2052 , \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 ,
         \2061 , \2062 , \2063 , \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 ,
         \2071 , \2072 , \2073 , \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 ,
         \2081 , \2082 , \2083 , \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 ,
         \2091 , \2092 , \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 ,
         \2101 , \2102 , \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 ,
         \2111 , \2112 , \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 ,
         \2121 , \2122 , \2123 , \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 ,
         \2131 , \2132 , \2133 , \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 ,
         \2141 , \2142 , \2143 , \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 ,
         \2151 , \2152 , \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 ,
         \2161 , \2162 , \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 ,
         \2171 , \2172 , \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 ,
         \2181 , \2182 , \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 ,
         \2191 , \2192 , \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 ,
         \2201 , \2202 , \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 ,
         \2211 , \2212 , \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 ,
         \2221 , \2222 , \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 ,
         \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 ,
         \2241 , \2242 , \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 ,
         \2251 , \2252 , \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 ,
         \2261 , \2262 , \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 ,
         \2271 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 ,
         \2281 , \2282 , \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 ,
         \2291 , \2292 , \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 ,
         \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 ,
         \2311 , \2312 , \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 ,
         \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 ,
         \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 ,
         \2341 , \2342 , \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 ,
         \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 ,
         \2361 , \2362 , \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 ,
         \2371 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 ,
         \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 ,
         \2391 , \2392 , \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 ,
         \2401 , \2402 , \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 ,
         \2411 , \2412 , \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 ,
         \2421 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 ,
         \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 ,
         \2441 , \2442 , \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 ,
         \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 ,
         \2461 , \2462 , \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 ,
         \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 ,
         \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 ,
         \2491 , \2492 , \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 ,
         \2501 , \2502 , \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 ,
         \2511 , \2512 , \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 ,
         \2521 , \2522 , \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 ,
         \2531 , \2532 , \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 ,
         \2541 , \2542 , \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 ,
         \2551 , \2552 , \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 ,
         \2561 , \2562 , \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 ,
         \2571 , \2572 , \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 ,
         \2581 , \2582 , \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 ,
         \2591 , \2592 , \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 ,
         \2601 , \2602 , \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 ,
         \2611 , \2612 , \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 ,
         \2621 , \2622 , \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 ,
         \2631 , \2632 , \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 ,
         \2641 , \2642 , \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 ,
         \2651 , \2652 , \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 ,
         \2661 , \2662 , \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 ,
         \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 ,
         \2681 , \2682 , \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 ,
         \2691 , \2692 , \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 ,
         \2701 , \2702 , \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 ,
         \2711 , \2712 , \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 ,
         \2721 , \2722 , \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 ,
         \2731 , \2732 , \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 ,
         \2741 , \2742 , \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 ,
         \2751 , \2752 , \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 ,
         \2761 , \2762 , \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 ,
         \2771 , \2772 , \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 ,
         \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 ,
         \2791 , \2792 , \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 ,
         \2801 , \2802 , \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 ,
         \2811 , \2812 , \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 ,
         \2821 , \2822 , \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 ,
         \2831 , \2832 , \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 ,
         \2841 , \2842 , \2843 , \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 ,
         \2851 , \2852 , \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 ,
         \2861 , \2862 , \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 ,
         \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 ,
         \2881 , \2882 , \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 ,
         \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 ,
         \2901 , \2902 , \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 ,
         \2911 , \2912 , \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 ,
         \2921 , \2922 , \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 ,
         \2931 , \2932 , \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 ,
         \2941 , \2942 , \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 ,
         \2951 , \2952 , \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 ,
         \2961 , \2962 , \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 ,
         \2971 , \2972 , \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 ,
         \2981 , \2982 , \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 ,
         \2991 , \2992 , \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 ,
         \3001 , \3002 , \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 ,
         \3011 , \3012 , \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 ,
         \3021 , \3022 , \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 ,
         \3031 , \3032 , \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 ,
         \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 ,
         \3051 , \3052 , \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 ,
         \3061 , \3062 , \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 ,
         \3071 , \3072 , \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 ,
         \3081 , \3082 , \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 ,
         \3091 , \3092 , \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 ,
         \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 ,
         \3111 , \3112 , \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 ,
         \3121 , \3122 , \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 ,
         \3131 , \3132 , \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 ,
         \3141 , \3142 , \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 ,
         \3151 , \3152 , \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 ,
         \3161 , \3162 , \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 ,
         \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 ,
         \3181 , \3182 , \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 ,
         \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 ,
         \3201 , \3202 , \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 ,
         \3211 , \3212 , \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 ,
         \3221 , \3222 , \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 ,
         \3231 , \3232 , \3233 , \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 ,
         \3241 , \3242 , \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 ,
         \3251 , \3252 , \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 ,
         \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 ,
         \3271 , \3272 , \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 ,
         \3281 , \3282 , \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 ,
         \3291 , \3292 , \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 ,
         \3301 , \3302 , \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 ,
         \3311 , \3312 , \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 ,
         \3321 , \3322 , \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 ,
         \3331 , \3332 , \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 ,
         \3341 , \3342 , \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 ,
         \3351 , \3352 , \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 ,
         \3361 , \3362 , \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 ,
         \3371 , \3372 , \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 ,
         \3381 , \3382 , \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 ,
         \3391 , \3392 , \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 ,
         \3401 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 ,
         \3411 , \3412 , \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 ,
         \3421 , \3422 , \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 ,
         \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 ,
         \3441 , \3442 , \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 ,
         \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 ,
         \3461 , \3462 , \3463 , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 ,
         \3471 , \3472 , \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 ,
         \3481 , \3482 , \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 ,
         \3491 , \3492 , \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 ,
         \3501 , \3502 , \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 ,
         \3511 , \3512 , \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 ,
         \3521 , \3522 , \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 ,
         \3531 , \3532 , \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 ,
         \3541 , \3542 , \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 ,
         \3551 , \3552 , \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 ,
         \3561 , \3562 , \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 ,
         \3571 , \3572 , \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 ,
         \3581 , \3582 , \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 ,
         \3591 , \3592 , \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 ,
         \3601 , \3602 , \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 ,
         \3611 , \3612 , \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 ,
         \3621 , \3622 , \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 ,
         \3631 , \3632 , \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 ,
         \3641 , \3642 , \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 ,
         \3651 , \3652 , \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 ,
         \3661 , \3662 , \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 ,
         \3671 , \3672 , \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 ,
         \3681 , \3682 , \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 ,
         \3691 , \3692 , \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 ,
         \3701 , \3702 , \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 ,
         \3711 , \3712 , \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 ,
         \3721 , \3722 , \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 ,
         \3731 , \3732 , \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 ,
         \3741 , \3742 , \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 ,
         \3751 , \3752 , \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 ,
         \3761 , \3762 , \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 ,
         \3771 , \3772 , \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 ,
         \3781 , \3782 , \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 ,
         \3791 , \3792 , \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 ,
         \3801 , \3802 , \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 ,
         \3811 , \3812 , \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 ,
         \3821 , \3822 , \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 ,
         \3831 , \3832 , \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 ,
         \3841 , \3842 , \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 ,
         \3851 , \3852 , \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 ,
         \3861 , \3862 , \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 ,
         \3871 , \3872 , \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 ,
         \3881 , \3882 , \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 ,
         \3891 , \3892 , \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 ,
         \3901 , \3902 , \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 ,
         \3911 , \3912 , \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 ,
         \3921 , \3922 , \3923 , \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 ,
         \3931 , \3932 , \3933 , \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 ,
         \3941 , \3942 , \3943 , \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 ,
         \3951 , \3952 , \3953 , \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 ,
         \3961 , \3962 , \3963 , \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 ,
         \3971 , \3972 , \3973 , \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 ,
         \3981 , \3982 , \3983 , \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 ,
         \3991 , \3992 , \3993 , \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 ,
         \4001 , \4002 , \4003 , \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 ,
         \4011 , \4012 , \4013 , \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 ,
         \4021 , \4022 , \4023 , \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 ,
         \4031 , \4032 , \4033 , \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 ,
         \4041 , \4042 , \4043 , \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 ,
         \4051 , \4052 , \4053 , \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 ,
         \4061 , \4062 , \4063 , \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 ,
         \4071 , \4072 , \4073 , \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 ,
         \4081 , \4082 , \4083 , \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 ,
         \4091 , \4092 , \4093 , \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 ,
         \4101 , \4102 , \4103 , \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 ,
         \4111 , \4112 , \4113 , \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 ,
         \4121 , \4122 , \4123 , \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 ,
         \4131 , \4132 , \4133 , \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 ,
         \4141 , \4142 , \4143 , \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 ,
         \4151 , \4152 , \4153 , \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 ,
         \4161 , \4162 , \4163 , \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 ,
         \4171 , \4172 , \4173 , \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 ,
         \4181 , \4182 , \4183 , \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 ,
         \4191 , \4192 , \4193 , \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 ,
         \4201 , \4202 , \4203 , \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 ,
         \4211 , \4212 , \4213 , \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 ,
         \4221 , \4222 , \4223 , \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 ,
         \4231 , \4232 , \4233 , \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 ,
         \4241 , \4242 , \4243 , \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 ,
         \4251 , \4252 , \4253 , \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 ,
         \4261 , \4262 , \4263 , \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 ,
         \4271 , \4272 , \4273 , \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 ,
         \4281 , \4282 , \4283 , \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 ,
         \4291 , \4292 , \4293 , \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 ,
         \4301 , \4302 , \4303 , \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 ,
         \4311 , \4312 , \4313 , \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 ,
         \4321 , \4322 , \4323 , \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 ,
         \4331 , \4332 , \4333 , \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 ,
         \4341 , \4342 , \4343 , \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 ,
         \4351 , \4352 , \4353 , \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 ,
         \4361 , \4362 , \4363 , \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 ,
         \4371 , \4372 , \4373 , \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 ,
         \4381 , \4382 , \4383 , \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 ,
         \4391 , \4392 , \4393 , \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 ,
         \4401 , \4402 , \4403 , \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 ,
         \4411 , \4412 , \4413 , \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 ,
         \4421 , \4422 , \4423 , \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 ,
         \4431 , \4432 , \4433 , \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 ,
         \4441 , \4442 , \4443 , \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 ,
         \4451 , \4452 , \4453 , \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 ,
         \4461 , \4462 , \4463 , \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 ,
         \4471 , \4472 , \4473 , \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 ,
         \4481 , \4482 , \4483 , \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 ,
         \4491 , \4492 , \4493 , \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 ,
         \4501 , \4502 , \4503 , \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 ,
         \4511 , \4512 , \4513 , \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 ,
         \4521 , \4522 , \4523 , \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 ,
         \4531 , \4532 , \4533 , \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 ,
         \4541 , \4542 , \4543 , \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 ,
         \4551 , \4552 , \4553 , \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 ,
         \4561 , \4562 , \4563 , \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 ,
         \4571 , \4572 , \4573 , \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 ,
         \4581 , \4582 , \4583 , \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 ,
         \4591 , \4592 , \4593 , \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 ,
         \4601 , \4602 , \4603 , \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 ,
         \4611 , \4612 , \4613 , \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 ,
         \4621 , \4622 , \4623 , \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 ,
         \4631 , \4632 , \4633 , \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 ,
         \4641 , \4642 , \4643 , \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 ,
         \4651 , \4652 , \4653 , \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 ,
         \4661 , \4662 , \4663 , \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 ,
         \4671 , \4672 , \4673 , \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 ,
         \4681 , \4682 , \4683 , \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 ,
         \4691 , \4692 , \4693 , \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 ,
         \4701 , \4702 , \4703 , \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 ,
         \4711 , \4712 , \4713 , \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 ,
         \4721 , \4722 , \4723 , \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 ,
         \4731 , \4732 , \4733 , \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 ,
         \4741 , \4742 , \4743 , \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 ,
         \4751 , \4752 , \4753 , \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 ,
         \4761 , \4762 , \4763 , \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 ,
         \4771 , \4772 , \4773 , \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 ,
         \4781 , \4782 , \4783 , \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 ,
         \4791 , \4792 , \4793 , \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 ,
         \4801 , \4802 , \4803 , \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 ,
         \4811 , \4812 , \4813 , \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 ,
         \4821 , \4822 , \4823 , \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 ,
         \4831 , \4832 , \4833 , \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 ,
         \4841 , \4842 , \4843 , \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 ,
         \4851 , \4852 , \4853 , \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 ,
         \4861 , \4862 , \4863 , \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 ,
         \4871 , \4872 , \4873 , \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 ,
         \4881 , \4882 , \4883 , \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 ,
         \4891 , \4892 , \4893 , \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 ,
         \4901 , \4902 , \4903 , \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 ,
         \4911 , \4912 , \4913 , \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 ,
         \4921 , \4922 , \4923 , \4924 , \4925 , \4926 , \4927 , \4928 , \4929 , \4930 ,
         \4931 , \4932 , \4933 , \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 ,
         \4941 , \4942 , \4943 , \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 ,
         \4951 , \4952 , \4953 , \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 ,
         \4961 , \4962 , \4963 , \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 ,
         \4971 , \4972 , \4973 , \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 ,
         \4981 , \4982 , \4983 , \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 ,
         \4991 , \4992 , \4993 , \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 ,
         \5001 , \5002 , \5003 , \5004 , \5005 , \5006 , \5007 , \5008 , \5009 , \5010 ,
         \5011 , \5012 , \5013 , \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 ,
         \5021 , \5022 , \5023 , \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 ,
         \5031 , \5032 , \5033 , \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 ,
         \5041 , \5042 , \5043 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 ,
         \5051 , \5052 , \5053 , \5054 , \5055 , \5056 , \5057 , \5058 , \5059 , \5060 ,
         \5061 , \5062 , \5063 , \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 ,
         \5071 , \5072 , \5073 , \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 ,
         \5081 , \5082 , \5083 , \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 ,
         \5091 , \5092 , \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 ,
         \5101 , \5102 , \5103 , \5104 , \5105 , \5106 , \5107 , \5108 , \5109 , \5110 ,
         \5111 , \5112 , \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 ,
         \5121 , \5122 , \5123 , \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 ,
         \5131 , \5132 , \5133 , \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 ,
         \5141 , \5142 , \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 ,
         \5151 , \5152 , \5153 , \5154 , \5155 , \5156 , \5157 , \5158 , \5159 , \5160 ,
         \5161 , \5162 , \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 ,
         \5171 , \5172 , \5173 , \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 ,
         \5181 , \5182 , \5183 , \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 ,
         \5191 , \5192 , \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 ,
         \5201 , \5202 , \5203 , \5204 , \5205 , \5206 , \5207 , \5208 , \5209 , \5210 ,
         \5211 , \5212 , \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 ,
         \5221 , \5222 , \5223 , \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 ,
         \5231 , \5232 , \5233 , \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 ,
         \5241 , \5242 , \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 ,
         \5251 , \5252 , \5253 , \5254 , \5255 , \5256 , \5257 , \5258 , \5259 , \5260 ,
         \5261 , \5262 , \5263 , \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 ,
         \5271 , \5272 , \5273 , \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 ,
         \5281 , \5282 , \5283 , \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 ,
         \5291 , \5292 , \5293 , \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 ,
         \5301 , \5302 , \5303 , \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 ,
         \5311 , \5312 , \5313 , \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 ,
         \5321 , \5322 , \5323 , \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 ,
         \5331 , \5332 , \5333 , \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 ,
         \5341 , \5342 , \5343 , \5344 , \5345 , \5346 , \5347 , \5348 , \5349 , \5350 ,
         \5351 , \5352 , \5353 , \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 ,
         \5361 , \5362 , \5363 , \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 ,
         \5371 , \5372 , \5373 , \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 ,
         \5381 , \5382 , \5383 , \5384 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 ,
         \5391 , \5392 , \5393 , \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 ,
         \5401 , \5402 , \5403 , \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 ,
         \5411 , \5412 , \5413 , \5414 , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 ,
         \5421 , \5422 , \5423 , \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 ,
         \5431 , \5432 , \5433 , \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 ,
         \5441 , \5442 , \5443 , \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 ,
         \5451 , \5452 , \5453 , \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 ,
         \5461 , \5462 , \5463 , \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 ,
         \5471 , \5472 , \5473 , \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 ,
         \5481 , \5482 , \5483 , \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 ,
         \5491 , \5492 , \5493 , \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 ,
         \5501 , \5502 , \5503 , \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510 ,
         \5511 , \5512 , \5513 , \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 ,
         \5521 , \5522 , \5523 , \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 ,
         \5531 , \5532 , \5533 , \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 ,
         \5541 , \5542 , \5543 , \5544 , \5545 , \5546 , \5547 , \5548 , \5549 , \5550 ,
         \5551 , \5552 , \5553 , \5554 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 ,
         \5561 , \5562 , \5563 , \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 ,
         \5571 , \5572 , \5573 , \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 ,
         \5581 , \5582 , \5583 , \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 ,
         \5591 , \5592 , \5593 , \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 ,
         \5601 , \5602 , \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 ,
         \5611 , \5612 , \5613 , \5614 , \5615 , \5616 , \5617 , \5618 , \5619 , \5620 ,
         \5621 , \5622 , \5623 , \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 ,
         \5631 , \5632 , \5633 , \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 ,
         \5641 , \5642 , \5643 , \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 ,
         \5651 , \5652 , \5653 , \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 ,
         \5661 , \5662 , \5663 , \5664 , \5665 , \5666 , \5667 , \5668 , \5669 , \5670 ,
         \5671 , \5672 , \5673 , \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 ,
         \5681 , \5682 , \5683 , \5684 , \5685 , \5686 , \5687 , \5688 , \5689 , \5690 ,
         \5691 , \5692 , \5693 , \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 ,
         \5701 , \5702 , \5703 , \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 ,
         \5711 , \5712 , \5713 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 ,
         \5721 , \5722 , \5723 , \5724 , \5725 , \5726 , \5727 , \5728 , \5729 , \5730 ,
         \5731 , \5732 , \5733 , \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 ,
         \5741 , \5742 , \5743 , \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 ,
         \5751 , \5752 , \5753 , \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760 ,
         \5761 , \5762 , \5763 , \5764 , \5765 , \5766 , \5767 , \5768 , \5769 , \5770 ,
         \5771 , \5772 , \5773 , \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 ,
         \5781 , \5782 , \5783 , \5784 , \5785 , \5786 , \5787 , \5788 , \5789 , \5790 ,
         \5791 , \5792 , \5793 , \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 ,
         \5801 , \5802 , \5803 , \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 ,
         \5811 , \5812 , \5813 , \5814 , \5815 , \5816 , \5817 , \5818 , \5819 , \5820 ,
         \5821 , \5822 , \5823 , \5824 , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 ,
         \5831 , \5832 , \5833 , \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 ,
         \5841 , \5842 , \5843 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 ,
         \5851 , \5852 , \5853 , \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 ,
         \5861 , \5862 , \5863 , \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 ,
         \5871 , \5872 , \5873 , \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880 ,
         \5881 , \5882 , \5883 , \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 ,
         \5891 , \5892 , \5893 , \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 ,
         \5901 , \5902 , \5903 , \5904 , \5905 , \5906 , \5907 , \5908 , \5909 , \5910 ,
         \5911 , \5912 , \5913 , \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 ,
         \5921 , \5922 , \5923 , \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 ,
         \5931 , \5932 , \5933 , \5934 , \5935 , \5936 , \5937 , \5938 , \5939 , \5940 ,
         \5941 , \5942 , \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 ,
         \5951 , \5952 , \5953 , \5954 , \5955 , \5956 , \5957 , \5958 , \5959 , \5960 ,
         \5961 , \5962 , \5963 , \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 ,
         \5971 , \5972 , \5973 , \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 ,
         \5981 , \5982 , \5983 , \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 ,
         \5991 , \5992 , \5993 , \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 ,
         \6001 , \6002 , \6003 , \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 ,
         \6011 , \6012 , \6013 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 ,
         \6021 , \6022 , \6023 , \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 ,
         \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 ,
         \6041 , \6042 , \6043 , \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050 ,
         \6051 , \6052 , \6053 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 ,
         \6061 , \6062 , \6063 , \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 ,
         \6071 , \6072 , \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 ,
         \6081 , \6082 , \6083 , \6084 , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 ,
         \6091 , \6092 , \6093 , \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 ,
         \6101 , \6102 , \6103 , \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 ,
         \6111 , \6112 , \6113 , \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 ,
         \6121 , \6122 , \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 ,
         \6131 , \6132 , \6133 , \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 ,
         \6141 , \6142 , \6143 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 ,
         \6151 , \6152 , \6153 , \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 ,
         \6161 , \6162 , \6163 , \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 ,
         \6171 , \6172 , \6173 , \6174 , \6175 , \6176 , \6177 , \6178 , \6179 , \6180 ,
         \6181 , \6182 , \6183 , \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 ,
         \6191 , \6192 , \6193 , \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 ,
         \6201 , \6202 , \6203 , \6204 , \6205 , \6206 , \6207 , \6208 , \6209 , \6210 ,
         \6211 , \6212 , \6213 , \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220 ,
         \6221 , \6222 , \6223 , \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 ,
         \6231 , \6232 , \6233 , \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 ,
         \6241 , \6242 , \6243 , \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 ,
         \6251 , \6252 , \6253 , \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 ,
         \6261 , \6262 , \6263 , \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 ,
         \6271 , \6272 , \6273 , \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 ,
         \6281 , \6282 , \6283 , \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 ,
         \6291 , \6292 , \6293 , \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 ,
         \6301 , \6302 , \6303 , \6304 , \6305 , \6306 , \6307 , \6308 , \6309 , \6310 ,
         \6311 , \6312 , \6313 , \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 ,
         \6321 , \6322 , \6323 , \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 ,
         \6331 , \6332 , \6333 , \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 ,
         \6341 , \6342 , \6343 , \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 ,
         \6351 , \6352 , \6353 , \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 ,
         \6361 , \6362 , \6363 , \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 ,
         \6371 , \6372 , \6373 , \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 ,
         \6381 , \6382 , \6383 , \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 ,
         \6391 , \6392 , \6393 , \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 ,
         \6401 , \6402 , \6403 , \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 ,
         \6411 , \6412 , \6413 , \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 ,
         \6421 , \6422 , \6423 , \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 ,
         \6431 , \6432 , \6433 , \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 ,
         \6441 , \6442 , \6443 , \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 ,
         \6451 , \6452 , \6453 , \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 ,
         \6461 , \6462 , \6463 , \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 ,
         \6471 , \6472 , \6473 , \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 ,
         \6481 , \6482 , \6483 , \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 ,
         \6491 , \6492 , \6493 , \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 ,
         \6501 , \6502 , \6503 , \6504 , \6505 , \6506 , \6507 , \6508 , \6509 , \6510 ,
         \6511 , \6512 , \6513 , \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 ,
         \6521 , \6522 , \6523 , \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 ,
         \6531 , \6532 , \6533 , \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 ,
         \6541 , \6542 , \6543 , \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 ,
         \6551 , \6552 , \6553 , \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 ,
         \6561 , \6562 , \6563 , \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 ,
         \6571 , \6572 , \6573 , \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 ,
         \6581 , \6582 , \6583 , \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 ,
         \6591 , \6592 , \6593 , \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 ,
         \6601 , \6602 , \6603 , \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 ,
         \6611 , \6612 , \6613 , \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 ,
         \6621 , \6622 , \6623 , \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 ,
         \6631 , \6632 , \6633 , \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 ,
         \6641 , \6642 , \6643 , \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 ,
         \6651 , \6652 , \6653 , \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 ,
         \6661 , \6662 , \6663 , \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 ,
         \6671 , \6672 , \6673 , \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 ,
         \6681 , \6682 , \6683 , \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 ,
         \6691 , \6692 , \6693 , \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 ,
         \6701 , \6702 , \6703 , \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 ,
         \6711 , \6712 , \6713 , \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 ,
         \6721 , \6722 , \6723 , \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 ,
         \6731 , \6732 , \6733 , \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 ,
         \6741 , \6742 , \6743 , \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 ,
         \6751 , \6752 , \6753 , \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 ,
         \6761 , \6762 , \6763 , \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 ,
         \6771 , \6772 , \6773 , \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 ,
         \6781 , \6782 , \6783 , \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 ,
         \6791 , \6792 , \6793 , \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 ,
         \6801 , \6802 , \6803 , \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 ,
         \6811 , \6812 , \6813 , \6814 , \6815 , \6816 , \6817 , \6818 , \6819 , \6820 ,
         \6821 , \6822 , \6823 , \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 ,
         \6831 , \6832 , \6833 , \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 ,
         \6841 , \6842 , \6843 , \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 ,
         \6851 , \6852 , \6853 , \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 ,
         \6861 , \6862 , \6863 , \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 ,
         \6871 , \6872 , \6873 , \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 ,
         \6881 , \6882 , \6883 , \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 ,
         \6891 , \6892 , \6893 , \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 ,
         \6901 , \6902 , \6903 , \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 ,
         \6911 , \6912 , \6913 , \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 ,
         \6921 , \6922 , \6923 , \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 ,
         \6931 , \6932 , \6933 , \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 ,
         \6941 , \6942 , \6943 , \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 ,
         \6951 , \6952 , \6953 , \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 ,
         \6961 , \6962 , \6963 , \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 ,
         \6971 , \6972 , \6973 , \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 ,
         \6981 , \6982 , \6983 , \6984 , \6985 , \6986 , \6987 , \6988 , \6989 , \6990 ,
         \6991 , \6992 , \6993 , \6994 , \6995 , \6996 , \6997 , \6998 , \6999 , \7000 ,
         \7001 , \7002 , \7003 , \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 ,
         \7011 , \7012 , \7013 , \7014 , \7015 , \7016 , \7017 , \7018 , \7019 , \7020 ,
         \7021 , \7022 , \7023 , \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 ,
         \7031 , \7032 , \7033 , \7034 , \7035 , \7036 , \7037 , \7038 , \7039 , \7040 ,
         \7041 , \7042 , \7043 , \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 ,
         \7051 , \7052 , \7053 , \7054 , \7055 , \7056 , \7057 , \7058 , \7059 , \7060 ,
         \7061 , \7062 , \7063 , \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 ,
         \7071 , \7072 , \7073 , \7074 , \7075 , \7076 , \7077 , \7078 , \7079 , \7080 ,
         \7081 , \7082 , \7083 , \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 ,
         \7091 , \7092 , \7093 , \7094 , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 ,
         \7101 , \7102 , \7103 , \7104 , \7105 , \7106 , \7107 , \7108 , \7109 , \7110 ,
         \7111 , \7112 , \7113 , \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 ,
         \7121 , \7122 , \7123 , \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 ,
         \7131 , \7132 , \7133 , \7134 , \7135 , \7136 , \7137 , \7138 , \7139 , \7140 ,
         \7141 , \7142 , \7143 , \7144 , \7145 , \7146 , \7147 , \7148 , \7149 , \7150 ,
         \7151 , \7152 , \7153 , \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 ,
         \7161 , \7162 , \7163 , \7164 , \7165 , \7166 , \7167 , \7168 , \7169 , \7170 ,
         \7171 , \7172 , \7173 , \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 ,
         \7181 , \7182 , \7183 , \7184 , \7185 , \7186 , \7187 , \7188 , \7189 , \7190 ,
         \7191 , \7192 , \7193 , \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 ,
         \7201 , \7202 , \7203 , \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 ,
         \7211 , \7212 , \7213 , \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 ,
         \7221 , \7222 , \7223 , \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 ,
         \7231 , \7232 , \7233 , \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 ,
         \7241 , \7242 , \7243 , \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 ,
         \7251 , \7252 , \7253 , \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 ,
         \7261 , \7262 , \7263 , \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 ,
         \7271 , \7272 , \7273 , \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 ,
         \7281 , \7282 , \7283 , \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 ,
         \7291 , \7292 , \7293 , \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 ,
         \7301 , \7302 , \7303 , \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 ,
         \7311 , \7312 , \7313 , \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 ,
         \7321 , \7322 , \7323 , \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 ,
         \7331 , \7332 , \7333 , \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 ,
         \7341 , \7342 , \7343 , \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 ,
         \7351 , \7352 , \7353 , \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 ,
         \7361 , \7362 , \7363 , \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 ,
         \7371 , \7372 , \7373 , \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 ,
         \7381 , \7382 , \7383 , \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 ,
         \7391 , \7392 , \7393 , \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 ,
         \7401 , \7402 , \7403 , \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 ,
         \7411 , \7412 , \7413 , \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 ,
         \7421 , \7422 , \7423 , \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 ,
         \7431 , \7432 , \7433 , \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 ,
         \7441 , \7442 , \7443 , \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 ,
         \7451 , \7452 , \7453 , \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 ,
         \7461 , \7462 , \7463 , \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 ,
         \7471 , \7472 , \7473 , \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 ,
         \7481 , \7482 , \7483 , \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 ,
         \7491 , \7492 , \7493 , \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 ,
         \7501 , \7502 , \7503 , \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 ,
         \7511 , \7512 , \7513 , \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 ,
         \7521 , \7522 , \7523 , \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 ,
         \7531 , \7532 , \7533 , \7534 , \7535 , \7536 , \7537 , \7538 , \7539 , \7540 ,
         \7541 , \7542 , \7543 , \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 ,
         \7551 , \7552 , \7553 , \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 ,
         \7561 , \7562 , \7563 , \7564 , \7565 , \7566 , \7567 , \7568 , \7569 , \7570 ,
         \7571 , \7572 , \7573 , \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 ,
         \7581 , \7582 , \7583 , \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 ,
         \7591 , \7592 , \7593 , \7594 , \7595 , \7596 , \7597 , \7598 , \7599 , \7600 ,
         \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 ,
         \7611 , \7612 , \7613 , \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 ,
         \7621 , \7622 , \7623 , \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 ,
         \7631 , \7632 , \7633 , \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 ,
         \7641 , \7642 , \7643 , \7644 , \7645 , \7646 , \7647 , \7648 , \7649 , \7650 ,
         \7651 , \7652 , \7653 , \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 ,
         \7661 , \7662 , \7663 , \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 ,
         \7671 , \7672 , \7673 , \7674 , \7675 , \7676 , \7677 , \7678 , \7679 , \7680 ,
         \7681 , \7682 , \7683 , \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 ,
         \7691 , \7692 , \7693 , \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 ,
         \7701 , \7702 , \7703 , \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 ,
         \7711 , \7712 , \7713 , \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 ,
         \7721 , \7722 , \7723 , \7724 , \7725 , \7726 , \7727 , \7728 , \7729 , \7730 ,
         \7731 , \7732 , \7733 , \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 ,
         \7741 , \7742 , \7743 , \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 ,
         \7751 , \7752 , \7753 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 ,
         \7761 , \7762 , \7763 , \7764 , \7765 , \7766 , \7767 , \7768 , \7769 , \7770 ,
         \7771 , \7772 , \7773 , \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 ,
         \7781 , \7782 , \7783 , \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 ,
         \7791 , \7792 , \7793 , \7794 , \7795 , \7796 , \7797 , \7798 , \7799 , \7800 ,
         \7801 , \7802 , \7803 , \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 ,
         \7811 , \7812 , \7813 , \7814 , \7815 , \7816 , \7817 , \7818 , \7819 , \7820 ,
         \7821 , \7822 , \7823 , \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 ,
         \7831 , \7832 , \7833 , \7834 , \7835 , \7836 , \7837 , \7838 , \7839 , \7840 ,
         \7841 , \7842 , \7843 , \7844 , \7845 , \7846 , \7847 , \7848 , \7849 , \7850 ,
         \7851 , \7852 , \7853 , \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 ,
         \7861 , \7862 , \7863 , \7864 , \7865 , \7866 , \7867 , \7868 , \7869 , \7870 ,
         \7871 , \7872 , \7873 , \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 ,
         \7881 , \7882 , \7883 , \7884 , \7885 , \7886 , \7887 , \7888 , \7889 , \7890 ,
         \7891 , \7892 , \7893 , \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 ,
         \7901 , \7902 , \7903 , \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 ,
         \7911 , \7912 , \7913 , \7914 , \7915 , \7916 , \7917 , \7918 , \7919 , \7920 ,
         \7921 , \7922 , \7923 , \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 ,
         \7931 , \7932 , \7933 , \7934 , \7935 , \7936 , \7937 , \7938 , \7939 , \7940 ,
         \7941 , \7942 , \7943 , \7944 , \7945 , \7946 , \7947 , \7948 , \7949 , \7950 ,
         \7951 , \7952 , \7953 , \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 ,
         \7961 , \7962 , \7963 , \7964 , \7965 , \7966 , \7967 , \7968 , \7969 , \7970 ,
         \7971 , \7972 , \7973 , \7974 , \7975 , \7976 , \7977 , \7978 , \7979 , \7980 ,
         \7981 , \7982 , \7983 , \7984 , \7985 , \7986 , \7987 , \7988 , \7989 , \7990 ,
         \7991 , \7992 , \7993 , \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 ,
         \8001 , \8002 , \8003 , \8004 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 ,
         \8011 , \8012 , \8013 , \8014 , \8015 , \8016 , \8017 , \8018 , \8019 , \8020 ,
         \8021 , \8022 , \8023 , \8024 , \8025 , \8026 , \8027 , \8028 , \8029 , \8030 ,
         \8031 , \8032 , \8033 , \8034 , \8035 , \8036 , \8037 , \8038 , \8039 , \8040 ,
         \8041 , \8042 , \8043 , \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 ,
         \8051 , \8052 , \8053 , \8054 , \8055 , \8056 , \8057 , \8058 , \8059 , \8060 ,
         \8061 , \8062 , \8063 , \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 ,
         \8071 , \8072 , \8073 , \8074 , \8075 , \8076 , \8077 , \8078 , \8079 , \8080 ,
         \8081 , \8082 , \8083 , \8084 , \8085 , \8086 , \8087 , \8088 , \8089 , \8090 ,
         \8091 , \8092 , \8093 , \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 ,
         \8101 , \8102 , \8103 , \8104 , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 ,
         \8111 , \8112 , \8113 , \8114 , \8115 , \8116 , \8117 , \8118 , \8119 , \8120 ,
         \8121 , \8122 , \8123 , \8124 , \8125 , \8126 , \8127 , \8128 , \8129 , \8130 ,
         \8131 , \8132 , \8133 , \8134 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 ,
         \8141 , \8142 , \8143 , \8144 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 ,
         \8151 , \8152 , \8153 , \8154 , \8155 , \8156 , \8157 , \8158 , \8159 , \8160 ,
         \8161 , \8162 , \8163 , \8164 , \8165 , \8166 , \8167 , \8168 , \8169 , \8170 ,
         \8171 , \8172 , \8173 , \8174 , \8175 , \8176 , \8177 , \8178 , \8179 , \8180 ,
         \8181 , \8182 , \8183 , \8184 , \8185 , \8186 , \8187 , \8188 , \8189 , \8190 ,
         \8191 , \8192 , \8193 , \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 ,
         \8201 , \8202 , \8203 , \8204 , \8205 , \8206 , \8207 , \8208 , \8209 , \8210 ,
         \8211 , \8212 , \8213 , \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 ,
         \8221 , \8222 , \8223 , \8224 , \8225 , \8226 , \8227 , \8228 , \8229 , \8230 ,
         \8231 , \8232 , \8233 , \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 ,
         \8241 , \8242 , \8243 , \8244 , \8245 , \8246 , \8247 , \8248 , \8249 , \8250 ,
         \8251 , \8252 , \8253 , \8254 , \8255 , \8256 , \8257 , \8258 , \8259 , \8260 ,
         \8261 , \8262 , \8263 , \8264 , \8265 , \8266 , \8267 , \8268 , \8269 , \8270 ,
         \8271 , \8272 , \8273 , \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 ,
         \8281 , \8282 , \8283 , \8284 , \8285 , \8286 , \8287 , \8288 , \8289 , \8290 ,
         \8291 , \8292 , \8293 , \8294 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 ,
         \8301 , \8302 , \8303 , \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 ,
         \8311 , \8312 , \8313 , \8314 , \8315 , \8316 , \8317 , \8318 , \8319 , \8320 ,
         \8321 , \8322 , \8323 , \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 ,
         \8331 , \8332 , \8333 , \8334 , \8335 , \8336 , \8337 , \8338 , \8339 , \8340 ,
         \8341 , \8342 , \8343 , \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 ,
         \8351 , \8352 , \8353 , \8354 , \8355 , \8356 , \8357 , \8358 , \8359 , \8360 ,
         \8361 , \8362 , \8363 , \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 ,
         \8371 , \8372 , \8373 , \8374 , \8375 , \8376 , \8377 , \8378 , \8379 , \8380 ,
         \8381 , \8382 , \8383 , \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 ,
         \8391 , \8392 , \8393 , \8394 , \8395 , \8396 , \8397 , \8398 , \8399 , \8400 ,
         \8401 , \8402 , \8403 , \8404 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 ,
         \8411 , \8412 , \8413 , \8414 , \8415 , \8416 , \8417 , \8418 , \8419 , \8420 ,
         \8421 , \8422 , \8423 , \8424 , \8425 , \8426 , \8427 , \8428 , \8429 , \8430 ,
         \8431 , \8432 , \8433 , \8434 , \8435 , \8436 , \8437 , \8438 , \8439 , \8440 ,
         \8441 , \8442 , \8443 , \8444 , \8445 , \8446 , \8447 , \8448 , \8449 , \8450 ,
         \8451 , \8452 , \8453 , \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460 ,
         \8461 , \8462 , \8463 , \8464 , \8465 , \8466 , \8467 , \8468 , \8469 , \8470 ,
         \8471 , \8472 , \8473 , \8474 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 ,
         \8481 , \8482 , \8483 , \8484 , \8485 , \8486 , \8487 , \8488 , \8489 , \8490 ,
         \8491 , \8492 , \8493 , \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 ,
         \8501 , \8502 , \8503 , \8504 , \8505 , \8506 , \8507 , \8508 , \8509 , \8510 ,
         \8511 , \8512 , \8513 , \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 ,
         \8521 , \8522 , \8523 , \8524 , \8525 , \8526 , \8527 , \8528 , \8529 , \8530 ,
         \8531 , \8532 , \8533 , \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 ,
         \8541 , \8542 , \8543 , \8544 , \8545 , \8546 , \8547 , \8548 , \8549 , \8550 ,
         \8551 , \8552 , \8553 , \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 ,
         \8561 , \8562 , \8563 , \8564 , \8565 , \8566 , \8567 , \8568 , \8569 , \8570 ,
         \8571 , \8572 , \8573 , \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 ,
         \8581 , \8582 , \8583 , \8584 , \8585 , \8586 , \8587 , \8588 , \8589 , \8590 ,
         \8591 , \8592 , \8593 , \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 ,
         \8601 , \8602 , \8603 , \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 ,
         \8611 , \8612 , \8613 , \8614 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 ,
         \8621 , \8622 , \8623 , \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 ,
         \8631 , \8632 , \8633 , \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 ,
         \8641 , \8642 , \8643 , \8644 , \8645 , \8646 , \8647 , \8648 , \8649 , \8650 ,
         \8651 , \8652 , \8653 , \8654 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 ,
         \8661 , \8662 , \8663 , \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 ,
         \8671 , \8672 , \8673 , \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 ,
         \8681 , \8682 , \8683 , \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 ,
         \8691 , \8692 , \8693 , \8694 , \8695 , \8696 , \8697 , \8698 , \8699 , \8700 ,
         \8701 , \8702 , \8703 , \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 ,
         \8711 , \8712 , \8713 , \8714 , \8715 , \8716 , \8717 , \8718 , \8719 , \8720 ,
         \8721 , \8722 , \8723 , \8724 , \8725 , \8726 , \8727 , \8728 , \8729 , \8730 ,
         \8731 , \8732 , \8733 , \8734 , \8735 , \8736 , \8737 , \8738 , \8739 , \8740 ,
         \8741 , \8742 , \8743 , \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 ,
         \8751 , \8752 , \8753 , \8754 , \8755 , \8756 , \8757 , \8758 , \8759 , \8760 ,
         \8761 , \8762 , \8763 , \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 ,
         \8771 , \8772 , \8773 , \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780 ,
         \8781 , \8782 , \8783 , \8784 , \8785 , \8786 , \8787 , \8788 , \8789 , \8790 ,
         \8791 , \8792 , \8793 , \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 ,
         \8801 , \8802 , \8803 , \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 ,
         \8811 , \8812 , \8813 , \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 ,
         \8821 , \8822 , \8823 , \8824 , \8825 , \8826 , \8827 , \8828 , \8829 , \8830 ,
         \8831 , \8832 , \8833 , \8834 , \8835 , \8836 , \8837 , \8838 , \8839 , \8840 ,
         \8841 , \8842 , \8843 , \8844 , \8845 , \8846 , \8847 , \8848 , \8849 , \8850 ,
         \8851 , \8852 , \8853 , \8854 , \8855 , \8856 , \8857 , \8858 , \8859 , \8860 ,
         \8861 , \8862 , \8863 , \8864 , \8865 , \8866 , \8867 , \8868 , \8869 , \8870 ,
         \8871 , \8872 , \8873 , \8874 , \8875 , \8876 , \8877 , \8878 , \8879 , \8880 ,
         \8881 , \8882 , \8883 , \8884 , \8885 , \8886 , \8887 , \8888 , \8889 , \8890 ,
         \8891 , \8892 , \8893 , \8894 , \8895 , \8896 , \8897 , \8898 , \8899 , \8900 ,
         \8901 , \8902 , \8903 , \8904 , \8905 , \8906 , \8907 , \8908 , \8909 , \8910 ,
         \8911 , \8912 , \8913 , \8914 , \8915 , \8916 , \8917 , \8918 , \8919 , \8920 ,
         \8921 , \8922 , \8923 , \8924 , \8925 , \8926 , \8927 , \8928 , \8929 , \8930 ,
         \8931 , \8932 , \8933 , \8934 , \8935 , \8936 , \8937 , \8938 , \8939 , \8940 ,
         \8941 , \8942 , \8943 , \8944 , \8945 , \8946 , \8947 , \8948 , \8949 , \8950 ,
         \8951 , \8952 , \8953 , \8954 , \8955 , \8956 , \8957 , \8958 , \8959 , \8960 ,
         \8961 , \8962 , \8963 , \8964 , \8965 , \8966 , \8967 , \8968 , \8969 , \8970 ,
         \8971 , \8972 , \8973 , \8974 , \8975 , \8976 , \8977 , \8978 , \8979 , \8980 ,
         \8981 , \8982 , \8983 , \8984 , \8985 , \8986 , \8987 , \8988 , \8989 , \8990 ,
         \8991 , \8992 , \8993 , \8994 , \8995 , \8996 , \8997 , \8998 , \8999 , \9000 ,
         \9001 , \9002 , \9003 , \9004 , \9005 , \9006 , \9007 , \9008 , \9009 , \9010 ,
         \9011 , \9012 , \9013 , \9014 , \9015 , \9016 , \9017 , \9018 , \9019 , \9020 ,
         \9021 , \9022 , \9023 , \9024 , \9025 , \9026 , \9027 , \9028 , \9029 , \9030 ,
         \9031 , \9032 , \9033 , \9034 , \9035 , \9036 , \9037 , \9038 , \9039 , \9040 ,
         \9041 , \9042 , \9043 , \9044 , \9045 , \9046 , \9047 , \9048 , \9049 , \9050 ,
         \9051 , \9052 , \9053 , \9054 , \9055 , \9056 , \9057 , \9058 , \9059 , \9060 ,
         \9061 , \9062 , \9063 , \9064 , \9065 , \9066 , \9067 , \9068 , \9069 , \9070 ,
         \9071 , \9072 , \9073 , \9074 , \9075 , \9076 , \9077 , \9078 , \9079 , \9080 ,
         \9081 , \9082 , \9083 , \9084 , \9085 , \9086 , \9087 , \9088 , \9089 , \9090 ,
         \9091 , \9092 , \9093 , \9094 , \9095 , \9096 , \9097 , \9098 , \9099 , \9100 ,
         \9101 , \9102 , \9103 , \9104 , \9105 , \9106 , \9107 , \9108 , \9109 , \9110 ,
         \9111 , \9112 , \9113 , \9114 , \9115 , \9116 , \9117 , \9118 , \9119 , \9120 ,
         \9121 , \9122 , \9123 , \9124 , \9125 , \9126 , \9127 , \9128 , \9129 , \9130 ,
         \9131 , \9132 , \9133 , \9134 , \9135 , \9136 , \9137 , \9138 , \9139 , \9140 ,
         \9141 , \9142 , \9143 , \9144 , \9145 , \9146 , \9147 , \9148 , \9149 , \9150 ,
         \9151 , \9152 , \9153 , \9154 , \9155 , \9156 , \9157 , \9158 , \9159 , \9160 ,
         \9161 , \9162 , \9163 , \9164 , \9165 , \9166 , \9167 , \9168 , \9169 , \9170 ,
         \9171 , \9172 , \9173 , \9174 , \9175 , \9176 , \9177 , \9178 , \9179 , \9180 ,
         \9181 , \9182 , \9183 , \9184 , \9185 , \9186 , \9187 , \9188 , \9189 , \9190 ,
         \9191 , \9192 , \9193 , \9194 , \9195 , \9196 , \9197 , \9198 , \9199 , \9200 ,
         \9201 , \9202 , \9203 , \9204 , \9205 , \9206 , \9207 , \9208 , \9209 , \9210 ,
         \9211 , \9212 , \9213 , \9214 , \9215 , \9216 , \9217 , \9218 , \9219 , \9220 ,
         \9221 , \9222 , \9223 , \9224 , \9225 , \9226 , \9227 , \9228 , \9229 , \9230 ,
         \9231 , \9232 , \9233 , \9234 , \9235 , \9236 , \9237 , \9238 , \9239 , \9240 ,
         \9241 , \9242 , \9243 , \9244 , \9245 , \9246 , \9247 , \9248 , \9249 , \9250 ,
         \9251 , \9252 , \9253 , \9254 , \9255 , \9256 , \9257 , \9258 , \9259 , \9260 ,
         \9261 , \9262 , \9263 , \9264 , \9265 , \9266 , \9267 , \9268 , \9269 , \9270 ,
         \9271 , \9272 , \9273 , \9274 , \9275 , \9276 , \9277 , \9278 , \9279 , \9280 ,
         \9281 , \9282 , \9283 , \9284 , \9285 , \9286 , \9287 , \9288 , \9289 , \9290 ,
         \9291 , \9292 , \9293 , \9294 , \9295 , \9296 , \9297 , \9298 , \9299 , \9300 ,
         \9301 , \9302 , \9303 , \9304 , \9305 , \9306 , \9307 , \9308 , \9309 , \9310 ,
         \9311 , \9312 , \9313 , \9314 , \9315 , \9316 , \9317 , \9318 , \9319 , \9320 ,
         \9321 , \9322 , \9323 , \9324 , \9325 , \9326 , \9327 , \9328 , \9329 , \9330 ,
         \9331 , \9332 , \9333 , \9334 , \9335 , \9336 , \9337 , \9338 , \9339 , \9340 ,
         \9341 , \9342 , \9343 , \9344 , \9345 , \9346 , \9347 , \9348 , \9349 , \9350 ,
         \9351 , \9352 , \9353 , \9354 , \9355 , \9356 , \9357 , \9358 , \9359 , \9360 ,
         \9361 , \9362 , \9363 , \9364 , \9365 , \9366 , \9367 , \9368 , \9369 , \9370 ,
         \9371 , \9372 , \9373 , \9374 , \9375 , \9376 , \9377 , \9378 , \9379 , \9380 ,
         \9381 , \9382 , \9383 , \9384 , \9385 , \9386 , \9387 , \9388 , \9389 , \9390 ,
         \9391 , \9392 , \9393 , \9394 , \9395 , \9396 , \9397 , \9398 , \9399 , \9400 ,
         \9401 , \9402 , \9403 , \9404 , \9405 , \9406 , \9407 , \9408 , \9409 , \9410 ,
         \9411 , \9412 , \9413 , \9414 , \9415 , \9416 , \9417 , \9418 , \9419 , \9420 ,
         \9421 , \9422 , \9423 , \9424 , \9425 , \9426 , \9427 , \9428 , \9429 , \9430 ,
         \9431 , \9432 , \9433 , \9434 , \9435 , \9436 , \9437 , \9438 , \9439 , \9440 ,
         \9441 , \9442 , \9443 , \9444 , \9445 , \9446 , \9447 , \9448 , \9449 , \9450 ,
         \9451 , \9452 , \9453 , \9454 , \9455 , \9456 , \9457 , \9458 , \9459 , \9460 ,
         \9461 , \9462 , \9463 , \9464 , \9465 , \9466 , \9467 , \9468 , \9469 , \9470 ,
         \9471 , \9472 , \9473 , \9474 , \9475 , \9476 , \9477 , \9478 , \9479 , \9480 ,
         \9481 , \9482 , \9483 , \9484 , \9485 , \9486 , \9487 , \9488 , \9489 , \9490 ,
         \9491 , \9492 , \9493 , \9494 , \9495 , \9496 , \9497 , \9498 , \9499 , \9500 ,
         \9501 , \9502 , \9503 , \9504 , \9505 , \9506 , \9507 , \9508 , \9509 , \9510 ,
         \9511 , \9512 , \9513 , \9514 , \9515 , \9516 , \9517 , \9518 , \9519 , \9520 ,
         \9521 , \9522 , \9523 , \9524 , \9525 , \9526 , \9527 , \9528 , \9529 , \9530 ,
         \9531 , \9532 , \9533 , \9534 , \9535 , \9536 , \9537 , \9538 , \9539 , \9540 ,
         \9541 , \9542 , \9543 , \9544 , \9545 , \9546 , \9547 , \9548 , \9549 , \9550 ,
         \9551 , \9552 , \9553 , \9554 , \9555 , \9556 , \9557 , \9558 , \9559 , \9560 ,
         \9561 , \9562 , \9563 , \9564 , \9565 , \9566 , \9567 , \9568 , \9569 , \9570 ,
         \9571 , \9572 , \9573 , \9574 , \9575 , \9576 , \9577 , \9578 , \9579 , \9580 ,
         \9581 , \9582 , \9583 , \9584 , \9585 , \9586 , \9587 , \9588 , \9589 , \9590 ,
         \9591 , \9592 , \9593 , \9594 , \9595 , \9596 , \9597 , \9598 , \9599 , \9600 ,
         \9601 , \9602 , \9603 , \9604 , \9605 , \9606 , \9607 , \9608 , \9609 , \9610 ,
         \9611 , \9612 , \9613 , \9614 , \9615 , \9616 , \9617 , \9618 , \9619 , \9620 ,
         \9621 , \9622 , \9623 , \9624 , \9625 , \9626 , \9627 , \9628 , \9629 , \9630 ,
         \9631 , \9632 , \9633 , \9634 , \9635 , \9636 , \9637 , \9638 , \9639 , \9640 ,
         \9641 , \9642 , \9643 , \9644 , \9645 , \9646 , \9647 , \9648 , \9649 , \9650 ,
         \9651 , \9652 , \9653 , \9654 , \9655 , \9656 , \9657 , \9658 , \9659 , \9660 ,
         \9661 , \9662 , \9663 , \9664 , \9665 , \9666 , \9667 , \9668 , \9669 , \9670 ,
         \9671 , \9672 , \9673 , \9674 , \9675 , \9676 , \9677 , \9678 , \9679 , \9680 ,
         \9681 , \9682 , \9683 , \9684 , \9685 , \9686 , \9687 , \9688 , \9689 , \9690 ,
         \9691 , \9692 , \9693 , \9694 , \9695 , \9696 , \9697 , \9698 , \9699 , \9700 ,
         \9701 , \9702 , \9703 , \9704 , \9705 , \9706 , \9707 , \9708 , \9709 , \9710 ,
         \9711 , \9712 , \9713 , \9714 , \9715 , \9716 , \9717 , \9718 , \9719 , \9720 ,
         \9721 , \9722 , \9723 , \9724 , \9725 , \9726 , \9727 , \9728 , \9729 , \9730 ,
         \9731 , \9732 , \9733 , \9734 , \9735 , \9736 , \9737 , \9738 , \9739 , \9740 ,
         \9741 , \9742 , \9743 , \9744 , \9745 , \9746 , \9747 , \9748 , \9749 , \9750 ,
         \9751 , \9752 , \9753 , \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 ,
         \9761 , \9762 , \9763 , \9764 , \9765 , \9766 , \9767 , \9768 , \9769 , \9770 ,
         \9771 , \9772 , \9773 , \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 ,
         \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 ,
         \9791 , \9792 , \9793 , \9794 , \9795 , \9796 , \9797 , \9798 , \9799 , \9800 ,
         \9801 , \9802 , \9803 , \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 ,
         \9811 , \9812 , \9813 , \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 ,
         \9821 , \9822 , \9823 , \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 ,
         \9831 , \9832 , \9833 , \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 ,
         \9841 , \9842 , \9843 , \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 ,
         \9851 , \9852 , \9853 , \9854 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 ,
         \9861 , \9862 , \9863 , \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 ,
         \9871 , \9872 , \9873 , \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 ,
         \9881 , \9882 , \9883 , \9884 , \9885 , \9886 , \9887 , \9888 , \9889 , \9890 ,
         \9891 , \9892 , \9893 , \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 ,
         \9901 , \9902 , \9903 , \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 ,
         \9911 , \9912 , \9913 , \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 ,
         \9921 , \9922 , \9923 , \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 ,
         \9931 , \9932 , \9933 , \9934 , \9935 , \9936 , \9937 , \9938 , \9939 , \9940 ,
         \9941 , \9942 , \9943 , \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 ,
         \9951 , \9952 , \9953 , \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 ,
         \9961 , \9962 , \9963 , \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 ,
         \9971 , \9972 , \9973 , \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 ,
         \9981 , \9982 , \9983 , \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 ,
         \9991 , \9992 , \9993 , \9994 , \9995 , \9996 , \9997 , \9998 , \9999 , \10000 ,
         \10001 , \10002 , \10003 , \10004 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 ,
         \10011 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 ,
         \10021 , \10022 , \10023 , \10024 , \10025 , \10026 , \10027 , \10028 , \10029 , \10030 ,
         \10031 , \10032 , \10033 , \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 ,
         \10041 , \10042 , \10043 , \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 ,
         \10051 , \10052 , \10053 , \10054 , \10055 , \10056 , \10057 , \10058 , \10059 , \10060 ,
         \10061 , \10062 , \10063 , \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 ,
         \10071 , \10072 , \10073 , \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080 ,
         \10081 , \10082 , \10083 , \10084 , \10085 , \10086 , \10087 , \10088 , \10089 , \10090 ,
         \10091 , \10092 , \10093 , \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 ,
         \10101 , \10102 , \10103 , \10104 , \10105 , \10106 , \10107 , \10108 , \10109 , \10110 ,
         \10111 , \10112 , \10113 , \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 ,
         \10121 , \10122 , \10123 , \10124 , \10125 , \10126 , \10127 , \10128 , \10129 , \10130 ,
         \10131 , \10132 , \10133 , \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 ,
         \10141 , \10142 , \10143 , \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 ,
         \10151 , \10152 , \10153 , \10154 , \10155 , \10156 , \10157 , \10158 , \10159 , \10160 ,
         \10161 , \10162 , \10163 , \10164 , \10165 , \10166 , \10167 , \10168 , \10169 , \10170 ,
         \10171 , \10172 , \10173 , \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 ,
         \10181 , \10182 , \10183 , \10184 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 ,
         \10191 , \10192 , \10193 , \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 ,
         \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10207 , \10208 , \10209 , \10210 ,
         \10211 , \10212 , \10213 , \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 ,
         \10221 , \10222 , \10223 , \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 ,
         \10231 , \10232 , \10233 , \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 ,
         \10241 , \10242 , \10243 , \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 ,
         \10251 , \10252 , \10253 , \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 ,
         \10261 , \10262 , \10263 , \10264 , \10265 , \10266 , \10267 , \10268 , \10269 , \10270 ,
         \10271 , \10272 , \10273 , \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 ,
         \10281 , \10282 , \10283 , \10284 , \10285 , \10286 , \10287 , \10288 , \10289 , \10290 ,
         \10291 , \10292 , \10293 , \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 ,
         \10301 , \10302 , \10303 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 ,
         \10311 , \10312 , \10313 , \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 ,
         \10321 , \10322 , \10323 , \10324 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 ,
         \10331 , \10332 , \10333 , \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 ,
         \10341 , \10342 , \10343 , \10344 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 ,
         \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 ,
         \10361 , \10362 , \10363 , \10364 , \10365 , \10366 , \10367 , \10368 , \10369 , \10370 ,
         \10371 , \10372 , \10373 , \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 ,
         \10381 , \10382 , \10383 , \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 ,
         \10391 , \10392 , \10393 , \10394 , \10395 , \10396 , \10397 , \10398 , \10399 , \10400 ,
         \10401 , \10402 , \10403 , \10404 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 ,
         \10411 , \10412 , \10413 , \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 ,
         \10421 , \10422 , \10423 , \10424 , \10425 , \10426 , \10427 , \10428 , \10429 , \10430 ,
         \10431 , \10432 , \10433 , \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 ,
         \10441 , \10442 , \10443 , \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 ,
         \10451 , \10452 , \10453 , \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 ,
         \10461 , \10462 , \10463 , \10464 , \10465 , \10466 , \10467 , \10468 , \10469 , \10470 ,
         \10471 , \10472 , \10473 , \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 ,
         \10481 , \10482 , \10483 , \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 ,
         \10491 , \10492 , \10493 , \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 ,
         \10501 , \10502 , \10503 , \10504 , \10505 , \10506 , \10507 , \10508 , \10509 , \10510 ,
         \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 ,
         \10521 , \10522 , \10523 , \10524 , \10525 , \10526 , \10527 , \10528 , \10529 , \10530 ,
         \10531 , \10532 , \10533 , \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 ,
         \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 ,
         \10551 , \10552 , \10553 , \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 ,
         \10561 , \10562 , \10563 , \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 ,
         \10571 , \10572 , \10573 , \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 ,
         \10581 , \10582 , \10583 , \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 ,
         \10591 , \10592 , \10593 , \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 ,
         \10601 , \10602 , \10603 , \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610 ,
         \10611 , \10612 , \10613 , \10614 , \10615 , \10616 , \10617 , \10618 , \10619 , \10620 ,
         \10621 , \10622 , \10623 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 ,
         \10631 , \10632 , \10633 , \10634 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 ,
         \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 ,
         \10651 , \10652 , \10653 , \10654 , \10655 , \10656 , \10657 , \10658 , \10659 , \10660 ,
         \10661 , \10662 , \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 ,
         \10671 , \10672 , \10673 , \10674 , \10675 , \10676 , \10677 , \10678 , \10679 , \10680 ,
         \10681 , \10682 , \10683 , \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 ,
         \10691 , \10692 , \10693 , \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 ,
         \10701 , \10702 , \10703 , \10704 , \10705 , \10706 , \10707 , \10708 , \10709 , \10710 ,
         \10711 , \10712 , \10713 , \10714 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 ,
         \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 ,
         \10731 , \10732 , \10733 , \10734 , \10735 , \10736 , \10737 , \10738 , \10739 , \10740 ,
         \10741 , \10742 , \10743 , \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750 ,
         \10751 , \10752 , \10753 , \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 ,
         \10761 , \10762 , \10763 , \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 ,
         \10771 , \10772 , \10773 , \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 ,
         \10781 , \10782 , \10783 , \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 ,
         \10791 , \10792 , \10793 , \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 ,
         \10801 , \10802 , \10803 , \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 ,
         \10811 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 ,
         \10821 , \10822 , \10823 , \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 ,
         \10831 , \10832 , \10833 , \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 ,
         \10841 , \10842 , \10843 , \10844 , \10845 , \10846 , \10847 , \10848 , \10849 , \10850 ,
         \10851 , \10852 , \10853 , \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 ,
         \10861 , \10862 , \10863 , \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 ,
         \10871 , \10872 , \10873 , \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 ,
         \10881 , \10882 , \10883 , \10884 , \10885 , \10886 , \10887 , \10888 , \10889 , \10890 ,
         \10891 , \10892 , \10893 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 ,
         \10901 , \10902 , \10903 , \10904 , \10905 , \10906 , \10907 , \10908 , \10909 , \10910 ,
         \10911 , \10912 , \10913 , \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 ,
         \10921 , \10922 , \10923 , \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 ,
         \10931 , \10932 , \10933 , \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 ,
         \10941 , \10942 , \10943 , \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 ,
         \10951 , \10952 , \10953 , \10954 , \10955 , \10956 , \10957 , \10958 , \10959 , \10960 ,
         \10961 , \10962 , \10963 , \10964 , \10965 , \10966 , \10967 , \10968 , \10969 , \10970 ,
         \10971 , \10972 , \10973 , \10974 , \10975 , \10976 , \10977 , \10978 , \10979 , \10980 ,
         \10981 , \10982 , \10983 , \10984 , \10985 , \10986 , \10987 , \10988 , \10989 , \10990 ,
         \10991 , \10992 , \10993 , \10994 , \10995 , \10996 , \10997 , \10998 , \10999 , \11000 ,
         \11001 , \11002 , \11003 , \11004 , \11005 , \11006 , \11007 , \11008 , \11009 , \11010 ,
         \11011 , \11012 , \11013 , \11014 , \11015 , \11016 , \11017 , \11018 , \11019 , \11020 ,
         \11021 , \11022 , \11023 , \11024 , \11025 , \11026 , \11027 , \11028 , \11029 , \11030 ,
         \11031 , \11032 , \11033 , \11034 , \11035 , \11036 , \11037 , \11038 , \11039 , \11040 ,
         \11041 , \11042 , \11043 , \11044 , \11045 , \11046 , \11047 , \11048 , \11049 , \11050 ,
         \11051 , \11052 , \11053 , \11054 , \11055 , \11056 , \11057 , \11058 , \11059 , \11060 ,
         \11061 , \11062 , \11063 , \11064 , \11065 , \11066 , \11067 , \11068 , \11069 , \11070 ,
         \11071 , \11072 , \11073 , \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 ,
         \11081 , \11082 , \11083 , \11084 , \11085 , \11086 , \11087 , \11088 , \11089 , \11090 ,
         \11091 , \11092 , \11093 , \11094 , \11095 , \11096 , \11097 , \11098 , \11099 , \11100 ,
         \11101 , \11102 , \11103 , \11104 , \11105 , \11106 , \11107 , \11108 , \11109 , \11110 ,
         \11111 , \11112 , \11113 , \11114 , \11115 , \11116 , \11117 , \11118 , \11119 , \11120 ,
         \11121 , \11122 , \11123 , \11124 , \11125 , \11126 , \11127 , \11128 , \11129 , \11130 ,
         \11131 , \11132 , \11133 , \11134 , \11135 , \11136 , \11137 , \11138 , \11139 , \11140 ,
         \11141 , \11142 , \11143 , \11144 , \11145 , \11146 , \11147 , \11148 , \11149 , \11150 ,
         \11151 , \11152 , \11153 , \11154 , \11155 , \11156 , \11157 , \11158 , \11159 , \11160 ,
         \11161 , \11162 , \11163 , \11164 , \11165 , \11166 , \11167 , \11168 , \11169 , \11170 ,
         \11171 , \11172 , \11173 , \11174 , \11175 , \11176 , \11177 , \11178 , \11179 , \11180 ,
         \11181 , \11182 , \11183 , \11184 , \11185 , \11186 , \11187 , \11188 , \11189 , \11190 ,
         \11191 , \11192 , \11193 , \11194 , \11195 , \11196 , \11197 , \11198 , \11199 , \11200 ,
         \11201 , \11202 , \11203 , \11204 , \11205 , \11206 , \11207 , \11208 , \11209 , \11210 ,
         \11211 , \11212 , \11213 , \11214 , \11215 , \11216 , \11217 , \11218 , \11219 , \11220 ,
         \11221 , \11222 , \11223 , \11224 , \11225 , \11226 , \11227 , \11228 , \11229 , \11230 ,
         \11231 , \11232 , \11233 , \11234 , \11235 , \11236 , \11237 , \11238 , \11239 , \11240 ,
         \11241 , \11242 , \11243 , \11244 , \11245 , \11246 , \11247 , \11248 , \11249 , \11250 ,
         \11251 , \11252 , \11253 , \11254 , \11255 , \11256 , \11257 , \11258 , \11259 , \11260 ,
         \11261 , \11262 , \11263 , \11264 , \11265 , \11266 , \11267 , \11268 , \11269 , \11270 ,
         \11271 , \11272 , \11273 , \11274 , \11275 , \11276 , \11277 , \11278 , \11279 , \11280 ,
         \11281 , \11282 , \11283 , \11284 , \11285 , \11286 , \11287 , \11288 , \11289 , \11290 ,
         \11291 , \11292 , \11293 , \11294 , \11295 , \11296 , \11297 , \11298 , \11299 , \11300 ,
         \11301 , \11302 , \11303 , \11304 , \11305 , \11306 , \11307 , \11308 , \11309 , \11310 ,
         \11311 , \11312 , \11313 , \11314 , \11315 , \11316 , \11317 , \11318 , \11319 , \11320 ,
         \11321 , \11322 , \11323 , \11324 , \11325 , \11326 , \11327 , \11328 , \11329 , \11330 ,
         \11331 , \11332 , \11333 , \11334 , \11335 , \11336 , \11337 , \11338 , \11339 , \11340 ,
         \11341 , \11342 , \11343 , \11344 , \11345 , \11346 , \11347 , \11348 , \11349 , \11350 ,
         \11351 , \11352 , \11353 , \11354 , \11355 , \11356 , \11357 , \11358 , \11359 , \11360 ,
         \11361 , \11362 , \11363 , \11364 , \11365 , \11366 , \11367 , \11368 , \11369 , \11370 ,
         \11371 , \11372 , \11373 , \11374 , \11375 , \11376 , \11377 , \11378 , \11379 , \11380 ,
         \11381 , \11382 , \11383 , \11384 , \11385 , \11386 , \11387 , \11388 , \11389 , \11390 ,
         \11391 , \11392 , \11393 , \11394 , \11395 , \11396 , \11397 , \11398 , \11399 , \11400 ,
         \11401 , \11402 , \11403 , \11404 , \11405 , \11406 , \11407 , \11408 , \11409 , \11410 ,
         \11411 , \11412 , \11413 , \11414 , \11415 , \11416 , \11417 , \11418 , \11419 , \11420 ,
         \11421 , \11422 , \11423 , \11424 , \11425 , \11426 , \11427 , \11428 , \11429 , \11430 ,
         \11431 , \11432 , \11433 , \11434 , \11435 , \11436 , \11437 , \11438 , \11439 , \11440 ,
         \11441 , \11442 , \11443 , \11444 , \11445 , \11446 , \11447 , \11448 , \11449 , \11450 ,
         \11451 , \11452 , \11453 , \11454 , \11455 , \11456 , \11457 , \11458 , \11459 , \11460 ,
         \11461 , \11462 , \11463 , \11464 , \11465 , \11466 , \11467 , \11468 , \11469 , \11470 ,
         \11471 , \11472 , \11473 , \11474 , \11475 , \11476 , \11477 , \11478 , \11479 , \11480 ,
         \11481 , \11482 , \11483 , \11484 , \11485 , \11486 , \11487 , \11488 , \11489 , \11490 ,
         \11491 , \11492 , \11493 , \11494 , \11495 , \11496 , \11497 , \11498 , \11499 , \11500 ,
         \11501 , \11502 , \11503 , \11504 , \11505 , \11506 , \11507 , \11508 , \11509 , \11510 ,
         \11511 , \11512 , \11513 , \11514 , \11515 , \11516 , \11517 , \11518 , \11519 , \11520 ,
         \11521 , \11522 , \11523 , \11524 , \11525 , \11526 , \11527 , \11528 , \11529 , \11530 ,
         \11531 , \11532 , \11533 , \11534 , \11535 , \11536 , \11537 , \11538 , \11539 , \11540 ,
         \11541 , \11542 , \11543 , \11544 , \11545 , \11546 , \11547 , \11548 , \11549 , \11550 ,
         \11551 , \11552 , \11553 , \11554 , \11555 , \11556 , \11557 , \11558 , \11559 , \11560 ,
         \11561 , \11562 , \11563 , \11564 , \11565 , \11566 , \11567 , \11568 , \11569 , \11570 ,
         \11571 , \11572 , \11573 , \11574 , \11575 , \11576 , \11577 , \11578 , \11579 , \11580 ,
         \11581 , \11582 , \11583 , \11584 , \11585 , \11586 , \11587 , \11588 , \11589 , \11590 ,
         \11591 , \11592 , \11593 , \11594 , \11595 , \11596 , \11597 , \11598 , \11599 , \11600 ,
         \11601 , \11602 , \11603 , \11604 , \11605 , \11606 , \11607 , \11608 , \11609 , \11610 ,
         \11611 , \11612 , \11613 , \11614 , \11615 , \11616 , \11617 , \11618 , \11619 , \11620 ,
         \11621 , \11622 , \11623 , \11624 , \11625 , \11626 , \11627 , \11628 , \11629 , \11630 ,
         \11631 , \11632 , \11633 , \11634 , \11635 , \11636 , \11637 , \11638 , \11639 , \11640 ,
         \11641 , \11642 , \11643 , \11644 , \11645 , \11646 , \11647 , \11648 , \11649 , \11650 ,
         \11651 , \11652 , \11653 , \11654 , \11655 , \11656 , \11657 , \11658 , \11659 , \11660 ,
         \11661 , \11662 , \11663 , \11664 , \11665 , \11666 , \11667 , \11668 , \11669 , \11670 ,
         \11671 , \11672 , \11673 , \11674 , \11675 , \11676 , \11677 , \11678 , \11679 , \11680 ,
         \11681 , \11682 , \11683 , \11684 , \11685 , \11686 , \11687 , \11688 , \11689 , \11690 ,
         \11691 , \11692 , \11693 , \11694 , \11695 , \11696 , \11697 , \11698 , \11699 , \11700 ,
         \11701 , \11702 , \11703 , \11704 , \11705 , \11706 , \11707 , \11708 , \11709 , \11710 ,
         \11711 , \11712 , \11713 , \11714 , \11715 , \11716 , \11717 , \11718 , \11719 , \11720 ,
         \11721 , \11722 , \11723 , \11724 , \11725 , \11726 , \11727 , \11728 , \11729 , \11730 ,
         \11731 , \11732 , \11733 , \11734 , \11735 , \11736 , \11737 , \11738 , \11739 , \11740 ,
         \11741 , \11742 , \11743 , \11744 , \11745 , \11746 , \11747 , \11748 , \11749 , \11750 ,
         \11751 , \11752 , \11753 , \11754 , \11755 , \11756 , \11757 , \11758 , \11759 , \11760 ,
         \11761 , \11762 , \11763 , \11764 , \11765 , \11766 , \11767 , \11768 , \11769 , \11770 ,
         \11771 , \11772 , \11773 , \11774 , \11775 , \11776 , \11777 , \11778 , \11779 , \11780 ,
         \11781 , \11782 , \11783 , \11784 , \11785 , \11786 , \11787 , \11788 , \11789 , \11790 ,
         \11791 , \11792 , \11793 , \11794 , \11795 , \11796 , \11797 , \11798 , \11799 , \11800 ,
         \11801 , \11802 , \11803 , \11804 , \11805 , \11806 , \11807 , \11808 , \11809 , \11810 ,
         \11811 , \11812 , \11813 , \11814 , \11815 , \11816 , \11817 , \11818 , \11819 , \11820 ,
         \11821 , \11822 , \11823 , \11824 , \11825 , \11826 , \11827 , \11828 , \11829 , \11830 ,
         \11831 , \11832 , \11833 , \11834 , \11835 , \11836 , \11837 , \11838 , \11839 , \11840 ,
         \11841 , \11842 , \11843 , \11844 , \11845 , \11846 , \11847 , \11848 , \11849 , \11850 ,
         \11851 , \11852 , \11853 , \11854 , \11855 , \11856 , \11857 , \11858 , \11859 , \11860 ,
         \11861 , \11862 , \11863 , \11864 , \11865 , \11866 , \11867 , \11868 , \11869 , \11870 ,
         \11871 , \11872 , \11873 , \11874 , \11875 , \11876 , \11877 , \11878 , \11879 , \11880 ,
         \11881 , \11882 , \11883 , \11884 , \11885 , \11886 , \11887 , \11888 , \11889 , \11890 ,
         \11891 , \11892 , \11893 , \11894 , \11895 , \11896 , \11897 , \11898 , \11899 , \11900 ,
         \11901 , \11902 , \11903 , \11904 , \11905 , \11906 , \11907 , \11908 , \11909 , \11910 ,
         \11911 , \11912 , \11913 , \11914 , \11915 , \11916 , \11917 , \11918 , \11919 , \11920 ,
         \11921 , \11922 , \11923 , \11924 , \11925 , \11926 , \11927 , \11928 , \11929 , \11930 ,
         \11931 , \11932 , \11933 , \11934 , \11935 , \11936 , \11937 , \11938 , \11939 , \11940 ,
         \11941 , \11942 , \11943 , \11944 , \11945 , \11946 , \11947 , \11948 , \11949 , \11950 ,
         \11951 , \11952 , \11953 , \11954 , \11955 , \11956 , \11957 , \11958 , \11959 , \11960 ,
         \11961 , \11962 , \11963 , \11964 , \11965 , \11966 , \11967 , \11968 , \11969 , \11970 ,
         \11971 , \11972 , \11973 , \11974 , \11975 , \11976 , \11977 , \11978 , \11979 , \11980 ,
         \11981 , \11982 , \11983 , \11984 , \11985 , \11986 , \11987 , \11988 , \11989 , \11990 ,
         \11991 , \11992 , \11993 , \11994 , \11995 , \11996 , \11997 , \11998 , \11999 , \12000 ,
         \12001 , \12002 , \12003 , \12004 , \12005 , \12006 , \12007 , \12008 , \12009 , \12010 ,
         \12011 , \12012 , \12013 , \12014 , \12015 , \12016 , \12017 , \12018 , \12019 , \12020 ,
         \12021 , \12022 , \12023 , \12024 , \12025 , \12026 , \12027 , \12028 , \12029 , \12030 ,
         \12031 , \12032 , \12033 , \12034 , \12035 , \12036 , \12037 , \12038 , \12039 , \12040 ,
         \12041 , \12042 , \12043 , \12044 , \12045 , \12046 , \12047 , \12048 , \12049 , \12050 ,
         \12051 , \12052 , \12053 , \12054 , \12055 , \12056 , \12057 , \12058 , \12059 , \12060 ,
         \12061 , \12062 , \12063 , \12064 , \12065 , \12066 , \12067 , \12068 , \12069 , \12070 ,
         \12071 , \12072 , \12073 , \12074 , \12075 , \12076 , \12077 , \12078 , \12079 , \12080 ,
         \12081 , \12082 , \12083 , \12084 , \12085 , \12086 , \12087 , \12088 , \12089 , \12090 ,
         \12091 , \12092 , \12093 , \12094 , \12095 , \12096 , \12097 , \12098 , \12099 , \12100 ,
         \12101 , \12102 , \12103 , \12104 , \12105 , \12106 , \12107 , \12108 , \12109 , \12110 ,
         \12111 , \12112 , \12113 , \12114 , \12115 , \12116 , \12117 , \12118 , \12119 , \12120 ,
         \12121 , \12122 , \12123 , \12124 , \12125 , \12126 , \12127 , \12128 , \12129 , \12130 ,
         \12131 , \12132 , \12133 , \12134 , \12135 , \12136 , \12137 , \12138 , \12139 , \12140 ,
         \12141 , \12142 , \12143 , \12144 , \12145 , \12146 , \12147 , \12148 , \12149 , \12150 ,
         \12151 , \12152 , \12153 , \12154 , \12155 , \12156 , \12157 , \12158 , \12159 , \12160 ,
         \12161 , \12162 , \12163 , \12164 , \12165 , \12166 , \12167 , \12168 , \12169 , \12170 ,
         \12171 , \12172 , \12173 , \12174 , \12175 , \12176 , \12177 , \12178 , \12179 , \12180 ,
         \12181 , \12182 , \12183 , \12184 , \12185 , \12186 , \12187 , \12188 , \12189 , \12190 ,
         \12191 , \12192 , \12193 , \12194 , \12195 , \12196 , \12197 , \12198 , \12199 , \12200 ,
         \12201 , \12202 , \12203 , \12204 , \12205 , \12206 , \12207 , \12208 , \12209 , \12210 ,
         \12211 , \12212 , \12213 , \12214 , \12215 , \12216 , \12217 , \12218 , \12219 , \12220 ,
         \12221 , \12222 , \12223 , \12224 , \12225 , \12226 , \12227 , \12228 , \12229 , \12230 ,
         \12231 , \12232 , \12233 , \12234 , \12235 , \12236 , \12237 , \12238 , \12239 , \12240 ,
         \12241 , \12242 , \12243 , \12244 , \12245 , \12246 , \12247 , \12248 , \12249 , \12250 ,
         \12251 , \12252 , \12253 , \12254 , \12255 , \12256 , \12257 , \12258 , \12259 , \12260 ,
         \12261 , \12262 , \12263 , \12264 , \12265 , \12266 , \12267 , \12268 , \12269 , \12270 ,
         \12271 , \12272 , \12273 , \12274 , \12275 , \12276 , \12277 , \12278 , \12279 , \12280 ,
         \12281 , \12282 , \12283 , \12284 , \12285 , \12286 , \12287 , \12288 , \12289 , \12290 ,
         \12291 , \12292 , \12293 , \12294 , \12295 , \12296 , \12297 , \12298 , \12299 , \12300 ,
         \12301 , \12302 , \12303 , \12304 , \12305 , \12306 , \12307 , \12308 , \12309 , \12310 ,
         \12311 , \12312 , \12313 , \12314 , \12315 , \12316 , \12317 , \12318 , \12319 , \12320 ,
         \12321 , \12322 , \12323 , \12324 , \12325 , \12326 , \12327 , \12328 , \12329 , \12330 ,
         \12331 , \12332 , \12333 , \12334 , \12335 , \12336 , \12337 , \12338 , \12339 , \12340 ,
         \12341 , \12342 , \12343 , \12344 , \12345 , \12346 , \12347 , \12348 , \12349 , \12350 ,
         \12351 , \12352 , \12353 , \12354 , \12355 , \12356 , \12357 , \12358 , \12359 , \12360 ,
         \12361 , \12362 , \12363 , \12364 , \12365 , \12366 , \12367 , \12368 , \12369 , \12370 ,
         \12371 , \12372 , \12373 , \12374 , \12375 , \12376 , \12377 , \12378 , \12379 , \12380 ,
         \12381 , \12382 , \12383 , \12384 , \12385 , \12386 , \12387 , \12388 , \12389 , \12390 ,
         \12391 , \12392 , \12393 , \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 ,
         \12401 , \12402 , \12403 , \12404 , \12405 , \12406 , \12407 , \12408 , \12409 , \12410 ,
         \12411 , \12412 , \12413 , \12414 , \12415 , \12416 , \12417 , \12418 , \12419 , \12420 ,
         \12421 , \12422 , \12423 , \12424 , \12425 , \12426 , \12427 , \12428 , \12429 , \12430 ,
         \12431 , \12432 , \12433 , \12434 , \12435 , \12436 , \12437 , \12438 , \12439 , \12440 ,
         \12441 , \12442 , \12443 , \12444 , \12445 , \12446 , \12447 , \12448 , \12449 , \12450 ,
         \12451 , \12452 , \12453 , \12454 , \12455 , \12456 , \12457 , \12458 , \12459 , \12460 ,
         \12461 , \12462 , \12463 , \12464 , \12465 , \12466 , \12467 , \12468 , \12469 , \12470 ,
         \12471 , \12472 , \12473 , \12474 , \12475 , \12476 , \12477 , \12478 , \12479 , \12480 ,
         \12481 , \12482 , \12483 , \12484 , \12485 , \12486 , \12487 , \12488 , \12489 , \12490 ,
         \12491 , \12492 , \12493 , \12494 , \12495 , \12496 , \12497 , \12498 , \12499 , \12500 ,
         \12501 , \12502 , \12503 , \12504 , \12505 , \12506 , \12507 , \12508 , \12509 , \12510 ,
         \12511 , \12512 , \12513 , \12514 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 ,
         \12521 , \12522 , \12523 , \12524 , \12525 , \12526 , \12527 , \12528 , \12529 , \12530 ,
         \12531 , \12532 , \12533 , \12534 , \12535 , \12536 , \12537 , \12538 , \12539 , \12540 ,
         \12541 , \12542 , \12543 , \12544 , \12545 , \12546 , \12547 , \12548 , \12549 , \12550 ,
         \12551 , \12552 , \12553 , \12554 , \12555 , \12556 , \12557 , \12558 , \12559 , \12560 ,
         \12561 , \12562 , \12563 , \12564 , \12565 , \12566 , \12567 , \12568 , \12569 , \12570 ,
         \12571 , \12572 , \12573 , \12574 , \12575 , \12576 , \12577 , \12578 , \12579 , \12580 ,
         \12581 , \12582 , \12583 , \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 ,
         \12591 , \12592 , \12593 , \12594 , \12595 , \12596 , \12597 , \12598 , \12599 , \12600 ,
         \12601 , \12602 , \12603 , \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12610 ,
         \12611 , \12612 , \12613 , \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 ,
         \12621 , \12622 , \12623 , \12624 , \12625 , \12626 , \12627 , \12628 , \12629 , \12630 ,
         \12631 , \12632 , \12633 , \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 ,
         \12641 , \12642 , \12643 , \12644 , \12645 , \12646 , \12647 , \12648 , \12649 , \12650 ,
         \12651 , \12652 , \12653 , \12654 , \12655 , \12656 , \12657 , \12658 , \12659 , \12660 ,
         \12661 , \12662 , \12663 , \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 ,
         \12671 , \12672 , \12673 , \12674 , \12675 , \12676 , \12677 , \12678 , \12679 , \12680 ,
         \12681 , \12682 , \12683 , \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 ,
         \12691 , \12692 , \12693 , \12694 , \12695 , \12696 , \12697 , \12698 , \12699 , \12700 ,
         \12701 , \12702 , \12703 , \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 ,
         \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 ,
         \12721 , \12722 , \12723 , \12724 , \12725 , \12726 , \12727 , \12728 , \12729 , \12730 ,
         \12731 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 ,
         \12741 , \12742 , \12743 , \12744 , \12745 , \12746 , \12747 , \12748 , \12749 , \12750 ,
         \12751 , \12752 , \12753 , \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 ,
         \12761 , \12762 , \12763 , \12764 , \12765 , \12766 , \12767 , \12768 , \12769 , \12770 ,
         \12771 , \12772 , \12773 , \12774 , \12775 , \12776 , \12777 , \12778 , \12779 , \12780 ,
         \12781 , \12782 , \12783 , \12784 , \12785 , \12786 , \12787 , \12788 , \12789 , \12790 ,
         \12791 , \12792 , \12793 , \12794 , \12795 , \12796 , \12797 , \12798 , \12799 , \12800 ,
         \12801 , \12802 , \12803 , \12804 , \12805 , \12806 , \12807 , \12808 , \12809 , \12810 ,
         \12811 , \12812 , \12813 , \12814 , \12815 , \12816 , \12817 , \12818 , \12819 , \12820 ,
         \12821 , \12822 , \12823 , \12824 , \12825 , \12826 , \12827 , \12828 , \12829 , \12830 ,
         \12831 , \12832 , \12833 , \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 ,
         \12841 , \12842 , \12843 , \12844 , \12845 , \12846 , \12847 , \12848 , \12849 , \12850 ,
         \12851 , \12852 , \12853 , \12854 , \12855 , \12856 , \12857 , \12858 , \12859 , \12860 ,
         \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 ,
         \12871 , \12872 , \12873 , \12874 , \12875 , \12876 , \12877 , \12878 , \12879 , \12880 ,
         \12881 , \12882 , \12883 , \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 ,
         \12891 , \12892 , \12893 , \12894 , \12895 , \12896 , \12897 , \12898 , \12899 , \12900 ,
         \12901 , \12902 , \12903 , \12904 , \12905 , \12906 , \12907 , \12908 , \12909 , \12910 ,
         \12911 , \12912 , \12913 , \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 ,
         \12921 , \12922 , \12923 , \12924 , \12925 , \12926 , \12927 , \12928 , \12929 , \12930 ,
         \12931 , \12932 , \12933 , \12934 , \12935 , \12936 , \12937 , \12938 , \12939 , \12940 ,
         \12941 , \12942 , \12943 , \12944 , \12945 , \12946 , \12947 , \12948 , \12949 , \12950 ,
         \12951 , \12952 , \12953 , \12954 , \12955 , \12956 , \12957 , \12958 , \12959 , \12960 ,
         \12961 , \12962 , \12963 , \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 ,
         \12971 , \12972 , \12973 , \12974 , \12975 , \12976 , \12977 , \12978 , \12979 , \12980 ,
         \12981 , \12982 , \12983 , \12984 , \12985 , \12986 , \12987 , \12988 , \12989 , \12990 ,
         \12991 , \12992 , \12993 , \12994 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 ,
         \13001 , \13002 , \13003 , \13004 , \13005 , \13006 , \13007 , \13008 , \13009 , \13010 ,
         \13011 , \13012 , \13013 , \13014 , \13015 , \13016 , \13017 , \13018 , \13019 , \13020 ,
         \13021 , \13022 , \13023 , \13024 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 ,
         \13031 , \13032 , \13033 , \13034 , \13035 , \13036 , \13037 , \13038 , \13039 , \13040 ,
         \13041 , \13042 , \13043 , \13044 , \13045 , \13046 , \13047 , \13048 , \13049 , \13050 ,
         \13051 , \13052 , \13053 , \13054 , \13055 , \13056 , \13057 , \13058 , \13059 , \13060 ,
         \13061 , \13062 , \13063 , \13064 , \13065 , \13066 , \13067 , \13068 , \13069 , \13070 ,
         \13071 , \13072 , \13073 , \13074 , \13075 , \13076 , \13077 , \13078 , \13079 , \13080 ,
         \13081 , \13082 , \13083 , \13084 , \13085 , \13086 , \13087 , \13088 , \13089 , \13090 ,
         \13091 , \13092 , \13093 , \13094 , \13095 , \13096 , \13097 , \13098 , \13099 , \13100 ,
         \13101 , \13102 , \13103 , \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 ,
         \13111 , \13112 , \13113 , \13114 , \13115 , \13116 , \13117 , \13118 , \13119 , \13120 ,
         \13121 , \13122 , \13123 , \13124 , \13125 , \13126 , \13127 , \13128 , \13129 , \13130 ,
         \13131 , \13132 , \13133 , \13134 , \13135 , \13136 , \13137 , \13138 , \13139 , \13140 ,
         \13141 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 ,
         \13151 , \13152 , \13153 , \13154 , \13155 , \13156 , \13157 , \13158 , \13159 , \13160 ,
         \13161 , \13162 , \13163 , \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 ,
         \13171 , \13172 , \13173 , \13174 , \13175 , \13176 , \13177 , \13178 , \13179 , \13180 ,
         \13181 , \13182 , \13183 , \13184 , \13185 , \13186 , \13187 , \13188 , \13189 , \13190 ,
         \13191 , \13192 , \13193 , \13194 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 ,
         \13201 , \13202 , \13203 , \13204 , \13205 , \13206 , \13207 , \13208 , \13209 , \13210 ,
         \13211 , \13212 , \13213 , \13214 , \13215 , \13216 , \13217 , \13218 , \13219 , \13220 ,
         \13221 , \13222 , \13223 , \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 ,
         \13231 , \13232 , \13233 , \13234 , \13235 , \13236 , \13237 , \13238 , \13239 , \13240 ,
         \13241 , \13242 , \13243 , \13244 , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 ,
         \13251 , \13252 , \13253 , \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 ,
         \13261 , \13262 , \13263 , \13264 , \13265 , \13266 , \13267 , \13268 , \13269 , \13270 ,
         \13271 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 ,
         \13281 , \13282 , \13283 , \13284 , \13285 , \13286 , \13287 , \13288 , \13289 , \13290 ,
         \13291 , \13292 , \13293 , \13294 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 ,
         \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 ,
         \13311 , \13312 , \13313 , \13314 , \13315 , \13316 , \13317 , \13318 , \13319 , \13320 ,
         \13321 , \13322 , \13323 , \13324 , \13325 , \13326 , \13327 , \13328 , \13329 , \13330 ,
         \13331 , \13332 , \13333 , \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 ,
         \13341 , \13342 , \13343 , \13344 , \13345 , \13346 , \13347 , \13348 , \13349 , \13350 ,
         \13351 , \13352 , \13353 , \13354 , \13355 , \13356 , \13357 , \13358 , \13359 , \13360 ,
         \13361 , \13362 , \13363 , \13364 , \13365 , \13366 , \13367 , \13368 , \13369 , \13370 ,
         \13371 , \13372 , \13373 , \13374 , \13375 , \13376 , \13377 , \13378 , \13379 , \13380 ,
         \13381 , \13382 , \13383 , \13384 , \13385 , \13386 , \13387 , \13388 , \13389 , \13390 ,
         \13391 , \13392 , \13393 , \13394 , \13395 , \13396 , \13397 , \13398 , \13399 , \13400 ,
         \13401 , \13402 , \13403 , \13404 , \13405 , \13406 , \13407 , \13408 , \13409 , \13410 ,
         \13411 , \13412 , \13413 , \13414 , \13415 , \13416 , \13417 , \13418 , \13419 , \13420 ,
         \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430 ,
         \13431 , \13432 , \13433 , \13434 , \13435 , \13436 , \13437 , \13438 , \13439 , \13440 ,
         \13441 , \13442 , \13443 , \13444 , \13445 , \13446 , \13447 , \13448 , \13449 , \13450 ,
         \13451 , \13452 , \13453 , \13454 , \13455 , \13456 , \13457 , \13458 , \13459 , \13460 ,
         \13461 , \13462 , \13463 , \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 ,
         \13471 , \13472 , \13473 , \13474 , \13475 , \13476 , \13477 , \13478 , \13479 , \13480 ,
         \13481 , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 ,
         \13491 , \13492 , \13493 , \13494 , \13495 , \13496 , \13497 , \13498 , \13499 , \13500 ,
         \13501 , \13502 , \13503 , \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 ,
         \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 ,
         \13521 , \13522 , \13523 , \13524 , \13525 , \13526 , \13527 , \13528 , \13529 , \13530 ,
         \13531 , \13532 , \13533 , \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 ,
         \13541 , \13542 , \13543 , \13544 , \13545 , \13546 , \13547 , \13548 , \13549 , \13550 ,
         \13551 , \13552 , \13553 , \13554 , \13555 , \13556 , \13557 , \13558 , \13559 , \13560 ,
         \13561 , \13562 , \13563 , \13564 , \13565 , \13566 , \13567 , \13568 , \13569 , \13570 ,
         \13571 , \13572 , \13573 , \13574 , \13575 , \13576 , \13577 , \13578 , \13579 , \13580 ,
         \13581 , \13582 , \13583 , \13584 , \13585 , \13586 , \13587 , \13588 , \13589 , \13590 ,
         \13591 , \13592 , \13593 , \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 ,
         \13601 , \13602 , \13603 , \13604 , \13605 , \13606 , \13607 , \13608 , \13609 , \13610 ,
         \13611 , \13612 , \13613 , \13614 , \13615 , \13616 , \13617 , \13618 , \13619 , \13620 ,
         \13621 , \13622 , \13623 , \13624 , \13625 , \13626 , \13627 , \13628 , \13629 , \13630 ,
         \13631 , \13632 , \13633 , \13634 , \13635 , \13636 , \13637 , \13638 , \13639 , \13640 ,
         \13641 , \13642 , \13643 , \13644 , \13645 , \13646 , \13647 , \13648 , \13649 , \13650 ,
         \13651 , \13652 , \13653 , \13654 , \13655 , \13656 , \13657 , \13658 , \13659 , \13660 ,
         \13661 , \13662 , \13663 , \13664 , \13665 , \13666 , \13667 , \13668 , \13669 , \13670 ,
         \13671 , \13672 , \13673 , \13674 , \13675 , \13676 , \13677 , \13678 , \13679 , \13680 ,
         \13681 , \13682 , \13683 , \13684 , \13685 , \13686 , \13687 , \13688 , \13689 , \13690 ,
         \13691 , \13692 , \13693 , \13694 , \13695 , \13696 , \13697 , \13698 , \13699 , \13700 ,
         \13701 , \13702 , \13703 , \13704 , \13705 , \13706 , \13707 , \13708 , \13709 , \13710 ,
         \13711 , \13712 , \13713 , \13714 , \13715 , \13716 , \13717 , \13718 , \13719 , \13720 ,
         \13721 , \13722 , \13723 , \13724 , \13725 , \13726 , \13727 , \13728 , \13729 , \13730 ,
         \13731 , \13732 , \13733 , \13734 , \13735 , \13736 , \13737 , \13738 , \13739 , \13740 ,
         \13741 , \13742 , \13743 , \13744 , \13745 , \13746 , \13747 , \13748 , \13749 , \13750 ,
         \13751 , \13752 , \13753 , \13754 , \13755 , \13756 , \13757 , \13758 , \13759 , \13760 ,
         \13761 , \13762 , \13763 , \13764 , \13765 , \13766 , \13767 , \13768 , \13769 , \13770 ,
         \13771 , \13772 , \13773 , \13774 , \13775 , \13776 , \13777 , \13778 , \13779 , \13780 ,
         \13781 , \13782 , \13783 , \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 ,
         \13791 , \13792 , \13793 , \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 ,
         \13801 , \13802 , \13803 , \13804 , \13805 , \13806 , \13807 , \13808 , \13809 , \13810 ,
         \13811 , \13812 , \13813 , \13814 , \13815 , \13816 , \13817 , \13818 , \13819 , \13820 ,
         \13821 , \13822 , \13823 , \13824 , \13825 , \13826 , \13827 , \13828 , \13829 , \13830 ,
         \13831 , \13832 , \13833 , \13834 , \13835 , \13836 , \13837 , \13838 , \13839 , \13840 ,
         \13841 , \13842 , \13843 , \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 ,
         \13851 , \13852 , \13853 , \13854 , \13855 , \13856 , \13857 , \13858 , \13859 , \13860 ,
         \13861 , \13862 , \13863 , \13864 , \13865 , \13866 , \13867 , \13868 , \13869 , \13870 ,
         \13871 , \13872 , \13873 , \13874 , \13875 , \13876 , \13877 , \13878 , \13879 , \13880 ,
         \13881 , \13882 , \13883 , \13884 , \13885 , \13886 , \13887 , \13888 , \13889 , \13890 ,
         \13891 , \13892 , \13893 , \13894 , \13895 , \13896 , \13897 , \13898 , \13899 , \13900 ,
         \13901 , \13902 , \13903 , \13904 , \13905 , \13906 , \13907 , \13908 , \13909 , \13910 ,
         \13911 , \13912 , \13913 , \13914 , \13915 , \13916 , \13917 , \13918 , \13919 , \13920 ,
         \13921 , \13922 , \13923 , \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 ,
         \13931 , \13932 , \13933 , \13934 , \13935 , \13936 , \13937 , \13938 , \13939 , \13940 ,
         \13941 , \13942 , \13943 , \13944 , \13945 , \13946 , \13947 , \13948 , \13949 , \13950 ,
         \13951 , \13952 , \13953 , \13954 , \13955 , \13956 , \13957 , \13958 , \13959 , \13960 ,
         \13961 , \13962 , \13963 , \13964 , \13965 , \13966 , \13967 , \13968 , \13969 , \13970 ,
         \13971 , \13972 , \13973 , \13974 , \13975 , \13976 , \13977 , \13978 , \13979 , \13980 ,
         \13981 , \13982 , \13983 , \13984 , \13985 , \13986 , \13987 , \13988 , \13989 , \13990 ,
         \13991 , \13992 , \13993 , \13994 , \13995 , \13996 , \13997 , \13998 , \13999 , \14000 ,
         \14001 , \14002 , \14003 , \14004 , \14005 , \14006 , \14007 , \14008 , \14009 , \14010 ,
         \14011 , \14012 , \14013 , \14014 , \14015 , \14016 , \14017 , \14018 , \14019 , \14020 ,
         \14021 , \14022 , \14023 , \14024 , \14025 , \14026 , \14027 , \14028 , \14029 , \14030 ,
         \14031 , \14032 , \14033 , \14034 , \14035 , \14036 , \14037 , \14038 , \14039 , \14040 ,
         \14041 , \14042 , \14043 , \14044 , \14045 , \14046 , \14047 , \14048 , \14049 , \14050 ,
         \14051 , \14052 , \14053 , \14054 , \14055 , \14056 , \14057 , \14058 , \14059 , \14060 ,
         \14061 , \14062 , \14063 , \14064 , \14065 , \14066 , \14067 , \14068 , \14069 , \14070 ,
         \14071 , \14072 , \14073 , \14074 , \14075 , \14076 , \14077 , \14078 , \14079 , \14080 ,
         \14081 , \14082 , \14083 , \14084 , \14085 , \14086 , \14087 , \14088 , \14089 , \14090 ,
         \14091 , \14092 , \14093 , \14094 , \14095 , \14096 , \14097 , \14098 , \14099 , \14100 ,
         \14101 , \14102 , \14103 , \14104 , \14105 , \14106 , \14107 , \14108 , \14109 , \14110 ,
         \14111 , \14112 , \14113 , \14114 , \14115 , \14116 , \14117 , \14118 , \14119 , \14120 ,
         \14121 , \14122 , \14123 , \14124 , \14125 , \14126 , \14127 , \14128 , \14129 , \14130 ,
         \14131 , \14132 , \14133 , \14134 , \14135 , \14136 , \14137 , \14138 , \14139 , \14140 ,
         \14141 , \14142 , \14143 , \14144 , \14145 , \14146 , \14147 , \14148 , \14149 , \14150 ,
         \14151 , \14152 , \14153 , \14154 , \14155 , \14156 , \14157 , \14158 , \14159 , \14160 ,
         \14161 , \14162 , \14163 , \14164 , \14165 , \14166 , \14167 , \14168 , \14169 , \14170 ,
         \14171 , \14172 , \14173 , \14174 , \14175 , \14176 , \14177 , \14178 , \14179 , \14180 ,
         \14181 , \14182 , \14183 , \14184 , \14185 , \14186 , \14187 , \14188 , \14189 , \14190 ,
         \14191 , \14192 , \14193 , \14194 , \14195 , \14196 , \14197 , \14198 , \14199 , \14200 ,
         \14201 , \14202 , \14203 , \14204 , \14205 , \14206 , \14207 , \14208 , \14209 , \14210 ,
         \14211 , \14212 , \14213 , \14214 , \14215 , \14216 , \14217 , \14218 , \14219 , \14220 ,
         \14221 , \14222 , \14223 , \14224 , \14225 , \14226 , \14227 , \14228 , \14229 , \14230 ,
         \14231 , \14232 , \14233 , \14234 , \14235 , \14236 , \14237 , \14238 , \14239 , \14240 ,
         \14241 , \14242 , \14243 , \14244 , \14245 , \14246 , \14247 , \14248 , \14249 , \14250 ,
         \14251 , \14252 , \14253 , \14254 , \14255 , \14256 , \14257 , \14258 , \14259 , \14260 ,
         \14261 , \14262 , \14263 , \14264 , \14265 , \14266 , \14267 , \14268 , \14269 , \14270 ,
         \14271 , \14272 , \14273 , \14274 , \14275 , \14276 , \14277 , \14278 , \14279 , \14280 ,
         \14281 , \14282 , \14283 , \14284 , \14285 , \14286 , \14287 , \14288 , \14289 , \14290 ,
         \14291 , \14292 , \14293 , \14294 , \14295 , \14296 , \14297 , \14298 , \14299 , \14300 ,
         \14301 , \14302 , \14303 , \14304 , \14305 , \14306 , \14307 , \14308 , \14309 , \14310 ,
         \14311 , \14312 , \14313 , \14314 , \14315 , \14316 , \14317 , \14318 , \14319 , \14320 ,
         \14321 , \14322 , \14323 , \14324 , \14325 , \14326 , \14327 , \14328 , \14329 , \14330 ,
         \14331 , \14332 , \14333 , \14334 , \14335 , \14336 , \14337 , \14338 , \14339 , \14340 ,
         \14341 , \14342 , \14343 , \14344 , \14345 , \14346 , \14347 , \14348 , \14349 , \14350 ,
         \14351 , \14352 , \14353 , \14354 , \14355 , \14356 , \14357 , \14358 , \14359 , \14360 ,
         \14361 , \14362 , \14363 , \14364 , \14365 , \14366 , \14367 , \14368 , \14369 , \14370 ,
         \14371 , \14372 , \14373 , \14374 , \14375 , \14376 , \14377 , \14378 , \14379 , \14380 ,
         \14381 , \14382 , \14383 , \14384 , \14385 , \14386 , \14387 , \14388 , \14389 , \14390 ,
         \14391 , \14392 , \14393 , \14394 , \14395 , \14396 , \14397 , \14398 , \14399 , \14400 ,
         \14401 , \14402 , \14403 , \14404 , \14405 , \14406 , \14407 , \14408 , \14409 , \14410 ,
         \14411 , \14412 , \14413 , \14414 , \14415 , \14416 , \14417 , \14418 , \14419 , \14420 ,
         \14421 , \14422 , \14423 , \14424 , \14425 , \14426 , \14427 , \14428 , \14429 , \14430 ,
         \14431 , \14432 , \14433 , \14434 , \14435 , \14436 , \14437 , \14438 , \14439 , \14440 ,
         \14441 , \14442 , \14443 , \14444 , \14445 , \14446 , \14447 , \14448 , \14449 , \14450 ,
         \14451 , \14452 , \14453 , \14454 , \14455 , \14456 , \14457 , \14458 , \14459 , \14460 ,
         \14461 , \14462 , \14463 , \14464 , \14465 , \14466 , \14467 , \14468 , \14469 , \14470 ,
         \14471 , \14472 , \14473 , \14474 , \14475 , \14476 , \14477 , \14478 , \14479 , \14480 ,
         \14481 , \14482 , \14483 , \14484 , \14485 , \14486 , \14487 , \14488 , \14489 , \14490 ,
         \14491 , \14492 , \14493 , \14494 , \14495 , \14496 , \14497 , \14498 , \14499 , \14500 ,
         \14501 , \14502 , \14503 , \14504 , \14505 , \14506 , \14507 , \14508 , \14509 , \14510 ,
         \14511 , \14512 , \14513 , \14514 , \14515 , \14516 , \14517 , \14518 , \14519 , \14520 ,
         \14521 , \14522 , \14523 , \14524 , \14525 , \14526 , \14527 , \14528 , \14529 , \14530 ,
         \14531 , \14532 , \14533 , \14534 , \14535 , \14536 , \14537 , \14538 , \14539 , \14540 ,
         \14541 , \14542 , \14543 , \14544 , \14545 , \14546 , \14547 , \14548 , \14549 , \14550 ,
         \14551 , \14552 , \14553 , \14554 , \14555 , \14556 , \14557 , \14558 , \14559 , \14560 ,
         \14561 , \14562 , \14563 , \14564 , \14565 , \14566 , \14567 , \14568 , \14569 , \14570 ,
         \14571 , \14572 , \14573 , \14574 , \14575 , \14576 , \14577 , \14578 , \14579 , \14580 ,
         \14581 , \14582 , \14583 , \14584 , \14585 , \14586 , \14587 , \14588 , \14589 , \14590 ,
         \14591 , \14592 , \14593 , \14594 , \14595 , \14596 , \14597 , \14598 , \14599 , \14600 ,
         \14601 , \14602 , \14603 , \14604 , \14605 , \14606 , \14607 , \14608 , \14609 , \14610 ,
         \14611 , \14612 , \14613 , \14614 , \14615 , \14616 , \14617 , \14618 , \14619 , \14620 ,
         \14621 , \14622 , \14623 , \14624 , \14625 , \14626 , \14627 , \14628 , \14629 , \14630 ,
         \14631 , \14632 , \14633 , \14634 , \14635 , \14636 , \14637 , \14638 , \14639 , \14640 ,
         \14641 , \14642 , \14643 , \14644 , \14645 , \14646 , \14647 , \14648 , \14649 , \14650 ,
         \14651 , \14652 , \14653 , \14654 , \14655 , \14656 , \14657 , \14658 , \14659 , \14660 ,
         \14661 , \14662 , \14663 , \14664 , \14665 , \14666 , \14667 , \14668 , \14669 , \14670 ,
         \14671 , \14672 , \14673 , \14674 , \14675 , \14676 , \14677 , \14678 , \14679 , \14680 ,
         \14681 , \14682 , \14683 , \14684 , \14685 , \14686 , \14687 , \14688 , \14689 , \14690 ,
         \14691 , \14692 , \14693 , \14694 , \14695 , \14696 , \14697 , \14698 , \14699 , \14700 ,
         \14701 , \14702 , \14703 , \14704 , \14705 , \14706 , \14707 , \14708 , \14709 , \14710 ,
         \14711 , \14712 , \14713 , \14714 , \14715 , \14716 , \14717 , \14718 , \14719 , \14720 ,
         \14721 , \14722 , \14723 , \14724 , \14725 , \14726 , \14727 , \14728 , \14729 , \14730 ,
         \14731 , \14732 , \14733 , \14734 , \14735 , \14736 , \14737 , \14738 , \14739 , \14740 ,
         \14741 , \14742 , \14743 , \14744 , \14745 , \14746 , \14747 , \14748 , \14749 , \14750 ,
         \14751 , \14752 , \14753 , \14754 , \14755 , \14756 , \14757 , \14758 , \14759 , \14760 ,
         \14761 , \14762 , \14763 , \14764 , \14765 , \14766 , \14767 , \14768 , \14769 , \14770 ,
         \14771 , \14772 , \14773 , \14774 , \14775 , \14776 , \14777 , \14778 , \14779 , \14780 ,
         \14781 , \14782 , \14783 , \14784 , \14785 , \14786 , \14787 , \14788 , \14789 , \14790 ,
         \14791 , \14792 , \14793 , \14794 , \14795 , \14796 , \14797 , \14798 , \14799 , \14800 ,
         \14801 , \14802 , \14803 , \14804 , \14805 , \14806 , \14807 , \14808 , \14809 , \14810 ,
         \14811 , \14812 , \14813 , \14814 , \14815 , \14816 , \14817 , \14818 , \14819 , \14820 ,
         \14821 , \14822 , \14823 , \14824 , \14825 , \14826 , \14827 , \14828 , \14829 , \14830 ,
         \14831 , \14832 , \14833 , \14834 , \14835 , \14836 , \14837 , \14838 , \14839 , \14840 ,
         \14841 , \14842 , \14843 , \14844 , \14845 , \14846 , \14847 , \14848 , \14849 , \14850 ,
         \14851 , \14852 , \14853 , \14854 , \14855 , \14856 , \14857 , \14858 , \14859 , \14860 ,
         \14861 , \14862 , \14863 , \14864 , \14865 , \14866 , \14867 , \14868 , \14869 , \14870 ,
         \14871 , \14872 , \14873 , \14874 , \14875 , \14876 , \14877 , \14878 , \14879 , \14880 ,
         \14881 , \14882 , \14883 , \14884 , \14885 , \14886 , \14887 , \14888 , \14889 , \14890 ,
         \14891 , \14892 , \14893 , \14894 , \14895 , \14896 , \14897 , \14898 , \14899 , \14900 ,
         \14901 , \14902 , \14903 , \14904 , \14905 , \14906 , \14907 , \14908 , \14909 , \14910 ,
         \14911 , \14912 , \14913 , \14914 , \14915 , \14916 , \14917 , \14918 , \14919 , \14920 ,
         \14921 , \14922 , \14923 , \14924 , \14925 , \14926 , \14927 , \14928 , \14929 , \14930 ,
         \14931 , \14932 , \14933 , \14934 , \14935 , \14936 , \14937 , \14938 , \14939 , \14940 ,
         \14941 , \14942 , \14943 , \14944 , \14945 , \14946 , \14947 , \14948 , \14949 , \14950 ,
         \14951 , \14952 , \14953 , \14954 , \14955 , \14956 , \14957 , \14958 , \14959 , \14960 ,
         \14961 , \14962 , \14963 , \14964 , \14965 , \14966 , \14967 , \14968 , \14969 , \14970 ,
         \14971 , \14972 , \14973 , \14974 , \14975 , \14976 , \14977 , \14978 , \14979 , \14980 ,
         \14981 , \14982 , \14983 , \14984 , \14985 , \14986 , \14987 , \14988 , \14989 , \14990 ,
         \14991 , \14992 , \14993 , \14994 , \14995 , \14996 , \14997 , \14998 , \14999 , \15000 ,
         \15001 , \15002 , \15003 , \15004 , \15005 , \15006 , \15007 , \15008 , \15009 , \15010 ,
         \15011 , \15012 , \15013 , \15014 , \15015 , \15016 , \15017 , \15018 , \15019 , \15020 ,
         \15021 , \15022 , \15023 , \15024 , \15025 , \15026 , \15027 , \15028 , \15029 , \15030 ,
         \15031 , \15032 , \15033 , \15034 , \15035 , \15036 , \15037 , \15038 , \15039 , \15040 ,
         \15041 , \15042 , \15043 , \15044 , \15045 , \15046 , \15047 , \15048 , \15049 , \15050 ,
         \15051 , \15052 , \15053 , \15054 , \15055 , \15056 , \15057 , \15058 , \15059 , \15060 ,
         \15061 , \15062 , \15063 , \15064 , \15065 , \15066 , \15067 , \15068 , \15069 , \15070 ,
         \15071 , \15072 , \15073 , \15074 , \15075 , \15076 , \15077 , \15078 , \15079 , \15080 ,
         \15081 , \15082 , \15083 , \15084 , \15085 , \15086 , \15087 , \15088 , \15089 , \15090 ,
         \15091 , \15092 , \15093 , \15094 , \15095 , \15096 , \15097 , \15098 , \15099 , \15100 ,
         \15101 , \15102 , \15103 , \15104 , \15105 , \15106 , \15107 , \15108 , \15109 , \15110 ,
         \15111 , \15112 , \15113 , \15114 , \15115 , \15116 , \15117 , \15118 , \15119 , \15120 ,
         \15121 , \15122 , \15123 , \15124 , \15125 , \15126 , \15127 , \15128 , \15129 , \15130 ,
         \15131 , \15132 , \15133 , \15134 , \15135 , \15136 , \15137 , \15138 , \15139 , \15140 ,
         \15141 , \15142 , \15143 , \15144 , \15145 , \15146 , \15147 , \15148 , \15149 , \15150 ,
         \15151 , \15152 , \15153 , \15154 , \15155 , \15156 , \15157 , \15158 , \15159 , \15160 ,
         \15161 , \15162 , \15163 , \15164 , \15165 , \15166 , \15167 , \15168 , \15169 , \15170 ,
         \15171 , \15172 , \15173 , \15174 , \15175 , \15176 , \15177 , \15178 , \15179 , \15180 ,
         \15181 , \15182 , \15183 , \15184 , \15185 , \15186 , \15187 , \15188 , \15189 , \15190 ,
         \15191 , \15192 , \15193 , \15194 , \15195 , \15196 , \15197 , \15198 , \15199 , \15200 ,
         \15201 , \15202 , \15203 , \15204 , \15205 , \15206 , \15207 , \15208 , \15209 , \15210 ,
         \15211 , \15212 , \15213 , \15214 , \15215 , \15216 , \15217 , \15218 , \15219 , \15220 ,
         \15221 , \15222 , \15223 , \15224 , \15225 , \15226 , \15227 , \15228 , \15229 , \15230 ,
         \15231 , \15232 , \15233 , \15234 , \15235 , \15236 , \15237 , \15238 , \15239 , \15240 ,
         \15241 , \15242 , \15243 , \15244 , \15245 , \15246 , \15247 , \15248 , \15249 , \15250 ,
         \15251 , \15252 , \15253 , \15254 , \15255 , \15256 , \15257 , \15258 , \15259 , \15260 ,
         \15261 , \15262 , \15263 , \15264 , \15265 , \15266 , \15267 , \15268 , \15269 , \15270 ,
         \15271 , \15272 , \15273 , \15274 , \15275 , \15276 , \15277 , \15278 , \15279 , \15280 ,
         \15281 , \15282 , \15283 , \15284 , \15285 , \15286 , \15287 , \15288 , \15289 , \15290 ,
         \15291 , \15292 , \15293 , \15294 , \15295 , \15296 , \15297 , \15298 , \15299 , \15300 ,
         \15301 , \15302 , \15303 , \15304 , \15305 , \15306 , \15307 , \15308 , \15309 , \15310 ,
         \15311 , \15312 , \15313 , \15314 , \15315 , \15316 , \15317 , \15318 , \15319 , \15320 ,
         \15321 , \15322 , \15323 , \15324 , \15325 , \15326 , \15327 , \15328 , \15329 , \15330 ,
         \15331 , \15332 , \15333 , \15334 , \15335 , \15336 , \15337 , \15338 , \15339 , \15340 ,
         \15341 , \15342 , \15343 , \15344 , \15345 , \15346 , \15347 , \15348 , \15349 , \15350 ,
         \15351 , \15352 , \15353 , \15354 , \15355 , \15356 , \15357 , \15358 , \15359 , \15360 ,
         \15361 , \15362 , \15363 , \15364 , \15365 , \15366 , \15367 , \15368 , \15369 , \15370 ,
         \15371 , \15372 , \15373 , \15374 , \15375 , \15376 , \15377 , \15378 , \15379 , \15380 ,
         \15381 , \15382 , \15383 , \15384 , \15385 , \15386 , \15387 , \15388 , \15389 , \15390 ,
         \15391 , \15392 , \15393 , \15394 , \15395 , \15396 , \15397 , \15398 , \15399 , \15400 ,
         \15401 , \15402 , \15403 , \15404 , \15405 , \15406 , \15407 , \15408 , \15409 , \15410 ,
         \15411 , \15412 , \15413 , \15414 , \15415 , \15416 , \15417 , \15418 , \15419 , \15420 ,
         \15421 , \15422 , \15423 , \15424 , \15425 , \15426 , \15427 , \15428 , \15429 , \15430 ,
         \15431 , \15432 , \15433 , \15434 , \15435 , \15436 , \15437 , \15438 , \15439 , \15440 ,
         \15441 , \15442 , \15443 , \15444 , \15445 , \15446 , \15447 , \15448 , \15449 , \15450 ,
         \15451 , \15452 , \15453 , \15454 , \15455 , \15456 , \15457 , \15458 , \15459 , \15460 ,
         \15461 , \15462 , \15463 , \15464 , \15465 , \15466 , \15467 , \15468 , \15469 , \15470 ,
         \15471 , \15472 , \15473 , \15474 , \15475 , \15476 , \15477 , \15478 , \15479 , \15480 ,
         \15481 , \15482 , \15483 , \15484 , \15485 , \15486 , \15487 , \15488 , \15489 , \15490 ,
         \15491 , \15492 , \15493 , \15494 , \15495 , \15496 , \15497 , \15498 , \15499 , \15500 ,
         \15501 , \15502 , \15503 , \15504 , \15505 , \15506 , \15507 , \15508 , \15509 , \15510 ,
         \15511 , \15512 , \15513 , \15514 , \15515 , \15516 , \15517 , \15518 , \15519 , \15520 ,
         \15521 , \15522 , \15523 , \15524 , \15525 , \15526 , \15527 , \15528 , \15529 , \15530 ,
         \15531 , \15532 , \15533 , \15534 , \15535 , \15536 , \15537 , \15538 , \15539 , \15540 ,
         \15541 , \15542 , \15543 , \15544 , \15545 , \15546 , \15547 , \15548 , \15549 , \15550 ,
         \15551 , \15552 , \15553 , \15554 , \15555 , \15556 , \15557 , \15558 , \15559 , \15560 ,
         \15561 , \15562 , \15563 , \15564 , \15565 , \15566 , \15567 , \15568 , \15569 , \15570 ,
         \15571 , \15572 , \15573 , \15574 , \15575 , \15576 , \15577 , \15578 , \15579 , \15580 ,
         \15581 , \15582 , \15583 , \15584 , \15585 , \15586 , \15587 , \15588 , \15589 , \15590 ,
         \15591 , \15592 , \15593 , \15594 , \15595 , \15596 , \15597 , \15598 , \15599 , \15600 ,
         \15601 , \15602 , \15603 , \15604 , \15605 , \15606 , \15607 , \15608 , \15609 , \15610 ,
         \15611 , \15612 , \15613 , \15614 , \15615 , \15616 , \15617 , \15618 , \15619 , \15620 ,
         \15621 , \15622 , \15623 , \15624 , \15625 , \15626 , \15627 , \15628 , \15629 , \15630 ,
         \15631 , \15632 , \15633 , \15634 , \15635 , \15636 , \15637 , \15638 , \15639 , \15640 ,
         \15641 , \15642 , \15643 , \15644 , \15645 , \15646 , \15647 , \15648 , \15649 , \15650 ,
         \15651 , \15652 , \15653 , \15654 , \15655 , \15656 , \15657 , \15658 , \15659 , \15660 ,
         \15661 , \15662 , \15663 , \15664 , \15665 , \15666 , \15667 , \15668 , \15669 , \15670 ,
         \15671 , \15672 , \15673 , \15674 , \15675 , \15676 , \15677 , \15678 , \15679 , \15680 ,
         \15681 , \15682 , \15683 , \15684 , \15685 , \15686 , \15687 , \15688 , \15689 , \15690 ,
         \15691 , \15692 , \15693 , \15694 , \15695 , \15696 , \15697 , \15698 , \15699 , \15700 ,
         \15701 , \15702 , \15703 , \15704 , \15705 , \15706 , \15707 , \15708 , \15709 , \15710 ,
         \15711 , \15712 , \15713 , \15714 , \15715 , \15716 , \15717 , \15718 , \15719 , \15720 ,
         \15721 , \15722 , \15723 , \15724 , \15725 , \15726 , \15727 , \15728 , \15729 , \15730 ,
         \15731 , \15732 , \15733 , \15734 , \15735 , \15736 , \15737 , \15738 , \15739 , \15740 ,
         \15741 , \15742 , \15743 , \15744 , \15745 , \15746 , \15747 , \15748 , \15749 , \15750 ,
         \15751 , \15752 , \15753 , \15754 , \15755 , \15756 , \15757 , \15758 , \15759 , \15760 ,
         \15761 , \15762 , \15763 , \15764 , \15765 , \15766 , \15767 , \15768 , \15769 , \15770 ,
         \15771 , \15772 , \15773 , \15774 , \15775 , \15776 , \15777 , \15778 , \15779 , \15780 ,
         \15781 , \15782 , \15783 , \15784 , \15785 , \15786 , \15787 , \15788 , \15789 , \15790 ,
         \15791 , \15792 , \15793 , \15794 , \15795 , \15796 , \15797 , \15798 , \15799 , \15800 ,
         \15801 , \15802 , \15803 , \15804 , \15805 , \15806 , \15807 , \15808 , \15809 , \15810 ,
         \15811 , \15812 , \15813 , \15814 , \15815 , \15816 , \15817 , \15818 , \15819 , \15820 ,
         \15821 , \15822 , \15823 , \15824 , \15825 , \15826 , \15827 , \15828 , \15829 , \15830 ,
         \15831 , \15832 , \15833 , \15834 , \15835 , \15836 , \15837 , \15838 , \15839 , \15840 ,
         \15841 , \15842 , \15843 , \15844 , \15845 , \15846 , \15847 , \15848 , \15849 , \15850 ,
         \15851 , \15852 , \15853 , \15854 , \15855 , \15856 , \15857 , \15858 , \15859 , \15860 ,
         \15861 , \15862 , \15863 , \15864 , \15865 , \15866 , \15867 , \15868 , \15869 , \15870 ,
         \15871 , \15872 , \15873 , \15874 , \15875 , \15876 , \15877 , \15878 , \15879 , \15880 ,
         \15881 , \15882 , \15883 , \15884 , \15885 , \15886 , \15887 , \15888 , \15889 , \15890 ,
         \15891 , \15892 , \15893 , \15894 , \15895 , \15896 , \15897 , \15898 , \15899 , \15900 ,
         \15901 , \15902 , \15903 , \15904 , \15905 , \15906 , \15907 , \15908 , \15909 , \15910 ,
         \15911 , \15912 , \15913 , \15914 , \15915 , \15916 , \15917 , \15918 , \15919 , \15920 ,
         \15921 , \15922 , \15923 , \15924 , \15925 , \15926 , \15927 , \15928 , \15929 , \15930 ,
         \15931 , \15932 , \15933 , \15934 , \15935 , \15936 , \15937 , \15938 , \15939 , \15940 ,
         \15941 , \15942 , \15943 , \15944 , \15945 , \15946 , \15947 , \15948 , \15949 , \15950 ,
         \15951 , \15952 , \15953 , \15954 , \15955 , \15956 , \15957 , \15958 , \15959 , \15960 ,
         \15961 , \15962 , \15963 , \15964 , \15965 , \15966 , \15967 , \15968 , \15969 , \15970 ,
         \15971 , \15972 , \15973 , \15974 , \15975 , \15976 , \15977 , \15978 , \15979 , \15980 ,
         \15981 , \15982 , \15983 , \15984 , \15985 , \15986 , \15987 , \15988 , \15989 , \15990 ,
         \15991 , \15992 , \15993 , \15994 , \15995 , \15996 , \15997 , \15998 , \15999 , \16000 ,
         \16001 , \16002 , \16003 , \16004 , \16005 , \16006 , \16007 , \16008 , \16009 , \16010 ,
         \16011 , \16012 , \16013 , \16014 , \16015 , \16016 , \16017 , \16018 , \16019 , \16020 ,
         \16021 , \16022 , \16023 , \16024 , \16025 , \16026 , \16027 , \16028 , \16029 , \16030 ,
         \16031 , \16032 , \16033 , \16034 , \16035 , \16036 , \16037 , \16038 , \16039 , \16040 ,
         \16041 , \16042 , \16043 , \16044 , \16045 , \16046 , \16047 , \16048 , \16049 , \16050 ,
         \16051 , \16052 , \16053 , \16054 , \16055 , \16056 , \16057 , \16058 , \16059 , \16060 ,
         \16061 , \16062 , \16063 , \16064 , \16065 , \16066 , \16067 , \16068 , \16069 , \16070 ,
         \16071 , \16072 , \16073 , \16074 , \16075 , \16076 , \16077 , \16078 , \16079 , \16080 ,
         \16081 , \16082 , \16083 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 , \16090 ,
         \16091 , \16092 , \16093 , \16094 , \16095 , \16096 , \16097 , \16098 , \16099 , \16100 ,
         \16101 , \16102 , \16103 , \16104 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 ,
         \16111 , \16112 , \16113 , \16114 , \16115 , \16116 , \16117 , \16118 , \16119 , \16120 ,
         \16121 , \16122 , \16123 , \16124 , \16125 , \16126 , \16127 , \16128 , \16129 , \16130 ,
         \16131 , \16132 , \16133 , \16134 , \16135 , \16136 , \16137 , \16138 , \16139 , \16140 ,
         \16141 , \16142 , \16143 , \16144 , \16145 , \16146 , \16147 , \16148 , \16149 , \16150 ,
         \16151 , \16152 , \16153 , \16154 , \16155 , \16156 , \16157 , \16158 , \16159 , \16160 ,
         \16161 , \16162 , \16163 , \16164 , \16165 , \16166 , \16167 , \16168 , \16169 , \16170 ,
         \16171 , \16172 , \16173 , \16174 , \16175 , \16176 , \16177 , \16178 , \16179 , \16180 ,
         \16181 , \16182 , \16183 , \16184 , \16185 , \16186 , \16187 , \16188 , \16189 , \16190 ,
         \16191 , \16192 , \16193 , \16194 , \16195 , \16196 , \16197 , \16198 , \16199 , \16200 ,
         \16201 , \16202 , \16203 , \16204 , \16205 , \16206 , \16207 , \16208 , \16209 , \16210 ,
         \16211 , \16212 , \16213 , \16214 , \16215 , \16216 , \16217 , \16218 , \16219 , \16220 ,
         \16221 , \16222 , \16223 , \16224 , \16225 , \16226 , \16227 , \16228 , \16229 , \16230 ,
         \16231 , \16232 , \16233 , \16234 , \16235 , \16236 , \16237 , \16238 , \16239 , \16240 ,
         \16241 , \16242 , \16243 , \16244 , \16245 , \16246 , \16247 , \16248 , \16249 , \16250 ,
         \16251 , \16252 , \16253 , \16254 , \16255 , \16256 , \16257 , \16258 , \16259 , \16260 ,
         \16261 , \16262 , \16263 , \16264 , \16265 , \16266 , \16267 , \16268 , \16269 , \16270 ,
         \16271 , \16272 , \16273 , \16274 , \16275 , \16276 , \16277 , \16278 , \16279 , \16280 ,
         \16281 , \16282 , \16283 , \16284 , \16285 , \16286 , \16287 , \16288 , \16289 , \16290 ,
         \16291 , \16292 , \16293 , \16294 , \16295 , \16296 , \16297 , \16298 , \16299 , \16300 ,
         \16301 , \16302 , \16303 , \16304 , \16305 , \16306 , \16307 , \16308 , \16309 , \16310 ,
         \16311 , \16312 , \16313 , \16314 , \16315 , \16316 , \16317 , \16318 , \16319 , \16320 ,
         \16321 , \16322 , \16323 , \16324 , \16325 , \16326 , \16327 , \16328 , \16329 , \16330 ,
         \16331 , \16332 , \16333 , \16334 , \16335 , \16336 , \16337 , \16338 , \16339 , \16340 ,
         \16341 , \16342 , \16343 , \16344 , \16345 , \16346 , \16347 , \16348 , \16349 , \16350 ,
         \16351 , \16352 , \16353 , \16354 , \16355 , \16356 , \16357 , \16358 , \16359 , \16360 ,
         \16361 , \16362 , \16363 , \16364 , \16365 , \16366 , \16367 , \16368 , \16369 , \16370 ,
         \16371 , \16372 , \16373 , \16374 , \16375 , \16376 , \16377 , \16378 , \16379 , \16380 ,
         \16381 , \16382 , \16383 , \16384 , \16385 , \16386 , \16387 , \16388 , \16389 , \16390 ,
         \16391 , \16392 , \16393 , \16394 , \16395 , \16396 , \16397 , \16398 , \16399 , \16400 ,
         \16401 , \16402 , \16403 , \16404 , \16405 , \16406 , \16407 , \16408 , \16409 , \16410 ,
         \16411 , \16412 , \16413 , \16414 , \16415 , \16416 , \16417 , \16418 , \16419 , \16420 ,
         \16421 , \16422 , \16423 , \16424 , \16425 , \16426 , \16427 , \16428 , \16429 , \16430 ,
         \16431 , \16432 , \16433 , \16434 , \16435 , \16436 , \16437 , \16438 , \16439 , \16440 ,
         \16441 , \16442 , \16443 , \16444 , \16445 , \16446 , \16447 , \16448 , \16449 , \16450 ,
         \16451 , \16452 , \16453 , \16454 , \16455 , \16456 , \16457 , \16458 , \16459 , \16460 ,
         \16461 , \16462 , \16463 , \16464 , \16465 , \16466 , \16467 , \16468 , \16469 , \16470 ,
         \16471 , \16472 , \16473 , \16474 , \16475 , \16476 , \16477 , \16478 , \16479 , \16480 ,
         \16481 , \16482 , \16483 , \16484 , \16485 , \16486 , \16487 , \16488 , \16489 , \16490 ,
         \16491 , \16492 , \16493 , \16494 , \16495 , \16496 , \16497 , \16498 , \16499 , \16500 ,
         \16501 , \16502 , \16503 , \16504 , \16505 , \16506 , \16507 , \16508 , \16509 , \16510 ,
         \16511 , \16512 , \16513 , \16514 , \16515 , \16516 , \16517 , \16518 , \16519 , \16520 ,
         \16521 , \16522 , \16523 , \16524 , \16525 , \16526 , \16527 , \16528 , \16529 , \16530 ,
         \16531 , \16532 , \16533 , \16534 , \16535 , \16536 , \16537 , \16538 , \16539 , \16540 ,
         \16541 , \16542 , \16543 , \16544 , \16545 , \16546 , \16547 , \16548 , \16549 , \16550 ,
         \16551 , \16552 , \16553 , \16554 , \16555 , \16556 , \16557 , \16558 , \16559 , \16560 ,
         \16561 , \16562 , \16563 , \16564 , \16565 , \16566 , \16567 , \16568 , \16569 , \16570 ,
         \16571 , \16572 , \16573 , \16574 , \16575 , \16576 , \16577 , \16578 , \16579 , \16580 ,
         \16581 , \16582 , \16583 , \16584 , \16585 , \16586 , \16587 , \16588 , \16589 , \16590 ,
         \16591 , \16592 , \16593 , \16594 , \16595 , \16596 , \16597 , \16598 , \16599 , \16600 ,
         \16601 , \16602 , \16603 , \16604 , \16605 , \16606 , \16607 , \16608 , \16609 , \16610 ,
         \16611 , \16612 , \16613 , \16614 , \16615 , \16616 , \16617 , \16618 , \16619 , \16620 ,
         \16621 , \16622 , \16623 , \16624 , \16625 , \16626 , \16627 , \16628 , \16629 , \16630 ,
         \16631 , \16632 , \16633 , \16634 , \16635 , \16636 , \16637 , \16638 , \16639 , \16640 ,
         \16641 , \16642 , \16643 , \16644 , \16645 , \16646 , \16647 , \16648 , \16649 , \16650 ,
         \16651 , \16652 , \16653 , \16654 , \16655 , \16656 , \16657 , \16658 , \16659 , \16660 ,
         \16661 , \16662 , \16663 , \16664 , \16665 , \16666 , \16667 , \16668 , \16669 , \16670 ,
         \16671 , \16672 , \16673 , \16674 , \16675 , \16676 , \16677 , \16678 , \16679 , \16680 ,
         \16681 , \16682 , \16683 , \16684 , \16685 , \16686 , \16687 , \16688 , \16689 , \16690 ,
         \16691 , \16692 , \16693 , \16694 , \16695 , \16696 , \16697 , \16698 , \16699 , \16700 ,
         \16701 , \16702 , \16703 , \16704 , \16705 , \16706 , \16707 , \16708 , \16709 , \16710 ,
         \16711 , \16712 , \16713 , \16714 , \16715 , \16716 , \16717 , \16718 , \16719 , \16720 ,
         \16721 , \16722 , \16723 , \16724 , \16725 , \16726 , \16727 , \16728 , \16729 , \16730 ,
         \16731 , \16732 , \16733 , \16734 , \16735 , \16736 , \16737 , \16738 , \16739 , \16740 ,
         \16741 , \16742 , \16743 , \16744 , \16745 , \16746 , \16747 , \16748 , \16749 , \16750 ,
         \16751 , \16752 , \16753 , \16754 , \16755 , \16756 , \16757 , \16758 , \16759 , \16760 ,
         \16761 , \16762 , \16763 , \16764 , \16765 , \16766 , \16767 , \16768 , \16769 , \16770 ,
         \16771 , \16772 , \16773 , \16774 , \16775 , \16776 , \16777 , \16778 , \16779 , \16780 ,
         \16781 , \16782 , \16783 , \16784 , \16785 , \16786 , \16787 , \16788 , \16789 , \16790 ,
         \16791 , \16792 , \16793 , \16794 , \16795 , \16796 , \16797 , \16798 , \16799 , \16800 ,
         \16801 , \16802 , \16803 , \16804 , \16805 , \16806 , \16807 , \16808 , \16809 , \16810 ,
         \16811 , \16812 , \16813 , \16814 , \16815 , \16816 , \16817 , \16818 , \16819 , \16820 ,
         \16821 , \16822 , \16823 , \16824 , \16825 , \16826 , \16827 , \16828 , \16829 , \16830 ,
         \16831 , \16832 , \16833 , \16834 , \16835 , \16836 , \16837 , \16838 , \16839 , \16840 ,
         \16841 , \16842 , \16843 , \16844 , \16845 , \16846 , \16847 , \16848 , \16849 , \16850 ,
         \16851 , \16852 , \16853 , \16854 , \16855 , \16856 , \16857 , \16858 , \16859 , \16860 ,
         \16861 , \16862 , \16863 , \16864 , \16865 , \16866 , \16867 , \16868 , \16869 , \16870 ,
         \16871 , \16872 , \16873 , \16874 , \16875 , \16876 , \16877 , \16878 , \16879 , \16880 ,
         \16881 , \16882 , \16883 , \16884 , \16885 , \16886 , \16887 , \16888 , \16889 , \16890 ,
         \16891 , \16892 , \16893 , \16894 , \16895 , \16896 , \16897 , \16898 , \16899 , \16900 ,
         \16901 , \16902 , \16903 , \16904 , \16905 , \16906 , \16907 , \16908 , \16909 , \16910 ,
         \16911 , \16912 , \16913 , \16914 , \16915 , \16916 , \16917 , \16918 , \16919 , \16920 ,
         \16921 , \16922 , \16923 , \16924 , \16925 , \16926 , \16927 , \16928 , \16929 , \16930 ,
         \16931 , \16932 , \16933 , \16934 , \16935 , \16936 , \16937 , \16938 , \16939 , \16940 ,
         \16941 , \16942 , \16943 , \16944 , \16945 , \16946 , \16947 , \16948 , \16949 , \16950 ,
         \16951 , \16952 , \16953 , \16954 , \16955 , \16956 , \16957 , \16958 , \16959 , \16960 ,
         \16961 , \16962 , \16963 , \16964 , \16965 , \16966 , \16967 , \16968 , \16969 , \16970 ,
         \16971 , \16972 , \16973 , \16974 , \16975 , \16976 , \16977 , \16978 , \16979 , \16980 ,
         \16981 , \16982 , \16983 , \16984 , \16985 , \16986 , \16987 , \16988 , \16989 , \16990 ,
         \16991 , \16992 , \16993 , \16994 , \16995 , \16996 , \16997 , \16998 , \16999 , \17000 ,
         \17001 , \17002 , \17003 , \17004 , \17005 , \17006 , \17007 , \17008 , \17009 , \17010 ,
         \17011 , \17012 , \17013 , \17014 , \17015 , \17016 , \17017 , \17018 , \17019 , \17020 ,
         \17021 , \17022 , \17023 , \17024 , \17025 , \17026 , \17027 , \17028 , \17029 , \17030 ,
         \17031 , \17032 , \17033 , \17034 , \17035 , \17036 , \17037 , \17038 , \17039 , \17040 ,
         \17041 , \17042 , \17043 , \17044 , \17045 , \17046 , \17047 , \17048 , \17049 , \17050 ,
         \17051 , \17052 , \17053 , \17054 , \17055 , \17056 , \17057 , \17058 , \17059 , \17060 ,
         \17061 , \17062 , \17063 , \17064 , \17065 , \17066 , \17067 , \17068 , \17069 , \17070 ,
         \17071 , \17072 , \17073 , \17074 , \17075 , \17076 , \17077 , \17078 , \17079 , \17080 ,
         \17081 , \17082 , \17083 , \17084 , \17085 , \17086 , \17087 , \17088 , \17089 , \17090 ,
         \17091 , \17092 , \17093 , \17094 , \17095 , \17096 , \17097 , \17098 , \17099 , \17100 ,
         \17101 , \17102 , \17103 , \17104 , \17105 , \17106 , \17107 , \17108 , \17109 , \17110 ,
         \17111 , \17112 , \17113 , \17114 , \17115 , \17116 , \17117 , \17118 , \17119 , \17120 ,
         \17121 , \17122 , \17123 , \17124 , \17125 , \17126 , \17127 , \17128 , \17129 , \17130 ,
         \17131 , \17132 , \17133 , \17134 , \17135 , \17136 , \17137 , \17138 , \17139 , \17140 ,
         \17141 , \17142 , \17143 , \17144 , \17145 , \17146 , \17147 , \17148 , \17149 , \17150 ,
         \17151 , \17152 , \17153 , \17154 , \17155 , \17156 , \17157 , \17158 , \17159 , \17160 ,
         \17161 , \17162 , \17163 , \17164 , \17165 , \17166 , \17167 , \17168 , \17169 , \17170 ,
         \17171 , \17172 , \17173 , \17174 , \17175 , \17176 , \17177 , \17178 , \17179 , \17180 ,
         \17181 , \17182 , \17183 , \17184 , \17185 , \17186 , \17187 , \17188 , \17189 , \17190 ,
         \17191 , \17192 , \17193 , \17194 , \17195 , \17196 , \17197 , \17198 , \17199 , \17200 ,
         \17201 , \17202 , \17203 , \17204 , \17205 , \17206 , \17207 , \17208 , \17209 , \17210 ,
         \17211 , \17212 , \17213 , \17214 , \17215 , \17216 , \17217 , \17218 , \17219 , \17220 ,
         \17221 , \17222 , \17223 , \17224 , \17225 , \17226 , \17227 , \17228 , \17229 , \17230 ,
         \17231 , \17232 , \17233 , \17234 , \17235 , \17236 , \17237 , \17238 , \17239 , \17240 ,
         \17241 , \17242 , \17243 , \17244 , \17245 , \17246 , \17247 , \17248 , \17249 , \17250 ,
         \17251 , \17252 , \17253 , \17254 , \17255 , \17256 , \17257 , \17258 , \17259 , \17260 ,
         \17261 , \17262 , \17263 , \17264 , \17265 , \17266 , \17267 , \17268 , \17269 , \17270 ,
         \17271 , \17272 , \17273 , \17274 , \17275 , \17276 , \17277 , \17278 , \17279 , \17280 ,
         \17281 , \17282 , \17283 , \17284 , \17285 , \17286 , \17287 , \17288 , \17289 , \17290 ,
         \17291 , \17292 , \17293 , \17294 , \17295 , \17296 , \17297 , \17298 , \17299 , \17300 ,
         \17301 , \17302 , \17303 , \17304 , \17305 , \17306 , \17307 , \17308 , \17309 , \17310 ,
         \17311 , \17312 , \17313 , \17314 , \17315 , \17316 , \17317 , \17318 , \17319 , \17320 ,
         \17321 , \17322 , \17323 , \17324 , \17325 , \17326 , \17327 , \17328 , \17329 , \17330 ,
         \17331 , \17332 , \17333 , \17334 , \17335 , \17336 , \17337 , \17338 , \17339 , \17340 ,
         \17341 , \17342 , \17343 , \17344 , \17345 , \17346 , \17347 , \17348 , \17349 , \17350 ,
         \17351 , \17352 , \17353 , \17354 , \17355 , \17356 , \17357 , \17358 , \17359 , \17360 ,
         \17361 , \17362 , \17363 , \17364 , \17365 , \17366 , \17367 , \17368 , \17369 , \17370 ,
         \17371 , \17372 , \17373 , \17374 , \17375 , \17376 , \17377 , \17378 , \17379 , \17380 ,
         \17381 , \17382 , \17383 , \17384 , \17385 , \17386 , \17387 , \17388 , \17389 , \17390 ,
         \17391 , \17392 , \17393 , \17394 , \17395 , \17396 , \17397 , \17398 , \17399 , \17400 ,
         \17401 , \17402 , \17403 , \17404 , \17405 , \17406 , \17407 , \17408 , \17409 , \17410 ,
         \17411 , \17412 , \17413 , \17414 , \17415 , \17416 , \17417 , \17418 , \17419 , \17420 ,
         \17421 , \17422 , \17423 , \17424 , \17425 , \17426 , \17427 , \17428 , \17429 , \17430 ,
         \17431 , \17432 , \17433 , \17434 , \17435 , \17436 , \17437 , \17438 , \17439 , \17440 ,
         \17441 , \17442 , \17443 , \17444 , \17445 , \17446 , \17447 , \17448 , \17449 , \17450 ,
         \17451 , \17452 , \17453 , \17454 , \17455 , \17456 , \17457 , \17458 , \17459 , \17460 ,
         \17461 , \17462 , \17463 , \17464 , \17465 , \17466 , \17467 , \17468 , \17469 , \17470 ,
         \17471 , \17472 , \17473 , \17474 , \17475 , \17476 , \17477 , \17478 , \17479 , \17480 ,
         \17481 , \17482 , \17483 , \17484 , \17485 , \17486 , \17487 , \17488 , \17489 , \17490 ,
         \17491 , \17492 , \17493 , \17494 , \17495 , \17496 , \17497 , \17498 , \17499 , \17500 ,
         \17501 , \17502 , \17503 , \17504 , \17505 , \17506 , \17507 , \17508 , \17509 , \17510 ,
         \17511 , \17512 , \17513 , \17514 , \17515 , \17516 , \17517 , \17518 , \17519 , \17520 ,
         \17521 , \17522 , \17523 , \17524 , \17525 , \17526 , \17527 , \17528 , \17529 , \17530 ,
         \17531 , \17532 , \17533 , \17534 , \17535 , \17536 , \17537 , \17538 , \17539 , \17540 ,
         \17541 , \17542 , \17543 , \17544 , \17545 , \17546 , \17547 , \17548 , \17549 , \17550 ,
         \17551 , \17552 , \17553 , \17554 , \17555 , \17556 , \17557 , \17558 , \17559 , \17560 ,
         \17561 , \17562 , \17563 , \17564 , \17565 , \17566 , \17567 , \17568 , \17569 , \17570 ,
         \17571 , \17572 , \17573 , \17574 , \17575 , \17576 , \17577 , \17578 , \17579 , \17580 ,
         \17581 , \17582 , \17583 , \17584 , \17585 , \17586 , \17587 , \17588 , \17589 , \17590 ,
         \17591 , \17592 , \17593 , \17594 , \17595 , \17596 , \17597 , \17598 , \17599 , \17600 ,
         \17601 , \17602 , \17603 , \17604 , \17605 , \17606 , \17607 , \17608 , \17609 , \17610 ,
         \17611 , \17612 , \17613 , \17614 , \17615 , \17616 , \17617 , \17618 , \17619 , \17620 ,
         \17621 , \17622 , \17623 , \17624 , \17625 , \17626 , \17627 , \17628 , \17629 , \17630 ,
         \17631 , \17632 , \17633 , \17634 , \17635 , \17636 , \17637 , \17638 , \17639 , \17640 ,
         \17641 , \17642 , \17643 , \17644 , \17645 , \17646 , \17647 , \17648 , \17649 , \17650 ,
         \17651 , \17652 , \17653 , \17654 , \17655 , \17656 , \17657 , \17658 , \17659 , \17660 ,
         \17661 , \17662 , \17663 , \17664 , \17665 , \17666 , \17667 , \17668 , \17669 , \17670 ,
         \17671 , \17672 , \17673 , \17674 , \17675 , \17676 , \17677 , \17678 , \17679 , \17680 ,
         \17681 , \17682 , \17683 , \17684 , \17685 , \17686 , \17687 , \17688 , \17689 , \17690 ,
         \17691 , \17692 , \17693 , \17694 , \17695 , \17696 , \17697 , \17698 , \17699 , \17700 ,
         \17701 , \17702 , \17703 , \17704 , \17705 , \17706 , \17707 , \17708 , \17709 , \17710 ,
         \17711 , \17712 , \17713 , \17714 , \17715 , \17716 , \17717 , \17718 , \17719 , \17720 ,
         \17721 , \17722 , \17723 , \17724 , \17725 , \17726 , \17727 , \17728 , \17729 , \17730 ,
         \17731 , \17732 , \17733 , \17734 , \17735 , \17736 , \17737 , \17738 , \17739 , \17740 ,
         \17741 , \17742 , \17743 , \17744 , \17745 , \17746 , \17747 , \17748 , \17749 , \17750 ,
         \17751 , \17752 , \17753 , \17754 , \17755 , \17756 , \17757 , \17758 , \17759 , \17760 ,
         \17761 , \17762 , \17763 , \17764 , \17765 , \17766 , \17767 , \17768 , \17769 , \17770 ,
         \17771 , \17772 , \17773 , \17774 , \17775 , \17776 , \17777 , \17778 , \17779 , \17780 ,
         \17781 , \17782 , \17783 , \17784 , \17785 , \17786 , \17787 , \17788 , \17789 , \17790 ,
         \17791 , \17792 , \17793 , \17794 , \17795 , \17796 , \17797 , \17798 , \17799 , \17800 ,
         \17801 , \17802 , \17803 , \17804 , \17805 , \17806 , \17807 , \17808 , \17809 , \17810 ,
         \17811 , \17812 , \17813 , \17814 , \17815 , \17816 , \17817 , \17818 , \17819 , \17820 ,
         \17821 , \17822 , \17823 , \17824 , \17825 , \17826 , \17827 , \17828 , \17829 , \17830 ,
         \17831 , \17832 , \17833 , \17834 , \17835 , \17836 , \17837 , \17838 , \17839 , \17840 ,
         \17841 , \17842 , \17843 , \17844 , \17845 , \17846 , \17847 , \17848 , \17849 , \17850 ,
         \17851 , \17852 , \17853 , \17854 , \17855 , \17856 , \17857 , \17858 , \17859 , \17860 ,
         \17861 , \17862 , \17863 , \17864 , \17865 , \17866 , \17867 , \17868 , \17869 , \17870 ,
         \17871 , \17872 , \17873 , \17874 , \17875 , \17876 , \17877 , \17878 , \17879 , \17880 ,
         \17881 , \17882 , \17883 , \17884 , \17885 , \17886 , \17887 , \17888 , \17889 , \17890 ,
         \17891 , \17892 , \17893 , \17894 , \17895 , \17896 , \17897 , \17898 , \17899 , \17900 ,
         \17901 , \17902 , \17903 , \17904 , \17905 , \17906 , \17907 , \17908 , \17909 , \17910 ,
         \17911 , \17912 , \17913 , \17914 , \17915 , \17916 , \17917 , \17918 , \17919 , \17920 ,
         \17921 , \17922 , \17923 , \17924 , \17925 , \17926 , \17927 , \17928 , \17929 , \17930 ,
         \17931 , \17932 , \17933 , \17934 , \17935 , \17936 , \17937 , \17938 , \17939 , \17940 ,
         \17941 , \17942 , \17943 , \17944 , \17945 , \17946 , \17947 , \17948 , \17949 , \17950 ,
         \17951 , \17952 , \17953 , \17954 , \17955 , \17956 , \17957 , \17958 , \17959 , \17960 ,
         \17961 , \17962 , \17963 , \17964 , \17965 , \17966 , \17967 , \17968 , \17969 , \17970 ,
         \17971 , \17972 , \17973 , \17974 , \17975 , \17976 , \17977 , \17978 , \17979 , \17980 ,
         \17981 , \17982 , \17983 , \17984 , \17985 , \17986 , \17987 , \17988 , \17989 , \17990 ,
         \17991 , \17992 , \17993 , \17994 , \17995 , \17996 , \17997 , \17998 , \17999 , \18000 ,
         \18001 , \18002 , \18003 , \18004 , \18005 , \18006 , \18007 , \18008 , \18009 , \18010 ,
         \18011 , \18012 , \18013 , \18014 , \18015 , \18016 , \18017 , \18018 , \18019 , \18020 ,
         \18021 , \18022 , \18023 , \18024 , \18025 , \18026 , \18027 , \18028 , \18029 , \18030 ,
         \18031 , \18032 , \18033 , \18034 , \18035 , \18036 , \18037 , \18038 , \18039 , \18040 ,
         \18041 , \18042 , \18043 , \18044 , \18045 , \18046 , \18047 , \18048 , \18049 , \18050 ,
         \18051 , \18052 , \18053 , \18054 , \18055 , \18056 , \18057 , \18058 , \18059 , \18060 ,
         \18061 , \18062 , \18063 , \18064 , \18065 , \18066 , \18067 , \18068 , \18069 , \18070 ,
         \18071 , \18072 , \18073 , \18074 , \18075 , \18076 , \18077 , \18078 , \18079 , \18080 ,
         \18081 , \18082 , \18083 , \18084 , \18085 , \18086 , \18087 , \18088 , \18089 , \18090 ,
         \18091 , \18092 , \18093 , \18094 , \18095 , \18096 , \18097 , \18098 , \18099 , \18100 ,
         \18101 , \18102 , \18103 , \18104 , \18105 , \18106 , \18107 , \18108 , \18109 , \18110 ,
         \18111 , \18112 , \18113 , \18114 , \18115 , \18116 , \18117 , \18118 , \18119 , \18120 ,
         \18121 , \18122 , \18123 , \18124 , \18125 , \18126 , \18127 , \18128 , \18129 , \18130 ,
         \18131 , \18132 , \18133 , \18134 , \18135 , \18136 , \18137 , \18138 , \18139 , \18140 ,
         \18141 , \18142 , \18143 , \18144 , \18145 , \18146 , \18147 , \18148 , \18149 , \18150 ,
         \18151 , \18152 , \18153 , \18154 , \18155 , \18156 , \18157 , \18158 , \18159 , \18160 ,
         \18161 , \18162 , \18163 , \18164 , \18165 , \18166 , \18167 , \18168 , \18169 , \18170 ,
         \18171 , \18172 , \18173 , \18174 , \18175 , \18176 , \18177 , \18178 , \18179 , \18180 ,
         \18181 , \18182 , \18183 , \18184 , \18185 , \18186 , \18187 , \18188 , \18189 , \18190 ,
         \18191 , \18192 , \18193 , \18194 , \18195 , \18196 , \18197 , \18198 , \18199 , \18200 ,
         \18201 , \18202 , \18203 , \18204 , \18205 , \18206 , \18207 , \18208 , \18209 , \18210 ,
         \18211 , \18212 , \18213 , \18214 , \18215 , \18216 , \18217 , \18218 , \18219 , \18220 ,
         \18221 , \18222 , \18223 , \18224 , \18225 , \18226 , \18227 , \18228 , \18229 , \18230 ,
         \18231 , \18232 , \18233 , \18234 , \18235 , \18236 , \18237 , \18238 , \18239 , \18240 ,
         \18241 , \18242 , \18243 , \18244 , \18245 , \18246 , \18247 , \18248 , \18249 , \18250 ,
         \18251 , \18252 , \18253 , \18254 , \18255 , \18256 , \18257 , \18258 , \18259 , \18260 ,
         \18261 , \18262 , \18263 , \18264 , \18265 , \18266 , \18267 , \18268 , \18269 , \18270 ,
         \18271 , \18272 , \18273 , \18274 , \18275 , \18276 , \18277 , \18278 , \18279 , \18280 ,
         \18281 , \18282 , \18283 , \18284 , \18285 , \18286 , \18287 , \18288 , \18289 , \18290 ,
         \18291 , \18292 , \18293 , \18294 , \18295 , \18296 , \18297 , \18298 , \18299 , \18300 ,
         \18301 , \18302 , \18303 , \18304 , \18305 , \18306 , \18307 , \18308 , \18309 , \18310 ,
         \18311 , \18312 , \18313 , \18314 , \18315 , \18316 , \18317 , \18318 , \18319 , \18320 ,
         \18321 , \18322 , \18323 , \18324 , \18325 , \18326 , \18327 , \18328 , \18329 , \18330 ,
         \18331 , \18332 , \18333 , \18334 , \18335 , \18336 , \18337 , \18338 , \18339 , \18340 ,
         \18341 , \18342 , \18343 , \18344 , \18345 , \18346 , \18347 , \18348 , \18349 , \18350 ,
         \18351 , \18352 , \18353 , \18354 , \18355 , \18356 , \18357 , \18358 , \18359 , \18360 ,
         \18361 , \18362 , \18363 , \18364 , \18365 , \18366 , \18367 , \18368 , \18369 , \18370 ,
         \18371 , \18372 , \18373 , \18374 , \18375 , \18376 , \18377 , \18378 , \18379 , \18380 ,
         \18381 , \18382 , \18383 , \18384 , \18385 , \18386 , \18387 , \18388 , \18389 , \18390 ,
         \18391 , \18392 , \18393 , \18394 , \18395 , \18396 , \18397 , \18398 , \18399 , \18400 ,
         \18401 , \18402 , \18403 , \18404 , \18405 , \18406 , \18407 , \18408 , \18409 , \18410 ,
         \18411 , \18412 , \18413 , \18414 , \18415 , \18416 , \18417 , \18418 , \18419 , \18420 ,
         \18421 , \18422 , \18423 , \18424 , \18425 , \18426 , \18427 , \18428 , \18429 , \18430 ,
         \18431 , \18432 , \18433 , \18434 , \18435 , \18436 , \18437 , \18438 , \18439 , \18440 ,
         \18441 , \18442 , \18443 , \18444 , \18445 , \18446 , \18447 , \18448 , \18449 , \18450 ,
         \18451 , \18452 , \18453 , \18454 , \18455 , \18456 , \18457 , \18458 , \18459 , \18460 ,
         \18461 , \18462 , \18463 , \18464 , \18465 , \18466 , \18467 , \18468 , \18469 , \18470 ,
         \18471 , \18472 , \18473 , \18474 , \18475 , \18476 , \18477 , \18478 , \18479 , \18480 ,
         \18481 , \18482 , \18483 , \18484 , \18485 , \18486 , \18487 , \18488 , \18489 , \18490 ,
         \18491 , \18492 , \18493 , \18494 , \18495 , \18496 , \18497 , \18498 , \18499 , \18500 ,
         \18501 , \18502 , \18503 , \18504 , \18505 , \18506 , \18507 , \18508 , \18509 , \18510 ,
         \18511 , \18512 , \18513 , \18514 , \18515 , \18516 , \18517 , \18518 , \18519 , \18520 ,
         \18521 , \18522 , \18523 , \18524 , \18525 , \18526 , \18527 , \18528 , \18529 , \18530 ,
         \18531 , \18532 , \18533 , \18534 , \18535 , \18536 , \18537 , \18538 , \18539 , \18540 ,
         \18541 , \18542 , \18543 , \18544 , \18545 , \18546 , \18547 , \18548 , \18549 , \18550 ,
         \18551 , \18552 , \18553 , \18554 , \18555 , \18556 , \18557 , \18558 , \18559 , \18560 ,
         \18561 , \18562 , \18563 , \18564 , \18565 , \18566 , \18567 , \18568 , \18569 , \18570 ,
         \18571 , \18572 , \18573 , \18574 , \18575 , \18576 , \18577 , \18578 , \18579 , \18580 ,
         \18581 , \18582 , \18583 , \18584 , \18585 , \18586 , \18587 , \18588 , \18589 , \18590 ,
         \18591 , \18592 , \18593 , \18594 , \18595 , \18596 , \18597 , \18598 , \18599 , \18600 ,
         \18601 , \18602 , \18603 , \18604 , \18605 , \18606 , \18607 , \18608 , \18609 , \18610 ,
         \18611 , \18612 , \18613 , \18614 , \18615 , \18616 , \18617 , \18618 , \18619 , \18620 ,
         \18621 , \18622 , \18623 , \18624 , \18625 , \18626 , \18627 , \18628 , \18629 , \18630 ,
         \18631 , \18632 , \18633 , \18634 , \18635 , \18636 , \18637 , \18638 , \18639 , \18640 ,
         \18641 , \18642 , \18643 , \18644 , \18645 , \18646 , \18647 , \18648 , \18649 , \18650 ,
         \18651 , \18652 , \18653 , \18654 , \18655 , \18656 , \18657 , \18658 , \18659 , \18660 ,
         \18661 , \18662 , \18663 , \18664 , \18665 , \18666 , \18667 , \18668 , \18669 , \18670 ,
         \18671 , \18672 , \18673 , \18674 , \18675 , \18676 , \18677 , \18678 , \18679 , \18680 ,
         \18681 , \18682 , \18683 , \18684 , \18685 , \18686 , \18687 , \18688 , \18689 , \18690 ,
         \18691 , \18692 , \18693 , \18694 , \18695 , \18696 , \18697 , \18698 , \18699 , \18700 ,
         \18701 , \18702 , \18703 , \18704 , \18705 , \18706 , \18707 , \18708 , \18709 , \18710 ,
         \18711 , \18712 , \18713 , \18714 , \18715 , \18716 , \18717 , \18718 , \18719 , \18720 ,
         \18721 , \18722 , \18723 , \18724 , \18725 , \18726 , \18727 , \18728 , \18729 , \18730 ,
         \18731 , \18732 , \18733 , \18734 , \18735 , \18736 , \18737 , \18738 , \18739 , \18740 ,
         \18741 , \18742 , \18743 , \18744 , \18745 , \18746 , \18747 , \18748 , \18749 , \18750 ,
         \18751 , \18752 , \18753 , \18754 , \18755 , \18756 , \18757 , \18758 , \18759 , \18760 ,
         \18761 , \18762 , \18763 , \18764 , \18765 , \18766 , \18767 , \18768 , \18769 , \18770 ,
         \18771 , \18772 , \18773 , \18774 , \18775 , \18776 , \18777 , \18778 , \18779 , \18780 ,
         \18781 , \18782 , \18783 , \18784 , \18785 , \18786 , \18787 , \18788 , \18789 , \18790 ,
         \18791 , \18792 , \18793 , \18794 , \18795 , \18796 , \18797 , \18798 , \18799 , \18800 ,
         \18801 , \18802 , \18803 , \18804 , \18805 , \18806 , \18807 , \18808 , \18809 , \18810 ,
         \18811 , \18812 , \18813 , \18814 , \18815 , \18816 , \18817 , \18818 , \18819 , \18820 ,
         \18821 , \18822 , \18823 , \18824 , \18825 , \18826 , \18827 , \18828 , \18829 , \18830 ,
         \18831 , \18832 , \18833 , \18834 , \18835 , \18836 , \18837 , \18838 , \18839 , \18840 ,
         \18841 , \18842 , \18843 , \18844 , \18845 , \18846 , \18847 , \18848 , \18849 , \18850 ,
         \18851 , \18852 , \18853 , \18854 , \18855 , \18856 , \18857 , \18858 , \18859 , \18860 ,
         \18861 , \18862 , \18863 , \18864 , \18865 , \18866 , \18867 , \18868 , \18869 , \18870 ,
         \18871 , \18872 , \18873 , \18874 , \18875 , \18876 , \18877 , \18878 , \18879 , \18880 ,
         \18881 , \18882 , \18883 , \18884 , \18885 , \18886 , \18887 , \18888 , \18889 , \18890 ,
         \18891 , \18892 , \18893 , \18894 , \18895 , \18896 , \18897 , \18898 , \18899 , \18900 ,
         \18901 , \18902 , \18903 , \18904 , \18905 , \18906 , \18907 , \18908 , \18909 , \18910 ,
         \18911 , \18912 , \18913 , \18914 , \18915 , \18916 , \18917 , \18918 , \18919 , \18920 ,
         \18921 , \18922 , \18923 , \18924 , \18925 , \18926 , \18927 , \18928 , \18929 , \18930 ,
         \18931 , \18932 , \18933 , \18934 , \18935 , \18936 , \18937 , \18938 , \18939 , \18940 ,
         \18941 , \18942 , \18943 , \18944 , \18945 , \18946 , \18947 , \18948 , \18949 , \18950 ,
         \18951 , \18952 , \18953 , \18954 , \18955 , \18956 , \18957 , \18958 , \18959 , \18960 ,
         \18961 , \18962 , \18963 , \18964 , \18965 , \18966 , \18967 , \18968 , \18969 , \18970 ,
         \18971 , \18972 , \18973 , \18974 , \18975 , \18976 , \18977 , \18978 , \18979 , \18980 ,
         \18981 , \18982 , \18983 , \18984 , \18985 , \18986 , \18987 , \18988 , \18989 , \18990 ,
         \18991 , \18992 , \18993 , \18994 , \18995 , \18996 , \18997 , \18998 , \18999 , \19000 ,
         \19001 , \19002 , \19003 , \19004 , \19005 , \19006 , \19007 , \19008 , \19009 , \19010 ,
         \19011 , \19012 , \19013 , \19014 , \19015 , \19016 , \19017 , \19018 , \19019 , \19020 ,
         \19021 , \19022 , \19023 , \19024 , \19025 , \19026 , \19027 , \19028 , \19029 , \19030 ,
         \19031 , \19032 , \19033 , \19034 , \19035 , \19036 , \19037 , \19038 , \19039 , \19040 ,
         \19041 , \19042 , \19043 , \19044 , \19045 , \19046 , \19047 , \19048 , \19049 , \19050 ,
         \19051 , \19052 , \19053 , \19054 , \19055 , \19056 , \19057 , \19058 , \19059 , \19060 ,
         \19061 , \19062 , \19063 , \19064 , \19065 , \19066 , \19067 , \19068 , \19069 , \19070 ,
         \19071 , \19072 , \19073 , \19074 , \19075 , \19076 , \19077 , \19078 , \19079 , \19080 ,
         \19081 , \19082 , \19083 , \19084 , \19085 , \19086 , \19087 , \19088 , \19089 , \19090 ,
         \19091 , \19092 , \19093 , \19094 , \19095 , \19096 , \19097 , \19098 , \19099 , \19100 ,
         \19101 , \19102 , \19103 , \19104 , \19105 , \19106 , \19107 , \19108 , \19109 , \19110 ,
         \19111 , \19112 , \19113 , \19114 , \19115 , \19116 , \19117 , \19118 , \19119 , \19120 ,
         \19121 , \19122 , \19123 , \19124 , \19125 , \19126 , \19127 , \19128 , \19129 , \19130 ,
         \19131 , \19132 , \19133 , \19134 , \19135 , \19136 , \19137 , \19138 , \19139 , \19140 ,
         \19141 , \19142 , \19143 , \19144 , \19145 , \19146 , \19147 , \19148 , \19149 , \19150 ,
         \19151 , \19152 , \19153 , \19154 , \19155 , \19156 , \19157 , \19158 , \19159 , \19160 ,
         \19161 , \19162 , \19163 , \19164 , \19165 , \19166 , \19167 , \19168 , \19169 , \19170 ,
         \19171 , \19172 , \19173 , \19174 , \19175 , \19176 , \19177 , \19178 , \19179 , \19180 ,
         \19181 , \19182 , \19183 , \19184 , \19185 , \19186 , \19187 , \19188 , \19189 , \19190 ,
         \19191 , \19192 , \19193 , \19194 , \19195 , \19196 , \19197 , \19198 , \19199 , \19200 ,
         \19201 , \19202 , \19203 , \19204 , \19205 , \19206 , \19207 , \19208 , \19209 , \19210 ,
         \19211 , \19212 , \19213 , \19214 , \19215 , \19216 , \19217 , \19218 , \19219 , \19220 ,
         \19221 , \19222 , \19223 , \19224 , \19225 , \19226 , \19227 , \19228 , \19229 , \19230 ,
         \19231 , \19232 , \19233 , \19234 , \19235 , \19236 , \19237 , \19238 , \19239 , \19240 ,
         \19241 , \19242 , \19243 , \19244 , \19245 , \19246 , \19247 , \19248 , \19249 , \19250 ,
         \19251 , \19252 , \19253 , \19254 , \19255 , \19256 , \19257 , \19258 , \19259 , \19260 ,
         \19261 , \19262 , \19263 , \19264 , \19265 , \19266 , \19267 , \19268 , \19269 , \19270 ,
         \19271 , \19272 , \19273 , \19274 , \19275 , \19276 , \19277 , \19278 , \19279 , \19280 ,
         \19281 , \19282 , \19283 , \19284 , \19285 , \19286 , \19287 , \19288 , \19289 , \19290 ,
         \19291 , \19292 , \19293 , \19294 , \19295 , \19296 , \19297 , \19298 , \19299 , \19300 ,
         \19301 , \19302 , \19303 , \19304 , \19305 , \19306 , \19307 , \19308 , \19309 , \19310 ,
         \19311 , \19312 , \19313 , \19314 , \19315 , \19316 , \19317 , \19318 , \19319 , \19320 ,
         \19321 , \19322 , \19323 , \19324 , \19325 , \19326 , \19327 , \19328 , \19329 , \19330 ,
         \19331 , \19332 , \19333 , \19334 , \19335 , \19336 , \19337 , \19338 , \19339 , \19340 ,
         \19341 , \19342 , \19343 , \19344 , \19345 , \19346 , \19347 , \19348 , \19349 , \19350 ,
         \19351 , \19352 , \19353 , \19354 , \19355 , \19356 , \19357 , \19358 , \19359 , \19360 ,
         \19361 , \19362 , \19363 , \19364 , \19365 , \19366 , \19367 , \19368 , \19369 , \19370 ,
         \19371 , \19372 , \19373 , \19374 , \19375 , \19376 , \19377 , \19378 , \19379 , \19380 ,
         \19381 , \19382 , \19383 , \19384 , \19385 , \19386 , \19387 , \19388 , \19389 , \19390 ,
         \19391 , \19392 , \19393 , \19394 , \19395 , \19396 , \19397 , \19398 , \19399 , \19400 ,
         \19401 , \19402 , \19403 , \19404 , \19405 , \19406 , \19407 , \19408 , \19409 , \19410 ,
         \19411 , \19412 , \19413 , \19414 , \19415 , \19416 , \19417 , \19418 , \19419 , \19420 ,
         \19421 , \19422 , \19423 , \19424 , \19425 , \19426 , \19427 , \19428 , \19429 , \19430 ,
         \19431 , \19432 , \19433 , \19434 , \19435 , \19436 , \19437 , \19438 , \19439 , \19440 ,
         \19441 , \19442 , \19443 , \19444 , \19445 , \19446 , \19447 , \19448 , \19449 , \19450 ,
         \19451 , \19452 , \19453 , \19454 , \19455 , \19456 , \19457 , \19458 , \19459 , \19460 ,
         \19461 , \19462 , \19463 , \19464 , \19465 , \19466 , \19467 , \19468 , \19469 , \19470 ,
         \19471 , \19472 , \19473 , \19474 , \19475 , \19476 , \19477 , \19478 , \19479 , \19480 ,
         \19481 , \19482 , \19483 , \19484 , \19485 , \19486 , \19487 , \19488 , \19489 , \19490 ,
         \19491 , \19492 , \19493 , \19494 , \19495 , \19496 , \19497 , \19498 , \19499 , \19500 ,
         \19501 , \19502 , \19503 , \19504 , \19505 , \19506 , \19507 , \19508 , \19509 , \19510 ,
         \19511 , \19512 , \19513 , \19514 , \19515 , \19516 , \19517 , \19518 , \19519 , \19520 ,
         \19521 , \19522 , \19523 , \19524 , \19525 , \19526 , \19527 , \19528 , \19529 , \19530 ,
         \19531 , \19532 , \19533 , \19534 , \19535 , \19536 , \19537 , \19538 , \19539 , \19540 ,
         \19541 , \19542 , \19543 , \19544 , \19545 , \19546 , \19547 , \19548 , \19549 , \19550 ,
         \19551 , \19552 , \19553 , \19554 , \19555 , \19556 , \19557 , \19558 , \19559 , \19560 ,
         \19561 , \19562 , \19563 , \19564 , \19565 , \19566 , \19567 , \19568 , \19569 , \19570 ,
         \19571 , \19572 , \19573 , \19574 , \19575 , \19576 , \19577 , \19578 , \19579 , \19580 ,
         \19581 , \19582 , \19583 , \19584 , \19585 , \19586 , \19587 , \19588 , \19589 , \19590 ,
         \19591 , \19592 , \19593 , \19594 , \19595 , \19596 , \19597 , \19598 , \19599 , \19600 ,
         \19601 , \19602 , \19603 , \19604 , \19605 , \19606 , \19607 , \19608 , \19609 , \19610 ,
         \19611 , \19612 , \19613 , \19614 , \19615 , \19616 , \19617 , \19618 , \19619 , \19620 ,
         \19621 , \19622 , \19623 , \19624 , \19625 , \19626 , \19627 , \19628 , \19629 , \19630 ,
         \19631 , \19632 , \19633 , \19634 , \19635 , \19636 , \19637 , \19638 , \19639 , \19640 ,
         \19641 , \19642 , \19643 , \19644 , \19645 , \19646 , \19647 , \19648 , \19649 , \19650 ,
         \19651 , \19652 , \19653 , \19654 , \19655 , \19656 , \19657 , \19658 , \19659 , \19660 ,
         \19661 , \19662 , \19663 , \19664 , \19665 , \19666 , \19667 , \19668 , \19669 , \19670 ,
         \19671 , \19672 , \19673 , \19674 , \19675 , \19676 , \19677 , \19678 , \19679 , \19680 ,
         \19681 , \19682 , \19683 , \19684 , \19685 , \19686 , \19687 , \19688 , \19689 , \19690 ,
         \19691 , \19692 , \19693 , \19694 , \19695 , \19696 , \19697 , \19698 , \19699 , \19700 ,
         \19701 , \19702 , \19703 , \19704 , \19705 , \19706 , \19707 , \19708 , \19709 , \19710 ,
         \19711 , \19712 , \19713 , \19714 , \19715 , \19716 , \19717 , \19718 , \19719 , \19720 ,
         \19721 , \19722 , \19723 , \19724 , \19725 , \19726 , \19727 , \19728 , \19729 , \19730 ,
         \19731 , \19732 , \19733 , \19734 , \19735 , \19736 , \19737 , \19738 , \19739 , \19740 ,
         \19741 , \19742 , \19743 , \19744 , \19745 , \19746 , \19747 , \19748 , \19749 , \19750 ,
         \19751 , \19752 , \19753 , \19754 , \19755 , \19756 , \19757 , \19758 , \19759 , \19760 ,
         \19761 , \19762 , \19763 , \19764 , \19765 , \19766 , \19767 , \19768 , \19769 , \19770 ,
         \19771 , \19772 , \19773 , \19774 , \19775 , \19776 , \19777 , \19778 , \19779 , \19780 ,
         \19781 , \19782 , \19783 , \19784 , \19785 , \19786 , \19787 , \19788 , \19789 , \19790 ,
         \19791 , \19792 , \19793 , \19794 , \19795 , \19796 , \19797 , \19798 , \19799 , \19800 ,
         \19801 , \19802 , \19803 , \19804 , \19805 , \19806 , \19807 , \19808 , \19809 , \19810 ,
         \19811 , \19812 , \19813 , \19814 , \19815 , \19816 , \19817 , \19818 , \19819 , \19820 ,
         \19821 , \19822 , \19823 , \19824 , \19825 , \19826 , \19827 , \19828 , \19829 , \19830 ,
         \19831 , \19832 , \19833 , \19834 , \19835 , \19836 , \19837 , \19838 , \19839 , \19840 ,
         \19841 , \19842 , \19843 , \19844 , \19845 , \19846 , \19847 , \19848 , \19849 , \19850 ,
         \19851 , \19852 , \19853 , \19854 , \19855 , \19856 , \19857 , \19858 , \19859 , \19860 ,
         \19861 , \19862 , \19863 , \19864 , \19865 , \19866 , \19867 , \19868 , \19869 , \19870 ,
         \19871 , \19872 , \19873 , \19874 , \19875 , \19876 , \19877 , \19878 , \19879 , \19880 ,
         \19881 , \19882 , \19883 , \19884 , \19885 , \19886 , \19887 , \19888 , \19889 , \19890 ,
         \19891 , \19892 , \19893 , \19894 , \19895 , \19896 , \19897 , \19898 , \19899 , \19900 ,
         \19901 , \19902 , \19903 , \19904 , \19905 , \19906 , \19907 , \19908 , \19909 , \19910 ,
         \19911 , \19912 , \19913 , \19914 , \19915 , \19916 , \19917 , \19918 , \19919 , \19920 ,
         \19921 , \19922 , \19923 , \19924 , \19925 , \19926 , \19927 , \19928 , \19929 , \19930 ,
         \19931 , \19932 , \19933 , \19934 , \19935 , \19936 , \19937 , \19938 , \19939 , \19940 ,
         \19941 , \19942 , \19943 , \19944 , \19945 , \19946 , \19947 , \19948 , \19949 , \19950 ,
         \19951 , \19952 , \19953 , \19954 , \19955 , \19956 , \19957 , \19958 , \19959 , \19960 ,
         \19961 , \19962 , \19963 , \19964 , \19965 , \19966 , \19967 , \19968 , \19969 , \19970 ,
         \19971 , \19972 , \19973 , \19974 , \19975 , \19976 , \19977 , \19978 , \19979 , \19980 ,
         \19981 , \19982 , \19983 , \19984 , \19985 , \19986 , \19987 , \19988 , \19989 , \19990 ,
         \19991 , \19992 , \19993 , \19994 , \19995 , \19996 , \19997 , \19998 , \19999 , \20000 ,
         \20001 , \20002 , \20003 , \20004 , \20005 , \20006 , \20007 , \20008 , \20009 , \20010 ,
         \20011 , \20012 , \20013 , \20014 , \20015 , \20016 , \20017 , \20018 , \20019 , \20020 ,
         \20021 , \20022 , \20023 , \20024 , \20025 , \20026 , \20027 , \20028 , \20029 , \20030 ,
         \20031 , \20032 , \20033 , \20034 , \20035 , \20036 , \20037 , \20038 , \20039 , \20040 ,
         \20041 , \20042 , \20043 , \20044 , \20045 , \20046 , \20047 , \20048 , \20049 , \20050 ,
         \20051 , \20052 , \20053 , \20054 , \20055 , \20056 , \20057 , \20058 , \20059 , \20060 ,
         \20061 , \20062 , \20063 , \20064 , \20065 , \20066 , \20067 , \20068 , \20069 , \20070 ,
         \20071 , \20072 , \20073 , \20074 , \20075 , \20076 , \20077 , \20078 , \20079 , \20080 ,
         \20081 , \20082 , \20083 , \20084 , \20085 , \20086 , \20087 , \20088 , \20089 , \20090 ,
         \20091 , \20092 , \20093 , \20094 , \20095 , \20096 , \20097 , \20098 , \20099 , \20100 ,
         \20101 , \20102 , \20103 , \20104 , \20105 , \20106 , \20107 , \20108 , \20109 , \20110 ,
         \20111 , \20112 , \20113 , \20114 , \20115 , \20116 , \20117 , \20118 , \20119 , \20120 ,
         \20121 , \20122 , \20123 , \20124 , \20125 , \20126 , \20127 , \20128 , \20129 , \20130 ,
         \20131 , \20132 , \20133 , \20134 , \20135 , \20136 , \20137 , \20138 , \20139 , \20140 ,
         \20141 , \20142 , \20143 , \20144 , \20145 , \20146 , \20147 , \20148 , \20149 , \20150 ,
         \20151 , \20152 , \20153 , \20154 , \20155 , \20156 , \20157 , \20158 , \20159 , \20160 ,
         \20161 , \20162 , \20163 , \20164 , \20165 , \20166 , \20167 , \20168 , \20169 , \20170 ,
         \20171 , \20172 , \20173 , \20174 , \20175 , \20176 , \20177 , \20178 , \20179 , \20180 ,
         \20181 , \20182 , \20183 , \20184 , \20185 , \20186 , \20187 , \20188 , \20189 , \20190 ,
         \20191 , \20192 , \20193 , \20194 , \20195 , \20196 , \20197 , \20198 , \20199 , \20200 ,
         \20201 , \20202 , \20203 , \20204 , \20205 , \20206 , \20207 , \20208 , \20209 , \20210 ,
         \20211 , \20212 , \20213 , \20214 , \20215 , \20216 , \20217 , \20218 , \20219 , \20220 ,
         \20221 , \20222 , \20223 , \20224 , \20225 , \20226 , \20227 , \20228 , \20229 , \20230 ,
         \20231 , \20232 , \20233 , \20234 , \20235 , \20236 , \20237 , \20238 , \20239 , \20240 ,
         \20241 , \20242 , \20243 , \20244 , \20245 , \20246 , \20247 , \20248 , \20249 , \20250 ,
         \20251 , \20252 , \20253 , \20254 , \20255 , \20256 , \20257 , \20258 , \20259 , \20260 ,
         \20261 , \20262 , \20263 , \20264 , \20265 , \20266 , \20267 , \20268 , \20269 , \20270 ,
         \20271 , \20272 , \20273 , \20274 , \20275 , \20276 , \20277 , \20278 , \20279 , \20280 ,
         \20281 , \20282 , \20283 , \20284 , \20285 , \20286 , \20287 , \20288 , \20289 , \20290 ,
         \20291 , \20292 , \20293 , \20294 , \20295 , \20296 , \20297 , \20298 , \20299 , \20300 ,
         \20301 , \20302 , \20303 , \20304 , \20305 , \20306 , \20307 , \20308 , \20309 , \20310 ,
         \20311 , \20312 , \20313 , \20314 , \20315 , \20316 , \20317 , \20318 , \20319 , \20320 ,
         \20321 , \20322 , \20323 , \20324 , \20325 , \20326 , \20327 , \20328 , \20329 , \20330 ,
         \20331 , \20332 , \20333 , \20334 , \20335 , \20336 , \20337 , \20338 , \20339 , \20340 ,
         \20341 , \20342 , \20343 , \20344 , \20345 , \20346 , \20347 , \20348 , \20349 , \20350 ,
         \20351 , \20352 , \20353 , \20354 , \20355 , \20356 , \20357 , \20358 , \20359 , \20360 ,
         \20361 , \20362 , \20363 , \20364 , \20365 , \20366 , \20367 , \20368 , \20369 , \20370 ,
         \20371 , \20372 , \20373 , \20374 , \20375 , \20376 , \20377 , \20378 , \20379 , \20380 ,
         \20381 , \20382 , \20383 , \20384 , \20385 , \20386 , \20387 , \20388 , \20389 , \20390 ,
         \20391 , \20392 , \20393 , \20394 , \20395 , \20396 , \20397 , \20398 , \20399 , \20400 ,
         \20401 , \20402 , \20403 , \20404 , \20405 , \20406 , \20407 , \20408 , \20409 , \20410 ,
         \20411 , \20412 , \20413 , \20414 , \20415 , \20416 , \20417 , \20418 , \20419 , \20420 ,
         \20421 , \20422 , \20423 , \20424 , \20425 , \20426 , \20427 , \20428 , \20429 , \20430 ,
         \20431 , \20432 , \20433 , \20434 , \20435 , \20436 , \20437 , \20438 , \20439 , \20440 ,
         \20441 , \20442 , \20443 , \20444 , \20445 , \20446 , \20447 , \20448 , \20449 , \20450 ,
         \20451 , \20452 , \20453 , \20454 , \20455 , \20456 , \20457 , \20458 , \20459 , \20460 ,
         \20461 , \20462 , \20463 , \20464 , \20465 , \20466 , \20467 , \20468 , \20469 , \20470 ,
         \20471 , \20472 , \20473 , \20474 , \20475 , \20476 , \20477 , \20478 , \20479 , \20480 ,
         \20481 , \20482 , \20483 , \20484 , \20485 , \20486 , \20487 , \20488 , \20489 , \20490 ,
         \20491 , \20492 , \20493 , \20494 , \20495 , \20496 , \20497 , \20498 , \20499 , \20500 ,
         \20501 , \20502 , \20503 , \20504 , \20505 , \20506 , \20507 , \20508 , \20509 , \20510 ,
         \20511 , \20512 , \20513 , \20514 , \20515 , \20516 , \20517 , \20518 , \20519 , \20520 ,
         \20521 , \20522 , \20523 , \20524 , \20525 , \20526 , \20527 , \20528 , \20529 , \20530 ,
         \20531 , \20532 , \20533 , \20534 , \20535 , \20536 , \20537 , \20538 , \20539 , \20540 ,
         \20541 , \20542 , \20543 , \20544 , \20545 , \20546 , \20547 , \20548 , \20549 , \20550 ,
         \20551 , \20552 , \20553 , \20554 , \20555 , \20556 , \20557 , \20558 , \20559 , \20560 ,
         \20561 , \20562 , \20563 , \20564 , \20565 , \20566 , \20567 , \20568 , \20569 , \20570 ,
         \20571 , \20572 , \20573 , \20574 , \20575 , \20576 , \20577 , \20578 , \20579 , \20580 ,
         \20581 , \20582 , \20583 , \20584 , \20585 , \20586 , \20587 , \20588 , \20589 , \20590 ,
         \20591 , \20592 , \20593 , \20594 , \20595 , \20596 , \20597 , \20598 , \20599 , \20600 ,
         \20601 , \20602 , \20603 , \20604 , \20605 , \20606 , \20607 , \20608 , \20609 , \20610 ,
         \20611 , \20612 , \20613 , \20614 , \20615 , \20616 , \20617 , \20618 , \20619 , \20620 ,
         \20621 , \20622 , \20623 , \20624 , \20625 , \20626 , \20627 , \20628 , \20629 , \20630 ,
         \20631 , \20632 , \20633 , \20634 , \20635 , \20636 , \20637 , \20638 , \20639 , \20640 ,
         \20641 , \20642 , \20643 , \20644 , \20645 , \20646 , \20647 , \20648 , \20649 , \20650 ,
         \20651 , \20652 , \20653 , \20654 , \20655 , \20656 , \20657 , \20658 , \20659 , \20660 ,
         \20661 , \20662 , \20663 , \20664 , \20665 , \20666 , \20667 , \20668 , \20669 , \20670 ,
         \20671 , \20672 , \20673 , \20674 , \20675 , \20676 , \20677 , \20678 , \20679 , \20680 ,
         \20681 , \20682 , \20683 , \20684 , \20685 , \20686 , \20687 , \20688 , \20689 , \20690 ,
         \20691 , \20692 , \20693 , \20694 , \20695 , \20696 , \20697 , \20698 , \20699 , \20700 ,
         \20701 , \20702 , \20703 , \20704 , \20705 , \20706 , \20707 , \20708 , \20709 , \20710 ,
         \20711 , \20712 , \20713 , \20714 , \20715 , \20716 , \20717 , \20718 , \20719 , \20720 ,
         \20721 , \20722 , \20723 , \20724 , \20725 , \20726 , \20727 , \20728 , \20729 , \20730 ,
         \20731 , \20732 , \20733 , \20734 , \20735 , \20736 , \20737 , \20738 , \20739 , \20740 ,
         \20741 , \20742 , \20743 , \20744 , \20745 , \20746 , \20747 , \20748 , \20749 , \20750 ,
         \20751 , \20752 , \20753 , \20754 , \20755 , \20756 , \20757 , \20758 , \20759 , \20760 ,
         \20761 , \20762 , \20763 , \20764 , \20765 , \20766 , \20767 , \20768 , \20769 , \20770 ,
         \20771 , \20772 , \20773 , \20774 , \20775 , \20776 , \20777 , \20778 , \20779 , \20780 ,
         \20781 , \20782 , \20783 , \20784 , \20785 , \20786 , \20787 , \20788 , \20789 , \20790 ,
         \20791 , \20792 , \20793 , \20794 , \20795 , \20796 , \20797 , \20798 , \20799 , \20800 ,
         \20801 , \20802 , \20803 , \20804 , \20805 , \20806 , \20807 , \20808 , \20809 , \20810 ,
         \20811 , \20812 , \20813 , \20814 , \20815 , \20816 , \20817 , \20818 , \20819 , \20820 ,
         \20821 , \20822 , \20823 , \20824 , \20825 , \20826 , \20827 , \20828 , \20829 , \20830 ,
         \20831 , \20832 , \20833 , \20834 , \20835 , \20836 , \20837 , \20838 , \20839 , \20840 ,
         \20841 , \20842 , \20843 , \20844 , \20845 , \20846 , \20847 , \20848 , \20849 , \20850 ,
         \20851 , \20852 , \20853 , \20854 , \20855 , \20856 , \20857 , \20858 , \20859 , \20860 ,
         \20861 , \20862 , \20863 , \20864 , \20865 , \20866 , \20867 , \20868 , \20869 , \20870 ,
         \20871 , \20872 , \20873 , \20874 , \20875 , \20876 , \20877 , \20878 , \20879 , \20880 ,
         \20881 , \20882 , \20883 , \20884 , \20885 , \20886 , \20887 , \20888 , \20889 , \20890 ,
         \20891 , \20892 , \20893 , \20894 , \20895 , \20896 , \20897 , \20898 , \20899 , \20900 ,
         \20901 , \20902 , \20903 , \20904 , \20905 , \20906 , \20907 , \20908 , \20909 , \20910 ,
         \20911 , \20912 , \20913 , \20914 , \20915 , \20916 , \20917 , \20918 , \20919 , \20920 ,
         \20921 , \20922 , \20923 , \20924 , \20925 , \20926 , \20927 , \20928 , \20929 , \20930 ,
         \20931 , \20932 , \20933 , \20934 , \20935 , \20936 , \20937 , \20938 , \20939 , \20940 ,
         \20941 , \20942 , \20943 , \20944 , \20945 , \20946 , \20947 , \20948 , \20949 , \20950 ,
         \20951 , \20952 , \20953 , \20954 , \20955 , \20956 , \20957 , \20958 , \20959 , \20960 ,
         \20961 , \20962 , \20963 , \20964 , \20965 , \20966 , \20967 , \20968 , \20969 , \20970 ,
         \20971 , \20972 , \20973 , \20974 , \20975 , \20976 , \20977 , \20978 , \20979 , \20980 ,
         \20981 , \20982 , \20983 , \20984 , \20985 , \20986 , \20987 , \20988 , \20989 , \20990 ,
         \20991 , \20992 , \20993 , \20994 , \20995 , \20996 , \20997 , \20998 , \20999 , \21000 ,
         \21001 , \21002 , \21003 , \21004 , \21005 , \21006 , \21007 , \21008 , \21009 , \21010 ,
         \21011 , \21012 , \21013 , \21014 , \21015 , \21016 , \21017 , \21018 , \21019 , \21020 ,
         \21021 , \21022 , \21023 , \21024 , \21025 , \21026 , \21027 , \21028 , \21029 , \21030 ,
         \21031 , \21032 , \21033 , \21034 , \21035 , \21036 , \21037 , \21038 , \21039 , \21040 ,
         \21041 , \21042 , \21043 , \21044 , \21045 , \21046 , \21047 , \21048 , \21049 , \21050 ,
         \21051 , \21052 , \21053 , \21054 , \21055 , \21056 , \21057 , \21058 , \21059 , \21060 ,
         \21061 , \21062 , \21063 , \21064 , \21065 , \21066 , \21067 , \21068 , \21069 , \21070 ,
         \21071 , \21072 , \21073 , \21074 , \21075 , \21076 , \21077 , \21078 , \21079 , \21080 ,
         \21081 , \21082 , \21083 , \21084 , \21085 , \21086 , \21087 , \21088 , \21089 , \21090 ,
         \21091 , \21092 , \21093 , \21094 , \21095 , \21096 , \21097 , \21098 , \21099 , \21100 ,
         \21101 , \21102 , \21103 , \21104 , \21105 , \21106 , \21107 , \21108 , \21109 , \21110 ,
         \21111 , \21112 , \21113 , \21114 , \21115 , \21116 , \21117 , \21118 , \21119 , \21120 ,
         \21121 , \21122 , \21123 , \21124 , \21125 , \21126 , \21127 , \21128 , \21129 , \21130 ,
         \21131 , \21132 , \21133 , \21134 , \21135 , \21136 , \21137 , \21138 , \21139 , \21140 ,
         \21141 , \21142 , \21143 , \21144 , \21145 , \21146 , \21147 , \21148 , \21149 , \21150 ,
         \21151 , \21152 , \21153 , \21154 , \21155 , \21156 , \21157 , \21158 , \21159 , \21160 ,
         \21161 , \21162 , \21163 , \21164 , \21165 , \21166 , \21167 , \21168 , \21169 , \21170 ,
         \21171 , \21172 , \21173 , \21174 , \21175 , \21176 , \21177 , \21178 , \21179 , \21180 ,
         \21181 , \21182 , \21183 , \21184 , \21185 , \21186 , \21187 , \21188 , \21189 , \21190 ,
         \21191 , \21192 , \21193 , \21194 , \21195 , \21196 , \21197 , \21198 , \21199 , \21200 ,
         \21201 , \21202 , \21203 , \21204 , \21205 , \21206 , \21207 , \21208 , \21209 , \21210 ,
         \21211 , \21212 , \21213 , \21214 , \21215 , \21216 , \21217 , \21218 , \21219 , \21220 ,
         \21221 , \21222 , \21223 , \21224 , \21225 , \21226 , \21227 , \21228 , \21229 , \21230 ,
         \21231 , \21232 , \21233 , \21234 , \21235 , \21236 , \21237 , \21238 , \21239 , \21240 ,
         \21241 , \21242 , \21243 , \21244 , \21245 , \21246 , \21247 , \21248 , \21249 , \21250 ,
         \21251 , \21252 , \21253 , \21254 , \21255 , \21256 , \21257 , \21258 , \21259 , \21260 ,
         \21261 , \21262 , \21263 , \21264 , \21265 , \21266 , \21267 , \21268 , \21269 , \21270 ,
         \21271 , \21272 , \21273 , \21274 , \21275 , \21276 , \21277 , \21278 , \21279 , \21280 ,
         \21281 , \21282 , \21283 , \21284 , \21285 , \21286 , \21287 , \21288 , \21289 , \21290 ,
         \21291 , \21292 , \21293 , \21294 , \21295 , \21296 , \21297 , \21298 , \21299 , \21300 ,
         \21301 , \21302 , \21303 , \21304 , \21305 , \21306 , \21307 , \21308 , \21309 , \21310 ,
         \21311 , \21312 , \21313 , \21314 , \21315 , \21316 , \21317 , \21318 , \21319 , \21320 ,
         \21321 , \21322 , \21323 , \21324 , \21325 , \21326 , \21327 , \21328 , \21329 , \21330 ,
         \21331 , \21332 , \21333 , \21334 , \21335 , \21336 , \21337 , \21338 , \21339 , \21340 ,
         \21341 , \21342 , \21343 , \21344 , \21345 , \21346 , \21347 , \21348 , \21349 , \21350 ,
         \21351 , \21352 , \21353 , \21354 , \21355 , \21356 , \21357 , \21358 , \21359 , \21360 ,
         \21361 , \21362 , \21363 , \21364 , \21365 , \21366 , \21367 , \21368 , \21369 , \21370_nGac4c ,
         \21371 , \21372 , \21373 , \21374 , \21375 , \21376 , \21377 , \21378 , \21379 , \21380 ,
         \21381 , \21382 , \21383 , \21384 , \21385 , \21386 , \21387 , \21388 , \21389 , \21390 ,
         \21391 , \21392 , \21393 , \21394 , \21395 , \21396 , \21397 , \21398 , \21399 , \21400 ,
         \21401 , \21402 , \21403 , \21404 , \21405 , \21406 , \21407 , \21408 , \21409 , \21410 ,
         \21411 , \21412 , \21413 , \21414 , \21415 , \21416 , \21417 , \21418 , \21419 , \21420 ,
         \21421 , \21422 , \21423 , \21424 , \21425 , \21426 , \21427 , \21428 , \21429 , \21430 ,
         \21431 , \21432 , \21433 , \21434 , \21435 , \21436 , \21437 , \21438 , \21439 , \21440 ,
         \21441 , \21442 , \21443 , \21444 , \21445 , \21446 , \21447 , \21448 , \21449 , \21450 ,
         \21451 , \21452 , \21453 , \21454 , \21455 , \21456 , \21457 , \21458 , \21459 , \21460 ,
         \21461 , \21462 , \21463 , \21464 , \21465 , \21466 , \21467 , \21468 , \21469 , \21470 ,
         \21471 , \21472 , \21473 , \21474 , \21475 , \21476 , \21477 , \21478 , \21479 , \21480 ,
         \21481 , \21482 , \21483 , \21484 , \21485 , \21486 , \21487 , \21488 , \21489 , \21490 ,
         \21491 , \21492 , \21493 , \21494 , \21495 , \21496 , \21497 , \21498 , \21499 , \21500 ,
         \21501 , \21502 , \21503 , \21504 , \21505 , \21506 , \21507 , \21508 , \21509 , \21510 ,
         \21511 , \21512 , \21513 , \21514 , \21515 , \21516 , \21517 , \21518 , \21519 , \21520 ,
         \21521 , \21522 , \21523 , \21524 , \21525 , \21526 , \21527 , \21528 , \21529 , \21530 ,
         \21531 , \21532 , \21533 , \21534 , \21535 , \21536 , \21537 , \21538 , \21539 , \21540 ,
         \21541 , \21542 , \21543 , \21544 , \21545 , \21546 , \21547 , \21548 , \21549 , \21550 ,
         \21551 , \21552 , \21553 , \21554 , \21555 , \21556 , \21557 , \21558 , \21559 , \21560 ,
         \21561 , \21562 , \21563 , \21564 , \21565 , \21566 , \21567 , \21568 , \21569 , \21570 ,
         \21571 , \21572 , \21573 , \21574 , \21575 , \21576 , \21577 , \21578 , \21579 , \21580 ,
         \21581 , \21582 , \21583 , \21584 , \21585 , \21586 , \21587 , \21588 , \21589 , \21590 ,
         \21591 , \21592 , \21593 , \21594 , \21595 , \21596 , \21597 , \21598 , \21599 , \21600 ,
         \21601 , \21602 , \21603 , \21604 , \21605 , \21606 , \21607 , \21608 , \21609 , \21610 ,
         \21611 , \21612 , \21613 , \21614 , \21615 , \21616 , \21617 , \21618 , \21619 , \21620 ,
         \21621 , \21622 , \21623 , \21624 , \21625 , \21626 , \21627 , \21628 , \21629 , \21630 ,
         \21631 , \21632 , \21633 , \21634 , \21635 , \21636 , \21637 , \21638 , \21639 , \21640 ,
         \21641 , \21642 , \21643 , \21644 , \21645 , \21646 , \21647 , \21648 , \21649 , \21650 ,
         \21651 , \21652 , \21653 , \21654 , \21655 , \21656 , \21657 , \21658 , \21659 , \21660 ,
         \21661 , \21662 , \21663 , \21664 , \21665 , \21666 , \21667 , \21668 , \21669 , \21670 ,
         \21671 , \21672 , \21673 , \21674 , \21675 , \21676 , \21677 , \21678 , \21679 , \21680 ,
         \21681 , \21682 , \21683 , \21684 , \21685 , \21686 , \21687 , \21688 , \21689 , \21690 ,
         \21691 , \21692 , \21693 , \21694 , \21695 , \21696 , \21697 , \21698 , \21699 , \21700 ,
         \21701 , \21702 , \21703 , \21704 , \21705 , \21706 , \21707 , \21708 , \21709 , \21710 ,
         \21711 , \21712 , \21713 , \21714 , \21715 , \21716 , \21717 , \21718 , \21719 , \21720 ,
         \21721 , \21722 , \21723 , \21724 , \21725 , \21726 , \21727 , \21728 , \21729 , \21730 ,
         \21731 , \21732 , \21733 , \21734 , \21735 , \21736 , \21737 , \21738 , \21739 , \21740 ,
         \21741 , \21742 , \21743 , \21744 , \21745 , \21746 , \21747 , \21748 , \21749 , \21750 ,
         \21751 , \21752 , \21753 , \21754 , \21755 , \21756 , \21757 , \21758 , \21759 , \21760 ,
         \21761 , \21762 , \21763 , \21764 , \21765 , \21766 , \21767 , \21768 , \21769 , \21770 ,
         \21771 , \21772 , \21773 , \21774 , \21775 , \21776 , \21777 , \21778 , \21779 , \21780 ,
         \21781 , \21782 , \21783 , \21784 , \21785 , \21786 , \21787 , \21788 , \21789 , \21790 ,
         \21791 , \21792 , \21793 , \21794 , \21795 , \21796 , \21797 , \21798 , \21799 , \21800 ,
         \21801 , \21802 , \21803 , \21804 , \21805 , \21806 , \21807 , \21808 , \21809 , \21810 ,
         \21811 , \21812 , \21813 , \21814 , \21815 , \21816 , \21817 , \21818 , \21819 , \21820 ,
         \21821 , \21822 , \21823 , \21824 , \21825 , \21826 , \21827 , \21828 , \21829 , \21830 ,
         \21831 , \21832 , \21833 , \21834 , \21835 , \21836 , \21837 , \21838 , \21839 , \21840 ,
         \21841 , \21842 , \21843 , \21844 , \21845 , \21846 , \21847 , \21848 , \21849 , \21850 ,
         \21851 , \21852 , \21853 , \21854 , \21855 , \21856 , \21857 , \21858 , \21859 , \21860 ,
         \21861 , \21862 , \21863 , \21864 , \21865 , \21866 , \21867 , \21868 , \21869 , \21870 ,
         \21871 , \21872 , \21873 , \21874 , \21875 , \21876 , \21877 , \21878 , \21879 , \21880 ,
         \21881 , \21882 , \21883 , \21884 , \21885 , \21886 , \21887 , \21888 , \21889 , \21890 ,
         \21891 , \21892 , \21893 , \21894 , \21895 , \21896 , \21897 , \21898 , \21899 , \21900 ,
         \21901 , \21902 , \21903 , \21904 , \21905 , \21906 , \21907 , \21908 , \21909 , \21910 ,
         \21911 , \21912 , \21913 , \21914 , \21915 , \21916 , \21917 , \21918 , \21919 , \21920 ,
         \21921 , \21922 , \21923 , \21924 , \21925 , \21926 , \21927 , \21928 , \21929 , \21930 ,
         \21931 , \21932 , \21933 , \21934 , \21935 , \21936 , \21937 , \21938 , \21939 , \21940 ,
         \21941 , \21942 , \21943 , \21944 , \21945 , \21946 , \21947 , \21948 , \21949 , \21950 ,
         \21951 , \21952 , \21953 , \21954 , \21955 , \21956 , \21957 , \21958 , \21959 , \21960 ,
         \21961 , \21962 , \21963 , \21964 , \21965 , \21966 , \21967 , \21968 , \21969 , \21970 ,
         \21971 , \21972 , \21973 , \21974 , \21975 , \21976 , \21977 , \21978 , \21979 , \21980 ,
         \21981 , \21982 , \21983 , \21984 , \21985 , \21986 , \21987 , \21988 , \21989 , \21990 ,
         \21991 , \21992 , \21993 , \21994 , \21995 , \21996 , \21997 , \21998 , \21999 , \22000 ,
         \22001 , \22002 , \22003 , \22004 , \22005 , \22006 , \22007 , \22008 , \22009 , \22010 ,
         \22011 , \22012 , \22013 , \22014 , \22015 , \22016 , \22017 , \22018 , \22019 , \22020 ,
         \22021 , \22022 , \22023 , \22024 , \22025 , \22026 , \22027 , \22028 , \22029 , \22030 ,
         \22031 , \22032 , \22033 , \22034 , \22035 , \22036 , \22037 , \22038 , \22039 , \22040 ,
         \22041 , \22042 , \22043 , \22044 , \22045 , \22046 , \22047 , \22048 , \22049 , \22050 ,
         \22051 , \22052 , \22053 , \22054 , \22055 , \22056 , \22057 , \22058 , \22059 , \22060 ,
         \22061 , \22062 , \22063 , \22064 , \22065 , \22066 , \22067 , \22068 , \22069 , \22070 ,
         \22071 , \22072 , \22073 , \22074 , \22075 , \22076 , \22077 , \22078 , \22079 , \22080 ,
         \22081 , \22082 , \22083 , \22084 , \22085 , \22086 , \22087 , \22088 , \22089 , \22090 ,
         \22091 , \22092 , \22093 , \22094 , \22095 , \22096 , \22097 , \22098 , \22099 , \22100 ,
         \22101 , \22102 , \22103 , \22104 , \22105 , \22106 , \22107 , \22108 , \22109 , \22110 ,
         \22111 , \22112 , \22113 , \22114 , \22115 , \22116 , \22117 , \22118 , \22119 , \22120 ,
         \22121 , \22122 , \22123 , \22124 , \22125 , \22126 , \22127 , \22128 , \22129 , \22130 ,
         \22131 , \22132 , \22133 , \22134 , \22135 , \22136 , \22137 , \22138 , \22139 , \22140 ,
         \22141 , \22142 , \22143 , \22144 , \22145 , \22146 , \22147 , \22148 , \22149 , \22150 ,
         \22151 , \22152 , \22153 , \22154 , \22155 , \22156 , \22157 , \22158 , \22159 , \22160 ,
         \22161 , \22162 , \22163 , \22164 , \22165 , \22166 , \22167 , \22168 , \22169 , \22170 ,
         \22171 , \22172 , \22173 , \22174 , \22175 , \22176 , \22177 , \22178 , \22179 , \22180 ,
         \22181 , \22182 , \22183 , \22184 , \22185 , \22186 , \22187 , \22188 , \22189 , \22190 ,
         \22191 , \22192 , \22193 , \22194 , \22195 , \22196 , \22197 , \22198 , \22199 , \22200 ,
         \22201 , \22202 , \22203 , \22204 , \22205 , \22206 , \22207 , \22208 , \22209 , \22210 ,
         \22211 , \22212 , \22213 , \22214 , \22215 , \22216 , \22217 , \22218 , \22219 , \22220 ,
         \22221 , \22222 , \22223 , \22224 , \22225 , \22226 , \22227 , \22228 , \22229 , \22230 ,
         \22231 , \22232 , \22233 , \22234 , \22235 , \22236 , \22237 , \22238 , \22239 , \22240 ,
         \22241 , \22242 , \22243 , \22244 , \22245 , \22246 , \22247 , \22248 , \22249 , \22250 ,
         \22251 , \22252 , \22253 , \22254 , \22255 , \22256 , \22257 , \22258 , \22259 , \22260 ,
         \22261 , \22262 , \22263 , \22264 , \22265 , \22266 , \22267 , \22268 , \22269 , \22270 ,
         \22271 , \22272 , \22273 , \22274 , \22275 , \22276 , \22277 , \22278 , \22279 , \22280 ,
         \22281 , \22282 , \22283 , \22284 , \22285 , \22286 , \22287 , \22288 , \22289 , \22290 ,
         \22291 , \22292 , \22293 , \22294 , \22295 , \22296 , \22297 , \22298 , \22299 , \22300 ,
         \22301 , \22302 , \22303 , \22304 , \22305 , \22306 , \22307 , \22308 , \22309 , \22310 ,
         \22311 , \22312 , \22313 , \22314 , \22315 , \22316 , \22317 , \22318 , \22319 , \22320 ,
         \22321 , \22322 , \22323 , \22324 , \22325 , \22326 , \22327 , \22328 , \22329 , \22330 ,
         \22331 , \22332 , \22333 , \22334 , \22335 , \22336 , \22337 , \22338 , \22339 , \22340 ,
         \22341 , \22342 , \22343 , \22344 , \22345 , \22346 , \22347 , \22348 , \22349 , \22350 ,
         \22351 , \22352 , \22353 , \22354 , \22355 , \22356 , \22357 , \22358 , \22359 , \22360 ,
         \22361 , \22362 , \22363 , \22364 , \22365 , \22366 , \22367 , \22368 , \22369 , \22370 ,
         \22371 , \22372 , \22373 , \22374 , \22375 , \22376 , \22377 , \22378 , \22379 , \22380 ,
         \22381 , \22382 , \22383 , \22384 , \22385 , \22386 , \22387 , \22388 , \22389 , \22390 ,
         \22391 , \22392 , \22393 , \22394 , \22395 , \22396 , \22397 , \22398 , \22399 , \22400 ,
         \22401 , \22402 , \22403 , \22404 , \22405 , \22406 , \22407 , \22408 , \22409 , \22410 ,
         \22411 , \22412 , \22413 , \22414 , \22415 , \22416 , \22417 , \22418 , \22419 , \22420 ,
         \22421 , \22422 , \22423 , \22424 , \22425 , \22426 , \22427 , \22428 , \22429 , \22430 ,
         \22431 , \22432 , \22433 , \22434 , \22435 , \22436 , \22437 , \22438 , \22439 , \22440 ,
         \22441 , \22442 , \22443 , \22444 , \22445 , \22446 , \22447 , \22448 , \22449 , \22450 ,
         \22451 , \22452 , \22453 , \22454 , \22455 , \22456 , \22457 , \22458 , \22459 , \22460 ,
         \22461 , \22462 , \22463 , \22464 , \22465 , \22466 , \22467 , \22468 , \22469 , \22470 ,
         \22471 , \22472 , \22473 , \22474 , \22475 , \22476 , \22477 , \22478 , \22479 , \22480 ,
         \22481 , \22482 , \22483 , \22484 , \22485 , \22486 , \22487 , \22488 , \22489 , \22490 ,
         \22491 , \22492 , \22493 , \22494 , \22495 , \22496 , \22497 , \22498 , \22499 , \22500 ,
         \22501 , \22502 , \22503 , \22504 , \22505 , \22506 , \22507 , \22508 , \22509 , \22510 ,
         \22511 , \22512 , \22513 , \22514 , \22515 , \22516 , \22517 , \22518 , \22519 , \22520 ,
         \22521 , \22522 , \22523 , \22524 , \22525 , \22526 , \22527 , \22528 , \22529 , \22530 ,
         \22531 , \22532 , \22533 , \22534 , \22535 , \22536 , \22537 , \22538 , \22539 , \22540 ,
         \22541 , \22542 , \22543 , \22544 , \22545 , \22546 , \22547 , \22548 , \22549 , \22550 ,
         \22551 , \22552 , \22553 , \22554 , \22555 , \22556 , \22557 , \22558 , \22559 , \22560 ,
         \22561 , \22562 , \22563 , \22564 , \22565 , \22566 , \22567 , \22568 , \22569 , \22570 ,
         \22571 , \22572 , \22573 , \22574 , \22575 , \22576 , \22577 , \22578 , \22579 , \22580 ,
         \22581 , \22582 , \22583 , \22584 , \22585 , \22586 , \22587 , \22588 , \22589 , \22590 ,
         \22591 , \22592 , \22593 , \22594 , \22595 , \22596 , \22597 , \22598 , \22599 , \22600 ,
         \22601 , \22602 , \22603 , \22604 , \22605 , \22606 , \22607 , \22608 , \22609 , \22610 ,
         \22611 , \22612 , \22613 , \22614 , \22615 , \22616 , \22617 , \22618 , \22619 , \22620 ,
         \22621 , \22622 , \22623 , \22624 , \22625 , \22626 , \22627 , \22628 , \22629 , \22630 ,
         \22631 , \22632 , \22633 , \22634 , \22635 , \22636 , \22637 , \22638 , \22639 , \22640 ,
         \22641 , \22642 , \22643 , \22644 , \22645 , \22646 , \22647 , \22648 , \22649 , \22650 ,
         \22651 , \22652 , \22653 , \22654 , \22655 , \22656 , \22657 , \22658 , \22659 , \22660 ,
         \22661 , \22662 , \22663 , \22664 , \22665 , \22666 , \22667 , \22668 , \22669 , \22670 ,
         \22671 , \22672 , \22673 , \22674 , \22675 , \22676 , \22677 , \22678 , \22679 , \22680 ,
         \22681 , \22682 , \22683 , \22684 , \22685 , \22686 , \22687 , \22688 , \22689 , \22690 ,
         \22691 , \22692 , \22693 , \22694 , \22695 , \22696 , \22697 , \22698 , \22699 , \22700 ,
         \22701 , \22702 , \22703 , \22704 , \22705 , \22706 , \22707 , \22708 , \22709 , \22710 ,
         \22711 , \22712 , \22713 , \22714 , \22715 , \22716 , \22717 , \22718 , \22719 , \22720 ,
         \22721 , \22722 , \22723 , \22724 , \22725 , \22726 , \22727 , \22728 , \22729 , \22730 ,
         \22731 , \22732 , \22733 , \22734 , \22735 , \22736 , \22737 , \22738 , \22739 , \22740 ,
         \22741 , \22742 , \22743 , \22744 , \22745 , \22746 , \22747 , \22748 , \22749 , \22750 ,
         \22751 , \22752 , \22753 , \22754 , \22755 , \22756 , \22757 , \22758 , \22759 , \22760 ,
         \22761 , \22762 , \22763 , \22764 , \22765 , \22766 , \22767 , \22768 , \22769 , \22770 ,
         \22771 , \22772 , \22773 , \22774 , \22775 , \22776 , \22777 , \22778 , \22779 , \22780 ,
         \22781 , \22782 , \22783 , \22784 , \22785 , \22786 , \22787 , \22788 , \22789 , \22790 ,
         \22791 , \22792 , \22793 , \22794 , \22795 , \22796 , \22797 , \22798 , \22799 , \22800 ,
         \22801 , \22802 , \22803 , \22804 , \22805 , \22806 , \22807 , \22808 , \22809 , \22810 ,
         \22811 , \22812 , \22813 , \22814 , \22815 , \22816 , \22817 , \22818 , \22819 , \22820 ,
         \22821 , \22822 , \22823 , \22824 , \22825 , \22826 , \22827 , \22828 , \22829 , \22830 ,
         \22831 , \22832 , \22833 , \22834 , \22835 , \22836 , \22837 , \22838 , \22839 , \22840 ,
         \22841 , \22842 , \22843 , \22844 , \22845 , \22846 , \22847 , \22848 , \22849 , \22850 ,
         \22851 , \22852 , \22853 , \22854 , \22855 , \22856 , \22857 , \22858 , \22859 , \22860 ,
         \22861 , \22862 , \22863 , \22864 , \22865 , \22866 , \22867 , \22868 , \22869 , \22870 ,
         \22871 , \22872 , \22873 , \22874 , \22875 , \22876 , \22877 , \22878 , \22879 , \22880 ,
         \22881 , \22882 , \22883 , \22884 , \22885 , \22886 , \22887 , \22888 , \22889 , \22890 ,
         \22891 , \22892 , \22893 , \22894 , \22895 , \22896 , \22897 , \22898 , \22899 , \22900 ,
         \22901 , \22902 , \22903 , \22904 , \22905 , \22906 , \22907 , \22908 , \22909 , \22910 ,
         \22911 , \22912 , \22913 , \22914 , \22915 , \22916 , \22917 , \22918 , \22919 , \22920 ,
         \22921 , \22922 , \22923 , \22924 , \22925 , \22926 , \22927 , \22928 , \22929 , \22930 ,
         \22931 , \22932 , \22933 , \22934 , \22935 , \22936 , \22937 , \22938 , \22939 , \22940 ,
         \22941 , \22942 , \22943 , \22944 , \22945 , \22946 , \22947 , \22948 , \22949 , \22950 ,
         \22951 , \22952 , \22953 , \22954 , \22955 , \22956 , \22957 , \22958 , \22959 , \22960 ,
         \22961 , \22962 , \22963 , \22964 , \22965 , \22966 , \22967 , \22968 , \22969 , \22970 ,
         \22971 , \22972 , \22973 , \22974 , \22975 , \22976 , \22977 , \22978 , \22979 , \22980 ,
         \22981 , \22982 , \22983 , \22984 , \22985 , \22986 , \22987 , \22988 , \22989 , \22990 ,
         \22991 , \22992 , \22993 , \22994 , \22995 , \22996 , \22997 , \22998 , \22999 , \23000 ,
         \23001 , \23002 , \23003 , \23004 , \23005 , \23006 , \23007 , \23008 , \23009 , \23010 ,
         \23011 , \23012 , \23013 , \23014 , \23015 , \23016 , \23017 , \23018 , \23019 , \23020 ,
         \23021 , \23022 , \23023 , \23024 , \23025 , \23026 , \23027 , \23028 , \23029 , \23030 ,
         \23031 , \23032 , \23033 , \23034 , \23035 , \23036 , \23037 , \23038 , \23039 , \23040 ,
         \23041 , \23042 , \23043 , \23044 , \23045 , \23046 , \23047 , \23048 , \23049 , \23050 ,
         \23051 , \23052 , \23053 , \23054 , \23055 , \23056 , \23057 , \23058 , \23059 , \23060 ,
         \23061 , \23062 , \23063 , \23064 , \23065 , \23066 , \23067 , \23068 , \23069 , \23070 ,
         \23071 , \23072 , \23073 , \23074 , \23075 , \23076 , \23077 , \23078 , \23079 , \23080 ,
         \23081 , \23082 , \23083 , \23084 , \23085 , \23086 , \23087 , \23088 , \23089 , \23090 ,
         \23091 , \23092 , \23093 , \23094 , \23095 , \23096 , \23097 , \23098 , \23099 , \23100 ,
         \23101 , \23102 , \23103 , \23104 , \23105 , \23106 , \23107 , \23108 , \23109 , \23110 ,
         \23111 , \23112 , \23113 , \23114 , \23115 , \23116 , \23117 , \23118 , \23119 , \23120 ,
         \23121 , \23122 , \23123 , \23124 , \23125 , \23126 , \23127 , \23128 , \23129 , \23130 ,
         \23131 , \23132 , \23133 , \23134 , \23135 , \23136 , \23137 , \23138 , \23139 , \23140 ,
         \23141 , \23142 , \23143 , \23144 , \23145 , \23146 , \23147 , \23148 , \23149 , \23150 ,
         \23151 , \23152 , \23153 , \23154 , \23155 , \23156 , \23157 , \23158 , \23159 , \23160 ,
         \23161 , \23162 , \23163 , \23164 , \23165 , \23166 , \23167 , \23168 , \23169 , \23170 ,
         \23171 , \23172 , \23173 , \23174 , \23175 , \23176 , \23177 , \23178 , \23179 , \23180 ,
         \23181 , \23182 , \23183 , \23184 , \23185 , \23186 , \23187 , \23188 , \23189 , \23190 ,
         \23191 , \23192 , \23193 , \23194 , \23195 , \23196 , \23197 , \23198 , \23199 , \23200 ,
         \23201 , \23202 , \23203 , \23204 , \23205 , \23206 , \23207 , \23208 , \23209 , \23210 ,
         \23211 , \23212 , \23213 , \23214 , \23215 , \23216 , \23217 , \23218 , \23219 , \23220 ,
         \23221 , \23222 , \23223 , \23224 , \23225 , \23226 , \23227 , \23228 , \23229 , \23230 ,
         \23231 , \23232 , \23233 , \23234 , \23235 , \23236 , \23237 , \23238 , \23239 , \23240 ,
         \23241 , \23242 , \23243 , \23244 , \23245 , \23246 , \23247 , \23248 , \23249 , \23250 ,
         \23251 , \23252 , \23253 , \23254 , \23255 , \23256 , \23257 , \23258 , \23259 , \23260 ,
         \23261 , \23262 , \23263 , \23264 , \23265 , \23266 , \23267 , \23268 , \23269 , \23270 ,
         \23271 , \23272 , \23273 , \23274 , \23275 , \23276 , \23277 , \23278 , \23279 , \23280 ,
         \23281 , \23282 , \23283 , \23284 , \23285 , \23286 , \23287 , \23288 , \23289 , \23290 ,
         \23291 , \23292 , \23293 , \23294 , \23295 , \23296 , \23297 , \23298 , \23299 , \23300 ,
         \23301 , \23302 , \23303 , \23304 , \23305 , \23306 , \23307 , \23308 , \23309 , \23310 ,
         \23311 , \23312 , \23313 , \23314 , \23315 , \23316 , \23317 , \23318 , \23319 , \23320 ,
         \23321 , \23322 , \23323 , \23324 , \23325 , \23326 , \23327 , \23328 , \23329 , \23330 ,
         \23331 , \23332 , \23333 , \23334 , \23335 , \23336 , \23337 , \23338 , \23339 , \23340 ,
         \23341 , \23342 , \23343 , \23344 , \23345 , \23346 , \23347 , \23348 , \23349 , \23350 ,
         \23351 , \23352 , \23353 , \23354 , \23355 , \23356 , \23357 , \23358 , \23359 , \23360 ,
         \23361 , \23362 , \23363 , \23364 , \23365 , \23366 , \23367 , \23368 , \23369 , \23370 ,
         \23371 , \23372 , \23373 , \23374 , \23375 , \23376 , \23377 , \23378 , \23379 , \23380 ,
         \23381 , \23382 , \23383 , \23384 , \23385 , \23386 , \23387 , \23388 , \23389 , \23390 ,
         \23391 , \23392 , \23393 , \23394 , \23395 , \23396 , \23397 , \23398 , \23399 , \23400 ,
         \23401 , \23402 , \23403 , \23404 , \23405 , \23406 , \23407 , \23408 , \23409 , \23410 ,
         \23411 , \23412 , \23413 , \23414 , \23415 , \23416 , \23417 , \23418 , \23419 , \23420 ,
         \23421 , \23422 , \23423 , \23424 , \23425 , \23426 , \23427 , \23428 , \23429 , \23430 ,
         \23431 , \23432 , \23433 , \23434 , \23435 , \23436 , \23437 , \23438 , \23439 , \23440 ,
         \23441 , \23442 , \23443 , \23444 , \23445 , \23446 , \23447 , \23448 , \23449 , \23450 ,
         \23451 , \23452 , \23453 , \23454 , \23455 , \23456 , \23457 , \23458 , \23459 , \23460 ,
         \23461 , \23462 , \23463 , \23464 , \23465 , \23466 , \23467 , \23468 , \23469 , \23470 ,
         \23471 , \23472 , \23473 , \23474 , \23475 , \23476 , \23477 , \23478 , \23479 , \23480 ,
         \23481 , \23482 , \23483 , \23484 , \23485 , \23486 , \23487 , \23488 , \23489 , \23490 ,
         \23491 , \23492 , \23493 , \23494 , \23495 , \23496 , \23497 , \23498 , \23499 , \23500 ,
         \23501 , \23502 , \23503 , \23504 , \23505 , \23506 , \23507 , \23508 , \23509 , \23510 ,
         \23511 , \23512 , \23513 , \23514 , \23515 , \23516 , \23517 , \23518 , \23519 , \23520 ,
         \23521 , \23522 , \23523 , \23524 , \23525 , \23526 , \23527 , \23528 , \23529 , \23530 ,
         \23531 , \23532 , \23533 , \23534 , \23535 , \23536 , \23537 , \23538 , \23539 , \23540 ,
         \23541 , \23542 , \23543 , \23544 , \23545 , \23546 , \23547 , \23548 , \23549 , \23550 ,
         \23551 , \23552 , \23553 , \23554 , \23555 , \23556 , \23557 , \23558 , \23559 , \23560 ,
         \23561 , \23562 , \23563 , \23564 , \23565 , \23566 , \23567 , \23568 , \23569 , \23570 ,
         \23571 , \23572 , \23573 , \23574 , \23575 , \23576 , \23577 , \23578 , \23579 , \23580 ,
         \23581 , \23582 , \23583 , \23584 , \23585 , \23586 , \23587 , \23588 , \23589 , \23590 ,
         \23591 , \23592 , \23593 , \23594 , \23595 , \23596 , \23597 , \23598 , \23599 , \23600 ,
         \23601 , \23602 , \23603 , \23604 , \23605 , \23606 , \23607 , \23608 , \23609 , \23610 ,
         \23611 , \23612 , \23613 , \23614 , \23615 , \23616 , \23617 , \23618 , \23619 , \23620 ,
         \23621 , \23622 , \23623 , \23624 , \23625 , \23626 , \23627 , \23628 , \23629 , \23630 ,
         \23631 , \23632 , \23633 , \23634 , \23635 , \23636 , \23637 , \23638 , \23639 , \23640 ,
         \23641 , \23642 , \23643 , \23644 , \23645 , \23646 , \23647 , \23648 , \23649 , \23650 ,
         \23651 , \23652 , \23653 , \23654 , \23655 , \23656 , \23657 , \23658 , \23659 , \23660 ,
         \23661 , \23662 , \23663 , \23664 , \23665 , \23666 , \23667 , \23668 , \23669 , \23670 ,
         \23671 , \23672 , \23673 , \23674 , \23675 , \23676 , \23677 , \23678 , \23679 , \23680 ,
         \23681 , \23682 , \23683 , \23684 , \23685 , \23686 , \23687 , \23688 , \23689 , \23690 ,
         \23691 , \23692 , \23693 , \23694 , \23695 , \23696 , \23697 , \23698 , \23699 , \23700 ,
         \23701 , \23702 , \23703 , \23704 , \23705 , \23706 , \23707 , \23708 , \23709 , \23710 ,
         \23711 , \23712 , \23713 , \23714 , \23715 , \23716 , \23717 , \23718 , \23719 , \23720 ,
         \23721 , \23722 , \23723 , \23724 , \23725 , \23726 , \23727 , \23728 , \23729 , \23730 ,
         \23731 , \23732 , \23733 , \23734 , \23735 , \23736 , \23737 , \23738 , \23739 , \23740 ,
         \23741 , \23742 , \23743 , \23744 , \23745 , \23746 , \23747 , \23748 , \23749 , \23750 ,
         \23751 , \23752 , \23753 , \23754 , \23755 , \23756 , \23757 , \23758 , \23759 , \23760 ,
         \23761 , \23762 , \23763 , \23764 , \23765 , \23766 , \23767 , \23768 , \23769 , \23770 ,
         \23771 , \23772 , \23773 , \23774 , \23775 , \23776 , \23777 , \23778 , \23779 , \23780 ,
         \23781 , \23782 , \23783 , \23784 , \23785 , \23786 , \23787 , \23788 , \23789 , \23790 ,
         \23791 , \23792 , \23793 , \23794 , \23795 , \23796 , \23797 , \23798 , \23799 , \23800 ,
         \23801 , \23802 , \23803 , \23804 , \23805 , \23806 , \23807 , \23808 , \23809 , \23810 ,
         \23811 , \23812 , \23813 , \23814 , \23815 , \23816 , \23817 , \23818 , \23819 , \23820 ,
         \23821 , \23822 , \23823 , \23824 , \23825 , \23826 , \23827 , \23828 , \23829 , \23830 ,
         \23831 , \23832 , \23833 , \23834 , \23835 , \23836 , \23837 , \23838 , \23839 , \23840 ,
         \23841 , \23842 , \23843 , \23844 , \23845 , \23846 , \23847 , \23848 , \23849 , \23850 ,
         \23851 , \23852 , \23853 , \23854 , \23855 , \23856 , \23857 , \23858 , \23859 , \23860 ,
         \23861 , \23862 , \23863 , \23864 , \23865 , \23866 , \23867 , \23868 , \23869 , \23870 ,
         \23871 , \23872 , \23873 , \23874 , \23875 , \23876 , \23877 , \23878 , \23879 , \23880 ,
         \23881 , \23882 , \23883 , \23884 , \23885 , \23886 , \23887 , \23888 , \23889 , \23890 ,
         \23891 , \23892 , \23893 , \23894 , \23895 , \23896 , \23897 , \23898 , \23899 , \23900 ,
         \23901 , \23902 , \23903 , \23904 , \23905 , \23906 , \23907 , \23908 , \23909 , \23910 ,
         \23911 , \23912 , \23913 , \23914 , \23915 , \23916 , \23917 , \23918 , \23919 , \23920 ,
         \23921 , \23922 , \23923 , \23924 , \23925 , \23926 , \23927 , \23928 , \23929 , \23930 ,
         \23931 , \23932 , \23933 , \23934 , \23935 , \23936 , \23937 , \23938 , \23939 , \23940 ,
         \23941 , \23942 , \23943 , \23944 , \23945 , \23946 , \23947 , \23948 , \23949 , \23950 ,
         \23951 , \23952 , \23953 , \23954 , \23955 , \23956 , \23957 , \23958 , \23959 , \23960 ,
         \23961 , \23962 , \23963 , \23964 , \23965 , \23966 , \23967 , \23968 , \23969 , \23970 ,
         \23971 , \23972 , \23973 , \23974 , \23975 , \23976 , \23977 , \23978 , \23979 , \23980 ,
         \23981 , \23982 , \23983 , \23984 , \23985 , \23986 , \23987 , \23988 , \23989 , \23990 ,
         \23991 , \23992 , \23993 , \23994 , \23995 , \23996 , \23997 , \23998 , \23999 , \24000 ,
         \24001 , \24002 , \24003 , \24004 , \24005 , \24006 , \24007 , \24008 , \24009 , \24010 ,
         \24011 , \24012 , \24013 , \24014 , \24015 , \24016 , \24017 , \24018 , \24019 , \24020 ,
         \24021 , \24022 , \24023 , \24024 , \24025 , \24026 , \24027 , \24028 , \24029 , \24030 ,
         \24031 , \24032 , \24033 , \24034 , \24035 , \24036 , \24037 , \24038 , \24039 , \24040 ,
         \24041 , \24042 , \24043 , \24044 , \24045 , \24046 , \24047 , \24048 , \24049 , \24050 ,
         \24051 , \24052 , \24053 , \24054 , \24055 , \24056 , \24057 , \24058 , \24059 , \24060 ,
         \24061 , \24062 , \24063 , \24064 , \24065 , \24066 , \24067 , \24068 , \24069 , \24070 ,
         \24071 , \24072 , \24073 , \24074 , \24075 , \24076 , \24077 , \24078 , \24079 , \24080 ,
         \24081 , \24082 , \24083 , \24084 , \24085 , \24086 , \24087 , \24088 , \24089 , \24090 ,
         \24091 , \24092 , \24093 , \24094 , \24095 , \24096 , \24097 , \24098 , \24099 , \24100 ,
         \24101 , \24102 , \24103 , \24104 , \24105 , \24106 , \24107 , \24108 , \24109 , \24110 ,
         \24111 , \24112 , \24113 , \24114 , \24115 , \24116 , \24117 , \24118 , \24119 , \24120 ,
         \24121 , \24122 , \24123 , \24124 , \24125 , \24126 , \24127 , \24128 , \24129 , \24130 ,
         \24131 , \24132 , \24133 , \24134 , \24135 , \24136 , \24137 , \24138 , \24139 , \24140 ,
         \24141 , \24142 , \24143 , \24144 , \24145 , \24146 , \24147 , \24148 , \24149 , \24150 ,
         \24151 , \24152 , \24153 , \24154 , \24155 , \24156 , \24157 , \24158 , \24159 , \24160 ,
         \24161 , \24162 , \24163 , \24164 , \24165 , \24166 , \24167 , \24168 , \24169 , \24170 ,
         \24171 , \24172 , \24173 , \24174 , \24175 , \24176 , \24177 , \24178 , \24179 , \24180 ,
         \24181 , \24182 , \24183 , \24184 , \24185 , \24186 , \24187 , \24188 , \24189 , \24190 ,
         \24191 , \24192 , \24193 , \24194 , \24195 , \24196 , \24197 , \24198 , \24199 , \24200 ,
         \24201 , \24202 , \24203 , \24204 , \24205 , \24206 , \24207 , \24208 , \24209 , \24210 ,
         \24211 , \24212 , \24213 , \24214 , \24215 , \24216 , \24217 , \24218 , \24219 , \24220 ,
         \24221 , \24222 , \24223 , \24224 , \24225 , \24226 , \24227 , \24228 , \24229 , \24230 ,
         \24231 , \24232 , \24233 , \24234 , \24235 , \24236 , \24237 , \24238 , \24239 , \24240 ,
         \24241 , \24242 , \24243 , \24244 , \24245 , \24246 , \24247 , \24248 , \24249 , \24250 ,
         \24251 , \24252 , \24253 , \24254 , \24255 , \24256 , \24257 , \24258 , \24259 , \24260 ,
         \24261 , \24262 , \24263 , \24264 , \24265 , \24266 , \24267 , \24268 , \24269 , \24270 ,
         \24271 , \24272 , \24273 , \24274 , \24275 , \24276 , \24277 , \24278 , \24279 , \24280 ,
         \24281 , \24282 , \24283 , \24284 , \24285 , \24286 , \24287 , \24288 , \24289 , \24290 ,
         \24291 , \24292 , \24293 , \24294 , \24295 , \24296 , \24297 , \24298 , \24299 , \24300 ,
         \24301 , \24302 , \24303 , \24304 , \24305 , \24306 , \24307 , \24308 , \24309 , \24310 ,
         \24311 , \24312 , \24313 , \24314 , \24315 , \24316 , \24317 , \24318 , \24319 , \24320 ,
         \24321 , \24322 , \24323 , \24324 , \24325 , \24326 , \24327 , \24328 , \24329 , \24330 ,
         \24331 , \24332 , \24333 , \24334 , \24335 , \24336 , \24337 , \24338 , \24339 , \24340 ,
         \24341 , \24342 , \24343 , \24344 , \24345 , \24346 , \24347 , \24348 , \24349 , \24350 ,
         \24351 , \24352 , \24353 , \24354 , \24355 , \24356 , \24357 , \24358 , \24359 , \24360 ,
         \24361 , \24362 , \24363 , \24364 , \24365 , \24366 , \24367 , \24368 , \24369 , \24370 ,
         \24371 , \24372 , \24373 , \24374 , \24375 , \24376 , \24377 , \24378 , \24379 , \24380 ,
         \24381 , \24382 , \24383 , \24384 , \24385 , \24386 , \24387 , \24388 , \24389 , \24390 ,
         \24391 , \24392 , \24393 , \24394 , \24395 , \24396 , \24397 , \24398 , \24399 , \24400 ,
         \24401 , \24402 , \24403 , \24404 , \24405 , \24406 , \24407 , \24408 , \24409 , \24410 ,
         \24411 , \24412 , \24413 , \24414 , \24415 , \24416 , \24417 , \24418 , \24419 , \24420 ,
         \24421 , \24422 , \24423 , \24424 , \24425 , \24426 , \24427 , \24428 , \24429 , \24430 ,
         \24431 , \24432 , \24433 , \24434 , \24435 , \24436 , \24437 , \24438 , \24439 , \24440 ,
         \24441 , \24442 , \24443 , \24444 , \24445 , \24446 , \24447 , \24448 , \24449 , \24450 ,
         \24451 , \24452 , \24453 , \24454 , \24455 , \24456 , \24457 , \24458 , \24459 , \24460 ,
         \24461 , \24462 , \24463 , \24464 , \24465 , \24466 , \24467 , \24468 , \24469 , \24470 ,
         \24471 , \24472 , \24473 , \24474 , \24475 , \24476 , \24477 , \24478 , \24479 , \24480 ,
         \24481 , \24482 , \24483 , \24484 , \24485 , \24486 , \24487 , \24488 , \24489 , \24490 ,
         \24491 , \24492 , \24493 , \24494 , \24495 , \24496 , \24497 , \24498 , \24499 , \24500 ,
         \24501 , \24502 , \24503 , \24504 , \24505 , \24506 , \24507 , \24508 , \24509 , \24510 ,
         \24511 , \24512 , \24513 , \24514 , \24515 , \24516 , \24517 , \24518 , \24519 , \24520 ,
         \24521 , \24522 , \24523 , \24524 , \24525 , \24526 , \24527 , \24528 , \24529 , \24530 ,
         \24531 , \24532 , \24533 , \24534 , \24535 , \24536 , \24537 , \24538 , \24539 , \24540 ,
         \24541 , \24542 , \24543 , \24544 , \24545 , \24546 , \24547 , \24548 , \24549 , \24550 ,
         \24551 , \24552 , \24553 , \24554 , \24555 , \24556 , \24557 , \24558 , \24559 , \24560 ,
         \24561 , \24562 , \24563 , \24564 , \24565 , \24566 , \24567 , \24568 , \24569 , \24570 ,
         \24571 , \24572 , \24573 , \24574 , \24575 , \24576 , \24577 , \24578 , \24579 , \24580 ,
         \24581 , \24582 , \24583 , \24584 , \24585 , \24586 , \24587 , \24588 , \24589 , \24590 ,
         \24591 , \24592 , \24593 , \24594 , \24595 , \24596 , \24597 , \24598 , \24599 , \24600 ,
         \24601 , \24602 , \24603 , \24604 , \24605 , \24606 , \24607 , \24608 , \24609 , \24610 ,
         \24611 , \24612 , \24613 , \24614 , \24615 , \24616 , \24617 , \24618 , \24619 , \24620 ,
         \24621 , \24622 , \24623 , \24624 , \24625 , \24626 , \24627 , \24628 , \24629 , \24630 ,
         \24631 , \24632 , \24633 , \24634 , \24635 , \24636 , \24637 , \24638 , \24639 , \24640 ,
         \24641 , \24642 , \24643 , \24644 , \24645 , \24646 , \24647 , \24648 , \24649 , \24650 ,
         \24651 , \24652 , \24653 , \24654 , \24655 , \24656 , \24657 , \24658 , \24659 , \24660 ,
         \24661 , \24662 , \24663 , \24664 , \24665 , \24666 , \24667 , \24668 , \24669 , \24670 ,
         \24671 , \24672 , \24673 , \24674 , \24675 , \24676 , \24677 , \24678 , \24679 , \24680 ,
         \24681 , \24682 , \24683 , \24684 , \24685 , \24686 , \24687 , \24688 , \24689 , \24690 ,
         \24691 , \24692 , \24693 , \24694 , \24695 , \24696 , \24697 , \24698 , \24699 , \24700 ,
         \24701 , \24702 , \24703 , \24704 , \24705 , \24706 , \24707 , \24708 , \24709 , \24710 ,
         \24711 , \24712 , \24713 , \24714 , \24715 , \24716 , \24717 , \24718 , \24719 , \24720 ,
         \24721 , \24722 , \24723 , \24724 , \24725 , \24726 , \24727 , \24728 , \24729 , \24730 ,
         \24731 , \24732 , \24733 , \24734 , \24735 , \24736 , \24737 , \24738 , \24739 , \24740 ,
         \24741 , \24742 , \24743 , \24744 , \24745 , \24746 , \24747 , \24748 , \24749 , \24750 ,
         \24751 , \24752 , \24753 , \24754 , \24755 , \24756 , \24757 , \24758 , \24759 , \24760 ,
         \24761 , \24762 , \24763 , \24764 , \24765 , \24766 , \24767 , \24768 , \24769 , \24770 ,
         \24771 , \24772 , \24773 , \24774 , \24775 , \24776 , \24777 , \24778 , \24779 , \24780 ,
         \24781 , \24782 , \24783 , \24784 , \24785 , \24786 , \24787 , \24788 , \24789 , \24790 ,
         \24791 , \24792 , \24793 , \24794 , \24795 , \24796 , \24797 , \24798 , \24799 , \24800 ,
         \24801 , \24802 , \24803 , \24804 , \24805 , \24806 , \24807 , \24808 , \24809 , \24810 ,
         \24811 , \24812 , \24813 , \24814 , \24815 , \24816 , \24817 , \24818 , \24819 , \24820 ,
         \24821 , \24822 , \24823 , \24824 , \24825 , \24826 , \24827 , \24828 , \24829 , \24830 ,
         \24831 , \24832 , \24833 , \24834 , \24835 , \24836 , \24837 , \24838 , \24839 , \24840 ,
         \24841 , \24842 , \24843 , \24844 , \24845 , \24846 , \24847 , \24848 , \24849 , \24850 ,
         \24851 , \24852 , \24853 , \24854 , \24855 , \24856 , \24857 , \24858 , \24859 , \24860 ,
         \24861 , \24862 , \24863 , \24864 , \24865 , \24866 , \24867 , \24868 , \24869 , \24870 ,
         \24871 , \24872 , \24873 , \24874 , \24875 , \24876 , \24877 , \24878 , \24879 , \24880 ,
         \24881 , \24882 , \24883 , \24884 , \24885 , \24886 , \24887 , \24888 , \24889 , \24890 ,
         \24891 , \24892 , \24893 , \24894 , \24895 , \24896 , \24897 , \24898 , \24899 , \24900 ,
         \24901 , \24902 , \24903 , \24904 , \24905 , \24906 , \24907 , \24908 , \24909 , \24910 ,
         \24911 , \24912 , \24913 , \24914 , \24915 , \24916 , \24917 , \24918 , \24919 , \24920 ,
         \24921 , \24922 , \24923 , \24924 , \24925 , \24926 , \24927 , \24928 , \24929 , \24930 ,
         \24931 , \24932 , \24933 , \24934 , \24935 , \24936 , \24937 , \24938 , \24939 , \24940 ,
         \24941 , \24942 , \24943 , \24944 , \24945 , \24946 , \24947 , \24948 , \24949 , \24950 ,
         \24951 , \24952 , \24953 , \24954 , \24955 , \24956 , \24957 , \24958 , \24959 , \24960 ,
         \24961 , \24962 , \24963 , \24964 , \24965 , \24966 , \24967 , \24968 , \24969 , \24970 ,
         \24971 , \24972 , \24973 , \24974 , \24975 , \24976 , \24977 , \24978 , \24979 , \24980 ,
         \24981 , \24982 , \24983 , \24984 , \24985 , \24986 , \24987 , \24988 , \24989 , \24990 ,
         \24991 , \24992 , \24993 , \24994 , \24995 , \24996 , \24997 , \24998 , \24999 , \25000 ,
         \25001 , \25002 , \25003 , \25004 , \25005 , \25006 , \25007 , \25008 , \25009 , \25010 ,
         \25011 , \25012 , \25013 , \25014 , \25015 , \25016 , \25017 , \25018 , \25019 , \25020 ,
         \25021 , \25022 , \25023 , \25024 , \25025 , \25026 , \25027 , \25028 , \25029 , \25030 ,
         \25031 , \25032 , \25033 , \25034 , \25035 , \25036 , \25037 , \25038 , \25039 , \25040 ,
         \25041 , \25042 , \25043 , \25044 , \25045 , \25046 , \25047 , \25048 , \25049 , \25050 ,
         \25051 , \25052 , \25053 , \25054 , \25055 , \25056 , \25057 , \25058 , \25059 , \25060 ,
         \25061 , \25062 , \25063 , \25064 , \25065 , \25066 , \25067 , \25068 , \25069 , \25070 ,
         \25071 , \25072 , \25073 , \25074 , \25075 , \25076 , \25077 , \25078 , \25079 , \25080 ,
         \25081 , \25082 , \25083 , \25084 , \25085 , \25086 , \25087 , \25088 , \25089 , \25090 ,
         \25091 , \25092 , \25093 , \25094 , \25095 , \25096 , \25097 , \25098 , \25099 , \25100 ,
         \25101 , \25102 , \25103 , \25104 , \25105 , \25106 , \25107 , \25108 , \25109 , \25110 ,
         \25111 , \25112 , \25113 , \25114 , \25115 , \25116 , \25117 , \25118 , \25119 , \25120 ,
         \25121 , \25122 , \25123 , \25124 , \25125 , \25126 , \25127 , \25128 , \25129 , \25130 ,
         \25131 , \25132 , \25133 , \25134 , \25135 , \25136 , \25137 , \25138 , \25139 , \25140 ,
         \25141 , \25142 , \25143 , \25144 , \25145 , \25146 , \25147 , \25148 , \25149 , \25150 ,
         \25151 , \25152 , \25153 , \25154 , \25155 , \25156 , \25157 , \25158 , \25159 , \25160 ,
         \25161 , \25162 , \25163 , \25164 , \25165 , \25166 , \25167 , \25168 , \25169 , \25170 ,
         \25171 , \25172 , \25173 , \25174 , \25175 , \25176 , \25177 , \25178 , \25179 , \25180 ,
         \25181 , \25182 , \25183 , \25184 , \25185 , \25186 , \25187 , \25188 , \25189 , \25190 ,
         \25191 , \25192 , \25193 , \25194 , \25195 , \25196 , \25197 , \25198 , \25199 , \25200 ,
         \25201 , \25202 , \25203 , \25204 , \25205 , \25206 , \25207 , \25208 , \25209 , \25210 ,
         \25211 , \25212 , \25213 , \25214 , \25215 , \25216 , \25217 , \25218 , \25219 , \25220 ,
         \25221 , \25222 , \25223 , \25224 , \25225 , \25226 , \25227 , \25228 , \25229 , \25230 ,
         \25231 , \25232 , \25233 , \25234 , \25235 , \25236 , \25237 , \25238 , \25239 , \25240 ,
         \25241 , \25242 , \25243 , \25244 , \25245 , \25246 , \25247 , \25248 , \25249 , \25250 ,
         \25251 , \25252 , \25253 , \25254 , \25255 , \25256 , \25257 , \25258 , \25259 , \25260 ,
         \25261 , \25262 , \25263 , \25264 , \25265 , \25266 , \25267 , \25268 , \25269 , \25270 ,
         \25271 , \25272 , \25273 , \25274 , \25275 , \25276 , \25277 , \25278 , \25279 , \25280 ,
         \25281 , \25282 , \25283 , \25284 , \25285 , \25286 , \25287 , \25288 , \25289 , \25290 ,
         \25291 , \25292 , \25293 , \25294 , \25295 , \25296 , \25297 , \25298 , \25299 , \25300 ,
         \25301 , \25302 , \25303 , \25304 , \25305 , \25306 , \25307 , \25308 , \25309 , \25310 ,
         \25311 , \25312 , \25313 , \25314 , \25315 , \25316 , \25317 , \25318 , \25319 , \25320 ,
         \25321 , \25322 , \25323 , \25324 , \25325 , \25326 , \25327 , \25328 , \25329 , \25330 ,
         \25331 , \25332 , \25333 , \25334 , \25335 , \25336 , \25337 , \25338 , \25339 , \25340 ,
         \25341 , \25342 , \25343 , \25344 , \25345 , \25346 , \25347 , \25348 , \25349 , \25350 ,
         \25351 , \25352 , \25353 , \25354 , \25355 , \25356 , \25357 , \25358 , \25359 , \25360 ,
         \25361 , \25362 , \25363 , \25364 , \25365 , \25366 , \25367 , \25368 , \25369 , \25370 ,
         \25371 , \25372 , \25373 , \25374 , \25375 , \25376 , \25377 , \25378 , \25379 , \25380 ,
         \25381 , \25382 , \25383 , \25384 , \25385 , \25386 , \25387 , \25388 , \25389 , \25390 ,
         \25391 , \25392 , \25393 , \25394 , \25395 , \25396 , \25397 , \25398 , \25399 , \25400 ,
         \25401 , \25402 , \25403 , \25404 , \25405 , \25406 , \25407 , \25408 , \25409 , \25410 ,
         \25411 , \25412 , \25413 , \25414 , \25415 , \25416 , \25417 , \25418 , \25419 , \25420 ,
         \25421 , \25422 , \25423 , \25424 , \25425 , \25426 , \25427 , \25428 , \25429 , \25430 ,
         \25431 , \25432 , \25433 , \25434 , \25435 , \25436 , \25437 , \25438 , \25439 , \25440 ,
         \25441 , \25442 , \25443 , \25444 , \25445 , \25446 , \25447 , \25448 , \25449 , \25450 ,
         \25451 , \25452 , \25453 , \25454 , \25455 , \25456 , \25457 , \25458 , \25459 , \25460 ,
         \25461 , \25462 , \25463 , \25464 , \25465 , \25466 , \25467 , \25468 , \25469 , \25470 ,
         \25471 , \25472 , \25473 , \25474 , \25475 , \25476 , \25477 , \25478 , \25479 , \25480 ,
         \25481 , \25482 , \25483 , \25484 , \25485 , \25486 , \25487 , \25488 , \25489 , \25490 ,
         \25491 , \25492 , \25493 , \25494 , \25495 , \25496 , \25497 , \25498 , \25499 , \25500 ,
         \25501 , \25502 , \25503 , \25504 , \25505 , \25506 , \25507 , \25508 , \25509 , \25510 ,
         \25511 , \25512 , \25513 , \25514 , \25515 , \25516 , \25517 , \25518 , \25519 , \25520 ,
         \25521 , \25522 , \25523 , \25524 , \25525 , \25526 , \25527 , \25528 , \25529 , \25530 ,
         \25531 , \25532 , \25533 , \25534 , \25535 , \25536 , \25537 , \25538 , \25539 , \25540 ,
         \25541 , \25542 , \25543 , \25544 , \25545 , \25546 , \25547 , \25548 , \25549 , \25550 ,
         \25551 , \25552 , \25553 , \25554 , \25555 , \25556 , \25557 , \25558 , \25559 , \25560 ,
         \25561 , \25562 , \25563 , \25564 , \25565 , \25566 , \25567 , \25568 , \25569 , \25570 ,
         \25571 , \25572 , \25573 , \25574 , \25575 , \25576 , \25577 , \25578 , \25579 , \25580 ,
         \25581 , \25582 , \25583 , \25584 , \25585 , \25586 , \25587 , \25588 , \25589 , \25590 ,
         \25591 , \25592 , \25593 , \25594 , \25595 , \25596 , \25597 , \25598 , \25599 , \25600 ,
         \25601 , \25602 , \25603 , \25604 , \25605 , \25606 , \25607 , \25608 , \25609 , \25610 ,
         \25611 , \25612 , \25613 , \25614 , \25615 , \25616 , \25617 , \25618 , \25619 , \25620 ,
         \25621 , \25622 , \25623 , \25624 , \25625 , \25626 , \25627 , \25628 , \25629 , \25630 ,
         \25631 , \25632 , \25633 , \25634 , \25635 , \25636 , \25637 , \25638 , \25639 , \25640 ,
         \25641 , \25642 , \25643 , \25644 , \25645 , \25646 , \25647 , \25648 , \25649 , \25650 ,
         \25651 , \25652 , \25653 , \25654 , \25655 , \25656 , \25657 , \25658 , \25659 , \25660 ,
         \25661 , \25662 , \25663 , \25664 , \25665 , \25666 , \25667 , \25668 , \25669 , \25670 ,
         \25671 , \25672 , \25673 , \25674 , \25675 , \25676 , \25677 , \25678 , \25679 , \25680 ,
         \25681 , \25682 , \25683 , \25684 , \25685 , \25686 , \25687 , \25688 , \25689 , \25690 ,
         \25691 , \25692 , \25693 , \25694 , \25695 , \25696 , \25697 , \25698 , \25699 , \25700 ,
         \25701 , \25702 , \25703 , \25704 , \25705 , \25706 , \25707 , \25708 , \25709 , \25710 ,
         \25711 , \25712 , \25713 , \25714 , \25715 , \25716 , \25717 , \25718 , \25719 , \25720 ,
         \25721 , \25722 , \25723 , \25724 , \25725 , \25726 , \25727 , \25728 , \25729 , \25730 ,
         \25731 , \25732 , \25733 , \25734 , \25735 , \25736 , \25737 , \25738 , \25739 , \25740 ,
         \25741 , \25742 , \25743 , \25744 , \25745 , \25746 , \25747 , \25748 , \25749 , \25750 ,
         \25751 , \25752 , \25753 , \25754 , \25755 , \25756 , \25757 , \25758 , \25759 , \25760 ,
         \25761 , \25762 , \25763 , \25764 , \25765 , \25766 , \25767 , \25768 , \25769 , \25770 ,
         \25771 , \25772 , \25773 , \25774 , \25775 , \25776 , \25777 , \25778 , \25779 , \25780 ,
         \25781 , \25782 , \25783 , \25784 , \25785 , \25786 , \25787 , \25788 , \25789 , \25790 ,
         \25791 , \25792 , \25793 , \25794 , \25795 , \25796 , \25797 , \25798 , \25799 , \25800 ,
         \25801 , \25802 , \25803 , \25804 , \25805 , \25806 , \25807 , \25808 , \25809 , \25810 ,
         \25811 , \25812 , \25813 , \25814 , \25815 , \25816 , \25817 , \25818 , \25819 , \25820 ,
         \25821 , \25822 , \25823 , \25824 , \25825 , \25826 , \25827 , \25828 , \25829 , \25830 ,
         \25831 , \25832 , \25833 , \25834 , \25835 , \25836 , \25837 , \25838 , \25839 , \25840 ,
         \25841 , \25842 , \25843 , \25844 , \25845 , \25846 , \25847 , \25848 , \25849 , \25850 ,
         \25851 , \25852 , \25853 , \25854 , \25855 , \25856 , \25857 , \25858 , \25859 , \25860 ,
         \25861 , \25862 , \25863 , \25864 , \25865 , \25866 , \25867 , \25868 , \25869 , \25870 ,
         \25871 , \25872 , \25873 , \25874 , \25875 , \25876 , \25877 , \25878 , \25879 , \25880 ,
         \25881 , \25882 , \25883 , \25884 , \25885 , \25886 , \25887 , \25888 , \25889 , \25890 ,
         \25891 , \25892 , \25893 , \25894 , \25895 , \25896 , \25897 , \25898 , \25899 , \25900 ,
         \25901 , \25902 , \25903 , \25904 , \25905 , \25906 , \25907 , \25908 , \25909 , \25910 ,
         \25911 , \25912 , \25913 , \25914 , \25915 , \25916 , \25917 , \25918 , \25919 , \25920 ,
         \25921 , \25922 , \25923 , \25924 , \25925 , \25926 , \25927 , \25928 , \25929 , \25930 ,
         \25931 , \25932 , \25933 , \25934 , \25935 , \25936 , \25937 , \25938 , \25939 , \25940 ,
         \25941 , \25942 , \25943 , \25944 , \25945 , \25946 , \25947 , \25948 , \25949 , \25950 ,
         \25951 , \25952 , \25953 , \25954 , \25955 , \25956 , \25957 , \25958 , \25959 , \25960 ,
         \25961 , \25962 , \25963 , \25964 , \25965 , \25966 , \25967 , \25968 , \25969 , \25970 ,
         \25971 , \25972 , \25973 , \25974 , \25975 , \25976 , \25977 , \25978 , \25979 , \25980 ,
         \25981 , \25982 , \25983 , \25984 , \25985 , \25986 , \25987 , \25988 , \25989 , \25990 ,
         \25991 , \25992 , \25993 , \25994 , \25995 , \25996 , \25997 , \25998 , \25999 , \26000 ,
         \26001 , \26002 , \26003 , \26004 , \26005 , \26006 , \26007 , \26008 , \26009 , \26010 ,
         \26011 , \26012 , \26013 , \26014 , \26015 , \26016 , \26017 , \26018 , \26019 , \26020 ,
         \26021 , \26022 , \26023 , \26024 , \26025 , \26026 , \26027 , \26028 , \26029 , \26030 ,
         \26031 , \26032 , \26033 , \26034 , \26035 , \26036 , \26037 , \26038 , \26039 , \26040 ,
         \26041 , \26042 , \26043 , \26044 , \26045 , \26046 , \26047 , \26048 , \26049 , \26050 ,
         \26051 , \26052 , \26053 , \26054 , \26055 , \26056 , \26057 , \26058 , \26059 , \26060 ,
         \26061 , \26062 , \26063 , \26064 , \26065 , \26066 , \26067 , \26068 , \26069 , \26070 ,
         \26071 , \26072 , \26073 , \26074 , \26075 , \26076 , \26077 , \26078 , \26079 , \26080 ,
         \26081 , \26082 , \26083 , \26084 , \26085 , \26086 , \26087 , \26088 , \26089 , \26090 ,
         \26091 , \26092 , \26093 , \26094 , \26095 , \26096 , \26097 , \26098 , \26099 , \26100 ,
         \26101 , \26102 , \26103 , \26104 , \26105 , \26106 , \26107 , \26108 , \26109 , \26110 ,
         \26111 , \26112 , \26113 , \26114 , \26115 , \26116 , \26117 , \26118 , \26119 , \26120 ,
         \26121 , \26122 , \26123 , \26124 , \26125 , \26126 , \26127 , \26128 , \26129 , \26130 ,
         \26131 , \26132 , \26133 , \26134 , \26135 , \26136 , \26137 , \26138 , \26139 , \26140 ,
         \26141 , \26142 , \26143 , \26144 , \26145 , \26146 , \26147 , \26148 , \26149 , \26150 ,
         \26151 , \26152 , \26153 , \26154 , \26155 , \26156 , \26157 , \26158 , \26159 , \26160 ,
         \26161 , \26162 , \26163 , \26164 , \26165 , \26166 , \26167 , \26168 , \26169 , \26170 ,
         \26171 , \26172 , \26173 , \26174 , \26175 , \26176 , \26177 , \26178 , \26179 , \26180 ,
         \26181 , \26182 , \26183 , \26184 , \26185 , \26186 , \26187 , \26188 , \26189 , \26190 ,
         \26191 , \26192 , \26193 , \26194 , \26195 , \26196 , \26197 , \26198 , \26199 , \26200 ,
         \26201 , \26202 , \26203 , \26204 , \26205 , \26206 , \26207 , \26208 , \26209 , \26210 ,
         \26211 , \26212 , \26213 , \26214 , \26215 , \26216 , \26217 , \26218 , \26219 , \26220 ,
         \26221 , \26222 , \26223 , \26224 , \26225 , \26226 , \26227 , \26228 , \26229 , \26230 ,
         \26231 , \26232 , \26233 , \26234 , \26235 , \26236 , \26237 , \26238 , \26239 , \26240 ,
         \26241 , \26242 , \26243 , \26244 , \26245 , \26246 , \26247 , \26248 , \26249 , \26250 ,
         \26251 , \26252 , \26253 , \26254 , \26255 , \26256 , \26257 , \26258 , \26259 , \26260 ,
         \26261 , \26262 , \26263 , \26264 , \26265 , \26266 , \26267 , \26268 , \26269 , \26270 ,
         \26271 , \26272 , \26273 , \26274 , \26275 , \26276 , \26277 , \26278 , \26279 , \26280 ,
         \26281 , \26282 , \26283 , \26284 , \26285 , \26286 , \26287 , \26288 , \26289 , \26290 ,
         \26291 , \26292 , \26293 , \26294 , \26295 , \26296 , \26297 , \26298 , \26299 , \26300 ,
         \26301 , \26302 , \26303 , \26304 , \26305 , \26306 , \26307 , \26308 , \26309 , \26310 ,
         \26311 , \26312 , \26313 , \26314 , \26315 , \26316 , \26317 , \26318 , \26319 , \26320 ,
         \26321 , \26322 , \26323 , \26324 , \26325 , \26326 , \26327 , \26328 , \26329 , \26330 ,
         \26331 , \26332 , \26333 , \26334 , \26335 , \26336 , \26337 , \26338 , \26339 , \26340 ,
         \26341 , \26342 , \26343 , \26344 , \26345 , \26346 , \26347 , \26348 , \26349 , \26350 ,
         \26351 , \26352 , \26353 , \26354 , \26355 , \26356 , \26357 , \26358 , \26359 , \26360 ,
         \26361 , \26362 , \26363 , \26364 , \26365 , \26366 , \26367 , \26368 , \26369 , \26370 ,
         \26371 , \26372 , \26373 , \26374 , \26375 , \26376 , \26377 , \26378 , \26379 , \26380 ,
         \26381 , \26382 , \26383 , \26384 , \26385 , \26386 , \26387 , \26388 , \26389 , \26390 ,
         \26391 , \26392 , \26393 , \26394 , \26395 , \26396 , \26397 , \26398 , \26399 , \26400 ,
         \26401 , \26402 , \26403 , \26404 , \26405 , \26406 , \26407 , \26408 , \26409 , \26410 ,
         \26411 , \26412 , \26413 , \26414 , \26415 , \26416 , \26417 , \26418 , \26419 , \26420 ,
         \26421 , \26422 , \26423 , \26424 , \26425 , \26426 , \26427 , \26428 , \26429 , \26430 ,
         \26431 , \26432 , \26433 , \26434 , \26435 , \26436 , \26437 , \26438 , \26439 , \26440 ,
         \26441 , \26442 , \26443 , \26444 , \26445 , \26446 , \26447 , \26448 , \26449 , \26450 ,
         \26451 , \26452 , \26453 , \26454 , \26455 , \26456 , \26457 , \26458 , \26459 , \26460 ,
         \26461 , \26462 , \26463 , \26464 , \26465 , \26466 , \26467 , \26468 , \26469 , \26470 ,
         \26471 , \26472 , \26473 , \26474 , \26475 , \26476 , \26477 , \26478 , \26479 , \26480 ,
         \26481 , \26482 , \26483 , \26484 , \26485 , \26486 , \26487 , \26488 , \26489 , \26490 ,
         \26491 , \26492 , \26493 , \26494 , \26495 , \26496 , \26497 , \26498 , \26499 , \26500 ,
         \26501 , \26502 , \26503 , \26504 , \26505 , \26506 , \26507 , \26508 , \26509 , \26510 ,
         \26511 , \26512 , \26513 , \26514 , \26515 , \26516 , \26517 , \26518 , \26519 , \26520 ,
         \26521 , \26522 , \26523 , \26524 , \26525 , \26526 , \26527 , \26528 , \26529 , \26530 ,
         \26531 , \26532 , \26533 , \26534 , \26535 , \26536 , \26537 , \26538 , \26539 , \26540 ,
         \26541 , \26542 , \26543 , \26544 , \26545 , \26546 , \26547 , \26548 , \26549 , \26550 ,
         \26551 , \26552 , \26553 , \26554 , \26555 , \26556 , \26557 , \26558 , \26559 , \26560 ,
         \26561 , \26562 , \26563 , \26564 , \26565 , \26566 , \26567 , \26568 , \26569 , \26570 ,
         \26571 , \26572 , \26573 , \26574 , \26575 , \26576 , \26577 , \26578 , \26579 , \26580 ,
         \26581 , \26582 , \26583 , \26584 , \26585 , \26586 , \26587 , \26588 , \26589 , \26590 ,
         \26591 , \26592 , \26593 , \26594 , \26595 , \26596 , \26597 , \26598 , \26599 , \26600 ,
         \26601 , \26602 , \26603 , \26604 , \26605 , \26606 , \26607 , \26608 , \26609 , \26610 ,
         \26611 , \26612 , \26613 , \26614 , \26615 , \26616 , \26617 , \26618 , \26619 , \26620 ,
         \26621 , \26622 , \26623 , \26624 , \26625 , \26626 , \26627 , \26628 , \26629 , \26630 ,
         \26631 , \26632 , \26633 , \26634 , \26635 , \26636 , \26637 , \26638 , \26639 , \26640 ,
         \26641 , \26642 , \26643 , \26644 , \26645 , \26646 , \26647 , \26648 , \26649 , \26650 ,
         \26651 , \26652 , \26653 , \26654 , \26655 , \26656 , \26657 , \26658 , \26659 , \26660 ,
         \26661 , \26662 , \26663 , \26664 , \26665 , \26666 , \26667 , \26668 , \26669 , \26670 ,
         \26671 , \26672 , \26673 , \26674 , \26675 , \26676 , \26677 , \26678 , \26679 , \26680 ,
         \26681 , \26682 , \26683 , \26684 , \26685 , \26686 , \26687 , \26688 , \26689 , \26690 ,
         \26691 , \26692 , \26693 , \26694 , \26695 , \26696 , \26697 , \26698 , \26699 , \26700 ,
         \26701 , \26702 , \26703 , \26704 , \26705 , \26706 , \26707 , \26708 , \26709 , \26710 ,
         \26711 , \26712 , \26713 , \26714 , \26715 , \26716 , \26717 , \26718 , \26719 , \26720 ,
         \26721 , \26722 , \26723 , \26724 , \26725 , \26726 , \26727 , \26728 , \26729 , \26730 ,
         \26731 , \26732 , \26733 , \26734 , \26735 , \26736 , \26737 , \26738 , \26739 , \26740 ,
         \26741 , \26742 , \26743 , \26744 , \26745 , \26746 , \26747 , \26748 , \26749 , \26750 ,
         \26751 , \26752 , \26753 , \26754 , \26755 , \26756 , \26757 , \26758 , \26759 , \26760 ,
         \26761 , \26762 , \26763 , \26764 , \26765 , \26766 , \26767 , \26768 , \26769 , \26770 ,
         \26771 , \26772 , \26773 , \26774 , \26775 , \26776 , \26777 , \26778 , \26779 , \26780 ,
         \26781 , \26782 , \26783 , \26784 , \26785 , \26786 , \26787 , \26788 , \26789 , \26790 ,
         \26791 , \26792 , \26793 , \26794 , \26795 , \26796 , \26797 , \26798 , \26799 , \26800 ,
         \26801 , \26802 , \26803 , \26804 , \26805 , \26806 , \26807 , \26808 , \26809 , \26810 ,
         \26811 , \26812 , \26813 , \26814 , \26815 , \26816 , \26817 , \26818 , \26819 , \26820 ,
         \26821 , \26822 , \26823 , \26824 , \26825 , \26826 , \26827 , \26828 , \26829 , \26830 ,
         \26831 , \26832 , \26833 , \26834 , \26835 , \26836 , \26837 , \26838 , \26839 , \26840 ,
         \26841 , \26842 , \26843 , \26844 , \26845 , \26846 , \26847 , \26848 , \26849 , \26850 ,
         \26851 , \26852 , \26853 , \26854 , \26855 , \26856 , \26857 , \26858 , \26859 , \26860 ,
         \26861 , \26862 , \26863 , \26864 , \26865 , \26866 , \26867 , \26868 , \26869 , \26870 ,
         \26871 , \26872 , \26873 , \26874 , \26875 , \26876 , \26877 , \26878 , \26879 , \26880 ,
         \26881 , \26882 , \26883 , \26884 , \26885 , \26886 , \26887 , \26888 , \26889 , \26890 ,
         \26891 , \26892 , \26893 , \26894 , \26895 , \26896 , \26897 , \26898 , \26899 , \26900 ,
         \26901 , \26902 , \26903 , \26904 , \26905 , \26906 , \26907 , \26908 , \26909 , \26910 ,
         \26911 , \26912 , \26913 , \26914 , \26915 , \26916 , \26917 , \26918 , \26919 , \26920 ,
         \26921 , \26922 , \26923 , \26924 , \26925 , \26926 , \26927 , \26928 , \26929 , \26930 ,
         \26931 , \26932 , \26933 , \26934 , \26935 , \26936 , \26937 , \26938 , \26939 , \26940 ,
         \26941 , \26942 , \26943 , \26944 , \26945 , \26946 , \26947 , \26948 , \26949 , \26950 ,
         \26951 , \26952 , \26953 , \26954 , \26955 , \26956 , \26957 , \26958 , \26959 , \26960 ,
         \26961 , \26962 , \26963 , \26964 , \26965 , \26966 , \26967 , \26968 , \26969 , \26970 ,
         \26971 , \26972 , \26973 , \26974 , \26975 , \26976 , \26977 , \26978 , \26979 , \26980 ,
         \26981 , \26982 , \26983 , \26984 , \26985 , \26986 , \26987 , \26988 , \26989 , \26990 ,
         \26991 , \26992 , \26993 , \26994 , \26995 , \26996 , \26997 , \26998 , \26999 , \27000 ,
         \27001 , \27002 , \27003 , \27004 , \27005 , \27006 , \27007 , \27008 , \27009 , \27010 ,
         \27011 , \27012 , \27013 , \27014 , \27015 , \27016 , \27017 , \27018 , \27019 , \27020 ,
         \27021 , \27022 , \27023 , \27024 , \27025 , \27026 , \27027 , \27028 , \27029 , \27030 ,
         \27031 , \27032 , \27033 , \27034 , \27035 , \27036 , \27037 , \27038 , \27039 , \27040 ,
         \27041 , \27042 , \27043 , \27044 , \27045 , \27046 , \27047 , \27048 , \27049 , \27050 ,
         \27051 , \27052 , \27053 , \27054 , \27055 , \27056 , \27057 , \27058 , \27059 , \27060 ,
         \27061 , \27062 , \27063 , \27064 , \27065 , \27066 , \27067 , \27068 , \27069 , \27070 ,
         \27071 , \27072 , \27073 , \27074 , \27075 , \27076 , \27077 , \27078 , \27079 , \27080 ,
         \27081 , \27082 , \27083 , \27084 , \27085 , \27086 , \27087 , \27088 , \27089 , \27090 ,
         \27091 , \27092 , \27093 , \27094 , \27095 , \27096 , \27097 , \27098 , \27099 , \27100 ,
         \27101 , \27102 , \27103 , \27104 , \27105 , \27106 , \27107 , \27108 , \27109 , \27110 ,
         \27111 , \27112 , \27113 , \27114 , \27115 , \27116 , \27117 , \27118 , \27119 , \27120 ,
         \27121 , \27122 , \27123 , \27124 , \27125 , \27126 , \27127 , \27128 , \27129 , \27130 ,
         \27131 , \27132 , \27133 , \27134 , \27135 , \27136 , \27137 , \27138 , \27139 , \27140 ,
         \27141 , \27142 , \27143 , \27144 , \27145 , \27146 , \27147 , \27148 , \27149 , \27150 ,
         \27151 , \27152 , \27153 , \27154 , \27155 , \27156 , \27157 , \27158 , \27159 , \27160 ,
         \27161 , \27162 , \27163 , \27164 , \27165 , \27166 , \27167 , \27168 , \27169 , \27170 ,
         \27171 , \27172 , \27173 , \27174 , \27175 , \27176 , \27177 , \27178 , \27179 , \27180 ,
         \27181 , \27182 , \27183 , \27184 , \27185 , \27186 , \27187 , \27188 , \27189 , \27190 ,
         \27191 , \27192 , \27193 , \27194 , \27195 , \27196 , \27197 , \27198 , \27199 , \27200 ,
         \27201 , \27202 , \27203 , \27204 , \27205 , \27206 , \27207 , \27208 , \27209 , \27210 ,
         \27211 , \27212 , \27213 , \27214 , \27215 , \27216 , \27217 , \27218 , \27219 , \27220 ,
         \27221 , \27222 , \27223 , \27224 , \27225 , \27226 , \27227 , \27228 , \27229 , \27230 ,
         \27231 , \27232 , \27233 , \27234 , \27235 , \27236 , \27237 , \27238 , \27239 , \27240 ,
         \27241 , \27242 , \27243 , \27244 , \27245 , \27246 , \27247 , \27248 , \27249 , \27250 ,
         \27251 , \27252 , \27253 , \27254 , \27255 , \27256 , \27257 , \27258 , \27259 , \27260 ,
         \27261 , \27262 , \27263 , \27264 , \27265 , \27266 , \27267 , \27268 , \27269 , \27270 ,
         \27271 , \27272 , \27273 , \27274 , \27275 , \27276 , \27277 , \27278 , \27279 , \27280 ,
         \27281 , \27282 , \27283 , \27284 , \27285 , \27286 , \27287 , \27288 , \27289 , \27290 ,
         \27291 , \27292 , \27293 , \27294 , \27295 , \27296 , \27297 , \27298 , \27299 , \27300 ,
         \27301 , \27302 , \27303 , \27304 , \27305 , \27306 , \27307 , \27308 , \27309 , \27310 ,
         \27311 , \27312 , \27313 , \27314 , \27315 , \27316 , \27317 , \27318 , \27319 , \27320 ,
         \27321 , \27322 , \27323 , \27324 , \27325 , \27326 , \27327 , \27328 , \27329 , \27330 ,
         \27331 , \27332 , \27333 , \27334 , \27335 , \27336 , \27337 , \27338 , \27339 , \27340 ,
         \27341 , \27342 , \27343 , \27344 , \27345 , \27346 , \27347 , \27348 , \27349 , \27350 ,
         \27351 , \27352 , \27353 , \27354 , \27355 , \27356 , \27357 , \27358 , \27359 , \27360 ,
         \27361 , \27362 , \27363 , \27364 , \27365 , \27366 , \27367 , \27368 , \27369 , \27370 ,
         \27371 , \27372 , \27373 , \27374 , \27375 , \27376 , \27377 , \27378 , \27379 , \27380 ,
         \27381 , \27382 , \27383 , \27384 , \27385 , \27386 , \27387 , \27388 , \27389 , \27390 ,
         \27391 , \27392 , \27393 , \27394 , \27395 , \27396 , \27397 , \27398 , \27399 , \27400 ,
         \27401 , \27402 , \27403 , \27404 , \27405 , \27406 , \27407 , \27408 , \27409 , \27410 ,
         \27411 , \27412 , \27413 , \27414 , \27415 , \27416 , \27417 , \27418 , \27419 , \27420 ,
         \27421 , \27422 , \27423 , \27424 , \27425 , \27426 , \27427 , \27428 , \27429 , \27430 ,
         \27431 , \27432 , \27433 , \27434 , \27435 , \27436 , \27437 , \27438 , \27439 , \27440 ,
         \27441 , \27442 , \27443 , \27444 , \27445 , \27446 , \27447 , \27448 , \27449 , \27450 ,
         \27451 , \27452 , \27453 , \27454 , \27455 , \27456 , \27457 , \27458 , \27459 , \27460 ,
         \27461 , \27462 , \27463 , \27464 , \27465 , \27466 , \27467 , \27468 , \27469 , \27470 ,
         \27471 , \27472 , \27473 , \27474 , \27475 , \27476 , \27477 , \27478 , \27479 , \27480 ,
         \27481 , \27482 , \27483 , \27484 , \27485 , \27486 , \27487 , \27488 , \27489 , \27490 ,
         \27491 , \27492 , \27493 , \27494 , \27495 , \27496 , \27497 , \27498 , \27499 , \27500 ,
         \27501 , \27502 , \27503 , \27504 , \27505 , \27506 , \27507 , \27508 , \27509 , \27510 ,
         \27511 , \27512 , \27513 , \27514 , \27515 , \27516 , \27517 , \27518 , \27519 , \27520 ,
         \27521 , \27522 , \27523 , \27524 , \27525 , \27526 , \27527 , \27528 , \27529 , \27530 ,
         \27531 , \27532 , \27533 , \27534 , \27535 , \27536 , \27537 , \27538 , \27539 , \27540 ,
         \27541 , \27542 , \27543 , \27544 , \27545 , \27546 , \27547 , \27548 , \27549 , \27550 ,
         \27551 , \27552 , \27553 , \27554 , \27555 , \27556 , \27557 , \27558 , \27559 , \27560 ,
         \27561 , \27562 , \27563 , \27564 , \27565 , \27566 , \27567 , \27568 , \27569 , \27570 ,
         \27571 , \27572 , \27573 , \27574 , \27575 , \27576 , \27577 , \27578 , \27579 , \27580 ,
         \27581 , \27582 , \27583 , \27584 , \27585 , \27586 , \27587 , \27588 , \27589 , \27590 ,
         \27591 , \27592 , \27593 , \27594 , \27595 , \27596 , \27597 , \27598 , \27599 , \27600 ,
         \27601 , \27602 , \27603 , \27604 , \27605 , \27606 , \27607 , \27608 , \27609 , \27610 ,
         \27611 , \27612 , \27613 , \27614 , \27615 , \27616 , \27617 , \27618 , \27619 , \27620 ,
         \27621 , \27622 , \27623 , \27624 , \27625 , \27626 , \27627 , \27628 , \27629 , \27630 ,
         \27631 , \27632 , \27633 , \27634 , \27635 , \27636 , \27637 , \27638 , \27639 , \27640 ,
         \27641 , \27642 , \27643 , \27644 , \27645 , \27646 , \27647 , \27648 , \27649 , \27650 ,
         \27651 , \27652 , \27653 , \27654 , \27655 , \27656 , \27657 , \27658 , \27659 , \27660 ,
         \27661 , \27662 , \27663 , \27664 , \27665 , \27666 , \27667 , \27668 , \27669 , \27670 ,
         \27671 , \27672 , \27673 , \27674 , \27675 , \27676 , \27677 , \27678 , \27679 , \27680 ,
         \27681 , \27682 , \27683 , \27684 , \27685 , \27686 , \27687 , \27688 , \27689 , \27690 ,
         \27691 , \27692 , \27693 , \27694 , \27695 , \27696 , \27697 , \27698 , \27699 , \27700 ,
         \27701 , \27702 , \27703 , \27704 , \27705 , \27706 , \27707 , \27708 , \27709 , \27710 ,
         \27711 , \27712 , \27713 , \27714 , \27715 , \27716 , \27717 , \27718 , \27719 , \27720 ,
         \27721 , \27722 , \27723 , \27724 , \27725 , \27726 , \27727 , \27728 , \27729 , \27730 ,
         \27731 , \27732 , \27733 , \27734 , \27735 , \27736 , \27737 , \27738 , \27739 , \27740 ,
         \27741 , \27742 , \27743 , \27744 , \27745 , \27746 , \27747 , \27748 , \27749 , \27750 ,
         \27751 , \27752 , \27753 , \27754 , \27755 , \27756 , \27757 , \27758 , \27759 , \27760 ,
         \27761 , \27762 , \27763 , \27764 , \27765 , \27766 , \27767 , \27768 , \27769 , \27770 ,
         \27771 , \27772 , \27773 , \27774 , \27775 , \27776 , \27777 , \27778 , \27779 , \27780 ,
         \27781 , \27782 , \27783 , \27784 , \27785 , \27786 , \27787 , \27788 , \27789 , \27790 ,
         \27791 , \27792 , \27793 , \27794 , \27795 , \27796 , \27797 , \27798 , \27799 , \27800 ,
         \27801 , \27802 , \27803 , \27804 , \27805 , \27806 , \27807 , \27808 , \27809 , \27810 ,
         \27811 , \27812 , \27813 , \27814 , \27815 , \27816 , \27817 , \27818 , \27819 , \27820 ,
         \27821 , \27822 , \27823 , \27824 , \27825 , \27826 , \27827 , \27828 , \27829 , \27830 ,
         \27831 , \27832 , \27833 , \27834 , \27835 , \27836 , \27837 , \27838 , \27839 , \27840 ,
         \27841 , \27842 , \27843 , \27844 , \27845 , \27846 , \27847 , \27848 , \27849 , \27850 ,
         \27851 , \27852 , \27853 , \27854 , \27855 , \27856 , \27857 , \27858 , \27859 , \27860 ,
         \27861 , \27862 , \27863 , \27864 , \27865 , \27866 , \27867 , \27868 , \27869 , \27870 ,
         \27871 , \27872 , \27873 , \27874 , \27875 , \27876 , \27877 , \27878 , \27879 , \27880 ,
         \27881 , \27882 , \27883 , \27884 , \27885 , \27886 , \27887 , \27888 , \27889 , \27890 ,
         \27891 , \27892 , \27893 , \27894 , \27895 , \27896 , \27897 , \27898 , \27899 , \27900 ,
         \27901 , \27902 , \27903 , \27904 , \27905 , \27906 , \27907 , \27908 , \27909 , \27910 ,
         \27911 , \27912 , \27913 , \27914 , \27915 , \27916 , \27917 , \27918 , \27919 , \27920 ,
         \27921 , \27922 , \27923 , \27924 , \27925 , \27926 , \27927 , \27928 , \27929 , \27930 ,
         \27931 , \27932 , \27933 , \27934 , \27935 , \27936 , \27937 , \27938 , \27939 , \27940 ,
         \27941 , \27942 , \27943 , \27944 , \27945 , \27946 , \27947 , \27948 , \27949 , \27950 ,
         \27951 , \27952 , \27953 , \27954 , \27955 , \27956 , \27957 , \27958 , \27959 , \27960 ,
         \27961 , \27962 , \27963 , \27964 , \27965 , \27966 , \27967 , \27968 , \27969 , \27970 ,
         \27971 , \27972 , \27973 , \27974 , \27975 , \27976 , \27977 , \27978 , \27979 , \27980 ,
         \27981 , \27982 , \27983 , \27984 , \27985 , \27986 , \27987 , \27988 , \27989 , \27990 ,
         \27991 , \27992 , \27993 , \27994 , \27995 , \27996 , \27997 , \27998 , \27999 , \28000 ,
         \28001 , \28002 , \28003 , \28004 , \28005 , \28006 , \28007 , \28008 , \28009 , \28010 ,
         \28011 , \28012 , \28013 , \28014 , \28015 , \28016 , \28017 , \28018 , \28019 , \28020 ,
         \28021 , \28022 , \28023 , \28024 , \28025 , \28026 , \28027 , \28028 , \28029 , \28030 ,
         \28031 , \28032 , \28033 , \28034 , \28035 , \28036 , \28037 , \28038 , \28039 , \28040 ,
         \28041 , \28042 , \28043 , \28044 , \28045 , \28046 , \28047 , \28048 , \28049 , \28050 ,
         \28051 , \28052 , \28053 , \28054 , \28055 , \28056 , \28057 , \28058 , \28059 , \28060 ,
         \28061 , \28062 , \28063 , \28064 , \28065 , \28066 , \28067 , \28068 , \28069 , \28070 ,
         \28071 , \28072 , \28073 , \28074 , \28075 , \28076 , \28077 , \28078 , \28079 , \28080 ,
         \28081 , \28082 , \28083 , \28084 , \28085 , \28086 , \28087 , \28088 , \28089 , \28090 ,
         \28091 , \28092 , \28093 , \28094 , \28095 , \28096 , \28097 , \28098 , \28099 , \28100 ,
         \28101 , \28102 , \28103 , \28104 , \28105 , \28106 , \28107 , \28108 , \28109 , \28110 ,
         \28111 , \28112 , \28113 , \28114 , \28115 , \28116 , \28117 , \28118 , \28119 , \28120 ,
         \28121 , \28122 , \28123 , \28124 , \28125 , \28126 , \28127 , \28128 , \28129 , \28130 ,
         \28131 , \28132 , \28133 , \28134 , \28135 , \28136 , \28137 , \28138 , \28139 , \28140 ,
         \28141 , \28142 , \28143 , \28144 , \28145 , \28146 , \28147 , \28148 , \28149 , \28150 ,
         \28151 , \28152 , \28153 , \28154 , \28155 , \28156 , \28157 , \28158 , \28159 , \28160 ,
         \28161 , \28162 , \28163 , \28164 , \28165 , \28166 , \28167 , \28168 , \28169 , \28170 ,
         \28171 , \28172 , \28173 , \28174 , \28175 , \28176 , \28177 , \28178 , \28179 , \28180 ,
         \28181 , \28182 , \28183 , \28184 , \28185 , \28186 , \28187 , \28188 , \28189 , \28190 ,
         \28191 , \28192 , \28193 , \28194 , \28195 , \28196 , \28197 , \28198 , \28199 , \28200 ,
         \28201 , \28202 , \28203 , \28204 , \28205 , \28206 , \28207 , \28208 , \28209 , \28210 ,
         \28211 , \28212 , \28213 , \28214 , \28215 , \28216 , \28217 , \28218 , \28219 , \28220 ,
         \28221 , \28222 , \28223 , \28224 , \28225 , \28226 , \28227 , \28228 , \28229 , \28230 ,
         \28231 , \28232 , \28233 , \28234 , \28235 , \28236 , \28237 , \28238 , \28239 , \28240 ,
         \28241 , \28242 , \28243 , \28244 , \28245 , \28246 , \28247 , \28248 , \28249 , \28250 ,
         \28251 , \28252 , \28253 , \28254 , \28255 , \28256 , \28257 , \28258 , \28259 , \28260 ,
         \28261 , \28262 , \28263 , \28264 , \28265 , \28266 , \28267 , \28268 , \28269 , \28270 ,
         \28271 , \28272 , \28273 , \28274 , \28275 , \28276 , \28277 , \28278 , \28279 , \28280 ,
         \28281 , \28282 , \28283 , \28284 , \28285 , \28286 , \28287 , \28288 , \28289 , \28290 ,
         \28291 , \28292 , \28293 , \28294 , \28295 , \28296 , \28297 , \28298 , \28299 , \28300 ,
         \28301 , \28302 , \28303 , \28304 , \28305 , \28306 , \28307 , \28308 , \28309 , \28310 ,
         \28311 , \28312 , \28313 , \28314 , \28315 , \28316 , \28317 , \28318 , \28319 , \28320 ,
         \28321 , \28322 , \28323 , \28324 , \28325 , \28326 , \28327 , \28328 , \28329 , \28330 ,
         \28331 , \28332 , \28333 , \28334 , \28335 , \28336 , \28337 , \28338 , \28339 , \28340 ,
         \28341 , \28342 , \28343 , \28344 , \28345 , \28346 , \28347 , \28348 , \28349 , \28350 ,
         \28351 , \28352 , \28353 , \28354 , \28355 , \28356 , \28357 , \28358 , \28359 , \28360 ,
         \28361 , \28362 , \28363 , \28364 , \28365 , \28366 , \28367 , \28368 , \28369 , \28370 ,
         \28371 , \28372 , \28373 , \28374 , \28375 , \28376 , \28377 , \28378 , \28379 , \28380 ,
         \28381 , \28382 , \28383 , \28384 , \28385 , \28386 , \28387 , \28388 , \28389 , \28390 ,
         \28391 , \28392 , \28393 , \28394 , \28395 , \28396 , \28397 , \28398 , \28399 , \28400 ,
         \28401 , \28402 , \28403 , \28404 , \28405 , \28406 , \28407 , \28408 , \28409 , \28410 ,
         \28411 , \28412 , \28413 , \28414 , \28415 , \28416 , \28417 , \28418 , \28419 , \28420 ,
         \28421 , \28422 , \28423 , \28424 , \28425 , \28426 , \28427 , \28428 , \28429 , \28430 ,
         \28431 , \28432 , \28433 , \28434 , \28435 , \28436 , \28437 , \28438 , \28439 , \28440 ,
         \28441 , \28442 , \28443 , \28444 , \28445 , \28446 , \28447 , \28448 , \28449 , \28450 ,
         \28451 , \28452 , \28453 , \28454 , \28455 , \28456 , \28457 , \28458 , \28459 , \28460 ,
         \28461 , \28462 , \28463 , \28464 , \28465 , \28466 , \28467 , \28468 , \28469 , \28470 ,
         \28471 , \28472 , \28473 , \28474 , \28475 , \28476 , \28477 , \28478 , \28479 , \28480 ,
         \28481 , \28482 , \28483 , \28484 , \28485 , \28486 , \28487 , \28488 , \28489 , \28490 ,
         \28491 , \28492 , \28493 , \28494 , \28495 , \28496 , \28497 , \28498 , \28499 , \28500 ,
         \28501 , \28502 , \28503 , \28504 , \28505 , \28506 , \28507 , \28508 , \28509 , \28510 ,
         \28511 , \28512 , \28513 , \28514 , \28515 , \28516 , \28517 , \28518 , \28519 , \28520 ,
         \28521 , \28522 , \28523 , \28524 , \28525 , \28526 , \28527 , \28528 , \28529 , \28530 ,
         \28531 , \28532 , \28533 , \28534 , \28535 , \28536 , \28537 , \28538 , \28539 , \28540 ,
         \28541 , \28542 , \28543 , \28544 , \28545 , \28546 , \28547 , \28548 , \28549 , \28550 ,
         \28551 , \28552 , \28553 , \28554 , \28555 , \28556 , \28557 , \28558 , \28559 , \28560 ,
         \28561 , \28562 , \28563 , \28564 , \28565 , \28566 , \28567 , \28568 , \28569 , \28570 ,
         \28571 , \28572 , \28573 , \28574 , \28575 , \28576 , \28577 , \28578 , \28579 , \28580 ,
         \28581 , \28582 , \28583 , \28584 , \28585 , \28586 , \28587 , \28588 , \28589 , \28590 ,
         \28591 , \28592 , \28593 , \28594 , \28595 , \28596 , \28597 , \28598 , \28599 , \28600 ,
         \28601 , \28602 , \28603 , \28604 , \28605 , \28606 , \28607 , \28608 , \28609 , \28610 ,
         \28611 , \28612 , \28613 , \28614 , \28615 , \28616 , \28617 , \28618 , \28619 , \28620 ,
         \28621 , \28622 , \28623 , \28624 , \28625 , \28626 , \28627 , \28628 , \28629 , \28630 ,
         \28631 , \28632 , \28633 , \28634 , \28635 , \28636 , \28637 , \28638 , \28639 , \28640 ,
         \28641 , \28642 , \28643 , \28644 , \28645 , \28646 , \28647 , \28648 , \28649 , \28650 ,
         \28651 , \28652 , \28653 , \28654 , \28655 , \28656 , \28657 , \28658 , \28659 , \28660 ,
         \28661 , \28662 , \28663 , \28664 , \28665 , \28666 , \28667 , \28668 , \28669 , \28670 ,
         \28671 , \28672 , \28673 , \28674 , \28675 , \28676 , \28677 , \28678 , \28679 , \28680 ,
         \28681 , \28682 , \28683 , \28684 , \28685 , \28686 , \28687 , \28688 , \28689 , \28690 ,
         \28691 , \28692 , \28693 , \28694 , \28695 , \28696 , \28697 , \28698 , \28699 , \28700 ,
         \28701 , \28702 , \28703 , \28704 , \28705 , \28706 , \28707 , \28708 , \28709 , \28710 ,
         \28711 , \28712 , \28713 , \28714 , \28715 , \28716 , \28717 , \28718 , \28719 , \28720 ,
         \28721 , \28722 , \28723 , \28724 , \28725 , \28726 , \28727 , \28728 , \28729 , \28730 ,
         \28731 , \28732 , \28733 , \28734 , \28735 , \28736 , \28737 , \28738 , \28739 , \28740 ,
         \28741 , \28742 , \28743 , \28744 , \28745 , \28746 , \28747 , \28748 , \28749 , \28750 ,
         \28751 , \28752 , \28753 , \28754 , \28755 , \28756 , \28757 , \28758 , \28759 , \28760 ,
         \28761 , \28762 , \28763 , \28764 , \28765 , \28766 , \28767 , \28768 , \28769 , \28770 ,
         \28771 , \28772 , \28773 , \28774 , \28775 , \28776 , \28777 , \28778 , \28779 , \28780 ,
         \28781 , \28782 , \28783 , \28784 , \28785 , \28786 , \28787 , \28788 , \28789 , \28790 ,
         \28791 , \28792 , \28793 , \28794 , \28795 , \28796 , \28797 , \28798 , \28799 , \28800 ,
         \28801 , \28802 , \28803 , \28804 , \28805 , \28806 , \28807 , \28808 , \28809 , \28810 ,
         \28811 , \28812 , \28813 , \28814 , \28815 , \28816 , \28817 , \28818 , \28819 , \28820 ,
         \28821 , \28822 , \28823 , \28824 , \28825 , \28826 , \28827 , \28828 , \28829 , \28830 ,
         \28831 , \28832 , \28833 , \28834 , \28835 , \28836 , \28837 , \28838 , \28839 , \28840 ,
         \28841 , \28842 , \28843 , \28844 , \28845 , \28846 , \28847 , \28848 , \28849 , \28850 ,
         \28851 , \28852 , \28853 , \28854 , \28855 , \28856 , \28857 , \28858 , \28859 , \28860 ,
         \28861 , \28862 , \28863 , \28864 , \28865 , \28866 , \28867 , \28868 , \28869 , \28870 ,
         \28871 , \28872 , \28873 , \28874 , \28875 , \28876 , \28877 , \28878 , \28879 , \28880 ,
         \28881 , \28882 , \28883 , \28884 , \28885 , \28886 , \28887 , \28888 , \28889 , \28890 ,
         \28891 , \28892 , \28893 , \28894 , \28895 , \28896 , \28897 , \28898 , \28899 , \28900 ,
         \28901 , \28902 , \28903 , \28904 , \28905 , \28906 , \28907 , \28908 , \28909 , \28910 ,
         \28911 , \28912 , \28913 , \28914 , \28915 , \28916 , \28917 , \28918 , \28919 , \28920 ,
         \28921 , \28922 , \28923 , \28924 , \28925 , \28926 , \28927 , \28928 , \28929 , \28930 ,
         \28931 , \28932 , \28933 , \28934 , \28935 , \28936 , \28937 , \28938 , \28939 , \28940 ,
         \28941 , \28942 , \28943 , \28944 , \28945 , \28946 , \28947 , \28948 , \28949 , \28950 ,
         \28951 , \28952 , \28953 , \28954 , \28955 , \28956 , \28957 , \28958 , \28959 , \28960 ,
         \28961 , \28962 , \28963 , \28964 , \28965 , \28966 , \28967 , \28968 , \28969 , \28970 ,
         \28971 , \28972 , \28973 , \28974 , \28975 , \28976 , \28977 , \28978 , \28979 , \28980 ,
         \28981 , \28982 , \28983 , \28984 , \28985 , \28986 , \28987 , \28988 , \28989 , \28990 ,
         \28991 , \28992 , \28993 , \28994 , \28995 , \28996 , \28997 , \28998 , \28999 , \29000 ,
         \29001 , \29002 , \29003 , \29004 , \29005 , \29006 , \29007 , \29008 , \29009 , \29010 ,
         \29011 , \29012 , \29013 , \29014 , \29015 , \29016 , \29017 , \29018 , \29019 , \29020 ,
         \29021 , \29022 , \29023 , \29024 , \29025 , \29026 , \29027 , \29028 , \29029 , \29030 ,
         \29031 , \29032 , \29033 , \29034 , \29035 , \29036 , \29037 , \29038 , \29039 , \29040 ,
         \29041 , \29042 , \29043 , \29044 , \29045 , \29046 , \29047 , \29048 , \29049 , \29050 ,
         \29051 , \29052 , \29053 , \29054 , \29055 , \29056 , \29057 , \29058 , \29059 , \29060 ,
         \29061 , \29062 , \29063 , \29064 , \29065 , \29066 , \29067 , \29068 , \29069 , \29070 ,
         \29071 , \29072 , \29073 , \29074 , \29075 , \29076 , \29077 , \29078 , \29079 , \29080 ,
         \29081 , \29082 , \29083 , \29084 , \29085 , \29086 , \29087 , \29088 , \29089 , \29090 ,
         \29091 , \29092 , \29093 , \29094 , \29095 , \29096 , \29097 , \29098 , \29099 , \29100 ,
         \29101 , \29102 , \29103 , \29104 , \29105 , \29106 , \29107 , \29108 , \29109 , \29110 ,
         \29111 , \29112 , \29113 , \29114 , \29115 , \29116 , \29117 , \29118 , \29119 , \29120 ,
         \29121 , \29122 , \29123 , \29124 , \29125 , \29126 , \29127 , \29128 , \29129 , \29130 ,
         \29131 , \29132 , \29133 , \29134 , \29135 , \29136 , \29137 , \29138 , \29139 , \29140 ,
         \29141 , \29142 , \29143 , \29144 , \29145 , \29146 , \29147 , \29148 , \29149 , \29150 ,
         \29151 , \29152 , \29153 , \29154 , \29155 , \29156 , \29157 , \29158 , \29159 , \29160 ,
         \29161 , \29162 , \29163 , \29164 , \29165 , \29166 , \29167 , \29168 , \29169 , \29170 ,
         \29171 , \29172 , \29173 , \29174 , \29175 , \29176 , \29177 , \29178 , \29179 , \29180 ,
         \29181 , \29182 , \29183 , \29184 , \29185 , \29186 , \29187 , \29188 , \29189 , \29190 ,
         \29191 , \29192 , \29193 , \29194 , \29195 , \29196 , \29197 , \29198 , \29199 , \29200 ,
         \29201 , \29202 , \29203 , \29204 , \29205 , \29206 , \29207 , \29208 , \29209 , \29210 ,
         \29211 , \29212 , \29213 , \29214 , \29215 , \29216 , \29217 , \29218 , \29219 , \29220 ,
         \29221 , \29222 , \29223 , \29224 , \29225 , \29226 , \29227 , \29228 , \29229 , \29230 ,
         \29231 , \29232 , \29233 , \29234 , \29235 , \29236 , \29237 , \29238 , \29239 , \29240 ,
         \29241 , \29242 , \29243 , \29244 , \29245 , \29246 , \29247 , \29248 , \29249 , \29250 ,
         \29251 , \29252 , \29253 , \29254 , \29255 , \29256 , \29257 , \29258 , \29259 , \29260 ,
         \29261 , \29262 , \29263 , \29264 , \29265 , \29266 , \29267 , \29268 , \29269 , \29270 ,
         \29271 , \29272 , \29273 , \29274 , \29275 , \29276 , \29277 , \29278 , \29279 , \29280 ,
         \29281 , \29282 , \29283 , \29284 , \29285 , \29286 , \29287 , \29288 , \29289 , \29290 ,
         \29291 , \29292 , \29293 , \29294 , \29295 , \29296 , \29297 , \29298 , \29299 , \29300 ,
         \29301 , \29302 , \29303 , \29304 , \29305 , \29306 , \29307 , \29308 , \29309 , \29310 ,
         \29311 , \29312 , \29313 , \29314 , \29315 , \29316 , \29317 , \29318 , \29319 , \29320 ,
         \29321 , \29322 , \29323 , \29324 , \29325 , \29326 , \29327 , \29328 , \29329 , \29330 ,
         \29331 , \29332 , \29333 , \29334 , \29335 , \29336 , \29337 , \29338 , \29339 , \29340 ,
         \29341 , \29342 , \29343 , \29344 , \29345 , \29346 , \29347 , \29348 , \29349 , \29350 ,
         \29351 , \29352 , \29353 , \29354 , \29355 , \29356 , \29357 , \29358 , \29359 , \29360 ,
         \29361 , \29362 , \29363 , \29364 , \29365 , \29366 , \29367 , \29368 , \29369 , \29370 ,
         \29371 , \29372 , \29373 , \29374 , \29375 , \29376 , \29377 , \29378 , \29379 , \29380 ,
         \29381 , \29382 , \29383 , \29384 , \29385 , \29386 , \29387 , \29388 , \29389 , \29390 ,
         \29391 , \29392 , \29393 , \29394 , \29395 , \29396 , \29397 , \29398 , \29399 , \29400 ,
         \29401 , \29402 , \29403 , \29404 , \29405 , \29406 , \29407 , \29408 , \29409 , \29410 ,
         \29411 , \29412 , \29413 , \29414 , \29415 , \29416 , \29417 , \29418 , \29419 , \29420 ,
         \29421 , \29422 , \29423 , \29424 , \29425 , \29426 , \29427 , \29428 , \29429 , \29430 ,
         \29431 , \29432 , \29433 , \29434 , \29435 , \29436 , \29437 , \29438 , \29439 , \29440 ,
         \29441 , \29442 , \29443 , \29444 , \29445 , \29446 , \29447 , \29448 , \29449 , \29450 ,
         \29451 , \29452 , \29453 , \29454 , \29455 , \29456 , \29457 , \29458 , \29459 , \29460 ,
         \29461 , \29462 , \29463 , \29464 , \29465 , \29466 , \29467 , \29468 , \29469 , \29470 ,
         \29471 , \29472 , \29473 , \29474 , \29475 , \29476 , \29477 , \29478 , \29479 , \29480 ,
         \29481 , \29482 , \29483 , \29484 , \29485 , \29486 , \29487 , \29488 , \29489 , \29490 ,
         \29491 , \29492 , \29493 , \29494 , \29495 , \29496 , \29497 , \29498 , \29499 , \29500 ,
         \29501 , \29502 , \29503 , \29504 , \29505 , \29506 , \29507 , \29508 , \29509 , \29510 ,
         \29511 , \29512 , \29513 , \29514 , \29515 , \29516 , \29517 , \29518 , \29519 , \29520 ,
         \29521 , \29522 , \29523 , \29524 , \29525 , \29526 , \29527 , \29528 , \29529 , \29530 ,
         \29531 , \29532 , \29533 , \29534 , \29535 , \29536 , \29537 , \29538 , \29539 , \29540 ,
         \29541 , \29542 , \29543 , \29544 , \29545 , \29546 , \29547 , \29548 , \29549 , \29550 ,
         \29551 , \29552 , \29553 , \29554 , \29555 , \29556 , \29557 , \29558 , \29559 , \29560 ,
         \29561 , \29562 , \29563 , \29564 , \29565 , \29566 , \29567 , \29568 , \29569 , \29570 ,
         \29571 , \29572 , \29573 , \29574 , \29575 , \29576 , \29577 , \29578 , \29579 , \29580 ,
         \29581 , \29582 , \29583 , \29584 , \29585 , \29586 , \29587 , \29588 , \29589 , \29590 ,
         \29591 , \29592 , \29593 , \29594 , \29595 , \29596 , \29597 , \29598 , \29599 , \29600 ,
         \29601 , \29602 , \29603 , \29604 , \29605 , \29606 , \29607 , \29608 , \29609 , \29610 ,
         \29611 , \29612 , \29613 , \29614 , \29615 , \29616 , \29617 , \29618 , \29619 , \29620 ,
         \29621 , \29622 , \29623 , \29624 , \29625 , \29626 , \29627 , \29628 , \29629 , \29630 ,
         \29631 , \29632 , \29633 , \29634 , \29635 , \29636 , \29637 , \29638 , \29639 , \29640 ,
         \29641 , \29642 , \29643 , \29644 , \29645 , \29646 , \29647 , \29648 , \29649 , \29650 ,
         \29651 , \29652 , \29653 , \29654 , \29655 , \29656 , \29657 , \29658 , \29659 , \29660 ,
         \29661 , \29662 , \29663 , \29664 , \29665 , \29666 , \29667 , \29668 , \29669 , \29670 ,
         \29671 , \29672 , \29673 , \29674 , \29675 , \29676 , \29677 , \29678 , \29679 , \29680 ,
         \29681 , \29682 , \29683 , \29684 , \29685 , \29686 , \29687 , \29688 , \29689 , \29690 ,
         \29691 , \29692 , \29693 , \29694 , \29695 , \29696 , \29697 , \29698 , \29699 , \29700 ,
         \29701 , \29702 , \29703 , \29704 , \29705 , \29706 , \29707 , \29708 , \29709 , \29710 ,
         \29711 , \29712 , \29713 , \29714 , \29715 , \29716 , \29717 , \29718 , \29719 , \29720 ,
         \29721 , \29722 , \29723 , \29724 , \29725 , \29726 , \29727 , \29728 , \29729 , \29730 ,
         \29731 , \29732 , \29733 , \29734 , \29735 , \29736 , \29737 , \29738 , \29739 , \29740 ,
         \29741 , \29742 , \29743 , \29744 , \29745 , \29746 , \29747 , \29748 , \29749 , \29750 ,
         \29751 , \29752 , \29753 , \29754 , \29755 , \29756 , \29757 , \29758 , \29759 , \29760 ,
         \29761 , \29762 , \29763 , \29764 , \29765 , \29766 , \29767 , \29768 , \29769 , \29770 ,
         \29771 , \29772 , \29773 , \29774 , \29775 , \29776 , \29777 , \29778 , \29779 , \29780 ,
         \29781 , \29782 , \29783 , \29784 , \29785 , \29786 , \29787 , \29788 , \29789 , \29790 ,
         \29791 , \29792 , \29793 , \29794 , \29795 , \29796 , \29797 , \29798 , \29799 , \29800 ,
         \29801 , \29802 , \29803 , \29804 , \29805 , \29806 , \29807 , \29808 , \29809 , \29810 ,
         \29811 , \29812 , \29813 , \29814 , \29815 , \29816 , \29817 , \29818 , \29819 , \29820 ,
         \29821 , \29822 , \29823 , \29824 , \29825 , \29826 , \29827 , \29828 , \29829 , \29830 ,
         \29831 , \29832 , \29833 , \29834 , \29835 , \29836 , \29837 , \29838 , \29839 , \29840 ,
         \29841 , \29842 , \29843 , \29844 , \29845 , \29846 , \29847 , \29848 , \29849 , \29850 ,
         \29851 , \29852 , \29853 , \29854 , \29855 , \29856 , \29857 , \29858 , \29859 , \29860 ,
         \29861 , \29862 , \29863 , \29864 , \29865 , \29866 , \29867 , \29868 , \29869 , \29870 ,
         \29871 , \29872 , \29873 , \29874 , \29875 , \29876 , \29877 , \29878 , \29879 , \29880 ,
         \29881 , \29882 , \29883 , \29884 , \29885 , \29886 , \29887 , \29888 , \29889 , \29890 ,
         \29891 , \29892 , \29893 , \29894 , \29895 , \29896 , \29897 , \29898 , \29899 , \29900 ,
         \29901 , \29902 , \29903 , \29904 , \29905 , \29906 , \29907 , \29908 , \29909 , \29910 ,
         \29911 , \29912 , \29913 , \29914 , \29915 , \29916 , \29917 , \29918 , \29919 , \29920 ,
         \29921 , \29922 , \29923 , \29924 , \29925 , \29926 , \29927 , \29928 , \29929 , \29930 ,
         \29931 , \29932 , \29933 , \29934 , \29935 , \29936 , \29937 , \29938 , \29939 , \29940 ,
         \29941 , \29942 , \29943 , \29944 , \29945 , \29946 , \29947 , \29948 , \29949 , \29950 ,
         \29951 , \29952 , \29953 , \29954 , \29955 , \29956 , \29957 , \29958 , \29959 , \29960 ,
         \29961 , \29962 , \29963 , \29964 , \29965 , \29966 , \29967 , \29968 , \29969 , \29970 ,
         \29971 , \29972 , \29973 , \29974 , \29975 , \29976 , \29977 , \29978 , \29979 , \29980 ,
         \29981 , \29982 , \29983 , \29984 , \29985 , \29986 , \29987 , \29988 , \29989 , \29990 ,
         \29991 , \29992 , \29993 , \29994 , \29995 , \29996 , \29997 , \29998 , \29999 , \30000 ,
         \30001 , \30002 , \30003 , \30004 , \30005 , \30006 , \30007 , \30008 , \30009 , \30010 ,
         \30011 , \30012 , \30013 , \30014 , \30015 , \30016 , \30017 , \30018 , \30019 , \30020 ,
         \30021 , \30022 , \30023 , \30024 , \30025 , \30026 , \30027 , \30028 , \30029 , \30030 ,
         \30031 , \30032 , \30033 , \30034 , \30035 , \30036 , \30037 , \30038 , \30039 , \30040 ,
         \30041 , \30042 , \30043 , \30044 , \30045 , \30046 , \30047 , \30048 , \30049 , \30050 ,
         \30051 , \30052 , \30053 , \30054 , \30055 , \30056 , \30057 , \30058 , \30059 , \30060 ,
         \30061 , \30062 , \30063 , \30064 , \30065 , \30066 , \30067 , \30068 , \30069 , \30070 ,
         \30071 , \30072 , \30073 , \30074 , \30075 , \30076 , \30077 , \30078 , \30079 , \30080 ,
         \30081 , \30082 , \30083 , \30084 , \30085 , \30086 , \30087 , \30088 , \30089 , \30090 ,
         \30091 , \30092 , \30093 , \30094 , \30095 , \30096 , \30097 , \30098 , \30099 , \30100 ,
         \30101 , \30102 , \30103 , \30104 , \30105 , \30106 , \30107 , \30108 , \30109 , \30110 ,
         \30111 , \30112 , \30113 , \30114 , \30115 , \30116 , \30117 , \30118 , \30119 , \30120 ,
         \30121 , \30122 , \30123 , \30124 , \30125 , \30126 , \30127 , \30128 , \30129 , \30130 ,
         \30131 , \30132 , \30133 , \30134 , \30135 , \30136 , \30137 , \30138 , \30139 , \30140 ,
         \30141 , \30142 , \30143 , \30144 , \30145 , \30146 , \30147 , \30148 , \30149 , \30150 ,
         \30151 , \30152 , \30153 , \30154 , \30155 , \30156 , \30157 , \30158 , \30159 , \30160 ,
         \30161 , \30162 , \30163 , \30164 , \30165 , \30166 , \30167 , \30168 , \30169 , \30170 ,
         \30171 , \30172 , \30173 , \30174 , \30175 , \30176 , \30177 , \30178 , \30179 , \30180 ,
         \30181 , \30182 , \30183 , \30184 , \30185 , \30186 , \30187 , \30188 , \30189 , \30190 ,
         \30191 , \30192 , \30193 , \30194 , \30195 , \30196 , \30197 , \30198 , \30199 , \30200 ,
         \30201 , \30202 , \30203 , \30204 , \30205 , \30206 , \30207 , \30208 , \30209 , \30210 ,
         \30211 , \30212 , \30213 , \30214 , \30215 , \30216 , \30217 , \30218 , \30219 , \30220 ,
         \30221 , \30222 , \30223 , \30224 , \30225 , \30226 , \30227 , \30228 , \30229 , \30230 ,
         \30231 , \30232 , \30233 , \30234 , \30235 , \30236 , \30237 , \30238 , \30239 , \30240 ,
         \30241 , \30242 , \30243 , \30244 , \30245 , \30246 , \30247 , \30248 , \30249 , \30250 ,
         \30251 , \30252 , \30253 , \30254 , \30255 , \30256 , \30257 , \30258 , \30259 , \30260 ,
         \30261 , \30262 , \30263 , \30264 , \30265 , \30266 , \30267 , \30268 , \30269 , \30270 ,
         \30271 , \30272 , \30273 , \30274 , \30275 , \30276 , \30277 , \30278 , \30279 , \30280 ,
         \30281 , \30282 , \30283 , \30284 , \30285 , \30286 , \30287 , \30288 , \30289 , \30290 ,
         \30291 , \30292 , \30293 , \30294 , \30295 , \30296 , \30297 , \30298 , \30299 , \30300 ,
         \30301 , \30302 , \30303 , \30304 , \30305 , \30306 , \30307 , \30308 , \30309 , \30310 ,
         \30311 , \30312 , \30313 , \30314 , \30315 , \30316 , \30317 , \30318 , \30319 , \30320 ,
         \30321 , \30322 , \30323 , \30324 , \30325 , \30326 , \30327 , \30328 , \30329 , \30330 ,
         \30331 , \30332 , \30333 , \30334 , \30335 , \30336 , \30337 , \30338 , \30339 , \30340 ,
         \30341 , \30342 , \30343 , \30344 , \30345 , \30346 , \30347 , \30348 , \30349 , \30350 ,
         \30351 , \30352 , \30353 , \30354 , \30355 , \30356 , \30357 , \30358 , \30359 , \30360 ,
         \30361 , \30362 , \30363 , \30364 , \30365 , \30366 , \30367 , \30368 , \30369 , \30370 ,
         \30371 , \30372 , \30373 , \30374 , \30375 , \30376 , \30377 , \30378 , \30379 , \30380 ,
         \30381 , \30382 , \30383 , \30384 , \30385 , \30386 , \30387 , \30388 , \30389 , \30390 ,
         \30391 , \30392 , \30393 , \30394 , \30395 , \30396 , \30397 , \30398 , \30399 , \30400 ,
         \30401 , \30402 , \30403 , \30404 , \30405 , \30406 , \30407 , \30408 , \30409 , \30410 ,
         \30411 , \30412 , \30413 , \30414 , \30415 , \30416 , \30417 , \30418 , \30419 , \30420 ,
         \30421 , \30422 , \30423 , \30424 , \30425 , \30426 , \30427 , \30428 , \30429 , \30430 ,
         \30431 , \30432 , \30433 , \30434 , \30435 , \30436 , \30437 , \30438 , \30439 , \30440 ,
         \30441 , \30442 , \30443 , \30444 , \30445 , \30446 , \30447 , \30448 , \30449 , \30450 ,
         \30451 , \30452 , \30453 , \30454 , \30455 , \30456 , \30457 , \30458 , \30459 , \30460 ,
         \30461 , \30462 , \30463 , \30464 , \30465 , \30466 , \30467 , \30468 , \30469 , \30470 ,
         \30471 , \30472 , \30473 , \30474 , \30475 , \30476 , \30477 , \30478 , \30479 , \30480 ,
         \30481 , \30482 , \30483 , \30484 , \30485 , \30486 , \30487 , \30488 , \30489 , \30490 ,
         \30491 , \30492 , \30493 , \30494 , \30495 , \30496 , \30497 , \30498 , \30499 , \30500 ,
         \30501 , \30502 , \30503 , \30504 , \30505 , \30506 , \30507 , \30508 , \30509 , \30510 ,
         \30511 , \30512 , \30513 , \30514 , \30515 , \30516 , \30517 , \30518 , \30519 , \30520 ,
         \30521 , \30522 , \30523 , \30524 , \30525 , \30526 , \30527 , \30528 , \30529 , \30530 ,
         \30531 , \30532 , \30533 , \30534 , \30535 , \30536 , \30537 , \30538 , \30539 , \30540 ,
         \30541 , \30542 , \30543 , \30544 , \30545 , \30546 , \30547 , \30548 , \30549 , \30550 ,
         \30551 , \30552 , \30553 , \30554 , \30555 , \30556 , \30557 , \30558 , \30559 , \30560 ,
         \30561 , \30562 , \30563 , \30564 , \30565 , \30566 , \30567 , \30568 , \30569 , \30570 ,
         \30571 , \30572 , \30573 , \30574 , \30575 , \30576 , \30577 , \30578 , \30579 , \30580 ,
         \30581 , \30582 , \30583 , \30584 , \30585 , \30586 , \30587 , \30588 , \30589 , \30590 ,
         \30591 , \30592 , \30593 , \30594 , \30595 , \30596 , \30597 , \30598 , \30599 , \30600 ,
         \30601 , \30602 , \30603 , \30604 , \30605 , \30606 , \30607 , \30608 , \30609 , \30610 ,
         \30611 , \30612 , \30613 , \30614 , \30615 , \30616 , \30617 , \30618 , \30619 , \30620 ,
         \30621 , \30622 , \30623 , \30624 , \30625 , \30626 , \30627 , \30628 , \30629 , \30630 ,
         \30631 , \30632 , \30633 , \30634 , \30635 , \30636 , \30637 , \30638 , \30639 , \30640 ,
         \30641 , \30642 , \30643 , \30644 , \30645 , \30646 , \30647 , \30648 , \30649 , \30650 ,
         \30651 , \30652 , \30653 , \30654 , \30655 , \30656 , \30657 , \30658 , \30659 , \30660 ,
         \30661 , \30662 , \30663 , \30664 , \30665 , \30666 , \30667 , \30668 , \30669 , \30670 ,
         \30671 , \30672 , \30673 , \30674 , \30675 , \30676 , \30677 , \30678 , \30679 , \30680 ,
         \30681 , \30682 , \30683 , \30684 , \30685 , \30686 , \30687 , \30688 , \30689 , \30690 ,
         \30691 , \30692 , \30693 , \30694 , \30695 , \30696 , \30697 , \30698 , \30699 , \30700 ,
         \30701 , \30702 , \30703 , \30704 , \30705 , \30706 , \30707 , \30708 , \30709 , \30710 ,
         \30711 , \30712 , \30713 , \30714 , \30715 , \30716 , \30717 , \30718 , \30719 , \30720 ,
         \30721 , \30722 , \30723 , \30724 , \30725 , \30726 , \30727 , \30728 , \30729 , \30730 ,
         \30731 , \30732 , \30733 , \30734 , \30735 , \30736 , \30737 , \30738 , \30739 , \30740 ,
         \30741 , \30742 , \30743 , \30744 , \30745 , \30746 , \30747 , \30748 , \30749 , \30750 ,
         \30751 , \30752 , \30753 , \30754 , \30755 , \30756 , \30757 , \30758 , \30759 , \30760 ,
         \30761 , \30762 , \30763 , \30764 , \30765 , \30766 , \30767 , \30768 , \30769 , \30770 ,
         \30771 , \30772 , \30773 , \30774 , \30775 , \30776 , \30777 , \30778 , \30779 , \30780 ,
         \30781 , \30782 , \30783 , \30784 , \30785 , \30786 , \30787 , \30788 , \30789 , \30790 ,
         \30791 , \30792 , \30793 , \30794 , \30795 , \30796 , \30797 , \30798 , \30799 , \30800 ,
         \30801 , \30802 , \30803 , \30804 , \30805 , \30806 , \30807 , \30808 , \30809 , \30810 ,
         \30811 , \30812 , \30813 , \30814 , \30815 , \30816 , \30817 , \30818 , \30819 , \30820 ,
         \30821 , \30822 , \30823 , \30824 , \30825 , \30826 , \30827 , \30828 , \30829 , \30830 ,
         \30831 , \30832 , \30833 , \30834 , \30835 , \30836 , \30837 , \30838 , \30839 , \30840 ,
         \30841 , \30842 , \30843 , \30844 , \30845 , \30846 , \30847 , \30848 , \30849 , \30850 ,
         \30851 , \30852 , \30853 , \30854 , \30855 , \30856 , \30857 , \30858 , \30859 , \30860 ,
         \30861 , \30862 , \30863 , \30864 , \30865 , \30866 , \30867 , \30868 , \30869 , \30870 ,
         \30871 , \30872 , \30873 , \30874 , \30875 , \30876 , \30877 , \30878 , \30879 , \30880 ,
         \30881 , \30882 , \30883 , \30884 , \30885 , \30886 , \30887 , \30888 , \30889 , \30890 ,
         \30891 , \30892 , \30893 , \30894 , \30895 , \30896 , \30897 , \30898 , \30899 , \30900 ,
         \30901 , \30902 , \30903 , \30904 , \30905 , \30906 , \30907 , \30908 , \30909 , \30910 ,
         \30911 , \30912 , \30913 , \30914 , \30915 , \30916 , \30917 , \30918 , \30919 , \30920 ,
         \30921 , \30922 , \30923 , \30924 , \30925 , \30926 , \30927 , \30928 , \30929 , \30930 ,
         \30931 , \30932 , \30933 , \30934 , \30935 , \30936 , \30937 , \30938 , \30939 , \30940 ,
         \30941 , \30942 , \30943 , \30944 , \30945 , \30946 , \30947 , \30948 , \30949 , \30950 ,
         \30951 , \30952 , \30953 , \30954 , \30955 , \30956 , \30957 , \30958 , \30959 , \30960 ,
         \30961 , \30962 , \30963 , \30964 , \30965 , \30966 , \30967 , \30968 , \30969 , \30970 ,
         \30971 , \30972 , \30973 , \30974 , \30975 , \30976 , \30977 , \30978 , \30979 , \30980 ,
         \30981 , \30982 , \30983 , \30984 , \30985 , \30986 , \30987 , \30988 , \30989 , \30990 ,
         \30991 , \30992 , \30993 , \30994 , \30995 , \30996 , \30997 , \30998 , \30999 , \31000 ,
         \31001 , \31002 , \31003 , \31004 , \31005 , \31006 , \31007 , \31008 , \31009 , \31010 ,
         \31011 , \31012 , \31013 , \31014 , \31015 , \31016 , \31017 , \31018 , \31019 , \31020 ,
         \31021 , \31022 , \31023 , \31024 , \31025 , \31026 , \31027 , \31028 , \31029 , \31030 ,
         \31031 , \31032 , \31033 , \31034 , \31035 , \31036 , \31037 , \31038 , \31039 , \31040 ,
         \31041 , \31042 , \31043 , \31044 , \31045 , \31046 , \31047 , \31048 , \31049 , \31050 ,
         \31051 , \31052 , \31053 , \31054 , \31055 , \31056 , \31057 , \31058 , \31059 , \31060 ,
         \31061 , \31062 , \31063 , \31064 , \31065 , \31066 , \31067 , \31068 , \31069 , \31070 ,
         \31071 , \31072 , \31073 , \31074 , \31075 , \31076 , \31077 , \31078 , \31079 , \31080 ,
         \31081 , \31082 , \31083 , \31084 , \31085 , \31086 , \31087 , \31088 , \31089 , \31090 ,
         \31091 , \31092 , \31093 , \31094 , \31095 , \31096 , \31097 , \31098 , \31099 , \31100 ,
         \31101 , \31102 , \31103 , \31104 , \31105 , \31106 , \31107 , \31108 , \31109 , \31110 ,
         \31111 , \31112 , \31113 , \31114 , \31115 , \31116 , \31117 , \31118 , \31119 , \31120 ,
         \31121 , \31122 , \31123 , \31124 , \31125 , \31126 , \31127 , \31128 , \31129 , \31130 ,
         \31131 , \31132 , \31133 , \31134 , \31135 , \31136 , \31137 , \31138 , \31139 , \31140 ,
         \31141 , \31142 , \31143 , \31144 , \31145 , \31146 , \31147 , \31148 , \31149 , \31150 ,
         \31151 , \31152 , \31153 , \31154 , \31155 , \31156 , \31157 , \31158 , \31159 , \31160 ,
         \31161 , \31162 , \31163 , \31164 , \31165 , \31166 , \31167 , \31168 , \31169 , \31170 ,
         \31171 , \31172 , \31173 , \31174 , \31175 , \31176 , \31177 , \31178 , \31179 , \31180 ,
         \31181 , \31182 , \31183 , \31184 , \31185 , \31186 , \31187 , \31188 , \31189 , \31190 ,
         \31191 , \31192 , \31193 , \31194 , \31195 , \31196 , \31197 , \31198 , \31199 , \31200 ,
         \31201 , \31202 , \31203 , \31204 , \31205 , \31206 , \31207 , \31208 , \31209 , \31210 ,
         \31211 , \31212 , \31213 , \31214 , \31215 , \31216 , \31217 , \31218 , \31219 , \31220 ,
         \31221 , \31222 , \31223 , \31224 , \31225 , \31226 , \31227 , \31228 , \31229 , \31230 ,
         \31231 , \31232 , \31233 , \31234 , \31235 , \31236 , \31237 , \31238 , \31239 , \31240 ,
         \31241 , \31242 , \31243 , \31244 , \31245 , \31246 , \31247 , \31248 , \31249 , \31250 ,
         \31251 , \31252 , \31253 , \31254 , \31255 , \31256 , \31257 , \31258 , \31259 , \31260 ,
         \31261 , \31262 , \31263 , \31264 , \31265 , \31266 , \31267 , \31268 , \31269 , \31270 ,
         \31271 , \31272 , \31273 , \31274 , \31275 , \31276 , \31277 , \31278 , \31279 , \31280 ,
         \31281 , \31282 , \31283 , \31284 , \31285 , \31286 , \31287 , \31288 , \31289 , \31290 ,
         \31291 , \31292 , \31293 , \31294 , \31295 , \31296 , \31297 , \31298 , \31299 , \31300 ,
         \31301 , \31302 , \31303 , \31304 , \31305 , \31306 , \31307 , \31308 , \31309 , \31310 ,
         \31311 , \31312 , \31313 , \31314 , \31315 , \31316 , \31317 , \31318 , \31319 , \31320 ,
         \31321 , \31322 , \31323 , \31324 , \31325 , \31326 , \31327 , \31328 , \31329 , \31330 ,
         \31331 , \31332 , \31333 , \31334 , \31335 , \31336 , \31337 , \31338 , \31339 , \31340 ,
         \31341 , \31342 , \31343 , \31344 , \31345 , \31346 , \31347 , \31348 , \31349 , \31350 ,
         \31351 , \31352 , \31353 , \31354 , \31355 , \31356 , \31357 , \31358 , \31359 , \31360 ,
         \31361 , \31362 , \31363 , \31364 , \31365 , \31366 , \31367 , \31368 , \31369 , \31370 ,
         \31371 , \31372 , \31373 , \31374 , \31375 , \31376 , \31377 , \31378 , \31379 , \31380 ,
         \31381 , \31382 , \31383 , \31384 , \31385 , \31386 , \31387 , \31388 , \31389 , \31390 ,
         \31391 , \31392 , \31393 , \31394 , \31395 , \31396 , \31397 , \31398 , \31399 , \31400 ,
         \31401 , \31402 , \31403 , \31404 , \31405 , \31406 , \31407 , \31408 , \31409 , \31410 ,
         \31411 , \31412 , \31413 , \31414 , \31415 , \31416 , \31417 , \31418 , \31419 , \31420 ,
         \31421 , \31422 , \31423 , \31424 , \31425 , \31426 , \31427 , \31428 , \31429 , \31430 ,
         \31431 , \31432 , \31433 , \31434 , \31435 , \31436 , \31437 , \31438 , \31439 , \31440 ,
         \31441 , \31442 , \31443 , \31444 , \31445 , \31446 , \31447 , \31448 , \31449 , \31450 ,
         \31451 , \31452 , \31453 , \31454 , \31455 , \31456 , \31457 , \31458 , \31459 , \31460 ,
         \31461 , \31462 , \31463 , \31464 , \31465 , \31466 , \31467 , \31468 , \31469 , \31470 ,
         \31471 , \31472 , \31473 , \31474 , \31475 , \31476 , \31477 , \31478 , \31479 , \31480 ,
         \31481 , \31482 , \31483 , \31484 , \31485 , \31486 , \31487 , \31488 , \31489 , \31490 ,
         \31491 , \31492 , \31493 , \31494 , \31495 , \31496 , \31497 , \31498 , \31499 , \31500 ,
         \31501 , \31502 , \31503 , \31504 , \31505 , \31506 , \31507 , \31508 , \31509 , \31510 ,
         \31511 , \31512 , \31513 , \31514 , \31515 , \31516 , \31517 , \31518 , \31519 , \31520 ,
         \31521 , \31522 , \31523 , \31524 , \31525 , \31526 , \31527 , \31528 , \31529 , \31530 ,
         \31531 , \31532 , \31533 , \31534 , \31535 , \31536 , \31537 , \31538 , \31539 , \31540 ,
         \31541 , \31542 , \31543 , \31544 , \31545 , \31546 , \31547 , \31548 , \31549 , \31550 ,
         \31551 , \31552 , \31553 , \31554 , \31555 , \31556 , \31557 , \31558 , \31559 , \31560 ,
         \31561 , \31562 , \31563 , \31564 , \31565 , \31566 , \31567 , \31568 , \31569 , \31570 ,
         \31571 , \31572 , \31573 , \31574 , \31575 , \31576 , \31577 , \31578 , \31579 , \31580 ,
         \31581 , \31582 , \31583 , \31584 , \31585 , \31586 , \31587 , \31588 , \31589 , \31590 ,
         \31591 , \31592 , \31593 , \31594 , \31595 , \31596 , \31597 , \31598 , \31599 , \31600 ,
         \31601 , \31602 , \31603 , \31604 , \31605 , \31606 , \31607 , \31608 , \31609 , \31610 ,
         \31611 , \31612 , \31613 , \31614 , \31615 , \31616 , \31617 , \31618 , \31619 , \31620 ,
         \31621 , \31622 , \31623 , \31624 , \31625 , \31626 , \31627 , \31628 , \31629 , \31630 ,
         \31631 , \31632 , \31633 , \31634 , \31635 , \31636 , \31637 , \31638 , \31639 , \31640 ,
         \31641 , \31642 , \31643 , \31644 , \31645 , \31646 , \31647 , \31648 , \31649 , \31650 ,
         \31651 , \31652 , \31653 , \31654 , \31655 , \31656 , \31657 , \31658 , \31659 , \31660 ,
         \31661 , \31662 , \31663 , \31664 , \31665 , \31666 , \31667 , \31668 , \31669 , \31670 ,
         \31671 , \31672 , \31673 , \31674 , \31675 , \31676 , \31677 , \31678 , \31679 , \31680 ,
         \31681 , \31682 , \31683 , \31684 , \31685 , \31686 , \31687 , \31688 , \31689 , \31690 ,
         \31691 , \31692 , \31693 , \31694 , \31695 , \31696 , \31697 , \31698 , \31699 , \31700 ,
         \31701 , \31702 , \31703 , \31704 , \31705 , \31706 , \31707 , \31708 , \31709 , \31710 ,
         \31711 , \31712 , \31713 , \31714 , \31715 , \31716 , \31717 , \31718 , \31719 , \31720 ,
         \31721 , \31722 , \31723 , \31724 , \31725 , \31726 , \31727 , \31728 , \31729 , \31730 ,
         \31731 , \31732 , \31733 , \31734 , \31735 , \31736 , \31737 , \31738 , \31739 , \31740 ,
         \31741 , \31742 , \31743 , \31744 , \31745 , \31746 , \31747 , \31748 , \31749 , \31750 ,
         \31751 , \31752 , \31753 , \31754 , \31755 , \31756 , \31757 , \31758 , \31759 , \31760 ,
         \31761 , \31762 , \31763 , \31764 , \31765 , \31766 , \31767 , \31768 , \31769 , \31770 ,
         \31771 , \31772 , \31773 , \31774 , \31775 , \31776 , \31777 , \31778 , \31779 , \31780 ,
         \31781 , \31782 , \31783 , \31784 , \31785 , \31786 , \31787 , \31788 , \31789 , \31790 ,
         \31791 , \31792 , \31793 , \31794 , \31795 , \31796 , \31797 , \31798 , \31799 , \31800 ,
         \31801 , \31802 , \31803 , \31804 , \31805 , \31806 , \31807 , \31808 , \31809 , \31810 ,
         \31811 , \31812 , \31813 , \31814 , \31815 , \31816 , \31817 , \31818 , \31819 , \31820 ,
         \31821 , \31822 , \31823 , \31824 , \31825 , \31826 , \31827 , \31828 , \31829 , \31830 ,
         \31831 , \31832 , \31833 , \31834 , \31835 , \31836 , \31837 , \31838 , \31839 , \31840 ,
         \31841 , \31842 , \31843 , \31844 , \31845 , \31846 , \31847 , \31848 , \31849 , \31850 ,
         \31851 , \31852 , \31853 , \31854 , \31855 , \31856 , \31857 , \31858 , \31859 , \31860 ,
         \31861 , \31862 , \31863 , \31864 , \31865 , \31866 , \31867 , \31868 , \31869 , \31870 ,
         \31871 , \31872 , \31873 , \31874 , \31875 , \31876 , \31877 , \31878 , \31879 , \31880 ,
         \31881 , \31882 , \31883 , \31884 , \31885 , \31886 , \31887 , \31888 , \31889 , \31890 ,
         \31891 , \31892 , \31893 , \31894 , \31895 , \31896 , \31897 , \31898 , \31899 , \31900 ,
         \31901 , \31902 , \31903 , \31904 , \31905 , \31906 , \31907 , \31908 , \31909 , \31910 ,
         \31911 , \31912 , \31913 , \31914 , \31915 , \31916 , \31917 , \31918 , \31919 , \31920 ,
         \31921 , \31922 , \31923 , \31924 , \31925 , \31926 , \31927 , \31928 , \31929 , \31930 ,
         \31931 , \31932 , \31933 , \31934 , \31935 , \31936 , \31937 , \31938 , \31939 , \31940 ,
         \31941 , \31942 , \31943 , \31944 , \31945 , \31946 , \31947 , \31948 , \31949 , \31950 ,
         \31951 , \31952 , \31953 , \31954 , \31955 , \31956 , \31957 , \31958 , \31959 , \31960 ,
         \31961 , \31962 , \31963 , \31964 , \31965 , \31966 , \31967 , \31968 , \31969 , \31970 ,
         \31971 , \31972 , \31973 , \31974 , \31975 , \31976 , \31977 , \31978 , \31979 , \31980 ,
         \31981 , \31982 , \31983 , \31984 , \31985 , \31986 , \31987 , \31988 , \31989 , \31990 ,
         \31991 , \31992 , \31993 , \31994 , \31995 , \31996 , \31997 , \31998 , \31999 , \32000 ,
         \32001 , \32002 , \32003 , \32004 , \32005 , \32006 , \32007 , \32008 , \32009 , \32010 ,
         \32011 , \32012 , \32013 , \32014 , \32015 , \32016 , \32017 , \32018 , \32019 , \32020 ,
         \32021 , \32022 , \32023 , \32024 , \32025 , \32026 , \32027 , \32028 , \32029 , \32030 ,
         \32031 , \32032 , \32033 , \32034 , \32035 , \32036 , \32037 , \32038 , \32039 , \32040 ,
         \32041 , \32042 , \32043 , \32044 , \32045 , \32046 , \32047 , \32048 , \32049 , \32050 ,
         \32051 , \32052 , \32053 , \32054 , \32055 , \32056 , \32057 , \32058 , \32059 , \32060 ,
         \32061 , \32062 , \32063 , \32064 , \32065 , \32066 , \32067 , \32068 , \32069 , \32070 ,
         \32071 , \32072 , \32073 , \32074 , \32075 , \32076 , \32077 , \32078 , \32079 , \32080 ,
         \32081 , \32082 , \32083 , \32084 , \32085 , \32086 , \32087 , \32088 , \32089 , \32090 ,
         \32091 , \32092 , \32093 , \32094 , \32095 , \32096 , \32097 , \32098 , \32099 , \32100 ,
         \32101 , \32102 , \32103 , \32104 , \32105 , \32106 , \32107 , \32108 , \32109 , \32110 ,
         \32111 , \32112 , \32113 , \32114 , \32115 , \32116 , \32117 , \32118 , \32119 , \32120 ,
         \32121 , \32122 , \32123 , \32124 , \32125 , \32126 , \32127 , \32128 , \32129 , \32130 ,
         \32131 , \32132 , \32133 , \32134 , \32135 , \32136 , \32137 , \32138 , \32139 , \32140 ,
         \32141 , \32142 , \32143 , \32144 , \32145 , \32146 , \32147 , \32148 , \32149 , \32150 ,
         \32151 , \32152 , \32153 , \32154 , \32155 , \32156 , \32157 , \32158 , \32159 , \32160 ,
         \32161 , \32162 , \32163 , \32164 , \32165 , \32166 , \32167 , \32168 , \32169 , \32170 ,
         \32171 , \32172 , \32173 , \32174 , \32175 , \32176 , \32177 , \32178 , \32179 , \32180 ,
         \32181 , \32182 , \32183 , \32184 , \32185 , \32186 , \32187 , \32188 , \32189 , \32190 ,
         \32191 , \32192 , \32193 , \32194 , \32195 , \32196 , \32197 , \32198 , \32199 , \32200 ,
         \32201 , \32202 , \32203 , \32204 , \32205 , \32206 , \32207 , \32208 , \32209 , \32210 ,
         \32211 , \32212 , \32213 , \32214 , \32215 , \32216 , \32217 , \32218 , \32219 , \32220 ,
         \32221 , \32222 , \32223 , \32224 , \32225 , \32226 , \32227 , \32228 , \32229 , \32230 ,
         \32231 , \32232 , \32233 , \32234 , \32235 , \32236 , \32237 , \32238 , \32239 , \32240 ,
         \32241 , \32242 , \32243 , \32244 , \32245 , \32246 , \32247 , \32248 , \32249 , \32250 ,
         \32251 , \32252 , \32253 , \32254 , \32255 , \32256 , \32257 , \32258 , \32259 , \32260 ,
         \32261 , \32262 , \32263 , \32264 , \32265 , \32266 , \32267 , \32268 , \32269 , \32270 ,
         \32271 , \32272 , \32273 , \32274 , \32275 , \32276 , \32277 , \32278 , \32279 , \32280 ,
         \32281 , \32282 , \32283 , \32284 , \32285 , \32286 , \32287 , \32288 , \32289 , \32290 ,
         \32291 , \32292 , \32293 , \32294 , \32295 , \32296 , \32297 , \32298 , \32299 , \32300 ,
         \32301 , \32302 , \32303 , \32304 , \32305 , \32306 , \32307 , \32308 , \32309 , \32310 ,
         \32311 , \32312 , \32313 , \32314 , \32315 , \32316 , \32317 , \32318 , \32319 , \32320 ,
         \32321 , \32322 , \32323 , \32324 , \32325 , \32326 , \32327 , \32328 , \32329 , \32330 ,
         \32331 , \32332 , \32333 , \32334 , \32335 , \32336 , \32337 , \32338 , \32339 , \32340 ,
         \32341 , \32342 , \32343 , \32344 , \32345 , \32346 , \32347 , \32348 , \32349 , \32350 ,
         \32351 , \32352 , \32353 , \32354 , \32355 , \32356 , \32357 , \32358 , \32359 , \32360 ,
         \32361 , \32362 , \32363 , \32364 , \32365 , \32366 , \32367 , \32368 , \32369 , \32370 ,
         \32371 , \32372 , \32373 , \32374 , \32375 , \32376 , \32377 , \32378 , \32379 , \32380 ,
         \32381 , \32382 , \32383 , \32384 , \32385 , \32386 , \32387 , \32388 , \32389 , \32390 ,
         \32391 , \32392 , \32393 , \32394 , \32395 , \32396 , \32397 , \32398 , \32399 , \32400 ,
         \32401 , \32402 , \32403 , \32404 , \32405 , \32406 , \32407 , \32408 , \32409 , \32410 ,
         \32411 , \32412 , \32413 , \32414 , \32415 , \32416 , \32417 , \32418 , \32419 , \32420 ,
         \32421 , \32422 , \32423 , \32424 , \32425 , \32426 , \32427 , \32428 , \32429 , \32430 ,
         \32431 , \32432 , \32433 , \32434 , \32435 , \32436 , \32437 , \32438 , \32439 , \32440 ,
         \32441 , \32442 , \32443 , \32444 , \32445 , \32446 , \32447 , \32448 , \32449 , \32450 ,
         \32451 , \32452 , \32453 , \32454 , \32455 , \32456 , \32457 , \32458 , \32459 , \32460 ,
         \32461 , \32462 , \32463 , \32464 , \32465 , \32466 , \32467 , \32468 , \32469 , \32470 ,
         \32471 , \32472 , \32473 , \32474 , \32475 , \32476 , \32477 , \32478 , \32479 , \32480 ,
         \32481 , \32482 , \32483 , \32484 , \32485 , \32486 , \32487 , \32488 , \32489 , \32490 ,
         \32491 , \32492 , \32493 , \32494 , \32495 , \32496 , \32497 , \32498 , \32499 , \32500 ,
         \32501 , \32502 , \32503 , \32504 , \32505 , \32506 , \32507 , \32508 , \32509 , \32510 ,
         \32511 , \32512 , \32513 , \32514 , \32515 , \32516 , \32517 , \32518 , \32519 , \32520 ,
         \32521 , \32522 , \32523 , \32524 , \32525 , \32526 , \32527 , \32528 , \32529 , \32530 ,
         \32531 , \32532 , \32533 , \32534 , \32535 , \32536 , \32537 , \32538 , \32539 , \32540 ,
         \32541 , \32542 , \32543 , \32544 , \32545 , \32546 , \32547 , \32548 , \32549 , \32550 ,
         \32551 , \32552 , \32553 , \32554 , \32555 , \32556 , \32557 , \32558 , \32559 , \32560 ,
         \32561 , \32562 , \32563 , \32564 , \32565 , \32566 , \32567 , \32568 , \32569 , \32570 ,
         \32571 , \32572 , \32573 , \32574 , \32575 , \32576 , \32577 , \32578 , \32579 , \32580 ,
         \32581 , \32582 , \32583 , \32584 , \32585 , \32586 , \32587 , \32588 , \32589 , \32590 ,
         \32591 , \32592 , \32593 , \32594 , \32595 , \32596 , \32597 , \32598 , \32599 , \32600 ,
         \32601 , \32602 , \32603 , \32604 , \32605 , \32606 , \32607 , \32608 , \32609 , \32610 ,
         \32611 , \32612 , \32613 , \32614 , \32615 , \32616 , \32617 , \32618 , \32619 , \32620 ,
         \32621 , \32622 , \32623 , \32624 , \32625 , \32626 , \32627 , \32628 , \32629 , \32630 ,
         \32631 , \32632 , \32633 , \32634 , \32635 , \32636 , \32637 , \32638 , \32639 , \32640 ,
         \32641 , \32642 , \32643 , \32644 , \32645 , \32646 , \32647 , \32648 , \32649 , \32650 ,
         \32651 , \32652 , \32653 , \32654 , \32655 , \32656 , \32657 , \32658 , \32659 , \32660 ,
         \32661 , \32662 , \32663 , \32664 , \32665 , \32666 , \32667 , \32668 , \32669 , \32670 ,
         \32671 , \32672 , \32673 , \32674 , \32675 , \32676 , \32677 , \32678 , \32679 , \32680 ,
         \32681 , \32682 , \32683 , \32684 , \32685 , \32686 , \32687 , \32688 , \32689 , \32690 ,
         \32691 , \32692 , \32693 , \32694 , \32695 , \32696 , \32697 , \32698 , \32699 , \32700 ,
         \32701 , \32702 , \32703 , \32704 , \32705 , \32706 , \32707 , \32708 , \32709 , \32710 ,
         \32711 , \32712 , \32713 , \32714 , \32715 , \32716 , \32717 , \32718 , \32719 , \32720 ,
         \32721 , \32722 , \32723 , \32724 , \32725 , \32726 , \32727 , \32728 , \32729 , \32730 ,
         \32731 , \32732 , \32733 , \32734 , \32735 , \32736 , \32737 , \32738 , \32739 , \32740 ,
         \32741 , \32742 , \32743 , \32744 , \32745 , \32746 , \32747 , \32748 , \32749 , \32750 ,
         \32751 , \32752 , \32753 , \32754 , \32755 , \32756 , \32757 , \32758 , \32759 , \32760 ,
         \32761 , \32762 , \32763 , \32764 , \32765 , \32766 , \32767 , \32768 , \32769 , \32770 ,
         \32771 , \32772 , \32773 , \32774 , \32775 , \32776 , \32777 , \32778 , \32779 , \32780 ,
         \32781 , \32782 , \32783 , \32784 , \32785 , \32786 , \32787 , \32788 , \32789 , \32790 ,
         \32791 , \32792 , \32793 , \32794 , \32795 , \32796 , \32797 , \32798 , \32799 , \32800 ,
         \32801 , \32802 , \32803 , \32804 , \32805 , \32806 , \32807 , \32808 , \32809 , \32810 ,
         \32811 , \32812 , \32813 , \32814 , \32815 , \32816 , \32817 , \32818 , \32819 , \32820 ,
         \32821 , \32822 , \32823 , \32824 , \32825 , \32826 , \32827 , \32828 , \32829 , \32830 ,
         \32831 , \32832 , \32833 , \32834 , \32835 , \32836 , \32837 , \32838 , \32839 , \32840 ,
         \32841 , \32842 , \32843 , \32844 , \32845 , \32846 , \32847 , \32848 , \32849 , \32850 ,
         \32851 , \32852 , \32853 , \32854 , \32855 , \32856 , \32857 , \32858 , \32859 , \32860 ,
         \32861 , \32862 , \32863 , \32864 , \32865 , \32866 , \32867 , \32868 , \32869 , \32870 ,
         \32871 , \32872 , \32873 , \32874 , \32875 , \32876 , \32877 , \32878 , \32879 , \32880 ,
         \32881 , \32882 , \32883 , \32884 , \32885 , \32886 , \32887 , \32888 , \32889 , \32890 ,
         \32891 , \32892 , \32893 , \32894 , \32895 , \32896 , \32897 , \32898 , \32899 , \32900 ,
         \32901 , \32902 , \32903 , \32904 , \32905 , \32906 , \32907 , \32908 , \32909 , \32910 ,
         \32911 , \32912 , \32913 , \32914 , \32915 , \32916 , \32917 , \32918 , \32919 , \32920 ,
         \32921 , \32922 , \32923 , \32924 , \32925 , \32926 , \32927 , \32928 , \32929 , \32930 ,
         \32931 , \32932 , \32933 , \32934 , \32935 , \32936 , \32937 , \32938 , \32939 , \32940 ,
         \32941 , \32942 , \32943 , \32944 , \32945 , \32946 , \32947 , \32948 , \32949 , \32950 ,
         \32951 , \32952 , \32953 , \32954 , \32955 , \32956 , \32957 , \32958 , \32959 , \32960 ,
         \32961 , \32962 , \32963 , \32964 , \32965 , \32966 , \32967 , \32968 , \32969 , \32970 ,
         \32971 , \32972 , \32973 , \32974 , \32975 , \32976 , \32977 , \32978 , \32979 , \32980 ,
         \32981 , \32982 , \32983 , \32984 , \32985 , \32986 , \32987 , \32988 , \32989 , \32990 ,
         \32991 , \32992 , \32993 , \32994 , \32995 , \32996 , \32997 , \32998 , \32999 , \33000 ,
         \33001 , \33002 , \33003 , \33004 , \33005 , \33006 , \33007 , \33008 , \33009 , \33010 ,
         \33011 , \33012 , \33013 , \33014 , \33015 , \33016 , \33017 , \33018 , \33019 , \33020 ,
         \33021 , \33022 , \33023 , \33024 , \33025 , \33026 , \33027 , \33028 , \33029 , \33030 ,
         \33031 , \33032 , \33033 , \33034 , \33035 , \33036 , \33037 , \33038 , \33039 , \33040 ,
         \33041 , \33042 , \33043 , \33044 , \33045 , \33046 , \33047 , \33048 , \33049 , \33050 ,
         \33051 , \33052 , \33053 , \33054 , \33055 , \33056 , \33057 , \33058 , \33059 , \33060 ,
         \33061 , \33062 , \33063 , \33064 , \33065 , \33066 , \33067 , \33068 , \33069 , \33070 ,
         \33071 , \33072 , \33073 , \33074 , \33075 , \33076 , \33077 , \33078 , \33079 , \33080 ,
         \33081 , \33082 , \33083 , \33084 , \33085 , \33086 , \33087 , \33088 , \33089 , \33090 ,
         \33091 , \33092 , \33093 , \33094 , \33095 , \33096 , \33097 , \33098 , \33099 , \33100 ,
         \33101 , \33102 , \33103 , \33104 , \33105 , \33106 , \33107 , \33108 , \33109 , \33110 ,
         \33111 , \33112 , \33113 , \33114 , \33115 , \33116 , \33117 , \33118 , \33119 , \33120 ,
         \33121 , \33122 , \33123 , \33124 , \33125 , \33126 , \33127 , \33128 , \33129 , \33130 ,
         \33131 , \33132 , \33133 , \33134 , \33135 , \33136 , \33137 , \33138 , \33139 , \33140 ,
         \33141 , \33142 , \33143 , \33144 , \33145 , \33146 , \33147 , \33148 , \33149 , \33150 ,
         \33151 , \33152 , \33153 , \33154 , \33155 , \33156 , \33157 , \33158 , \33159 , \33160 ,
         \33161 , \33162 , \33163 , \33164 , \33165 , \33166 , \33167 , \33168 , \33169 , \33170 ,
         \33171 , \33172 , \33173 , \33174 , \33175 , \33176 , \33177 , \33178 , \33179 , \33180 ,
         \33181 , \33182 , \33183 , \33184 , \33185 , \33186 , \33187 , \33188 , \33189 , \33190 ,
         \33191 , \33192 , \33193 , \33194 , \33195 , \33196 , \33197 , \33198 , \33199 , \33200 ,
         \33201 , \33202 , \33203 , \33204 , \33205 , \33206 , \33207 , \33208 , \33209 , \33210 ,
         \33211 , \33212 , \33213 , \33214 , \33215 , \33216 , \33217 , \33218 , \33219 , \33220 ,
         \33221 , \33222 , \33223 , \33224 , \33225 , \33226 , \33227 , \33228 , \33229 , \33230 ,
         \33231 , \33232 , \33233 , \33234 , \33235 , \33236 , \33237 , \33238 , \33239 , \33240 ,
         \33241 , \33242 , \33243 , \33244 , \33245 , \33246 , \33247 , \33248 , \33249 , \33250 ,
         \33251 , \33252 , \33253 , \33254 , \33255 , \33256 , \33257 , \33258 , \33259 , \33260 ,
         \33261 , \33262 , \33263 , \33264 , \33265 , \33266 , \33267 , \33268 , \33269 , \33270 ,
         \33271 , \33272 , \33273 , \33274 , \33275 , \33276 , \33277 , \33278 , \33279 , \33280 ,
         \33281 , \33282 , \33283 , \33284 , \33285 , \33286 , \33287 , \33288 , \33289 , \33290 ,
         \33291 , \33292 , \33293 , \33294 , \33295 , \33296 , \33297 , \33298 , \33299 , \33300 ,
         \33301 , \33302 , \33303 , \33304 , \33305 , \33306 , \33307 , \33308 , \33309 , \33310 ,
         \33311 , \33312 , \33313 , \33314 , \33315 , \33316 , \33317 , \33318 , \33319 , \33320 ,
         \33321 , \33322 , \33323 , \33324 , \33325 , \33326 , \33327 , \33328 , \33329 , \33330 ,
         \33331 , \33332 , \33333 , \33334 , \33335 , \33336 , \33337 , \33338 , \33339 , \33340 ,
         \33341 , \33342 , \33343 , \33344 , \33345 , \33346 , \33347 , \33348 , \33349 , \33350 ,
         \33351 , \33352 , \33353 , \33354 , \33355 , \33356 , \33357 , \33358 , \33359 , \33360 ,
         \33361 , \33362 , \33363 , \33364 , \33365 , \33366 , \33367 , \33368 , \33369 , \33370 ,
         \33371 , \33372 , \33373 , \33374 , \33375 , \33376 , \33377 , \33378 , \33379 , \33380 ,
         \33381 , \33382 , \33383 , \33384 , \33385 , \33386 , \33387 , \33388 , \33389 , \33390 ,
         \33391 , \33392 , \33393 , \33394 , \33395 , \33396 , \33397 , \33398 , \33399 , \33400 ,
         \33401 , \33402 , \33403 , \33404 , \33405 , \33406 , \33407 , \33408 , \33409 , \33410 ,
         \33411 , \33412 , \33413 , \33414 , \33415 , \33416 , \33417 , \33418 , \33419 , \33420 ,
         \33421 , \33422 , \33423 , \33424 , \33425 , \33426 , \33427 , \33428 , \33429 , \33430 ,
         \33431 , \33432 , \33433 , \33434 , \33435 , \33436 , \33437 , \33438 , \33439 , \33440 ,
         \33441 , \33442 , \33443 , \33444 , \33445 , \33446 , \33447 , \33448 , \33449 , \33450 ,
         \33451 , \33452 , \33453 , \33454 , \33455 , \33456 , \33457 , \33458 , \33459 , \33460 ,
         \33461 , \33462 , \33463 , \33464 , \33465 , \33466 , \33467 , \33468 , \33469 , \33470 ,
         \33471 , \33472 , \33473 , \33474 , \33475 , \33476 , \33477 , \33478 , \33479 , \33480 ,
         \33481 , \33482 , \33483 , \33484 , \33485 , \33486 , \33487 , \33488 , \33489 , \33490 ,
         \33491 , \33492 , \33493 , \33494 , \33495 , \33496 , \33497 , \33498 , \33499 , \33500 ,
         \33501 , \33502 , \33503 , \33504 , \33505 , \33506 , \33507 , \33508 , \33509 , \33510 ,
         \33511 , \33512 , \33513 , \33514 , \33515 , \33516 , \33517 , \33518 , \33519 , \33520 ,
         \33521 , \33522 , \33523 , \33524 , \33525 , \33526 , \33527 , \33528 , \33529 , \33530 ,
         \33531 , \33532 , \33533 , \33534 , \33535 , \33536 , \33537 , \33538 , \33539 , \33540 ,
         \33541 , \33542 , \33543 , \33544 , \33545 , \33546 , \33547 , \33548 , \33549 , \33550 ,
         \33551 , \33552 , \33553 , \33554 , \33555 , \33556 , \33557 , \33558 , \33559 , \33560 ,
         \33561 , \33562 , \33563 , \33564 , \33565 , \33566 , \33567 , \33568 , \33569 , \33570 ,
         \33571 , \33572 , \33573 , \33574 , \33575 , \33576 , \33577 , \33578 , \33579 , \33580 ,
         \33581 , \33582 , \33583 , \33584 , \33585 , \33586 , \33587 , \33588 , \33589 , \33590 ,
         \33591 , \33592 , \33593 , \33594 , \33595 , \33596 , \33597 , \33598 , \33599 , \33600 ,
         \33601 , \33602 , \33603 , \33604 , \33605 , \33606 , \33607 , \33608 , \33609 , \33610 ,
         \33611 , \33612 , \33613 , \33614 , \33615 , \33616 , \33617 , \33618 , \33619 , \33620 ,
         \33621 , \33622 , \33623 , \33624 , \33625 , \33626 , \33627 , \33628 , \33629 , \33630 ,
         \33631 , \33632 , \33633 , \33634 , \33635 , \33636 , \33637 , \33638 , \33639 , \33640 ,
         \33641 , \33642 , \33643 , \33644 , \33645 , \33646 , \33647 , \33648 , \33649 , \33650 ,
         \33651 , \33652 , \33653 , \33654 , \33655 , \33656 , \33657 , \33658 , \33659 , \33660 ,
         \33661 , \33662 , \33663 , \33664 , \33665 , \33666 , \33667 , \33668 , \33669 , \33670 ,
         \33671 , \33672 , \33673 , \33674 , \33675 , \33676 , \33677 , \33678 , \33679 , \33680 ,
         \33681 , \33682 , \33683 , \33684 , \33685 , \33686 , \33687 , \33688 , \33689 , \33690 ,
         \33691 , \33692 , \33693 , \33694 , \33695 , \33696 , \33697 , \33698 , \33699 , \33700 ,
         \33701 , \33702 , \33703 , \33704 , \33705 , \33706 , \33707 , \33708 , \33709 , \33710 ,
         \33711 , \33712 , \33713 , \33714 , \33715 , \33716 , \33717 , \33718 , \33719 , \33720 ,
         \33721 , \33722 , \33723 , \33724 , \33725 , \33726 , \33727 , \33728 , \33729 , \33730 ,
         \33731 , \33732 , \33733 , \33734 , \33735 , \33736 , \33737 , \33738 , \33739 , \33740 ,
         \33741 , \33742 , \33743 , \33744 , \33745 , \33746 , \33747 , \33748 , \33749 , \33750 ,
         \33751 , \33752 , \33753 , \33754 , \33755 , \33756 , \33757 , \33758 , \33759 , \33760 ,
         \33761 , \33762 , \33763 , \33764 , \33765 , \33766 , \33767 , \33768 , \33769 , \33770 ,
         \33771 , \33772 , \33773 , \33774 , \33775 , \33776 , \33777 , \33778 , \33779 , \33780 ,
         \33781 , \33782 , \33783 , \33784 , \33785 , \33786 , \33787 , \33788 , \33789 , \33790 ,
         \33791 , \33792 , \33793 , \33794 , \33795 , \33796 , \33797 , \33798 , \33799 , \33800 ,
         \33801 , \33802 , \33803 , \33804 , \33805 , \33806 , \33807 , \33808 , \33809 , \33810 ,
         \33811 , \33812 , \33813 , \33814 , \33815 , \33816 , \33817 , \33818 , \33819 , \33820 ,
         \33821 , \33822 , \33823 , \33824 , \33825 , \33826 , \33827 , \33828 , \33829 , \33830 ,
         \33831 , \33832 , \33833 , \33834 , \33835 , \33836 , \33837 , \33838 , \33839 , \33840 ,
         \33841 , \33842 , \33843 , \33844 , \33845 , \33846 , \33847 , \33848 , \33849 , \33850 ,
         \33851 , \33852 , \33853 , \33854 , \33855 , \33856 , \33857 , \33858 , \33859 , \33860 ,
         \33861 , \33862 , \33863 , \33864 , \33865 , \33866 , \33867 , \33868 , \33869 , \33870 ,
         \33871 , \33872 , \33873 , \33874 , \33875 , \33876 , \33877 , \33878 , \33879 , \33880 ,
         \33881 , \33882 , \33883 , \33884 , \33885 , \33886 , \33887 , \33888 , \33889 , \33890 ,
         \33891 , \33892 , \33893 , \33894 , \33895 , \33896 , \33897 , \33898 , \33899 , \33900 ,
         \33901 , \33902 , \33903 , \33904 , \33905 , \33906 , \33907 , \33908 , \33909 , \33910 ,
         \33911 , \33912 , \33913 , \33914 , \33915 , \33916 , \33917 , \33918 , \33919 , \33920 ,
         \33921 , \33922 , \33923 , \33924 , \33925 , \33926 , \33927 , \33928 , \33929 , \33930 ,
         \33931 , \33932 , \33933 , \33934 , \33935 , \33936 , \33937 , \33938 , \33939 , \33940 ,
         \33941 , \33942 , \33943 , \33944 , \33945 , \33946 , \33947 , \33948 , \33949 , \33950 ,
         \33951 , \33952 , \33953 , \33954 , \33955 , \33956 , \33957 , \33958 , \33959 , \33960 ,
         \33961 , \33962 , \33963 , \33964 , \33965 , \33966 , \33967 , \33968 , \33969 , \33970 ,
         \33971 , \33972 , \33973 , \33974 , \33975 , \33976 , \33977 , \33978 , \33979 , \33980 ,
         \33981 , \33982 , \33983 , \33984 , \33985 , \33986 , \33987 , \33988 , \33989 , \33990 ,
         \33991 , \33992 , \33993 , \33994 , \33995 , \33996 , \33997 , \33998 , \33999 , \34000 ,
         \34001 , \34002 , \34003 , \34004 , \34005 , \34006 , \34007 , \34008 , \34009 , \34010 ,
         \34011 , \34012 , \34013 , \34014 , \34015 , \34016 , \34017 , \34018 , \34019 , \34020 ,
         \34021 , \34022 , \34023 , \34024 , \34025 , \34026 , \34027 , \34028 , \34029 , \34030 ,
         \34031 , \34032 , \34033 , \34034 , \34035 , \34036 , \34037 , \34038 , \34039 , \34040 ,
         \34041 , \34042 , \34043 , \34044 , \34045 , \34046 , \34047 , \34048 , \34049 , \34050 ,
         \34051 , \34052 , \34053 , \34054 , \34055 , \34056 , \34057 , \34058 , \34059 , \34060 ,
         \34061 , \34062 , \34063 , \34064 , \34065 , \34066 , \34067 , \34068 , \34069 , \34070 ,
         \34071 , \34072 , \34073 , \34074 , \34075 , \34076 , \34077 , \34078 , \34079 , \34080 ,
         \34081 , \34082 , \34083 , \34084 , \34085 , \34086 , \34087 , \34088 , \34089 , \34090 ,
         \34091 , \34092 , \34093 , \34094 , \34095 , \34096 , \34097 , \34098 , \34099 , \34100 ,
         \34101 , \34102 , \34103 , \34104 , \34105 , \34106 , \34107 , \34108 , \34109 , \34110 ,
         \34111 , \34112 , \34113 , \34114 , \34115 , \34116 , \34117 , \34118 , \34119 , \34120 ,
         \34121 , \34122 , \34123 , \34124 , \34125 , \34126 , \34127 , \34128 , \34129 , \34130 ,
         \34131 , \34132 , \34133 , \34134 , \34135 , \34136 , \34137 , \34138 , \34139 , \34140 ,
         \34141 , \34142 , \34143 , \34144 , \34145 , \34146 , \34147 , \34148 , \34149 , \34150 ,
         \34151 , \34152 , \34153 , \34154 , \34155 , \34156 , \34157 , \34158 , \34159 , \34160 ,
         \34161 , \34162 , \34163 , \34164 , \34165 , \34166 , \34167 , \34168 , \34169 , \34170 ,
         \34171 , \34172 , \34173 , \34174 , \34175 , \34176 , \34177 , \34178 , \34179 , \34180 ,
         \34181 , \34182 , \34183 , \34184 , \34185 , \34186 , \34187 , \34188 , \34189 , \34190 ,
         \34191 , \34192 , \34193 , \34194 , \34195 , \34196 , \34197 , \34198 , \34199 , \34200 ,
         \34201 , \34202 , \34203 , \34204 , \34205 , \34206 , \34207 , \34208 , \34209 , \34210 ,
         \34211 , \34212 , \34213 , \34214 , \34215 , \34216 , \34217 , \34218 , \34219 , \34220 ,
         \34221 , \34222 , \34223 , \34224 , \34225 , \34226 , \34227 , \34228 , \34229 , \34230 ,
         \34231 , \34232 , \34233 , \34234 , \34235 , \34236 , \34237 , \34238 , \34239 , \34240 ,
         \34241 , \34242 , \34243 , \34244 , \34245 , \34246 , \34247 , \34248 , \34249 , \34250 ,
         \34251 , \34252 , \34253 , \34254 , \34255 , \34256 , \34257 , \34258 , \34259 , \34260 ,
         \34261 , \34262 , \34263 , \34264 , \34265 , \34266 , \34267 , \34268 , \34269 , \34270 ,
         \34271 , \34272 , \34273 , \34274 , \34275 , \34276 , \34277 , \34278 , \34279 , \34280 ,
         \34281 , \34282 , \34283 , \34284 , \34285 , \34286 , \34287 , \34288 , \34289 , \34290 ,
         \34291 , \34292 , \34293 , \34294 , \34295 , \34296 , \34297 , \34298 , \34299 , \34300 ,
         \34301 , \34302 , \34303 , \34304 , \34305 , \34306 , \34307 , \34308 , \34309 , \34310 ,
         \34311 , \34312 , \34313 , \34314 , \34315 , \34316 , \34317 , \34318 , \34319 , \34320 ,
         \34321 , \34322 , \34323 , \34324 , \34325 , \34326 , \34327 , \34328 , \34329 , \34330 ,
         \34331 , \34332 , \34333 , \34334 , \34335 , \34336 , \34337 , \34338 , \34339 , \34340 ,
         \34341 , \34342 , \34343 , \34344 , \34345 , \34346 , \34347 , \34348 , \34349 , \34350 ,
         \34351 , \34352 , \34353 , \34354 , \34355 , \34356 , \34357 , \34358 , \34359 , \34360 ,
         \34361 , \34362 , \34363 , \34364 , \34365 , \34366 , \34367 , \34368 , \34369 , \34370 ,
         \34371 , \34372 , \34373 , \34374 , \34375 , \34376 , \34377 , \34378 , \34379 , \34380 ,
         \34381 , \34382 , \34383 , \34384 , \34385 , \34386 , \34387 , \34388 , \34389 , \34390 ,
         \34391 , \34392 , \34393 , \34394 , \34395 , \34396 , \34397 , \34398 , \34399 , \34400 ,
         \34401 , \34402 , \34403 , \34404 , \34405 , \34406 , \34407 , \34408 , \34409 , \34410 ,
         \34411 , \34412 , \34413 , \34414 , \34415 , \34416 , \34417 , \34418 , \34419 , \34420 ,
         \34421 , \34422 , \34423 , \34424 , \34425 , \34426 , \34427 , \34428 , \34429 , \34430 ,
         \34431 , \34432 , \34433 , \34434 , \34435 , \34436 , \34437 , \34438 , \34439 , \34440 ,
         \34441 , \34442 , \34443 , \34444 , \34445 , \34446 , \34447 , \34448 , \34449 , \34450 ,
         \34451 , \34452 , \34453 , \34454 , \34455 , \34456 , \34457 , \34458 , \34459 , \34460 ,
         \34461 , \34462 , \34463 , \34464 , \34465 , \34466 , \34467 , \34468 , \34469 , \34470 ,
         \34471 , \34472 , \34473 , \34474 , \34475 , \34476 , \34477 , \34478 , \34479 , \34480 ,
         \34481 , \34482 , \34483 , \34484 , \34485 , \34486 , \34487 , \34488 , \34489 , \34490 ,
         \34491 , \34492 , \34493 , \34494 , \34495 , \34496 , \34497 , \34498 , \34499 , \34500 ,
         \34501 , \34502 , \34503 , \34504 , \34505 , \34506 , \34507 , \34508 , \34509 , \34510 ,
         \34511 , \34512 , \34513 , \34514 , \34515 , \34516 , \34517 , \34518 , \34519 , \34520 ,
         \34521 , \34522 , \34523 , \34524 , \34525 , \34526 , \34527 , \34528 , \34529 , \34530 ,
         \34531 , \34532 , \34533 , \34534 , \34535 , \34536 , \34537 , \34538 , \34539 , \34540 ,
         \34541 , \34542 , \34543 , \34544 , \34545 , \34546 , \34547 , \34548 , \34549 , \34550 ,
         \34551 , \34552 , \34553 , \34554 , \34555 , \34556 , \34557 , \34558 , \34559 , \34560 ,
         \34561 , \34562 , \34563 , \34564 , \34565 , \34566 , \34567 , \34568 , \34569 , \34570 ,
         \34571 , \34572 , \34573 , \34574 , \34575 , \34576 , \34577 , \34578 , \34579 , \34580 ,
         \34581 , \34582 , \34583 , \34584 , \34585 , \34586 , \34587 , \34588 , \34589 , \34590 ,
         \34591 , \34592 , \34593 , \34594 , \34595 , \34596 , \34597 , \34598 , \34599 , \34600 ,
         \34601 , \34602 , \34603 , \34604 , \34605 , \34606 , \34607 , \34608 , \34609 , \34610 ,
         \34611 , \34612 , \34613 , \34614 , \34615 , \34616 , \34617 , \34618 , \34619 , \34620 ,
         \34621 , \34622 , \34623 , \34624 , \34625 , \34626 , \34627 , \34628 , \34629 , \34630 ,
         \34631 , \34632 , \34633 , \34634 , \34635 , \34636 , \34637 , \34638 , \34639 , \34640 ,
         \34641 , \34642 , \34643 , \34644 , \34645 , \34646 , \34647 , \34648 , \34649 , \34650 ,
         \34651 , \34652 , \34653 , \34654 , \34655 , \34656 , \34657 , \34658 , \34659 , \34660 ,
         \34661 , \34662 , \34663 , \34664 , \34665 , \34666 , \34667 , \34668 , \34669 , \34670 ,
         \34671 , \34672 , \34673 , \34674 , \34675 , \34676 , \34677 , \34678 , \34679 , \34680 ,
         \34681 , \34682 , \34683 , \34684 , \34685 , \34686 , \34687 , \34688 , \34689 , \34690 ,
         \34691 , \34692 , \34693 , \34694 , \34695 , \34696 , \34697 , \34698 , \34699 , \34700 ,
         \34701 , \34702 , \34703 , \34704 , \34705 , \34706 , \34707 , \34708 , \34709 , \34710 ,
         \34711 , \34712 , \34713 , \34714 , \34715 , \34716 , \34717 , \34718 , \34719 , \34720 ,
         \34721 , \34722 , \34723 , \34724 , \34725 , \34726 , \34727 , \34728 , \34729 , \34730 ,
         \34731 , \34732 , \34733 , \34734 , \34735 , \34736 , \34737 , \34738 , \34739 , \34740 ,
         \34741 , \34742 , \34743 , \34744 , \34745 , \34746 , \34747 , \34748 , \34749 , \34750 ,
         \34751 , \34752 , \34753 , \34754 , \34755 , \34756 , \34757 , \34758 , \34759 , \34760 ,
         \34761 , \34762 , \34763 , \34764 , \34765 , \34766 , \34767 , \34768 , \34769 , \34770 ,
         \34771 , \34772 , \34773 , \34774 , \34775 , \34776 , \34777 , \34778 , \34779 , \34780 ,
         \34781 , \34782 , \34783 , \34784 , \34785 , \34786 , \34787 , \34788 , \34789 , \34790 ,
         \34791 , \34792 , \34793 , \34794 , \34795 , \34796 , \34797 , \34798 , \34799 , \34800 ,
         \34801 , \34802 , \34803 , \34804 , \34805 , \34806 , \34807 , \34808 , \34809 , \34810 ,
         \34811 , \34812 , \34813 , \34814 , \34815 , \34816 , \34817 , \34818 , \34819 , \34820 ,
         \34821 , \34822 , \34823 , \34824 , \34825 , \34826 , \34827 , \34828 , \34829 , \34830 ,
         \34831 , \34832 , \34833 , \34834 , \34835 , \34836 , \34837 , \34838 , \34839 , \34840 ,
         \34841 , \34842 , \34843 , \34844 , \34845 , \34846 , \34847 , \34848 , \34849 , \34850 ,
         \34851 , \34852 , \34853 , \34854 , \34855 , \34856 , \34857 , \34858 , \34859 , \34860 ,
         \34861 , \34862 , \34863 , \34864 , \34865 , \34866 , \34867 , \34868 , \34869 , \34870 ,
         \34871 , \34872 , \34873 , \34874 , \34875 , \34876 , \34877 , \34878 , \34879 , \34880 ,
         \34881 , \34882 , \34883 , \34884 , \34885 , \34886 , \34887 , \34888 , \34889 , \34890 ,
         \34891 , \34892 , \34893 , \34894 , \34895 , \34896 , \34897 , \34898 , \34899 , \34900 ,
         \34901 , \34902 , \34903 , \34904 , \34905 , \34906 , \34907 , \34908 , \34909 , \34910 ,
         \34911 , \34912 , \34913 , \34914 , \34915 , \34916 , \34917 , \34918 , \34919 , \34920 ,
         \34921 , \34922 , \34923 , \34924 , \34925 , \34926 , \34927 , \34928 , \34929 , \34930 ,
         \34931 , \34932 , \34933 , \34934 , \34935 , \34936 , \34937 , \34938 , \34939 , \34940 ,
         \34941 , \34942 , \34943 , \34944 , \34945 , \34946 , \34947 , \34948 , \34949 , \34950 ,
         \34951 , \34952 , \34953 , \34954 , \34955 , \34956 , \34957 , \34958 , \34959 , \34960 ,
         \34961 , \34962 , \34963 , \34964 , \34965 , \34966 , \34967 , \34968 , \34969 , \34970 ,
         \34971 , \34972 , \34973 , \34974 , \34975 , \34976 , \34977 , \34978 , \34979 , \34980 ,
         \34981 , \34982 , \34983 , \34984 , \34985 , \34986 , \34987 , \34988 , \34989 , \34990 ,
         \34991 , \34992 , \34993 , \34994 , \34995 , \34996 , \34997 , \34998 , \34999 , \35000 ,
         \35001 , \35002 , \35003 , \35004 , \35005 , \35006 , \35007 , \35008 , \35009 , \35010 ,
         \35011 , \35012 , \35013 , \35014 , \35015 , \35016 , \35017 , \35018 , \35019 , \35020 ,
         \35021 , \35022 , \35023 , \35024 , \35025 , \35026 , \35027 , \35028 , \35029 , \35030 ,
         \35031 , \35032 , \35033 , \35034 , \35035 , \35036 , \35037 , \35038 , \35039 , \35040 ,
         \35041 , \35042 , \35043 , \35044 , \35045 , \35046 , \35047 , \35048 , \35049 , \35050 ,
         \35051 , \35052 , \35053 , \35054 , \35055 , \35056 , \35057 , \35058 , \35059 , \35060 ,
         \35061 , \35062 , \35063 , \35064 , \35065 , \35066 , \35067 , \35068 , \35069 , \35070 ,
         \35071 , \35072 , \35073 , \35074 , \35075 , \35076 , \35077 , \35078 , \35079 , \35080 ,
         \35081 , \35082 , \35083 , \35084 , \35085 , \35086 , \35087 , \35088 , \35089 , \35090 ,
         \35091 , \35092 , \35093 , \35094 , \35095 , \35096 , \35097 , \35098 , \35099 , \35100 ,
         \35101 , \35102 , \35103 , \35104 , \35105 , \35106 , \35107 , \35108 , \35109 , \35110 ,
         \35111 , \35112 , \35113 , \35114 , \35115 , \35116 , \35117 , \35118 , \35119 , \35120 ,
         \35121 , \35122 , \35123 , \35124 , \35125 , \35126 , \35127 , \35128 , \35129 , \35130 ,
         \35131 , \35132 , \35133 , \35134 , \35135 , \35136 , \35137 , \35138 , \35139 , \35140 ,
         \35141 , \35142 , \35143 , \35144 , \35145 , \35146 , \35147 , \35148 , \35149 , \35150 ,
         \35151 , \35152 , \35153 , \35154 , \35155 , \35156 , \35157 , \35158 , \35159 , \35160 ,
         \35161 , \35162 , \35163 , \35164 , \35165 , \35166 , \35167 , \35168 , \35169 , \35170 ,
         \35171 , \35172 , \35173 , \35174 , \35175 , \35176 , \35177 , \35178 , \35179 , \35180 ,
         \35181 , \35182 , \35183 , \35184 , \35185 , \35186 , \35187 , \35188 , \35189 , \35190 ,
         \35191 , \35192 , \35193 , \35194 , \35195 , \35196 , \35197 , \35198 , \35199 , \35200 ,
         \35201 , \35202 , \35203 , \35204 , \35205 , \35206 , \35207 , \35208 , \35209 , \35210 ,
         \35211 , \35212 , \35213 , \35214 , \35215 , \35216 , \35217 , \35218 , \35219 , \35220 ,
         \35221 , \35222 , \35223 , \35224 , \35225 , \35226 , \35227 , \35228 , \35229 , \35230 ,
         \35231 , \35232 , \35233 , \35234 , \35235 , \35236 , \35237 , \35238 , \35239 , \35240 ,
         \35241 , \35242 , \35243 , \35244 , \35245 , \35246 , \35247 , \35248 , \35249 , \35250 ,
         \35251 , \35252 , \35253 , \35254 , \35255 , \35256 , \35257 , \35258 , \35259 , \35260 ,
         \35261 , \35262 , \35263 , \35264 , \35265 , \35266 , \35267 , \35268 , \35269 , \35270 ,
         \35271 , \35272 , \35273 , \35274 , \35275 , \35276 , \35277 , \35278 , \35279 , \35280 ,
         \35281 , \35282 , \35283 , \35284 , \35285 , \35286 , \35287 , \35288 , \35289 , \35290 ,
         \35291 , \35292 , \35293 , \35294 , \35295 , \35296 , \35297 , \35298 , \35299 , \35300 ,
         \35301 , \35302 , \35303 , \35304 , \35305 , \35306 , \35307 , \35308 , \35309 , \35310 ,
         \35311 , \35312 , \35313 , \35314 , \35315 , \35316 , \35317 , \35318 , \35319 , \35320 ,
         \35321 , \35322 , \35323 , \35324 , \35325 , \35326 , \35327 , \35328 , \35329 , \35330 ,
         \35331 , \35332 , \35333 , \35334 , \35335 , \35336 , \35337 , \35338 , \35339 , \35340 ,
         \35341 , \35342 , \35343 , \35344 , \35345 , \35346 , \35347 , \35348 , \35349 , \35350 ,
         \35351 , \35352 , \35353 , \35354 , \35355 , \35356 , \35357 , \35358 , \35359 , \35360 ,
         \35361 , \35362 , \35363 , \35364 , \35365 , \35366 , \35367 , \35368 , \35369 , \35370 ,
         \35371 , \35372 , \35373 , \35374 , \35375 , \35376 , \35377 , \35378 , \35379 , \35380 ,
         \35381 , \35382 , \35383 , \35384 , \35385 , \35386 , \35387 , \35388 , \35389 , \35390 ,
         \35391 , \35392 , \35393 , \35394 , \35395 , \35396 , \35397 , \35398 , \35399 , \35400 ,
         \35401 , \35402 , \35403 , \35404 , \35405 , \35406 , \35407 , \35408 , \35409 , \35410 ,
         \35411 , \35412 , \35413 , \35414 , \35415 , \35416 , \35417 , \35418 , \35419 , \35420 ,
         \35421 , \35422 , \35423 , \35424 , \35425 , \35426 , \35427 , \35428 , \35429 , \35430 ,
         \35431 , \35432 , \35433 , \35434 , \35435 , \35436 , \35437 , \35438 , \35439 , \35440 ,
         \35441 , \35442 , \35443 , \35444 , \35445 , \35446 , \35447 , \35448 , \35449 , \35450 ,
         \35451 , \35452 , \35453 , \35454 , \35455 , \35456 , \35457 , \35458 , \35459 , \35460 ,
         \35461 , \35462 , \35463 , \35464 , \35465 , \35466 , \35467 , \35468 , \35469 , \35470 ,
         \35471 , \35472 , \35473 , \35474 , \35475 , \35476 , \35477 , \35478 , \35479 , \35480 ,
         \35481 , \35482 , \35483 , \35484 , \35485 , \35486 , \35487 , \35488 , \35489 , \35490 ,
         \35491 , \35492 , \35493 , \35494 , \35495 , \35496 , \35497 , \35498 , \35499 , \35500 ,
         \35501 , \35502 , \35503 , \35504 , \35505 , \35506 , \35507 , \35508 , \35509 , \35510 ,
         \35511 , \35512 , \35513 , \35514 , \35515 , \35516 , \35517 , \35518 , \35519 , \35520 ,
         \35521 , \35522 , \35523 , \35524 , \35525 , \35526 , \35527 , \35528 , \35529 , \35530 ,
         \35531 , \35532 , \35533 , \35534 , \35535 , \35536 , \35537 , \35538 , \35539 , \35540 ,
         \35541 , \35542 , \35543 , \35544 , \35545 , \35546 , \35547 , \35548 , \35549 , \35550 ,
         \35551 , \35552 , \35553 , \35554 , \35555 , \35556 , \35557 , \35558 , \35559 , \35560 ,
         \35561 , \35562 , \35563 , \35564 , \35565 , \35566 , \35567 , \35568 , \35569 , \35570 ,
         \35571 , \35572 , \35573 , \35574 , \35575 , \35576 , \35577 , \35578 , \35579 , \35580 ,
         \35581 , \35582 , \35583 , \35584 , \35585 , \35586 , \35587 , \35588 , \35589 , \35590 ,
         \35591 , \35592 , \35593 , \35594 , \35595 , \35596 , \35597 , \35598 , \35599 , \35600 ,
         \35601 , \35602 , \35603 , \35604 , \35605 , \35606 , \35607 , \35608 , \35609 , \35610 ,
         \35611 , \35612 , \35613 , \35614 , \35615 , \35616 , \35617 , \35618 , \35619 , \35620 ,
         \35621 , \35622 , \35623 , \35624 , \35625 , \35626 , \35627 , \35628 , \35629 , \35630 ,
         \35631 , \35632 , \35633 , \35634 , \35635 , \35636 , \35637 , \35638 , \35639 , \35640 ,
         \35641 , \35642 , \35643 , \35644 , \35645 , \35646 , \35647 , \35648 , \35649 , \35650 ,
         \35651 , \35652 , \35653 , \35654 , \35655 , \35656 , \35657 , \35658 , \35659 , \35660 ,
         \35661 , \35662 , \35663 , \35664 , \35665 , \35666 , \35667 , \35668 , \35669 , \35670 ,
         \35671 , \35672 , \35673 , \35674 , \35675 , \35676 , \35677 , \35678 , \35679 , \35680 ,
         \35681 , \35682 , \35683 , \35684 , \35685 , \35686 , \35687 , \35688 , \35689 , \35690 ,
         \35691 , \35692 , \35693 , \35694 , \35695 , \35696 , \35697 , \35698 , \35699 , \35700 ,
         \35701 , \35702 , \35703 , \35704 , \35705 , \35706 , \35707 , \35708 , \35709 , \35710 ,
         \35711 , \35712 , \35713 , \35714 , \35715 , \35716 , \35717 , \35718 , \35719 , \35720 ,
         \35721 , \35722 , \35723 , \35724 , \35725 , \35726 , \35727 , \35728 , \35729 , \35730 ,
         \35731 , \35732 , \35733 , \35734 , \35735 , \35736 , \35737 , \35738 , \35739 , \35740 ,
         \35741 , \35742 , \35743 , \35744 , \35745 , \35746 , \35747 , \35748 , \35749 , \35750 ,
         \35751 , \35752 , \35753 , \35754 , \35755 , \35756 , \35757 , \35758 , \35759 , \35760 ,
         \35761 , \35762 , \35763 , \35764 , \35765 , \35766 , \35767 , \35768 , \35769 , \35770 ,
         \35771 , \35772 , \35773 , \35774 , \35775 , \35776 , \35777 , \35778 , \35779 , \35780 ,
         \35781 , \35782 , \35783 , \35784 , \35785 , \35786 , \35787 , \35788 , \35789 , \35790 ,
         \35791 , \35792 , \35793 , \35794 , \35795 , \35796 , \35797 , \35798 , \35799 , \35800 ,
         \35801 , \35802 , \35803 , \35804 , \35805 , \35806 , \35807 , \35808 , \35809 , \35810 ,
         \35811 , \35812 , \35813 , \35814 , \35815 , \35816 , \35817 , \35818 , \35819 , \35820 ,
         \35821 , \35822 , \35823 , \35824 , \35825 , \35826 , \35827 , \35828 , \35829 , \35830 ,
         \35831 , \35832 , \35833 , \35834 , \35835 , \35836 , \35837 , \35838 , \35839 , \35840 ,
         \35841 , \35842 , \35843 , \35844 , \35845 , \35846 , \35847 , \35848 , \35849 , \35850 ,
         \35851 , \35852 , \35853 , \35854 , \35855 , \35856 , \35857 , \35858 , \35859 , \35860 ,
         \35861 , \35862 , \35863 , \35864 , \35865 , \35866 , \35867 , \35868 , \35869 , \35870 ,
         \35871 , \35872 , \35873 , \35874 , \35875 , \35876 , \35877 , \35878 , \35879 , \35880 ,
         \35881 , \35882 , \35883 , \35884 , \35885 , \35886 , \35887 , \35888 , \35889 , \35890 ,
         \35891 , \35892 , \35893 , \35894 , \35895 , \35896 , \35897 , \35898 , \35899 , \35900 ,
         \35901 , \35902 , \35903 , \35904 , \35905 , \35906 , \35907 , \35908 , \35909 , \35910 ,
         \35911 , \35912 , \35913 , \35914 , \35915 , \35916 , \35917 , \35918 , \35919 , \35920 ,
         \35921 , \35922 , \35923 , \35924 , \35925 , \35926 , \35927 , \35928 , \35929 , \35930 ,
         \35931 , \35932 , \35933 , \35934 , \35935 , \35936 , \35937 , \35938 , \35939 , \35940 ,
         \35941 , \35942 , \35943 , \35944 , \35945 , \35946 , \35947 , \35948 , \35949 , \35950 ,
         \35951 , \35952 , \35953 , \35954 , \35955 , \35956 , \35957 , \35958 , \35959 , \35960 ,
         \35961 , \35962 , \35963 , \35964 , \35965 , \35966 , \35967 , \35968 , \35969 , \35970 ,
         \35971 , \35972 , \35973 , \35974 , \35975 , \35976 , \35977 , \35978 , \35979 , \35980 ,
         \35981 , \35982 , \35983 , \35984 , \35985 , \35986 , \35987 , \35988 , \35989 , \35990 ,
         \35991 , \35992 , \35993 , \35994 , \35995 , \35996 , \35997 , \35998 , \35999 , \36000 ,
         \36001 , \36002 , \36003 , \36004 , \36005 , \36006 , \36007 , \36008 , \36009 , \36010 ,
         \36011 , \36012 , \36013 , \36014 , \36015 , \36016 , \36017 , \36018 , \36019 , \36020 ,
         \36021 , \36022 , \36023 , \36024 , \36025 , \36026 , \36027 , \36028 , \36029 , \36030 ,
         \36031 , \36032 , \36033 , \36034 , \36035 , \36036 , \36037 , \36038 , \36039 , \36040 ,
         \36041 , \36042 , \36043 , \36044 , \36045 , \36046 , \36047 , \36048 , \36049 , \36050 ,
         \36051 , \36052 , \36053 , \36054 , \36055 , \36056 , \36057 , \36058 , \36059 , \36060 ,
         \36061 , \36062 , \36063 , \36064 , \36065 , \36066 , \36067 , \36068 , \36069 , \36070 ,
         \36071 , \36072 , \36073 , \36074 , \36075 , \36076 , \36077 , \36078 , \36079 , \36080 ,
         \36081 , \36082 , \36083 , \36084 , \36085 , \36086 , \36087 , \36088 , \36089 , \36090 ,
         \36091 , \36092 , \36093 , \36094 , \36095 , \36096 , \36097 , \36098 , \36099 , \36100 ,
         \36101 , \36102 , \36103 , \36104 , \36105 , \36106 , \36107 , \36108 , \36109 , \36110 ,
         \36111 , \36112 , \36113 , \36114 , \36115 , \36116 , \36117 , \36118 , \36119 , \36120 ,
         \36121 , \36122 , \36123 , \36124 , \36125 , \36126 , \36127 , \36128 , \36129 , \36130 ,
         \36131 , \36132 , \36133 , \36134 , \36135 , \36136 , \36137 , \36138 , \36139 , \36140 ,
         \36141 , \36142 , \36143 , \36144 , \36145 , \36146 , \36147 , \36148 , \36149 , \36150 ,
         \36151 , \36152 , \36153 , \36154 , \36155 , \36156 , \36157 , \36158 , \36159 , \36160 ,
         \36161 , \36162 , \36163 , \36164 , \36165 , \36166 , \36167 , \36168 , \36169 , \36170 ,
         \36171 , \36172 , \36173 , \36174 , \36175 , \36176 , \36177 , \36178 , \36179 , \36180 ,
         \36181 , \36182 , \36183 , \36184 , \36185 , \36186 , \36187 , \36188 , \36189 , \36190 ,
         \36191 , \36192 , \36193 , \36194 , \36195 , \36196 , \36197 , \36198 , \36199 , \36200 ,
         \36201 , \36202 , \36203 , \36204 , \36205 , \36206 , \36207 , \36208 , \36209 , \36210 ,
         \36211 , \36212 , \36213 , \36214 , \36215 , \36216 , \36217 , \36218 , \36219 , \36220 ,
         \36221 , \36222 , \36223 , \36224 , \36225 , \36226 , \36227 , \36228 , \36229 , \36230 ,
         \36231 , \36232 , \36233 , \36234 , \36235 , \36236 , \36237 , \36238 , \36239 , \36240 ,
         \36241 , \36242 , \36243 , \36244 , \36245 , \36246 , \36247 , \36248 , \36249 , \36250 ,
         \36251 , \36252 , \36253 , \36254 , \36255 , \36256 , \36257 , \36258 , \36259 , \36260 ,
         \36261 , \36262 , \36263 , \36264 , \36265 , \36266 , \36267 , \36268 , \36269 , \36270 ,
         \36271 , \36272 , \36273 , \36274 , \36275 , \36276 , \36277 , \36278 , \36279 , \36280 ,
         \36281 , \36282 , \36283 , \36284 , \36285 , \36286 , \36287 , \36288 , \36289 , \36290 ,
         \36291 , \36292 , \36293 , \36294 , \36295 , \36296 , \36297 , \36298 , \36299 , \36300 ,
         \36301 , \36302 , \36303 , \36304 , \36305 , \36306 , \36307 , \36308 , \36309 , \36310 ,
         \36311 , \36312 , \36313 , \36314 , \36315 , \36316 , \36317 , \36318 , \36319 , \36320 ,
         \36321 , \36322 , \36323 , \36324 , \36325 , \36326 , \36327 , \36328 , \36329 , \36330 ,
         \36331 , \36332 , \36333 , \36334 , \36335 , \36336 , \36337 , \36338 , \36339 , \36340 ,
         \36341 , \36342 , \36343 , \36344 , \36345 , \36346 , \36347 , \36348 , \36349 , \36350 ,
         \36351 , \36352 , \36353 , \36354 , \36355 , \36356 , \36357 , \36358 , \36359 , \36360 ,
         \36361 , \36362 , \36363 , \36364 , \36365 , \36366 , \36367 , \36368 , \36369 , \36370 ,
         \36371 , \36372 , \36373 , \36374 , \36375 , \36376 , \36377 , \36378 , \36379 , \36380 ,
         \36381 , \36382 , \36383 , \36384 , \36385 , \36386 , \36387 , \36388 , \36389 , \36390 ,
         \36391 , \36392 , \36393 , \36394 , \36395 , \36396 , \36397 , \36398 , \36399 , \36400 ,
         \36401 , \36402 , \36403 , \36404 , \36405 , \36406 , \36407 , \36408 , \36409 , \36410 ,
         \36411 , \36412 , \36413 , \36414 , \36415 , \36416 , \36417 , \36418 , \36419 , \36420 ,
         \36421 , \36422 , \36423 , \36424 , \36425 , \36426 , \36427 , \36428 , \36429 , \36430 ,
         \36431 , \36432 , \36433 , \36434 , \36435 , \36436 , \36437 , \36438 , \36439 , \36440 ,
         \36441 , \36442 , \36443 , \36444 , \36445 , \36446 , \36447 , \36448 , \36449 , \36450 ,
         \36451 , \36452 , \36453 , \36454 , \36455 , \36456 , \36457 , \36458 , \36459 , \36460 ,
         \36461 , \36462 , \36463 , \36464 , \36465 , \36466 , \36467 , \36468 , \36469 , \36470 ,
         \36471 , \36472 , \36473 , \36474 , \36475 , \36476 , \36477 , \36478 , \36479 , \36480 ,
         \36481 , \36482 , \36483 , \36484 , \36485 , \36486 , \36487 , \36488 , \36489 , \36490 ,
         \36491 , \36492 , \36493 , \36494 , \36495 , \36496 , \36497 , \36498 , \36499 , \36500 ,
         \36501 , \36502 , \36503 , \36504 , \36505 , \36506 , \36507 , \36508 , \36509 , \36510 ,
         \36511 , \36512 , \36513 , \36514 , \36515 , \36516 , \36517 , \36518 , \36519 , \36520 ,
         \36521 , \36522 , \36523 , \36524 , \36525 , \36526 , \36527 , \36528 , \36529 , \36530 ,
         \36531 , \36532 , \36533 , \36534 , \36535 , \36536 , \36537 , \36538 , \36539 , \36540 ,
         \36541 , \36542 , \36543 , \36544 , \36545 , \36546 , \36547 , \36548 , \36549 , \36550 ,
         \36551 , \36552 , \36553 , \36554 , \36555 , \36556 , \36557 , \36558 , \36559 , \36560 ,
         \36561 , \36562 , \36563 , \36564 , \36565 , \36566 , \36567 , \36568 , \36569 , \36570 ,
         \36571 , \36572 , \36573 , \36574 , \36575 , \36576 , \36577 , \36578 , \36579 , \36580 ,
         \36581 , \36582 , \36583 , \36584 , \36585 , \36586 , \36587 , \36588 , \36589 , \36590 ,
         \36591 , \36592 , \36593 , \36594 , \36595 , \36596 , \36597 , \36598 , \36599 , \36600 ,
         \36601 , \36602 , \36603 , \36604 , \36605 , \36606 , \36607 , \36608 , \36609 , \36610 ,
         \36611 , \36612 , \36613 , \36614 , \36615 , \36616 , \36617 , \36618 , \36619 , \36620 ,
         \36621 , \36622 , \36623 , \36624 , \36625 , \36626 , \36627 , \36628 , \36629 , \36630 ,
         \36631 , \36632 , \36633 , \36634 , \36635 , \36636 , \36637 , \36638 , \36639 , \36640 ,
         \36641 , \36642 , \36643 , \36644 , \36645 , \36646 , \36647 , \36648 , \36649 , \36650 ,
         \36651 , \36652 , \36653 , \36654 , \36655 , \36656 , \36657 , \36658 , \36659 , \36660 ,
         \36661 , \36662 , \36663 , \36664 , \36665 , \36666 , \36667 , \36668 , \36669 , \36670 ,
         \36671 , \36672 , \36673 , \36674 , \36675 , \36676 , \36677 , \36678 , \36679 , \36680 ,
         \36681 , \36682 , \36683 , \36684 , \36685 , \36686 , \36687 , \36688 , \36689 , \36690 ,
         \36691 , \36692 , \36693 , \36694 , \36695 , \36696 , \36697 , \36698 , \36699 , \36700 ,
         \36701 , \36702 , \36703 , \36704 , \36705 , \36706 , \36707 , \36708 , \36709 , \36710 ,
         \36711 , \36712 , \36713 , \36714 , \36715 , \36716 , \36717 , \36718 , \36719 , \36720 ,
         \36721 , \36722 , \36723 , \36724 , \36725 , \36726 , \36727 , \36728 , \36729 , \36730 ,
         \36731 , \36732 , \36733 , \36734 , \36735 , \36736 , \36737 , \36738 , \36739 , \36740 ,
         \36741 , \36742 , \36743 , \36744 , \36745 , \36746 , \36747 , \36748 , \36749 , \36750 ,
         \36751 , \36752 , \36753 , \36754 , \36755 , \36756 , \36757 , \36758 , \36759 , \36760 ,
         \36761 , \36762 , \36763 , \36764 , \36765 , \36766 , \36767 , \36768 , \36769 , \36770 ,
         \36771 , \36772 , \36773 , \36774 , \36775 , \36776 , \36777 , \36778 , \36779 , \36780 ,
         \36781 , \36782 , \36783 , \36784 , \36785 , \36786 , \36787 , \36788 , \36789 , \36790 ,
         \36791 , \36792 , \36793 , \36794 , \36795 , \36796 , \36797 , \36798 , \36799 , \36800 ,
         \36801 , \36802 , \36803 , \36804 , \36805 , \36806 , \36807 , \36808 , \36809 , \36810 ,
         \36811 , \36812 , \36813 , \36814 , \36815 , \36816 , \36817 , \36818 , \36819 , \36820 ,
         \36821 , \36822 , \36823 , \36824 , \36825 , \36826 , \36827 , \36828 , \36829 , \36830 ,
         \36831 , \36832 , \36833 , \36834 , \36835 , \36836 , \36837 , \36838 , \36839 , \36840 ,
         \36841 , \36842 , \36843 , \36844 , \36845 , \36846 , \36847 , \36848 , \36849 , \36850 ,
         \36851 , \36852 , \36853 , \36854 , \36855 , \36856 , \36857 , \36858 , \36859 , \36860 ,
         \36861 , \36862 , \36863 , \36864 , \36865 , \36866 , \36867 , \36868 , \36869 , \36870 ,
         \36871 , \36872 , \36873 , \36874 , \36875 , \36876 , \36877 , \36878 , \36879 , \36880 ,
         \36881 , \36882 , \36883 , \36884 , \36885 , \36886 , \36887 , \36888 , \36889 , \36890 ,
         \36891 , \36892 , \36893 , \36894 , \36895 , \36896 , \36897 , \36898 , \36899 , \36900 ,
         \36901 , \36902 , \36903 , \36904 , \36905 , \36906 , \36907 , \36908 , \36909 , \36910 ,
         \36911 , \36912 , \36913 , \36914 , \36915 , \36916 , \36917 , \36918 , \36919 , \36920 ,
         \36921 , \36922 , \36923 , \36924 , \36925 , \36926 , \36927 , \36928 , \36929 , \36930 ,
         \36931 , \36932 , \36933 , \36934 , \36935 , \36936 , \36937 , \36938 , \36939 , \36940 ,
         \36941 , \36942 , \36943 , \36944 , \36945 , \36946 , \36947 , \36948 , \36949 , \36950 ,
         \36951 , \36952 , \36953 , \36954 , \36955 , \36956 , \36957 , \36958 , \36959 , \36960 ,
         \36961 , \36962 , \36963 , \36964 , \36965 , \36966 , \36967 , \36968 , \36969 , \36970 ,
         \36971 , \36972 , \36973 , \36974 , \36975 , \36976 , \36977 , \36978 , \36979 , \36980 ,
         \36981 , \36982 , \36983 , \36984 , \36985 , \36986 , \36987 , \36988 , \36989 , \36990 ,
         \36991 , \36992 , \36993 , \36994 , \36995 , \36996 , \36997 , \36998 , \36999 , \37000 ,
         \37001 , \37002 , \37003 , \37004 , \37005 , \37006 , \37007 , \37008 , \37009 , \37010 ,
         \37011 , \37012 , \37013 , \37014 , \37015 , \37016 , \37017 , \37018 , \37019 , \37020 ,
         \37021 , \37022 , \37023 , \37024 , \37025 , \37026 , \37027 , \37028 , \37029 , \37030 ,
         \37031 , \37032 , \37033 , \37034 , \37035 , \37036 , \37037 , \37038 , \37039 , \37040 ,
         \37041 , \37042 , \37043 , \37044 , \37045 , \37046 , \37047 , \37048 , \37049 , \37050 ,
         \37051 , \37052 , \37053 , \37054 , \37055 , \37056 , \37057 , \37058 , \37059 , \37060 ,
         \37061 , \37062 , \37063 , \37064 , \37065 , \37066 , \37067 , \37068 , \37069 , \37070 ,
         \37071 , \37072 , \37073 , \37074 , \37075 , \37076 , \37077 , \37078 , \37079 , \37080 ,
         \37081 , \37082 , \37083 , \37084 , \37085 , \37086 , \37087 , \37088 , \37089 , \37090 ,
         \37091 , \37092 , \37093 , \37094 , \37095 , \37096 , \37097 , \37098 , \37099 , \37100 ,
         \37101 , \37102 , \37103 , \37104 , \37105 , \37106 , \37107 , \37108 , \37109 , \37110 ,
         \37111 , \37112 , \37113 , \37114 , \37115 , \37116 , \37117 , \37118 , \37119 , \37120 ,
         \37121 , \37122 , \37123 , \37124 , \37125 , \37126 , \37127 , \37128 , \37129 , \37130 ,
         \37131 , \37132 , \37133 , \37134 , \37135 , \37136 , \37137 , \37138 , \37139 , \37140 ,
         \37141 , \37142 , \37143 , \37144 , \37145 , \37146 , \37147 , \37148 , \37149 , \37150 ,
         \37151 , \37152 , \37153 , \37154 , \37155 , \37156 , \37157 , \37158 , \37159 , \37160 ,
         \37161 , \37162 , \37163 , \37164 , \37165 , \37166 , \37167 , \37168 , \37169 , \37170 ,
         \37171 , \37172 , \37173 , \37174 , \37175 , \37176 , \37177 , \37178 , \37179 , \37180 ,
         \37181 , \37182 , \37183 , \37184 , \37185 , \37186 , \37187 , \37188 , \37189 , \37190 ,
         \37191 , \37192 , \37193 , \37194 , \37195 , \37196 , \37197 , \37198 , \37199 , \37200 ,
         \37201 , \37202 , \37203 , \37204 , \37205 , \37206 , \37207 , \37208 , \37209 , \37210 ,
         \37211 , \37212 , \37213 , \37214 , \37215 , \37216 , \37217 , \37218 , \37219 , \37220 ,
         \37221 , \37222 , \37223 , \37224 , \37225 , \37226 , \37227 , \37228 , \37229 , \37230 ,
         \37231 , \37232 , \37233 , \37234 , \37235 , \37236 , \37237 , \37238 , \37239 , \37240 ,
         \37241 , \37242 , \37243 , \37244 , \37245 , \37246 , \37247 , \37248 , \37249 , \37250 ,
         \37251 , \37252 , \37253 , \37254 , \37255 , \37256 , \37257 , \37258 , \37259 , \37260 ,
         \37261 , \37262 , \37263 , \37264 , \37265 , \37266 , \37267 , \37268 , \37269 , \37270 ,
         \37271 , \37272 , \37273 , \37274 , \37275 , \37276 , \37277 , \37278 , \37279 , \37280 ,
         \37281 , \37282 , \37283 , \37284 , \37285 , \37286 , \37287 , \37288 , \37289 , \37290 ,
         \37291 , \37292 , \37293 , \37294 , \37295 , \37296 , \37297 , \37298 , \37299 , \37300 ,
         \37301 , \37302 , \37303 , \37304 , \37305 , \37306 , \37307 , \37308 , \37309 , \37310 ,
         \37311 , \37312 , \37313 , \37314 , \37315 , \37316 , \37317 , \37318 , \37319 , \37320 ,
         \37321 , \37322 , \37323 , \37324 , \37325 , \37326 , \37327 , \37328 , \37329 , \37330 ,
         \37331 , \37332 , \37333 , \37334 , \37335 , \37336 , \37337 , \37338 , \37339 , \37340 ,
         \37341 , \37342 , \37343 , \37344 , \37345 , \37346 , \37347 , \37348 , \37349 , \37350 ,
         \37351 , \37352 , \37353 , \37354 , \37355 , \37356 , \37357 , \37358 , \37359 , \37360 ,
         \37361 , \37362 , \37363 , \37364 , \37365 , \37366 , \37367 , \37368 , \37369 , \37370 ,
         \37371 , \37372 , \37373 , \37374 , \37375 , \37376 , \37377 , \37378 , \37379 , \37380 ,
         \37381 , \37382 , \37383 , \37384 , \37385 , \37386 , \37387 , \37388 , \37389 , \37390 ,
         \37391 , \37392 , \37393 , \37394 , \37395 , \37396 , \37397 , \37398 , \37399 , \37400 ,
         \37401 , \37402 , \37403 , \37404 , \37405 , \37406 , \37407 , \37408 , \37409 , \37410 ,
         \37411 , \37412 , \37413 , \37414 , \37415 , \37416 , \37417 , \37418 , \37419 , \37420 ,
         \37421 , \37422 , \37423 , \37424 , \37425 , \37426 , \37427 , \37428 , \37429 , \37430 ,
         \37431 , \37432 , \37433 , \37434 , \37435 , \37436 , \37437 , \37438 , \37439 , \37440 ,
         \37441 , \37442 , \37443 , \37444 , \37445 , \37446 , \37447 , \37448 , \37449 , \37450 ,
         \37451 , \37452 , \37453 , \37454 , \37455 , \37456 , \37457 , \37458 , \37459 , \37460 ,
         \37461 , \37462 , \37463 , \37464 , \37465 , \37466 , \37467 , \37468 , \37469 , \37470 ,
         \37471 , \37472 , \37473 , \37474 , \37475 , \37476 , \37477 , \37478 , \37479 , \37480 ,
         \37481 , \37482 , \37483 , \37484 , \37485 , \37486 , \37487 , \37488 , \37489 , \37490 ,
         \37491 , \37492 , \37493 , \37494 , \37495 , \37496 , \37497 , \37498 , \37499 , \37500 ,
         \37501 , \37502 , \37503 , \37504 , \37505 , \37506 , \37507 , \37508 , \37509 , \37510 ,
         \37511 , \37512 , \37513 , \37514 , \37515 , \37516 , \37517 , \37518 , \37519 , \37520 ,
         \37521 , \37522 , \37523 , \37524 , \37525 , \37526 , \37527 , \37528 , \37529 , \37530 ,
         \37531 , \37532 , \37533 , \37534 , \37535 , \37536 , \37537 , \37538 , \37539 , \37540 ,
         \37541 , \37542 , \37543 , \37544 , \37545 , \37546 , \37547 , \37548 , \37549 , \37550 ,
         \37551 , \37552 , \37553 , \37554 , \37555 , \37556 , \37557 , \37558 , \37559 , \37560 ,
         \37561 , \37562 , \37563 , \37564 , \37565 , \37566 , \37567 , \37568 , \37569 , \37570 ,
         \37571 , \37572 , \37573 , \37574 , \37575 , \37576 , \37577 , \37578 , \37579 , \37580 ,
         \37581 , \37582 , \37583 , \37584 , \37585 , \37586 , \37587 , \37588 , \37589 , \37590 ,
         \37591 , \37592 , \37593 , \37594 , \37595 , \37596 , \37597 , \37598 , \37599 , \37600 ,
         \37601 , \37602 , \37603 , \37604 , \37605 , \37606 , \37607 , \37608 , \37609 , \37610 ,
         \37611 , \37612 , \37613 , \37614 , \37615 , \37616 , \37617 , \37618 , \37619 , \37620 ,
         \37621 , \37622 , \37623 , \37624 , \37625 , \37626 , \37627 , \37628 , \37629 , \37630 ,
         \37631 , \37632 , \37633 , \37634 , \37635 , \37636 , \37637 , \37638 , \37639 , \37640 ,
         \37641 , \37642 , \37643 , \37644 , \37645 , \37646 , \37647 , \37648 , \37649 , \37650 ,
         \37651 , \37652 , \37653 , \37654 , \37655 , \37656 , \37657 , \37658 , \37659 , \37660 ,
         \37661 , \37662 , \37663 , \37664 , \37665 , \37666 , \37667 , \37668 , \37669 , \37670 ,
         \37671 , \37672 , \37673 , \37674 , \37675 , \37676 , \37677 , \37678 , \37679 , \37680 ,
         \37681 , \37682 , \37683 , \37684 , \37685 , \37686 , \37687 , \37688 , \37689 , \37690 ,
         \37691 , \37692 , \37693 , \37694 , \37695 , \37696 , \37697 , \37698 , \37699 , \37700 ,
         \37701 , \37702 , \37703 , \37704 , \37705 , \37706 , \37707 , \37708 , \37709 , \37710 ,
         \37711 , \37712 , \37713 , \37714 , \37715 , \37716 , \37717 , \37718 , \37719 , \37720 ,
         \37721 , \37722 , \37723 , \37724 , \37725 , \37726 , \37727 , \37728 , \37729 , \37730 ,
         \37731 , \37732 , \37733 , \37734 , \37735 , \37736 , \37737 , \37738 , \37739 , \37740 ,
         \37741 , \37742 , \37743 , \37744 , \37745 , \37746 , \37747 , \37748 , \37749 , \37750 ,
         \37751 , \37752 , \37753 , \37754 , \37755 , \37756 , \37757 , \37758 , \37759 , \37760 ,
         \37761 , \37762 , \37763 , \37764 , \37765 , \37766 , \37767 , \37768 , \37769 , \37770 ,
         \37771 , \37772 , \37773 , \37774 , \37775 , \37776 , \37777 , \37778 , \37779 , \37780 ,
         \37781 , \37782 , \37783 , \37784 , \37785 , \37786 , \37787 , \37788 , \37789 , \37790 ,
         \37791 , \37792 , \37793 , \37794 , \37795 , \37796 , \37797 , \37798 , \37799 , \37800 ,
         \37801 , \37802 , \37803 , \37804 , \37805 , \37806 , \37807 , \37808 , \37809 , \37810 ,
         \37811 , \37812 , \37813 , \37814 , \37815 , \37816 , \37817 , \37818 , \37819 , \37820 ,
         \37821 , \37822 , \37823 , \37824 , \37825 , \37826 , \37827 , \37828 , \37829 , \37830 ,
         \37831 , \37832 , \37833 , \37834 , \37835 , \37836 , \37837 , \37838 , \37839 , \37840 ,
         \37841 , \37842 , \37843 , \37844 , \37845 , \37846 , \37847 , \37848 , \37849 , \37850 ,
         \37851 , \37852 , \37853 , \37854 , \37855 , \37856 , \37857 , \37858 , \37859 , \37860 ,
         \37861 , \37862 , \37863 , \37864 , \37865 , \37866 , \37867 , \37868 , \37869 , \37870 ,
         \37871 , \37872 , \37873 , \37874 , \37875 , \37876 , \37877 , \37878 , \37879 , \37880 ,
         \37881 , \37882 , \37883 , \37884 , \37885 , \37886 , \37887 , \37888 , \37889 , \37890 ,
         \37891 , \37892 , \37893 , \37894 , \37895 , \37896 , \37897 , \37898 , \37899 , \37900 ,
         \37901 , \37902 , \37903 , \37904 , \37905 , \37906 , \37907 , \37908 , \37909 , \37910 ,
         \37911 , \37912 , \37913 , \37914 , \37915 , \37916 , \37917 , \37918 , \37919 , \37920 ,
         \37921 , \37922 , \37923 , \37924 , \37925 , \37926 , \37927 , \37928 , \37929 , \37930 ,
         \37931 , \37932 , \37933 , \37934 , \37935 , \37936 , \37937 , \37938 , \37939 , \37940 ,
         \37941 , \37942 , \37943 , \37944 , \37945 , \37946 , \37947 , \37948 , \37949 , \37950 ,
         \37951 , \37952 , \37953 , \37954 , \37955 , \37956 , \37957 , \37958 , \37959 , \37960 ,
         \37961 , \37962 , \37963 , \37964 , \37965 , \37966 , \37967 , \37968 , \37969 , \37970 ,
         \37971 , \37972 , \37973 , \37974 , \37975 , \37976 , \37977 , \37978 , \37979 , \37980 ,
         \37981 , \37982 , \37983 , \37984 , \37985 , \37986 , \37987 , \37988 , \37989 , \37990 ,
         \37991 , \37992 , \37993 , \37994 , \37995 , \37996 , \37997 , \37998 , \37999 , \38000 ,
         \38001 , \38002 , \38003 , \38004 , \38005 , \38006 , \38007 , \38008 , \38009 , \38010 ,
         \38011 , \38012 , \38013 , \38014 , \38015 , \38016 , \38017 , \38018 , \38019 , \38020 ,
         \38021 , \38022 , \38023 , \38024 , \38025 , \38026 , \38027 , \38028 , \38029 , \38030 ,
         \38031 , \38032 , \38033 , \38034 , \38035 , \38036 , \38037 , \38038 , \38039 , \38040 ,
         \38041 , \38042 , \38043 , \38044 , \38045 , \38046 , \38047 , \38048 , \38049 , \38050 ,
         \38051 , \38052 , \38053 , \38054 , \38055 , \38056 , \38057 , \38058 , \38059 , \38060 ,
         \38061 , \38062 , \38063 , \38064 , \38065 , \38066 , \38067 , \38068 , \38069 , \38070 ,
         \38071 , \38072 , \38073 , \38074 , \38075 , \38076 , \38077 , \38078 , \38079 , \38080 ,
         \38081 , \38082 , \38083 , \38084 , \38085 , \38086 , \38087 , \38088 , \38089 , \38090 ,
         \38091 , \38092 , \38093 , \38094 , \38095 , \38096 , \38097 , \38098 , \38099 , \38100 ,
         \38101 , \38102 , \38103 , \38104 , \38105 , \38106 , \38107 , \38108 , \38109 , \38110 ,
         \38111 , \38112 , \38113 , \38114 , \38115 , \38116 , \38117 , \38118 , \38119 , \38120 ,
         \38121 , \38122 , \38123 , \38124 , \38125 , \38126 , \38127 , \38128 , \38129 , \38130 ,
         \38131 , \38132 , \38133 , \38134 , \38135 , \38136 , \38137 , \38138 , \38139 , \38140 ,
         \38141 , \38142 , \38143 , \38144 , \38145 , \38146 , \38147 , \38148 , \38149 , \38150 ,
         \38151 , \38152 , \38153 , \38154 , \38155 , \38156 , \38157 , \38158 , \38159 , \38160 ,
         \38161 , \38162 , \38163 , \38164 , \38165 , \38166 , \38167 , \38168 , \38169 , \38170 ,
         \38171 , \38172 , \38173 , \38174 , \38175 , \38176 , \38177 , \38178 , \38179 , \38180 ,
         \38181 , \38182 , \38183 , \38184 , \38185 , \38186 , \38187 , \38188 , \38189 , \38190 ,
         \38191 , \38192 , \38193 , \38194 , \38195 , \38196 , \38197 , \38198 , \38199 , \38200 ,
         \38201 , \38202 , \38203 , \38204 , \38205 , \38206 , \38207 , \38208 , \38209 , \38210 ,
         \38211 , \38212 , \38213 , \38214 , \38215 , \38216 , \38217 , \38218 , \38219 , \38220 ,
         \38221 , \38222 , \38223 , \38224 , \38225 , \38226 , \38227 , \38228 , \38229 , \38230 ,
         \38231 , \38232 , \38233 , \38234 , \38235 , \38236 , \38237 , \38238 , \38239 , \38240 ,
         \38241 , \38242 , \38243 , \38244 , \38245 , \38246 , \38247 , \38248 , \38249 , \38250 ,
         \38251 , \38252 , \38253 , \38254 , \38255 , \38256 , \38257 , \38258 , \38259 , \38260 ,
         \38261 , \38262 , \38263 , \38264 , \38265 , \38266 , \38267 , \38268 , \38269 , \38270 ,
         \38271 , \38272 , \38273 , \38274 , \38275 , \38276 , \38277 , \38278 , \38279 , \38280 ,
         \38281 , \38282 , \38283 , \38284 , \38285 , \38286 , \38287 , \38288 , \38289 , \38290 ,
         \38291 , \38292 , \38293 , \38294 , \38295 , \38296 , \38297 , \38298 , \38299 , \38300 ,
         \38301 , \38302 , \38303 , \38304 , \38305 , \38306 , \38307 , \38308 , \38309 , \38310 ,
         \38311 , \38312 , \38313 , \38314 , \38315 , \38316 , \38317 , \38318 , \38319 , \38320 ,
         \38321 , \38322 , \38323 , \38324 , \38325 , \38326 , \38327 , \38328 , \38329 , \38330 ,
         \38331 , \38332 , \38333 , \38334 , \38335 , \38336 , \38337 , \38338 , \38339 , \38340 ,
         \38341 , \38342 , \38343 , \38344 , \38345 , \38346 , \38347 , \38348 , \38349 , \38350 ,
         \38351 , \38352 , \38353 , \38354 , \38355 , \38356 , \38357 , \38358 , \38359 , \38360 ,
         \38361 , \38362 , \38363 , \38364 , \38365 , \38366 , \38367 , \38368 , \38369 , \38370 ,
         \38371 , \38372 , \38373 , \38374 , \38375 , \38376 , \38377 , \38378 , \38379 , \38380 ,
         \38381 , \38382 , \38383 , \38384 , \38385 , \38386 , \38387 , \38388 , \38389 , \38390 ,
         \38391 , \38392 , \38393 , \38394 , \38395 , \38396 , \38397 , \38398 , \38399 , \38400 ,
         \38401 , \38402 , \38403 , \38404 , \38405 , \38406 , \38407 , \38408 , \38409 , \38410 ,
         \38411 , \38412 , \38413 , \38414 , \38415 , \38416 , \38417 , \38418 , \38419 , \38420 ,
         \38421 , \38422 , \38423 , \38424 , \38425 , \38426 , \38427 , \38428 , \38429 , \38430 ,
         \38431 , \38432 , \38433 , \38434 , \38435 , \38436 , \38437 , \38438 , \38439 , \38440 ,
         \38441 , \38442 , \38443 , \38444 , \38445 , \38446 , \38447 , \38448 , \38449 , \38450 ,
         \38451 , \38452 , \38453 , \38454 , \38455 , \38456 , \38457 , \38458 , \38459 , \38460 ,
         \38461 , \38462 , \38463 , \38464 , \38465 , \38466 , \38467 , \38468 , \38469 , \38470 ,
         \38471 , \38472 , \38473 , \38474 , \38475 , \38476 , \38477 , \38478 , \38479 , \38480 ,
         \38481 , \38482 , \38483 , \38484 , \38485 , \38486 , \38487 , \38488 , \38489 , \38490 ,
         \38491 , \38492 , \38493 , \38494 , \38495 , \38496 , \38497 , \38498 , \38499 , \38500 ,
         \38501 , \38502 , \38503 , \38504 , \38505 , \38506 , \38507 , \38508 , \38509 , \38510 ,
         \38511 , \38512 , \38513 , \38514 , \38515 , \38516 , \38517 , \38518 , \38519 , \38520 ,
         \38521 , \38522 , \38523 , \38524 , \38525 , \38526 , \38527 , \38528 , \38529 , \38530 ,
         \38531 , \38532 , \38533 , \38534 , \38535 , \38536 , \38537 , \38538 , \38539 , \38540 ,
         \38541 , \38542 , \38543 , \38544 , \38545 , \38546 , \38547 , \38548 , \38549 , \38550 ,
         \38551 , \38552 , \38553 , \38554 , \38555 , \38556 , \38557 , \38558 , \38559 , \38560 ,
         \38561 , \38562 , \38563 , \38564 , \38565 , \38566 , \38567 , \38568 , \38569 , \38570 ,
         \38571 , \38572 , \38573 , \38574 , \38575 , \38576 , \38577 , \38578 , \38579 , \38580 ,
         \38581 , \38582 , \38583 , \38584 , \38585 , \38586 , \38587 , \38588 , \38589 , \38590 ,
         \38591 , \38592 , \38593 , \38594 , \38595 , \38596 , \38597 , \38598 , \38599 , \38600 ,
         \38601 , \38602 , \38603 , \38604 , \38605 , \38606 , \38607 , \38608 , \38609 , \38610 ,
         \38611 , \38612 , \38613 , \38614 , \38615 , \38616 , \38617 , \38618 , \38619 , \38620 ,
         \38621 , \38622 , \38623 , \38624 , \38625 , \38626 , \38627 , \38628 , \38629 , \38630 ,
         \38631 , \38632 , \38633 , \38634 , \38635 , \38636 , \38637 , \38638 , \38639 , \38640 ,
         \38641 , \38642 , \38643 , \38644 , \38645 , \38646 , \38647 , \38648 , \38649 , \38650 ,
         \38651 , \38652 , \38653 , \38654 , \38655 , \38656 , \38657 , \38658 , \38659 , \38660 ,
         \38661 , \38662 , \38663 , \38664 , \38665 , \38666 , \38667 , \38668 , \38669 , \38670 ,
         \38671 , \38672 , \38673 , \38674 , \38675 , \38676 , \38677 , \38678 , \38679 , \38680 ,
         \38681 , \38682 , \38683 , \38684 , \38685 , \38686 , \38687 , \38688 , \38689 , \38690 ,
         \38691 , \38692 , \38693 , \38694 , \38695 , \38696 , \38697 , \38698 , \38699 , \38700 ,
         \38701 , \38702 , \38703 , \38704 , \38705 , \38706 , \38707 , \38708 , \38709 , \38710 ,
         \38711 , \38712 , \38713 , \38714 , \38715 , \38716 , \38717 , \38718 , \38719 , \38720 ,
         \38721 , \38722 , \38723 , \38724 , \38725 , \38726 , \38727 , \38728 , \38729 , \38730 ,
         \38731 , \38732 , \38733 , \38734 , \38735 , \38736 , \38737 , \38738 , \38739 , \38740 ,
         \38741 , \38742 , \38743 , \38744 , \38745 , \38746 , \38747 , \38748 , \38749 , \38750 ,
         \38751 , \38752 , \38753 , \38754 , \38755 , \38756 , \38757 , \38758 , \38759 , \38760 ,
         \38761 , \38762 , \38763 , \38764 , \38765 , \38766 , \38767 , \38768 , \38769 , \38770 ,
         \38771 , \38772 , \38773 , \38774 , \38775 , \38776 , \38777 , \38778 , \38779 , \38780 ,
         \38781 , \38782 , \38783 , \38784 , \38785 , \38786 , \38787 , \38788 , \38789 , \38790 ,
         \38791 , \38792 , \38793 , \38794 , \38795 , \38796 , \38797 , \38798 , \38799 , \38800 ,
         \38801 , \38802 , \38803 , \38804 , \38805 , \38806 , \38807 , \38808 , \38809 , \38810 ,
         \38811 , \38812 , \38813 , \38814 , \38815 , \38816 , \38817 , \38818 , \38819 , \38820 ,
         \38821 , \38822 , \38823 , \38824 , \38825 , \38826 , \38827 , \38828 , \38829 , \38830 ,
         \38831 , \38832 , \38833 , \38834 , \38835 , \38836 , \38837 , \38838 , \38839 , \38840 ,
         \38841 , \38842 , \38843 , \38844 , \38845 , \38846 , \38847 , \38848 , \38849 , \38850 ,
         \38851 , \38852 , \38853 , \38854 , \38855 , \38856 , \38857 , \38858 , \38859 , \38860 ,
         \38861 , \38862 , \38863 , \38864 , \38865 , \38866 , \38867 , \38868 , \38869 , \38870 ,
         \38871 , \38872 , \38873 , \38874 , \38875 , \38876 , \38877 , \38878 , \38879 , \38880 ,
         \38881 , \38882 , \38883 , \38884 , \38885 , \38886 , \38887 , \38888 , \38889 , \38890 ,
         \38891 , \38892 , \38893 , \38894 , \38895 , \38896 , \38897 , \38898 , \38899 , \38900 ,
         \38901 , \38902 , \38903 , \38904 , \38905 , \38906 , \38907 , \38908 , \38909 , \38910 ,
         \38911 , \38912 , \38913 , \38914 , \38915 , \38916 , \38917 , \38918 , \38919 , \38920 ,
         \38921 , \38922 , \38923 , \38924 , \38925 , \38926 , \38927 , \38928 , \38929 , \38930 ,
         \38931 , \38932 , \38933 , \38934 , \38935 , \38936 , \38937 , \38938 , \38939 , \38940 ,
         \38941 , \38942 , \38943 , \38944 , \38945 , \38946 , \38947 , \38948 , \38949 , \38950 ,
         \38951 , \38952 , \38953 , \38954 , \38955 , \38956 , \38957 , \38958 , \38959 , \38960 ,
         \38961 , \38962 , \38963 , \38964 , \38965 , \38966 , \38967 , \38968 , \38969 , \38970 ,
         \38971 , \38972 , \38973 , \38974 , \38975 , \38976 , \38977 , \38978 , \38979 , \38980 ,
         \38981 , \38982 , \38983 , \38984 , \38985 , \38986 , \38987 , \38988 , \38989 , \38990 ,
         \38991 , \38992 , \38993 , \38994 , \38995 , \38996 , \38997 , \38998 , \38999 , \39000 ,
         \39001 , \39002 , \39003 , \39004 , \39005 , \39006 , \39007 , \39008 , \39009 , \39010 ,
         \39011 , \39012 , \39013 , \39014 , \39015 , \39016 , \39017 , \39018 , \39019 , \39020 ,
         \39021 , \39022 , \39023 , \39024 , \39025 , \39026 , \39027 , \39028 , \39029 , \39030 ,
         \39031 , \39032 , \39033 , \39034 , \39035 , \39036 , \39037 , \39038 , \39039 , \39040 ,
         \39041 , \39042 , \39043 , \39044 , \39045 , \39046 , \39047 , \39048 , \39049 , \39050 ,
         \39051 , \39052 , \39053 , \39054 , \39055 , \39056 , \39057 , \39058 , \39059 , \39060 ,
         \39061 , \39062 , \39063 , \39064 , \39065 , \39066 , \39067 , \39068 , \39069 , \39070 ,
         \39071 , \39072 , \39073 , \39074 , \39075 , \39076 , \39077 , \39078 , \39079 , \39080 ,
         \39081 , \39082 , \39083 , \39084 , \39085 , \39086 , \39087 , \39088 , \39089 , \39090 ,
         \39091 , \39092 , \39093 , \39094 , \39095 , \39096 , \39097 , \39098 , \39099 , \39100 ,
         \39101 , \39102 , \39103 , \39104 , \39105 , \39106 , \39107 , \39108 , \39109 , \39110 ,
         \39111 , \39112 , \39113 , \39114 , \39115 , \39116 , \39117 , \39118 , \39119 , \39120 ,
         \39121 , \39122 , \39123 , \39124 , \39125 , \39126 , \39127 , \39128 , \39129 , \39130 ,
         \39131 , \39132 , \39133 , \39134 , \39135 , \39136 , \39137 , \39138 , \39139 , \39140 ,
         \39141 , \39142 , \39143 , \39144 , \39145 , \39146 , \39147 , \39148 , \39149 , \39150 ,
         \39151 , \39152 , \39153 , \39154 , \39155 , \39156 , \39157 , \39158 , \39159 , \39160 ,
         \39161 , \39162 , \39163 , \39164 , \39165 , \39166 , \39167 , \39168 , \39169 , \39170 ,
         \39171 , \39172 , \39173 , \39174 , \39175 , \39176 , \39177 , \39178 , \39179 , \39180 ,
         \39181 , \39182 , \39183 , \39184 , \39185 , \39186 , \39187 , \39188 , \39189 , \39190 ,
         \39191 , \39192 , \39193 , \39194 , \39195 , \39196 , \39197 , \39198 , \39199 , \39200 ,
         \39201 , \39202 , \39203 , \39204 , \39205 , \39206 , \39207 , \39208 , \39209 , \39210 ,
         \39211 , \39212 , \39213 , \39214 , \39215 , \39216 , \39217 , \39218 , \39219 , \39220 ,
         \39221 , \39222 , \39223 , \39224 , \39225 , \39226 , \39227 , \39228 , \39229 , \39230 ,
         \39231 , \39232 , \39233 , \39234 , \39235 , \39236 , \39237 , \39238 , \39239 , \39240 ,
         \39241 , \39242 , \39243 , \39244 , \39245 , \39246 , \39247 , \39248 , \39249 , \39250 ,
         \39251 , \39252 , \39253 , \39254 , \39255 , \39256 , \39257 , \39258 , \39259 , \39260 ,
         \39261 , \39262 , \39263 , \39264 , \39265 , \39266 , \39267 , \39268 , \39269 , \39270 ,
         \39271 , \39272 , \39273 , \39274 , \39275 , \39276 , \39277 , \39278 , \39279 , \39280 ,
         \39281 , \39282 , \39283 , \39284 , \39285 , \39286 , \39287 , \39288 , \39289 , \39290 ,
         \39291 , \39292 , \39293 , \39294 , \39295 , \39296 , \39297 , \39298 , \39299 , \39300 ,
         \39301 , \39302 , \39303 , \39304 , \39305 , \39306 , \39307 , \39308 , \39309 , \39310 ,
         \39311 , \39312 , \39313 , \39314 , \39315 , \39316 , \39317 , \39318 , \39319 , \39320 ,
         \39321 , \39322 , \39323 , \39324 , \39325 , \39326 , \39327 , \39328 , \39329 , \39330 ,
         \39331 , \39332 , \39333 , \39334 , \39335 , \39336 , \39337 , \39338 , \39339 , \39340 ,
         \39341 , \39342 , \39343 , \39344 , \39345 , \39346 , \39347 , \39348 , \39349 , \39350 ,
         \39351 , \39352 , \39353 , \39354 , \39355 , \39356 , \39357 , \39358 , \39359 , \39360 ,
         \39361 , \39362 , \39363 , \39364 , \39365 , \39366 , \39367 , \39368 , \39369 , \39370 ,
         \39371 , \39372 , \39373 , \39374 , \39375 , \39376 , \39377 , \39378 , \39379 , \39380 ,
         \39381 , \39382 , \39383 , \39384 , \39385 , \39386 , \39387 , \39388 , \39389 , \39390 ,
         \39391 , \39392 , \39393 , \39394 , \39395 , \39396 , \39397 , \39398 , \39399 , \39400 ,
         \39401 , \39402 , \39403 , \39404 , \39405 , \39406 , \39407 , \39408 , \39409 , \39410 ,
         \39411 , \39412 , \39413 , \39414 , \39415 , \39416 , \39417 , \39418 , \39419 , \39420 ,
         \39421 , \39422 , \39423 , \39424 , \39425 , \39426 , \39427 , \39428 , \39429 , \39430 ,
         \39431 , \39432 , \39433 , \39434 , \39435 , \39436 , \39437 , \39438 , \39439 , \39440 ,
         \39441 , \39442 , \39443 , \39444 , \39445 , \39446 , \39447 , \39448 , \39449 , \39450 ,
         \39451 , \39452 , \39453 , \39454 , \39455 , \39456 , \39457 , \39458 , \39459 , \39460 ,
         \39461 , \39462 , \39463 , \39464 , \39465 , \39466 , \39467 , \39468 , \39469 , \39470 ,
         \39471 , \39472 , \39473 , \39474 , \39475 , \39476 , \39477 , \39478 , \39479 , \39480 ,
         \39481 , \39482 , \39483 , \39484 , \39485 , \39486 , \39487 , \39488 , \39489 , \39490 ,
         \39491 , \39492 , \39493 , \39494 , \39495 , \39496 , \39497 , \39498 , \39499 , \39500 ,
         \39501 , \39502 , \39503 , \39504 , \39505 , \39506 , \39507 , \39508 , \39509 , \39510 ,
         \39511 , \39512 , \39513 , \39514 , \39515 , \39516 , \39517 , \39518 , \39519 , \39520 ,
         \39521 , \39522 , \39523 , \39524 , \39525 , \39526 , \39527 , \39528 , \39529 , \39530 ,
         \39531 , \39532 , \39533 , \39534 , \39535 , \39536 , \39537 , \39538 , \39539 , \39540 ,
         \39541 , \39542 , \39543 , \39544 , \39545 , \39546 , \39547 , \39548 , \39549 , \39550 ,
         \39551 , \39552 , \39553 , \39554 , \39555 , \39556 , \39557 , \39558 , \39559 , \39560 ,
         \39561 , \39562 , \39563 , \39564 , \39565 , \39566 , \39567 , \39568 , \39569 , \39570 ,
         \39571 , \39572 , \39573 , \39574 , \39575 , \39576 , \39577 , \39578 , \39579 , \39580 ,
         \39581 , \39582 , \39583 , \39584 , \39585 , \39586 , \39587 , \39588 , \39589 , \39590 ,
         \39591 , \39592 , \39593 , \39594 , \39595 , \39596 , \39597 , \39598 , \39599 , \39600 ,
         \39601 , \39602 , \39603 , \39604 , \39605 , \39606 , \39607 , \39608 , \39609 , \39610 ,
         \39611 , \39612 , \39613 , \39614 , \39615 , \39616 , \39617 , \39618 , \39619 , \39620 ,
         \39621 , \39622 , \39623 , \39624 , \39625 , \39626 , \39627 , \39628 , \39629 , \39630 ,
         \39631 , \39632 , \39633 , \39634 , \39635 , \39636 , \39637 , \39638 , \39639 , \39640 ,
         \39641 , \39642 , \39643 , \39644 , \39645 , \39646 , \39647 , \39648 , \39649 , \39650 ,
         \39651 , \39652 , \39653 , \39654 , \39655 , \39656 , \39657 , \39658 , \39659 , \39660 ,
         \39661 , \39662 , \39663 , \39664 , \39665 , \39666 , \39667 , \39668 , \39669 , \39670 ,
         \39671 , \39672 , \39673 , \39674 , \39675 , \39676 , \39677 , \39678 , \39679 , \39680 ,
         \39681 , \39682 , \39683 , \39684 , \39685 , \39686 , \39687 , \39688 , \39689 , \39690 ,
         \39691 , \39692 , \39693 , \39694 , \39695 , \39696 , \39697 , \39698 , \39699 , \39700 ,
         \39701 , \39702 , \39703 , \39704 , \39705 , \39706 , \39707 , \39708 , \39709 , \39710 ,
         \39711 , \39712 , \39713 , \39714 , \39715 , \39716 , \39717 , \39718 , \39719 , \39720 ,
         \39721 , \39722 , \39723 , \39724 , \39725 , \39726 , \39727 , \39728 , \39729 , \39730 ,
         \39731 , \39732 , \39733 , \39734 , \39735 , \39736 , \39737 , \39738 , \39739 , \39740 ,
         \39741 , \39742 , \39743 , \39744 , \39745 , \39746 , \39747 , \39748 , \39749 , \39750 ,
         \39751 , \39752 , \39753 , \39754 , \39755 , \39756 , \39757 , \39758 , \39759 , \39760 ,
         \39761 , \39762 , \39763 , \39764 , \39765 , \39766 , \39767 , \39768 , \39769 , \39770 ,
         \39771 , \39772 , \39773 , \39774 , \39775 , \39776 , \39777 , \39778 , \39779 , \39780 ,
         \39781 , \39782 , \39783 , \39784 , \39785 , \39786 , \39787 , \39788 , \39789 , \39790 ,
         \39791 , \39792 , \39793 , \39794 , \39795 , \39796 , \39797 , \39798 , \39799 , \39800 ,
         \39801 , \39802 , \39803 , \39804 , \39805 , \39806 , \39807 , \39808 , \39809 , \39810 ,
         \39811 , \39812 , \39813 , \39814 , \39815 , \39816 , \39817 , \39818 , \39819 , \39820 ,
         \39821 , \39822 , \39823 , \39824 , \39825 , \39826 , \39827 , \39828 , \39829 , \39830 ,
         \39831 , \39832 , \39833 , \39834 , \39835 , \39836 , \39837 , \39838 , \39839 , \39840 ,
         \39841 , \39842 , \39843 , \39844 , \39845 , \39846 , \39847 , \39848 , \39849 , \39850 ,
         \39851 , \39852 , \39853 , \39854 , \39855 , \39856 , \39857 , \39858 , \39859 , \39860 ,
         \39861 , \39862 , \39863 , \39864 , \39865 , \39866 , \39867 , \39868 , \39869 , \39870 ,
         \39871 , \39872 , \39873 , \39874 , \39875 , \39876 , \39877 , \39878 , \39879 , \39880 ,
         \39881 , \39882 , \39883 , \39884 , \39885 , \39886 , \39887 , \39888 , \39889 , \39890 ,
         \39891 , \39892 , \39893 , \39894 , \39895 , \39896 , \39897 , \39898 , \39899 , \39900 ,
         \39901 , \39902 , \39903 , \39904 , \39905 , \39906 , \39907 , \39908 , \39909 , \39910 ,
         \39911 , \39912 , \39913 , \39914 , \39915 , \39916 , \39917 , \39918 , \39919 , \39920 ,
         \39921 , \39922 , \39923 , \39924 , \39925 , \39926 , \39927 , \39928 , \39929 , \39930 ,
         \39931 , \39932 , \39933 , \39934 , \39935 , \39936 , \39937 , \39938 , \39939 , \39940 ,
         \39941 , \39942 , \39943 , \39944 , \39945 , \39946 , \39947 , \39948 , \39949 , \39950 ,
         \39951 , \39952 , \39953 , \39954 , \39955 , \39956 , \39957 , \39958 , \39959 , \39960 ,
         \39961 , \39962 , \39963 , \39964 , \39965 , \39966 , \39967 , \39968 , \39969 , \39970 ,
         \39971 , \39972 , \39973 , \39974 , \39975 , \39976 , \39977 , \39978 , \39979 , \39980 ,
         \39981 , \39982 , \39983 , \39984 , \39985 , \39986 , \39987 , \39988 , \39989 , \39990 ,
         \39991 , \39992 , \39993 , \39994 , \39995 , \39996 , \39997 , \39998 , \39999 , \40000 ,
         \40001 , \40002 , \40003 , \40004 , \40005 , \40006 , \40007 , \40008 , \40009 , \40010 ,
         \40011 , \40012 , \40013 , \40014 , \40015 , \40016 , \40017 , \40018 , \40019 , \40020 ,
         \40021 , \40022 , \40023 , \40024 , \40025 , \40026 , \40027 , \40028 , \40029 , \40030 ,
         \40031 , \40032 , \40033 , \40034 , \40035 , \40036 , \40037 , \40038 , \40039 , \40040 ,
         \40041 , \40042 , \40043 , \40044 , \40045 , \40046 , \40047 , \40048 , \40049 , \40050 ,
         \40051 , \40052 , \40053 , \40054 , \40055 , \40056 , \40057 , \40058 , \40059 , \40060 ,
         \40061 , \40062 , \40063 , \40064 , \40065 , \40066 , \40067 , \40068 , \40069 , \40070 ,
         \40071 , \40072 , \40073 , \40074 , \40075 , \40076 , \40077 , \40078 , \40079 , \40080 ,
         \40081 , \40082 , \40083 , \40084 , \40085 , \40086 , \40087 , \40088 , \40089 , \40090 ,
         \40091 , \40092 , \40093 , \40094 , \40095 , \40096 , \40097 , \40098 , \40099 , \40100 ,
         \40101 , \40102 , \40103 , \40104 , \40105 , \40106 , \40107 , \40108 , \40109 , \40110 ,
         \40111 , \40112 , \40113 , \40114 , \40115 , \40116 , \40117 , \40118 , \40119 , \40120 ,
         \40121 , \40122 , \40123 , \40124 , \40125 , \40126 , \40127 , \40128 , \40129 , \40130 ,
         \40131 , \40132 , \40133 , \40134 , \40135 , \40136 , \40137 , \40138 , \40139 , \40140 ,
         \40141 , \40142 , \40143 , \40144 , \40145 , \40146 , \40147 , \40148 , \40149 , \40150 ,
         \40151 , \40152 , \40153 , \40154 , \40155 , \40156 , \40157 , \40158 , \40159 , \40160 ,
         \40161 , \40162 , \40163 , \40164 , \40165 , \40166 , \40167 , \40168 , \40169 , \40170 ,
         \40171 , \40172 , \40173 , \40174 , \40175 , \40176 , \40177 , \40178 , \40179 , \40180 ,
         \40181 , \40182 , \40183 , \40184 , \40185 , \40186 , \40187 , \40188 , \40189 , \40190 ,
         \40191 , \40192 , \40193 , \40194 , \40195 , \40196 , \40197 , \40198 , \40199 , \40200 ,
         \40201 , \40202 , \40203 , \40204 , \40205 , \40206 , \40207 , \40208 , \40209 , \40210 ,
         \40211 , \40212 , \40213 , \40214 , \40215 , \40216 , \40217 , \40218 , \40219 , \40220 ,
         \40221 , \40222 , \40223 , \40224 , \40225 , \40226 , \40227 , \40228 , \40229 , \40230 ,
         \40231 , \40232 , \40233 , \40234 , \40235 , \40236 , \40237 , \40238 , \40239 , \40240 ,
         \40241 , \40242 , \40243 , \40244 , \40245 , \40246 , \40247 , \40248 , \40249 , \40250 ,
         \40251 , \40252 , \40253 , \40254 , \40255 , \40256 , \40257 , \40258 , \40259 , \40260 ,
         \40261 , \40262 , \40263 , \40264 , \40265 , \40266 , \40267 , \40268 , \40269 , \40270 ,
         \40271 , \40272 , \40273 , \40274 , \40275 , \40276 , \40277 , \40278 , \40279 , \40280 ,
         \40281 , \40282 , \40283 , \40284 , \40285 , \40286 , \40287 , \40288 , \40289 , \40290 ,
         \40291 , \40292 , \40293 , \40294 , \40295 , \40296 , \40297 , \40298 , \40299 , \40300 ,
         \40301 , \40302 , \40303 , \40304 , \40305 , \40306 , \40307 , \40308 , \40309 , \40310 ,
         \40311 , \40312 , \40313 , \40314 , \40315 , \40316 , \40317 , \40318 , \40319 , \40320 ,
         \40321 , \40322 , \40323 , \40324 , \40325 , \40326 , \40327 , \40328 , \40329 , \40330 ,
         \40331 , \40332 , \40333 , \40334 , \40335 , \40336 , \40337 , \40338 , \40339 , \40340 ,
         \40341 , \40342 , \40343 , \40344 , \40345 , \40346 , \40347 , \40348 , \40349 , \40350 ,
         \40351 , \40352 , \40353 , \40354 , \40355 , \40356 , \40357 , \40358 , \40359 , \40360 ,
         \40361 , \40362 , \40363 , \40364 , \40365 , \40366 , \40367 , \40368 , \40369 , \40370 ,
         \40371 , \40372 , \40373 , \40374 , \40375 , \40376 , \40377 , \40378 , \40379 , \40380 ,
         \40381 , \40382 , \40383 , \40384 , \40385 , \40386 , \40387 , \40388 , \40389 , \40390 ,
         \40391 , \40392 , \40393 , \40394 , \40395 , \40396 , \40397 , \40398 , \40399 , \40400 ,
         \40401 , \40402 , \40403 , \40404 , \40405 , \40406 , \40407 , \40408 , \40409 , \40410 ,
         \40411 , \40412 , \40413 , \40414 , \40415 , \40416 , \40417 , \40418 , \40419 , \40420 ,
         \40421 , \40422 , \40423 , \40424 , \40425 , \40426 , \40427 , \40428 , \40429 , \40430 ,
         \40431 , \40432 , \40433 , \40434 , \40435 , \40436 , \40437 , \40438 , \40439 , \40440 ,
         \40441 , \40442 , \40443 , \40444 , \40445 , \40446 , \40447 , \40448 , \40449 , \40450 ,
         \40451 , \40452 , \40453 , \40454 , \40455 , \40456 , \40457 , \40458 , \40459 , \40460 ,
         \40461 , \40462 , \40463 , \40464 , \40465 , \40466 , \40467 , \40468 , \40469 , \40470 ,
         \40471 , \40472 , \40473 , \40474 , \40475 , \40476 , \40477 , \40478 , \40479 , \40480 ,
         \40481 , \40482 , \40483 , \40484 , \40485 , \40486 , \40487 , \40488 , \40489 , \40490 ,
         \40491 , \40492 , \40493 , \40494 , \40495 , \40496 , \40497 , \40498 , \40499 , \40500 ,
         \40501 , \40502 , \40503 , \40504 , \40505 , \40506 , \40507 , \40508 , \40509 , \40510 ,
         \40511 , \40512 , \40513 , \40514 , \40515 , \40516 , \40517 , \40518 , \40519 , \40520 ,
         \40521 , \40522 , \40523 , \40524 , \40525 , \40526 , \40527 , \40528 , \40529 , \40530 ,
         \40531 , \40532 , \40533 , \40534 , \40535 , \40536 , \40537 , \40538 , \40539 , \40540 ,
         \40541 , \40542 , \40543 , \40544 , \40545 , \40546 , \40547 , \40548 , \40549 , \40550 ,
         \40551 , \40552 , \40553 , \40554 , \40555 , \40556 , \40557 , \40558 , \40559 , \40560 ,
         \40561 , \40562 , \40563 , \40564 , \40565 , \40566 , \40567 , \40568 , \40569 , \40570 ,
         \40571 , \40572 , \40573 , \40574 , \40575 , \40576 , \40577 , \40578 , \40579 , \40580 ,
         \40581 , \40582 , \40583 , \40584 , \40585 , \40586 , \40587 , \40588 , \40589 , \40590 ,
         \40591 , \40592 , \40593 , \40594 , \40595 , \40596 , \40597 , \40598 , \40599 , \40600 ,
         \40601 , \40602 , \40603 , \40604 , \40605 , \40606 , \40607 , \40608 , \40609 , \40610 ,
         \40611 , \40612 , \40613 , \40614 , \40615 , \40616 , \40617 , \40618 , \40619 , \40620 ,
         \40621 , \40622 , \40623 , \40624 , \40625 , \40626 , \40627 , \40628 , \40629 , \40630 ,
         \40631 , \40632 , \40633 , \40634 , \40635 , \40636 , \40637 , \40638 , \40639 , \40640 ,
         \40641 , \40642 , \40643 , \40644 , \40645 , \40646 , \40647 , \40648 , \40649 , \40650 ,
         \40651 , \40652 , \40653 , \40654 , \40655 , \40656 , \40657 , \40658 , \40659 , \40660 ,
         \40661 , \40662 , \40663 , \40664 , \40665 , \40666 , \40667 , \40668 , \40669 , \40670 ,
         \40671 , \40672 , \40673 , \40674 , \40675 , \40676 , \40677 , \40678 , \40679 , \40680 ,
         \40681 , \40682 , \40683 , \40684 , \40685 , \40686 , \40687 , \40688 , \40689 , \40690 ,
         \40691 , \40692 , \40693 , \40694 , \40695 , \40696 , \40697 , \40698 , \40699 , \40700 ,
         \40701 , \40702 , \40703 , \40704 , \40705 , \40706 , \40707 , \40708 , \40709 , \40710 ,
         \40711 , \40712 , \40713 , \40714 , \40715 , \40716 , \40717 , \40718 , \40719 , \40720 ,
         \40721 , \40722 , \40723 , \40724 , \40725 , \40726 , \40727 , \40728 , \40729 , \40730 ,
         \40731 , \40732 , \40733 , \40734 , \40735 , \40736 , \40737 , \40738 , \40739 , \40740 ,
         \40741 , \40742 , \40743 , \40744 , \40745 , \40746 , \40747 , \40748 , \40749 , \40750 ,
         \40751 , \40752 , \40753 , \40754 , \40755 , \40756 , \40757 , \40758 , \40759 , \40760 ,
         \40761 , \40762 , \40763 , \40764 , \40765 , \40766 , \40767 , \40768 , \40769 , \40770 ,
         \40771 , \40772 , \40773 , \40774 , \40775 , \40776 , \40777 , \40778 , \40779 , \40780 ,
         \40781 , \40782 , \40783 , \40784 , \40785 , \40786 , \40787 , \40788 , \40789 , \40790 ,
         \40791 , \40792 , \40793 , \40794 , \40795 , \40796 , \40797 , \40798 , \40799 , \40800 ,
         \40801 , \40802 , \40803 , \40804 , \40805 , \40806 , \40807 , \40808 , \40809 , \40810 ,
         \40811 , \40812 , \40813 , \40814 , \40815 , \40816 , \40817 , \40818 , \40819 , \40820 ,
         \40821 , \40822 , \40823 , \40824 , \40825 , \40826 , \40827 , \40828 , \40829 , \40830 ,
         \40831 , \40832 , \40833 , \40834 , \40835 , \40836 , \40837 , \40838 , \40839 , \40840 ,
         \40841 , \40842 , \40843 , \40844 , \40845 , \40846 , \40847 , \40848 , \40849 , \40850 ,
         \40851 , \40852 , \40853 , \40854 , \40855 , \40856 , \40857 , \40858 , \40859 , \40860 ,
         \40861 , \40862 , \40863 , \40864 , \40865 , \40866 , \40867 , \40868 , \40869 , \40870 ,
         \40871 , \40872 , \40873 , \40874 , \40875 , \40876 , \40877 , \40878 , \40879 , \40880 ,
         \40881 , \40882 , \40883 , \40884 , \40885 , \40886 , \40887 , \40888 , \40889 , \40890 ,
         \40891 , \40892 , \40893 , \40894 , \40895 , \40896 , \40897 , \40898 , \40899 , \40900 ,
         \40901 , \40902 , \40903 , \40904 , \40905 , \40906 , \40907 , \40908 , \40909 , \40910 ,
         \40911 , \40912 , \40913 , \40914 , \40915 , \40916 , \40917 , \40918 , \40919 , \40920 ,
         \40921 , \40922 , \40923 , \40924 , \40925 , \40926 , \40927 , \40928 , \40929 , \40930 ,
         \40931 , \40932 , \40933 , \40934 , \40935 , \40936 , \40937 , \40938 , \40939 , \40940 ,
         \40941 , \40942 , \40943 , \40944 , \40945 , \40946 , \40947 , \40948 , \40949 , \40950 ,
         \40951 , \40952 , \40953 , \40954 , \40955 , \40956 , \40957 , \40958 , \40959 , \40960 ,
         \40961 , \40962 , \40963 , \40964 , \40965 , \40966 , \40967 , \40968 , \40969 , \40970 ,
         \40971 , \40972 , \40973 , \40974 , \40975 , \40976 , \40977 , \40978 , \40979 , \40980 ,
         \40981 , \40982 , \40983 , \40984 , \40985 , \40986 , \40987 , \40988 , \40989 , \40990 ,
         \40991 , \40992 , \40993 , \40994 , \40995 , \40996 , \40997 , \40998 , \40999 , \41000 ,
         \41001 , \41002 , \41003 , \41004 , \41005 , \41006 , \41007 , \41008 , \41009 , \41010 ,
         \41011 , \41012 , \41013 , \41014 , \41015 , \41016 , \41017 , \41018 , \41019 , \41020 ,
         \41021 , \41022 , \41023 , \41024 , \41025 , \41026 , \41027 , \41028 , \41029 , \41030 ,
         \41031 , \41032 , \41033 , \41034 , \41035 , \41036 , \41037 , \41038 , \41039 , \41040 ,
         \41041 , \41042 , \41043 , \41044 , \41045 , \41046 , \41047 , \41048 , \41049 , \41050 ,
         \41051 , \41052 , \41053 , \41054 , \41055 , \41056 , \41057 , \41058 , \41059 , \41060 ,
         \41061 , \41062 , \41063 , \41064 , \41065 , \41066 , \41067 , \41068 , \41069 , \41070 ,
         \41071 , \41072 , \41073 , \41074 , \41075 , \41076 , \41077 , \41078 , \41079 , \41080 ,
         \41081 , \41082 , \41083 , \41084 , \41085 , \41086 , \41087 , \41088 , \41089 , \41090 ,
         \41091 , \41092 , \41093 , \41094 , \41095 , \41096 , \41097 , \41098 , \41099 , \41100 ,
         \41101 , \41102 , \41103 , \41104 , \41105 , \41106 , \41107 , \41108 , \41109 , \41110 ,
         \41111 , \41112 , \41113 , \41114 , \41115 , \41116 , \41117 , \41118 , \41119 , \41120 ,
         \41121 , \41122 , \41123 , \41124 , \41125 , \41126 , \41127 , \41128 , \41129 , \41130 ,
         \41131 , \41132 , \41133 , \41134 , \41135 , \41136 , \41137 , \41138 , \41139 , \41140 ,
         \41141 , \41142 , \41143 , \41144 , \41145 , \41146 , \41147 , \41148 , \41149 , \41150 ,
         \41151 , \41152 , \41153 , \41154 , \41155 , \41156 , \41157 , \41158 , \41159 , \41160 ,
         \41161 , \41162 , \41163 , \41164 , \41165 , \41166 , \41167 , \41168 , \41169 , \41170 ,
         \41171 , \41172 , \41173 , \41174 , \41175 , \41176 , \41177 , \41178 , \41179 , \41180 ,
         \41181 , \41182 , \41183 , \41184 , \41185 , \41186 , \41187 , \41188 , \41189 , \41190 ,
         \41191 , \41192 , \41193 , \41194 , \41195 , \41196 , \41197 , \41198 , \41199 , \41200 ,
         \41201 , \41202 , \41203 , \41204 , \41205 , \41206 , \41207 , \41208 , \41209 , \41210 ,
         \41211 , \41212 , \41213 , \41214 , \41215 , \41216 , \41217 , \41218 , \41219 , \41220 ,
         \41221 , \41222 , \41223 , \41224 , \41225 , \41226 , \41227 , \41228 , \41229 , \41230 ,
         \41231 , \41232 , \41233 , \41234 , \41235 , \41236 , \41237 , \41238 , \41239 , \41240 ,
         \41241 , \41242 , \41243 , \41244 , \41245 , \41246 , \41247 , \41248 , \41249 , \41250 ,
         \41251 , \41252 , \41253 , \41254 , \41255 , \41256 , \41257 , \41258 , \41259 , \41260 ,
         \41261 , \41262 , \41263 , \41264 , \41265 , \41266 , \41267 , \41268 , \41269 , \41270 ,
         \41271 , \41272 , \41273 , \41274 , \41275 , \41276 , \41277 , \41278 , \41279 , \41280 ,
         \41281 , \41282 , \41283 , \41284 , \41285 , \41286 , \41287 , \41288 , \41289 , \41290 ,
         \41291 , \41292 , \41293 , \41294 , \41295 , \41296 , \41297 , \41298 , \41299 , \41300 ,
         \41301 , \41302 , \41303 , \41304 , \41305 , \41306 , \41307 , \41308 , \41309 , \41310 ,
         \41311 , \41312 , \41313 , \41314 , \41315 , \41316 , \41317 , \41318 , \41319 , \41320 ,
         \41321 , \41322 , \41323 , \41324 , \41325 , \41326 , \41327 , \41328 , \41329 , \41330 ,
         \41331 , \41332 , \41333 , \41334 , \41335 , \41336 , \41337 , \41338 , \41339 , \41340 ,
         \41341 , \41342 , \41343 , \41344 , \41345 , \41346 , \41347 , \41348 , \41349 , \41350 ,
         \41351 , \41352 , \41353 , \41354 , \41355 , \41356 , \41357 , \41358 , \41359 , \41360 ,
         \41361 , \41362 , \41363 , \41364 , \41365 , \41366 , \41367 , \41368 , \41369 , \41370 ,
         \41371 , \41372 , \41373 , \41374 , \41375 , \41376 , \41377 , \41378 , \41379 , \41380 ,
         \41381 , \41382 , \41383 , \41384 , \41385 , \41386 , \41387 , \41388 , \41389 , \41390 ,
         \41391 , \41392 , \41393 , \41394 , \41395 , \41396 , \41397 , \41398 , \41399 , \41400 ,
         \41401 , \41402 , \41403 , \41404 , \41405 , \41406 , \41407 , \41408 , \41409 , \41410 ,
         \41411 , \41412 , \41413 , \41414 , \41415 , \41416 , \41417 , \41418 , \41419 , \41420 ,
         \41421 , \41422 , \41423 , \41424 , \41425 , \41426 , \41427 , \41428 , \41429 , \41430 ,
         \41431 , \41432 , \41433 , \41434 , \41435 , \41436 , \41437 , \41438 , \41439 , \41440 ,
         \41441 , \41442 , \41443 , \41444 , \41445 , \41446 , \41447 , \41448 , \41449 , \41450 ,
         \41451 , \41452 , \41453 , \41454 , \41455 , \41456 , \41457 , \41458 , \41459 , \41460 ,
         \41461 , \41462 , \41463 , \41464 , \41465 , \41466 , \41467 , \41468 , \41469 , \41470 ,
         \41471 , \41472 , \41473 , \41474 , \41475 , \41476 , \41477 , \41478 , \41479 , \41480 ,
         \41481 , \41482 , \41483 , \41484 , \41485 , \41486 , \41487 , \41488 , \41489 , \41490 ,
         \41491 , \41492 , \41493 , \41494 , \41495 , \41496 , \41497 , \41498 , \41499 , \41500 ,
         \41501 , \41502 , \41503 , \41504 , \41505 , \41506 , \41507 , \41508 , \41509 , \41510 ,
         \41511 , \41512 , \41513 , \41514 , \41515 , \41516 , \41517 , \41518 , \41519 , \41520 ,
         \41521 , \41522 , \41523 , \41524 , \41525 , \41526 , \41527 , \41528 , \41529 , \41530 ,
         \41531 , \41532 , \41533 , \41534 , \41535 , \41536 , \41537 , \41538 , \41539 , \41540 ,
         \41541 , \41542 , \41543 , \41544 , \41545 , \41546 , \41547 , \41548 , \41549 , \41550 ,
         \41551 , \41552 , \41553 , \41554 , \41555 , \41556 , \41557 , \41558 , \41559 , \41560 ,
         \41561 , \41562 , \41563 , \41564 , \41565 , \41566 , \41567 , \41568 , \41569 , \41570 ,
         \41571 , \41572 , \41573 , \41574 , \41575 , \41576 , \41577 , \41578 , \41579 , \41580 ,
         \41581 , \41582 , \41583 , \41584 , \41585 , \41586 , \41587 , \41588 , \41589 , \41590 ,
         \41591 , \41592 , \41593 , \41594 , \41595 , \41596 , \41597 , \41598 , \41599 , \41600 ,
         \41601 , \41602 , \41603 , \41604 , \41605 , \41606 , \41607 , \41608 , \41609 , \41610 ,
         \41611 , \41612 , \41613 , \41614 , \41615 , \41616 , \41617 , \41618 , \41619 , \41620 ,
         \41621 , \41622 , \41623 , \41624 , \41625 , \41626 , \41627 , \41628 , \41629 , \41630 ,
         \41631 , \41632 , \41633 , \41634 , \41635 , \41636 , \41637 , \41638 , \41639 , \41640 ,
         \41641 , \41642 , \41643 , \41644 , \41645 , \41646 , \41647 , \41648 , \41649 , \41650 ,
         \41651 , \41652 , \41653 , \41654 , \41655 , \41656 , \41657 , \41658 , \41659 , \41660 ,
         \41661 , \41662 , \41663 , \41664 , \41665 , \41666 , \41667 , \41668 , \41669 , \41670 ,
         \41671 , \41672 , \41673 , \41674 , \41675 , \41676 , \41677 , \41678 , \41679 , \41680 ,
         \41681 , \41682 , \41683 , \41684 , \41685 , \41686 , \41687 , \41688 , \41689 , \41690 ,
         \41691 , \41692 , \41693 , \41694 , \41695 , \41696 , \41697 , \41698 , \41699 , \41700 ,
         \41701 , \41702 , \41703 , \41704 , \41705 , \41706 , \41707 , \41708 , \41709 , \41710 ,
         \41711 , \41712 , \41713 , \41714 , \41715 , \41716 , \41717 , \41718 , \41719 , \41720 ,
         \41721 , \41722 , \41723 , \41724 , \41725 , \41726 , \41727 , \41728 , \41729 , \41730 ,
         \41731 , \41732 , \41733 , \41734 , \41735 , \41736 , \41737 , \41738 , \41739 , \41740 ,
         \41741 , \41742 , \41743 , \41744 , \41745 , \41746 , \41747 , \41748 , \41749 , \41750 ,
         \41751 , \41752 , \41753 , \41754 , \41755 , \41756 , \41757 , \41758 , \41759 , \41760 ,
         \41761 , \41762 , \41763 , \41764 , \41765 , \41766 , \41767 , \41768 , \41769 , \41770 ,
         \41771 , \41772 , \41773 , \41774 , \41775 , \41776 , \41777 , \41778 , \41779 , \41780 ,
         \41781 , \41782 , \41783 , \41784 , \41785 , \41786 , \41787 , \41788 , \41789 , \41790 ,
         \41791 , \41792 , \41793 , \41794 , \41795 , \41796 , \41797 , \41798 , \41799 , \41800 ,
         \41801 , \41802 , \41803 , \41804 , \41805 , \41806 , \41807 , \41808 , \41809 , \41810 ,
         \41811 , \41812 , \41813 , \41814 , \41815 , \41816 , \41817 , \41818 , \41819 , \41820 ,
         \41821 , \41822 , \41823 , \41824 , \41825 , \41826 , \41827 , \41828 , \41829 , \41830 ,
         \41831 , \41832 , \41833 , \41834 , \41835 , \41836 , \41837 , \41838 , \41839 , \41840 ,
         \41841 , \41842 , \41843 , \41844 , \41845 , \41846 , \41847 , \41848 , \41849 , \41850 ,
         \41851 , \41852 , \41853 , \41854 , \41855 , \41856 , \41857 , \41858 , \41859 , \41860 ,
         \41861 , \41862 , \41863 , \41864 , \41865 , \41866 , \41867 , \41868 , \41869 , \41870 ,
         \41871 , \41872 , \41873 , \41874 , \41875 , \41876 , \41877 , \41878 , \41879 , \41880 ,
         \41881 , \41882 , \41883 , \41884 , \41885 , \41886 , \41887 , \41888 , \41889 , \41890 ,
         \41891 , \41892 , \41893 , \41894 , \41895 , \41896 , \41897 , \41898 , \41899 , \41900 ,
         \41901 , \41902 , \41903 , \41904 , \41905 , \41906 , \41907 , \41908 , \41909 , \41910 ,
         \41911 , \41912 , \41913 , \41914 , \41915 , \41916 , \41917 , \41918 , \41919 , \41920 ,
         \41921 , \41922 , \41923 , \41924 , \41925 , \41926 , \41927 , \41928 , \41929 , \41930 ,
         \41931 , \41932 , \41933 , \41934 , \41935 , \41936 , \41937 , \41938 , \41939 , \41940 ,
         \41941 , \41942 , \41943 , \41944 , \41945 , \41946 , \41947 , \41948 , \41949 , \41950 ,
         \41951 , \41952 , \41953 , \41954 , \41955 , \41956 , \41957 , \41958 , \41959 , \41960 ,
         \41961 , \41962 , \41963 , \41964 , \41965 , \41966 , \41967 , \41968 , \41969 , \41970 ,
         \41971 , \41972 , \41973 , \41974 , \41975 , \41976 , \41977 , \41978 , \41979 , \41980 ,
         \41981 , \41982 , \41983 , \41984 , \41985 , \41986 , \41987 , \41988 , \41989 , \41990 ,
         \41991 , \41992 , \41993 , \41994 , \41995 , \41996 , \41997 , \41998 , \41999 , \42000 ,
         \42001 , \42002 , \42003 , \42004 , \42005 , \42006 , \42007 , \42008 , \42009 , \42010 ,
         \42011 , \42012 , \42013 , \42014 , \42015 , \42016 , \42017 , \42018 , \42019 , \42020 ,
         \42021 , \42022 , \42023 , \42024 , \42025 , \42026 , \42027 , \42028 , \42029 , \42030 ,
         \42031 , \42032 , \42033 , \42034 , \42035 , \42036 , \42037 , \42038 , \42039 , \42040 ,
         \42041 , \42042 , \42043 , \42044 , \42045 , \42046 , \42047 , \42048 , \42049 , \42050 ,
         \42051 , \42052 , \42053 , \42054 , \42055 , \42056 , \42057 , \42058 , \42059 , \42060 ,
         \42061 , \42062 , \42063 , \42064 , \42065 , \42066 , \42067 , \42068 , \42069 , \42070 ,
         \42071 , \42072 , \42073 , \42074 , \42075 , \42076 , \42077 , \42078 , \42079 , \42080 ,
         \42081 , \42082 , \42083 , \42084 , \42085 , \42086 , \42087 , \42088 , \42089 , \42090 ,
         \42091 , \42092 , \42093 , \42094 , \42095 , \42096 , \42097 , \42098 , \42099 , \42100 ,
         \42101 , \42102 , \42103 , \42104 , \42105 , \42106 , \42107 , \42108 , \42109 , \42110 ,
         \42111 , \42112 , \42113 , \42114 , \42115 , \42116 , \42117 , \42118 , \42119 , \42120 ,
         \42121 , \42122 , \42123 , \42124 , \42125 , \42126 , \42127 , \42128 , \42129 , \42130 ,
         \42131 , \42132 , \42133 , \42134 , \42135 , \42136 , \42137 , \42138 , \42139 , \42140 ,
         \42141 , \42142 , \42143 , \42144 , \42145 , \42146 , \42147 , \42148 , \42149 , \42150 ,
         \42151 , \42152 , \42153 , \42154 , \42155 , \42156 , \42157 , \42158 , \42159 , \42160 ,
         \42161 , \42162 , \42163 , \42164 , \42165 , \42166 , \42167 , \42168 , \42169 , \42170 ,
         \42171 , \42172 , \42173 , \42174 , \42175 , \42176 , \42177 , \42178 , \42179 , \42180 ,
         \42181 , \42182 , \42183 , \42184 , \42185 , \42186 , \42187 , \42188 , \42189 , \42190 ,
         \42191 , \42192 , \42193 , \42194 , \42195 , \42196 , \42197 , \42198 , \42199 , \42200 ,
         \42201 , \42202 , \42203 , \42204 , \42205 , \42206 , \42207 , \42208 , \42209 , \42210 ,
         \42211 , \42212 , \42213 , \42214 , \42215 , \42216 , \42217 , \42218 , \42219 , \42220 ,
         \42221 , \42222 , \42223 , \42224 , \42225 , \42226 , \42227 , \42228 , \42229 , \42230 ,
         \42231 , \42232 , \42233 , \42234 , \42235 , \42236 , \42237 , \42238 , \42239 , \42240 ,
         \42241 , \42242 , \42243 , \42244 , \42245 , \42246 , \42247 , \42248 , \42249 , \42250 ,
         \42251 , \42252 , \42253 , \42254 , \42255 , \42256 , \42257 , \42258 , \42259 , \42260 ,
         \42261 , \42262 , \42263 , \42264 , \42265 , \42266 , \42267 , \42268 , \42269 , \42270 ,
         \42271 , \42272 , \42273 , \42274 , \42275 , \42276 , \42277 , \42278 , \42279 , \42280 ,
         \42281 , \42282 , \42283 , \42284 , \42285 , \42286 , \42287 , \42288 , \42289 , \42290 ,
         \42291 , \42292 , \42293 , \42294 , \42295 , \42296 , \42297 , \42298 , \42299 , \42300 ,
         \42301 , \42302 , \42303 , \42304 , \42305 , \42306 , \42307 , \42308 , \42309 , \42310 ,
         \42311 , \42312 , \42313 , \42314 , \42315 , \42316 , \42317 , \42318 , \42319 , \42320 ,
         \42321 , \42322 , \42323 , \42324 , \42325 , \42326 , \42327 , \42328 , \42329 , \42330 ,
         \42331 , \42332 , \42333 , \42334 , \42335 , \42336 , \42337 , \42338 , \42339 , \42340 ,
         \42341 , \42342 , \42343 , \42344 , \42345 , \42346 , \42347 , \42348 , \42349 , \42350 ,
         \42351 , \42352 , \42353 , \42354 , \42355 , \42356 , \42357 , \42358 , \42359 , \42360 ,
         \42361 , \42362 , \42363 , \42364 , \42365 , \42366 , \42367 , \42368 , \42369 , \42370 ,
         \42371 , \42372 , \42373 , \42374 , \42375 , \42376 , \42377 , \42378 , \42379 , \42380 ,
         \42381 , \42382 , \42383 , \42384 , \42385 , \42386 , \42387 , \42388 , \42389 , \42390 ,
         \42391 , \42392 , \42393 , \42394 , \42395 , \42396 , \42397 , \42398_nGac83 , \42399 , \42400 ,
         \42401 , \42402_nGabce , \42403 , \42404 , \42405_nGac0d , \42406 , \42407 , \42408 , \42409_nGab43 , \42410 ,
         \42411 , \42412_nGab87 , \42413 , \42414 , \42415 , \42416_nGaab0 , \42417 , \42418 , \42419_nGaaf7 , \42420 ,
         \42421 , \42422 , \42423_nGaa15 , \42424 , \42425 , \42426_nGaa61 , \42427 , \42428 , \42429 , \42430_nGa96e ,
         \42431 , \42432 , \42433_nGa9c1 , \42434 , \42435 , \42436 , \42437_nGa8be , \42438 , \42439 , \42440_nGa913 ,
         \42441 , \42442 , \42443 , \42444_nGa804 , \42445 , \42446 , \42447_nGa861 , \42448 , \42449 , \42450 ,
         \42451_nGa740 , \42452 , \42453 , \42454_nGa79f , \42455 , \42456 , \42457 , \42458_nGa672 , \42459 , \42460 ,
         \42461_nGa6d9 , \42462 , \42463 , \42464 , \42465_nGa59a , \42466 , \42467 , \42468_nGa603 , \42469 , \42470 ,
         \42471 , \42472_nGa4bb , \42473 , \42474 , \42475_nGa529 , \42476 , \42477 , \42478 , \42479_nGa3d1 , \42480 ,
         \42481 , \42482_nGa445 , \42483 , \42484 , \42485 , \42486_nGa2da , \42487 , \42488 , \42489_nGa355 , \42490 ,
         \42491 , \42492 , \42493_nGa1d7 , \42494 , \42495 , \42496_nGa257 , \42497 , \42498 , \42499 , \42500_nGa0c9 ,
         \42501 , \42502 , \42503_nGa14f , \42504 , \42505 , \42506 , \42507_nG9fb4 , \42508 , \42509 , \42510_nGa03b ,
         \42511 , \42512 , \42513 , \42514_nG9e96 , \42515 , \42516 , \42517_nG9f25 , \42518 , \42519 , \42520 ,
         \42521_nG9d6b , \42522 , \42523 , \42524_nG9dff , \42525 , \42526 , \42527 , \42528_nG9c34 , \42529 , \42530 ,
         \42531_nG9ccf , \42532 , \42533 , \42534 , \42535_nG9af1 , \42536 , \42537 , \42538_nG9b91 , \42539 , \42540 ,
         \42541 , \42542_nG99a6 , \42543 , \42544 , \42545_nG9a49 , \42546 , \42547 , \42548 , \42549_nG9856 , \42550 ,
         \42551 , \42552_nG98fb , \42553 , \42554 , \42555 , \42556_nG96ff , \42557 , \42558 , \42559_nG97a9 , \42560 ,
         \42561 , \42562 , \42563_nG95a0 , \42564 , \42565 , \42566_nG964d , \42567 , \42568 , \42569 , \42570_nG9436 ,
         \42571 , \42572 , \42573_nG94eb , \42574 , \42575 , \42576 , \42577_nG92bf , \42578 , \42579 , \42580_nG9379 ,
         \42581 , \42582 , \42583 , \42584_nG913c , \42585 , \42586 , \42587_nG91fd , \42588 , \42589 , \42590 ,
         \42591_nG8fb0 , \42592 , \42593 , \42594_nG9073 , \42595 , \42596 , \42597 , \42598_nG8e1a , \42599 , \42600 ,
         \42601_nG8ee5 , \42602 , \42603 , \42604 , \42605_nG8c7a , \42606 , \42607 , \42608_nG8d47 , \42609 , \42610 ,
         \42611 , \42612_nG8ad0 , \42613 , \42614 , \42615_nG8ba5 , \42616 , \42617 , \42618 , \42619_nG8919 , \42620 ,
         \42621 , \42622_nG89f3 , \42623 , \42624 , \42625 , \42626_nG8757 , \42627 , \42628 , \42629_nG8837 , \42630 ,
         \42631 , \42632 , \42633_nG858b , \42634 , \42635 , \42636_nG866f , \42637 , \42638 , \42639 , \42640_nG83b4 ,
         \42641 , \42642 , \42643_nG849f , \42644 , \42645 , \42646 , \42647_nG81d4 , \42648 , \42649 , \42650_nG82c1 ,
         \42651 , \42652 , \42653 , \42654_nG7fea , \42655 , \42656 , \42657_nG80df , \42658 , \42659 , \42660 ,
         \42661_nG7df3 , \42662 , \42663 , \42664_nG7eed , \42665 , \42666 , \42667 , \42668_nG7bf4 , \42669 , \42670 ,
         \42671_nG7cf1 , \42672 , \42673 , \42674 , \42675_nG79f0 , \42676 , \42677 , \42678_nG7aef , \42679 , \42680 ,
         \42681 , \42682_nG77e5 , \42683 , \42684 , \42685_nG78e9 , \42686 , \42687 , \42688 , \42689_nG75cf , \42690 ,
         \42691 , \42692_nG76d9 , \42693 , \42694 , \42695 , \42696_nG73af , \42697 , \42698 , \42699_nG74bd , \42700 ,
         \42701 , \42702 , \42703_nG7188 , \42704 , \42705 , \42706_nG7299 , \42707 , \42708 , \42709 , \42710_nG6f56 ,
         \42711 , \42712 , \42713_nG706f , \42714 , \42715 , \42716 , \42717_nG6d1a , \42718 , \42719 , \42720_nG6e35 ,
         \42721 , \42722 , \42723 , \42724_nG6ad4 , \42725 , \42726 , \42727_nG6bf7 , \42728 , \42729 , \42730 ,
         \42731_nG6881 , \42732 , \42733 , \42734_nG69a9 , \42735 , \42736 , \42737 , \42738_nG6622 , \42739 , \42740 ,
         \42741_nG6751 , \42742 , \42743 , \42744 , \42745_nG63b7 , \42746 , \42747 , \42748_nG64eb , \42749 , \42750 ,
         \42751 , \42752_nG6144 , \42753 , \42754 , \42755_nG627b , \42756 , \42757 , \42758 , \42759_nG5ec9 , \42760 ,
         \42761 , \42762_nG6005 , \42763 , \42764 , \42765 , \42766_nG5c48 , \42767 , \42768 , \42769_nG5d85 , \42770 ,
         \42771 , \42772 , \42773_nG59c5 , \42774 , \42775 , \42776_nG5b03 , \42777 , \42778 , \42779 , \42780_nG5740 ,
         \42781 , \42782 , \42783_nG587f , \42784 , \42785 , \42786 , \42787_nG54b8 , \42788 , \42789 , \42790_nG55f9 ,
         \42791 , \42792 , \42793 , \42794_nG5231 , \42795 , \42796 , \42797_nG536f , \42798 , \42799 , \42800 ,
         \42801_nG4fb4 , \42802 , \42803 , \42804_nG50eb , \42805 , \42806 , \42807 , \42808_nG4d41 , \42809 , \42810 ,
         \42811_nG4e75 , \42812 , \42813 , \42814 , \42815_nG4ad8 , \42816 , \42817 , \42818_nG4c05 , \42819 , \42820 ,
         \42821 , \42822_nG4879 , \42823 , \42824 , \42825_nG49a3 , \42826 , \42827 , \42828 , \42829_nG4624 , \42830 ,
         \42831 , \42832_nG4747 , \42833 , \42834 , \42835 , \42836_nG43d9 , \42837 , \42838 , \42839_nG44f9 , \42840 ,
         \42841 , \42842 , \42843_nG4198 , \42844 , \42845 , \42846_nG42b1 , \42847 , \42848 , \42849 , \42850_nG3f61 ,
         \42851 , \42852 , \42853_nG4077 , \42854 , \42855 , \42856 , \42857_nG3d34 , \42858 , \42859 , \42860_nG3e43 ,
         \42861 , \42862 , \42863 , \42864_nG3b11 , \42865 , \42866 , \42867_nG3c1d , \42868 , \42869 , \42870 ,
         \42871_nG38f8 , \42872 , \42873 , \42874_nG39fd , \42875 , \42876 , \42877 , \42878_nG36e9 , \42879 , \42880 ,
         \42881_nG37eb , \42882 , \42883 , \42884 , \42885_nG34e4 , \42886 , \42887 , \42888_nG35df , \42889 , \42890 ,
         \42891 , \42892_nG32e9 , \42893 , \42894 , \42895_nG33e1 , \42896 , \42897 , \42898 , \42899_nG30f8 , \42900 ,
         \42901 , \42902_nG31e9 , \42903 , \42904 , \42905 , \42906_nG2f11 , \42907 , \42908 , \42909_nG2fff , \42910 ,
         \42911 , \42912 , \42913_nG2d34 , \42914 , \42915 , \42916_nG2e1b , \42917 , \42918 , \42919 , \42920_nG2b5e ,
         \42921 , \42922 , \42923_nG2c45 , \42924 , \42925 , \42926 , \42927_nG2993 , \42928 , \42929 , \42930_nG2a6f ,
         \42931 , \42932 , \42933 , \42934_nG27d5 , \42935 , \42936 , \42937_nG28af , \42938 , \42939 , \42940 ,
         \42941_nG2620 , \42942 , \42943 , \42944_nG26f3 , \42945 , \42946 , \42947 , \42948_nG2475 , \42949 , \42950 ,
         \42951_nG2545 , \42952 , \42953 , \42954 , \42955_nG22d4 , \42956 , \42957 , \42958_nG239d , \42959 , \42960 ,
         \42961 , \42962_nG213d , \42963 , \42964 , \42965_nG2203 , \42966 , \42967 , \42968 , \42969_nG1fb0 , \42970 ,
         \42971 , \42972_nG206f , \42973 , \42974 , \42975 , \42976_nG1e2d , \42977 , \42978 , \42979_nG1ee9 , \42980 ,
         \42981 , \42982 , \42983_nG1cb4 , \42984 , \42985 , \42986_nG1d69 , \42987 , \42988 , \42989 , \42990_nG1b45 ,
         \42991 , \42992 , \42993_nG1bf7 , \42994 , \42995 , \42996 , \42997_nG19e0 , \42998 , \42999 , \43000_nG1a8b ,
         \43001 , \43002 , \43003 , \43004_nG1885 , \43005 , \43006 , \43007_nG192d , \43008 , \43009 , \43010 ,
         \43011_nG1734 , \43012 , \43013 , \43014_nG17d5 , \43015 , \43016 , \43017 , \43018_nG15ed , \43019 , \43020 ,
         \43021_nG168b , \43022 , \43023 , \43024 , \43025_nG14b0 , \43026 , \43027 , \43028_nG1547 , \43029 , \43030 ,
         \43031 , \43032_nG137d , \43033 , \43034 , \43035_nG1411 , \43036 , \43037 , \43038 , \43039_nG1254 , \43040 ,
         \43041 , \43042_nG12e1 , \43043 , \43044 , \43045 , \43046_nG1135 , \43047 , \43048 , \43049_nG11bf , \43050 ,
         \43051 , \43052 , \43053_nG1020 , \43054 , \43055 , \43056_nG10a3 , \43057 , \43058 , \43059 , \43060_nGf15 ,
         \43061 , \43062 , \43063_nGf95 , \43064 , \43065 , \43066 , \43067_nGe14 , \43068 , \43069 , \43070_nGe8d ,
         \43071 , \43072 , \43073 , \43074_nGd1d , \43075 , \43076 , \43077_nGd93 , \43078 , \43079 , \43080 ,
         \43081_nGc30 , \43082 , \43083 , \43084_nGc9f , \43085 , \43086 , \43087 , \43088_nGb4d , \43089 , \43090 ,
         \43091_nGbb9 , \43092 , \43093 , \43094 , \43095_nGa74 , \43096 , \43097 , \43098_nGad9 , \43099 , \43100 ,
         \43101 , \43102_nG9a5 , \43103 , \43104 , \43105_nGa07 , \43106 , \43107 , \43108 , \43109_nG8e0 , \43110 ,
         \43111 , \43112_nG93b , \43113 , \43114 , \43115 , \43116_nG825 , \43117 , \43118 , \43119_nG87d , \43120 ,
         \43121 , \43122 , \43123_nG774 , \43124 , \43125 , \43126_nG7c5 , \43127 , \43128 , \43129 , \43130_nG6cd ,
         \43131 , \43132 , \43133_nG71b , \43134 , \43135 , \43136 , \43137_nG630 , \43138 , \43139 , \43140_nG677 ,
         \43141 , \43142 , \43143 , \43144_nG59d , \43145 , \43146 , \43147_nG5e1 , \43148 , \43149 , \43150 ,
         \43151_nG514 , \43152 , \43153 , \43154_nG551 , \43155 , \43156 , \43157 , \43158_nG495 , \43159 , \43160 ,
         \43161_nG4cf , \43162 , \43163 , \43164 , \43165_nG420 , \43166 , \43167 , \43168_nG453 , \43169 , \43170 ,
         \43171 , \43172_nG3b5 , \43173 , \43174 , \43175_nG3e5 , \43176 , \43177 , \43178 , \43179_nG354 , \43180 ,
         \43181 , \43182_nG37d , \43183 , \43184 , \43185 , \43186_nG2fd , \43187 , \43188 , \43189_nG323 , \43190 ,
         \43191 , \43192 , \43193_nG2b0 , \43194 , \43195 , \43196_nG2cf , \43197 , \43198 , \43199 , \43200_nG26d ,
         \43201 , \43202 , \43203_nG289 , \43204 , \43205 , \43206 , \43207_nG234 , \43208 , \43209 , \43210_nG249 ,
         \43211 , \43212 , \43213 , \43214_nG204 , \43215 , \43216 , \43217_nG217 , \43218 , \43219 , \43220 ,
         \43221_nG1e0 , \43222 , \43223 , \43224_nG1ec , \43225 , \43226 , \43227 , \43228_nG189 , \43229 , \43230 ,
         \43231_nG191 , \43232 , \43233 , \43234 , \43235 , \43236 , \43237 , \43238 , \43239 , \43240 ,
         \43241 , \43242 , \43243 , \43244 , \43245 , \43246 , \43247 , \43248 , \43249 , \43250 ,
         \43251 , \43252 , \43253 , \43254 , \43255 , \43256 , \43257 , \43258 , \43259 , \43260 ,
         \43261 , \43262 , \43263 , \43264 , \43265 , \43266 , \43267 , \43268 , \43269 , \43270 ,
         \43271 , \43272 , \43273 , \43274 , \43275 , \43276 , \43277 , \43278 , \43279 , \43280 ,
         \43281 , \43282 , \43283 , \43284 , \43285 , \43286 , \43287 , \43288 , \43289 , \43290 ,
         \43291 , \43292 , \43293 , \43294 , \43295 , \43296 , \43297 , \43298 , \43299 , \43300 ,
         \43301 , \43302 , \43303 , \43304 , \43305 , \43306 , \43307 , \43308 , \43309 , \43310 ,
         \43311 , \43312 , \43313 , \43314 , \43315 , \43316 , \43317 , \43318 , \43319 , \43320 ,
         \43321 , \43322 , \43323 , \43324 , \43325 , \43326 , \43327 , \43328 , \43329 , \43330 ,
         \43331 , \43332 , \43333 , \43334 , \43335 , \43336 , \43337 , \43338 , \43339 , \43340 ,
         \43341 , \43342 , \43343 , \43344 , \43345 , \43346 , \43347 , \43348 , \43349 , \43350 ,
         \43351 , \43352 , \43353 , \43354 , \43355 , \43356 , \43357 , \43358 , \43359 , \43360 ,
         \43361 , \43362 , \43363 , \43364 , \43365 , \43366 , \43367 , \43368 , \43369 , \43370 ,
         \43371 , \43372 , \43373 , \43374 , \43375 , \43376 , \43377 , \43378 , \43379 , \43380 ,
         \43381 , \43382 , \43383 , \43384 , \43385 , \43386 , \43387 , \43388 , \43389 , \43390 ,
         \43391 , \43392 , \43393 , \43394 , \43395 , \43396 , \43397 , \43398 , \43399 , \43400 ,
         \43401 , \43402 , \43403 , \43404 , \43405 , \43406 , \43407 , \43408 , \43409 , \43410 ,
         \43411 , \43412 , \43413 , \43414 , \43415 , \43416 , \43417 , \43418 , \43419 , \43420 ,
         \43421 , \43422 , \43423 , \43424 , \43425 , \43426 , \43427 , \43428 , \43429 , \43430 ,
         \43431 , \43432 , \43433 , \43434 , \43435 , \43436 , \43437 , \43438 , \43439 , \43440 ,
         \43441 , \43442 , \43443 , \43444 , \43445 , \43446 , \43447 , \43448 , \43449 , \43450 ,
         \43451 , \43452 , \43453 , \43454 , \43455 , \43456 , \43457 , \43458 , \43459 , \43460 ,
         \43461 , \43462 , \43463 , \43464 , \43465 , \43466 , \43467 , \43468 , \43469 , \43470 ,
         \43471 , \43472 , \43473 , \43474 , \43475 , \43476 , \43477 , \43478 , \43479 , \43480 ,
         \43481 , \43482 , \43483 , \43484 , \43485 , \43486 , \43487 , \43488 , \43489 , \43490 ,
         \43491 , \43492 , \43493 , \43494 , \43495 , \43496 , \43497 , \43498 , \43499 , \43500 ,
         \43501 , \43502 , \43503 , \43504 , \43505 , \43506 , \43507 , \43508 , \43509 , \43510 ,
         \43511 , \43512 , \43513 , \43514 , \43515 , \43516 , \43517 , \43518 , \43519 , \43520 ,
         \43521 , \43522 , \43523 , \43524 , \43525 , \43526 , \43527 , \43528 , \43529 , \43530 ,
         \43531 , \43532 , \43533 , \43534 , \43535 , \43536 , \43537 , \43538 , \43539 , \43540 ,
         \43541 , \43542 , \43543 , \43544 , \43545 , \43546 , \43547 , \43548 , \43549 , \43550 ,
         \43551 , \43552 , \43553 , \43554 , \43555 , \43556 , \43557 , \43558 , \43559 , \43560 ,
         \43561 , \43562 , \43563 , \43564 , \43565 , \43566 , \43567 , \43568 , \43569 , \43570 ,
         \43571 , \43572 , \43573 , \43574 , \43575 , \43576 , \43577 , \43578 , \43579 , \43580 ,
         \43581 , \43582 , \43583 , \43584 , \43585 , \43586 , \43587 , \43588 , \43589_nGac8b , \43590 ,
         \43591 , \43592 , \43593 , \43594 , \43595 , \43596 , \43597 , \43598 , \43599 , \43600 ,
         \43601 , \43602 , \43603 , \43604 , \43605 , \43606 , \43607 , \43608 , \43609 , \43610 ,
         \43611 , \43612 , \43613 , \43614 , \43615 , \43616 , \43617 , \43618 , \43619 , \43620 ,
         \43621 , \43622 , \43623 , \43624 , \43625 , \43626 , \43627 , \43628 , \43629 , \43630 ,
         \43631 , \43632 , \43633 , \43634 , \43635 , \43636 , \43637 , \43638 , \43639 , \43640 ,
         \43641 , \43642 , \43643 , \43644 , \43645 , \43646 , \43647 , \43648 , \43649 , \43650 ,
         \43651 , \43652 , \43653 , \43654_nGac8c , \43655 , \43656 , \43657 , \43658_nGac15 , \43659_nGac16 , \43660 ,
         \43661 , \43662 , \43663_nGaaff , \43664_nGab00 , \43665 , \43666 , \43667 , \43668_nGa91b , \43669_nGa91c , \43670 ,
         \43671 , \43672 , \43673_nGa7a7 , \43674_nGa7a8 , \43675 , \43676 , \43677 , \43678_nGa043 , \43679_nGa044 , \43680 ,
         \43681 , \43682 , \43683_nG9cd7 , \43684_nG9cd8 , \43685 , \43686 , \43687 , \43688_nG9b99 , \43689_nG9b9a , \43690 ,
         \43691 , \43692 , \43693_nG9903 , \43694_nG9904 , \43695 , \43696 , \43697 , \43698_nG94f3 , \43699_nG94f4 , \43700 ,
         \43701 , \43702 , \43703_nG9381 , \43704_nG9382 , \43705 , \43706 , \43707 , \43708_nG9205 , \43709_nG9206 , \43710 ,
         \43711 , \43712 , \43713_nG907b , \43714_nG907c , \43715 , \43716 , \43717 , \43718_nG8d4f , \43719_nG8d50 , \43720 ,
         \43721 , \43722 , \43723_nG8bad , \43724_nG8bae , \43725 , \43726 , \43727 , \43728_nG89fb , \43729_nG89fc , \43730 ,
         \43731 , \43732 , \43733_nG8677 , \43734_nG8678 , \43735 , \43736 , \43737 , \43738_nG84a7 , \43739_nG84a8 , \43740 ,
         \43741 , \43742 , \43743_nG80e7 , \43744_nG80e8 , \43745 , \43746 , \43747 , \43748_nG7ef5 , \43749_nG7ef6 , \43750 ,
         \43751 , \43752 , \43753_nG7cf9 , \43754_nG7cfa , \43755 , \43756 , \43757 , \43758_nG7af7 , \43759_nG7af8 , \43760 ,
         \43761 , \43762 , \43763_nG72a1 , \43764_nG72a2 , \43765 , \43766 , \43767 , \43768_nG7077 , \43769_nG7078 , \43770 ,
         \43771 , \43772 , \43773_nG6e3d , \43774_nG6e3e , \43775 , \43776 , \43777 , \43778_nG6bff , \43779_nG6c00 , \43780 ,
         \43781 , \43782 , \43783_nG69b1 , \43784_nG69b2 , \43785 , \43786 , \43787 , \43788_nG64f3 , \43789_nG64f4 , \43790 ,
         \43791 , \43792 , \43793_nG600d , \43794_nG600e , \43795 , \43796 , \43797 , \43798_nG5d8d , \43799_nG5d8e , \43800 ,
         \43801 , \43802 , \43803_nG5b0b , \43804_nG5b0c , \43805 , \43806 , \43807 , \43808_nG5887 , \43809_nG5888 , \43810 ,
         \43811 , \43812 , \43813_nG5601 , \43814_nG5602 , \43815 , \43816 , \43817 , \43818_nG50f3 , \43819_nG50f4 , \43820 ,
         \43821 , \43822 , \43823_nG4e7d , \43824_nG4e7e , \43825 , \43826 , \43827 , \43828_nG4c0d , \43829_nG4c0e , \43830 ,
         \43831 , \43832 , \43833_nG49ab , \43834_nG49ac , \43835 , \43836 , \43837 , \43838_nG474f , \43839_nG4750 , \43840 ,
         \43841 , \43842 , \43843_nG4501 , \43844_nG4502 , \43845 , \43846 , \43847 , \43848_nG42b9 , \43849_nG42ba , \43850 ,
         \43851 , \43852 , \43853_nG407f , \43854_nG4080 , \43855 , \43856 , \43857 , \43858_nG3e4b , \43859_nG3e4c , \43860 ,
         \43861 , \43862 , \43863_nG3c25 , \43864_nG3c26 , \43865 , \43866 , \43867 , \43868_nG3a05 , \43869_nG3a06 , \43870 ,
         \43871 , \43872 , \43873_nG37f3 , \43874_nG37f4 , \43875 , \43876 , \43877 , \43878_nG35e7 , \43879_nG35e8 , \43880 ,
         \43881 , \43882 , \43883_nG33e9 , \43884_nG33ea , \43885 , \43886 , \43887 , \43888_nG31f1 , \43889_nG31f2 , \43890 ,
         \43891 , \43892 , \43893_nG3007 , \43894_nG3008 , \43895 , \43896 , \43897 , \43898_nG2e23 , \43899_nG2e24 , \43900 ,
         \43901 , \43902 , \43903_nG2c4d , \43904_nG2c4e , \43905 , \43906 , \43907 , \43908_nG2a77 , \43909_nG2a78 , \43910 ,
         \43911 , \43912 , \43913_nG28b7 , \43914_nG28b8 , \43915 , \43916 , \43917 , \43918_nG26fb , \43919_nG26fc , \43920 ,
         \43921 , \43922 , \43923_nG254d , \43924_nG254e , \43925 , \43926 , \43927 , \43928_nG23a5 , \43929_nG23a6 , \43930 ,
         \43931 , \43932 , \43933_nG220b , \43934_nG220c , \43935 , \43936 , \43937 , \43938_nG2077 , \43939_nG2078 , \43940 ,
         \43941 , \43942 , \43943_nG1ef1 , \43944_nG1ef2 , \43945 , \43946 , \43947 , \43948_nG1d71 , \43949_nG1d72 , \43950 ,
         \43951 , \43952 , \43953_nG1bff , \43954_nG1c00 , \43955 , \43956 , \43957 , \43958_nG1a93 , \43959_nG1a94 , \43960 ,
         \43961 , \43962 , \43963_nG1935 , \43964_nG1936 , \43965 , \43966 , \43967 , \43968_nG17dd , \43969_nG17de , \43970 ,
         \43971 , \43972 , \43973_nG1693 , \43974_nG1694 , \43975 , \43976 , \43977 , \43978_nG154f , \43979_nG1550 , \43980 ,
         \43981 , \43982 , \43983_nG1419 , \43984_nG141a , \43985 , \43986 , \43987 , \43988_nG12e9 , \43989_nG12ea , \43990 ,
         \43991 , \43992 , \43993_nG11c7 , \43994_nG11c8 , \43995 , \43996 , \43997 , \43998_nG10ab , \43999_nG10ac , \44000 ,
         \44001 , \44002 , \44003_nGf9d , \44004_nGf9e , \44005 , \44006 , \44007 , \44008_nGe95 , \44009_nGe96 , \44010 ,
         \44011 , \44012 , \44013_nGd9b , \44014_nGd9c , \44015 , \44016 , \44017 , \44018_nGca7 , \44019_nGca8 , \44020 ,
         \44021 , \44022 , \44023_nGbc1 , \44024_nGbc2 , \44025 , \44026 , \44027 , \44028_nGae1 , \44029_nGae2 , \44030 ,
         \44031 , \44032 , \44033_nGa0f , \44034_nGa10 , \44035 , \44036 , \44037 , \44038_nG943 , \44039_nG944 , \44040 ,
         \44041 , \44042 , \44043_nG885 , \44044_nG886 , \44045 , \44046 , \44047 , \44048_nG7cd , \44049_nG7ce , \44050 ,
         \44051 , \44052 , \44053_nG723 , \44054_nG724 , \44055 , \44056 , \44057 , \44058_nG67f , \44059_nG680 , \44060 ,
         \44061 , \44062 , \44063_nG5e9 , \44064_nG5ea , \44065 , \44066 , \44067 , \44068_nG559 , \44069_nG55a , \44070 ,
         \44071 , \44072 , \44073_nG4d7 , \44074_nG4d8 , \44075 ;
buf \U$labaj4449 ( R_109_95e4d78, \43655 );
buf \U$labaj4450 ( R_10a_95e4e20, \43660 );
buf \U$labaj4451 ( R_10c_95e4f70, \43665 );
buf \U$labaj4452 ( R_10f_95e5168, \43670 );
buf \U$labaj4453 ( R_111_95e52b8, \43675 );
buf \U$labaj4454 ( R_119_95e57f8, \43680 );
buf \U$labaj4455 ( R_11c_95e59f0, \43685 );
buf \U$labaj4456 ( R_11d_95e5a98, \43690 );
buf \U$labaj4457 ( R_11f_95e5be8, \43695 );
buf \U$labaj4458 ( R_122_95e5de0, \43700 );
buf \U$labaj4459 ( R_123_95e5e88, \43705 );
buf \U$labaj4460 ( R_124_95e5f30, \43710 );
buf \U$labaj4461 ( R_125_95e5fd8, \43715 );
buf \U$labaj4462 ( R_127_95e6128, \43720 );
buf \U$labaj4463 ( R_128_95e61d0, \43725 );
buf \U$labaj4464 ( R_129_95e6278, \43730 );
buf \U$labaj4465 ( R_12b_95e63c8, \43735 );
buf \U$labaj4466 ( R_12c_95e6470, \43740 );
buf \U$labaj4467 ( R_12e_95e65c0, \43745 );
buf \U$labaj4468 ( R_12f_95e6668, \43750 );
buf \U$labaj4469 ( R_130_95e6710, \43755 );
buf \U$labaj4470 ( R_131_95e67b8, \43760 );
buf \U$labaj4471 ( R_135_95e6a58, \43765 );
buf \U$labaj4472 ( R_136_95e6b00, \43770 );
buf \U$labaj4473 ( R_137_95e6ba8, \43775 );
buf \U$labaj4474 ( R_138_95e6c50, \43780 );
buf \U$labaj4475 ( R_139_95e6cf8, \43785 );
buf \U$labaj4476 ( R_13b_95e6e48, \43790 );
buf \U$labaj4477 ( R_13d_95e6f98, \43795 );
buf \U$labaj4478 ( R_13e_95e7040, \43800 );
buf \U$labaj4479 ( R_13f_95e70e8, \43805 );
buf \U$labaj4480 ( R_140_95e7190, \43810 );
buf \U$labaj4481 ( R_141_95e7238, \43815 );
buf \U$labaj4482 ( R_143_95e7388, \43820 );
buf \U$labaj4483 ( R_144_95e7430, \43825 );
buf \U$labaj4484 ( R_145_95e74d8, \43830 );
buf \U$labaj4485 ( R_146_95e7580, \43835 );
buf \U$labaj4486 ( R_147_95e7628, \43840 );
buf \U$labaj4487 ( R_148_95e76d0, \43845 );
buf \U$labaj4488 ( R_149_95e7778, \43850 );
buf \U$labaj4489 ( R_14a_95e7820, \43855 );
buf \U$labaj4490 ( R_14b_95e78c8, \43860 );
buf \U$labaj4491 ( R_14c_95e7970, \43865 );
buf \U$labaj4492 ( R_14d_95e7a18, \43870 );
buf \U$labaj4493 ( R_14e_95e7ac0, \43875 );
buf \U$labaj4494 ( R_14f_95e7b68, \43880 );
buf \U$labaj4495 ( R_150_95e7c10, \43885 );
buf \U$labaj4496 ( R_151_95e7cb8, \43890 );
buf \U$labaj4497 ( R_152_95e7d60, \43895 );
buf \U$labaj4498 ( R_153_95e7e08, \43900 );
buf \U$labaj4499 ( R_154_95e7eb0, \43905 );
buf \U$labaj4500 ( R_155_95e7f58, \43910 );
buf \U$labaj4501 ( R_156_95e8000, \43915 );
buf \U$labaj4502 ( R_157_95e80a8, \43920 );
buf \U$labaj4503 ( R_158_95e8150, \43925 );
buf \U$labaj4504 ( R_159_95e81f8, \43930 );
buf \U$labaj4505 ( R_15a_95e82a0, \43935 );
buf \U$labaj4506 ( R_15b_95e8348, \43940 );
buf \U$labaj4507 ( R_15c_95e83f0, \43945 );
buf \U$labaj4508 ( R_15d_95e8498, \43950 );
buf \U$labaj4509 ( R_15e_95e8540, \43955 );
buf \U$labaj4510 ( R_15f_95e85e8, \43960 );
buf \U$labaj4511 ( R_160_95e8690, \43965 );
buf \U$labaj4512 ( R_161_95e8738, \43970 );
buf \U$labaj4513 ( R_162_95e87e0, \43975 );
buf \U$labaj4514 ( R_163_95e8888, \43980 );
buf \U$labaj4515 ( R_164_95e8930, \43985 );
buf \U$labaj4516 ( R_165_95e89d8, \43990 );
buf \U$labaj4517 ( R_166_95e8a80, \43995 );
buf \U$labaj4518 ( R_167_95e8b28, \44000 );
buf \U$labaj4519 ( R_168_95e8bd0, \44005 );
buf \U$labaj4520 ( R_169_95e8c78, \44010 );
buf \U$labaj4521 ( R_16a_95e8d20, \44015 );
buf \U$labaj4522 ( R_16b_95e8dc8, \44020 );
buf \U$labaj4523 ( R_16c_95e8e70, \44025 );
buf \U$labaj4524 ( R_16d_95e8f18, \44030 );
buf \U$labaj4525 ( R_16e_95e8fc0, \44035 );
buf \U$labaj4526 ( R_16f_95e9068, \44040 );
buf \U$labaj4527 ( R_170_95e9110, \44045 );
buf \U$labaj4528 ( R_171_95e91b8, \44050 );
buf \U$labaj4529 ( R_172_95e9260, \44055 );
buf \U$labaj4530 ( R_173_95e9308, \44060 );
buf \U$labaj4531 ( R_174_95e93b0, \44065 );
buf \U$labaj4532 ( R_175_95e9458, \44070 );
buf \U$labaj4533 ( R_176_95e9500, \44075 );
buf \U$1 ( \344 , RIbb2f070_13);
buf \U$2 ( \345 , RIbb2eff8_14);
buf \U$3 ( \346 , RIbb2ef80_15);
and \U$4 ( \347 , \345 , \346 );
not \U$5 ( \348 , \347 );
and \U$6 ( \349 , \344 , \348 );
not \U$7 ( \350 , \349 );
buf \U$8 ( \351 , RIbb2d798_66);
buf \U$9 ( \352 , RIbb2f160_11);
buf \U$10 ( \353 , RIbb2f0e8_12);
xor \U$11 ( \354 , \352 , \353 );
xor \U$12 ( \355 , \353 , \344 );
not \U$13 ( \356 , \355 );
and \U$14 ( \357 , \354 , \356 );
and \U$15 ( \358 , \351 , \357 );
buf \U$16 ( \359 , RIbb2d810_65);
and \U$17 ( \360 , \359 , \355 );
nor \U$18 ( \361 , \358 , \360 );
and \U$19 ( \362 , \353 , \344 );
not \U$20 ( \363 , \362 );
and \U$21 ( \364 , \352 , \363 );
xnor \U$22 ( \365 , \361 , \364 );
and \U$23 ( \366 , \350 , \365 );
buf \U$24 ( \367 , RIbb2d6a8_68);
buf \U$25 ( \368 , RIbb2f250_9);
buf \U$26 ( \369 , RIbb2f1d8_10);
xor \U$27 ( \370 , \368 , \369 );
xor \U$28 ( \371 , \369 , \352 );
not \U$29 ( \372 , \371 );
and \U$30 ( \373 , \370 , \372 );
and \U$31 ( \374 , \367 , \373 );
buf \U$32 ( \375 , RIbb2d720_67);
and \U$33 ( \376 , \375 , \371 );
nor \U$34 ( \377 , \374 , \376 );
and \U$35 ( \378 , \369 , \352 );
not \U$36 ( \379 , \378 );
and \U$37 ( \380 , \368 , \379 );
xnor \U$38 ( \381 , \377 , \380 );
and \U$39 ( \382 , \365 , \381 );
and \U$40 ( \383 , \350 , \381 );
or \U$41 ( \384 , \366 , \382 , \383 );
buf \U$42 ( \385 , RIbb2d5b8_70);
buf \U$43 ( \386 , RIbb2f340_7);
buf \U$44 ( \387 , RIbb2f2c8_8);
xor \U$45 ( \388 , \386 , \387 );
xor \U$46 ( \389 , \387 , \368 );
not \U$47 ( \390 , \389 );
and \U$48 ( \391 , \388 , \390 );
and \U$49 ( \392 , \385 , \391 );
buf \U$50 ( \393 , RIbb2d630_69);
and \U$51 ( \394 , \393 , \389 );
nor \U$52 ( \395 , \392 , \394 );
and \U$53 ( \396 , \387 , \368 );
not \U$54 ( \397 , \396 );
and \U$55 ( \398 , \386 , \397 );
xnor \U$56 ( \399 , \395 , \398 );
buf \U$57 ( \400 , RIbb2d4c8_72);
buf \U$58 ( \401 , RIbb2f430_5);
buf \U$59 ( \402 , RIbb2f3b8_6);
xor \U$60 ( \403 , \401 , \402 );
xor \U$61 ( \404 , \402 , \386 );
not \U$62 ( \405 , \404 );
and \U$63 ( \406 , \403 , \405 );
and \U$64 ( \407 , \400 , \406 );
buf \U$65 ( \408 , RIbb2d540_71);
and \U$66 ( \409 , \408 , \404 );
nor \U$67 ( \410 , \407 , \409 );
and \U$68 ( \411 , \402 , \386 );
not \U$69 ( \412 , \411 );
and \U$70 ( \413 , \401 , \412 );
xnor \U$71 ( \414 , \410 , \413 );
and \U$72 ( \415 , \399 , \414 );
buf \U$73 ( \416 , RIbb2d3d8_74);
buf \U$74 ( \417 , RIbb2f520_3);
buf \U$75 ( \418 , RIbb2f4a8_4);
xor \U$76 ( \419 , \417 , \418 );
xor \U$77 ( \420 , \418 , \401 );
not \U$78 ( \421 , \420 );
and \U$79 ( \422 , \419 , \421 );
and \U$80 ( \423 , \416 , \422 );
buf \U$81 ( \424 , RIbb2d450_73);
and \U$82 ( \425 , \424 , \420 );
nor \U$83 ( \426 , \423 , \425 );
and \U$84 ( \427 , \418 , \401 );
not \U$85 ( \428 , \427 );
and \U$86 ( \429 , \417 , \428 );
xnor \U$87 ( \430 , \426 , \429 );
and \U$88 ( \431 , \414 , \430 );
and \U$89 ( \432 , \399 , \430 );
or \U$90 ( \433 , \415 , \431 , \432 );
and \U$91 ( \434 , \384 , \433 );
buf \U$92 ( \435 , RIbb2d2e8_76);
buf \U$93 ( \436 , RIbb2f610_1);
buf \U$94 ( \437 , RIbb2f598_2);
xor \U$95 ( \438 , \436 , \437 );
xor \U$96 ( \439 , \437 , \417 );
not \U$97 ( \440 , \439 );
and \U$98 ( \441 , \438 , \440 );
and \U$99 ( \442 , \435 , \441 );
buf \U$100 ( \443 , RIbb2d360_75);
and \U$101 ( \444 , \443 , \439 );
nor \U$102 ( \445 , \442 , \444 );
and \U$103 ( \446 , \437 , \417 );
not \U$104 ( \447 , \446 );
and \U$105 ( \448 , \436 , \447 );
xnor \U$106 ( \449 , \445 , \448 );
buf \U$107 ( \450 , RIbb2d270_77);
and \U$108 ( \451 , \450 , \436 );
and \U$109 ( \452 , \449 , \451 );
and \U$110 ( \453 , \433 , \452 );
and \U$111 ( \454 , \384 , \452 );
or \U$112 ( \455 , \434 , \453 , \454 );
and \U$113 ( \456 , \408 , \406 );
and \U$114 ( \457 , \385 , \404 );
nor \U$115 ( \458 , \456 , \457 );
xnor \U$116 ( \459 , \458 , \413 );
and \U$117 ( \460 , \424 , \422 );
and \U$118 ( \461 , \400 , \420 );
nor \U$119 ( \462 , \460 , \461 );
xnor \U$120 ( \463 , \462 , \429 );
xor \U$121 ( \464 , \459 , \463 );
and \U$122 ( \465 , \443 , \441 );
and \U$123 ( \466 , \416 , \439 );
nor \U$124 ( \467 , \465 , \466 );
xnor \U$125 ( \468 , \467 , \448 );
xor \U$126 ( \469 , \464 , \468 );
and \U$127 ( \470 , \359 , \357 );
not \U$128 ( \471 , \470 );
xnor \U$129 ( \472 , \471 , \364 );
and \U$130 ( \473 , \375 , \373 );
and \U$131 ( \474 , \351 , \371 );
nor \U$132 ( \475 , \473 , \474 );
xnor \U$133 ( \476 , \475 , \380 );
xor \U$134 ( \477 , \472 , \476 );
and \U$135 ( \478 , \393 , \391 );
and \U$136 ( \479 , \367 , \389 );
nor \U$137 ( \480 , \478 , \479 );
xnor \U$138 ( \481 , \480 , \398 );
xor \U$139 ( \482 , \477 , \481 );
and \U$140 ( \483 , \469 , \482 );
and \U$141 ( \484 , \435 , \436 );
not \U$142 ( \485 , \484 );
and \U$143 ( \486 , \482 , \485 );
and \U$144 ( \487 , \469 , \485 );
or \U$145 ( \488 , \483 , \486 , \487 );
and \U$146 ( \489 , \455 , \488 );
and \U$147 ( \490 , \443 , \436 );
and \U$148 ( \491 , \385 , \406 );
and \U$149 ( \492 , \393 , \404 );
nor \U$150 ( \493 , \491 , \492 );
xnor \U$151 ( \494 , \493 , \413 );
and \U$152 ( \495 , \400 , \422 );
and \U$153 ( \496 , \408 , \420 );
nor \U$154 ( \497 , \495 , \496 );
xnor \U$155 ( \498 , \497 , \429 );
xor \U$156 ( \499 , \494 , \498 );
and \U$157 ( \500 , \416 , \441 );
and \U$158 ( \501 , \424 , \439 );
nor \U$159 ( \502 , \500 , \501 );
xnor \U$160 ( \503 , \502 , \448 );
xor \U$161 ( \504 , \499 , \503 );
xor \U$162 ( \505 , \490 , \504 );
not \U$163 ( \506 , \364 );
and \U$164 ( \507 , \351 , \373 );
and \U$165 ( \508 , \359 , \371 );
nor \U$166 ( \509 , \507 , \508 );
xnor \U$167 ( \510 , \509 , \380 );
xor \U$168 ( \511 , \506 , \510 );
and \U$169 ( \512 , \367 , \391 );
and \U$170 ( \513 , \375 , \389 );
nor \U$171 ( \514 , \512 , \513 );
xnor \U$172 ( \515 , \514 , \398 );
xor \U$173 ( \516 , \511 , \515 );
xor \U$174 ( \517 , \505 , \516 );
and \U$175 ( \518 , \488 , \517 );
and \U$176 ( \519 , \455 , \517 );
or \U$177 ( \520 , \489 , \518 , \519 );
and \U$178 ( \521 , \459 , \463 );
and \U$179 ( \522 , \463 , \468 );
and \U$180 ( \523 , \459 , \468 );
or \U$181 ( \524 , \521 , \522 , \523 );
and \U$182 ( \525 , \472 , \476 );
and \U$183 ( \526 , \476 , \481 );
and \U$184 ( \527 , \472 , \481 );
or \U$185 ( \528 , \525 , \526 , \527 );
and \U$186 ( \529 , \524 , \528 );
buf \U$187 ( \530 , \484 );
and \U$188 ( \531 , \528 , \530 );
and \U$189 ( \532 , \524 , \530 );
or \U$190 ( \533 , \529 , \531 , \532 );
and \U$191 ( \534 , \490 , \504 );
and \U$192 ( \535 , \504 , \516 );
and \U$193 ( \536 , \490 , \516 );
or \U$194 ( \537 , \534 , \535 , \536 );
xor \U$195 ( \538 , \533 , \537 );
and \U$196 ( \539 , \408 , \422 );
and \U$197 ( \540 , \385 , \420 );
nor \U$198 ( \541 , \539 , \540 );
xnor \U$199 ( \542 , \541 , \429 );
and \U$200 ( \543 , \424 , \441 );
and \U$201 ( \544 , \400 , \439 );
nor \U$202 ( \545 , \543 , \544 );
xnor \U$203 ( \546 , \545 , \448 );
xor \U$204 ( \547 , \542 , \546 );
and \U$205 ( \548 , \416 , \436 );
xor \U$206 ( \549 , \547 , \548 );
xor \U$207 ( \550 , \538 , \549 );
and \U$208 ( \551 , \520 , \550 );
and \U$209 ( \552 , \359 , \373 );
not \U$210 ( \553 , \552 );
xnor \U$211 ( \554 , \553 , \380 );
and \U$212 ( \555 , \375 , \391 );
and \U$213 ( \556 , \351 , \389 );
nor \U$214 ( \557 , \555 , \556 );
xnor \U$215 ( \558 , \557 , \398 );
xor \U$216 ( \559 , \554 , \558 );
and \U$217 ( \560 , \393 , \406 );
and \U$218 ( \561 , \367 , \404 );
nor \U$219 ( \562 , \560 , \561 );
xnor \U$220 ( \563 , \562 , \413 );
xor \U$221 ( \564 , \559 , \563 );
and \U$222 ( \565 , \494 , \498 );
and \U$223 ( \566 , \498 , \503 );
and \U$224 ( \567 , \494 , \503 );
or \U$225 ( \568 , \565 , \566 , \567 );
and \U$226 ( \569 , \506 , \510 );
and \U$227 ( \570 , \510 , \515 );
and \U$228 ( \571 , \506 , \515 );
or \U$229 ( \572 , \569 , \570 , \571 );
xnor \U$230 ( \573 , \568 , \572 );
xor \U$231 ( \574 , \564 , \573 );
and \U$232 ( \575 , \550 , \574 );
and \U$233 ( \576 , \520 , \574 );
or \U$234 ( \577 , \551 , \575 , \576 );
and \U$235 ( \578 , \533 , \537 );
and \U$236 ( \579 , \537 , \549 );
and \U$237 ( \580 , \533 , \549 );
or \U$238 ( \581 , \578 , \579 , \580 );
and \U$239 ( \582 , \564 , \573 );
xor \U$240 ( \583 , \581 , \582 );
or \U$241 ( \584 , \568 , \572 );
not \U$242 ( \585 , \380 );
and \U$243 ( \586 , \351 , \391 );
and \U$244 ( \587 , \359 , \389 );
nor \U$245 ( \588 , \586 , \587 );
xnor \U$246 ( \589 , \588 , \398 );
xor \U$247 ( \590 , \585 , \589 );
and \U$248 ( \591 , \367 , \406 );
and \U$249 ( \592 , \375 , \404 );
nor \U$250 ( \593 , \591 , \592 );
xnor \U$251 ( \594 , \593 , \413 );
xor \U$252 ( \595 , \590 , \594 );
xor \U$253 ( \596 , \584 , \595 );
and \U$254 ( \597 , \554 , \558 );
and \U$255 ( \598 , \558 , \563 );
and \U$256 ( \599 , \554 , \563 );
or \U$257 ( \600 , \597 , \598 , \599 );
and \U$258 ( \601 , \542 , \546 );
and \U$259 ( \602 , \546 , \548 );
and \U$260 ( \603 , \542 , \548 );
or \U$261 ( \604 , \601 , \602 , \603 );
xor \U$262 ( \605 , \600 , \604 );
and \U$263 ( \606 , \385 , \422 );
and \U$264 ( \607 , \393 , \420 );
nor \U$265 ( \608 , \606 , \607 );
xnor \U$266 ( \609 , \608 , \429 );
and \U$267 ( \610 , \400 , \441 );
and \U$268 ( \611 , \408 , \439 );
nor \U$269 ( \612 , \610 , \611 );
xnor \U$270 ( \613 , \612 , \448 );
xor \U$271 ( \614 , \609 , \613 );
and \U$272 ( \615 , \424 , \436 );
xor \U$273 ( \616 , \614 , \615 );
xor \U$274 ( \617 , \605 , \616 );
xor \U$275 ( \618 , \596 , \617 );
xor \U$276 ( \619 , \583 , \618 );
xor \U$277 ( \620 , \577 , \619 );
xor \U$278 ( \621 , \344 , \345 );
xor \U$279 ( \622 , \345 , \346 );
not \U$280 ( \623 , \622 );
and \U$281 ( \624 , \621 , \623 );
and \U$282 ( \625 , \359 , \624 );
not \U$283 ( \626 , \625 );
xnor \U$284 ( \627 , \626 , \349 );
and \U$285 ( \628 , \375 , \357 );
and \U$286 ( \629 , \351 , \355 );
nor \U$287 ( \630 , \628 , \629 );
xnor \U$288 ( \631 , \630 , \364 );
and \U$289 ( \632 , \627 , \631 );
and \U$290 ( \633 , \393 , \373 );
and \U$291 ( \634 , \367 , \371 );
nor \U$292 ( \635 , \633 , \634 );
xnor \U$293 ( \636 , \635 , \380 );
and \U$294 ( \637 , \631 , \636 );
and \U$295 ( \638 , \627 , \636 );
or \U$296 ( \639 , \632 , \637 , \638 );
and \U$297 ( \640 , \408 , \391 );
and \U$298 ( \641 , \385 , \389 );
nor \U$299 ( \642 , \640 , \641 );
xnor \U$300 ( \643 , \642 , \398 );
and \U$301 ( \644 , \424 , \406 );
and \U$302 ( \645 , \400 , \404 );
nor \U$303 ( \646 , \644 , \645 );
xnor \U$304 ( \647 , \646 , \413 );
and \U$305 ( \648 , \643 , \647 );
and \U$306 ( \649 , \443 , \422 );
and \U$307 ( \650 , \416 , \420 );
nor \U$308 ( \651 , \649 , \650 );
xnor \U$309 ( \652 , \651 , \429 );
and \U$310 ( \653 , \647 , \652 );
and \U$311 ( \654 , \643 , \652 );
or \U$312 ( \655 , \648 , \653 , \654 );
and \U$313 ( \656 , \639 , \655 );
and \U$314 ( \657 , \450 , \441 );
and \U$315 ( \658 , \435 , \439 );
nor \U$316 ( \659 , \657 , \658 );
xnor \U$317 ( \660 , \659 , \448 );
buf \U$318 ( \661 , RIbb2d1f8_78);
and \U$319 ( \662 , \661 , \436 );
or \U$320 ( \663 , \660 , \662 );
and \U$321 ( \664 , \655 , \663 );
and \U$322 ( \665 , \639 , \663 );
or \U$323 ( \666 , \656 , \664 , \665 );
xor \U$324 ( \667 , \350 , \365 );
xor \U$325 ( \668 , \667 , \381 );
xor \U$326 ( \669 , \399 , \414 );
xor \U$327 ( \670 , \669 , \430 );
and \U$328 ( \671 , \668 , \670 );
xor \U$329 ( \672 , \449 , \451 );
and \U$330 ( \673 , \670 , \672 );
and \U$331 ( \674 , \668 , \672 );
or \U$332 ( \675 , \671 , \673 , \674 );
and \U$333 ( \676 , \666 , \675 );
xor \U$334 ( \677 , \469 , \482 );
xor \U$335 ( \678 , \677 , \485 );
and \U$336 ( \679 , \675 , \678 );
and \U$337 ( \680 , \666 , \678 );
or \U$338 ( \681 , \676 , \679 , \680 );
xor \U$339 ( \682 , \524 , \528 );
xor \U$340 ( \683 , \682 , \530 );
and \U$341 ( \684 , \681 , \683 );
xor \U$342 ( \685 , \455 , \488 );
xor \U$343 ( \686 , \685 , \517 );
and \U$344 ( \687 , \683 , \686 );
and \U$345 ( \688 , \681 , \686 );
or \U$346 ( \689 , \684 , \687 , \688 );
xor \U$347 ( \690 , \520 , \550 );
xor \U$348 ( \691 , \690 , \574 );
and \U$349 ( \692 , \689 , \691 );
xor \U$350 ( \693 , \620 , \692 );
xor \U$351 ( \694 , \689 , \691 );
buf \U$352 ( \695 , RIbb2ef08_16);
buf \U$353 ( \696 , RIbb2ee90_17);
and \U$354 ( \697 , \695 , \696 );
not \U$355 ( \698 , \697 );
and \U$356 ( \699 , \346 , \698 );
not \U$357 ( \700 , \699 );
and \U$358 ( \701 , \351 , \624 );
and \U$359 ( \702 , \359 , \622 );
nor \U$360 ( \703 , \701 , \702 );
xnor \U$361 ( \704 , \703 , \349 );
and \U$362 ( \705 , \700 , \704 );
and \U$363 ( \706 , \367 , \357 );
and \U$364 ( \707 , \375 , \355 );
nor \U$365 ( \708 , \706 , \707 );
xnor \U$366 ( \709 , \708 , \364 );
and \U$367 ( \710 , \704 , \709 );
and \U$368 ( \711 , \700 , \709 );
or \U$369 ( \712 , \705 , \710 , \711 );
and \U$370 ( \713 , \435 , \422 );
and \U$371 ( \714 , \443 , \420 );
nor \U$372 ( \715 , \713 , \714 );
xnor \U$373 ( \716 , \715 , \429 );
and \U$374 ( \717 , \661 , \441 );
and \U$375 ( \718 , \450 , \439 );
nor \U$376 ( \719 , \717 , \718 );
xnor \U$377 ( \720 , \719 , \448 );
and \U$378 ( \721 , \716 , \720 );
buf \U$379 ( \722 , RIbb2d180_79);
and \U$380 ( \723 , \722 , \436 );
and \U$381 ( \724 , \720 , \723 );
and \U$382 ( \725 , \716 , \723 );
or \U$383 ( \726 , \721 , \724 , \725 );
and \U$384 ( \727 , \712 , \726 );
and \U$385 ( \728 , \385 , \373 );
and \U$386 ( \729 , \393 , \371 );
nor \U$387 ( \730 , \728 , \729 );
xnor \U$388 ( \731 , \730 , \380 );
and \U$389 ( \732 , \400 , \391 );
and \U$390 ( \733 , \408 , \389 );
nor \U$391 ( \734 , \732 , \733 );
xnor \U$392 ( \735 , \734 , \398 );
and \U$393 ( \736 , \731 , \735 );
and \U$394 ( \737 , \416 , \406 );
and \U$395 ( \738 , \424 , \404 );
nor \U$396 ( \739 , \737 , \738 );
xnor \U$397 ( \740 , \739 , \413 );
and \U$398 ( \741 , \735 , \740 );
and \U$399 ( \742 , \731 , \740 );
or \U$400 ( \743 , \736 , \741 , \742 );
and \U$401 ( \744 , \726 , \743 );
and \U$402 ( \745 , \712 , \743 );
or \U$403 ( \746 , \727 , \744 , \745 );
xor \U$404 ( \747 , \627 , \631 );
xor \U$405 ( \748 , \747 , \636 );
xor \U$406 ( \749 , \643 , \647 );
xor \U$407 ( \750 , \749 , \652 );
and \U$408 ( \751 , \748 , \750 );
xnor \U$409 ( \752 , \660 , \662 );
and \U$410 ( \753 , \750 , \752 );
and \U$411 ( \754 , \748 , \752 );
or \U$412 ( \755 , \751 , \753 , \754 );
and \U$413 ( \756 , \746 , \755 );
xor \U$414 ( \757 , \668 , \670 );
xor \U$415 ( \758 , \757 , \672 );
and \U$416 ( \759 , \755 , \758 );
and \U$417 ( \760 , \746 , \758 );
or \U$418 ( \761 , \756 , \759 , \760 );
xor \U$419 ( \762 , \384 , \433 );
xor \U$420 ( \763 , \762 , \452 );
and \U$421 ( \764 , \761 , \763 );
xor \U$422 ( \765 , \666 , \675 );
xor \U$423 ( \766 , \765 , \678 );
and \U$424 ( \767 , \763 , \766 );
and \U$425 ( \768 , \761 , \766 );
or \U$426 ( \769 , \764 , \767 , \768 );
xor \U$427 ( \770 , \681 , \683 );
xor \U$428 ( \771 , \770 , \686 );
and \U$429 ( \772 , \769 , \771 );
and \U$430 ( \773 , \694 , \772 );
xor \U$431 ( \774 , \694 , \772 );
xor \U$432 ( \775 , \769 , \771 );
and \U$433 ( \776 , \450 , \422 );
and \U$434 ( \777 , \435 , \420 );
nor \U$435 ( \778 , \776 , \777 );
xnor \U$436 ( \779 , \778 , \429 );
and \U$437 ( \780 , \722 , \441 );
and \U$438 ( \781 , \661 , \439 );
nor \U$439 ( \782 , \780 , \781 );
xnor \U$440 ( \783 , \782 , \448 );
and \U$441 ( \784 , \779 , \783 );
buf \U$442 ( \785 , RIbb2d108_80);
and \U$443 ( \786 , \785 , \436 );
and \U$444 ( \787 , \783 , \786 );
and \U$445 ( \788 , \779 , \786 );
or \U$446 ( \789 , \784 , \787 , \788 );
xor \U$447 ( \790 , \346 , \695 );
xor \U$448 ( \791 , \695 , \696 );
not \U$449 ( \792 , \791 );
and \U$450 ( \793 , \790 , \792 );
and \U$451 ( \794 , \359 , \793 );
not \U$452 ( \795 , \794 );
xnor \U$453 ( \796 , \795 , \699 );
and \U$454 ( \797 , \375 , \624 );
and \U$455 ( \798 , \351 , \622 );
nor \U$456 ( \799 , \797 , \798 );
xnor \U$457 ( \800 , \799 , \349 );
and \U$458 ( \801 , \796 , \800 );
and \U$459 ( \802 , \393 , \357 );
and \U$460 ( \803 , \367 , \355 );
nor \U$461 ( \804 , \802 , \803 );
xnor \U$462 ( \805 , \804 , \364 );
and \U$463 ( \806 , \800 , \805 );
and \U$464 ( \807 , \796 , \805 );
or \U$465 ( \808 , \801 , \806 , \807 );
and \U$466 ( \809 , \789 , \808 );
and \U$467 ( \810 , \408 , \373 );
and \U$468 ( \811 , \385 , \371 );
nor \U$469 ( \812 , \810 , \811 );
xnor \U$470 ( \813 , \812 , \380 );
and \U$471 ( \814 , \424 , \391 );
and \U$472 ( \815 , \400 , \389 );
nor \U$473 ( \816 , \814 , \815 );
xnor \U$474 ( \817 , \816 , \398 );
and \U$475 ( \818 , \813 , \817 );
and \U$476 ( \819 , \443 , \406 );
and \U$477 ( \820 , \416 , \404 );
nor \U$478 ( \821 , \819 , \820 );
xnor \U$479 ( \822 , \821 , \413 );
and \U$480 ( \823 , \817 , \822 );
and \U$481 ( \824 , \813 , \822 );
or \U$482 ( \825 , \818 , \823 , \824 );
and \U$483 ( \826 , \808 , \825 );
and \U$484 ( \827 , \789 , \825 );
or \U$485 ( \828 , \809 , \826 , \827 );
xor \U$486 ( \829 , \700 , \704 );
xor \U$487 ( \830 , \829 , \709 );
xor \U$488 ( \831 , \716 , \720 );
xor \U$489 ( \832 , \831 , \723 );
and \U$490 ( \833 , \830 , \832 );
xor \U$491 ( \834 , \731 , \735 );
xor \U$492 ( \835 , \834 , \740 );
and \U$493 ( \836 , \832 , \835 );
and \U$494 ( \837 , \830 , \835 );
or \U$495 ( \838 , \833 , \836 , \837 );
and \U$496 ( \839 , \828 , \838 );
xor \U$497 ( \840 , \748 , \750 );
xor \U$498 ( \841 , \840 , \752 );
and \U$499 ( \842 , \838 , \841 );
and \U$500 ( \843 , \828 , \841 );
or \U$501 ( \844 , \839 , \842 , \843 );
xor \U$502 ( \845 , \639 , \655 );
xor \U$503 ( \846 , \845 , \663 );
and \U$504 ( \847 , \844 , \846 );
xor \U$505 ( \848 , \746 , \755 );
xor \U$506 ( \849 , \848 , \758 );
and \U$507 ( \850 , \846 , \849 );
and \U$508 ( \851 , \844 , \849 );
or \U$509 ( \852 , \847 , \850 , \851 );
xor \U$510 ( \853 , \761 , \763 );
xor \U$511 ( \854 , \853 , \766 );
and \U$512 ( \855 , \852 , \854 );
and \U$513 ( \856 , \775 , \855 );
xor \U$514 ( \857 , \775 , \855 );
xor \U$515 ( \858 , \852 , \854 );
and \U$516 ( \859 , \385 , \357 );
and \U$517 ( \860 , \393 , \355 );
nor \U$518 ( \861 , \859 , \860 );
xnor \U$519 ( \862 , \861 , \364 );
and \U$520 ( \863 , \400 , \373 );
and \U$521 ( \864 , \408 , \371 );
nor \U$522 ( \865 , \863 , \864 );
xnor \U$523 ( \866 , \865 , \380 );
and \U$524 ( \867 , \862 , \866 );
and \U$525 ( \868 , \416 , \391 );
and \U$526 ( \869 , \424 , \389 );
nor \U$527 ( \870 , \868 , \869 );
xnor \U$528 ( \871 , \870 , \398 );
and \U$529 ( \872 , \866 , \871 );
and \U$530 ( \873 , \862 , \871 );
or \U$531 ( \874 , \867 , \872 , \873 );
buf \U$532 ( \875 , RIbb2ee18_18);
buf \U$533 ( \876 , RIbb2eda0_19);
and \U$534 ( \877 , \875 , \876 );
not \U$535 ( \878 , \877 );
and \U$536 ( \879 , \696 , \878 );
not \U$537 ( \880 , \879 );
and \U$538 ( \881 , \351 , \793 );
and \U$539 ( \882 , \359 , \791 );
nor \U$540 ( \883 , \881 , \882 );
xnor \U$541 ( \884 , \883 , \699 );
and \U$542 ( \885 , \880 , \884 );
and \U$543 ( \886 , \367 , \624 );
and \U$544 ( \887 , \375 , \622 );
nor \U$545 ( \888 , \886 , \887 );
xnor \U$546 ( \889 , \888 , \349 );
and \U$547 ( \890 , \884 , \889 );
and \U$548 ( \891 , \880 , \889 );
or \U$549 ( \892 , \885 , \890 , \891 );
and \U$550 ( \893 , \874 , \892 );
and \U$551 ( \894 , \435 , \406 );
and \U$552 ( \895 , \443 , \404 );
nor \U$553 ( \896 , \894 , \895 );
xnor \U$554 ( \897 , \896 , \413 );
and \U$555 ( \898 , \661 , \422 );
and \U$556 ( \899 , \450 , \420 );
nor \U$557 ( \900 , \898 , \899 );
xnor \U$558 ( \901 , \900 , \429 );
and \U$559 ( \902 , \897 , \901 );
and \U$560 ( \903 , \785 , \441 );
and \U$561 ( \904 , \722 , \439 );
nor \U$562 ( \905 , \903 , \904 );
xnor \U$563 ( \906 , \905 , \448 );
and \U$564 ( \907 , \901 , \906 );
and \U$565 ( \908 , \897 , \906 );
or \U$566 ( \909 , \902 , \907 , \908 );
and \U$567 ( \910 , \892 , \909 );
and \U$568 ( \911 , \874 , \909 );
or \U$569 ( \912 , \893 , \910 , \911 );
xor \U$570 ( \913 , \779 , \783 );
xor \U$571 ( \914 , \913 , \786 );
xor \U$572 ( \915 , \813 , \817 );
xor \U$573 ( \916 , \915 , \822 );
or \U$574 ( \917 , \914 , \916 );
and \U$575 ( \918 , \912 , \917 );
xor \U$576 ( \919 , \830 , \832 );
xor \U$577 ( \920 , \919 , \835 );
and \U$578 ( \921 , \917 , \920 );
and \U$579 ( \922 , \912 , \920 );
or \U$580 ( \923 , \918 , \921 , \922 );
xor \U$581 ( \924 , \712 , \726 );
xor \U$582 ( \925 , \924 , \743 );
and \U$583 ( \926 , \923 , \925 );
xor \U$584 ( \927 , \828 , \838 );
xor \U$585 ( \928 , \927 , \841 );
and \U$586 ( \929 , \925 , \928 );
and \U$587 ( \930 , \923 , \928 );
or \U$588 ( \931 , \926 , \929 , \930 );
xor \U$589 ( \932 , \844 , \846 );
xor \U$590 ( \933 , \932 , \849 );
and \U$591 ( \934 , \931 , \933 );
and \U$592 ( \935 , \858 , \934 );
xor \U$593 ( \936 , \858 , \934 );
xor \U$594 ( \937 , \931 , \933 );
and \U$595 ( \938 , \408 , \357 );
and \U$596 ( \939 , \385 , \355 );
nor \U$597 ( \940 , \938 , \939 );
xnor \U$598 ( \941 , \940 , \364 );
and \U$599 ( \942 , \424 , \373 );
and \U$600 ( \943 , \400 , \371 );
nor \U$601 ( \944 , \942 , \943 );
xnor \U$602 ( \945 , \944 , \380 );
and \U$603 ( \946 , \941 , \945 );
and \U$604 ( \947 , \443 , \391 );
and \U$605 ( \948 , \416 , \389 );
nor \U$606 ( \949 , \947 , \948 );
xnor \U$607 ( \950 , \949 , \398 );
and \U$608 ( \951 , \945 , \950 );
and \U$609 ( \952 , \941 , \950 );
or \U$610 ( \953 , \946 , \951 , \952 );
xor \U$611 ( \954 , \696 , \875 );
xor \U$612 ( \955 , \875 , \876 );
not \U$613 ( \956 , \955 );
and \U$614 ( \957 , \954 , \956 );
and \U$615 ( \958 , \359 , \957 );
not \U$616 ( \959 , \958 );
xnor \U$617 ( \960 , \959 , \879 );
and \U$618 ( \961 , \375 , \793 );
and \U$619 ( \962 , \351 , \791 );
nor \U$620 ( \963 , \961 , \962 );
xnor \U$621 ( \964 , \963 , \699 );
and \U$622 ( \965 , \960 , \964 );
and \U$623 ( \966 , \393 , \624 );
and \U$624 ( \967 , \367 , \622 );
nor \U$625 ( \968 , \966 , \967 );
xnor \U$626 ( \969 , \968 , \349 );
and \U$627 ( \970 , \964 , \969 );
and \U$628 ( \971 , \960 , \969 );
or \U$629 ( \972 , \965 , \970 , \971 );
and \U$630 ( \973 , \953 , \972 );
and \U$631 ( \974 , \450 , \406 );
and \U$632 ( \975 , \435 , \404 );
nor \U$633 ( \976 , \974 , \975 );
xnor \U$634 ( \977 , \976 , \413 );
and \U$635 ( \978 , \722 , \422 );
and \U$636 ( \979 , \661 , \420 );
nor \U$637 ( \980 , \978 , \979 );
xnor \U$638 ( \981 , \980 , \429 );
and \U$639 ( \982 , \977 , \981 );
buf \U$640 ( \983 , RIbb2d090_81);
and \U$641 ( \984 , \983 , \441 );
and \U$642 ( \985 , \785 , \439 );
nor \U$643 ( \986 , \984 , \985 );
xnor \U$644 ( \987 , \986 , \448 );
and \U$645 ( \988 , \981 , \987 );
and \U$646 ( \989 , \977 , \987 );
or \U$647 ( \990 , \982 , \988 , \989 );
and \U$648 ( \991 , \972 , \990 );
and \U$649 ( \992 , \953 , \990 );
or \U$650 ( \993 , \973 , \991 , \992 );
and \U$651 ( \994 , \983 , \436 );
xor \U$652 ( \995 , \862 , \866 );
xor \U$653 ( \996 , \995 , \871 );
and \U$654 ( \997 , \994 , \996 );
xor \U$655 ( \998 , \897 , \901 );
xor \U$656 ( \999 , \998 , \906 );
and \U$657 ( \1000 , \996 , \999 );
and \U$658 ( \1001 , \994 , \999 );
or \U$659 ( \1002 , \997 , \1000 , \1001 );
and \U$660 ( \1003 , \993 , \1002 );
xor \U$661 ( \1004 , \796 , \800 );
xor \U$662 ( \1005 , \1004 , \805 );
and \U$663 ( \1006 , \1002 , \1005 );
and \U$664 ( \1007 , \993 , \1005 );
or \U$665 ( \1008 , \1003 , \1006 , \1007 );
xor \U$666 ( \1009 , \789 , \808 );
xor \U$667 ( \1010 , \1009 , \825 );
and \U$668 ( \1011 , \1008 , \1010 );
xor \U$669 ( \1012 , \912 , \917 );
xor \U$670 ( \1013 , \1012 , \920 );
and \U$671 ( \1014 , \1010 , \1013 );
and \U$672 ( \1015 , \1008 , \1013 );
or \U$673 ( \1016 , \1011 , \1014 , \1015 );
buf \U$674 ( \1017 , RIbb2ed28_20);
buf \U$675 ( \1018 , RIbb2ecb0_21);
and \U$676 ( \1019 , \1017 , \1018 );
not \U$677 ( \1020 , \1019 );
and \U$678 ( \1021 , \876 , \1020 );
not \U$679 ( \1022 , \1021 );
and \U$680 ( \1023 , \351 , \957 );
and \U$681 ( \1024 , \359 , \955 );
nor \U$682 ( \1025 , \1023 , \1024 );
xnor \U$683 ( \1026 , \1025 , \879 );
and \U$684 ( \1027 , \1022 , \1026 );
and \U$685 ( \1028 , \367 , \793 );
and \U$686 ( \1029 , \375 , \791 );
nor \U$687 ( \1030 , \1028 , \1029 );
xnor \U$688 ( \1031 , \1030 , \699 );
and \U$689 ( \1032 , \1026 , \1031 );
and \U$690 ( \1033 , \1022 , \1031 );
or \U$691 ( \1034 , \1027 , \1032 , \1033 );
and \U$692 ( \1035 , \385 , \624 );
and \U$693 ( \1036 , \393 , \622 );
nor \U$694 ( \1037 , \1035 , \1036 );
xnor \U$695 ( \1038 , \1037 , \349 );
and \U$696 ( \1039 , \400 , \357 );
and \U$697 ( \1040 , \408 , \355 );
nor \U$698 ( \1041 , \1039 , \1040 );
xnor \U$699 ( \1042 , \1041 , \364 );
and \U$700 ( \1043 , \1038 , \1042 );
and \U$701 ( \1044 , \416 , \373 );
and \U$702 ( \1045 , \424 , \371 );
nor \U$703 ( \1046 , \1044 , \1045 );
xnor \U$704 ( \1047 , \1046 , \380 );
and \U$705 ( \1048 , \1042 , \1047 );
and \U$706 ( \1049 , \1038 , \1047 );
or \U$707 ( \1050 , \1043 , \1048 , \1049 );
and \U$708 ( \1051 , \1034 , \1050 );
and \U$709 ( \1052 , \435 , \391 );
and \U$710 ( \1053 , \443 , \389 );
nor \U$711 ( \1054 , \1052 , \1053 );
xnor \U$712 ( \1055 , \1054 , \398 );
and \U$713 ( \1056 , \661 , \406 );
and \U$714 ( \1057 , \450 , \404 );
nor \U$715 ( \1058 , \1056 , \1057 );
xnor \U$716 ( \1059 , \1058 , \413 );
and \U$717 ( \1060 , \1055 , \1059 );
and \U$718 ( \1061 , \785 , \422 );
and \U$719 ( \1062 , \722 , \420 );
nor \U$720 ( \1063 , \1061 , \1062 );
xnor \U$721 ( \1064 , \1063 , \429 );
and \U$722 ( \1065 , \1059 , \1064 );
and \U$723 ( \1066 , \1055 , \1064 );
or \U$724 ( \1067 , \1060 , \1065 , \1066 );
and \U$725 ( \1068 , \1050 , \1067 );
and \U$726 ( \1069 , \1034 , \1067 );
or \U$727 ( \1070 , \1051 , \1068 , \1069 );
buf \U$728 ( \1071 , RIbb2d018_82);
and \U$729 ( \1072 , \1071 , \436 );
xor \U$730 ( \1073 , \977 , \981 );
xor \U$731 ( \1074 , \1073 , \987 );
or \U$732 ( \1075 , \1072 , \1074 );
and \U$733 ( \1076 , \1070 , \1075 );
xor \U$734 ( \1077 , \941 , \945 );
xor \U$735 ( \1078 , \1077 , \950 );
xor \U$736 ( \1079 , \960 , \964 );
xor \U$737 ( \1080 , \1079 , \969 );
and \U$738 ( \1081 , \1078 , \1080 );
and \U$739 ( \1082 , \1075 , \1081 );
and \U$740 ( \1083 , \1070 , \1081 );
or \U$741 ( \1084 , \1076 , \1082 , \1083 );
xor \U$742 ( \1085 , \880 , \884 );
xor \U$743 ( \1086 , \1085 , \889 );
xor \U$744 ( \1087 , \953 , \972 );
xor \U$745 ( \1088 , \1087 , \990 );
and \U$746 ( \1089 , \1086 , \1088 );
xor \U$747 ( \1090 , \994 , \996 );
xor \U$748 ( \1091 , \1090 , \999 );
and \U$749 ( \1092 , \1088 , \1091 );
and \U$750 ( \1093 , \1086 , \1091 );
or \U$751 ( \1094 , \1089 , \1092 , \1093 );
and \U$752 ( \1095 , \1084 , \1094 );
xnor \U$753 ( \1096 , \914 , \916 );
and \U$754 ( \1097 , \1094 , \1096 );
and \U$755 ( \1098 , \1084 , \1096 );
or \U$756 ( \1099 , \1095 , \1097 , \1098 );
xor \U$757 ( \1100 , \874 , \892 );
xor \U$758 ( \1101 , \1100 , \909 );
xor \U$759 ( \1102 , \993 , \1002 );
xor \U$760 ( \1103 , \1102 , \1005 );
and \U$761 ( \1104 , \1101 , \1103 );
and \U$762 ( \1105 , \1099 , \1104 );
xor \U$763 ( \1106 , \1008 , \1010 );
xor \U$764 ( \1107 , \1106 , \1013 );
and \U$765 ( \1108 , \1104 , \1107 );
and \U$766 ( \1109 , \1099 , \1107 );
or \U$767 ( \1110 , \1105 , \1108 , \1109 );
and \U$768 ( \1111 , \1016 , \1110 );
xor \U$769 ( \1112 , \923 , \925 );
xor \U$770 ( \1113 , \1112 , \928 );
and \U$771 ( \1114 , \1110 , \1113 );
and \U$772 ( \1115 , \1016 , \1113 );
or \U$773 ( \1116 , \1111 , \1114 , \1115 );
and \U$774 ( \1117 , \937 , \1116 );
xor \U$775 ( \1118 , \937 , \1116 );
xor \U$776 ( \1119 , \1016 , \1110 );
xor \U$777 ( \1120 , \1119 , \1113 );
and \U$778 ( \1121 , \450 , \391 );
and \U$779 ( \1122 , \435 , \389 );
nor \U$780 ( \1123 , \1121 , \1122 );
xnor \U$781 ( \1124 , \1123 , \398 );
and \U$782 ( \1125 , \722 , \406 );
and \U$783 ( \1126 , \661 , \404 );
nor \U$784 ( \1127 , \1125 , \1126 );
xnor \U$785 ( \1128 , \1127 , \413 );
and \U$786 ( \1129 , \1124 , \1128 );
and \U$787 ( \1130 , \983 , \422 );
and \U$788 ( \1131 , \785 , \420 );
nor \U$789 ( \1132 , \1130 , \1131 );
xnor \U$790 ( \1133 , \1132 , \429 );
and \U$791 ( \1134 , \1128 , \1133 );
and \U$792 ( \1135 , \1124 , \1133 );
or \U$793 ( \1136 , \1129 , \1134 , \1135 );
and \U$794 ( \1137 , \408 , \624 );
and \U$795 ( \1138 , \385 , \622 );
nor \U$796 ( \1139 , \1137 , \1138 );
xnor \U$797 ( \1140 , \1139 , \349 );
and \U$798 ( \1141 , \424 , \357 );
and \U$799 ( \1142 , \400 , \355 );
nor \U$800 ( \1143 , \1141 , \1142 );
xnor \U$801 ( \1144 , \1143 , \364 );
and \U$802 ( \1145 , \1140 , \1144 );
and \U$803 ( \1146 , \443 , \373 );
and \U$804 ( \1147 , \416 , \371 );
nor \U$805 ( \1148 , \1146 , \1147 );
xnor \U$806 ( \1149 , \1148 , \380 );
and \U$807 ( \1150 , \1144 , \1149 );
and \U$808 ( \1151 , \1140 , \1149 );
or \U$809 ( \1152 , \1145 , \1150 , \1151 );
and \U$810 ( \1153 , \1136 , \1152 );
xor \U$811 ( \1154 , \876 , \1017 );
xor \U$812 ( \1155 , \1017 , \1018 );
not \U$813 ( \1156 , \1155 );
and \U$814 ( \1157 , \1154 , \1156 );
and \U$815 ( \1158 , \359 , \1157 );
not \U$816 ( \1159 , \1158 );
xnor \U$817 ( \1160 , \1159 , \1021 );
and \U$818 ( \1161 , \375 , \957 );
and \U$819 ( \1162 , \351 , \955 );
nor \U$820 ( \1163 , \1161 , \1162 );
xnor \U$821 ( \1164 , \1163 , \879 );
and \U$822 ( \1165 , \1160 , \1164 );
and \U$823 ( \1166 , \393 , \793 );
and \U$824 ( \1167 , \367 , \791 );
nor \U$825 ( \1168 , \1166 , \1167 );
xnor \U$826 ( \1169 , \1168 , \699 );
and \U$827 ( \1170 , \1164 , \1169 );
and \U$828 ( \1171 , \1160 , \1169 );
or \U$829 ( \1172 , \1165 , \1170 , \1171 );
and \U$830 ( \1173 , \1152 , \1172 );
and \U$831 ( \1174 , \1136 , \1172 );
or \U$832 ( \1175 , \1153 , \1173 , \1174 );
buf \U$833 ( \1176 , RIbb2cfa0_83);
and \U$834 ( \1177 , \1176 , \441 );
and \U$835 ( \1178 , \1071 , \439 );
nor \U$836 ( \1179 , \1177 , \1178 );
xnor \U$837 ( \1180 , \1179 , \448 );
buf \U$838 ( \1181 , RIbb2cf28_84);
and \U$839 ( \1182 , \1181 , \436 );
or \U$840 ( \1183 , \1180 , \1182 );
and \U$841 ( \1184 , \1071 , \441 );
and \U$842 ( \1185 , \983 , \439 );
nor \U$843 ( \1186 , \1184 , \1185 );
xnor \U$844 ( \1187 , \1186 , \448 );
and \U$845 ( \1188 , \1183 , \1187 );
and \U$846 ( \1189 , \1176 , \436 );
and \U$847 ( \1190 , \1187 , \1189 );
and \U$848 ( \1191 , \1183 , \1189 );
or \U$849 ( \1192 , \1188 , \1190 , \1191 );
and \U$850 ( \1193 , \1175 , \1192 );
xor \U$851 ( \1194 , \1022 , \1026 );
xor \U$852 ( \1195 , \1194 , \1031 );
xor \U$853 ( \1196 , \1038 , \1042 );
xor \U$854 ( \1197 , \1196 , \1047 );
and \U$855 ( \1198 , \1195 , \1197 );
xor \U$856 ( \1199 , \1055 , \1059 );
xor \U$857 ( \1200 , \1199 , \1064 );
and \U$858 ( \1201 , \1197 , \1200 );
and \U$859 ( \1202 , \1195 , \1200 );
or \U$860 ( \1203 , \1198 , \1201 , \1202 );
and \U$861 ( \1204 , \1192 , \1203 );
and \U$862 ( \1205 , \1175 , \1203 );
or \U$863 ( \1206 , \1193 , \1204 , \1205 );
xor \U$864 ( \1207 , \1034 , \1050 );
xor \U$865 ( \1208 , \1207 , \1067 );
xnor \U$866 ( \1209 , \1072 , \1074 );
and \U$867 ( \1210 , \1208 , \1209 );
xor \U$868 ( \1211 , \1078 , \1080 );
and \U$869 ( \1212 , \1209 , \1211 );
and \U$870 ( \1213 , \1208 , \1211 );
or \U$871 ( \1214 , \1210 , \1212 , \1213 );
and \U$872 ( \1215 , \1206 , \1214 );
xor \U$873 ( \1216 , \1086 , \1088 );
xor \U$874 ( \1217 , \1216 , \1091 );
and \U$875 ( \1218 , \1214 , \1217 );
and \U$876 ( \1219 , \1206 , \1217 );
or \U$877 ( \1220 , \1215 , \1218 , \1219 );
xor \U$878 ( \1221 , \1084 , \1094 );
xor \U$879 ( \1222 , \1221 , \1096 );
and \U$880 ( \1223 , \1220 , \1222 );
xor \U$881 ( \1224 , \1101 , \1103 );
and \U$882 ( \1225 , \1222 , \1224 );
and \U$883 ( \1226 , \1220 , \1224 );
or \U$884 ( \1227 , \1223 , \1225 , \1226 );
xor \U$885 ( \1228 , \1099 , \1104 );
xor \U$886 ( \1229 , \1228 , \1107 );
and \U$887 ( \1230 , \1227 , \1229 );
and \U$888 ( \1231 , \1120 , \1230 );
xor \U$889 ( \1232 , \1120 , \1230 );
xor \U$890 ( \1233 , \1227 , \1229 );
buf \U$891 ( \1234 , RIbb2ec38_22);
buf \U$892 ( \1235 , RIbb2ebc0_23);
and \U$893 ( \1236 , \1234 , \1235 );
not \U$894 ( \1237 , \1236 );
and \U$895 ( \1238 , \1018 , \1237 );
not \U$896 ( \1239 , \1238 );
and \U$897 ( \1240 , \351 , \1157 );
and \U$898 ( \1241 , \359 , \1155 );
nor \U$899 ( \1242 , \1240 , \1241 );
xnor \U$900 ( \1243 , \1242 , \1021 );
and \U$901 ( \1244 , \1239 , \1243 );
and \U$902 ( \1245 , \367 , \957 );
and \U$903 ( \1246 , \375 , \955 );
nor \U$904 ( \1247 , \1245 , \1246 );
xnor \U$905 ( \1248 , \1247 , \879 );
and \U$906 ( \1249 , \1243 , \1248 );
and \U$907 ( \1250 , \1239 , \1248 );
or \U$908 ( \1251 , \1244 , \1249 , \1250 );
and \U$909 ( \1252 , \435 , \373 );
and \U$910 ( \1253 , \443 , \371 );
nor \U$911 ( \1254 , \1252 , \1253 );
xnor \U$912 ( \1255 , \1254 , \380 );
and \U$913 ( \1256 , \661 , \391 );
and \U$914 ( \1257 , \450 , \389 );
nor \U$915 ( \1258 , \1256 , \1257 );
xnor \U$916 ( \1259 , \1258 , \398 );
and \U$917 ( \1260 , \1255 , \1259 );
and \U$918 ( \1261 , \785 , \406 );
and \U$919 ( \1262 , \722 , \404 );
nor \U$920 ( \1263 , \1261 , \1262 );
xnor \U$921 ( \1264 , \1263 , \413 );
and \U$922 ( \1265 , \1259 , \1264 );
and \U$923 ( \1266 , \1255 , \1264 );
or \U$924 ( \1267 , \1260 , \1265 , \1266 );
and \U$925 ( \1268 , \1251 , \1267 );
and \U$926 ( \1269 , \385 , \793 );
and \U$927 ( \1270 , \393 , \791 );
nor \U$928 ( \1271 , \1269 , \1270 );
xnor \U$929 ( \1272 , \1271 , \699 );
and \U$930 ( \1273 , \400 , \624 );
and \U$931 ( \1274 , \408 , \622 );
nor \U$932 ( \1275 , \1273 , \1274 );
xnor \U$933 ( \1276 , \1275 , \349 );
and \U$934 ( \1277 , \1272 , \1276 );
and \U$935 ( \1278 , \416 , \357 );
and \U$936 ( \1279 , \424 , \355 );
nor \U$937 ( \1280 , \1278 , \1279 );
xnor \U$938 ( \1281 , \1280 , \364 );
and \U$939 ( \1282 , \1276 , \1281 );
and \U$940 ( \1283 , \1272 , \1281 );
or \U$941 ( \1284 , \1277 , \1282 , \1283 );
and \U$942 ( \1285 , \1267 , \1284 );
and \U$943 ( \1286 , \1251 , \1284 );
or \U$944 ( \1287 , \1268 , \1285 , \1286 );
and \U$945 ( \1288 , \1071 , \422 );
and \U$946 ( \1289 , \983 , \420 );
nor \U$947 ( \1290 , \1288 , \1289 );
xnor \U$948 ( \1291 , \1290 , \429 );
and \U$949 ( \1292 , \1181 , \441 );
and \U$950 ( \1293 , \1176 , \439 );
nor \U$951 ( \1294 , \1292 , \1293 );
xnor \U$952 ( \1295 , \1294 , \448 );
and \U$953 ( \1296 , \1291 , \1295 );
buf \U$954 ( \1297 , RIbb2ceb0_85);
and \U$955 ( \1298 , \1297 , \436 );
and \U$956 ( \1299 , \1295 , \1298 );
and \U$957 ( \1300 , \1291 , \1298 );
or \U$958 ( \1301 , \1296 , \1299 , \1300 );
xor \U$959 ( \1302 , \1124 , \1128 );
xor \U$960 ( \1303 , \1302 , \1133 );
and \U$961 ( \1304 , \1301 , \1303 );
xnor \U$962 ( \1305 , \1180 , \1182 );
and \U$963 ( \1306 , \1303 , \1305 );
and \U$964 ( \1307 , \1301 , \1305 );
or \U$965 ( \1308 , \1304 , \1306 , \1307 );
and \U$966 ( \1309 , \1287 , \1308 );
xor \U$967 ( \1310 , \1140 , \1144 );
xor \U$968 ( \1311 , \1310 , \1149 );
xor \U$969 ( \1312 , \1160 , \1164 );
xor \U$970 ( \1313 , \1312 , \1169 );
and \U$971 ( \1314 , \1311 , \1313 );
and \U$972 ( \1315 , \1308 , \1314 );
and \U$973 ( \1316 , \1287 , \1314 );
or \U$974 ( \1317 , \1309 , \1315 , \1316 );
xor \U$975 ( \1318 , \1136 , \1152 );
xor \U$976 ( \1319 , \1318 , \1172 );
xor \U$977 ( \1320 , \1183 , \1187 );
xor \U$978 ( \1321 , \1320 , \1189 );
and \U$979 ( \1322 , \1319 , \1321 );
xor \U$980 ( \1323 , \1195 , \1197 );
xor \U$981 ( \1324 , \1323 , \1200 );
and \U$982 ( \1325 , \1321 , \1324 );
and \U$983 ( \1326 , \1319 , \1324 );
or \U$984 ( \1327 , \1322 , \1325 , \1326 );
and \U$985 ( \1328 , \1317 , \1327 );
xor \U$986 ( \1329 , \1208 , \1209 );
xor \U$987 ( \1330 , \1329 , \1211 );
and \U$988 ( \1331 , \1327 , \1330 );
and \U$989 ( \1332 , \1317 , \1330 );
or \U$990 ( \1333 , \1328 , \1331 , \1332 );
xor \U$991 ( \1334 , \1070 , \1075 );
xor \U$992 ( \1335 , \1334 , \1081 );
and \U$993 ( \1336 , \1333 , \1335 );
xor \U$994 ( \1337 , \1206 , \1214 );
xor \U$995 ( \1338 , \1337 , \1217 );
and \U$996 ( \1339 , \1335 , \1338 );
and \U$997 ( \1340 , \1333 , \1338 );
or \U$998 ( \1341 , \1336 , \1339 , \1340 );
xor \U$999 ( \1342 , \1220 , \1222 );
xor \U$1000 ( \1343 , \1342 , \1224 );
and \U$1001 ( \1344 , \1341 , \1343 );
and \U$1002 ( \1345 , \1233 , \1344 );
xor \U$1003 ( \1346 , \1233 , \1344 );
xor \U$1004 ( \1347 , \1341 , \1343 );
xor \U$1005 ( \1348 , \1018 , \1234 );
xor \U$1006 ( \1349 , \1234 , \1235 );
not \U$1007 ( \1350 , \1349 );
and \U$1008 ( \1351 , \1348 , \1350 );
and \U$1009 ( \1352 , \359 , \1351 );
not \U$1010 ( \1353 , \1352 );
xnor \U$1011 ( \1354 , \1353 , \1238 );
and \U$1012 ( \1355 , \375 , \1157 );
and \U$1013 ( \1356 , \351 , \1155 );
nor \U$1014 ( \1357 , \1355 , \1356 );
xnor \U$1015 ( \1358 , \1357 , \1021 );
and \U$1016 ( \1359 , \1354 , \1358 );
and \U$1017 ( \1360 , \393 , \957 );
and \U$1018 ( \1361 , \367 , \955 );
nor \U$1019 ( \1362 , \1360 , \1361 );
xnor \U$1020 ( \1363 , \1362 , \879 );
and \U$1021 ( \1364 , \1358 , \1363 );
and \U$1022 ( \1365 , \1354 , \1363 );
or \U$1023 ( \1366 , \1359 , \1364 , \1365 );
and \U$1024 ( \1367 , \450 , \373 );
and \U$1025 ( \1368 , \435 , \371 );
nor \U$1026 ( \1369 , \1367 , \1368 );
xnor \U$1027 ( \1370 , \1369 , \380 );
and \U$1028 ( \1371 , \722 , \391 );
and \U$1029 ( \1372 , \661 , \389 );
nor \U$1030 ( \1373 , \1371 , \1372 );
xnor \U$1031 ( \1374 , \1373 , \398 );
and \U$1032 ( \1375 , \1370 , \1374 );
and \U$1033 ( \1376 , \983 , \406 );
and \U$1034 ( \1377 , \785 , \404 );
nor \U$1035 ( \1378 , \1376 , \1377 );
xnor \U$1036 ( \1379 , \1378 , \413 );
and \U$1037 ( \1380 , \1374 , \1379 );
and \U$1038 ( \1381 , \1370 , \1379 );
or \U$1039 ( \1382 , \1375 , \1380 , \1381 );
and \U$1040 ( \1383 , \1366 , \1382 );
and \U$1041 ( \1384 , \408 , \793 );
and \U$1042 ( \1385 , \385 , \791 );
nor \U$1043 ( \1386 , \1384 , \1385 );
xnor \U$1044 ( \1387 , \1386 , \699 );
and \U$1045 ( \1388 , \424 , \624 );
and \U$1046 ( \1389 , \400 , \622 );
nor \U$1047 ( \1390 , \1388 , \1389 );
xnor \U$1048 ( \1391 , \1390 , \349 );
and \U$1049 ( \1392 , \1387 , \1391 );
and \U$1050 ( \1393 , \443 , \357 );
and \U$1051 ( \1394 , \416 , \355 );
nor \U$1052 ( \1395 , \1393 , \1394 );
xnor \U$1053 ( \1396 , \1395 , \364 );
and \U$1054 ( \1397 , \1391 , \1396 );
and \U$1055 ( \1398 , \1387 , \1396 );
or \U$1056 ( \1399 , \1392 , \1397 , \1398 );
and \U$1057 ( \1400 , \1382 , \1399 );
and \U$1058 ( \1401 , \1366 , \1399 );
or \U$1059 ( \1402 , \1383 , \1400 , \1401 );
and \U$1060 ( \1403 , \1176 , \422 );
and \U$1061 ( \1404 , \1071 , \420 );
nor \U$1062 ( \1405 , \1403 , \1404 );
xnor \U$1063 ( \1406 , \1405 , \429 );
and \U$1064 ( \1407 , \1297 , \441 );
and \U$1065 ( \1408 , \1181 , \439 );
nor \U$1066 ( \1409 , \1407 , \1408 );
xnor \U$1067 ( \1410 , \1409 , \448 );
and \U$1068 ( \1411 , \1406 , \1410 );
buf \U$1069 ( \1412 , RIbb2ce38_86);
and \U$1070 ( \1413 , \1412 , \436 );
and \U$1071 ( \1414 , \1410 , \1413 );
and \U$1072 ( \1415 , \1406 , \1413 );
or \U$1073 ( \1416 , \1411 , \1414 , \1415 );
xor \U$1074 ( \1417 , \1291 , \1295 );
xor \U$1075 ( \1418 , \1417 , \1298 );
and \U$1076 ( \1419 , \1416 , \1418 );
xor \U$1077 ( \1420 , \1255 , \1259 );
xor \U$1078 ( \1421 , \1420 , \1264 );
and \U$1079 ( \1422 , \1418 , \1421 );
and \U$1080 ( \1423 , \1416 , \1421 );
or \U$1081 ( \1424 , \1419 , \1422 , \1423 );
and \U$1082 ( \1425 , \1402 , \1424 );
xor \U$1083 ( \1426 , \1239 , \1243 );
xor \U$1084 ( \1427 , \1426 , \1248 );
xor \U$1085 ( \1428 , \1272 , \1276 );
xor \U$1086 ( \1429 , \1428 , \1281 );
and \U$1087 ( \1430 , \1427 , \1429 );
and \U$1088 ( \1431 , \1424 , \1430 );
and \U$1089 ( \1432 , \1402 , \1430 );
or \U$1090 ( \1433 , \1425 , \1431 , \1432 );
xor \U$1091 ( \1434 , \1251 , \1267 );
xor \U$1092 ( \1435 , \1434 , \1284 );
xor \U$1093 ( \1436 , \1301 , \1303 );
xor \U$1094 ( \1437 , \1436 , \1305 );
and \U$1095 ( \1438 , \1435 , \1437 );
xor \U$1096 ( \1439 , \1311 , \1313 );
and \U$1097 ( \1440 , \1437 , \1439 );
and \U$1098 ( \1441 , \1435 , \1439 );
or \U$1099 ( \1442 , \1438 , \1440 , \1441 );
and \U$1100 ( \1443 , \1433 , \1442 );
xor \U$1101 ( \1444 , \1319 , \1321 );
xor \U$1102 ( \1445 , \1444 , \1324 );
and \U$1103 ( \1446 , \1442 , \1445 );
and \U$1104 ( \1447 , \1433 , \1445 );
or \U$1105 ( \1448 , \1443 , \1446 , \1447 );
xor \U$1106 ( \1449 , \1175 , \1192 );
xor \U$1107 ( \1450 , \1449 , \1203 );
and \U$1108 ( \1451 , \1448 , \1450 );
xor \U$1109 ( \1452 , \1317 , \1327 );
xor \U$1110 ( \1453 , \1452 , \1330 );
and \U$1111 ( \1454 , \1450 , \1453 );
and \U$1112 ( \1455 , \1448 , \1453 );
or \U$1113 ( \1456 , \1451 , \1454 , \1455 );
xor \U$1114 ( \1457 , \1333 , \1335 );
xor \U$1115 ( \1458 , \1457 , \1338 );
and \U$1116 ( \1459 , \1456 , \1458 );
and \U$1117 ( \1460 , \1347 , \1459 );
xor \U$1118 ( \1461 , \1347 , \1459 );
xor \U$1119 ( \1462 , \1456 , \1458 );
buf \U$1120 ( \1463 , RIbb2eb48_24);
buf \U$1121 ( \1464 , RIbb2ead0_25);
and \U$1122 ( \1465 , \1463 , \1464 );
not \U$1123 ( \1466 , \1465 );
and \U$1124 ( \1467 , \1235 , \1466 );
not \U$1125 ( \1468 , \1467 );
and \U$1126 ( \1469 , \351 , \1351 );
and \U$1127 ( \1470 , \359 , \1349 );
nor \U$1128 ( \1471 , \1469 , \1470 );
xnor \U$1129 ( \1472 , \1471 , \1238 );
and \U$1130 ( \1473 , \1468 , \1472 );
and \U$1131 ( \1474 , \367 , \1157 );
and \U$1132 ( \1475 , \375 , \1155 );
nor \U$1133 ( \1476 , \1474 , \1475 );
xnor \U$1134 ( \1477 , \1476 , \1021 );
and \U$1135 ( \1478 , \1472 , \1477 );
and \U$1136 ( \1479 , \1468 , \1477 );
or \U$1137 ( \1480 , \1473 , \1478 , \1479 );
and \U$1138 ( \1481 , \385 , \957 );
and \U$1139 ( \1482 , \393 , \955 );
nor \U$1140 ( \1483 , \1481 , \1482 );
xnor \U$1141 ( \1484 , \1483 , \879 );
and \U$1142 ( \1485 , \400 , \793 );
and \U$1143 ( \1486 , \408 , \791 );
nor \U$1144 ( \1487 , \1485 , \1486 );
xnor \U$1145 ( \1488 , \1487 , \699 );
and \U$1146 ( \1489 , \1484 , \1488 );
and \U$1147 ( \1490 , \416 , \624 );
and \U$1148 ( \1491 , \424 , \622 );
nor \U$1149 ( \1492 , \1490 , \1491 );
xnor \U$1150 ( \1493 , \1492 , \349 );
and \U$1151 ( \1494 , \1488 , \1493 );
and \U$1152 ( \1495 , \1484 , \1493 );
or \U$1153 ( \1496 , \1489 , \1494 , \1495 );
and \U$1154 ( \1497 , \1480 , \1496 );
and \U$1155 ( \1498 , \435 , \357 );
and \U$1156 ( \1499 , \443 , \355 );
nor \U$1157 ( \1500 , \1498 , \1499 );
xnor \U$1158 ( \1501 , \1500 , \364 );
and \U$1159 ( \1502 , \661 , \373 );
and \U$1160 ( \1503 , \450 , \371 );
nor \U$1161 ( \1504 , \1502 , \1503 );
xnor \U$1162 ( \1505 , \1504 , \380 );
and \U$1163 ( \1506 , \1501 , \1505 );
and \U$1164 ( \1507 , \785 , \391 );
and \U$1165 ( \1508 , \722 , \389 );
nor \U$1166 ( \1509 , \1507 , \1508 );
xnor \U$1167 ( \1510 , \1509 , \398 );
and \U$1168 ( \1511 , \1505 , \1510 );
and \U$1169 ( \1512 , \1501 , \1510 );
or \U$1170 ( \1513 , \1506 , \1511 , \1512 );
and \U$1171 ( \1514 , \1496 , \1513 );
and \U$1172 ( \1515 , \1480 , \1513 );
or \U$1173 ( \1516 , \1497 , \1514 , \1515 );
xor \U$1174 ( \1517 , \1354 , \1358 );
xor \U$1175 ( \1518 , \1517 , \1363 );
xor \U$1176 ( \1519 , \1370 , \1374 );
xor \U$1177 ( \1520 , \1519 , \1379 );
and \U$1178 ( \1521 , \1518 , \1520 );
xor \U$1179 ( \1522 , \1387 , \1391 );
xor \U$1180 ( \1523 , \1522 , \1396 );
and \U$1181 ( \1524 , \1520 , \1523 );
and \U$1182 ( \1525 , \1518 , \1523 );
or \U$1183 ( \1526 , \1521 , \1524 , \1525 );
and \U$1184 ( \1527 , \1516 , \1526 );
and \U$1185 ( \1528 , \1071 , \406 );
and \U$1186 ( \1529 , \983 , \404 );
nor \U$1187 ( \1530 , \1528 , \1529 );
xnor \U$1188 ( \1531 , \1530 , \413 );
and \U$1189 ( \1532 , \1181 , \422 );
and \U$1190 ( \1533 , \1176 , \420 );
nor \U$1191 ( \1534 , \1532 , \1533 );
xnor \U$1192 ( \1535 , \1534 , \429 );
and \U$1193 ( \1536 , \1531 , \1535 );
and \U$1194 ( \1537 , \1412 , \441 );
and \U$1195 ( \1538 , \1297 , \439 );
nor \U$1196 ( \1539 , \1537 , \1538 );
xnor \U$1197 ( \1540 , \1539 , \448 );
and \U$1198 ( \1541 , \1535 , \1540 );
and \U$1199 ( \1542 , \1531 , \1540 );
or \U$1200 ( \1543 , \1536 , \1541 , \1542 );
xor \U$1201 ( \1544 , \1406 , \1410 );
xor \U$1202 ( \1545 , \1544 , \1413 );
or \U$1203 ( \1546 , \1543 , \1545 );
and \U$1204 ( \1547 , \1526 , \1546 );
and \U$1205 ( \1548 , \1516 , \1546 );
or \U$1206 ( \1549 , \1527 , \1547 , \1548 );
xor \U$1207 ( \1550 , \1366 , \1382 );
xor \U$1208 ( \1551 , \1550 , \1399 );
xor \U$1209 ( \1552 , \1416 , \1418 );
xor \U$1210 ( \1553 , \1552 , \1421 );
and \U$1211 ( \1554 , \1551 , \1553 );
xor \U$1212 ( \1555 , \1427 , \1429 );
and \U$1213 ( \1556 , \1553 , \1555 );
and \U$1214 ( \1557 , \1551 , \1555 );
or \U$1215 ( \1558 , \1554 , \1556 , \1557 );
and \U$1216 ( \1559 , \1549 , \1558 );
xor \U$1217 ( \1560 , \1435 , \1437 );
xor \U$1218 ( \1561 , \1560 , \1439 );
and \U$1219 ( \1562 , \1558 , \1561 );
and \U$1220 ( \1563 , \1549 , \1561 );
or \U$1221 ( \1564 , \1559 , \1562 , \1563 );
xor \U$1222 ( \1565 , \1287 , \1308 );
xor \U$1223 ( \1566 , \1565 , \1314 );
and \U$1224 ( \1567 , \1564 , \1566 );
xor \U$1225 ( \1568 , \1433 , \1442 );
xor \U$1226 ( \1569 , \1568 , \1445 );
and \U$1227 ( \1570 , \1566 , \1569 );
and \U$1228 ( \1571 , \1564 , \1569 );
or \U$1229 ( \1572 , \1567 , \1570 , \1571 );
xor \U$1230 ( \1573 , \1448 , \1450 );
xor \U$1231 ( \1574 , \1573 , \1453 );
and \U$1232 ( \1575 , \1572 , \1574 );
and \U$1233 ( \1576 , \1462 , \1575 );
xor \U$1234 ( \1577 , \1462 , \1575 );
xor \U$1235 ( \1578 , \1572 , \1574 );
and \U$1236 ( \1579 , \1176 , \406 );
and \U$1237 ( \1580 , \1071 , \404 );
nor \U$1238 ( \1581 , \1579 , \1580 );
xnor \U$1239 ( \1582 , \1581 , \413 );
and \U$1240 ( \1583 , \1297 , \422 );
and \U$1241 ( \1584 , \1181 , \420 );
nor \U$1242 ( \1585 , \1583 , \1584 );
xnor \U$1243 ( \1586 , \1585 , \429 );
and \U$1244 ( \1587 , \1582 , \1586 );
buf \U$1245 ( \1588 , RIbb2cdc0_87);
and \U$1246 ( \1589 , \1588 , \441 );
and \U$1247 ( \1590 , \1412 , \439 );
nor \U$1248 ( \1591 , \1589 , \1590 );
xnor \U$1249 ( \1592 , \1591 , \448 );
and \U$1250 ( \1593 , \1586 , \1592 );
and \U$1251 ( \1594 , \1582 , \1592 );
or \U$1252 ( \1595 , \1587 , \1593 , \1594 );
buf \U$1253 ( \1596 , RIbb2cd48_88);
and \U$1254 ( \1597 , \1596 , \436 );
buf \U$1255 ( \1598 , \1597 );
and \U$1256 ( \1599 , \1595 , \1598 );
and \U$1257 ( \1600 , \1588 , \436 );
and \U$1258 ( \1601 , \1598 , \1600 );
and \U$1259 ( \1602 , \1595 , \1600 );
or \U$1260 ( \1603 , \1599 , \1601 , \1602 );
and \U$1261 ( \1604 , \408 , \957 );
and \U$1262 ( \1605 , \385 , \955 );
nor \U$1263 ( \1606 , \1604 , \1605 );
xnor \U$1264 ( \1607 , \1606 , \879 );
and \U$1265 ( \1608 , \424 , \793 );
and \U$1266 ( \1609 , \400 , \791 );
nor \U$1267 ( \1610 , \1608 , \1609 );
xnor \U$1268 ( \1611 , \1610 , \699 );
and \U$1269 ( \1612 , \1607 , \1611 );
and \U$1270 ( \1613 , \443 , \624 );
and \U$1271 ( \1614 , \416 , \622 );
nor \U$1272 ( \1615 , \1613 , \1614 );
xnor \U$1273 ( \1616 , \1615 , \349 );
and \U$1274 ( \1617 , \1611 , \1616 );
and \U$1275 ( \1618 , \1607 , \1616 );
or \U$1276 ( \1619 , \1612 , \1617 , \1618 );
xor \U$1277 ( \1620 , \1235 , \1463 );
xor \U$1278 ( \1621 , \1463 , \1464 );
not \U$1279 ( \1622 , \1621 );
and \U$1280 ( \1623 , \1620 , \1622 );
and \U$1281 ( \1624 , \359 , \1623 );
not \U$1282 ( \1625 , \1624 );
xnor \U$1283 ( \1626 , \1625 , \1467 );
and \U$1284 ( \1627 , \375 , \1351 );
and \U$1285 ( \1628 , \351 , \1349 );
nor \U$1286 ( \1629 , \1627 , \1628 );
xnor \U$1287 ( \1630 , \1629 , \1238 );
and \U$1288 ( \1631 , \1626 , \1630 );
and \U$1289 ( \1632 , \393 , \1157 );
and \U$1290 ( \1633 , \367 , \1155 );
nor \U$1291 ( \1634 , \1632 , \1633 );
xnor \U$1292 ( \1635 , \1634 , \1021 );
and \U$1293 ( \1636 , \1630 , \1635 );
and \U$1294 ( \1637 , \1626 , \1635 );
or \U$1295 ( \1638 , \1631 , \1636 , \1637 );
and \U$1296 ( \1639 , \1619 , \1638 );
and \U$1297 ( \1640 , \450 , \357 );
and \U$1298 ( \1641 , \435 , \355 );
nor \U$1299 ( \1642 , \1640 , \1641 );
xnor \U$1300 ( \1643 , \1642 , \364 );
and \U$1301 ( \1644 , \722 , \373 );
and \U$1302 ( \1645 , \661 , \371 );
nor \U$1303 ( \1646 , \1644 , \1645 );
xnor \U$1304 ( \1647 , \1646 , \380 );
and \U$1305 ( \1648 , \1643 , \1647 );
and \U$1306 ( \1649 , \983 , \391 );
and \U$1307 ( \1650 , \785 , \389 );
nor \U$1308 ( \1651 , \1649 , \1650 );
xnor \U$1309 ( \1652 , \1651 , \398 );
and \U$1310 ( \1653 , \1647 , \1652 );
and \U$1311 ( \1654 , \1643 , \1652 );
or \U$1312 ( \1655 , \1648 , \1653 , \1654 );
and \U$1313 ( \1656 , \1638 , \1655 );
and \U$1314 ( \1657 , \1619 , \1655 );
or \U$1315 ( \1658 , \1639 , \1656 , \1657 );
and \U$1316 ( \1659 , \1603 , \1658 );
xor \U$1317 ( \1660 , \1484 , \1488 );
xor \U$1318 ( \1661 , \1660 , \1493 );
xor \U$1319 ( \1662 , \1531 , \1535 );
xor \U$1320 ( \1663 , \1662 , \1540 );
and \U$1321 ( \1664 , \1661 , \1663 );
xor \U$1322 ( \1665 , \1501 , \1505 );
xor \U$1323 ( \1666 , \1665 , \1510 );
and \U$1324 ( \1667 , \1663 , \1666 );
and \U$1325 ( \1668 , \1661 , \1666 );
or \U$1326 ( \1669 , \1664 , \1667 , \1668 );
and \U$1327 ( \1670 , \1658 , \1669 );
and \U$1328 ( \1671 , \1603 , \1669 );
or \U$1329 ( \1672 , \1659 , \1670 , \1671 );
xor \U$1330 ( \1673 , \1480 , \1496 );
xor \U$1331 ( \1674 , \1673 , \1513 );
xor \U$1332 ( \1675 , \1518 , \1520 );
xor \U$1333 ( \1676 , \1675 , \1523 );
and \U$1334 ( \1677 , \1674 , \1676 );
xnor \U$1335 ( \1678 , \1543 , \1545 );
and \U$1336 ( \1679 , \1676 , \1678 );
and \U$1337 ( \1680 , \1674 , \1678 );
or \U$1338 ( \1681 , \1677 , \1679 , \1680 );
and \U$1339 ( \1682 , \1672 , \1681 );
xor \U$1340 ( \1683 , \1551 , \1553 );
xor \U$1341 ( \1684 , \1683 , \1555 );
and \U$1342 ( \1685 , \1681 , \1684 );
and \U$1343 ( \1686 , \1672 , \1684 );
or \U$1344 ( \1687 , \1682 , \1685 , \1686 );
xor \U$1345 ( \1688 , \1402 , \1424 );
xor \U$1346 ( \1689 , \1688 , \1430 );
and \U$1347 ( \1690 , \1687 , \1689 );
xor \U$1348 ( \1691 , \1549 , \1558 );
xor \U$1349 ( \1692 , \1691 , \1561 );
and \U$1350 ( \1693 , \1689 , \1692 );
and \U$1351 ( \1694 , \1687 , \1692 );
or \U$1352 ( \1695 , \1690 , \1693 , \1694 );
xor \U$1353 ( \1696 , \1564 , \1566 );
xor \U$1354 ( \1697 , \1696 , \1569 );
and \U$1355 ( \1698 , \1695 , \1697 );
and \U$1356 ( \1699 , \1578 , \1698 );
xor \U$1357 ( \1700 , \1578 , \1698 );
xor \U$1358 ( \1701 , \1695 , \1697 );
and \U$1359 ( \1702 , \435 , \624 );
and \U$1360 ( \1703 , \443 , \622 );
nor \U$1361 ( \1704 , \1702 , \1703 );
xnor \U$1362 ( \1705 , \1704 , \349 );
and \U$1363 ( \1706 , \661 , \357 );
and \U$1364 ( \1707 , \450 , \355 );
nor \U$1365 ( \1708 , \1706 , \1707 );
xnor \U$1366 ( \1709 , \1708 , \364 );
and \U$1367 ( \1710 , \1705 , \1709 );
and \U$1368 ( \1711 , \785 , \373 );
and \U$1369 ( \1712 , \722 , \371 );
nor \U$1370 ( \1713 , \1711 , \1712 );
xnor \U$1371 ( \1714 , \1713 , \380 );
and \U$1372 ( \1715 , \1709 , \1714 );
and \U$1373 ( \1716 , \1705 , \1714 );
or \U$1374 ( \1717 , \1710 , \1715 , \1716 );
and \U$1375 ( \1718 , \385 , \1157 );
and \U$1376 ( \1719 , \393 , \1155 );
nor \U$1377 ( \1720 , \1718 , \1719 );
xnor \U$1378 ( \1721 , \1720 , \1021 );
and \U$1379 ( \1722 , \400 , \957 );
and \U$1380 ( \1723 , \408 , \955 );
nor \U$1381 ( \1724 , \1722 , \1723 );
xnor \U$1382 ( \1725 , \1724 , \879 );
and \U$1383 ( \1726 , \1721 , \1725 );
and \U$1384 ( \1727 , \416 , \793 );
and \U$1385 ( \1728 , \424 , \791 );
nor \U$1386 ( \1729 , \1727 , \1728 );
xnor \U$1387 ( \1730 , \1729 , \699 );
and \U$1388 ( \1731 , \1725 , \1730 );
and \U$1389 ( \1732 , \1721 , \1730 );
or \U$1390 ( \1733 , \1726 , \1731 , \1732 );
and \U$1391 ( \1734 , \1717 , \1733 );
buf \U$1392 ( \1735 , RIbb2ea58_26);
buf \U$1393 ( \1736 , RIbb2e9e0_27);
and \U$1394 ( \1737 , \1735 , \1736 );
not \U$1395 ( \1738 , \1737 );
and \U$1396 ( \1739 , \1464 , \1738 );
not \U$1397 ( \1740 , \1739 );
and \U$1398 ( \1741 , \351 , \1623 );
and \U$1399 ( \1742 , \359 , \1621 );
nor \U$1400 ( \1743 , \1741 , \1742 );
xnor \U$1401 ( \1744 , \1743 , \1467 );
and \U$1402 ( \1745 , \1740 , \1744 );
and \U$1403 ( \1746 , \367 , \1351 );
and \U$1404 ( \1747 , \375 , \1349 );
nor \U$1405 ( \1748 , \1746 , \1747 );
xnor \U$1406 ( \1749 , \1748 , \1238 );
and \U$1407 ( \1750 , \1744 , \1749 );
and \U$1408 ( \1751 , \1740 , \1749 );
or \U$1409 ( \1752 , \1745 , \1750 , \1751 );
and \U$1410 ( \1753 , \1733 , \1752 );
and \U$1411 ( \1754 , \1717 , \1752 );
or \U$1412 ( \1755 , \1734 , \1753 , \1754 );
xor \U$1413 ( \1756 , \1607 , \1611 );
xor \U$1414 ( \1757 , \1756 , \1616 );
xor \U$1415 ( \1758 , \1626 , \1630 );
xor \U$1416 ( \1759 , \1758 , \1635 );
and \U$1417 ( \1760 , \1757 , \1759 );
xor \U$1418 ( \1761 , \1643 , \1647 );
xor \U$1419 ( \1762 , \1761 , \1652 );
and \U$1420 ( \1763 , \1759 , \1762 );
and \U$1421 ( \1764 , \1757 , \1762 );
or \U$1422 ( \1765 , \1760 , \1763 , \1764 );
and \U$1423 ( \1766 , \1755 , \1765 );
and \U$1424 ( \1767 , \1071 , \391 );
and \U$1425 ( \1768 , \983 , \389 );
nor \U$1426 ( \1769 , \1767 , \1768 );
xnor \U$1427 ( \1770 , \1769 , \398 );
and \U$1428 ( \1771 , \1181 , \406 );
and \U$1429 ( \1772 , \1176 , \404 );
nor \U$1430 ( \1773 , \1771 , \1772 );
xnor \U$1431 ( \1774 , \1773 , \413 );
and \U$1432 ( \1775 , \1770 , \1774 );
and \U$1433 ( \1776 , \1412 , \422 );
and \U$1434 ( \1777 , \1297 , \420 );
nor \U$1435 ( \1778 , \1776 , \1777 );
xnor \U$1436 ( \1779 , \1778 , \429 );
and \U$1437 ( \1780 , \1774 , \1779 );
and \U$1438 ( \1781 , \1770 , \1779 );
or \U$1439 ( \1782 , \1775 , \1780 , \1781 );
xor \U$1440 ( \1783 , \1582 , \1586 );
xor \U$1441 ( \1784 , \1783 , \1592 );
and \U$1442 ( \1785 , \1782 , \1784 );
not \U$1443 ( \1786 , \1597 );
and \U$1444 ( \1787 , \1784 , \1786 );
and \U$1445 ( \1788 , \1782 , \1786 );
or \U$1446 ( \1789 , \1785 , \1787 , \1788 );
and \U$1447 ( \1790 , \1765 , \1789 );
and \U$1448 ( \1791 , \1755 , \1789 );
or \U$1449 ( \1792 , \1766 , \1790 , \1791 );
xor \U$1450 ( \1793 , \1468 , \1472 );
xor \U$1451 ( \1794 , \1793 , \1477 );
xor \U$1452 ( \1795 , \1595 , \1598 );
xor \U$1453 ( \1796 , \1795 , \1600 );
and \U$1454 ( \1797 , \1794 , \1796 );
xor \U$1455 ( \1798 , \1661 , \1663 );
xor \U$1456 ( \1799 , \1798 , \1666 );
and \U$1457 ( \1800 , \1796 , \1799 );
and \U$1458 ( \1801 , \1794 , \1799 );
or \U$1459 ( \1802 , \1797 , \1800 , \1801 );
and \U$1460 ( \1803 , \1792 , \1802 );
xor \U$1461 ( \1804 , \1674 , \1676 );
xor \U$1462 ( \1805 , \1804 , \1678 );
and \U$1463 ( \1806 , \1802 , \1805 );
and \U$1464 ( \1807 , \1792 , \1805 );
or \U$1465 ( \1808 , \1803 , \1806 , \1807 );
xor \U$1466 ( \1809 , \1516 , \1526 );
xor \U$1467 ( \1810 , \1809 , \1546 );
and \U$1468 ( \1811 , \1808 , \1810 );
xor \U$1469 ( \1812 , \1672 , \1681 );
xor \U$1470 ( \1813 , \1812 , \1684 );
and \U$1471 ( \1814 , \1810 , \1813 );
and \U$1472 ( \1815 , \1808 , \1813 );
or \U$1473 ( \1816 , \1811 , \1814 , \1815 );
xor \U$1474 ( \1817 , \1687 , \1689 );
xor \U$1475 ( \1818 , \1817 , \1692 );
and \U$1476 ( \1819 , \1816 , \1818 );
and \U$1477 ( \1820 , \1701 , \1819 );
xor \U$1478 ( \1821 , \1701 , \1819 );
xor \U$1479 ( \1822 , \1816 , \1818 );
and \U$1480 ( \1823 , \1176 , \391 );
and \U$1481 ( \1824 , \1071 , \389 );
nor \U$1482 ( \1825 , \1823 , \1824 );
xnor \U$1483 ( \1826 , \1825 , \398 );
and \U$1484 ( \1827 , \1297 , \406 );
and \U$1485 ( \1828 , \1181 , \404 );
nor \U$1486 ( \1829 , \1827 , \1828 );
xnor \U$1487 ( \1830 , \1829 , \413 );
and \U$1488 ( \1831 , \1826 , \1830 );
and \U$1489 ( \1832 , \1588 , \422 );
and \U$1490 ( \1833 , \1412 , \420 );
nor \U$1491 ( \1834 , \1832 , \1833 );
xnor \U$1492 ( \1835 , \1834 , \429 );
and \U$1493 ( \1836 , \1830 , \1835 );
and \U$1494 ( \1837 , \1826 , \1835 );
or \U$1495 ( \1838 , \1831 , \1836 , \1837 );
buf \U$1496 ( \1839 , RIbb2ccd0_89);
and \U$1497 ( \1840 , \1839 , \441 );
and \U$1498 ( \1841 , \1596 , \439 );
nor \U$1499 ( \1842 , \1840 , \1841 );
xnor \U$1500 ( \1843 , \1842 , \448 );
buf \U$1501 ( \1844 , RIbb2cc58_90);
and \U$1502 ( \1845 , \1844 , \436 );
or \U$1503 ( \1846 , \1843 , \1845 );
and \U$1504 ( \1847 , \1838 , \1846 );
and \U$1505 ( \1848 , \1596 , \441 );
and \U$1506 ( \1849 , \1588 , \439 );
nor \U$1507 ( \1850 , \1848 , \1849 );
xnor \U$1508 ( \1851 , \1850 , \448 );
and \U$1509 ( \1852 , \1846 , \1851 );
and \U$1510 ( \1853 , \1838 , \1851 );
or \U$1511 ( \1854 , \1847 , \1852 , \1853 );
and \U$1512 ( \1855 , \450 , \624 );
and \U$1513 ( \1856 , \435 , \622 );
nor \U$1514 ( \1857 , \1855 , \1856 );
xnor \U$1515 ( \1858 , \1857 , \349 );
and \U$1516 ( \1859 , \722 , \357 );
and \U$1517 ( \1860 , \661 , \355 );
nor \U$1518 ( \1861 , \1859 , \1860 );
xnor \U$1519 ( \1862 , \1861 , \364 );
and \U$1520 ( \1863 , \1858 , \1862 );
and \U$1521 ( \1864 , \983 , \373 );
and \U$1522 ( \1865 , \785 , \371 );
nor \U$1523 ( \1866 , \1864 , \1865 );
xnor \U$1524 ( \1867 , \1866 , \380 );
and \U$1525 ( \1868 , \1862 , \1867 );
and \U$1526 ( \1869 , \1858 , \1867 );
or \U$1527 ( \1870 , \1863 , \1868 , \1869 );
and \U$1528 ( \1871 , \408 , \1157 );
and \U$1529 ( \1872 , \385 , \1155 );
nor \U$1530 ( \1873 , \1871 , \1872 );
xnor \U$1531 ( \1874 , \1873 , \1021 );
and \U$1532 ( \1875 , \424 , \957 );
and \U$1533 ( \1876 , \400 , \955 );
nor \U$1534 ( \1877 , \1875 , \1876 );
xnor \U$1535 ( \1878 , \1877 , \879 );
and \U$1536 ( \1879 , \1874 , \1878 );
and \U$1537 ( \1880 , \443 , \793 );
and \U$1538 ( \1881 , \416 , \791 );
nor \U$1539 ( \1882 , \1880 , \1881 );
xnor \U$1540 ( \1883 , \1882 , \699 );
and \U$1541 ( \1884 , \1878 , \1883 );
and \U$1542 ( \1885 , \1874 , \1883 );
or \U$1543 ( \1886 , \1879 , \1884 , \1885 );
and \U$1544 ( \1887 , \1870 , \1886 );
xor \U$1545 ( \1888 , \1464 , \1735 );
xor \U$1546 ( \1889 , \1735 , \1736 );
not \U$1547 ( \1890 , \1889 );
and \U$1548 ( \1891 , \1888 , \1890 );
and \U$1549 ( \1892 , \359 , \1891 );
not \U$1550 ( \1893 , \1892 );
xnor \U$1551 ( \1894 , \1893 , \1739 );
and \U$1552 ( \1895 , \375 , \1623 );
and \U$1553 ( \1896 , \351 , \1621 );
nor \U$1554 ( \1897 , \1895 , \1896 );
xnor \U$1555 ( \1898 , \1897 , \1467 );
and \U$1556 ( \1899 , \1894 , \1898 );
and \U$1557 ( \1900 , \393 , \1351 );
and \U$1558 ( \1901 , \367 , \1349 );
nor \U$1559 ( \1902 , \1900 , \1901 );
xnor \U$1560 ( \1903 , \1902 , \1238 );
and \U$1561 ( \1904 , \1898 , \1903 );
and \U$1562 ( \1905 , \1894 , \1903 );
or \U$1563 ( \1906 , \1899 , \1904 , \1905 );
and \U$1564 ( \1907 , \1886 , \1906 );
and \U$1565 ( \1908 , \1870 , \1906 );
or \U$1566 ( \1909 , \1887 , \1907 , \1908 );
and \U$1567 ( \1910 , \1854 , \1909 );
and \U$1568 ( \1911 , \1839 , \436 );
xor \U$1569 ( \1912 , \1705 , \1709 );
xor \U$1570 ( \1913 , \1912 , \1714 );
and \U$1571 ( \1914 , \1911 , \1913 );
xor \U$1572 ( \1915 , \1770 , \1774 );
xor \U$1573 ( \1916 , \1915 , \1779 );
and \U$1574 ( \1917 , \1913 , \1916 );
and \U$1575 ( \1918 , \1911 , \1916 );
or \U$1576 ( \1919 , \1914 , \1917 , \1918 );
and \U$1577 ( \1920 , \1909 , \1919 );
and \U$1578 ( \1921 , \1854 , \1919 );
or \U$1579 ( \1922 , \1910 , \1920 , \1921 );
xor \U$1580 ( \1923 , \1717 , \1733 );
xor \U$1581 ( \1924 , \1923 , \1752 );
xor \U$1582 ( \1925 , \1757 , \1759 );
xor \U$1583 ( \1926 , \1925 , \1762 );
and \U$1584 ( \1927 , \1924 , \1926 );
xor \U$1585 ( \1928 , \1782 , \1784 );
xor \U$1586 ( \1929 , \1928 , \1786 );
and \U$1587 ( \1930 , \1926 , \1929 );
and \U$1588 ( \1931 , \1924 , \1929 );
or \U$1589 ( \1932 , \1927 , \1930 , \1931 );
and \U$1590 ( \1933 , \1922 , \1932 );
xor \U$1591 ( \1934 , \1619 , \1638 );
xor \U$1592 ( \1935 , \1934 , \1655 );
and \U$1593 ( \1936 , \1932 , \1935 );
and \U$1594 ( \1937 , \1922 , \1935 );
or \U$1595 ( \1938 , \1933 , \1936 , \1937 );
xor \U$1596 ( \1939 , \1755 , \1765 );
xor \U$1597 ( \1940 , \1939 , \1789 );
xor \U$1598 ( \1941 , \1794 , \1796 );
xor \U$1599 ( \1942 , \1941 , \1799 );
and \U$1600 ( \1943 , \1940 , \1942 );
and \U$1601 ( \1944 , \1938 , \1943 );
xor \U$1602 ( \1945 , \1603 , \1658 );
xor \U$1603 ( \1946 , \1945 , \1669 );
and \U$1604 ( \1947 , \1943 , \1946 );
and \U$1605 ( \1948 , \1938 , \1946 );
or \U$1606 ( \1949 , \1944 , \1947 , \1948 );
xor \U$1607 ( \1950 , \1808 , \1810 );
xor \U$1608 ( \1951 , \1950 , \1813 );
and \U$1609 ( \1952 , \1949 , \1951 );
and \U$1610 ( \1953 , \1822 , \1952 );
xor \U$1611 ( \1954 , \1822 , \1952 );
xor \U$1612 ( \1955 , \1949 , \1951 );
buf \U$1613 ( \1956 , RIbb2e968_28);
buf \U$1614 ( \1957 , RIbb2e8f0_29);
and \U$1615 ( \1958 , \1956 , \1957 );
not \U$1616 ( \1959 , \1958 );
and \U$1617 ( \1960 , \1736 , \1959 );
not \U$1618 ( \1961 , \1960 );
and \U$1619 ( \1962 , \351 , \1891 );
and \U$1620 ( \1963 , \359 , \1889 );
nor \U$1621 ( \1964 , \1962 , \1963 );
xnor \U$1622 ( \1965 , \1964 , \1739 );
and \U$1623 ( \1966 , \1961 , \1965 );
and \U$1624 ( \1967 , \367 , \1623 );
and \U$1625 ( \1968 , \375 , \1621 );
nor \U$1626 ( \1969 , \1967 , \1968 );
xnor \U$1627 ( \1970 , \1969 , \1467 );
and \U$1628 ( \1971 , \1965 , \1970 );
and \U$1629 ( \1972 , \1961 , \1970 );
or \U$1630 ( \1973 , \1966 , \1971 , \1972 );
and \U$1631 ( \1974 , \385 , \1351 );
and \U$1632 ( \1975 , \393 , \1349 );
nor \U$1633 ( \1976 , \1974 , \1975 );
xnor \U$1634 ( \1977 , \1976 , \1238 );
and \U$1635 ( \1978 , \400 , \1157 );
and \U$1636 ( \1979 , \408 , \1155 );
nor \U$1637 ( \1980 , \1978 , \1979 );
xnor \U$1638 ( \1981 , \1980 , \1021 );
and \U$1639 ( \1982 , \1977 , \1981 );
and \U$1640 ( \1983 , \416 , \957 );
and \U$1641 ( \1984 , \424 , \955 );
nor \U$1642 ( \1985 , \1983 , \1984 );
xnor \U$1643 ( \1986 , \1985 , \879 );
and \U$1644 ( \1987 , \1981 , \1986 );
and \U$1645 ( \1988 , \1977 , \1986 );
or \U$1646 ( \1989 , \1982 , \1987 , \1988 );
and \U$1647 ( \1990 , \1973 , \1989 );
and \U$1648 ( \1991 , \435 , \793 );
and \U$1649 ( \1992 , \443 , \791 );
nor \U$1650 ( \1993 , \1991 , \1992 );
xnor \U$1651 ( \1994 , \1993 , \699 );
and \U$1652 ( \1995 , \661 , \624 );
and \U$1653 ( \1996 , \450 , \622 );
nor \U$1654 ( \1997 , \1995 , \1996 );
xnor \U$1655 ( \1998 , \1997 , \349 );
and \U$1656 ( \1999 , \1994 , \1998 );
and \U$1657 ( \2000 , \785 , \357 );
and \U$1658 ( \2001 , \722 , \355 );
nor \U$1659 ( \2002 , \2000 , \2001 );
xnor \U$1660 ( \2003 , \2002 , \364 );
and \U$1661 ( \2004 , \1998 , \2003 );
and \U$1662 ( \2005 , \1994 , \2003 );
or \U$1663 ( \2006 , \1999 , \2004 , \2005 );
and \U$1664 ( \2007 , \1989 , \2006 );
and \U$1665 ( \2008 , \1973 , \2006 );
or \U$1666 ( \2009 , \1990 , \2007 , \2008 );
xor \U$1667 ( \2010 , \1858 , \1862 );
xor \U$1668 ( \2011 , \2010 , \1867 );
xor \U$1669 ( \2012 , \1874 , \1878 );
xor \U$1670 ( \2013 , \2012 , \1883 );
and \U$1671 ( \2014 , \2011 , \2013 );
xor \U$1672 ( \2015 , \1826 , \1830 );
xor \U$1673 ( \2016 , \2015 , \1835 );
and \U$1674 ( \2017 , \2013 , \2016 );
and \U$1675 ( \2018 , \2011 , \2016 );
or \U$1676 ( \2019 , \2014 , \2017 , \2018 );
and \U$1677 ( \2020 , \2009 , \2019 );
and \U$1678 ( \2021 , \1596 , \422 );
and \U$1679 ( \2022 , \1588 , \420 );
nor \U$1680 ( \2023 , \2021 , \2022 );
xnor \U$1681 ( \2024 , \2023 , \429 );
and \U$1682 ( \2025 , \1844 , \441 );
and \U$1683 ( \2026 , \1839 , \439 );
nor \U$1684 ( \2027 , \2025 , \2026 );
xnor \U$1685 ( \2028 , \2027 , \448 );
and \U$1686 ( \2029 , \2024 , \2028 );
buf \U$1687 ( \2030 , RIbb2cbe0_91);
and \U$1688 ( \2031 , \2030 , \436 );
and \U$1689 ( \2032 , \2028 , \2031 );
and \U$1690 ( \2033 , \2024 , \2031 );
or \U$1691 ( \2034 , \2029 , \2032 , \2033 );
and \U$1692 ( \2035 , \1071 , \373 );
and \U$1693 ( \2036 , \983 , \371 );
nor \U$1694 ( \2037 , \2035 , \2036 );
xnor \U$1695 ( \2038 , \2037 , \380 );
and \U$1696 ( \2039 , \1181 , \391 );
and \U$1697 ( \2040 , \1176 , \389 );
nor \U$1698 ( \2041 , \2039 , \2040 );
xnor \U$1699 ( \2042 , \2041 , \398 );
and \U$1700 ( \2043 , \2038 , \2042 );
and \U$1701 ( \2044 , \1412 , \406 );
and \U$1702 ( \2045 , \1297 , \404 );
nor \U$1703 ( \2046 , \2044 , \2045 );
xnor \U$1704 ( \2047 , \2046 , \413 );
and \U$1705 ( \2048 , \2042 , \2047 );
and \U$1706 ( \2049 , \2038 , \2047 );
or \U$1707 ( \2050 , \2043 , \2048 , \2049 );
and \U$1708 ( \2051 , \2034 , \2050 );
xnor \U$1709 ( \2052 , \1843 , \1845 );
and \U$1710 ( \2053 , \2050 , \2052 );
and \U$1711 ( \2054 , \2034 , \2052 );
or \U$1712 ( \2055 , \2051 , \2053 , \2054 );
and \U$1713 ( \2056 , \2019 , \2055 );
and \U$1714 ( \2057 , \2009 , \2055 );
or \U$1715 ( \2058 , \2020 , \2056 , \2057 );
xor \U$1716 ( \2059 , \1721 , \1725 );
xor \U$1717 ( \2060 , \2059 , \1730 );
xor \U$1718 ( \2061 , \1740 , \1744 );
xor \U$1719 ( \2062 , \2061 , \1749 );
and \U$1720 ( \2063 , \2060 , \2062 );
xor \U$1721 ( \2064 , \1911 , \1913 );
xor \U$1722 ( \2065 , \2064 , \1916 );
and \U$1723 ( \2066 , \2062 , \2065 );
and \U$1724 ( \2067 , \2060 , \2065 );
or \U$1725 ( \2068 , \2063 , \2066 , \2067 );
and \U$1726 ( \2069 , \2058 , \2068 );
xor \U$1727 ( \2070 , \1924 , \1926 );
xor \U$1728 ( \2071 , \2070 , \1929 );
and \U$1729 ( \2072 , \2068 , \2071 );
and \U$1730 ( \2073 , \2058 , \2071 );
or \U$1731 ( \2074 , \2069 , \2072 , \2073 );
xor \U$1732 ( \2075 , \1922 , \1932 );
xor \U$1733 ( \2076 , \2075 , \1935 );
and \U$1734 ( \2077 , \2074 , \2076 );
xor \U$1735 ( \2078 , \1940 , \1942 );
and \U$1736 ( \2079 , \2076 , \2078 );
and \U$1737 ( \2080 , \2074 , \2078 );
or \U$1738 ( \2081 , \2077 , \2079 , \2080 );
xor \U$1739 ( \2082 , \1938 , \1943 );
xor \U$1740 ( \2083 , \2082 , \1946 );
and \U$1741 ( \2084 , \2081 , \2083 );
xor \U$1742 ( \2085 , \1792 , \1802 );
xor \U$1743 ( \2086 , \2085 , \1805 );
and \U$1744 ( \2087 , \2083 , \2086 );
and \U$1745 ( \2088 , \2081 , \2086 );
or \U$1746 ( \2089 , \2084 , \2087 , \2088 );
and \U$1747 ( \2090 , \1955 , \2089 );
xor \U$1748 ( \2091 , \1955 , \2089 );
xor \U$1749 ( \2092 , \2081 , \2083 );
xor \U$1750 ( \2093 , \2092 , \2086 );
xor \U$1751 ( \2094 , \1736 , \1956 );
xor \U$1752 ( \2095 , \1956 , \1957 );
not \U$1753 ( \2096 , \2095 );
and \U$1754 ( \2097 , \2094 , \2096 );
and \U$1755 ( \2098 , \359 , \2097 );
not \U$1756 ( \2099 , \2098 );
xnor \U$1757 ( \2100 , \2099 , \1960 );
and \U$1758 ( \2101 , \375 , \1891 );
and \U$1759 ( \2102 , \351 , \1889 );
nor \U$1760 ( \2103 , \2101 , \2102 );
xnor \U$1761 ( \2104 , \2103 , \1739 );
and \U$1762 ( \2105 , \2100 , \2104 );
and \U$1763 ( \2106 , \393 , \1623 );
and \U$1764 ( \2107 , \367 , \1621 );
nor \U$1765 ( \2108 , \2106 , \2107 );
xnor \U$1766 ( \2109 , \2108 , \1467 );
and \U$1767 ( \2110 , \2104 , \2109 );
and \U$1768 ( \2111 , \2100 , \2109 );
or \U$1769 ( \2112 , \2105 , \2110 , \2111 );
and \U$1770 ( \2113 , \408 , \1351 );
and \U$1771 ( \2114 , \385 , \1349 );
nor \U$1772 ( \2115 , \2113 , \2114 );
xnor \U$1773 ( \2116 , \2115 , \1238 );
and \U$1774 ( \2117 , \424 , \1157 );
and \U$1775 ( \2118 , \400 , \1155 );
nor \U$1776 ( \2119 , \2117 , \2118 );
xnor \U$1777 ( \2120 , \2119 , \1021 );
and \U$1778 ( \2121 , \2116 , \2120 );
and \U$1779 ( \2122 , \443 , \957 );
and \U$1780 ( \2123 , \416 , \955 );
nor \U$1781 ( \2124 , \2122 , \2123 );
xnor \U$1782 ( \2125 , \2124 , \879 );
and \U$1783 ( \2126 , \2120 , \2125 );
and \U$1784 ( \2127 , \2116 , \2125 );
or \U$1785 ( \2128 , \2121 , \2126 , \2127 );
and \U$1786 ( \2129 , \2112 , \2128 );
and \U$1787 ( \2130 , \450 , \793 );
and \U$1788 ( \2131 , \435 , \791 );
nor \U$1789 ( \2132 , \2130 , \2131 );
xnor \U$1790 ( \2133 , \2132 , \699 );
and \U$1791 ( \2134 , \722 , \624 );
and \U$1792 ( \2135 , \661 , \622 );
nor \U$1793 ( \2136 , \2134 , \2135 );
xnor \U$1794 ( \2137 , \2136 , \349 );
and \U$1795 ( \2138 , \2133 , \2137 );
and \U$1796 ( \2139 , \983 , \357 );
and \U$1797 ( \2140 , \785 , \355 );
nor \U$1798 ( \2141 , \2139 , \2140 );
xnor \U$1799 ( \2142 , \2141 , \364 );
and \U$1800 ( \2143 , \2137 , \2142 );
and \U$1801 ( \2144 , \2133 , \2142 );
or \U$1802 ( \2145 , \2138 , \2143 , \2144 );
and \U$1803 ( \2146 , \2128 , \2145 );
and \U$1804 ( \2147 , \2112 , \2145 );
or \U$1805 ( \2148 , \2129 , \2146 , \2147 );
and \U$1806 ( \2149 , \1176 , \373 );
and \U$1807 ( \2150 , \1071 , \371 );
nor \U$1808 ( \2151 , \2149 , \2150 );
xnor \U$1809 ( \2152 , \2151 , \380 );
and \U$1810 ( \2153 , \1297 , \391 );
and \U$1811 ( \2154 , \1181 , \389 );
nor \U$1812 ( \2155 , \2153 , \2154 );
xnor \U$1813 ( \2156 , \2155 , \398 );
and \U$1814 ( \2157 , \2152 , \2156 );
and \U$1815 ( \2158 , \1588 , \406 );
and \U$1816 ( \2159 , \1412 , \404 );
nor \U$1817 ( \2160 , \2158 , \2159 );
xnor \U$1818 ( \2161 , \2160 , \413 );
and \U$1819 ( \2162 , \2156 , \2161 );
and \U$1820 ( \2163 , \2152 , \2161 );
or \U$1821 ( \2164 , \2157 , \2162 , \2163 );
and \U$1822 ( \2165 , \1839 , \422 );
and \U$1823 ( \2166 , \1596 , \420 );
nor \U$1824 ( \2167 , \2165 , \2166 );
xnor \U$1825 ( \2168 , \2167 , \429 );
and \U$1826 ( \2169 , \2030 , \441 );
and \U$1827 ( \2170 , \1844 , \439 );
nor \U$1828 ( \2171 , \2169 , \2170 );
xnor \U$1829 ( \2172 , \2171 , \448 );
and \U$1830 ( \2173 , \2168 , \2172 );
buf \U$1831 ( \2174 , RIbb2cb68_92);
and \U$1832 ( \2175 , \2174 , \436 );
and \U$1833 ( \2176 , \2172 , \2175 );
and \U$1834 ( \2177 , \2168 , \2175 );
or \U$1835 ( \2178 , \2173 , \2176 , \2177 );
and \U$1836 ( \2179 , \2164 , \2178 );
xor \U$1837 ( \2180 , \2024 , \2028 );
xor \U$1838 ( \2181 , \2180 , \2031 );
and \U$1839 ( \2182 , \2178 , \2181 );
and \U$1840 ( \2183 , \2164 , \2181 );
or \U$1841 ( \2184 , \2179 , \2182 , \2183 );
and \U$1842 ( \2185 , \2148 , \2184 );
xor \U$1843 ( \2186 , \1977 , \1981 );
xor \U$1844 ( \2187 , \2186 , \1986 );
xor \U$1845 ( \2188 , \2038 , \2042 );
xor \U$1846 ( \2189 , \2188 , \2047 );
and \U$1847 ( \2190 , \2187 , \2189 );
xor \U$1848 ( \2191 , \1994 , \1998 );
xor \U$1849 ( \2192 , \2191 , \2003 );
and \U$1850 ( \2193 , \2189 , \2192 );
and \U$1851 ( \2194 , \2187 , \2192 );
or \U$1852 ( \2195 , \2190 , \2193 , \2194 );
and \U$1853 ( \2196 , \2184 , \2195 );
and \U$1854 ( \2197 , \2148 , \2195 );
or \U$1855 ( \2198 , \2185 , \2196 , \2197 );
xor \U$1856 ( \2199 , \1894 , \1898 );
xor \U$1857 ( \2200 , \2199 , \1903 );
xor \U$1858 ( \2201 , \2011 , \2013 );
xor \U$1859 ( \2202 , \2201 , \2016 );
and \U$1860 ( \2203 , \2200 , \2202 );
xor \U$1861 ( \2204 , \2034 , \2050 );
xor \U$1862 ( \2205 , \2204 , \2052 );
and \U$1863 ( \2206 , \2202 , \2205 );
and \U$1864 ( \2207 , \2200 , \2205 );
or \U$1865 ( \2208 , \2203 , \2206 , \2207 );
and \U$1866 ( \2209 , \2198 , \2208 );
xor \U$1867 ( \2210 , \1838 , \1846 );
xor \U$1868 ( \2211 , \2210 , \1851 );
and \U$1869 ( \2212 , \2208 , \2211 );
and \U$1870 ( \2213 , \2198 , \2211 );
or \U$1871 ( \2214 , \2209 , \2212 , \2213 );
xor \U$1872 ( \2215 , \1870 , \1886 );
xor \U$1873 ( \2216 , \2215 , \1906 );
xor \U$1874 ( \2217 , \2009 , \2019 );
xor \U$1875 ( \2218 , \2217 , \2055 );
and \U$1876 ( \2219 , \2216 , \2218 );
xor \U$1877 ( \2220 , \2060 , \2062 );
xor \U$1878 ( \2221 , \2220 , \2065 );
and \U$1879 ( \2222 , \2218 , \2221 );
and \U$1880 ( \2223 , \2216 , \2221 );
or \U$1881 ( \2224 , \2219 , \2222 , \2223 );
and \U$1882 ( \2225 , \2214 , \2224 );
xor \U$1883 ( \2226 , \1854 , \1909 );
xor \U$1884 ( \2227 , \2226 , \1919 );
and \U$1885 ( \2228 , \2224 , \2227 );
and \U$1886 ( \2229 , \2214 , \2227 );
or \U$1887 ( \2230 , \2225 , \2228 , \2229 );
and \U$1888 ( \2231 , \385 , \1623 );
and \U$1889 ( \2232 , \393 , \1621 );
nor \U$1890 ( \2233 , \2231 , \2232 );
xnor \U$1891 ( \2234 , \2233 , \1467 );
and \U$1892 ( \2235 , \400 , \1351 );
and \U$1893 ( \2236 , \408 , \1349 );
nor \U$1894 ( \2237 , \2235 , \2236 );
xnor \U$1895 ( \2238 , \2237 , \1238 );
and \U$1896 ( \2239 , \2234 , \2238 );
and \U$1897 ( \2240 , \416 , \1157 );
and \U$1898 ( \2241 , \424 , \1155 );
nor \U$1899 ( \2242 , \2240 , \2241 );
xnor \U$1900 ( \2243 , \2242 , \1021 );
and \U$1901 ( \2244 , \2238 , \2243 );
and \U$1902 ( \2245 , \2234 , \2243 );
or \U$1903 ( \2246 , \2239 , \2244 , \2245 );
buf \U$1904 ( \2247 , RIbb2e878_30);
buf \U$1905 ( \2248 , RIbb2e800_31);
and \U$1906 ( \2249 , \2247 , \2248 );
not \U$1907 ( \2250 , \2249 );
and \U$1908 ( \2251 , \1957 , \2250 );
not \U$1909 ( \2252 , \2251 );
and \U$1910 ( \2253 , \351 , \2097 );
and \U$1911 ( \2254 , \359 , \2095 );
nor \U$1912 ( \2255 , \2253 , \2254 );
xnor \U$1913 ( \2256 , \2255 , \1960 );
and \U$1914 ( \2257 , \2252 , \2256 );
and \U$1915 ( \2258 , \367 , \1891 );
and \U$1916 ( \2259 , \375 , \1889 );
nor \U$1917 ( \2260 , \2258 , \2259 );
xnor \U$1918 ( \2261 , \2260 , \1739 );
and \U$1919 ( \2262 , \2256 , \2261 );
and \U$1920 ( \2263 , \2252 , \2261 );
or \U$1921 ( \2264 , \2257 , \2262 , \2263 );
and \U$1922 ( \2265 , \2246 , \2264 );
and \U$1923 ( \2266 , \435 , \957 );
and \U$1924 ( \2267 , \443 , \955 );
nor \U$1925 ( \2268 , \2266 , \2267 );
xnor \U$1926 ( \2269 , \2268 , \879 );
and \U$1927 ( \2270 , \661 , \793 );
and \U$1928 ( \2271 , \450 , \791 );
nor \U$1929 ( \2272 , \2270 , \2271 );
xnor \U$1930 ( \2273 , \2272 , \699 );
and \U$1931 ( \2274 , \2269 , \2273 );
and \U$1932 ( \2275 , \785 , \624 );
and \U$1933 ( \2276 , \722 , \622 );
nor \U$1934 ( \2277 , \2275 , \2276 );
xnor \U$1935 ( \2278 , \2277 , \349 );
and \U$1936 ( \2279 , \2273 , \2278 );
and \U$1937 ( \2280 , \2269 , \2278 );
or \U$1938 ( \2281 , \2274 , \2279 , \2280 );
and \U$1939 ( \2282 , \2264 , \2281 );
and \U$1940 ( \2283 , \2246 , \2281 );
or \U$1941 ( \2284 , \2265 , \2282 , \2283 );
xor \U$1942 ( \2285 , \2152 , \2156 );
xor \U$1943 ( \2286 , \2285 , \2161 );
xor \U$1944 ( \2287 , \2168 , \2172 );
xor \U$1945 ( \2288 , \2287 , \2175 );
and \U$1946 ( \2289 , \2286 , \2288 );
xor \U$1947 ( \2290 , \2133 , \2137 );
xor \U$1948 ( \2291 , \2290 , \2142 );
and \U$1949 ( \2292 , \2288 , \2291 );
and \U$1950 ( \2293 , \2286 , \2291 );
or \U$1951 ( \2294 , \2289 , \2292 , \2293 );
and \U$1952 ( \2295 , \2284 , \2294 );
and \U$1953 ( \2296 , \1596 , \406 );
and \U$1954 ( \2297 , \1588 , \404 );
nor \U$1955 ( \2298 , \2296 , \2297 );
xnor \U$1956 ( \2299 , \2298 , \413 );
and \U$1957 ( \2300 , \1844 , \422 );
and \U$1958 ( \2301 , \1839 , \420 );
nor \U$1959 ( \2302 , \2300 , \2301 );
xnor \U$1960 ( \2303 , \2302 , \429 );
and \U$1961 ( \2304 , \2299 , \2303 );
and \U$1962 ( \2305 , \2174 , \441 );
and \U$1963 ( \2306 , \2030 , \439 );
nor \U$1964 ( \2307 , \2305 , \2306 );
xnor \U$1965 ( \2308 , \2307 , \448 );
and \U$1966 ( \2309 , \2303 , \2308 );
and \U$1967 ( \2310 , \2299 , \2308 );
or \U$1968 ( \2311 , \2304 , \2309 , \2310 );
and \U$1969 ( \2312 , \1071 , \357 );
and \U$1970 ( \2313 , \983 , \355 );
nor \U$1971 ( \2314 , \2312 , \2313 );
xnor \U$1972 ( \2315 , \2314 , \364 );
and \U$1973 ( \2316 , \1181 , \373 );
and \U$1974 ( \2317 , \1176 , \371 );
nor \U$1975 ( \2318 , \2316 , \2317 );
xnor \U$1976 ( \2319 , \2318 , \380 );
and \U$1977 ( \2320 , \2315 , \2319 );
and \U$1978 ( \2321 , \1412 , \391 );
and \U$1979 ( \2322 , \1297 , \389 );
nor \U$1980 ( \2323 , \2321 , \2322 );
xnor \U$1981 ( \2324 , \2323 , \398 );
and \U$1982 ( \2325 , \2319 , \2324 );
and \U$1983 ( \2326 , \2315 , \2324 );
or \U$1984 ( \2327 , \2320 , \2325 , \2326 );
or \U$1985 ( \2328 , \2311 , \2327 );
and \U$1986 ( \2329 , \2294 , \2328 );
and \U$1987 ( \2330 , \2284 , \2328 );
or \U$1988 ( \2331 , \2295 , \2329 , \2330 );
xor \U$1989 ( \2332 , \1961 , \1965 );
xor \U$1990 ( \2333 , \2332 , \1970 );
xor \U$1991 ( \2334 , \2164 , \2178 );
xor \U$1992 ( \2335 , \2334 , \2181 );
and \U$1993 ( \2336 , \2333 , \2335 );
xor \U$1994 ( \2337 , \2187 , \2189 );
xor \U$1995 ( \2338 , \2337 , \2192 );
and \U$1996 ( \2339 , \2335 , \2338 );
and \U$1997 ( \2340 , \2333 , \2338 );
or \U$1998 ( \2341 , \2336 , \2339 , \2340 );
and \U$1999 ( \2342 , \2331 , \2341 );
xor \U$2000 ( \2343 , \1973 , \1989 );
xor \U$2001 ( \2344 , \2343 , \2006 );
and \U$2002 ( \2345 , \2341 , \2344 );
and \U$2003 ( \2346 , \2331 , \2344 );
or \U$2004 ( \2347 , \2342 , \2345 , \2346 );
xor \U$2005 ( \2348 , \2198 , \2208 );
xor \U$2006 ( \2349 , \2348 , \2211 );
and \U$2007 ( \2350 , \2347 , \2349 );
xor \U$2008 ( \2351 , \2216 , \2218 );
xor \U$2009 ( \2352 , \2351 , \2221 );
and \U$2010 ( \2353 , \2349 , \2352 );
and \U$2011 ( \2354 , \2347 , \2352 );
or \U$2012 ( \2355 , \2350 , \2353 , \2354 );
xor \U$2013 ( \2356 , \2214 , \2224 );
xor \U$2014 ( \2357 , \2356 , \2227 );
and \U$2015 ( \2358 , \2355 , \2357 );
xor \U$2016 ( \2359 , \2058 , \2068 );
xor \U$2017 ( \2360 , \2359 , \2071 );
and \U$2018 ( \2361 , \2357 , \2360 );
and \U$2019 ( \2362 , \2355 , \2360 );
or \U$2020 ( \2363 , \2358 , \2361 , \2362 );
and \U$2021 ( \2364 , \2230 , \2363 );
xor \U$2022 ( \2365 , \2074 , \2076 );
xor \U$2023 ( \2366 , \2365 , \2078 );
and \U$2024 ( \2367 , \2363 , \2366 );
and \U$2025 ( \2368 , \2230 , \2366 );
or \U$2026 ( \2369 , \2364 , \2367 , \2368 );
and \U$2027 ( \2370 , \2093 , \2369 );
xor \U$2028 ( \2371 , \2093 , \2369 );
xor \U$2029 ( \2372 , \2230 , \2363 );
xor \U$2030 ( \2373 , \2372 , \2366 );
and \U$2031 ( \2374 , \408 , \1623 );
and \U$2032 ( \2375 , \385 , \1621 );
nor \U$2033 ( \2376 , \2374 , \2375 );
xnor \U$2034 ( \2377 , \2376 , \1467 );
and \U$2035 ( \2378 , \424 , \1351 );
and \U$2036 ( \2379 , \400 , \1349 );
nor \U$2037 ( \2380 , \2378 , \2379 );
xnor \U$2038 ( \2381 , \2380 , \1238 );
and \U$2039 ( \2382 , \2377 , \2381 );
and \U$2040 ( \2383 , \443 , \1157 );
and \U$2041 ( \2384 , \416 , \1155 );
nor \U$2042 ( \2385 , \2383 , \2384 );
xnor \U$2043 ( \2386 , \2385 , \1021 );
and \U$2044 ( \2387 , \2381 , \2386 );
and \U$2045 ( \2388 , \2377 , \2386 );
or \U$2046 ( \2389 , \2382 , \2387 , \2388 );
xor \U$2047 ( \2390 , \1957 , \2247 );
xor \U$2048 ( \2391 , \2247 , \2248 );
not \U$2049 ( \2392 , \2391 );
and \U$2050 ( \2393 , \2390 , \2392 );
and \U$2051 ( \2394 , \359 , \2393 );
not \U$2052 ( \2395 , \2394 );
xnor \U$2053 ( \2396 , \2395 , \2251 );
and \U$2054 ( \2397 , \375 , \2097 );
and \U$2055 ( \2398 , \351 , \2095 );
nor \U$2056 ( \2399 , \2397 , \2398 );
xnor \U$2057 ( \2400 , \2399 , \1960 );
and \U$2058 ( \2401 , \2396 , \2400 );
and \U$2059 ( \2402 , \393 , \1891 );
and \U$2060 ( \2403 , \367 , \1889 );
nor \U$2061 ( \2404 , \2402 , \2403 );
xnor \U$2062 ( \2405 , \2404 , \1739 );
and \U$2063 ( \2406 , \2400 , \2405 );
and \U$2064 ( \2407 , \2396 , \2405 );
or \U$2065 ( \2408 , \2401 , \2406 , \2407 );
and \U$2066 ( \2409 , \2389 , \2408 );
and \U$2067 ( \2410 , \450 , \957 );
and \U$2068 ( \2411 , \435 , \955 );
nor \U$2069 ( \2412 , \2410 , \2411 );
xnor \U$2070 ( \2413 , \2412 , \879 );
and \U$2071 ( \2414 , \722 , \793 );
and \U$2072 ( \2415 , \661 , \791 );
nor \U$2073 ( \2416 , \2414 , \2415 );
xnor \U$2074 ( \2417 , \2416 , \699 );
and \U$2075 ( \2418 , \2413 , \2417 );
and \U$2076 ( \2419 , \983 , \624 );
and \U$2077 ( \2420 , \785 , \622 );
nor \U$2078 ( \2421 , \2419 , \2420 );
xnor \U$2079 ( \2422 , \2421 , \349 );
and \U$2080 ( \2423 , \2417 , \2422 );
and \U$2081 ( \2424 , \2413 , \2422 );
or \U$2082 ( \2425 , \2418 , \2423 , \2424 );
and \U$2083 ( \2426 , \2408 , \2425 );
and \U$2084 ( \2427 , \2389 , \2425 );
or \U$2085 ( \2428 , \2409 , \2426 , \2427 );
and \U$2086 ( \2429 , \1839 , \406 );
and \U$2087 ( \2430 , \1596 , \404 );
nor \U$2088 ( \2431 , \2429 , \2430 );
xnor \U$2089 ( \2432 , \2431 , \413 );
and \U$2090 ( \2433 , \2030 , \422 );
and \U$2091 ( \2434 , \1844 , \420 );
nor \U$2092 ( \2435 , \2433 , \2434 );
xnor \U$2093 ( \2436 , \2435 , \429 );
and \U$2094 ( \2437 , \2432 , \2436 );
buf \U$2095 ( \2438 , RIbb2caf0_93);
and \U$2096 ( \2439 , \2438 , \441 );
and \U$2097 ( \2440 , \2174 , \439 );
nor \U$2098 ( \2441 , \2439 , \2440 );
xnor \U$2099 ( \2442 , \2441 , \448 );
and \U$2100 ( \2443 , \2436 , \2442 );
and \U$2101 ( \2444 , \2432 , \2442 );
or \U$2102 ( \2445 , \2437 , \2443 , \2444 );
and \U$2103 ( \2446 , \1176 , \357 );
and \U$2104 ( \2447 , \1071 , \355 );
nor \U$2105 ( \2448 , \2446 , \2447 );
xnor \U$2106 ( \2449 , \2448 , \364 );
and \U$2107 ( \2450 , \1297 , \373 );
and \U$2108 ( \2451 , \1181 , \371 );
nor \U$2109 ( \2452 , \2450 , \2451 );
xnor \U$2110 ( \2453 , \2452 , \380 );
and \U$2111 ( \2454 , \2449 , \2453 );
and \U$2112 ( \2455 , \1588 , \391 );
and \U$2113 ( \2456 , \1412 , \389 );
nor \U$2114 ( \2457 , \2455 , \2456 );
xnor \U$2115 ( \2458 , \2457 , \398 );
and \U$2116 ( \2459 , \2453 , \2458 );
and \U$2117 ( \2460 , \2449 , \2458 );
or \U$2118 ( \2461 , \2454 , \2459 , \2460 );
and \U$2119 ( \2462 , \2445 , \2461 );
buf \U$2120 ( \2463 , RIbb2ca78_94);
and \U$2121 ( \2464 , \2463 , \436 );
buf \U$2122 ( \2465 , \2464 );
and \U$2123 ( \2466 , \2461 , \2465 );
and \U$2124 ( \2467 , \2445 , \2465 );
or \U$2125 ( \2468 , \2462 , \2466 , \2467 );
and \U$2126 ( \2469 , \2428 , \2468 );
and \U$2127 ( \2470 , \2438 , \436 );
xor \U$2128 ( \2471 , \2299 , \2303 );
xor \U$2129 ( \2472 , \2471 , \2308 );
and \U$2130 ( \2473 , \2470 , \2472 );
xor \U$2131 ( \2474 , \2315 , \2319 );
xor \U$2132 ( \2475 , \2474 , \2324 );
and \U$2133 ( \2476 , \2472 , \2475 );
and \U$2134 ( \2477 , \2470 , \2475 );
or \U$2135 ( \2478 , \2473 , \2476 , \2477 );
and \U$2136 ( \2479 , \2468 , \2478 );
and \U$2137 ( \2480 , \2428 , \2478 );
or \U$2138 ( \2481 , \2469 , \2479 , \2480 );
xor \U$2139 ( \2482 , \2234 , \2238 );
xor \U$2140 ( \2483 , \2482 , \2243 );
xor \U$2141 ( \2484 , \2252 , \2256 );
xor \U$2142 ( \2485 , \2484 , \2261 );
and \U$2143 ( \2486 , \2483 , \2485 );
xor \U$2144 ( \2487 , \2269 , \2273 );
xor \U$2145 ( \2488 , \2487 , \2278 );
and \U$2146 ( \2489 , \2485 , \2488 );
and \U$2147 ( \2490 , \2483 , \2488 );
or \U$2148 ( \2491 , \2486 , \2489 , \2490 );
xor \U$2149 ( \2492 , \2100 , \2104 );
xor \U$2150 ( \2493 , \2492 , \2109 );
and \U$2151 ( \2494 , \2491 , \2493 );
xor \U$2152 ( \2495 , \2116 , \2120 );
xor \U$2153 ( \2496 , \2495 , \2125 );
and \U$2154 ( \2497 , \2493 , \2496 );
and \U$2155 ( \2498 , \2491 , \2496 );
or \U$2156 ( \2499 , \2494 , \2497 , \2498 );
and \U$2157 ( \2500 , \2481 , \2499 );
xor \U$2158 ( \2501 , \2246 , \2264 );
xor \U$2159 ( \2502 , \2501 , \2281 );
xor \U$2160 ( \2503 , \2286 , \2288 );
xor \U$2161 ( \2504 , \2503 , \2291 );
and \U$2162 ( \2505 , \2502 , \2504 );
xnor \U$2163 ( \2506 , \2311 , \2327 );
and \U$2164 ( \2507 , \2504 , \2506 );
and \U$2165 ( \2508 , \2502 , \2506 );
or \U$2166 ( \2509 , \2505 , \2507 , \2508 );
and \U$2167 ( \2510 , \2499 , \2509 );
and \U$2168 ( \2511 , \2481 , \2509 );
or \U$2169 ( \2512 , \2500 , \2510 , \2511 );
xor \U$2170 ( \2513 , \2112 , \2128 );
xor \U$2171 ( \2514 , \2513 , \2145 );
xor \U$2172 ( \2515 , \2284 , \2294 );
xor \U$2173 ( \2516 , \2515 , \2328 );
and \U$2174 ( \2517 , \2514 , \2516 );
xor \U$2175 ( \2518 , \2333 , \2335 );
xor \U$2176 ( \2519 , \2518 , \2338 );
and \U$2177 ( \2520 , \2516 , \2519 );
and \U$2178 ( \2521 , \2514 , \2519 );
or \U$2179 ( \2522 , \2517 , \2520 , \2521 );
and \U$2180 ( \2523 , \2512 , \2522 );
xor \U$2181 ( \2524 , \2200 , \2202 );
xor \U$2182 ( \2525 , \2524 , \2205 );
and \U$2183 ( \2526 , \2522 , \2525 );
and \U$2184 ( \2527 , \2512 , \2525 );
or \U$2185 ( \2528 , \2523 , \2526 , \2527 );
xor \U$2186 ( \2529 , \2148 , \2184 );
xor \U$2187 ( \2530 , \2529 , \2195 );
xor \U$2188 ( \2531 , \2331 , \2341 );
xor \U$2189 ( \2532 , \2531 , \2344 );
and \U$2190 ( \2533 , \2530 , \2532 );
and \U$2191 ( \2534 , \2528 , \2533 );
xor \U$2192 ( \2535 , \2347 , \2349 );
xor \U$2193 ( \2536 , \2535 , \2352 );
and \U$2194 ( \2537 , \2533 , \2536 );
and \U$2195 ( \2538 , \2528 , \2536 );
or \U$2196 ( \2539 , \2534 , \2537 , \2538 );
xor \U$2197 ( \2540 , \2355 , \2357 );
xor \U$2198 ( \2541 , \2540 , \2360 );
and \U$2199 ( \2542 , \2539 , \2541 );
and \U$2200 ( \2543 , \2373 , \2542 );
xor \U$2201 ( \2544 , \2373 , \2542 );
xor \U$2202 ( \2545 , \2539 , \2541 );
and \U$2203 ( \2546 , \435 , \1157 );
and \U$2204 ( \2547 , \443 , \1155 );
nor \U$2205 ( \2548 , \2546 , \2547 );
xnor \U$2206 ( \2549 , \2548 , \1021 );
and \U$2207 ( \2550 , \661 , \957 );
and \U$2208 ( \2551 , \450 , \955 );
nor \U$2209 ( \2552 , \2550 , \2551 );
xnor \U$2210 ( \2553 , \2552 , \879 );
and \U$2211 ( \2554 , \2549 , \2553 );
and \U$2212 ( \2555 , \785 , \793 );
and \U$2213 ( \2556 , \722 , \791 );
nor \U$2214 ( \2557 , \2555 , \2556 );
xnor \U$2215 ( \2558 , \2557 , \699 );
and \U$2216 ( \2559 , \2553 , \2558 );
and \U$2217 ( \2560 , \2549 , \2558 );
or \U$2218 ( \2561 , \2554 , \2559 , \2560 );
buf \U$2219 ( \2562 , RIbb2e788_32);
buf \U$2220 ( \2563 , RIbb2e710_33);
and \U$2221 ( \2564 , \2562 , \2563 );
not \U$2222 ( \2565 , \2564 );
and \U$2223 ( \2566 , \2248 , \2565 );
not \U$2224 ( \2567 , \2566 );
and \U$2225 ( \2568 , \351 , \2393 );
and \U$2226 ( \2569 , \359 , \2391 );
nor \U$2227 ( \2570 , \2568 , \2569 );
xnor \U$2228 ( \2571 , \2570 , \2251 );
and \U$2229 ( \2572 , \2567 , \2571 );
and \U$2230 ( \2573 , \367 , \2097 );
and \U$2231 ( \2574 , \375 , \2095 );
nor \U$2232 ( \2575 , \2573 , \2574 );
xnor \U$2233 ( \2576 , \2575 , \1960 );
and \U$2234 ( \2577 , \2571 , \2576 );
and \U$2235 ( \2578 , \2567 , \2576 );
or \U$2236 ( \2579 , \2572 , \2577 , \2578 );
and \U$2237 ( \2580 , \2561 , \2579 );
and \U$2238 ( \2581 , \385 , \1891 );
and \U$2239 ( \2582 , \393 , \1889 );
nor \U$2240 ( \2583 , \2581 , \2582 );
xnor \U$2241 ( \2584 , \2583 , \1739 );
and \U$2242 ( \2585 , \400 , \1623 );
and \U$2243 ( \2586 , \408 , \1621 );
nor \U$2244 ( \2587 , \2585 , \2586 );
xnor \U$2245 ( \2588 , \2587 , \1467 );
and \U$2246 ( \2589 , \2584 , \2588 );
and \U$2247 ( \2590 , \416 , \1351 );
and \U$2248 ( \2591 , \424 , \1349 );
nor \U$2249 ( \2592 , \2590 , \2591 );
xnor \U$2250 ( \2593 , \2592 , \1238 );
and \U$2251 ( \2594 , \2588 , \2593 );
and \U$2252 ( \2595 , \2584 , \2593 );
or \U$2253 ( \2596 , \2589 , \2594 , \2595 );
and \U$2254 ( \2597 , \2579 , \2596 );
and \U$2255 ( \2598 , \2561 , \2596 );
or \U$2256 ( \2599 , \2580 , \2597 , \2598 );
and \U$2257 ( \2600 , \1596 , \391 );
and \U$2258 ( \2601 , \1588 , \389 );
nor \U$2259 ( \2602 , \2600 , \2601 );
xnor \U$2260 ( \2603 , \2602 , \398 );
and \U$2261 ( \2604 , \1844 , \406 );
and \U$2262 ( \2605 , \1839 , \404 );
nor \U$2263 ( \2606 , \2604 , \2605 );
xnor \U$2264 ( \2607 , \2606 , \413 );
and \U$2265 ( \2608 , \2603 , \2607 );
and \U$2266 ( \2609 , \2174 , \422 );
and \U$2267 ( \2610 , \2030 , \420 );
nor \U$2268 ( \2611 , \2609 , \2610 );
xnor \U$2269 ( \2612 , \2611 , \429 );
and \U$2270 ( \2613 , \2607 , \2612 );
and \U$2271 ( \2614 , \2603 , \2612 );
or \U$2272 ( \2615 , \2608 , \2613 , \2614 );
and \U$2273 ( \2616 , \1071 , \624 );
and \U$2274 ( \2617 , \983 , \622 );
nor \U$2275 ( \2618 , \2616 , \2617 );
xnor \U$2276 ( \2619 , \2618 , \349 );
and \U$2277 ( \2620 , \1181 , \357 );
and \U$2278 ( \2621 , \1176 , \355 );
nor \U$2279 ( \2622 , \2620 , \2621 );
xnor \U$2280 ( \2623 , \2622 , \364 );
and \U$2281 ( \2624 , \2619 , \2623 );
and \U$2282 ( \2625 , \1412 , \373 );
and \U$2283 ( \2626 , \1297 , \371 );
nor \U$2284 ( \2627 , \2625 , \2626 );
xnor \U$2285 ( \2628 , \2627 , \380 );
and \U$2286 ( \2629 , \2623 , \2628 );
and \U$2287 ( \2630 , \2619 , \2628 );
or \U$2288 ( \2631 , \2624 , \2629 , \2630 );
and \U$2289 ( \2632 , \2615 , \2631 );
and \U$2290 ( \2633 , \2463 , \441 );
and \U$2291 ( \2634 , \2438 , \439 );
nor \U$2292 ( \2635 , \2633 , \2634 );
xnor \U$2293 ( \2636 , \2635 , \448 );
buf \U$2294 ( \2637 , RIbb2ca00_95);
and \U$2295 ( \2638 , \2637 , \436 );
and \U$2296 ( \2639 , \2636 , \2638 );
and \U$2297 ( \2640 , \2631 , \2639 );
and \U$2298 ( \2641 , \2615 , \2639 );
or \U$2299 ( \2642 , \2632 , \2640 , \2641 );
and \U$2300 ( \2643 , \2599 , \2642 );
xor \U$2301 ( \2644 , \2432 , \2436 );
xor \U$2302 ( \2645 , \2644 , \2442 );
xor \U$2303 ( \2646 , \2449 , \2453 );
xor \U$2304 ( \2647 , \2646 , \2458 );
and \U$2305 ( \2648 , \2645 , \2647 );
not \U$2306 ( \2649 , \2464 );
and \U$2307 ( \2650 , \2647 , \2649 );
and \U$2308 ( \2651 , \2645 , \2649 );
or \U$2309 ( \2652 , \2648 , \2650 , \2651 );
and \U$2310 ( \2653 , \2642 , \2652 );
and \U$2311 ( \2654 , \2599 , \2652 );
or \U$2312 ( \2655 , \2643 , \2653 , \2654 );
xor \U$2313 ( \2656 , \2377 , \2381 );
xor \U$2314 ( \2657 , \2656 , \2386 );
xor \U$2315 ( \2658 , \2396 , \2400 );
xor \U$2316 ( \2659 , \2658 , \2405 );
and \U$2317 ( \2660 , \2657 , \2659 );
xor \U$2318 ( \2661 , \2413 , \2417 );
xor \U$2319 ( \2662 , \2661 , \2422 );
and \U$2320 ( \2663 , \2659 , \2662 );
and \U$2321 ( \2664 , \2657 , \2662 );
or \U$2322 ( \2665 , \2660 , \2663 , \2664 );
xor \U$2323 ( \2666 , \2483 , \2485 );
xor \U$2324 ( \2667 , \2666 , \2488 );
and \U$2325 ( \2668 , \2665 , \2667 );
xor \U$2326 ( \2669 , \2470 , \2472 );
xor \U$2327 ( \2670 , \2669 , \2475 );
and \U$2328 ( \2671 , \2667 , \2670 );
and \U$2329 ( \2672 , \2665 , \2670 );
or \U$2330 ( \2673 , \2668 , \2671 , \2672 );
and \U$2331 ( \2674 , \2655 , \2673 );
xor \U$2332 ( \2675 , \2389 , \2408 );
xor \U$2333 ( \2676 , \2675 , \2425 );
xor \U$2334 ( \2677 , \2445 , \2461 );
xor \U$2335 ( \2678 , \2677 , \2465 );
and \U$2336 ( \2679 , \2676 , \2678 );
and \U$2337 ( \2680 , \2673 , \2679 );
and \U$2338 ( \2681 , \2655 , \2679 );
or \U$2339 ( \2682 , \2674 , \2680 , \2681 );
xor \U$2340 ( \2683 , \2428 , \2468 );
xor \U$2341 ( \2684 , \2683 , \2478 );
xor \U$2342 ( \2685 , \2491 , \2493 );
xor \U$2343 ( \2686 , \2685 , \2496 );
and \U$2344 ( \2687 , \2684 , \2686 );
xor \U$2345 ( \2688 , \2502 , \2504 );
xor \U$2346 ( \2689 , \2688 , \2506 );
and \U$2347 ( \2690 , \2686 , \2689 );
and \U$2348 ( \2691 , \2684 , \2689 );
or \U$2349 ( \2692 , \2687 , \2690 , \2691 );
and \U$2350 ( \2693 , \2682 , \2692 );
xor \U$2351 ( \2694 , \2514 , \2516 );
xor \U$2352 ( \2695 , \2694 , \2519 );
and \U$2353 ( \2696 , \2692 , \2695 );
and \U$2354 ( \2697 , \2682 , \2695 );
or \U$2355 ( \2698 , \2693 , \2696 , \2697 );
xor \U$2356 ( \2699 , \2512 , \2522 );
xor \U$2357 ( \2700 , \2699 , \2525 );
and \U$2358 ( \2701 , \2698 , \2700 );
xor \U$2359 ( \2702 , \2530 , \2532 );
and \U$2360 ( \2703 , \2700 , \2702 );
and \U$2361 ( \2704 , \2698 , \2702 );
or \U$2362 ( \2705 , \2701 , \2703 , \2704 );
xor \U$2363 ( \2706 , \2528 , \2533 );
xor \U$2364 ( \2707 , \2706 , \2536 );
and \U$2365 ( \2708 , \2705 , \2707 );
and \U$2366 ( \2709 , \2545 , \2708 );
xor \U$2367 ( \2710 , \2545 , \2708 );
xor \U$2368 ( \2711 , \2705 , \2707 );
xor \U$2369 ( \2712 , \2248 , \2562 );
xor \U$2370 ( \2713 , \2562 , \2563 );
not \U$2371 ( \2714 , \2713 );
and \U$2372 ( \2715 , \2712 , \2714 );
and \U$2373 ( \2716 , \359 , \2715 );
not \U$2374 ( \2717 , \2716 );
xnor \U$2375 ( \2718 , \2717 , \2566 );
and \U$2376 ( \2719 , \375 , \2393 );
and \U$2377 ( \2720 , \351 , \2391 );
nor \U$2378 ( \2721 , \2719 , \2720 );
xnor \U$2379 ( \2722 , \2721 , \2251 );
and \U$2380 ( \2723 , \2718 , \2722 );
and \U$2381 ( \2724 , \393 , \2097 );
and \U$2382 ( \2725 , \367 , \2095 );
nor \U$2383 ( \2726 , \2724 , \2725 );
xnor \U$2384 ( \2727 , \2726 , \1960 );
and \U$2385 ( \2728 , \2722 , \2727 );
and \U$2386 ( \2729 , \2718 , \2727 );
or \U$2387 ( \2730 , \2723 , \2728 , \2729 );
and \U$2388 ( \2731 , \450 , \1157 );
and \U$2389 ( \2732 , \435 , \1155 );
nor \U$2390 ( \2733 , \2731 , \2732 );
xnor \U$2391 ( \2734 , \2733 , \1021 );
and \U$2392 ( \2735 , \722 , \957 );
and \U$2393 ( \2736 , \661 , \955 );
nor \U$2394 ( \2737 , \2735 , \2736 );
xnor \U$2395 ( \2738 , \2737 , \879 );
and \U$2396 ( \2739 , \2734 , \2738 );
and \U$2397 ( \2740 , \983 , \793 );
and \U$2398 ( \2741 , \785 , \791 );
nor \U$2399 ( \2742 , \2740 , \2741 );
xnor \U$2400 ( \2743 , \2742 , \699 );
and \U$2401 ( \2744 , \2738 , \2743 );
and \U$2402 ( \2745 , \2734 , \2743 );
or \U$2403 ( \2746 , \2739 , \2744 , \2745 );
and \U$2404 ( \2747 , \2730 , \2746 );
and \U$2405 ( \2748 , \408 , \1891 );
and \U$2406 ( \2749 , \385 , \1889 );
nor \U$2407 ( \2750 , \2748 , \2749 );
xnor \U$2408 ( \2751 , \2750 , \1739 );
and \U$2409 ( \2752 , \424 , \1623 );
and \U$2410 ( \2753 , \400 , \1621 );
nor \U$2411 ( \2754 , \2752 , \2753 );
xnor \U$2412 ( \2755 , \2754 , \1467 );
and \U$2413 ( \2756 , \2751 , \2755 );
and \U$2414 ( \2757 , \443 , \1351 );
and \U$2415 ( \2758 , \416 , \1349 );
nor \U$2416 ( \2759 , \2757 , \2758 );
xnor \U$2417 ( \2760 , \2759 , \1238 );
and \U$2418 ( \2761 , \2755 , \2760 );
and \U$2419 ( \2762 , \2751 , \2760 );
or \U$2420 ( \2763 , \2756 , \2761 , \2762 );
and \U$2421 ( \2764 , \2746 , \2763 );
and \U$2422 ( \2765 , \2730 , \2763 );
or \U$2423 ( \2766 , \2747 , \2764 , \2765 );
and \U$2424 ( \2767 , \1839 , \391 );
and \U$2425 ( \2768 , \1596 , \389 );
nor \U$2426 ( \2769 , \2767 , \2768 );
xnor \U$2427 ( \2770 , \2769 , \398 );
and \U$2428 ( \2771 , \2030 , \406 );
and \U$2429 ( \2772 , \1844 , \404 );
nor \U$2430 ( \2773 , \2771 , \2772 );
xnor \U$2431 ( \2774 , \2773 , \413 );
and \U$2432 ( \2775 , \2770 , \2774 );
and \U$2433 ( \2776 , \2438 , \422 );
and \U$2434 ( \2777 , \2174 , \420 );
nor \U$2435 ( \2778 , \2776 , \2777 );
xnor \U$2436 ( \2779 , \2778 , \429 );
and \U$2437 ( \2780 , \2774 , \2779 );
and \U$2438 ( \2781 , \2770 , \2779 );
or \U$2439 ( \2782 , \2775 , \2780 , \2781 );
and \U$2440 ( \2783 , \1176 , \624 );
and \U$2441 ( \2784 , \1071 , \622 );
nor \U$2442 ( \2785 , \2783 , \2784 );
xnor \U$2443 ( \2786 , \2785 , \349 );
and \U$2444 ( \2787 , \1297 , \357 );
and \U$2445 ( \2788 , \1181 , \355 );
nor \U$2446 ( \2789 , \2787 , \2788 );
xnor \U$2447 ( \2790 , \2789 , \364 );
and \U$2448 ( \2791 , \2786 , \2790 );
and \U$2449 ( \2792 , \1588 , \373 );
and \U$2450 ( \2793 , \1412 , \371 );
nor \U$2451 ( \2794 , \2792 , \2793 );
xnor \U$2452 ( \2795 , \2794 , \380 );
and \U$2453 ( \2796 , \2790 , \2795 );
and \U$2454 ( \2797 , \2786 , \2795 );
or \U$2455 ( \2798 , \2791 , \2796 , \2797 );
and \U$2456 ( \2799 , \2782 , \2798 );
and \U$2457 ( \2800 , \2637 , \441 );
and \U$2458 ( \2801 , \2463 , \439 );
nor \U$2459 ( \2802 , \2800 , \2801 );
xnor \U$2460 ( \2803 , \2802 , \448 );
buf \U$2461 ( \2804 , RIbb2c988_96);
and \U$2462 ( \2805 , \2804 , \436 );
or \U$2463 ( \2806 , \2803 , \2805 );
and \U$2464 ( \2807 , \2798 , \2806 );
and \U$2465 ( \2808 , \2782 , \2806 );
or \U$2466 ( \2809 , \2799 , \2807 , \2808 );
and \U$2467 ( \2810 , \2766 , \2809 );
xor \U$2468 ( \2811 , \2603 , \2607 );
xor \U$2469 ( \2812 , \2811 , \2612 );
xor \U$2470 ( \2813 , \2619 , \2623 );
xor \U$2471 ( \2814 , \2813 , \2628 );
and \U$2472 ( \2815 , \2812 , \2814 );
xor \U$2473 ( \2816 , \2636 , \2638 );
and \U$2474 ( \2817 , \2814 , \2816 );
and \U$2475 ( \2818 , \2812 , \2816 );
or \U$2476 ( \2819 , \2815 , \2817 , \2818 );
and \U$2477 ( \2820 , \2809 , \2819 );
and \U$2478 ( \2821 , \2766 , \2819 );
or \U$2479 ( \2822 , \2810 , \2820 , \2821 );
xor \U$2480 ( \2823 , \2549 , \2553 );
xor \U$2481 ( \2824 , \2823 , \2558 );
xor \U$2482 ( \2825 , \2567 , \2571 );
xor \U$2483 ( \2826 , \2825 , \2576 );
and \U$2484 ( \2827 , \2824 , \2826 );
xor \U$2485 ( \2828 , \2584 , \2588 );
xor \U$2486 ( \2829 , \2828 , \2593 );
and \U$2487 ( \2830 , \2826 , \2829 );
and \U$2488 ( \2831 , \2824 , \2829 );
or \U$2489 ( \2832 , \2827 , \2830 , \2831 );
xor \U$2490 ( \2833 , \2657 , \2659 );
xor \U$2491 ( \2834 , \2833 , \2662 );
and \U$2492 ( \2835 , \2832 , \2834 );
xor \U$2493 ( \2836 , \2645 , \2647 );
xor \U$2494 ( \2837 , \2836 , \2649 );
and \U$2495 ( \2838 , \2834 , \2837 );
and \U$2496 ( \2839 , \2832 , \2837 );
or \U$2497 ( \2840 , \2835 , \2838 , \2839 );
and \U$2498 ( \2841 , \2822 , \2840 );
xor \U$2499 ( \2842 , \2561 , \2579 );
xor \U$2500 ( \2843 , \2842 , \2596 );
xor \U$2501 ( \2844 , \2615 , \2631 );
xor \U$2502 ( \2845 , \2844 , \2639 );
and \U$2503 ( \2846 , \2843 , \2845 );
and \U$2504 ( \2847 , \2840 , \2846 );
and \U$2505 ( \2848 , \2822 , \2846 );
or \U$2506 ( \2849 , \2841 , \2847 , \2848 );
xor \U$2507 ( \2850 , \2599 , \2642 );
xor \U$2508 ( \2851 , \2850 , \2652 );
xor \U$2509 ( \2852 , \2665 , \2667 );
xor \U$2510 ( \2853 , \2852 , \2670 );
and \U$2511 ( \2854 , \2851 , \2853 );
xor \U$2512 ( \2855 , \2676 , \2678 );
and \U$2513 ( \2856 , \2853 , \2855 );
and \U$2514 ( \2857 , \2851 , \2855 );
or \U$2515 ( \2858 , \2854 , \2856 , \2857 );
and \U$2516 ( \2859 , \2849 , \2858 );
xor \U$2517 ( \2860 , \2684 , \2686 );
xor \U$2518 ( \2861 , \2860 , \2689 );
and \U$2519 ( \2862 , \2858 , \2861 );
and \U$2520 ( \2863 , \2849 , \2861 );
or \U$2521 ( \2864 , \2859 , \2862 , \2863 );
xor \U$2522 ( \2865 , \2481 , \2499 );
xor \U$2523 ( \2866 , \2865 , \2509 );
and \U$2524 ( \2867 , \2864 , \2866 );
xor \U$2525 ( \2868 , \2682 , \2692 );
xor \U$2526 ( \2869 , \2868 , \2695 );
and \U$2527 ( \2870 , \2866 , \2869 );
and \U$2528 ( \2871 , \2864 , \2869 );
or \U$2529 ( \2872 , \2867 , \2870 , \2871 );
xor \U$2530 ( \2873 , \2698 , \2700 );
xor \U$2531 ( \2874 , \2873 , \2702 );
and \U$2532 ( \2875 , \2872 , \2874 );
and \U$2533 ( \2876 , \2711 , \2875 );
xor \U$2534 ( \2877 , \2711 , \2875 );
xor \U$2535 ( \2878 , \2872 , \2874 );
and \U$2536 ( \2879 , \385 , \2097 );
and \U$2537 ( \2880 , \393 , \2095 );
nor \U$2538 ( \2881 , \2879 , \2880 );
xnor \U$2539 ( \2882 , \2881 , \1960 );
and \U$2540 ( \2883 , \400 , \1891 );
and \U$2541 ( \2884 , \408 , \1889 );
nor \U$2542 ( \2885 , \2883 , \2884 );
xnor \U$2543 ( \2886 , \2885 , \1739 );
and \U$2544 ( \2887 , \2882 , \2886 );
and \U$2545 ( \2888 , \416 , \1623 );
and \U$2546 ( \2889 , \424 , \1621 );
nor \U$2547 ( \2890 , \2888 , \2889 );
xnor \U$2548 ( \2891 , \2890 , \1467 );
and \U$2549 ( \2892 , \2886 , \2891 );
and \U$2550 ( \2893 , \2882 , \2891 );
or \U$2551 ( \2894 , \2887 , \2892 , \2893 );
and \U$2552 ( \2895 , \435 , \1351 );
and \U$2553 ( \2896 , \443 , \1349 );
nor \U$2554 ( \2897 , \2895 , \2896 );
xnor \U$2555 ( \2898 , \2897 , \1238 );
and \U$2556 ( \2899 , \661 , \1157 );
and \U$2557 ( \2900 , \450 , \1155 );
nor \U$2558 ( \2901 , \2899 , \2900 );
xnor \U$2559 ( \2902 , \2901 , \1021 );
and \U$2560 ( \2903 , \2898 , \2902 );
and \U$2561 ( \2904 , \785 , \957 );
and \U$2562 ( \2905 , \722 , \955 );
nor \U$2563 ( \2906 , \2904 , \2905 );
xnor \U$2564 ( \2907 , \2906 , \879 );
and \U$2565 ( \2908 , \2902 , \2907 );
and \U$2566 ( \2909 , \2898 , \2907 );
or \U$2567 ( \2910 , \2903 , \2908 , \2909 );
and \U$2568 ( \2911 , \2894 , \2910 );
buf \U$2569 ( \2912 , RIbb2e698_34);
buf \U$2570 ( \2913 , RIbb2e620_35);
and \U$2571 ( \2914 , \2912 , \2913 );
not \U$2572 ( \2915 , \2914 );
and \U$2573 ( \2916 , \2563 , \2915 );
not \U$2574 ( \2917 , \2916 );
and \U$2575 ( \2918 , \351 , \2715 );
and \U$2576 ( \2919 , \359 , \2713 );
nor \U$2577 ( \2920 , \2918 , \2919 );
xnor \U$2578 ( \2921 , \2920 , \2566 );
and \U$2579 ( \2922 , \2917 , \2921 );
and \U$2580 ( \2923 , \367 , \2393 );
and \U$2581 ( \2924 , \375 , \2391 );
nor \U$2582 ( \2925 , \2923 , \2924 );
xnor \U$2583 ( \2926 , \2925 , \2251 );
and \U$2584 ( \2927 , \2921 , \2926 );
and \U$2585 ( \2928 , \2917 , \2926 );
or \U$2586 ( \2929 , \2922 , \2927 , \2928 );
and \U$2587 ( \2930 , \2910 , \2929 );
and \U$2588 ( \2931 , \2894 , \2929 );
or \U$2589 ( \2932 , \2911 , \2930 , \2931 );
and \U$2590 ( \2933 , \2463 , \422 );
and \U$2591 ( \2934 , \2438 , \420 );
nor \U$2592 ( \2935 , \2933 , \2934 );
xnor \U$2593 ( \2936 , \2935 , \429 );
and \U$2594 ( \2937 , \2804 , \441 );
and \U$2595 ( \2938 , \2637 , \439 );
nor \U$2596 ( \2939 , \2937 , \2938 );
xnor \U$2597 ( \2940 , \2939 , \448 );
and \U$2598 ( \2941 , \2936 , \2940 );
buf \U$2599 ( \2942 , RIbb2c910_97);
and \U$2600 ( \2943 , \2942 , \436 );
and \U$2601 ( \2944 , \2940 , \2943 );
and \U$2602 ( \2945 , \2936 , \2943 );
or \U$2603 ( \2946 , \2941 , \2944 , \2945 );
and \U$2604 ( \2947 , \1596 , \373 );
and \U$2605 ( \2948 , \1588 , \371 );
nor \U$2606 ( \2949 , \2947 , \2948 );
xnor \U$2607 ( \2950 , \2949 , \380 );
and \U$2608 ( \2951 , \1844 , \391 );
and \U$2609 ( \2952 , \1839 , \389 );
nor \U$2610 ( \2953 , \2951 , \2952 );
xnor \U$2611 ( \2954 , \2953 , \398 );
and \U$2612 ( \2955 , \2950 , \2954 );
and \U$2613 ( \2956 , \2174 , \406 );
and \U$2614 ( \2957 , \2030 , \404 );
nor \U$2615 ( \2958 , \2956 , \2957 );
xnor \U$2616 ( \2959 , \2958 , \413 );
and \U$2617 ( \2960 , \2954 , \2959 );
and \U$2618 ( \2961 , \2950 , \2959 );
or \U$2619 ( \2962 , \2955 , \2960 , \2961 );
and \U$2620 ( \2963 , \2946 , \2962 );
and \U$2621 ( \2964 , \1071 , \793 );
and \U$2622 ( \2965 , \983 , \791 );
nor \U$2623 ( \2966 , \2964 , \2965 );
xnor \U$2624 ( \2967 , \2966 , \699 );
and \U$2625 ( \2968 , \1181 , \624 );
and \U$2626 ( \2969 , \1176 , \622 );
nor \U$2627 ( \2970 , \2968 , \2969 );
xnor \U$2628 ( \2971 , \2970 , \349 );
and \U$2629 ( \2972 , \2967 , \2971 );
and \U$2630 ( \2973 , \1412 , \357 );
and \U$2631 ( \2974 , \1297 , \355 );
nor \U$2632 ( \2975 , \2973 , \2974 );
xnor \U$2633 ( \2976 , \2975 , \364 );
and \U$2634 ( \2977 , \2971 , \2976 );
and \U$2635 ( \2978 , \2967 , \2976 );
or \U$2636 ( \2979 , \2972 , \2977 , \2978 );
and \U$2637 ( \2980 , \2962 , \2979 );
and \U$2638 ( \2981 , \2946 , \2979 );
or \U$2639 ( \2982 , \2963 , \2980 , \2981 );
and \U$2640 ( \2983 , \2932 , \2982 );
xor \U$2641 ( \2984 , \2770 , \2774 );
xor \U$2642 ( \2985 , \2984 , \2779 );
xor \U$2643 ( \2986 , \2786 , \2790 );
xor \U$2644 ( \2987 , \2986 , \2795 );
and \U$2645 ( \2988 , \2985 , \2987 );
xnor \U$2646 ( \2989 , \2803 , \2805 );
and \U$2647 ( \2990 , \2987 , \2989 );
and \U$2648 ( \2991 , \2985 , \2989 );
or \U$2649 ( \2992 , \2988 , \2990 , \2991 );
and \U$2650 ( \2993 , \2982 , \2992 );
and \U$2651 ( \2994 , \2932 , \2992 );
or \U$2652 ( \2995 , \2983 , \2993 , \2994 );
xor \U$2653 ( \2996 , \2718 , \2722 );
xor \U$2654 ( \2997 , \2996 , \2727 );
xor \U$2655 ( \2998 , \2734 , \2738 );
xor \U$2656 ( \2999 , \2998 , \2743 );
and \U$2657 ( \3000 , \2997 , \2999 );
xor \U$2658 ( \3001 , \2751 , \2755 );
xor \U$2659 ( \3002 , \3001 , \2760 );
and \U$2660 ( \3003 , \2999 , \3002 );
and \U$2661 ( \3004 , \2997 , \3002 );
or \U$2662 ( \3005 , \3000 , \3003 , \3004 );
xor \U$2663 ( \3006 , \2824 , \2826 );
xor \U$2664 ( \3007 , \3006 , \2829 );
and \U$2665 ( \3008 , \3005 , \3007 );
xor \U$2666 ( \3009 , \2812 , \2814 );
xor \U$2667 ( \3010 , \3009 , \2816 );
and \U$2668 ( \3011 , \3007 , \3010 );
and \U$2669 ( \3012 , \3005 , \3010 );
or \U$2670 ( \3013 , \3008 , \3011 , \3012 );
and \U$2671 ( \3014 , \2995 , \3013 );
xor \U$2672 ( \3015 , \2730 , \2746 );
xor \U$2673 ( \3016 , \3015 , \2763 );
xor \U$2674 ( \3017 , \2782 , \2798 );
xor \U$2675 ( \3018 , \3017 , \2806 );
and \U$2676 ( \3019 , \3016 , \3018 );
and \U$2677 ( \3020 , \3013 , \3019 );
and \U$2678 ( \3021 , \2995 , \3019 );
or \U$2679 ( \3022 , \3014 , \3020 , \3021 );
xor \U$2680 ( \3023 , \2766 , \2809 );
xor \U$2681 ( \3024 , \3023 , \2819 );
xor \U$2682 ( \3025 , \2832 , \2834 );
xor \U$2683 ( \3026 , \3025 , \2837 );
and \U$2684 ( \3027 , \3024 , \3026 );
xor \U$2685 ( \3028 , \2843 , \2845 );
and \U$2686 ( \3029 , \3026 , \3028 );
and \U$2687 ( \3030 , \3024 , \3028 );
or \U$2688 ( \3031 , \3027 , \3029 , \3030 );
and \U$2689 ( \3032 , \3022 , \3031 );
xor \U$2690 ( \3033 , \2851 , \2853 );
xor \U$2691 ( \3034 , \3033 , \2855 );
and \U$2692 ( \3035 , \3031 , \3034 );
and \U$2693 ( \3036 , \3022 , \3034 );
or \U$2694 ( \3037 , \3032 , \3035 , \3036 );
xor \U$2695 ( \3038 , \2655 , \2673 );
xor \U$2696 ( \3039 , \3038 , \2679 );
and \U$2697 ( \3040 , \3037 , \3039 );
xor \U$2698 ( \3041 , \2849 , \2858 );
xor \U$2699 ( \3042 , \3041 , \2861 );
and \U$2700 ( \3043 , \3039 , \3042 );
and \U$2701 ( \3044 , \3037 , \3042 );
or \U$2702 ( \3045 , \3040 , \3043 , \3044 );
xor \U$2703 ( \3046 , \2864 , \2866 );
xor \U$2704 ( \3047 , \3046 , \2869 );
and \U$2705 ( \3048 , \3045 , \3047 );
and \U$2706 ( \3049 , \2878 , \3048 );
xor \U$2707 ( \3050 , \2878 , \3048 );
xor \U$2708 ( \3051 , \3045 , \3047 );
and \U$2709 ( \3052 , \2637 , \422 );
and \U$2710 ( \3053 , \2463 , \420 );
nor \U$2711 ( \3054 , \3052 , \3053 );
xnor \U$2712 ( \3055 , \3054 , \429 );
and \U$2713 ( \3056 , \2942 , \441 );
and \U$2714 ( \3057 , \2804 , \439 );
nor \U$2715 ( \3058 , \3056 , \3057 );
xnor \U$2716 ( \3059 , \3058 , \448 );
and \U$2717 ( \3060 , \3055 , \3059 );
buf \U$2718 ( \3061 , RIbb2c898_98);
and \U$2719 ( \3062 , \3061 , \436 );
and \U$2720 ( \3063 , \3059 , \3062 );
and \U$2721 ( \3064 , \3055 , \3062 );
or \U$2722 ( \3065 , \3060 , \3063 , \3064 );
and \U$2723 ( \3066 , \1839 , \373 );
and \U$2724 ( \3067 , \1596 , \371 );
nor \U$2725 ( \3068 , \3066 , \3067 );
xnor \U$2726 ( \3069 , \3068 , \380 );
and \U$2727 ( \3070 , \2030 , \391 );
and \U$2728 ( \3071 , \1844 , \389 );
nor \U$2729 ( \3072 , \3070 , \3071 );
xnor \U$2730 ( \3073 , \3072 , \398 );
and \U$2731 ( \3074 , \3069 , \3073 );
and \U$2732 ( \3075 , \2438 , \406 );
and \U$2733 ( \3076 , \2174 , \404 );
nor \U$2734 ( \3077 , \3075 , \3076 );
xnor \U$2735 ( \3078 , \3077 , \413 );
and \U$2736 ( \3079 , \3073 , \3078 );
and \U$2737 ( \3080 , \3069 , \3078 );
or \U$2738 ( \3081 , \3074 , \3079 , \3080 );
and \U$2739 ( \3082 , \3065 , \3081 );
and \U$2740 ( \3083 , \1176 , \793 );
and \U$2741 ( \3084 , \1071 , \791 );
nor \U$2742 ( \3085 , \3083 , \3084 );
xnor \U$2743 ( \3086 , \3085 , \699 );
and \U$2744 ( \3087 , \1297 , \624 );
and \U$2745 ( \3088 , \1181 , \622 );
nor \U$2746 ( \3089 , \3087 , \3088 );
xnor \U$2747 ( \3090 , \3089 , \349 );
and \U$2748 ( \3091 , \3086 , \3090 );
and \U$2749 ( \3092 , \1588 , \357 );
and \U$2750 ( \3093 , \1412 , \355 );
nor \U$2751 ( \3094 , \3092 , \3093 );
xnor \U$2752 ( \3095 , \3094 , \364 );
and \U$2753 ( \3096 , \3090 , \3095 );
and \U$2754 ( \3097 , \3086 , \3095 );
or \U$2755 ( \3098 , \3091 , \3096 , \3097 );
and \U$2756 ( \3099 , \3081 , \3098 );
and \U$2757 ( \3100 , \3065 , \3098 );
or \U$2758 ( \3101 , \3082 , \3099 , \3100 );
and \U$2759 ( \3102 , \408 , \2097 );
and \U$2760 ( \3103 , \385 , \2095 );
nor \U$2761 ( \3104 , \3102 , \3103 );
xnor \U$2762 ( \3105 , \3104 , \1960 );
and \U$2763 ( \3106 , \424 , \1891 );
and \U$2764 ( \3107 , \400 , \1889 );
nor \U$2765 ( \3108 , \3106 , \3107 );
xnor \U$2766 ( \3109 , \3108 , \1739 );
and \U$2767 ( \3110 , \3105 , \3109 );
and \U$2768 ( \3111 , \443 , \1623 );
and \U$2769 ( \3112 , \416 , \1621 );
nor \U$2770 ( \3113 , \3111 , \3112 );
xnor \U$2771 ( \3114 , \3113 , \1467 );
and \U$2772 ( \3115 , \3109 , \3114 );
and \U$2773 ( \3116 , \3105 , \3114 );
or \U$2774 ( \3117 , \3110 , \3115 , \3116 );
xor \U$2775 ( \3118 , \2563 , \2912 );
xor \U$2776 ( \3119 , \2912 , \2913 );
not \U$2777 ( \3120 , \3119 );
and \U$2778 ( \3121 , \3118 , \3120 );
and \U$2779 ( \3122 , \359 , \3121 );
not \U$2780 ( \3123 , \3122 );
xnor \U$2781 ( \3124 , \3123 , \2916 );
and \U$2782 ( \3125 , \375 , \2715 );
and \U$2783 ( \3126 , \351 , \2713 );
nor \U$2784 ( \3127 , \3125 , \3126 );
xnor \U$2785 ( \3128 , \3127 , \2566 );
and \U$2786 ( \3129 , \3124 , \3128 );
and \U$2787 ( \3130 , \393 , \2393 );
and \U$2788 ( \3131 , \367 , \2391 );
nor \U$2789 ( \3132 , \3130 , \3131 );
xnor \U$2790 ( \3133 , \3132 , \2251 );
and \U$2791 ( \3134 , \3128 , \3133 );
and \U$2792 ( \3135 , \3124 , \3133 );
or \U$2793 ( \3136 , \3129 , \3134 , \3135 );
and \U$2794 ( \3137 , \3117 , \3136 );
and \U$2795 ( \3138 , \450 , \1351 );
and \U$2796 ( \3139 , \435 , \1349 );
nor \U$2797 ( \3140 , \3138 , \3139 );
xnor \U$2798 ( \3141 , \3140 , \1238 );
and \U$2799 ( \3142 , \722 , \1157 );
and \U$2800 ( \3143 , \661 , \1155 );
nor \U$2801 ( \3144 , \3142 , \3143 );
xnor \U$2802 ( \3145 , \3144 , \1021 );
and \U$2803 ( \3146 , \3141 , \3145 );
and \U$2804 ( \3147 , \983 , \957 );
and \U$2805 ( \3148 , \785 , \955 );
nor \U$2806 ( \3149 , \3147 , \3148 );
xnor \U$2807 ( \3150 , \3149 , \879 );
and \U$2808 ( \3151 , \3145 , \3150 );
and \U$2809 ( \3152 , \3141 , \3150 );
or \U$2810 ( \3153 , \3146 , \3151 , \3152 );
and \U$2811 ( \3154 , \3136 , \3153 );
and \U$2812 ( \3155 , \3117 , \3153 );
or \U$2813 ( \3156 , \3137 , \3154 , \3155 );
and \U$2814 ( \3157 , \3101 , \3156 );
xor \U$2815 ( \3158 , \2936 , \2940 );
xor \U$2816 ( \3159 , \3158 , \2943 );
xor \U$2817 ( \3160 , \2950 , \2954 );
xor \U$2818 ( \3161 , \3160 , \2959 );
and \U$2819 ( \3162 , \3159 , \3161 );
xor \U$2820 ( \3163 , \2967 , \2971 );
xor \U$2821 ( \3164 , \3163 , \2976 );
and \U$2822 ( \3165 , \3161 , \3164 );
and \U$2823 ( \3166 , \3159 , \3164 );
or \U$2824 ( \3167 , \3162 , \3165 , \3166 );
and \U$2825 ( \3168 , \3156 , \3167 );
and \U$2826 ( \3169 , \3101 , \3167 );
or \U$2827 ( \3170 , \3157 , \3168 , \3169 );
xor \U$2828 ( \3171 , \2882 , \2886 );
xor \U$2829 ( \3172 , \3171 , \2891 );
xor \U$2830 ( \3173 , \2898 , \2902 );
xor \U$2831 ( \3174 , \3173 , \2907 );
and \U$2832 ( \3175 , \3172 , \3174 );
xor \U$2833 ( \3176 , \2917 , \2921 );
xor \U$2834 ( \3177 , \3176 , \2926 );
and \U$2835 ( \3178 , \3174 , \3177 );
and \U$2836 ( \3179 , \3172 , \3177 );
or \U$2837 ( \3180 , \3175 , \3178 , \3179 );
xor \U$2838 ( \3181 , \2997 , \2999 );
xor \U$2839 ( \3182 , \3181 , \3002 );
and \U$2840 ( \3183 , \3180 , \3182 );
xor \U$2841 ( \3184 , \2985 , \2987 );
xor \U$2842 ( \3185 , \3184 , \2989 );
and \U$2843 ( \3186 , \3182 , \3185 );
and \U$2844 ( \3187 , \3180 , \3185 );
or \U$2845 ( \3188 , \3183 , \3186 , \3187 );
and \U$2846 ( \3189 , \3170 , \3188 );
xor \U$2847 ( \3190 , \2894 , \2910 );
xor \U$2848 ( \3191 , \3190 , \2929 );
xor \U$2849 ( \3192 , \2946 , \2962 );
xor \U$2850 ( \3193 , \3192 , \2979 );
and \U$2851 ( \3194 , \3191 , \3193 );
and \U$2852 ( \3195 , \3188 , \3194 );
and \U$2853 ( \3196 , \3170 , \3194 );
or \U$2854 ( \3197 , \3189 , \3195 , \3196 );
xor \U$2855 ( \3198 , \2932 , \2982 );
xor \U$2856 ( \3199 , \3198 , \2992 );
xor \U$2857 ( \3200 , \3005 , \3007 );
xor \U$2858 ( \3201 , \3200 , \3010 );
and \U$2859 ( \3202 , \3199 , \3201 );
xor \U$2860 ( \3203 , \3016 , \3018 );
and \U$2861 ( \3204 , \3201 , \3203 );
and \U$2862 ( \3205 , \3199 , \3203 );
or \U$2863 ( \3206 , \3202 , \3204 , \3205 );
and \U$2864 ( \3207 , \3197 , \3206 );
xor \U$2865 ( \3208 , \3024 , \3026 );
xor \U$2866 ( \3209 , \3208 , \3028 );
and \U$2867 ( \3210 , \3206 , \3209 );
and \U$2868 ( \3211 , \3197 , \3209 );
or \U$2869 ( \3212 , \3207 , \3210 , \3211 );
xor \U$2870 ( \3213 , \2822 , \2840 );
xor \U$2871 ( \3214 , \3213 , \2846 );
and \U$2872 ( \3215 , \3212 , \3214 );
xor \U$2873 ( \3216 , \3022 , \3031 );
xor \U$2874 ( \3217 , \3216 , \3034 );
and \U$2875 ( \3218 , \3214 , \3217 );
and \U$2876 ( \3219 , \3212 , \3217 );
or \U$2877 ( \3220 , \3215 , \3218 , \3219 );
xor \U$2878 ( \3221 , \3037 , \3039 );
xor \U$2879 ( \3222 , \3221 , \3042 );
and \U$2880 ( \3223 , \3220 , \3222 );
and \U$2881 ( \3224 , \3051 , \3223 );
xor \U$2882 ( \3225 , \3051 , \3223 );
xor \U$2883 ( \3226 , \3220 , \3222 );
and \U$2884 ( \3227 , \435 , \1623 );
and \U$2885 ( \3228 , \443 , \1621 );
nor \U$2886 ( \3229 , \3227 , \3228 );
xnor \U$2887 ( \3230 , \3229 , \1467 );
and \U$2888 ( \3231 , \661 , \1351 );
and \U$2889 ( \3232 , \450 , \1349 );
nor \U$2890 ( \3233 , \3231 , \3232 );
xnor \U$2891 ( \3234 , \3233 , \1238 );
and \U$2892 ( \3235 , \3230 , \3234 );
and \U$2893 ( \3236 , \785 , \1157 );
and \U$2894 ( \3237 , \722 , \1155 );
nor \U$2895 ( \3238 , \3236 , \3237 );
xnor \U$2896 ( \3239 , \3238 , \1021 );
and \U$2897 ( \3240 , \3234 , \3239 );
and \U$2898 ( \3241 , \3230 , \3239 );
or \U$2899 ( \3242 , \3235 , \3240 , \3241 );
buf \U$2900 ( \3243 , RIbb2e5a8_36);
buf \U$2901 ( \3244 , RIbb2e530_37);
and \U$2902 ( \3245 , \3243 , \3244 );
not \U$2903 ( \3246 , \3245 );
and \U$2904 ( \3247 , \2913 , \3246 );
not \U$2905 ( \3248 , \3247 );
and \U$2906 ( \3249 , \351 , \3121 );
and \U$2907 ( \3250 , \359 , \3119 );
nor \U$2908 ( \3251 , \3249 , \3250 );
xnor \U$2909 ( \3252 , \3251 , \2916 );
and \U$2910 ( \3253 , \3248 , \3252 );
and \U$2911 ( \3254 , \367 , \2715 );
and \U$2912 ( \3255 , \375 , \2713 );
nor \U$2913 ( \3256 , \3254 , \3255 );
xnor \U$2914 ( \3257 , \3256 , \2566 );
and \U$2915 ( \3258 , \3252 , \3257 );
and \U$2916 ( \3259 , \3248 , \3257 );
or \U$2917 ( \3260 , \3253 , \3258 , \3259 );
and \U$2918 ( \3261 , \3242 , \3260 );
and \U$2919 ( \3262 , \385 , \2393 );
and \U$2920 ( \3263 , \393 , \2391 );
nor \U$2921 ( \3264 , \3262 , \3263 );
xnor \U$2922 ( \3265 , \3264 , \2251 );
and \U$2923 ( \3266 , \400 , \2097 );
and \U$2924 ( \3267 , \408 , \2095 );
nor \U$2925 ( \3268 , \3266 , \3267 );
xnor \U$2926 ( \3269 , \3268 , \1960 );
and \U$2927 ( \3270 , \3265 , \3269 );
and \U$2928 ( \3271 , \416 , \1891 );
and \U$2929 ( \3272 , \424 , \1889 );
nor \U$2930 ( \3273 , \3271 , \3272 );
xnor \U$2931 ( \3274 , \3273 , \1739 );
and \U$2932 ( \3275 , \3269 , \3274 );
and \U$2933 ( \3276 , \3265 , \3274 );
or \U$2934 ( \3277 , \3270 , \3275 , \3276 );
and \U$2935 ( \3278 , \3260 , \3277 );
and \U$2936 ( \3279 , \3242 , \3277 );
or \U$2937 ( \3280 , \3261 , \3278 , \3279 );
and \U$2938 ( \3281 , \2463 , \406 );
and \U$2939 ( \3282 , \2438 , \404 );
nor \U$2940 ( \3283 , \3281 , \3282 );
xnor \U$2941 ( \3284 , \3283 , \413 );
and \U$2942 ( \3285 , \2804 , \422 );
and \U$2943 ( \3286 , \2637 , \420 );
nor \U$2944 ( \3287 , \3285 , \3286 );
xnor \U$2945 ( \3288 , \3287 , \429 );
and \U$2946 ( \3289 , \3284 , \3288 );
and \U$2947 ( \3290 , \3061 , \441 );
and \U$2948 ( \3291 , \2942 , \439 );
nor \U$2949 ( \3292 , \3290 , \3291 );
xnor \U$2950 ( \3293 , \3292 , \448 );
and \U$2951 ( \3294 , \3288 , \3293 );
and \U$2952 ( \3295 , \3284 , \3293 );
or \U$2953 ( \3296 , \3289 , \3294 , \3295 );
and \U$2954 ( \3297 , \1071 , \957 );
and \U$2955 ( \3298 , \983 , \955 );
nor \U$2956 ( \3299 , \3297 , \3298 );
xnor \U$2957 ( \3300 , \3299 , \879 );
and \U$2958 ( \3301 , \1181 , \793 );
and \U$2959 ( \3302 , \1176 , \791 );
nor \U$2960 ( \3303 , \3301 , \3302 );
xnor \U$2961 ( \3304 , \3303 , \699 );
and \U$2962 ( \3305 , \3300 , \3304 );
and \U$2963 ( \3306 , \1412 , \624 );
and \U$2964 ( \3307 , \1297 , \622 );
nor \U$2965 ( \3308 , \3306 , \3307 );
xnor \U$2966 ( \3309 , \3308 , \349 );
and \U$2967 ( \3310 , \3304 , \3309 );
and \U$2968 ( \3311 , \3300 , \3309 );
or \U$2969 ( \3312 , \3305 , \3310 , \3311 );
and \U$2970 ( \3313 , \3296 , \3312 );
and \U$2971 ( \3314 , \1596 , \357 );
and \U$2972 ( \3315 , \1588 , \355 );
nor \U$2973 ( \3316 , \3314 , \3315 );
xnor \U$2974 ( \3317 , \3316 , \364 );
and \U$2975 ( \3318 , \1844 , \373 );
and \U$2976 ( \3319 , \1839 , \371 );
nor \U$2977 ( \3320 , \3318 , \3319 );
xnor \U$2978 ( \3321 , \3320 , \380 );
and \U$2979 ( \3322 , \3317 , \3321 );
and \U$2980 ( \3323 , \2174 , \391 );
and \U$2981 ( \3324 , \2030 , \389 );
nor \U$2982 ( \3325 , \3323 , \3324 );
xnor \U$2983 ( \3326 , \3325 , \398 );
and \U$2984 ( \3327 , \3321 , \3326 );
and \U$2985 ( \3328 , \3317 , \3326 );
or \U$2986 ( \3329 , \3322 , \3327 , \3328 );
and \U$2987 ( \3330 , \3312 , \3329 );
and \U$2988 ( \3331 , \3296 , \3329 );
or \U$2989 ( \3332 , \3313 , \3330 , \3331 );
and \U$2990 ( \3333 , \3280 , \3332 );
xor \U$2991 ( \3334 , \3055 , \3059 );
xor \U$2992 ( \3335 , \3334 , \3062 );
xor \U$2993 ( \3336 , \3069 , \3073 );
xor \U$2994 ( \3337 , \3336 , \3078 );
or \U$2995 ( \3338 , \3335 , \3337 );
and \U$2996 ( \3339 , \3332 , \3338 );
and \U$2997 ( \3340 , \3280 , \3338 );
or \U$2998 ( \3341 , \3333 , \3339 , \3340 );
xor \U$2999 ( \3342 , \3105 , \3109 );
xor \U$3000 ( \3343 , \3342 , \3114 );
xor \U$3001 ( \3344 , \3141 , \3145 );
xor \U$3002 ( \3345 , \3344 , \3150 );
and \U$3003 ( \3346 , \3343 , \3345 );
xor \U$3004 ( \3347 , \3086 , \3090 );
xor \U$3005 ( \3348 , \3347 , \3095 );
and \U$3006 ( \3349 , \3345 , \3348 );
and \U$3007 ( \3350 , \3343 , \3348 );
or \U$3008 ( \3351 , \3346 , \3349 , \3350 );
xor \U$3009 ( \3352 , \3159 , \3161 );
xor \U$3010 ( \3353 , \3352 , \3164 );
and \U$3011 ( \3354 , \3351 , \3353 );
xor \U$3012 ( \3355 , \3172 , \3174 );
xor \U$3013 ( \3356 , \3355 , \3177 );
and \U$3014 ( \3357 , \3353 , \3356 );
and \U$3015 ( \3358 , \3351 , \3356 );
or \U$3016 ( \3359 , \3354 , \3357 , \3358 );
and \U$3017 ( \3360 , \3341 , \3359 );
xor \U$3018 ( \3361 , \3065 , \3081 );
xor \U$3019 ( \3362 , \3361 , \3098 );
xor \U$3020 ( \3363 , \3117 , \3136 );
xor \U$3021 ( \3364 , \3363 , \3153 );
and \U$3022 ( \3365 , \3362 , \3364 );
and \U$3023 ( \3366 , \3359 , \3365 );
and \U$3024 ( \3367 , \3341 , \3365 );
or \U$3025 ( \3368 , \3360 , \3366 , \3367 );
xor \U$3026 ( \3369 , \3101 , \3156 );
xor \U$3027 ( \3370 , \3369 , \3167 );
xor \U$3028 ( \3371 , \3180 , \3182 );
xor \U$3029 ( \3372 , \3371 , \3185 );
and \U$3030 ( \3373 , \3370 , \3372 );
xor \U$3031 ( \3374 , \3191 , \3193 );
and \U$3032 ( \3375 , \3372 , \3374 );
and \U$3033 ( \3376 , \3370 , \3374 );
or \U$3034 ( \3377 , \3373 , \3375 , \3376 );
and \U$3035 ( \3378 , \3368 , \3377 );
xor \U$3036 ( \3379 , \3199 , \3201 );
xor \U$3037 ( \3380 , \3379 , \3203 );
and \U$3038 ( \3381 , \3377 , \3380 );
and \U$3039 ( \3382 , \3368 , \3380 );
or \U$3040 ( \3383 , \3378 , \3381 , \3382 );
xor \U$3041 ( \3384 , \2995 , \3013 );
xor \U$3042 ( \3385 , \3384 , \3019 );
and \U$3043 ( \3386 , \3383 , \3385 );
xor \U$3044 ( \3387 , \3197 , \3206 );
xor \U$3045 ( \3388 , \3387 , \3209 );
and \U$3046 ( \3389 , \3385 , \3388 );
and \U$3047 ( \3390 , \3383 , \3388 );
or \U$3048 ( \3391 , \3386 , \3389 , \3390 );
xor \U$3049 ( \3392 , \3212 , \3214 );
xor \U$3050 ( \3393 , \3392 , \3217 );
and \U$3051 ( \3394 , \3391 , \3393 );
and \U$3052 ( \3395 , \3226 , \3394 );
xor \U$3053 ( \3396 , \3226 , \3394 );
xor \U$3054 ( \3397 , \3391 , \3393 );
and \U$3055 ( \3398 , \450 , \1623 );
and \U$3056 ( \3399 , \435 , \1621 );
nor \U$3057 ( \3400 , \3398 , \3399 );
xnor \U$3058 ( \3401 , \3400 , \1467 );
and \U$3059 ( \3402 , \722 , \1351 );
and \U$3060 ( \3403 , \661 , \1349 );
nor \U$3061 ( \3404 , \3402 , \3403 );
xnor \U$3062 ( \3405 , \3404 , \1238 );
and \U$3063 ( \3406 , \3401 , \3405 );
and \U$3064 ( \3407 , \983 , \1157 );
and \U$3065 ( \3408 , \785 , \1155 );
nor \U$3066 ( \3409 , \3407 , \3408 );
xnor \U$3067 ( \3410 , \3409 , \1021 );
and \U$3068 ( \3411 , \3405 , \3410 );
and \U$3069 ( \3412 , \3401 , \3410 );
or \U$3070 ( \3413 , \3406 , \3411 , \3412 );
and \U$3071 ( \3414 , \408 , \2393 );
and \U$3072 ( \3415 , \385 , \2391 );
nor \U$3073 ( \3416 , \3414 , \3415 );
xnor \U$3074 ( \3417 , \3416 , \2251 );
and \U$3075 ( \3418 , \424 , \2097 );
and \U$3076 ( \3419 , \400 , \2095 );
nor \U$3077 ( \3420 , \3418 , \3419 );
xnor \U$3078 ( \3421 , \3420 , \1960 );
and \U$3079 ( \3422 , \3417 , \3421 );
and \U$3080 ( \3423 , \443 , \1891 );
and \U$3081 ( \3424 , \416 , \1889 );
nor \U$3082 ( \3425 , \3423 , \3424 );
xnor \U$3083 ( \3426 , \3425 , \1739 );
and \U$3084 ( \3427 , \3421 , \3426 );
and \U$3085 ( \3428 , \3417 , \3426 );
or \U$3086 ( \3429 , \3422 , \3427 , \3428 );
and \U$3087 ( \3430 , \3413 , \3429 );
xor \U$3088 ( \3431 , \2913 , \3243 );
xor \U$3089 ( \3432 , \3243 , \3244 );
not \U$3090 ( \3433 , \3432 );
and \U$3091 ( \3434 , \3431 , \3433 );
and \U$3092 ( \3435 , \359 , \3434 );
not \U$3093 ( \3436 , \3435 );
xnor \U$3094 ( \3437 , \3436 , \3247 );
and \U$3095 ( \3438 , \375 , \3121 );
and \U$3096 ( \3439 , \351 , \3119 );
nor \U$3097 ( \3440 , \3438 , \3439 );
xnor \U$3098 ( \3441 , \3440 , \2916 );
and \U$3099 ( \3442 , \3437 , \3441 );
and \U$3100 ( \3443 , \393 , \2715 );
and \U$3101 ( \3444 , \367 , \2713 );
nor \U$3102 ( \3445 , \3443 , \3444 );
xnor \U$3103 ( \3446 , \3445 , \2566 );
and \U$3104 ( \3447 , \3441 , \3446 );
and \U$3105 ( \3448 , \3437 , \3446 );
or \U$3106 ( \3449 , \3442 , \3447 , \3448 );
and \U$3107 ( \3450 , \3429 , \3449 );
and \U$3108 ( \3451 , \3413 , \3449 );
or \U$3109 ( \3452 , \3430 , \3450 , \3451 );
and \U$3110 ( \3453 , \1176 , \957 );
and \U$3111 ( \3454 , \1071 , \955 );
nor \U$3112 ( \3455 , \3453 , \3454 );
xnor \U$3113 ( \3456 , \3455 , \879 );
and \U$3114 ( \3457 , \1297 , \793 );
and \U$3115 ( \3458 , \1181 , \791 );
nor \U$3116 ( \3459 , \3457 , \3458 );
xnor \U$3117 ( \3460 , \3459 , \699 );
and \U$3118 ( \3461 , \3456 , \3460 );
and \U$3119 ( \3462 , \1588 , \624 );
and \U$3120 ( \3463 , \1412 , \622 );
nor \U$3121 ( \3464 , \3462 , \3463 );
xnor \U$3122 ( \3465 , \3464 , \349 );
and \U$3123 ( \3466 , \3460 , \3465 );
and \U$3124 ( \3467 , \3456 , \3465 );
or \U$3125 ( \3468 , \3461 , \3466 , \3467 );
and \U$3126 ( \3469 , \2637 , \406 );
and \U$3127 ( \3470 , \2463 , \404 );
nor \U$3128 ( \3471 , \3469 , \3470 );
xnor \U$3129 ( \3472 , \3471 , \413 );
and \U$3130 ( \3473 , \2942 , \422 );
and \U$3131 ( \3474 , \2804 , \420 );
nor \U$3132 ( \3475 , \3473 , \3474 );
xnor \U$3133 ( \3476 , \3475 , \429 );
and \U$3134 ( \3477 , \3472 , \3476 );
buf \U$3135 ( \3478 , RIbb2c820_99);
and \U$3136 ( \3479 , \3478 , \441 );
and \U$3137 ( \3480 , \3061 , \439 );
nor \U$3138 ( \3481 , \3479 , \3480 );
xnor \U$3139 ( \3482 , \3481 , \448 );
and \U$3140 ( \3483 , \3476 , \3482 );
and \U$3141 ( \3484 , \3472 , \3482 );
or \U$3142 ( \3485 , \3477 , \3483 , \3484 );
and \U$3143 ( \3486 , \3468 , \3485 );
and \U$3144 ( \3487 , \1839 , \357 );
and \U$3145 ( \3488 , \1596 , \355 );
nor \U$3146 ( \3489 , \3487 , \3488 );
xnor \U$3147 ( \3490 , \3489 , \364 );
and \U$3148 ( \3491 , \2030 , \373 );
and \U$3149 ( \3492 , \1844 , \371 );
nor \U$3150 ( \3493 , \3491 , \3492 );
xnor \U$3151 ( \3494 , \3493 , \380 );
and \U$3152 ( \3495 , \3490 , \3494 );
and \U$3153 ( \3496 , \2438 , \391 );
and \U$3154 ( \3497 , \2174 , \389 );
nor \U$3155 ( \3498 , \3496 , \3497 );
xnor \U$3156 ( \3499 , \3498 , \398 );
and \U$3157 ( \3500 , \3494 , \3499 );
and \U$3158 ( \3501 , \3490 , \3499 );
or \U$3159 ( \3502 , \3495 , \3500 , \3501 );
and \U$3160 ( \3503 , \3485 , \3502 );
and \U$3161 ( \3504 , \3468 , \3502 );
or \U$3162 ( \3505 , \3486 , \3503 , \3504 );
and \U$3163 ( \3506 , \3452 , \3505 );
and \U$3164 ( \3507 , \3478 , \436 );
xor \U$3165 ( \3508 , \3284 , \3288 );
xor \U$3166 ( \3509 , \3508 , \3293 );
and \U$3167 ( \3510 , \3507 , \3509 );
xor \U$3168 ( \3511 , \3317 , \3321 );
xor \U$3169 ( \3512 , \3511 , \3326 );
and \U$3170 ( \3513 , \3509 , \3512 );
and \U$3171 ( \3514 , \3507 , \3512 );
or \U$3172 ( \3515 , \3510 , \3513 , \3514 );
and \U$3173 ( \3516 , \3505 , \3515 );
and \U$3174 ( \3517 , \3452 , \3515 );
or \U$3175 ( \3518 , \3506 , \3516 , \3517 );
xor \U$3176 ( \3519 , \3230 , \3234 );
xor \U$3177 ( \3520 , \3519 , \3239 );
xor \U$3178 ( \3521 , \3300 , \3304 );
xor \U$3179 ( \3522 , \3521 , \3309 );
and \U$3180 ( \3523 , \3520 , \3522 );
xor \U$3181 ( \3524 , \3265 , \3269 );
xor \U$3182 ( \3525 , \3524 , \3274 );
and \U$3183 ( \3526 , \3522 , \3525 );
and \U$3184 ( \3527 , \3520 , \3525 );
or \U$3185 ( \3528 , \3523 , \3526 , \3527 );
xor \U$3186 ( \3529 , \3124 , \3128 );
xor \U$3187 ( \3530 , \3529 , \3133 );
and \U$3188 ( \3531 , \3528 , \3530 );
xor \U$3189 ( \3532 , \3343 , \3345 );
xor \U$3190 ( \3533 , \3532 , \3348 );
and \U$3191 ( \3534 , \3530 , \3533 );
and \U$3192 ( \3535 , \3528 , \3533 );
or \U$3193 ( \3536 , \3531 , \3534 , \3535 );
and \U$3194 ( \3537 , \3518 , \3536 );
xor \U$3195 ( \3538 , \3242 , \3260 );
xor \U$3196 ( \3539 , \3538 , \3277 );
xor \U$3197 ( \3540 , \3296 , \3312 );
xor \U$3198 ( \3541 , \3540 , \3329 );
and \U$3199 ( \3542 , \3539 , \3541 );
xnor \U$3200 ( \3543 , \3335 , \3337 );
and \U$3201 ( \3544 , \3541 , \3543 );
and \U$3202 ( \3545 , \3539 , \3543 );
or \U$3203 ( \3546 , \3542 , \3544 , \3545 );
and \U$3204 ( \3547 , \3536 , \3546 );
and \U$3205 ( \3548 , \3518 , \3546 );
or \U$3206 ( \3549 , \3537 , \3547 , \3548 );
xor \U$3207 ( \3550 , \3280 , \3332 );
xor \U$3208 ( \3551 , \3550 , \3338 );
xor \U$3209 ( \3552 , \3351 , \3353 );
xor \U$3210 ( \3553 , \3552 , \3356 );
and \U$3211 ( \3554 , \3551 , \3553 );
xor \U$3212 ( \3555 , \3362 , \3364 );
and \U$3213 ( \3556 , \3553 , \3555 );
and \U$3214 ( \3557 , \3551 , \3555 );
or \U$3215 ( \3558 , \3554 , \3556 , \3557 );
and \U$3216 ( \3559 , \3549 , \3558 );
xor \U$3217 ( \3560 , \3370 , \3372 );
xor \U$3218 ( \3561 , \3560 , \3374 );
and \U$3219 ( \3562 , \3558 , \3561 );
and \U$3220 ( \3563 , \3549 , \3561 );
or \U$3221 ( \3564 , \3559 , \3562 , \3563 );
xor \U$3222 ( \3565 , \3170 , \3188 );
xor \U$3223 ( \3566 , \3565 , \3194 );
and \U$3224 ( \3567 , \3564 , \3566 );
xor \U$3225 ( \3568 , \3368 , \3377 );
xor \U$3226 ( \3569 , \3568 , \3380 );
and \U$3227 ( \3570 , \3566 , \3569 );
and \U$3228 ( \3571 , \3564 , \3569 );
or \U$3229 ( \3572 , \3567 , \3570 , \3571 );
xor \U$3230 ( \3573 , \3383 , \3385 );
xor \U$3231 ( \3574 , \3573 , \3388 );
and \U$3232 ( \3575 , \3572 , \3574 );
and \U$3233 ( \3576 , \3397 , \3575 );
xor \U$3234 ( \3577 , \3397 , \3575 );
xor \U$3235 ( \3578 , \3572 , \3574 );
buf \U$3236 ( \3579 , RIbb2e4b8_38);
buf \U$3237 ( \3580 , RIbb2e440_39);
and \U$3238 ( \3581 , \3579 , \3580 );
not \U$3239 ( \3582 , \3581 );
and \U$3240 ( \3583 , \3244 , \3582 );
not \U$3241 ( \3584 , \3583 );
and \U$3242 ( \3585 , \351 , \3434 );
and \U$3243 ( \3586 , \359 , \3432 );
nor \U$3244 ( \3587 , \3585 , \3586 );
xnor \U$3245 ( \3588 , \3587 , \3247 );
and \U$3246 ( \3589 , \3584 , \3588 );
and \U$3247 ( \3590 , \367 , \3121 );
and \U$3248 ( \3591 , \375 , \3119 );
nor \U$3249 ( \3592 , \3590 , \3591 );
xnor \U$3250 ( \3593 , \3592 , \2916 );
and \U$3251 ( \3594 , \3588 , \3593 );
and \U$3252 ( \3595 , \3584 , \3593 );
or \U$3253 ( \3596 , \3589 , \3594 , \3595 );
and \U$3254 ( \3597 , \385 , \2715 );
and \U$3255 ( \3598 , \393 , \2713 );
nor \U$3256 ( \3599 , \3597 , \3598 );
xnor \U$3257 ( \3600 , \3599 , \2566 );
and \U$3258 ( \3601 , \400 , \2393 );
and \U$3259 ( \3602 , \408 , \2391 );
nor \U$3260 ( \3603 , \3601 , \3602 );
xnor \U$3261 ( \3604 , \3603 , \2251 );
and \U$3262 ( \3605 , \3600 , \3604 );
and \U$3263 ( \3606 , \416 , \2097 );
and \U$3264 ( \3607 , \424 , \2095 );
nor \U$3265 ( \3608 , \3606 , \3607 );
xnor \U$3266 ( \3609 , \3608 , \1960 );
and \U$3267 ( \3610 , \3604 , \3609 );
and \U$3268 ( \3611 , \3600 , \3609 );
or \U$3269 ( \3612 , \3605 , \3610 , \3611 );
and \U$3270 ( \3613 , \3596 , \3612 );
and \U$3271 ( \3614 , \435 , \1891 );
and \U$3272 ( \3615 , \443 , \1889 );
nor \U$3273 ( \3616 , \3614 , \3615 );
xnor \U$3274 ( \3617 , \3616 , \1739 );
and \U$3275 ( \3618 , \661 , \1623 );
and \U$3276 ( \3619 , \450 , \1621 );
nor \U$3277 ( \3620 , \3618 , \3619 );
xnor \U$3278 ( \3621 , \3620 , \1467 );
and \U$3279 ( \3622 , \3617 , \3621 );
and \U$3280 ( \3623 , \785 , \1351 );
and \U$3281 ( \3624 , \722 , \1349 );
nor \U$3282 ( \3625 , \3623 , \3624 );
xnor \U$3283 ( \3626 , \3625 , \1238 );
and \U$3284 ( \3627 , \3621 , \3626 );
and \U$3285 ( \3628 , \3617 , \3626 );
or \U$3286 ( \3629 , \3622 , \3627 , \3628 );
and \U$3287 ( \3630 , \3612 , \3629 );
and \U$3288 ( \3631 , \3596 , \3629 );
or \U$3289 ( \3632 , \3613 , \3630 , \3631 );
and \U$3290 ( \3633 , \1596 , \624 );
and \U$3291 ( \3634 , \1588 , \622 );
nor \U$3292 ( \3635 , \3633 , \3634 );
xnor \U$3293 ( \3636 , \3635 , \349 );
and \U$3294 ( \3637 , \1844 , \357 );
and \U$3295 ( \3638 , \1839 , \355 );
nor \U$3296 ( \3639 , \3637 , \3638 );
xnor \U$3297 ( \3640 , \3639 , \364 );
and \U$3298 ( \3641 , \3636 , \3640 );
and \U$3299 ( \3642 , \2174 , \373 );
and \U$3300 ( \3643 , \2030 , \371 );
nor \U$3301 ( \3644 , \3642 , \3643 );
xnor \U$3302 ( \3645 , \3644 , \380 );
and \U$3303 ( \3646 , \3640 , \3645 );
and \U$3304 ( \3647 , \3636 , \3645 );
or \U$3305 ( \3648 , \3641 , \3646 , \3647 );
and \U$3306 ( \3649 , \1071 , \1157 );
and \U$3307 ( \3650 , \983 , \1155 );
nor \U$3308 ( \3651 , \3649 , \3650 );
xnor \U$3309 ( \3652 , \3651 , \1021 );
and \U$3310 ( \3653 , \1181 , \957 );
and \U$3311 ( \3654 , \1176 , \955 );
nor \U$3312 ( \3655 , \3653 , \3654 );
xnor \U$3313 ( \3656 , \3655 , \879 );
and \U$3314 ( \3657 , \3652 , \3656 );
and \U$3315 ( \3658 , \1412 , \793 );
and \U$3316 ( \3659 , \1297 , \791 );
nor \U$3317 ( \3660 , \3658 , \3659 );
xnor \U$3318 ( \3661 , \3660 , \699 );
and \U$3319 ( \3662 , \3656 , \3661 );
and \U$3320 ( \3663 , \3652 , \3661 );
or \U$3321 ( \3664 , \3657 , \3662 , \3663 );
and \U$3322 ( \3665 , \3648 , \3664 );
and \U$3323 ( \3666 , \2463 , \391 );
and \U$3324 ( \3667 , \2438 , \389 );
nor \U$3325 ( \3668 , \3666 , \3667 );
xnor \U$3326 ( \3669 , \3668 , \398 );
and \U$3327 ( \3670 , \2804 , \406 );
and \U$3328 ( \3671 , \2637 , \404 );
nor \U$3329 ( \3672 , \3670 , \3671 );
xnor \U$3330 ( \3673 , \3672 , \413 );
and \U$3331 ( \3674 , \3669 , \3673 );
and \U$3332 ( \3675 , \3061 , \422 );
and \U$3333 ( \3676 , \2942 , \420 );
nor \U$3334 ( \3677 , \3675 , \3676 );
xnor \U$3335 ( \3678 , \3677 , \429 );
and \U$3336 ( \3679 , \3673 , \3678 );
and \U$3337 ( \3680 , \3669 , \3678 );
or \U$3338 ( \3681 , \3674 , \3679 , \3680 );
and \U$3339 ( \3682 , \3664 , \3681 );
and \U$3340 ( \3683 , \3648 , \3681 );
or \U$3341 ( \3684 , \3665 , \3682 , \3683 );
and \U$3342 ( \3685 , \3632 , \3684 );
buf \U$3343 ( \3686 , RIbb2c7a8_100);
and \U$3344 ( \3687 , \3686 , \436 );
xor \U$3345 ( \3688 , \3472 , \3476 );
xor \U$3346 ( \3689 , \3688 , \3482 );
or \U$3347 ( \3690 , \3687 , \3689 );
and \U$3348 ( \3691 , \3684 , \3690 );
and \U$3349 ( \3692 , \3632 , \3690 );
or \U$3350 ( \3693 , \3685 , \3691 , \3692 );
xor \U$3351 ( \3694 , \3401 , \3405 );
xor \U$3352 ( \3695 , \3694 , \3410 );
xor \U$3353 ( \3696 , \3456 , \3460 );
xor \U$3354 ( \3697 , \3696 , \3465 );
and \U$3355 ( \3698 , \3695 , \3697 );
xor \U$3356 ( \3699 , \3490 , \3494 );
xor \U$3357 ( \3700 , \3699 , \3499 );
and \U$3358 ( \3701 , \3697 , \3700 );
and \U$3359 ( \3702 , \3695 , \3700 );
or \U$3360 ( \3703 , \3698 , \3701 , \3702 );
xor \U$3361 ( \3704 , \3248 , \3252 );
xor \U$3362 ( \3705 , \3704 , \3257 );
and \U$3363 ( \3706 , \3703 , \3705 );
xor \U$3364 ( \3707 , \3520 , \3522 );
xor \U$3365 ( \3708 , \3707 , \3525 );
and \U$3366 ( \3709 , \3705 , \3708 );
and \U$3367 ( \3710 , \3703 , \3708 );
or \U$3368 ( \3711 , \3706 , \3709 , \3710 );
and \U$3369 ( \3712 , \3693 , \3711 );
xor \U$3370 ( \3713 , \3413 , \3429 );
xor \U$3371 ( \3714 , \3713 , \3449 );
xor \U$3372 ( \3715 , \3468 , \3485 );
xor \U$3373 ( \3716 , \3715 , \3502 );
and \U$3374 ( \3717 , \3714 , \3716 );
xor \U$3375 ( \3718 , \3507 , \3509 );
xor \U$3376 ( \3719 , \3718 , \3512 );
and \U$3377 ( \3720 , \3716 , \3719 );
and \U$3378 ( \3721 , \3714 , \3719 );
or \U$3379 ( \3722 , \3717 , \3720 , \3721 );
and \U$3380 ( \3723 , \3711 , \3722 );
and \U$3381 ( \3724 , \3693 , \3722 );
or \U$3382 ( \3725 , \3712 , \3723 , \3724 );
xor \U$3383 ( \3726 , \3452 , \3505 );
xor \U$3384 ( \3727 , \3726 , \3515 );
xor \U$3385 ( \3728 , \3528 , \3530 );
xor \U$3386 ( \3729 , \3728 , \3533 );
and \U$3387 ( \3730 , \3727 , \3729 );
xor \U$3388 ( \3731 , \3539 , \3541 );
xor \U$3389 ( \3732 , \3731 , \3543 );
and \U$3390 ( \3733 , \3729 , \3732 );
and \U$3391 ( \3734 , \3727 , \3732 );
or \U$3392 ( \3735 , \3730 , \3733 , \3734 );
and \U$3393 ( \3736 , \3725 , \3735 );
xor \U$3394 ( \3737 , \3551 , \3553 );
xor \U$3395 ( \3738 , \3737 , \3555 );
and \U$3396 ( \3739 , \3735 , \3738 );
and \U$3397 ( \3740 , \3725 , \3738 );
or \U$3398 ( \3741 , \3736 , \3739 , \3740 );
xor \U$3399 ( \3742 , \3341 , \3359 );
xor \U$3400 ( \3743 , \3742 , \3365 );
and \U$3401 ( \3744 , \3741 , \3743 );
xor \U$3402 ( \3745 , \3549 , \3558 );
xor \U$3403 ( \3746 , \3745 , \3561 );
and \U$3404 ( \3747 , \3743 , \3746 );
and \U$3405 ( \3748 , \3741 , \3746 );
or \U$3406 ( \3749 , \3744 , \3747 , \3748 );
xor \U$3407 ( \3750 , \3564 , \3566 );
xor \U$3408 ( \3751 , \3750 , \3569 );
and \U$3409 ( \3752 , \3749 , \3751 );
and \U$3410 ( \3753 , \3578 , \3752 );
xor \U$3411 ( \3754 , \3578 , \3752 );
xor \U$3412 ( \3755 , \3749 , \3751 );
and \U$3413 ( \3756 , \1176 , \1157 );
and \U$3414 ( \3757 , \1071 , \1155 );
nor \U$3415 ( \3758 , \3756 , \3757 );
xnor \U$3416 ( \3759 , \3758 , \1021 );
and \U$3417 ( \3760 , \1297 , \957 );
and \U$3418 ( \3761 , \1181 , \955 );
nor \U$3419 ( \3762 , \3760 , \3761 );
xnor \U$3420 ( \3763 , \3762 , \879 );
and \U$3421 ( \3764 , \3759 , \3763 );
and \U$3422 ( \3765 , \1588 , \793 );
and \U$3423 ( \3766 , \1412 , \791 );
nor \U$3424 ( \3767 , \3765 , \3766 );
xnor \U$3425 ( \3768 , \3767 , \699 );
and \U$3426 ( \3769 , \3763 , \3768 );
and \U$3427 ( \3770 , \3759 , \3768 );
or \U$3428 ( \3771 , \3764 , \3769 , \3770 );
and \U$3429 ( \3772 , \1839 , \624 );
and \U$3430 ( \3773 , \1596 , \622 );
nor \U$3431 ( \3774 , \3772 , \3773 );
xnor \U$3432 ( \3775 , \3774 , \349 );
and \U$3433 ( \3776 , \2030 , \357 );
and \U$3434 ( \3777 , \1844 , \355 );
nor \U$3435 ( \3778 , \3776 , \3777 );
xnor \U$3436 ( \3779 , \3778 , \364 );
and \U$3437 ( \3780 , \3775 , \3779 );
and \U$3438 ( \3781 , \2438 , \373 );
and \U$3439 ( \3782 , \2174 , \371 );
nor \U$3440 ( \3783 , \3781 , \3782 );
xnor \U$3441 ( \3784 , \3783 , \380 );
and \U$3442 ( \3785 , \3779 , \3784 );
and \U$3443 ( \3786 , \3775 , \3784 );
or \U$3444 ( \3787 , \3780 , \3785 , \3786 );
and \U$3445 ( \3788 , \3771 , \3787 );
and \U$3446 ( \3789 , \2637 , \391 );
and \U$3447 ( \3790 , \2463 , \389 );
nor \U$3448 ( \3791 , \3789 , \3790 );
xnor \U$3449 ( \3792 , \3791 , \398 );
and \U$3450 ( \3793 , \2942 , \406 );
and \U$3451 ( \3794 , \2804 , \404 );
nor \U$3452 ( \3795 , \3793 , \3794 );
xnor \U$3453 ( \3796 , \3795 , \413 );
and \U$3454 ( \3797 , \3792 , \3796 );
and \U$3455 ( \3798 , \3478 , \422 );
and \U$3456 ( \3799 , \3061 , \420 );
nor \U$3457 ( \3800 , \3798 , \3799 );
xnor \U$3458 ( \3801 , \3800 , \429 );
and \U$3459 ( \3802 , \3796 , \3801 );
and \U$3460 ( \3803 , \3792 , \3801 );
or \U$3461 ( \3804 , \3797 , \3802 , \3803 );
and \U$3462 ( \3805 , \3787 , \3804 );
and \U$3463 ( \3806 , \3771 , \3804 );
or \U$3464 ( \3807 , \3788 , \3805 , \3806 );
buf \U$3465 ( \3808 , RIbb2c730_101);
and \U$3466 ( \3809 , \3808 , \441 );
and \U$3467 ( \3810 , \3686 , \439 );
nor \U$3468 ( \3811 , \3809 , \3810 );
xnor \U$3469 ( \3812 , \3811 , \448 );
buf \U$3470 ( \3813 , RIbb2c6b8_102);
and \U$3471 ( \3814 , \3813 , \436 );
or \U$3472 ( \3815 , \3812 , \3814 );
and \U$3473 ( \3816 , \3686 , \441 );
and \U$3474 ( \3817 , \3478 , \439 );
nor \U$3475 ( \3818 , \3816 , \3817 );
xnor \U$3476 ( \3819 , \3818 , \448 );
and \U$3477 ( \3820 , \3815 , \3819 );
and \U$3478 ( \3821 , \3808 , \436 );
and \U$3479 ( \3822 , \3819 , \3821 );
and \U$3480 ( \3823 , \3815 , \3821 );
or \U$3481 ( \3824 , \3820 , \3822 , \3823 );
and \U$3482 ( \3825 , \3807 , \3824 );
xor \U$3483 ( \3826 , \3244 , \3579 );
xor \U$3484 ( \3827 , \3579 , \3580 );
not \U$3485 ( \3828 , \3827 );
and \U$3486 ( \3829 , \3826 , \3828 );
and \U$3487 ( \3830 , \359 , \3829 );
not \U$3488 ( \3831 , \3830 );
xnor \U$3489 ( \3832 , \3831 , \3583 );
and \U$3490 ( \3833 , \375 , \3434 );
and \U$3491 ( \3834 , \351 , \3432 );
nor \U$3492 ( \3835 , \3833 , \3834 );
xnor \U$3493 ( \3836 , \3835 , \3247 );
and \U$3494 ( \3837 , \3832 , \3836 );
and \U$3495 ( \3838 , \393 , \3121 );
and \U$3496 ( \3839 , \367 , \3119 );
nor \U$3497 ( \3840 , \3838 , \3839 );
xnor \U$3498 ( \3841 , \3840 , \2916 );
and \U$3499 ( \3842 , \3836 , \3841 );
and \U$3500 ( \3843 , \3832 , \3841 );
or \U$3501 ( \3844 , \3837 , \3842 , \3843 );
and \U$3502 ( \3845 , \408 , \2715 );
and \U$3503 ( \3846 , \385 , \2713 );
nor \U$3504 ( \3847 , \3845 , \3846 );
xnor \U$3505 ( \3848 , \3847 , \2566 );
and \U$3506 ( \3849 , \424 , \2393 );
and \U$3507 ( \3850 , \400 , \2391 );
nor \U$3508 ( \3851 , \3849 , \3850 );
xnor \U$3509 ( \3852 , \3851 , \2251 );
and \U$3510 ( \3853 , \3848 , \3852 );
and \U$3511 ( \3854 , \443 , \2097 );
and \U$3512 ( \3855 , \416 , \2095 );
nor \U$3513 ( \3856 , \3854 , \3855 );
xnor \U$3514 ( \3857 , \3856 , \1960 );
and \U$3515 ( \3858 , \3852 , \3857 );
and \U$3516 ( \3859 , \3848 , \3857 );
or \U$3517 ( \3860 , \3853 , \3858 , \3859 );
and \U$3518 ( \3861 , \3844 , \3860 );
and \U$3519 ( \3862 , \450 , \1891 );
and \U$3520 ( \3863 , \435 , \1889 );
nor \U$3521 ( \3864 , \3862 , \3863 );
xnor \U$3522 ( \3865 , \3864 , \1739 );
and \U$3523 ( \3866 , \722 , \1623 );
and \U$3524 ( \3867 , \661 , \1621 );
nor \U$3525 ( \3868 , \3866 , \3867 );
xnor \U$3526 ( \3869 , \3868 , \1467 );
and \U$3527 ( \3870 , \3865 , \3869 );
and \U$3528 ( \3871 , \983 , \1351 );
and \U$3529 ( \3872 , \785 , \1349 );
nor \U$3530 ( \3873 , \3871 , \3872 );
xnor \U$3531 ( \3874 , \3873 , \1238 );
and \U$3532 ( \3875 , \3869 , \3874 );
and \U$3533 ( \3876 , \3865 , \3874 );
or \U$3534 ( \3877 , \3870 , \3875 , \3876 );
and \U$3535 ( \3878 , \3860 , \3877 );
and \U$3536 ( \3879 , \3844 , \3877 );
or \U$3537 ( \3880 , \3861 , \3878 , \3879 );
and \U$3538 ( \3881 , \3824 , \3880 );
and \U$3539 ( \3882 , \3807 , \3880 );
or \U$3540 ( \3883 , \3825 , \3881 , \3882 );
xor \U$3541 ( \3884 , \3636 , \3640 );
xor \U$3542 ( \3885 , \3884 , \3645 );
xor \U$3543 ( \3886 , \3652 , \3656 );
xor \U$3544 ( \3887 , \3886 , \3661 );
and \U$3545 ( \3888 , \3885 , \3887 );
xor \U$3546 ( \3889 , \3669 , \3673 );
xor \U$3547 ( \3890 , \3889 , \3678 );
and \U$3548 ( \3891 , \3887 , \3890 );
and \U$3549 ( \3892 , \3885 , \3890 );
or \U$3550 ( \3893 , \3888 , \3891 , \3892 );
xor \U$3551 ( \3894 , \3584 , \3588 );
xor \U$3552 ( \3895 , \3894 , \3593 );
xor \U$3553 ( \3896 , \3600 , \3604 );
xor \U$3554 ( \3897 , \3896 , \3609 );
and \U$3555 ( \3898 , \3895 , \3897 );
xor \U$3556 ( \3899 , \3617 , \3621 );
xor \U$3557 ( \3900 , \3899 , \3626 );
and \U$3558 ( \3901 , \3897 , \3900 );
and \U$3559 ( \3902 , \3895 , \3900 );
or \U$3560 ( \3903 , \3898 , \3901 , \3902 );
and \U$3561 ( \3904 , \3893 , \3903 );
xor \U$3562 ( \3905 , \3417 , \3421 );
xor \U$3563 ( \3906 , \3905 , \3426 );
and \U$3564 ( \3907 , \3903 , \3906 );
and \U$3565 ( \3908 , \3893 , \3906 );
or \U$3566 ( \3909 , \3904 , \3907 , \3908 );
and \U$3567 ( \3910 , \3883 , \3909 );
xor \U$3568 ( \3911 , \3437 , \3441 );
xor \U$3569 ( \3912 , \3911 , \3446 );
xor \U$3570 ( \3913 , \3695 , \3697 );
xor \U$3571 ( \3914 , \3913 , \3700 );
and \U$3572 ( \3915 , \3912 , \3914 );
xnor \U$3573 ( \3916 , \3687 , \3689 );
and \U$3574 ( \3917 , \3914 , \3916 );
and \U$3575 ( \3918 , \3912 , \3916 );
or \U$3576 ( \3919 , \3915 , \3917 , \3918 );
and \U$3577 ( \3920 , \3909 , \3919 );
and \U$3578 ( \3921 , \3883 , \3919 );
or \U$3579 ( \3922 , \3910 , \3920 , \3921 );
xor \U$3580 ( \3923 , \3632 , \3684 );
xor \U$3581 ( \3924 , \3923 , \3690 );
xor \U$3582 ( \3925 , \3703 , \3705 );
xor \U$3583 ( \3926 , \3925 , \3708 );
and \U$3584 ( \3927 , \3924 , \3926 );
xor \U$3585 ( \3928 , \3714 , \3716 );
xor \U$3586 ( \3929 , \3928 , \3719 );
and \U$3587 ( \3930 , \3926 , \3929 );
and \U$3588 ( \3931 , \3924 , \3929 );
or \U$3589 ( \3932 , \3927 , \3930 , \3931 );
and \U$3590 ( \3933 , \3922 , \3932 );
xor \U$3591 ( \3934 , \3727 , \3729 );
xor \U$3592 ( \3935 , \3934 , \3732 );
and \U$3593 ( \3936 , \3932 , \3935 );
and \U$3594 ( \3937 , \3922 , \3935 );
or \U$3595 ( \3938 , \3933 , \3936 , \3937 );
xor \U$3596 ( \3939 , \3518 , \3536 );
xor \U$3597 ( \3940 , \3939 , \3546 );
and \U$3598 ( \3941 , \3938 , \3940 );
xor \U$3599 ( \3942 , \3725 , \3735 );
xor \U$3600 ( \3943 , \3942 , \3738 );
and \U$3601 ( \3944 , \3940 , \3943 );
and \U$3602 ( \3945 , \3938 , \3943 );
or \U$3603 ( \3946 , \3941 , \3944 , \3945 );
xor \U$3604 ( \3947 , \3741 , \3743 );
xor \U$3605 ( \3948 , \3947 , \3746 );
and \U$3606 ( \3949 , \3946 , \3948 );
and \U$3607 ( \3950 , \3755 , \3949 );
xor \U$3608 ( \3951 , \3755 , \3949 );
xor \U$3609 ( \3952 , \3946 , \3948 );
and \U$3610 ( \3953 , \1596 , \793 );
and \U$3611 ( \3954 , \1588 , \791 );
nor \U$3612 ( \3955 , \3953 , \3954 );
xnor \U$3613 ( \3956 , \3955 , \699 );
and \U$3614 ( \3957 , \1844 , \624 );
and \U$3615 ( \3958 , \1839 , \622 );
nor \U$3616 ( \3959 , \3957 , \3958 );
xnor \U$3617 ( \3960 , \3959 , \349 );
and \U$3618 ( \3961 , \3956 , \3960 );
and \U$3619 ( \3962 , \2174 , \357 );
and \U$3620 ( \3963 , \2030 , \355 );
nor \U$3621 ( \3964 , \3962 , \3963 );
xnor \U$3622 ( \3965 , \3964 , \364 );
and \U$3623 ( \3966 , \3960 , \3965 );
and \U$3624 ( \3967 , \3956 , \3965 );
or \U$3625 ( \3968 , \3961 , \3966 , \3967 );
and \U$3626 ( \3969 , \1071 , \1351 );
and \U$3627 ( \3970 , \983 , \1349 );
nor \U$3628 ( \3971 , \3969 , \3970 );
xnor \U$3629 ( \3972 , \3971 , \1238 );
and \U$3630 ( \3973 , \1181 , \1157 );
and \U$3631 ( \3974 , \1176 , \1155 );
nor \U$3632 ( \3975 , \3973 , \3974 );
xnor \U$3633 ( \3976 , \3975 , \1021 );
and \U$3634 ( \3977 , \3972 , \3976 );
and \U$3635 ( \3978 , \1412 , \957 );
and \U$3636 ( \3979 , \1297 , \955 );
nor \U$3637 ( \3980 , \3978 , \3979 );
xnor \U$3638 ( \3981 , \3980 , \879 );
and \U$3639 ( \3982 , \3976 , \3981 );
and \U$3640 ( \3983 , \3972 , \3981 );
or \U$3641 ( \3984 , \3977 , \3982 , \3983 );
and \U$3642 ( \3985 , \3968 , \3984 );
and \U$3643 ( \3986 , \2463 , \373 );
and \U$3644 ( \3987 , \2438 , \371 );
nor \U$3645 ( \3988 , \3986 , \3987 );
xnor \U$3646 ( \3989 , \3988 , \380 );
and \U$3647 ( \3990 , \2804 , \391 );
and \U$3648 ( \3991 , \2637 , \389 );
nor \U$3649 ( \3992 , \3990 , \3991 );
xnor \U$3650 ( \3993 , \3992 , \398 );
and \U$3651 ( \3994 , \3989 , \3993 );
and \U$3652 ( \3995 , \3061 , \406 );
and \U$3653 ( \3996 , \2942 , \404 );
nor \U$3654 ( \3997 , \3995 , \3996 );
xnor \U$3655 ( \3998 , \3997 , \413 );
and \U$3656 ( \3999 , \3993 , \3998 );
and \U$3657 ( \4000 , \3989 , \3998 );
or \U$3658 ( \4001 , \3994 , \3999 , \4000 );
and \U$3659 ( \4002 , \3984 , \4001 );
and \U$3660 ( \4003 , \3968 , \4001 );
or \U$3661 ( \4004 , \3985 , \4002 , \4003 );
buf \U$3662 ( \4005 , RIbb2e3c8_40);
buf \U$3663 ( \4006 , RIbb2e350_41);
and \U$3664 ( \4007 , \4005 , \4006 );
not \U$3665 ( \4008 , \4007 );
and \U$3666 ( \4009 , \3580 , \4008 );
not \U$3667 ( \4010 , \4009 );
and \U$3668 ( \4011 , \351 , \3829 );
and \U$3669 ( \4012 , \359 , \3827 );
nor \U$3670 ( \4013 , \4011 , \4012 );
xnor \U$3671 ( \4014 , \4013 , \3583 );
and \U$3672 ( \4015 , \4010 , \4014 );
and \U$3673 ( \4016 , \367 , \3434 );
and \U$3674 ( \4017 , \375 , \3432 );
nor \U$3675 ( \4018 , \4016 , \4017 );
xnor \U$3676 ( \4019 , \4018 , \3247 );
and \U$3677 ( \4020 , \4014 , \4019 );
and \U$3678 ( \4021 , \4010 , \4019 );
or \U$3679 ( \4022 , \4015 , \4020 , \4021 );
and \U$3680 ( \4023 , \385 , \3121 );
and \U$3681 ( \4024 , \393 , \3119 );
nor \U$3682 ( \4025 , \4023 , \4024 );
xnor \U$3683 ( \4026 , \4025 , \2916 );
and \U$3684 ( \4027 , \400 , \2715 );
and \U$3685 ( \4028 , \408 , \2713 );
nor \U$3686 ( \4029 , \4027 , \4028 );
xnor \U$3687 ( \4030 , \4029 , \2566 );
and \U$3688 ( \4031 , \4026 , \4030 );
and \U$3689 ( \4032 , \416 , \2393 );
and \U$3690 ( \4033 , \424 , \2391 );
nor \U$3691 ( \4034 , \4032 , \4033 );
xnor \U$3692 ( \4035 , \4034 , \2251 );
and \U$3693 ( \4036 , \4030 , \4035 );
and \U$3694 ( \4037 , \4026 , \4035 );
or \U$3695 ( \4038 , \4031 , \4036 , \4037 );
and \U$3696 ( \4039 , \4022 , \4038 );
and \U$3697 ( \4040 , \435 , \2097 );
and \U$3698 ( \4041 , \443 , \2095 );
nor \U$3699 ( \4042 , \4040 , \4041 );
xnor \U$3700 ( \4043 , \4042 , \1960 );
and \U$3701 ( \4044 , \661 , \1891 );
and \U$3702 ( \4045 , \450 , \1889 );
nor \U$3703 ( \4046 , \4044 , \4045 );
xnor \U$3704 ( \4047 , \4046 , \1739 );
and \U$3705 ( \4048 , \4043 , \4047 );
and \U$3706 ( \4049 , \785 , \1623 );
and \U$3707 ( \4050 , \722 , \1621 );
nor \U$3708 ( \4051 , \4049 , \4050 );
xnor \U$3709 ( \4052 , \4051 , \1467 );
and \U$3710 ( \4053 , \4047 , \4052 );
and \U$3711 ( \4054 , \4043 , \4052 );
or \U$3712 ( \4055 , \4048 , \4053 , \4054 );
and \U$3713 ( \4056 , \4038 , \4055 );
and \U$3714 ( \4057 , \4022 , \4055 );
or \U$3715 ( \4058 , \4039 , \4056 , \4057 );
and \U$3716 ( \4059 , \4004 , \4058 );
and \U$3717 ( \4060 , \3686 , \422 );
and \U$3718 ( \4061 , \3478 , \420 );
nor \U$3719 ( \4062 , \4060 , \4061 );
xnor \U$3720 ( \4063 , \4062 , \429 );
and \U$3721 ( \4064 , \3813 , \441 );
and \U$3722 ( \4065 , \3808 , \439 );
nor \U$3723 ( \4066 , \4064 , \4065 );
xnor \U$3724 ( \4067 , \4066 , \448 );
and \U$3725 ( \4068 , \4063 , \4067 );
buf \U$3726 ( \4069 , RIbb2c640_103);
and \U$3727 ( \4070 , \4069 , \436 );
and \U$3728 ( \4071 , \4067 , \4070 );
and \U$3729 ( \4072 , \4063 , \4070 );
or \U$3730 ( \4073 , \4068 , \4071 , \4072 );
xor \U$3731 ( \4074 , \3792 , \3796 );
xor \U$3732 ( \4075 , \4074 , \3801 );
and \U$3733 ( \4076 , \4073 , \4075 );
xnor \U$3734 ( \4077 , \3812 , \3814 );
and \U$3735 ( \4078 , \4075 , \4077 );
and \U$3736 ( \4079 , \4073 , \4077 );
or \U$3737 ( \4080 , \4076 , \4078 , \4079 );
and \U$3738 ( \4081 , \4058 , \4080 );
and \U$3739 ( \4082 , \4004 , \4080 );
or \U$3740 ( \4083 , \4059 , \4081 , \4082 );
xor \U$3741 ( \4084 , \3759 , \3763 );
xor \U$3742 ( \4085 , \4084 , \3768 );
xor \U$3743 ( \4086 , \3775 , \3779 );
xor \U$3744 ( \4087 , \4086 , \3784 );
and \U$3745 ( \4088 , \4085 , \4087 );
xor \U$3746 ( \4089 , \3865 , \3869 );
xor \U$3747 ( \4090 , \4089 , \3874 );
and \U$3748 ( \4091 , \4087 , \4090 );
and \U$3749 ( \4092 , \4085 , \4090 );
or \U$3750 ( \4093 , \4088 , \4091 , \4092 );
xor \U$3751 ( \4094 , \3832 , \3836 );
xor \U$3752 ( \4095 , \4094 , \3841 );
xor \U$3753 ( \4096 , \3848 , \3852 );
xor \U$3754 ( \4097 , \4096 , \3857 );
and \U$3755 ( \4098 , \4095 , \4097 );
and \U$3756 ( \4099 , \4093 , \4098 );
xor \U$3757 ( \4100 , \3895 , \3897 );
xor \U$3758 ( \4101 , \4100 , \3900 );
and \U$3759 ( \4102 , \4098 , \4101 );
and \U$3760 ( \4103 , \4093 , \4101 );
or \U$3761 ( \4104 , \4099 , \4102 , \4103 );
and \U$3762 ( \4105 , \4083 , \4104 );
xor \U$3763 ( \4106 , \3771 , \3787 );
xor \U$3764 ( \4107 , \4106 , \3804 );
xor \U$3765 ( \4108 , \3815 , \3819 );
xor \U$3766 ( \4109 , \4108 , \3821 );
and \U$3767 ( \4110 , \4107 , \4109 );
xor \U$3768 ( \4111 , \3885 , \3887 );
xor \U$3769 ( \4112 , \4111 , \3890 );
and \U$3770 ( \4113 , \4109 , \4112 );
and \U$3771 ( \4114 , \4107 , \4112 );
or \U$3772 ( \4115 , \4110 , \4113 , \4114 );
and \U$3773 ( \4116 , \4104 , \4115 );
and \U$3774 ( \4117 , \4083 , \4115 );
or \U$3775 ( \4118 , \4105 , \4116 , \4117 );
xor \U$3776 ( \4119 , \3596 , \3612 );
xor \U$3777 ( \4120 , \4119 , \3629 );
xor \U$3778 ( \4121 , \3648 , \3664 );
xor \U$3779 ( \4122 , \4121 , \3681 );
and \U$3780 ( \4123 , \4120 , \4122 );
xor \U$3781 ( \4124 , \3912 , \3914 );
xor \U$3782 ( \4125 , \4124 , \3916 );
and \U$3783 ( \4126 , \4122 , \4125 );
and \U$3784 ( \4127 , \4120 , \4125 );
or \U$3785 ( \4128 , \4123 , \4126 , \4127 );
and \U$3786 ( \4129 , \4118 , \4128 );
xor \U$3787 ( \4130 , \3924 , \3926 );
xor \U$3788 ( \4131 , \4130 , \3929 );
and \U$3789 ( \4132 , \4128 , \4131 );
and \U$3790 ( \4133 , \4118 , \4131 );
or \U$3791 ( \4134 , \4129 , \4132 , \4133 );
xor \U$3792 ( \4135 , \3693 , \3711 );
xor \U$3793 ( \4136 , \4135 , \3722 );
and \U$3794 ( \4137 , \4134 , \4136 );
xor \U$3795 ( \4138 , \3922 , \3932 );
xor \U$3796 ( \4139 , \4138 , \3935 );
and \U$3797 ( \4140 , \4136 , \4139 );
and \U$3798 ( \4141 , \4134 , \4139 );
or \U$3799 ( \4142 , \4137 , \4140 , \4141 );
xor \U$3800 ( \4143 , \3938 , \3940 );
xor \U$3801 ( \4144 , \4143 , \3943 );
and \U$3802 ( \4145 , \4142 , \4144 );
and \U$3803 ( \4146 , \3952 , \4145 );
xor \U$3804 ( \4147 , \3952 , \4145 );
xor \U$3805 ( \4148 , \4142 , \4144 );
xor \U$3806 ( \4149 , \3580 , \4005 );
xor \U$3807 ( \4150 , \4005 , \4006 );
not \U$3808 ( \4151 , \4150 );
and \U$3809 ( \4152 , \4149 , \4151 );
and \U$3810 ( \4153 , \359 , \4152 );
not \U$3811 ( \4154 , \4153 );
xnor \U$3812 ( \4155 , \4154 , \4009 );
and \U$3813 ( \4156 , \375 , \3829 );
and \U$3814 ( \4157 , \351 , \3827 );
nor \U$3815 ( \4158 , \4156 , \4157 );
xnor \U$3816 ( \4159 , \4158 , \3583 );
and \U$3817 ( \4160 , \4155 , \4159 );
and \U$3818 ( \4161 , \393 , \3434 );
and \U$3819 ( \4162 , \367 , \3432 );
nor \U$3820 ( \4163 , \4161 , \4162 );
xnor \U$3821 ( \4164 , \4163 , \3247 );
and \U$3822 ( \4165 , \4159 , \4164 );
and \U$3823 ( \4166 , \4155 , \4164 );
or \U$3824 ( \4167 , \4160 , \4165 , \4166 );
and \U$3825 ( \4168 , \408 , \3121 );
and \U$3826 ( \4169 , \385 , \3119 );
nor \U$3827 ( \4170 , \4168 , \4169 );
xnor \U$3828 ( \4171 , \4170 , \2916 );
and \U$3829 ( \4172 , \424 , \2715 );
and \U$3830 ( \4173 , \400 , \2713 );
nor \U$3831 ( \4174 , \4172 , \4173 );
xnor \U$3832 ( \4175 , \4174 , \2566 );
and \U$3833 ( \4176 , \4171 , \4175 );
and \U$3834 ( \4177 , \443 , \2393 );
and \U$3835 ( \4178 , \416 , \2391 );
nor \U$3836 ( \4179 , \4177 , \4178 );
xnor \U$3837 ( \4180 , \4179 , \2251 );
and \U$3838 ( \4181 , \4175 , \4180 );
and \U$3839 ( \4182 , \4171 , \4180 );
or \U$3840 ( \4183 , \4176 , \4181 , \4182 );
and \U$3841 ( \4184 , \4167 , \4183 );
and \U$3842 ( \4185 , \450 , \2097 );
and \U$3843 ( \4186 , \435 , \2095 );
nor \U$3844 ( \4187 , \4185 , \4186 );
xnor \U$3845 ( \4188 , \4187 , \1960 );
and \U$3846 ( \4189 , \722 , \1891 );
and \U$3847 ( \4190 , \661 , \1889 );
nor \U$3848 ( \4191 , \4189 , \4190 );
xnor \U$3849 ( \4192 , \4191 , \1739 );
and \U$3850 ( \4193 , \4188 , \4192 );
and \U$3851 ( \4194 , \983 , \1623 );
and \U$3852 ( \4195 , \785 , \1621 );
nor \U$3853 ( \4196 , \4194 , \4195 );
xnor \U$3854 ( \4197 , \4196 , \1467 );
and \U$3855 ( \4198 , \4192 , \4197 );
and \U$3856 ( \4199 , \4188 , \4197 );
or \U$3857 ( \4200 , \4193 , \4198 , \4199 );
and \U$3858 ( \4201 , \4183 , \4200 );
and \U$3859 ( \4202 , \4167 , \4200 );
or \U$3860 ( \4203 , \4184 , \4201 , \4202 );
and \U$3861 ( \4204 , \2637 , \373 );
and \U$3862 ( \4205 , \2463 , \371 );
nor \U$3863 ( \4206 , \4204 , \4205 );
xnor \U$3864 ( \4207 , \4206 , \380 );
and \U$3865 ( \4208 , \2942 , \391 );
and \U$3866 ( \4209 , \2804 , \389 );
nor \U$3867 ( \4210 , \4208 , \4209 );
xnor \U$3868 ( \4211 , \4210 , \398 );
and \U$3869 ( \4212 , \4207 , \4211 );
and \U$3870 ( \4213 , \3478 , \406 );
and \U$3871 ( \4214 , \3061 , \404 );
nor \U$3872 ( \4215 , \4213 , \4214 );
xnor \U$3873 ( \4216 , \4215 , \413 );
and \U$3874 ( \4217 , \4211 , \4216 );
and \U$3875 ( \4218 , \4207 , \4216 );
or \U$3876 ( \4219 , \4212 , \4217 , \4218 );
and \U$3877 ( \4220 , \1176 , \1351 );
and \U$3878 ( \4221 , \1071 , \1349 );
nor \U$3879 ( \4222 , \4220 , \4221 );
xnor \U$3880 ( \4223 , \4222 , \1238 );
and \U$3881 ( \4224 , \1297 , \1157 );
and \U$3882 ( \4225 , \1181 , \1155 );
nor \U$3883 ( \4226 , \4224 , \4225 );
xnor \U$3884 ( \4227 , \4226 , \1021 );
and \U$3885 ( \4228 , \4223 , \4227 );
and \U$3886 ( \4229 , \1588 , \957 );
and \U$3887 ( \4230 , \1412 , \955 );
nor \U$3888 ( \4231 , \4229 , \4230 );
xnor \U$3889 ( \4232 , \4231 , \879 );
and \U$3890 ( \4233 , \4227 , \4232 );
and \U$3891 ( \4234 , \4223 , \4232 );
or \U$3892 ( \4235 , \4228 , \4233 , \4234 );
and \U$3893 ( \4236 , \4219 , \4235 );
and \U$3894 ( \4237 , \1839 , \793 );
and \U$3895 ( \4238 , \1596 , \791 );
nor \U$3896 ( \4239 , \4237 , \4238 );
xnor \U$3897 ( \4240 , \4239 , \699 );
and \U$3898 ( \4241 , \2030 , \624 );
and \U$3899 ( \4242 , \1844 , \622 );
nor \U$3900 ( \4243 , \4241 , \4242 );
xnor \U$3901 ( \4244 , \4243 , \349 );
and \U$3902 ( \4245 , \4240 , \4244 );
and \U$3903 ( \4246 , \2438 , \357 );
and \U$3904 ( \4247 , \2174 , \355 );
nor \U$3905 ( \4248 , \4246 , \4247 );
xnor \U$3906 ( \4249 , \4248 , \364 );
and \U$3907 ( \4250 , \4244 , \4249 );
and \U$3908 ( \4251 , \4240 , \4249 );
or \U$3909 ( \4252 , \4245 , \4250 , \4251 );
and \U$3910 ( \4253 , \4235 , \4252 );
and \U$3911 ( \4254 , \4219 , \4252 );
or \U$3912 ( \4255 , \4236 , \4253 , \4254 );
and \U$3913 ( \4256 , \4203 , \4255 );
and \U$3914 ( \4257 , \3808 , \422 );
and \U$3915 ( \4258 , \3686 , \420 );
nor \U$3916 ( \4259 , \4257 , \4258 );
xnor \U$3917 ( \4260 , \4259 , \429 );
and \U$3918 ( \4261 , \4069 , \441 );
and \U$3919 ( \4262 , \3813 , \439 );
nor \U$3920 ( \4263 , \4261 , \4262 );
xnor \U$3921 ( \4264 , \4263 , \448 );
and \U$3922 ( \4265 , \4260 , \4264 );
buf \U$3923 ( \4266 , RIbb2c5c8_104);
and \U$3924 ( \4267 , \4266 , \436 );
and \U$3925 ( \4268 , \4264 , \4267 );
and \U$3926 ( \4269 , \4260 , \4267 );
or \U$3927 ( \4270 , \4265 , \4268 , \4269 );
xor \U$3928 ( \4271 , \4063 , \4067 );
xor \U$3929 ( \4272 , \4271 , \4070 );
and \U$3930 ( \4273 , \4270 , \4272 );
xor \U$3931 ( \4274 , \3989 , \3993 );
xor \U$3932 ( \4275 , \4274 , \3998 );
and \U$3933 ( \4276 , \4272 , \4275 );
and \U$3934 ( \4277 , \4270 , \4275 );
or \U$3935 ( \4278 , \4273 , \4276 , \4277 );
and \U$3936 ( \4279 , \4255 , \4278 );
and \U$3937 ( \4280 , \4203 , \4278 );
or \U$3938 ( \4281 , \4256 , \4279 , \4280 );
xor \U$3939 ( \4282 , \3968 , \3984 );
xor \U$3940 ( \4283 , \4282 , \4001 );
xor \U$3941 ( \4284 , \4022 , \4038 );
xor \U$3942 ( \4285 , \4284 , \4055 );
and \U$3943 ( \4286 , \4283 , \4285 );
xor \U$3944 ( \4287 , \4073 , \4075 );
xor \U$3945 ( \4288 , \4287 , \4077 );
and \U$3946 ( \4289 , \4285 , \4288 );
and \U$3947 ( \4290 , \4283 , \4288 );
or \U$3948 ( \4291 , \4286 , \4289 , \4290 );
and \U$3949 ( \4292 , \4281 , \4291 );
xor \U$3950 ( \4293 , \3956 , \3960 );
xor \U$3951 ( \4294 , \4293 , \3965 );
xor \U$3952 ( \4295 , \3972 , \3976 );
xor \U$3953 ( \4296 , \4295 , \3981 );
and \U$3954 ( \4297 , \4294 , \4296 );
xor \U$3955 ( \4298 , \4043 , \4047 );
xor \U$3956 ( \4299 , \4298 , \4052 );
and \U$3957 ( \4300 , \4296 , \4299 );
and \U$3958 ( \4301 , \4294 , \4299 );
or \U$3959 ( \4302 , \4297 , \4300 , \4301 );
xor \U$3960 ( \4303 , \4085 , \4087 );
xor \U$3961 ( \4304 , \4303 , \4090 );
and \U$3962 ( \4305 , \4302 , \4304 );
xor \U$3963 ( \4306 , \4095 , \4097 );
and \U$3964 ( \4307 , \4304 , \4306 );
and \U$3965 ( \4308 , \4302 , \4306 );
or \U$3966 ( \4309 , \4305 , \4307 , \4308 );
and \U$3967 ( \4310 , \4291 , \4309 );
and \U$3968 ( \4311 , \4281 , \4309 );
or \U$3969 ( \4312 , \4292 , \4310 , \4311 );
xor \U$3970 ( \4313 , \3844 , \3860 );
xor \U$3971 ( \4314 , \4313 , \3877 );
xor \U$3972 ( \4315 , \4093 , \4098 );
xor \U$3973 ( \4316 , \4315 , \4101 );
and \U$3974 ( \4317 , \4314 , \4316 );
xor \U$3975 ( \4318 , \4107 , \4109 );
xor \U$3976 ( \4319 , \4318 , \4112 );
and \U$3977 ( \4320 , \4316 , \4319 );
and \U$3978 ( \4321 , \4314 , \4319 );
or \U$3979 ( \4322 , \4317 , \4320 , \4321 );
and \U$3980 ( \4323 , \4312 , \4322 );
xor \U$3981 ( \4324 , \3893 , \3903 );
xor \U$3982 ( \4325 , \4324 , \3906 );
and \U$3983 ( \4326 , \4322 , \4325 );
and \U$3984 ( \4327 , \4312 , \4325 );
or \U$3985 ( \4328 , \4323 , \4326 , \4327 );
xor \U$3986 ( \4329 , \3807 , \3824 );
xor \U$3987 ( \4330 , \4329 , \3880 );
xor \U$3988 ( \4331 , \4083 , \4104 );
xor \U$3989 ( \4332 , \4331 , \4115 );
and \U$3990 ( \4333 , \4330 , \4332 );
xor \U$3991 ( \4334 , \4120 , \4122 );
xor \U$3992 ( \4335 , \4334 , \4125 );
and \U$3993 ( \4336 , \4332 , \4335 );
and \U$3994 ( \4337 , \4330 , \4335 );
or \U$3995 ( \4338 , \4333 , \4336 , \4337 );
and \U$3996 ( \4339 , \4328 , \4338 );
xor \U$3997 ( \4340 , \3883 , \3909 );
xor \U$3998 ( \4341 , \4340 , \3919 );
and \U$3999 ( \4342 , \4338 , \4341 );
and \U$4000 ( \4343 , \4328 , \4341 );
or \U$4001 ( \4344 , \4339 , \4342 , \4343 );
xor \U$4002 ( \4345 , \4134 , \4136 );
xor \U$4003 ( \4346 , \4345 , \4139 );
and \U$4004 ( \4347 , \4344 , \4346 );
and \U$4005 ( \4348 , \4148 , \4347 );
xor \U$4006 ( \4349 , \4148 , \4347 );
xor \U$4007 ( \4350 , \4344 , \4346 );
and \U$4008 ( \4351 , \435 , \2393 );
and \U$4009 ( \4352 , \443 , \2391 );
nor \U$4010 ( \4353 , \4351 , \4352 );
xnor \U$4011 ( \4354 , \4353 , \2251 );
and \U$4012 ( \4355 , \661 , \2097 );
and \U$4013 ( \4356 , \450 , \2095 );
nor \U$4014 ( \4357 , \4355 , \4356 );
xnor \U$4015 ( \4358 , \4357 , \1960 );
and \U$4016 ( \4359 , \4354 , \4358 );
and \U$4017 ( \4360 , \785 , \1891 );
and \U$4018 ( \4361 , \722 , \1889 );
nor \U$4019 ( \4362 , \4360 , \4361 );
xnor \U$4020 ( \4363 , \4362 , \1739 );
and \U$4021 ( \4364 , \4358 , \4363 );
and \U$4022 ( \4365 , \4354 , \4363 );
or \U$4023 ( \4366 , \4359 , \4364 , \4365 );
buf \U$4024 ( \4367 , RIbb2e2d8_42);
buf \U$4025 ( \4368 , RIbb2e260_43);
and \U$4026 ( \4369 , \4367 , \4368 );
not \U$4027 ( \4370 , \4369 );
and \U$4028 ( \4371 , \4006 , \4370 );
not \U$4029 ( \4372 , \4371 );
and \U$4030 ( \4373 , \351 , \4152 );
and \U$4031 ( \4374 , \359 , \4150 );
nor \U$4032 ( \4375 , \4373 , \4374 );
xnor \U$4033 ( \4376 , \4375 , \4009 );
and \U$4034 ( \4377 , \4372 , \4376 );
and \U$4035 ( \4378 , \367 , \3829 );
and \U$4036 ( \4379 , \375 , \3827 );
nor \U$4037 ( \4380 , \4378 , \4379 );
xnor \U$4038 ( \4381 , \4380 , \3583 );
and \U$4039 ( \4382 , \4376 , \4381 );
and \U$4040 ( \4383 , \4372 , \4381 );
or \U$4041 ( \4384 , \4377 , \4382 , \4383 );
and \U$4042 ( \4385 , \4366 , \4384 );
and \U$4043 ( \4386 , \385 , \3434 );
and \U$4044 ( \4387 , \393 , \3432 );
nor \U$4045 ( \4388 , \4386 , \4387 );
xnor \U$4046 ( \4389 , \4388 , \3247 );
and \U$4047 ( \4390 , \400 , \3121 );
and \U$4048 ( \4391 , \408 , \3119 );
nor \U$4049 ( \4392 , \4390 , \4391 );
xnor \U$4050 ( \4393 , \4392 , \2916 );
and \U$4051 ( \4394 , \4389 , \4393 );
and \U$4052 ( \4395 , \416 , \2715 );
and \U$4053 ( \4396 , \424 , \2713 );
nor \U$4054 ( \4397 , \4395 , \4396 );
xnor \U$4055 ( \4398 , \4397 , \2566 );
and \U$4056 ( \4399 , \4393 , \4398 );
and \U$4057 ( \4400 , \4389 , \4398 );
or \U$4058 ( \4401 , \4394 , \4399 , \4400 );
and \U$4059 ( \4402 , \4384 , \4401 );
and \U$4060 ( \4403 , \4366 , \4401 );
or \U$4061 ( \4404 , \4385 , \4402 , \4403 );
and \U$4062 ( \4405 , \2463 , \357 );
and \U$4063 ( \4406 , \2438 , \355 );
nor \U$4064 ( \4407 , \4405 , \4406 );
xnor \U$4065 ( \4408 , \4407 , \364 );
and \U$4066 ( \4409 , \2804 , \373 );
and \U$4067 ( \4410 , \2637 , \371 );
nor \U$4068 ( \4411 , \4409 , \4410 );
xnor \U$4069 ( \4412 , \4411 , \380 );
and \U$4070 ( \4413 , \4408 , \4412 );
and \U$4071 ( \4414 , \3061 , \391 );
and \U$4072 ( \4415 , \2942 , \389 );
nor \U$4073 ( \4416 , \4414 , \4415 );
xnor \U$4074 ( \4417 , \4416 , \398 );
and \U$4075 ( \4418 , \4412 , \4417 );
and \U$4076 ( \4419 , \4408 , \4417 );
or \U$4077 ( \4420 , \4413 , \4418 , \4419 );
and \U$4078 ( \4421 , \1071 , \1623 );
and \U$4079 ( \4422 , \983 , \1621 );
nor \U$4080 ( \4423 , \4421 , \4422 );
xnor \U$4081 ( \4424 , \4423 , \1467 );
and \U$4082 ( \4425 , \1181 , \1351 );
and \U$4083 ( \4426 , \1176 , \1349 );
nor \U$4084 ( \4427 , \4425 , \4426 );
xnor \U$4085 ( \4428 , \4427 , \1238 );
and \U$4086 ( \4429 , \4424 , \4428 );
and \U$4087 ( \4430 , \1412 , \1157 );
and \U$4088 ( \4431 , \1297 , \1155 );
nor \U$4089 ( \4432 , \4430 , \4431 );
xnor \U$4090 ( \4433 , \4432 , \1021 );
and \U$4091 ( \4434 , \4428 , \4433 );
and \U$4092 ( \4435 , \4424 , \4433 );
or \U$4093 ( \4436 , \4429 , \4434 , \4435 );
and \U$4094 ( \4437 , \4420 , \4436 );
and \U$4095 ( \4438 , \1596 , \957 );
and \U$4096 ( \4439 , \1588 , \955 );
nor \U$4097 ( \4440 , \4438 , \4439 );
xnor \U$4098 ( \4441 , \4440 , \879 );
and \U$4099 ( \4442 , \1844 , \793 );
and \U$4100 ( \4443 , \1839 , \791 );
nor \U$4101 ( \4444 , \4442 , \4443 );
xnor \U$4102 ( \4445 , \4444 , \699 );
and \U$4103 ( \4446 , \4441 , \4445 );
and \U$4104 ( \4447 , \2174 , \624 );
and \U$4105 ( \4448 , \2030 , \622 );
nor \U$4106 ( \4449 , \4447 , \4448 );
xnor \U$4107 ( \4450 , \4449 , \349 );
and \U$4108 ( \4451 , \4445 , \4450 );
and \U$4109 ( \4452 , \4441 , \4450 );
or \U$4110 ( \4453 , \4446 , \4451 , \4452 );
and \U$4111 ( \4454 , \4436 , \4453 );
and \U$4112 ( \4455 , \4420 , \4453 );
or \U$4113 ( \4456 , \4437 , \4454 , \4455 );
and \U$4114 ( \4457 , \4404 , \4456 );
and \U$4115 ( \4458 , \3686 , \406 );
and \U$4116 ( \4459 , \3478 , \404 );
nor \U$4117 ( \4460 , \4458 , \4459 );
xnor \U$4118 ( \4461 , \4460 , \413 );
and \U$4119 ( \4462 , \3813 , \422 );
and \U$4120 ( \4463 , \3808 , \420 );
nor \U$4121 ( \4464 , \4462 , \4463 );
xnor \U$4122 ( \4465 , \4464 , \429 );
and \U$4123 ( \4466 , \4461 , \4465 );
and \U$4124 ( \4467 , \4266 , \441 );
and \U$4125 ( \4468 , \4069 , \439 );
nor \U$4126 ( \4469 , \4467 , \4468 );
xnor \U$4127 ( \4470 , \4469 , \448 );
and \U$4128 ( \4471 , \4465 , \4470 );
and \U$4129 ( \4472 , \4461 , \4470 );
or \U$4130 ( \4473 , \4466 , \4471 , \4472 );
xor \U$4131 ( \4474 , \4260 , \4264 );
xor \U$4132 ( \4475 , \4474 , \4267 );
or \U$4133 ( \4476 , \4473 , \4475 );
and \U$4134 ( \4477 , \4456 , \4476 );
and \U$4135 ( \4478 , \4404 , \4476 );
or \U$4136 ( \4479 , \4457 , \4477 , \4478 );
xor \U$4137 ( \4480 , \4207 , \4211 );
xor \U$4138 ( \4481 , \4480 , \4216 );
xor \U$4139 ( \4482 , \4223 , \4227 );
xor \U$4140 ( \4483 , \4482 , \4232 );
and \U$4141 ( \4484 , \4481 , \4483 );
xor \U$4142 ( \4485 , \4240 , \4244 );
xor \U$4143 ( \4486 , \4485 , \4249 );
and \U$4144 ( \4487 , \4483 , \4486 );
and \U$4145 ( \4488 , \4481 , \4486 );
or \U$4146 ( \4489 , \4484 , \4487 , \4488 );
xor \U$4147 ( \4490 , \4155 , \4159 );
xor \U$4148 ( \4491 , \4490 , \4164 );
xor \U$4149 ( \4492 , \4171 , \4175 );
xor \U$4150 ( \4493 , \4492 , \4180 );
and \U$4151 ( \4494 , \4491 , \4493 );
xor \U$4152 ( \4495 , \4188 , \4192 );
xor \U$4153 ( \4496 , \4495 , \4197 );
and \U$4154 ( \4497 , \4493 , \4496 );
and \U$4155 ( \4498 , \4491 , \4496 );
or \U$4156 ( \4499 , \4494 , \4497 , \4498 );
and \U$4157 ( \4500 , \4489 , \4499 );
xor \U$4158 ( \4501 , \4026 , \4030 );
xor \U$4159 ( \4502 , \4501 , \4035 );
and \U$4160 ( \4503 , \4499 , \4502 );
and \U$4161 ( \4504 , \4489 , \4502 );
or \U$4162 ( \4505 , \4500 , \4503 , \4504 );
and \U$4163 ( \4506 , \4479 , \4505 );
xor \U$4164 ( \4507 , \4010 , \4014 );
xor \U$4165 ( \4508 , \4507 , \4019 );
xor \U$4166 ( \4509 , \4294 , \4296 );
xor \U$4167 ( \4510 , \4509 , \4299 );
and \U$4168 ( \4511 , \4508 , \4510 );
xor \U$4169 ( \4512 , \4270 , \4272 );
xor \U$4170 ( \4513 , \4512 , \4275 );
and \U$4171 ( \4514 , \4510 , \4513 );
and \U$4172 ( \4515 , \4508 , \4513 );
or \U$4173 ( \4516 , \4511 , \4514 , \4515 );
and \U$4174 ( \4517 , \4505 , \4516 );
and \U$4175 ( \4518 , \4479 , \4516 );
or \U$4176 ( \4519 , \4506 , \4517 , \4518 );
xor \U$4177 ( \4520 , \4203 , \4255 );
xor \U$4178 ( \4521 , \4520 , \4278 );
xor \U$4179 ( \4522 , \4283 , \4285 );
xor \U$4180 ( \4523 , \4522 , \4288 );
and \U$4181 ( \4524 , \4521 , \4523 );
xor \U$4182 ( \4525 , \4302 , \4304 );
xor \U$4183 ( \4526 , \4525 , \4306 );
and \U$4184 ( \4527 , \4523 , \4526 );
and \U$4185 ( \4528 , \4521 , \4526 );
or \U$4186 ( \4529 , \4524 , \4527 , \4528 );
and \U$4187 ( \4530 , \4519 , \4529 );
xor \U$4188 ( \4531 , \4004 , \4058 );
xor \U$4189 ( \4532 , \4531 , \4080 );
and \U$4190 ( \4533 , \4529 , \4532 );
and \U$4191 ( \4534 , \4519 , \4532 );
or \U$4192 ( \4535 , \4530 , \4533 , \4534 );
xor \U$4193 ( \4536 , \4281 , \4291 );
xor \U$4194 ( \4537 , \4536 , \4309 );
xor \U$4195 ( \4538 , \4314 , \4316 );
xor \U$4196 ( \4539 , \4538 , \4319 );
and \U$4197 ( \4540 , \4537 , \4539 );
and \U$4198 ( \4541 , \4535 , \4540 );
xor \U$4199 ( \4542 , \4330 , \4332 );
xor \U$4200 ( \4543 , \4542 , \4335 );
and \U$4201 ( \4544 , \4540 , \4543 );
and \U$4202 ( \4545 , \4535 , \4543 );
or \U$4203 ( \4546 , \4541 , \4544 , \4545 );
xor \U$4204 ( \4547 , \4328 , \4338 );
xor \U$4205 ( \4548 , \4547 , \4341 );
and \U$4206 ( \4549 , \4546 , \4548 );
xor \U$4207 ( \4550 , \4118 , \4128 );
xor \U$4208 ( \4551 , \4550 , \4131 );
and \U$4209 ( \4552 , \4548 , \4551 );
and \U$4210 ( \4553 , \4546 , \4551 );
or \U$4211 ( \4554 , \4549 , \4552 , \4553 );
and \U$4212 ( \4555 , \4350 , \4554 );
xor \U$4213 ( \4556 , \4350 , \4554 );
xor \U$4214 ( \4557 , \4546 , \4548 );
xor \U$4215 ( \4558 , \4557 , \4551 );
and \U$4216 ( \4559 , \3808 , \406 );
and \U$4217 ( \4560 , \3686 , \404 );
nor \U$4218 ( \4561 , \4559 , \4560 );
xnor \U$4219 ( \4562 , \4561 , \413 );
and \U$4220 ( \4563 , \4069 , \422 );
and \U$4221 ( \4564 , \3813 , \420 );
nor \U$4222 ( \4565 , \4563 , \4564 );
xnor \U$4223 ( \4566 , \4565 , \429 );
and \U$4224 ( \4567 , \4562 , \4566 );
buf \U$4225 ( \4568 , RIbb2c550_105);
and \U$4226 ( \4569 , \4568 , \441 );
and \U$4227 ( \4570 , \4266 , \439 );
nor \U$4228 ( \4571 , \4569 , \4570 );
xnor \U$4229 ( \4572 , \4571 , \448 );
and \U$4230 ( \4573 , \4566 , \4572 );
and \U$4231 ( \4574 , \4562 , \4572 );
or \U$4232 ( \4575 , \4567 , \4573 , \4574 );
buf \U$4233 ( \4576 , RIbb2c4d8_106);
and \U$4234 ( \4577 , \4576 , \436 );
buf \U$4235 ( \4578 , \4577 );
and \U$4236 ( \4579 , \4575 , \4578 );
and \U$4237 ( \4580 , \4568 , \436 );
and \U$4238 ( \4581 , \4578 , \4580 );
and \U$4239 ( \4582 , \4575 , \4580 );
or \U$4240 ( \4583 , \4579 , \4581 , \4582 );
and \U$4241 ( \4584 , \450 , \2393 );
and \U$4242 ( \4585 , \435 , \2391 );
nor \U$4243 ( \4586 , \4584 , \4585 );
xnor \U$4244 ( \4587 , \4586 , \2251 );
and \U$4245 ( \4588 , \722 , \2097 );
and \U$4246 ( \4589 , \661 , \2095 );
nor \U$4247 ( \4590 , \4588 , \4589 );
xnor \U$4248 ( \4591 , \4590 , \1960 );
and \U$4249 ( \4592 , \4587 , \4591 );
and \U$4250 ( \4593 , \983 , \1891 );
and \U$4251 ( \4594 , \785 , \1889 );
nor \U$4252 ( \4595 , \4593 , \4594 );
xnor \U$4253 ( \4596 , \4595 , \1739 );
and \U$4254 ( \4597 , \4591 , \4596 );
and \U$4255 ( \4598 , \4587 , \4596 );
or \U$4256 ( \4599 , \4592 , \4597 , \4598 );
xor \U$4257 ( \4600 , \4006 , \4367 );
xor \U$4258 ( \4601 , \4367 , \4368 );
not \U$4259 ( \4602 , \4601 );
and \U$4260 ( \4603 , \4600 , \4602 );
and \U$4261 ( \4604 , \359 , \4603 );
not \U$4262 ( \4605 , \4604 );
xnor \U$4263 ( \4606 , \4605 , \4371 );
and \U$4264 ( \4607 , \375 , \4152 );
and \U$4265 ( \4608 , \351 , \4150 );
nor \U$4266 ( \4609 , \4607 , \4608 );
xnor \U$4267 ( \4610 , \4609 , \4009 );
and \U$4268 ( \4611 , \4606 , \4610 );
and \U$4269 ( \4612 , \393 , \3829 );
and \U$4270 ( \4613 , \367 , \3827 );
nor \U$4271 ( \4614 , \4612 , \4613 );
xnor \U$4272 ( \4615 , \4614 , \3583 );
and \U$4273 ( \4616 , \4610 , \4615 );
and \U$4274 ( \4617 , \4606 , \4615 );
or \U$4275 ( \4618 , \4611 , \4616 , \4617 );
and \U$4276 ( \4619 , \4599 , \4618 );
and \U$4277 ( \4620 , \408 , \3434 );
and \U$4278 ( \4621 , \385 , \3432 );
nor \U$4279 ( \4622 , \4620 , \4621 );
xnor \U$4280 ( \4623 , \4622 , \3247 );
and \U$4281 ( \4624 , \424 , \3121 );
and \U$4282 ( \4625 , \400 , \3119 );
nor \U$4283 ( \4626 , \4624 , \4625 );
xnor \U$4284 ( \4627 , \4626 , \2916 );
and \U$4285 ( \4628 , \4623 , \4627 );
and \U$4286 ( \4629 , \443 , \2715 );
and \U$4287 ( \4630 , \416 , \2713 );
nor \U$4288 ( \4631 , \4629 , \4630 );
xnor \U$4289 ( \4632 , \4631 , \2566 );
and \U$4290 ( \4633 , \4627 , \4632 );
and \U$4291 ( \4634 , \4623 , \4632 );
or \U$4292 ( \4635 , \4628 , \4633 , \4634 );
and \U$4293 ( \4636 , \4618 , \4635 );
and \U$4294 ( \4637 , \4599 , \4635 );
or \U$4295 ( \4638 , \4619 , \4636 , \4637 );
and \U$4296 ( \4639 , \4583 , \4638 );
and \U$4297 ( \4640 , \2637 , \357 );
and \U$4298 ( \4641 , \2463 , \355 );
nor \U$4299 ( \4642 , \4640 , \4641 );
xnor \U$4300 ( \4643 , \4642 , \364 );
and \U$4301 ( \4644 , \2942 , \373 );
and \U$4302 ( \4645 , \2804 , \371 );
nor \U$4303 ( \4646 , \4644 , \4645 );
xnor \U$4304 ( \4647 , \4646 , \380 );
and \U$4305 ( \4648 , \4643 , \4647 );
and \U$4306 ( \4649 , \3478 , \391 );
and \U$4307 ( \4650 , \3061 , \389 );
nor \U$4308 ( \4651 , \4649 , \4650 );
xnor \U$4309 ( \4652 , \4651 , \398 );
and \U$4310 ( \4653 , \4647 , \4652 );
and \U$4311 ( \4654 , \4643 , \4652 );
or \U$4312 ( \4655 , \4648 , \4653 , \4654 );
and \U$4313 ( \4656 , \1839 , \957 );
and \U$4314 ( \4657 , \1596 , \955 );
nor \U$4315 ( \4658 , \4656 , \4657 );
xnor \U$4316 ( \4659 , \4658 , \879 );
and \U$4317 ( \4660 , \2030 , \793 );
and \U$4318 ( \4661 , \1844 , \791 );
nor \U$4319 ( \4662 , \4660 , \4661 );
xnor \U$4320 ( \4663 , \4662 , \699 );
and \U$4321 ( \4664 , \4659 , \4663 );
and \U$4322 ( \4665 , \2438 , \624 );
and \U$4323 ( \4666 , \2174 , \622 );
nor \U$4324 ( \4667 , \4665 , \4666 );
xnor \U$4325 ( \4668 , \4667 , \349 );
and \U$4326 ( \4669 , \4663 , \4668 );
and \U$4327 ( \4670 , \4659 , \4668 );
or \U$4328 ( \4671 , \4664 , \4669 , \4670 );
and \U$4329 ( \4672 , \4655 , \4671 );
and \U$4330 ( \4673 , \1176 , \1623 );
and \U$4331 ( \4674 , \1071 , \1621 );
nor \U$4332 ( \4675 , \4673 , \4674 );
xnor \U$4333 ( \4676 , \4675 , \1467 );
and \U$4334 ( \4677 , \1297 , \1351 );
and \U$4335 ( \4678 , \1181 , \1349 );
nor \U$4336 ( \4679 , \4677 , \4678 );
xnor \U$4337 ( \4680 , \4679 , \1238 );
and \U$4338 ( \4681 , \4676 , \4680 );
and \U$4339 ( \4682 , \1588 , \1157 );
and \U$4340 ( \4683 , \1412 , \1155 );
nor \U$4341 ( \4684 , \4682 , \4683 );
xnor \U$4342 ( \4685 , \4684 , \1021 );
and \U$4343 ( \4686 , \4680 , \4685 );
and \U$4344 ( \4687 , \4676 , \4685 );
or \U$4345 ( \4688 , \4681 , \4686 , \4687 );
and \U$4346 ( \4689 , \4671 , \4688 );
and \U$4347 ( \4690 , \4655 , \4688 );
or \U$4348 ( \4691 , \4672 , \4689 , \4690 );
and \U$4349 ( \4692 , \4638 , \4691 );
and \U$4350 ( \4693 , \4583 , \4691 );
or \U$4351 ( \4694 , \4639 , \4692 , \4693 );
xor \U$4352 ( \4695 , \4408 , \4412 );
xor \U$4353 ( \4696 , \4695 , \4417 );
xor \U$4354 ( \4697 , \4441 , \4445 );
xor \U$4355 ( \4698 , \4697 , \4450 );
and \U$4356 ( \4699 , \4696 , \4698 );
xor \U$4357 ( \4700 , \4461 , \4465 );
xor \U$4358 ( \4701 , \4700 , \4470 );
and \U$4359 ( \4702 , \4698 , \4701 );
and \U$4360 ( \4703 , \4696 , \4701 );
or \U$4361 ( \4704 , \4699 , \4702 , \4703 );
xor \U$4362 ( \4705 , \4354 , \4358 );
xor \U$4363 ( \4706 , \4705 , \4363 );
xor \U$4364 ( \4707 , \4424 , \4428 );
xor \U$4365 ( \4708 , \4707 , \4433 );
and \U$4366 ( \4709 , \4706 , \4708 );
xor \U$4367 ( \4710 , \4389 , \4393 );
xor \U$4368 ( \4711 , \4710 , \4398 );
and \U$4369 ( \4712 , \4708 , \4711 );
and \U$4370 ( \4713 , \4706 , \4711 );
or \U$4371 ( \4714 , \4709 , \4712 , \4713 );
and \U$4372 ( \4715 , \4704 , \4714 );
xor \U$4373 ( \4716 , \4491 , \4493 );
xor \U$4374 ( \4717 , \4716 , \4496 );
and \U$4375 ( \4718 , \4714 , \4717 );
and \U$4376 ( \4719 , \4704 , \4717 );
or \U$4377 ( \4720 , \4715 , \4718 , \4719 );
and \U$4378 ( \4721 , \4694 , \4720 );
xor \U$4379 ( \4722 , \4420 , \4436 );
xor \U$4380 ( \4723 , \4722 , \4453 );
xor \U$4381 ( \4724 , \4481 , \4483 );
xor \U$4382 ( \4725 , \4724 , \4486 );
and \U$4383 ( \4726 , \4723 , \4725 );
xnor \U$4384 ( \4727 , \4473 , \4475 );
and \U$4385 ( \4728 , \4725 , \4727 );
and \U$4386 ( \4729 , \4723 , \4727 );
or \U$4387 ( \4730 , \4726 , \4728 , \4729 );
and \U$4388 ( \4731 , \4720 , \4730 );
and \U$4389 ( \4732 , \4694 , \4730 );
or \U$4390 ( \4733 , \4721 , \4731 , \4732 );
xor \U$4391 ( \4734 , \4167 , \4183 );
xor \U$4392 ( \4735 , \4734 , \4200 );
xor \U$4393 ( \4736 , \4219 , \4235 );
xor \U$4394 ( \4737 , \4736 , \4252 );
and \U$4395 ( \4738 , \4735 , \4737 );
xor \U$4396 ( \4739 , \4508 , \4510 );
xor \U$4397 ( \4740 , \4739 , \4513 );
and \U$4398 ( \4741 , \4737 , \4740 );
and \U$4399 ( \4742 , \4735 , \4740 );
or \U$4400 ( \4743 , \4738 , \4741 , \4742 );
and \U$4401 ( \4744 , \4733 , \4743 );
xor \U$4402 ( \4745 , \4521 , \4523 );
xor \U$4403 ( \4746 , \4745 , \4526 );
and \U$4404 ( \4747 , \4743 , \4746 );
and \U$4405 ( \4748 , \4733 , \4746 );
or \U$4406 ( \4749 , \4744 , \4747 , \4748 );
xor \U$4407 ( \4750 , \4519 , \4529 );
xor \U$4408 ( \4751 , \4750 , \4532 );
and \U$4409 ( \4752 , \4749 , \4751 );
xor \U$4410 ( \4753 , \4537 , \4539 );
and \U$4411 ( \4754 , \4751 , \4753 );
and \U$4412 ( \4755 , \4749 , \4753 );
or \U$4413 ( \4756 , \4752 , \4754 , \4755 );
xor \U$4414 ( \4757 , \4312 , \4322 );
xor \U$4415 ( \4758 , \4757 , \4325 );
and \U$4416 ( \4759 , \4756 , \4758 );
xor \U$4417 ( \4760 , \4535 , \4540 );
xor \U$4418 ( \4761 , \4760 , \4543 );
and \U$4419 ( \4762 , \4758 , \4761 );
and \U$4420 ( \4763 , \4756 , \4761 );
or \U$4421 ( \4764 , \4759 , \4762 , \4763 );
and \U$4422 ( \4765 , \4558 , \4764 );
xor \U$4423 ( \4766 , \4558 , \4764 );
xor \U$4424 ( \4767 , \4756 , \4758 );
xor \U$4425 ( \4768 , \4767 , \4761 );
and \U$4426 ( \4769 , \435 , \2715 );
and \U$4427 ( \4770 , \443 , \2713 );
nor \U$4428 ( \4771 , \4769 , \4770 );
xnor \U$4429 ( \4772 , \4771 , \2566 );
and \U$4430 ( \4773 , \661 , \2393 );
and \U$4431 ( \4774 , \450 , \2391 );
nor \U$4432 ( \4775 , \4773 , \4774 );
xnor \U$4433 ( \4776 , \4775 , \2251 );
and \U$4434 ( \4777 , \4772 , \4776 );
and \U$4435 ( \4778 , \785 , \2097 );
and \U$4436 ( \4779 , \722 , \2095 );
nor \U$4437 ( \4780 , \4778 , \4779 );
xnor \U$4438 ( \4781 , \4780 , \1960 );
and \U$4439 ( \4782 , \4776 , \4781 );
and \U$4440 ( \4783 , \4772 , \4781 );
or \U$4441 ( \4784 , \4777 , \4782 , \4783 );
buf \U$4442 ( \4785 , RIbb2e1e8_44);
buf \U$4443 ( \4786 , RIbb2e170_45);
and \U$4444 ( \4787 , \4785 , \4786 );
not \U$4445 ( \4788 , \4787 );
and \U$4446 ( \4789 , \4368 , \4788 );
not \U$4447 ( \4790 , \4789 );
and \U$4448 ( \4791 , \351 , \4603 );
and \U$4449 ( \4792 , \359 , \4601 );
nor \U$4450 ( \4793 , \4791 , \4792 );
xnor \U$4451 ( \4794 , \4793 , \4371 );
and \U$4452 ( \4795 , \4790 , \4794 );
and \U$4453 ( \4796 , \367 , \4152 );
and \U$4454 ( \4797 , \375 , \4150 );
nor \U$4455 ( \4798 , \4796 , \4797 );
xnor \U$4456 ( \4799 , \4798 , \4009 );
and \U$4457 ( \4800 , \4794 , \4799 );
and \U$4458 ( \4801 , \4790 , \4799 );
or \U$4459 ( \4802 , \4795 , \4800 , \4801 );
and \U$4460 ( \4803 , \4784 , \4802 );
and \U$4461 ( \4804 , \385 , \3829 );
and \U$4462 ( \4805 , \393 , \3827 );
nor \U$4463 ( \4806 , \4804 , \4805 );
xnor \U$4464 ( \4807 , \4806 , \3583 );
and \U$4465 ( \4808 , \400 , \3434 );
and \U$4466 ( \4809 , \408 , \3432 );
nor \U$4467 ( \4810 , \4808 , \4809 );
xnor \U$4468 ( \4811 , \4810 , \3247 );
and \U$4469 ( \4812 , \4807 , \4811 );
and \U$4470 ( \4813 , \416 , \3121 );
and \U$4471 ( \4814 , \424 , \3119 );
nor \U$4472 ( \4815 , \4813 , \4814 );
xnor \U$4473 ( \4816 , \4815 , \2916 );
and \U$4474 ( \4817 , \4811 , \4816 );
and \U$4475 ( \4818 , \4807 , \4816 );
or \U$4476 ( \4819 , \4812 , \4817 , \4818 );
and \U$4477 ( \4820 , \4802 , \4819 );
and \U$4478 ( \4821 , \4784 , \4819 );
or \U$4479 ( \4822 , \4803 , \4820 , \4821 );
and \U$4480 ( \4823 , \1071 , \1891 );
and \U$4481 ( \4824 , \983 , \1889 );
nor \U$4482 ( \4825 , \4823 , \4824 );
xnor \U$4483 ( \4826 , \4825 , \1739 );
and \U$4484 ( \4827 , \1181 , \1623 );
and \U$4485 ( \4828 , \1176 , \1621 );
nor \U$4486 ( \4829 , \4827 , \4828 );
xnor \U$4487 ( \4830 , \4829 , \1467 );
and \U$4488 ( \4831 , \4826 , \4830 );
and \U$4489 ( \4832 , \1412 , \1351 );
and \U$4490 ( \4833 , \1297 , \1349 );
nor \U$4491 ( \4834 , \4832 , \4833 );
xnor \U$4492 ( \4835 , \4834 , \1238 );
and \U$4493 ( \4836 , \4830 , \4835 );
and \U$4494 ( \4837 , \4826 , \4835 );
or \U$4495 ( \4838 , \4831 , \4836 , \4837 );
and \U$4496 ( \4839 , \2463 , \624 );
and \U$4497 ( \4840 , \2438 , \622 );
nor \U$4498 ( \4841 , \4839 , \4840 );
xnor \U$4499 ( \4842 , \4841 , \349 );
and \U$4500 ( \4843 , \2804 , \357 );
and \U$4501 ( \4844 , \2637 , \355 );
nor \U$4502 ( \4845 , \4843 , \4844 );
xnor \U$4503 ( \4846 , \4845 , \364 );
and \U$4504 ( \4847 , \4842 , \4846 );
and \U$4505 ( \4848 , \3061 , \373 );
and \U$4506 ( \4849 , \2942 , \371 );
nor \U$4507 ( \4850 , \4848 , \4849 );
xnor \U$4508 ( \4851 , \4850 , \380 );
and \U$4509 ( \4852 , \4846 , \4851 );
and \U$4510 ( \4853 , \4842 , \4851 );
or \U$4511 ( \4854 , \4847 , \4852 , \4853 );
and \U$4512 ( \4855 , \4838 , \4854 );
and \U$4513 ( \4856 , \1596 , \1157 );
and \U$4514 ( \4857 , \1588 , \1155 );
nor \U$4515 ( \4858 , \4856 , \4857 );
xnor \U$4516 ( \4859 , \4858 , \1021 );
and \U$4517 ( \4860 , \1844 , \957 );
and \U$4518 ( \4861 , \1839 , \955 );
nor \U$4519 ( \4862 , \4860 , \4861 );
xnor \U$4520 ( \4863 , \4862 , \879 );
and \U$4521 ( \4864 , \4859 , \4863 );
and \U$4522 ( \4865 , \2174 , \793 );
and \U$4523 ( \4866 , \2030 , \791 );
nor \U$4524 ( \4867 , \4865 , \4866 );
xnor \U$4525 ( \4868 , \4867 , \699 );
and \U$4526 ( \4869 , \4863 , \4868 );
and \U$4527 ( \4870 , \4859 , \4868 );
or \U$4528 ( \4871 , \4864 , \4869 , \4870 );
and \U$4529 ( \4872 , \4854 , \4871 );
and \U$4530 ( \4873 , \4838 , \4871 );
or \U$4531 ( \4874 , \4855 , \4872 , \4873 );
and \U$4532 ( \4875 , \4822 , \4874 );
and \U$4533 ( \4876 , \3686 , \391 );
and \U$4534 ( \4877 , \3478 , \389 );
nor \U$4535 ( \4878 , \4876 , \4877 );
xnor \U$4536 ( \4879 , \4878 , \398 );
and \U$4537 ( \4880 , \3813 , \406 );
and \U$4538 ( \4881 , \3808 , \404 );
nor \U$4539 ( \4882 , \4880 , \4881 );
xnor \U$4540 ( \4883 , \4882 , \413 );
and \U$4541 ( \4884 , \4879 , \4883 );
and \U$4542 ( \4885 , \4266 , \422 );
and \U$4543 ( \4886 , \4069 , \420 );
nor \U$4544 ( \4887 , \4885 , \4886 );
xnor \U$4545 ( \4888 , \4887 , \429 );
and \U$4546 ( \4889 , \4883 , \4888 );
and \U$4547 ( \4890 , \4879 , \4888 );
or \U$4548 ( \4891 , \4884 , \4889 , \4890 );
xor \U$4549 ( \4892 , \4562 , \4566 );
xor \U$4550 ( \4893 , \4892 , \4572 );
and \U$4551 ( \4894 , \4891 , \4893 );
not \U$4552 ( \4895 , \4577 );
and \U$4553 ( \4896 , \4893 , \4895 );
and \U$4554 ( \4897 , \4891 , \4895 );
or \U$4555 ( \4898 , \4894 , \4896 , \4897 );
and \U$4556 ( \4899 , \4874 , \4898 );
and \U$4557 ( \4900 , \4822 , \4898 );
or \U$4558 ( \4901 , \4875 , \4899 , \4900 );
xor \U$4559 ( \4902 , \4643 , \4647 );
xor \U$4560 ( \4903 , \4902 , \4652 );
xor \U$4561 ( \4904 , \4659 , \4663 );
xor \U$4562 ( \4905 , \4904 , \4668 );
and \U$4563 ( \4906 , \4903 , \4905 );
xor \U$4564 ( \4907 , \4676 , \4680 );
xor \U$4565 ( \4908 , \4907 , \4685 );
and \U$4566 ( \4909 , \4905 , \4908 );
and \U$4567 ( \4910 , \4903 , \4908 );
or \U$4568 ( \4911 , \4906 , \4909 , \4910 );
xor \U$4569 ( \4912 , \4587 , \4591 );
xor \U$4570 ( \4913 , \4912 , \4596 );
xor \U$4571 ( \4914 , \4606 , \4610 );
xor \U$4572 ( \4915 , \4914 , \4615 );
and \U$4573 ( \4916 , \4913 , \4915 );
xor \U$4574 ( \4917 , \4623 , \4627 );
xor \U$4575 ( \4918 , \4917 , \4632 );
and \U$4576 ( \4919 , \4915 , \4918 );
and \U$4577 ( \4920 , \4913 , \4918 );
or \U$4578 ( \4921 , \4916 , \4919 , \4920 );
and \U$4579 ( \4922 , \4911 , \4921 );
xor \U$4580 ( \4923 , \4372 , \4376 );
xor \U$4581 ( \4924 , \4923 , \4381 );
and \U$4582 ( \4925 , \4921 , \4924 );
and \U$4583 ( \4926 , \4911 , \4924 );
or \U$4584 ( \4927 , \4922 , \4925 , \4926 );
and \U$4585 ( \4928 , \4901 , \4927 );
xor \U$4586 ( \4929 , \4575 , \4578 );
xor \U$4587 ( \4930 , \4929 , \4580 );
xor \U$4588 ( \4931 , \4696 , \4698 );
xor \U$4589 ( \4932 , \4931 , \4701 );
and \U$4590 ( \4933 , \4930 , \4932 );
xor \U$4591 ( \4934 , \4706 , \4708 );
xor \U$4592 ( \4935 , \4934 , \4711 );
and \U$4593 ( \4936 , \4932 , \4935 );
and \U$4594 ( \4937 , \4930 , \4935 );
or \U$4595 ( \4938 , \4933 , \4936 , \4937 );
and \U$4596 ( \4939 , \4927 , \4938 );
and \U$4597 ( \4940 , \4901 , \4938 );
or \U$4598 ( \4941 , \4928 , \4939 , \4940 );
xor \U$4599 ( \4942 , \4366 , \4384 );
xor \U$4600 ( \4943 , \4942 , \4401 );
xor \U$4601 ( \4944 , \4704 , \4714 );
xor \U$4602 ( \4945 , \4944 , \4717 );
and \U$4603 ( \4946 , \4943 , \4945 );
xor \U$4604 ( \4947 , \4723 , \4725 );
xor \U$4605 ( \4948 , \4947 , \4727 );
and \U$4606 ( \4949 , \4945 , \4948 );
and \U$4607 ( \4950 , \4943 , \4948 );
or \U$4608 ( \4951 , \4946 , \4949 , \4950 );
and \U$4609 ( \4952 , \4941 , \4951 );
xor \U$4610 ( \4953 , \4489 , \4499 );
xor \U$4611 ( \4954 , \4953 , \4502 );
and \U$4612 ( \4955 , \4951 , \4954 );
and \U$4613 ( \4956 , \4941 , \4954 );
or \U$4614 ( \4957 , \4952 , \4955 , \4956 );
xor \U$4615 ( \4958 , \4404 , \4456 );
xor \U$4616 ( \4959 , \4958 , \4476 );
xor \U$4617 ( \4960 , \4694 , \4720 );
xor \U$4618 ( \4961 , \4960 , \4730 );
and \U$4619 ( \4962 , \4959 , \4961 );
xor \U$4620 ( \4963 , \4735 , \4737 );
xor \U$4621 ( \4964 , \4963 , \4740 );
and \U$4622 ( \4965 , \4961 , \4964 );
and \U$4623 ( \4966 , \4959 , \4964 );
or \U$4624 ( \4967 , \4962 , \4965 , \4966 );
and \U$4625 ( \4968 , \4957 , \4967 );
xor \U$4626 ( \4969 , \4479 , \4505 );
xor \U$4627 ( \4970 , \4969 , \4516 );
and \U$4628 ( \4971 , \4967 , \4970 );
and \U$4629 ( \4972 , \4957 , \4970 );
or \U$4630 ( \4973 , \4968 , \4971 , \4972 );
xor \U$4631 ( \4974 , \4368 , \4785 );
xor \U$4632 ( \4975 , \4785 , \4786 );
not \U$4633 ( \4976 , \4975 );
and \U$4634 ( \4977 , \4974 , \4976 );
and \U$4635 ( \4978 , \359 , \4977 );
not \U$4636 ( \4979 , \4978 );
xnor \U$4637 ( \4980 , \4979 , \4789 );
and \U$4638 ( \4981 , \375 , \4603 );
and \U$4639 ( \4982 , \351 , \4601 );
nor \U$4640 ( \4983 , \4981 , \4982 );
xnor \U$4641 ( \4984 , \4983 , \4371 );
and \U$4642 ( \4985 , \4980 , \4984 );
and \U$4643 ( \4986 , \393 , \4152 );
and \U$4644 ( \4987 , \367 , \4150 );
nor \U$4645 ( \4988 , \4986 , \4987 );
xnor \U$4646 ( \4989 , \4988 , \4009 );
and \U$4647 ( \4990 , \4984 , \4989 );
and \U$4648 ( \4991 , \4980 , \4989 );
or \U$4649 ( \4992 , \4985 , \4990 , \4991 );
and \U$4650 ( \4993 , \450 , \2715 );
and \U$4651 ( \4994 , \435 , \2713 );
nor \U$4652 ( \4995 , \4993 , \4994 );
xnor \U$4653 ( \4996 , \4995 , \2566 );
and \U$4654 ( \4997 , \722 , \2393 );
and \U$4655 ( \4998 , \661 , \2391 );
nor \U$4656 ( \4999 , \4997 , \4998 );
xnor \U$4657 ( \5000 , \4999 , \2251 );
and \U$4658 ( \5001 , \4996 , \5000 );
and \U$4659 ( \5002 , \983 , \2097 );
and \U$4660 ( \5003 , \785 , \2095 );
nor \U$4661 ( \5004 , \5002 , \5003 );
xnor \U$4662 ( \5005 , \5004 , \1960 );
and \U$4663 ( \5006 , \5000 , \5005 );
and \U$4664 ( \5007 , \4996 , \5005 );
or \U$4665 ( \5008 , \5001 , \5006 , \5007 );
and \U$4666 ( \5009 , \4992 , \5008 );
and \U$4667 ( \5010 , \408 , \3829 );
and \U$4668 ( \5011 , \385 , \3827 );
nor \U$4669 ( \5012 , \5010 , \5011 );
xnor \U$4670 ( \5013 , \5012 , \3583 );
and \U$4671 ( \5014 , \424 , \3434 );
and \U$4672 ( \5015 , \400 , \3432 );
nor \U$4673 ( \5016 , \5014 , \5015 );
xnor \U$4674 ( \5017 , \5016 , \3247 );
and \U$4675 ( \5018 , \5013 , \5017 );
and \U$4676 ( \5019 , \443 , \3121 );
and \U$4677 ( \5020 , \416 , \3119 );
nor \U$4678 ( \5021 , \5019 , \5020 );
xnor \U$4679 ( \5022 , \5021 , \2916 );
and \U$4680 ( \5023 , \5017 , \5022 );
and \U$4681 ( \5024 , \5013 , \5022 );
or \U$4682 ( \5025 , \5018 , \5023 , \5024 );
and \U$4683 ( \5026 , \5008 , \5025 );
and \U$4684 ( \5027 , \4992 , \5025 );
or \U$4685 ( \5028 , \5009 , \5026 , \5027 );
and \U$4686 ( \5029 , \3808 , \391 );
and \U$4687 ( \5030 , \3686 , \389 );
nor \U$4688 ( \5031 , \5029 , \5030 );
xnor \U$4689 ( \5032 , \5031 , \398 );
and \U$4690 ( \5033 , \4069 , \406 );
and \U$4691 ( \5034 , \3813 , \404 );
nor \U$4692 ( \5035 , \5033 , \5034 );
xnor \U$4693 ( \5036 , \5035 , \413 );
and \U$4694 ( \5037 , \5032 , \5036 );
and \U$4695 ( \5038 , \4568 , \422 );
and \U$4696 ( \5039 , \4266 , \420 );
nor \U$4697 ( \5040 , \5038 , \5039 );
xnor \U$4698 ( \5041 , \5040 , \429 );
and \U$4699 ( \5042 , \5036 , \5041 );
and \U$4700 ( \5043 , \5032 , \5041 );
or \U$4701 ( \5044 , \5037 , \5042 , \5043 );
buf \U$4702 ( \5045 , RIbb2c460_107);
and \U$4703 ( \5046 , \5045 , \441 );
and \U$4704 ( \5047 , \4576 , \439 );
nor \U$4705 ( \5048 , \5046 , \5047 );
xnor \U$4706 ( \5049 , \5048 , \448 );
buf \U$4707 ( \5050 , RIbb2c3e8_108);
and \U$4708 ( \5051 , \5050 , \436 );
or \U$4709 ( \5052 , \5049 , \5051 );
and \U$4710 ( \5053 , \5044 , \5052 );
and \U$4711 ( \5054 , \4576 , \441 );
and \U$4712 ( \5055 , \4568 , \439 );
nor \U$4713 ( \5056 , \5054 , \5055 );
xnor \U$4714 ( \5057 , \5056 , \448 );
and \U$4715 ( \5058 , \5052 , \5057 );
and \U$4716 ( \5059 , \5044 , \5057 );
or \U$4717 ( \5060 , \5053 , \5058 , \5059 );
and \U$4718 ( \5061 , \5028 , \5060 );
and \U$4719 ( \5062 , \1176 , \1891 );
and \U$4720 ( \5063 , \1071 , \1889 );
nor \U$4721 ( \5064 , \5062 , \5063 );
xnor \U$4722 ( \5065 , \5064 , \1739 );
and \U$4723 ( \5066 , \1297 , \1623 );
and \U$4724 ( \5067 , \1181 , \1621 );
nor \U$4725 ( \5068 , \5066 , \5067 );
xnor \U$4726 ( \5069 , \5068 , \1467 );
and \U$4727 ( \5070 , \5065 , \5069 );
and \U$4728 ( \5071 , \1588 , \1351 );
and \U$4729 ( \5072 , \1412 , \1349 );
nor \U$4730 ( \5073 , \5071 , \5072 );
xnor \U$4731 ( \5074 , \5073 , \1238 );
and \U$4732 ( \5075 , \5069 , \5074 );
and \U$4733 ( \5076 , \5065 , \5074 );
or \U$4734 ( \5077 , \5070 , \5075 , \5076 );
and \U$4735 ( \5078 , \1839 , \1157 );
and \U$4736 ( \5079 , \1596 , \1155 );
nor \U$4737 ( \5080 , \5078 , \5079 );
xnor \U$4738 ( \5081 , \5080 , \1021 );
and \U$4739 ( \5082 , \2030 , \957 );
and \U$4740 ( \5083 , \1844 , \955 );
nor \U$4741 ( \5084 , \5082 , \5083 );
xnor \U$4742 ( \5085 , \5084 , \879 );
and \U$4743 ( \5086 , \5081 , \5085 );
and \U$4744 ( \5087 , \2438 , \793 );
and \U$4745 ( \5088 , \2174 , \791 );
nor \U$4746 ( \5089 , \5087 , \5088 );
xnor \U$4747 ( \5090 , \5089 , \699 );
and \U$4748 ( \5091 , \5085 , \5090 );
and \U$4749 ( \5092 , \5081 , \5090 );
or \U$4750 ( \5093 , \5086 , \5091 , \5092 );
and \U$4751 ( \5094 , \5077 , \5093 );
and \U$4752 ( \5095 , \2637 , \624 );
and \U$4753 ( \5096 , \2463 , \622 );
nor \U$4754 ( \5097 , \5095 , \5096 );
xnor \U$4755 ( \5098 , \5097 , \349 );
and \U$4756 ( \5099 , \2942 , \357 );
and \U$4757 ( \5100 , \2804 , \355 );
nor \U$4758 ( \5101 , \5099 , \5100 );
xnor \U$4759 ( \5102 , \5101 , \364 );
and \U$4760 ( \5103 , \5098 , \5102 );
and \U$4761 ( \5104 , \3478 , \373 );
and \U$4762 ( \5105 , \3061 , \371 );
nor \U$4763 ( \5106 , \5104 , \5105 );
xnor \U$4764 ( \5107 , \5106 , \380 );
and \U$4765 ( \5108 , \5102 , \5107 );
and \U$4766 ( \5109 , \5098 , \5107 );
or \U$4767 ( \5110 , \5103 , \5108 , \5109 );
and \U$4768 ( \5111 , \5093 , \5110 );
and \U$4769 ( \5112 , \5077 , \5110 );
or \U$4770 ( \5113 , \5094 , \5111 , \5112 );
and \U$4771 ( \5114 , \5060 , \5113 );
and \U$4772 ( \5115 , \5028 , \5113 );
or \U$4773 ( \5116 , \5061 , \5114 , \5115 );
and \U$4774 ( \5117 , \5045 , \436 );
xor \U$4775 ( \5118 , \4879 , \4883 );
xor \U$4776 ( \5119 , \5118 , \4888 );
and \U$4777 ( \5120 , \5117 , \5119 );
xor \U$4778 ( \5121 , \4842 , \4846 );
xor \U$4779 ( \5122 , \5121 , \4851 );
and \U$4780 ( \5123 , \5119 , \5122 );
and \U$4781 ( \5124 , \5117 , \5122 );
or \U$4782 ( \5125 , \5120 , \5123 , \5124 );
xor \U$4783 ( \5126 , \4826 , \4830 );
xor \U$4784 ( \5127 , \5126 , \4835 );
xor \U$4785 ( \5128 , \4772 , \4776 );
xor \U$4786 ( \5129 , \5128 , \4781 );
and \U$4787 ( \5130 , \5127 , \5129 );
xor \U$4788 ( \5131 , \4859 , \4863 );
xor \U$4789 ( \5132 , \5131 , \4868 );
and \U$4790 ( \5133 , \5129 , \5132 );
and \U$4791 ( \5134 , \5127 , \5132 );
or \U$4792 ( \5135 , \5130 , \5133 , \5134 );
and \U$4793 ( \5136 , \5125 , \5135 );
xor \U$4794 ( \5137 , \4913 , \4915 );
xor \U$4795 ( \5138 , \5137 , \4918 );
and \U$4796 ( \5139 , \5135 , \5138 );
and \U$4797 ( \5140 , \5125 , \5138 );
or \U$4798 ( \5141 , \5136 , \5139 , \5140 );
and \U$4799 ( \5142 , \5116 , \5141 );
xor \U$4800 ( \5143 , \4838 , \4854 );
xor \U$4801 ( \5144 , \5143 , \4871 );
xor \U$4802 ( \5145 , \4903 , \4905 );
xor \U$4803 ( \5146 , \5145 , \4908 );
and \U$4804 ( \5147 , \5144 , \5146 );
xor \U$4805 ( \5148 , \4891 , \4893 );
xor \U$4806 ( \5149 , \5148 , \4895 );
and \U$4807 ( \5150 , \5146 , \5149 );
and \U$4808 ( \5151 , \5144 , \5149 );
or \U$4809 ( \5152 , \5147 , \5150 , \5151 );
and \U$4810 ( \5153 , \5141 , \5152 );
and \U$4811 ( \5154 , \5116 , \5152 );
or \U$4812 ( \5155 , \5142 , \5153 , \5154 );
xor \U$4813 ( \5156 , \4599 , \4618 );
xor \U$4814 ( \5157 , \5156 , \4635 );
xor \U$4815 ( \5158 , \4655 , \4671 );
xor \U$4816 ( \5159 , \5158 , \4688 );
and \U$4817 ( \5160 , \5157 , \5159 );
xor \U$4818 ( \5161 , \4930 , \4932 );
xor \U$4819 ( \5162 , \5161 , \4935 );
and \U$4820 ( \5163 , \5159 , \5162 );
and \U$4821 ( \5164 , \5157 , \5162 );
or \U$4822 ( \5165 , \5160 , \5163 , \5164 );
and \U$4823 ( \5166 , \5155 , \5165 );
xor \U$4824 ( \5167 , \4583 , \4638 );
xor \U$4825 ( \5168 , \5167 , \4691 );
and \U$4826 ( \5169 , \5165 , \5168 );
and \U$4827 ( \5170 , \5155 , \5168 );
or \U$4828 ( \5171 , \5166 , \5169 , \5170 );
xor \U$4829 ( \5172 , \4941 , \4951 );
xor \U$4830 ( \5173 , \5172 , \4954 );
and \U$4831 ( \5174 , \5171 , \5173 );
xor \U$4832 ( \5175 , \4959 , \4961 );
xor \U$4833 ( \5176 , \5175 , \4964 );
and \U$4834 ( \5177 , \5173 , \5176 );
and \U$4835 ( \5178 , \5171 , \5176 );
or \U$4836 ( \5179 , \5174 , \5177 , \5178 );
xor \U$4837 ( \5180 , \4957 , \4967 );
xor \U$4838 ( \5181 , \5180 , \4970 );
and \U$4839 ( \5182 , \5179 , \5181 );
xor \U$4840 ( \5183 , \4733 , \4743 );
xor \U$4841 ( \5184 , \5183 , \4746 );
and \U$4842 ( \5185 , \5181 , \5184 );
and \U$4843 ( \5186 , \5179 , \5184 );
or \U$4844 ( \5187 , \5182 , \5185 , \5186 );
and \U$4845 ( \5188 , \4973 , \5187 );
xor \U$4846 ( \5189 , \4749 , \4751 );
xor \U$4847 ( \5190 , \5189 , \4753 );
and \U$4848 ( \5191 , \5187 , \5190 );
and \U$4849 ( \5192 , \4973 , \5190 );
or \U$4850 ( \5193 , \5188 , \5191 , \5192 );
and \U$4851 ( \5194 , \4768 , \5193 );
xor \U$4852 ( \5195 , \4768 , \5193 );
xor \U$4853 ( \5196 , \4973 , \5187 );
xor \U$4854 ( \5197 , \5196 , \5190 );
buf \U$4855 ( \5198 , RIbb2e0f8_46);
buf \U$4856 ( \5199 , RIbb2e080_47);
and \U$4857 ( \5200 , \5198 , \5199 );
not \U$4858 ( \5201 , \5200 );
and \U$4859 ( \5202 , \4786 , \5201 );
not \U$4860 ( \5203 , \5202 );
and \U$4861 ( \5204 , \351 , \4977 );
and \U$4862 ( \5205 , \359 , \4975 );
nor \U$4863 ( \5206 , \5204 , \5205 );
xnor \U$4864 ( \5207 , \5206 , \4789 );
and \U$4865 ( \5208 , \5203 , \5207 );
and \U$4866 ( \5209 , \367 , \4603 );
and \U$4867 ( \5210 , \375 , \4601 );
nor \U$4868 ( \5211 , \5209 , \5210 );
xnor \U$4869 ( \5212 , \5211 , \4371 );
and \U$4870 ( \5213 , \5207 , \5212 );
and \U$4871 ( \5214 , \5203 , \5212 );
or \U$4872 ( \5215 , \5208 , \5213 , \5214 );
and \U$4873 ( \5216 , \385 , \4152 );
and \U$4874 ( \5217 , \393 , \4150 );
nor \U$4875 ( \5218 , \5216 , \5217 );
xnor \U$4876 ( \5219 , \5218 , \4009 );
and \U$4877 ( \5220 , \400 , \3829 );
and \U$4878 ( \5221 , \408 , \3827 );
nor \U$4879 ( \5222 , \5220 , \5221 );
xnor \U$4880 ( \5223 , \5222 , \3583 );
and \U$4881 ( \5224 , \5219 , \5223 );
and \U$4882 ( \5225 , \416 , \3434 );
and \U$4883 ( \5226 , \424 , \3432 );
nor \U$4884 ( \5227 , \5225 , \5226 );
xnor \U$4885 ( \5228 , \5227 , \3247 );
and \U$4886 ( \5229 , \5223 , \5228 );
and \U$4887 ( \5230 , \5219 , \5228 );
or \U$4888 ( \5231 , \5224 , \5229 , \5230 );
and \U$4889 ( \5232 , \5215 , \5231 );
and \U$4890 ( \5233 , \435 , \3121 );
and \U$4891 ( \5234 , \443 , \3119 );
nor \U$4892 ( \5235 , \5233 , \5234 );
xnor \U$4893 ( \5236 , \5235 , \2916 );
and \U$4894 ( \5237 , \661 , \2715 );
and \U$4895 ( \5238 , \450 , \2713 );
nor \U$4896 ( \5239 , \5237 , \5238 );
xnor \U$4897 ( \5240 , \5239 , \2566 );
and \U$4898 ( \5241 , \5236 , \5240 );
and \U$4899 ( \5242 , \785 , \2393 );
and \U$4900 ( \5243 , \722 , \2391 );
nor \U$4901 ( \5244 , \5242 , \5243 );
xnor \U$4902 ( \5245 , \5244 , \2251 );
and \U$4903 ( \5246 , \5240 , \5245 );
and \U$4904 ( \5247 , \5236 , \5245 );
or \U$4905 ( \5248 , \5241 , \5246 , \5247 );
and \U$4906 ( \5249 , \5231 , \5248 );
and \U$4907 ( \5250 , \5215 , \5248 );
or \U$4908 ( \5251 , \5232 , \5249 , \5250 );
and \U$4909 ( \5252 , \1071 , \2097 );
and \U$4910 ( \5253 , \983 , \2095 );
nor \U$4911 ( \5254 , \5252 , \5253 );
xnor \U$4912 ( \5255 , \5254 , \1960 );
and \U$4913 ( \5256 , \1181 , \1891 );
and \U$4914 ( \5257 , \1176 , \1889 );
nor \U$4915 ( \5258 , \5256 , \5257 );
xnor \U$4916 ( \5259 , \5258 , \1739 );
and \U$4917 ( \5260 , \5255 , \5259 );
and \U$4918 ( \5261 , \1412 , \1623 );
and \U$4919 ( \5262 , \1297 , \1621 );
nor \U$4920 ( \5263 , \5261 , \5262 );
xnor \U$4921 ( \5264 , \5263 , \1467 );
and \U$4922 ( \5265 , \5259 , \5264 );
and \U$4923 ( \5266 , \5255 , \5264 );
or \U$4924 ( \5267 , \5260 , \5265 , \5266 );
and \U$4925 ( \5268 , \1596 , \1351 );
and \U$4926 ( \5269 , \1588 , \1349 );
nor \U$4927 ( \5270 , \5268 , \5269 );
xnor \U$4928 ( \5271 , \5270 , \1238 );
and \U$4929 ( \5272 , \1844 , \1157 );
and \U$4930 ( \5273 , \1839 , \1155 );
nor \U$4931 ( \5274 , \5272 , \5273 );
xnor \U$4932 ( \5275 , \5274 , \1021 );
and \U$4933 ( \5276 , \5271 , \5275 );
and \U$4934 ( \5277 , \2174 , \957 );
and \U$4935 ( \5278 , \2030 , \955 );
nor \U$4936 ( \5279 , \5277 , \5278 );
xnor \U$4937 ( \5280 , \5279 , \879 );
and \U$4938 ( \5281 , \5275 , \5280 );
and \U$4939 ( \5282 , \5271 , \5280 );
or \U$4940 ( \5283 , \5276 , \5281 , \5282 );
and \U$4941 ( \5284 , \5267 , \5283 );
and \U$4942 ( \5285 , \2463 , \793 );
and \U$4943 ( \5286 , \2438 , \791 );
nor \U$4944 ( \5287 , \5285 , \5286 );
xnor \U$4945 ( \5288 , \5287 , \699 );
and \U$4946 ( \5289 , \2804 , \624 );
and \U$4947 ( \5290 , \2637 , \622 );
nor \U$4948 ( \5291 , \5289 , \5290 );
xnor \U$4949 ( \5292 , \5291 , \349 );
and \U$4950 ( \5293 , \5288 , \5292 );
and \U$4951 ( \5294 , \3061 , \357 );
and \U$4952 ( \5295 , \2942 , \355 );
nor \U$4953 ( \5296 , \5294 , \5295 );
xnor \U$4954 ( \5297 , \5296 , \364 );
and \U$4955 ( \5298 , \5292 , \5297 );
and \U$4956 ( \5299 , \5288 , \5297 );
or \U$4957 ( \5300 , \5293 , \5298 , \5299 );
and \U$4958 ( \5301 , \5283 , \5300 );
and \U$4959 ( \5302 , \5267 , \5300 );
or \U$4960 ( \5303 , \5284 , \5301 , \5302 );
and \U$4961 ( \5304 , \5251 , \5303 );
and \U$4962 ( \5305 , \4576 , \422 );
and \U$4963 ( \5306 , \4568 , \420 );
nor \U$4964 ( \5307 , \5305 , \5306 );
xnor \U$4965 ( \5308 , \5307 , \429 );
and \U$4966 ( \5309 , \5050 , \441 );
and \U$4967 ( \5310 , \5045 , \439 );
nor \U$4968 ( \5311 , \5309 , \5310 );
xnor \U$4969 ( \5312 , \5311 , \448 );
and \U$4970 ( \5313 , \5308 , \5312 );
buf \U$4971 ( \5314 , RIbb2c370_109);
and \U$4972 ( \5315 , \5314 , \436 );
and \U$4973 ( \5316 , \5312 , \5315 );
and \U$4974 ( \5317 , \5308 , \5315 );
or \U$4975 ( \5318 , \5313 , \5316 , \5317 );
and \U$4976 ( \5319 , \3686 , \373 );
and \U$4977 ( \5320 , \3478 , \371 );
nor \U$4978 ( \5321 , \5319 , \5320 );
xnor \U$4979 ( \5322 , \5321 , \380 );
and \U$4980 ( \5323 , \3813 , \391 );
and \U$4981 ( \5324 , \3808 , \389 );
nor \U$4982 ( \5325 , \5323 , \5324 );
xnor \U$4983 ( \5326 , \5325 , \398 );
and \U$4984 ( \5327 , \5322 , \5326 );
and \U$4985 ( \5328 , \4266 , \406 );
and \U$4986 ( \5329 , \4069 , \404 );
nor \U$4987 ( \5330 , \5328 , \5329 );
xnor \U$4988 ( \5331 , \5330 , \413 );
and \U$4989 ( \5332 , \5326 , \5331 );
and \U$4990 ( \5333 , \5322 , \5331 );
or \U$4991 ( \5334 , \5327 , \5332 , \5333 );
and \U$4992 ( \5335 , \5318 , \5334 );
xnor \U$4993 ( \5336 , \5049 , \5051 );
and \U$4994 ( \5337 , \5334 , \5336 );
and \U$4995 ( \5338 , \5318 , \5336 );
or \U$4996 ( \5339 , \5335 , \5337 , \5338 );
and \U$4997 ( \5340 , \5303 , \5339 );
and \U$4998 ( \5341 , \5251 , \5339 );
or \U$4999 ( \5342 , \5304 , \5340 , \5341 );
xor \U$5000 ( \5343 , \5032 , \5036 );
xor \U$5001 ( \5344 , \5343 , \5041 );
xor \U$5002 ( \5345 , \5081 , \5085 );
xor \U$5003 ( \5346 , \5345 , \5090 );
and \U$5004 ( \5347 , \5344 , \5346 );
xor \U$5005 ( \5348 , \5098 , \5102 );
xor \U$5006 ( \5349 , \5348 , \5107 );
and \U$5007 ( \5350 , \5346 , \5349 );
and \U$5008 ( \5351 , \5344 , \5349 );
or \U$5009 ( \5352 , \5347 , \5350 , \5351 );
xor \U$5010 ( \5353 , \5065 , \5069 );
xor \U$5011 ( \5354 , \5353 , \5074 );
xor \U$5012 ( \5355 , \4996 , \5000 );
xor \U$5013 ( \5356 , \5355 , \5005 );
and \U$5014 ( \5357 , \5354 , \5356 );
xor \U$5015 ( \5358 , \5013 , \5017 );
xor \U$5016 ( \5359 , \5358 , \5022 );
and \U$5017 ( \5360 , \5356 , \5359 );
and \U$5018 ( \5361 , \5354 , \5359 );
or \U$5019 ( \5362 , \5357 , \5360 , \5361 );
and \U$5020 ( \5363 , \5352 , \5362 );
xor \U$5021 ( \5364 , \4807 , \4811 );
xor \U$5022 ( \5365 , \5364 , \4816 );
and \U$5023 ( \5366 , \5362 , \5365 );
and \U$5024 ( \5367 , \5352 , \5365 );
or \U$5025 ( \5368 , \5363 , \5366 , \5367 );
and \U$5026 ( \5369 , \5342 , \5368 );
xor \U$5027 ( \5370 , \4790 , \4794 );
xor \U$5028 ( \5371 , \5370 , \4799 );
xor \U$5029 ( \5372 , \5117 , \5119 );
xor \U$5030 ( \5373 , \5372 , \5122 );
and \U$5031 ( \5374 , \5371 , \5373 );
xor \U$5032 ( \5375 , \5127 , \5129 );
xor \U$5033 ( \5376 , \5375 , \5132 );
and \U$5034 ( \5377 , \5373 , \5376 );
and \U$5035 ( \5378 , \5371 , \5376 );
or \U$5036 ( \5379 , \5374 , \5377 , \5378 );
and \U$5037 ( \5380 , \5368 , \5379 );
and \U$5038 ( \5381 , \5342 , \5379 );
or \U$5039 ( \5382 , \5369 , \5380 , \5381 );
xor \U$5040 ( \5383 , \4992 , \5008 );
xor \U$5041 ( \5384 , \5383 , \5025 );
xor \U$5042 ( \5385 , \5044 , \5052 );
xor \U$5043 ( \5386 , \5385 , \5057 );
and \U$5044 ( \5387 , \5384 , \5386 );
xor \U$5045 ( \5388 , \5077 , \5093 );
xor \U$5046 ( \5389 , \5388 , \5110 );
and \U$5047 ( \5390 , \5386 , \5389 );
and \U$5048 ( \5391 , \5384 , \5389 );
or \U$5049 ( \5392 , \5387 , \5390 , \5391 );
xor \U$5050 ( \5393 , \4784 , \4802 );
xor \U$5051 ( \5394 , \5393 , \4819 );
and \U$5052 ( \5395 , \5392 , \5394 );
xor \U$5053 ( \5396 , \5144 , \5146 );
xor \U$5054 ( \5397 , \5396 , \5149 );
and \U$5055 ( \5398 , \5394 , \5397 );
and \U$5056 ( \5399 , \5392 , \5397 );
or \U$5057 ( \5400 , \5395 , \5398 , \5399 );
and \U$5058 ( \5401 , \5382 , \5400 );
xor \U$5059 ( \5402 , \4911 , \4921 );
xor \U$5060 ( \5403 , \5402 , \4924 );
and \U$5061 ( \5404 , \5400 , \5403 );
and \U$5062 ( \5405 , \5382 , \5403 );
or \U$5063 ( \5406 , \5401 , \5404 , \5405 );
xor \U$5064 ( \5407 , \4822 , \4874 );
xor \U$5065 ( \5408 , \5407 , \4898 );
xor \U$5066 ( \5409 , \5116 , \5141 );
xor \U$5067 ( \5410 , \5409 , \5152 );
and \U$5068 ( \5411 , \5408 , \5410 );
xor \U$5069 ( \5412 , \5157 , \5159 );
xor \U$5070 ( \5413 , \5412 , \5162 );
and \U$5071 ( \5414 , \5410 , \5413 );
and \U$5072 ( \5415 , \5408 , \5413 );
or \U$5073 ( \5416 , \5411 , \5414 , \5415 );
and \U$5074 ( \5417 , \5406 , \5416 );
xor \U$5075 ( \5418 , \4943 , \4945 );
xor \U$5076 ( \5419 , \5418 , \4948 );
and \U$5077 ( \5420 , \5416 , \5419 );
and \U$5078 ( \5421 , \5406 , \5419 );
or \U$5079 ( \5422 , \5417 , \5420 , \5421 );
xor \U$5080 ( \5423 , \4901 , \4927 );
xor \U$5081 ( \5424 , \5423 , \4938 );
xor \U$5082 ( \5425 , \5155 , \5165 );
xor \U$5083 ( \5426 , \5425 , \5168 );
and \U$5084 ( \5427 , \5424 , \5426 );
and \U$5085 ( \5428 , \5422 , \5427 );
xor \U$5086 ( \5429 , \5171 , \5173 );
xor \U$5087 ( \5430 , \5429 , \5176 );
and \U$5088 ( \5431 , \5427 , \5430 );
and \U$5089 ( \5432 , \5422 , \5430 );
or \U$5090 ( \5433 , \5428 , \5431 , \5432 );
xor \U$5091 ( \5434 , \5179 , \5181 );
xor \U$5092 ( \5435 , \5434 , \5184 );
and \U$5093 ( \5436 , \5433 , \5435 );
and \U$5094 ( \5437 , \5197 , \5436 );
xor \U$5095 ( \5438 , \5197 , \5436 );
xor \U$5096 ( \5439 , \5433 , \5435 );
xor \U$5097 ( \5440 , \4786 , \5198 );
xor \U$5098 ( \5441 , \5198 , \5199 );
not \U$5099 ( \5442 , \5441 );
and \U$5100 ( \5443 , \5440 , \5442 );
and \U$5101 ( \5444 , \359 , \5443 );
not \U$5102 ( \5445 , \5444 );
xnor \U$5103 ( \5446 , \5445 , \5202 );
and \U$5104 ( \5447 , \375 , \4977 );
and \U$5105 ( \5448 , \351 , \4975 );
nor \U$5106 ( \5449 , \5447 , \5448 );
xnor \U$5107 ( \5450 , \5449 , \4789 );
and \U$5108 ( \5451 , \5446 , \5450 );
and \U$5109 ( \5452 , \393 , \4603 );
and \U$5110 ( \5453 , \367 , \4601 );
nor \U$5111 ( \5454 , \5452 , \5453 );
xnor \U$5112 ( \5455 , \5454 , \4371 );
and \U$5113 ( \5456 , \5450 , \5455 );
and \U$5114 ( \5457 , \5446 , \5455 );
or \U$5115 ( \5458 , \5451 , \5456 , \5457 );
and \U$5116 ( \5459 , \408 , \4152 );
and \U$5117 ( \5460 , \385 , \4150 );
nor \U$5118 ( \5461 , \5459 , \5460 );
xnor \U$5119 ( \5462 , \5461 , \4009 );
and \U$5120 ( \5463 , \424 , \3829 );
and \U$5121 ( \5464 , \400 , \3827 );
nor \U$5122 ( \5465 , \5463 , \5464 );
xnor \U$5123 ( \5466 , \5465 , \3583 );
and \U$5124 ( \5467 , \5462 , \5466 );
and \U$5125 ( \5468 , \443 , \3434 );
and \U$5126 ( \5469 , \416 , \3432 );
nor \U$5127 ( \5470 , \5468 , \5469 );
xnor \U$5128 ( \5471 , \5470 , \3247 );
and \U$5129 ( \5472 , \5466 , \5471 );
and \U$5130 ( \5473 , \5462 , \5471 );
or \U$5131 ( \5474 , \5467 , \5472 , \5473 );
and \U$5132 ( \5475 , \5458 , \5474 );
and \U$5133 ( \5476 , \450 , \3121 );
and \U$5134 ( \5477 , \435 , \3119 );
nor \U$5135 ( \5478 , \5476 , \5477 );
xnor \U$5136 ( \5479 , \5478 , \2916 );
and \U$5137 ( \5480 , \722 , \2715 );
and \U$5138 ( \5481 , \661 , \2713 );
nor \U$5139 ( \5482 , \5480 , \5481 );
xnor \U$5140 ( \5483 , \5482 , \2566 );
and \U$5141 ( \5484 , \5479 , \5483 );
and \U$5142 ( \5485 , \983 , \2393 );
and \U$5143 ( \5486 , \785 , \2391 );
nor \U$5144 ( \5487 , \5485 , \5486 );
xnor \U$5145 ( \5488 , \5487 , \2251 );
and \U$5146 ( \5489 , \5483 , \5488 );
and \U$5147 ( \5490 , \5479 , \5488 );
or \U$5148 ( \5491 , \5484 , \5489 , \5490 );
and \U$5149 ( \5492 , \5474 , \5491 );
and \U$5150 ( \5493 , \5458 , \5491 );
or \U$5151 ( \5494 , \5475 , \5492 , \5493 );
and \U$5152 ( \5495 , \1176 , \2097 );
and \U$5153 ( \5496 , \1071 , \2095 );
nor \U$5154 ( \5497 , \5495 , \5496 );
xnor \U$5155 ( \5498 , \5497 , \1960 );
and \U$5156 ( \5499 , \1297 , \1891 );
and \U$5157 ( \5500 , \1181 , \1889 );
nor \U$5158 ( \5501 , \5499 , \5500 );
xnor \U$5159 ( \5502 , \5501 , \1739 );
and \U$5160 ( \5503 , \5498 , \5502 );
and \U$5161 ( \5504 , \1588 , \1623 );
and \U$5162 ( \5505 , \1412 , \1621 );
nor \U$5163 ( \5506 , \5504 , \5505 );
xnor \U$5164 ( \5507 , \5506 , \1467 );
and \U$5165 ( \5508 , \5502 , \5507 );
and \U$5166 ( \5509 , \5498 , \5507 );
or \U$5167 ( \5510 , \5503 , \5508 , \5509 );
and \U$5168 ( \5511 , \1839 , \1351 );
and \U$5169 ( \5512 , \1596 , \1349 );
nor \U$5170 ( \5513 , \5511 , \5512 );
xnor \U$5171 ( \5514 , \5513 , \1238 );
and \U$5172 ( \5515 , \2030 , \1157 );
and \U$5173 ( \5516 , \1844 , \1155 );
nor \U$5174 ( \5517 , \5515 , \5516 );
xnor \U$5175 ( \5518 , \5517 , \1021 );
and \U$5176 ( \5519 , \5514 , \5518 );
and \U$5177 ( \5520 , \2438 , \957 );
and \U$5178 ( \5521 , \2174 , \955 );
nor \U$5179 ( \5522 , \5520 , \5521 );
xnor \U$5180 ( \5523 , \5522 , \879 );
and \U$5181 ( \5524 , \5518 , \5523 );
and \U$5182 ( \5525 , \5514 , \5523 );
or \U$5183 ( \5526 , \5519 , \5524 , \5525 );
and \U$5184 ( \5527 , \5510 , \5526 );
and \U$5185 ( \5528 , \2637 , \793 );
and \U$5186 ( \5529 , \2463 , \791 );
nor \U$5187 ( \5530 , \5528 , \5529 );
xnor \U$5188 ( \5531 , \5530 , \699 );
and \U$5189 ( \5532 , \2942 , \624 );
and \U$5190 ( \5533 , \2804 , \622 );
nor \U$5191 ( \5534 , \5532 , \5533 );
xnor \U$5192 ( \5535 , \5534 , \349 );
and \U$5193 ( \5536 , \5531 , \5535 );
and \U$5194 ( \5537 , \3478 , \357 );
and \U$5195 ( \5538 , \3061 , \355 );
nor \U$5196 ( \5539 , \5537 , \5538 );
xnor \U$5197 ( \5540 , \5539 , \364 );
and \U$5198 ( \5541 , \5535 , \5540 );
and \U$5199 ( \5542 , \5531 , \5540 );
or \U$5200 ( \5543 , \5536 , \5541 , \5542 );
and \U$5201 ( \5544 , \5526 , \5543 );
and \U$5202 ( \5545 , \5510 , \5543 );
or \U$5203 ( \5546 , \5527 , \5544 , \5545 );
and \U$5204 ( \5547 , \5494 , \5546 );
and \U$5205 ( \5548 , \3808 , \373 );
and \U$5206 ( \5549 , \3686 , \371 );
nor \U$5207 ( \5550 , \5548 , \5549 );
xnor \U$5208 ( \5551 , \5550 , \380 );
and \U$5209 ( \5552 , \4069 , \391 );
and \U$5210 ( \5553 , \3813 , \389 );
nor \U$5211 ( \5554 , \5552 , \5553 );
xnor \U$5212 ( \5555 , \5554 , \398 );
and \U$5213 ( \5556 , \5551 , \5555 );
and \U$5214 ( \5557 , \4568 , \406 );
and \U$5215 ( \5558 , \4266 , \404 );
nor \U$5216 ( \5559 , \5557 , \5558 );
xnor \U$5217 ( \5560 , \5559 , \413 );
and \U$5218 ( \5561 , \5555 , \5560 );
and \U$5219 ( \5562 , \5551 , \5560 );
or \U$5220 ( \5563 , \5556 , \5561 , \5562 );
and \U$5221 ( \5564 , \5045 , \422 );
and \U$5222 ( \5565 , \4576 , \420 );
nor \U$5223 ( \5566 , \5564 , \5565 );
xnor \U$5224 ( \5567 , \5566 , \429 );
and \U$5225 ( \5568 , \5314 , \441 );
and \U$5226 ( \5569 , \5050 , \439 );
nor \U$5227 ( \5570 , \5568 , \5569 );
xnor \U$5228 ( \5571 , \5570 , \448 );
and \U$5229 ( \5572 , \5567 , \5571 );
buf \U$5230 ( \5573 , RIbb2c2f8_110);
and \U$5231 ( \5574 , \5573 , \436 );
and \U$5232 ( \5575 , \5571 , \5574 );
and \U$5233 ( \5576 , \5567 , \5574 );
or \U$5234 ( \5577 , \5572 , \5575 , \5576 );
and \U$5235 ( \5578 , \5563 , \5577 );
xor \U$5236 ( \5579 , \5308 , \5312 );
xor \U$5237 ( \5580 , \5579 , \5315 );
and \U$5238 ( \5581 , \5577 , \5580 );
and \U$5239 ( \5582 , \5563 , \5580 );
or \U$5240 ( \5583 , \5578 , \5581 , \5582 );
and \U$5241 ( \5584 , \5546 , \5583 );
and \U$5242 ( \5585 , \5494 , \5583 );
or \U$5243 ( \5586 , \5547 , \5584 , \5585 );
xor \U$5244 ( \5587 , \5255 , \5259 );
xor \U$5245 ( \5588 , \5587 , \5264 );
xor \U$5246 ( \5589 , \5219 , \5223 );
xor \U$5247 ( \5590 , \5589 , \5228 );
and \U$5248 ( \5591 , \5588 , \5590 );
xor \U$5249 ( \5592 , \5236 , \5240 );
xor \U$5250 ( \5593 , \5592 , \5245 );
and \U$5251 ( \5594 , \5590 , \5593 );
and \U$5252 ( \5595 , \5588 , \5593 );
or \U$5253 ( \5596 , \5591 , \5594 , \5595 );
xor \U$5254 ( \5597 , \5271 , \5275 );
xor \U$5255 ( \5598 , \5597 , \5280 );
xor \U$5256 ( \5599 , \5288 , \5292 );
xor \U$5257 ( \5600 , \5599 , \5297 );
and \U$5258 ( \5601 , \5598 , \5600 );
xor \U$5259 ( \5602 , \5322 , \5326 );
xor \U$5260 ( \5603 , \5602 , \5331 );
and \U$5261 ( \5604 , \5600 , \5603 );
and \U$5262 ( \5605 , \5598 , \5603 );
or \U$5263 ( \5606 , \5601 , \5604 , \5605 );
and \U$5264 ( \5607 , \5596 , \5606 );
xor \U$5265 ( \5608 , \4980 , \4984 );
xor \U$5266 ( \5609 , \5608 , \4989 );
and \U$5267 ( \5610 , \5606 , \5609 );
and \U$5268 ( \5611 , \5596 , \5609 );
or \U$5269 ( \5612 , \5607 , \5610 , \5611 );
and \U$5270 ( \5613 , \5586 , \5612 );
xor \U$5271 ( \5614 , \5344 , \5346 );
xor \U$5272 ( \5615 , \5614 , \5349 );
xor \U$5273 ( \5616 , \5354 , \5356 );
xor \U$5274 ( \5617 , \5616 , \5359 );
and \U$5275 ( \5618 , \5615 , \5617 );
xor \U$5276 ( \5619 , \5318 , \5334 );
xor \U$5277 ( \5620 , \5619 , \5336 );
and \U$5278 ( \5621 , \5617 , \5620 );
and \U$5279 ( \5622 , \5615 , \5620 );
or \U$5280 ( \5623 , \5618 , \5621 , \5622 );
and \U$5281 ( \5624 , \5612 , \5623 );
and \U$5282 ( \5625 , \5586 , \5623 );
or \U$5283 ( \5626 , \5613 , \5624 , \5625 );
xor \U$5284 ( \5627 , \5352 , \5362 );
xor \U$5285 ( \5628 , \5627 , \5365 );
xor \U$5286 ( \5629 , \5384 , \5386 );
xor \U$5287 ( \5630 , \5629 , \5389 );
and \U$5288 ( \5631 , \5628 , \5630 );
xor \U$5289 ( \5632 , \5371 , \5373 );
xor \U$5290 ( \5633 , \5632 , \5376 );
and \U$5291 ( \5634 , \5630 , \5633 );
and \U$5292 ( \5635 , \5628 , \5633 );
or \U$5293 ( \5636 , \5631 , \5634 , \5635 );
and \U$5294 ( \5637 , \5626 , \5636 );
xor \U$5295 ( \5638 , \5125 , \5135 );
xor \U$5296 ( \5639 , \5638 , \5138 );
and \U$5297 ( \5640 , \5636 , \5639 );
and \U$5298 ( \5641 , \5626 , \5639 );
or \U$5299 ( \5642 , \5637 , \5640 , \5641 );
xor \U$5300 ( \5643 , \5028 , \5060 );
xor \U$5301 ( \5644 , \5643 , \5113 );
xor \U$5302 ( \5645 , \5342 , \5368 );
xor \U$5303 ( \5646 , \5645 , \5379 );
and \U$5304 ( \5647 , \5644 , \5646 );
xor \U$5305 ( \5648 , \5392 , \5394 );
xor \U$5306 ( \5649 , \5648 , \5397 );
and \U$5307 ( \5650 , \5646 , \5649 );
and \U$5308 ( \5651 , \5644 , \5649 );
or \U$5309 ( \5652 , \5647 , \5650 , \5651 );
and \U$5310 ( \5653 , \5642 , \5652 );
xor \U$5311 ( \5654 , \5408 , \5410 );
xor \U$5312 ( \5655 , \5654 , \5413 );
and \U$5313 ( \5656 , \5652 , \5655 );
and \U$5314 ( \5657 , \5642 , \5655 );
or \U$5315 ( \5658 , \5653 , \5656 , \5657 );
xor \U$5316 ( \5659 , \5406 , \5416 );
xor \U$5317 ( \5660 , \5659 , \5419 );
and \U$5318 ( \5661 , \5658 , \5660 );
xor \U$5319 ( \5662 , \5424 , \5426 );
and \U$5320 ( \5663 , \5660 , \5662 );
and \U$5321 ( \5664 , \5658 , \5662 );
or \U$5322 ( \5665 , \5661 , \5663 , \5664 );
xor \U$5323 ( \5666 , \5422 , \5427 );
xor \U$5324 ( \5667 , \5666 , \5430 );
and \U$5325 ( \5668 , \5665 , \5667 );
and \U$5326 ( \5669 , \5439 , \5668 );
xor \U$5327 ( \5670 , \5439 , \5668 );
xor \U$5328 ( \5671 , \5665 , \5667 );
and \U$5329 ( \5672 , \385 , \4603 );
and \U$5330 ( \5673 , \393 , \4601 );
nor \U$5331 ( \5674 , \5672 , \5673 );
xnor \U$5332 ( \5675 , \5674 , \4371 );
and \U$5333 ( \5676 , \400 , \4152 );
and \U$5334 ( \5677 , \408 , \4150 );
nor \U$5335 ( \5678 , \5676 , \5677 );
xnor \U$5336 ( \5679 , \5678 , \4009 );
and \U$5337 ( \5680 , \5675 , \5679 );
and \U$5338 ( \5681 , \416 , \3829 );
and \U$5339 ( \5682 , \424 , \3827 );
nor \U$5340 ( \5683 , \5681 , \5682 );
xnor \U$5341 ( \5684 , \5683 , \3583 );
and \U$5342 ( \5685 , \5679 , \5684 );
and \U$5343 ( \5686 , \5675 , \5684 );
or \U$5344 ( \5687 , \5680 , \5685 , \5686 );
buf \U$5345 ( \5688 , RIbb2e008_48);
buf \U$5346 ( \5689 , RIbb2df90_49);
and \U$5347 ( \5690 , \5688 , \5689 );
not \U$5348 ( \5691 , \5690 );
and \U$5349 ( \5692 , \5199 , \5691 );
not \U$5350 ( \5693 , \5692 );
and \U$5351 ( \5694 , \351 , \5443 );
and \U$5352 ( \5695 , \359 , \5441 );
nor \U$5353 ( \5696 , \5694 , \5695 );
xnor \U$5354 ( \5697 , \5696 , \5202 );
and \U$5355 ( \5698 , \5693 , \5697 );
and \U$5356 ( \5699 , \367 , \4977 );
and \U$5357 ( \5700 , \375 , \4975 );
nor \U$5358 ( \5701 , \5699 , \5700 );
xnor \U$5359 ( \5702 , \5701 , \4789 );
and \U$5360 ( \5703 , \5697 , \5702 );
and \U$5361 ( \5704 , \5693 , \5702 );
or \U$5362 ( \5705 , \5698 , \5703 , \5704 );
and \U$5363 ( \5706 , \5687 , \5705 );
and \U$5364 ( \5707 , \435 , \3434 );
and \U$5365 ( \5708 , \443 , \3432 );
nor \U$5366 ( \5709 , \5707 , \5708 );
xnor \U$5367 ( \5710 , \5709 , \3247 );
and \U$5368 ( \5711 , \661 , \3121 );
and \U$5369 ( \5712 , \450 , \3119 );
nor \U$5370 ( \5713 , \5711 , \5712 );
xnor \U$5371 ( \5714 , \5713 , \2916 );
and \U$5372 ( \5715 , \5710 , \5714 );
and \U$5373 ( \5716 , \785 , \2715 );
and \U$5374 ( \5717 , \722 , \2713 );
nor \U$5375 ( \5718 , \5716 , \5717 );
xnor \U$5376 ( \5719 , \5718 , \2566 );
and \U$5377 ( \5720 , \5714 , \5719 );
and \U$5378 ( \5721 , \5710 , \5719 );
or \U$5379 ( \5722 , \5715 , \5720 , \5721 );
and \U$5380 ( \5723 , \5705 , \5722 );
and \U$5381 ( \5724 , \5687 , \5722 );
or \U$5382 ( \5725 , \5706 , \5723 , \5724 );
and \U$5383 ( \5726 , \2463 , \957 );
and \U$5384 ( \5727 , \2438 , \955 );
nor \U$5385 ( \5728 , \5726 , \5727 );
xnor \U$5386 ( \5729 , \5728 , \879 );
and \U$5387 ( \5730 , \2804 , \793 );
and \U$5388 ( \5731 , \2637 , \791 );
nor \U$5389 ( \5732 , \5730 , \5731 );
xnor \U$5390 ( \5733 , \5732 , \699 );
and \U$5391 ( \5734 , \5729 , \5733 );
and \U$5392 ( \5735 , \3061 , \624 );
and \U$5393 ( \5736 , \2942 , \622 );
nor \U$5394 ( \5737 , \5735 , \5736 );
xnor \U$5395 ( \5738 , \5737 , \349 );
and \U$5396 ( \5739 , \5733 , \5738 );
and \U$5397 ( \5740 , \5729 , \5738 );
or \U$5398 ( \5741 , \5734 , \5739 , \5740 );
and \U$5399 ( \5742 , \1596 , \1623 );
and \U$5400 ( \5743 , \1588 , \1621 );
nor \U$5401 ( \5744 , \5742 , \5743 );
xnor \U$5402 ( \5745 , \5744 , \1467 );
and \U$5403 ( \5746 , \1844 , \1351 );
and \U$5404 ( \5747 , \1839 , \1349 );
nor \U$5405 ( \5748 , \5746 , \5747 );
xnor \U$5406 ( \5749 , \5748 , \1238 );
and \U$5407 ( \5750 , \5745 , \5749 );
and \U$5408 ( \5751 , \2174 , \1157 );
and \U$5409 ( \5752 , \2030 , \1155 );
nor \U$5410 ( \5753 , \5751 , \5752 );
xnor \U$5411 ( \5754 , \5753 , \1021 );
and \U$5412 ( \5755 , \5749 , \5754 );
and \U$5413 ( \5756 , \5745 , \5754 );
or \U$5414 ( \5757 , \5750 , \5755 , \5756 );
and \U$5415 ( \5758 , \5741 , \5757 );
and \U$5416 ( \5759 , \1071 , \2393 );
and \U$5417 ( \5760 , \983 , \2391 );
nor \U$5418 ( \5761 , \5759 , \5760 );
xnor \U$5419 ( \5762 , \5761 , \2251 );
and \U$5420 ( \5763 , \1181 , \2097 );
and \U$5421 ( \5764 , \1176 , \2095 );
nor \U$5422 ( \5765 , \5763 , \5764 );
xnor \U$5423 ( \5766 , \5765 , \1960 );
and \U$5424 ( \5767 , \5762 , \5766 );
and \U$5425 ( \5768 , \1412 , \1891 );
and \U$5426 ( \5769 , \1297 , \1889 );
nor \U$5427 ( \5770 , \5768 , \5769 );
xnor \U$5428 ( \5771 , \5770 , \1739 );
and \U$5429 ( \5772 , \5766 , \5771 );
and \U$5430 ( \5773 , \5762 , \5771 );
or \U$5431 ( \5774 , \5767 , \5772 , \5773 );
and \U$5432 ( \5775 , \5757 , \5774 );
and \U$5433 ( \5776 , \5741 , \5774 );
or \U$5434 ( \5777 , \5758 , \5775 , \5776 );
and \U$5435 ( \5778 , \5725 , \5777 );
and \U$5436 ( \5779 , \3686 , \357 );
and \U$5437 ( \5780 , \3478 , \355 );
nor \U$5438 ( \5781 , \5779 , \5780 );
xnor \U$5439 ( \5782 , \5781 , \364 );
and \U$5440 ( \5783 , \3813 , \373 );
and \U$5441 ( \5784 , \3808 , \371 );
nor \U$5442 ( \5785 , \5783 , \5784 );
xnor \U$5443 ( \5786 , \5785 , \380 );
and \U$5444 ( \5787 , \5782 , \5786 );
and \U$5445 ( \5788 , \4266 , \391 );
and \U$5446 ( \5789 , \4069 , \389 );
nor \U$5447 ( \5790 , \5788 , \5789 );
xnor \U$5448 ( \5791 , \5790 , \398 );
and \U$5449 ( \5792 , \5786 , \5791 );
and \U$5450 ( \5793 , \5782 , \5791 );
or \U$5451 ( \5794 , \5787 , \5792 , \5793 );
and \U$5452 ( \5795 , \4576 , \406 );
and \U$5453 ( \5796 , \4568 , \404 );
nor \U$5454 ( \5797 , \5795 , \5796 );
xnor \U$5455 ( \5798 , \5797 , \413 );
and \U$5456 ( \5799 , \5050 , \422 );
and \U$5457 ( \5800 , \5045 , \420 );
nor \U$5458 ( \5801 , \5799 , \5800 );
xnor \U$5459 ( \5802 , \5801 , \429 );
and \U$5460 ( \5803 , \5798 , \5802 );
and \U$5461 ( \5804 , \5573 , \441 );
and \U$5462 ( \5805 , \5314 , \439 );
nor \U$5463 ( \5806 , \5804 , \5805 );
xnor \U$5464 ( \5807 , \5806 , \448 );
and \U$5465 ( \5808 , \5802 , \5807 );
and \U$5466 ( \5809 , \5798 , \5807 );
or \U$5467 ( \5810 , \5803 , \5808 , \5809 );
or \U$5468 ( \5811 , \5794 , \5810 );
and \U$5469 ( \5812 , \5777 , \5811 );
and \U$5470 ( \5813 , \5725 , \5811 );
or \U$5471 ( \5814 , \5778 , \5812 , \5813 );
xor \U$5472 ( \5815 , \5498 , \5502 );
xor \U$5473 ( \5816 , \5815 , \5507 );
xor \U$5474 ( \5817 , \5514 , \5518 );
xor \U$5475 ( \5818 , \5817 , \5523 );
and \U$5476 ( \5819 , \5816 , \5818 );
xor \U$5477 ( \5820 , \5479 , \5483 );
xor \U$5478 ( \5821 , \5820 , \5488 );
and \U$5479 ( \5822 , \5818 , \5821 );
and \U$5480 ( \5823 , \5816 , \5821 );
or \U$5481 ( \5824 , \5819 , \5822 , \5823 );
xor \U$5482 ( \5825 , \5531 , \5535 );
xor \U$5483 ( \5826 , \5825 , \5540 );
xor \U$5484 ( \5827 , \5551 , \5555 );
xor \U$5485 ( \5828 , \5827 , \5560 );
and \U$5486 ( \5829 , \5826 , \5828 );
xor \U$5487 ( \5830 , \5567 , \5571 );
xor \U$5488 ( \5831 , \5830 , \5574 );
and \U$5489 ( \5832 , \5828 , \5831 );
and \U$5490 ( \5833 , \5826 , \5831 );
or \U$5491 ( \5834 , \5829 , \5832 , \5833 );
and \U$5492 ( \5835 , \5824 , \5834 );
xor \U$5493 ( \5836 , \5446 , \5450 );
xor \U$5494 ( \5837 , \5836 , \5455 );
xor \U$5495 ( \5838 , \5462 , \5466 );
xor \U$5496 ( \5839 , \5838 , \5471 );
and \U$5497 ( \5840 , \5837 , \5839 );
and \U$5498 ( \5841 , \5834 , \5840 );
and \U$5499 ( \5842 , \5824 , \5840 );
or \U$5500 ( \5843 , \5835 , \5841 , \5842 );
and \U$5501 ( \5844 , \5814 , \5843 );
xor \U$5502 ( \5845 , \5203 , \5207 );
xor \U$5503 ( \5846 , \5845 , \5212 );
xor \U$5504 ( \5847 , \5588 , \5590 );
xor \U$5505 ( \5848 , \5847 , \5593 );
and \U$5506 ( \5849 , \5846 , \5848 );
xor \U$5507 ( \5850 , \5598 , \5600 );
xor \U$5508 ( \5851 , \5850 , \5603 );
and \U$5509 ( \5852 , \5848 , \5851 );
and \U$5510 ( \5853 , \5846 , \5851 );
or \U$5511 ( \5854 , \5849 , \5852 , \5853 );
and \U$5512 ( \5855 , \5843 , \5854 );
and \U$5513 ( \5856 , \5814 , \5854 );
or \U$5514 ( \5857 , \5844 , \5855 , \5856 );
xor \U$5515 ( \5858 , \5458 , \5474 );
xor \U$5516 ( \5859 , \5858 , \5491 );
xor \U$5517 ( \5860 , \5510 , \5526 );
xor \U$5518 ( \5861 , \5860 , \5543 );
and \U$5519 ( \5862 , \5859 , \5861 );
xor \U$5520 ( \5863 , \5563 , \5577 );
xor \U$5521 ( \5864 , \5863 , \5580 );
and \U$5522 ( \5865 , \5861 , \5864 );
and \U$5523 ( \5866 , \5859 , \5864 );
or \U$5524 ( \5867 , \5862 , \5865 , \5866 );
xor \U$5525 ( \5868 , \5215 , \5231 );
xor \U$5526 ( \5869 , \5868 , \5248 );
and \U$5527 ( \5870 , \5867 , \5869 );
xor \U$5528 ( \5871 , \5267 , \5283 );
xor \U$5529 ( \5872 , \5871 , \5300 );
and \U$5530 ( \5873 , \5869 , \5872 );
and \U$5531 ( \5874 , \5867 , \5872 );
or \U$5532 ( \5875 , \5870 , \5873 , \5874 );
and \U$5533 ( \5876 , \5857 , \5875 );
xor \U$5534 ( \5877 , \5494 , \5546 );
xor \U$5535 ( \5878 , \5877 , \5583 );
xor \U$5536 ( \5879 , \5596 , \5606 );
xor \U$5537 ( \5880 , \5879 , \5609 );
and \U$5538 ( \5881 , \5878 , \5880 );
xor \U$5539 ( \5882 , \5615 , \5617 );
xor \U$5540 ( \5883 , \5882 , \5620 );
and \U$5541 ( \5884 , \5880 , \5883 );
and \U$5542 ( \5885 , \5878 , \5883 );
or \U$5543 ( \5886 , \5881 , \5884 , \5885 );
and \U$5544 ( \5887 , \5875 , \5886 );
and \U$5545 ( \5888 , \5857 , \5886 );
or \U$5546 ( \5889 , \5876 , \5887 , \5888 );
xor \U$5547 ( \5890 , \5251 , \5303 );
xor \U$5548 ( \5891 , \5890 , \5339 );
xor \U$5549 ( \5892 , \5586 , \5612 );
xor \U$5550 ( \5893 , \5892 , \5623 );
and \U$5551 ( \5894 , \5891 , \5893 );
xor \U$5552 ( \5895 , \5628 , \5630 );
xor \U$5553 ( \5896 , \5895 , \5633 );
and \U$5554 ( \5897 , \5893 , \5896 );
and \U$5555 ( \5898 , \5891 , \5896 );
or \U$5556 ( \5899 , \5894 , \5897 , \5898 );
and \U$5557 ( \5900 , \5889 , \5899 );
xor \U$5558 ( \5901 , \5644 , \5646 );
xor \U$5559 ( \5902 , \5901 , \5649 );
and \U$5560 ( \5903 , \5899 , \5902 );
and \U$5561 ( \5904 , \5889 , \5902 );
or \U$5562 ( \5905 , \5900 , \5903 , \5904 );
xor \U$5563 ( \5906 , \5382 , \5400 );
xor \U$5564 ( \5907 , \5906 , \5403 );
and \U$5565 ( \5908 , \5905 , \5907 );
xor \U$5566 ( \5909 , \5642 , \5652 );
xor \U$5567 ( \5910 , \5909 , \5655 );
and \U$5568 ( \5911 , \5907 , \5910 );
and \U$5569 ( \5912 , \5905 , \5910 );
or \U$5570 ( \5913 , \5908 , \5911 , \5912 );
xor \U$5571 ( \5914 , \5658 , \5660 );
xor \U$5572 ( \5915 , \5914 , \5662 );
and \U$5573 ( \5916 , \5913 , \5915 );
and \U$5574 ( \5917 , \5671 , \5916 );
xor \U$5575 ( \5918 , \5671 , \5916 );
xor \U$5576 ( \5919 , \5913 , \5915 );
and \U$5577 ( \5920 , \3808 , \357 );
and \U$5578 ( \5921 , \3686 , \355 );
nor \U$5579 ( \5922 , \5920 , \5921 );
xnor \U$5580 ( \5923 , \5922 , \364 );
and \U$5581 ( \5924 , \4069 , \373 );
and \U$5582 ( \5925 , \3813 , \371 );
nor \U$5583 ( \5926 , \5924 , \5925 );
xnor \U$5584 ( \5927 , \5926 , \380 );
and \U$5585 ( \5928 , \5923 , \5927 );
and \U$5586 ( \5929 , \4568 , \391 );
and \U$5587 ( \5930 , \4266 , \389 );
nor \U$5588 ( \5931 , \5929 , \5930 );
xnor \U$5589 ( \5932 , \5931 , \398 );
and \U$5590 ( \5933 , \5927 , \5932 );
and \U$5591 ( \5934 , \5923 , \5932 );
or \U$5592 ( \5935 , \5928 , \5933 , \5934 );
and \U$5593 ( \5936 , \5045 , \406 );
and \U$5594 ( \5937 , \4576 , \404 );
nor \U$5595 ( \5938 , \5936 , \5937 );
xnor \U$5596 ( \5939 , \5938 , \413 );
and \U$5597 ( \5940 , \5314 , \422 );
and \U$5598 ( \5941 , \5050 , \420 );
nor \U$5599 ( \5942 , \5940 , \5941 );
xnor \U$5600 ( \5943 , \5942 , \429 );
and \U$5601 ( \5944 , \5939 , \5943 );
buf \U$5602 ( \5945 , RIbb2c280_111);
and \U$5603 ( \5946 , \5945 , \441 );
and \U$5604 ( \5947 , \5573 , \439 );
nor \U$5605 ( \5948 , \5946 , \5947 );
xnor \U$5606 ( \5949 , \5948 , \448 );
and \U$5607 ( \5950 , \5943 , \5949 );
and \U$5608 ( \5951 , \5939 , \5949 );
or \U$5609 ( \5952 , \5944 , \5950 , \5951 );
and \U$5610 ( \5953 , \5935 , \5952 );
buf \U$5611 ( \5954 , RIbb2c208_112);
and \U$5612 ( \5955 , \5954 , \436 );
buf \U$5613 ( \5956 , \5955 );
and \U$5614 ( \5957 , \5952 , \5956 );
and \U$5615 ( \5958 , \5935 , \5956 );
or \U$5616 ( \5959 , \5953 , \5957 , \5958 );
and \U$5617 ( \5960 , \1839 , \1623 );
and \U$5618 ( \5961 , \1596 , \1621 );
nor \U$5619 ( \5962 , \5960 , \5961 );
xnor \U$5620 ( \5963 , \5962 , \1467 );
and \U$5621 ( \5964 , \2030 , \1351 );
and \U$5622 ( \5965 , \1844 , \1349 );
nor \U$5623 ( \5966 , \5964 , \5965 );
xnor \U$5624 ( \5967 , \5966 , \1238 );
and \U$5625 ( \5968 , \5963 , \5967 );
and \U$5626 ( \5969 , \2438 , \1157 );
and \U$5627 ( \5970 , \2174 , \1155 );
nor \U$5628 ( \5971 , \5969 , \5970 );
xnor \U$5629 ( \5972 , \5971 , \1021 );
and \U$5630 ( \5973 , \5967 , \5972 );
and \U$5631 ( \5974 , \5963 , \5972 );
or \U$5632 ( \5975 , \5968 , \5973 , \5974 );
and \U$5633 ( \5976 , \1176 , \2393 );
and \U$5634 ( \5977 , \1071 , \2391 );
nor \U$5635 ( \5978 , \5976 , \5977 );
xnor \U$5636 ( \5979 , \5978 , \2251 );
and \U$5637 ( \5980 , \1297 , \2097 );
and \U$5638 ( \5981 , \1181 , \2095 );
nor \U$5639 ( \5982 , \5980 , \5981 );
xnor \U$5640 ( \5983 , \5982 , \1960 );
and \U$5641 ( \5984 , \5979 , \5983 );
and \U$5642 ( \5985 , \1588 , \1891 );
and \U$5643 ( \5986 , \1412 , \1889 );
nor \U$5644 ( \5987 , \5985 , \5986 );
xnor \U$5645 ( \5988 , \5987 , \1739 );
and \U$5646 ( \5989 , \5983 , \5988 );
and \U$5647 ( \5990 , \5979 , \5988 );
or \U$5648 ( \5991 , \5984 , \5989 , \5990 );
and \U$5649 ( \5992 , \5975 , \5991 );
and \U$5650 ( \5993 , \2637 , \957 );
and \U$5651 ( \5994 , \2463 , \955 );
nor \U$5652 ( \5995 , \5993 , \5994 );
xnor \U$5653 ( \5996 , \5995 , \879 );
and \U$5654 ( \5997 , \2942 , \793 );
and \U$5655 ( \5998 , \2804 , \791 );
nor \U$5656 ( \5999 , \5997 , \5998 );
xnor \U$5657 ( \6000 , \5999 , \699 );
and \U$5658 ( \6001 , \5996 , \6000 );
and \U$5659 ( \6002 , \3478 , \624 );
and \U$5660 ( \6003 , \3061 , \622 );
nor \U$5661 ( \6004 , \6002 , \6003 );
xnor \U$5662 ( \6005 , \6004 , \349 );
and \U$5663 ( \6006 , \6000 , \6005 );
and \U$5664 ( \6007 , \5996 , \6005 );
or \U$5665 ( \6008 , \6001 , \6006 , \6007 );
and \U$5666 ( \6009 , \5991 , \6008 );
and \U$5667 ( \6010 , \5975 , \6008 );
or \U$5668 ( \6011 , \5992 , \6009 , \6010 );
and \U$5669 ( \6012 , \5959 , \6011 );
and \U$5670 ( \6013 , \408 , \4603 );
and \U$5671 ( \6014 , \385 , \4601 );
nor \U$5672 ( \6015 , \6013 , \6014 );
xnor \U$5673 ( \6016 , \6015 , \4371 );
and \U$5674 ( \6017 , \424 , \4152 );
and \U$5675 ( \6018 , \400 , \4150 );
nor \U$5676 ( \6019 , \6017 , \6018 );
xnor \U$5677 ( \6020 , \6019 , \4009 );
and \U$5678 ( \6021 , \6016 , \6020 );
and \U$5679 ( \6022 , \443 , \3829 );
and \U$5680 ( \6023 , \416 , \3827 );
nor \U$5681 ( \6024 , \6022 , \6023 );
xnor \U$5682 ( \6025 , \6024 , \3583 );
and \U$5683 ( \6026 , \6020 , \6025 );
and \U$5684 ( \6027 , \6016 , \6025 );
or \U$5685 ( \6028 , \6021 , \6026 , \6027 );
xor \U$5686 ( \6029 , \5199 , \5688 );
xor \U$5687 ( \6030 , \5688 , \5689 );
not \U$5688 ( \6031 , \6030 );
and \U$5689 ( \6032 , \6029 , \6031 );
and \U$5690 ( \6033 , \359 , \6032 );
not \U$5691 ( \6034 , \6033 );
xnor \U$5692 ( \6035 , \6034 , \5692 );
and \U$5693 ( \6036 , \375 , \5443 );
and \U$5694 ( \6037 , \351 , \5441 );
nor \U$5695 ( \6038 , \6036 , \6037 );
xnor \U$5696 ( \6039 , \6038 , \5202 );
and \U$5697 ( \6040 , \6035 , \6039 );
and \U$5698 ( \6041 , \393 , \4977 );
and \U$5699 ( \6042 , \367 , \4975 );
nor \U$5700 ( \6043 , \6041 , \6042 );
xnor \U$5701 ( \6044 , \6043 , \4789 );
and \U$5702 ( \6045 , \6039 , \6044 );
and \U$5703 ( \6046 , \6035 , \6044 );
or \U$5704 ( \6047 , \6040 , \6045 , \6046 );
and \U$5705 ( \6048 , \6028 , \6047 );
and \U$5706 ( \6049 , \450 , \3434 );
and \U$5707 ( \6050 , \435 , \3432 );
nor \U$5708 ( \6051 , \6049 , \6050 );
xnor \U$5709 ( \6052 , \6051 , \3247 );
and \U$5710 ( \6053 , \722 , \3121 );
and \U$5711 ( \6054 , \661 , \3119 );
nor \U$5712 ( \6055 , \6053 , \6054 );
xnor \U$5713 ( \6056 , \6055 , \2916 );
and \U$5714 ( \6057 , \6052 , \6056 );
and \U$5715 ( \6058 , \983 , \2715 );
and \U$5716 ( \6059 , \785 , \2713 );
nor \U$5717 ( \6060 , \6058 , \6059 );
xnor \U$5718 ( \6061 , \6060 , \2566 );
and \U$5719 ( \6062 , \6056 , \6061 );
and \U$5720 ( \6063 , \6052 , \6061 );
or \U$5721 ( \6064 , \6057 , \6062 , \6063 );
and \U$5722 ( \6065 , \6047 , \6064 );
and \U$5723 ( \6066 , \6028 , \6064 );
or \U$5724 ( \6067 , \6048 , \6065 , \6066 );
and \U$5725 ( \6068 , \6011 , \6067 );
and \U$5726 ( \6069 , \5959 , \6067 );
or \U$5727 ( \6070 , \6012 , \6068 , \6069 );
xor \U$5728 ( \6071 , \5675 , \5679 );
xor \U$5729 ( \6072 , \6071 , \5684 );
xor \U$5730 ( \6073 , \5693 , \5697 );
xor \U$5731 ( \6074 , \6073 , \5702 );
and \U$5732 ( \6075 , \6072 , \6074 );
xor \U$5733 ( \6076 , \5710 , \5714 );
xor \U$5734 ( \6077 , \6076 , \5719 );
and \U$5735 ( \6078 , \6074 , \6077 );
and \U$5736 ( \6079 , \6072 , \6077 );
or \U$5737 ( \6080 , \6075 , \6078 , \6079 );
xor \U$5738 ( \6081 , \5729 , \5733 );
xor \U$5739 ( \6082 , \6081 , \5738 );
xor \U$5740 ( \6083 , \5745 , \5749 );
xor \U$5741 ( \6084 , \6083 , \5754 );
and \U$5742 ( \6085 , \6082 , \6084 );
xor \U$5743 ( \6086 , \5762 , \5766 );
xor \U$5744 ( \6087 , \6086 , \5771 );
and \U$5745 ( \6088 , \6084 , \6087 );
and \U$5746 ( \6089 , \6082 , \6087 );
or \U$5747 ( \6090 , \6085 , \6088 , \6089 );
and \U$5748 ( \6091 , \6080 , \6090 );
and \U$5749 ( \6092 , \5945 , \436 );
xor \U$5750 ( \6093 , \5782 , \5786 );
xor \U$5751 ( \6094 , \6093 , \5791 );
and \U$5752 ( \6095 , \6092 , \6094 );
xor \U$5753 ( \6096 , \5798 , \5802 );
xor \U$5754 ( \6097 , \6096 , \5807 );
and \U$5755 ( \6098 , \6094 , \6097 );
and \U$5756 ( \6099 , \6092 , \6097 );
or \U$5757 ( \6100 , \6095 , \6098 , \6099 );
and \U$5758 ( \6101 , \6090 , \6100 );
and \U$5759 ( \6102 , \6080 , \6100 );
or \U$5760 ( \6103 , \6091 , \6101 , \6102 );
and \U$5761 ( \6104 , \6070 , \6103 );
xor \U$5762 ( \6105 , \5816 , \5818 );
xor \U$5763 ( \6106 , \6105 , \5821 );
xor \U$5764 ( \6107 , \5826 , \5828 );
xor \U$5765 ( \6108 , \6107 , \5831 );
and \U$5766 ( \6109 , \6106 , \6108 );
xor \U$5767 ( \6110 , \5837 , \5839 );
and \U$5768 ( \6111 , \6108 , \6110 );
and \U$5769 ( \6112 , \6106 , \6110 );
or \U$5770 ( \6113 , \6109 , \6111 , \6112 );
and \U$5771 ( \6114 , \6103 , \6113 );
and \U$5772 ( \6115 , \6070 , \6113 );
or \U$5773 ( \6116 , \6104 , \6114 , \6115 );
xor \U$5774 ( \6117 , \5687 , \5705 );
xor \U$5775 ( \6118 , \6117 , \5722 );
xor \U$5776 ( \6119 , \5741 , \5757 );
xor \U$5777 ( \6120 , \6119 , \5774 );
and \U$5778 ( \6121 , \6118 , \6120 );
xnor \U$5779 ( \6122 , \5794 , \5810 );
and \U$5780 ( \6123 , \6120 , \6122 );
and \U$5781 ( \6124 , \6118 , \6122 );
or \U$5782 ( \6125 , \6121 , \6123 , \6124 );
xor \U$5783 ( \6126 , \5846 , \5848 );
xor \U$5784 ( \6127 , \6126 , \5851 );
and \U$5785 ( \6128 , \6125 , \6127 );
xor \U$5786 ( \6129 , \5859 , \5861 );
xor \U$5787 ( \6130 , \6129 , \5864 );
and \U$5788 ( \6131 , \6127 , \6130 );
and \U$5789 ( \6132 , \6125 , \6130 );
or \U$5790 ( \6133 , \6128 , \6131 , \6132 );
and \U$5791 ( \6134 , \6116 , \6133 );
xor \U$5792 ( \6135 , \5725 , \5777 );
xor \U$5793 ( \6136 , \6135 , \5811 );
xor \U$5794 ( \6137 , \5824 , \5834 );
xor \U$5795 ( \6138 , \6137 , \5840 );
and \U$5796 ( \6139 , \6136 , \6138 );
and \U$5797 ( \6140 , \6133 , \6139 );
and \U$5798 ( \6141 , \6116 , \6139 );
or \U$5799 ( \6142 , \6134 , \6140 , \6141 );
xor \U$5800 ( \6143 , \5814 , \5843 );
xor \U$5801 ( \6144 , \6143 , \5854 );
xor \U$5802 ( \6145 , \5867 , \5869 );
xor \U$5803 ( \6146 , \6145 , \5872 );
and \U$5804 ( \6147 , \6144 , \6146 );
xor \U$5805 ( \6148 , \5878 , \5880 );
xor \U$5806 ( \6149 , \6148 , \5883 );
and \U$5807 ( \6150 , \6146 , \6149 );
and \U$5808 ( \6151 , \6144 , \6149 );
or \U$5809 ( \6152 , \6147 , \6150 , \6151 );
and \U$5810 ( \6153 , \6142 , \6152 );
xor \U$5811 ( \6154 , \5891 , \5893 );
xor \U$5812 ( \6155 , \6154 , \5896 );
and \U$5813 ( \6156 , \6152 , \6155 );
and \U$5814 ( \6157 , \6142 , \6155 );
or \U$5815 ( \6158 , \6153 , \6156 , \6157 );
xor \U$5816 ( \6159 , \5626 , \5636 );
xor \U$5817 ( \6160 , \6159 , \5639 );
and \U$5818 ( \6161 , \6158 , \6160 );
xor \U$5819 ( \6162 , \5889 , \5899 );
xor \U$5820 ( \6163 , \6162 , \5902 );
and \U$5821 ( \6164 , \6160 , \6163 );
and \U$5822 ( \6165 , \6158 , \6163 );
or \U$5823 ( \6166 , \6161 , \6164 , \6165 );
xor \U$5824 ( \6167 , \5905 , \5907 );
xor \U$5825 ( \6168 , \6167 , \5910 );
and \U$5826 ( \6169 , \6166 , \6168 );
and \U$5827 ( \6170 , \5919 , \6169 );
xor \U$5828 ( \6171 , \5919 , \6169 );
xor \U$5829 ( \6172 , \6166 , \6168 );
xor \U$5830 ( \6173 , \5963 , \5967 );
xor \U$5831 ( \6174 , \6173 , \5972 );
xor \U$5832 ( \6175 , \5979 , \5983 );
xor \U$5833 ( \6176 , \6175 , \5988 );
and \U$5834 ( \6177 , \6174 , \6176 );
xor \U$5835 ( \6178 , \5996 , \6000 );
xor \U$5836 ( \6179 , \6178 , \6005 );
and \U$5837 ( \6180 , \6176 , \6179 );
and \U$5838 ( \6181 , \6174 , \6179 );
or \U$5839 ( \6182 , \6177 , \6180 , \6181 );
xor \U$5840 ( \6183 , \6016 , \6020 );
xor \U$5841 ( \6184 , \6183 , \6025 );
xor \U$5842 ( \6185 , \6035 , \6039 );
xor \U$5843 ( \6186 , \6185 , \6044 );
and \U$5844 ( \6187 , \6184 , \6186 );
xor \U$5845 ( \6188 , \6052 , \6056 );
xor \U$5846 ( \6189 , \6188 , \6061 );
and \U$5847 ( \6190 , \6186 , \6189 );
and \U$5848 ( \6191 , \6184 , \6189 );
or \U$5849 ( \6192 , \6187 , \6190 , \6191 );
and \U$5850 ( \6193 , \6182 , \6192 );
xor \U$5851 ( \6194 , \5923 , \5927 );
xor \U$5852 ( \6195 , \6194 , \5932 );
xor \U$5853 ( \6196 , \5939 , \5943 );
xor \U$5854 ( \6197 , \6196 , \5949 );
and \U$5855 ( \6198 , \6195 , \6197 );
not \U$5856 ( \6199 , \5955 );
and \U$5857 ( \6200 , \6197 , \6199 );
and \U$5858 ( \6201 , \6195 , \6199 );
or \U$5859 ( \6202 , \6198 , \6200 , \6201 );
and \U$5860 ( \6203 , \6192 , \6202 );
and \U$5861 ( \6204 , \6182 , \6202 );
or \U$5862 ( \6205 , \6193 , \6203 , \6204 );
and \U$5863 ( \6206 , \385 , \4977 );
and \U$5864 ( \6207 , \393 , \4975 );
nor \U$5865 ( \6208 , \6206 , \6207 );
xnor \U$5866 ( \6209 , \6208 , \4789 );
and \U$5867 ( \6210 , \400 , \4603 );
and \U$5868 ( \6211 , \408 , \4601 );
nor \U$5869 ( \6212 , \6210 , \6211 );
xnor \U$5870 ( \6213 , \6212 , \4371 );
and \U$5871 ( \6214 , \6209 , \6213 );
and \U$5872 ( \6215 , \416 , \4152 );
and \U$5873 ( \6216 , \424 , \4150 );
nor \U$5874 ( \6217 , \6215 , \6216 );
xnor \U$5875 ( \6218 , \6217 , \4009 );
and \U$5876 ( \6219 , \6213 , \6218 );
and \U$5877 ( \6220 , \6209 , \6218 );
or \U$5878 ( \6221 , \6214 , \6219 , \6220 );
buf \U$5879 ( \6222 , RIbb2df18_50);
buf \U$5880 ( \6223 , RIbb2dea0_51);
and \U$5881 ( \6224 , \6222 , \6223 );
not \U$5882 ( \6225 , \6224 );
and \U$5883 ( \6226 , \5689 , \6225 );
not \U$5884 ( \6227 , \6226 );
and \U$5885 ( \6228 , \351 , \6032 );
and \U$5886 ( \6229 , \359 , \6030 );
nor \U$5887 ( \6230 , \6228 , \6229 );
xnor \U$5888 ( \6231 , \6230 , \5692 );
and \U$5889 ( \6232 , \6227 , \6231 );
and \U$5890 ( \6233 , \367 , \5443 );
and \U$5891 ( \6234 , \375 , \5441 );
nor \U$5892 ( \6235 , \6233 , \6234 );
xnor \U$5893 ( \6236 , \6235 , \5202 );
and \U$5894 ( \6237 , \6231 , \6236 );
and \U$5895 ( \6238 , \6227 , \6236 );
or \U$5896 ( \6239 , \6232 , \6237 , \6238 );
and \U$5897 ( \6240 , \6221 , \6239 );
and \U$5898 ( \6241 , \435 , \3829 );
and \U$5899 ( \6242 , \443 , \3827 );
nor \U$5900 ( \6243 , \6241 , \6242 );
xnor \U$5901 ( \6244 , \6243 , \3583 );
and \U$5902 ( \6245 , \661 , \3434 );
and \U$5903 ( \6246 , \450 , \3432 );
nor \U$5904 ( \6247 , \6245 , \6246 );
xnor \U$5905 ( \6248 , \6247 , \3247 );
and \U$5906 ( \6249 , \6244 , \6248 );
and \U$5907 ( \6250 , \785 , \3121 );
and \U$5908 ( \6251 , \722 , \3119 );
nor \U$5909 ( \6252 , \6250 , \6251 );
xnor \U$5910 ( \6253 , \6252 , \2916 );
and \U$5911 ( \6254 , \6248 , \6253 );
and \U$5912 ( \6255 , \6244 , \6253 );
or \U$5913 ( \6256 , \6249 , \6254 , \6255 );
and \U$5914 ( \6257 , \6239 , \6256 );
and \U$5915 ( \6258 , \6221 , \6256 );
or \U$5916 ( \6259 , \6240 , \6257 , \6258 );
and \U$5917 ( \6260 , \3686 , \624 );
and \U$5918 ( \6261 , \3478 , \622 );
nor \U$5919 ( \6262 , \6260 , \6261 );
xnor \U$5920 ( \6263 , \6262 , \349 );
and \U$5921 ( \6264 , \3813 , \357 );
and \U$5922 ( \6265 , \3808 , \355 );
nor \U$5923 ( \6266 , \6264 , \6265 );
xnor \U$5924 ( \6267 , \6266 , \364 );
and \U$5925 ( \6268 , \6263 , \6267 );
and \U$5926 ( \6269 , \4266 , \373 );
and \U$5927 ( \6270 , \4069 , \371 );
nor \U$5928 ( \6271 , \6269 , \6270 );
xnor \U$5929 ( \6272 , \6271 , \380 );
and \U$5930 ( \6273 , \6267 , \6272 );
and \U$5931 ( \6274 , \6263 , \6272 );
or \U$5932 ( \6275 , \6268 , \6273 , \6274 );
and \U$5933 ( \6276 , \4576 , \391 );
and \U$5934 ( \6277 , \4568 , \389 );
nor \U$5935 ( \6278 , \6276 , \6277 );
xnor \U$5936 ( \6279 , \6278 , \398 );
and \U$5937 ( \6280 , \5050 , \406 );
and \U$5938 ( \6281 , \5045 , \404 );
nor \U$5939 ( \6282 , \6280 , \6281 );
xnor \U$5940 ( \6283 , \6282 , \413 );
and \U$5941 ( \6284 , \6279 , \6283 );
and \U$5942 ( \6285 , \5573 , \422 );
and \U$5943 ( \6286 , \5314 , \420 );
nor \U$5944 ( \6287 , \6285 , \6286 );
xnor \U$5945 ( \6288 , \6287 , \429 );
and \U$5946 ( \6289 , \6283 , \6288 );
and \U$5947 ( \6290 , \6279 , \6288 );
or \U$5948 ( \6291 , \6284 , \6289 , \6290 );
and \U$5949 ( \6292 , \6275 , \6291 );
and \U$5950 ( \6293 , \5954 , \441 );
and \U$5951 ( \6294 , \5945 , \439 );
nor \U$5952 ( \6295 , \6293 , \6294 );
xnor \U$5953 ( \6296 , \6295 , \448 );
buf \U$5954 ( \6297 , RIbb2c190_113);
and \U$5955 ( \6298 , \6297 , \436 );
and \U$5956 ( \6299 , \6296 , \6298 );
and \U$5957 ( \6300 , \6291 , \6299 );
and \U$5958 ( \6301 , \6275 , \6299 );
or \U$5959 ( \6302 , \6292 , \6300 , \6301 );
and \U$5960 ( \6303 , \6259 , \6302 );
and \U$5961 ( \6304 , \1071 , \2715 );
and \U$5962 ( \6305 , \983 , \2713 );
nor \U$5963 ( \6306 , \6304 , \6305 );
xnor \U$5964 ( \6307 , \6306 , \2566 );
and \U$5965 ( \6308 , \1181 , \2393 );
and \U$5966 ( \6309 , \1176 , \2391 );
nor \U$5967 ( \6310 , \6308 , \6309 );
xnor \U$5968 ( \6311 , \6310 , \2251 );
and \U$5969 ( \6312 , \6307 , \6311 );
and \U$5970 ( \6313 , \1412 , \2097 );
and \U$5971 ( \6314 , \1297 , \2095 );
nor \U$5972 ( \6315 , \6313 , \6314 );
xnor \U$5973 ( \6316 , \6315 , \1960 );
and \U$5974 ( \6317 , \6311 , \6316 );
and \U$5975 ( \6318 , \6307 , \6316 );
or \U$5976 ( \6319 , \6312 , \6317 , \6318 );
and \U$5977 ( \6320 , \1596 , \1891 );
and \U$5978 ( \6321 , \1588 , \1889 );
nor \U$5979 ( \6322 , \6320 , \6321 );
xnor \U$5980 ( \6323 , \6322 , \1739 );
and \U$5981 ( \6324 , \1844 , \1623 );
and \U$5982 ( \6325 , \1839 , \1621 );
nor \U$5983 ( \6326 , \6324 , \6325 );
xnor \U$5984 ( \6327 , \6326 , \1467 );
and \U$5985 ( \6328 , \6323 , \6327 );
and \U$5986 ( \6329 , \2174 , \1351 );
and \U$5987 ( \6330 , \2030 , \1349 );
nor \U$5988 ( \6331 , \6329 , \6330 );
xnor \U$5989 ( \6332 , \6331 , \1238 );
and \U$5990 ( \6333 , \6327 , \6332 );
and \U$5991 ( \6334 , \6323 , \6332 );
or \U$5992 ( \6335 , \6328 , \6333 , \6334 );
and \U$5993 ( \6336 , \6319 , \6335 );
and \U$5994 ( \6337 , \2463 , \1157 );
and \U$5995 ( \6338 , \2438 , \1155 );
nor \U$5996 ( \6339 , \6337 , \6338 );
xnor \U$5997 ( \6340 , \6339 , \1021 );
and \U$5998 ( \6341 , \2804 , \957 );
and \U$5999 ( \6342 , \2637 , \955 );
nor \U$6000 ( \6343 , \6341 , \6342 );
xnor \U$6001 ( \6344 , \6343 , \879 );
and \U$6002 ( \6345 , \6340 , \6344 );
and \U$6003 ( \6346 , \3061 , \793 );
and \U$6004 ( \6347 , \2942 , \791 );
nor \U$6005 ( \6348 , \6346 , \6347 );
xnor \U$6006 ( \6349 , \6348 , \699 );
and \U$6007 ( \6350 , \6344 , \6349 );
and \U$6008 ( \6351 , \6340 , \6349 );
or \U$6009 ( \6352 , \6345 , \6350 , \6351 );
and \U$6010 ( \6353 , \6335 , \6352 );
and \U$6011 ( \6354 , \6319 , \6352 );
or \U$6012 ( \6355 , \6336 , \6353 , \6354 );
and \U$6013 ( \6356 , \6302 , \6355 );
and \U$6014 ( \6357 , \6259 , \6355 );
or \U$6015 ( \6358 , \6303 , \6356 , \6357 );
and \U$6016 ( \6359 , \6205 , \6358 );
xor \U$6017 ( \6360 , \6072 , \6074 );
xor \U$6018 ( \6361 , \6360 , \6077 );
xor \U$6019 ( \6362 , \6082 , \6084 );
xor \U$6020 ( \6363 , \6362 , \6087 );
and \U$6021 ( \6364 , \6361 , \6363 );
xor \U$6022 ( \6365 , \6092 , \6094 );
xor \U$6023 ( \6366 , \6365 , \6097 );
and \U$6024 ( \6367 , \6363 , \6366 );
and \U$6025 ( \6368 , \6361 , \6366 );
or \U$6026 ( \6369 , \6364 , \6367 , \6368 );
and \U$6027 ( \6370 , \6358 , \6369 );
and \U$6028 ( \6371 , \6205 , \6369 );
or \U$6029 ( \6372 , \6359 , \6370 , \6371 );
xor \U$6030 ( \6373 , \5935 , \5952 );
xor \U$6031 ( \6374 , \6373 , \5956 );
xor \U$6032 ( \6375 , \5975 , \5991 );
xor \U$6033 ( \6376 , \6375 , \6008 );
and \U$6034 ( \6377 , \6374 , \6376 );
xor \U$6035 ( \6378 , \6028 , \6047 );
xor \U$6036 ( \6379 , \6378 , \6064 );
and \U$6037 ( \6380 , \6376 , \6379 );
and \U$6038 ( \6381 , \6374 , \6379 );
or \U$6039 ( \6382 , \6377 , \6380 , \6381 );
xor \U$6040 ( \6383 , \6118 , \6120 );
xor \U$6041 ( \6384 , \6383 , \6122 );
and \U$6042 ( \6385 , \6382 , \6384 );
xor \U$6043 ( \6386 , \6106 , \6108 );
xor \U$6044 ( \6387 , \6386 , \6110 );
and \U$6045 ( \6388 , \6384 , \6387 );
and \U$6046 ( \6389 , \6382 , \6387 );
or \U$6047 ( \6390 , \6385 , \6388 , \6389 );
and \U$6048 ( \6391 , \6372 , \6390 );
xor \U$6049 ( \6392 , \5959 , \6011 );
xor \U$6050 ( \6393 , \6392 , \6067 );
xor \U$6051 ( \6394 , \6080 , \6090 );
xor \U$6052 ( \6395 , \6394 , \6100 );
and \U$6053 ( \6396 , \6393 , \6395 );
and \U$6054 ( \6397 , \6390 , \6396 );
and \U$6055 ( \6398 , \6372 , \6396 );
or \U$6056 ( \6399 , \6391 , \6397 , \6398 );
xor \U$6057 ( \6400 , \6070 , \6103 );
xor \U$6058 ( \6401 , \6400 , \6113 );
xor \U$6059 ( \6402 , \6125 , \6127 );
xor \U$6060 ( \6403 , \6402 , \6130 );
and \U$6061 ( \6404 , \6401 , \6403 );
xor \U$6062 ( \6405 , \6136 , \6138 );
and \U$6063 ( \6406 , \6403 , \6405 );
and \U$6064 ( \6407 , \6401 , \6405 );
or \U$6065 ( \6408 , \6404 , \6406 , \6407 );
and \U$6066 ( \6409 , \6399 , \6408 );
xor \U$6067 ( \6410 , \6144 , \6146 );
xor \U$6068 ( \6411 , \6410 , \6149 );
and \U$6069 ( \6412 , \6408 , \6411 );
and \U$6070 ( \6413 , \6399 , \6411 );
or \U$6071 ( \6414 , \6409 , \6412 , \6413 );
xor \U$6072 ( \6415 , \5857 , \5875 );
xor \U$6073 ( \6416 , \6415 , \5886 );
and \U$6074 ( \6417 , \6414 , \6416 );
xor \U$6075 ( \6418 , \6142 , \6152 );
xor \U$6076 ( \6419 , \6418 , \6155 );
and \U$6077 ( \6420 , \6416 , \6419 );
and \U$6078 ( \6421 , \6414 , \6419 );
or \U$6079 ( \6422 , \6417 , \6420 , \6421 );
xor \U$6080 ( \6423 , \6158 , \6160 );
xor \U$6081 ( \6424 , \6423 , \6163 );
and \U$6082 ( \6425 , \6422 , \6424 );
and \U$6083 ( \6426 , \6172 , \6425 );
xor \U$6084 ( \6427 , \6172 , \6425 );
xor \U$6085 ( \6428 , \6422 , \6424 );
xor \U$6086 ( \6429 , \6307 , \6311 );
xor \U$6087 ( \6430 , \6429 , \6316 );
xor \U$6088 ( \6431 , \6323 , \6327 );
xor \U$6089 ( \6432 , \6431 , \6332 );
and \U$6090 ( \6433 , \6430 , \6432 );
xor \U$6091 ( \6434 , \6340 , \6344 );
xor \U$6092 ( \6435 , \6434 , \6349 );
and \U$6093 ( \6436 , \6432 , \6435 );
and \U$6094 ( \6437 , \6430 , \6435 );
or \U$6095 ( \6438 , \6433 , \6436 , \6437 );
xor \U$6096 ( \6439 , \6209 , \6213 );
xor \U$6097 ( \6440 , \6439 , \6218 );
xor \U$6098 ( \6441 , \6227 , \6231 );
xor \U$6099 ( \6442 , \6441 , \6236 );
and \U$6100 ( \6443 , \6440 , \6442 );
xor \U$6101 ( \6444 , \6244 , \6248 );
xor \U$6102 ( \6445 , \6444 , \6253 );
and \U$6103 ( \6446 , \6442 , \6445 );
and \U$6104 ( \6447 , \6440 , \6445 );
or \U$6105 ( \6448 , \6443 , \6446 , \6447 );
and \U$6106 ( \6449 , \6438 , \6448 );
xor \U$6107 ( \6450 , \6263 , \6267 );
xor \U$6108 ( \6451 , \6450 , \6272 );
xor \U$6109 ( \6452 , \6279 , \6283 );
xor \U$6110 ( \6453 , \6452 , \6288 );
and \U$6111 ( \6454 , \6451 , \6453 );
xor \U$6112 ( \6455 , \6296 , \6298 );
and \U$6113 ( \6456 , \6453 , \6455 );
and \U$6114 ( \6457 , \6451 , \6455 );
or \U$6115 ( \6458 , \6454 , \6456 , \6457 );
and \U$6116 ( \6459 , \6448 , \6458 );
and \U$6117 ( \6460 , \6438 , \6458 );
or \U$6118 ( \6461 , \6449 , \6459 , \6460 );
and \U$6119 ( \6462 , \3808 , \624 );
and \U$6120 ( \6463 , \3686 , \622 );
nor \U$6121 ( \6464 , \6462 , \6463 );
xnor \U$6122 ( \6465 , \6464 , \349 );
and \U$6123 ( \6466 , \4069 , \357 );
and \U$6124 ( \6467 , \3813 , \355 );
nor \U$6125 ( \6468 , \6466 , \6467 );
xnor \U$6126 ( \6469 , \6468 , \364 );
and \U$6127 ( \6470 , \6465 , \6469 );
and \U$6128 ( \6471 , \4568 , \373 );
and \U$6129 ( \6472 , \4266 , \371 );
nor \U$6130 ( \6473 , \6471 , \6472 );
xnor \U$6131 ( \6474 , \6473 , \380 );
and \U$6132 ( \6475 , \6469 , \6474 );
and \U$6133 ( \6476 , \6465 , \6474 );
or \U$6134 ( \6477 , \6470 , \6475 , \6476 );
and \U$6135 ( \6478 , \5045 , \391 );
and \U$6136 ( \6479 , \4576 , \389 );
nor \U$6137 ( \6480 , \6478 , \6479 );
xnor \U$6138 ( \6481 , \6480 , \398 );
and \U$6139 ( \6482 , \5314 , \406 );
and \U$6140 ( \6483 , \5050 , \404 );
nor \U$6141 ( \6484 , \6482 , \6483 );
xnor \U$6142 ( \6485 , \6484 , \413 );
and \U$6143 ( \6486 , \6481 , \6485 );
and \U$6144 ( \6487 , \5945 , \422 );
and \U$6145 ( \6488 , \5573 , \420 );
nor \U$6146 ( \6489 , \6487 , \6488 );
xnor \U$6147 ( \6490 , \6489 , \429 );
and \U$6148 ( \6491 , \6485 , \6490 );
and \U$6149 ( \6492 , \6481 , \6490 );
or \U$6150 ( \6493 , \6486 , \6491 , \6492 );
and \U$6151 ( \6494 , \6477 , \6493 );
and \U$6152 ( \6495 , \6297 , \441 );
and \U$6153 ( \6496 , \5954 , \439 );
nor \U$6154 ( \6497 , \6495 , \6496 );
xnor \U$6155 ( \6498 , \6497 , \448 );
buf \U$6156 ( \6499 , RIbb2c118_114);
and \U$6157 ( \6500 , \6499 , \436 );
or \U$6158 ( \6501 , \6498 , \6500 );
and \U$6159 ( \6502 , \6493 , \6501 );
and \U$6160 ( \6503 , \6477 , \6501 );
or \U$6161 ( \6504 , \6494 , \6502 , \6503 );
and \U$6162 ( \6505 , \450 , \3829 );
and \U$6163 ( \6506 , \435 , \3827 );
nor \U$6164 ( \6507 , \6505 , \6506 );
xnor \U$6165 ( \6508 , \6507 , \3583 );
and \U$6166 ( \6509 , \722 , \3434 );
and \U$6167 ( \6510 , \661 , \3432 );
nor \U$6168 ( \6511 , \6509 , \6510 );
xnor \U$6169 ( \6512 , \6511 , \3247 );
and \U$6170 ( \6513 , \6508 , \6512 );
and \U$6171 ( \6514 , \983 , \3121 );
and \U$6172 ( \6515 , \785 , \3119 );
nor \U$6173 ( \6516 , \6514 , \6515 );
xnor \U$6174 ( \6517 , \6516 , \2916 );
and \U$6175 ( \6518 , \6512 , \6517 );
and \U$6176 ( \6519 , \6508 , \6517 );
or \U$6177 ( \6520 , \6513 , \6518 , \6519 );
and \U$6178 ( \6521 , \408 , \4977 );
and \U$6179 ( \6522 , \385 , \4975 );
nor \U$6180 ( \6523 , \6521 , \6522 );
xnor \U$6181 ( \6524 , \6523 , \4789 );
and \U$6182 ( \6525 , \424 , \4603 );
and \U$6183 ( \6526 , \400 , \4601 );
nor \U$6184 ( \6527 , \6525 , \6526 );
xnor \U$6185 ( \6528 , \6527 , \4371 );
and \U$6186 ( \6529 , \6524 , \6528 );
and \U$6187 ( \6530 , \443 , \4152 );
and \U$6188 ( \6531 , \416 , \4150 );
nor \U$6189 ( \6532 , \6530 , \6531 );
xnor \U$6190 ( \6533 , \6532 , \4009 );
and \U$6191 ( \6534 , \6528 , \6533 );
and \U$6192 ( \6535 , \6524 , \6533 );
or \U$6193 ( \6536 , \6529 , \6534 , \6535 );
and \U$6194 ( \6537 , \6520 , \6536 );
xor \U$6195 ( \6538 , \5689 , \6222 );
xor \U$6196 ( \6539 , \6222 , \6223 );
not \U$6197 ( \6540 , \6539 );
and \U$6198 ( \6541 , \6538 , \6540 );
and \U$6199 ( \6542 , \359 , \6541 );
not \U$6200 ( \6543 , \6542 );
xnor \U$6201 ( \6544 , \6543 , \6226 );
and \U$6202 ( \6545 , \375 , \6032 );
and \U$6203 ( \6546 , \351 , \6030 );
nor \U$6204 ( \6547 , \6545 , \6546 );
xnor \U$6205 ( \6548 , \6547 , \5692 );
and \U$6206 ( \6549 , \6544 , \6548 );
and \U$6207 ( \6550 , \393 , \5443 );
and \U$6208 ( \6551 , \367 , \5441 );
nor \U$6209 ( \6552 , \6550 , \6551 );
xnor \U$6210 ( \6553 , \6552 , \5202 );
and \U$6211 ( \6554 , \6548 , \6553 );
and \U$6212 ( \6555 , \6544 , \6553 );
or \U$6213 ( \6556 , \6549 , \6554 , \6555 );
and \U$6214 ( \6557 , \6536 , \6556 );
and \U$6215 ( \6558 , \6520 , \6556 );
or \U$6216 ( \6559 , \6537 , \6557 , \6558 );
and \U$6217 ( \6560 , \6504 , \6559 );
and \U$6218 ( \6561 , \1839 , \1891 );
and \U$6219 ( \6562 , \1596 , \1889 );
nor \U$6220 ( \6563 , \6561 , \6562 );
xnor \U$6221 ( \6564 , \6563 , \1739 );
and \U$6222 ( \6565 , \2030 , \1623 );
and \U$6223 ( \6566 , \1844 , \1621 );
nor \U$6224 ( \6567 , \6565 , \6566 );
xnor \U$6225 ( \6568 , \6567 , \1467 );
and \U$6226 ( \6569 , \6564 , \6568 );
and \U$6227 ( \6570 , \2438 , \1351 );
and \U$6228 ( \6571 , \2174 , \1349 );
nor \U$6229 ( \6572 , \6570 , \6571 );
xnor \U$6230 ( \6573 , \6572 , \1238 );
and \U$6231 ( \6574 , \6568 , \6573 );
and \U$6232 ( \6575 , \6564 , \6573 );
or \U$6233 ( \6576 , \6569 , \6574 , \6575 );
and \U$6234 ( \6577 , \2637 , \1157 );
and \U$6235 ( \6578 , \2463 , \1155 );
nor \U$6236 ( \6579 , \6577 , \6578 );
xnor \U$6237 ( \6580 , \6579 , \1021 );
and \U$6238 ( \6581 , \2942 , \957 );
and \U$6239 ( \6582 , \2804 , \955 );
nor \U$6240 ( \6583 , \6581 , \6582 );
xnor \U$6241 ( \6584 , \6583 , \879 );
and \U$6242 ( \6585 , \6580 , \6584 );
and \U$6243 ( \6586 , \3478 , \793 );
and \U$6244 ( \6587 , \3061 , \791 );
nor \U$6245 ( \6588 , \6586 , \6587 );
xnor \U$6246 ( \6589 , \6588 , \699 );
and \U$6247 ( \6590 , \6584 , \6589 );
and \U$6248 ( \6591 , \6580 , \6589 );
or \U$6249 ( \6592 , \6585 , \6590 , \6591 );
and \U$6250 ( \6593 , \6576 , \6592 );
and \U$6251 ( \6594 , \1176 , \2715 );
and \U$6252 ( \6595 , \1071 , \2713 );
nor \U$6253 ( \6596 , \6594 , \6595 );
xnor \U$6254 ( \6597 , \6596 , \2566 );
and \U$6255 ( \6598 , \1297 , \2393 );
and \U$6256 ( \6599 , \1181 , \2391 );
nor \U$6257 ( \6600 , \6598 , \6599 );
xnor \U$6258 ( \6601 , \6600 , \2251 );
and \U$6259 ( \6602 , \6597 , \6601 );
and \U$6260 ( \6603 , \1588 , \2097 );
and \U$6261 ( \6604 , \1412 , \2095 );
nor \U$6262 ( \6605 , \6603 , \6604 );
xnor \U$6263 ( \6606 , \6605 , \1960 );
and \U$6264 ( \6607 , \6601 , \6606 );
and \U$6265 ( \6608 , \6597 , \6606 );
or \U$6266 ( \6609 , \6602 , \6607 , \6608 );
and \U$6267 ( \6610 , \6592 , \6609 );
and \U$6268 ( \6611 , \6576 , \6609 );
or \U$6269 ( \6612 , \6593 , \6610 , \6611 );
and \U$6270 ( \6613 , \6559 , \6612 );
and \U$6271 ( \6614 , \6504 , \6612 );
or \U$6272 ( \6615 , \6560 , \6613 , \6614 );
and \U$6273 ( \6616 , \6461 , \6615 );
xor \U$6274 ( \6617 , \6174 , \6176 );
xor \U$6275 ( \6618 , \6617 , \6179 );
xor \U$6276 ( \6619 , \6184 , \6186 );
xor \U$6277 ( \6620 , \6619 , \6189 );
and \U$6278 ( \6621 , \6618 , \6620 );
xor \U$6279 ( \6622 , \6195 , \6197 );
xor \U$6280 ( \6623 , \6622 , \6199 );
and \U$6281 ( \6624 , \6620 , \6623 );
and \U$6282 ( \6625 , \6618 , \6623 );
or \U$6283 ( \6626 , \6621 , \6624 , \6625 );
and \U$6284 ( \6627 , \6615 , \6626 );
and \U$6285 ( \6628 , \6461 , \6626 );
or \U$6286 ( \6629 , \6616 , \6627 , \6628 );
xor \U$6287 ( \6630 , \6221 , \6239 );
xor \U$6288 ( \6631 , \6630 , \6256 );
xor \U$6289 ( \6632 , \6275 , \6291 );
xor \U$6290 ( \6633 , \6632 , \6299 );
and \U$6291 ( \6634 , \6631 , \6633 );
xor \U$6292 ( \6635 , \6319 , \6335 );
xor \U$6293 ( \6636 , \6635 , \6352 );
and \U$6294 ( \6637 , \6633 , \6636 );
and \U$6295 ( \6638 , \6631 , \6636 );
or \U$6296 ( \6639 , \6634 , \6637 , \6638 );
xor \U$6297 ( \6640 , \6374 , \6376 );
xor \U$6298 ( \6641 , \6640 , \6379 );
and \U$6299 ( \6642 , \6639 , \6641 );
xor \U$6300 ( \6643 , \6361 , \6363 );
xor \U$6301 ( \6644 , \6643 , \6366 );
and \U$6302 ( \6645 , \6641 , \6644 );
and \U$6303 ( \6646 , \6639 , \6644 );
or \U$6304 ( \6647 , \6642 , \6645 , \6646 );
and \U$6305 ( \6648 , \6629 , \6647 );
xor \U$6306 ( \6649 , \6182 , \6192 );
xor \U$6307 ( \6650 , \6649 , \6202 );
xor \U$6308 ( \6651 , \6259 , \6302 );
xor \U$6309 ( \6652 , \6651 , \6355 );
and \U$6310 ( \6653 , \6650 , \6652 );
and \U$6311 ( \6654 , \6647 , \6653 );
and \U$6312 ( \6655 , \6629 , \6653 );
or \U$6313 ( \6656 , \6648 , \6654 , \6655 );
xor \U$6314 ( \6657 , \6205 , \6358 );
xor \U$6315 ( \6658 , \6657 , \6369 );
xor \U$6316 ( \6659 , \6382 , \6384 );
xor \U$6317 ( \6660 , \6659 , \6387 );
and \U$6318 ( \6661 , \6658 , \6660 );
xor \U$6319 ( \6662 , \6393 , \6395 );
and \U$6320 ( \6663 , \6660 , \6662 );
and \U$6321 ( \6664 , \6658 , \6662 );
or \U$6322 ( \6665 , \6661 , \6663 , \6664 );
and \U$6323 ( \6666 , \6656 , \6665 );
xor \U$6324 ( \6667 , \6401 , \6403 );
xor \U$6325 ( \6668 , \6667 , \6405 );
and \U$6326 ( \6669 , \6665 , \6668 );
and \U$6327 ( \6670 , \6656 , \6668 );
or \U$6328 ( \6671 , \6666 , \6669 , \6670 );
xor \U$6329 ( \6672 , \6116 , \6133 );
xor \U$6330 ( \6673 , \6672 , \6139 );
and \U$6331 ( \6674 , \6671 , \6673 );
xor \U$6332 ( \6675 , \6399 , \6408 );
xor \U$6333 ( \6676 , \6675 , \6411 );
and \U$6334 ( \6677 , \6673 , \6676 );
and \U$6335 ( \6678 , \6671 , \6676 );
or \U$6336 ( \6679 , \6674 , \6677 , \6678 );
xor \U$6337 ( \6680 , \6414 , \6416 );
xor \U$6338 ( \6681 , \6680 , \6419 );
and \U$6339 ( \6682 , \6679 , \6681 );
and \U$6340 ( \6683 , \6428 , \6682 );
xor \U$6341 ( \6684 , \6428 , \6682 );
xor \U$6342 ( \6685 , \6679 , \6681 );
and \U$6343 ( \6686 , \1071 , \3121 );
and \U$6344 ( \6687 , \983 , \3119 );
nor \U$6345 ( \6688 , \6686 , \6687 );
xnor \U$6346 ( \6689 , \6688 , \2916 );
and \U$6347 ( \6690 , \1181 , \2715 );
and \U$6348 ( \6691 , \1176 , \2713 );
nor \U$6349 ( \6692 , \6690 , \6691 );
xnor \U$6350 ( \6693 , \6692 , \2566 );
and \U$6351 ( \6694 , \6689 , \6693 );
and \U$6352 ( \6695 , \1412 , \2393 );
and \U$6353 ( \6696 , \1297 , \2391 );
nor \U$6354 ( \6697 , \6695 , \6696 );
xnor \U$6355 ( \6698 , \6697 , \2251 );
and \U$6356 ( \6699 , \6693 , \6698 );
and \U$6357 ( \6700 , \6689 , \6698 );
or \U$6358 ( \6701 , \6694 , \6699 , \6700 );
and \U$6359 ( \6702 , \1596 , \2097 );
and \U$6360 ( \6703 , \1588 , \2095 );
nor \U$6361 ( \6704 , \6702 , \6703 );
xnor \U$6362 ( \6705 , \6704 , \1960 );
and \U$6363 ( \6706 , \1844 , \1891 );
and \U$6364 ( \6707 , \1839 , \1889 );
nor \U$6365 ( \6708 , \6706 , \6707 );
xnor \U$6366 ( \6709 , \6708 , \1739 );
and \U$6367 ( \6710 , \6705 , \6709 );
and \U$6368 ( \6711 , \2174 , \1623 );
and \U$6369 ( \6712 , \2030 , \1621 );
nor \U$6370 ( \6713 , \6711 , \6712 );
xnor \U$6371 ( \6714 , \6713 , \1467 );
and \U$6372 ( \6715 , \6709 , \6714 );
and \U$6373 ( \6716 , \6705 , \6714 );
or \U$6374 ( \6717 , \6710 , \6715 , \6716 );
and \U$6375 ( \6718 , \6701 , \6717 );
and \U$6376 ( \6719 , \2463 , \1351 );
and \U$6377 ( \6720 , \2438 , \1349 );
nor \U$6378 ( \6721 , \6719 , \6720 );
xnor \U$6379 ( \6722 , \6721 , \1238 );
and \U$6380 ( \6723 , \2804 , \1157 );
and \U$6381 ( \6724 , \2637 , \1155 );
nor \U$6382 ( \6725 , \6723 , \6724 );
xnor \U$6383 ( \6726 , \6725 , \1021 );
and \U$6384 ( \6727 , \6722 , \6726 );
and \U$6385 ( \6728 , \3061 , \957 );
and \U$6386 ( \6729 , \2942 , \955 );
nor \U$6387 ( \6730 , \6728 , \6729 );
xnor \U$6388 ( \6731 , \6730 , \879 );
and \U$6389 ( \6732 , \6726 , \6731 );
and \U$6390 ( \6733 , \6722 , \6731 );
or \U$6391 ( \6734 , \6727 , \6732 , \6733 );
and \U$6392 ( \6735 , \6717 , \6734 );
and \U$6393 ( \6736 , \6701 , \6734 );
or \U$6394 ( \6737 , \6718 , \6735 , \6736 );
and \U$6395 ( \6738 , \385 , \5443 );
and \U$6396 ( \6739 , \393 , \5441 );
nor \U$6397 ( \6740 , \6738 , \6739 );
xnor \U$6398 ( \6741 , \6740 , \5202 );
and \U$6399 ( \6742 , \400 , \4977 );
and \U$6400 ( \6743 , \408 , \4975 );
nor \U$6401 ( \6744 , \6742 , \6743 );
xnor \U$6402 ( \6745 , \6744 , \4789 );
and \U$6403 ( \6746 , \6741 , \6745 );
and \U$6404 ( \6747 , \416 , \4603 );
and \U$6405 ( \6748 , \424 , \4601 );
nor \U$6406 ( \6749 , \6747 , \6748 );
xnor \U$6407 ( \6750 , \6749 , \4371 );
and \U$6408 ( \6751 , \6745 , \6750 );
and \U$6409 ( \6752 , \6741 , \6750 );
or \U$6410 ( \6753 , \6746 , \6751 , \6752 );
and \U$6411 ( \6754 , \435 , \4152 );
and \U$6412 ( \6755 , \443 , \4150 );
nor \U$6413 ( \6756 , \6754 , \6755 );
xnor \U$6414 ( \6757 , \6756 , \4009 );
and \U$6415 ( \6758 , \661 , \3829 );
and \U$6416 ( \6759 , \450 , \3827 );
nor \U$6417 ( \6760 , \6758 , \6759 );
xnor \U$6418 ( \6761 , \6760 , \3583 );
and \U$6419 ( \6762 , \6757 , \6761 );
and \U$6420 ( \6763 , \785 , \3434 );
and \U$6421 ( \6764 , \722 , \3432 );
nor \U$6422 ( \6765 , \6763 , \6764 );
xnor \U$6423 ( \6766 , \6765 , \3247 );
and \U$6424 ( \6767 , \6761 , \6766 );
and \U$6425 ( \6768 , \6757 , \6766 );
or \U$6426 ( \6769 , \6762 , \6767 , \6768 );
and \U$6427 ( \6770 , \6753 , \6769 );
buf \U$6428 ( \6771 , RIbb2de28_52);
buf \U$6429 ( \6772 , RIbb2ddb0_53);
and \U$6430 ( \6773 , \6771 , \6772 );
not \U$6431 ( \6774 , \6773 );
and \U$6432 ( \6775 , \6223 , \6774 );
not \U$6433 ( \6776 , \6775 );
and \U$6434 ( \6777 , \351 , \6541 );
and \U$6435 ( \6778 , \359 , \6539 );
nor \U$6436 ( \6779 , \6777 , \6778 );
xnor \U$6437 ( \6780 , \6779 , \6226 );
and \U$6438 ( \6781 , \6776 , \6780 );
and \U$6439 ( \6782 , \367 , \6032 );
and \U$6440 ( \6783 , \375 , \6030 );
nor \U$6441 ( \6784 , \6782 , \6783 );
xnor \U$6442 ( \6785 , \6784 , \5692 );
and \U$6443 ( \6786 , \6780 , \6785 );
and \U$6444 ( \6787 , \6776 , \6785 );
or \U$6445 ( \6788 , \6781 , \6786 , \6787 );
and \U$6446 ( \6789 , \6769 , \6788 );
and \U$6447 ( \6790 , \6753 , \6788 );
or \U$6448 ( \6791 , \6770 , \6789 , \6790 );
and \U$6449 ( \6792 , \6737 , \6791 );
and \U$6450 ( \6793 , \5954 , \422 );
and \U$6451 ( \6794 , \5945 , \420 );
nor \U$6452 ( \6795 , \6793 , \6794 );
xnor \U$6453 ( \6796 , \6795 , \429 );
and \U$6454 ( \6797 , \6499 , \441 );
and \U$6455 ( \6798 , \6297 , \439 );
nor \U$6456 ( \6799 , \6797 , \6798 );
xnor \U$6457 ( \6800 , \6799 , \448 );
and \U$6458 ( \6801 , \6796 , \6800 );
buf \U$6459 ( \6802 , RIbb2c0a0_115);
and \U$6460 ( \6803 , \6802 , \436 );
and \U$6461 ( \6804 , \6800 , \6803 );
and \U$6462 ( \6805 , \6796 , \6803 );
or \U$6463 ( \6806 , \6801 , \6804 , \6805 );
and \U$6464 ( \6807 , \3686 , \793 );
and \U$6465 ( \6808 , \3478 , \791 );
nor \U$6466 ( \6809 , \6807 , \6808 );
xnor \U$6467 ( \6810 , \6809 , \699 );
and \U$6468 ( \6811 , \3813 , \624 );
and \U$6469 ( \6812 , \3808 , \622 );
nor \U$6470 ( \6813 , \6811 , \6812 );
xnor \U$6471 ( \6814 , \6813 , \349 );
and \U$6472 ( \6815 , \6810 , \6814 );
and \U$6473 ( \6816 , \4266 , \357 );
and \U$6474 ( \6817 , \4069 , \355 );
nor \U$6475 ( \6818 , \6816 , \6817 );
xnor \U$6476 ( \6819 , \6818 , \364 );
and \U$6477 ( \6820 , \6814 , \6819 );
and \U$6478 ( \6821 , \6810 , \6819 );
or \U$6479 ( \6822 , \6815 , \6820 , \6821 );
and \U$6480 ( \6823 , \6806 , \6822 );
and \U$6481 ( \6824 , \4576 , \373 );
and \U$6482 ( \6825 , \4568 , \371 );
nor \U$6483 ( \6826 , \6824 , \6825 );
xnor \U$6484 ( \6827 , \6826 , \380 );
and \U$6485 ( \6828 , \5050 , \391 );
and \U$6486 ( \6829 , \5045 , \389 );
nor \U$6487 ( \6830 , \6828 , \6829 );
xnor \U$6488 ( \6831 , \6830 , \398 );
and \U$6489 ( \6832 , \6827 , \6831 );
and \U$6490 ( \6833 , \5573 , \406 );
and \U$6491 ( \6834 , \5314 , \404 );
nor \U$6492 ( \6835 , \6833 , \6834 );
xnor \U$6493 ( \6836 , \6835 , \413 );
and \U$6494 ( \6837 , \6831 , \6836 );
and \U$6495 ( \6838 , \6827 , \6836 );
or \U$6496 ( \6839 , \6832 , \6837 , \6838 );
and \U$6497 ( \6840 , \6822 , \6839 );
and \U$6498 ( \6841 , \6806 , \6839 );
or \U$6499 ( \6842 , \6823 , \6840 , \6841 );
and \U$6500 ( \6843 , \6791 , \6842 );
and \U$6501 ( \6844 , \6737 , \6842 );
or \U$6502 ( \6845 , \6792 , \6843 , \6844 );
xor \U$6503 ( \6846 , \6564 , \6568 );
xor \U$6504 ( \6847 , \6846 , \6573 );
xor \U$6505 ( \6848 , \6580 , \6584 );
xor \U$6506 ( \6849 , \6848 , \6589 );
and \U$6507 ( \6850 , \6847 , \6849 );
xor \U$6508 ( \6851 , \6597 , \6601 );
xor \U$6509 ( \6852 , \6851 , \6606 );
and \U$6510 ( \6853 , \6849 , \6852 );
and \U$6511 ( \6854 , \6847 , \6852 );
or \U$6512 ( \6855 , \6850 , \6853 , \6854 );
xor \U$6513 ( \6856 , \6508 , \6512 );
xor \U$6514 ( \6857 , \6856 , \6517 );
xor \U$6515 ( \6858 , \6524 , \6528 );
xor \U$6516 ( \6859 , \6858 , \6533 );
and \U$6517 ( \6860 , \6857 , \6859 );
xor \U$6518 ( \6861 , \6544 , \6548 );
xor \U$6519 ( \6862 , \6861 , \6553 );
and \U$6520 ( \6863 , \6859 , \6862 );
and \U$6521 ( \6864 , \6857 , \6862 );
or \U$6522 ( \6865 , \6860 , \6863 , \6864 );
and \U$6523 ( \6866 , \6855 , \6865 );
xor \U$6524 ( \6867 , \6465 , \6469 );
xor \U$6525 ( \6868 , \6867 , \6474 );
xor \U$6526 ( \6869 , \6481 , \6485 );
xor \U$6527 ( \6870 , \6869 , \6490 );
and \U$6528 ( \6871 , \6868 , \6870 );
xnor \U$6529 ( \6872 , \6498 , \6500 );
and \U$6530 ( \6873 , \6870 , \6872 );
and \U$6531 ( \6874 , \6868 , \6872 );
or \U$6532 ( \6875 , \6871 , \6873 , \6874 );
and \U$6533 ( \6876 , \6865 , \6875 );
and \U$6534 ( \6877 , \6855 , \6875 );
or \U$6535 ( \6878 , \6866 , \6876 , \6877 );
and \U$6536 ( \6879 , \6845 , \6878 );
xor \U$6537 ( \6880 , \6430 , \6432 );
xor \U$6538 ( \6881 , \6880 , \6435 );
xor \U$6539 ( \6882 , \6440 , \6442 );
xor \U$6540 ( \6883 , \6882 , \6445 );
and \U$6541 ( \6884 , \6881 , \6883 );
xor \U$6542 ( \6885 , \6451 , \6453 );
xor \U$6543 ( \6886 , \6885 , \6455 );
and \U$6544 ( \6887 , \6883 , \6886 );
and \U$6545 ( \6888 , \6881 , \6886 );
or \U$6546 ( \6889 , \6884 , \6887 , \6888 );
and \U$6547 ( \6890 , \6878 , \6889 );
and \U$6548 ( \6891 , \6845 , \6889 );
or \U$6549 ( \6892 , \6879 , \6890 , \6891 );
xor \U$6550 ( \6893 , \6477 , \6493 );
xor \U$6551 ( \6894 , \6893 , \6501 );
xor \U$6552 ( \6895 , \6520 , \6536 );
xor \U$6553 ( \6896 , \6895 , \6556 );
and \U$6554 ( \6897 , \6894 , \6896 );
xor \U$6555 ( \6898 , \6576 , \6592 );
xor \U$6556 ( \6899 , \6898 , \6609 );
and \U$6557 ( \6900 , \6896 , \6899 );
and \U$6558 ( \6901 , \6894 , \6899 );
or \U$6559 ( \6902 , \6897 , \6900 , \6901 );
xor \U$6560 ( \6903 , \6631 , \6633 );
xor \U$6561 ( \6904 , \6903 , \6636 );
and \U$6562 ( \6905 , \6902 , \6904 );
xor \U$6563 ( \6906 , \6618 , \6620 );
xor \U$6564 ( \6907 , \6906 , \6623 );
and \U$6565 ( \6908 , \6904 , \6907 );
and \U$6566 ( \6909 , \6902 , \6907 );
or \U$6567 ( \6910 , \6905 , \6908 , \6909 );
and \U$6568 ( \6911 , \6892 , \6910 );
xor \U$6569 ( \6912 , \6438 , \6448 );
xor \U$6570 ( \6913 , \6912 , \6458 );
xor \U$6571 ( \6914 , \6504 , \6559 );
xor \U$6572 ( \6915 , \6914 , \6612 );
and \U$6573 ( \6916 , \6913 , \6915 );
and \U$6574 ( \6917 , \6910 , \6916 );
and \U$6575 ( \6918 , \6892 , \6916 );
or \U$6576 ( \6919 , \6911 , \6917 , \6918 );
xor \U$6577 ( \6920 , \6461 , \6615 );
xor \U$6578 ( \6921 , \6920 , \6626 );
xor \U$6579 ( \6922 , \6639 , \6641 );
xor \U$6580 ( \6923 , \6922 , \6644 );
and \U$6581 ( \6924 , \6921 , \6923 );
xor \U$6582 ( \6925 , \6650 , \6652 );
and \U$6583 ( \6926 , \6923 , \6925 );
and \U$6584 ( \6927 , \6921 , \6925 );
or \U$6585 ( \6928 , \6924 , \6926 , \6927 );
and \U$6586 ( \6929 , \6919 , \6928 );
xor \U$6587 ( \6930 , \6658 , \6660 );
xor \U$6588 ( \6931 , \6930 , \6662 );
and \U$6589 ( \6932 , \6928 , \6931 );
and \U$6590 ( \6933 , \6919 , \6931 );
or \U$6591 ( \6934 , \6929 , \6932 , \6933 );
xor \U$6592 ( \6935 , \6372 , \6390 );
xor \U$6593 ( \6936 , \6935 , \6396 );
and \U$6594 ( \6937 , \6934 , \6936 );
xor \U$6595 ( \6938 , \6656 , \6665 );
xor \U$6596 ( \6939 , \6938 , \6668 );
and \U$6597 ( \6940 , \6936 , \6939 );
and \U$6598 ( \6941 , \6934 , \6939 );
or \U$6599 ( \6942 , \6937 , \6940 , \6941 );
xor \U$6600 ( \6943 , \6671 , \6673 );
xor \U$6601 ( \6944 , \6943 , \6676 );
and \U$6602 ( \6945 , \6942 , \6944 );
and \U$6603 ( \6946 , \6685 , \6945 );
xor \U$6604 ( \6947 , \6685 , \6945 );
xor \U$6605 ( \6948 , \6942 , \6944 );
and \U$6606 ( \6949 , \3808 , \793 );
and \U$6607 ( \6950 , \3686 , \791 );
nor \U$6608 ( \6951 , \6949 , \6950 );
xnor \U$6609 ( \6952 , \6951 , \699 );
and \U$6610 ( \6953 , \4069 , \624 );
and \U$6611 ( \6954 , \3813 , \622 );
nor \U$6612 ( \6955 , \6953 , \6954 );
xnor \U$6613 ( \6956 , \6955 , \349 );
and \U$6614 ( \6957 , \6952 , \6956 );
and \U$6615 ( \6958 , \4568 , \357 );
and \U$6616 ( \6959 , \4266 , \355 );
nor \U$6617 ( \6960 , \6958 , \6959 );
xnor \U$6618 ( \6961 , \6960 , \364 );
and \U$6619 ( \6962 , \6956 , \6961 );
and \U$6620 ( \6963 , \6952 , \6961 );
or \U$6621 ( \6964 , \6957 , \6962 , \6963 );
and \U$6622 ( \6965 , \6297 , \422 );
and \U$6623 ( \6966 , \5954 , \420 );
nor \U$6624 ( \6967 , \6965 , \6966 );
xnor \U$6625 ( \6968 , \6967 , \429 );
and \U$6626 ( \6969 , \6802 , \441 );
and \U$6627 ( \6970 , \6499 , \439 );
nor \U$6628 ( \6971 , \6969 , \6970 );
xnor \U$6629 ( \6972 , \6971 , \448 );
and \U$6630 ( \6973 , \6968 , \6972 );
buf \U$6631 ( \6974 , RIbb2c028_116);
and \U$6632 ( \6975 , \6974 , \436 );
and \U$6633 ( \6976 , \6972 , \6975 );
and \U$6634 ( \6977 , \6968 , \6975 );
or \U$6635 ( \6978 , \6973 , \6976 , \6977 );
and \U$6636 ( \6979 , \6964 , \6978 );
and \U$6637 ( \6980 , \5045 , \373 );
and \U$6638 ( \6981 , \4576 , \371 );
nor \U$6639 ( \6982 , \6980 , \6981 );
xnor \U$6640 ( \6983 , \6982 , \380 );
and \U$6641 ( \6984 , \5314 , \391 );
and \U$6642 ( \6985 , \5050 , \389 );
nor \U$6643 ( \6986 , \6984 , \6985 );
xnor \U$6644 ( \6987 , \6986 , \398 );
and \U$6645 ( \6988 , \6983 , \6987 );
and \U$6646 ( \6989 , \5945 , \406 );
and \U$6647 ( \6990 , \5573 , \404 );
nor \U$6648 ( \6991 , \6989 , \6990 );
xnor \U$6649 ( \6992 , \6991 , \413 );
and \U$6650 ( \6993 , \6987 , \6992 );
and \U$6651 ( \6994 , \6983 , \6992 );
or \U$6652 ( \6995 , \6988 , \6993 , \6994 );
and \U$6653 ( \6996 , \6978 , \6995 );
and \U$6654 ( \6997 , \6964 , \6995 );
or \U$6655 ( \6998 , \6979 , \6996 , \6997 );
and \U$6656 ( \6999 , \408 , \5443 );
and \U$6657 ( \7000 , \385 , \5441 );
nor \U$6658 ( \7001 , \6999 , \7000 );
xnor \U$6659 ( \7002 , \7001 , \5202 );
and \U$6660 ( \7003 , \424 , \4977 );
and \U$6661 ( \7004 , \400 , \4975 );
nor \U$6662 ( \7005 , \7003 , \7004 );
xnor \U$6663 ( \7006 , \7005 , \4789 );
and \U$6664 ( \7007 , \7002 , \7006 );
and \U$6665 ( \7008 , \443 , \4603 );
and \U$6666 ( \7009 , \416 , \4601 );
nor \U$6667 ( \7010 , \7008 , \7009 );
xnor \U$6668 ( \7011 , \7010 , \4371 );
and \U$6669 ( \7012 , \7006 , \7011 );
and \U$6670 ( \7013 , \7002 , \7011 );
or \U$6671 ( \7014 , \7007 , \7012 , \7013 );
and \U$6672 ( \7015 , \450 , \4152 );
and \U$6673 ( \7016 , \435 , \4150 );
nor \U$6674 ( \7017 , \7015 , \7016 );
xnor \U$6675 ( \7018 , \7017 , \4009 );
and \U$6676 ( \7019 , \722 , \3829 );
and \U$6677 ( \7020 , \661 , \3827 );
nor \U$6678 ( \7021 , \7019 , \7020 );
xnor \U$6679 ( \7022 , \7021 , \3583 );
and \U$6680 ( \7023 , \7018 , \7022 );
and \U$6681 ( \7024 , \983 , \3434 );
and \U$6682 ( \7025 , \785 , \3432 );
nor \U$6683 ( \7026 , \7024 , \7025 );
xnor \U$6684 ( \7027 , \7026 , \3247 );
and \U$6685 ( \7028 , \7022 , \7027 );
and \U$6686 ( \7029 , \7018 , \7027 );
or \U$6687 ( \7030 , \7023 , \7028 , \7029 );
and \U$6688 ( \7031 , \7014 , \7030 );
xor \U$6689 ( \7032 , \6223 , \6771 );
xor \U$6690 ( \7033 , \6771 , \6772 );
not \U$6691 ( \7034 , \7033 );
and \U$6692 ( \7035 , \7032 , \7034 );
and \U$6693 ( \7036 , \359 , \7035 );
not \U$6694 ( \7037 , \7036 );
xnor \U$6695 ( \7038 , \7037 , \6775 );
and \U$6696 ( \7039 , \375 , \6541 );
and \U$6697 ( \7040 , \351 , \6539 );
nor \U$6698 ( \7041 , \7039 , \7040 );
xnor \U$6699 ( \7042 , \7041 , \6226 );
and \U$6700 ( \7043 , \7038 , \7042 );
and \U$6701 ( \7044 , \393 , \6032 );
and \U$6702 ( \7045 , \367 , \6030 );
nor \U$6703 ( \7046 , \7044 , \7045 );
xnor \U$6704 ( \7047 , \7046 , \5692 );
and \U$6705 ( \7048 , \7042 , \7047 );
and \U$6706 ( \7049 , \7038 , \7047 );
or \U$6707 ( \7050 , \7043 , \7048 , \7049 );
and \U$6708 ( \7051 , \7030 , \7050 );
and \U$6709 ( \7052 , \7014 , \7050 );
or \U$6710 ( \7053 , \7031 , \7051 , \7052 );
and \U$6711 ( \7054 , \6998 , \7053 );
and \U$6712 ( \7055 , \1176 , \3121 );
and \U$6713 ( \7056 , \1071 , \3119 );
nor \U$6714 ( \7057 , \7055 , \7056 );
xnor \U$6715 ( \7058 , \7057 , \2916 );
and \U$6716 ( \7059 , \1297 , \2715 );
and \U$6717 ( \7060 , \1181 , \2713 );
nor \U$6718 ( \7061 , \7059 , \7060 );
xnor \U$6719 ( \7062 , \7061 , \2566 );
and \U$6720 ( \7063 , \7058 , \7062 );
and \U$6721 ( \7064 , \1588 , \2393 );
and \U$6722 ( \7065 , \1412 , \2391 );
nor \U$6723 ( \7066 , \7064 , \7065 );
xnor \U$6724 ( \7067 , \7066 , \2251 );
and \U$6725 ( \7068 , \7062 , \7067 );
and \U$6726 ( \7069 , \7058 , \7067 );
or \U$6727 ( \7070 , \7063 , \7068 , \7069 );
and \U$6728 ( \7071 , \1839 , \2097 );
and \U$6729 ( \7072 , \1596 , \2095 );
nor \U$6730 ( \7073 , \7071 , \7072 );
xnor \U$6731 ( \7074 , \7073 , \1960 );
and \U$6732 ( \7075 , \2030 , \1891 );
and \U$6733 ( \7076 , \1844 , \1889 );
nor \U$6734 ( \7077 , \7075 , \7076 );
xnor \U$6735 ( \7078 , \7077 , \1739 );
and \U$6736 ( \7079 , \7074 , \7078 );
and \U$6737 ( \7080 , \2438 , \1623 );
and \U$6738 ( \7081 , \2174 , \1621 );
nor \U$6739 ( \7082 , \7080 , \7081 );
xnor \U$6740 ( \7083 , \7082 , \1467 );
and \U$6741 ( \7084 , \7078 , \7083 );
and \U$6742 ( \7085 , \7074 , \7083 );
or \U$6743 ( \7086 , \7079 , \7084 , \7085 );
and \U$6744 ( \7087 , \7070 , \7086 );
and \U$6745 ( \7088 , \2637 , \1351 );
and \U$6746 ( \7089 , \2463 , \1349 );
nor \U$6747 ( \7090 , \7088 , \7089 );
xnor \U$6748 ( \7091 , \7090 , \1238 );
and \U$6749 ( \7092 , \2942 , \1157 );
and \U$6750 ( \7093 , \2804 , \1155 );
nor \U$6751 ( \7094 , \7092 , \7093 );
xnor \U$6752 ( \7095 , \7094 , \1021 );
and \U$6753 ( \7096 , \7091 , \7095 );
and \U$6754 ( \7097 , \3478 , \957 );
and \U$6755 ( \7098 , \3061 , \955 );
nor \U$6756 ( \7099 , \7097 , \7098 );
xnor \U$6757 ( \7100 , \7099 , \879 );
and \U$6758 ( \7101 , \7095 , \7100 );
and \U$6759 ( \7102 , \7091 , \7100 );
or \U$6760 ( \7103 , \7096 , \7101 , \7102 );
and \U$6761 ( \7104 , \7086 , \7103 );
and \U$6762 ( \7105 , \7070 , \7103 );
or \U$6763 ( \7106 , \7087 , \7104 , \7105 );
and \U$6764 ( \7107 , \7053 , \7106 );
and \U$6765 ( \7108 , \6998 , \7106 );
or \U$6766 ( \7109 , \7054 , \7107 , \7108 );
xor \U$6767 ( \7110 , \6796 , \6800 );
xor \U$6768 ( \7111 , \7110 , \6803 );
xor \U$6769 ( \7112 , \6810 , \6814 );
xor \U$6770 ( \7113 , \7112 , \6819 );
and \U$6771 ( \7114 , \7111 , \7113 );
xor \U$6772 ( \7115 , \6827 , \6831 );
xor \U$6773 ( \7116 , \7115 , \6836 );
and \U$6774 ( \7117 , \7113 , \7116 );
and \U$6775 ( \7118 , \7111 , \7116 );
or \U$6776 ( \7119 , \7114 , \7117 , \7118 );
xor \U$6777 ( \7120 , \6689 , \6693 );
xor \U$6778 ( \7121 , \7120 , \6698 );
xor \U$6779 ( \7122 , \6705 , \6709 );
xor \U$6780 ( \7123 , \7122 , \6714 );
and \U$6781 ( \7124 , \7121 , \7123 );
xor \U$6782 ( \7125 , \6722 , \6726 );
xor \U$6783 ( \7126 , \7125 , \6731 );
and \U$6784 ( \7127 , \7123 , \7126 );
and \U$6785 ( \7128 , \7121 , \7126 );
or \U$6786 ( \7129 , \7124 , \7127 , \7128 );
and \U$6787 ( \7130 , \7119 , \7129 );
xor \U$6788 ( \7131 , \6741 , \6745 );
xor \U$6789 ( \7132 , \7131 , \6750 );
xor \U$6790 ( \7133 , \6757 , \6761 );
xor \U$6791 ( \7134 , \7133 , \6766 );
and \U$6792 ( \7135 , \7132 , \7134 );
xor \U$6793 ( \7136 , \6776 , \6780 );
xor \U$6794 ( \7137 , \7136 , \6785 );
and \U$6795 ( \7138 , \7134 , \7137 );
and \U$6796 ( \7139 , \7132 , \7137 );
or \U$6797 ( \7140 , \7135 , \7138 , \7139 );
and \U$6798 ( \7141 , \7129 , \7140 );
and \U$6799 ( \7142 , \7119 , \7140 );
or \U$6800 ( \7143 , \7130 , \7141 , \7142 );
and \U$6801 ( \7144 , \7109 , \7143 );
xor \U$6802 ( \7145 , \6847 , \6849 );
xor \U$6803 ( \7146 , \7145 , \6852 );
xor \U$6804 ( \7147 , \6857 , \6859 );
xor \U$6805 ( \7148 , \7147 , \6862 );
and \U$6806 ( \7149 , \7146 , \7148 );
xor \U$6807 ( \7150 , \6868 , \6870 );
xor \U$6808 ( \7151 , \7150 , \6872 );
and \U$6809 ( \7152 , \7148 , \7151 );
and \U$6810 ( \7153 , \7146 , \7151 );
or \U$6811 ( \7154 , \7149 , \7152 , \7153 );
and \U$6812 ( \7155 , \7143 , \7154 );
and \U$6813 ( \7156 , \7109 , \7154 );
or \U$6814 ( \7157 , \7144 , \7155 , \7156 );
xor \U$6815 ( \7158 , \6701 , \6717 );
xor \U$6816 ( \7159 , \7158 , \6734 );
xor \U$6817 ( \7160 , \6753 , \6769 );
xor \U$6818 ( \7161 , \7160 , \6788 );
and \U$6819 ( \7162 , \7159 , \7161 );
xor \U$6820 ( \7163 , \6806 , \6822 );
xor \U$6821 ( \7164 , \7163 , \6839 );
and \U$6822 ( \7165 , \7161 , \7164 );
and \U$6823 ( \7166 , \7159 , \7164 );
or \U$6824 ( \7167 , \7162 , \7165 , \7166 );
xor \U$6825 ( \7168 , \6894 , \6896 );
xor \U$6826 ( \7169 , \7168 , \6899 );
and \U$6827 ( \7170 , \7167 , \7169 );
xor \U$6828 ( \7171 , \6881 , \6883 );
xor \U$6829 ( \7172 , \7171 , \6886 );
and \U$6830 ( \7173 , \7169 , \7172 );
and \U$6831 ( \7174 , \7167 , \7172 );
or \U$6832 ( \7175 , \7170 , \7173 , \7174 );
and \U$6833 ( \7176 , \7157 , \7175 );
xor \U$6834 ( \7177 , \6737 , \6791 );
xor \U$6835 ( \7178 , \7177 , \6842 );
xor \U$6836 ( \7179 , \6855 , \6865 );
xor \U$6837 ( \7180 , \7179 , \6875 );
and \U$6838 ( \7181 , \7178 , \7180 );
and \U$6839 ( \7182 , \7175 , \7181 );
and \U$6840 ( \7183 , \7157 , \7181 );
or \U$6841 ( \7184 , \7176 , \7182 , \7183 );
xor \U$6842 ( \7185 , \6845 , \6878 );
xor \U$6843 ( \7186 , \7185 , \6889 );
xor \U$6844 ( \7187 , \6902 , \6904 );
xor \U$6845 ( \7188 , \7187 , \6907 );
and \U$6846 ( \7189 , \7186 , \7188 );
xor \U$6847 ( \7190 , \6913 , \6915 );
and \U$6848 ( \7191 , \7188 , \7190 );
and \U$6849 ( \7192 , \7186 , \7190 );
or \U$6850 ( \7193 , \7189 , \7191 , \7192 );
and \U$6851 ( \7194 , \7184 , \7193 );
xor \U$6852 ( \7195 , \6921 , \6923 );
xor \U$6853 ( \7196 , \7195 , \6925 );
and \U$6854 ( \7197 , \7193 , \7196 );
and \U$6855 ( \7198 , \7184 , \7196 );
or \U$6856 ( \7199 , \7194 , \7197 , \7198 );
xor \U$6857 ( \7200 , \6629 , \6647 );
xor \U$6858 ( \7201 , \7200 , \6653 );
and \U$6859 ( \7202 , \7199 , \7201 );
xor \U$6860 ( \7203 , \6919 , \6928 );
xor \U$6861 ( \7204 , \7203 , \6931 );
and \U$6862 ( \7205 , \7201 , \7204 );
and \U$6863 ( \7206 , \7199 , \7204 );
or \U$6864 ( \7207 , \7202 , \7205 , \7206 );
xor \U$6865 ( \7208 , \6934 , \6936 );
xor \U$6866 ( \7209 , \7208 , \6939 );
and \U$6867 ( \7210 , \7207 , \7209 );
and \U$6868 ( \7211 , \6948 , \7210 );
xor \U$6869 ( \7212 , \6948 , \7210 );
xor \U$6870 ( \7213 , \7207 , \7209 );
xor \U$6871 ( \7214 , \7002 , \7006 );
xor \U$6872 ( \7215 , \7214 , \7011 );
xor \U$6873 ( \7216 , \7058 , \7062 );
xor \U$6874 ( \7217 , \7216 , \7067 );
and \U$6875 ( \7218 , \7215 , \7217 );
xor \U$6876 ( \7219 , \7018 , \7022 );
xor \U$6877 ( \7220 , \7219 , \7027 );
and \U$6878 ( \7221 , \7217 , \7220 );
and \U$6879 ( \7222 , \7215 , \7220 );
or \U$6880 ( \7223 , \7218 , \7221 , \7222 );
xor \U$6881 ( \7224 , \7074 , \7078 );
xor \U$6882 ( \7225 , \7224 , \7083 );
xor \U$6883 ( \7226 , \6952 , \6956 );
xor \U$6884 ( \7227 , \7226 , \6961 );
and \U$6885 ( \7228 , \7225 , \7227 );
xor \U$6886 ( \7229 , \7091 , \7095 );
xor \U$6887 ( \7230 , \7229 , \7100 );
and \U$6888 ( \7231 , \7227 , \7230 );
and \U$6889 ( \7232 , \7225 , \7230 );
or \U$6890 ( \7233 , \7228 , \7231 , \7232 );
and \U$6891 ( \7234 , \7223 , \7233 );
xor \U$6892 ( \7235 , \6968 , \6972 );
xor \U$6893 ( \7236 , \7235 , \6975 );
xor \U$6894 ( \7237 , \6983 , \6987 );
xor \U$6895 ( \7238 , \7237 , \6992 );
or \U$6896 ( \7239 , \7236 , \7238 );
and \U$6897 ( \7240 , \7233 , \7239 );
and \U$6898 ( \7241 , \7223 , \7239 );
or \U$6899 ( \7242 , \7234 , \7240 , \7241 );
and \U$6900 ( \7243 , \1596 , \2393 );
and \U$6901 ( \7244 , \1588 , \2391 );
nor \U$6902 ( \7245 , \7243 , \7244 );
xnor \U$6903 ( \7246 , \7245 , \2251 );
and \U$6904 ( \7247 , \1844 , \2097 );
and \U$6905 ( \7248 , \1839 , \2095 );
nor \U$6906 ( \7249 , \7247 , \7248 );
xnor \U$6907 ( \7250 , \7249 , \1960 );
and \U$6908 ( \7251 , \7246 , \7250 );
and \U$6909 ( \7252 , \2174 , \1891 );
and \U$6910 ( \7253 , \2030 , \1889 );
nor \U$6911 ( \7254 , \7252 , \7253 );
xnor \U$6912 ( \7255 , \7254 , \1739 );
and \U$6913 ( \7256 , \7250 , \7255 );
and \U$6914 ( \7257 , \7246 , \7255 );
or \U$6915 ( \7258 , \7251 , \7256 , \7257 );
and \U$6916 ( \7259 , \1071 , \3434 );
and \U$6917 ( \7260 , \983 , \3432 );
nor \U$6918 ( \7261 , \7259 , \7260 );
xnor \U$6919 ( \7262 , \7261 , \3247 );
and \U$6920 ( \7263 , \1181 , \3121 );
and \U$6921 ( \7264 , \1176 , \3119 );
nor \U$6922 ( \7265 , \7263 , \7264 );
xnor \U$6923 ( \7266 , \7265 , \2916 );
and \U$6924 ( \7267 , \7262 , \7266 );
and \U$6925 ( \7268 , \1412 , \2715 );
and \U$6926 ( \7269 , \1297 , \2713 );
nor \U$6927 ( \7270 , \7268 , \7269 );
xnor \U$6928 ( \7271 , \7270 , \2566 );
and \U$6929 ( \7272 , \7266 , \7271 );
and \U$6930 ( \7273 , \7262 , \7271 );
or \U$6931 ( \7274 , \7267 , \7272 , \7273 );
and \U$6932 ( \7275 , \7258 , \7274 );
and \U$6933 ( \7276 , \2463 , \1623 );
and \U$6934 ( \7277 , \2438 , \1621 );
nor \U$6935 ( \7278 , \7276 , \7277 );
xnor \U$6936 ( \7279 , \7278 , \1467 );
and \U$6937 ( \7280 , \2804 , \1351 );
and \U$6938 ( \7281 , \2637 , \1349 );
nor \U$6939 ( \7282 , \7280 , \7281 );
xnor \U$6940 ( \7283 , \7282 , \1238 );
and \U$6941 ( \7284 , \7279 , \7283 );
and \U$6942 ( \7285 , \3061 , \1157 );
and \U$6943 ( \7286 , \2942 , \1155 );
nor \U$6944 ( \7287 , \7285 , \7286 );
xnor \U$6945 ( \7288 , \7287 , \1021 );
and \U$6946 ( \7289 , \7283 , \7288 );
and \U$6947 ( \7290 , \7279 , \7288 );
or \U$6948 ( \7291 , \7284 , \7289 , \7290 );
and \U$6949 ( \7292 , \7274 , \7291 );
and \U$6950 ( \7293 , \7258 , \7291 );
or \U$6951 ( \7294 , \7275 , \7292 , \7293 );
and \U$6952 ( \7295 , \385 , \6032 );
and \U$6953 ( \7296 , \393 , \6030 );
nor \U$6954 ( \7297 , \7295 , \7296 );
xnor \U$6955 ( \7298 , \7297 , \5692 );
and \U$6956 ( \7299 , \400 , \5443 );
and \U$6957 ( \7300 , \408 , \5441 );
nor \U$6958 ( \7301 , \7299 , \7300 );
xnor \U$6959 ( \7302 , \7301 , \5202 );
and \U$6960 ( \7303 , \7298 , \7302 );
and \U$6961 ( \7304 , \416 , \4977 );
and \U$6962 ( \7305 , \424 , \4975 );
nor \U$6963 ( \7306 , \7304 , \7305 );
xnor \U$6964 ( \7307 , \7306 , \4789 );
and \U$6965 ( \7308 , \7302 , \7307 );
and \U$6966 ( \7309 , \7298 , \7307 );
or \U$6967 ( \7310 , \7303 , \7308 , \7309 );
buf \U$6968 ( \7311 , RIbb2dd38_54);
buf \U$6969 ( \7312 , RIbb2dcc0_55);
and \U$6970 ( \7313 , \7311 , \7312 );
not \U$6971 ( \7314 , \7313 );
and \U$6972 ( \7315 , \6772 , \7314 );
not \U$6973 ( \7316 , \7315 );
and \U$6974 ( \7317 , \351 , \7035 );
and \U$6975 ( \7318 , \359 , \7033 );
nor \U$6976 ( \7319 , \7317 , \7318 );
xnor \U$6977 ( \7320 , \7319 , \6775 );
and \U$6978 ( \7321 , \7316 , \7320 );
and \U$6979 ( \7322 , \367 , \6541 );
and \U$6980 ( \7323 , \375 , \6539 );
nor \U$6981 ( \7324 , \7322 , \7323 );
xnor \U$6982 ( \7325 , \7324 , \6226 );
and \U$6983 ( \7326 , \7320 , \7325 );
and \U$6984 ( \7327 , \7316 , \7325 );
or \U$6985 ( \7328 , \7321 , \7326 , \7327 );
and \U$6986 ( \7329 , \7310 , \7328 );
and \U$6987 ( \7330 , \435 , \4603 );
and \U$6988 ( \7331 , \443 , \4601 );
nor \U$6989 ( \7332 , \7330 , \7331 );
xnor \U$6990 ( \7333 , \7332 , \4371 );
and \U$6991 ( \7334 , \661 , \4152 );
and \U$6992 ( \7335 , \450 , \4150 );
nor \U$6993 ( \7336 , \7334 , \7335 );
xnor \U$6994 ( \7337 , \7336 , \4009 );
and \U$6995 ( \7338 , \7333 , \7337 );
and \U$6996 ( \7339 , \785 , \3829 );
and \U$6997 ( \7340 , \722 , \3827 );
nor \U$6998 ( \7341 , \7339 , \7340 );
xnor \U$6999 ( \7342 , \7341 , \3583 );
and \U$7000 ( \7343 , \7337 , \7342 );
and \U$7001 ( \7344 , \7333 , \7342 );
or \U$7002 ( \7345 , \7338 , \7343 , \7344 );
and \U$7003 ( \7346 , \7328 , \7345 );
and \U$7004 ( \7347 , \7310 , \7345 );
or \U$7005 ( \7348 , \7329 , \7346 , \7347 );
and \U$7006 ( \7349 , \7294 , \7348 );
and \U$7007 ( \7350 , \3686 , \957 );
and \U$7008 ( \7351 , \3478 , \955 );
nor \U$7009 ( \7352 , \7350 , \7351 );
xnor \U$7010 ( \7353 , \7352 , \879 );
and \U$7011 ( \7354 , \3813 , \793 );
and \U$7012 ( \7355 , \3808 , \791 );
nor \U$7013 ( \7356 , \7354 , \7355 );
xnor \U$7014 ( \7357 , \7356 , \699 );
and \U$7015 ( \7358 , \7353 , \7357 );
and \U$7016 ( \7359 , \4266 , \624 );
and \U$7017 ( \7360 , \4069 , \622 );
nor \U$7018 ( \7361 , \7359 , \7360 );
xnor \U$7019 ( \7362 , \7361 , \349 );
and \U$7020 ( \7363 , \7357 , \7362 );
and \U$7021 ( \7364 , \7353 , \7362 );
or \U$7022 ( \7365 , \7358 , \7363 , \7364 );
and \U$7023 ( \7366 , \4576 , \357 );
and \U$7024 ( \7367 , \4568 , \355 );
nor \U$7025 ( \7368 , \7366 , \7367 );
xnor \U$7026 ( \7369 , \7368 , \364 );
and \U$7027 ( \7370 , \5050 , \373 );
and \U$7028 ( \7371 , \5045 , \371 );
nor \U$7029 ( \7372 , \7370 , \7371 );
xnor \U$7030 ( \7373 , \7372 , \380 );
and \U$7031 ( \7374 , \7369 , \7373 );
and \U$7032 ( \7375 , \5573 , \391 );
and \U$7033 ( \7376 , \5314 , \389 );
nor \U$7034 ( \7377 , \7375 , \7376 );
xnor \U$7035 ( \7378 , \7377 , \398 );
and \U$7036 ( \7379 , \7373 , \7378 );
and \U$7037 ( \7380 , \7369 , \7378 );
or \U$7038 ( \7381 , \7374 , \7379 , \7380 );
and \U$7039 ( \7382 , \7365 , \7381 );
and \U$7040 ( \7383 , \5954 , \406 );
and \U$7041 ( \7384 , \5945 , \404 );
nor \U$7042 ( \7385 , \7383 , \7384 );
xnor \U$7043 ( \7386 , \7385 , \413 );
and \U$7044 ( \7387 , \6499 , \422 );
and \U$7045 ( \7388 , \6297 , \420 );
nor \U$7046 ( \7389 , \7387 , \7388 );
xnor \U$7047 ( \7390 , \7389 , \429 );
and \U$7048 ( \7391 , \7386 , \7390 );
and \U$7049 ( \7392 , \6974 , \441 );
and \U$7050 ( \7393 , \6802 , \439 );
nor \U$7051 ( \7394 , \7392 , \7393 );
xnor \U$7052 ( \7395 , \7394 , \448 );
and \U$7053 ( \7396 , \7390 , \7395 );
and \U$7054 ( \7397 , \7386 , \7395 );
or \U$7055 ( \7398 , \7391 , \7396 , \7397 );
and \U$7056 ( \7399 , \7381 , \7398 );
and \U$7057 ( \7400 , \7365 , \7398 );
or \U$7058 ( \7401 , \7382 , \7399 , \7400 );
and \U$7059 ( \7402 , \7348 , \7401 );
and \U$7060 ( \7403 , \7294 , \7401 );
or \U$7061 ( \7404 , \7349 , \7402 , \7403 );
and \U$7062 ( \7405 , \7242 , \7404 );
xor \U$7063 ( \7406 , \7111 , \7113 );
xor \U$7064 ( \7407 , \7406 , \7116 );
xor \U$7065 ( \7408 , \7121 , \7123 );
xor \U$7066 ( \7409 , \7408 , \7126 );
and \U$7067 ( \7410 , \7407 , \7409 );
xor \U$7068 ( \7411 , \7132 , \7134 );
xor \U$7069 ( \7412 , \7411 , \7137 );
and \U$7070 ( \7413 , \7409 , \7412 );
and \U$7071 ( \7414 , \7407 , \7412 );
or \U$7072 ( \7415 , \7410 , \7413 , \7414 );
and \U$7073 ( \7416 , \7404 , \7415 );
and \U$7074 ( \7417 , \7242 , \7415 );
or \U$7075 ( \7418 , \7405 , \7416 , \7417 );
xor \U$7076 ( \7419 , \6964 , \6978 );
xor \U$7077 ( \7420 , \7419 , \6995 );
xor \U$7078 ( \7421 , \7014 , \7030 );
xor \U$7079 ( \7422 , \7421 , \7050 );
and \U$7080 ( \7423 , \7420 , \7422 );
xor \U$7081 ( \7424 , \7070 , \7086 );
xor \U$7082 ( \7425 , \7424 , \7103 );
and \U$7083 ( \7426 , \7422 , \7425 );
and \U$7084 ( \7427 , \7420 , \7425 );
or \U$7085 ( \7428 , \7423 , \7426 , \7427 );
xor \U$7086 ( \7429 , \7159 , \7161 );
xor \U$7087 ( \7430 , \7429 , \7164 );
and \U$7088 ( \7431 , \7428 , \7430 );
xor \U$7089 ( \7432 , \7146 , \7148 );
xor \U$7090 ( \7433 , \7432 , \7151 );
and \U$7091 ( \7434 , \7430 , \7433 );
and \U$7092 ( \7435 , \7428 , \7433 );
or \U$7093 ( \7436 , \7431 , \7434 , \7435 );
and \U$7094 ( \7437 , \7418 , \7436 );
xor \U$7095 ( \7438 , \6998 , \7053 );
xor \U$7096 ( \7439 , \7438 , \7106 );
xor \U$7097 ( \7440 , \7119 , \7129 );
xor \U$7098 ( \7441 , \7440 , \7140 );
and \U$7099 ( \7442 , \7439 , \7441 );
and \U$7100 ( \7443 , \7436 , \7442 );
and \U$7101 ( \7444 , \7418 , \7442 );
or \U$7102 ( \7445 , \7437 , \7443 , \7444 );
xor \U$7103 ( \7446 , \7109 , \7143 );
xor \U$7104 ( \7447 , \7446 , \7154 );
xor \U$7105 ( \7448 , \7167 , \7169 );
xor \U$7106 ( \7449 , \7448 , \7172 );
and \U$7107 ( \7450 , \7447 , \7449 );
xor \U$7108 ( \7451 , \7178 , \7180 );
and \U$7109 ( \7452 , \7449 , \7451 );
and \U$7110 ( \7453 , \7447 , \7451 );
or \U$7111 ( \7454 , \7450 , \7452 , \7453 );
and \U$7112 ( \7455 , \7445 , \7454 );
xor \U$7113 ( \7456 , \7186 , \7188 );
xor \U$7114 ( \7457 , \7456 , \7190 );
and \U$7115 ( \7458 , \7454 , \7457 );
and \U$7116 ( \7459 , \7445 , \7457 );
or \U$7117 ( \7460 , \7455 , \7458 , \7459 );
xor \U$7118 ( \7461 , \6892 , \6910 );
xor \U$7119 ( \7462 , \7461 , \6916 );
and \U$7120 ( \7463 , \7460 , \7462 );
xor \U$7121 ( \7464 , \7184 , \7193 );
xor \U$7122 ( \7465 , \7464 , \7196 );
and \U$7123 ( \7466 , \7462 , \7465 );
and \U$7124 ( \7467 , \7460 , \7465 );
or \U$7125 ( \7468 , \7463 , \7466 , \7467 );
xor \U$7126 ( \7469 , \7199 , \7201 );
xor \U$7127 ( \7470 , \7469 , \7204 );
and \U$7128 ( \7471 , \7468 , \7470 );
and \U$7129 ( \7472 , \7213 , \7471 );
xor \U$7130 ( \7473 , \7213 , \7471 );
xor \U$7131 ( \7474 , \7468 , \7470 );
and \U$7132 ( \7475 , \3808 , \957 );
and \U$7133 ( \7476 , \3686 , \955 );
nor \U$7134 ( \7477 , \7475 , \7476 );
xnor \U$7135 ( \7478 , \7477 , \879 );
and \U$7136 ( \7479 , \4069 , \793 );
and \U$7137 ( \7480 , \3813 , \791 );
nor \U$7138 ( \7481 , \7479 , \7480 );
xnor \U$7139 ( \7482 , \7481 , \699 );
and \U$7140 ( \7483 , \7478 , \7482 );
and \U$7141 ( \7484 , \4568 , \624 );
and \U$7142 ( \7485 , \4266 , \622 );
nor \U$7143 ( \7486 , \7484 , \7485 );
xnor \U$7144 ( \7487 , \7486 , \349 );
and \U$7145 ( \7488 , \7482 , \7487 );
and \U$7146 ( \7489 , \7478 , \7487 );
or \U$7147 ( \7490 , \7483 , \7488 , \7489 );
and \U$7148 ( \7491 , \6297 , \406 );
and \U$7149 ( \7492 , \5954 , \404 );
nor \U$7150 ( \7493 , \7491 , \7492 );
xnor \U$7151 ( \7494 , \7493 , \413 );
and \U$7152 ( \7495 , \6802 , \422 );
and \U$7153 ( \7496 , \6499 , \420 );
nor \U$7154 ( \7497 , \7495 , \7496 );
xnor \U$7155 ( \7498 , \7497 , \429 );
and \U$7156 ( \7499 , \7494 , \7498 );
buf \U$7157 ( \7500 , RIbb2bfb0_117);
and \U$7158 ( \7501 , \7500 , \441 );
and \U$7159 ( \7502 , \6974 , \439 );
nor \U$7160 ( \7503 , \7501 , \7502 );
xnor \U$7161 ( \7504 , \7503 , \448 );
and \U$7162 ( \7505 , \7498 , \7504 );
and \U$7163 ( \7506 , \7494 , \7504 );
or \U$7164 ( \7507 , \7499 , \7505 , \7506 );
and \U$7165 ( \7508 , \7490 , \7507 );
and \U$7166 ( \7509 , \5045 , \357 );
and \U$7167 ( \7510 , \4576 , \355 );
nor \U$7168 ( \7511 , \7509 , \7510 );
xnor \U$7169 ( \7512 , \7511 , \364 );
and \U$7170 ( \7513 , \5314 , \373 );
and \U$7171 ( \7514 , \5050 , \371 );
nor \U$7172 ( \7515 , \7513 , \7514 );
xnor \U$7173 ( \7516 , \7515 , \380 );
and \U$7174 ( \7517 , \7512 , \7516 );
and \U$7175 ( \7518 , \5945 , \391 );
and \U$7176 ( \7519 , \5573 , \389 );
nor \U$7177 ( \7520 , \7518 , \7519 );
xnor \U$7178 ( \7521 , \7520 , \398 );
and \U$7179 ( \7522 , \7516 , \7521 );
and \U$7180 ( \7523 , \7512 , \7521 );
or \U$7181 ( \7524 , \7517 , \7522 , \7523 );
and \U$7182 ( \7525 , \7507 , \7524 );
and \U$7183 ( \7526 , \7490 , \7524 );
or \U$7184 ( \7527 , \7508 , \7525 , \7526 );
and \U$7185 ( \7528 , \408 , \6032 );
and \U$7186 ( \7529 , \385 , \6030 );
nor \U$7187 ( \7530 , \7528 , \7529 );
xnor \U$7188 ( \7531 , \7530 , \5692 );
and \U$7189 ( \7532 , \424 , \5443 );
and \U$7190 ( \7533 , \400 , \5441 );
nor \U$7191 ( \7534 , \7532 , \7533 );
xnor \U$7192 ( \7535 , \7534 , \5202 );
and \U$7193 ( \7536 , \7531 , \7535 );
and \U$7194 ( \7537 , \443 , \4977 );
and \U$7195 ( \7538 , \416 , \4975 );
nor \U$7196 ( \7539 , \7537 , \7538 );
xnor \U$7197 ( \7540 , \7539 , \4789 );
and \U$7198 ( \7541 , \7535 , \7540 );
and \U$7199 ( \7542 , \7531 , \7540 );
or \U$7200 ( \7543 , \7536 , \7541 , \7542 );
and \U$7201 ( \7544 , \450 , \4603 );
and \U$7202 ( \7545 , \435 , \4601 );
nor \U$7203 ( \7546 , \7544 , \7545 );
xnor \U$7204 ( \7547 , \7546 , \4371 );
and \U$7205 ( \7548 , \722 , \4152 );
and \U$7206 ( \7549 , \661 , \4150 );
nor \U$7207 ( \7550 , \7548 , \7549 );
xnor \U$7208 ( \7551 , \7550 , \4009 );
and \U$7209 ( \7552 , \7547 , \7551 );
and \U$7210 ( \7553 , \983 , \3829 );
and \U$7211 ( \7554 , \785 , \3827 );
nor \U$7212 ( \7555 , \7553 , \7554 );
xnor \U$7213 ( \7556 , \7555 , \3583 );
and \U$7214 ( \7557 , \7551 , \7556 );
and \U$7215 ( \7558 , \7547 , \7556 );
or \U$7216 ( \7559 , \7552 , \7557 , \7558 );
and \U$7217 ( \7560 , \7543 , \7559 );
xor \U$7218 ( \7561 , \6772 , \7311 );
xor \U$7219 ( \7562 , \7311 , \7312 );
not \U$7220 ( \7563 , \7562 );
and \U$7221 ( \7564 , \7561 , \7563 );
and \U$7222 ( \7565 , \359 , \7564 );
not \U$7223 ( \7566 , \7565 );
xnor \U$7224 ( \7567 , \7566 , \7315 );
and \U$7225 ( \7568 , \375 , \7035 );
and \U$7226 ( \7569 , \351 , \7033 );
nor \U$7227 ( \7570 , \7568 , \7569 );
xnor \U$7228 ( \7571 , \7570 , \6775 );
and \U$7229 ( \7572 , \7567 , \7571 );
and \U$7230 ( \7573 , \393 , \6541 );
and \U$7231 ( \7574 , \367 , \6539 );
nor \U$7232 ( \7575 , \7573 , \7574 );
xnor \U$7233 ( \7576 , \7575 , \6226 );
and \U$7234 ( \7577 , \7571 , \7576 );
and \U$7235 ( \7578 , \7567 , \7576 );
or \U$7236 ( \7579 , \7572 , \7577 , \7578 );
and \U$7237 ( \7580 , \7559 , \7579 );
and \U$7238 ( \7581 , \7543 , \7579 );
or \U$7239 ( \7582 , \7560 , \7580 , \7581 );
and \U$7240 ( \7583 , \7527 , \7582 );
and \U$7241 ( \7584 , \2637 , \1623 );
and \U$7242 ( \7585 , \2463 , \1621 );
nor \U$7243 ( \7586 , \7584 , \7585 );
xnor \U$7244 ( \7587 , \7586 , \1467 );
and \U$7245 ( \7588 , \2942 , \1351 );
and \U$7246 ( \7589 , \2804 , \1349 );
nor \U$7247 ( \7590 , \7588 , \7589 );
xnor \U$7248 ( \7591 , \7590 , \1238 );
and \U$7249 ( \7592 , \7587 , \7591 );
and \U$7250 ( \7593 , \3478 , \1157 );
and \U$7251 ( \7594 , \3061 , \1155 );
nor \U$7252 ( \7595 , \7593 , \7594 );
xnor \U$7253 ( \7596 , \7595 , \1021 );
and \U$7254 ( \7597 , \7591 , \7596 );
and \U$7255 ( \7598 , \7587 , \7596 );
or \U$7256 ( \7599 , \7592 , \7597 , \7598 );
and \U$7257 ( \7600 , \1176 , \3434 );
and \U$7258 ( \7601 , \1071 , \3432 );
nor \U$7259 ( \7602 , \7600 , \7601 );
xnor \U$7260 ( \7603 , \7602 , \3247 );
and \U$7261 ( \7604 , \1297 , \3121 );
and \U$7262 ( \7605 , \1181 , \3119 );
nor \U$7263 ( \7606 , \7604 , \7605 );
xnor \U$7264 ( \7607 , \7606 , \2916 );
and \U$7265 ( \7608 , \7603 , \7607 );
and \U$7266 ( \7609 , \1588 , \2715 );
and \U$7267 ( \7610 , \1412 , \2713 );
nor \U$7268 ( \7611 , \7609 , \7610 );
xnor \U$7269 ( \7612 , \7611 , \2566 );
and \U$7270 ( \7613 , \7607 , \7612 );
and \U$7271 ( \7614 , \7603 , \7612 );
or \U$7272 ( \7615 , \7608 , \7613 , \7614 );
and \U$7273 ( \7616 , \7599 , \7615 );
and \U$7274 ( \7617 , \1839 , \2393 );
and \U$7275 ( \7618 , \1596 , \2391 );
nor \U$7276 ( \7619 , \7617 , \7618 );
xnor \U$7277 ( \7620 , \7619 , \2251 );
and \U$7278 ( \7621 , \2030 , \2097 );
and \U$7279 ( \7622 , \1844 , \2095 );
nor \U$7280 ( \7623 , \7621 , \7622 );
xnor \U$7281 ( \7624 , \7623 , \1960 );
and \U$7282 ( \7625 , \7620 , \7624 );
and \U$7283 ( \7626 , \2438 , \1891 );
and \U$7284 ( \7627 , \2174 , \1889 );
nor \U$7285 ( \7628 , \7626 , \7627 );
xnor \U$7286 ( \7629 , \7628 , \1739 );
and \U$7287 ( \7630 , \7624 , \7629 );
and \U$7288 ( \7631 , \7620 , \7629 );
or \U$7289 ( \7632 , \7625 , \7630 , \7631 );
and \U$7290 ( \7633 , \7615 , \7632 );
and \U$7291 ( \7634 , \7599 , \7632 );
or \U$7292 ( \7635 , \7616 , \7633 , \7634 );
and \U$7293 ( \7636 , \7582 , \7635 );
and \U$7294 ( \7637 , \7527 , \7635 );
or \U$7295 ( \7638 , \7583 , \7636 , \7637 );
xor \U$7296 ( \7639 , \7298 , \7302 );
xor \U$7297 ( \7640 , \7639 , \7307 );
xor \U$7298 ( \7641 , \7262 , \7266 );
xor \U$7299 ( \7642 , \7641 , \7271 );
and \U$7300 ( \7643 , \7640 , \7642 );
xor \U$7301 ( \7644 , \7333 , \7337 );
xor \U$7302 ( \7645 , \7644 , \7342 );
and \U$7303 ( \7646 , \7642 , \7645 );
and \U$7304 ( \7647 , \7640 , \7645 );
or \U$7305 ( \7648 , \7643 , \7646 , \7647 );
and \U$7306 ( \7649 , \7500 , \436 );
xor \U$7307 ( \7650 , \7369 , \7373 );
xor \U$7308 ( \7651 , \7650 , \7378 );
and \U$7309 ( \7652 , \7649 , \7651 );
xor \U$7310 ( \7653 , \7386 , \7390 );
xor \U$7311 ( \7654 , \7653 , \7395 );
and \U$7312 ( \7655 , \7651 , \7654 );
and \U$7313 ( \7656 , \7649 , \7654 );
or \U$7314 ( \7657 , \7652 , \7655 , \7656 );
and \U$7315 ( \7658 , \7648 , \7657 );
xor \U$7316 ( \7659 , \7353 , \7357 );
xor \U$7317 ( \7660 , \7659 , \7362 );
xor \U$7318 ( \7661 , \7246 , \7250 );
xor \U$7319 ( \7662 , \7661 , \7255 );
and \U$7320 ( \7663 , \7660 , \7662 );
xor \U$7321 ( \7664 , \7279 , \7283 );
xor \U$7322 ( \7665 , \7664 , \7288 );
and \U$7323 ( \7666 , \7662 , \7665 );
and \U$7324 ( \7667 , \7660 , \7665 );
or \U$7325 ( \7668 , \7663 , \7666 , \7667 );
and \U$7326 ( \7669 , \7657 , \7668 );
and \U$7327 ( \7670 , \7648 , \7668 );
or \U$7328 ( \7671 , \7658 , \7669 , \7670 );
and \U$7329 ( \7672 , \7638 , \7671 );
xor \U$7330 ( \7673 , \7038 , \7042 );
xor \U$7331 ( \7674 , \7673 , \7047 );
xor \U$7332 ( \7675 , \7215 , \7217 );
xor \U$7333 ( \7676 , \7675 , \7220 );
and \U$7334 ( \7677 , \7674 , \7676 );
xor \U$7335 ( \7678 , \7225 , \7227 );
xor \U$7336 ( \7679 , \7678 , \7230 );
and \U$7337 ( \7680 , \7676 , \7679 );
and \U$7338 ( \7681 , \7674 , \7679 );
or \U$7339 ( \7682 , \7677 , \7680 , \7681 );
and \U$7340 ( \7683 , \7671 , \7682 );
and \U$7341 ( \7684 , \7638 , \7682 );
or \U$7342 ( \7685 , \7672 , \7683 , \7684 );
xor \U$7343 ( \7686 , \7258 , \7274 );
xor \U$7344 ( \7687 , \7686 , \7291 );
xor \U$7345 ( \7688 , \7365 , \7381 );
xor \U$7346 ( \7689 , \7688 , \7398 );
and \U$7347 ( \7690 , \7687 , \7689 );
xnor \U$7348 ( \7691 , \7236 , \7238 );
and \U$7349 ( \7692 , \7689 , \7691 );
and \U$7350 ( \7693 , \7687 , \7691 );
or \U$7351 ( \7694 , \7690 , \7692 , \7693 );
xor \U$7352 ( \7695 , \7420 , \7422 );
xor \U$7353 ( \7696 , \7695 , \7425 );
and \U$7354 ( \7697 , \7694 , \7696 );
xor \U$7355 ( \7698 , \7407 , \7409 );
xor \U$7356 ( \7699 , \7698 , \7412 );
and \U$7357 ( \7700 , \7696 , \7699 );
and \U$7358 ( \7701 , \7694 , \7699 );
or \U$7359 ( \7702 , \7697 , \7700 , \7701 );
and \U$7360 ( \7703 , \7685 , \7702 );
xor \U$7361 ( \7704 , \7223 , \7233 );
xor \U$7362 ( \7705 , \7704 , \7239 );
xor \U$7363 ( \7706 , \7294 , \7348 );
xor \U$7364 ( \7707 , \7706 , \7401 );
and \U$7365 ( \7708 , \7705 , \7707 );
and \U$7366 ( \7709 , \7702 , \7708 );
and \U$7367 ( \7710 , \7685 , \7708 );
or \U$7368 ( \7711 , \7703 , \7709 , \7710 );
xor \U$7369 ( \7712 , \7242 , \7404 );
xor \U$7370 ( \7713 , \7712 , \7415 );
xor \U$7371 ( \7714 , \7428 , \7430 );
xor \U$7372 ( \7715 , \7714 , \7433 );
and \U$7373 ( \7716 , \7713 , \7715 );
xor \U$7374 ( \7717 , \7439 , \7441 );
and \U$7375 ( \7718 , \7715 , \7717 );
and \U$7376 ( \7719 , \7713 , \7717 );
or \U$7377 ( \7720 , \7716 , \7718 , \7719 );
and \U$7378 ( \7721 , \7711 , \7720 );
xor \U$7379 ( \7722 , \7447 , \7449 );
xor \U$7380 ( \7723 , \7722 , \7451 );
and \U$7381 ( \7724 , \7720 , \7723 );
and \U$7382 ( \7725 , \7711 , \7723 );
or \U$7383 ( \7726 , \7721 , \7724 , \7725 );
xor \U$7384 ( \7727 , \7157 , \7175 );
xor \U$7385 ( \7728 , \7727 , \7181 );
and \U$7386 ( \7729 , \7726 , \7728 );
xor \U$7387 ( \7730 , \7445 , \7454 );
xor \U$7388 ( \7731 , \7730 , \7457 );
and \U$7389 ( \7732 , \7728 , \7731 );
and \U$7390 ( \7733 , \7726 , \7731 );
or \U$7391 ( \7734 , \7729 , \7732 , \7733 );
xor \U$7392 ( \7735 , \7460 , \7462 );
xor \U$7393 ( \7736 , \7735 , \7465 );
and \U$7394 ( \7737 , \7734 , \7736 );
and \U$7395 ( \7738 , \7474 , \7737 );
xor \U$7396 ( \7739 , \7474 , \7737 );
xor \U$7397 ( \7740 , \7734 , \7736 );
and \U$7398 ( \7741 , \2463 , \1891 );
and \U$7399 ( \7742 , \2438 , \1889 );
nor \U$7400 ( \7743 , \7741 , \7742 );
xnor \U$7401 ( \7744 , \7743 , \1739 );
and \U$7402 ( \7745 , \2804 , \1623 );
and \U$7403 ( \7746 , \2637 , \1621 );
nor \U$7404 ( \7747 , \7745 , \7746 );
xnor \U$7405 ( \7748 , \7747 , \1467 );
and \U$7406 ( \7749 , \7744 , \7748 );
and \U$7407 ( \7750 , \3061 , \1351 );
and \U$7408 ( \7751 , \2942 , \1349 );
nor \U$7409 ( \7752 , \7750 , \7751 );
xnor \U$7410 ( \7753 , \7752 , \1238 );
and \U$7411 ( \7754 , \7748 , \7753 );
and \U$7412 ( \7755 , \7744 , \7753 );
or \U$7413 ( \7756 , \7749 , \7754 , \7755 );
and \U$7414 ( \7757 , \1071 , \3829 );
and \U$7415 ( \7758 , \983 , \3827 );
nor \U$7416 ( \7759 , \7757 , \7758 );
xnor \U$7417 ( \7760 , \7759 , \3583 );
and \U$7418 ( \7761 , \1181 , \3434 );
and \U$7419 ( \7762 , \1176 , \3432 );
nor \U$7420 ( \7763 , \7761 , \7762 );
xnor \U$7421 ( \7764 , \7763 , \3247 );
and \U$7422 ( \7765 , \7760 , \7764 );
and \U$7423 ( \7766 , \1412 , \3121 );
and \U$7424 ( \7767 , \1297 , \3119 );
nor \U$7425 ( \7768 , \7766 , \7767 );
xnor \U$7426 ( \7769 , \7768 , \2916 );
and \U$7427 ( \7770 , \7764 , \7769 );
and \U$7428 ( \7771 , \7760 , \7769 );
or \U$7429 ( \7772 , \7765 , \7770 , \7771 );
and \U$7430 ( \7773 , \7756 , \7772 );
and \U$7431 ( \7774 , \1596 , \2715 );
and \U$7432 ( \7775 , \1588 , \2713 );
nor \U$7433 ( \7776 , \7774 , \7775 );
xnor \U$7434 ( \7777 , \7776 , \2566 );
and \U$7435 ( \7778 , \1844 , \2393 );
and \U$7436 ( \7779 , \1839 , \2391 );
nor \U$7437 ( \7780 , \7778 , \7779 );
xnor \U$7438 ( \7781 , \7780 , \2251 );
and \U$7439 ( \7782 , \7777 , \7781 );
and \U$7440 ( \7783 , \2174 , \2097 );
and \U$7441 ( \7784 , \2030 , \2095 );
nor \U$7442 ( \7785 , \7783 , \7784 );
xnor \U$7443 ( \7786 , \7785 , \1960 );
and \U$7444 ( \7787 , \7781 , \7786 );
and \U$7445 ( \7788 , \7777 , \7786 );
or \U$7446 ( \7789 , \7782 , \7787 , \7788 );
and \U$7447 ( \7790 , \7772 , \7789 );
and \U$7448 ( \7791 , \7756 , \7789 );
or \U$7449 ( \7792 , \7773 , \7790 , \7791 );
and \U$7450 ( \7793 , \435 , \4977 );
and \U$7451 ( \7794 , \443 , \4975 );
nor \U$7452 ( \7795 , \7793 , \7794 );
xnor \U$7453 ( \7796 , \7795 , \4789 );
and \U$7454 ( \7797 , \661 , \4603 );
and \U$7455 ( \7798 , \450 , \4601 );
nor \U$7456 ( \7799 , \7797 , \7798 );
xnor \U$7457 ( \7800 , \7799 , \4371 );
and \U$7458 ( \7801 , \7796 , \7800 );
and \U$7459 ( \7802 , \785 , \4152 );
and \U$7460 ( \7803 , \722 , \4150 );
nor \U$7461 ( \7804 , \7802 , \7803 );
xnor \U$7462 ( \7805 , \7804 , \4009 );
and \U$7463 ( \7806 , \7800 , \7805 );
and \U$7464 ( \7807 , \7796 , \7805 );
or \U$7465 ( \7808 , \7801 , \7806 , \7807 );
buf \U$7466 ( \7809 , RIbb2dc48_56);
buf \U$7467 ( \7810 , RIbb2dbd0_57);
and \U$7468 ( \7811 , \7809 , \7810 );
not \U$7469 ( \7812 , \7811 );
and \U$7470 ( \7813 , \7312 , \7812 );
not \U$7471 ( \7814 , \7813 );
and \U$7472 ( \7815 , \351 , \7564 );
and \U$7473 ( \7816 , \359 , \7562 );
nor \U$7474 ( \7817 , \7815 , \7816 );
xnor \U$7475 ( \7818 , \7817 , \7315 );
and \U$7476 ( \7819 , \7814 , \7818 );
and \U$7477 ( \7820 , \367 , \7035 );
and \U$7478 ( \7821 , \375 , \7033 );
nor \U$7479 ( \7822 , \7820 , \7821 );
xnor \U$7480 ( \7823 , \7822 , \6775 );
and \U$7481 ( \7824 , \7818 , \7823 );
and \U$7482 ( \7825 , \7814 , \7823 );
or \U$7483 ( \7826 , \7819 , \7824 , \7825 );
and \U$7484 ( \7827 , \7808 , \7826 );
and \U$7485 ( \7828 , \385 , \6541 );
and \U$7486 ( \7829 , \393 , \6539 );
nor \U$7487 ( \7830 , \7828 , \7829 );
xnor \U$7488 ( \7831 , \7830 , \6226 );
and \U$7489 ( \7832 , \400 , \6032 );
and \U$7490 ( \7833 , \408 , \6030 );
nor \U$7491 ( \7834 , \7832 , \7833 );
xnor \U$7492 ( \7835 , \7834 , \5692 );
and \U$7493 ( \7836 , \7831 , \7835 );
and \U$7494 ( \7837 , \416 , \5443 );
and \U$7495 ( \7838 , \424 , \5441 );
nor \U$7496 ( \7839 , \7837 , \7838 );
xnor \U$7497 ( \7840 , \7839 , \5202 );
and \U$7498 ( \7841 , \7835 , \7840 );
and \U$7499 ( \7842 , \7831 , \7840 );
or \U$7500 ( \7843 , \7836 , \7841 , \7842 );
and \U$7501 ( \7844 , \7826 , \7843 );
and \U$7502 ( \7845 , \7808 , \7843 );
or \U$7503 ( \7846 , \7827 , \7844 , \7845 );
and \U$7504 ( \7847 , \7792 , \7846 );
and \U$7505 ( \7848 , \4576 , \624 );
and \U$7506 ( \7849 , \4568 , \622 );
nor \U$7507 ( \7850 , \7848 , \7849 );
xnor \U$7508 ( \7851 , \7850 , \349 );
and \U$7509 ( \7852 , \5050 , \357 );
and \U$7510 ( \7853 , \5045 , \355 );
nor \U$7511 ( \7854 , \7852 , \7853 );
xnor \U$7512 ( \7855 , \7854 , \364 );
and \U$7513 ( \7856 , \7851 , \7855 );
and \U$7514 ( \7857 , \5573 , \373 );
and \U$7515 ( \7858 , \5314 , \371 );
nor \U$7516 ( \7859 , \7857 , \7858 );
xnor \U$7517 ( \7860 , \7859 , \380 );
and \U$7518 ( \7861 , \7855 , \7860 );
and \U$7519 ( \7862 , \7851 , \7860 );
or \U$7520 ( \7863 , \7856 , \7861 , \7862 );
and \U$7521 ( \7864 , \5954 , \391 );
and \U$7522 ( \7865 , \5945 , \389 );
nor \U$7523 ( \7866 , \7864 , \7865 );
xnor \U$7524 ( \7867 , \7866 , \398 );
and \U$7525 ( \7868 , \6499 , \406 );
and \U$7526 ( \7869 , \6297 , \404 );
nor \U$7527 ( \7870 , \7868 , \7869 );
xnor \U$7528 ( \7871 , \7870 , \413 );
and \U$7529 ( \7872 , \7867 , \7871 );
and \U$7530 ( \7873 , \6974 , \422 );
and \U$7531 ( \7874 , \6802 , \420 );
nor \U$7532 ( \7875 , \7873 , \7874 );
xnor \U$7533 ( \7876 , \7875 , \429 );
and \U$7534 ( \7877 , \7871 , \7876 );
and \U$7535 ( \7878 , \7867 , \7876 );
or \U$7536 ( \7879 , \7872 , \7877 , \7878 );
and \U$7537 ( \7880 , \7863 , \7879 );
and \U$7538 ( \7881 , \3686 , \1157 );
and \U$7539 ( \7882 , \3478 , \1155 );
nor \U$7540 ( \7883 , \7881 , \7882 );
xnor \U$7541 ( \7884 , \7883 , \1021 );
and \U$7542 ( \7885 , \3813 , \957 );
and \U$7543 ( \7886 , \3808 , \955 );
nor \U$7544 ( \7887 , \7885 , \7886 );
xnor \U$7545 ( \7888 , \7887 , \879 );
and \U$7546 ( \7889 , \7884 , \7888 );
and \U$7547 ( \7890 , \4266 , \793 );
and \U$7548 ( \7891 , \4069 , \791 );
nor \U$7549 ( \7892 , \7890 , \7891 );
xnor \U$7550 ( \7893 , \7892 , \699 );
and \U$7551 ( \7894 , \7888 , \7893 );
and \U$7552 ( \7895 , \7884 , \7893 );
or \U$7553 ( \7896 , \7889 , \7894 , \7895 );
and \U$7554 ( \7897 , \7879 , \7896 );
and \U$7555 ( \7898 , \7863 , \7896 );
or \U$7556 ( \7899 , \7880 , \7897 , \7898 );
and \U$7557 ( \7900 , \7846 , \7899 );
and \U$7558 ( \7901 , \7792 , \7899 );
or \U$7559 ( \7902 , \7847 , \7900 , \7901 );
xor \U$7560 ( \7903 , \7478 , \7482 );
xor \U$7561 ( \7904 , \7903 , \7487 );
xor \U$7562 ( \7905 , \7587 , \7591 );
xor \U$7563 ( \7906 , \7905 , \7596 );
and \U$7564 ( \7907 , \7904 , \7906 );
xor \U$7565 ( \7908 , \7512 , \7516 );
xor \U$7566 ( \7909 , \7908 , \7521 );
and \U$7567 ( \7910 , \7906 , \7909 );
and \U$7568 ( \7911 , \7904 , \7909 );
or \U$7569 ( \7912 , \7907 , \7910 , \7911 );
xor \U$7570 ( \7913 , \7547 , \7551 );
xor \U$7571 ( \7914 , \7913 , \7556 );
xor \U$7572 ( \7915 , \7603 , \7607 );
xor \U$7573 ( \7916 , \7915 , \7612 );
and \U$7574 ( \7917 , \7914 , \7916 );
xor \U$7575 ( \7918 , \7620 , \7624 );
xor \U$7576 ( \7919 , \7918 , \7629 );
and \U$7577 ( \7920 , \7916 , \7919 );
and \U$7578 ( \7921 , \7914 , \7919 );
or \U$7579 ( \7922 , \7917 , \7920 , \7921 );
and \U$7580 ( \7923 , \7912 , \7922 );
buf \U$7581 ( \7924 , RIbb2bf38_118);
and \U$7582 ( \7925 , \7924 , \436 );
xor \U$7583 ( \7926 , \7494 , \7498 );
xor \U$7584 ( \7927 , \7926 , \7504 );
or \U$7585 ( \7928 , \7925 , \7927 );
and \U$7586 ( \7929 , \7922 , \7928 );
and \U$7587 ( \7930 , \7912 , \7928 );
or \U$7588 ( \7931 , \7923 , \7929 , \7930 );
and \U$7589 ( \7932 , \7902 , \7931 );
xor \U$7590 ( \7933 , \7316 , \7320 );
xor \U$7591 ( \7934 , \7933 , \7325 );
xor \U$7592 ( \7935 , \7640 , \7642 );
xor \U$7593 ( \7936 , \7935 , \7645 );
and \U$7594 ( \7937 , \7934 , \7936 );
xor \U$7595 ( \7938 , \7660 , \7662 );
xor \U$7596 ( \7939 , \7938 , \7665 );
and \U$7597 ( \7940 , \7936 , \7939 );
and \U$7598 ( \7941 , \7934 , \7939 );
or \U$7599 ( \7942 , \7937 , \7940 , \7941 );
and \U$7600 ( \7943 , \7931 , \7942 );
and \U$7601 ( \7944 , \7902 , \7942 );
or \U$7602 ( \7945 , \7932 , \7943 , \7944 );
xor \U$7603 ( \7946 , \7527 , \7582 );
xor \U$7604 ( \7947 , \7946 , \7635 );
xor \U$7605 ( \7948 , \7648 , \7657 );
xor \U$7606 ( \7949 , \7948 , \7668 );
and \U$7607 ( \7950 , \7947 , \7949 );
xor \U$7608 ( \7951 , \7674 , \7676 );
xor \U$7609 ( \7952 , \7951 , \7679 );
and \U$7610 ( \7953 , \7949 , \7952 );
and \U$7611 ( \7954 , \7947 , \7952 );
or \U$7612 ( \7955 , \7950 , \7953 , \7954 );
and \U$7613 ( \7956 , \7945 , \7955 );
xor \U$7614 ( \7957 , \7490 , \7507 );
xor \U$7615 ( \7958 , \7957 , \7524 );
xor \U$7616 ( \7959 , \7599 , \7615 );
xor \U$7617 ( \7960 , \7959 , \7632 );
and \U$7618 ( \7961 , \7958 , \7960 );
xor \U$7619 ( \7962 , \7649 , \7651 );
xor \U$7620 ( \7963 , \7962 , \7654 );
and \U$7621 ( \7964 , \7960 , \7963 );
and \U$7622 ( \7965 , \7958 , \7963 );
or \U$7623 ( \7966 , \7961 , \7964 , \7965 );
xor \U$7624 ( \7967 , \7310 , \7328 );
xor \U$7625 ( \7968 , \7967 , \7345 );
and \U$7626 ( \7969 , \7966 , \7968 );
xor \U$7627 ( \7970 , \7687 , \7689 );
xor \U$7628 ( \7971 , \7970 , \7691 );
and \U$7629 ( \7972 , \7968 , \7971 );
and \U$7630 ( \7973 , \7966 , \7971 );
or \U$7631 ( \7974 , \7969 , \7972 , \7973 );
and \U$7632 ( \7975 , \7955 , \7974 );
and \U$7633 ( \7976 , \7945 , \7974 );
or \U$7634 ( \7977 , \7956 , \7975 , \7976 );
xor \U$7635 ( \7978 , \7638 , \7671 );
xor \U$7636 ( \7979 , \7978 , \7682 );
xor \U$7637 ( \7980 , \7694 , \7696 );
xor \U$7638 ( \7981 , \7980 , \7699 );
and \U$7639 ( \7982 , \7979 , \7981 );
xor \U$7640 ( \7983 , \7705 , \7707 );
and \U$7641 ( \7984 , \7981 , \7983 );
and \U$7642 ( \7985 , \7979 , \7983 );
or \U$7643 ( \7986 , \7982 , \7984 , \7985 );
and \U$7644 ( \7987 , \7977 , \7986 );
xor \U$7645 ( \7988 , \7713 , \7715 );
xor \U$7646 ( \7989 , \7988 , \7717 );
and \U$7647 ( \7990 , \7986 , \7989 );
and \U$7648 ( \7991 , \7977 , \7989 );
or \U$7649 ( \7992 , \7987 , \7990 , \7991 );
xor \U$7650 ( \7993 , \7418 , \7436 );
xor \U$7651 ( \7994 , \7993 , \7442 );
and \U$7652 ( \7995 , \7992 , \7994 );
xor \U$7653 ( \7996 , \7711 , \7720 );
xor \U$7654 ( \7997 , \7996 , \7723 );
and \U$7655 ( \7998 , \7994 , \7997 );
and \U$7656 ( \7999 , \7992 , \7997 );
or \U$7657 ( \8000 , \7995 , \7998 , \7999 );
xor \U$7658 ( \8001 , \7726 , \7728 );
xor \U$7659 ( \8002 , \8001 , \7731 );
and \U$7660 ( \8003 , \8000 , \8002 );
and \U$7661 ( \8004 , \7740 , \8003 );
xor \U$7662 ( \8005 , \7740 , \8003 );
xor \U$7663 ( \8006 , \8000 , \8002 );
and \U$7664 ( \8007 , \1839 , \2715 );
and \U$7665 ( \8008 , \1596 , \2713 );
nor \U$7666 ( \8009 , \8007 , \8008 );
xnor \U$7667 ( \8010 , \8009 , \2566 );
and \U$7668 ( \8011 , \2030 , \2393 );
and \U$7669 ( \8012 , \1844 , \2391 );
nor \U$7670 ( \8013 , \8011 , \8012 );
xnor \U$7671 ( \8014 , \8013 , \2251 );
and \U$7672 ( \8015 , \8010 , \8014 );
and \U$7673 ( \8016 , \2438 , \2097 );
and \U$7674 ( \8017 , \2174 , \2095 );
nor \U$7675 ( \8018 , \8016 , \8017 );
xnor \U$7676 ( \8019 , \8018 , \1960 );
and \U$7677 ( \8020 , \8014 , \8019 );
and \U$7678 ( \8021 , \8010 , \8019 );
or \U$7679 ( \8022 , \8015 , \8020 , \8021 );
and \U$7680 ( \8023 , \2637 , \1891 );
and \U$7681 ( \8024 , \2463 , \1889 );
nor \U$7682 ( \8025 , \8023 , \8024 );
xnor \U$7683 ( \8026 , \8025 , \1739 );
and \U$7684 ( \8027 , \2942 , \1623 );
and \U$7685 ( \8028 , \2804 , \1621 );
nor \U$7686 ( \8029 , \8027 , \8028 );
xnor \U$7687 ( \8030 , \8029 , \1467 );
and \U$7688 ( \8031 , \8026 , \8030 );
and \U$7689 ( \8032 , \3478 , \1351 );
and \U$7690 ( \8033 , \3061 , \1349 );
nor \U$7691 ( \8034 , \8032 , \8033 );
xnor \U$7692 ( \8035 , \8034 , \1238 );
and \U$7693 ( \8036 , \8030 , \8035 );
and \U$7694 ( \8037 , \8026 , \8035 );
or \U$7695 ( \8038 , \8031 , \8036 , \8037 );
and \U$7696 ( \8039 , \8022 , \8038 );
and \U$7697 ( \8040 , \1176 , \3829 );
and \U$7698 ( \8041 , \1071 , \3827 );
nor \U$7699 ( \8042 , \8040 , \8041 );
xnor \U$7700 ( \8043 , \8042 , \3583 );
and \U$7701 ( \8044 , \1297 , \3434 );
and \U$7702 ( \8045 , \1181 , \3432 );
nor \U$7703 ( \8046 , \8044 , \8045 );
xnor \U$7704 ( \8047 , \8046 , \3247 );
and \U$7705 ( \8048 , \8043 , \8047 );
and \U$7706 ( \8049 , \1588 , \3121 );
and \U$7707 ( \8050 , \1412 , \3119 );
nor \U$7708 ( \8051 , \8049 , \8050 );
xnor \U$7709 ( \8052 , \8051 , \2916 );
and \U$7710 ( \8053 , \8047 , \8052 );
and \U$7711 ( \8054 , \8043 , \8052 );
or \U$7712 ( \8055 , \8048 , \8053 , \8054 );
and \U$7713 ( \8056 , \8038 , \8055 );
and \U$7714 ( \8057 , \8022 , \8055 );
or \U$7715 ( \8058 , \8039 , \8056 , \8057 );
and \U$7716 ( \8059 , \5045 , \624 );
and \U$7717 ( \8060 , \4576 , \622 );
nor \U$7718 ( \8061 , \8059 , \8060 );
xnor \U$7719 ( \8062 , \8061 , \349 );
and \U$7720 ( \8063 , \5314 , \357 );
and \U$7721 ( \8064 , \5050 , \355 );
nor \U$7722 ( \8065 , \8063 , \8064 );
xnor \U$7723 ( \8066 , \8065 , \364 );
and \U$7724 ( \8067 , \8062 , \8066 );
and \U$7725 ( \8068 , \5945 , \373 );
and \U$7726 ( \8069 , \5573 , \371 );
nor \U$7727 ( \8070 , \8068 , \8069 );
xnor \U$7728 ( \8071 , \8070 , \380 );
and \U$7729 ( \8072 , \8066 , \8071 );
and \U$7730 ( \8073 , \8062 , \8071 );
or \U$7731 ( \8074 , \8067 , \8072 , \8073 );
and \U$7732 ( \8075 , \3808 , \1157 );
and \U$7733 ( \8076 , \3686 , \1155 );
nor \U$7734 ( \8077 , \8075 , \8076 );
xnor \U$7735 ( \8078 , \8077 , \1021 );
and \U$7736 ( \8079 , \4069 , \957 );
and \U$7737 ( \8080 , \3813 , \955 );
nor \U$7738 ( \8081 , \8079 , \8080 );
xnor \U$7739 ( \8082 , \8081 , \879 );
and \U$7740 ( \8083 , \8078 , \8082 );
and \U$7741 ( \8084 , \4568 , \793 );
and \U$7742 ( \8085 , \4266 , \791 );
nor \U$7743 ( \8086 , \8084 , \8085 );
xnor \U$7744 ( \8087 , \8086 , \699 );
and \U$7745 ( \8088 , \8082 , \8087 );
and \U$7746 ( \8089 , \8078 , \8087 );
or \U$7747 ( \8090 , \8083 , \8088 , \8089 );
and \U$7748 ( \8091 , \8074 , \8090 );
and \U$7749 ( \8092 , \6297 , \391 );
and \U$7750 ( \8093 , \5954 , \389 );
nor \U$7751 ( \8094 , \8092 , \8093 );
xnor \U$7752 ( \8095 , \8094 , \398 );
and \U$7753 ( \8096 , \6802 , \406 );
and \U$7754 ( \8097 , \6499 , \404 );
nor \U$7755 ( \8098 , \8096 , \8097 );
xnor \U$7756 ( \8099 , \8098 , \413 );
and \U$7757 ( \8100 , \8095 , \8099 );
and \U$7758 ( \8101 , \7500 , \422 );
and \U$7759 ( \8102 , \6974 , \420 );
nor \U$7760 ( \8103 , \8101 , \8102 );
xnor \U$7761 ( \8104 , \8103 , \429 );
and \U$7762 ( \8105 , \8099 , \8104 );
and \U$7763 ( \8106 , \8095 , \8104 );
or \U$7764 ( \8107 , \8100 , \8105 , \8106 );
and \U$7765 ( \8108 , \8090 , \8107 );
and \U$7766 ( \8109 , \8074 , \8107 );
or \U$7767 ( \8110 , \8091 , \8108 , \8109 );
and \U$7768 ( \8111 , \8058 , \8110 );
and \U$7769 ( \8112 , \450 , \4977 );
and \U$7770 ( \8113 , \435 , \4975 );
nor \U$7771 ( \8114 , \8112 , \8113 );
xnor \U$7772 ( \8115 , \8114 , \4789 );
and \U$7773 ( \8116 , \722 , \4603 );
and \U$7774 ( \8117 , \661 , \4601 );
nor \U$7775 ( \8118 , \8116 , \8117 );
xnor \U$7776 ( \8119 , \8118 , \4371 );
and \U$7777 ( \8120 , \8115 , \8119 );
and \U$7778 ( \8121 , \983 , \4152 );
and \U$7779 ( \8122 , \785 , \4150 );
nor \U$7780 ( \8123 , \8121 , \8122 );
xnor \U$7781 ( \8124 , \8123 , \4009 );
and \U$7782 ( \8125 , \8119 , \8124 );
and \U$7783 ( \8126 , \8115 , \8124 );
or \U$7784 ( \8127 , \8120 , \8125 , \8126 );
xor \U$7785 ( \8128 , \7312 , \7809 );
xor \U$7786 ( \8129 , \7809 , \7810 );
not \U$7787 ( \8130 , \8129 );
and \U$7788 ( \8131 , \8128 , \8130 );
and \U$7789 ( \8132 , \359 , \8131 );
not \U$7790 ( \8133 , \8132 );
xnor \U$7791 ( \8134 , \8133 , \7813 );
and \U$7792 ( \8135 , \375 , \7564 );
and \U$7793 ( \8136 , \351 , \7562 );
nor \U$7794 ( \8137 , \8135 , \8136 );
xnor \U$7795 ( \8138 , \8137 , \7315 );
and \U$7796 ( \8139 , \8134 , \8138 );
and \U$7797 ( \8140 , \393 , \7035 );
and \U$7798 ( \8141 , \367 , \7033 );
nor \U$7799 ( \8142 , \8140 , \8141 );
xnor \U$7800 ( \8143 , \8142 , \6775 );
and \U$7801 ( \8144 , \8138 , \8143 );
and \U$7802 ( \8145 , \8134 , \8143 );
or \U$7803 ( \8146 , \8139 , \8144 , \8145 );
and \U$7804 ( \8147 , \8127 , \8146 );
and \U$7805 ( \8148 , \408 , \6541 );
and \U$7806 ( \8149 , \385 , \6539 );
nor \U$7807 ( \8150 , \8148 , \8149 );
xnor \U$7808 ( \8151 , \8150 , \6226 );
and \U$7809 ( \8152 , \424 , \6032 );
and \U$7810 ( \8153 , \400 , \6030 );
nor \U$7811 ( \8154 , \8152 , \8153 );
xnor \U$7812 ( \8155 , \8154 , \5692 );
and \U$7813 ( \8156 , \8151 , \8155 );
and \U$7814 ( \8157 , \443 , \5443 );
and \U$7815 ( \8158 , \416 , \5441 );
nor \U$7816 ( \8159 , \8157 , \8158 );
xnor \U$7817 ( \8160 , \8159 , \5202 );
and \U$7818 ( \8161 , \8155 , \8160 );
and \U$7819 ( \8162 , \8151 , \8160 );
or \U$7820 ( \8163 , \8156 , \8161 , \8162 );
and \U$7821 ( \8164 , \8146 , \8163 );
and \U$7822 ( \8165 , \8127 , \8163 );
or \U$7823 ( \8166 , \8147 , \8164 , \8165 );
and \U$7824 ( \8167 , \8110 , \8166 );
and \U$7825 ( \8168 , \8058 , \8166 );
or \U$7826 ( \8169 , \8111 , \8167 , \8168 );
buf \U$7827 ( \8170 , RIbb2bec0_119);
and \U$7828 ( \8171 , \8170 , \441 );
and \U$7829 ( \8172 , \7924 , \439 );
nor \U$7830 ( \8173 , \8171 , \8172 );
xnor \U$7831 ( \8174 , \8173 , \448 );
buf \U$7832 ( \8175 , RIbb2be48_120);
and \U$7833 ( \8176 , \8175 , \436 );
or \U$7834 ( \8177 , \8174 , \8176 );
and \U$7835 ( \8178 , \7924 , \441 );
and \U$7836 ( \8179 , \7500 , \439 );
nor \U$7837 ( \8180 , \8178 , \8179 );
xnor \U$7838 ( \8181 , \8180 , \448 );
and \U$7839 ( \8182 , \8177 , \8181 );
and \U$7840 ( \8183 , \8170 , \436 );
and \U$7841 ( \8184 , \8181 , \8183 );
and \U$7842 ( \8185 , \8177 , \8183 );
or \U$7843 ( \8186 , \8182 , \8184 , \8185 );
xor \U$7844 ( \8187 , \7851 , \7855 );
xor \U$7845 ( \8188 , \8187 , \7860 );
xor \U$7846 ( \8189 , \7867 , \7871 );
xor \U$7847 ( \8190 , \8189 , \7876 );
and \U$7848 ( \8191 , \8188 , \8190 );
xor \U$7849 ( \8192 , \7884 , \7888 );
xor \U$7850 ( \8193 , \8192 , \7893 );
and \U$7851 ( \8194 , \8190 , \8193 );
and \U$7852 ( \8195 , \8188 , \8193 );
or \U$7853 ( \8196 , \8191 , \8194 , \8195 );
and \U$7854 ( \8197 , \8186 , \8196 );
xor \U$7855 ( \8198 , \7744 , \7748 );
xor \U$7856 ( \8199 , \8198 , \7753 );
xor \U$7857 ( \8200 , \7760 , \7764 );
xor \U$7858 ( \8201 , \8200 , \7769 );
and \U$7859 ( \8202 , \8199 , \8201 );
xor \U$7860 ( \8203 , \7777 , \7781 );
xor \U$7861 ( \8204 , \8203 , \7786 );
and \U$7862 ( \8205 , \8201 , \8204 );
and \U$7863 ( \8206 , \8199 , \8204 );
or \U$7864 ( \8207 , \8202 , \8205 , \8206 );
and \U$7865 ( \8208 , \8196 , \8207 );
and \U$7866 ( \8209 , \8186 , \8207 );
or \U$7867 ( \8210 , \8197 , \8208 , \8209 );
and \U$7868 ( \8211 , \8169 , \8210 );
xor \U$7869 ( \8212 , \7796 , \7800 );
xor \U$7870 ( \8213 , \8212 , \7805 );
xor \U$7871 ( \8214 , \7814 , \7818 );
xor \U$7872 ( \8215 , \8214 , \7823 );
and \U$7873 ( \8216 , \8213 , \8215 );
xor \U$7874 ( \8217 , \7831 , \7835 );
xor \U$7875 ( \8218 , \8217 , \7840 );
and \U$7876 ( \8219 , \8215 , \8218 );
and \U$7877 ( \8220 , \8213 , \8218 );
or \U$7878 ( \8221 , \8216 , \8219 , \8220 );
xor \U$7879 ( \8222 , \7531 , \7535 );
xor \U$7880 ( \8223 , \8222 , \7540 );
and \U$7881 ( \8224 , \8221 , \8223 );
xor \U$7882 ( \8225 , \7567 , \7571 );
xor \U$7883 ( \8226 , \8225 , \7576 );
and \U$7884 ( \8227 , \8223 , \8226 );
and \U$7885 ( \8228 , \8221 , \8226 );
or \U$7886 ( \8229 , \8224 , \8227 , \8228 );
and \U$7887 ( \8230 , \8210 , \8229 );
and \U$7888 ( \8231 , \8169 , \8229 );
or \U$7889 ( \8232 , \8211 , \8230 , \8231 );
xor \U$7890 ( \8233 , \7756 , \7772 );
xor \U$7891 ( \8234 , \8233 , \7789 );
xor \U$7892 ( \8235 , \7808 , \7826 );
xor \U$7893 ( \8236 , \8235 , \7843 );
and \U$7894 ( \8237 , \8234 , \8236 );
xor \U$7895 ( \8238 , \7863 , \7879 );
xor \U$7896 ( \8239 , \8238 , \7896 );
and \U$7897 ( \8240 , \8236 , \8239 );
and \U$7898 ( \8241 , \8234 , \8239 );
or \U$7899 ( \8242 , \8237 , \8240 , \8241 );
xor \U$7900 ( \8243 , \7904 , \7906 );
xor \U$7901 ( \8244 , \8243 , \7909 );
xor \U$7902 ( \8245 , \7914 , \7916 );
xor \U$7903 ( \8246 , \8245 , \7919 );
and \U$7904 ( \8247 , \8244 , \8246 );
xnor \U$7905 ( \8248 , \7925 , \7927 );
and \U$7906 ( \8249 , \8246 , \8248 );
and \U$7907 ( \8250 , \8244 , \8248 );
or \U$7908 ( \8251 , \8247 , \8249 , \8250 );
and \U$7909 ( \8252 , \8242 , \8251 );
xor \U$7910 ( \8253 , \7543 , \7559 );
xor \U$7911 ( \8254 , \8253 , \7579 );
and \U$7912 ( \8255 , \8251 , \8254 );
and \U$7913 ( \8256 , \8242 , \8254 );
or \U$7914 ( \8257 , \8252 , \8255 , \8256 );
and \U$7915 ( \8258 , \8232 , \8257 );
xor \U$7916 ( \8259 , \7912 , \7922 );
xor \U$7917 ( \8260 , \8259 , \7928 );
xor \U$7918 ( \8261 , \7958 , \7960 );
xor \U$7919 ( \8262 , \8261 , \7963 );
and \U$7920 ( \8263 , \8260 , \8262 );
xor \U$7921 ( \8264 , \7934 , \7936 );
xor \U$7922 ( \8265 , \8264 , \7939 );
and \U$7923 ( \8266 , \8262 , \8265 );
and \U$7924 ( \8267 , \8260 , \8265 );
or \U$7925 ( \8268 , \8263 , \8266 , \8267 );
and \U$7926 ( \8269 , \8257 , \8268 );
and \U$7927 ( \8270 , \8232 , \8268 );
or \U$7928 ( \8271 , \8258 , \8269 , \8270 );
xor \U$7929 ( \8272 , \7902 , \7931 );
xor \U$7930 ( \8273 , \8272 , \7942 );
xor \U$7931 ( \8274 , \7947 , \7949 );
xor \U$7932 ( \8275 , \8274 , \7952 );
and \U$7933 ( \8276 , \8273 , \8275 );
xor \U$7934 ( \8277 , \7966 , \7968 );
xor \U$7935 ( \8278 , \8277 , \7971 );
and \U$7936 ( \8279 , \8275 , \8278 );
and \U$7937 ( \8280 , \8273 , \8278 );
or \U$7938 ( \8281 , \8276 , \8279 , \8280 );
and \U$7939 ( \8282 , \8271 , \8281 );
xor \U$7940 ( \8283 , \7979 , \7981 );
xor \U$7941 ( \8284 , \8283 , \7983 );
and \U$7942 ( \8285 , \8281 , \8284 );
and \U$7943 ( \8286 , \8271 , \8284 );
or \U$7944 ( \8287 , \8282 , \8285 , \8286 );
xor \U$7945 ( \8288 , \7685 , \7702 );
xor \U$7946 ( \8289 , \8288 , \7708 );
and \U$7947 ( \8290 , \8287 , \8289 );
xor \U$7948 ( \8291 , \7977 , \7986 );
xor \U$7949 ( \8292 , \8291 , \7989 );
and \U$7950 ( \8293 , \8289 , \8292 );
and \U$7951 ( \8294 , \8287 , \8292 );
or \U$7952 ( \8295 , \8290 , \8293 , \8294 );
xor \U$7953 ( \8296 , \7992 , \7994 );
xor \U$7954 ( \8297 , \8296 , \7997 );
and \U$7955 ( \8298 , \8295 , \8297 );
and \U$7956 ( \8299 , \8006 , \8298 );
xor \U$7957 ( \8300 , \8006 , \8298 );
xor \U$7958 ( \8301 , \8295 , \8297 );
and \U$7959 ( \8302 , \385 , \7035 );
and \U$7960 ( \8303 , \393 , \7033 );
nor \U$7961 ( \8304 , \8302 , \8303 );
xnor \U$7962 ( \8305 , \8304 , \6775 );
and \U$7963 ( \8306 , \400 , \6541 );
and \U$7964 ( \8307 , \408 , \6539 );
nor \U$7965 ( \8308 , \8306 , \8307 );
xnor \U$7966 ( \8309 , \8308 , \6226 );
and \U$7967 ( \8310 , \8305 , \8309 );
and \U$7968 ( \8311 , \416 , \6032 );
and \U$7969 ( \8312 , \424 , \6030 );
nor \U$7970 ( \8313 , \8311 , \8312 );
xnor \U$7971 ( \8314 , \8313 , \5692 );
and \U$7972 ( \8315 , \8309 , \8314 );
and \U$7973 ( \8316 , \8305 , \8314 );
or \U$7974 ( \8317 , \8310 , \8315 , \8316 );
buf \U$7975 ( \8318 , RIbb2db58_58);
buf \U$7976 ( \8319 , RIbb2dae0_59);
and \U$7977 ( \8320 , \8318 , \8319 );
not \U$7978 ( \8321 , \8320 );
and \U$7979 ( \8322 , \7810 , \8321 );
not \U$7980 ( \8323 , \8322 );
and \U$7981 ( \8324 , \351 , \8131 );
and \U$7982 ( \8325 , \359 , \8129 );
nor \U$7983 ( \8326 , \8324 , \8325 );
xnor \U$7984 ( \8327 , \8326 , \7813 );
and \U$7985 ( \8328 , \8323 , \8327 );
and \U$7986 ( \8329 , \367 , \7564 );
and \U$7987 ( \8330 , \375 , \7562 );
nor \U$7988 ( \8331 , \8329 , \8330 );
xnor \U$7989 ( \8332 , \8331 , \7315 );
and \U$7990 ( \8333 , \8327 , \8332 );
and \U$7991 ( \8334 , \8323 , \8332 );
or \U$7992 ( \8335 , \8328 , \8333 , \8334 );
and \U$7993 ( \8336 , \8317 , \8335 );
and \U$7994 ( \8337 , \435 , \5443 );
and \U$7995 ( \8338 , \443 , \5441 );
nor \U$7996 ( \8339 , \8337 , \8338 );
xnor \U$7997 ( \8340 , \8339 , \5202 );
and \U$7998 ( \8341 , \661 , \4977 );
and \U$7999 ( \8342 , \450 , \4975 );
nor \U$8000 ( \8343 , \8341 , \8342 );
xnor \U$8001 ( \8344 , \8343 , \4789 );
and \U$8002 ( \8345 , \8340 , \8344 );
and \U$8003 ( \8346 , \785 , \4603 );
and \U$8004 ( \8347 , \722 , \4601 );
nor \U$8005 ( \8348 , \8346 , \8347 );
xnor \U$8006 ( \8349 , \8348 , \4371 );
and \U$8007 ( \8350 , \8344 , \8349 );
and \U$8008 ( \8351 , \8340 , \8349 );
or \U$8009 ( \8352 , \8345 , \8350 , \8351 );
and \U$8010 ( \8353 , \8335 , \8352 );
and \U$8011 ( \8354 , \8317 , \8352 );
or \U$8012 ( \8355 , \8336 , \8353 , \8354 );
and \U$8013 ( \8356 , \2463 , \2097 );
and \U$8014 ( \8357 , \2438 , \2095 );
nor \U$8015 ( \8358 , \8356 , \8357 );
xnor \U$8016 ( \8359 , \8358 , \1960 );
and \U$8017 ( \8360 , \2804 , \1891 );
and \U$8018 ( \8361 , \2637 , \1889 );
nor \U$8019 ( \8362 , \8360 , \8361 );
xnor \U$8020 ( \8363 , \8362 , \1739 );
and \U$8021 ( \8364 , \8359 , \8363 );
and \U$8022 ( \8365 , \3061 , \1623 );
and \U$8023 ( \8366 , \2942 , \1621 );
nor \U$8024 ( \8367 , \8365 , \8366 );
xnor \U$8025 ( \8368 , \8367 , \1467 );
and \U$8026 ( \8369 , \8363 , \8368 );
and \U$8027 ( \8370 , \8359 , \8368 );
or \U$8028 ( \8371 , \8364 , \8369 , \8370 );
and \U$8029 ( \8372 , \1596 , \3121 );
and \U$8030 ( \8373 , \1588 , \3119 );
nor \U$8031 ( \8374 , \8372 , \8373 );
xnor \U$8032 ( \8375 , \8374 , \2916 );
and \U$8033 ( \8376 , \1844 , \2715 );
and \U$8034 ( \8377 , \1839 , \2713 );
nor \U$8035 ( \8378 , \8376 , \8377 );
xnor \U$8036 ( \8379 , \8378 , \2566 );
and \U$8037 ( \8380 , \8375 , \8379 );
and \U$8038 ( \8381 , \2174 , \2393 );
and \U$8039 ( \8382 , \2030 , \2391 );
nor \U$8040 ( \8383 , \8381 , \8382 );
xnor \U$8041 ( \8384 , \8383 , \2251 );
and \U$8042 ( \8385 , \8379 , \8384 );
and \U$8043 ( \8386 , \8375 , \8384 );
or \U$8044 ( \8387 , \8380 , \8385 , \8386 );
and \U$8045 ( \8388 , \8371 , \8387 );
and \U$8046 ( \8389 , \1071 , \4152 );
and \U$8047 ( \8390 , \983 , \4150 );
nor \U$8048 ( \8391 , \8389 , \8390 );
xnor \U$8049 ( \8392 , \8391 , \4009 );
and \U$8050 ( \8393 , \1181 , \3829 );
and \U$8051 ( \8394 , \1176 , \3827 );
nor \U$8052 ( \8395 , \8393 , \8394 );
xnor \U$8053 ( \8396 , \8395 , \3583 );
and \U$8054 ( \8397 , \8392 , \8396 );
and \U$8055 ( \8398 , \1412 , \3434 );
and \U$8056 ( \8399 , \1297 , \3432 );
nor \U$8057 ( \8400 , \8398 , \8399 );
xnor \U$8058 ( \8401 , \8400 , \3247 );
and \U$8059 ( \8402 , \8396 , \8401 );
and \U$8060 ( \8403 , \8392 , \8401 );
or \U$8061 ( \8404 , \8397 , \8402 , \8403 );
and \U$8062 ( \8405 , \8387 , \8404 );
and \U$8063 ( \8406 , \8371 , \8404 );
or \U$8064 ( \8407 , \8388 , \8405 , \8406 );
and \U$8065 ( \8408 , \8355 , \8407 );
and \U$8066 ( \8409 , \4576 , \793 );
and \U$8067 ( \8410 , \4568 , \791 );
nor \U$8068 ( \8411 , \8409 , \8410 );
xnor \U$8069 ( \8412 , \8411 , \699 );
and \U$8070 ( \8413 , \5050 , \624 );
and \U$8071 ( \8414 , \5045 , \622 );
nor \U$8072 ( \8415 , \8413 , \8414 );
xnor \U$8073 ( \8416 , \8415 , \349 );
and \U$8074 ( \8417 , \8412 , \8416 );
and \U$8075 ( \8418 , \5573 , \357 );
and \U$8076 ( \8419 , \5314 , \355 );
nor \U$8077 ( \8420 , \8418 , \8419 );
xnor \U$8078 ( \8421 , \8420 , \364 );
and \U$8079 ( \8422 , \8416 , \8421 );
and \U$8080 ( \8423 , \8412 , \8421 );
or \U$8081 ( \8424 , \8417 , \8422 , \8423 );
and \U$8082 ( \8425 , \3686 , \1351 );
and \U$8083 ( \8426 , \3478 , \1349 );
nor \U$8084 ( \8427 , \8425 , \8426 );
xnor \U$8085 ( \8428 , \8427 , \1238 );
and \U$8086 ( \8429 , \3813 , \1157 );
and \U$8087 ( \8430 , \3808 , \1155 );
nor \U$8088 ( \8431 , \8429 , \8430 );
xnor \U$8089 ( \8432 , \8431 , \1021 );
and \U$8090 ( \8433 , \8428 , \8432 );
and \U$8091 ( \8434 , \4266 , \957 );
and \U$8092 ( \8435 , \4069 , \955 );
nor \U$8093 ( \8436 , \8434 , \8435 );
xnor \U$8094 ( \8437 , \8436 , \879 );
and \U$8095 ( \8438 , \8432 , \8437 );
and \U$8096 ( \8439 , \8428 , \8437 );
or \U$8097 ( \8440 , \8433 , \8438 , \8439 );
and \U$8098 ( \8441 , \8424 , \8440 );
and \U$8099 ( \8442 , \5954 , \373 );
and \U$8100 ( \8443 , \5945 , \371 );
nor \U$8101 ( \8444 , \8442 , \8443 );
xnor \U$8102 ( \8445 , \8444 , \380 );
and \U$8103 ( \8446 , \6499 , \391 );
and \U$8104 ( \8447 , \6297 , \389 );
nor \U$8105 ( \8448 , \8446 , \8447 );
xnor \U$8106 ( \8449 , \8448 , \398 );
and \U$8107 ( \8450 , \8445 , \8449 );
and \U$8108 ( \8451 , \6974 , \406 );
and \U$8109 ( \8452 , \6802 , \404 );
nor \U$8110 ( \8453 , \8451 , \8452 );
xnor \U$8111 ( \8454 , \8453 , \413 );
and \U$8112 ( \8455 , \8449 , \8454 );
and \U$8113 ( \8456 , \8445 , \8454 );
or \U$8114 ( \8457 , \8450 , \8455 , \8456 );
and \U$8115 ( \8458 , \8440 , \8457 );
and \U$8116 ( \8459 , \8424 , \8457 );
or \U$8117 ( \8460 , \8441 , \8458 , \8459 );
and \U$8118 ( \8461 , \8407 , \8460 );
and \U$8119 ( \8462 , \8355 , \8460 );
or \U$8120 ( \8463 , \8408 , \8461 , \8462 );
xor \U$8121 ( \8464 , \8010 , \8014 );
xor \U$8122 ( \8465 , \8464 , \8019 );
xor \U$8123 ( \8466 , \8115 , \8119 );
xor \U$8124 ( \8467 , \8466 , \8124 );
and \U$8125 ( \8468 , \8465 , \8467 );
xor \U$8126 ( \8469 , \8043 , \8047 );
xor \U$8127 ( \8470 , \8469 , \8052 );
and \U$8128 ( \8471 , \8467 , \8470 );
and \U$8129 ( \8472 , \8465 , \8470 );
or \U$8130 ( \8473 , \8468 , \8471 , \8472 );
xor \U$8131 ( \8474 , \8026 , \8030 );
xor \U$8132 ( \8475 , \8474 , \8035 );
xor \U$8133 ( \8476 , \8062 , \8066 );
xor \U$8134 ( \8477 , \8476 , \8071 );
and \U$8135 ( \8478 , \8475 , \8477 );
xor \U$8136 ( \8479 , \8078 , \8082 );
xor \U$8137 ( \8480 , \8479 , \8087 );
and \U$8138 ( \8481 , \8477 , \8480 );
and \U$8139 ( \8482 , \8475 , \8480 );
or \U$8140 ( \8483 , \8478 , \8481 , \8482 );
and \U$8141 ( \8484 , \8473 , \8483 );
and \U$8142 ( \8485 , \7924 , \422 );
and \U$8143 ( \8486 , \7500 , \420 );
nor \U$8144 ( \8487 , \8485 , \8486 );
xnor \U$8145 ( \8488 , \8487 , \429 );
and \U$8146 ( \8489 , \8175 , \441 );
and \U$8147 ( \8490 , \8170 , \439 );
nor \U$8148 ( \8491 , \8489 , \8490 );
xnor \U$8149 ( \8492 , \8491 , \448 );
and \U$8150 ( \8493 , \8488 , \8492 );
buf \U$8151 ( \8494 , RIbb2bdd0_121);
and \U$8152 ( \8495 , \8494 , \436 );
and \U$8153 ( \8496 , \8492 , \8495 );
and \U$8154 ( \8497 , \8488 , \8495 );
or \U$8155 ( \8498 , \8493 , \8496 , \8497 );
xor \U$8156 ( \8499 , \8095 , \8099 );
xor \U$8157 ( \8500 , \8499 , \8104 );
and \U$8158 ( \8501 , \8498 , \8500 );
xnor \U$8159 ( \8502 , \8174 , \8176 );
and \U$8160 ( \8503 , \8500 , \8502 );
and \U$8161 ( \8504 , \8498 , \8502 );
or \U$8162 ( \8505 , \8501 , \8503 , \8504 );
and \U$8163 ( \8506 , \8483 , \8505 );
and \U$8164 ( \8507 , \8473 , \8505 );
or \U$8165 ( \8508 , \8484 , \8506 , \8507 );
and \U$8166 ( \8509 , \8463 , \8508 );
xor \U$8167 ( \8510 , \8188 , \8190 );
xor \U$8168 ( \8511 , \8510 , \8193 );
xor \U$8169 ( \8512 , \8199 , \8201 );
xor \U$8170 ( \8513 , \8512 , \8204 );
and \U$8171 ( \8514 , \8511 , \8513 );
xor \U$8172 ( \8515 , \8213 , \8215 );
xor \U$8173 ( \8516 , \8515 , \8218 );
and \U$8174 ( \8517 , \8513 , \8516 );
and \U$8175 ( \8518 , \8511 , \8516 );
or \U$8176 ( \8519 , \8514 , \8517 , \8518 );
and \U$8177 ( \8520 , \8508 , \8519 );
and \U$8178 ( \8521 , \8463 , \8519 );
or \U$8179 ( \8522 , \8509 , \8520 , \8521 );
xor \U$8180 ( \8523 , \8058 , \8110 );
xor \U$8181 ( \8524 , \8523 , \8166 );
xor \U$8182 ( \8525 , \8186 , \8196 );
xor \U$8183 ( \8526 , \8525 , \8207 );
and \U$8184 ( \8527 , \8524 , \8526 );
xor \U$8185 ( \8528 , \8221 , \8223 );
xor \U$8186 ( \8529 , \8528 , \8226 );
and \U$8187 ( \8530 , \8526 , \8529 );
and \U$8188 ( \8531 , \8524 , \8529 );
or \U$8189 ( \8532 , \8527 , \8530 , \8531 );
and \U$8190 ( \8533 , \8522 , \8532 );
xor \U$8191 ( \8534 , \8022 , \8038 );
xor \U$8192 ( \8535 , \8534 , \8055 );
xor \U$8193 ( \8536 , \8074 , \8090 );
xor \U$8194 ( \8537 , \8536 , \8107 );
and \U$8195 ( \8538 , \8535 , \8537 );
xor \U$8196 ( \8539 , \8177 , \8181 );
xor \U$8197 ( \8540 , \8539 , \8183 );
and \U$8198 ( \8541 , \8537 , \8540 );
and \U$8199 ( \8542 , \8535 , \8540 );
or \U$8200 ( \8543 , \8538 , \8541 , \8542 );
xor \U$8201 ( \8544 , \8234 , \8236 );
xor \U$8202 ( \8545 , \8544 , \8239 );
and \U$8203 ( \8546 , \8543 , \8545 );
xor \U$8204 ( \8547 , \8244 , \8246 );
xor \U$8205 ( \8548 , \8547 , \8248 );
and \U$8206 ( \8549 , \8545 , \8548 );
and \U$8207 ( \8550 , \8543 , \8548 );
or \U$8208 ( \8551 , \8546 , \8549 , \8550 );
and \U$8209 ( \8552 , \8532 , \8551 );
and \U$8210 ( \8553 , \8522 , \8551 );
or \U$8211 ( \8554 , \8533 , \8552 , \8553 );
xor \U$8212 ( \8555 , \7792 , \7846 );
xor \U$8213 ( \8556 , \8555 , \7899 );
xor \U$8214 ( \8557 , \8242 , \8251 );
xor \U$8215 ( \8558 , \8557 , \8254 );
and \U$8216 ( \8559 , \8556 , \8558 );
xor \U$8217 ( \8560 , \8260 , \8262 );
xor \U$8218 ( \8561 , \8560 , \8265 );
and \U$8219 ( \8562 , \8558 , \8561 );
and \U$8220 ( \8563 , \8556 , \8561 );
or \U$8221 ( \8564 , \8559 , \8562 , \8563 );
and \U$8222 ( \8565 , \8554 , \8564 );
xor \U$8223 ( \8566 , \8273 , \8275 );
xor \U$8224 ( \8567 , \8566 , \8278 );
and \U$8225 ( \8568 , \8564 , \8567 );
and \U$8226 ( \8569 , \8554 , \8567 );
or \U$8227 ( \8570 , \8565 , \8568 , \8569 );
xor \U$8228 ( \8571 , \7945 , \7955 );
xor \U$8229 ( \8572 , \8571 , \7974 );
and \U$8230 ( \8573 , \8570 , \8572 );
xor \U$8231 ( \8574 , \8271 , \8281 );
xor \U$8232 ( \8575 , \8574 , \8284 );
and \U$8233 ( \8576 , \8572 , \8575 );
and \U$8234 ( \8577 , \8570 , \8575 );
or \U$8235 ( \8578 , \8573 , \8576 , \8577 );
xor \U$8236 ( \8579 , \8287 , \8289 );
xor \U$8237 ( \8580 , \8579 , \8292 );
and \U$8238 ( \8581 , \8578 , \8580 );
and \U$8239 ( \8582 , \8301 , \8581 );
xor \U$8240 ( \8583 , \8301 , \8581 );
xor \U$8241 ( \8584 , \8578 , \8580 );
and \U$8242 ( \8585 , \2637 , \2097 );
and \U$8243 ( \8586 , \2463 , \2095 );
nor \U$8244 ( \8587 , \8585 , \8586 );
xnor \U$8245 ( \8588 , \8587 , \1960 );
and \U$8246 ( \8589 , \2942 , \1891 );
and \U$8247 ( \8590 , \2804 , \1889 );
nor \U$8248 ( \8591 , \8589 , \8590 );
xnor \U$8249 ( \8592 , \8591 , \1739 );
and \U$8250 ( \8593 , \8588 , \8592 );
and \U$8251 ( \8594 , \3478 , \1623 );
and \U$8252 ( \8595 , \3061 , \1621 );
nor \U$8253 ( \8596 , \8594 , \8595 );
xnor \U$8254 ( \8597 , \8596 , \1467 );
and \U$8255 ( \8598 , \8592 , \8597 );
and \U$8256 ( \8599 , \8588 , \8597 );
or \U$8257 ( \8600 , \8593 , \8598 , \8599 );
and \U$8258 ( \8601 , \1176 , \4152 );
and \U$8259 ( \8602 , \1071 , \4150 );
nor \U$8260 ( \8603 , \8601 , \8602 );
xnor \U$8261 ( \8604 , \8603 , \4009 );
and \U$8262 ( \8605 , \1297 , \3829 );
and \U$8263 ( \8606 , \1181 , \3827 );
nor \U$8264 ( \8607 , \8605 , \8606 );
xnor \U$8265 ( \8608 , \8607 , \3583 );
and \U$8266 ( \8609 , \8604 , \8608 );
and \U$8267 ( \8610 , \1588 , \3434 );
and \U$8268 ( \8611 , \1412 , \3432 );
nor \U$8269 ( \8612 , \8610 , \8611 );
xnor \U$8270 ( \8613 , \8612 , \3247 );
and \U$8271 ( \8614 , \8608 , \8613 );
and \U$8272 ( \8615 , \8604 , \8613 );
or \U$8273 ( \8616 , \8609 , \8614 , \8615 );
and \U$8274 ( \8617 , \8600 , \8616 );
and \U$8275 ( \8618 , \1839 , \3121 );
and \U$8276 ( \8619 , \1596 , \3119 );
nor \U$8277 ( \8620 , \8618 , \8619 );
xnor \U$8278 ( \8621 , \8620 , \2916 );
and \U$8279 ( \8622 , \2030 , \2715 );
and \U$8280 ( \8623 , \1844 , \2713 );
nor \U$8281 ( \8624 , \8622 , \8623 );
xnor \U$8282 ( \8625 , \8624 , \2566 );
and \U$8283 ( \8626 , \8621 , \8625 );
and \U$8284 ( \8627 , \2438 , \2393 );
and \U$8285 ( \8628 , \2174 , \2391 );
nor \U$8286 ( \8629 , \8627 , \8628 );
xnor \U$8287 ( \8630 , \8629 , \2251 );
and \U$8288 ( \8631 , \8625 , \8630 );
and \U$8289 ( \8632 , \8621 , \8630 );
or \U$8290 ( \8633 , \8626 , \8631 , \8632 );
and \U$8291 ( \8634 , \8616 , \8633 );
and \U$8292 ( \8635 , \8600 , \8633 );
or \U$8293 ( \8636 , \8617 , \8634 , \8635 );
and \U$8294 ( \8637 , \6297 , \373 );
and \U$8295 ( \8638 , \5954 , \371 );
nor \U$8296 ( \8639 , \8637 , \8638 );
xnor \U$8297 ( \8640 , \8639 , \380 );
and \U$8298 ( \8641 , \6802 , \391 );
and \U$8299 ( \8642 , \6499 , \389 );
nor \U$8300 ( \8643 , \8641 , \8642 );
xnor \U$8301 ( \8644 , \8643 , \398 );
and \U$8302 ( \8645 , \8640 , \8644 );
and \U$8303 ( \8646 , \7500 , \406 );
and \U$8304 ( \8647 , \6974 , \404 );
nor \U$8305 ( \8648 , \8646 , \8647 );
xnor \U$8306 ( \8649 , \8648 , \413 );
and \U$8307 ( \8650 , \8644 , \8649 );
and \U$8308 ( \8651 , \8640 , \8649 );
or \U$8309 ( \8652 , \8645 , \8650 , \8651 );
and \U$8310 ( \8653 , \5045 , \793 );
and \U$8311 ( \8654 , \4576 , \791 );
nor \U$8312 ( \8655 , \8653 , \8654 );
xnor \U$8313 ( \8656 , \8655 , \699 );
and \U$8314 ( \8657 , \5314 , \624 );
and \U$8315 ( \8658 , \5050 , \622 );
nor \U$8316 ( \8659 , \8657 , \8658 );
xnor \U$8317 ( \8660 , \8659 , \349 );
and \U$8318 ( \8661 , \8656 , \8660 );
and \U$8319 ( \8662 , \5945 , \357 );
and \U$8320 ( \8663 , \5573 , \355 );
nor \U$8321 ( \8664 , \8662 , \8663 );
xnor \U$8322 ( \8665 , \8664 , \364 );
and \U$8323 ( \8666 , \8660 , \8665 );
and \U$8324 ( \8667 , \8656 , \8665 );
or \U$8325 ( \8668 , \8661 , \8666 , \8667 );
and \U$8326 ( \8669 , \8652 , \8668 );
and \U$8327 ( \8670 , \3808 , \1351 );
and \U$8328 ( \8671 , \3686 , \1349 );
nor \U$8329 ( \8672 , \8670 , \8671 );
xnor \U$8330 ( \8673 , \8672 , \1238 );
and \U$8331 ( \8674 , \4069 , \1157 );
and \U$8332 ( \8675 , \3813 , \1155 );
nor \U$8333 ( \8676 , \8674 , \8675 );
xnor \U$8334 ( \8677 , \8676 , \1021 );
and \U$8335 ( \8678 , \8673 , \8677 );
and \U$8336 ( \8679 , \4568 , \957 );
and \U$8337 ( \8680 , \4266 , \955 );
nor \U$8338 ( \8681 , \8679 , \8680 );
xnor \U$8339 ( \8682 , \8681 , \879 );
and \U$8340 ( \8683 , \8677 , \8682 );
and \U$8341 ( \8684 , \8673 , \8682 );
or \U$8342 ( \8685 , \8678 , \8683 , \8684 );
and \U$8343 ( \8686 , \8668 , \8685 );
and \U$8344 ( \8687 , \8652 , \8685 );
or \U$8345 ( \8688 , \8669 , \8686 , \8687 );
and \U$8346 ( \8689 , \8636 , \8688 );
xor \U$8347 ( \8690 , \7810 , \8318 );
xor \U$8348 ( \8691 , \8318 , \8319 );
not \U$8349 ( \8692 , \8691 );
and \U$8350 ( \8693 , \8690 , \8692 );
and \U$8351 ( \8694 , \359 , \8693 );
not \U$8352 ( \8695 , \8694 );
xnor \U$8353 ( \8696 , \8695 , \8322 );
and \U$8354 ( \8697 , \375 , \8131 );
and \U$8355 ( \8698 , \351 , \8129 );
nor \U$8356 ( \8699 , \8697 , \8698 );
xnor \U$8357 ( \8700 , \8699 , \7813 );
and \U$8358 ( \8701 , \8696 , \8700 );
and \U$8359 ( \8702 , \393 , \7564 );
and \U$8360 ( \8703 , \367 , \7562 );
nor \U$8361 ( \8704 , \8702 , \8703 );
xnor \U$8362 ( \8705 , \8704 , \7315 );
and \U$8363 ( \8706 , \8700 , \8705 );
and \U$8364 ( \8707 , \8696 , \8705 );
or \U$8365 ( \8708 , \8701 , \8706 , \8707 );
and \U$8366 ( \8709 , \450 , \5443 );
and \U$8367 ( \8710 , \435 , \5441 );
nor \U$8368 ( \8711 , \8709 , \8710 );
xnor \U$8369 ( \8712 , \8711 , \5202 );
and \U$8370 ( \8713 , \722 , \4977 );
and \U$8371 ( \8714 , \661 , \4975 );
nor \U$8372 ( \8715 , \8713 , \8714 );
xnor \U$8373 ( \8716 , \8715 , \4789 );
and \U$8374 ( \8717 , \8712 , \8716 );
and \U$8375 ( \8718 , \983 , \4603 );
and \U$8376 ( \8719 , \785 , \4601 );
nor \U$8377 ( \8720 , \8718 , \8719 );
xnor \U$8378 ( \8721 , \8720 , \4371 );
and \U$8379 ( \8722 , \8716 , \8721 );
and \U$8380 ( \8723 , \8712 , \8721 );
or \U$8381 ( \8724 , \8717 , \8722 , \8723 );
and \U$8382 ( \8725 , \8708 , \8724 );
and \U$8383 ( \8726 , \408 , \7035 );
and \U$8384 ( \8727 , \385 , \7033 );
nor \U$8385 ( \8728 , \8726 , \8727 );
xnor \U$8386 ( \8729 , \8728 , \6775 );
and \U$8387 ( \8730 , \424 , \6541 );
and \U$8388 ( \8731 , \400 , \6539 );
nor \U$8389 ( \8732 , \8730 , \8731 );
xnor \U$8390 ( \8733 , \8732 , \6226 );
and \U$8391 ( \8734 , \8729 , \8733 );
and \U$8392 ( \8735 , \443 , \6032 );
and \U$8393 ( \8736 , \416 , \6030 );
nor \U$8394 ( \8737 , \8735 , \8736 );
xnor \U$8395 ( \8738 , \8737 , \5692 );
and \U$8396 ( \8739 , \8733 , \8738 );
and \U$8397 ( \8740 , \8729 , \8738 );
or \U$8398 ( \8741 , \8734 , \8739 , \8740 );
and \U$8399 ( \8742 , \8724 , \8741 );
and \U$8400 ( \8743 , \8708 , \8741 );
or \U$8401 ( \8744 , \8725 , \8742 , \8743 );
and \U$8402 ( \8745 , \8688 , \8744 );
and \U$8403 ( \8746 , \8636 , \8744 );
or \U$8404 ( \8747 , \8689 , \8745 , \8746 );
xor \U$8405 ( \8748 , \8340 , \8344 );
xor \U$8406 ( \8749 , \8748 , \8349 );
xor \U$8407 ( \8750 , \8375 , \8379 );
xor \U$8408 ( \8751 , \8750 , \8384 );
and \U$8409 ( \8752 , \8749 , \8751 );
xor \U$8410 ( \8753 , \8392 , \8396 );
xor \U$8411 ( \8754 , \8753 , \8401 );
and \U$8412 ( \8755 , \8751 , \8754 );
and \U$8413 ( \8756 , \8749 , \8754 );
or \U$8414 ( \8757 , \8752 , \8755 , \8756 );
xor \U$8415 ( \8758 , \8359 , \8363 );
xor \U$8416 ( \8759 , \8758 , \8368 );
xor \U$8417 ( \8760 , \8412 , \8416 );
xor \U$8418 ( \8761 , \8760 , \8421 );
and \U$8419 ( \8762 , \8759 , \8761 );
xor \U$8420 ( \8763 , \8428 , \8432 );
xor \U$8421 ( \8764 , \8763 , \8437 );
and \U$8422 ( \8765 , \8761 , \8764 );
and \U$8423 ( \8766 , \8759 , \8764 );
or \U$8424 ( \8767 , \8762 , \8765 , \8766 );
and \U$8425 ( \8768 , \8757 , \8767 );
and \U$8426 ( \8769 , \8170 , \422 );
and \U$8427 ( \8770 , \7924 , \420 );
nor \U$8428 ( \8771 , \8769 , \8770 );
xnor \U$8429 ( \8772 , \8771 , \429 );
and \U$8430 ( \8773 , \8494 , \441 );
and \U$8431 ( \8774 , \8175 , \439 );
nor \U$8432 ( \8775 , \8773 , \8774 );
xnor \U$8433 ( \8776 , \8775 , \448 );
and \U$8434 ( \8777 , \8772 , \8776 );
buf \U$8435 ( \8778 , RIbb2bd58_122);
and \U$8436 ( \8779 , \8778 , \436 );
and \U$8437 ( \8780 , \8776 , \8779 );
and \U$8438 ( \8781 , \8772 , \8779 );
or \U$8439 ( \8782 , \8777 , \8780 , \8781 );
xor \U$8440 ( \8783 , \8488 , \8492 );
xor \U$8441 ( \8784 , \8783 , \8495 );
and \U$8442 ( \8785 , \8782 , \8784 );
xor \U$8443 ( \8786 , \8445 , \8449 );
xor \U$8444 ( \8787 , \8786 , \8454 );
and \U$8445 ( \8788 , \8784 , \8787 );
and \U$8446 ( \8789 , \8782 , \8787 );
or \U$8447 ( \8790 , \8785 , \8788 , \8789 );
and \U$8448 ( \8791 , \8767 , \8790 );
and \U$8449 ( \8792 , \8757 , \8790 );
or \U$8450 ( \8793 , \8768 , \8791 , \8792 );
and \U$8451 ( \8794 , \8747 , \8793 );
xor \U$8452 ( \8795 , \8134 , \8138 );
xor \U$8453 ( \8796 , \8795 , \8143 );
xor \U$8454 ( \8797 , \8151 , \8155 );
xor \U$8455 ( \8798 , \8797 , \8160 );
and \U$8456 ( \8799 , \8796 , \8798 );
xor \U$8457 ( \8800 , \8465 , \8467 );
xor \U$8458 ( \8801 , \8800 , \8470 );
and \U$8459 ( \8802 , \8798 , \8801 );
and \U$8460 ( \8803 , \8796 , \8801 );
or \U$8461 ( \8804 , \8799 , \8802 , \8803 );
and \U$8462 ( \8805 , \8793 , \8804 );
and \U$8463 ( \8806 , \8747 , \8804 );
or \U$8464 ( \8807 , \8794 , \8805 , \8806 );
xor \U$8465 ( \8808 , \8424 , \8440 );
xor \U$8466 ( \8809 , \8808 , \8457 );
xor \U$8467 ( \8810 , \8475 , \8477 );
xor \U$8468 ( \8811 , \8810 , \8480 );
and \U$8469 ( \8812 , \8809 , \8811 );
xor \U$8470 ( \8813 , \8498 , \8500 );
xor \U$8471 ( \8814 , \8813 , \8502 );
and \U$8472 ( \8815 , \8811 , \8814 );
and \U$8473 ( \8816 , \8809 , \8814 );
or \U$8474 ( \8817 , \8812 , \8815 , \8816 );
xor \U$8475 ( \8818 , \8127 , \8146 );
xor \U$8476 ( \8819 , \8818 , \8163 );
and \U$8477 ( \8820 , \8817 , \8819 );
xor \U$8478 ( \8821 , \8535 , \8537 );
xor \U$8479 ( \8822 , \8821 , \8540 );
and \U$8480 ( \8823 , \8819 , \8822 );
and \U$8481 ( \8824 , \8817 , \8822 );
or \U$8482 ( \8825 , \8820 , \8823 , \8824 );
and \U$8483 ( \8826 , \8807 , \8825 );
xor \U$8484 ( \8827 , \8355 , \8407 );
xor \U$8485 ( \8828 , \8827 , \8460 );
xor \U$8486 ( \8829 , \8473 , \8483 );
xor \U$8487 ( \8830 , \8829 , \8505 );
and \U$8488 ( \8831 , \8828 , \8830 );
xor \U$8489 ( \8832 , \8511 , \8513 );
xor \U$8490 ( \8833 , \8832 , \8516 );
and \U$8491 ( \8834 , \8830 , \8833 );
and \U$8492 ( \8835 , \8828 , \8833 );
or \U$8493 ( \8836 , \8831 , \8834 , \8835 );
and \U$8494 ( \8837 , \8825 , \8836 );
and \U$8495 ( \8838 , \8807 , \8836 );
or \U$8496 ( \8839 , \8826 , \8837 , \8838 );
xor \U$8497 ( \8840 , \8463 , \8508 );
xor \U$8498 ( \8841 , \8840 , \8519 );
xor \U$8499 ( \8842 , \8524 , \8526 );
xor \U$8500 ( \8843 , \8842 , \8529 );
and \U$8501 ( \8844 , \8841 , \8843 );
xor \U$8502 ( \8845 , \8543 , \8545 );
xor \U$8503 ( \8846 , \8845 , \8548 );
and \U$8504 ( \8847 , \8843 , \8846 );
and \U$8505 ( \8848 , \8841 , \8846 );
or \U$8506 ( \8849 , \8844 , \8847 , \8848 );
and \U$8507 ( \8850 , \8839 , \8849 );
xor \U$8508 ( \8851 , \8169 , \8210 );
xor \U$8509 ( \8852 , \8851 , \8229 );
and \U$8510 ( \8853 , \8849 , \8852 );
and \U$8511 ( \8854 , \8839 , \8852 );
or \U$8512 ( \8855 , \8850 , \8853 , \8854 );
xor \U$8513 ( \8856 , \8522 , \8532 );
xor \U$8514 ( \8857 , \8856 , \8551 );
xor \U$8515 ( \8858 , \8556 , \8558 );
xor \U$8516 ( \8859 , \8858 , \8561 );
and \U$8517 ( \8860 , \8857 , \8859 );
and \U$8518 ( \8861 , \8855 , \8860 );
xor \U$8519 ( \8862 , \8232 , \8257 );
xor \U$8520 ( \8863 , \8862 , \8268 );
and \U$8521 ( \8864 , \8860 , \8863 );
and \U$8522 ( \8865 , \8855 , \8863 );
or \U$8523 ( \8866 , \8861 , \8864 , \8865 );
xor \U$8524 ( \8867 , \8570 , \8572 );
xor \U$8525 ( \8868 , \8867 , \8575 );
and \U$8526 ( \8869 , \8866 , \8868 );
and \U$8527 ( \8870 , \8584 , \8869 );
xor \U$8528 ( \8871 , \8584 , \8869 );
xor \U$8529 ( \8872 , \8866 , \8868 );
xor \U$8530 ( \8873 , \8640 , \8644 );
xor \U$8531 ( \8874 , \8873 , \8649 );
xor \U$8532 ( \8875 , \8656 , \8660 );
xor \U$8533 ( \8876 , \8875 , \8665 );
and \U$8534 ( \8877 , \8874 , \8876 );
xor \U$8535 ( \8878 , \8673 , \8677 );
xor \U$8536 ( \8879 , \8878 , \8682 );
and \U$8537 ( \8880 , \8876 , \8879 );
and \U$8538 ( \8881 , \8874 , \8879 );
or \U$8539 ( \8882 , \8877 , \8880 , \8881 );
xor \U$8540 ( \8883 , \8588 , \8592 );
xor \U$8541 ( \8884 , \8883 , \8597 );
xor \U$8542 ( \8885 , \8604 , \8608 );
xor \U$8543 ( \8886 , \8885 , \8613 );
and \U$8544 ( \8887 , \8884 , \8886 );
xor \U$8545 ( \8888 , \8621 , \8625 );
xor \U$8546 ( \8889 , \8888 , \8630 );
and \U$8547 ( \8890 , \8886 , \8889 );
and \U$8548 ( \8891 , \8884 , \8889 );
or \U$8549 ( \8892 , \8887 , \8890 , \8891 );
and \U$8550 ( \8893 , \8882 , \8892 );
and \U$8551 ( \8894 , \7924 , \406 );
and \U$8552 ( \8895 , \7500 , \404 );
nor \U$8553 ( \8896 , \8894 , \8895 );
xnor \U$8554 ( \8897 , \8896 , \413 );
and \U$8555 ( \8898 , \8175 , \422 );
and \U$8556 ( \8899 , \8170 , \420 );
nor \U$8557 ( \8900 , \8898 , \8899 );
xnor \U$8558 ( \8901 , \8900 , \429 );
and \U$8559 ( \8902 , \8897 , \8901 );
and \U$8560 ( \8903 , \8778 , \441 );
and \U$8561 ( \8904 , \8494 , \439 );
nor \U$8562 ( \8905 , \8903 , \8904 );
xnor \U$8563 ( \8906 , \8905 , \448 );
and \U$8564 ( \8907 , \8901 , \8906 );
and \U$8565 ( \8908 , \8897 , \8906 );
or \U$8566 ( \8909 , \8902 , \8907 , \8908 );
xor \U$8567 ( \8910 , \8772 , \8776 );
xor \U$8568 ( \8911 , \8910 , \8779 );
or \U$8569 ( \8912 , \8909 , \8911 );
and \U$8570 ( \8913 , \8892 , \8912 );
and \U$8571 ( \8914 , \8882 , \8912 );
or \U$8572 ( \8915 , \8893 , \8913 , \8914 );
buf \U$8573 ( \8916 , RIbb2da68_60);
buf \U$8574 ( \8917 , RIbb2d9f0_61);
and \U$8575 ( \8918 , \8916 , \8917 );
not \U$8576 ( \8919 , \8918 );
and \U$8577 ( \8920 , \8319 , \8919 );
not \U$8578 ( \8921 , \8920 );
and \U$8579 ( \8922 , \351 , \8693 );
and \U$8580 ( \8923 , \359 , \8691 );
nor \U$8581 ( \8924 , \8922 , \8923 );
xnor \U$8582 ( \8925 , \8924 , \8322 );
and \U$8583 ( \8926 , \8921 , \8925 );
and \U$8584 ( \8927 , \367 , \8131 );
and \U$8585 ( \8928 , \375 , \8129 );
nor \U$8586 ( \8929 , \8927 , \8928 );
xnor \U$8587 ( \8930 , \8929 , \7813 );
and \U$8588 ( \8931 , \8925 , \8930 );
and \U$8589 ( \8932 , \8921 , \8930 );
or \U$8590 ( \8933 , \8926 , \8931 , \8932 );
and \U$8591 ( \8934 , \435 , \6032 );
and \U$8592 ( \8935 , \443 , \6030 );
nor \U$8593 ( \8936 , \8934 , \8935 );
xnor \U$8594 ( \8937 , \8936 , \5692 );
and \U$8595 ( \8938 , \661 , \5443 );
and \U$8596 ( \8939 , \450 , \5441 );
nor \U$8597 ( \8940 , \8938 , \8939 );
xnor \U$8598 ( \8941 , \8940 , \5202 );
and \U$8599 ( \8942 , \8937 , \8941 );
and \U$8600 ( \8943 , \785 , \4977 );
and \U$8601 ( \8944 , \722 , \4975 );
nor \U$8602 ( \8945 , \8943 , \8944 );
xnor \U$8603 ( \8946 , \8945 , \4789 );
and \U$8604 ( \8947 , \8941 , \8946 );
and \U$8605 ( \8948 , \8937 , \8946 );
or \U$8606 ( \8949 , \8942 , \8947 , \8948 );
and \U$8607 ( \8950 , \8933 , \8949 );
and \U$8608 ( \8951 , \385 , \7564 );
and \U$8609 ( \8952 , \393 , \7562 );
nor \U$8610 ( \8953 , \8951 , \8952 );
xnor \U$8611 ( \8954 , \8953 , \7315 );
and \U$8612 ( \8955 , \400 , \7035 );
and \U$8613 ( \8956 , \408 , \7033 );
nor \U$8614 ( \8957 , \8955 , \8956 );
xnor \U$8615 ( \8958 , \8957 , \6775 );
and \U$8616 ( \8959 , \8954 , \8958 );
and \U$8617 ( \8960 , \416 , \6541 );
and \U$8618 ( \8961 , \424 , \6539 );
nor \U$8619 ( \8962 , \8960 , \8961 );
xnor \U$8620 ( \8963 , \8962 , \6226 );
and \U$8621 ( \8964 , \8958 , \8963 );
and \U$8622 ( \8965 , \8954 , \8963 );
or \U$8623 ( \8966 , \8959 , \8964 , \8965 );
and \U$8624 ( \8967 , \8949 , \8966 );
and \U$8625 ( \8968 , \8933 , \8966 );
or \U$8626 ( \8969 , \8950 , \8967 , \8968 );
and \U$8627 ( \8970 , \1596 , \3434 );
and \U$8628 ( \8971 , \1588 , \3432 );
nor \U$8629 ( \8972 , \8970 , \8971 );
xnor \U$8630 ( \8973 , \8972 , \3247 );
and \U$8631 ( \8974 , \1844 , \3121 );
and \U$8632 ( \8975 , \1839 , \3119 );
nor \U$8633 ( \8976 , \8974 , \8975 );
xnor \U$8634 ( \8977 , \8976 , \2916 );
and \U$8635 ( \8978 , \8973 , \8977 );
and \U$8636 ( \8979 , \2174 , \2715 );
and \U$8637 ( \8980 , \2030 , \2713 );
nor \U$8638 ( \8981 , \8979 , \8980 );
xnor \U$8639 ( \8982 , \8981 , \2566 );
and \U$8640 ( \8983 , \8977 , \8982 );
and \U$8641 ( \8984 , \8973 , \8982 );
or \U$8642 ( \8985 , \8978 , \8983 , \8984 );
and \U$8643 ( \8986 , \2463 , \2393 );
and \U$8644 ( \8987 , \2438 , \2391 );
nor \U$8645 ( \8988 , \8986 , \8987 );
xnor \U$8646 ( \8989 , \8988 , \2251 );
and \U$8647 ( \8990 , \2804 , \2097 );
and \U$8648 ( \8991 , \2637 , \2095 );
nor \U$8649 ( \8992 , \8990 , \8991 );
xnor \U$8650 ( \8993 , \8992 , \1960 );
and \U$8651 ( \8994 , \8989 , \8993 );
and \U$8652 ( \8995 , \3061 , \1891 );
and \U$8653 ( \8996 , \2942 , \1889 );
nor \U$8654 ( \8997 , \8995 , \8996 );
xnor \U$8655 ( \8998 , \8997 , \1739 );
and \U$8656 ( \8999 , \8993 , \8998 );
and \U$8657 ( \9000 , \8989 , \8998 );
or \U$8658 ( \9001 , \8994 , \8999 , \9000 );
and \U$8659 ( \9002 , \8985 , \9001 );
and \U$8660 ( \9003 , \1071 , \4603 );
and \U$8661 ( \9004 , \983 , \4601 );
nor \U$8662 ( \9005 , \9003 , \9004 );
xnor \U$8663 ( \9006 , \9005 , \4371 );
and \U$8664 ( \9007 , \1181 , \4152 );
and \U$8665 ( \9008 , \1176 , \4150 );
nor \U$8666 ( \9009 , \9007 , \9008 );
xnor \U$8667 ( \9010 , \9009 , \4009 );
and \U$8668 ( \9011 , \9006 , \9010 );
and \U$8669 ( \9012 , \1412 , \3829 );
and \U$8670 ( \9013 , \1297 , \3827 );
nor \U$8671 ( \9014 , \9012 , \9013 );
xnor \U$8672 ( \9015 , \9014 , \3583 );
and \U$8673 ( \9016 , \9010 , \9015 );
and \U$8674 ( \9017 , \9006 , \9015 );
or \U$8675 ( \9018 , \9011 , \9016 , \9017 );
and \U$8676 ( \9019 , \9001 , \9018 );
and \U$8677 ( \9020 , \8985 , \9018 );
or \U$8678 ( \9021 , \9002 , \9019 , \9020 );
and \U$8679 ( \9022 , \8969 , \9021 );
and \U$8680 ( \9023 , \5954 , \357 );
and \U$8681 ( \9024 , \5945 , \355 );
nor \U$8682 ( \9025 , \9023 , \9024 );
xnor \U$8683 ( \9026 , \9025 , \364 );
and \U$8684 ( \9027 , \6499 , \373 );
and \U$8685 ( \9028 , \6297 , \371 );
nor \U$8686 ( \9029 , \9027 , \9028 );
xnor \U$8687 ( \9030 , \9029 , \380 );
and \U$8688 ( \9031 , \9026 , \9030 );
and \U$8689 ( \9032 , \6974 , \391 );
and \U$8690 ( \9033 , \6802 , \389 );
nor \U$8691 ( \9034 , \9032 , \9033 );
xnor \U$8692 ( \9035 , \9034 , \398 );
and \U$8693 ( \9036 , \9030 , \9035 );
and \U$8694 ( \9037 , \9026 , \9035 );
or \U$8695 ( \9038 , \9031 , \9036 , \9037 );
and \U$8696 ( \9039 , \4576 , \957 );
and \U$8697 ( \9040 , \4568 , \955 );
nor \U$8698 ( \9041 , \9039 , \9040 );
xnor \U$8699 ( \9042 , \9041 , \879 );
and \U$8700 ( \9043 , \5050 , \793 );
and \U$8701 ( \9044 , \5045 , \791 );
nor \U$8702 ( \9045 , \9043 , \9044 );
xnor \U$8703 ( \9046 , \9045 , \699 );
and \U$8704 ( \9047 , \9042 , \9046 );
and \U$8705 ( \9048 , \5573 , \624 );
and \U$8706 ( \9049 , \5314 , \622 );
nor \U$8707 ( \9050 , \9048 , \9049 );
xnor \U$8708 ( \9051 , \9050 , \349 );
and \U$8709 ( \9052 , \9046 , \9051 );
and \U$8710 ( \9053 , \9042 , \9051 );
or \U$8711 ( \9054 , \9047 , \9052 , \9053 );
and \U$8712 ( \9055 , \9038 , \9054 );
and \U$8713 ( \9056 , \3686 , \1623 );
and \U$8714 ( \9057 , \3478 , \1621 );
nor \U$8715 ( \9058 , \9056 , \9057 );
xnor \U$8716 ( \9059 , \9058 , \1467 );
and \U$8717 ( \9060 , \3813 , \1351 );
and \U$8718 ( \9061 , \3808 , \1349 );
nor \U$8719 ( \9062 , \9060 , \9061 );
xnor \U$8720 ( \9063 , \9062 , \1238 );
and \U$8721 ( \9064 , \9059 , \9063 );
and \U$8722 ( \9065 , \4266 , \1157 );
and \U$8723 ( \9066 , \4069 , \1155 );
nor \U$8724 ( \9067 , \9065 , \9066 );
xnor \U$8725 ( \9068 , \9067 , \1021 );
and \U$8726 ( \9069 , \9063 , \9068 );
and \U$8727 ( \9070 , \9059 , \9068 );
or \U$8728 ( \9071 , \9064 , \9069 , \9070 );
and \U$8729 ( \9072 , \9054 , \9071 );
and \U$8730 ( \9073 , \9038 , \9071 );
or \U$8731 ( \9074 , \9055 , \9072 , \9073 );
and \U$8732 ( \9075 , \9021 , \9074 );
and \U$8733 ( \9076 , \8969 , \9074 );
or \U$8734 ( \9077 , \9022 , \9075 , \9076 );
and \U$8735 ( \9078 , \8915 , \9077 );
xor \U$8736 ( \9079 , \8696 , \8700 );
xor \U$8737 ( \9080 , \9079 , \8705 );
xor \U$8738 ( \9081 , \8712 , \8716 );
xor \U$8739 ( \9082 , \9081 , \8721 );
and \U$8740 ( \9083 , \9080 , \9082 );
xor \U$8741 ( \9084 , \8729 , \8733 );
xor \U$8742 ( \9085 , \9084 , \8738 );
and \U$8743 ( \9086 , \9082 , \9085 );
and \U$8744 ( \9087 , \9080 , \9085 );
or \U$8745 ( \9088 , \9083 , \9086 , \9087 );
xor \U$8746 ( \9089 , \8305 , \8309 );
xor \U$8747 ( \9090 , \9089 , \8314 );
and \U$8748 ( \9091 , \9088 , \9090 );
xor \U$8749 ( \9092 , \8323 , \8327 );
xor \U$8750 ( \9093 , \9092 , \8332 );
and \U$8751 ( \9094 , \9090 , \9093 );
and \U$8752 ( \9095 , \9088 , \9093 );
or \U$8753 ( \9096 , \9091 , \9094 , \9095 );
and \U$8754 ( \9097 , \9077 , \9096 );
and \U$8755 ( \9098 , \8915 , \9096 );
or \U$8756 ( \9099 , \9078 , \9097 , \9098 );
xor \U$8757 ( \9100 , \8600 , \8616 );
xor \U$8758 ( \9101 , \9100 , \8633 );
xor \U$8759 ( \9102 , \8652 , \8668 );
xor \U$8760 ( \9103 , \9102 , \8685 );
and \U$8761 ( \9104 , \9101 , \9103 );
xor \U$8762 ( \9105 , \8708 , \8724 );
xor \U$8763 ( \9106 , \9105 , \8741 );
and \U$8764 ( \9107 , \9103 , \9106 );
and \U$8765 ( \9108 , \9101 , \9106 );
or \U$8766 ( \9109 , \9104 , \9107 , \9108 );
xor \U$8767 ( \9110 , \8749 , \8751 );
xor \U$8768 ( \9111 , \9110 , \8754 );
xor \U$8769 ( \9112 , \8759 , \8761 );
xor \U$8770 ( \9113 , \9112 , \8764 );
and \U$8771 ( \9114 , \9111 , \9113 );
xor \U$8772 ( \9115 , \8782 , \8784 );
xor \U$8773 ( \9116 , \9115 , \8787 );
and \U$8774 ( \9117 , \9113 , \9116 );
and \U$8775 ( \9118 , \9111 , \9116 );
or \U$8776 ( \9119 , \9114 , \9117 , \9118 );
and \U$8777 ( \9120 , \9109 , \9119 );
xor \U$8778 ( \9121 , \8371 , \8387 );
xor \U$8779 ( \9122 , \9121 , \8404 );
and \U$8780 ( \9123 , \9119 , \9122 );
and \U$8781 ( \9124 , \9109 , \9122 );
or \U$8782 ( \9125 , \9120 , \9123 , \9124 );
and \U$8783 ( \9126 , \9099 , \9125 );
xor \U$8784 ( \9127 , \8317 , \8335 );
xor \U$8785 ( \9128 , \9127 , \8352 );
xor \U$8786 ( \9129 , \8796 , \8798 );
xor \U$8787 ( \9130 , \9129 , \8801 );
and \U$8788 ( \9131 , \9128 , \9130 );
xor \U$8789 ( \9132 , \8809 , \8811 );
xor \U$8790 ( \9133 , \9132 , \8814 );
and \U$8791 ( \9134 , \9130 , \9133 );
and \U$8792 ( \9135 , \9128 , \9133 );
or \U$8793 ( \9136 , \9131 , \9134 , \9135 );
and \U$8794 ( \9137 , \9125 , \9136 );
and \U$8795 ( \9138 , \9099 , \9136 );
or \U$8796 ( \9139 , \9126 , \9137 , \9138 );
xor \U$8797 ( \9140 , \8747 , \8793 );
xor \U$8798 ( \9141 , \9140 , \8804 );
xor \U$8799 ( \9142 , \8817 , \8819 );
xor \U$8800 ( \9143 , \9142 , \8822 );
and \U$8801 ( \9144 , \9141 , \9143 );
xor \U$8802 ( \9145 , \8828 , \8830 );
xor \U$8803 ( \9146 , \9145 , \8833 );
and \U$8804 ( \9147 , \9143 , \9146 );
and \U$8805 ( \9148 , \9141 , \9146 );
or \U$8806 ( \9149 , \9144 , \9147 , \9148 );
and \U$8807 ( \9150 , \9139 , \9149 );
xor \U$8808 ( \9151 , \8841 , \8843 );
xor \U$8809 ( \9152 , \9151 , \8846 );
and \U$8810 ( \9153 , \9149 , \9152 );
and \U$8811 ( \9154 , \9139 , \9152 );
or \U$8812 ( \9155 , \9150 , \9153 , \9154 );
xor \U$8813 ( \9156 , \8839 , \8849 );
xor \U$8814 ( \9157 , \9156 , \8852 );
and \U$8815 ( \9158 , \9155 , \9157 );
xor \U$8816 ( \9159 , \8857 , \8859 );
and \U$8817 ( \9160 , \9157 , \9159 );
and \U$8818 ( \9161 , \9155 , \9159 );
or \U$8819 ( \9162 , \9158 , \9160 , \9161 );
xor \U$8820 ( \9163 , \8855 , \8860 );
xor \U$8821 ( \9164 , \9163 , \8863 );
and \U$8822 ( \9165 , \9162 , \9164 );
xor \U$8823 ( \9166 , \8554 , \8564 );
xor \U$8824 ( \9167 , \9166 , \8567 );
and \U$8825 ( \9168 , \9164 , \9167 );
and \U$8826 ( \9169 , \9162 , \9167 );
or \U$8827 ( \9170 , \9165 , \9168 , \9169 );
and \U$8828 ( \9171 , \8872 , \9170 );
xor \U$8829 ( \9172 , \8872 , \9170 );
xor \U$8830 ( \9173 , \9162 , \9164 );
xor \U$8831 ( \9174 , \9173 , \9167 );
and \U$8832 ( \9175 , \5045 , \957 );
and \U$8833 ( \9176 , \4576 , \955 );
nor \U$8834 ( \9177 , \9175 , \9176 );
xnor \U$8835 ( \9178 , \9177 , \879 );
and \U$8836 ( \9179 , \5314 , \793 );
and \U$8837 ( \9180 , \5050 , \791 );
nor \U$8838 ( \9181 , \9179 , \9180 );
xnor \U$8839 ( \9182 , \9181 , \699 );
and \U$8840 ( \9183 , \9178 , \9182 );
and \U$8841 ( \9184 , \5945 , \624 );
and \U$8842 ( \9185 , \5573 , \622 );
nor \U$8843 ( \9186 , \9184 , \9185 );
xnor \U$8844 ( \9187 , \9186 , \349 );
and \U$8845 ( \9188 , \9182 , \9187 );
and \U$8846 ( \9189 , \9178 , \9187 );
or \U$8847 ( \9190 , \9183 , \9188 , \9189 );
and \U$8848 ( \9191 , \3808 , \1623 );
and \U$8849 ( \9192 , \3686 , \1621 );
nor \U$8850 ( \9193 , \9191 , \9192 );
xnor \U$8851 ( \9194 , \9193 , \1467 );
and \U$8852 ( \9195 , \4069 , \1351 );
and \U$8853 ( \9196 , \3813 , \1349 );
nor \U$8854 ( \9197 , \9195 , \9196 );
xnor \U$8855 ( \9198 , \9197 , \1238 );
and \U$8856 ( \9199 , \9194 , \9198 );
and \U$8857 ( \9200 , \4568 , \1157 );
and \U$8858 ( \9201 , \4266 , \1155 );
nor \U$8859 ( \9202 , \9200 , \9201 );
xnor \U$8860 ( \9203 , \9202 , \1021 );
and \U$8861 ( \9204 , \9198 , \9203 );
and \U$8862 ( \9205 , \9194 , \9203 );
or \U$8863 ( \9206 , \9199 , \9204 , \9205 );
and \U$8864 ( \9207 , \9190 , \9206 );
and \U$8865 ( \9208 , \6297 , \357 );
and \U$8866 ( \9209 , \5954 , \355 );
nor \U$8867 ( \9210 , \9208 , \9209 );
xnor \U$8868 ( \9211 , \9210 , \364 );
and \U$8869 ( \9212 , \6802 , \373 );
and \U$8870 ( \9213 , \6499 , \371 );
nor \U$8871 ( \9214 , \9212 , \9213 );
xnor \U$8872 ( \9215 , \9214 , \380 );
and \U$8873 ( \9216 , \9211 , \9215 );
and \U$8874 ( \9217 , \7500 , \391 );
and \U$8875 ( \9218 , \6974 , \389 );
nor \U$8876 ( \9219 , \9217 , \9218 );
xnor \U$8877 ( \9220 , \9219 , \398 );
and \U$8878 ( \9221 , \9215 , \9220 );
and \U$8879 ( \9222 , \9211 , \9220 );
or \U$8880 ( \9223 , \9216 , \9221 , \9222 );
and \U$8881 ( \9224 , \9206 , \9223 );
and \U$8882 ( \9225 , \9190 , \9223 );
or \U$8883 ( \9226 , \9207 , \9224 , \9225 );
xor \U$8884 ( \9227 , \8319 , \8916 );
xor \U$8885 ( \9228 , \8916 , \8917 );
not \U$8886 ( \9229 , \9228 );
and \U$8887 ( \9230 , \9227 , \9229 );
and \U$8888 ( \9231 , \359 , \9230 );
not \U$8889 ( \9232 , \9231 );
xnor \U$8890 ( \9233 , \9232 , \8920 );
and \U$8891 ( \9234 , \375 , \8693 );
and \U$8892 ( \9235 , \351 , \8691 );
nor \U$8893 ( \9236 , \9234 , \9235 );
xnor \U$8894 ( \9237 , \9236 , \8322 );
and \U$8895 ( \9238 , \9233 , \9237 );
and \U$8896 ( \9239 , \393 , \8131 );
and \U$8897 ( \9240 , \367 , \8129 );
nor \U$8898 ( \9241 , \9239 , \9240 );
xnor \U$8899 ( \9242 , \9241 , \7813 );
and \U$8900 ( \9243 , \9237 , \9242 );
and \U$8901 ( \9244 , \9233 , \9242 );
or \U$8902 ( \9245 , \9238 , \9243 , \9244 );
and \U$8903 ( \9246 , \450 , \6032 );
and \U$8904 ( \9247 , \435 , \6030 );
nor \U$8905 ( \9248 , \9246 , \9247 );
xnor \U$8906 ( \9249 , \9248 , \5692 );
and \U$8907 ( \9250 , \722 , \5443 );
and \U$8908 ( \9251 , \661 , \5441 );
nor \U$8909 ( \9252 , \9250 , \9251 );
xnor \U$8910 ( \9253 , \9252 , \5202 );
and \U$8911 ( \9254 , \9249 , \9253 );
and \U$8912 ( \9255 , \983 , \4977 );
and \U$8913 ( \9256 , \785 , \4975 );
nor \U$8914 ( \9257 , \9255 , \9256 );
xnor \U$8915 ( \9258 , \9257 , \4789 );
and \U$8916 ( \9259 , \9253 , \9258 );
and \U$8917 ( \9260 , \9249 , \9258 );
or \U$8918 ( \9261 , \9254 , \9259 , \9260 );
and \U$8919 ( \9262 , \9245 , \9261 );
and \U$8920 ( \9263 , \408 , \7564 );
and \U$8921 ( \9264 , \385 , \7562 );
nor \U$8922 ( \9265 , \9263 , \9264 );
xnor \U$8923 ( \9266 , \9265 , \7315 );
and \U$8924 ( \9267 , \424 , \7035 );
and \U$8925 ( \9268 , \400 , \7033 );
nor \U$8926 ( \9269 , \9267 , \9268 );
xnor \U$8927 ( \9270 , \9269 , \6775 );
and \U$8928 ( \9271 , \9266 , \9270 );
and \U$8929 ( \9272 , \443 , \6541 );
and \U$8930 ( \9273 , \416 , \6539 );
nor \U$8931 ( \9274 , \9272 , \9273 );
xnor \U$8932 ( \9275 , \9274 , \6226 );
and \U$8933 ( \9276 , \9270 , \9275 );
and \U$8934 ( \9277 , \9266 , \9275 );
or \U$8935 ( \9278 , \9271 , \9276 , \9277 );
and \U$8936 ( \9279 , \9261 , \9278 );
and \U$8937 ( \9280 , \9245 , \9278 );
or \U$8938 ( \9281 , \9262 , \9279 , \9280 );
and \U$8939 ( \9282 , \9226 , \9281 );
and \U$8940 ( \9283 , \1176 , \4603 );
and \U$8941 ( \9284 , \1071 , \4601 );
nor \U$8942 ( \9285 , \9283 , \9284 );
xnor \U$8943 ( \9286 , \9285 , \4371 );
and \U$8944 ( \9287 , \1297 , \4152 );
and \U$8945 ( \9288 , \1181 , \4150 );
nor \U$8946 ( \9289 , \9287 , \9288 );
xnor \U$8947 ( \9290 , \9289 , \4009 );
and \U$8948 ( \9291 , \9286 , \9290 );
and \U$8949 ( \9292 , \1588 , \3829 );
and \U$8950 ( \9293 , \1412 , \3827 );
nor \U$8951 ( \9294 , \9292 , \9293 );
xnor \U$8952 ( \9295 , \9294 , \3583 );
and \U$8953 ( \9296 , \9290 , \9295 );
and \U$8954 ( \9297 , \9286 , \9295 );
or \U$8955 ( \9298 , \9291 , \9296 , \9297 );
and \U$8956 ( \9299 , \2637 , \2393 );
and \U$8957 ( \9300 , \2463 , \2391 );
nor \U$8958 ( \9301 , \9299 , \9300 );
xnor \U$8959 ( \9302 , \9301 , \2251 );
and \U$8960 ( \9303 , \2942 , \2097 );
and \U$8961 ( \9304 , \2804 , \2095 );
nor \U$8962 ( \9305 , \9303 , \9304 );
xnor \U$8963 ( \9306 , \9305 , \1960 );
and \U$8964 ( \9307 , \9302 , \9306 );
and \U$8965 ( \9308 , \3478 , \1891 );
and \U$8966 ( \9309 , \3061 , \1889 );
nor \U$8967 ( \9310 , \9308 , \9309 );
xnor \U$8968 ( \9311 , \9310 , \1739 );
and \U$8969 ( \9312 , \9306 , \9311 );
and \U$8970 ( \9313 , \9302 , \9311 );
or \U$8971 ( \9314 , \9307 , \9312 , \9313 );
and \U$8972 ( \9315 , \9298 , \9314 );
and \U$8973 ( \9316 , \1839 , \3434 );
and \U$8974 ( \9317 , \1596 , \3432 );
nor \U$8975 ( \9318 , \9316 , \9317 );
xnor \U$8976 ( \9319 , \9318 , \3247 );
and \U$8977 ( \9320 , \2030 , \3121 );
and \U$8978 ( \9321 , \1844 , \3119 );
nor \U$8979 ( \9322 , \9320 , \9321 );
xnor \U$8980 ( \9323 , \9322 , \2916 );
and \U$8981 ( \9324 , \9319 , \9323 );
and \U$8982 ( \9325 , \2438 , \2715 );
and \U$8983 ( \9326 , \2174 , \2713 );
nor \U$8984 ( \9327 , \9325 , \9326 );
xnor \U$8985 ( \9328 , \9327 , \2566 );
and \U$8986 ( \9329 , \9323 , \9328 );
and \U$8987 ( \9330 , \9319 , \9328 );
or \U$8988 ( \9331 , \9324 , \9329 , \9330 );
and \U$8989 ( \9332 , \9314 , \9331 );
and \U$8990 ( \9333 , \9298 , \9331 );
or \U$8991 ( \9334 , \9315 , \9332 , \9333 );
and \U$8992 ( \9335 , \9281 , \9334 );
and \U$8993 ( \9336 , \9226 , \9334 );
or \U$8994 ( \9337 , \9282 , \9335 , \9336 );
and \U$8995 ( \9338 , \8170 , \406 );
and \U$8996 ( \9339 , \7924 , \404 );
nor \U$8997 ( \9340 , \9338 , \9339 );
xnor \U$8998 ( \9341 , \9340 , \413 );
and \U$8999 ( \9342 , \8494 , \422 );
and \U$9000 ( \9343 , \8175 , \420 );
nor \U$9001 ( \9344 , \9342 , \9343 );
xnor \U$9002 ( \9345 , \9344 , \429 );
and \U$9003 ( \9346 , \9341 , \9345 );
buf \U$9004 ( \9347 , RIbb2bce0_123);
and \U$9005 ( \9348 , \9347 , \441 );
and \U$9006 ( \9349 , \8778 , \439 );
nor \U$9007 ( \9350 , \9348 , \9349 );
xnor \U$9008 ( \9351 , \9350 , \448 );
and \U$9009 ( \9352 , \9345 , \9351 );
and \U$9010 ( \9353 , \9341 , \9351 );
or \U$9011 ( \9354 , \9346 , \9352 , \9353 );
buf \U$9012 ( \9355 , RIbb2bc68_124);
and \U$9013 ( \9356 , \9355 , \436 );
buf \U$9014 ( \9357 , \9356 );
and \U$9015 ( \9358 , \9354 , \9357 );
and \U$9016 ( \9359 , \9347 , \436 );
and \U$9017 ( \9360 , \9357 , \9359 );
and \U$9018 ( \9361 , \9354 , \9359 );
or \U$9019 ( \9362 , \9358 , \9360 , \9361 );
xor \U$9020 ( \9363 , \8897 , \8901 );
xor \U$9021 ( \9364 , \9363 , \8906 );
xor \U$9022 ( \9365 , \9026 , \9030 );
xor \U$9023 ( \9366 , \9365 , \9035 );
and \U$9024 ( \9367 , \9364 , \9366 );
xor \U$9025 ( \9368 , \9042 , \9046 );
xor \U$9026 ( \9369 , \9368 , \9051 );
and \U$9027 ( \9370 , \9366 , \9369 );
and \U$9028 ( \9371 , \9364 , \9369 );
or \U$9029 ( \9372 , \9367 , \9370 , \9371 );
and \U$9030 ( \9373 , \9362 , \9372 );
xor \U$9031 ( \9374 , \9059 , \9063 );
xor \U$9032 ( \9375 , \9374 , \9068 );
xor \U$9033 ( \9376 , \8973 , \8977 );
xor \U$9034 ( \9377 , \9376 , \8982 );
and \U$9035 ( \9378 , \9375 , \9377 );
xor \U$9036 ( \9379 , \8989 , \8993 );
xor \U$9037 ( \9380 , \9379 , \8998 );
and \U$9038 ( \9381 , \9377 , \9380 );
and \U$9039 ( \9382 , \9375 , \9380 );
or \U$9040 ( \9383 , \9378 , \9381 , \9382 );
and \U$9041 ( \9384 , \9372 , \9383 );
and \U$9042 ( \9385 , \9362 , \9383 );
or \U$9043 ( \9386 , \9373 , \9384 , \9385 );
and \U$9044 ( \9387 , \9337 , \9386 );
xor \U$9045 ( \9388 , \8937 , \8941 );
xor \U$9046 ( \9389 , \9388 , \8946 );
xor \U$9047 ( \9390 , \8954 , \8958 );
xor \U$9048 ( \9391 , \9390 , \8963 );
and \U$9049 ( \9392 , \9389 , \9391 );
xor \U$9050 ( \9393 , \9006 , \9010 );
xor \U$9051 ( \9394 , \9393 , \9015 );
and \U$9052 ( \9395 , \9391 , \9394 );
and \U$9053 ( \9396 , \9389 , \9394 );
or \U$9054 ( \9397 , \9392 , \9395 , \9396 );
xor \U$9055 ( \9398 , \9080 , \9082 );
xor \U$9056 ( \9399 , \9398 , \9085 );
and \U$9057 ( \9400 , \9397 , \9399 );
xor \U$9058 ( \9401 , \8884 , \8886 );
xor \U$9059 ( \9402 , \9401 , \8889 );
and \U$9060 ( \9403 , \9399 , \9402 );
and \U$9061 ( \9404 , \9397 , \9402 );
or \U$9062 ( \9405 , \9400 , \9403 , \9404 );
and \U$9063 ( \9406 , \9386 , \9405 );
and \U$9064 ( \9407 , \9337 , \9405 );
or \U$9065 ( \9408 , \9387 , \9406 , \9407 );
xor \U$9066 ( \9409 , \8882 , \8892 );
xor \U$9067 ( \9410 , \9409 , \8912 );
xor \U$9068 ( \9411 , \8969 , \9021 );
xor \U$9069 ( \9412 , \9411 , \9074 );
and \U$9070 ( \9413 , \9410 , \9412 );
xor \U$9071 ( \9414 , \9088 , \9090 );
xor \U$9072 ( \9415 , \9414 , \9093 );
and \U$9073 ( \9416 , \9412 , \9415 );
and \U$9074 ( \9417 , \9410 , \9415 );
or \U$9075 ( \9418 , \9413 , \9416 , \9417 );
and \U$9076 ( \9419 , \9408 , \9418 );
xor \U$9077 ( \9420 , \9038 , \9054 );
xor \U$9078 ( \9421 , \9420 , \9071 );
xor \U$9079 ( \9422 , \8874 , \8876 );
xor \U$9080 ( \9423 , \9422 , \8879 );
and \U$9081 ( \9424 , \9421 , \9423 );
xnor \U$9082 ( \9425 , \8909 , \8911 );
and \U$9083 ( \9426 , \9423 , \9425 );
and \U$9084 ( \9427 , \9421 , \9425 );
or \U$9085 ( \9428 , \9424 , \9426 , \9427 );
xor \U$9086 ( \9429 , \9101 , \9103 );
xor \U$9087 ( \9430 , \9429 , \9106 );
and \U$9088 ( \9431 , \9428 , \9430 );
xor \U$9089 ( \9432 , \9111 , \9113 );
xor \U$9090 ( \9433 , \9432 , \9116 );
and \U$9091 ( \9434 , \9430 , \9433 );
and \U$9092 ( \9435 , \9428 , \9433 );
or \U$9093 ( \9436 , \9431 , \9434 , \9435 );
and \U$9094 ( \9437 , \9418 , \9436 );
and \U$9095 ( \9438 , \9408 , \9436 );
or \U$9096 ( \9439 , \9419 , \9437 , \9438 );
xor \U$9097 ( \9440 , \8636 , \8688 );
xor \U$9098 ( \9441 , \9440 , \8744 );
xor \U$9099 ( \9442 , \8757 , \8767 );
xor \U$9100 ( \9443 , \9442 , \8790 );
and \U$9101 ( \9444 , \9441 , \9443 );
xor \U$9102 ( \9445 , \9128 , \9130 );
xor \U$9103 ( \9446 , \9445 , \9133 );
and \U$9104 ( \9447 , \9443 , \9446 );
and \U$9105 ( \9448 , \9441 , \9446 );
or \U$9106 ( \9449 , \9444 , \9447 , \9448 );
and \U$9107 ( \9450 , \9439 , \9449 );
xor \U$9108 ( \9451 , \9141 , \9143 );
xor \U$9109 ( \9452 , \9451 , \9146 );
and \U$9110 ( \9453 , \9449 , \9452 );
and \U$9111 ( \9454 , \9439 , \9452 );
or \U$9112 ( \9455 , \9450 , \9453 , \9454 );
xor \U$9113 ( \9456 , \8807 , \8825 );
xor \U$9114 ( \9457 , \9456 , \8836 );
and \U$9115 ( \9458 , \9455 , \9457 );
xor \U$9116 ( \9459 , \9139 , \9149 );
xor \U$9117 ( \9460 , \9459 , \9152 );
and \U$9118 ( \9461 , \9457 , \9460 );
and \U$9119 ( \9462 , \9455 , \9460 );
or \U$9120 ( \9463 , \9458 , \9461 , \9462 );
xor \U$9121 ( \9464 , \9155 , \9157 );
xor \U$9122 ( \9465 , \9464 , \9159 );
and \U$9123 ( \9466 , \9463 , \9465 );
and \U$9124 ( \9467 , \9174 , \9466 );
xor \U$9125 ( \9468 , \9174 , \9466 );
xor \U$9126 ( \9469 , \9463 , \9465 );
and \U$9127 ( \9470 , \2463 , \2715 );
and \U$9128 ( \9471 , \2438 , \2713 );
nor \U$9129 ( \9472 , \9470 , \9471 );
xnor \U$9130 ( \9473 , \9472 , \2566 );
and \U$9131 ( \9474 , \2804 , \2393 );
and \U$9132 ( \9475 , \2637 , \2391 );
nor \U$9133 ( \9476 , \9474 , \9475 );
xnor \U$9134 ( \9477 , \9476 , \2251 );
and \U$9135 ( \9478 , \9473 , \9477 );
and \U$9136 ( \9479 , \3061 , \2097 );
and \U$9137 ( \9480 , \2942 , \2095 );
nor \U$9138 ( \9481 , \9479 , \9480 );
xnor \U$9139 ( \9482 , \9481 , \1960 );
and \U$9140 ( \9483 , \9477 , \9482 );
and \U$9141 ( \9484 , \9473 , \9482 );
or \U$9142 ( \9485 , \9478 , \9483 , \9484 );
and \U$9143 ( \9486 , \1596 , \3829 );
and \U$9144 ( \9487 , \1588 , \3827 );
nor \U$9145 ( \9488 , \9486 , \9487 );
xnor \U$9146 ( \9489 , \9488 , \3583 );
and \U$9147 ( \9490 , \1844 , \3434 );
and \U$9148 ( \9491 , \1839 , \3432 );
nor \U$9149 ( \9492 , \9490 , \9491 );
xnor \U$9150 ( \9493 , \9492 , \3247 );
and \U$9151 ( \9494 , \9489 , \9493 );
and \U$9152 ( \9495 , \2174 , \3121 );
and \U$9153 ( \9496 , \2030 , \3119 );
nor \U$9154 ( \9497 , \9495 , \9496 );
xnor \U$9155 ( \9498 , \9497 , \2916 );
and \U$9156 ( \9499 , \9493 , \9498 );
and \U$9157 ( \9500 , \9489 , \9498 );
or \U$9158 ( \9501 , \9494 , \9499 , \9500 );
and \U$9159 ( \9502 , \9485 , \9501 );
and \U$9160 ( \9503 , \1071 , \4977 );
and \U$9161 ( \9504 , \983 , \4975 );
nor \U$9162 ( \9505 , \9503 , \9504 );
xnor \U$9163 ( \9506 , \9505 , \4789 );
and \U$9164 ( \9507 , \1181 , \4603 );
and \U$9165 ( \9508 , \1176 , \4601 );
nor \U$9166 ( \9509 , \9507 , \9508 );
xnor \U$9167 ( \9510 , \9509 , \4371 );
and \U$9168 ( \9511 , \9506 , \9510 );
and \U$9169 ( \9512 , \1412 , \4152 );
and \U$9170 ( \9513 , \1297 , \4150 );
nor \U$9171 ( \9514 , \9512 , \9513 );
xnor \U$9172 ( \9515 , \9514 , \4009 );
and \U$9173 ( \9516 , \9510 , \9515 );
and \U$9174 ( \9517 , \9506 , \9515 );
or \U$9175 ( \9518 , \9511 , \9516 , \9517 );
and \U$9176 ( \9519 , \9501 , \9518 );
and \U$9177 ( \9520 , \9485 , \9518 );
or \U$9178 ( \9521 , \9502 , \9519 , \9520 );
and \U$9179 ( \9522 , \435 , \6541 );
and \U$9180 ( \9523 , \443 , \6539 );
nor \U$9181 ( \9524 , \9522 , \9523 );
xnor \U$9182 ( \9525 , \9524 , \6226 );
and \U$9183 ( \9526 , \661 , \6032 );
and \U$9184 ( \9527 , \450 , \6030 );
nor \U$9185 ( \9528 , \9526 , \9527 );
xnor \U$9186 ( \9529 , \9528 , \5692 );
and \U$9187 ( \9530 , \9525 , \9529 );
and \U$9188 ( \9531 , \785 , \5443 );
and \U$9189 ( \9532 , \722 , \5441 );
nor \U$9190 ( \9533 , \9531 , \9532 );
xnor \U$9191 ( \9534 , \9533 , \5202 );
and \U$9192 ( \9535 , \9529 , \9534 );
and \U$9193 ( \9536 , \9525 , \9534 );
or \U$9194 ( \9537 , \9530 , \9535 , \9536 );
and \U$9195 ( \9538 , \385 , \8131 );
and \U$9196 ( \9539 , \393 , \8129 );
nor \U$9197 ( \9540 , \9538 , \9539 );
xnor \U$9198 ( \9541 , \9540 , \7813 );
and \U$9199 ( \9542 , \400 , \7564 );
and \U$9200 ( \9543 , \408 , \7562 );
nor \U$9201 ( \9544 , \9542 , \9543 );
xnor \U$9202 ( \9545 , \9544 , \7315 );
and \U$9203 ( \9546 , \9541 , \9545 );
and \U$9204 ( \9547 , \416 , \7035 );
and \U$9205 ( \9548 , \424 , \7033 );
nor \U$9206 ( \9549 , \9547 , \9548 );
xnor \U$9207 ( \9550 , \9549 , \6775 );
and \U$9208 ( \9551 , \9545 , \9550 );
and \U$9209 ( \9552 , \9541 , \9550 );
or \U$9210 ( \9553 , \9546 , \9551 , \9552 );
and \U$9211 ( \9554 , \9537 , \9553 );
buf \U$9212 ( \9555 , RIbb2d978_62);
buf \U$9213 ( \9556 , RIbb2d900_63);
and \U$9214 ( \9557 , \9555 , \9556 );
not \U$9215 ( \9558 , \9557 );
and \U$9216 ( \9559 , \8917 , \9558 );
not \U$9217 ( \9560 , \9559 );
and \U$9218 ( \9561 , \351 , \9230 );
and \U$9219 ( \9562 , \359 , \9228 );
nor \U$9220 ( \9563 , \9561 , \9562 );
xnor \U$9221 ( \9564 , \9563 , \8920 );
and \U$9222 ( \9565 , \9560 , \9564 );
and \U$9223 ( \9566 , \367 , \8693 );
and \U$9224 ( \9567 , \375 , \8691 );
nor \U$9225 ( \9568 , \9566 , \9567 );
xnor \U$9226 ( \9569 , \9568 , \8322 );
and \U$9227 ( \9570 , \9564 , \9569 );
and \U$9228 ( \9571 , \9560 , \9569 );
or \U$9229 ( \9572 , \9565 , \9570 , \9571 );
and \U$9230 ( \9573 , \9553 , \9572 );
and \U$9231 ( \9574 , \9537 , \9572 );
or \U$9232 ( \9575 , \9554 , \9573 , \9574 );
and \U$9233 ( \9576 , \9521 , \9575 );
and \U$9234 ( \9577 , \5954 , \624 );
and \U$9235 ( \9578 , \5945 , \622 );
nor \U$9236 ( \9579 , \9577 , \9578 );
xnor \U$9237 ( \9580 , \9579 , \349 );
and \U$9238 ( \9581 , \6499 , \357 );
and \U$9239 ( \9582 , \6297 , \355 );
nor \U$9240 ( \9583 , \9581 , \9582 );
xnor \U$9241 ( \9584 , \9583 , \364 );
and \U$9242 ( \9585 , \9580 , \9584 );
and \U$9243 ( \9586 , \6974 , \373 );
and \U$9244 ( \9587 , \6802 , \371 );
nor \U$9245 ( \9588 , \9586 , \9587 );
xnor \U$9246 ( \9589 , \9588 , \380 );
and \U$9247 ( \9590 , \9584 , \9589 );
and \U$9248 ( \9591 , \9580 , \9589 );
or \U$9249 ( \9592 , \9585 , \9590 , \9591 );
and \U$9250 ( \9593 , \4576 , \1157 );
and \U$9251 ( \9594 , \4568 , \1155 );
nor \U$9252 ( \9595 , \9593 , \9594 );
xnor \U$9253 ( \9596 , \9595 , \1021 );
and \U$9254 ( \9597 , \5050 , \957 );
and \U$9255 ( \9598 , \5045 , \955 );
nor \U$9256 ( \9599 , \9597 , \9598 );
xnor \U$9257 ( \9600 , \9599 , \879 );
and \U$9258 ( \9601 , \9596 , \9600 );
and \U$9259 ( \9602 , \5573 , \793 );
and \U$9260 ( \9603 , \5314 , \791 );
nor \U$9261 ( \9604 , \9602 , \9603 );
xnor \U$9262 ( \9605 , \9604 , \699 );
and \U$9263 ( \9606 , \9600 , \9605 );
and \U$9264 ( \9607 , \9596 , \9605 );
or \U$9265 ( \9608 , \9601 , \9606 , \9607 );
and \U$9266 ( \9609 , \9592 , \9608 );
and \U$9267 ( \9610 , \3686 , \1891 );
and \U$9268 ( \9611 , \3478 , \1889 );
nor \U$9269 ( \9612 , \9610 , \9611 );
xnor \U$9270 ( \9613 , \9612 , \1739 );
and \U$9271 ( \9614 , \3813 , \1623 );
and \U$9272 ( \9615 , \3808 , \1621 );
nor \U$9273 ( \9616 , \9614 , \9615 );
xnor \U$9274 ( \9617 , \9616 , \1467 );
and \U$9275 ( \9618 , \9613 , \9617 );
and \U$9276 ( \9619 , \4266 , \1351 );
and \U$9277 ( \9620 , \4069 , \1349 );
nor \U$9278 ( \9621 , \9619 , \9620 );
xnor \U$9279 ( \9622 , \9621 , \1238 );
and \U$9280 ( \9623 , \9617 , \9622 );
and \U$9281 ( \9624 , \9613 , \9622 );
or \U$9282 ( \9625 , \9618 , \9623 , \9624 );
and \U$9283 ( \9626 , \9608 , \9625 );
and \U$9284 ( \9627 , \9592 , \9625 );
or \U$9285 ( \9628 , \9609 , \9626 , \9627 );
and \U$9286 ( \9629 , \9575 , \9628 );
and \U$9287 ( \9630 , \9521 , \9628 );
or \U$9288 ( \9631 , \9576 , \9629 , \9630 );
xor \U$9289 ( \9632 , \9286 , \9290 );
xor \U$9290 ( \9633 , \9632 , \9295 );
xor \U$9291 ( \9634 , \9302 , \9306 );
xor \U$9292 ( \9635 , \9634 , \9311 );
and \U$9293 ( \9636 , \9633 , \9635 );
xor \U$9294 ( \9637 , \9319 , \9323 );
xor \U$9295 ( \9638 , \9637 , \9328 );
and \U$9296 ( \9639 , \9635 , \9638 );
and \U$9297 ( \9640 , \9633 , \9638 );
or \U$9298 ( \9641 , \9636 , \9639 , \9640 );
xor \U$9299 ( \9642 , \9178 , \9182 );
xor \U$9300 ( \9643 , \9642 , \9187 );
xor \U$9301 ( \9644 , \9194 , \9198 );
xor \U$9302 ( \9645 , \9644 , \9203 );
and \U$9303 ( \9646 , \9643 , \9645 );
xor \U$9304 ( \9647 , \9211 , \9215 );
xor \U$9305 ( \9648 , \9647 , \9220 );
and \U$9306 ( \9649 , \9645 , \9648 );
and \U$9307 ( \9650 , \9643 , \9648 );
or \U$9308 ( \9651 , \9646 , \9649 , \9650 );
and \U$9309 ( \9652 , \9641 , \9651 );
and \U$9310 ( \9653 , \7924 , \391 );
and \U$9311 ( \9654 , \7500 , \389 );
nor \U$9312 ( \9655 , \9653 , \9654 );
xnor \U$9313 ( \9656 , \9655 , \398 );
and \U$9314 ( \9657 , \8175 , \406 );
and \U$9315 ( \9658 , \8170 , \404 );
nor \U$9316 ( \9659 , \9657 , \9658 );
xnor \U$9317 ( \9660 , \9659 , \413 );
and \U$9318 ( \9661 , \9656 , \9660 );
and \U$9319 ( \9662 , \8778 , \422 );
and \U$9320 ( \9663 , \8494 , \420 );
nor \U$9321 ( \9664 , \9662 , \9663 );
xnor \U$9322 ( \9665 , \9664 , \429 );
and \U$9323 ( \9666 , \9660 , \9665 );
and \U$9324 ( \9667 , \9656 , \9665 );
or \U$9325 ( \9668 , \9661 , \9666 , \9667 );
xor \U$9326 ( \9669 , \9341 , \9345 );
xor \U$9327 ( \9670 , \9669 , \9351 );
and \U$9328 ( \9671 , \9668 , \9670 );
not \U$9329 ( \9672 , \9356 );
and \U$9330 ( \9673 , \9670 , \9672 );
and \U$9331 ( \9674 , \9668 , \9672 );
or \U$9332 ( \9675 , \9671 , \9673 , \9674 );
and \U$9333 ( \9676 , \9651 , \9675 );
and \U$9334 ( \9677 , \9641 , \9675 );
or \U$9335 ( \9678 , \9652 , \9676 , \9677 );
and \U$9336 ( \9679 , \9631 , \9678 );
xor \U$9337 ( \9680 , \9233 , \9237 );
xor \U$9338 ( \9681 , \9680 , \9242 );
xor \U$9339 ( \9682 , \9249 , \9253 );
xor \U$9340 ( \9683 , \9682 , \9258 );
and \U$9341 ( \9684 , \9681 , \9683 );
xor \U$9342 ( \9685 , \9266 , \9270 );
xor \U$9343 ( \9686 , \9685 , \9275 );
and \U$9344 ( \9687 , \9683 , \9686 );
and \U$9345 ( \9688 , \9681 , \9686 );
or \U$9346 ( \9689 , \9684 , \9687 , \9688 );
xor \U$9347 ( \9690 , \8921 , \8925 );
xor \U$9348 ( \9691 , \9690 , \8930 );
and \U$9349 ( \9692 , \9689 , \9691 );
xor \U$9350 ( \9693 , \9389 , \9391 );
xor \U$9351 ( \9694 , \9693 , \9394 );
and \U$9352 ( \9695 , \9691 , \9694 );
and \U$9353 ( \9696 , \9689 , \9694 );
or \U$9354 ( \9697 , \9692 , \9695 , \9696 );
and \U$9355 ( \9698 , \9678 , \9697 );
and \U$9356 ( \9699 , \9631 , \9697 );
or \U$9357 ( \9700 , \9679 , \9698 , \9699 );
xor \U$9358 ( \9701 , \9190 , \9206 );
xor \U$9359 ( \9702 , \9701 , \9223 );
xor \U$9360 ( \9703 , \9245 , \9261 );
xor \U$9361 ( \9704 , \9703 , \9278 );
and \U$9362 ( \9705 , \9702 , \9704 );
xor \U$9363 ( \9706 , \9298 , \9314 );
xor \U$9364 ( \9707 , \9706 , \9331 );
and \U$9365 ( \9708 , \9704 , \9707 );
and \U$9366 ( \9709 , \9702 , \9707 );
or \U$9367 ( \9710 , \9705 , \9708 , \9709 );
xor \U$9368 ( \9711 , \9354 , \9357 );
xor \U$9369 ( \9712 , \9711 , \9359 );
xor \U$9370 ( \9713 , \9364 , \9366 );
xor \U$9371 ( \9714 , \9713 , \9369 );
and \U$9372 ( \9715 , \9712 , \9714 );
xor \U$9373 ( \9716 , \9375 , \9377 );
xor \U$9374 ( \9717 , \9716 , \9380 );
and \U$9375 ( \9718 , \9714 , \9717 );
and \U$9376 ( \9719 , \9712 , \9717 );
or \U$9377 ( \9720 , \9715 , \9718 , \9719 );
and \U$9378 ( \9721 , \9710 , \9720 );
xor \U$9379 ( \9722 , \8985 , \9001 );
xor \U$9380 ( \9723 , \9722 , \9018 );
and \U$9381 ( \9724 , \9720 , \9723 );
and \U$9382 ( \9725 , \9710 , \9723 );
or \U$9383 ( \9726 , \9721 , \9724 , \9725 );
and \U$9384 ( \9727 , \9700 , \9726 );
xor \U$9385 ( \9728 , \8933 , \8949 );
xor \U$9386 ( \9729 , \9728 , \8966 );
xor \U$9387 ( \9730 , \9397 , \9399 );
xor \U$9388 ( \9731 , \9730 , \9402 );
and \U$9389 ( \9732 , \9729 , \9731 );
xor \U$9390 ( \9733 , \9421 , \9423 );
xor \U$9391 ( \9734 , \9733 , \9425 );
and \U$9392 ( \9735 , \9731 , \9734 );
and \U$9393 ( \9736 , \9729 , \9734 );
or \U$9394 ( \9737 , \9732 , \9735 , \9736 );
and \U$9395 ( \9738 , \9726 , \9737 );
and \U$9396 ( \9739 , \9700 , \9737 );
or \U$9397 ( \9740 , \9727 , \9738 , \9739 );
xor \U$9398 ( \9741 , \9337 , \9386 );
xor \U$9399 ( \9742 , \9741 , \9405 );
xor \U$9400 ( \9743 , \9410 , \9412 );
xor \U$9401 ( \9744 , \9743 , \9415 );
and \U$9402 ( \9745 , \9742 , \9744 );
xor \U$9403 ( \9746 , \9428 , \9430 );
xor \U$9404 ( \9747 , \9746 , \9433 );
and \U$9405 ( \9748 , \9744 , \9747 );
and \U$9406 ( \9749 , \9742 , \9747 );
or \U$9407 ( \9750 , \9745 , \9748 , \9749 );
and \U$9408 ( \9751 , \9740 , \9750 );
xor \U$9409 ( \9752 , \9109 , \9119 );
xor \U$9410 ( \9753 , \9752 , \9122 );
and \U$9411 ( \9754 , \9750 , \9753 );
and \U$9412 ( \9755 , \9740 , \9753 );
or \U$9413 ( \9756 , \9751 , \9754 , \9755 );
xor \U$9414 ( \9757 , \8915 , \9077 );
xor \U$9415 ( \9758 , \9757 , \9096 );
xor \U$9416 ( \9759 , \9408 , \9418 );
xor \U$9417 ( \9760 , \9759 , \9436 );
and \U$9418 ( \9761 , \9758 , \9760 );
xor \U$9419 ( \9762 , \9441 , \9443 );
xor \U$9420 ( \9763 , \9762 , \9446 );
and \U$9421 ( \9764 , \9760 , \9763 );
and \U$9422 ( \9765 , \9758 , \9763 );
or \U$9423 ( \9766 , \9761 , \9764 , \9765 );
and \U$9424 ( \9767 , \9756 , \9766 );
xor \U$9425 ( \9768 , \9099 , \9125 );
xor \U$9426 ( \9769 , \9768 , \9136 );
and \U$9427 ( \9770 , \9766 , \9769 );
and \U$9428 ( \9771 , \9756 , \9769 );
or \U$9429 ( \9772 , \9767 , \9770 , \9771 );
xor \U$9430 ( \9773 , \9455 , \9457 );
xor \U$9431 ( \9774 , \9773 , \9460 );
and \U$9432 ( \9775 , \9772 , \9774 );
and \U$9433 ( \9776 , \9469 , \9775 );
xor \U$9434 ( \9777 , \9469 , \9775 );
xor \U$9435 ( \9778 , \9772 , \9774 );
and \U$9436 ( \9779 , \450 , \6541 );
and \U$9437 ( \9780 , \435 , \6539 );
nor \U$9438 ( \9781 , \9779 , \9780 );
xnor \U$9439 ( \9782 , \9781 , \6226 );
and \U$9440 ( \9783 , \722 , \6032 );
and \U$9441 ( \9784 , \661 , \6030 );
nor \U$9442 ( \9785 , \9783 , \9784 );
xnor \U$9443 ( \9786 , \9785 , \5692 );
and \U$9444 ( \9787 , \9782 , \9786 );
and \U$9445 ( \9788 , \983 , \5443 );
and \U$9446 ( \9789 , \785 , \5441 );
nor \U$9447 ( \9790 , \9788 , \9789 );
xnor \U$9448 ( \9791 , \9790 , \5202 );
and \U$9449 ( \9792 , \9786 , \9791 );
and \U$9450 ( \9793 , \9782 , \9791 );
or \U$9451 ( \9794 , \9787 , \9792 , \9793 );
xor \U$9452 ( \9795 , \8917 , \9555 );
xor \U$9453 ( \9796 , \9555 , \9556 );
not \U$9454 ( \9797 , \9796 );
and \U$9455 ( \9798 , \9795 , \9797 );
and \U$9456 ( \9799 , \359 , \9798 );
not \U$9457 ( \9800 , \9799 );
xnor \U$9458 ( \9801 , \9800 , \9559 );
and \U$9459 ( \9802 , \375 , \9230 );
and \U$9460 ( \9803 , \351 , \9228 );
nor \U$9461 ( \9804 , \9802 , \9803 );
xnor \U$9462 ( \9805 , \9804 , \8920 );
and \U$9463 ( \9806 , \9801 , \9805 );
and \U$9464 ( \9807 , \393 , \8693 );
and \U$9465 ( \9808 , \367 , \8691 );
nor \U$9466 ( \9809 , \9807 , \9808 );
xnor \U$9467 ( \9810 , \9809 , \8322 );
and \U$9468 ( \9811 , \9805 , \9810 );
and \U$9469 ( \9812 , \9801 , \9810 );
or \U$9470 ( \9813 , \9806 , \9811 , \9812 );
and \U$9471 ( \9814 , \9794 , \9813 );
and \U$9472 ( \9815 , \408 , \8131 );
and \U$9473 ( \9816 , \385 , \8129 );
nor \U$9474 ( \9817 , \9815 , \9816 );
xnor \U$9475 ( \9818 , \9817 , \7813 );
and \U$9476 ( \9819 , \424 , \7564 );
and \U$9477 ( \9820 , \400 , \7562 );
nor \U$9478 ( \9821 , \9819 , \9820 );
xnor \U$9479 ( \9822 , \9821 , \7315 );
and \U$9480 ( \9823 , \9818 , \9822 );
and \U$9481 ( \9824 , \443 , \7035 );
and \U$9482 ( \9825 , \416 , \7033 );
nor \U$9483 ( \9826 , \9824 , \9825 );
xnor \U$9484 ( \9827 , \9826 , \6775 );
and \U$9485 ( \9828 , \9822 , \9827 );
and \U$9486 ( \9829 , \9818 , \9827 );
or \U$9487 ( \9830 , \9823 , \9828 , \9829 );
and \U$9488 ( \9831 , \9813 , \9830 );
and \U$9489 ( \9832 , \9794 , \9830 );
or \U$9490 ( \9833 , \9814 , \9831 , \9832 );
and \U$9491 ( \9834 , \6297 , \624 );
and \U$9492 ( \9835 , \5954 , \622 );
nor \U$9493 ( \9836 , \9834 , \9835 );
xnor \U$9494 ( \9837 , \9836 , \349 );
and \U$9495 ( \9838 , \6802 , \357 );
and \U$9496 ( \9839 , \6499 , \355 );
nor \U$9497 ( \9840 , \9838 , \9839 );
xnor \U$9498 ( \9841 , \9840 , \364 );
and \U$9499 ( \9842 , \9837 , \9841 );
and \U$9500 ( \9843 , \7500 , \373 );
and \U$9501 ( \9844 , \6974 , \371 );
nor \U$9502 ( \9845 , \9843 , \9844 );
xnor \U$9503 ( \9846 , \9845 , \380 );
and \U$9504 ( \9847 , \9841 , \9846 );
and \U$9505 ( \9848 , \9837 , \9846 );
or \U$9506 ( \9849 , \9842 , \9847 , \9848 );
and \U$9507 ( \9850 , \3808 , \1891 );
and \U$9508 ( \9851 , \3686 , \1889 );
nor \U$9509 ( \9852 , \9850 , \9851 );
xnor \U$9510 ( \9853 , \9852 , \1739 );
and \U$9511 ( \9854 , \4069 , \1623 );
and \U$9512 ( \9855 , \3813 , \1621 );
nor \U$9513 ( \9856 , \9854 , \9855 );
xnor \U$9514 ( \9857 , \9856 , \1467 );
and \U$9515 ( \9858 , \9853 , \9857 );
and \U$9516 ( \9859 , \4568 , \1351 );
and \U$9517 ( \9860 , \4266 , \1349 );
nor \U$9518 ( \9861 , \9859 , \9860 );
xnor \U$9519 ( \9862 , \9861 , \1238 );
and \U$9520 ( \9863 , \9857 , \9862 );
and \U$9521 ( \9864 , \9853 , \9862 );
or \U$9522 ( \9865 , \9858 , \9863 , \9864 );
and \U$9523 ( \9866 , \9849 , \9865 );
and \U$9524 ( \9867 , \5045 , \1157 );
and \U$9525 ( \9868 , \4576 , \1155 );
nor \U$9526 ( \9869 , \9867 , \9868 );
xnor \U$9527 ( \9870 , \9869 , \1021 );
and \U$9528 ( \9871 , \5314 , \957 );
and \U$9529 ( \9872 , \5050 , \955 );
nor \U$9530 ( \9873 , \9871 , \9872 );
xnor \U$9531 ( \9874 , \9873 , \879 );
and \U$9532 ( \9875 , \9870 , \9874 );
and \U$9533 ( \9876 , \5945 , \793 );
and \U$9534 ( \9877 , \5573 , \791 );
nor \U$9535 ( \9878 , \9876 , \9877 );
xnor \U$9536 ( \9879 , \9878 , \699 );
and \U$9537 ( \9880 , \9874 , \9879 );
and \U$9538 ( \9881 , \9870 , \9879 );
or \U$9539 ( \9882 , \9875 , \9880 , \9881 );
and \U$9540 ( \9883 , \9865 , \9882 );
and \U$9541 ( \9884 , \9849 , \9882 );
or \U$9542 ( \9885 , \9866 , \9883 , \9884 );
and \U$9543 ( \9886 , \9833 , \9885 );
and \U$9544 ( \9887 , \1176 , \4977 );
and \U$9545 ( \9888 , \1071 , \4975 );
nor \U$9546 ( \9889 , \9887 , \9888 );
xnor \U$9547 ( \9890 , \9889 , \4789 );
and \U$9548 ( \9891 , \1297 , \4603 );
and \U$9549 ( \9892 , \1181 , \4601 );
nor \U$9550 ( \9893 , \9891 , \9892 );
xnor \U$9551 ( \9894 , \9893 , \4371 );
and \U$9552 ( \9895 , \9890 , \9894 );
and \U$9553 ( \9896 , \1588 , \4152 );
and \U$9554 ( \9897 , \1412 , \4150 );
nor \U$9555 ( \9898 , \9896 , \9897 );
xnor \U$9556 ( \9899 , \9898 , \4009 );
and \U$9557 ( \9900 , \9894 , \9899 );
and \U$9558 ( \9901 , \9890 , \9899 );
or \U$9559 ( \9902 , \9895 , \9900 , \9901 );
and \U$9560 ( \9903 , \2637 , \2715 );
and \U$9561 ( \9904 , \2463 , \2713 );
nor \U$9562 ( \9905 , \9903 , \9904 );
xnor \U$9563 ( \9906 , \9905 , \2566 );
and \U$9564 ( \9907 , \2942 , \2393 );
and \U$9565 ( \9908 , \2804 , \2391 );
nor \U$9566 ( \9909 , \9907 , \9908 );
xnor \U$9567 ( \9910 , \9909 , \2251 );
and \U$9568 ( \9911 , \9906 , \9910 );
and \U$9569 ( \9912 , \3478 , \2097 );
and \U$9570 ( \9913 , \3061 , \2095 );
nor \U$9571 ( \9914 , \9912 , \9913 );
xnor \U$9572 ( \9915 , \9914 , \1960 );
and \U$9573 ( \9916 , \9910 , \9915 );
and \U$9574 ( \9917 , \9906 , \9915 );
or \U$9575 ( \9918 , \9911 , \9916 , \9917 );
and \U$9576 ( \9919 , \9902 , \9918 );
and \U$9577 ( \9920 , \1839 , \3829 );
and \U$9578 ( \9921 , \1596 , \3827 );
nor \U$9579 ( \9922 , \9920 , \9921 );
xnor \U$9580 ( \9923 , \9922 , \3583 );
and \U$9581 ( \9924 , \2030 , \3434 );
and \U$9582 ( \9925 , \1844 , \3432 );
nor \U$9583 ( \9926 , \9924 , \9925 );
xnor \U$9584 ( \9927 , \9926 , \3247 );
and \U$9585 ( \9928 , \9923 , \9927 );
and \U$9586 ( \9929 , \2438 , \3121 );
and \U$9587 ( \9930 , \2174 , \3119 );
nor \U$9588 ( \9931 , \9929 , \9930 );
xnor \U$9589 ( \9932 , \9931 , \2916 );
and \U$9590 ( \9933 , \9927 , \9932 );
and \U$9591 ( \9934 , \9923 , \9932 );
or \U$9592 ( \9935 , \9928 , \9933 , \9934 );
and \U$9593 ( \9936 , \9918 , \9935 );
and \U$9594 ( \9937 , \9902 , \9935 );
or \U$9595 ( \9938 , \9919 , \9936 , \9937 );
and \U$9596 ( \9939 , \9885 , \9938 );
and \U$9597 ( \9940 , \9833 , \9938 );
or \U$9598 ( \9941 , \9886 , \9939 , \9940 );
and \U$9599 ( \9942 , \8170 , \391 );
and \U$9600 ( \9943 , \7924 , \389 );
nor \U$9601 ( \9944 , \9942 , \9943 );
xnor \U$9602 ( \9945 , \9944 , \398 );
and \U$9603 ( \9946 , \8494 , \406 );
and \U$9604 ( \9947 , \8175 , \404 );
nor \U$9605 ( \9948 , \9946 , \9947 );
xnor \U$9606 ( \9949 , \9948 , \413 );
and \U$9607 ( \9950 , \9945 , \9949 );
and \U$9608 ( \9951 , \9347 , \422 );
and \U$9609 ( \9952 , \8778 , \420 );
nor \U$9610 ( \9953 , \9951 , \9952 );
xnor \U$9611 ( \9954 , \9953 , \429 );
and \U$9612 ( \9955 , \9949 , \9954 );
and \U$9613 ( \9956 , \9945 , \9954 );
or \U$9614 ( \9957 , \9950 , \9955 , \9956 );
buf \U$9615 ( \9958 , RIbb2bbf0_125);
and \U$9616 ( \9959 , \9958 , \441 );
and \U$9617 ( \9960 , \9355 , \439 );
nor \U$9618 ( \9961 , \9959 , \9960 );
xnor \U$9619 ( \9962 , \9961 , \448 );
buf \U$9620 ( \9963 , RIbb2bb78_126);
and \U$9621 ( \9964 , \9963 , \436 );
or \U$9622 ( \9965 , \9962 , \9964 );
and \U$9623 ( \9966 , \9957 , \9965 );
and \U$9624 ( \9967 , \9355 , \441 );
and \U$9625 ( \9968 , \9347 , \439 );
nor \U$9626 ( \9969 , \9967 , \9968 );
xnor \U$9627 ( \9970 , \9969 , \448 );
and \U$9628 ( \9971 , \9965 , \9970 );
and \U$9629 ( \9972 , \9957 , \9970 );
or \U$9630 ( \9973 , \9966 , \9971 , \9972 );
and \U$9631 ( \9974 , \9958 , \436 );
xor \U$9632 ( \9975 , \9580 , \9584 );
xor \U$9633 ( \9976 , \9975 , \9589 );
and \U$9634 ( \9977 , \9974 , \9976 );
xor \U$9635 ( \9978 , \9656 , \9660 );
xor \U$9636 ( \9979 , \9978 , \9665 );
and \U$9637 ( \9980 , \9976 , \9979 );
and \U$9638 ( \9981 , \9974 , \9979 );
or \U$9639 ( \9982 , \9977 , \9980 , \9981 );
and \U$9640 ( \9983 , \9973 , \9982 );
xor \U$9641 ( \9984 , \9473 , \9477 );
xor \U$9642 ( \9985 , \9984 , \9482 );
xor \U$9643 ( \9986 , \9596 , \9600 );
xor \U$9644 ( \9987 , \9986 , \9605 );
and \U$9645 ( \9988 , \9985 , \9987 );
xor \U$9646 ( \9989 , \9613 , \9617 );
xor \U$9647 ( \9990 , \9989 , \9622 );
and \U$9648 ( \9991 , \9987 , \9990 );
and \U$9649 ( \9992 , \9985 , \9990 );
or \U$9650 ( \9993 , \9988 , \9991 , \9992 );
and \U$9651 ( \9994 , \9982 , \9993 );
and \U$9652 ( \9995 , \9973 , \9993 );
or \U$9653 ( \9996 , \9983 , \9994 , \9995 );
and \U$9654 ( \9997 , \9941 , \9996 );
xor \U$9655 ( \9998 , \9525 , \9529 );
xor \U$9656 ( \9999 , \9998 , \9534 );
xor \U$9657 ( \10000 , \9489 , \9493 );
xor \U$9658 ( \10001 , \10000 , \9498 );
and \U$9659 ( \10002 , \9999 , \10001 );
xor \U$9660 ( \10003 , \9506 , \9510 );
xor \U$9661 ( \10004 , \10003 , \9515 );
and \U$9662 ( \10005 , \10001 , \10004 );
and \U$9663 ( \10006 , \9999 , \10004 );
or \U$9664 ( \10007 , \10002 , \10005 , \10006 );
xor \U$9665 ( \10008 , \9541 , \9545 );
xor \U$9666 ( \10009 , \10008 , \9550 );
xor \U$9667 ( \10010 , \9560 , \9564 );
xor \U$9668 ( \10011 , \10010 , \9569 );
and \U$9669 ( \10012 , \10009 , \10011 );
and \U$9670 ( \10013 , \10007 , \10012 );
xor \U$9671 ( \10014 , \9681 , \9683 );
xor \U$9672 ( \10015 , \10014 , \9686 );
and \U$9673 ( \10016 , \10012 , \10015 );
and \U$9674 ( \10017 , \10007 , \10015 );
or \U$9675 ( \10018 , \10013 , \10016 , \10017 );
and \U$9676 ( \10019 , \9996 , \10018 );
and \U$9677 ( \10020 , \9941 , \10018 );
or \U$9678 ( \10021 , \9997 , \10019 , \10020 );
xor \U$9679 ( \10022 , \9485 , \9501 );
xor \U$9680 ( \10023 , \10022 , \9518 );
xor \U$9681 ( \10024 , \9537 , \9553 );
xor \U$9682 ( \10025 , \10024 , \9572 );
and \U$9683 ( \10026 , \10023 , \10025 );
xor \U$9684 ( \10027 , \9592 , \9608 );
xor \U$9685 ( \10028 , \10027 , \9625 );
and \U$9686 ( \10029 , \10025 , \10028 );
and \U$9687 ( \10030 , \10023 , \10028 );
or \U$9688 ( \10031 , \10026 , \10029 , \10030 );
xor \U$9689 ( \10032 , \9633 , \9635 );
xor \U$9690 ( \10033 , \10032 , \9638 );
xor \U$9691 ( \10034 , \9643 , \9645 );
xor \U$9692 ( \10035 , \10034 , \9648 );
and \U$9693 ( \10036 , \10033 , \10035 );
xor \U$9694 ( \10037 , \9668 , \9670 );
xor \U$9695 ( \10038 , \10037 , \9672 );
and \U$9696 ( \10039 , \10035 , \10038 );
and \U$9697 ( \10040 , \10033 , \10038 );
or \U$9698 ( \10041 , \10036 , \10039 , \10040 );
and \U$9699 ( \10042 , \10031 , \10041 );
xor \U$9700 ( \10043 , \9702 , \9704 );
xor \U$9701 ( \10044 , \10043 , \9707 );
and \U$9702 ( \10045 , \10041 , \10044 );
and \U$9703 ( \10046 , \10031 , \10044 );
or \U$9704 ( \10047 , \10042 , \10045 , \10046 );
and \U$9705 ( \10048 , \10021 , \10047 );
xor \U$9706 ( \10049 , \9641 , \9651 );
xor \U$9707 ( \10050 , \10049 , \9675 );
xor \U$9708 ( \10051 , \9712 , \9714 );
xor \U$9709 ( \10052 , \10051 , \9717 );
and \U$9710 ( \10053 , \10050 , \10052 );
xor \U$9711 ( \10054 , \9689 , \9691 );
xor \U$9712 ( \10055 , \10054 , \9694 );
and \U$9713 ( \10056 , \10052 , \10055 );
and \U$9714 ( \10057 , \10050 , \10055 );
or \U$9715 ( \10058 , \10053 , \10056 , \10057 );
and \U$9716 ( \10059 , \10047 , \10058 );
and \U$9717 ( \10060 , \10021 , \10058 );
or \U$9718 ( \10061 , \10048 , \10059 , \10060 );
xor \U$9719 ( \10062 , \9226 , \9281 );
xor \U$9720 ( \10063 , \10062 , \9334 );
xor \U$9721 ( \10064 , \9362 , \9372 );
xor \U$9722 ( \10065 , \10064 , \9383 );
and \U$9723 ( \10066 , \10063 , \10065 );
xor \U$9724 ( \10067 , \9729 , \9731 );
xor \U$9725 ( \10068 , \10067 , \9734 );
and \U$9726 ( \10069 , \10065 , \10068 );
and \U$9727 ( \10070 , \10063 , \10068 );
or \U$9728 ( \10071 , \10066 , \10069 , \10070 );
and \U$9729 ( \10072 , \10061 , \10071 );
xor \U$9730 ( \10073 , \9742 , \9744 );
xor \U$9731 ( \10074 , \10073 , \9747 );
and \U$9732 ( \10075 , \10071 , \10074 );
and \U$9733 ( \10076 , \10061 , \10074 );
or \U$9734 ( \10077 , \10072 , \10075 , \10076 );
xor \U$9735 ( \10078 , \9740 , \9750 );
xor \U$9736 ( \10079 , \10078 , \9753 );
and \U$9737 ( \10080 , \10077 , \10079 );
xor \U$9738 ( \10081 , \9758 , \9760 );
xor \U$9739 ( \10082 , \10081 , \9763 );
and \U$9740 ( \10083 , \10079 , \10082 );
and \U$9741 ( \10084 , \10077 , \10082 );
or \U$9742 ( \10085 , \10080 , \10083 , \10084 );
xor \U$9743 ( \10086 , \9756 , \9766 );
xor \U$9744 ( \10087 , \10086 , \9769 );
and \U$9745 ( \10088 , \10085 , \10087 );
xor \U$9746 ( \10089 , \9439 , \9449 );
xor \U$9747 ( \10090 , \10089 , \9452 );
and \U$9748 ( \10091 , \10087 , \10090 );
and \U$9749 ( \10092 , \10085 , \10090 );
or \U$9750 ( \10093 , \10088 , \10091 , \10092 );
and \U$9751 ( \10094 , \9778 , \10093 );
xor \U$9752 ( \10095 , \9778 , \10093 );
xor \U$9753 ( \10096 , \10085 , \10087 );
xor \U$9754 ( \10097 , \10096 , \10090 );
xor \U$9755 ( \10098 , \9906 , \9910 );
xor \U$9756 ( \10099 , \10098 , \9915 );
xor \U$9757 ( \10100 , \9923 , \9927 );
xor \U$9758 ( \10101 , \10100 , \9932 );
and \U$9759 ( \10102 , \10099 , \10101 );
xor \U$9760 ( \10103 , \9853 , \9857 );
xor \U$9761 ( \10104 , \10103 , \9862 );
and \U$9762 ( \10105 , \10101 , \10104 );
and \U$9763 ( \10106 , \10099 , \10104 );
or \U$9764 ( \10107 , \10102 , \10105 , \10106 );
xor \U$9765 ( \10108 , \9837 , \9841 );
xor \U$9766 ( \10109 , \10108 , \9846 );
xor \U$9767 ( \10110 , \9945 , \9949 );
xor \U$9768 ( \10111 , \10110 , \9954 );
and \U$9769 ( \10112 , \10109 , \10111 );
xor \U$9770 ( \10113 , \9870 , \9874 );
xor \U$9771 ( \10114 , \10113 , \9879 );
and \U$9772 ( \10115 , \10111 , \10114 );
and \U$9773 ( \10116 , \10109 , \10114 );
or \U$9774 ( \10117 , \10112 , \10115 , \10116 );
and \U$9775 ( \10118 , \10107 , \10117 );
and \U$9776 ( \10119 , \7924 , \373 );
and \U$9777 ( \10120 , \7500 , \371 );
nor \U$9778 ( \10121 , \10119 , \10120 );
xnor \U$9779 ( \10122 , \10121 , \380 );
and \U$9780 ( \10123 , \8175 , \391 );
and \U$9781 ( \10124 , \8170 , \389 );
nor \U$9782 ( \10125 , \10123 , \10124 );
xnor \U$9783 ( \10126 , \10125 , \398 );
and \U$9784 ( \10127 , \10122 , \10126 );
and \U$9785 ( \10128 , \8778 , \406 );
and \U$9786 ( \10129 , \8494 , \404 );
nor \U$9787 ( \10130 , \10128 , \10129 );
xnor \U$9788 ( \10131 , \10130 , \413 );
and \U$9789 ( \10132 , \10126 , \10131 );
and \U$9790 ( \10133 , \10122 , \10131 );
or \U$9791 ( \10134 , \10127 , \10132 , \10133 );
and \U$9792 ( \10135 , \9355 , \422 );
and \U$9793 ( \10136 , \9347 , \420 );
nor \U$9794 ( \10137 , \10135 , \10136 );
xnor \U$9795 ( \10138 , \10137 , \429 );
and \U$9796 ( \10139 , \9963 , \441 );
and \U$9797 ( \10140 , \9958 , \439 );
nor \U$9798 ( \10141 , \10139 , \10140 );
xnor \U$9799 ( \10142 , \10141 , \448 );
and \U$9800 ( \10143 , \10138 , \10142 );
buf \U$9801 ( \10144 , RIbb31500_127);
and \U$9802 ( \10145 , \10144 , \436 );
and \U$9803 ( \10146 , \10142 , \10145 );
and \U$9804 ( \10147 , \10138 , \10145 );
or \U$9805 ( \10148 , \10143 , \10146 , \10147 );
and \U$9806 ( \10149 , \10134 , \10148 );
xnor \U$9807 ( \10150 , \9962 , \9964 );
and \U$9808 ( \10151 , \10148 , \10150 );
and \U$9809 ( \10152 , \10134 , \10150 );
or \U$9810 ( \10153 , \10149 , \10151 , \10152 );
and \U$9811 ( \10154 , \10117 , \10153 );
and \U$9812 ( \10155 , \10107 , \10153 );
or \U$9813 ( \10156 , \10118 , \10154 , \10155 );
not \U$9814 ( \10157 , \9556 );
and \U$9815 ( \10158 , \351 , \9798 );
and \U$9816 ( \10159 , \359 , \9796 );
nor \U$9817 ( \10160 , \10158 , \10159 );
xnor \U$9818 ( \10161 , \10160 , \9559 );
and \U$9819 ( \10162 , \10157 , \10161 );
and \U$9820 ( \10163 , \367 , \9230 );
and \U$9821 ( \10164 , \375 , \9228 );
nor \U$9822 ( \10165 , \10163 , \10164 );
xnor \U$9823 ( \10166 , \10165 , \8920 );
and \U$9824 ( \10167 , \10161 , \10166 );
and \U$9825 ( \10168 , \10157 , \10166 );
or \U$9826 ( \10169 , \10162 , \10167 , \10168 );
and \U$9827 ( \10170 , \385 , \8693 );
and \U$9828 ( \10171 , \393 , \8691 );
nor \U$9829 ( \10172 , \10170 , \10171 );
xnor \U$9830 ( \10173 , \10172 , \8322 );
and \U$9831 ( \10174 , \400 , \8131 );
and \U$9832 ( \10175 , \408 , \8129 );
nor \U$9833 ( \10176 , \10174 , \10175 );
xnor \U$9834 ( \10177 , \10176 , \7813 );
and \U$9835 ( \10178 , \10173 , \10177 );
and \U$9836 ( \10179 , \416 , \7564 );
and \U$9837 ( \10180 , \424 , \7562 );
nor \U$9838 ( \10181 , \10179 , \10180 );
xnor \U$9839 ( \10182 , \10181 , \7315 );
and \U$9840 ( \10183 , \10177 , \10182 );
and \U$9841 ( \10184 , \10173 , \10182 );
or \U$9842 ( \10185 , \10178 , \10183 , \10184 );
and \U$9843 ( \10186 , \10169 , \10185 );
and \U$9844 ( \10187 , \435 , \7035 );
and \U$9845 ( \10188 , \443 , \7033 );
nor \U$9846 ( \10189 , \10187 , \10188 );
xnor \U$9847 ( \10190 , \10189 , \6775 );
and \U$9848 ( \10191 , \661 , \6541 );
and \U$9849 ( \10192 , \450 , \6539 );
nor \U$9850 ( \10193 , \10191 , \10192 );
xnor \U$9851 ( \10194 , \10193 , \6226 );
and \U$9852 ( \10195 , \10190 , \10194 );
and \U$9853 ( \10196 , \785 , \6032 );
and \U$9854 ( \10197 , \722 , \6030 );
nor \U$9855 ( \10198 , \10196 , \10197 );
xnor \U$9856 ( \10199 , \10198 , \5692 );
and \U$9857 ( \10200 , \10194 , \10199 );
and \U$9858 ( \10201 , \10190 , \10199 );
or \U$9859 ( \10202 , \10195 , \10200 , \10201 );
and \U$9860 ( \10203 , \10185 , \10202 );
and \U$9861 ( \10204 , \10169 , \10202 );
or \U$9862 ( \10205 , \10186 , \10203 , \10204 );
and \U$9863 ( \10206 , \4576 , \1351 );
and \U$9864 ( \10207 , \4568 , \1349 );
nor \U$9865 ( \10208 , \10206 , \10207 );
xnor \U$9866 ( \10209 , \10208 , \1238 );
and \U$9867 ( \10210 , \5050 , \1157 );
and \U$9868 ( \10211 , \5045 , \1155 );
nor \U$9869 ( \10212 , \10210 , \10211 );
xnor \U$9870 ( \10213 , \10212 , \1021 );
and \U$9871 ( \10214 , \10209 , \10213 );
and \U$9872 ( \10215 , \5573 , \957 );
and \U$9873 ( \10216 , \5314 , \955 );
nor \U$9874 ( \10217 , \10215 , \10216 );
xnor \U$9875 ( \10218 , \10217 , \879 );
and \U$9876 ( \10219 , \10213 , \10218 );
and \U$9877 ( \10220 , \10209 , \10218 );
or \U$9878 ( \10221 , \10214 , \10219 , \10220 );
and \U$9879 ( \10222 , \3686 , \2097 );
and \U$9880 ( \10223 , \3478 , \2095 );
nor \U$9881 ( \10224 , \10222 , \10223 );
xnor \U$9882 ( \10225 , \10224 , \1960 );
and \U$9883 ( \10226 , \3813 , \1891 );
and \U$9884 ( \10227 , \3808 , \1889 );
nor \U$9885 ( \10228 , \10226 , \10227 );
xnor \U$9886 ( \10229 , \10228 , \1739 );
and \U$9887 ( \10230 , \10225 , \10229 );
and \U$9888 ( \10231 , \4266 , \1623 );
and \U$9889 ( \10232 , \4069 , \1621 );
nor \U$9890 ( \10233 , \10231 , \10232 );
xnor \U$9891 ( \10234 , \10233 , \1467 );
and \U$9892 ( \10235 , \10229 , \10234 );
and \U$9893 ( \10236 , \10225 , \10234 );
or \U$9894 ( \10237 , \10230 , \10235 , \10236 );
and \U$9895 ( \10238 , \10221 , \10237 );
and \U$9896 ( \10239 , \5954 , \793 );
and \U$9897 ( \10240 , \5945 , \791 );
nor \U$9898 ( \10241 , \10239 , \10240 );
xnor \U$9899 ( \10242 , \10241 , \699 );
and \U$9900 ( \10243 , \6499 , \624 );
and \U$9901 ( \10244 , \6297 , \622 );
nor \U$9902 ( \10245 , \10243 , \10244 );
xnor \U$9903 ( \10246 , \10245 , \349 );
and \U$9904 ( \10247 , \10242 , \10246 );
and \U$9905 ( \10248 , \6974 , \357 );
and \U$9906 ( \10249 , \6802 , \355 );
nor \U$9907 ( \10250 , \10248 , \10249 );
xnor \U$9908 ( \10251 , \10250 , \364 );
and \U$9909 ( \10252 , \10246 , \10251 );
and \U$9910 ( \10253 , \10242 , \10251 );
or \U$9911 ( \10254 , \10247 , \10252 , \10253 );
and \U$9912 ( \10255 , \10237 , \10254 );
and \U$9913 ( \10256 , \10221 , \10254 );
or \U$9914 ( \10257 , \10238 , \10255 , \10256 );
and \U$9915 ( \10258 , \10205 , \10257 );
and \U$9916 ( \10259 , \1596 , \4152 );
and \U$9917 ( \10260 , \1588 , \4150 );
nor \U$9918 ( \10261 , \10259 , \10260 );
xnor \U$9919 ( \10262 , \10261 , \4009 );
and \U$9920 ( \10263 , \1844 , \3829 );
and \U$9921 ( \10264 , \1839 , \3827 );
nor \U$9922 ( \10265 , \10263 , \10264 );
xnor \U$9923 ( \10266 , \10265 , \3583 );
and \U$9924 ( \10267 , \10262 , \10266 );
and \U$9925 ( \10268 , \2174 , \3434 );
and \U$9926 ( \10269 , \2030 , \3432 );
nor \U$9927 ( \10270 , \10268 , \10269 );
xnor \U$9928 ( \10271 , \10270 , \3247 );
and \U$9929 ( \10272 , \10266 , \10271 );
and \U$9930 ( \10273 , \10262 , \10271 );
or \U$9931 ( \10274 , \10267 , \10272 , \10273 );
and \U$9932 ( \10275 , \2463 , \3121 );
and \U$9933 ( \10276 , \2438 , \3119 );
nor \U$9934 ( \10277 , \10275 , \10276 );
xnor \U$9935 ( \10278 , \10277 , \2916 );
and \U$9936 ( \10279 , \2804 , \2715 );
and \U$9937 ( \10280 , \2637 , \2713 );
nor \U$9938 ( \10281 , \10279 , \10280 );
xnor \U$9939 ( \10282 , \10281 , \2566 );
and \U$9940 ( \10283 , \10278 , \10282 );
and \U$9941 ( \10284 , \3061 , \2393 );
and \U$9942 ( \10285 , \2942 , \2391 );
nor \U$9943 ( \10286 , \10284 , \10285 );
xnor \U$9944 ( \10287 , \10286 , \2251 );
and \U$9945 ( \10288 , \10282 , \10287 );
and \U$9946 ( \10289 , \10278 , \10287 );
or \U$9947 ( \10290 , \10283 , \10288 , \10289 );
and \U$9948 ( \10291 , \10274 , \10290 );
and \U$9949 ( \10292 , \1071 , \5443 );
and \U$9950 ( \10293 , \983 , \5441 );
nor \U$9951 ( \10294 , \10292 , \10293 );
xnor \U$9952 ( \10295 , \10294 , \5202 );
and \U$9953 ( \10296 , \1181 , \4977 );
and \U$9954 ( \10297 , \1176 , \4975 );
nor \U$9955 ( \10298 , \10296 , \10297 );
xnor \U$9956 ( \10299 , \10298 , \4789 );
and \U$9957 ( \10300 , \10295 , \10299 );
and \U$9958 ( \10301 , \1412 , \4603 );
and \U$9959 ( \10302 , \1297 , \4601 );
nor \U$9960 ( \10303 , \10301 , \10302 );
xnor \U$9961 ( \10304 , \10303 , \4371 );
and \U$9962 ( \10305 , \10299 , \10304 );
and \U$9963 ( \10306 , \10295 , \10304 );
or \U$9964 ( \10307 , \10300 , \10305 , \10306 );
and \U$9965 ( \10308 , \10290 , \10307 );
and \U$9966 ( \10309 , \10274 , \10307 );
or \U$9967 ( \10310 , \10291 , \10308 , \10309 );
and \U$9968 ( \10311 , \10257 , \10310 );
and \U$9969 ( \10312 , \10205 , \10310 );
or \U$9970 ( \10313 , \10258 , \10311 , \10312 );
and \U$9971 ( \10314 , \10156 , \10313 );
xor \U$9972 ( \10315 , \9890 , \9894 );
xor \U$9973 ( \10316 , \10315 , \9899 );
xor \U$9974 ( \10317 , \9782 , \9786 );
xor \U$9975 ( \10318 , \10317 , \9791 );
and \U$9976 ( \10319 , \10316 , \10318 );
xor \U$9977 ( \10320 , \9818 , \9822 );
xor \U$9978 ( \10321 , \10320 , \9827 );
and \U$9979 ( \10322 , \10318 , \10321 );
and \U$9980 ( \10323 , \10316 , \10321 );
or \U$9981 ( \10324 , \10319 , \10322 , \10323 );
xor \U$9982 ( \10325 , \9999 , \10001 );
xor \U$9983 ( \10326 , \10325 , \10004 );
and \U$9984 ( \10327 , \10324 , \10326 );
xor \U$9985 ( \10328 , \10009 , \10011 );
and \U$9986 ( \10329 , \10326 , \10328 );
and \U$9987 ( \10330 , \10324 , \10328 );
or \U$9988 ( \10331 , \10327 , \10329 , \10330 );
and \U$9989 ( \10332 , \10313 , \10331 );
and \U$9990 ( \10333 , \10156 , \10331 );
or \U$9991 ( \10334 , \10314 , \10332 , \10333 );
xor \U$9992 ( \10335 , \9794 , \9813 );
xor \U$9993 ( \10336 , \10335 , \9830 );
xor \U$9994 ( \10337 , \9849 , \9865 );
xor \U$9995 ( \10338 , \10337 , \9882 );
and \U$9996 ( \10339 , \10336 , \10338 );
xor \U$9997 ( \10340 , \9902 , \9918 );
xor \U$9998 ( \10341 , \10340 , \9935 );
and \U$9999 ( \10342 , \10338 , \10341 );
and \U$10000 ( \10343 , \10336 , \10341 );
or \U$10001 ( \10344 , \10339 , \10342 , \10343 );
xor \U$10002 ( \10345 , \9957 , \9965 );
xor \U$10003 ( \10346 , \10345 , \9970 );
xor \U$10004 ( \10347 , \9974 , \9976 );
xor \U$10005 ( \10348 , \10347 , \9979 );
and \U$10006 ( \10349 , \10346 , \10348 );
xor \U$10007 ( \10350 , \9985 , \9987 );
xor \U$10008 ( \10351 , \10350 , \9990 );
and \U$10009 ( \10352 , \10348 , \10351 );
and \U$10010 ( \10353 , \10346 , \10351 );
or \U$10011 ( \10354 , \10349 , \10352 , \10353 );
and \U$10012 ( \10355 , \10344 , \10354 );
xor \U$10013 ( \10356 , \10023 , \10025 );
xor \U$10014 ( \10357 , \10356 , \10028 );
and \U$10015 ( \10358 , \10354 , \10357 );
and \U$10016 ( \10359 , \10344 , \10357 );
or \U$10017 ( \10360 , \10355 , \10358 , \10359 );
and \U$10018 ( \10361 , \10334 , \10360 );
xor \U$10019 ( \10362 , \9973 , \9982 );
xor \U$10020 ( \10363 , \10362 , \9993 );
xor \U$10021 ( \10364 , \10007 , \10012 );
xor \U$10022 ( \10365 , \10364 , \10015 );
and \U$10023 ( \10366 , \10363 , \10365 );
xor \U$10024 ( \10367 , \10033 , \10035 );
xor \U$10025 ( \10368 , \10367 , \10038 );
and \U$10026 ( \10369 , \10365 , \10368 );
and \U$10027 ( \10370 , \10363 , \10368 );
or \U$10028 ( \10371 , \10366 , \10369 , \10370 );
and \U$10029 ( \10372 , \10360 , \10371 );
and \U$10030 ( \10373 , \10334 , \10371 );
or \U$10031 ( \10374 , \10361 , \10372 , \10373 );
xor \U$10032 ( \10375 , \9521 , \9575 );
xor \U$10033 ( \10376 , \10375 , \9628 );
xor \U$10034 ( \10377 , \10031 , \10041 );
xor \U$10035 ( \10378 , \10377 , \10044 );
and \U$10036 ( \10379 , \10376 , \10378 );
xor \U$10037 ( \10380 , \10050 , \10052 );
xor \U$10038 ( \10381 , \10380 , \10055 );
and \U$10039 ( \10382 , \10378 , \10381 );
and \U$10040 ( \10383 , \10376 , \10381 );
or \U$10041 ( \10384 , \10379 , \10382 , \10383 );
and \U$10042 ( \10385 , \10374 , \10384 );
xor \U$10043 ( \10386 , \9710 , \9720 );
xor \U$10044 ( \10387 , \10386 , \9723 );
and \U$10045 ( \10388 , \10384 , \10387 );
and \U$10046 ( \10389 , \10374 , \10387 );
or \U$10047 ( \10390 , \10385 , \10388 , \10389 );
xor \U$10048 ( \10391 , \9631 , \9678 );
xor \U$10049 ( \10392 , \10391 , \9697 );
xor \U$10050 ( \10393 , \10021 , \10047 );
xor \U$10051 ( \10394 , \10393 , \10058 );
and \U$10052 ( \10395 , \10392 , \10394 );
xor \U$10053 ( \10396 , \10063 , \10065 );
xor \U$10054 ( \10397 , \10396 , \10068 );
and \U$10055 ( \10398 , \10394 , \10397 );
and \U$10056 ( \10399 , \10392 , \10397 );
or \U$10057 ( \10400 , \10395 , \10398 , \10399 );
and \U$10058 ( \10401 , \10390 , \10400 );
xor \U$10059 ( \10402 , \9700 , \9726 );
xor \U$10060 ( \10403 , \10402 , \9737 );
and \U$10061 ( \10404 , \10400 , \10403 );
and \U$10062 ( \10405 , \10390 , \10403 );
or \U$10063 ( \10406 , \10401 , \10404 , \10405 );
xor \U$10064 ( \10407 , \10077 , \10079 );
xor \U$10065 ( \10408 , \10407 , \10082 );
and \U$10066 ( \10409 , \10406 , \10408 );
and \U$10067 ( \10410 , \10097 , \10409 );
xor \U$10068 ( \10411 , \10097 , \10409 );
xor \U$10069 ( \10412 , \10406 , \10408 );
xor \U$10070 ( \10413 , \10209 , \10213 );
xor \U$10071 ( \10414 , \10413 , \10218 );
xor \U$10072 ( \10415 , \10225 , \10229 );
xor \U$10073 ( \10416 , \10415 , \10234 );
and \U$10074 ( \10417 , \10414 , \10416 );
xor \U$10075 ( \10418 , \10278 , \10282 );
xor \U$10076 ( \10419 , \10418 , \10287 );
and \U$10077 ( \10420 , \10416 , \10419 );
and \U$10078 ( \10421 , \10414 , \10419 );
or \U$10079 ( \10422 , \10417 , \10420 , \10421 );
xor \U$10080 ( \10423 , \10122 , \10126 );
xor \U$10081 ( \10424 , \10423 , \10131 );
xor \U$10082 ( \10425 , \10138 , \10142 );
xor \U$10083 ( \10426 , \10425 , \10145 );
and \U$10084 ( \10427 , \10424 , \10426 );
xor \U$10085 ( \10428 , \10242 , \10246 );
xor \U$10086 ( \10429 , \10428 , \10251 );
and \U$10087 ( \10430 , \10426 , \10429 );
and \U$10088 ( \10431 , \10424 , \10429 );
or \U$10089 ( \10432 , \10427 , \10430 , \10431 );
and \U$10090 ( \10433 , \10422 , \10432 );
and \U$10091 ( \10434 , \7500 , \357 );
and \U$10092 ( \10435 , \6974 , \355 );
nor \U$10093 ( \10436 , \10434 , \10435 );
xnor \U$10094 ( \10437 , \10436 , \364 );
and \U$10095 ( \10438 , \8170 , \373 );
and \U$10096 ( \10439 , \7924 , \371 );
nor \U$10097 ( \10440 , \10438 , \10439 );
xnor \U$10098 ( \10441 , \10440 , \380 );
and \U$10099 ( \10442 , \10437 , \10441 );
and \U$10100 ( \10443 , \8494 , \391 );
and \U$10101 ( \10444 , \8175 , \389 );
nor \U$10102 ( \10445 , \10443 , \10444 );
xnor \U$10103 ( \10446 , \10445 , \398 );
and \U$10104 ( \10447 , \10441 , \10446 );
and \U$10105 ( \10448 , \10437 , \10446 );
or \U$10106 ( \10449 , \10442 , \10447 , \10448 );
and \U$10107 ( \10450 , \9347 , \406 );
and \U$10108 ( \10451 , \8778 , \404 );
nor \U$10109 ( \10452 , \10450 , \10451 );
xnor \U$10110 ( \10453 , \10452 , \413 );
and \U$10111 ( \10454 , \9958 , \422 );
and \U$10112 ( \10455 , \9355 , \420 );
nor \U$10113 ( \10456 , \10454 , \10455 );
xnor \U$10114 ( \10457 , \10456 , \429 );
and \U$10115 ( \10458 , \10453 , \10457 );
and \U$10116 ( \10459 , \10144 , \441 );
and \U$10117 ( \10460 , \9963 , \439 );
nor \U$10118 ( \10461 , \10459 , \10460 );
xnor \U$10119 ( \10462 , \10461 , \448 );
and \U$10120 ( \10463 , \10457 , \10462 );
and \U$10121 ( \10464 , \10453 , \10462 );
or \U$10122 ( \10465 , \10458 , \10463 , \10464 );
or \U$10123 ( \10466 , \10449 , \10465 );
and \U$10124 ( \10467 , \10432 , \10466 );
and \U$10125 ( \10468 , \10422 , \10466 );
or \U$10126 ( \10469 , \10433 , \10467 , \10468 );
and \U$10127 ( \10470 , \4568 , \1623 );
and \U$10128 ( \10471 , \4266 , \1621 );
nor \U$10129 ( \10472 , \10470 , \10471 );
xnor \U$10130 ( \10473 , \10472 , \1467 );
and \U$10131 ( \10474 , \5045 , \1351 );
and \U$10132 ( \10475 , \4576 , \1349 );
nor \U$10133 ( \10476 , \10474 , \10475 );
xnor \U$10134 ( \10477 , \10476 , \1238 );
and \U$10135 ( \10478 , \10473 , \10477 );
and \U$10136 ( \10479 , \5314 , \1157 );
and \U$10137 ( \10480 , \5050 , \1155 );
nor \U$10138 ( \10481 , \10479 , \10480 );
xnor \U$10139 ( \10482 , \10481 , \1021 );
and \U$10140 ( \10483 , \10477 , \10482 );
and \U$10141 ( \10484 , \10473 , \10482 );
or \U$10142 ( \10485 , \10478 , \10483 , \10484 );
and \U$10143 ( \10486 , \5945 , \957 );
and \U$10144 ( \10487 , \5573 , \955 );
nor \U$10145 ( \10488 , \10486 , \10487 );
xnor \U$10146 ( \10489 , \10488 , \879 );
and \U$10147 ( \10490 , \6297 , \793 );
and \U$10148 ( \10491 , \5954 , \791 );
nor \U$10149 ( \10492 , \10490 , \10491 );
xnor \U$10150 ( \10493 , \10492 , \699 );
and \U$10151 ( \10494 , \10489 , \10493 );
and \U$10152 ( \10495 , \6802 , \624 );
and \U$10153 ( \10496 , \6499 , \622 );
nor \U$10154 ( \10497 , \10495 , \10496 );
xnor \U$10155 ( \10498 , \10497 , \349 );
and \U$10156 ( \10499 , \10493 , \10498 );
and \U$10157 ( \10500 , \10489 , \10498 );
or \U$10158 ( \10501 , \10494 , \10499 , \10500 );
and \U$10159 ( \10502 , \10485 , \10501 );
and \U$10160 ( \10503 , \3478 , \2393 );
and \U$10161 ( \10504 , \3061 , \2391 );
nor \U$10162 ( \10505 , \10503 , \10504 );
xnor \U$10163 ( \10506 , \10505 , \2251 );
and \U$10164 ( \10507 , \3808 , \2097 );
and \U$10165 ( \10508 , \3686 , \2095 );
nor \U$10166 ( \10509 , \10507 , \10508 );
xnor \U$10167 ( \10510 , \10509 , \1960 );
and \U$10168 ( \10511 , \10506 , \10510 );
and \U$10169 ( \10512 , \4069 , \1891 );
and \U$10170 ( \10513 , \3813 , \1889 );
nor \U$10171 ( \10514 , \10512 , \10513 );
xnor \U$10172 ( \10515 , \10514 , \1739 );
and \U$10173 ( \10516 , \10510 , \10515 );
and \U$10174 ( \10517 , \10506 , \10515 );
or \U$10175 ( \10518 , \10511 , \10516 , \10517 );
and \U$10176 ( \10519 , \10501 , \10518 );
and \U$10177 ( \10520 , \10485 , \10518 );
or \U$10178 ( \10521 , \10502 , \10519 , \10520 );
and \U$10179 ( \10522 , \1588 , \4603 );
and \U$10180 ( \10523 , \1412 , \4601 );
nor \U$10181 ( \10524 , \10522 , \10523 );
xnor \U$10182 ( \10525 , \10524 , \4371 );
and \U$10183 ( \10526 , \1839 , \4152 );
and \U$10184 ( \10527 , \1596 , \4150 );
nor \U$10185 ( \10528 , \10526 , \10527 );
xnor \U$10186 ( \10529 , \10528 , \4009 );
and \U$10187 ( \10530 , \10525 , \10529 );
and \U$10188 ( \10531 , \2030 , \3829 );
and \U$10189 ( \10532 , \1844 , \3827 );
nor \U$10190 ( \10533 , \10531 , \10532 );
xnor \U$10191 ( \10534 , \10533 , \3583 );
and \U$10192 ( \10535 , \10529 , \10534 );
and \U$10193 ( \10536 , \10525 , \10534 );
or \U$10194 ( \10537 , \10530 , \10535 , \10536 );
and \U$10195 ( \10538 , \2438 , \3434 );
and \U$10196 ( \10539 , \2174 , \3432 );
nor \U$10197 ( \10540 , \10538 , \10539 );
xnor \U$10198 ( \10541 , \10540 , \3247 );
and \U$10199 ( \10542 , \2637 , \3121 );
and \U$10200 ( \10543 , \2463 , \3119 );
nor \U$10201 ( \10544 , \10542 , \10543 );
xnor \U$10202 ( \10545 , \10544 , \2916 );
and \U$10203 ( \10546 , \10541 , \10545 );
and \U$10204 ( \10547 , \2942 , \2715 );
and \U$10205 ( \10548 , \2804 , \2713 );
nor \U$10206 ( \10549 , \10547 , \10548 );
xnor \U$10207 ( \10550 , \10549 , \2566 );
and \U$10208 ( \10551 , \10545 , \10550 );
and \U$10209 ( \10552 , \10541 , \10550 );
or \U$10210 ( \10553 , \10546 , \10551 , \10552 );
and \U$10211 ( \10554 , \10537 , \10553 );
and \U$10212 ( \10555 , \983 , \6032 );
and \U$10213 ( \10556 , \785 , \6030 );
nor \U$10214 ( \10557 , \10555 , \10556 );
xnor \U$10215 ( \10558 , \10557 , \5692 );
and \U$10216 ( \10559 , \1176 , \5443 );
and \U$10217 ( \10560 , \1071 , \5441 );
nor \U$10218 ( \10561 , \10559 , \10560 );
xnor \U$10219 ( \10562 , \10561 , \5202 );
and \U$10220 ( \10563 , \10558 , \10562 );
and \U$10221 ( \10564 , \1297 , \4977 );
and \U$10222 ( \10565 , \1181 , \4975 );
nor \U$10223 ( \10566 , \10564 , \10565 );
xnor \U$10224 ( \10567 , \10566 , \4789 );
and \U$10225 ( \10568 , \10562 , \10567 );
and \U$10226 ( \10569 , \10558 , \10567 );
or \U$10227 ( \10570 , \10563 , \10568 , \10569 );
and \U$10228 ( \10571 , \10553 , \10570 );
and \U$10229 ( \10572 , \10537 , \10570 );
or \U$10230 ( \10573 , \10554 , \10571 , \10572 );
and \U$10231 ( \10574 , \10521 , \10573 );
and \U$10232 ( \10575 , \393 , \9230 );
and \U$10233 ( \10576 , \367 , \9228 );
nor \U$10234 ( \10577 , \10575 , \10576 );
xnor \U$10235 ( \10578 , \10577 , \8920 );
and \U$10236 ( \10579 , \408 , \8693 );
and \U$10237 ( \10580 , \385 , \8691 );
nor \U$10238 ( \10581 , \10579 , \10580 );
xnor \U$10239 ( \10582 , \10581 , \8322 );
and \U$10240 ( \10583 , \10578 , \10582 );
and \U$10241 ( \10584 , \424 , \8131 );
and \U$10242 ( \10585 , \400 , \8129 );
nor \U$10243 ( \10586 , \10584 , \10585 );
xnor \U$10244 ( \10587 , \10586 , \7813 );
and \U$10245 ( \10588 , \10582 , \10587 );
and \U$10246 ( \10589 , \10578 , \10587 );
or \U$10247 ( \10590 , \10583 , \10588 , \10589 );
and \U$10248 ( \10591 , \443 , \7564 );
and \U$10249 ( \10592 , \416 , \7562 );
nor \U$10250 ( \10593 , \10591 , \10592 );
xnor \U$10251 ( \10594 , \10593 , \7315 );
and \U$10252 ( \10595 , \450 , \7035 );
and \U$10253 ( \10596 , \435 , \7033 );
nor \U$10254 ( \10597 , \10595 , \10596 );
xnor \U$10255 ( \10598 , \10597 , \6775 );
and \U$10256 ( \10599 , \10594 , \10598 );
and \U$10257 ( \10600 , \722 , \6541 );
and \U$10258 ( \10601 , \661 , \6539 );
nor \U$10259 ( \10602 , \10600 , \10601 );
xnor \U$10260 ( \10603 , \10602 , \6226 );
and \U$10261 ( \10604 , \10598 , \10603 );
and \U$10262 ( \10605 , \10594 , \10603 );
or \U$10263 ( \10606 , \10599 , \10604 , \10605 );
and \U$10264 ( \10607 , \10590 , \10606 );
buf \U$10265 ( \10608 , RIbb2d888_64);
xor \U$10266 ( \10609 , \9556 , \10608 );
not \U$10267 ( \10610 , \10608 );
and \U$10268 ( \10611 , \10609 , \10610 );
and \U$10269 ( \10612 , \359 , \10611 );
not \U$10270 ( \10613 , \10612 );
xnor \U$10271 ( \10614 , \10613 , \9556 );
and \U$10272 ( \10615 , \375 , \9798 );
and \U$10273 ( \10616 , \351 , \9796 );
nor \U$10274 ( \10617 , \10615 , \10616 );
xnor \U$10275 ( \10618 , \10617 , \9559 );
and \U$10276 ( \10619 , \10614 , \10618 );
and \U$10277 ( \10620 , \10606 , \10619 );
and \U$10278 ( \10621 , \10590 , \10619 );
or \U$10279 ( \10622 , \10607 , \10620 , \10621 );
and \U$10280 ( \10623 , \10573 , \10622 );
and \U$10281 ( \10624 , \10521 , \10622 );
or \U$10282 ( \10625 , \10574 , \10623 , \10624 );
and \U$10283 ( \10626 , \10469 , \10625 );
xor \U$10284 ( \10627 , \10262 , \10266 );
xor \U$10285 ( \10628 , \10627 , \10271 );
xor \U$10286 ( \10629 , \10190 , \10194 );
xor \U$10287 ( \10630 , \10629 , \10199 );
and \U$10288 ( \10631 , \10628 , \10630 );
xor \U$10289 ( \10632 , \10295 , \10299 );
xor \U$10290 ( \10633 , \10632 , \10304 );
and \U$10291 ( \10634 , \10630 , \10633 );
and \U$10292 ( \10635 , \10628 , \10633 );
or \U$10293 ( \10636 , \10631 , \10634 , \10635 );
xor \U$10294 ( \10637 , \10157 , \10161 );
xor \U$10295 ( \10638 , \10637 , \10166 );
xor \U$10296 ( \10639 , \10173 , \10177 );
xor \U$10297 ( \10640 , \10639 , \10182 );
and \U$10298 ( \10641 , \10638 , \10640 );
and \U$10299 ( \10642 , \10636 , \10641 );
xor \U$10300 ( \10643 , \9801 , \9805 );
xor \U$10301 ( \10644 , \10643 , \9810 );
and \U$10302 ( \10645 , \10641 , \10644 );
and \U$10303 ( \10646 , \10636 , \10644 );
or \U$10304 ( \10647 , \10642 , \10645 , \10646 );
and \U$10305 ( \10648 , \10625 , \10647 );
and \U$10306 ( \10649 , \10469 , \10647 );
or \U$10307 ( \10650 , \10626 , \10648 , \10649 );
xor \U$10308 ( \10651 , \10316 , \10318 );
xor \U$10309 ( \10652 , \10651 , \10321 );
xor \U$10310 ( \10653 , \10099 , \10101 );
xor \U$10311 ( \10654 , \10653 , \10104 );
and \U$10312 ( \10655 , \10652 , \10654 );
xor \U$10313 ( \10656 , \10109 , \10111 );
xor \U$10314 ( \10657 , \10656 , \10114 );
and \U$10315 ( \10658 , \10654 , \10657 );
and \U$10316 ( \10659 , \10652 , \10657 );
or \U$10317 ( \10660 , \10655 , \10658 , \10659 );
xor \U$10318 ( \10661 , \10221 , \10237 );
xor \U$10319 ( \10662 , \10661 , \10254 );
xor \U$10320 ( \10663 , \10274 , \10290 );
xor \U$10321 ( \10664 , \10663 , \10307 );
and \U$10322 ( \10665 , \10662 , \10664 );
xor \U$10323 ( \10666 , \10134 , \10148 );
xor \U$10324 ( \10667 , \10666 , \10150 );
and \U$10325 ( \10668 , \10664 , \10667 );
and \U$10326 ( \10669 , \10662 , \10667 );
or \U$10327 ( \10670 , \10665 , \10668 , \10669 );
and \U$10328 ( \10671 , \10660 , \10670 );
xor \U$10329 ( \10672 , \10336 , \10338 );
xor \U$10330 ( \10673 , \10672 , \10341 );
and \U$10331 ( \10674 , \10670 , \10673 );
and \U$10332 ( \10675 , \10660 , \10673 );
or \U$10333 ( \10676 , \10671 , \10674 , \10675 );
and \U$10334 ( \10677 , \10650 , \10676 );
xor \U$10335 ( \10678 , \10107 , \10117 );
xor \U$10336 ( \10679 , \10678 , \10153 );
xor \U$10337 ( \10680 , \10346 , \10348 );
xor \U$10338 ( \10681 , \10680 , \10351 );
and \U$10339 ( \10682 , \10679 , \10681 );
xor \U$10340 ( \10683 , \10324 , \10326 );
xor \U$10341 ( \10684 , \10683 , \10328 );
and \U$10342 ( \10685 , \10681 , \10684 );
and \U$10343 ( \10686 , \10679 , \10684 );
or \U$10344 ( \10687 , \10682 , \10685 , \10686 );
and \U$10345 ( \10688 , \10676 , \10687 );
and \U$10346 ( \10689 , \10650 , \10687 );
or \U$10347 ( \10690 , \10677 , \10688 , \10689 );
xor \U$10348 ( \10691 , \9833 , \9885 );
xor \U$10349 ( \10692 , \10691 , \9938 );
xor \U$10350 ( \10693 , \10344 , \10354 );
xor \U$10351 ( \10694 , \10693 , \10357 );
and \U$10352 ( \10695 , \10692 , \10694 );
xor \U$10353 ( \10696 , \10363 , \10365 );
xor \U$10354 ( \10697 , \10696 , \10368 );
and \U$10355 ( \10698 , \10694 , \10697 );
and \U$10356 ( \10699 , \10692 , \10697 );
or \U$10357 ( \10700 , \10695 , \10698 , \10699 );
and \U$10358 ( \10701 , \10690 , \10700 );
xor \U$10359 ( \10702 , \9941 , \9996 );
xor \U$10360 ( \10703 , \10702 , \10018 );
and \U$10361 ( \10704 , \10700 , \10703 );
and \U$10362 ( \10705 , \10690 , \10703 );
or \U$10363 ( \10706 , \10701 , \10704 , \10705 );
xor \U$10364 ( \10707 , \10374 , \10384 );
xor \U$10365 ( \10708 , \10707 , \10387 );
and \U$10366 ( \10709 , \10706 , \10708 );
xor \U$10367 ( \10710 , \10392 , \10394 );
xor \U$10368 ( \10711 , \10710 , \10397 );
and \U$10369 ( \10712 , \10708 , \10711 );
and \U$10370 ( \10713 , \10706 , \10711 );
or \U$10371 ( \10714 , \10709 , \10712 , \10713 );
xor \U$10372 ( \10715 , \10390 , \10400 );
xor \U$10373 ( \10716 , \10715 , \10403 );
and \U$10374 ( \10717 , \10714 , \10716 );
xor \U$10375 ( \10718 , \10061 , \10071 );
xor \U$10376 ( \10719 , \10718 , \10074 );
and \U$10377 ( \10720 , \10716 , \10719 );
and \U$10378 ( \10721 , \10714 , \10719 );
or \U$10379 ( \10722 , \10717 , \10720 , \10721 );
and \U$10380 ( \10723 , \10412 , \10722 );
xor \U$10381 ( \10724 , \10412 , \10722 );
xor \U$10382 ( \10725 , \10714 , \10716 );
xor \U$10383 ( \10726 , \10725 , \10719 );
xor \U$10384 ( \10727 , \10473 , \10477 );
xor \U$10385 ( \10728 , \10727 , \10482 );
xor \U$10386 ( \10729 , \10437 , \10441 );
xor \U$10387 ( \10730 , \10729 , \10446 );
and \U$10388 ( \10731 , \10728 , \10730 );
xor \U$10389 ( \10732 , \10489 , \10493 );
xor \U$10390 ( \10733 , \10732 , \10498 );
and \U$10391 ( \10734 , \10730 , \10733 );
and \U$10392 ( \10735 , \10728 , \10733 );
or \U$10393 ( \10736 , \10731 , \10734 , \10735 );
xor \U$10394 ( \10737 , \10525 , \10529 );
xor \U$10395 ( \10738 , \10737 , \10534 );
xor \U$10396 ( \10739 , \10541 , \10545 );
xor \U$10397 ( \10740 , \10739 , \10550 );
and \U$10398 ( \10741 , \10738 , \10740 );
xor \U$10399 ( \10742 , \10506 , \10510 );
xor \U$10400 ( \10743 , \10742 , \10515 );
and \U$10401 ( \10744 , \10740 , \10743 );
and \U$10402 ( \10745 , \10738 , \10743 );
or \U$10403 ( \10746 , \10741 , \10744 , \10745 );
and \U$10404 ( \10747 , \10736 , \10746 );
and \U$10405 ( \10748 , \8175 , \373 );
and \U$10406 ( \10749 , \8170 , \371 );
nor \U$10407 ( \10750 , \10748 , \10749 );
xnor \U$10408 ( \10751 , \10750 , \380 );
and \U$10409 ( \10752 , \8778 , \391 );
and \U$10410 ( \10753 , \8494 , \389 );
nor \U$10411 ( \10754 , \10752 , \10753 );
xnor \U$10412 ( \10755 , \10754 , \398 );
and \U$10413 ( \10756 , \10751 , \10755 );
and \U$10414 ( \10757 , \9355 , \406 );
and \U$10415 ( \10758 , \9347 , \404 );
nor \U$10416 ( \10759 , \10757 , \10758 );
xnor \U$10417 ( \10760 , \10759 , \413 );
and \U$10418 ( \10761 , \10755 , \10760 );
and \U$10419 ( \10762 , \10751 , \10760 );
or \U$10420 ( \10763 , \10756 , \10761 , \10762 );
buf \U$10421 ( \10764 , RIbb31578_128);
nand \U$10422 ( \10765 , \10764 , \436 );
not \U$10423 ( \10766 , \10765 );
and \U$10424 ( \10767 , \10763 , \10766 );
xor \U$10425 ( \10768 , \10453 , \10457 );
xor \U$10426 ( \10769 , \10768 , \10462 );
and \U$10427 ( \10770 , \10766 , \10769 );
and \U$10428 ( \10771 , \10763 , \10769 );
or \U$10429 ( \10772 , \10767 , \10770 , \10771 );
and \U$10430 ( \10773 , \10746 , \10772 );
and \U$10431 ( \10774 , \10736 , \10772 );
or \U$10432 ( \10775 , \10747 , \10773 , \10774 );
and \U$10433 ( \10776 , \1844 , \4152 );
and \U$10434 ( \10777 , \1839 , \4150 );
nor \U$10435 ( \10778 , \10776 , \10777 );
xnor \U$10436 ( \10779 , \10778 , \4009 );
and \U$10437 ( \10780 , \2174 , \3829 );
and \U$10438 ( \10781 , \2030 , \3827 );
nor \U$10439 ( \10782 , \10780 , \10781 );
xnor \U$10440 ( \10783 , \10782 , \3583 );
and \U$10441 ( \10784 , \10779 , \10783 );
and \U$10442 ( \10785 , \2463 , \3434 );
and \U$10443 ( \10786 , \2438 , \3432 );
nor \U$10444 ( \10787 , \10785 , \10786 );
xnor \U$10445 ( \10788 , \10787 , \3247 );
and \U$10446 ( \10789 , \10783 , \10788 );
and \U$10447 ( \10790 , \10779 , \10788 );
or \U$10448 ( \10791 , \10784 , \10789 , \10790 );
and \U$10449 ( \10792 , \1181 , \5443 );
and \U$10450 ( \10793 , \1176 , \5441 );
nor \U$10451 ( \10794 , \10792 , \10793 );
xnor \U$10452 ( \10795 , \10794 , \5202 );
and \U$10453 ( \10796 , \1412 , \4977 );
and \U$10454 ( \10797 , \1297 , \4975 );
nor \U$10455 ( \10798 , \10796 , \10797 );
xnor \U$10456 ( \10799 , \10798 , \4789 );
and \U$10457 ( \10800 , \10795 , \10799 );
and \U$10458 ( \10801 , \1596 , \4603 );
and \U$10459 ( \10802 , \1588 , \4601 );
nor \U$10460 ( \10803 , \10801 , \10802 );
xnor \U$10461 ( \10804 , \10803 , \4371 );
and \U$10462 ( \10805 , \10799 , \10804 );
and \U$10463 ( \10806 , \10795 , \10804 );
or \U$10464 ( \10807 , \10800 , \10805 , \10806 );
and \U$10465 ( \10808 , \10791 , \10807 );
and \U$10466 ( \10809 , \2804 , \3121 );
and \U$10467 ( \10810 , \2637 , \3119 );
nor \U$10468 ( \10811 , \10809 , \10810 );
xnor \U$10469 ( \10812 , \10811 , \2916 );
and \U$10470 ( \10813 , \3061 , \2715 );
and \U$10471 ( \10814 , \2942 , \2713 );
nor \U$10472 ( \10815 , \10813 , \10814 );
xnor \U$10473 ( \10816 , \10815 , \2566 );
and \U$10474 ( \10817 , \10812 , \10816 );
and \U$10475 ( \10818 , \3686 , \2393 );
and \U$10476 ( \10819 , \3478 , \2391 );
nor \U$10477 ( \10820 , \10818 , \10819 );
xnor \U$10478 ( \10821 , \10820 , \2251 );
and \U$10479 ( \10822 , \10816 , \10821 );
and \U$10480 ( \10823 , \10812 , \10821 );
or \U$10481 ( \10824 , \10817 , \10822 , \10823 );
and \U$10482 ( \10825 , \10807 , \10824 );
and \U$10483 ( \10826 , \10791 , \10824 );
or \U$10484 ( \10827 , \10808 , \10825 , \10826 );
and \U$10485 ( \10828 , \661 , \7035 );
and \U$10486 ( \10829 , \450 , \7033 );
nor \U$10487 ( \10830 , \10828 , \10829 );
xnor \U$10488 ( \10831 , \10830 , \6775 );
and \U$10489 ( \10832 , \785 , \6541 );
and \U$10490 ( \10833 , \722 , \6539 );
nor \U$10491 ( \10834 , \10832 , \10833 );
xnor \U$10492 ( \10835 , \10834 , \6226 );
and \U$10493 ( \10836 , \10831 , \10835 );
and \U$10494 ( \10837 , \1071 , \6032 );
and \U$10495 ( \10838 , \983 , \6030 );
nor \U$10496 ( \10839 , \10837 , \10838 );
xnor \U$10497 ( \10840 , \10839 , \5692 );
and \U$10498 ( \10841 , \10835 , \10840 );
and \U$10499 ( \10842 , \10831 , \10840 );
or \U$10500 ( \10843 , \10836 , \10841 , \10842 );
and \U$10501 ( \10844 , \400 , \8693 );
and \U$10502 ( \10845 , \408 , \8691 );
nor \U$10503 ( \10846 , \10844 , \10845 );
xnor \U$10504 ( \10847 , \10846 , \8322 );
and \U$10505 ( \10848 , \416 , \8131 );
and \U$10506 ( \10849 , \424 , \8129 );
nor \U$10507 ( \10850 , \10848 , \10849 );
xnor \U$10508 ( \10851 , \10850 , \7813 );
and \U$10509 ( \10852 , \10847 , \10851 );
and \U$10510 ( \10853 , \435 , \7564 );
and \U$10511 ( \10854 , \443 , \7562 );
nor \U$10512 ( \10855 , \10853 , \10854 );
xnor \U$10513 ( \10856 , \10855 , \7315 );
and \U$10514 ( \10857 , \10851 , \10856 );
and \U$10515 ( \10858 , \10847 , \10856 );
or \U$10516 ( \10859 , \10852 , \10857 , \10858 );
and \U$10517 ( \10860 , \10843 , \10859 );
and \U$10518 ( \10861 , \351 , \10611 );
and \U$10519 ( \10862 , \359 , \10608 );
nor \U$10520 ( \10863 , \10861 , \10862 );
xnor \U$10521 ( \10864 , \10863 , \9556 );
and \U$10522 ( \10865 , \367 , \9798 );
and \U$10523 ( \10866 , \375 , \9796 );
nor \U$10524 ( \10867 , \10865 , \10866 );
xnor \U$10525 ( \10868 , \10867 , \9559 );
and \U$10526 ( \10869 , \10864 , \10868 );
and \U$10527 ( \10870 , \385 , \9230 );
and \U$10528 ( \10871 , \393 , \9228 );
nor \U$10529 ( \10872 , \10870 , \10871 );
xnor \U$10530 ( \10873 , \10872 , \8920 );
and \U$10531 ( \10874 , \10868 , \10873 );
and \U$10532 ( \10875 , \10864 , \10873 );
or \U$10533 ( \10876 , \10869 , \10874 , \10875 );
and \U$10534 ( \10877 , \10859 , \10876 );
and \U$10535 ( \10878 , \10843 , \10876 );
or \U$10536 ( \10879 , \10860 , \10877 , \10878 );
and \U$10537 ( \10880 , \10827 , \10879 );
and \U$10538 ( \10881 , \5050 , \1351 );
and \U$10539 ( \10882 , \5045 , \1349 );
nor \U$10540 ( \10883 , \10881 , \10882 );
xnor \U$10541 ( \10884 , \10883 , \1238 );
and \U$10542 ( \10885 , \5573 , \1157 );
and \U$10543 ( \10886 , \5314 , \1155 );
nor \U$10544 ( \10887 , \10885 , \10886 );
xnor \U$10545 ( \10888 , \10887 , \1021 );
and \U$10546 ( \10889 , \10884 , \10888 );
and \U$10547 ( \10890 , \5954 , \957 );
and \U$10548 ( \10891 , \5945 , \955 );
nor \U$10549 ( \10892 , \10890 , \10891 );
xnor \U$10550 ( \10893 , \10892 , \879 );
and \U$10551 ( \10894 , \10888 , \10893 );
and \U$10552 ( \10895 , \10884 , \10893 );
or \U$10553 ( \10896 , \10889 , \10894 , \10895 );
and \U$10554 ( \10897 , \3813 , \2097 );
and \U$10555 ( \10898 , \3808 , \2095 );
nor \U$10556 ( \10899 , \10897 , \10898 );
xnor \U$10557 ( \10900 , \10899 , \1960 );
and \U$10558 ( \10901 , \4266 , \1891 );
and \U$10559 ( \10902 , \4069 , \1889 );
nor \U$10560 ( \10903 , \10901 , \10902 );
xnor \U$10561 ( \10904 , \10903 , \1739 );
and \U$10562 ( \10905 , \10900 , \10904 );
and \U$10563 ( \10906 , \4576 , \1623 );
and \U$10564 ( \10907 , \4568 , \1621 );
nor \U$10565 ( \10908 , \10906 , \10907 );
xnor \U$10566 ( \10909 , \10908 , \1467 );
and \U$10567 ( \10910 , \10904 , \10909 );
and \U$10568 ( \10911 , \10900 , \10909 );
or \U$10569 ( \10912 , \10905 , \10910 , \10911 );
and \U$10570 ( \10913 , \10896 , \10912 );
and \U$10571 ( \10914 , \6499 , \793 );
and \U$10572 ( \10915 , \6297 , \791 );
nor \U$10573 ( \10916 , \10914 , \10915 );
xnor \U$10574 ( \10917 , \10916 , \699 );
and \U$10575 ( \10918 , \6974 , \624 );
and \U$10576 ( \10919 , \6802 , \622 );
nor \U$10577 ( \10920 , \10918 , \10919 );
xnor \U$10578 ( \10921 , \10920 , \349 );
and \U$10579 ( \10922 , \10917 , \10921 );
and \U$10580 ( \10923 , \7924 , \357 );
and \U$10581 ( \10924 , \7500 , \355 );
nor \U$10582 ( \10925 , \10923 , \10924 );
xnor \U$10583 ( \10926 , \10925 , \364 );
and \U$10584 ( \10927 , \10921 , \10926 );
and \U$10585 ( \10928 , \10917 , \10926 );
or \U$10586 ( \10929 , \10922 , \10927 , \10928 );
and \U$10587 ( \10930 , \10912 , \10929 );
and \U$10588 ( \10931 , \10896 , \10929 );
or \U$10589 ( \10932 , \10913 , \10930 , \10931 );
and \U$10590 ( \10933 , \10879 , \10932 );
and \U$10591 ( \10934 , \10827 , \10932 );
or \U$10592 ( \10935 , \10880 , \10933 , \10934 );
and \U$10593 ( \10936 , \10775 , \10935 );
xor \U$10594 ( \10937 , \10578 , \10582 );
xor \U$10595 ( \10938 , \10937 , \10587 );
xor \U$10596 ( \10939 , \10594 , \10598 );
xor \U$10597 ( \10940 , \10939 , \10603 );
and \U$10598 ( \10941 , \10938 , \10940 );
xor \U$10599 ( \10942 , \10558 , \10562 );
xor \U$10600 ( \10943 , \10942 , \10567 );
and \U$10601 ( \10944 , \10940 , \10943 );
and \U$10602 ( \10945 , \10938 , \10943 );
or \U$10603 ( \10946 , \10941 , \10944 , \10945 );
xor \U$10604 ( \10947 , \10628 , \10630 );
xor \U$10605 ( \10948 , \10947 , \10633 );
and \U$10606 ( \10949 , \10946 , \10948 );
xor \U$10607 ( \10950 , \10638 , \10640 );
and \U$10608 ( \10951 , \10948 , \10950 );
and \U$10609 ( \10952 , \10946 , \10950 );
or \U$10610 ( \10953 , \10949 , \10951 , \10952 );
and \U$10611 ( \10954 , \10935 , \10953 );
and \U$10612 ( \10955 , \10775 , \10953 );
or \U$10613 ( \10956 , \10936 , \10954 , \10955 );
xor \U$10614 ( \10957 , \10485 , \10501 );
xor \U$10615 ( \10958 , \10957 , \10518 );
xor \U$10616 ( \10959 , \10537 , \10553 );
xor \U$10617 ( \10960 , \10959 , \10570 );
and \U$10618 ( \10961 , \10958 , \10960 );
xor \U$10619 ( \10962 , \10590 , \10606 );
xor \U$10620 ( \10963 , \10962 , \10619 );
and \U$10621 ( \10964 , \10960 , \10963 );
and \U$10622 ( \10965 , \10958 , \10963 );
or \U$10623 ( \10966 , \10961 , \10964 , \10965 );
xor \U$10624 ( \10967 , \10414 , \10416 );
xor \U$10625 ( \10968 , \10967 , \10419 );
xor \U$10626 ( \10969 , \10424 , \10426 );
xor \U$10627 ( \10970 , \10969 , \10429 );
and \U$10628 ( \10971 , \10968 , \10970 );
xnor \U$10629 ( \10972 , \10449 , \10465 );
and \U$10630 ( \10973 , \10970 , \10972 );
and \U$10631 ( \10974 , \10968 , \10972 );
or \U$10632 ( \10975 , \10971 , \10973 , \10974 );
and \U$10633 ( \10976 , \10966 , \10975 );
xor \U$10634 ( \10977 , \10169 , \10185 );
xor \U$10635 ( \10978 , \10977 , \10202 );
and \U$10636 ( \10979 , \10975 , \10978 );
and \U$10637 ( \10980 , \10966 , \10978 );
or \U$10638 ( \10981 , \10976 , \10979 , \10980 );
and \U$10639 ( \10982 , \10956 , \10981 );
xor \U$10640 ( \10983 , \10636 , \10641 );
xor \U$10641 ( \10984 , \10983 , \10644 );
xor \U$10642 ( \10985 , \10652 , \10654 );
xor \U$10643 ( \10986 , \10985 , \10657 );
and \U$10644 ( \10987 , \10984 , \10986 );
xor \U$10645 ( \10988 , \10662 , \10664 );
xor \U$10646 ( \10989 , \10988 , \10667 );
and \U$10647 ( \10990 , \10986 , \10989 );
and \U$10648 ( \10991 , \10984 , \10989 );
or \U$10649 ( \10992 , \10987 , \10990 , \10991 );
and \U$10650 ( \10993 , \10981 , \10992 );
and \U$10651 ( \10994 , \10956 , \10992 );
or \U$10652 ( \10995 , \10982 , \10993 , \10994 );
xor \U$10653 ( \10996 , \10205 , \10257 );
xor \U$10654 ( \10997 , \10996 , \10310 );
xor \U$10655 ( \10998 , \10660 , \10670 );
xor \U$10656 ( \10999 , \10998 , \10673 );
and \U$10657 ( \11000 , \10997 , \10999 );
xor \U$10658 ( \11001 , \10679 , \10681 );
xor \U$10659 ( \11002 , \11001 , \10684 );
and \U$10660 ( \11003 , \10999 , \11002 );
and \U$10661 ( \11004 , \10997 , \11002 );
or \U$10662 ( \11005 , \11000 , \11003 , \11004 );
and \U$10663 ( \11006 , \10995 , \11005 );
xor \U$10664 ( \11007 , \10156 , \10313 );
xor \U$10665 ( \11008 , \11007 , \10331 );
and \U$10666 ( \11009 , \11005 , \11008 );
and \U$10667 ( \11010 , \10995 , \11008 );
or \U$10668 ( \11011 , \11006 , \11009 , \11010 );
xor \U$10669 ( \11012 , \10650 , \10676 );
xor \U$10670 ( \11013 , \11012 , \10687 );
xor \U$10671 ( \11014 , \10692 , \10694 );
xor \U$10672 ( \11015 , \11014 , \10697 );
and \U$10673 ( \11016 , \11013 , \11015 );
and \U$10674 ( \11017 , \11011 , \11016 );
xor \U$10675 ( \11018 , \10376 , \10378 );
xor \U$10676 ( \11019 , \11018 , \10381 );
and \U$10677 ( \11020 , \11016 , \11019 );
and \U$10678 ( \11021 , \11011 , \11019 );
or \U$10679 ( \11022 , \11017 , \11020 , \11021 );
xor \U$10680 ( \11023 , \10334 , \10360 );
xor \U$10681 ( \11024 , \11023 , \10371 );
xor \U$10682 ( \11025 , \10690 , \10700 );
xor \U$10683 ( \11026 , \11025 , \10703 );
and \U$10684 ( \11027 , \11024 , \11026 );
and \U$10685 ( \11028 , \11022 , \11027 );
xor \U$10686 ( \11029 , \10706 , \10708 );
xor \U$10687 ( \11030 , \11029 , \10711 );
and \U$10688 ( \11031 , \11027 , \11030 );
and \U$10689 ( \11032 , \11022 , \11030 );
or \U$10690 ( \11033 , \11028 , \11031 , \11032 );
and \U$10691 ( \11034 , \10726 , \11033 );
xor \U$10692 ( \11035 , \10726 , \11033 );
xor \U$10693 ( \11036 , \11022 , \11027 );
xor \U$10694 ( \11037 , \11036 , \11030 );
and \U$10695 ( \11038 , \9958 , \406 );
and \U$10696 ( \11039 , \9355 , \404 );
nor \U$10697 ( \11040 , \11038 , \11039 );
xnor \U$10698 ( \11041 , \11040 , \413 );
and \U$10699 ( \11042 , \10144 , \422 );
and \U$10700 ( \11043 , \9963 , \420 );
nor \U$10701 ( \11044 , \11042 , \11043 );
xnor \U$10702 ( \11045 , \11044 , \429 );
and \U$10703 ( \11046 , \11041 , \11045 );
nand \U$10704 ( \11047 , \10764 , \439 );
xnor \U$10705 ( \11048 , \11047 , \448 );
and \U$10706 ( \11049 , \11045 , \11048 );
and \U$10707 ( \11050 , \11041 , \11048 );
or \U$10708 ( \11051 , \11046 , \11049 , \11050 );
and \U$10709 ( \11052 , \8170 , \357 );
and \U$10710 ( \11053 , \7924 , \355 );
nor \U$10711 ( \11054 , \11052 , \11053 );
xnor \U$10712 ( \11055 , \11054 , \364 );
and \U$10713 ( \11056 , \8494 , \373 );
and \U$10714 ( \11057 , \8175 , \371 );
nor \U$10715 ( \11058 , \11056 , \11057 );
xnor \U$10716 ( \11059 , \11058 , \380 );
and \U$10717 ( \11060 , \11055 , \11059 );
and \U$10718 ( \11061 , \9347 , \391 );
and \U$10719 ( \11062 , \8778 , \389 );
nor \U$10720 ( \11063 , \11061 , \11062 );
xnor \U$10721 ( \11064 , \11063 , \398 );
and \U$10722 ( \11065 , \11059 , \11064 );
and \U$10723 ( \11066 , \11055 , \11064 );
or \U$10724 ( \11067 , \11060 , \11065 , \11066 );
and \U$10725 ( \11068 , \11051 , \11067 );
and \U$10726 ( \11069 , \9963 , \422 );
and \U$10727 ( \11070 , \9958 , \420 );
nor \U$10728 ( \11071 , \11069 , \11070 );
xnor \U$10729 ( \11072 , \11071 , \429 );
and \U$10730 ( \11073 , \11067 , \11072 );
and \U$10731 ( \11074 , \11051 , \11072 );
or \U$10732 ( \11075 , \11068 , \11073 , \11074 );
and \U$10733 ( \11076 , \10764 , \441 );
and \U$10734 ( \11077 , \10144 , \439 );
nor \U$10735 ( \11078 , \11076 , \11077 );
xnor \U$10736 ( \11079 , \11078 , \448 );
xor \U$10737 ( \11080 , \10917 , \10921 );
xor \U$10738 ( \11081 , \11080 , \10926 );
and \U$10739 ( \11082 , \11079 , \11081 );
xor \U$10740 ( \11083 , \10751 , \10755 );
xor \U$10741 ( \11084 , \11083 , \10760 );
and \U$10742 ( \11085 , \11081 , \11084 );
and \U$10743 ( \11086 , \11079 , \11084 );
or \U$10744 ( \11087 , \11082 , \11085 , \11086 );
and \U$10745 ( \11088 , \11075 , \11087 );
xor \U$10746 ( \11089 , \10884 , \10888 );
xor \U$10747 ( \11090 , \11089 , \10893 );
xor \U$10748 ( \11091 , \10900 , \10904 );
xor \U$10749 ( \11092 , \11091 , \10909 );
and \U$10750 ( \11093 , \11090 , \11092 );
xor \U$10751 ( \11094 , \10812 , \10816 );
xor \U$10752 ( \11095 , \11094 , \10821 );
and \U$10753 ( \11096 , \11092 , \11095 );
and \U$10754 ( \11097 , \11090 , \11095 );
or \U$10755 ( \11098 , \11093 , \11096 , \11097 );
and \U$10756 ( \11099 , \11087 , \11098 );
and \U$10757 ( \11100 , \11075 , \11098 );
or \U$10758 ( \11101 , \11088 , \11099 , \11100 );
and \U$10759 ( \11102 , \5045 , \1623 );
and \U$10760 ( \11103 , \4576 , \1621 );
nor \U$10761 ( \11104 , \11102 , \11103 );
xnor \U$10762 ( \11105 , \11104 , \1467 );
and \U$10763 ( \11106 , \5314 , \1351 );
and \U$10764 ( \11107 , \5050 , \1349 );
nor \U$10765 ( \11108 , \11106 , \11107 );
xnor \U$10766 ( \11109 , \11108 , \1238 );
and \U$10767 ( \11110 , \11105 , \11109 );
and \U$10768 ( \11111 , \5945 , \1157 );
and \U$10769 ( \11112 , \5573 , \1155 );
nor \U$10770 ( \11113 , \11111 , \11112 );
xnor \U$10771 ( \11114 , \11113 , \1021 );
and \U$10772 ( \11115 , \11109 , \11114 );
and \U$10773 ( \11116 , \11105 , \11114 );
or \U$10774 ( \11117 , \11110 , \11115 , \11116 );
and \U$10775 ( \11118 , \3808 , \2393 );
and \U$10776 ( \11119 , \3686 , \2391 );
nor \U$10777 ( \11120 , \11118 , \11119 );
xnor \U$10778 ( \11121 , \11120 , \2251 );
and \U$10779 ( \11122 , \4069 , \2097 );
and \U$10780 ( \11123 , \3813 , \2095 );
nor \U$10781 ( \11124 , \11122 , \11123 );
xnor \U$10782 ( \11125 , \11124 , \1960 );
and \U$10783 ( \11126 , \11121 , \11125 );
and \U$10784 ( \11127 , \4568 , \1891 );
and \U$10785 ( \11128 , \4266 , \1889 );
nor \U$10786 ( \11129 , \11127 , \11128 );
xnor \U$10787 ( \11130 , \11129 , \1739 );
and \U$10788 ( \11131 , \11125 , \11130 );
and \U$10789 ( \11132 , \11121 , \11130 );
or \U$10790 ( \11133 , \11126 , \11131 , \11132 );
and \U$10791 ( \11134 , \11117 , \11133 );
and \U$10792 ( \11135 , \6297 , \957 );
and \U$10793 ( \11136 , \5954 , \955 );
nor \U$10794 ( \11137 , \11135 , \11136 );
xnor \U$10795 ( \11138 , \11137 , \879 );
and \U$10796 ( \11139 , \6802 , \793 );
and \U$10797 ( \11140 , \6499 , \791 );
nor \U$10798 ( \11141 , \11139 , \11140 );
xnor \U$10799 ( \11142 , \11141 , \699 );
and \U$10800 ( \11143 , \11138 , \11142 );
and \U$10801 ( \11144 , \7500 , \624 );
and \U$10802 ( \11145 , \6974 , \622 );
nor \U$10803 ( \11146 , \11144 , \11145 );
xnor \U$10804 ( \11147 , \11146 , \349 );
and \U$10805 ( \11148 , \11142 , \11147 );
and \U$10806 ( \11149 , \11138 , \11147 );
or \U$10807 ( \11150 , \11143 , \11148 , \11149 );
and \U$10808 ( \11151 , \11133 , \11150 );
and \U$10809 ( \11152 , \11117 , \11150 );
or \U$10810 ( \11153 , \11134 , \11151 , \11152 );
and \U$10811 ( \11154 , \450 , \7564 );
and \U$10812 ( \11155 , \435 , \7562 );
nor \U$10813 ( \11156 , \11154 , \11155 );
xnor \U$10814 ( \11157 , \11156 , \7315 );
and \U$10815 ( \11158 , \722 , \7035 );
and \U$10816 ( \11159 , \661 , \7033 );
nor \U$10817 ( \11160 , \11158 , \11159 );
xnor \U$10818 ( \11161 , \11160 , \6775 );
and \U$10819 ( \11162 , \11157 , \11161 );
and \U$10820 ( \11163 , \983 , \6541 );
and \U$10821 ( \11164 , \785 , \6539 );
nor \U$10822 ( \11165 , \11163 , \11164 );
xnor \U$10823 ( \11166 , \11165 , \6226 );
and \U$10824 ( \11167 , \11161 , \11166 );
and \U$10825 ( \11168 , \11157 , \11166 );
or \U$10826 ( \11169 , \11162 , \11167 , \11168 );
and \U$10827 ( \11170 , \375 , \10611 );
and \U$10828 ( \11171 , \351 , \10608 );
nor \U$10829 ( \11172 , \11170 , \11171 );
xnor \U$10830 ( \11173 , \11172 , \9556 );
and \U$10831 ( \11174 , \393 , \9798 );
and \U$10832 ( \11175 , \367 , \9796 );
nor \U$10833 ( \11176 , \11174 , \11175 );
xnor \U$10834 ( \11177 , \11176 , \9559 );
and \U$10835 ( \11178 , \11173 , \11177 );
and \U$10836 ( \11179 , \11177 , \448 );
and \U$10837 ( \11180 , \11173 , \448 );
or \U$10838 ( \11181 , \11178 , \11179 , \11180 );
and \U$10839 ( \11182 , \11169 , \11181 );
and \U$10840 ( \11183 , \408 , \9230 );
and \U$10841 ( \11184 , \385 , \9228 );
nor \U$10842 ( \11185 , \11183 , \11184 );
xnor \U$10843 ( \11186 , \11185 , \8920 );
and \U$10844 ( \11187 , \424 , \8693 );
and \U$10845 ( \11188 , \400 , \8691 );
nor \U$10846 ( \11189 , \11187 , \11188 );
xnor \U$10847 ( \11190 , \11189 , \8322 );
and \U$10848 ( \11191 , \11186 , \11190 );
and \U$10849 ( \11192 , \443 , \8131 );
and \U$10850 ( \11193 , \416 , \8129 );
nor \U$10851 ( \11194 , \11192 , \11193 );
xnor \U$10852 ( \11195 , \11194 , \7813 );
and \U$10853 ( \11196 , \11190 , \11195 );
and \U$10854 ( \11197 , \11186 , \11195 );
or \U$10855 ( \11198 , \11191 , \11196 , \11197 );
and \U$10856 ( \11199 , \11181 , \11198 );
and \U$10857 ( \11200 , \11169 , \11198 );
or \U$10858 ( \11201 , \11182 , \11199 , \11200 );
and \U$10859 ( \11202 , \11153 , \11201 );
and \U$10860 ( \11203 , \1839 , \4603 );
and \U$10861 ( \11204 , \1596 , \4601 );
nor \U$10862 ( \11205 , \11203 , \11204 );
xnor \U$10863 ( \11206 , \11205 , \4371 );
and \U$10864 ( \11207 , \2030 , \4152 );
and \U$10865 ( \11208 , \1844 , \4150 );
nor \U$10866 ( \11209 , \11207 , \11208 );
xnor \U$10867 ( \11210 , \11209 , \4009 );
and \U$10868 ( \11211 , \11206 , \11210 );
and \U$10869 ( \11212 , \2438 , \3829 );
and \U$10870 ( \11213 , \2174 , \3827 );
nor \U$10871 ( \11214 , \11212 , \11213 );
xnor \U$10872 ( \11215 , \11214 , \3583 );
and \U$10873 ( \11216 , \11210 , \11215 );
and \U$10874 ( \11217 , \11206 , \11215 );
or \U$10875 ( \11218 , \11211 , \11216 , \11217 );
and \U$10876 ( \11219 , \1176 , \6032 );
and \U$10877 ( \11220 , \1071 , \6030 );
nor \U$10878 ( \11221 , \11219 , \11220 );
xnor \U$10879 ( \11222 , \11221 , \5692 );
and \U$10880 ( \11223 , \1297 , \5443 );
and \U$10881 ( \11224 , \1181 , \5441 );
nor \U$10882 ( \11225 , \11223 , \11224 );
xnor \U$10883 ( \11226 , \11225 , \5202 );
and \U$10884 ( \11227 , \11222 , \11226 );
and \U$10885 ( \11228 , \1588 , \4977 );
and \U$10886 ( \11229 , \1412 , \4975 );
nor \U$10887 ( \11230 , \11228 , \11229 );
xnor \U$10888 ( \11231 , \11230 , \4789 );
and \U$10889 ( \11232 , \11226 , \11231 );
and \U$10890 ( \11233 , \11222 , \11231 );
or \U$10891 ( \11234 , \11227 , \11232 , \11233 );
and \U$10892 ( \11235 , \11218 , \11234 );
and \U$10893 ( \11236 , \2637 , \3434 );
and \U$10894 ( \11237 , \2463 , \3432 );
nor \U$10895 ( \11238 , \11236 , \11237 );
xnor \U$10896 ( \11239 , \11238 , \3247 );
and \U$10897 ( \11240 , \2942 , \3121 );
and \U$10898 ( \11241 , \2804 , \3119 );
nor \U$10899 ( \11242 , \11240 , \11241 );
xnor \U$10900 ( \11243 , \11242 , \2916 );
and \U$10901 ( \11244 , \11239 , \11243 );
and \U$10902 ( \11245 , \3478 , \2715 );
and \U$10903 ( \11246 , \3061 , \2713 );
nor \U$10904 ( \11247 , \11245 , \11246 );
xnor \U$10905 ( \11248 , \11247 , \2566 );
and \U$10906 ( \11249 , \11243 , \11248 );
and \U$10907 ( \11250 , \11239 , \11248 );
or \U$10908 ( \11251 , \11244 , \11249 , \11250 );
and \U$10909 ( \11252 , \11234 , \11251 );
and \U$10910 ( \11253 , \11218 , \11251 );
or \U$10911 ( \11254 , \11235 , \11252 , \11253 );
and \U$10912 ( \11255 , \11201 , \11254 );
and \U$10913 ( \11256 , \11153 , \11254 );
or \U$10914 ( \11257 , \11202 , \11255 , \11256 );
and \U$10915 ( \11258 , \11101 , \11257 );
xor \U$10916 ( \11259 , \10779 , \10783 );
xor \U$10917 ( \11260 , \11259 , \10788 );
xor \U$10918 ( \11261 , \10795 , \10799 );
xor \U$10919 ( \11262 , \11261 , \10804 );
and \U$10920 ( \11263 , \11260 , \11262 );
xor \U$10921 ( \11264 , \10831 , \10835 );
xor \U$10922 ( \11265 , \11264 , \10840 );
and \U$10923 ( \11266 , \11262 , \11265 );
and \U$10924 ( \11267 , \11260 , \11265 );
or \U$10925 ( \11268 , \11263 , \11266 , \11267 );
xor \U$10926 ( \11269 , \10847 , \10851 );
xor \U$10927 ( \11270 , \11269 , \10856 );
xor \U$10928 ( \11271 , \10864 , \10868 );
xor \U$10929 ( \11272 , \11271 , \10873 );
and \U$10930 ( \11273 , \11270 , \11272 );
and \U$10931 ( \11274 , \11268 , \11273 );
xor \U$10932 ( \11275 , \10614 , \10618 );
and \U$10933 ( \11276 , \11273 , \11275 );
and \U$10934 ( \11277 , \11268 , \11275 );
or \U$10935 ( \11278 , \11274 , \11276 , \11277 );
and \U$10936 ( \11279 , \11257 , \11278 );
and \U$10937 ( \11280 , \11101 , \11278 );
or \U$10938 ( \11281 , \11258 , \11279 , \11280 );
xor \U$10939 ( \11282 , \10791 , \10807 );
xor \U$10940 ( \11283 , \11282 , \10824 );
xor \U$10941 ( \11284 , \10896 , \10912 );
xor \U$10942 ( \11285 , \11284 , \10929 );
and \U$10943 ( \11286 , \11283 , \11285 );
xor \U$10944 ( \11287 , \10763 , \10766 );
xor \U$10945 ( \11288 , \11287 , \10769 );
and \U$10946 ( \11289 , \11285 , \11288 );
and \U$10947 ( \11290 , \11283 , \11288 );
or \U$10948 ( \11291 , \11286 , \11289 , \11290 );
xor \U$10949 ( \11292 , \10938 , \10940 );
xor \U$10950 ( \11293 , \11292 , \10943 );
xor \U$10951 ( \11294 , \10728 , \10730 );
xor \U$10952 ( \11295 , \11294 , \10733 );
and \U$10953 ( \11296 , \11293 , \11295 );
xor \U$10954 ( \11297 , \10738 , \10740 );
xor \U$10955 ( \11298 , \11297 , \10743 );
and \U$10956 ( \11299 , \11295 , \11298 );
and \U$10957 ( \11300 , \11293 , \11298 );
or \U$10958 ( \11301 , \11296 , \11299 , \11300 );
and \U$10959 ( \11302 , \11291 , \11301 );
xor \U$10960 ( \11303 , \10958 , \10960 );
xor \U$10961 ( \11304 , \11303 , \10963 );
and \U$10962 ( \11305 , \11301 , \11304 );
and \U$10963 ( \11306 , \11291 , \11304 );
or \U$10964 ( \11307 , \11302 , \11305 , \11306 );
and \U$10965 ( \11308 , \11281 , \11307 );
xor \U$10966 ( \11309 , \10736 , \10746 );
xor \U$10967 ( \11310 , \11309 , \10772 );
xor \U$10968 ( \11311 , \10968 , \10970 );
xor \U$10969 ( \11312 , \11311 , \10972 );
and \U$10970 ( \11313 , \11310 , \11312 );
xor \U$10971 ( \11314 , \10946 , \10948 );
xor \U$10972 ( \11315 , \11314 , \10950 );
and \U$10973 ( \11316 , \11312 , \11315 );
and \U$10974 ( \11317 , \11310 , \11315 );
or \U$10975 ( \11318 , \11313 , \11316 , \11317 );
and \U$10976 ( \11319 , \11307 , \11318 );
and \U$10977 ( \11320 , \11281 , \11318 );
or \U$10978 ( \11321 , \11308 , \11319 , \11320 );
xor \U$10979 ( \11322 , \10422 , \10432 );
xor \U$10980 ( \11323 , \11322 , \10466 );
xor \U$10981 ( \11324 , \10521 , \10573 );
xor \U$10982 ( \11325 , \11324 , \10622 );
and \U$10983 ( \11326 , \11323 , \11325 );
xor \U$10984 ( \11327 , \10984 , \10986 );
xor \U$10985 ( \11328 , \11327 , \10989 );
and \U$10986 ( \11329 , \11325 , \11328 );
and \U$10987 ( \11330 , \11323 , \11328 );
or \U$10988 ( \11331 , \11326 , \11329 , \11330 );
and \U$10989 ( \11332 , \11321 , \11331 );
xor \U$10990 ( \11333 , \10469 , \10625 );
xor \U$10991 ( \11334 , \11333 , \10647 );
and \U$10992 ( \11335 , \11331 , \11334 );
and \U$10993 ( \11336 , \11321 , \11334 );
or \U$10994 ( \11337 , \11332 , \11335 , \11336 );
xor \U$10995 ( \11338 , \10995 , \11005 );
xor \U$10996 ( \11339 , \11338 , \11008 );
and \U$10997 ( \11340 , \11337 , \11339 );
xor \U$10998 ( \11341 , \11013 , \11015 );
and \U$10999 ( \11342 , \11339 , \11341 );
and \U$11000 ( \11343 , \11337 , \11341 );
or \U$11001 ( \11344 , \11340 , \11342 , \11343 );
xor \U$11002 ( \11345 , \11011 , \11016 );
xor \U$11003 ( \11346 , \11345 , \11019 );
and \U$11004 ( \11347 , \11344 , \11346 );
xor \U$11005 ( \11348 , \11024 , \11026 );
and \U$11006 ( \11349 , \11346 , \11348 );
and \U$11007 ( \11350 , \11344 , \11348 );
or \U$11008 ( \11351 , \11347 , \11349 , \11350 );
and \U$11009 ( \11352 , \11037 , \11351 );
xor \U$11010 ( \11353 , \11037 , \11351 );
xor \U$11011 ( \11354 , \11344 , \11346 );
xor \U$11012 ( \11355 , \11354 , \11348 );
and \U$11013 ( \11356 , \416 , \8693 );
and \U$11014 ( \11357 , \424 , \8691 );
nor \U$11015 ( \11358 , \11356 , \11357 );
xnor \U$11016 ( \11359 , \11358 , \8322 );
and \U$11017 ( \11360 , \435 , \8131 );
and \U$11018 ( \11361 , \443 , \8129 );
nor \U$11019 ( \11362 , \11360 , \11361 );
xnor \U$11020 ( \11363 , \11362 , \7813 );
and \U$11021 ( \11364 , \11359 , \11363 );
and \U$11022 ( \11365 , \661 , \7564 );
and \U$11023 ( \11366 , \450 , \7562 );
nor \U$11024 ( \11367 , \11365 , \11366 );
xnor \U$11025 ( \11368 , \11367 , \7315 );
and \U$11026 ( \11369 , \11363 , \11368 );
and \U$11027 ( \11370 , \11359 , \11368 );
or \U$11028 ( \11371 , \11364 , \11369 , \11370 );
and \U$11029 ( \11372 , \367 , \10611 );
and \U$11030 ( \11373 , \375 , \10608 );
nor \U$11031 ( \11374 , \11372 , \11373 );
xnor \U$11032 ( \11375 , \11374 , \9556 );
and \U$11033 ( \11376 , \385 , \9798 );
and \U$11034 ( \11377 , \393 , \9796 );
nor \U$11035 ( \11378 , \11376 , \11377 );
xnor \U$11036 ( \11379 , \11378 , \9559 );
and \U$11037 ( \11380 , \11375 , \11379 );
and \U$11038 ( \11381 , \400 , \9230 );
and \U$11039 ( \11382 , \408 , \9228 );
nor \U$11040 ( \11383 , \11381 , \11382 );
xnor \U$11041 ( \11384 , \11383 , \8920 );
and \U$11042 ( \11385 , \11379 , \11384 );
and \U$11043 ( \11386 , \11375 , \11384 );
or \U$11044 ( \11387 , \11380 , \11385 , \11386 );
and \U$11045 ( \11388 , \11371 , \11387 );
and \U$11046 ( \11389 , \785 , \7035 );
and \U$11047 ( \11390 , \722 , \7033 );
nor \U$11048 ( \11391 , \11389 , \11390 );
xnor \U$11049 ( \11392 , \11391 , \6775 );
and \U$11050 ( \11393 , \1071 , \6541 );
and \U$11051 ( \11394 , \983 , \6539 );
nor \U$11052 ( \11395 , \11393 , \11394 );
xnor \U$11053 ( \11396 , \11395 , \6226 );
and \U$11054 ( \11397 , \11392 , \11396 );
and \U$11055 ( \11398 , \1181 , \6032 );
and \U$11056 ( \11399 , \1176 , \6030 );
nor \U$11057 ( \11400 , \11398 , \11399 );
xnor \U$11058 ( \11401 , \11400 , \5692 );
and \U$11059 ( \11402 , \11396 , \11401 );
and \U$11060 ( \11403 , \11392 , \11401 );
or \U$11061 ( \11404 , \11397 , \11402 , \11403 );
and \U$11062 ( \11405 , \11387 , \11404 );
and \U$11063 ( \11406 , \11371 , \11404 );
or \U$11064 ( \11407 , \11388 , \11405 , \11406 );
and \U$11065 ( \11408 , \5573 , \1351 );
and \U$11066 ( \11409 , \5314 , \1349 );
nor \U$11067 ( \11410 , \11408 , \11409 );
xnor \U$11068 ( \11411 , \11410 , \1238 );
and \U$11069 ( \11412 , \5954 , \1157 );
and \U$11070 ( \11413 , \5945 , \1155 );
nor \U$11071 ( \11414 , \11412 , \11413 );
xnor \U$11072 ( \11415 , \11414 , \1021 );
and \U$11073 ( \11416 , \11411 , \11415 );
and \U$11074 ( \11417 , \6499 , \957 );
and \U$11075 ( \11418 , \6297 , \955 );
nor \U$11076 ( \11419 , \11417 , \11418 );
xnor \U$11077 ( \11420 , \11419 , \879 );
and \U$11078 ( \11421 , \11415 , \11420 );
and \U$11079 ( \11422 , \11411 , \11420 );
or \U$11080 ( \11423 , \11416 , \11421 , \11422 );
and \U$11081 ( \11424 , \6974 , \793 );
and \U$11082 ( \11425 , \6802 , \791 );
nor \U$11083 ( \11426 , \11424 , \11425 );
xnor \U$11084 ( \11427 , \11426 , \699 );
and \U$11085 ( \11428 , \7924 , \624 );
and \U$11086 ( \11429 , \7500 , \622 );
nor \U$11087 ( \11430 , \11428 , \11429 );
xnor \U$11088 ( \11431 , \11430 , \349 );
and \U$11089 ( \11432 , \11427 , \11431 );
and \U$11090 ( \11433 , \8175 , \357 );
and \U$11091 ( \11434 , \8170 , \355 );
nor \U$11092 ( \11435 , \11433 , \11434 );
xnor \U$11093 ( \11436 , \11435 , \364 );
and \U$11094 ( \11437 , \11431 , \11436 );
and \U$11095 ( \11438 , \11427 , \11436 );
or \U$11096 ( \11439 , \11432 , \11437 , \11438 );
and \U$11097 ( \11440 , \11423 , \11439 );
and \U$11098 ( \11441 , \4266 , \2097 );
and \U$11099 ( \11442 , \4069 , \2095 );
nor \U$11100 ( \11443 , \11441 , \11442 );
xnor \U$11101 ( \11444 , \11443 , \1960 );
and \U$11102 ( \11445 , \4576 , \1891 );
and \U$11103 ( \11446 , \4568 , \1889 );
nor \U$11104 ( \11447 , \11445 , \11446 );
xnor \U$11105 ( \11448 , \11447 , \1739 );
and \U$11106 ( \11449 , \11444 , \11448 );
and \U$11107 ( \11450 , \5050 , \1623 );
and \U$11108 ( \11451 , \5045 , \1621 );
nor \U$11109 ( \11452 , \11450 , \11451 );
xnor \U$11110 ( \11453 , \11452 , \1467 );
and \U$11111 ( \11454 , \11448 , \11453 );
and \U$11112 ( \11455 , \11444 , \11453 );
or \U$11113 ( \11456 , \11449 , \11454 , \11455 );
and \U$11114 ( \11457 , \11439 , \11456 );
and \U$11115 ( \11458 , \11423 , \11456 );
or \U$11116 ( \11459 , \11440 , \11457 , \11458 );
and \U$11117 ( \11460 , \11407 , \11459 );
and \U$11118 ( \11461 , \1412 , \5443 );
and \U$11119 ( \11462 , \1297 , \5441 );
nor \U$11120 ( \11463 , \11461 , \11462 );
xnor \U$11121 ( \11464 , \11463 , \5202 );
and \U$11122 ( \11465 , \1596 , \4977 );
and \U$11123 ( \11466 , \1588 , \4975 );
nor \U$11124 ( \11467 , \11465 , \11466 );
xnor \U$11125 ( \11468 , \11467 , \4789 );
and \U$11126 ( \11469 , \11464 , \11468 );
and \U$11127 ( \11470 , \1844 , \4603 );
and \U$11128 ( \11471 , \1839 , \4601 );
nor \U$11129 ( \11472 , \11470 , \11471 );
xnor \U$11130 ( \11473 , \11472 , \4371 );
and \U$11131 ( \11474 , \11468 , \11473 );
and \U$11132 ( \11475 , \11464 , \11473 );
or \U$11133 ( \11476 , \11469 , \11474 , \11475 );
and \U$11134 ( \11477 , \3061 , \3121 );
and \U$11135 ( \11478 , \2942 , \3119 );
nor \U$11136 ( \11479 , \11477 , \11478 );
xnor \U$11137 ( \11480 , \11479 , \2916 );
and \U$11138 ( \11481 , \3686 , \2715 );
and \U$11139 ( \11482 , \3478 , \2713 );
nor \U$11140 ( \11483 , \11481 , \11482 );
xnor \U$11141 ( \11484 , \11483 , \2566 );
and \U$11142 ( \11485 , \11480 , \11484 );
and \U$11143 ( \11486 , \3813 , \2393 );
and \U$11144 ( \11487 , \3808 , \2391 );
nor \U$11145 ( \11488 , \11486 , \11487 );
xnor \U$11146 ( \11489 , \11488 , \2251 );
and \U$11147 ( \11490 , \11484 , \11489 );
and \U$11148 ( \11491 , \11480 , \11489 );
or \U$11149 ( \11492 , \11485 , \11490 , \11491 );
and \U$11150 ( \11493 , \11476 , \11492 );
and \U$11151 ( \11494 , \2174 , \4152 );
and \U$11152 ( \11495 , \2030 , \4150 );
nor \U$11153 ( \11496 , \11494 , \11495 );
xnor \U$11154 ( \11497 , \11496 , \4009 );
and \U$11155 ( \11498 , \2463 , \3829 );
and \U$11156 ( \11499 , \2438 , \3827 );
nor \U$11157 ( \11500 , \11498 , \11499 );
xnor \U$11158 ( \11501 , \11500 , \3583 );
and \U$11159 ( \11502 , \11497 , \11501 );
and \U$11160 ( \11503 , \2804 , \3434 );
and \U$11161 ( \11504 , \2637 , \3432 );
nor \U$11162 ( \11505 , \11503 , \11504 );
xnor \U$11163 ( \11506 , \11505 , \3247 );
and \U$11164 ( \11507 , \11501 , \11506 );
and \U$11165 ( \11508 , \11497 , \11506 );
or \U$11166 ( \11509 , \11502 , \11507 , \11508 );
and \U$11167 ( \11510 , \11492 , \11509 );
and \U$11168 ( \11511 , \11476 , \11509 );
or \U$11169 ( \11512 , \11493 , \11510 , \11511 );
and \U$11170 ( \11513 , \11459 , \11512 );
and \U$11171 ( \11514 , \11407 , \11512 );
or \U$11172 ( \11515 , \11460 , \11513 , \11514 );
xor \U$11173 ( \11516 , \11206 , \11210 );
xor \U$11174 ( \11517 , \11516 , \11215 );
xor \U$11175 ( \11518 , \11222 , \11226 );
xor \U$11176 ( \11519 , \11518 , \11231 );
and \U$11177 ( \11520 , \11517 , \11519 );
xor \U$11178 ( \11521 , \11239 , \11243 );
xor \U$11179 ( \11522 , \11521 , \11248 );
and \U$11180 ( \11523 , \11519 , \11522 );
and \U$11181 ( \11524 , \11517 , \11522 );
or \U$11182 ( \11525 , \11520 , \11523 , \11524 );
and \U$11183 ( \11526 , \8778 , \373 );
and \U$11184 ( \11527 , \8494 , \371 );
nor \U$11185 ( \11528 , \11526 , \11527 );
xnor \U$11186 ( \11529 , \11528 , \380 );
and \U$11187 ( \11530 , \9355 , \391 );
and \U$11188 ( \11531 , \9347 , \389 );
nor \U$11189 ( \11532 , \11530 , \11531 );
xnor \U$11190 ( \11533 , \11532 , \398 );
and \U$11191 ( \11534 , \11529 , \11533 );
and \U$11192 ( \11535 , \9963 , \406 );
and \U$11193 ( \11536 , \9958 , \404 );
nor \U$11194 ( \11537 , \11535 , \11536 );
xnor \U$11195 ( \11538 , \11537 , \413 );
and \U$11196 ( \11539 , \11533 , \11538 );
and \U$11197 ( \11540 , \11529 , \11538 );
or \U$11198 ( \11541 , \11534 , \11539 , \11540 );
xor \U$11199 ( \11542 , \11041 , \11045 );
xor \U$11200 ( \11543 , \11542 , \11048 );
and \U$11201 ( \11544 , \11541 , \11543 );
xor \U$11202 ( \11545 , \11055 , \11059 );
xor \U$11203 ( \11546 , \11545 , \11064 );
and \U$11204 ( \11547 , \11543 , \11546 );
and \U$11205 ( \11548 , \11541 , \11546 );
or \U$11206 ( \11549 , \11544 , \11547 , \11548 );
and \U$11207 ( \11550 , \11525 , \11549 );
xor \U$11208 ( \11551 , \11105 , \11109 );
xor \U$11209 ( \11552 , \11551 , \11114 );
xor \U$11210 ( \11553 , \11121 , \11125 );
xor \U$11211 ( \11554 , \11553 , \11130 );
and \U$11212 ( \11555 , \11552 , \11554 );
xor \U$11213 ( \11556 , \11138 , \11142 );
xor \U$11214 ( \11557 , \11556 , \11147 );
and \U$11215 ( \11558 , \11554 , \11557 );
and \U$11216 ( \11559 , \11552 , \11557 );
or \U$11217 ( \11560 , \11555 , \11558 , \11559 );
and \U$11218 ( \11561 , \11549 , \11560 );
and \U$11219 ( \11562 , \11525 , \11560 );
or \U$11220 ( \11563 , \11550 , \11561 , \11562 );
and \U$11221 ( \11564 , \11515 , \11563 );
xor \U$11222 ( \11565 , \11157 , \11161 );
xor \U$11223 ( \11566 , \11565 , \11166 );
xor \U$11224 ( \11567 , \11173 , \11177 );
xor \U$11225 ( \11568 , \11567 , \448 );
and \U$11226 ( \11569 , \11566 , \11568 );
xor \U$11227 ( \11570 , \11186 , \11190 );
xor \U$11228 ( \11571 , \11570 , \11195 );
and \U$11229 ( \11572 , \11568 , \11571 );
and \U$11230 ( \11573 , \11566 , \11571 );
or \U$11231 ( \11574 , \11569 , \11572 , \11573 );
xor \U$11232 ( \11575 , \11260 , \11262 );
xor \U$11233 ( \11576 , \11575 , \11265 );
and \U$11234 ( \11577 , \11574 , \11576 );
xor \U$11235 ( \11578 , \11270 , \11272 );
and \U$11236 ( \11579 , \11576 , \11578 );
and \U$11237 ( \11580 , \11574 , \11578 );
or \U$11238 ( \11581 , \11577 , \11579 , \11580 );
and \U$11239 ( \11582 , \11563 , \11581 );
and \U$11240 ( \11583 , \11515 , \11581 );
or \U$11241 ( \11584 , \11564 , \11582 , \11583 );
xor \U$11242 ( \11585 , \11117 , \11133 );
xor \U$11243 ( \11586 , \11585 , \11150 );
xor \U$11244 ( \11587 , \11169 , \11181 );
xor \U$11245 ( \11588 , \11587 , \11198 );
and \U$11246 ( \11589 , \11586 , \11588 );
xor \U$11247 ( \11590 , \11218 , \11234 );
xor \U$11248 ( \11591 , \11590 , \11251 );
and \U$11249 ( \11592 , \11588 , \11591 );
and \U$11250 ( \11593 , \11586 , \11591 );
or \U$11251 ( \11594 , \11589 , \11592 , \11593 );
xor \U$11252 ( \11595 , \11051 , \11067 );
xor \U$11253 ( \11596 , \11595 , \11072 );
xor \U$11254 ( \11597 , \11079 , \11081 );
xor \U$11255 ( \11598 , \11597 , \11084 );
and \U$11256 ( \11599 , \11596 , \11598 );
xor \U$11257 ( \11600 , \11090 , \11092 );
xor \U$11258 ( \11601 , \11600 , \11095 );
and \U$11259 ( \11602 , \11598 , \11601 );
and \U$11260 ( \11603 , \11596 , \11601 );
or \U$11261 ( \11604 , \11599 , \11602 , \11603 );
and \U$11262 ( \11605 , \11594 , \11604 );
xor \U$11263 ( \11606 , \10843 , \10859 );
xor \U$11264 ( \11607 , \11606 , \10876 );
and \U$11265 ( \11608 , \11604 , \11607 );
and \U$11266 ( \11609 , \11594 , \11607 );
or \U$11267 ( \11610 , \11605 , \11608 , \11609 );
and \U$11268 ( \11611 , \11584 , \11610 );
xor \U$11269 ( \11612 , \11283 , \11285 );
xor \U$11270 ( \11613 , \11612 , \11288 );
xor \U$11271 ( \11614 , \11293 , \11295 );
xor \U$11272 ( \11615 , \11614 , \11298 );
and \U$11273 ( \11616 , \11613 , \11615 );
xor \U$11274 ( \11617 , \11268 , \11273 );
xor \U$11275 ( \11618 , \11617 , \11275 );
and \U$11276 ( \11619 , \11615 , \11618 );
and \U$11277 ( \11620 , \11613 , \11618 );
or \U$11278 ( \11621 , \11616 , \11619 , \11620 );
and \U$11279 ( \11622 , \11610 , \11621 );
and \U$11280 ( \11623 , \11584 , \11621 );
or \U$11281 ( \11624 , \11611 , \11622 , \11623 );
xor \U$11282 ( \11625 , \10827 , \10879 );
xor \U$11283 ( \11626 , \11625 , \10932 );
xor \U$11284 ( \11627 , \11291 , \11301 );
xor \U$11285 ( \11628 , \11627 , \11304 );
and \U$11286 ( \11629 , \11626 , \11628 );
xor \U$11287 ( \11630 , \11310 , \11312 );
xor \U$11288 ( \11631 , \11630 , \11315 );
and \U$11289 ( \11632 , \11628 , \11631 );
and \U$11290 ( \11633 , \11626 , \11631 );
or \U$11291 ( \11634 , \11629 , \11632 , \11633 );
and \U$11292 ( \11635 , \11624 , \11634 );
xor \U$11293 ( \11636 , \10966 , \10975 );
xor \U$11294 ( \11637 , \11636 , \10978 );
and \U$11295 ( \11638 , \11634 , \11637 );
and \U$11296 ( \11639 , \11624 , \11637 );
or \U$11297 ( \11640 , \11635 , \11638 , \11639 );
xor \U$11298 ( \11641 , \10775 , \10935 );
xor \U$11299 ( \11642 , \11641 , \10953 );
xor \U$11300 ( \11643 , \11281 , \11307 );
xor \U$11301 ( \11644 , \11643 , \11318 );
and \U$11302 ( \11645 , \11642 , \11644 );
xor \U$11303 ( \11646 , \11323 , \11325 );
xor \U$11304 ( \11647 , \11646 , \11328 );
and \U$11305 ( \11648 , \11644 , \11647 );
and \U$11306 ( \11649 , \11642 , \11647 );
or \U$11307 ( \11650 , \11645 , \11648 , \11649 );
and \U$11308 ( \11651 , \11640 , \11650 );
xor \U$11309 ( \11652 , \10997 , \10999 );
xor \U$11310 ( \11653 , \11652 , \11002 );
and \U$11311 ( \11654 , \11650 , \11653 );
and \U$11312 ( \11655 , \11640 , \11653 );
or \U$11313 ( \11656 , \11651 , \11654 , \11655 );
xor \U$11314 ( \11657 , \10956 , \10981 );
xor \U$11315 ( \11658 , \11657 , \10992 );
xor \U$11316 ( \11659 , \11321 , \11331 );
xor \U$11317 ( \11660 , \11659 , \11334 );
and \U$11318 ( \11661 , \11658 , \11660 );
and \U$11319 ( \11662 , \11656 , \11661 );
xor \U$11320 ( \11663 , \11337 , \11339 );
xor \U$11321 ( \11664 , \11663 , \11341 );
and \U$11322 ( \11665 , \11661 , \11664 );
and \U$11323 ( \11666 , \11656 , \11664 );
or \U$11324 ( \11667 , \11662 , \11665 , \11666 );
and \U$11325 ( \11668 , \11355 , \11667 );
xor \U$11326 ( \11669 , \11355 , \11667 );
xor \U$11327 ( \11670 , \11656 , \11661 );
xor \U$11328 ( \11671 , \11670 , \11664 );
and \U$11329 ( \11672 , \6802 , \957 );
and \U$11330 ( \11673 , \6499 , \955 );
nor \U$11331 ( \11674 , \11672 , \11673 );
xnor \U$11332 ( \11675 , \11674 , \879 );
and \U$11333 ( \11676 , \7500 , \793 );
and \U$11334 ( \11677 , \6974 , \791 );
nor \U$11335 ( \11678 , \11676 , \11677 );
xnor \U$11336 ( \11679 , \11678 , \699 );
and \U$11337 ( \11680 , \11675 , \11679 );
and \U$11338 ( \11681 , \8170 , \624 );
and \U$11339 ( \11682 , \7924 , \622 );
nor \U$11340 ( \11683 , \11681 , \11682 );
xnor \U$11341 ( \11684 , \11683 , \349 );
and \U$11342 ( \11685 , \11679 , \11684 );
and \U$11343 ( \11686 , \11675 , \11684 );
or \U$11344 ( \11687 , \11680 , \11685 , \11686 );
and \U$11345 ( \11688 , \4069 , \2393 );
and \U$11346 ( \11689 , \3813 , \2391 );
nor \U$11347 ( \11690 , \11688 , \11689 );
xnor \U$11348 ( \11691 , \11690 , \2251 );
and \U$11349 ( \11692 , \4568 , \2097 );
and \U$11350 ( \11693 , \4266 , \2095 );
nor \U$11351 ( \11694 , \11692 , \11693 );
xnor \U$11352 ( \11695 , \11694 , \1960 );
and \U$11353 ( \11696 , \11691 , \11695 );
and \U$11354 ( \11697 , \5045 , \1891 );
and \U$11355 ( \11698 , \4576 , \1889 );
nor \U$11356 ( \11699 , \11697 , \11698 );
xnor \U$11357 ( \11700 , \11699 , \1739 );
and \U$11358 ( \11701 , \11695 , \11700 );
and \U$11359 ( \11702 , \11691 , \11700 );
or \U$11360 ( \11703 , \11696 , \11701 , \11702 );
and \U$11361 ( \11704 , \11687 , \11703 );
and \U$11362 ( \11705 , \5314 , \1623 );
and \U$11363 ( \11706 , \5050 , \1621 );
nor \U$11364 ( \11707 , \11705 , \11706 );
xnor \U$11365 ( \11708 , \11707 , \1467 );
and \U$11366 ( \11709 , \5945 , \1351 );
and \U$11367 ( \11710 , \5573 , \1349 );
nor \U$11368 ( \11711 , \11709 , \11710 );
xnor \U$11369 ( \11712 , \11711 , \1238 );
and \U$11370 ( \11713 , \11708 , \11712 );
and \U$11371 ( \11714 , \6297 , \1157 );
and \U$11372 ( \11715 , \5954 , \1155 );
nor \U$11373 ( \11716 , \11714 , \11715 );
xnor \U$11374 ( \11717 , \11716 , \1021 );
and \U$11375 ( \11718 , \11712 , \11717 );
and \U$11376 ( \11719 , \11708 , \11717 );
or \U$11377 ( \11720 , \11713 , \11718 , \11719 );
and \U$11378 ( \11721 , \11703 , \11720 );
and \U$11379 ( \11722 , \11687 , \11720 );
or \U$11380 ( \11723 , \11704 , \11721 , \11722 );
and \U$11381 ( \11724 , \722 , \7564 );
and \U$11382 ( \11725 , \661 , \7562 );
nor \U$11383 ( \11726 , \11724 , \11725 );
xnor \U$11384 ( \11727 , \11726 , \7315 );
and \U$11385 ( \11728 , \983 , \7035 );
and \U$11386 ( \11729 , \785 , \7033 );
nor \U$11387 ( \11730 , \11728 , \11729 );
xnor \U$11388 ( \11731 , \11730 , \6775 );
and \U$11389 ( \11732 , \11727 , \11731 );
and \U$11390 ( \11733 , \1176 , \6541 );
and \U$11391 ( \11734 , \1071 , \6539 );
nor \U$11392 ( \11735 , \11733 , \11734 );
xnor \U$11393 ( \11736 , \11735 , \6226 );
and \U$11394 ( \11737 , \11731 , \11736 );
and \U$11395 ( \11738 , \11727 , \11736 );
or \U$11396 ( \11739 , \11732 , \11737 , \11738 );
and \U$11397 ( \11740 , \424 , \9230 );
and \U$11398 ( \11741 , \400 , \9228 );
nor \U$11399 ( \11742 , \11740 , \11741 );
xnor \U$11400 ( \11743 , \11742 , \8920 );
and \U$11401 ( \11744 , \443 , \8693 );
and \U$11402 ( \11745 , \416 , \8691 );
nor \U$11403 ( \11746 , \11744 , \11745 );
xnor \U$11404 ( \11747 , \11746 , \8322 );
and \U$11405 ( \11748 , \11743 , \11747 );
and \U$11406 ( \11749 , \450 , \8131 );
and \U$11407 ( \11750 , \435 , \8129 );
nor \U$11408 ( \11751 , \11749 , \11750 );
xnor \U$11409 ( \11752 , \11751 , \7813 );
and \U$11410 ( \11753 , \11747 , \11752 );
and \U$11411 ( \11754 , \11743 , \11752 );
or \U$11412 ( \11755 , \11748 , \11753 , \11754 );
and \U$11413 ( \11756 , \11739 , \11755 );
and \U$11414 ( \11757 , \393 , \10611 );
and \U$11415 ( \11758 , \367 , \10608 );
nor \U$11416 ( \11759 , \11757 , \11758 );
xnor \U$11417 ( \11760 , \11759 , \9556 );
and \U$11418 ( \11761 , \408 , \9798 );
and \U$11419 ( \11762 , \385 , \9796 );
nor \U$11420 ( \11763 , \11761 , \11762 );
xnor \U$11421 ( \11764 , \11763 , \9559 );
and \U$11422 ( \11765 , \11760 , \11764 );
and \U$11423 ( \11766 , \11764 , \429 );
and \U$11424 ( \11767 , \11760 , \429 );
or \U$11425 ( \11768 , \11765 , \11766 , \11767 );
and \U$11426 ( \11769 , \11755 , \11768 );
and \U$11427 ( \11770 , \11739 , \11768 );
or \U$11428 ( \11771 , \11756 , \11769 , \11770 );
and \U$11429 ( \11772 , \11723 , \11771 );
and \U$11430 ( \11773 , \1297 , \6032 );
and \U$11431 ( \11774 , \1181 , \6030 );
nor \U$11432 ( \11775 , \11773 , \11774 );
xnor \U$11433 ( \11776 , \11775 , \5692 );
and \U$11434 ( \11777 , \1588 , \5443 );
and \U$11435 ( \11778 , \1412 , \5441 );
nor \U$11436 ( \11779 , \11777 , \11778 );
xnor \U$11437 ( \11780 , \11779 , \5202 );
and \U$11438 ( \11781 , \11776 , \11780 );
and \U$11439 ( \11782 , \1839 , \4977 );
and \U$11440 ( \11783 , \1596 , \4975 );
nor \U$11441 ( \11784 , \11782 , \11783 );
xnor \U$11442 ( \11785 , \11784 , \4789 );
and \U$11443 ( \11786 , \11780 , \11785 );
and \U$11444 ( \11787 , \11776 , \11785 );
or \U$11445 ( \11788 , \11781 , \11786 , \11787 );
and \U$11446 ( \11789 , \2030 , \4603 );
and \U$11447 ( \11790 , \1844 , \4601 );
nor \U$11448 ( \11791 , \11789 , \11790 );
xnor \U$11449 ( \11792 , \11791 , \4371 );
and \U$11450 ( \11793 , \2438 , \4152 );
and \U$11451 ( \11794 , \2174 , \4150 );
nor \U$11452 ( \11795 , \11793 , \11794 );
xnor \U$11453 ( \11796 , \11795 , \4009 );
and \U$11454 ( \11797 , \11792 , \11796 );
and \U$11455 ( \11798 , \2637 , \3829 );
and \U$11456 ( \11799 , \2463 , \3827 );
nor \U$11457 ( \11800 , \11798 , \11799 );
xnor \U$11458 ( \11801 , \11800 , \3583 );
and \U$11459 ( \11802 , \11796 , \11801 );
and \U$11460 ( \11803 , \11792 , \11801 );
or \U$11461 ( \11804 , \11797 , \11802 , \11803 );
and \U$11462 ( \11805 , \11788 , \11804 );
and \U$11463 ( \11806 , \2942 , \3434 );
and \U$11464 ( \11807 , \2804 , \3432 );
nor \U$11465 ( \11808 , \11806 , \11807 );
xnor \U$11466 ( \11809 , \11808 , \3247 );
and \U$11467 ( \11810 , \3478 , \3121 );
and \U$11468 ( \11811 , \3061 , \3119 );
nor \U$11469 ( \11812 , \11810 , \11811 );
xnor \U$11470 ( \11813 , \11812 , \2916 );
and \U$11471 ( \11814 , \11809 , \11813 );
and \U$11472 ( \11815 , \3808 , \2715 );
and \U$11473 ( \11816 , \3686 , \2713 );
nor \U$11474 ( \11817 , \11815 , \11816 );
xnor \U$11475 ( \11818 , \11817 , \2566 );
and \U$11476 ( \11819 , \11813 , \11818 );
and \U$11477 ( \11820 , \11809 , \11818 );
or \U$11478 ( \11821 , \11814 , \11819 , \11820 );
and \U$11479 ( \11822 , \11804 , \11821 );
and \U$11480 ( \11823 , \11788 , \11821 );
or \U$11481 ( \11824 , \11805 , \11822 , \11823 );
and \U$11482 ( \11825 , \11771 , \11824 );
and \U$11483 ( \11826 , \11723 , \11824 );
or \U$11484 ( \11827 , \11772 , \11825 , \11826 );
and \U$11485 ( \11828 , \8494 , \357 );
and \U$11486 ( \11829 , \8175 , \355 );
nor \U$11487 ( \11830 , \11828 , \11829 );
xnor \U$11488 ( \11831 , \11830 , \364 );
and \U$11489 ( \11832 , \9347 , \373 );
and \U$11490 ( \11833 , \8778 , \371 );
nor \U$11491 ( \11834 , \11832 , \11833 );
xnor \U$11492 ( \11835 , \11834 , \380 );
and \U$11493 ( \11836 , \11831 , \11835 );
and \U$11494 ( \11837 , \9958 , \391 );
and \U$11495 ( \11838 , \9355 , \389 );
nor \U$11496 ( \11839 , \11837 , \11838 );
xnor \U$11497 ( \11840 , \11839 , \398 );
and \U$11498 ( \11841 , \11835 , \11840 );
and \U$11499 ( \11842 , \11831 , \11840 );
or \U$11500 ( \11843 , \11836 , \11841 , \11842 );
and \U$11501 ( \11844 , \10144 , \406 );
and \U$11502 ( \11845 , \9963 , \404 );
nor \U$11503 ( \11846 , \11844 , \11845 );
xnor \U$11504 ( \11847 , \11846 , \413 );
nand \U$11505 ( \11848 , \10764 , \420 );
xnor \U$11506 ( \11849 , \11848 , \429 );
and \U$11507 ( \11850 , \11847 , \11849 );
and \U$11508 ( \11851 , \11843 , \11850 );
and \U$11509 ( \11852 , \10764 , \422 );
and \U$11510 ( \11853 , \10144 , \420 );
nor \U$11511 ( \11854 , \11852 , \11853 );
xnor \U$11512 ( \11855 , \11854 , \429 );
and \U$11513 ( \11856 , \11850 , \11855 );
and \U$11514 ( \11857 , \11843 , \11855 );
or \U$11515 ( \11858 , \11851 , \11856 , \11857 );
xor \U$11516 ( \11859 , \11444 , \11448 );
xor \U$11517 ( \11860 , \11859 , \11453 );
xor \U$11518 ( \11861 , \11480 , \11484 );
xor \U$11519 ( \11862 , \11861 , \11489 );
and \U$11520 ( \11863 , \11860 , \11862 );
xor \U$11521 ( \11864 , \11497 , \11501 );
xor \U$11522 ( \11865 , \11864 , \11506 );
and \U$11523 ( \11866 , \11862 , \11865 );
and \U$11524 ( \11867 , \11860 , \11865 );
or \U$11525 ( \11868 , \11863 , \11866 , \11867 );
and \U$11526 ( \11869 , \11858 , \11868 );
xor \U$11527 ( \11870 , \11411 , \11415 );
xor \U$11528 ( \11871 , \11870 , \11420 );
xor \U$11529 ( \11872 , \11427 , \11431 );
xor \U$11530 ( \11873 , \11872 , \11436 );
and \U$11531 ( \11874 , \11871 , \11873 );
xor \U$11532 ( \11875 , \11529 , \11533 );
xor \U$11533 ( \11876 , \11875 , \11538 );
and \U$11534 ( \11877 , \11873 , \11876 );
and \U$11535 ( \11878 , \11871 , \11876 );
or \U$11536 ( \11879 , \11874 , \11877 , \11878 );
and \U$11537 ( \11880 , \11868 , \11879 );
and \U$11538 ( \11881 , \11858 , \11879 );
or \U$11539 ( \11882 , \11869 , \11880 , \11881 );
and \U$11540 ( \11883 , \11827 , \11882 );
xor \U$11541 ( \11884 , \11359 , \11363 );
xor \U$11542 ( \11885 , \11884 , \11368 );
xor \U$11543 ( \11886 , \11464 , \11468 );
xor \U$11544 ( \11887 , \11886 , \11473 );
and \U$11545 ( \11888 , \11885 , \11887 );
xor \U$11546 ( \11889 , \11392 , \11396 );
xor \U$11547 ( \11890 , \11889 , \11401 );
and \U$11548 ( \11891 , \11887 , \11890 );
and \U$11549 ( \11892 , \11885 , \11890 );
or \U$11550 ( \11893 , \11888 , \11891 , \11892 );
xor \U$11551 ( \11894 , \11566 , \11568 );
xor \U$11552 ( \11895 , \11894 , \11571 );
and \U$11553 ( \11896 , \11893 , \11895 );
xor \U$11554 ( \11897 , \11517 , \11519 );
xor \U$11555 ( \11898 , \11897 , \11522 );
and \U$11556 ( \11899 , \11895 , \11898 );
and \U$11557 ( \11900 , \11893 , \11898 );
or \U$11558 ( \11901 , \11896 , \11899 , \11900 );
and \U$11559 ( \11902 , \11882 , \11901 );
and \U$11560 ( \11903 , \11827 , \11901 );
or \U$11561 ( \11904 , \11883 , \11902 , \11903 );
xor \U$11562 ( \11905 , \11423 , \11439 );
xor \U$11563 ( \11906 , \11905 , \11456 );
xor \U$11564 ( \11907 , \11541 , \11543 );
xor \U$11565 ( \11908 , \11907 , \11546 );
and \U$11566 ( \11909 , \11906 , \11908 );
xor \U$11567 ( \11910 , \11552 , \11554 );
xor \U$11568 ( \11911 , \11910 , \11557 );
and \U$11569 ( \11912 , \11908 , \11911 );
and \U$11570 ( \11913 , \11906 , \11911 );
or \U$11571 ( \11914 , \11909 , \11912 , \11913 );
xor \U$11572 ( \11915 , \11586 , \11588 );
xor \U$11573 ( \11916 , \11915 , \11591 );
and \U$11574 ( \11917 , \11914 , \11916 );
xor \U$11575 ( \11918 , \11596 , \11598 );
xor \U$11576 ( \11919 , \11918 , \11601 );
and \U$11577 ( \11920 , \11916 , \11919 );
and \U$11578 ( \11921 , \11914 , \11919 );
or \U$11579 ( \11922 , \11917 , \11920 , \11921 );
and \U$11580 ( \11923 , \11904 , \11922 );
xor \U$11581 ( \11924 , \11407 , \11459 );
xor \U$11582 ( \11925 , \11924 , \11512 );
xor \U$11583 ( \11926 , \11525 , \11549 );
xor \U$11584 ( \11927 , \11926 , \11560 );
and \U$11585 ( \11928 , \11925 , \11927 );
xor \U$11586 ( \11929 , \11574 , \11576 );
xor \U$11587 ( \11930 , \11929 , \11578 );
and \U$11588 ( \11931 , \11927 , \11930 );
and \U$11589 ( \11932 , \11925 , \11930 );
or \U$11590 ( \11933 , \11928 , \11931 , \11932 );
and \U$11591 ( \11934 , \11922 , \11933 );
and \U$11592 ( \11935 , \11904 , \11933 );
or \U$11593 ( \11936 , \11923 , \11934 , \11935 );
xor \U$11594 ( \11937 , \11075 , \11087 );
xor \U$11595 ( \11938 , \11937 , \11098 );
xor \U$11596 ( \11939 , \11153 , \11201 );
xor \U$11597 ( \11940 , \11939 , \11254 );
and \U$11598 ( \11941 , \11938 , \11940 );
xor \U$11599 ( \11942 , \11613 , \11615 );
xor \U$11600 ( \11943 , \11942 , \11618 );
and \U$11601 ( \11944 , \11940 , \11943 );
and \U$11602 ( \11945 , \11938 , \11943 );
or \U$11603 ( \11946 , \11941 , \11944 , \11945 );
and \U$11604 ( \11947 , \11936 , \11946 );
xor \U$11605 ( \11948 , \11101 , \11257 );
xor \U$11606 ( \11949 , \11948 , \11278 );
and \U$11607 ( \11950 , \11946 , \11949 );
and \U$11608 ( \11951 , \11936 , \11949 );
or \U$11609 ( \11952 , \11947 , \11950 , \11951 );
xor \U$11610 ( \11953 , \11624 , \11634 );
xor \U$11611 ( \11954 , \11953 , \11637 );
and \U$11612 ( \11955 , \11952 , \11954 );
xor \U$11613 ( \11956 , \11642 , \11644 );
xor \U$11614 ( \11957 , \11956 , \11647 );
and \U$11615 ( \11958 , \11954 , \11957 );
and \U$11616 ( \11959 , \11952 , \11957 );
or \U$11617 ( \11960 , \11955 , \11958 , \11959 );
xor \U$11618 ( \11961 , \11640 , \11650 );
xor \U$11619 ( \11962 , \11961 , \11653 );
and \U$11620 ( \11963 , \11960 , \11962 );
xor \U$11621 ( \11964 , \11658 , \11660 );
and \U$11622 ( \11965 , \11962 , \11964 );
and \U$11623 ( \11966 , \11960 , \11964 );
or \U$11624 ( \11967 , \11963 , \11965 , \11966 );
and \U$11625 ( \11968 , \11671 , \11967 );
xor \U$11626 ( \11969 , \11671 , \11967 );
xor \U$11627 ( \11970 , \11960 , \11962 );
xor \U$11628 ( \11971 , \11970 , \11964 );
xor \U$11629 ( \11972 , \11675 , \11679 );
xor \U$11630 ( \11973 , \11972 , \11684 );
xor \U$11631 ( \11974 , \11691 , \11695 );
xor \U$11632 ( \11975 , \11974 , \11700 );
and \U$11633 ( \11976 , \11973 , \11975 );
xor \U$11634 ( \11977 , \11708 , \11712 );
xor \U$11635 ( \11978 , \11977 , \11717 );
and \U$11636 ( \11979 , \11975 , \11978 );
and \U$11637 ( \11980 , \11973 , \11978 );
or \U$11638 ( \11981 , \11976 , \11979 , \11980 );
xor \U$11639 ( \11982 , \11776 , \11780 );
xor \U$11640 ( \11983 , \11982 , \11785 );
xor \U$11641 ( \11984 , \11792 , \11796 );
xor \U$11642 ( \11985 , \11984 , \11801 );
and \U$11643 ( \11986 , \11983 , \11985 );
xor \U$11644 ( \11987 , \11809 , \11813 );
xor \U$11645 ( \11988 , \11987 , \11818 );
and \U$11646 ( \11989 , \11985 , \11988 );
and \U$11647 ( \11990 , \11983 , \11988 );
or \U$11648 ( \11991 , \11986 , \11989 , \11990 );
and \U$11649 ( \11992 , \11981 , \11991 );
and \U$11650 ( \11993 , \9355 , \373 );
and \U$11651 ( \11994 , \9347 , \371 );
nor \U$11652 ( \11995 , \11993 , \11994 );
xnor \U$11653 ( \11996 , \11995 , \380 );
and \U$11654 ( \11997 , \9963 , \391 );
and \U$11655 ( \11998 , \9958 , \389 );
nor \U$11656 ( \11999 , \11997 , \11998 );
xnor \U$11657 ( \12000 , \11999 , \398 );
and \U$11658 ( \12001 , \11996 , \12000 );
and \U$11659 ( \12002 , \10764 , \406 );
and \U$11660 ( \12003 , \10144 , \404 );
nor \U$11661 ( \12004 , \12002 , \12003 );
xnor \U$11662 ( \12005 , \12004 , \413 );
and \U$11663 ( \12006 , \12000 , \12005 );
and \U$11664 ( \12007 , \11996 , \12005 );
or \U$11665 ( \12008 , \12001 , \12006 , \12007 );
xor \U$11666 ( \12009 , \11831 , \11835 );
xor \U$11667 ( \12010 , \12009 , \11840 );
and \U$11668 ( \12011 , \12008 , \12010 );
xor \U$11669 ( \12012 , \11847 , \11849 );
and \U$11670 ( \12013 , \12010 , \12012 );
and \U$11671 ( \12014 , \12008 , \12012 );
or \U$11672 ( \12015 , \12011 , \12013 , \12014 );
and \U$11673 ( \12016 , \11991 , \12015 );
and \U$11674 ( \12017 , \11981 , \12015 );
or \U$11675 ( \12018 , \11992 , \12016 , \12017 );
and \U$11676 ( \12019 , \3686 , \3121 );
and \U$11677 ( \12020 , \3478 , \3119 );
nor \U$11678 ( \12021 , \12019 , \12020 );
xnor \U$11679 ( \12022 , \12021 , \2916 );
and \U$11680 ( \12023 , \3813 , \2715 );
and \U$11681 ( \12024 , \3808 , \2713 );
nor \U$11682 ( \12025 , \12023 , \12024 );
xnor \U$11683 ( \12026 , \12025 , \2566 );
and \U$11684 ( \12027 , \12022 , \12026 );
and \U$11685 ( \12028 , \4266 , \2393 );
and \U$11686 ( \12029 , \4069 , \2391 );
nor \U$11687 ( \12030 , \12028 , \12029 );
xnor \U$11688 ( \12031 , \12030 , \2251 );
and \U$11689 ( \12032 , \12026 , \12031 );
and \U$11690 ( \12033 , \12022 , \12031 );
or \U$11691 ( \12034 , \12027 , \12032 , \12033 );
and \U$11692 ( \12035 , \1596 , \5443 );
and \U$11693 ( \12036 , \1588 , \5441 );
nor \U$11694 ( \12037 , \12035 , \12036 );
xnor \U$11695 ( \12038 , \12037 , \5202 );
and \U$11696 ( \12039 , \1844 , \4977 );
and \U$11697 ( \12040 , \1839 , \4975 );
nor \U$11698 ( \12041 , \12039 , \12040 );
xnor \U$11699 ( \12042 , \12041 , \4789 );
and \U$11700 ( \12043 , \12038 , \12042 );
and \U$11701 ( \12044 , \2174 , \4603 );
and \U$11702 ( \12045 , \2030 , \4601 );
nor \U$11703 ( \12046 , \12044 , \12045 );
xnor \U$11704 ( \12047 , \12046 , \4371 );
and \U$11705 ( \12048 , \12042 , \12047 );
and \U$11706 ( \12049 , \12038 , \12047 );
or \U$11707 ( \12050 , \12043 , \12048 , \12049 );
and \U$11708 ( \12051 , \12034 , \12050 );
and \U$11709 ( \12052 , \2463 , \4152 );
and \U$11710 ( \12053 , \2438 , \4150 );
nor \U$11711 ( \12054 , \12052 , \12053 );
xnor \U$11712 ( \12055 , \12054 , \4009 );
and \U$11713 ( \12056 , \2804 , \3829 );
and \U$11714 ( \12057 , \2637 , \3827 );
nor \U$11715 ( \12058 , \12056 , \12057 );
xnor \U$11716 ( \12059 , \12058 , \3583 );
and \U$11717 ( \12060 , \12055 , \12059 );
and \U$11718 ( \12061 , \3061 , \3434 );
and \U$11719 ( \12062 , \2942 , \3432 );
nor \U$11720 ( \12063 , \12061 , \12062 );
xnor \U$11721 ( \12064 , \12063 , \3247 );
and \U$11722 ( \12065 , \12059 , \12064 );
and \U$11723 ( \12066 , \12055 , \12064 );
or \U$11724 ( \12067 , \12060 , \12065 , \12066 );
and \U$11725 ( \12068 , \12050 , \12067 );
and \U$11726 ( \12069 , \12034 , \12067 );
or \U$11727 ( \12070 , \12051 , \12068 , \12069 );
and \U$11728 ( \12071 , \1071 , \7035 );
and \U$11729 ( \12072 , \983 , \7033 );
nor \U$11730 ( \12073 , \12071 , \12072 );
xnor \U$11731 ( \12074 , \12073 , \6775 );
and \U$11732 ( \12075 , \1181 , \6541 );
and \U$11733 ( \12076 , \1176 , \6539 );
nor \U$11734 ( \12077 , \12075 , \12076 );
xnor \U$11735 ( \12078 , \12077 , \6226 );
and \U$11736 ( \12079 , \12074 , \12078 );
and \U$11737 ( \12080 , \1412 , \6032 );
and \U$11738 ( \12081 , \1297 , \6030 );
nor \U$11739 ( \12082 , \12080 , \12081 );
xnor \U$11740 ( \12083 , \12082 , \5692 );
and \U$11741 ( \12084 , \12078 , \12083 );
and \U$11742 ( \12085 , \12074 , \12083 );
or \U$11743 ( \12086 , \12079 , \12084 , \12085 );
and \U$11744 ( \12087 , \385 , \10611 );
and \U$11745 ( \12088 , \393 , \10608 );
nor \U$11746 ( \12089 , \12087 , \12088 );
xnor \U$11747 ( \12090 , \12089 , \9556 );
and \U$11748 ( \12091 , \400 , \9798 );
and \U$11749 ( \12092 , \408 , \9796 );
nor \U$11750 ( \12093 , \12091 , \12092 );
xnor \U$11751 ( \12094 , \12093 , \9559 );
and \U$11752 ( \12095 , \12090 , \12094 );
and \U$11753 ( \12096 , \416 , \9230 );
and \U$11754 ( \12097 , \424 , \9228 );
nor \U$11755 ( \12098 , \12096 , \12097 );
xnor \U$11756 ( \12099 , \12098 , \8920 );
and \U$11757 ( \12100 , \12094 , \12099 );
and \U$11758 ( \12101 , \12090 , \12099 );
or \U$11759 ( \12102 , \12095 , \12100 , \12101 );
and \U$11760 ( \12103 , \12086 , \12102 );
and \U$11761 ( \12104 , \435 , \8693 );
and \U$11762 ( \12105 , \443 , \8691 );
nor \U$11763 ( \12106 , \12104 , \12105 );
xnor \U$11764 ( \12107 , \12106 , \8322 );
and \U$11765 ( \12108 , \661 , \8131 );
and \U$11766 ( \12109 , \450 , \8129 );
nor \U$11767 ( \12110 , \12108 , \12109 );
xnor \U$11768 ( \12111 , \12110 , \7813 );
and \U$11769 ( \12112 , \12107 , \12111 );
and \U$11770 ( \12113 , \785 , \7564 );
and \U$11771 ( \12114 , \722 , \7562 );
nor \U$11772 ( \12115 , \12113 , \12114 );
xnor \U$11773 ( \12116 , \12115 , \7315 );
and \U$11774 ( \12117 , \12111 , \12116 );
and \U$11775 ( \12118 , \12107 , \12116 );
or \U$11776 ( \12119 , \12112 , \12117 , \12118 );
and \U$11777 ( \12120 , \12102 , \12119 );
and \U$11778 ( \12121 , \12086 , \12119 );
or \U$11779 ( \12122 , \12103 , \12120 , \12121 );
and \U$11780 ( \12123 , \12070 , \12122 );
and \U$11781 ( \12124 , \4576 , \2097 );
and \U$11782 ( \12125 , \4568 , \2095 );
nor \U$11783 ( \12126 , \12124 , \12125 );
xnor \U$11784 ( \12127 , \12126 , \1960 );
and \U$11785 ( \12128 , \5050 , \1891 );
and \U$11786 ( \12129 , \5045 , \1889 );
nor \U$11787 ( \12130 , \12128 , \12129 );
xnor \U$11788 ( \12131 , \12130 , \1739 );
and \U$11789 ( \12132 , \12127 , \12131 );
and \U$11790 ( \12133 , \5573 , \1623 );
and \U$11791 ( \12134 , \5314 , \1621 );
nor \U$11792 ( \12135 , \12133 , \12134 );
xnor \U$11793 ( \12136 , \12135 , \1467 );
and \U$11794 ( \12137 , \12131 , \12136 );
and \U$11795 ( \12138 , \12127 , \12136 );
or \U$11796 ( \12139 , \12132 , \12137 , \12138 );
and \U$11797 ( \12140 , \7924 , \793 );
and \U$11798 ( \12141 , \7500 , \791 );
nor \U$11799 ( \12142 , \12140 , \12141 );
xnor \U$11800 ( \12143 , \12142 , \699 );
and \U$11801 ( \12144 , \8175 , \624 );
and \U$11802 ( \12145 , \8170 , \622 );
nor \U$11803 ( \12146 , \12144 , \12145 );
xnor \U$11804 ( \12147 , \12146 , \349 );
and \U$11805 ( \12148 , \12143 , \12147 );
and \U$11806 ( \12149 , \8778 , \357 );
and \U$11807 ( \12150 , \8494 , \355 );
nor \U$11808 ( \12151 , \12149 , \12150 );
xnor \U$11809 ( \12152 , \12151 , \364 );
and \U$11810 ( \12153 , \12147 , \12152 );
and \U$11811 ( \12154 , \12143 , \12152 );
or \U$11812 ( \12155 , \12148 , \12153 , \12154 );
and \U$11813 ( \12156 , \12139 , \12155 );
and \U$11814 ( \12157 , \5954 , \1351 );
and \U$11815 ( \12158 , \5945 , \1349 );
nor \U$11816 ( \12159 , \12157 , \12158 );
xnor \U$11817 ( \12160 , \12159 , \1238 );
and \U$11818 ( \12161 , \6499 , \1157 );
and \U$11819 ( \12162 , \6297 , \1155 );
nor \U$11820 ( \12163 , \12161 , \12162 );
xnor \U$11821 ( \12164 , \12163 , \1021 );
and \U$11822 ( \12165 , \12160 , \12164 );
and \U$11823 ( \12166 , \6974 , \957 );
and \U$11824 ( \12167 , \6802 , \955 );
nor \U$11825 ( \12168 , \12166 , \12167 );
xnor \U$11826 ( \12169 , \12168 , \879 );
and \U$11827 ( \12170 , \12164 , \12169 );
and \U$11828 ( \12171 , \12160 , \12169 );
or \U$11829 ( \12172 , \12165 , \12170 , \12171 );
and \U$11830 ( \12173 , \12155 , \12172 );
and \U$11831 ( \12174 , \12139 , \12172 );
or \U$11832 ( \12175 , \12156 , \12173 , \12174 );
and \U$11833 ( \12176 , \12122 , \12175 );
and \U$11834 ( \12177 , \12070 , \12175 );
or \U$11835 ( \12178 , \12123 , \12176 , \12177 );
and \U$11836 ( \12179 , \12018 , \12178 );
xor \U$11837 ( \12180 , \11727 , \11731 );
xor \U$11838 ( \12181 , \12180 , \11736 );
xor \U$11839 ( \12182 , \11743 , \11747 );
xor \U$11840 ( \12183 , \12182 , \11752 );
and \U$11841 ( \12184 , \12181 , \12183 );
xor \U$11842 ( \12185 , \11760 , \11764 );
xor \U$11843 ( \12186 , \12185 , \429 );
and \U$11844 ( \12187 , \12183 , \12186 );
and \U$11845 ( \12188 , \12181 , \12186 );
or \U$11846 ( \12189 , \12184 , \12187 , \12188 );
xor \U$11847 ( \12190 , \11375 , \11379 );
xor \U$11848 ( \12191 , \12190 , \11384 );
and \U$11849 ( \12192 , \12189 , \12191 );
xor \U$11850 ( \12193 , \11885 , \11887 );
xor \U$11851 ( \12194 , \12193 , \11890 );
and \U$11852 ( \12195 , \12191 , \12194 );
and \U$11853 ( \12196 , \12189 , \12194 );
or \U$11854 ( \12197 , \12192 , \12195 , \12196 );
and \U$11855 ( \12198 , \12178 , \12197 );
and \U$11856 ( \12199 , \12018 , \12197 );
or \U$11857 ( \12200 , \12179 , \12198 , \12199 );
xor \U$11858 ( \12201 , \11687 , \11703 );
xor \U$11859 ( \12202 , \12201 , \11720 );
xor \U$11860 ( \12203 , \11739 , \11755 );
xor \U$11861 ( \12204 , \12203 , \11768 );
and \U$11862 ( \12205 , \12202 , \12204 );
xor \U$11863 ( \12206 , \11788 , \11804 );
xor \U$11864 ( \12207 , \12206 , \11821 );
and \U$11865 ( \12208 , \12204 , \12207 );
and \U$11866 ( \12209 , \12202 , \12207 );
or \U$11867 ( \12210 , \12205 , \12208 , \12209 );
xor \U$11868 ( \12211 , \11843 , \11850 );
xor \U$11869 ( \12212 , \12211 , \11855 );
xor \U$11870 ( \12213 , \11860 , \11862 );
xor \U$11871 ( \12214 , \12213 , \11865 );
and \U$11872 ( \12215 , \12212 , \12214 );
xor \U$11873 ( \12216 , \11871 , \11873 );
xor \U$11874 ( \12217 , \12216 , \11876 );
and \U$11875 ( \12218 , \12214 , \12217 );
and \U$11876 ( \12219 , \12212 , \12217 );
or \U$11877 ( \12220 , \12215 , \12218 , \12219 );
and \U$11878 ( \12221 , \12210 , \12220 );
xor \U$11879 ( \12222 , \11476 , \11492 );
xor \U$11880 ( \12223 , \12222 , \11509 );
and \U$11881 ( \12224 , \12220 , \12223 );
and \U$11882 ( \12225 , \12210 , \12223 );
or \U$11883 ( \12226 , \12221 , \12224 , \12225 );
and \U$11884 ( \12227 , \12200 , \12226 );
xor \U$11885 ( \12228 , \11371 , \11387 );
xor \U$11886 ( \12229 , \12228 , \11404 );
xor \U$11887 ( \12230 , \11906 , \11908 );
xor \U$11888 ( \12231 , \12230 , \11911 );
and \U$11889 ( \12232 , \12229 , \12231 );
xor \U$11890 ( \12233 , \11893 , \11895 );
xor \U$11891 ( \12234 , \12233 , \11898 );
and \U$11892 ( \12235 , \12231 , \12234 );
and \U$11893 ( \12236 , \12229 , \12234 );
or \U$11894 ( \12237 , \12232 , \12235 , \12236 );
and \U$11895 ( \12238 , \12226 , \12237 );
and \U$11896 ( \12239 , \12200 , \12237 );
or \U$11897 ( \12240 , \12227 , \12238 , \12239 );
xor \U$11898 ( \12241 , \11827 , \11882 );
xor \U$11899 ( \12242 , \12241 , \11901 );
xor \U$11900 ( \12243 , \11914 , \11916 );
xor \U$11901 ( \12244 , \12243 , \11919 );
and \U$11902 ( \12245 , \12242 , \12244 );
xor \U$11903 ( \12246 , \11925 , \11927 );
xor \U$11904 ( \12247 , \12246 , \11930 );
and \U$11905 ( \12248 , \12244 , \12247 );
and \U$11906 ( \12249 , \12242 , \12247 );
or \U$11907 ( \12250 , \12245 , \12248 , \12249 );
and \U$11908 ( \12251 , \12240 , \12250 );
xor \U$11909 ( \12252 , \11594 , \11604 );
xor \U$11910 ( \12253 , \12252 , \11607 );
and \U$11911 ( \12254 , \12250 , \12253 );
and \U$11912 ( \12255 , \12240 , \12253 );
or \U$11913 ( \12256 , \12251 , \12254 , \12255 );
xor \U$11914 ( \12257 , \11515 , \11563 );
xor \U$11915 ( \12258 , \12257 , \11581 );
xor \U$11916 ( \12259 , \11904 , \11922 );
xor \U$11917 ( \12260 , \12259 , \11933 );
and \U$11918 ( \12261 , \12258 , \12260 );
xor \U$11919 ( \12262 , \11938 , \11940 );
xor \U$11920 ( \12263 , \12262 , \11943 );
and \U$11921 ( \12264 , \12260 , \12263 );
and \U$11922 ( \12265 , \12258 , \12263 );
or \U$11923 ( \12266 , \12261 , \12264 , \12265 );
and \U$11924 ( \12267 , \12256 , \12266 );
xor \U$11925 ( \12268 , \11626 , \11628 );
xor \U$11926 ( \12269 , \12268 , \11631 );
and \U$11927 ( \12270 , \12266 , \12269 );
and \U$11928 ( \12271 , \12256 , \12269 );
or \U$11929 ( \12272 , \12267 , \12270 , \12271 );
xor \U$11930 ( \12273 , \11584 , \11610 );
xor \U$11931 ( \12274 , \12273 , \11621 );
xor \U$11932 ( \12275 , \11936 , \11946 );
xor \U$11933 ( \12276 , \12275 , \11949 );
and \U$11934 ( \12277 , \12274 , \12276 );
and \U$11935 ( \12278 , \12272 , \12277 );
xor \U$11936 ( \12279 , \11952 , \11954 );
xor \U$11937 ( \12280 , \12279 , \11957 );
and \U$11938 ( \12281 , \12277 , \12280 );
and \U$11939 ( \12282 , \12272 , \12280 );
or \U$11940 ( \12283 , \12278 , \12281 , \12282 );
and \U$11941 ( \12284 , \11971 , \12283 );
xor \U$11942 ( \12285 , \11971 , \12283 );
xor \U$11943 ( \12286 , \12272 , \12277 );
xor \U$11944 ( \12287 , \12286 , \12280 );
xor \U$11945 ( \12288 , \12022 , \12026 );
xor \U$11946 ( \12289 , \12288 , \12031 );
xor \U$11947 ( \12290 , \12127 , \12131 );
xor \U$11948 ( \12291 , \12290 , \12136 );
and \U$11949 ( \12292 , \12289 , \12291 );
xor \U$11950 ( \12293 , \12160 , \12164 );
xor \U$11951 ( \12294 , \12293 , \12169 );
and \U$11952 ( \12295 , \12291 , \12294 );
and \U$11953 ( \12296 , \12289 , \12294 );
or \U$11954 ( \12297 , \12292 , \12295 , \12296 );
and \U$11955 ( \12298 , \9347 , \357 );
and \U$11956 ( \12299 , \8778 , \355 );
nor \U$11957 ( \12300 , \12298 , \12299 );
xnor \U$11958 ( \12301 , \12300 , \364 );
and \U$11959 ( \12302 , \9958 , \373 );
and \U$11960 ( \12303 , \9355 , \371 );
nor \U$11961 ( \12304 , \12302 , \12303 );
xnor \U$11962 ( \12305 , \12304 , \380 );
and \U$11963 ( \12306 , \12301 , \12305 );
and \U$11964 ( \12307 , \10144 , \391 );
and \U$11965 ( \12308 , \9963 , \389 );
nor \U$11966 ( \12309 , \12307 , \12308 );
xnor \U$11967 ( \12310 , \12309 , \398 );
and \U$11968 ( \12311 , \12305 , \12310 );
and \U$11969 ( \12312 , \12301 , \12310 );
or \U$11970 ( \12313 , \12306 , \12311 , \12312 );
xor \U$11971 ( \12314 , \12143 , \12147 );
xor \U$11972 ( \12315 , \12314 , \12152 );
and \U$11973 ( \12316 , \12313 , \12315 );
xor \U$11974 ( \12317 , \11996 , \12000 );
xor \U$11975 ( \12318 , \12317 , \12005 );
and \U$11976 ( \12319 , \12315 , \12318 );
and \U$11977 ( \12320 , \12313 , \12318 );
or \U$11978 ( \12321 , \12316 , \12319 , \12320 );
and \U$11979 ( \12322 , \12297 , \12321 );
xor \U$11980 ( \12323 , \12074 , \12078 );
xor \U$11981 ( \12324 , \12323 , \12083 );
xor \U$11982 ( \12325 , \12038 , \12042 );
xor \U$11983 ( \12326 , \12325 , \12047 );
and \U$11984 ( \12327 , \12324 , \12326 );
xor \U$11985 ( \12328 , \12055 , \12059 );
xor \U$11986 ( \12329 , \12328 , \12064 );
and \U$11987 ( \12330 , \12326 , \12329 );
and \U$11988 ( \12331 , \12324 , \12329 );
or \U$11989 ( \12332 , \12327 , \12330 , \12331 );
and \U$11990 ( \12333 , \12321 , \12332 );
and \U$11991 ( \12334 , \12297 , \12332 );
or \U$11992 ( \12335 , \12322 , \12333 , \12334 );
and \U$11993 ( \12336 , \983 , \7564 );
and \U$11994 ( \12337 , \785 , \7562 );
nor \U$11995 ( \12338 , \12336 , \12337 );
xnor \U$11996 ( \12339 , \12338 , \7315 );
and \U$11997 ( \12340 , \1176 , \7035 );
and \U$11998 ( \12341 , \1071 , \7033 );
nor \U$11999 ( \12342 , \12340 , \12341 );
xnor \U$12000 ( \12343 , \12342 , \6775 );
and \U$12001 ( \12344 , \12339 , \12343 );
and \U$12002 ( \12345 , \1297 , \6541 );
and \U$12003 ( \12346 , \1181 , \6539 );
nor \U$12004 ( \12347 , \12345 , \12346 );
xnor \U$12005 ( \12348 , \12347 , \6226 );
and \U$12006 ( \12349 , \12343 , \12348 );
and \U$12007 ( \12350 , \12339 , \12348 );
or \U$12008 ( \12351 , \12344 , \12349 , \12350 );
and \U$12009 ( \12352 , \408 , \10611 );
and \U$12010 ( \12353 , \385 , \10608 );
nor \U$12011 ( \12354 , \12352 , \12353 );
xnor \U$12012 ( \12355 , \12354 , \9556 );
and \U$12013 ( \12356 , \424 , \9798 );
and \U$12014 ( \12357 , \400 , \9796 );
nor \U$12015 ( \12358 , \12356 , \12357 );
xnor \U$12016 ( \12359 , \12358 , \9559 );
and \U$12017 ( \12360 , \12355 , \12359 );
and \U$12018 ( \12361 , \12359 , \413 );
and \U$12019 ( \12362 , \12355 , \413 );
or \U$12020 ( \12363 , \12360 , \12361 , \12362 );
and \U$12021 ( \12364 , \12351 , \12363 );
and \U$12022 ( \12365 , \443 , \9230 );
and \U$12023 ( \12366 , \416 , \9228 );
nor \U$12024 ( \12367 , \12365 , \12366 );
xnor \U$12025 ( \12368 , \12367 , \8920 );
and \U$12026 ( \12369 , \450 , \8693 );
and \U$12027 ( \12370 , \435 , \8691 );
nor \U$12028 ( \12371 , \12369 , \12370 );
xnor \U$12029 ( \12372 , \12371 , \8322 );
and \U$12030 ( \12373 , \12368 , \12372 );
and \U$12031 ( \12374 , \722 , \8131 );
and \U$12032 ( \12375 , \661 , \8129 );
nor \U$12033 ( \12376 , \12374 , \12375 );
xnor \U$12034 ( \12377 , \12376 , \7813 );
and \U$12035 ( \12378 , \12372 , \12377 );
and \U$12036 ( \12379 , \12368 , \12377 );
or \U$12037 ( \12380 , \12373 , \12378 , \12379 );
and \U$12038 ( \12381 , \12363 , \12380 );
and \U$12039 ( \12382 , \12351 , \12380 );
or \U$12040 ( \12383 , \12364 , \12381 , \12382 );
and \U$12041 ( \12384 , \3478 , \3434 );
and \U$12042 ( \12385 , \3061 , \3432 );
nor \U$12043 ( \12386 , \12384 , \12385 );
xnor \U$12044 ( \12387 , \12386 , \3247 );
and \U$12045 ( \12388 , \3808 , \3121 );
and \U$12046 ( \12389 , \3686 , \3119 );
nor \U$12047 ( \12390 , \12388 , \12389 );
xnor \U$12048 ( \12391 , \12390 , \2916 );
and \U$12049 ( \12392 , \12387 , \12391 );
and \U$12050 ( \12393 , \4069 , \2715 );
and \U$12051 ( \12394 , \3813 , \2713 );
nor \U$12052 ( \12395 , \12393 , \12394 );
xnor \U$12053 ( \12396 , \12395 , \2566 );
and \U$12054 ( \12397 , \12391 , \12396 );
and \U$12055 ( \12398 , \12387 , \12396 );
or \U$12056 ( \12399 , \12392 , \12397 , \12398 );
and \U$12057 ( \12400 , \2438 , \4603 );
and \U$12058 ( \12401 , \2174 , \4601 );
nor \U$12059 ( \12402 , \12400 , \12401 );
xnor \U$12060 ( \12403 , \12402 , \4371 );
and \U$12061 ( \12404 , \2637 , \4152 );
and \U$12062 ( \12405 , \2463 , \4150 );
nor \U$12063 ( \12406 , \12404 , \12405 );
xnor \U$12064 ( \12407 , \12406 , \4009 );
and \U$12065 ( \12408 , \12403 , \12407 );
and \U$12066 ( \12409 , \2942 , \3829 );
and \U$12067 ( \12410 , \2804 , \3827 );
nor \U$12068 ( \12411 , \12409 , \12410 );
xnor \U$12069 ( \12412 , \12411 , \3583 );
and \U$12070 ( \12413 , \12407 , \12412 );
and \U$12071 ( \12414 , \12403 , \12412 );
or \U$12072 ( \12415 , \12408 , \12413 , \12414 );
and \U$12073 ( \12416 , \12399 , \12415 );
and \U$12074 ( \12417 , \1588 , \6032 );
and \U$12075 ( \12418 , \1412 , \6030 );
nor \U$12076 ( \12419 , \12417 , \12418 );
xnor \U$12077 ( \12420 , \12419 , \5692 );
and \U$12078 ( \12421 , \1839 , \5443 );
and \U$12079 ( \12422 , \1596 , \5441 );
nor \U$12080 ( \12423 , \12421 , \12422 );
xnor \U$12081 ( \12424 , \12423 , \5202 );
and \U$12082 ( \12425 , \12420 , \12424 );
and \U$12083 ( \12426 , \2030 , \4977 );
and \U$12084 ( \12427 , \1844 , \4975 );
nor \U$12085 ( \12428 , \12426 , \12427 );
xnor \U$12086 ( \12429 , \12428 , \4789 );
and \U$12087 ( \12430 , \12424 , \12429 );
and \U$12088 ( \12431 , \12420 , \12429 );
or \U$12089 ( \12432 , \12425 , \12430 , \12431 );
and \U$12090 ( \12433 , \12415 , \12432 );
and \U$12091 ( \12434 , \12399 , \12432 );
or \U$12092 ( \12435 , \12416 , \12433 , \12434 );
and \U$12093 ( \12436 , \12383 , \12435 );
and \U$12094 ( \12437 , \4568 , \2393 );
and \U$12095 ( \12438 , \4266 , \2391 );
nor \U$12096 ( \12439 , \12437 , \12438 );
xnor \U$12097 ( \12440 , \12439 , \2251 );
and \U$12098 ( \12441 , \5045 , \2097 );
and \U$12099 ( \12442 , \4576 , \2095 );
nor \U$12100 ( \12443 , \12441 , \12442 );
xnor \U$12101 ( \12444 , \12443 , \1960 );
and \U$12102 ( \12445 , \12440 , \12444 );
and \U$12103 ( \12446 , \5314 , \1891 );
and \U$12104 ( \12447 , \5050 , \1889 );
nor \U$12105 ( \12448 , \12446 , \12447 );
xnor \U$12106 ( \12449 , \12448 , \1739 );
and \U$12107 ( \12450 , \12444 , \12449 );
and \U$12108 ( \12451 , \12440 , \12449 );
or \U$12109 ( \12452 , \12445 , \12450 , \12451 );
and \U$12110 ( \12453 , \5945 , \1623 );
and \U$12111 ( \12454 , \5573 , \1621 );
nor \U$12112 ( \12455 , \12453 , \12454 );
xnor \U$12113 ( \12456 , \12455 , \1467 );
and \U$12114 ( \12457 , \6297 , \1351 );
and \U$12115 ( \12458 , \5954 , \1349 );
nor \U$12116 ( \12459 , \12457 , \12458 );
xnor \U$12117 ( \12460 , \12459 , \1238 );
and \U$12118 ( \12461 , \12456 , \12460 );
and \U$12119 ( \12462 , \6802 , \1157 );
and \U$12120 ( \12463 , \6499 , \1155 );
nor \U$12121 ( \12464 , \12462 , \12463 );
xnor \U$12122 ( \12465 , \12464 , \1021 );
and \U$12123 ( \12466 , \12460 , \12465 );
and \U$12124 ( \12467 , \12456 , \12465 );
or \U$12125 ( \12468 , \12461 , \12466 , \12467 );
and \U$12126 ( \12469 , \12452 , \12468 );
and \U$12127 ( \12470 , \7500 , \957 );
and \U$12128 ( \12471 , \6974 , \955 );
nor \U$12129 ( \12472 , \12470 , \12471 );
xnor \U$12130 ( \12473 , \12472 , \879 );
and \U$12131 ( \12474 , \8170 , \793 );
and \U$12132 ( \12475 , \7924 , \791 );
nor \U$12133 ( \12476 , \12474 , \12475 );
xnor \U$12134 ( \12477 , \12476 , \699 );
and \U$12135 ( \12478 , \12473 , \12477 );
and \U$12136 ( \12479 , \8494 , \624 );
and \U$12137 ( \12480 , \8175 , \622 );
nor \U$12138 ( \12481 , \12479 , \12480 );
xnor \U$12139 ( \12482 , \12481 , \349 );
and \U$12140 ( \12483 , \12477 , \12482 );
and \U$12141 ( \12484 , \12473 , \12482 );
or \U$12142 ( \12485 , \12478 , \12483 , \12484 );
and \U$12143 ( \12486 , \12468 , \12485 );
and \U$12144 ( \12487 , \12452 , \12485 );
or \U$12145 ( \12488 , \12469 , \12486 , \12487 );
and \U$12146 ( \12489 , \12435 , \12488 );
and \U$12147 ( \12490 , \12383 , \12488 );
or \U$12148 ( \12491 , \12436 , \12489 , \12490 );
and \U$12149 ( \12492 , \12335 , \12491 );
xor \U$12150 ( \12493 , \12181 , \12183 );
xor \U$12151 ( \12494 , \12493 , \12186 );
xor \U$12152 ( \12495 , \11973 , \11975 );
xor \U$12153 ( \12496 , \12495 , \11978 );
and \U$12154 ( \12497 , \12494 , \12496 );
xor \U$12155 ( \12498 , \11983 , \11985 );
xor \U$12156 ( \12499 , \12498 , \11988 );
and \U$12157 ( \12500 , \12496 , \12499 );
and \U$12158 ( \12501 , \12494 , \12499 );
or \U$12159 ( \12502 , \12497 , \12500 , \12501 );
and \U$12160 ( \12503 , \12491 , \12502 );
and \U$12161 ( \12504 , \12335 , \12502 );
or \U$12162 ( \12505 , \12492 , \12503 , \12504 );
xor \U$12163 ( \12506 , \12034 , \12050 );
xor \U$12164 ( \12507 , \12506 , \12067 );
xor \U$12165 ( \12508 , \12139 , \12155 );
xor \U$12166 ( \12509 , \12508 , \12172 );
and \U$12167 ( \12510 , \12507 , \12509 );
xor \U$12168 ( \12511 , \12008 , \12010 );
xor \U$12169 ( \12512 , \12511 , \12012 );
and \U$12170 ( \12513 , \12509 , \12512 );
and \U$12171 ( \12514 , \12507 , \12512 );
or \U$12172 ( \12515 , \12510 , \12513 , \12514 );
xor \U$12173 ( \12516 , \12202 , \12204 );
xor \U$12174 ( \12517 , \12516 , \12207 );
and \U$12175 ( \12518 , \12515 , \12517 );
xor \U$12176 ( \12519 , \12212 , \12214 );
xor \U$12177 ( \12520 , \12519 , \12217 );
and \U$12178 ( \12521 , \12517 , \12520 );
and \U$12179 ( \12522 , \12515 , \12520 );
or \U$12180 ( \12523 , \12518 , \12521 , \12522 );
and \U$12181 ( \12524 , \12505 , \12523 );
xor \U$12182 ( \12525 , \11981 , \11991 );
xor \U$12183 ( \12526 , \12525 , \12015 );
xor \U$12184 ( \12527 , \12070 , \12122 );
xor \U$12185 ( \12528 , \12527 , \12175 );
and \U$12186 ( \12529 , \12526 , \12528 );
xor \U$12187 ( \12530 , \12189 , \12191 );
xor \U$12188 ( \12531 , \12530 , \12194 );
and \U$12189 ( \12532 , \12528 , \12531 );
and \U$12190 ( \12533 , \12526 , \12531 );
or \U$12191 ( \12534 , \12529 , \12532 , \12533 );
and \U$12192 ( \12535 , \12523 , \12534 );
and \U$12193 ( \12536 , \12505 , \12534 );
or \U$12194 ( \12537 , \12524 , \12535 , \12536 );
xor \U$12195 ( \12538 , \11723 , \11771 );
xor \U$12196 ( \12539 , \12538 , \11824 );
xor \U$12197 ( \12540 , \11858 , \11868 );
xor \U$12198 ( \12541 , \12540 , \11879 );
and \U$12199 ( \12542 , \12539 , \12541 );
xor \U$12200 ( \12543 , \12229 , \12231 );
xor \U$12201 ( \12544 , \12543 , \12234 );
and \U$12202 ( \12545 , \12541 , \12544 );
and \U$12203 ( \12546 , \12539 , \12544 );
or \U$12204 ( \12547 , \12542 , \12545 , \12546 );
and \U$12205 ( \12548 , \12537 , \12547 );
xor \U$12206 ( \12549 , \12242 , \12244 );
xor \U$12207 ( \12550 , \12549 , \12247 );
and \U$12208 ( \12551 , \12547 , \12550 );
and \U$12209 ( \12552 , \12537 , \12550 );
or \U$12210 ( \12553 , \12548 , \12551 , \12552 );
xor \U$12211 ( \12554 , \12240 , \12250 );
xor \U$12212 ( \12555 , \12554 , \12253 );
and \U$12213 ( \12556 , \12553 , \12555 );
xor \U$12214 ( \12557 , \12258 , \12260 );
xor \U$12215 ( \12558 , \12557 , \12263 );
and \U$12216 ( \12559 , \12555 , \12558 );
and \U$12217 ( \12560 , \12553 , \12558 );
or \U$12218 ( \12561 , \12556 , \12559 , \12560 );
xor \U$12219 ( \12562 , \12256 , \12266 );
xor \U$12220 ( \12563 , \12562 , \12269 );
and \U$12221 ( \12564 , \12561 , \12563 );
xor \U$12222 ( \12565 , \12274 , \12276 );
and \U$12223 ( \12566 , \12563 , \12565 );
and \U$12224 ( \12567 , \12561 , \12565 );
or \U$12225 ( \12568 , \12564 , \12566 , \12567 );
and \U$12226 ( \12569 , \12287 , \12568 );
xor \U$12227 ( \12570 , \12287 , \12568 );
xor \U$12228 ( \12571 , \12561 , \12563 );
xor \U$12229 ( \12572 , \12571 , \12565 );
and \U$12230 ( \12573 , \2804 , \4152 );
and \U$12231 ( \12574 , \2637 , \4150 );
nor \U$12232 ( \12575 , \12573 , \12574 );
xnor \U$12233 ( \12576 , \12575 , \4009 );
and \U$12234 ( \12577 , \3061 , \3829 );
and \U$12235 ( \12578 , \2942 , \3827 );
nor \U$12236 ( \12579 , \12577 , \12578 );
xnor \U$12237 ( \12580 , \12579 , \3583 );
and \U$12238 ( \12581 , \12576 , \12580 );
and \U$12239 ( \12582 , \3686 , \3434 );
and \U$12240 ( \12583 , \3478 , \3432 );
nor \U$12241 ( \12584 , \12582 , \12583 );
xnor \U$12242 ( \12585 , \12584 , \3247 );
and \U$12243 ( \12586 , \12580 , \12585 );
and \U$12244 ( \12587 , \12576 , \12585 );
or \U$12245 ( \12588 , \12581 , \12586 , \12587 );
and \U$12246 ( \12589 , \3813 , \3121 );
and \U$12247 ( \12590 , \3808 , \3119 );
nor \U$12248 ( \12591 , \12589 , \12590 );
xnor \U$12249 ( \12592 , \12591 , \2916 );
and \U$12250 ( \12593 , \4266 , \2715 );
and \U$12251 ( \12594 , \4069 , \2713 );
nor \U$12252 ( \12595 , \12593 , \12594 );
xnor \U$12253 ( \12596 , \12595 , \2566 );
and \U$12254 ( \12597 , \12592 , \12596 );
and \U$12255 ( \12598 , \4576 , \2393 );
and \U$12256 ( \12599 , \4568 , \2391 );
nor \U$12257 ( \12600 , \12598 , \12599 );
xnor \U$12258 ( \12601 , \12600 , \2251 );
and \U$12259 ( \12602 , \12596 , \12601 );
and \U$12260 ( \12603 , \12592 , \12601 );
or \U$12261 ( \12604 , \12597 , \12602 , \12603 );
and \U$12262 ( \12605 , \12588 , \12604 );
and \U$12263 ( \12606 , \1844 , \5443 );
and \U$12264 ( \12607 , \1839 , \5441 );
nor \U$12265 ( \12608 , \12606 , \12607 );
xnor \U$12266 ( \12609 , \12608 , \5202 );
and \U$12267 ( \12610 , \2174 , \4977 );
and \U$12268 ( \12611 , \2030 , \4975 );
nor \U$12269 ( \12612 , \12610 , \12611 );
xnor \U$12270 ( \12613 , \12612 , \4789 );
and \U$12271 ( \12614 , \12609 , \12613 );
and \U$12272 ( \12615 , \2463 , \4603 );
and \U$12273 ( \12616 , \2438 , \4601 );
nor \U$12274 ( \12617 , \12615 , \12616 );
xnor \U$12275 ( \12618 , \12617 , \4371 );
and \U$12276 ( \12619 , \12613 , \12618 );
and \U$12277 ( \12620 , \12609 , \12618 );
or \U$12278 ( \12621 , \12614 , \12619 , \12620 );
and \U$12279 ( \12622 , \12604 , \12621 );
and \U$12280 ( \12623 , \12588 , \12621 );
or \U$12281 ( \12624 , \12605 , \12622 , \12623 );
and \U$12282 ( \12625 , \6499 , \1351 );
and \U$12283 ( \12626 , \6297 , \1349 );
nor \U$12284 ( \12627 , \12625 , \12626 );
xnor \U$12285 ( \12628 , \12627 , \1238 );
and \U$12286 ( \12629 , \6974 , \1157 );
and \U$12287 ( \12630 , \6802 , \1155 );
nor \U$12288 ( \12631 , \12629 , \12630 );
xnor \U$12289 ( \12632 , \12631 , \1021 );
and \U$12290 ( \12633 , \12628 , \12632 );
and \U$12291 ( \12634 , \7924 , \957 );
and \U$12292 ( \12635 , \7500 , \955 );
nor \U$12293 ( \12636 , \12634 , \12635 );
xnor \U$12294 ( \12637 , \12636 , \879 );
and \U$12295 ( \12638 , \12632 , \12637 );
and \U$12296 ( \12639 , \12628 , \12637 );
or \U$12297 ( \12640 , \12633 , \12638 , \12639 );
and \U$12298 ( \12641 , \8175 , \793 );
and \U$12299 ( \12642 , \8170 , \791 );
nor \U$12300 ( \12643 , \12641 , \12642 );
xnor \U$12301 ( \12644 , \12643 , \699 );
and \U$12302 ( \12645 , \8778 , \624 );
and \U$12303 ( \12646 , \8494 , \622 );
nor \U$12304 ( \12647 , \12645 , \12646 );
xnor \U$12305 ( \12648 , \12647 , \349 );
and \U$12306 ( \12649 , \12644 , \12648 );
and \U$12307 ( \12650 , \9355 , \357 );
and \U$12308 ( \12651 , \9347 , \355 );
nor \U$12309 ( \12652 , \12650 , \12651 );
xnor \U$12310 ( \12653 , \12652 , \364 );
and \U$12311 ( \12654 , \12648 , \12653 );
and \U$12312 ( \12655 , \12644 , \12653 );
or \U$12313 ( \12656 , \12649 , \12654 , \12655 );
and \U$12314 ( \12657 , \12640 , \12656 );
and \U$12315 ( \12658 , \5050 , \2097 );
and \U$12316 ( \12659 , \5045 , \2095 );
nor \U$12317 ( \12660 , \12658 , \12659 );
xnor \U$12318 ( \12661 , \12660 , \1960 );
and \U$12319 ( \12662 , \5573 , \1891 );
and \U$12320 ( \12663 , \5314 , \1889 );
nor \U$12321 ( \12664 , \12662 , \12663 );
xnor \U$12322 ( \12665 , \12664 , \1739 );
and \U$12323 ( \12666 , \12661 , \12665 );
and \U$12324 ( \12667 , \5954 , \1623 );
and \U$12325 ( \12668 , \5945 , \1621 );
nor \U$12326 ( \12669 , \12667 , \12668 );
xnor \U$12327 ( \12670 , \12669 , \1467 );
and \U$12328 ( \12671 , \12665 , \12670 );
and \U$12329 ( \12672 , \12661 , \12670 );
or \U$12330 ( \12673 , \12666 , \12671 , \12672 );
and \U$12331 ( \12674 , \12656 , \12673 );
and \U$12332 ( \12675 , \12640 , \12673 );
or \U$12333 ( \12676 , \12657 , \12674 , \12675 );
and \U$12334 ( \12677 , \12624 , \12676 );
and \U$12335 ( \12678 , \400 , \10611 );
and \U$12336 ( \12679 , \408 , \10608 );
nor \U$12337 ( \12680 , \12678 , \12679 );
xnor \U$12338 ( \12681 , \12680 , \9556 );
and \U$12339 ( \12682 , \416 , \9798 );
and \U$12340 ( \12683 , \424 , \9796 );
nor \U$12341 ( \12684 , \12682 , \12683 );
xnor \U$12342 ( \12685 , \12684 , \9559 );
and \U$12343 ( \12686 , \12681 , \12685 );
and \U$12344 ( \12687 , \435 , \9230 );
and \U$12345 ( \12688 , \443 , \9228 );
nor \U$12346 ( \12689 , \12687 , \12688 );
xnor \U$12347 ( \12690 , \12689 , \8920 );
and \U$12348 ( \12691 , \12685 , \12690 );
and \U$12349 ( \12692 , \12681 , \12690 );
or \U$12350 ( \12693 , \12686 , \12691 , \12692 );
and \U$12351 ( \12694 , \661 , \8693 );
and \U$12352 ( \12695 , \450 , \8691 );
nor \U$12353 ( \12696 , \12694 , \12695 );
xnor \U$12354 ( \12697 , \12696 , \8322 );
and \U$12355 ( \12698 , \785 , \8131 );
and \U$12356 ( \12699 , \722 , \8129 );
nor \U$12357 ( \12700 , \12698 , \12699 );
xnor \U$12358 ( \12701 , \12700 , \7813 );
and \U$12359 ( \12702 , \12697 , \12701 );
and \U$12360 ( \12703 , \1071 , \7564 );
and \U$12361 ( \12704 , \983 , \7562 );
nor \U$12362 ( \12705 , \12703 , \12704 );
xnor \U$12363 ( \12706 , \12705 , \7315 );
and \U$12364 ( \12707 , \12701 , \12706 );
and \U$12365 ( \12708 , \12697 , \12706 );
or \U$12366 ( \12709 , \12702 , \12707 , \12708 );
and \U$12367 ( \12710 , \12693 , \12709 );
and \U$12368 ( \12711 , \1181 , \7035 );
and \U$12369 ( \12712 , \1176 , \7033 );
nor \U$12370 ( \12713 , \12711 , \12712 );
xnor \U$12371 ( \12714 , \12713 , \6775 );
and \U$12372 ( \12715 , \1412 , \6541 );
and \U$12373 ( \12716 , \1297 , \6539 );
nor \U$12374 ( \12717 , \12715 , \12716 );
xnor \U$12375 ( \12718 , \12717 , \6226 );
and \U$12376 ( \12719 , \12714 , \12718 );
and \U$12377 ( \12720 , \1596 , \6032 );
and \U$12378 ( \12721 , \1588 , \6030 );
nor \U$12379 ( \12722 , \12720 , \12721 );
xnor \U$12380 ( \12723 , \12722 , \5692 );
and \U$12381 ( \12724 , \12718 , \12723 );
and \U$12382 ( \12725 , \12714 , \12723 );
or \U$12383 ( \12726 , \12719 , \12724 , \12725 );
and \U$12384 ( \12727 , \12709 , \12726 );
and \U$12385 ( \12728 , \12693 , \12726 );
or \U$12386 ( \12729 , \12710 , \12727 , \12728 );
and \U$12387 ( \12730 , \12676 , \12729 );
and \U$12388 ( \12731 , \12624 , \12729 );
or \U$12389 ( \12732 , \12677 , \12730 , \12731 );
xor \U$12390 ( \12733 , \12339 , \12343 );
xor \U$12391 ( \12734 , \12733 , \12348 );
xor \U$12392 ( \12735 , \12403 , \12407 );
xor \U$12393 ( \12736 , \12735 , \12412 );
and \U$12394 ( \12737 , \12734 , \12736 );
xor \U$12395 ( \12738 , \12420 , \12424 );
xor \U$12396 ( \12739 , \12738 , \12429 );
and \U$12397 ( \12740 , \12736 , \12739 );
and \U$12398 ( \12741 , \12734 , \12739 );
or \U$12399 ( \12742 , \12737 , \12740 , \12741 );
xor \U$12400 ( \12743 , \12387 , \12391 );
xor \U$12401 ( \12744 , \12743 , \12396 );
xor \U$12402 ( \12745 , \12440 , \12444 );
xor \U$12403 ( \12746 , \12745 , \12449 );
and \U$12404 ( \12747 , \12744 , \12746 );
xor \U$12405 ( \12748 , \12456 , \12460 );
xor \U$12406 ( \12749 , \12748 , \12465 );
and \U$12407 ( \12750 , \12746 , \12749 );
and \U$12408 ( \12751 , \12744 , \12749 );
or \U$12409 ( \12752 , \12747 , \12750 , \12751 );
and \U$12410 ( \12753 , \12742 , \12752 );
nand \U$12411 ( \12754 , \10764 , \404 );
xnor \U$12412 ( \12755 , \12754 , \413 );
xor \U$12413 ( \12756 , \12473 , \12477 );
xor \U$12414 ( \12757 , \12756 , \12482 );
and \U$12415 ( \12758 , \12755 , \12757 );
xor \U$12416 ( \12759 , \12301 , \12305 );
xor \U$12417 ( \12760 , \12759 , \12310 );
and \U$12418 ( \12761 , \12757 , \12760 );
and \U$12419 ( \12762 , \12755 , \12760 );
or \U$12420 ( \12763 , \12758 , \12761 , \12762 );
and \U$12421 ( \12764 , \12752 , \12763 );
and \U$12422 ( \12765 , \12742 , \12763 );
or \U$12423 ( \12766 , \12753 , \12764 , \12765 );
and \U$12424 ( \12767 , \12732 , \12766 );
xor \U$12425 ( \12768 , \12090 , \12094 );
xor \U$12426 ( \12769 , \12768 , \12099 );
xor \U$12427 ( \12770 , \12107 , \12111 );
xor \U$12428 ( \12771 , \12770 , \12116 );
and \U$12429 ( \12772 , \12769 , \12771 );
xor \U$12430 ( \12773 , \12324 , \12326 );
xor \U$12431 ( \12774 , \12773 , \12329 );
and \U$12432 ( \12775 , \12771 , \12774 );
and \U$12433 ( \12776 , \12769 , \12774 );
or \U$12434 ( \12777 , \12772 , \12775 , \12776 );
and \U$12435 ( \12778 , \12766 , \12777 );
and \U$12436 ( \12779 , \12732 , \12777 );
or \U$12437 ( \12780 , \12767 , \12778 , \12779 );
xor \U$12438 ( \12781 , \12297 , \12321 );
xor \U$12439 ( \12782 , \12781 , \12332 );
xor \U$12440 ( \12783 , \12383 , \12435 );
xor \U$12441 ( \12784 , \12783 , \12488 );
and \U$12442 ( \12785 , \12782 , \12784 );
xor \U$12443 ( \12786 , \12494 , \12496 );
xor \U$12444 ( \12787 , \12786 , \12499 );
and \U$12445 ( \12788 , \12784 , \12787 );
and \U$12446 ( \12789 , \12782 , \12787 );
or \U$12447 ( \12790 , \12785 , \12788 , \12789 );
and \U$12448 ( \12791 , \12780 , \12790 );
xor \U$12449 ( \12792 , \12452 , \12468 );
xor \U$12450 ( \12793 , \12792 , \12485 );
xor \U$12451 ( \12794 , \12289 , \12291 );
xor \U$12452 ( \12795 , \12794 , \12294 );
and \U$12453 ( \12796 , \12793 , \12795 );
xor \U$12454 ( \12797 , \12313 , \12315 );
xor \U$12455 ( \12798 , \12797 , \12318 );
and \U$12456 ( \12799 , \12795 , \12798 );
and \U$12457 ( \12800 , \12793 , \12798 );
or \U$12458 ( \12801 , \12796 , \12799 , \12800 );
xor \U$12459 ( \12802 , \12086 , \12102 );
xor \U$12460 ( \12803 , \12802 , \12119 );
and \U$12461 ( \12804 , \12801 , \12803 );
xor \U$12462 ( \12805 , \12507 , \12509 );
xor \U$12463 ( \12806 , \12805 , \12512 );
and \U$12464 ( \12807 , \12803 , \12806 );
and \U$12465 ( \12808 , \12801 , \12806 );
or \U$12466 ( \12809 , \12804 , \12807 , \12808 );
and \U$12467 ( \12810 , \12790 , \12809 );
and \U$12468 ( \12811 , \12780 , \12809 );
or \U$12469 ( \12812 , \12791 , \12810 , \12811 );
xor \U$12470 ( \12813 , \12335 , \12491 );
xor \U$12471 ( \12814 , \12813 , \12502 );
xor \U$12472 ( \12815 , \12515 , \12517 );
xor \U$12473 ( \12816 , \12815 , \12520 );
and \U$12474 ( \12817 , \12814 , \12816 );
xor \U$12475 ( \12818 , \12526 , \12528 );
xor \U$12476 ( \12819 , \12818 , \12531 );
and \U$12477 ( \12820 , \12816 , \12819 );
and \U$12478 ( \12821 , \12814 , \12819 );
or \U$12479 ( \12822 , \12817 , \12820 , \12821 );
and \U$12480 ( \12823 , \12812 , \12822 );
xor \U$12481 ( \12824 , \12210 , \12220 );
xor \U$12482 ( \12825 , \12824 , \12223 );
and \U$12483 ( \12826 , \12822 , \12825 );
and \U$12484 ( \12827 , \12812 , \12825 );
or \U$12485 ( \12828 , \12823 , \12826 , \12827 );
xor \U$12486 ( \12829 , \12018 , \12178 );
xor \U$12487 ( \12830 , \12829 , \12197 );
xor \U$12488 ( \12831 , \12505 , \12523 );
xor \U$12489 ( \12832 , \12831 , \12534 );
and \U$12490 ( \12833 , \12830 , \12832 );
xor \U$12491 ( \12834 , \12539 , \12541 );
xor \U$12492 ( \12835 , \12834 , \12544 );
and \U$12493 ( \12836 , \12832 , \12835 );
and \U$12494 ( \12837 , \12830 , \12835 );
or \U$12495 ( \12838 , \12833 , \12836 , \12837 );
and \U$12496 ( \12839 , \12828 , \12838 );
xor \U$12497 ( \12840 , \12200 , \12226 );
xor \U$12498 ( \12841 , \12840 , \12237 );
and \U$12499 ( \12842 , \12838 , \12841 );
and \U$12500 ( \12843 , \12828 , \12841 );
or \U$12501 ( \12844 , \12839 , \12842 , \12843 );
xor \U$12502 ( \12845 , \12553 , \12555 );
xor \U$12503 ( \12846 , \12845 , \12558 );
and \U$12504 ( \12847 , \12844 , \12846 );
and \U$12505 ( \12848 , \12572 , \12847 );
xor \U$12506 ( \12849 , \12572 , \12847 );
xor \U$12507 ( \12850 , \12844 , \12846 );
and \U$12508 ( \12851 , \9958 , \357 );
and \U$12509 ( \12852 , \9355 , \355 );
nor \U$12510 ( \12853 , \12851 , \12852 );
xnor \U$12511 ( \12854 , \12853 , \364 );
and \U$12512 ( \12855 , \10144 , \373 );
and \U$12513 ( \12856 , \9963 , \371 );
nor \U$12514 ( \12857 , \12855 , \12856 );
xnor \U$12515 ( \12858 , \12857 , \380 );
and \U$12516 ( \12859 , \12854 , \12858 );
nand \U$12517 ( \12860 , \10764 , \389 );
xnor \U$12518 ( \12861 , \12860 , \398 );
and \U$12519 ( \12862 , \12858 , \12861 );
and \U$12520 ( \12863 , \12854 , \12861 );
or \U$12521 ( \12864 , \12859 , \12862 , \12863 );
and \U$12522 ( \12865 , \9963 , \373 );
and \U$12523 ( \12866 , \9958 , \371 );
nor \U$12524 ( \12867 , \12865 , \12866 );
xnor \U$12525 ( \12868 , \12867 , \380 );
and \U$12526 ( \12869 , \12864 , \12868 );
and \U$12527 ( \12870 , \10764 , \391 );
and \U$12528 ( \12871 , \10144 , \389 );
nor \U$12529 ( \12872 , \12870 , \12871 );
xnor \U$12530 ( \12873 , \12872 , \398 );
and \U$12531 ( \12874 , \12868 , \12873 );
and \U$12532 ( \12875 , \12864 , \12873 );
or \U$12533 ( \12876 , \12869 , \12874 , \12875 );
xor \U$12534 ( \12877 , \12628 , \12632 );
xor \U$12535 ( \12878 , \12877 , \12637 );
xor \U$12536 ( \12879 , \12644 , \12648 );
xor \U$12537 ( \12880 , \12879 , \12653 );
and \U$12538 ( \12881 , \12878 , \12880 );
xor \U$12539 ( \12882 , \12661 , \12665 );
xor \U$12540 ( \12883 , \12882 , \12670 );
and \U$12541 ( \12884 , \12880 , \12883 );
and \U$12542 ( \12885 , \12878 , \12883 );
or \U$12543 ( \12886 , \12881 , \12884 , \12885 );
and \U$12544 ( \12887 , \12876 , \12886 );
xor \U$12545 ( \12888 , \12576 , \12580 );
xor \U$12546 ( \12889 , \12888 , \12585 );
xor \U$12547 ( \12890 , \12592 , \12596 );
xor \U$12548 ( \12891 , \12890 , \12601 );
and \U$12549 ( \12892 , \12889 , \12891 );
xor \U$12550 ( \12893 , \12609 , \12613 );
xor \U$12551 ( \12894 , \12893 , \12618 );
and \U$12552 ( \12895 , \12891 , \12894 );
and \U$12553 ( \12896 , \12889 , \12894 );
or \U$12554 ( \12897 , \12892 , \12895 , \12896 );
and \U$12555 ( \12898 , \12886 , \12897 );
and \U$12556 ( \12899 , \12876 , \12897 );
or \U$12557 ( \12900 , \12887 , \12898 , \12899 );
and \U$12558 ( \12901 , \450 , \9230 );
and \U$12559 ( \12902 , \435 , \9228 );
nor \U$12560 ( \12903 , \12901 , \12902 );
xnor \U$12561 ( \12904 , \12903 , \8920 );
and \U$12562 ( \12905 , \722 , \8693 );
and \U$12563 ( \12906 , \661 , \8691 );
nor \U$12564 ( \12907 , \12905 , \12906 );
xnor \U$12565 ( \12908 , \12907 , \8322 );
and \U$12566 ( \12909 , \12904 , \12908 );
and \U$12567 ( \12910 , \983 , \8131 );
and \U$12568 ( \12911 , \785 , \8129 );
nor \U$12569 ( \12912 , \12910 , \12911 );
xnor \U$12570 ( \12913 , \12912 , \7813 );
and \U$12571 ( \12914 , \12908 , \12913 );
and \U$12572 ( \12915 , \12904 , \12913 );
or \U$12573 ( \12916 , \12909 , \12914 , \12915 );
and \U$12574 ( \12917 , \1176 , \7564 );
and \U$12575 ( \12918 , \1071 , \7562 );
nor \U$12576 ( \12919 , \12917 , \12918 );
xnor \U$12577 ( \12920 , \12919 , \7315 );
and \U$12578 ( \12921 , \1297 , \7035 );
and \U$12579 ( \12922 , \1181 , \7033 );
nor \U$12580 ( \12923 , \12921 , \12922 );
xnor \U$12581 ( \12924 , \12923 , \6775 );
and \U$12582 ( \12925 , \12920 , \12924 );
and \U$12583 ( \12926 , \1588 , \6541 );
and \U$12584 ( \12927 , \1412 , \6539 );
nor \U$12585 ( \12928 , \12926 , \12927 );
xnor \U$12586 ( \12929 , \12928 , \6226 );
and \U$12587 ( \12930 , \12924 , \12929 );
and \U$12588 ( \12931 , \12920 , \12929 );
or \U$12589 ( \12932 , \12925 , \12930 , \12931 );
and \U$12590 ( \12933 , \12916 , \12932 );
and \U$12591 ( \12934 , \424 , \10611 );
and \U$12592 ( \12935 , \400 , \10608 );
nor \U$12593 ( \12936 , \12934 , \12935 );
xnor \U$12594 ( \12937 , \12936 , \9556 );
and \U$12595 ( \12938 , \443 , \9798 );
and \U$12596 ( \12939 , \416 , \9796 );
nor \U$12597 ( \12940 , \12938 , \12939 );
xnor \U$12598 ( \12941 , \12940 , \9559 );
and \U$12599 ( \12942 , \12937 , \12941 );
and \U$12600 ( \12943 , \12941 , \398 );
and \U$12601 ( \12944 , \12937 , \398 );
or \U$12602 ( \12945 , \12942 , \12943 , \12944 );
and \U$12603 ( \12946 , \12932 , \12945 );
and \U$12604 ( \12947 , \12916 , \12945 );
or \U$12605 ( \12948 , \12933 , \12946 , \12947 );
and \U$12606 ( \12949 , \3808 , \3434 );
and \U$12607 ( \12950 , \3686 , \3432 );
nor \U$12608 ( \12951 , \12949 , \12950 );
xnor \U$12609 ( \12952 , \12951 , \3247 );
and \U$12610 ( \12953 , \4069 , \3121 );
and \U$12611 ( \12954 , \3813 , \3119 );
nor \U$12612 ( \12955 , \12953 , \12954 );
xnor \U$12613 ( \12956 , \12955 , \2916 );
and \U$12614 ( \12957 , \12952 , \12956 );
and \U$12615 ( \12958 , \4568 , \2715 );
and \U$12616 ( \12959 , \4266 , \2713 );
nor \U$12617 ( \12960 , \12958 , \12959 );
xnor \U$12618 ( \12961 , \12960 , \2566 );
and \U$12619 ( \12962 , \12956 , \12961 );
and \U$12620 ( \12963 , \12952 , \12961 );
or \U$12621 ( \12964 , \12957 , \12962 , \12963 );
and \U$12622 ( \12965 , \1839 , \6032 );
and \U$12623 ( \12966 , \1596 , \6030 );
nor \U$12624 ( \12967 , \12965 , \12966 );
xnor \U$12625 ( \12968 , \12967 , \5692 );
and \U$12626 ( \12969 , \2030 , \5443 );
and \U$12627 ( \12970 , \1844 , \5441 );
nor \U$12628 ( \12971 , \12969 , \12970 );
xnor \U$12629 ( \12972 , \12971 , \5202 );
and \U$12630 ( \12973 , \12968 , \12972 );
and \U$12631 ( \12974 , \2438 , \4977 );
and \U$12632 ( \12975 , \2174 , \4975 );
nor \U$12633 ( \12976 , \12974 , \12975 );
xnor \U$12634 ( \12977 , \12976 , \4789 );
and \U$12635 ( \12978 , \12972 , \12977 );
and \U$12636 ( \12979 , \12968 , \12977 );
or \U$12637 ( \12980 , \12973 , \12978 , \12979 );
and \U$12638 ( \12981 , \12964 , \12980 );
and \U$12639 ( \12982 , \2637 , \4603 );
and \U$12640 ( \12983 , \2463 , \4601 );
nor \U$12641 ( \12984 , \12982 , \12983 );
xnor \U$12642 ( \12985 , \12984 , \4371 );
and \U$12643 ( \12986 , \2942 , \4152 );
and \U$12644 ( \12987 , \2804 , \4150 );
nor \U$12645 ( \12988 , \12986 , \12987 );
xnor \U$12646 ( \12989 , \12988 , \4009 );
and \U$12647 ( \12990 , \12985 , \12989 );
and \U$12648 ( \12991 , \3478 , \3829 );
and \U$12649 ( \12992 , \3061 , \3827 );
nor \U$12650 ( \12993 , \12991 , \12992 );
xnor \U$12651 ( \12994 , \12993 , \3583 );
and \U$12652 ( \12995 , \12989 , \12994 );
and \U$12653 ( \12996 , \12985 , \12994 );
or \U$12654 ( \12997 , \12990 , \12995 , \12996 );
and \U$12655 ( \12998 , \12980 , \12997 );
and \U$12656 ( \12999 , \12964 , \12997 );
or \U$12657 ( \13000 , \12981 , \12998 , \12999 );
and \U$12658 ( \13001 , \12948 , \13000 );
and \U$12659 ( \13002 , \6297 , \1623 );
and \U$12660 ( \13003 , \5954 , \1621 );
nor \U$12661 ( \13004 , \13002 , \13003 );
xnor \U$12662 ( \13005 , \13004 , \1467 );
and \U$12663 ( \13006 , \6802 , \1351 );
and \U$12664 ( \13007 , \6499 , \1349 );
nor \U$12665 ( \13008 , \13006 , \13007 );
xnor \U$12666 ( \13009 , \13008 , \1238 );
and \U$12667 ( \13010 , \13005 , \13009 );
and \U$12668 ( \13011 , \7500 , \1157 );
and \U$12669 ( \13012 , \6974 , \1155 );
nor \U$12670 ( \13013 , \13011 , \13012 );
xnor \U$12671 ( \13014 , \13013 , \1021 );
and \U$12672 ( \13015 , \13009 , \13014 );
and \U$12673 ( \13016 , \13005 , \13014 );
or \U$12674 ( \13017 , \13010 , \13015 , \13016 );
and \U$12675 ( \13018 , \8170 , \957 );
and \U$12676 ( \13019 , \7924 , \955 );
nor \U$12677 ( \13020 , \13018 , \13019 );
xnor \U$12678 ( \13021 , \13020 , \879 );
and \U$12679 ( \13022 , \8494 , \793 );
and \U$12680 ( \13023 , \8175 , \791 );
nor \U$12681 ( \13024 , \13022 , \13023 );
xnor \U$12682 ( \13025 , \13024 , \699 );
and \U$12683 ( \13026 , \13021 , \13025 );
and \U$12684 ( \13027 , \9347 , \624 );
and \U$12685 ( \13028 , \8778 , \622 );
nor \U$12686 ( \13029 , \13027 , \13028 );
xnor \U$12687 ( \13030 , \13029 , \349 );
and \U$12688 ( \13031 , \13025 , \13030 );
and \U$12689 ( \13032 , \13021 , \13030 );
or \U$12690 ( \13033 , \13026 , \13031 , \13032 );
and \U$12691 ( \13034 , \13017 , \13033 );
and \U$12692 ( \13035 , \5045 , \2393 );
and \U$12693 ( \13036 , \4576 , \2391 );
nor \U$12694 ( \13037 , \13035 , \13036 );
xnor \U$12695 ( \13038 , \13037 , \2251 );
and \U$12696 ( \13039 , \5314 , \2097 );
and \U$12697 ( \13040 , \5050 , \2095 );
nor \U$12698 ( \13041 , \13039 , \13040 );
xnor \U$12699 ( \13042 , \13041 , \1960 );
and \U$12700 ( \13043 , \13038 , \13042 );
and \U$12701 ( \13044 , \5945 , \1891 );
and \U$12702 ( \13045 , \5573 , \1889 );
nor \U$12703 ( \13046 , \13044 , \13045 );
xnor \U$12704 ( \13047 , \13046 , \1739 );
and \U$12705 ( \13048 , \13042 , \13047 );
and \U$12706 ( \13049 , \13038 , \13047 );
or \U$12707 ( \13050 , \13043 , \13048 , \13049 );
and \U$12708 ( \13051 , \13033 , \13050 );
and \U$12709 ( \13052 , \13017 , \13050 );
or \U$12710 ( \13053 , \13034 , \13051 , \13052 );
and \U$12711 ( \13054 , \13000 , \13053 );
and \U$12712 ( \13055 , \12948 , \13053 );
or \U$12713 ( \13056 , \13001 , \13054 , \13055 );
and \U$12714 ( \13057 , \12900 , \13056 );
xor \U$12715 ( \13058 , \12681 , \12685 );
xor \U$12716 ( \13059 , \13058 , \12690 );
xor \U$12717 ( \13060 , \12697 , \12701 );
xor \U$12718 ( \13061 , \13060 , \12706 );
and \U$12719 ( \13062 , \13059 , \13061 );
xor \U$12720 ( \13063 , \12714 , \12718 );
xor \U$12721 ( \13064 , \13063 , \12723 );
and \U$12722 ( \13065 , \13061 , \13064 );
and \U$12723 ( \13066 , \13059 , \13064 );
or \U$12724 ( \13067 , \13062 , \13065 , \13066 );
xor \U$12725 ( \13068 , \12355 , \12359 );
xor \U$12726 ( \13069 , \13068 , \413 );
and \U$12727 ( \13070 , \13067 , \13069 );
xor \U$12728 ( \13071 , \12368 , \12372 );
xor \U$12729 ( \13072 , \13071 , \12377 );
and \U$12730 ( \13073 , \13069 , \13072 );
and \U$12731 ( \13074 , \13067 , \13072 );
or \U$12732 ( \13075 , \13070 , \13073 , \13074 );
and \U$12733 ( \13076 , \13056 , \13075 );
and \U$12734 ( \13077 , \12900 , \13075 );
or \U$12735 ( \13078 , \13057 , \13076 , \13077 );
xor \U$12736 ( \13079 , \12588 , \12604 );
xor \U$12737 ( \13080 , \13079 , \12621 );
xor \U$12738 ( \13081 , \12640 , \12656 );
xor \U$12739 ( \13082 , \13081 , \12673 );
and \U$12740 ( \13083 , \13080 , \13082 );
xor \U$12741 ( \13084 , \12693 , \12709 );
xor \U$12742 ( \13085 , \13084 , \12726 );
and \U$12743 ( \13086 , \13082 , \13085 );
and \U$12744 ( \13087 , \13080 , \13085 );
or \U$12745 ( \13088 , \13083 , \13086 , \13087 );
xor \U$12746 ( \13089 , \12734 , \12736 );
xor \U$12747 ( \13090 , \13089 , \12739 );
xor \U$12748 ( \13091 , \12744 , \12746 );
xor \U$12749 ( \13092 , \13091 , \12749 );
and \U$12750 ( \13093 , \13090 , \13092 );
xor \U$12751 ( \13094 , \12755 , \12757 );
xor \U$12752 ( \13095 , \13094 , \12760 );
and \U$12753 ( \13096 , \13092 , \13095 );
and \U$12754 ( \13097 , \13090 , \13095 );
or \U$12755 ( \13098 , \13093 , \13096 , \13097 );
and \U$12756 ( \13099 , \13088 , \13098 );
xor \U$12757 ( \13100 , \12399 , \12415 );
xor \U$12758 ( \13101 , \13100 , \12432 );
and \U$12759 ( \13102 , \13098 , \13101 );
and \U$12760 ( \13103 , \13088 , \13101 );
or \U$12761 ( \13104 , \13099 , \13102 , \13103 );
and \U$12762 ( \13105 , \13078 , \13104 );
xor \U$12763 ( \13106 , \12351 , \12363 );
xor \U$12764 ( \13107 , \13106 , \12380 );
xor \U$12765 ( \13108 , \12769 , \12771 );
xor \U$12766 ( \13109 , \13108 , \12774 );
and \U$12767 ( \13110 , \13107 , \13109 );
xor \U$12768 ( \13111 , \12793 , \12795 );
xor \U$12769 ( \13112 , \13111 , \12798 );
and \U$12770 ( \13113 , \13109 , \13112 );
and \U$12771 ( \13114 , \13107 , \13112 );
or \U$12772 ( \13115 , \13110 , \13113 , \13114 );
and \U$12773 ( \13116 , \13104 , \13115 );
and \U$12774 ( \13117 , \13078 , \13115 );
or \U$12775 ( \13118 , \13105 , \13116 , \13117 );
xor \U$12776 ( \13119 , \12732 , \12766 );
xor \U$12777 ( \13120 , \13119 , \12777 );
xor \U$12778 ( \13121 , \12782 , \12784 );
xor \U$12779 ( \13122 , \13121 , \12787 );
and \U$12780 ( \13123 , \13120 , \13122 );
xor \U$12781 ( \13124 , \12801 , \12803 );
xor \U$12782 ( \13125 , \13124 , \12806 );
and \U$12783 ( \13126 , \13122 , \13125 );
and \U$12784 ( \13127 , \13120 , \13125 );
or \U$12785 ( \13128 , \13123 , \13126 , \13127 );
and \U$12786 ( \13129 , \13118 , \13128 );
xor \U$12787 ( \13130 , \12814 , \12816 );
xor \U$12788 ( \13131 , \13130 , \12819 );
and \U$12789 ( \13132 , \13128 , \13131 );
and \U$12790 ( \13133 , \13118 , \13131 );
or \U$12791 ( \13134 , \13129 , \13132 , \13133 );
xor \U$12792 ( \13135 , \12812 , \12822 );
xor \U$12793 ( \13136 , \13135 , \12825 );
and \U$12794 ( \13137 , \13134 , \13136 );
xor \U$12795 ( \13138 , \12830 , \12832 );
xor \U$12796 ( \13139 , \13138 , \12835 );
and \U$12797 ( \13140 , \13136 , \13139 );
and \U$12798 ( \13141 , \13134 , \13139 );
or \U$12799 ( \13142 , \13137 , \13140 , \13141 );
xor \U$12800 ( \13143 , \12828 , \12838 );
xor \U$12801 ( \13144 , \13143 , \12841 );
and \U$12802 ( \13145 , \13142 , \13144 );
xor \U$12803 ( \13146 , \12537 , \12547 );
xor \U$12804 ( \13147 , \13146 , \12550 );
and \U$12805 ( \13148 , \13144 , \13147 );
and \U$12806 ( \13149 , \13142 , \13147 );
or \U$12807 ( \13150 , \13145 , \13148 , \13149 );
and \U$12808 ( \13151 , \12850 , \13150 );
xor \U$12809 ( \13152 , \12850 , \13150 );
xor \U$12810 ( \13153 , \13142 , \13144 );
xor \U$12811 ( \13154 , \13153 , \13147 );
xor \U$12812 ( \13155 , \12904 , \12908 );
xor \U$12813 ( \13156 , \13155 , \12913 );
xor \U$12814 ( \13157 , \12920 , \12924 );
xor \U$12815 ( \13158 , \13157 , \12929 );
and \U$12816 ( \13159 , \13156 , \13158 );
xor \U$12817 ( \13160 , \12968 , \12972 );
xor \U$12818 ( \13161 , \13160 , \12977 );
and \U$12819 ( \13162 , \13158 , \13161 );
and \U$12820 ( \13163 , \13156 , \13161 );
or \U$12821 ( \13164 , \13159 , \13162 , \13163 );
xor \U$12822 ( \13165 , \12952 , \12956 );
xor \U$12823 ( \13166 , \13165 , \12961 );
xor \U$12824 ( \13167 , \12985 , \12989 );
xor \U$12825 ( \13168 , \13167 , \12994 );
and \U$12826 ( \13169 , \13166 , \13168 );
xor \U$12827 ( \13170 , \13038 , \13042 );
xor \U$12828 ( \13171 , \13170 , \13047 );
and \U$12829 ( \13172 , \13168 , \13171 );
and \U$12830 ( \13173 , \13166 , \13171 );
or \U$12831 ( \13174 , \13169 , \13172 , \13173 );
and \U$12832 ( \13175 , \13164 , \13174 );
xor \U$12833 ( \13176 , \13005 , \13009 );
xor \U$12834 ( \13177 , \13176 , \13014 );
xor \U$12835 ( \13178 , \12854 , \12858 );
xor \U$12836 ( \13179 , \13178 , \12861 );
and \U$12837 ( \13180 , \13177 , \13179 );
xor \U$12838 ( \13181 , \13021 , \13025 );
xor \U$12839 ( \13182 , \13181 , \13030 );
and \U$12840 ( \13183 , \13179 , \13182 );
and \U$12841 ( \13184 , \13177 , \13182 );
or \U$12842 ( \13185 , \13180 , \13183 , \13184 );
and \U$12843 ( \13186 , \13174 , \13185 );
and \U$12844 ( \13187 , \13164 , \13185 );
or \U$12845 ( \13188 , \13175 , \13186 , \13187 );
and \U$12846 ( \13189 , \2174 , \5443 );
and \U$12847 ( \13190 , \2030 , \5441 );
nor \U$12848 ( \13191 , \13189 , \13190 );
xnor \U$12849 ( \13192 , \13191 , \5202 );
and \U$12850 ( \13193 , \2463 , \4977 );
and \U$12851 ( \13194 , \2438 , \4975 );
nor \U$12852 ( \13195 , \13193 , \13194 );
xnor \U$12853 ( \13196 , \13195 , \4789 );
and \U$12854 ( \13197 , \13192 , \13196 );
and \U$12855 ( \13198 , \2804 , \4603 );
and \U$12856 ( \13199 , \2637 , \4601 );
nor \U$12857 ( \13200 , \13198 , \13199 );
xnor \U$12858 ( \13201 , \13200 , \4371 );
and \U$12859 ( \13202 , \13196 , \13201 );
and \U$12860 ( \13203 , \13192 , \13201 );
or \U$12861 ( \13204 , \13197 , \13202 , \13203 );
and \U$12862 ( \13205 , \4266 , \3121 );
and \U$12863 ( \13206 , \4069 , \3119 );
nor \U$12864 ( \13207 , \13205 , \13206 );
xnor \U$12865 ( \13208 , \13207 , \2916 );
and \U$12866 ( \13209 , \4576 , \2715 );
and \U$12867 ( \13210 , \4568 , \2713 );
nor \U$12868 ( \13211 , \13209 , \13210 );
xnor \U$12869 ( \13212 , \13211 , \2566 );
and \U$12870 ( \13213 , \13208 , \13212 );
and \U$12871 ( \13214 , \5050 , \2393 );
and \U$12872 ( \13215 , \5045 , \2391 );
nor \U$12873 ( \13216 , \13214 , \13215 );
xnor \U$12874 ( \13217 , \13216 , \2251 );
and \U$12875 ( \13218 , \13212 , \13217 );
and \U$12876 ( \13219 , \13208 , \13217 );
or \U$12877 ( \13220 , \13213 , \13218 , \13219 );
and \U$12878 ( \13221 , \13204 , \13220 );
and \U$12879 ( \13222 , \3061 , \4152 );
and \U$12880 ( \13223 , \2942 , \4150 );
nor \U$12881 ( \13224 , \13222 , \13223 );
xnor \U$12882 ( \13225 , \13224 , \4009 );
and \U$12883 ( \13226 , \3686 , \3829 );
and \U$12884 ( \13227 , \3478 , \3827 );
nor \U$12885 ( \13228 , \13226 , \13227 );
xnor \U$12886 ( \13229 , \13228 , \3583 );
and \U$12887 ( \13230 , \13225 , \13229 );
and \U$12888 ( \13231 , \3813 , \3434 );
and \U$12889 ( \13232 , \3808 , \3432 );
nor \U$12890 ( \13233 , \13231 , \13232 );
xnor \U$12891 ( \13234 , \13233 , \3247 );
and \U$12892 ( \13235 , \13229 , \13234 );
and \U$12893 ( \13236 , \13225 , \13234 );
or \U$12894 ( \13237 , \13230 , \13235 , \13236 );
and \U$12895 ( \13238 , \13220 , \13237 );
and \U$12896 ( \13239 , \13204 , \13237 );
or \U$12897 ( \13240 , \13221 , \13238 , \13239 );
and \U$12898 ( \13241 , \8778 , \793 );
and \U$12899 ( \13242 , \8494 , \791 );
nor \U$12900 ( \13243 , \13241 , \13242 );
xnor \U$12901 ( \13244 , \13243 , \699 );
and \U$12902 ( \13245 , \9355 , \624 );
and \U$12903 ( \13246 , \9347 , \622 );
nor \U$12904 ( \13247 , \13245 , \13246 );
xnor \U$12905 ( \13248 , \13247 , \349 );
and \U$12906 ( \13249 , \13244 , \13248 );
and \U$12907 ( \13250 , \9963 , \357 );
and \U$12908 ( \13251 , \9958 , \355 );
nor \U$12909 ( \13252 , \13250 , \13251 );
xnor \U$12910 ( \13253 , \13252 , \364 );
and \U$12911 ( \13254 , \13248 , \13253 );
and \U$12912 ( \13255 , \13244 , \13253 );
or \U$12913 ( \13256 , \13249 , \13254 , \13255 );
and \U$12914 ( \13257 , \6974 , \1351 );
and \U$12915 ( \13258 , \6802 , \1349 );
nor \U$12916 ( \13259 , \13257 , \13258 );
xnor \U$12917 ( \13260 , \13259 , \1238 );
and \U$12918 ( \13261 , \7924 , \1157 );
and \U$12919 ( \13262 , \7500 , \1155 );
nor \U$12920 ( \13263 , \13261 , \13262 );
xnor \U$12921 ( \13264 , \13263 , \1021 );
and \U$12922 ( \13265 , \13260 , \13264 );
and \U$12923 ( \13266 , \8175 , \957 );
and \U$12924 ( \13267 , \8170 , \955 );
nor \U$12925 ( \13268 , \13266 , \13267 );
xnor \U$12926 ( \13269 , \13268 , \879 );
and \U$12927 ( \13270 , \13264 , \13269 );
and \U$12928 ( \13271 , \13260 , \13269 );
or \U$12929 ( \13272 , \13265 , \13270 , \13271 );
and \U$12930 ( \13273 , \13256 , \13272 );
and \U$12931 ( \13274 , \5573 , \2097 );
and \U$12932 ( \13275 , \5314 , \2095 );
nor \U$12933 ( \13276 , \13274 , \13275 );
xnor \U$12934 ( \13277 , \13276 , \1960 );
and \U$12935 ( \13278 , \5954 , \1891 );
and \U$12936 ( \13279 , \5945 , \1889 );
nor \U$12937 ( \13280 , \13278 , \13279 );
xnor \U$12938 ( \13281 , \13280 , \1739 );
and \U$12939 ( \13282 , \13277 , \13281 );
and \U$12940 ( \13283 , \6499 , \1623 );
and \U$12941 ( \13284 , \6297 , \1621 );
nor \U$12942 ( \13285 , \13283 , \13284 );
xnor \U$12943 ( \13286 , \13285 , \1467 );
and \U$12944 ( \13287 , \13281 , \13286 );
and \U$12945 ( \13288 , \13277 , \13286 );
or \U$12946 ( \13289 , \13282 , \13287 , \13288 );
and \U$12947 ( \13290 , \13272 , \13289 );
and \U$12948 ( \13291 , \13256 , \13289 );
or \U$12949 ( \13292 , \13273 , \13290 , \13291 );
and \U$12950 ( \13293 , \13240 , \13292 );
and \U$12951 ( \13294 , \1412 , \7035 );
and \U$12952 ( \13295 , \1297 , \7033 );
nor \U$12953 ( \13296 , \13294 , \13295 );
xnor \U$12954 ( \13297 , \13296 , \6775 );
and \U$12955 ( \13298 , \1596 , \6541 );
and \U$12956 ( \13299 , \1588 , \6539 );
nor \U$12957 ( \13300 , \13298 , \13299 );
xnor \U$12958 ( \13301 , \13300 , \6226 );
and \U$12959 ( \13302 , \13297 , \13301 );
and \U$12960 ( \13303 , \1844 , \6032 );
and \U$12961 ( \13304 , \1839 , \6030 );
nor \U$12962 ( \13305 , \13303 , \13304 );
xnor \U$12963 ( \13306 , \13305 , \5692 );
and \U$12964 ( \13307 , \13301 , \13306 );
and \U$12965 ( \13308 , \13297 , \13306 );
or \U$12966 ( \13309 , \13302 , \13307 , \13308 );
and \U$12967 ( \13310 , \416 , \10611 );
and \U$12968 ( \13311 , \424 , \10608 );
nor \U$12969 ( \13312 , \13310 , \13311 );
xnor \U$12970 ( \13313 , \13312 , \9556 );
and \U$12971 ( \13314 , \435 , \9798 );
and \U$12972 ( \13315 , \443 , \9796 );
nor \U$12973 ( \13316 , \13314 , \13315 );
xnor \U$12974 ( \13317 , \13316 , \9559 );
and \U$12975 ( \13318 , \13313 , \13317 );
and \U$12976 ( \13319 , \661 , \9230 );
and \U$12977 ( \13320 , \450 , \9228 );
nor \U$12978 ( \13321 , \13319 , \13320 );
xnor \U$12979 ( \13322 , \13321 , \8920 );
and \U$12980 ( \13323 , \13317 , \13322 );
and \U$12981 ( \13324 , \13313 , \13322 );
or \U$12982 ( \13325 , \13318 , \13323 , \13324 );
and \U$12983 ( \13326 , \13309 , \13325 );
and \U$12984 ( \13327 , \785 , \8693 );
and \U$12985 ( \13328 , \722 , \8691 );
nor \U$12986 ( \13329 , \13327 , \13328 );
xnor \U$12987 ( \13330 , \13329 , \8322 );
and \U$12988 ( \13331 , \1071 , \8131 );
and \U$12989 ( \13332 , \983 , \8129 );
nor \U$12990 ( \13333 , \13331 , \13332 );
xnor \U$12991 ( \13334 , \13333 , \7813 );
and \U$12992 ( \13335 , \13330 , \13334 );
and \U$12993 ( \13336 , \1181 , \7564 );
and \U$12994 ( \13337 , \1176 , \7562 );
nor \U$12995 ( \13338 , \13336 , \13337 );
xnor \U$12996 ( \13339 , \13338 , \7315 );
and \U$12997 ( \13340 , \13334 , \13339 );
and \U$12998 ( \13341 , \13330 , \13339 );
or \U$12999 ( \13342 , \13335 , \13340 , \13341 );
and \U$13000 ( \13343 , \13325 , \13342 );
and \U$13001 ( \13344 , \13309 , \13342 );
or \U$13002 ( \13345 , \13326 , \13343 , \13344 );
and \U$13003 ( \13346 , \13292 , \13345 );
and \U$13004 ( \13347 , \13240 , \13345 );
or \U$13005 ( \13348 , \13293 , \13346 , \13347 );
and \U$13006 ( \13349 , \13188 , \13348 );
xor \U$13007 ( \13350 , \12878 , \12880 );
xor \U$13008 ( \13351 , \13350 , \12883 );
xor \U$13009 ( \13352 , \13059 , \13061 );
xor \U$13010 ( \13353 , \13352 , \13064 );
and \U$13011 ( \13354 , \13351 , \13353 );
xor \U$13012 ( \13355 , \12889 , \12891 );
xor \U$13013 ( \13356 , \13355 , \12894 );
and \U$13014 ( \13357 , \13353 , \13356 );
and \U$13015 ( \13358 , \13351 , \13356 );
or \U$13016 ( \13359 , \13354 , \13357 , \13358 );
and \U$13017 ( \13360 , \13348 , \13359 );
and \U$13018 ( \13361 , \13188 , \13359 );
or \U$13019 ( \13362 , \13349 , \13360 , \13361 );
xor \U$13020 ( \13363 , \12876 , \12886 );
xor \U$13021 ( \13364 , \13363 , \12897 );
xor \U$13022 ( \13365 , \12948 , \13000 );
xor \U$13023 ( \13366 , \13365 , \13053 );
and \U$13024 ( \13367 , \13364 , \13366 );
xor \U$13025 ( \13368 , \13067 , \13069 );
xor \U$13026 ( \13369 , \13368 , \13072 );
and \U$13027 ( \13370 , \13366 , \13369 );
and \U$13028 ( \13371 , \13364 , \13369 );
or \U$13029 ( \13372 , \13367 , \13370 , \13371 );
and \U$13030 ( \13373 , \13362 , \13372 );
xor \U$13031 ( \13374 , \12864 , \12868 );
xor \U$13032 ( \13375 , \13374 , \12873 );
xor \U$13033 ( \13376 , \12964 , \12980 );
xor \U$13034 ( \13377 , \13376 , \12997 );
and \U$13035 ( \13378 , \13375 , \13377 );
xor \U$13036 ( \13379 , \13017 , \13033 );
xor \U$13037 ( \13380 , \13379 , \13050 );
and \U$13038 ( \13381 , \13377 , \13380 );
and \U$13039 ( \13382 , \13375 , \13380 );
or \U$13040 ( \13383 , \13378 , \13381 , \13382 );
xor \U$13041 ( \13384 , \13080 , \13082 );
xor \U$13042 ( \13385 , \13384 , \13085 );
and \U$13043 ( \13386 , \13383 , \13385 );
xor \U$13044 ( \13387 , \13090 , \13092 );
xor \U$13045 ( \13388 , \13387 , \13095 );
and \U$13046 ( \13389 , \13385 , \13388 );
and \U$13047 ( \13390 , \13383 , \13388 );
or \U$13048 ( \13391 , \13386 , \13389 , \13390 );
and \U$13049 ( \13392 , \13372 , \13391 );
and \U$13050 ( \13393 , \13362 , \13391 );
or \U$13051 ( \13394 , \13373 , \13392 , \13393 );
xor \U$13052 ( \13395 , \12624 , \12676 );
xor \U$13053 ( \13396 , \13395 , \12729 );
xor \U$13054 ( \13397 , \12742 , \12752 );
xor \U$13055 ( \13398 , \13397 , \12763 );
and \U$13056 ( \13399 , \13396 , \13398 );
xor \U$13057 ( \13400 , \13107 , \13109 );
xor \U$13058 ( \13401 , \13400 , \13112 );
and \U$13059 ( \13402 , \13398 , \13401 );
and \U$13060 ( \13403 , \13396 , \13401 );
or \U$13061 ( \13404 , \13399 , \13402 , \13403 );
and \U$13062 ( \13405 , \13394 , \13404 );
xor \U$13063 ( \13406 , \13120 , \13122 );
xor \U$13064 ( \13407 , \13406 , \13125 );
and \U$13065 ( \13408 , \13404 , \13407 );
and \U$13066 ( \13409 , \13394 , \13407 );
or \U$13067 ( \13410 , \13405 , \13408 , \13409 );
xor \U$13068 ( \13411 , \12780 , \12790 );
xor \U$13069 ( \13412 , \13411 , \12809 );
and \U$13070 ( \13413 , \13410 , \13412 );
xor \U$13071 ( \13414 , \13118 , \13128 );
xor \U$13072 ( \13415 , \13414 , \13131 );
and \U$13073 ( \13416 , \13412 , \13415 );
and \U$13074 ( \13417 , \13410 , \13415 );
or \U$13075 ( \13418 , \13413 , \13416 , \13417 );
xor \U$13076 ( \13419 , \13134 , \13136 );
xor \U$13077 ( \13420 , \13419 , \13139 );
and \U$13078 ( \13421 , \13418 , \13420 );
and \U$13079 ( \13422 , \13154 , \13421 );
xor \U$13080 ( \13423 , \13154 , \13421 );
xor \U$13081 ( \13424 , \13418 , \13420 );
xor \U$13082 ( \13425 , \13208 , \13212 );
xor \U$13083 ( \13426 , \13425 , \13217 );
xor \U$13084 ( \13427 , \13225 , \13229 );
xor \U$13085 ( \13428 , \13427 , \13234 );
and \U$13086 ( \13429 , \13426 , \13428 );
xor \U$13087 ( \13430 , \13277 , \13281 );
xor \U$13088 ( \13431 , \13430 , \13286 );
and \U$13089 ( \13432 , \13428 , \13431 );
and \U$13090 ( \13433 , \13426 , \13431 );
or \U$13091 ( \13434 , \13429 , \13432 , \13433 );
xor \U$13092 ( \13435 , \13192 , \13196 );
xor \U$13093 ( \13436 , \13435 , \13201 );
xor \U$13094 ( \13437 , \13297 , \13301 );
xor \U$13095 ( \13438 , \13437 , \13306 );
and \U$13096 ( \13439 , \13436 , \13438 );
xor \U$13097 ( \13440 , \13330 , \13334 );
xor \U$13098 ( \13441 , \13440 , \13339 );
and \U$13099 ( \13442 , \13438 , \13441 );
and \U$13100 ( \13443 , \13436 , \13441 );
or \U$13101 ( \13444 , \13439 , \13442 , \13443 );
and \U$13102 ( \13445 , \13434 , \13444 );
and \U$13103 ( \13446 , \10764 , \373 );
and \U$13104 ( \13447 , \10144 , \371 );
nor \U$13105 ( \13448 , \13446 , \13447 );
xnor \U$13106 ( \13449 , \13448 , \380 );
xor \U$13107 ( \13450 , \13244 , \13248 );
xor \U$13108 ( \13451 , \13450 , \13253 );
and \U$13109 ( \13452 , \13449 , \13451 );
xor \U$13110 ( \13453 , \13260 , \13264 );
xor \U$13111 ( \13454 , \13453 , \13269 );
and \U$13112 ( \13455 , \13451 , \13454 );
and \U$13113 ( \13456 , \13449 , \13454 );
or \U$13114 ( \13457 , \13452 , \13455 , \13456 );
and \U$13115 ( \13458 , \13444 , \13457 );
and \U$13116 ( \13459 , \13434 , \13457 );
or \U$13117 ( \13460 , \13445 , \13458 , \13459 );
and \U$13118 ( \13461 , \1297 , \7564 );
and \U$13119 ( \13462 , \1181 , \7562 );
nor \U$13120 ( \13463 , \13461 , \13462 );
xnor \U$13121 ( \13464 , \13463 , \7315 );
and \U$13122 ( \13465 , \1588 , \7035 );
and \U$13123 ( \13466 , \1412 , \7033 );
nor \U$13124 ( \13467 , \13465 , \13466 );
xnor \U$13125 ( \13468 , \13467 , \6775 );
and \U$13126 ( \13469 , \13464 , \13468 );
and \U$13127 ( \13470 , \1839 , \6541 );
and \U$13128 ( \13471 , \1596 , \6539 );
nor \U$13129 ( \13472 , \13470 , \13471 );
xnor \U$13130 ( \13473 , \13472 , \6226 );
and \U$13131 ( \13474 , \13468 , \13473 );
and \U$13132 ( \13475 , \13464 , \13473 );
or \U$13133 ( \13476 , \13469 , \13474 , \13475 );
and \U$13134 ( \13477 , \722 , \9230 );
and \U$13135 ( \13478 , \661 , \9228 );
nor \U$13136 ( \13479 , \13477 , \13478 );
xnor \U$13137 ( \13480 , \13479 , \8920 );
and \U$13138 ( \13481 , \983 , \8693 );
and \U$13139 ( \13482 , \785 , \8691 );
nor \U$13140 ( \13483 , \13481 , \13482 );
xnor \U$13141 ( \13484 , \13483 , \8322 );
and \U$13142 ( \13485 , \13480 , \13484 );
and \U$13143 ( \13486 , \1176 , \8131 );
and \U$13144 ( \13487 , \1071 , \8129 );
nor \U$13145 ( \13488 , \13486 , \13487 );
xnor \U$13146 ( \13489 , \13488 , \7813 );
and \U$13147 ( \13490 , \13484 , \13489 );
and \U$13148 ( \13491 , \13480 , \13489 );
or \U$13149 ( \13492 , \13485 , \13490 , \13491 );
and \U$13150 ( \13493 , \13476 , \13492 );
and \U$13151 ( \13494 , \443 , \10611 );
and \U$13152 ( \13495 , \416 , \10608 );
nor \U$13153 ( \13496 , \13494 , \13495 );
xnor \U$13154 ( \13497 , \13496 , \9556 );
and \U$13155 ( \13498 , \450 , \9798 );
and \U$13156 ( \13499 , \435 , \9796 );
nor \U$13157 ( \13500 , \13498 , \13499 );
xnor \U$13158 ( \13501 , \13500 , \9559 );
and \U$13159 ( \13502 , \13497 , \13501 );
and \U$13160 ( \13503 , \13501 , \380 );
and \U$13161 ( \13504 , \13497 , \380 );
or \U$13162 ( \13505 , \13502 , \13503 , \13504 );
and \U$13163 ( \13506 , \13492 , \13505 );
and \U$13164 ( \13507 , \13476 , \13505 );
or \U$13165 ( \13508 , \13493 , \13506 , \13507 );
and \U$13166 ( \13509 , \8494 , \957 );
and \U$13167 ( \13510 , \8175 , \955 );
nor \U$13168 ( \13511 , \13509 , \13510 );
xnor \U$13169 ( \13512 , \13511 , \879 );
and \U$13170 ( \13513 , \9347 , \793 );
and \U$13171 ( \13514 , \8778 , \791 );
nor \U$13172 ( \13515 , \13513 , \13514 );
xnor \U$13173 ( \13516 , \13515 , \699 );
and \U$13174 ( \13517 , \13512 , \13516 );
and \U$13175 ( \13518 , \9958 , \624 );
and \U$13176 ( \13519 , \9355 , \622 );
nor \U$13177 ( \13520 , \13518 , \13519 );
xnor \U$13178 ( \13521 , \13520 , \349 );
and \U$13179 ( \13522 , \13516 , \13521 );
and \U$13180 ( \13523 , \13512 , \13521 );
or \U$13181 ( \13524 , \13517 , \13522 , \13523 );
and \U$13182 ( \13525 , \5314 , \2393 );
and \U$13183 ( \13526 , \5050 , \2391 );
nor \U$13184 ( \13527 , \13525 , \13526 );
xnor \U$13185 ( \13528 , \13527 , \2251 );
and \U$13186 ( \13529 , \5945 , \2097 );
and \U$13187 ( \13530 , \5573 , \2095 );
nor \U$13188 ( \13531 , \13529 , \13530 );
xnor \U$13189 ( \13532 , \13531 , \1960 );
and \U$13190 ( \13533 , \13528 , \13532 );
and \U$13191 ( \13534 , \6297 , \1891 );
and \U$13192 ( \13535 , \5954 , \1889 );
nor \U$13193 ( \13536 , \13534 , \13535 );
xnor \U$13194 ( \13537 , \13536 , \1739 );
and \U$13195 ( \13538 , \13532 , \13537 );
and \U$13196 ( \13539 , \13528 , \13537 );
or \U$13197 ( \13540 , \13533 , \13538 , \13539 );
and \U$13198 ( \13541 , \13524 , \13540 );
and \U$13199 ( \13542 , \6802 , \1623 );
and \U$13200 ( \13543 , \6499 , \1621 );
nor \U$13201 ( \13544 , \13542 , \13543 );
xnor \U$13202 ( \13545 , \13544 , \1467 );
and \U$13203 ( \13546 , \7500 , \1351 );
and \U$13204 ( \13547 , \6974 , \1349 );
nor \U$13205 ( \13548 , \13546 , \13547 );
xnor \U$13206 ( \13549 , \13548 , \1238 );
and \U$13207 ( \13550 , \13545 , \13549 );
and \U$13208 ( \13551 , \8170 , \1157 );
and \U$13209 ( \13552 , \7924 , \1155 );
nor \U$13210 ( \13553 , \13551 , \13552 );
xnor \U$13211 ( \13554 , \13553 , \1021 );
and \U$13212 ( \13555 , \13549 , \13554 );
and \U$13213 ( \13556 , \13545 , \13554 );
or \U$13214 ( \13557 , \13550 , \13555 , \13556 );
and \U$13215 ( \13558 , \13540 , \13557 );
and \U$13216 ( \13559 , \13524 , \13557 );
or \U$13217 ( \13560 , \13541 , \13558 , \13559 );
and \U$13218 ( \13561 , \13508 , \13560 );
and \U$13219 ( \13562 , \4069 , \3434 );
and \U$13220 ( \13563 , \3813 , \3432 );
nor \U$13221 ( \13564 , \13562 , \13563 );
xnor \U$13222 ( \13565 , \13564 , \3247 );
and \U$13223 ( \13566 , \4568 , \3121 );
and \U$13224 ( \13567 , \4266 , \3119 );
nor \U$13225 ( \13568 , \13566 , \13567 );
xnor \U$13226 ( \13569 , \13568 , \2916 );
and \U$13227 ( \13570 , \13565 , \13569 );
and \U$13228 ( \13571 , \5045 , \2715 );
and \U$13229 ( \13572 , \4576 , \2713 );
nor \U$13230 ( \13573 , \13571 , \13572 );
xnor \U$13231 ( \13574 , \13573 , \2566 );
and \U$13232 ( \13575 , \13569 , \13574 );
and \U$13233 ( \13576 , \13565 , \13574 );
or \U$13234 ( \13577 , \13570 , \13575 , \13576 );
and \U$13235 ( \13578 , \2942 , \4603 );
and \U$13236 ( \13579 , \2804 , \4601 );
nor \U$13237 ( \13580 , \13578 , \13579 );
xnor \U$13238 ( \13581 , \13580 , \4371 );
and \U$13239 ( \13582 , \3478 , \4152 );
and \U$13240 ( \13583 , \3061 , \4150 );
nor \U$13241 ( \13584 , \13582 , \13583 );
xnor \U$13242 ( \13585 , \13584 , \4009 );
and \U$13243 ( \13586 , \13581 , \13585 );
and \U$13244 ( \13587 , \3808 , \3829 );
and \U$13245 ( \13588 , \3686 , \3827 );
nor \U$13246 ( \13589 , \13587 , \13588 );
xnor \U$13247 ( \13590 , \13589 , \3583 );
and \U$13248 ( \13591 , \13585 , \13590 );
and \U$13249 ( \13592 , \13581 , \13590 );
or \U$13250 ( \13593 , \13586 , \13591 , \13592 );
and \U$13251 ( \13594 , \13577 , \13593 );
and \U$13252 ( \13595 , \2030 , \6032 );
and \U$13253 ( \13596 , \1844 , \6030 );
nor \U$13254 ( \13597 , \13595 , \13596 );
xnor \U$13255 ( \13598 , \13597 , \5692 );
and \U$13256 ( \13599 , \2438 , \5443 );
and \U$13257 ( \13600 , \2174 , \5441 );
nor \U$13258 ( \13601 , \13599 , \13600 );
xnor \U$13259 ( \13602 , \13601 , \5202 );
and \U$13260 ( \13603 , \13598 , \13602 );
and \U$13261 ( \13604 , \2637 , \4977 );
and \U$13262 ( \13605 , \2463 , \4975 );
nor \U$13263 ( \13606 , \13604 , \13605 );
xnor \U$13264 ( \13607 , \13606 , \4789 );
and \U$13265 ( \13608 , \13602 , \13607 );
and \U$13266 ( \13609 , \13598 , \13607 );
or \U$13267 ( \13610 , \13603 , \13608 , \13609 );
and \U$13268 ( \13611 , \13593 , \13610 );
and \U$13269 ( \13612 , \13577 , \13610 );
or \U$13270 ( \13613 , \13594 , \13611 , \13612 );
and \U$13271 ( \13614 , \13560 , \13613 );
and \U$13272 ( \13615 , \13508 , \13613 );
or \U$13273 ( \13616 , \13561 , \13614 , \13615 );
and \U$13274 ( \13617 , \13460 , \13616 );
xor \U$13275 ( \13618 , \12937 , \12941 );
xor \U$13276 ( \13619 , \13618 , \398 );
xor \U$13277 ( \13620 , \13156 , \13158 );
xor \U$13278 ( \13621 , \13620 , \13161 );
and \U$13279 ( \13622 , \13619 , \13621 );
xor \U$13280 ( \13623 , \13166 , \13168 );
xor \U$13281 ( \13624 , \13623 , \13171 );
and \U$13282 ( \13625 , \13621 , \13624 );
and \U$13283 ( \13626 , \13619 , \13624 );
or \U$13284 ( \13627 , \13622 , \13625 , \13626 );
and \U$13285 ( \13628 , \13616 , \13627 );
and \U$13286 ( \13629 , \13460 , \13627 );
or \U$13287 ( \13630 , \13617 , \13628 , \13629 );
xor \U$13288 ( \13631 , \13204 , \13220 );
xor \U$13289 ( \13632 , \13631 , \13237 );
xor \U$13290 ( \13633 , \13256 , \13272 );
xor \U$13291 ( \13634 , \13633 , \13289 );
and \U$13292 ( \13635 , \13632 , \13634 );
xor \U$13293 ( \13636 , \13177 , \13179 );
xor \U$13294 ( \13637 , \13636 , \13182 );
and \U$13295 ( \13638 , \13634 , \13637 );
and \U$13296 ( \13639 , \13632 , \13637 );
or \U$13297 ( \13640 , \13635 , \13638 , \13639 );
xor \U$13298 ( \13641 , \12916 , \12932 );
xor \U$13299 ( \13642 , \13641 , \12945 );
and \U$13300 ( \13643 , \13640 , \13642 );
xor \U$13301 ( \13644 , \13375 , \13377 );
xor \U$13302 ( \13645 , \13644 , \13380 );
and \U$13303 ( \13646 , \13642 , \13645 );
and \U$13304 ( \13647 , \13640 , \13645 );
or \U$13305 ( \13648 , \13643 , \13646 , \13647 );
and \U$13306 ( \13649 , \13630 , \13648 );
xor \U$13307 ( \13650 , \13164 , \13174 );
xor \U$13308 ( \13651 , \13650 , \13185 );
xor \U$13309 ( \13652 , \13240 , \13292 );
xor \U$13310 ( \13653 , \13652 , \13345 );
and \U$13311 ( \13654 , \13651 , \13653 );
xor \U$13312 ( \13655 , \13351 , \13353 );
xor \U$13313 ( \13656 , \13655 , \13356 );
and \U$13314 ( \13657 , \13653 , \13656 );
and \U$13315 ( \13658 , \13651 , \13656 );
or \U$13316 ( \13659 , \13654 , \13657 , \13658 );
and \U$13317 ( \13660 , \13648 , \13659 );
and \U$13318 ( \13661 , \13630 , \13659 );
or \U$13319 ( \13662 , \13649 , \13660 , \13661 );
xor \U$13320 ( \13663 , \13188 , \13348 );
xor \U$13321 ( \13664 , \13663 , \13359 );
xor \U$13322 ( \13665 , \13364 , \13366 );
xor \U$13323 ( \13666 , \13665 , \13369 );
and \U$13324 ( \13667 , \13664 , \13666 );
xor \U$13325 ( \13668 , \13383 , \13385 );
xor \U$13326 ( \13669 , \13668 , \13388 );
and \U$13327 ( \13670 , \13666 , \13669 );
and \U$13328 ( \13671 , \13664 , \13669 );
or \U$13329 ( \13672 , \13667 , \13670 , \13671 );
and \U$13330 ( \13673 , \13662 , \13672 );
xor \U$13331 ( \13674 , \13088 , \13098 );
xor \U$13332 ( \13675 , \13674 , \13101 );
and \U$13333 ( \13676 , \13672 , \13675 );
and \U$13334 ( \13677 , \13662 , \13675 );
or \U$13335 ( \13678 , \13673 , \13676 , \13677 );
xor \U$13336 ( \13679 , \12900 , \13056 );
xor \U$13337 ( \13680 , \13679 , \13075 );
xor \U$13338 ( \13681 , \13362 , \13372 );
xor \U$13339 ( \13682 , \13681 , \13391 );
and \U$13340 ( \13683 , \13680 , \13682 );
xor \U$13341 ( \13684 , \13396 , \13398 );
xor \U$13342 ( \13685 , \13684 , \13401 );
and \U$13343 ( \13686 , \13682 , \13685 );
and \U$13344 ( \13687 , \13680 , \13685 );
or \U$13345 ( \13688 , \13683 , \13686 , \13687 );
and \U$13346 ( \13689 , \13678 , \13688 );
xor \U$13347 ( \13690 , \13078 , \13104 );
xor \U$13348 ( \13691 , \13690 , \13115 );
and \U$13349 ( \13692 , \13688 , \13691 );
and \U$13350 ( \13693 , \13678 , \13691 );
or \U$13351 ( \13694 , \13689 , \13692 , \13693 );
xor \U$13352 ( \13695 , \13410 , \13412 );
xor \U$13353 ( \13696 , \13695 , \13415 );
and \U$13354 ( \13697 , \13694 , \13696 );
and \U$13355 ( \13698 , \13424 , \13697 );
xor \U$13356 ( \13699 , \13424 , \13697 );
xor \U$13357 ( \13700 , \13694 , \13696 );
xor \U$13358 ( \13701 , \13565 , \13569 );
xor \U$13359 ( \13702 , \13701 , \13574 );
xor \U$13360 ( \13703 , \13528 , \13532 );
xor \U$13361 ( \13704 , \13703 , \13537 );
and \U$13362 ( \13705 , \13702 , \13704 );
xor \U$13363 ( \13706 , \13545 , \13549 );
xor \U$13364 ( \13707 , \13706 , \13554 );
and \U$13365 ( \13708 , \13704 , \13707 );
and \U$13366 ( \13709 , \13702 , \13707 );
or \U$13367 ( \13710 , \13705 , \13708 , \13709 );
and \U$13368 ( \13711 , \10144 , \357 );
and \U$13369 ( \13712 , \9963 , \355 );
nor \U$13370 ( \13713 , \13711 , \13712 );
xnor \U$13371 ( \13714 , \13713 , \364 );
nand \U$13372 ( \13715 , \10764 , \371 );
xnor \U$13373 ( \13716 , \13715 , \380 );
and \U$13374 ( \13717 , \13714 , \13716 );
xor \U$13375 ( \13718 , \13512 , \13516 );
xor \U$13376 ( \13719 , \13718 , \13521 );
and \U$13377 ( \13720 , \13716 , \13719 );
and \U$13378 ( \13721 , \13714 , \13719 );
or \U$13379 ( \13722 , \13717 , \13720 , \13721 );
and \U$13380 ( \13723 , \13710 , \13722 );
xor \U$13381 ( \13724 , \13464 , \13468 );
xor \U$13382 ( \13725 , \13724 , \13473 );
xor \U$13383 ( \13726 , \13581 , \13585 );
xor \U$13384 ( \13727 , \13726 , \13590 );
and \U$13385 ( \13728 , \13725 , \13727 );
xor \U$13386 ( \13729 , \13598 , \13602 );
xor \U$13387 ( \13730 , \13729 , \13607 );
and \U$13388 ( \13731 , \13727 , \13730 );
and \U$13389 ( \13732 , \13725 , \13730 );
or \U$13390 ( \13733 , \13728 , \13731 , \13732 );
and \U$13391 ( \13734 , \13722 , \13733 );
and \U$13392 ( \13735 , \13710 , \13733 );
or \U$13393 ( \13736 , \13723 , \13734 , \13735 );
and \U$13394 ( \13737 , \9355 , \793 );
and \U$13395 ( \13738 , \9347 , \791 );
nor \U$13396 ( \13739 , \13737 , \13738 );
xnor \U$13397 ( \13740 , \13739 , \699 );
and \U$13398 ( \13741 , \9963 , \624 );
and \U$13399 ( \13742 , \9958 , \622 );
nor \U$13400 ( \13743 , \13741 , \13742 );
xnor \U$13401 ( \13744 , \13743 , \349 );
and \U$13402 ( \13745 , \13740 , \13744 );
and \U$13403 ( \13746 , \10764 , \357 );
and \U$13404 ( \13747 , \10144 , \355 );
nor \U$13405 ( \13748 , \13746 , \13747 );
xnor \U$13406 ( \13749 , \13748 , \364 );
and \U$13407 ( \13750 , \13744 , \13749 );
and \U$13408 ( \13751 , \13740 , \13749 );
or \U$13409 ( \13752 , \13745 , \13750 , \13751 );
and \U$13410 ( \13753 , \5954 , \2097 );
and \U$13411 ( \13754 , \5945 , \2095 );
nor \U$13412 ( \13755 , \13753 , \13754 );
xnor \U$13413 ( \13756 , \13755 , \1960 );
and \U$13414 ( \13757 , \6499 , \1891 );
and \U$13415 ( \13758 , \6297 , \1889 );
nor \U$13416 ( \13759 , \13757 , \13758 );
xnor \U$13417 ( \13760 , \13759 , \1739 );
and \U$13418 ( \13761 , \13756 , \13760 );
and \U$13419 ( \13762 , \6974 , \1623 );
and \U$13420 ( \13763 , \6802 , \1621 );
nor \U$13421 ( \13764 , \13762 , \13763 );
xnor \U$13422 ( \13765 , \13764 , \1467 );
and \U$13423 ( \13766 , \13760 , \13765 );
and \U$13424 ( \13767 , \13756 , \13765 );
or \U$13425 ( \13768 , \13761 , \13766 , \13767 );
and \U$13426 ( \13769 , \13752 , \13768 );
and \U$13427 ( \13770 , \7924 , \1351 );
and \U$13428 ( \13771 , \7500 , \1349 );
nor \U$13429 ( \13772 , \13770 , \13771 );
xnor \U$13430 ( \13773 , \13772 , \1238 );
and \U$13431 ( \13774 , \8175 , \1157 );
and \U$13432 ( \13775 , \8170 , \1155 );
nor \U$13433 ( \13776 , \13774 , \13775 );
xnor \U$13434 ( \13777 , \13776 , \1021 );
and \U$13435 ( \13778 , \13773 , \13777 );
and \U$13436 ( \13779 , \8778 , \957 );
and \U$13437 ( \13780 , \8494 , \955 );
nor \U$13438 ( \13781 , \13779 , \13780 );
xnor \U$13439 ( \13782 , \13781 , \879 );
and \U$13440 ( \13783 , \13777 , \13782 );
and \U$13441 ( \13784 , \13773 , \13782 );
or \U$13442 ( \13785 , \13778 , \13783 , \13784 );
and \U$13443 ( \13786 , \13768 , \13785 );
and \U$13444 ( \13787 , \13752 , \13785 );
or \U$13445 ( \13788 , \13769 , \13786 , \13787 );
and \U$13446 ( \13789 , \1071 , \8693 );
and \U$13447 ( \13790 , \983 , \8691 );
nor \U$13448 ( \13791 , \13789 , \13790 );
xnor \U$13449 ( \13792 , \13791 , \8322 );
and \U$13450 ( \13793 , \1181 , \8131 );
and \U$13451 ( \13794 , \1176 , \8129 );
nor \U$13452 ( \13795 , \13793 , \13794 );
xnor \U$13453 ( \13796 , \13795 , \7813 );
and \U$13454 ( \13797 , \13792 , \13796 );
and \U$13455 ( \13798 , \1412 , \7564 );
and \U$13456 ( \13799 , \1297 , \7562 );
nor \U$13457 ( \13800 , \13798 , \13799 );
xnor \U$13458 ( \13801 , \13800 , \7315 );
and \U$13459 ( \13802 , \13796 , \13801 );
and \U$13460 ( \13803 , \13792 , \13801 );
or \U$13461 ( \13804 , \13797 , \13802 , \13803 );
and \U$13462 ( \13805 , \1596 , \7035 );
and \U$13463 ( \13806 , \1588 , \7033 );
nor \U$13464 ( \13807 , \13805 , \13806 );
xnor \U$13465 ( \13808 , \13807 , \6775 );
and \U$13466 ( \13809 , \1844 , \6541 );
and \U$13467 ( \13810 , \1839 , \6539 );
nor \U$13468 ( \13811 , \13809 , \13810 );
xnor \U$13469 ( \13812 , \13811 , \6226 );
and \U$13470 ( \13813 , \13808 , \13812 );
and \U$13471 ( \13814 , \2174 , \6032 );
and \U$13472 ( \13815 , \2030 , \6030 );
nor \U$13473 ( \13816 , \13814 , \13815 );
xnor \U$13474 ( \13817 , \13816 , \5692 );
and \U$13475 ( \13818 , \13812 , \13817 );
and \U$13476 ( \13819 , \13808 , \13817 );
or \U$13477 ( \13820 , \13813 , \13818 , \13819 );
and \U$13478 ( \13821 , \13804 , \13820 );
and \U$13479 ( \13822 , \435 , \10611 );
and \U$13480 ( \13823 , \443 , \10608 );
nor \U$13481 ( \13824 , \13822 , \13823 );
xnor \U$13482 ( \13825 , \13824 , \9556 );
and \U$13483 ( \13826 , \661 , \9798 );
and \U$13484 ( \13827 , \450 , \9796 );
nor \U$13485 ( \13828 , \13826 , \13827 );
xnor \U$13486 ( \13829 , \13828 , \9559 );
and \U$13487 ( \13830 , \13825 , \13829 );
and \U$13488 ( \13831 , \785 , \9230 );
and \U$13489 ( \13832 , \722 , \9228 );
nor \U$13490 ( \13833 , \13831 , \13832 );
xnor \U$13491 ( \13834 , \13833 , \8920 );
and \U$13492 ( \13835 , \13829 , \13834 );
and \U$13493 ( \13836 , \13825 , \13834 );
or \U$13494 ( \13837 , \13830 , \13835 , \13836 );
and \U$13495 ( \13838 , \13820 , \13837 );
and \U$13496 ( \13839 , \13804 , \13837 );
or \U$13497 ( \13840 , \13821 , \13838 , \13839 );
and \U$13498 ( \13841 , \13788 , \13840 );
and \U$13499 ( \13842 , \4576 , \3121 );
and \U$13500 ( \13843 , \4568 , \3119 );
nor \U$13501 ( \13844 , \13842 , \13843 );
xnor \U$13502 ( \13845 , \13844 , \2916 );
and \U$13503 ( \13846 , \5050 , \2715 );
and \U$13504 ( \13847 , \5045 , \2713 );
nor \U$13505 ( \13848 , \13846 , \13847 );
xnor \U$13506 ( \13849 , \13848 , \2566 );
and \U$13507 ( \13850 , \13845 , \13849 );
and \U$13508 ( \13851 , \5573 , \2393 );
and \U$13509 ( \13852 , \5314 , \2391 );
nor \U$13510 ( \13853 , \13851 , \13852 );
xnor \U$13511 ( \13854 , \13853 , \2251 );
and \U$13512 ( \13855 , \13849 , \13854 );
and \U$13513 ( \13856 , \13845 , \13854 );
or \U$13514 ( \13857 , \13850 , \13855 , \13856 );
and \U$13515 ( \13858 , \3686 , \4152 );
and \U$13516 ( \13859 , \3478 , \4150 );
nor \U$13517 ( \13860 , \13858 , \13859 );
xnor \U$13518 ( \13861 , \13860 , \4009 );
and \U$13519 ( \13862 , \3813 , \3829 );
and \U$13520 ( \13863 , \3808 , \3827 );
nor \U$13521 ( \13864 , \13862 , \13863 );
xnor \U$13522 ( \13865 , \13864 , \3583 );
and \U$13523 ( \13866 , \13861 , \13865 );
and \U$13524 ( \13867 , \4266 , \3434 );
and \U$13525 ( \13868 , \4069 , \3432 );
nor \U$13526 ( \13869 , \13867 , \13868 );
xnor \U$13527 ( \13870 , \13869 , \3247 );
and \U$13528 ( \13871 , \13865 , \13870 );
and \U$13529 ( \13872 , \13861 , \13870 );
or \U$13530 ( \13873 , \13866 , \13871 , \13872 );
and \U$13531 ( \13874 , \13857 , \13873 );
and \U$13532 ( \13875 , \2463 , \5443 );
and \U$13533 ( \13876 , \2438 , \5441 );
nor \U$13534 ( \13877 , \13875 , \13876 );
xnor \U$13535 ( \13878 , \13877 , \5202 );
and \U$13536 ( \13879 , \2804 , \4977 );
and \U$13537 ( \13880 , \2637 , \4975 );
nor \U$13538 ( \13881 , \13879 , \13880 );
xnor \U$13539 ( \13882 , \13881 , \4789 );
and \U$13540 ( \13883 , \13878 , \13882 );
and \U$13541 ( \13884 , \3061 , \4603 );
and \U$13542 ( \13885 , \2942 , \4601 );
nor \U$13543 ( \13886 , \13884 , \13885 );
xnor \U$13544 ( \13887 , \13886 , \4371 );
and \U$13545 ( \13888 , \13882 , \13887 );
and \U$13546 ( \13889 , \13878 , \13887 );
or \U$13547 ( \13890 , \13883 , \13888 , \13889 );
and \U$13548 ( \13891 , \13873 , \13890 );
and \U$13549 ( \13892 , \13857 , \13890 );
or \U$13550 ( \13893 , \13874 , \13891 , \13892 );
and \U$13551 ( \13894 , \13840 , \13893 );
and \U$13552 ( \13895 , \13788 , \13893 );
or \U$13553 ( \13896 , \13841 , \13894 , \13895 );
and \U$13554 ( \13897 , \13736 , \13896 );
xor \U$13555 ( \13898 , \13313 , \13317 );
xor \U$13556 ( \13899 , \13898 , \13322 );
xor \U$13557 ( \13900 , \13426 , \13428 );
xor \U$13558 ( \13901 , \13900 , \13431 );
and \U$13559 ( \13902 , \13899 , \13901 );
xor \U$13560 ( \13903 , \13436 , \13438 );
xor \U$13561 ( \13904 , \13903 , \13441 );
and \U$13562 ( \13905 , \13901 , \13904 );
and \U$13563 ( \13906 , \13899 , \13904 );
or \U$13564 ( \13907 , \13902 , \13905 , \13906 );
and \U$13565 ( \13908 , \13896 , \13907 );
and \U$13566 ( \13909 , \13736 , \13907 );
or \U$13567 ( \13910 , \13897 , \13908 , \13909 );
xor \U$13568 ( \13911 , \13524 , \13540 );
xor \U$13569 ( \13912 , \13911 , \13557 );
xor \U$13570 ( \13913 , \13577 , \13593 );
xor \U$13571 ( \13914 , \13913 , \13610 );
and \U$13572 ( \13915 , \13912 , \13914 );
xor \U$13573 ( \13916 , \13449 , \13451 );
xor \U$13574 ( \13917 , \13916 , \13454 );
and \U$13575 ( \13918 , \13914 , \13917 );
and \U$13576 ( \13919 , \13912 , \13917 );
or \U$13577 ( \13920 , \13915 , \13918 , \13919 );
xor \U$13578 ( \13921 , \13309 , \13325 );
xor \U$13579 ( \13922 , \13921 , \13342 );
and \U$13580 ( \13923 , \13920 , \13922 );
xor \U$13581 ( \13924 , \13632 , \13634 );
xor \U$13582 ( \13925 , \13924 , \13637 );
and \U$13583 ( \13926 , \13922 , \13925 );
and \U$13584 ( \13927 , \13920 , \13925 );
or \U$13585 ( \13928 , \13923 , \13926 , \13927 );
and \U$13586 ( \13929 , \13910 , \13928 );
xor \U$13587 ( \13930 , \13434 , \13444 );
xor \U$13588 ( \13931 , \13930 , \13457 );
xor \U$13589 ( \13932 , \13508 , \13560 );
xor \U$13590 ( \13933 , \13932 , \13613 );
and \U$13591 ( \13934 , \13931 , \13933 );
xor \U$13592 ( \13935 , \13619 , \13621 );
xor \U$13593 ( \13936 , \13935 , \13624 );
and \U$13594 ( \13937 , \13933 , \13936 );
and \U$13595 ( \13938 , \13931 , \13936 );
or \U$13596 ( \13939 , \13934 , \13937 , \13938 );
and \U$13597 ( \13940 , \13928 , \13939 );
and \U$13598 ( \13941 , \13910 , \13939 );
or \U$13599 ( \13942 , \13929 , \13940 , \13941 );
xor \U$13600 ( \13943 , \13460 , \13616 );
xor \U$13601 ( \13944 , \13943 , \13627 );
xor \U$13602 ( \13945 , \13640 , \13642 );
xor \U$13603 ( \13946 , \13945 , \13645 );
and \U$13604 ( \13947 , \13944 , \13946 );
xor \U$13605 ( \13948 , \13651 , \13653 );
xor \U$13606 ( \13949 , \13948 , \13656 );
and \U$13607 ( \13950 , \13946 , \13949 );
and \U$13608 ( \13951 , \13944 , \13949 );
or \U$13609 ( \13952 , \13947 , \13950 , \13951 );
and \U$13610 ( \13953 , \13942 , \13952 );
xor \U$13611 ( \13954 , \13664 , \13666 );
xor \U$13612 ( \13955 , \13954 , \13669 );
and \U$13613 ( \13956 , \13952 , \13955 );
and \U$13614 ( \13957 , \13942 , \13955 );
or \U$13615 ( \13958 , \13953 , \13956 , \13957 );
xor \U$13616 ( \13959 , \13662 , \13672 );
xor \U$13617 ( \13960 , \13959 , \13675 );
and \U$13618 ( \13961 , \13958 , \13960 );
xor \U$13619 ( \13962 , \13680 , \13682 );
xor \U$13620 ( \13963 , \13962 , \13685 );
and \U$13621 ( \13964 , \13960 , \13963 );
and \U$13622 ( \13965 , \13958 , \13963 );
or \U$13623 ( \13966 , \13961 , \13964 , \13965 );
xor \U$13624 ( \13967 , \13678 , \13688 );
xor \U$13625 ( \13968 , \13967 , \13691 );
and \U$13626 ( \13969 , \13966 , \13968 );
xor \U$13627 ( \13970 , \13394 , \13404 );
xor \U$13628 ( \13971 , \13970 , \13407 );
and \U$13629 ( \13972 , \13968 , \13971 );
and \U$13630 ( \13973 , \13966 , \13971 );
or \U$13631 ( \13974 , \13969 , \13972 , \13973 );
and \U$13632 ( \13975 , \13700 , \13974 );
xor \U$13633 ( \13976 , \13700 , \13974 );
xor \U$13634 ( \13977 , \13966 , \13968 );
xor \U$13635 ( \13978 , \13977 , \13971 );
xor \U$13636 ( \13979 , \13845 , \13849 );
xor \U$13637 ( \13980 , \13979 , \13854 );
xor \U$13638 ( \13981 , \13861 , \13865 );
xor \U$13639 ( \13982 , \13981 , \13870 );
and \U$13640 ( \13983 , \13980 , \13982 );
xor \U$13641 ( \13984 , \13878 , \13882 );
xor \U$13642 ( \13985 , \13984 , \13887 );
and \U$13643 ( \13986 , \13982 , \13985 );
and \U$13644 ( \13987 , \13980 , \13985 );
or \U$13645 ( \13988 , \13983 , \13986 , \13987 );
xor \U$13646 ( \13989 , \13740 , \13744 );
xor \U$13647 ( \13990 , \13989 , \13749 );
xor \U$13648 ( \13991 , \13756 , \13760 );
xor \U$13649 ( \13992 , \13991 , \13765 );
and \U$13650 ( \13993 , \13990 , \13992 );
xor \U$13651 ( \13994 , \13773 , \13777 );
xor \U$13652 ( \13995 , \13994 , \13782 );
and \U$13653 ( \13996 , \13992 , \13995 );
and \U$13654 ( \13997 , \13990 , \13995 );
or \U$13655 ( \13998 , \13993 , \13996 , \13997 );
and \U$13656 ( \13999 , \13988 , \13998 );
xor \U$13657 ( \14000 , \13792 , \13796 );
xor \U$13658 ( \14001 , \14000 , \13801 );
xor \U$13659 ( \14002 , \13808 , \13812 );
xor \U$13660 ( \14003 , \14002 , \13817 );
and \U$13661 ( \14004 , \14001 , \14003 );
xor \U$13662 ( \14005 , \13825 , \13829 );
xor \U$13663 ( \14006 , \14005 , \13834 );
and \U$13664 ( \14007 , \14003 , \14006 );
and \U$13665 ( \14008 , \14001 , \14006 );
or \U$13666 ( \14009 , \14004 , \14007 , \14008 );
and \U$13667 ( \14010 , \13998 , \14009 );
and \U$13668 ( \14011 , \13988 , \14009 );
or \U$13669 ( \14012 , \13999 , \14010 , \14011 );
and \U$13670 ( \14013 , \4568 , \3434 );
and \U$13671 ( \14014 , \4266 , \3432 );
nor \U$13672 ( \14015 , \14013 , \14014 );
xnor \U$13673 ( \14016 , \14015 , \3247 );
and \U$13674 ( \14017 , \5045 , \3121 );
and \U$13675 ( \14018 , \4576 , \3119 );
nor \U$13676 ( \14019 , \14017 , \14018 );
xnor \U$13677 ( \14020 , \14019 , \2916 );
and \U$13678 ( \14021 , \14016 , \14020 );
and \U$13679 ( \14022 , \5314 , \2715 );
and \U$13680 ( \14023 , \5050 , \2713 );
nor \U$13681 ( \14024 , \14022 , \14023 );
xnor \U$13682 ( \14025 , \14024 , \2566 );
and \U$13683 ( \14026 , \14020 , \14025 );
and \U$13684 ( \14027 , \14016 , \14025 );
or \U$13685 ( \14028 , \14021 , \14026 , \14027 );
and \U$13686 ( \14029 , \2438 , \6032 );
and \U$13687 ( \14030 , \2174 , \6030 );
nor \U$13688 ( \14031 , \14029 , \14030 );
xnor \U$13689 ( \14032 , \14031 , \5692 );
and \U$13690 ( \14033 , \2637 , \5443 );
and \U$13691 ( \14034 , \2463 , \5441 );
nor \U$13692 ( \14035 , \14033 , \14034 );
xnor \U$13693 ( \14036 , \14035 , \5202 );
and \U$13694 ( \14037 , \14032 , \14036 );
and \U$13695 ( \14038 , \2942 , \4977 );
and \U$13696 ( \14039 , \2804 , \4975 );
nor \U$13697 ( \14040 , \14038 , \14039 );
xnor \U$13698 ( \14041 , \14040 , \4789 );
and \U$13699 ( \14042 , \14036 , \14041 );
and \U$13700 ( \14043 , \14032 , \14041 );
or \U$13701 ( \14044 , \14037 , \14042 , \14043 );
and \U$13702 ( \14045 , \14028 , \14044 );
and \U$13703 ( \14046 , \3478 , \4603 );
and \U$13704 ( \14047 , \3061 , \4601 );
nor \U$13705 ( \14048 , \14046 , \14047 );
xnor \U$13706 ( \14049 , \14048 , \4371 );
and \U$13707 ( \14050 , \3808 , \4152 );
and \U$13708 ( \14051 , \3686 , \4150 );
nor \U$13709 ( \14052 , \14050 , \14051 );
xnor \U$13710 ( \14053 , \14052 , \4009 );
and \U$13711 ( \14054 , \14049 , \14053 );
and \U$13712 ( \14055 , \4069 , \3829 );
and \U$13713 ( \14056 , \3813 , \3827 );
nor \U$13714 ( \14057 , \14055 , \14056 );
xnor \U$13715 ( \14058 , \14057 , \3583 );
and \U$13716 ( \14059 , \14053 , \14058 );
and \U$13717 ( \14060 , \14049 , \14058 );
or \U$13718 ( \14061 , \14054 , \14059 , \14060 );
and \U$13719 ( \14062 , \14044 , \14061 );
and \U$13720 ( \14063 , \14028 , \14061 );
or \U$13721 ( \14064 , \14045 , \14062 , \14063 );
and \U$13722 ( \14065 , \983 , \9230 );
and \U$13723 ( \14066 , \785 , \9228 );
nor \U$13724 ( \14067 , \14065 , \14066 );
xnor \U$13725 ( \14068 , \14067 , \8920 );
and \U$13726 ( \14069 , \1176 , \8693 );
and \U$13727 ( \14070 , \1071 , \8691 );
nor \U$13728 ( \14071 , \14069 , \14070 );
xnor \U$13729 ( \14072 , \14071 , \8322 );
and \U$13730 ( \14073 , \14068 , \14072 );
and \U$13731 ( \14074 , \1297 , \8131 );
and \U$13732 ( \14075 , \1181 , \8129 );
nor \U$13733 ( \14076 , \14074 , \14075 );
xnor \U$13734 ( \14077 , \14076 , \7813 );
and \U$13735 ( \14078 , \14072 , \14077 );
and \U$13736 ( \14079 , \14068 , \14077 );
or \U$13737 ( \14080 , \14073 , \14078 , \14079 );
and \U$13738 ( \14081 , \450 , \10611 );
and \U$13739 ( \14082 , \435 , \10608 );
nor \U$13740 ( \14083 , \14081 , \14082 );
xnor \U$13741 ( \14084 , \14083 , \9556 );
and \U$13742 ( \14085 , \722 , \9798 );
and \U$13743 ( \14086 , \661 , \9796 );
nor \U$13744 ( \14087 , \14085 , \14086 );
xnor \U$13745 ( \14088 , \14087 , \9559 );
and \U$13746 ( \14089 , \14084 , \14088 );
and \U$13747 ( \14090 , \14088 , \364 );
and \U$13748 ( \14091 , \14084 , \364 );
or \U$13749 ( \14092 , \14089 , \14090 , \14091 );
and \U$13750 ( \14093 , \14080 , \14092 );
and \U$13751 ( \14094 , \1588 , \7564 );
and \U$13752 ( \14095 , \1412 , \7562 );
nor \U$13753 ( \14096 , \14094 , \14095 );
xnor \U$13754 ( \14097 , \14096 , \7315 );
and \U$13755 ( \14098 , \1839 , \7035 );
and \U$13756 ( \14099 , \1596 , \7033 );
nor \U$13757 ( \14100 , \14098 , \14099 );
xnor \U$13758 ( \14101 , \14100 , \6775 );
and \U$13759 ( \14102 , \14097 , \14101 );
and \U$13760 ( \14103 , \2030 , \6541 );
and \U$13761 ( \14104 , \1844 , \6539 );
nor \U$13762 ( \14105 , \14103 , \14104 );
xnor \U$13763 ( \14106 , \14105 , \6226 );
and \U$13764 ( \14107 , \14101 , \14106 );
and \U$13765 ( \14108 , \14097 , \14106 );
or \U$13766 ( \14109 , \14102 , \14107 , \14108 );
and \U$13767 ( \14110 , \14092 , \14109 );
and \U$13768 ( \14111 , \14080 , \14109 );
or \U$13769 ( \14112 , \14093 , \14110 , \14111 );
and \U$13770 ( \14113 , \14064 , \14112 );
and \U$13771 ( \14114 , \9347 , \957 );
and \U$13772 ( \14115 , \8778 , \955 );
nor \U$13773 ( \14116 , \14114 , \14115 );
xnor \U$13774 ( \14117 , \14116 , \879 );
and \U$13775 ( \14118 , \9958 , \793 );
and \U$13776 ( \14119 , \9355 , \791 );
nor \U$13777 ( \14120 , \14118 , \14119 );
xnor \U$13778 ( \14121 , \14120 , \699 );
and \U$13779 ( \14122 , \14117 , \14121 );
and \U$13780 ( \14123 , \10144 , \624 );
and \U$13781 ( \14124 , \9963 , \622 );
nor \U$13782 ( \14125 , \14123 , \14124 );
xnor \U$13783 ( \14126 , \14125 , \349 );
and \U$13784 ( \14127 , \14121 , \14126 );
and \U$13785 ( \14128 , \14117 , \14126 );
or \U$13786 ( \14129 , \14122 , \14127 , \14128 );
and \U$13787 ( \14130 , \5945 , \2393 );
and \U$13788 ( \14131 , \5573 , \2391 );
nor \U$13789 ( \14132 , \14130 , \14131 );
xnor \U$13790 ( \14133 , \14132 , \2251 );
and \U$13791 ( \14134 , \6297 , \2097 );
and \U$13792 ( \14135 , \5954 , \2095 );
nor \U$13793 ( \14136 , \14134 , \14135 );
xnor \U$13794 ( \14137 , \14136 , \1960 );
and \U$13795 ( \14138 , \14133 , \14137 );
and \U$13796 ( \14139 , \6802 , \1891 );
and \U$13797 ( \14140 , \6499 , \1889 );
nor \U$13798 ( \14141 , \14139 , \14140 );
xnor \U$13799 ( \14142 , \14141 , \1739 );
and \U$13800 ( \14143 , \14137 , \14142 );
and \U$13801 ( \14144 , \14133 , \14142 );
or \U$13802 ( \14145 , \14138 , \14143 , \14144 );
and \U$13803 ( \14146 , \14129 , \14145 );
and \U$13804 ( \14147 , \7500 , \1623 );
and \U$13805 ( \14148 , \6974 , \1621 );
nor \U$13806 ( \14149 , \14147 , \14148 );
xnor \U$13807 ( \14150 , \14149 , \1467 );
and \U$13808 ( \14151 , \8170 , \1351 );
and \U$13809 ( \14152 , \7924 , \1349 );
nor \U$13810 ( \14153 , \14151 , \14152 );
xnor \U$13811 ( \14154 , \14153 , \1238 );
and \U$13812 ( \14155 , \14150 , \14154 );
and \U$13813 ( \14156 , \8494 , \1157 );
and \U$13814 ( \14157 , \8175 , \1155 );
nor \U$13815 ( \14158 , \14156 , \14157 );
xnor \U$13816 ( \14159 , \14158 , \1021 );
and \U$13817 ( \14160 , \14154 , \14159 );
and \U$13818 ( \14161 , \14150 , \14159 );
or \U$13819 ( \14162 , \14155 , \14160 , \14161 );
and \U$13820 ( \14163 , \14145 , \14162 );
and \U$13821 ( \14164 , \14129 , \14162 );
or \U$13822 ( \14165 , \14146 , \14163 , \14164 );
and \U$13823 ( \14166 , \14112 , \14165 );
and \U$13824 ( \14167 , \14064 , \14165 );
or \U$13825 ( \14168 , \14113 , \14166 , \14167 );
and \U$13826 ( \14169 , \14012 , \14168 );
xor \U$13827 ( \14170 , \13480 , \13484 );
xor \U$13828 ( \14171 , \14170 , \13489 );
xor \U$13829 ( \14172 , \13497 , \13501 );
xor \U$13830 ( \14173 , \14172 , \380 );
and \U$13831 ( \14174 , \14171 , \14173 );
xor \U$13832 ( \14175 , \13725 , \13727 );
xor \U$13833 ( \14176 , \14175 , \13730 );
and \U$13834 ( \14177 , \14173 , \14176 );
and \U$13835 ( \14178 , \14171 , \14176 );
or \U$13836 ( \14179 , \14174 , \14177 , \14178 );
and \U$13837 ( \14180 , \14168 , \14179 );
and \U$13838 ( \14181 , \14012 , \14179 );
or \U$13839 ( \14182 , \14169 , \14180 , \14181 );
xor \U$13840 ( \14183 , \13752 , \13768 );
xor \U$13841 ( \14184 , \14183 , \13785 );
xor \U$13842 ( \14185 , \13702 , \13704 );
xor \U$13843 ( \14186 , \14185 , \13707 );
and \U$13844 ( \14187 , \14184 , \14186 );
xor \U$13845 ( \14188 , \13714 , \13716 );
xor \U$13846 ( \14189 , \14188 , \13719 );
and \U$13847 ( \14190 , \14186 , \14189 );
and \U$13848 ( \14191 , \14184 , \14189 );
or \U$13849 ( \14192 , \14187 , \14190 , \14191 );
xor \U$13850 ( \14193 , \13804 , \13820 );
xor \U$13851 ( \14194 , \14193 , \13837 );
xor \U$13852 ( \14195 , \13857 , \13873 );
xor \U$13853 ( \14196 , \14195 , \13890 );
and \U$13854 ( \14197 , \14194 , \14196 );
and \U$13855 ( \14198 , \14192 , \14197 );
xor \U$13856 ( \14199 , \13476 , \13492 );
xor \U$13857 ( \14200 , \14199 , \13505 );
and \U$13858 ( \14201 , \14197 , \14200 );
and \U$13859 ( \14202 , \14192 , \14200 );
or \U$13860 ( \14203 , \14198 , \14201 , \14202 );
and \U$13861 ( \14204 , \14182 , \14203 );
xor \U$13862 ( \14205 , \13710 , \13722 );
xor \U$13863 ( \14206 , \14205 , \13733 );
xor \U$13864 ( \14207 , \13912 , \13914 );
xor \U$13865 ( \14208 , \14207 , \13917 );
and \U$13866 ( \14209 , \14206 , \14208 );
xor \U$13867 ( \14210 , \13899 , \13901 );
xor \U$13868 ( \14211 , \14210 , \13904 );
and \U$13869 ( \14212 , \14208 , \14211 );
and \U$13870 ( \14213 , \14206 , \14211 );
or \U$13871 ( \14214 , \14209 , \14212 , \14213 );
and \U$13872 ( \14215 , \14203 , \14214 );
and \U$13873 ( \14216 , \14182 , \14214 );
or \U$13874 ( \14217 , \14204 , \14215 , \14216 );
xor \U$13875 ( \14218 , \13736 , \13896 );
xor \U$13876 ( \14219 , \14218 , \13907 );
xor \U$13877 ( \14220 , \13920 , \13922 );
xor \U$13878 ( \14221 , \14220 , \13925 );
and \U$13879 ( \14222 , \14219 , \14221 );
xor \U$13880 ( \14223 , \13931 , \13933 );
xor \U$13881 ( \14224 , \14223 , \13936 );
and \U$13882 ( \14225 , \14221 , \14224 );
and \U$13883 ( \14226 , \14219 , \14224 );
or \U$13884 ( \14227 , \14222 , \14225 , \14226 );
and \U$13885 ( \14228 , \14217 , \14227 );
xor \U$13886 ( \14229 , \13944 , \13946 );
xor \U$13887 ( \14230 , \14229 , \13949 );
and \U$13888 ( \14231 , \14227 , \14230 );
and \U$13889 ( \14232 , \14217 , \14230 );
or \U$13890 ( \14233 , \14228 , \14231 , \14232 );
xor \U$13891 ( \14234 , \13630 , \13648 );
xor \U$13892 ( \14235 , \14234 , \13659 );
and \U$13893 ( \14236 , \14233 , \14235 );
xor \U$13894 ( \14237 , \13942 , \13952 );
xor \U$13895 ( \14238 , \14237 , \13955 );
and \U$13896 ( \14239 , \14235 , \14238 );
and \U$13897 ( \14240 , \14233 , \14238 );
or \U$13898 ( \14241 , \14236 , \14239 , \14240 );
xor \U$13899 ( \14242 , \13958 , \13960 );
xor \U$13900 ( \14243 , \14242 , \13963 );
and \U$13901 ( \14244 , \14241 , \14243 );
and \U$13902 ( \14245 , \13978 , \14244 );
xor \U$13903 ( \14246 , \13978 , \14244 );
xor \U$13904 ( \14247 , \14241 , \14243 );
and \U$13905 ( \14248 , \3813 , \4152 );
and \U$13906 ( \14249 , \3808 , \4150 );
nor \U$13907 ( \14250 , \14248 , \14249 );
xnor \U$13908 ( \14251 , \14250 , \4009 );
and \U$13909 ( \14252 , \4266 , \3829 );
and \U$13910 ( \14253 , \4069 , \3827 );
nor \U$13911 ( \14254 , \14252 , \14253 );
xnor \U$13912 ( \14255 , \14254 , \3583 );
and \U$13913 ( \14256 , \14251 , \14255 );
and \U$13914 ( \14257 , \4576 , \3434 );
and \U$13915 ( \14258 , \4568 , \3432 );
nor \U$13916 ( \14259 , \14257 , \14258 );
xnor \U$13917 ( \14260 , \14259 , \3247 );
and \U$13918 ( \14261 , \14255 , \14260 );
and \U$13919 ( \14262 , \14251 , \14260 );
or \U$13920 ( \14263 , \14256 , \14261 , \14262 );
and \U$13921 ( \14264 , \2804 , \5443 );
and \U$13922 ( \14265 , \2637 , \5441 );
nor \U$13923 ( \14266 , \14264 , \14265 );
xnor \U$13924 ( \14267 , \14266 , \5202 );
and \U$13925 ( \14268 , \3061 , \4977 );
and \U$13926 ( \14269 , \2942 , \4975 );
nor \U$13927 ( \14270 , \14268 , \14269 );
xnor \U$13928 ( \14271 , \14270 , \4789 );
and \U$13929 ( \14272 , \14267 , \14271 );
and \U$13930 ( \14273 , \3686 , \4603 );
and \U$13931 ( \14274 , \3478 , \4601 );
nor \U$13932 ( \14275 , \14273 , \14274 );
xnor \U$13933 ( \14276 , \14275 , \4371 );
and \U$13934 ( \14277 , \14271 , \14276 );
and \U$13935 ( \14278 , \14267 , \14276 );
or \U$13936 ( \14279 , \14272 , \14277 , \14278 );
and \U$13937 ( \14280 , \14263 , \14279 );
and \U$13938 ( \14281 , \5050 , \3121 );
and \U$13939 ( \14282 , \5045 , \3119 );
nor \U$13940 ( \14283 , \14281 , \14282 );
xnor \U$13941 ( \14284 , \14283 , \2916 );
and \U$13942 ( \14285 , \5573 , \2715 );
and \U$13943 ( \14286 , \5314 , \2713 );
nor \U$13944 ( \14287 , \14285 , \14286 );
xnor \U$13945 ( \14288 , \14287 , \2566 );
and \U$13946 ( \14289 , \14284 , \14288 );
and \U$13947 ( \14290 , \5954 , \2393 );
and \U$13948 ( \14291 , \5945 , \2391 );
nor \U$13949 ( \14292 , \14290 , \14291 );
xnor \U$13950 ( \14293 , \14292 , \2251 );
and \U$13951 ( \14294 , \14288 , \14293 );
and \U$13952 ( \14295 , \14284 , \14293 );
or \U$13953 ( \14296 , \14289 , \14294 , \14295 );
and \U$13954 ( \14297 , \14279 , \14296 );
and \U$13955 ( \14298 , \14263 , \14296 );
or \U$13956 ( \14299 , \14280 , \14297 , \14298 );
and \U$13957 ( \14300 , \8175 , \1351 );
and \U$13958 ( \14301 , \8170 , \1349 );
nor \U$13959 ( \14302 , \14300 , \14301 );
xnor \U$13960 ( \14303 , \14302 , \1238 );
and \U$13961 ( \14304 , \8778 , \1157 );
and \U$13962 ( \14305 , \8494 , \1155 );
nor \U$13963 ( \14306 , \14304 , \14305 );
xnor \U$13964 ( \14307 , \14306 , \1021 );
and \U$13965 ( \14308 , \14303 , \14307 );
and \U$13966 ( \14309 , \9355 , \957 );
and \U$13967 ( \14310 , \9347 , \955 );
nor \U$13968 ( \14311 , \14309 , \14310 );
xnor \U$13969 ( \14312 , \14311 , \879 );
and \U$13970 ( \14313 , \14307 , \14312 );
and \U$13971 ( \14314 , \14303 , \14312 );
or \U$13972 ( \14315 , \14308 , \14313 , \14314 );
and \U$13973 ( \14316 , \6499 , \2097 );
and \U$13974 ( \14317 , \6297 , \2095 );
nor \U$13975 ( \14318 , \14316 , \14317 );
xnor \U$13976 ( \14319 , \14318 , \1960 );
and \U$13977 ( \14320 , \6974 , \1891 );
and \U$13978 ( \14321 , \6802 , \1889 );
nor \U$13979 ( \14322 , \14320 , \14321 );
xnor \U$13980 ( \14323 , \14322 , \1739 );
and \U$13981 ( \14324 , \14319 , \14323 );
and \U$13982 ( \14325 , \7924 , \1623 );
and \U$13983 ( \14326 , \7500 , \1621 );
nor \U$13984 ( \14327 , \14325 , \14326 );
xnor \U$13985 ( \14328 , \14327 , \1467 );
and \U$13986 ( \14329 , \14323 , \14328 );
and \U$13987 ( \14330 , \14319 , \14328 );
or \U$13988 ( \14331 , \14324 , \14329 , \14330 );
and \U$13989 ( \14332 , \14315 , \14331 );
and \U$13990 ( \14333 , \9963 , \793 );
and \U$13991 ( \14334 , \9958 , \791 );
nor \U$13992 ( \14335 , \14333 , \14334 );
xnor \U$13993 ( \14336 , \14335 , \699 );
and \U$13994 ( \14337 , \10764 , \624 );
and \U$13995 ( \14338 , \10144 , \622 );
nor \U$13996 ( \14339 , \14337 , \14338 );
xnor \U$13997 ( \14340 , \14339 , \349 );
and \U$13998 ( \14341 , \14336 , \14340 );
and \U$13999 ( \14342 , \14331 , \14341 );
and \U$14000 ( \14343 , \14315 , \14341 );
or \U$14001 ( \14344 , \14332 , \14342 , \14343 );
and \U$14002 ( \14345 , \14299 , \14344 );
and \U$14003 ( \14346 , \1844 , \7035 );
and \U$14004 ( \14347 , \1839 , \7033 );
nor \U$14005 ( \14348 , \14346 , \14347 );
xnor \U$14006 ( \14349 , \14348 , \6775 );
and \U$14007 ( \14350 , \2174 , \6541 );
and \U$14008 ( \14351 , \2030 , \6539 );
nor \U$14009 ( \14352 , \14350 , \14351 );
xnor \U$14010 ( \14353 , \14352 , \6226 );
and \U$14011 ( \14354 , \14349 , \14353 );
and \U$14012 ( \14355 , \2463 , \6032 );
and \U$14013 ( \14356 , \2438 , \6030 );
nor \U$14014 ( \14357 , \14355 , \14356 );
xnor \U$14015 ( \14358 , \14357 , \5692 );
and \U$14016 ( \14359 , \14353 , \14358 );
and \U$14017 ( \14360 , \14349 , \14358 );
or \U$14018 ( \14361 , \14354 , \14359 , \14360 );
and \U$14019 ( \14362 , \661 , \10611 );
and \U$14020 ( \14363 , \450 , \10608 );
nor \U$14021 ( \14364 , \14362 , \14363 );
xnor \U$14022 ( \14365 , \14364 , \9556 );
and \U$14023 ( \14366 , \785 , \9798 );
and \U$14024 ( \14367 , \722 , \9796 );
nor \U$14025 ( \14368 , \14366 , \14367 );
xnor \U$14026 ( \14369 , \14368 , \9559 );
and \U$14027 ( \14370 , \14365 , \14369 );
and \U$14028 ( \14371 , \1071 , \9230 );
and \U$14029 ( \14372 , \983 , \9228 );
nor \U$14030 ( \14373 , \14371 , \14372 );
xnor \U$14031 ( \14374 , \14373 , \8920 );
and \U$14032 ( \14375 , \14369 , \14374 );
and \U$14033 ( \14376 , \14365 , \14374 );
or \U$14034 ( \14377 , \14370 , \14375 , \14376 );
and \U$14035 ( \14378 , \14361 , \14377 );
and \U$14036 ( \14379 , \1181 , \8693 );
and \U$14037 ( \14380 , \1176 , \8691 );
nor \U$14038 ( \14381 , \14379 , \14380 );
xnor \U$14039 ( \14382 , \14381 , \8322 );
and \U$14040 ( \14383 , \1412 , \8131 );
and \U$14041 ( \14384 , \1297 , \8129 );
nor \U$14042 ( \14385 , \14383 , \14384 );
xnor \U$14043 ( \14386 , \14385 , \7813 );
and \U$14044 ( \14387 , \14382 , \14386 );
and \U$14045 ( \14388 , \1596 , \7564 );
and \U$14046 ( \14389 , \1588 , \7562 );
nor \U$14047 ( \14390 , \14388 , \14389 );
xnor \U$14048 ( \14391 , \14390 , \7315 );
and \U$14049 ( \14392 , \14386 , \14391 );
and \U$14050 ( \14393 , \14382 , \14391 );
or \U$14051 ( \14394 , \14387 , \14392 , \14393 );
and \U$14052 ( \14395 , \14377 , \14394 );
and \U$14053 ( \14396 , \14361 , \14394 );
or \U$14054 ( \14397 , \14378 , \14395 , \14396 );
and \U$14055 ( \14398 , \14344 , \14397 );
and \U$14056 ( \14399 , \14299 , \14397 );
or \U$14057 ( \14400 , \14345 , \14398 , \14399 );
xor \U$14058 ( \14401 , \14068 , \14072 );
xor \U$14059 ( \14402 , \14401 , \14077 );
xor \U$14060 ( \14403 , \14097 , \14101 );
xor \U$14061 ( \14404 , \14403 , \14106 );
and \U$14062 ( \14405 , \14402 , \14404 );
xor \U$14063 ( \14406 , \14032 , \14036 );
xor \U$14064 ( \14407 , \14406 , \14041 );
and \U$14065 ( \14408 , \14404 , \14407 );
and \U$14066 ( \14409 , \14402 , \14407 );
or \U$14067 ( \14410 , \14405 , \14408 , \14409 );
nand \U$14068 ( \14411 , \10764 , \355 );
xnor \U$14069 ( \14412 , \14411 , \364 );
xor \U$14070 ( \14413 , \14117 , \14121 );
xor \U$14071 ( \14414 , \14413 , \14126 );
and \U$14072 ( \14415 , \14412 , \14414 );
xor \U$14073 ( \14416 , \14150 , \14154 );
xor \U$14074 ( \14417 , \14416 , \14159 );
and \U$14075 ( \14418 , \14414 , \14417 );
and \U$14076 ( \14419 , \14412 , \14417 );
or \U$14077 ( \14420 , \14415 , \14418 , \14419 );
and \U$14078 ( \14421 , \14410 , \14420 );
xor \U$14079 ( \14422 , \14133 , \14137 );
xor \U$14080 ( \14423 , \14422 , \14142 );
xor \U$14081 ( \14424 , \14016 , \14020 );
xor \U$14082 ( \14425 , \14424 , \14025 );
and \U$14083 ( \14426 , \14423 , \14425 );
xor \U$14084 ( \14427 , \14049 , \14053 );
xor \U$14085 ( \14428 , \14427 , \14058 );
and \U$14086 ( \14429 , \14425 , \14428 );
and \U$14087 ( \14430 , \14423 , \14428 );
or \U$14088 ( \14431 , \14426 , \14429 , \14430 );
and \U$14089 ( \14432 , \14420 , \14431 );
and \U$14090 ( \14433 , \14410 , \14431 );
or \U$14091 ( \14434 , \14421 , \14432 , \14433 );
and \U$14092 ( \14435 , \14400 , \14434 );
xor \U$14093 ( \14436 , \13980 , \13982 );
xor \U$14094 ( \14437 , \14436 , \13985 );
xor \U$14095 ( \14438 , \13990 , \13992 );
xor \U$14096 ( \14439 , \14438 , \13995 );
and \U$14097 ( \14440 , \14437 , \14439 );
xor \U$14098 ( \14441 , \14001 , \14003 );
xor \U$14099 ( \14442 , \14441 , \14006 );
and \U$14100 ( \14443 , \14439 , \14442 );
and \U$14101 ( \14444 , \14437 , \14442 );
or \U$14102 ( \14445 , \14440 , \14443 , \14444 );
and \U$14103 ( \14446 , \14434 , \14445 );
and \U$14104 ( \14447 , \14400 , \14445 );
or \U$14105 ( \14448 , \14435 , \14446 , \14447 );
xor \U$14106 ( \14449 , \13988 , \13998 );
xor \U$14107 ( \14450 , \14449 , \14009 );
xor \U$14108 ( \14451 , \14064 , \14112 );
xor \U$14109 ( \14452 , \14451 , \14165 );
and \U$14110 ( \14453 , \14450 , \14452 );
xor \U$14111 ( \14454 , \14171 , \14173 );
xor \U$14112 ( \14455 , \14454 , \14176 );
and \U$14113 ( \14456 , \14452 , \14455 );
and \U$14114 ( \14457 , \14450 , \14455 );
or \U$14115 ( \14458 , \14453 , \14456 , \14457 );
and \U$14116 ( \14459 , \14448 , \14458 );
xor \U$14117 ( \14460 , \14028 , \14044 );
xor \U$14118 ( \14461 , \14460 , \14061 );
xor \U$14119 ( \14462 , \14080 , \14092 );
xor \U$14120 ( \14463 , \14462 , \14109 );
and \U$14121 ( \14464 , \14461 , \14463 );
xor \U$14122 ( \14465 , \14129 , \14145 );
xor \U$14123 ( \14466 , \14465 , \14162 );
and \U$14124 ( \14467 , \14463 , \14466 );
and \U$14125 ( \14468 , \14461 , \14466 );
or \U$14126 ( \14469 , \14464 , \14467 , \14468 );
xor \U$14127 ( \14470 , \14184 , \14186 );
xor \U$14128 ( \14471 , \14470 , \14189 );
and \U$14129 ( \14472 , \14469 , \14471 );
xor \U$14130 ( \14473 , \14194 , \14196 );
and \U$14131 ( \14474 , \14471 , \14473 );
and \U$14132 ( \14475 , \14469 , \14473 );
or \U$14133 ( \14476 , \14472 , \14474 , \14475 );
and \U$14134 ( \14477 , \14458 , \14476 );
and \U$14135 ( \14478 , \14448 , \14476 );
or \U$14136 ( \14479 , \14459 , \14477 , \14478 );
xor \U$14137 ( \14480 , \13788 , \13840 );
xor \U$14138 ( \14481 , \14480 , \13893 );
xor \U$14139 ( \14482 , \14192 , \14197 );
xor \U$14140 ( \14483 , \14482 , \14200 );
and \U$14141 ( \14484 , \14481 , \14483 );
xor \U$14142 ( \14485 , \14206 , \14208 );
xor \U$14143 ( \14486 , \14485 , \14211 );
and \U$14144 ( \14487 , \14483 , \14486 );
and \U$14145 ( \14488 , \14481 , \14486 );
or \U$14146 ( \14489 , \14484 , \14487 , \14488 );
and \U$14147 ( \14490 , \14479 , \14489 );
xor \U$14148 ( \14491 , \14219 , \14221 );
xor \U$14149 ( \14492 , \14491 , \14224 );
and \U$14150 ( \14493 , \14489 , \14492 );
and \U$14151 ( \14494 , \14479 , \14492 );
or \U$14152 ( \14495 , \14490 , \14493 , \14494 );
xor \U$14153 ( \14496 , \13910 , \13928 );
xor \U$14154 ( \14497 , \14496 , \13939 );
and \U$14155 ( \14498 , \14495 , \14497 );
xor \U$14156 ( \14499 , \14217 , \14227 );
xor \U$14157 ( \14500 , \14499 , \14230 );
and \U$14158 ( \14501 , \14497 , \14500 );
and \U$14159 ( \14502 , \14495 , \14500 );
or \U$14160 ( \14503 , \14498 , \14501 , \14502 );
xor \U$14161 ( \14504 , \14233 , \14235 );
xor \U$14162 ( \14505 , \14504 , \14238 );
and \U$14163 ( \14506 , \14503 , \14505 );
and \U$14164 ( \14507 , \14247 , \14506 );
xor \U$14165 ( \14508 , \14247 , \14506 );
xor \U$14166 ( \14509 , \14503 , \14505 );
and \U$14167 ( \14510 , \3808 , \4603 );
and \U$14168 ( \14511 , \3686 , \4601 );
nor \U$14169 ( \14512 , \14510 , \14511 );
xnor \U$14170 ( \14513 , \14512 , \4371 );
and \U$14171 ( \14514 , \4069 , \4152 );
and \U$14172 ( \14515 , \3813 , \4150 );
nor \U$14173 ( \14516 , \14514 , \14515 );
xnor \U$14174 ( \14517 , \14516 , \4009 );
and \U$14175 ( \14518 , \14513 , \14517 );
and \U$14176 ( \14519 , \4568 , \3829 );
and \U$14177 ( \14520 , \4266 , \3827 );
nor \U$14178 ( \14521 , \14519 , \14520 );
xnor \U$14179 ( \14522 , \14521 , \3583 );
and \U$14180 ( \14523 , \14517 , \14522 );
and \U$14181 ( \14524 , \14513 , \14522 );
or \U$14182 ( \14525 , \14518 , \14523 , \14524 );
and \U$14183 ( \14526 , \2637 , \6032 );
and \U$14184 ( \14527 , \2463 , \6030 );
nor \U$14185 ( \14528 , \14526 , \14527 );
xnor \U$14186 ( \14529 , \14528 , \5692 );
and \U$14187 ( \14530 , \2942 , \5443 );
and \U$14188 ( \14531 , \2804 , \5441 );
nor \U$14189 ( \14532 , \14530 , \14531 );
xnor \U$14190 ( \14533 , \14532 , \5202 );
and \U$14191 ( \14534 , \14529 , \14533 );
and \U$14192 ( \14535 , \3478 , \4977 );
and \U$14193 ( \14536 , \3061 , \4975 );
nor \U$14194 ( \14537 , \14535 , \14536 );
xnor \U$14195 ( \14538 , \14537 , \4789 );
and \U$14196 ( \14539 , \14533 , \14538 );
and \U$14197 ( \14540 , \14529 , \14538 );
or \U$14198 ( \14541 , \14534 , \14539 , \14540 );
and \U$14199 ( \14542 , \14525 , \14541 );
and \U$14200 ( \14543 , \5045 , \3434 );
and \U$14201 ( \14544 , \4576 , \3432 );
nor \U$14202 ( \14545 , \14543 , \14544 );
xnor \U$14203 ( \14546 , \14545 , \3247 );
and \U$14204 ( \14547 , \5314 , \3121 );
and \U$14205 ( \14548 , \5050 , \3119 );
nor \U$14206 ( \14549 , \14547 , \14548 );
xnor \U$14207 ( \14550 , \14549 , \2916 );
and \U$14208 ( \14551 , \14546 , \14550 );
and \U$14209 ( \14552 , \5945 , \2715 );
and \U$14210 ( \14553 , \5573 , \2713 );
nor \U$14211 ( \14554 , \14552 , \14553 );
xnor \U$14212 ( \14555 , \14554 , \2566 );
and \U$14213 ( \14556 , \14550 , \14555 );
and \U$14214 ( \14557 , \14546 , \14555 );
or \U$14215 ( \14558 , \14551 , \14556 , \14557 );
and \U$14216 ( \14559 , \14541 , \14558 );
and \U$14217 ( \14560 , \14525 , \14558 );
or \U$14218 ( \14561 , \14542 , \14559 , \14560 );
and \U$14219 ( \14562 , \1839 , \7564 );
and \U$14220 ( \14563 , \1596 , \7562 );
nor \U$14221 ( \14564 , \14562 , \14563 );
xnor \U$14222 ( \14565 , \14564 , \7315 );
and \U$14223 ( \14566 , \2030 , \7035 );
and \U$14224 ( \14567 , \1844 , \7033 );
nor \U$14225 ( \14568 , \14566 , \14567 );
xnor \U$14226 ( \14569 , \14568 , \6775 );
and \U$14227 ( \14570 , \14565 , \14569 );
and \U$14228 ( \14571 , \2438 , \6541 );
and \U$14229 ( \14572 , \2174 , \6539 );
nor \U$14230 ( \14573 , \14571 , \14572 );
xnor \U$14231 ( \14574 , \14573 , \6226 );
and \U$14232 ( \14575 , \14569 , \14574 );
and \U$14233 ( \14576 , \14565 , \14574 );
or \U$14234 ( \14577 , \14570 , \14575 , \14576 );
and \U$14235 ( \14578 , \1176 , \9230 );
and \U$14236 ( \14579 , \1071 , \9228 );
nor \U$14237 ( \14580 , \14578 , \14579 );
xnor \U$14238 ( \14581 , \14580 , \8920 );
and \U$14239 ( \14582 , \1297 , \8693 );
and \U$14240 ( \14583 , \1181 , \8691 );
nor \U$14241 ( \14584 , \14582 , \14583 );
xnor \U$14242 ( \14585 , \14584 , \8322 );
and \U$14243 ( \14586 , \14581 , \14585 );
and \U$14244 ( \14587 , \1588 , \8131 );
and \U$14245 ( \14588 , \1412 , \8129 );
nor \U$14246 ( \14589 , \14587 , \14588 );
xnor \U$14247 ( \14590 , \14589 , \7813 );
and \U$14248 ( \14591 , \14585 , \14590 );
and \U$14249 ( \14592 , \14581 , \14590 );
or \U$14250 ( \14593 , \14586 , \14591 , \14592 );
and \U$14251 ( \14594 , \14577 , \14593 );
and \U$14252 ( \14595 , \722 , \10611 );
and \U$14253 ( \14596 , \661 , \10608 );
nor \U$14254 ( \14597 , \14595 , \14596 );
xnor \U$14255 ( \14598 , \14597 , \9556 );
and \U$14256 ( \14599 , \983 , \9798 );
and \U$14257 ( \14600 , \785 , \9796 );
nor \U$14258 ( \14601 , \14599 , \14600 );
xnor \U$14259 ( \14602 , \14601 , \9559 );
and \U$14260 ( \14603 , \14598 , \14602 );
and \U$14261 ( \14604 , \14602 , \349 );
and \U$14262 ( \14605 , \14598 , \349 );
or \U$14263 ( \14606 , \14603 , \14604 , \14605 );
and \U$14264 ( \14607 , \14593 , \14606 );
and \U$14265 ( \14608 , \14577 , \14606 );
or \U$14266 ( \14609 , \14594 , \14607 , \14608 );
and \U$14267 ( \14610 , \14561 , \14609 );
and \U$14268 ( \14611 , \6297 , \2393 );
and \U$14269 ( \14612 , \5954 , \2391 );
nor \U$14270 ( \14613 , \14611 , \14612 );
xnor \U$14271 ( \14614 , \14613 , \2251 );
and \U$14272 ( \14615 , \6802 , \2097 );
and \U$14273 ( \14616 , \6499 , \2095 );
nor \U$14274 ( \14617 , \14615 , \14616 );
xnor \U$14275 ( \14618 , \14617 , \1960 );
and \U$14276 ( \14619 , \14614 , \14618 );
and \U$14277 ( \14620 , \7500 , \1891 );
and \U$14278 ( \14621 , \6974 , \1889 );
nor \U$14279 ( \14622 , \14620 , \14621 );
xnor \U$14280 ( \14623 , \14622 , \1739 );
and \U$14281 ( \14624 , \14618 , \14623 );
and \U$14282 ( \14625 , \14614 , \14623 );
or \U$14283 ( \14626 , \14619 , \14624 , \14625 );
and \U$14284 ( \14627 , \9958 , \957 );
and \U$14285 ( \14628 , \9355 , \955 );
nor \U$14286 ( \14629 , \14627 , \14628 );
xnor \U$14287 ( \14630 , \14629 , \879 );
and \U$14288 ( \14631 , \10144 , \793 );
and \U$14289 ( \14632 , \9963 , \791 );
nor \U$14290 ( \14633 , \14631 , \14632 );
xnor \U$14291 ( \14634 , \14633 , \699 );
and \U$14292 ( \14635 , \14630 , \14634 );
nand \U$14293 ( \14636 , \10764 , \622 );
xnor \U$14294 ( \14637 , \14636 , \349 );
and \U$14295 ( \14638 , \14634 , \14637 );
and \U$14296 ( \14639 , \14630 , \14637 );
or \U$14297 ( \14640 , \14635 , \14638 , \14639 );
and \U$14298 ( \14641 , \14626 , \14640 );
and \U$14299 ( \14642 , \8170 , \1623 );
and \U$14300 ( \14643 , \7924 , \1621 );
nor \U$14301 ( \14644 , \14642 , \14643 );
xnor \U$14302 ( \14645 , \14644 , \1467 );
and \U$14303 ( \14646 , \8494 , \1351 );
and \U$14304 ( \14647 , \8175 , \1349 );
nor \U$14305 ( \14648 , \14646 , \14647 );
xnor \U$14306 ( \14649 , \14648 , \1238 );
and \U$14307 ( \14650 , \14645 , \14649 );
and \U$14308 ( \14651 , \9347 , \1157 );
and \U$14309 ( \14652 , \8778 , \1155 );
nor \U$14310 ( \14653 , \14651 , \14652 );
xnor \U$14311 ( \14654 , \14653 , \1021 );
and \U$14312 ( \14655 , \14649 , \14654 );
and \U$14313 ( \14656 , \14645 , \14654 );
or \U$14314 ( \14657 , \14650 , \14655 , \14656 );
and \U$14315 ( \14658 , \14640 , \14657 );
and \U$14316 ( \14659 , \14626 , \14657 );
or \U$14317 ( \14660 , \14641 , \14658 , \14659 );
and \U$14318 ( \14661 , \14609 , \14660 );
and \U$14319 ( \14662 , \14561 , \14660 );
or \U$14320 ( \14663 , \14610 , \14661 , \14662 );
xor \U$14321 ( \14664 , \14349 , \14353 );
xor \U$14322 ( \14665 , \14664 , \14358 );
xor \U$14323 ( \14666 , \14365 , \14369 );
xor \U$14324 ( \14667 , \14666 , \14374 );
and \U$14325 ( \14668 , \14665 , \14667 );
xor \U$14326 ( \14669 , \14382 , \14386 );
xor \U$14327 ( \14670 , \14669 , \14391 );
and \U$14328 ( \14671 , \14667 , \14670 );
and \U$14329 ( \14672 , \14665 , \14670 );
or \U$14330 ( \14673 , \14668 , \14671 , \14672 );
xor \U$14331 ( \14674 , \14251 , \14255 );
xor \U$14332 ( \14675 , \14674 , \14260 );
xor \U$14333 ( \14676 , \14267 , \14271 );
xor \U$14334 ( \14677 , \14676 , \14276 );
and \U$14335 ( \14678 , \14675 , \14677 );
xor \U$14336 ( \14679 , \14284 , \14288 );
xor \U$14337 ( \14680 , \14679 , \14293 );
and \U$14338 ( \14681 , \14677 , \14680 );
and \U$14339 ( \14682 , \14675 , \14680 );
or \U$14340 ( \14683 , \14678 , \14681 , \14682 );
and \U$14341 ( \14684 , \14673 , \14683 );
xor \U$14342 ( \14685 , \14303 , \14307 );
xor \U$14343 ( \14686 , \14685 , \14312 );
xor \U$14344 ( \14687 , \14319 , \14323 );
xor \U$14345 ( \14688 , \14687 , \14328 );
and \U$14346 ( \14689 , \14686 , \14688 );
xor \U$14347 ( \14690 , \14336 , \14340 );
and \U$14348 ( \14691 , \14688 , \14690 );
and \U$14349 ( \14692 , \14686 , \14690 );
or \U$14350 ( \14693 , \14689 , \14691 , \14692 );
and \U$14351 ( \14694 , \14683 , \14693 );
and \U$14352 ( \14695 , \14673 , \14693 );
or \U$14353 ( \14696 , \14684 , \14694 , \14695 );
and \U$14354 ( \14697 , \14663 , \14696 );
xor \U$14355 ( \14698 , \14084 , \14088 );
xor \U$14356 ( \14699 , \14698 , \364 );
xor \U$14357 ( \14700 , \14402 , \14404 );
xor \U$14358 ( \14701 , \14700 , \14407 );
and \U$14359 ( \14702 , \14699 , \14701 );
xor \U$14360 ( \14703 , \14423 , \14425 );
xor \U$14361 ( \14704 , \14703 , \14428 );
and \U$14362 ( \14705 , \14701 , \14704 );
and \U$14363 ( \14706 , \14699 , \14704 );
or \U$14364 ( \14707 , \14702 , \14705 , \14706 );
and \U$14365 ( \14708 , \14696 , \14707 );
and \U$14366 ( \14709 , \14663 , \14707 );
or \U$14367 ( \14710 , \14697 , \14708 , \14709 );
xor \U$14368 ( \14711 , \14263 , \14279 );
xor \U$14369 ( \14712 , \14711 , \14296 );
xor \U$14370 ( \14713 , \14315 , \14331 );
xor \U$14371 ( \14714 , \14713 , \14341 );
and \U$14372 ( \14715 , \14712 , \14714 );
xor \U$14373 ( \14716 , \14412 , \14414 );
xor \U$14374 ( \14717 , \14716 , \14417 );
and \U$14375 ( \14718 , \14714 , \14717 );
and \U$14376 ( \14719 , \14712 , \14717 );
or \U$14377 ( \14720 , \14715 , \14718 , \14719 );
xor \U$14378 ( \14721 , \14461 , \14463 );
xor \U$14379 ( \14722 , \14721 , \14466 );
and \U$14380 ( \14723 , \14720 , \14722 );
xor \U$14381 ( \14724 , \14437 , \14439 );
xor \U$14382 ( \14725 , \14724 , \14442 );
and \U$14383 ( \14726 , \14722 , \14725 );
and \U$14384 ( \14727 , \14720 , \14725 );
or \U$14385 ( \14728 , \14723 , \14726 , \14727 );
and \U$14386 ( \14729 , \14710 , \14728 );
xor \U$14387 ( \14730 , \14299 , \14344 );
xor \U$14388 ( \14731 , \14730 , \14397 );
xor \U$14389 ( \14732 , \14410 , \14420 );
xor \U$14390 ( \14733 , \14732 , \14431 );
and \U$14391 ( \14734 , \14731 , \14733 );
and \U$14392 ( \14735 , \14728 , \14734 );
and \U$14393 ( \14736 , \14710 , \14734 );
or \U$14394 ( \14737 , \14729 , \14735 , \14736 );
xor \U$14395 ( \14738 , \14400 , \14434 );
xor \U$14396 ( \14739 , \14738 , \14445 );
xor \U$14397 ( \14740 , \14450 , \14452 );
xor \U$14398 ( \14741 , \14740 , \14455 );
and \U$14399 ( \14742 , \14739 , \14741 );
xor \U$14400 ( \14743 , \14469 , \14471 );
xor \U$14401 ( \14744 , \14743 , \14473 );
and \U$14402 ( \14745 , \14741 , \14744 );
and \U$14403 ( \14746 , \14739 , \14744 );
or \U$14404 ( \14747 , \14742 , \14745 , \14746 );
and \U$14405 ( \14748 , \14737 , \14747 );
xor \U$14406 ( \14749 , \14012 , \14168 );
xor \U$14407 ( \14750 , \14749 , \14179 );
and \U$14408 ( \14751 , \14747 , \14750 );
and \U$14409 ( \14752 , \14737 , \14750 );
or \U$14410 ( \14753 , \14748 , \14751 , \14752 );
xor \U$14411 ( \14754 , \14448 , \14458 );
xor \U$14412 ( \14755 , \14754 , \14476 );
xor \U$14413 ( \14756 , \14481 , \14483 );
xor \U$14414 ( \14757 , \14756 , \14486 );
and \U$14415 ( \14758 , \14755 , \14757 );
and \U$14416 ( \14759 , \14753 , \14758 );
xor \U$14417 ( \14760 , \14182 , \14203 );
xor \U$14418 ( \14761 , \14760 , \14214 );
and \U$14419 ( \14762 , \14758 , \14761 );
and \U$14420 ( \14763 , \14753 , \14761 );
or \U$14421 ( \14764 , \14759 , \14762 , \14763 );
xor \U$14422 ( \14765 , \14495 , \14497 );
xor \U$14423 ( \14766 , \14765 , \14500 );
and \U$14424 ( \14767 , \14764 , \14766 );
and \U$14425 ( \14768 , \14509 , \14767 );
xor \U$14426 ( \14769 , \14509 , \14767 );
xor \U$14427 ( \14770 , \14764 , \14766 );
xor \U$14428 ( \14771 , \14753 , \14758 );
xor \U$14429 ( \14772 , \14771 , \14761 );
xor \U$14430 ( \14773 , \14479 , \14489 );
xor \U$14431 ( \14774 , \14773 , \14492 );
and \U$14432 ( \14775 , \14772 , \14774 );
and \U$14433 ( \14776 , \14770 , \14775 );
xor \U$14434 ( \14777 , \14770 , \14775 );
xor \U$14435 ( \14778 , \14772 , \14774 );
and \U$14436 ( \14779 , \2174 , \7035 );
and \U$14437 ( \14780 , \2030 , \7033 );
nor \U$14438 ( \14781 , \14779 , \14780 );
xnor \U$14439 ( \14782 , \14781 , \6775 );
and \U$14440 ( \14783 , \2463 , \6541 );
and \U$14441 ( \14784 , \2438 , \6539 );
nor \U$14442 ( \14785 , \14783 , \14784 );
xnor \U$14443 ( \14786 , \14785 , \6226 );
and \U$14444 ( \14787 , \14782 , \14786 );
and \U$14445 ( \14788 , \2804 , \6032 );
and \U$14446 ( \14789 , \2637 , \6030 );
nor \U$14447 ( \14790 , \14788 , \14789 );
xnor \U$14448 ( \14791 , \14790 , \5692 );
and \U$14449 ( \14792 , \14786 , \14791 );
and \U$14450 ( \14793 , \14782 , \14791 );
or \U$14451 ( \14794 , \14787 , \14792 , \14793 );
and \U$14452 ( \14795 , \785 , \10611 );
and \U$14453 ( \14796 , \722 , \10608 );
nor \U$14454 ( \14797 , \14795 , \14796 );
xnor \U$14455 ( \14798 , \14797 , \9556 );
and \U$14456 ( \14799 , \1071 , \9798 );
and \U$14457 ( \14800 , \983 , \9796 );
nor \U$14458 ( \14801 , \14799 , \14800 );
xnor \U$14459 ( \14802 , \14801 , \9559 );
and \U$14460 ( \14803 , \14798 , \14802 );
and \U$14461 ( \14804 , \1181 , \9230 );
and \U$14462 ( \14805 , \1176 , \9228 );
nor \U$14463 ( \14806 , \14804 , \14805 );
xnor \U$14464 ( \14807 , \14806 , \8920 );
and \U$14465 ( \14808 , \14802 , \14807 );
and \U$14466 ( \14809 , \14798 , \14807 );
or \U$14467 ( \14810 , \14803 , \14808 , \14809 );
and \U$14468 ( \14811 , \14794 , \14810 );
and \U$14469 ( \14812 , \1412 , \8693 );
and \U$14470 ( \14813 , \1297 , \8691 );
nor \U$14471 ( \14814 , \14812 , \14813 );
xnor \U$14472 ( \14815 , \14814 , \8322 );
and \U$14473 ( \14816 , \1596 , \8131 );
and \U$14474 ( \14817 , \1588 , \8129 );
nor \U$14475 ( \14818 , \14816 , \14817 );
xnor \U$14476 ( \14819 , \14818 , \7813 );
and \U$14477 ( \14820 , \14815 , \14819 );
and \U$14478 ( \14821 , \1844 , \7564 );
and \U$14479 ( \14822 , \1839 , \7562 );
nor \U$14480 ( \14823 , \14821 , \14822 );
xnor \U$14481 ( \14824 , \14823 , \7315 );
and \U$14482 ( \14825 , \14819 , \14824 );
and \U$14483 ( \14826 , \14815 , \14824 );
or \U$14484 ( \14827 , \14820 , \14825 , \14826 );
and \U$14485 ( \14828 , \14810 , \14827 );
and \U$14486 ( \14829 , \14794 , \14827 );
or \U$14487 ( \14830 , \14811 , \14828 , \14829 );
and \U$14488 ( \14831 , \4266 , \4152 );
and \U$14489 ( \14832 , \4069 , \4150 );
nor \U$14490 ( \14833 , \14831 , \14832 );
xnor \U$14491 ( \14834 , \14833 , \4009 );
and \U$14492 ( \14835 , \4576 , \3829 );
and \U$14493 ( \14836 , \4568 , \3827 );
nor \U$14494 ( \14837 , \14835 , \14836 );
xnor \U$14495 ( \14838 , \14837 , \3583 );
and \U$14496 ( \14839 , \14834 , \14838 );
and \U$14497 ( \14840 , \5050 , \3434 );
and \U$14498 ( \14841 , \5045 , \3432 );
nor \U$14499 ( \14842 , \14840 , \14841 );
xnor \U$14500 ( \14843 , \14842 , \3247 );
and \U$14501 ( \14844 , \14838 , \14843 );
and \U$14502 ( \14845 , \14834 , \14843 );
or \U$14503 ( \14846 , \14839 , \14844 , \14845 );
and \U$14504 ( \14847 , \3061 , \5443 );
and \U$14505 ( \14848 , \2942 , \5441 );
nor \U$14506 ( \14849 , \14847 , \14848 );
xnor \U$14507 ( \14850 , \14849 , \5202 );
and \U$14508 ( \14851 , \3686 , \4977 );
and \U$14509 ( \14852 , \3478 , \4975 );
nor \U$14510 ( \14853 , \14851 , \14852 );
xnor \U$14511 ( \14854 , \14853 , \4789 );
and \U$14512 ( \14855 , \14850 , \14854 );
and \U$14513 ( \14856 , \3813 , \4603 );
and \U$14514 ( \14857 , \3808 , \4601 );
nor \U$14515 ( \14858 , \14856 , \14857 );
xnor \U$14516 ( \14859 , \14858 , \4371 );
and \U$14517 ( \14860 , \14854 , \14859 );
and \U$14518 ( \14861 , \14850 , \14859 );
or \U$14519 ( \14862 , \14855 , \14860 , \14861 );
and \U$14520 ( \14863 , \14846 , \14862 );
and \U$14521 ( \14864 , \5573 , \3121 );
and \U$14522 ( \14865 , \5314 , \3119 );
nor \U$14523 ( \14866 , \14864 , \14865 );
xnor \U$14524 ( \14867 , \14866 , \2916 );
and \U$14525 ( \14868 , \5954 , \2715 );
and \U$14526 ( \14869 , \5945 , \2713 );
nor \U$14527 ( \14870 , \14868 , \14869 );
xnor \U$14528 ( \14871 , \14870 , \2566 );
and \U$14529 ( \14872 , \14867 , \14871 );
and \U$14530 ( \14873 , \6499 , \2393 );
and \U$14531 ( \14874 , \6297 , \2391 );
nor \U$14532 ( \14875 , \14873 , \14874 );
xnor \U$14533 ( \14876 , \14875 , \2251 );
and \U$14534 ( \14877 , \14871 , \14876 );
and \U$14535 ( \14878 , \14867 , \14876 );
or \U$14536 ( \14879 , \14872 , \14877 , \14878 );
and \U$14537 ( \14880 , \14862 , \14879 );
and \U$14538 ( \14881 , \14846 , \14879 );
or \U$14539 ( \14882 , \14863 , \14880 , \14881 );
and \U$14540 ( \14883 , \14830 , \14882 );
and \U$14541 ( \14884 , \8778 , \1351 );
and \U$14542 ( \14885 , \8494 , \1349 );
nor \U$14543 ( \14886 , \14884 , \14885 );
xnor \U$14544 ( \14887 , \14886 , \1238 );
and \U$14545 ( \14888 , \9355 , \1157 );
and \U$14546 ( \14889 , \9347 , \1155 );
nor \U$14547 ( \14890 , \14888 , \14889 );
xnor \U$14548 ( \14891 , \14890 , \1021 );
and \U$14549 ( \14892 , \14887 , \14891 );
and \U$14550 ( \14893 , \9963 , \957 );
and \U$14551 ( \14894 , \9958 , \955 );
nor \U$14552 ( \14895 , \14893 , \14894 );
xnor \U$14553 ( \14896 , \14895 , \879 );
and \U$14554 ( \14897 , \14891 , \14896 );
and \U$14555 ( \14898 , \14887 , \14896 );
or \U$14556 ( \14899 , \14892 , \14897 , \14898 );
and \U$14557 ( \14900 , \6974 , \2097 );
and \U$14558 ( \14901 , \6802 , \2095 );
nor \U$14559 ( \14902 , \14900 , \14901 );
xnor \U$14560 ( \14903 , \14902 , \1960 );
and \U$14561 ( \14904 , \7924 , \1891 );
and \U$14562 ( \14905 , \7500 , \1889 );
nor \U$14563 ( \14906 , \14904 , \14905 );
xnor \U$14564 ( \14907 , \14906 , \1739 );
and \U$14565 ( \14908 , \14903 , \14907 );
and \U$14566 ( \14909 , \8175 , \1623 );
and \U$14567 ( \14910 , \8170 , \1621 );
nor \U$14568 ( \14911 , \14909 , \14910 );
xnor \U$14569 ( \14912 , \14911 , \1467 );
and \U$14570 ( \14913 , \14907 , \14912 );
and \U$14571 ( \14914 , \14903 , \14912 );
or \U$14572 ( \14915 , \14908 , \14913 , \14914 );
and \U$14573 ( \14916 , \14899 , \14915 );
xor \U$14574 ( \14917 , \14630 , \14634 );
xor \U$14575 ( \14918 , \14917 , \14637 );
and \U$14576 ( \14919 , \14915 , \14918 );
and \U$14577 ( \14920 , \14899 , \14918 );
or \U$14578 ( \14921 , \14916 , \14919 , \14920 );
and \U$14579 ( \14922 , \14882 , \14921 );
and \U$14580 ( \14923 , \14830 , \14921 );
or \U$14581 ( \14924 , \14883 , \14922 , \14923 );
xor \U$14582 ( \14925 , \14614 , \14618 );
xor \U$14583 ( \14926 , \14925 , \14623 );
xor \U$14584 ( \14927 , \14546 , \14550 );
xor \U$14585 ( \14928 , \14927 , \14555 );
and \U$14586 ( \14929 , \14926 , \14928 );
xor \U$14587 ( \14930 , \14645 , \14649 );
xor \U$14588 ( \14931 , \14930 , \14654 );
and \U$14589 ( \14932 , \14928 , \14931 );
and \U$14590 ( \14933 , \14926 , \14931 );
or \U$14591 ( \14934 , \14929 , \14932 , \14933 );
xor \U$14592 ( \14935 , \14513 , \14517 );
xor \U$14593 ( \14936 , \14935 , \14522 );
xor \U$14594 ( \14937 , \14529 , \14533 );
xor \U$14595 ( \14938 , \14937 , \14538 );
and \U$14596 ( \14939 , \14936 , \14938 );
xor \U$14597 ( \14940 , \14565 , \14569 );
xor \U$14598 ( \14941 , \14940 , \14574 );
and \U$14599 ( \14942 , \14938 , \14941 );
and \U$14600 ( \14943 , \14936 , \14941 );
or \U$14601 ( \14944 , \14939 , \14942 , \14943 );
and \U$14602 ( \14945 , \14934 , \14944 );
xor \U$14603 ( \14946 , \14581 , \14585 );
xor \U$14604 ( \14947 , \14946 , \14590 );
xor \U$14605 ( \14948 , \14598 , \14602 );
xor \U$14606 ( \14949 , \14948 , \349 );
and \U$14607 ( \14950 , \14947 , \14949 );
and \U$14608 ( \14951 , \14944 , \14950 );
and \U$14609 ( \14952 , \14934 , \14950 );
or \U$14610 ( \14953 , \14945 , \14951 , \14952 );
and \U$14611 ( \14954 , \14924 , \14953 );
xor \U$14612 ( \14955 , \14665 , \14667 );
xor \U$14613 ( \14956 , \14955 , \14670 );
xor \U$14614 ( \14957 , \14675 , \14677 );
xor \U$14615 ( \14958 , \14957 , \14680 );
and \U$14616 ( \14959 , \14956 , \14958 );
xor \U$14617 ( \14960 , \14686 , \14688 );
xor \U$14618 ( \14961 , \14960 , \14690 );
and \U$14619 ( \14962 , \14958 , \14961 );
and \U$14620 ( \14963 , \14956 , \14961 );
or \U$14621 ( \14964 , \14959 , \14962 , \14963 );
and \U$14622 ( \14965 , \14953 , \14964 );
and \U$14623 ( \14966 , \14924 , \14964 );
or \U$14624 ( \14967 , \14954 , \14965 , \14966 );
xor \U$14625 ( \14968 , \14525 , \14541 );
xor \U$14626 ( \14969 , \14968 , \14558 );
xor \U$14627 ( \14970 , \14577 , \14593 );
xor \U$14628 ( \14971 , \14970 , \14606 );
and \U$14629 ( \14972 , \14969 , \14971 );
xor \U$14630 ( \14973 , \14626 , \14640 );
xor \U$14631 ( \14974 , \14973 , \14657 );
and \U$14632 ( \14975 , \14971 , \14974 );
and \U$14633 ( \14976 , \14969 , \14974 );
or \U$14634 ( \14977 , \14972 , \14975 , \14976 );
xor \U$14635 ( \14978 , \14361 , \14377 );
xor \U$14636 ( \14979 , \14978 , \14394 );
and \U$14637 ( \14980 , \14977 , \14979 );
xor \U$14638 ( \14981 , \14712 , \14714 );
xor \U$14639 ( \14982 , \14981 , \14717 );
and \U$14640 ( \14983 , \14979 , \14982 );
and \U$14641 ( \14984 , \14977 , \14982 );
or \U$14642 ( \14985 , \14980 , \14983 , \14984 );
and \U$14643 ( \14986 , \14967 , \14985 );
xor \U$14644 ( \14987 , \14561 , \14609 );
xor \U$14645 ( \14988 , \14987 , \14660 );
xor \U$14646 ( \14989 , \14673 , \14683 );
xor \U$14647 ( \14990 , \14989 , \14693 );
and \U$14648 ( \14991 , \14988 , \14990 );
xor \U$14649 ( \14992 , \14699 , \14701 );
xor \U$14650 ( \14993 , \14992 , \14704 );
and \U$14651 ( \14994 , \14990 , \14993 );
and \U$14652 ( \14995 , \14988 , \14993 );
or \U$14653 ( \14996 , \14991 , \14994 , \14995 );
and \U$14654 ( \14997 , \14985 , \14996 );
and \U$14655 ( \14998 , \14967 , \14996 );
or \U$14656 ( \14999 , \14986 , \14997 , \14998 );
xor \U$14657 ( \15000 , \14663 , \14696 );
xor \U$14658 ( \15001 , \15000 , \14707 );
xor \U$14659 ( \15002 , \14720 , \14722 );
xor \U$14660 ( \15003 , \15002 , \14725 );
and \U$14661 ( \15004 , \15001 , \15003 );
xor \U$14662 ( \15005 , \14731 , \14733 );
and \U$14663 ( \15006 , \15003 , \15005 );
and \U$14664 ( \15007 , \15001 , \15005 );
or \U$14665 ( \15008 , \15004 , \15006 , \15007 );
and \U$14666 ( \15009 , \14999 , \15008 );
xor \U$14667 ( \15010 , \14739 , \14741 );
xor \U$14668 ( \15011 , \15010 , \14744 );
and \U$14669 ( \15012 , \15008 , \15011 );
and \U$14670 ( \15013 , \14999 , \15011 );
or \U$14671 ( \15014 , \15009 , \15012 , \15013 );
xor \U$14672 ( \15015 , \14737 , \14747 );
xor \U$14673 ( \15016 , \15015 , \14750 );
and \U$14674 ( \15017 , \15014 , \15016 );
xor \U$14675 ( \15018 , \14755 , \14757 );
and \U$14676 ( \15019 , \15016 , \15018 );
and \U$14677 ( \15020 , \15014 , \15018 );
or \U$14678 ( \15021 , \15017 , \15019 , \15020 );
and \U$14679 ( \15022 , \14778 , \15021 );
xor \U$14680 ( \15023 , \14778 , \15021 );
xor \U$14681 ( \15024 , \15014 , \15016 );
xor \U$14682 ( \15025 , \15024 , \15018 );
and \U$14683 ( \15026 , \2030 , \7564 );
and \U$14684 ( \15027 , \1844 , \7562 );
nor \U$14685 ( \15028 , \15026 , \15027 );
xnor \U$14686 ( \15029 , \15028 , \7315 );
and \U$14687 ( \15030 , \2438 , \7035 );
and \U$14688 ( \15031 , \2174 , \7033 );
nor \U$14689 ( \15032 , \15030 , \15031 );
xnor \U$14690 ( \15033 , \15032 , \6775 );
and \U$14691 ( \15034 , \15029 , \15033 );
and \U$14692 ( \15035 , \2637 , \6541 );
and \U$14693 ( \15036 , \2463 , \6539 );
nor \U$14694 ( \15037 , \15035 , \15036 );
xnor \U$14695 ( \15038 , \15037 , \6226 );
and \U$14696 ( \15039 , \15033 , \15038 );
and \U$14697 ( \15040 , \15029 , \15038 );
or \U$14698 ( \15041 , \15034 , \15039 , \15040 );
and \U$14699 ( \15042 , \1297 , \9230 );
and \U$14700 ( \15043 , \1181 , \9228 );
nor \U$14701 ( \15044 , \15042 , \15043 );
xnor \U$14702 ( \15045 , \15044 , \8920 );
and \U$14703 ( \15046 , \1588 , \8693 );
and \U$14704 ( \15047 , \1412 , \8691 );
nor \U$14705 ( \15048 , \15046 , \15047 );
xnor \U$14706 ( \15049 , \15048 , \8322 );
and \U$14707 ( \15050 , \15045 , \15049 );
and \U$14708 ( \15051 , \1839 , \8131 );
and \U$14709 ( \15052 , \1596 , \8129 );
nor \U$14710 ( \15053 , \15051 , \15052 );
xnor \U$14711 ( \15054 , \15053 , \7813 );
and \U$14712 ( \15055 , \15049 , \15054 );
and \U$14713 ( \15056 , \15045 , \15054 );
or \U$14714 ( \15057 , \15050 , \15055 , \15056 );
and \U$14715 ( \15058 , \15041 , \15057 );
and \U$14716 ( \15059 , \983 , \10611 );
and \U$14717 ( \15060 , \785 , \10608 );
nor \U$14718 ( \15061 , \15059 , \15060 );
xnor \U$14719 ( \15062 , \15061 , \9556 );
and \U$14720 ( \15063 , \1176 , \9798 );
and \U$14721 ( \15064 , \1071 , \9796 );
nor \U$14722 ( \15065 , \15063 , \15064 );
xnor \U$14723 ( \15066 , \15065 , \9559 );
and \U$14724 ( \15067 , \15062 , \15066 );
and \U$14725 ( \15068 , \15066 , \699 );
and \U$14726 ( \15069 , \15062 , \699 );
or \U$14727 ( \15070 , \15067 , \15068 , \15069 );
and \U$14728 ( \15071 , \15057 , \15070 );
and \U$14729 ( \15072 , \15041 , \15070 );
or \U$14730 ( \15073 , \15058 , \15071 , \15072 );
and \U$14731 ( \15074 , \6802 , \2393 );
and \U$14732 ( \15075 , \6499 , \2391 );
nor \U$14733 ( \15076 , \15074 , \15075 );
xnor \U$14734 ( \15077 , \15076 , \2251 );
and \U$14735 ( \15078 , \7500 , \2097 );
and \U$14736 ( \15079 , \6974 , \2095 );
nor \U$14737 ( \15080 , \15078 , \15079 );
xnor \U$14738 ( \15081 , \15080 , \1960 );
and \U$14739 ( \15082 , \15077 , \15081 );
and \U$14740 ( \15083 , \8170 , \1891 );
and \U$14741 ( \15084 , \7924 , \1889 );
nor \U$14742 ( \15085 , \15083 , \15084 );
xnor \U$14743 ( \15086 , \15085 , \1739 );
and \U$14744 ( \15087 , \15081 , \15086 );
and \U$14745 ( \15088 , \15077 , \15086 );
or \U$14746 ( \15089 , \15082 , \15087 , \15088 );
and \U$14747 ( \15090 , \8494 , \1623 );
and \U$14748 ( \15091 , \8175 , \1621 );
nor \U$14749 ( \15092 , \15090 , \15091 );
xnor \U$14750 ( \15093 , \15092 , \1467 );
and \U$14751 ( \15094 , \9347 , \1351 );
and \U$14752 ( \15095 , \8778 , \1349 );
nor \U$14753 ( \15096 , \15094 , \15095 );
xnor \U$14754 ( \15097 , \15096 , \1238 );
and \U$14755 ( \15098 , \15093 , \15097 );
and \U$14756 ( \15099 , \9958 , \1157 );
and \U$14757 ( \15100 , \9355 , \1155 );
nor \U$14758 ( \15101 , \15099 , \15100 );
xnor \U$14759 ( \15102 , \15101 , \1021 );
and \U$14760 ( \15103 , \15097 , \15102 );
and \U$14761 ( \15104 , \15093 , \15102 );
or \U$14762 ( \15105 , \15098 , \15103 , \15104 );
and \U$14763 ( \15106 , \15089 , \15105 );
and \U$14764 ( \15107 , \10764 , \793 );
and \U$14765 ( \15108 , \10144 , \791 );
nor \U$14766 ( \15109 , \15107 , \15108 );
xnor \U$14767 ( \15110 , \15109 , \699 );
and \U$14768 ( \15111 , \15105 , \15110 );
and \U$14769 ( \15112 , \15089 , \15110 );
or \U$14770 ( \15113 , \15106 , \15111 , \15112 );
and \U$14771 ( \15114 , \15073 , \15113 );
and \U$14772 ( \15115 , \4069 , \4603 );
and \U$14773 ( \15116 , \3813 , \4601 );
nor \U$14774 ( \15117 , \15115 , \15116 );
xnor \U$14775 ( \15118 , \15117 , \4371 );
and \U$14776 ( \15119 , \4568 , \4152 );
and \U$14777 ( \15120 , \4266 , \4150 );
nor \U$14778 ( \15121 , \15119 , \15120 );
xnor \U$14779 ( \15122 , \15121 , \4009 );
and \U$14780 ( \15123 , \15118 , \15122 );
and \U$14781 ( \15124 , \5045 , \3829 );
and \U$14782 ( \15125 , \4576 , \3827 );
nor \U$14783 ( \15126 , \15124 , \15125 );
xnor \U$14784 ( \15127 , \15126 , \3583 );
and \U$14785 ( \15128 , \15122 , \15127 );
and \U$14786 ( \15129 , \15118 , \15127 );
or \U$14787 ( \15130 , \15123 , \15128 , \15129 );
and \U$14788 ( \15131 , \2942 , \6032 );
and \U$14789 ( \15132 , \2804 , \6030 );
nor \U$14790 ( \15133 , \15131 , \15132 );
xnor \U$14791 ( \15134 , \15133 , \5692 );
and \U$14792 ( \15135 , \3478 , \5443 );
and \U$14793 ( \15136 , \3061 , \5441 );
nor \U$14794 ( \15137 , \15135 , \15136 );
xnor \U$14795 ( \15138 , \15137 , \5202 );
and \U$14796 ( \15139 , \15134 , \15138 );
and \U$14797 ( \15140 , \3808 , \4977 );
and \U$14798 ( \15141 , \3686 , \4975 );
nor \U$14799 ( \15142 , \15140 , \15141 );
xnor \U$14800 ( \15143 , \15142 , \4789 );
and \U$14801 ( \15144 , \15138 , \15143 );
and \U$14802 ( \15145 , \15134 , \15143 );
or \U$14803 ( \15146 , \15139 , \15144 , \15145 );
and \U$14804 ( \15147 , \15130 , \15146 );
and \U$14805 ( \15148 , \5314 , \3434 );
and \U$14806 ( \15149 , \5050 , \3432 );
nor \U$14807 ( \15150 , \15148 , \15149 );
xnor \U$14808 ( \15151 , \15150 , \3247 );
and \U$14809 ( \15152 , \5945 , \3121 );
and \U$14810 ( \15153 , \5573 , \3119 );
nor \U$14811 ( \15154 , \15152 , \15153 );
xnor \U$14812 ( \15155 , \15154 , \2916 );
and \U$14813 ( \15156 , \15151 , \15155 );
and \U$14814 ( \15157 , \6297 , \2715 );
and \U$14815 ( \15158 , \5954 , \2713 );
nor \U$14816 ( \15159 , \15157 , \15158 );
xnor \U$14817 ( \15160 , \15159 , \2566 );
and \U$14818 ( \15161 , \15155 , \15160 );
and \U$14819 ( \15162 , \15151 , \15160 );
or \U$14820 ( \15163 , \15156 , \15161 , \15162 );
and \U$14821 ( \15164 , \15146 , \15163 );
and \U$14822 ( \15165 , \15130 , \15163 );
or \U$14823 ( \15166 , \15147 , \15164 , \15165 );
and \U$14824 ( \15167 , \15113 , \15166 );
and \U$14825 ( \15168 , \15073 , \15166 );
or \U$14826 ( \15169 , \15114 , \15167 , \15168 );
xor \U$14827 ( \15170 , \14887 , \14891 );
xor \U$14828 ( \15171 , \15170 , \14896 );
xor \U$14829 ( \15172 , \14867 , \14871 );
xor \U$14830 ( \15173 , \15172 , \14876 );
and \U$14831 ( \15174 , \15171 , \15173 );
xor \U$14832 ( \15175 , \14903 , \14907 );
xor \U$14833 ( \15176 , \15175 , \14912 );
and \U$14834 ( \15177 , \15173 , \15176 );
and \U$14835 ( \15178 , \15171 , \15176 );
or \U$14836 ( \15179 , \15174 , \15177 , \15178 );
xor \U$14837 ( \15180 , \14834 , \14838 );
xor \U$14838 ( \15181 , \15180 , \14843 );
xor \U$14839 ( \15182 , \14850 , \14854 );
xor \U$14840 ( \15183 , \15182 , \14859 );
and \U$14841 ( \15184 , \15181 , \15183 );
xor \U$14842 ( \15185 , \14782 , \14786 );
xor \U$14843 ( \15186 , \15185 , \14791 );
and \U$14844 ( \15187 , \15183 , \15186 );
and \U$14845 ( \15188 , \15181 , \15186 );
or \U$14846 ( \15189 , \15184 , \15187 , \15188 );
and \U$14847 ( \15190 , \15179 , \15189 );
xor \U$14848 ( \15191 , \14798 , \14802 );
xor \U$14849 ( \15192 , \15191 , \14807 );
xor \U$14850 ( \15193 , \14815 , \14819 );
xor \U$14851 ( \15194 , \15193 , \14824 );
and \U$14852 ( \15195 , \15192 , \15194 );
and \U$14853 ( \15196 , \15189 , \15195 );
and \U$14854 ( \15197 , \15179 , \15195 );
or \U$14855 ( \15198 , \15190 , \15196 , \15197 );
and \U$14856 ( \15199 , \15169 , \15198 );
xor \U$14857 ( \15200 , \14926 , \14928 );
xor \U$14858 ( \15201 , \15200 , \14931 );
xor \U$14859 ( \15202 , \14936 , \14938 );
xor \U$14860 ( \15203 , \15202 , \14941 );
and \U$14861 ( \15204 , \15201 , \15203 );
xor \U$14862 ( \15205 , \14947 , \14949 );
and \U$14863 ( \15206 , \15203 , \15205 );
and \U$14864 ( \15207 , \15201 , \15205 );
or \U$14865 ( \15208 , \15204 , \15206 , \15207 );
and \U$14866 ( \15209 , \15198 , \15208 );
and \U$14867 ( \15210 , \15169 , \15208 );
or \U$14868 ( \15211 , \15199 , \15209 , \15210 );
xor \U$14869 ( \15212 , \14794 , \14810 );
xor \U$14870 ( \15213 , \15212 , \14827 );
xor \U$14871 ( \15214 , \14846 , \14862 );
xor \U$14872 ( \15215 , \15214 , \14879 );
and \U$14873 ( \15216 , \15213 , \15215 );
xor \U$14874 ( \15217 , \14899 , \14915 );
xor \U$14875 ( \15218 , \15217 , \14918 );
and \U$14876 ( \15219 , \15215 , \15218 );
and \U$14877 ( \15220 , \15213 , \15218 );
or \U$14878 ( \15221 , \15216 , \15219 , \15220 );
xor \U$14879 ( \15222 , \14969 , \14971 );
xor \U$14880 ( \15223 , \15222 , \14974 );
and \U$14881 ( \15224 , \15221 , \15223 );
xor \U$14882 ( \15225 , \14956 , \14958 );
xor \U$14883 ( \15226 , \15225 , \14961 );
and \U$14884 ( \15227 , \15223 , \15226 );
and \U$14885 ( \15228 , \15221 , \15226 );
or \U$14886 ( \15229 , \15224 , \15227 , \15228 );
and \U$14887 ( \15230 , \15211 , \15229 );
xor \U$14888 ( \15231 , \14988 , \14990 );
xor \U$14889 ( \15232 , \15231 , \14993 );
and \U$14890 ( \15233 , \15229 , \15232 );
and \U$14891 ( \15234 , \15211 , \15232 );
or \U$14892 ( \15235 , \15230 , \15233 , \15234 );
xor \U$14893 ( \15236 , \14967 , \14985 );
xor \U$14894 ( \15237 , \15236 , \14996 );
and \U$14895 ( \15238 , \15235 , \15237 );
xor \U$14896 ( \15239 , \15001 , \15003 );
xor \U$14897 ( \15240 , \15239 , \15005 );
and \U$14898 ( \15241 , \15237 , \15240 );
and \U$14899 ( \15242 , \15235 , \15240 );
or \U$14900 ( \15243 , \15238 , \15241 , \15242 );
xor \U$14901 ( \15244 , \14710 , \14728 );
xor \U$14902 ( \15245 , \15244 , \14734 );
and \U$14903 ( \15246 , \15243 , \15245 );
xor \U$14904 ( \15247 , \14999 , \15008 );
xor \U$14905 ( \15248 , \15247 , \15011 );
and \U$14906 ( \15249 , \15245 , \15248 );
and \U$14907 ( \15250 , \15243 , \15248 );
or \U$14908 ( \15251 , \15246 , \15249 , \15250 );
and \U$14909 ( \15252 , \15025 , \15251 );
xor \U$14910 ( \15253 , \15025 , \15251 );
xor \U$14911 ( \15254 , \15243 , \15245 );
xor \U$14912 ( \15255 , \15254 , \15248 );
xor \U$14913 ( \15256 , \15029 , \15033 );
xor \U$14914 ( \15257 , \15256 , \15038 );
xor \U$14915 ( \15258 , \15045 , \15049 );
xor \U$14916 ( \15259 , \15258 , \15054 );
and \U$14917 ( \15260 , \15257 , \15259 );
xor \U$14918 ( \15261 , \15062 , \15066 );
xor \U$14919 ( \15262 , \15261 , \699 );
and \U$14920 ( \15263 , \15259 , \15262 );
and \U$14921 ( \15264 , \15257 , \15262 );
or \U$14922 ( \15265 , \15260 , \15263 , \15264 );
nand \U$14923 ( \15266 , \10764 , \791 );
xnor \U$14924 ( \15267 , \15266 , \699 );
xor \U$14925 ( \15268 , \15077 , \15081 );
xor \U$14926 ( \15269 , \15268 , \15086 );
and \U$14927 ( \15270 , \15267 , \15269 );
xor \U$14928 ( \15271 , \15093 , \15097 );
xor \U$14929 ( \15272 , \15271 , \15102 );
and \U$14930 ( \15273 , \15269 , \15272 );
and \U$14931 ( \15274 , \15267 , \15272 );
or \U$14932 ( \15275 , \15270 , \15273 , \15274 );
and \U$14933 ( \15276 , \15265 , \15275 );
xor \U$14934 ( \15277 , \15118 , \15122 );
xor \U$14935 ( \15278 , \15277 , \15127 );
xor \U$14936 ( \15279 , \15134 , \15138 );
xor \U$14937 ( \15280 , \15279 , \15143 );
and \U$14938 ( \15281 , \15278 , \15280 );
xor \U$14939 ( \15282 , \15151 , \15155 );
xor \U$14940 ( \15283 , \15282 , \15160 );
and \U$14941 ( \15284 , \15280 , \15283 );
and \U$14942 ( \15285 , \15278 , \15283 );
or \U$14943 ( \15286 , \15281 , \15284 , \15285 );
and \U$14944 ( \15287 , \15275 , \15286 );
and \U$14945 ( \15288 , \15265 , \15286 );
or \U$14946 ( \15289 , \15276 , \15287 , \15288 );
and \U$14947 ( \15290 , \7924 , \2097 );
and \U$14948 ( \15291 , \7500 , \2095 );
nor \U$14949 ( \15292 , \15290 , \15291 );
xnor \U$14950 ( \15293 , \15292 , \1960 );
and \U$14951 ( \15294 , \8175 , \1891 );
and \U$14952 ( \15295 , \8170 , \1889 );
nor \U$14953 ( \15296 , \15294 , \15295 );
xnor \U$14954 ( \15297 , \15296 , \1739 );
and \U$14955 ( \15298 , \15293 , \15297 );
and \U$14956 ( \15299 , \8778 , \1623 );
and \U$14957 ( \15300 , \8494 , \1621 );
nor \U$14958 ( \15301 , \15299 , \15300 );
xnor \U$14959 ( \15302 , \15301 , \1467 );
and \U$14960 ( \15303 , \15297 , \15302 );
and \U$14961 ( \15304 , \15293 , \15302 );
or \U$14962 ( \15305 , \15298 , \15303 , \15304 );
and \U$14963 ( \15306 , \9355 , \1351 );
and \U$14964 ( \15307 , \9347 , \1349 );
nor \U$14965 ( \15308 , \15306 , \15307 );
xnor \U$14966 ( \15309 , \15308 , \1238 );
and \U$14967 ( \15310 , \9963 , \1157 );
and \U$14968 ( \15311 , \9958 , \1155 );
nor \U$14969 ( \15312 , \15310 , \15311 );
xnor \U$14970 ( \15313 , \15312 , \1021 );
and \U$14971 ( \15314 , \15309 , \15313 );
and \U$14972 ( \15315 , \10764 , \957 );
and \U$14973 ( \15316 , \10144 , \955 );
nor \U$14974 ( \15317 , \15315 , \15316 );
xnor \U$14975 ( \15318 , \15317 , \879 );
and \U$14976 ( \15319 , \15313 , \15318 );
and \U$14977 ( \15320 , \15309 , \15318 );
or \U$14978 ( \15321 , \15314 , \15319 , \15320 );
and \U$14979 ( \15322 , \15305 , \15321 );
and \U$14980 ( \15323 , \10144 , \957 );
and \U$14981 ( \15324 , \9963 , \955 );
nor \U$14982 ( \15325 , \15323 , \15324 );
xnor \U$14983 ( \15326 , \15325 , \879 );
and \U$14984 ( \15327 , \15321 , \15326 );
and \U$14985 ( \15328 , \15305 , \15326 );
or \U$14986 ( \15329 , \15322 , \15327 , \15328 );
and \U$14987 ( \15330 , \1071 , \10611 );
and \U$14988 ( \15331 , \983 , \10608 );
nor \U$14989 ( \15332 , \15330 , \15331 );
xnor \U$14990 ( \15333 , \15332 , \9556 );
and \U$14991 ( \15334 , \1181 , \9798 );
and \U$14992 ( \15335 , \1176 , \9796 );
nor \U$14993 ( \15336 , \15334 , \15335 );
xnor \U$14994 ( \15337 , \15336 , \9559 );
and \U$14995 ( \15338 , \15333 , \15337 );
and \U$14996 ( \15339 , \1412 , \9230 );
and \U$14997 ( \15340 , \1297 , \9228 );
nor \U$14998 ( \15341 , \15339 , \15340 );
xnor \U$14999 ( \15342 , \15341 , \8920 );
and \U$15000 ( \15343 , \15337 , \15342 );
and \U$15001 ( \15344 , \15333 , \15342 );
or \U$15002 ( \15345 , \15338 , \15343 , \15344 );
and \U$15003 ( \15346 , \1596 , \8693 );
and \U$15004 ( \15347 , \1588 , \8691 );
nor \U$15005 ( \15348 , \15346 , \15347 );
xnor \U$15006 ( \15349 , \15348 , \8322 );
and \U$15007 ( \15350 , \1844 , \8131 );
and \U$15008 ( \15351 , \1839 , \8129 );
nor \U$15009 ( \15352 , \15350 , \15351 );
xnor \U$15010 ( \15353 , \15352 , \7813 );
and \U$15011 ( \15354 , \15349 , \15353 );
and \U$15012 ( \15355 , \2174 , \7564 );
and \U$15013 ( \15356 , \2030 , \7562 );
nor \U$15014 ( \15357 , \15355 , \15356 );
xnor \U$15015 ( \15358 , \15357 , \7315 );
and \U$15016 ( \15359 , \15353 , \15358 );
and \U$15017 ( \15360 , \15349 , \15358 );
or \U$15018 ( \15361 , \15354 , \15359 , \15360 );
and \U$15019 ( \15362 , \15345 , \15361 );
and \U$15020 ( \15363 , \2463 , \7035 );
and \U$15021 ( \15364 , \2438 , \7033 );
nor \U$15022 ( \15365 , \15363 , \15364 );
xnor \U$15023 ( \15366 , \15365 , \6775 );
and \U$15024 ( \15367 , \2804 , \6541 );
and \U$15025 ( \15368 , \2637 , \6539 );
nor \U$15026 ( \15369 , \15367 , \15368 );
xnor \U$15027 ( \15370 , \15369 , \6226 );
and \U$15028 ( \15371 , \15366 , \15370 );
and \U$15029 ( \15372 , \3061 , \6032 );
and \U$15030 ( \15373 , \2942 , \6030 );
nor \U$15031 ( \15374 , \15372 , \15373 );
xnor \U$15032 ( \15375 , \15374 , \5692 );
and \U$15033 ( \15376 , \15370 , \15375 );
and \U$15034 ( \15377 , \15366 , \15375 );
or \U$15035 ( \15378 , \15371 , \15376 , \15377 );
and \U$15036 ( \15379 , \15361 , \15378 );
and \U$15037 ( \15380 , \15345 , \15378 );
or \U$15038 ( \15381 , \15362 , \15379 , \15380 );
and \U$15039 ( \15382 , \15329 , \15381 );
and \U$15040 ( \15383 , \4576 , \4152 );
and \U$15041 ( \15384 , \4568 , \4150 );
nor \U$15042 ( \15385 , \15383 , \15384 );
xnor \U$15043 ( \15386 , \15385 , \4009 );
and \U$15044 ( \15387 , \5050 , \3829 );
and \U$15045 ( \15388 , \5045 , \3827 );
nor \U$15046 ( \15389 , \15387 , \15388 );
xnor \U$15047 ( \15390 , \15389 , \3583 );
and \U$15048 ( \15391 , \15386 , \15390 );
and \U$15049 ( \15392 , \5573 , \3434 );
and \U$15050 ( \15393 , \5314 , \3432 );
nor \U$15051 ( \15394 , \15392 , \15393 );
xnor \U$15052 ( \15395 , \15394 , \3247 );
and \U$15053 ( \15396 , \15390 , \15395 );
and \U$15054 ( \15397 , \15386 , \15395 );
or \U$15055 ( \15398 , \15391 , \15396 , \15397 );
and \U$15056 ( \15399 , \5954 , \3121 );
and \U$15057 ( \15400 , \5945 , \3119 );
nor \U$15058 ( \15401 , \15399 , \15400 );
xnor \U$15059 ( \15402 , \15401 , \2916 );
and \U$15060 ( \15403 , \6499 , \2715 );
and \U$15061 ( \15404 , \6297 , \2713 );
nor \U$15062 ( \15405 , \15403 , \15404 );
xnor \U$15063 ( \15406 , \15405 , \2566 );
and \U$15064 ( \15407 , \15402 , \15406 );
and \U$15065 ( \15408 , \6974 , \2393 );
and \U$15066 ( \15409 , \6802 , \2391 );
nor \U$15067 ( \15410 , \15408 , \15409 );
xnor \U$15068 ( \15411 , \15410 , \2251 );
and \U$15069 ( \15412 , \15406 , \15411 );
and \U$15070 ( \15413 , \15402 , \15411 );
or \U$15071 ( \15414 , \15407 , \15412 , \15413 );
and \U$15072 ( \15415 , \15398 , \15414 );
and \U$15073 ( \15416 , \3686 , \5443 );
and \U$15074 ( \15417 , \3478 , \5441 );
nor \U$15075 ( \15418 , \15416 , \15417 );
xnor \U$15076 ( \15419 , \15418 , \5202 );
and \U$15077 ( \15420 , \3813 , \4977 );
and \U$15078 ( \15421 , \3808 , \4975 );
nor \U$15079 ( \15422 , \15420 , \15421 );
xnor \U$15080 ( \15423 , \15422 , \4789 );
and \U$15081 ( \15424 , \15419 , \15423 );
and \U$15082 ( \15425 , \4266 , \4603 );
and \U$15083 ( \15426 , \4069 , \4601 );
nor \U$15084 ( \15427 , \15425 , \15426 );
xnor \U$15085 ( \15428 , \15427 , \4371 );
and \U$15086 ( \15429 , \15423 , \15428 );
and \U$15087 ( \15430 , \15419 , \15428 );
or \U$15088 ( \15431 , \15424 , \15429 , \15430 );
and \U$15089 ( \15432 , \15414 , \15431 );
and \U$15090 ( \15433 , \15398 , \15431 );
or \U$15091 ( \15434 , \15415 , \15432 , \15433 );
and \U$15092 ( \15435 , \15381 , \15434 );
and \U$15093 ( \15436 , \15329 , \15434 );
or \U$15094 ( \15437 , \15382 , \15435 , \15436 );
and \U$15095 ( \15438 , \15289 , \15437 );
xor \U$15096 ( \15439 , \15171 , \15173 );
xor \U$15097 ( \15440 , \15439 , \15176 );
xor \U$15098 ( \15441 , \15181 , \15183 );
xor \U$15099 ( \15442 , \15441 , \15186 );
and \U$15100 ( \15443 , \15440 , \15442 );
xor \U$15101 ( \15444 , \15192 , \15194 );
and \U$15102 ( \15445 , \15442 , \15444 );
and \U$15103 ( \15446 , \15440 , \15444 );
or \U$15104 ( \15447 , \15443 , \15445 , \15446 );
and \U$15105 ( \15448 , \15437 , \15447 );
and \U$15106 ( \15449 , \15289 , \15447 );
or \U$15107 ( \15450 , \15438 , \15448 , \15449 );
xor \U$15108 ( \15451 , \15041 , \15057 );
xor \U$15109 ( \15452 , \15451 , \15070 );
xor \U$15110 ( \15453 , \15089 , \15105 );
xor \U$15111 ( \15454 , \15453 , \15110 );
and \U$15112 ( \15455 , \15452 , \15454 );
xor \U$15113 ( \15456 , \15130 , \15146 );
xor \U$15114 ( \15457 , \15456 , \15163 );
and \U$15115 ( \15458 , \15454 , \15457 );
and \U$15116 ( \15459 , \15452 , \15457 );
or \U$15117 ( \15460 , \15455 , \15458 , \15459 );
xor \U$15118 ( \15461 , \15213 , \15215 );
xor \U$15119 ( \15462 , \15461 , \15218 );
and \U$15120 ( \15463 , \15460 , \15462 );
xor \U$15121 ( \15464 , \15201 , \15203 );
xor \U$15122 ( \15465 , \15464 , \15205 );
and \U$15123 ( \15466 , \15462 , \15465 );
and \U$15124 ( \15467 , \15460 , \15465 );
or \U$15125 ( \15468 , \15463 , \15466 , \15467 );
and \U$15126 ( \15469 , \15450 , \15468 );
xor \U$15127 ( \15470 , \14934 , \14944 );
xor \U$15128 ( \15471 , \15470 , \14950 );
and \U$15129 ( \15472 , \15468 , \15471 );
and \U$15130 ( \15473 , \15450 , \15471 );
or \U$15131 ( \15474 , \15469 , \15472 , \15473 );
xor \U$15132 ( \15475 , \14830 , \14882 );
xor \U$15133 ( \15476 , \15475 , \14921 );
xor \U$15134 ( \15477 , \15169 , \15198 );
xor \U$15135 ( \15478 , \15477 , \15208 );
and \U$15136 ( \15479 , \15476 , \15478 );
xor \U$15137 ( \15480 , \15221 , \15223 );
xor \U$15138 ( \15481 , \15480 , \15226 );
and \U$15139 ( \15482 , \15478 , \15481 );
and \U$15140 ( \15483 , \15476 , \15481 );
or \U$15141 ( \15484 , \15479 , \15482 , \15483 );
and \U$15142 ( \15485 , \15474 , \15484 );
xor \U$15143 ( \15486 , \14977 , \14979 );
xor \U$15144 ( \15487 , \15486 , \14982 );
and \U$15145 ( \15488 , \15484 , \15487 );
and \U$15146 ( \15489 , \15474 , \15487 );
or \U$15147 ( \15490 , \15485 , \15488 , \15489 );
xor \U$15148 ( \15491 , \14924 , \14953 );
xor \U$15149 ( \15492 , \15491 , \14964 );
xor \U$15150 ( \15493 , \15211 , \15229 );
xor \U$15151 ( \15494 , \15493 , \15232 );
and \U$15152 ( \15495 , \15492 , \15494 );
and \U$15153 ( \15496 , \15490 , \15495 );
xor \U$15154 ( \15497 , \15235 , \15237 );
xor \U$15155 ( \15498 , \15497 , \15240 );
and \U$15156 ( \15499 , \15495 , \15498 );
and \U$15157 ( \15500 , \15490 , \15498 );
or \U$15158 ( \15501 , \15496 , \15499 , \15500 );
and \U$15159 ( \15502 , \15255 , \15501 );
xor \U$15160 ( \15503 , \15255 , \15501 );
xor \U$15161 ( \15504 , \15490 , \15495 );
xor \U$15162 ( \15505 , \15504 , \15498 );
and \U$15163 ( \15506 , \5945 , \3434 );
and \U$15164 ( \15507 , \5573 , \3432 );
nor \U$15165 ( \15508 , \15506 , \15507 );
xnor \U$15166 ( \15509 , \15508 , \3247 );
and \U$15167 ( \15510 , \6297 , \3121 );
and \U$15168 ( \15511 , \5954 , \3119 );
nor \U$15169 ( \15512 , \15510 , \15511 );
xnor \U$15170 ( \15513 , \15512 , \2916 );
and \U$15171 ( \15514 , \15509 , \15513 );
and \U$15172 ( \15515 , \6802 , \2715 );
and \U$15173 ( \15516 , \6499 , \2713 );
nor \U$15174 ( \15517 , \15515 , \15516 );
xnor \U$15175 ( \15518 , \15517 , \2566 );
and \U$15176 ( \15519 , \15513 , \15518 );
and \U$15177 ( \15520 , \15509 , \15518 );
or \U$15178 ( \15521 , \15514 , \15519 , \15520 );
and \U$15179 ( \15522 , \4568 , \4603 );
and \U$15180 ( \15523 , \4266 , \4601 );
nor \U$15181 ( \15524 , \15522 , \15523 );
xnor \U$15182 ( \15525 , \15524 , \4371 );
and \U$15183 ( \15526 , \5045 , \4152 );
and \U$15184 ( \15527 , \4576 , \4150 );
nor \U$15185 ( \15528 , \15526 , \15527 );
xnor \U$15186 ( \15529 , \15528 , \4009 );
and \U$15187 ( \15530 , \15525 , \15529 );
and \U$15188 ( \15531 , \5314 , \3829 );
and \U$15189 ( \15532 , \5050 , \3827 );
nor \U$15190 ( \15533 , \15531 , \15532 );
xnor \U$15191 ( \15534 , \15533 , \3583 );
and \U$15192 ( \15535 , \15529 , \15534 );
and \U$15193 ( \15536 , \15525 , \15534 );
or \U$15194 ( \15537 , \15530 , \15535 , \15536 );
and \U$15195 ( \15538 , \15521 , \15537 );
and \U$15196 ( \15539 , \3478 , \6032 );
and \U$15197 ( \15540 , \3061 , \6030 );
nor \U$15198 ( \15541 , \15539 , \15540 );
xnor \U$15199 ( \15542 , \15541 , \5692 );
and \U$15200 ( \15543 , \3808 , \5443 );
and \U$15201 ( \15544 , \3686 , \5441 );
nor \U$15202 ( \15545 , \15543 , \15544 );
xnor \U$15203 ( \15546 , \15545 , \5202 );
and \U$15204 ( \15547 , \15542 , \15546 );
and \U$15205 ( \15548 , \4069 , \4977 );
and \U$15206 ( \15549 , \3813 , \4975 );
nor \U$15207 ( \15550 , \15548 , \15549 );
xnor \U$15208 ( \15551 , \15550 , \4789 );
and \U$15209 ( \15552 , \15546 , \15551 );
and \U$15210 ( \15553 , \15542 , \15551 );
or \U$15211 ( \15554 , \15547 , \15552 , \15553 );
and \U$15212 ( \15555 , \15537 , \15554 );
and \U$15213 ( \15556 , \15521 , \15554 );
or \U$15214 ( \15557 , \15538 , \15555 , \15556 );
and \U$15215 ( \15558 , \1588 , \9230 );
and \U$15216 ( \15559 , \1412 , \9228 );
nor \U$15217 ( \15560 , \15558 , \15559 );
xnor \U$15218 ( \15561 , \15560 , \8920 );
and \U$15219 ( \15562 , \1839 , \8693 );
and \U$15220 ( \15563 , \1596 , \8691 );
nor \U$15221 ( \15564 , \15562 , \15563 );
xnor \U$15222 ( \15565 , \15564 , \8322 );
and \U$15223 ( \15566 , \15561 , \15565 );
and \U$15224 ( \15567 , \2030 , \8131 );
and \U$15225 ( \15568 , \1844 , \8129 );
nor \U$15226 ( \15569 , \15567 , \15568 );
xnor \U$15227 ( \15570 , \15569 , \7813 );
and \U$15228 ( \15571 , \15565 , \15570 );
and \U$15229 ( \15572 , \15561 , \15570 );
or \U$15230 ( \15573 , \15566 , \15571 , \15572 );
and \U$15231 ( \15574 , \1176 , \10611 );
and \U$15232 ( \15575 , \1071 , \10608 );
nor \U$15233 ( \15576 , \15574 , \15575 );
xnor \U$15234 ( \15577 , \15576 , \9556 );
and \U$15235 ( \15578 , \1297 , \9798 );
and \U$15236 ( \15579 , \1181 , \9796 );
nor \U$15237 ( \15580 , \15578 , \15579 );
xnor \U$15238 ( \15581 , \15580 , \9559 );
and \U$15239 ( \15582 , \15577 , \15581 );
and \U$15240 ( \15583 , \15581 , \879 );
and \U$15241 ( \15584 , \15577 , \879 );
or \U$15242 ( \15585 , \15582 , \15583 , \15584 );
and \U$15243 ( \15586 , \15573 , \15585 );
and \U$15244 ( \15587 , \2438 , \7564 );
and \U$15245 ( \15588 , \2174 , \7562 );
nor \U$15246 ( \15589 , \15587 , \15588 );
xnor \U$15247 ( \15590 , \15589 , \7315 );
and \U$15248 ( \15591 , \2637 , \7035 );
and \U$15249 ( \15592 , \2463 , \7033 );
nor \U$15250 ( \15593 , \15591 , \15592 );
xnor \U$15251 ( \15594 , \15593 , \6775 );
and \U$15252 ( \15595 , \15590 , \15594 );
and \U$15253 ( \15596 , \2942 , \6541 );
and \U$15254 ( \15597 , \2804 , \6539 );
nor \U$15255 ( \15598 , \15596 , \15597 );
xnor \U$15256 ( \15599 , \15598 , \6226 );
and \U$15257 ( \15600 , \15594 , \15599 );
and \U$15258 ( \15601 , \15590 , \15599 );
or \U$15259 ( \15602 , \15595 , \15600 , \15601 );
and \U$15260 ( \15603 , \15585 , \15602 );
and \U$15261 ( \15604 , \15573 , \15602 );
or \U$15262 ( \15605 , \15586 , \15603 , \15604 );
and \U$15263 ( \15606 , \15557 , \15605 );
and \U$15264 ( \15607 , \7500 , \2393 );
and \U$15265 ( \15608 , \6974 , \2391 );
nor \U$15266 ( \15609 , \15607 , \15608 );
xnor \U$15267 ( \15610 , \15609 , \2251 );
and \U$15268 ( \15611 , \8170 , \2097 );
and \U$15269 ( \15612 , \7924 , \2095 );
nor \U$15270 ( \15613 , \15611 , \15612 );
xnor \U$15271 ( \15614 , \15613 , \1960 );
and \U$15272 ( \15615 , \15610 , \15614 );
and \U$15273 ( \15616 , \8494 , \1891 );
and \U$15274 ( \15617 , \8175 , \1889 );
nor \U$15275 ( \15618 , \15616 , \15617 );
xnor \U$15276 ( \15619 , \15618 , \1739 );
and \U$15277 ( \15620 , \15614 , \15619 );
and \U$15278 ( \15621 , \15610 , \15619 );
or \U$15279 ( \15622 , \15615 , \15620 , \15621 );
and \U$15280 ( \15623 , \9347 , \1623 );
and \U$15281 ( \15624 , \8778 , \1621 );
nor \U$15282 ( \15625 , \15623 , \15624 );
xnor \U$15283 ( \15626 , \15625 , \1467 );
and \U$15284 ( \15627 , \9958 , \1351 );
and \U$15285 ( \15628 , \9355 , \1349 );
nor \U$15286 ( \15629 , \15627 , \15628 );
xnor \U$15287 ( \15630 , \15629 , \1238 );
and \U$15288 ( \15631 , \15626 , \15630 );
and \U$15289 ( \15632 , \10144 , \1157 );
and \U$15290 ( \15633 , \9963 , \1155 );
nor \U$15291 ( \15634 , \15632 , \15633 );
xnor \U$15292 ( \15635 , \15634 , \1021 );
and \U$15293 ( \15636 , \15630 , \15635 );
and \U$15294 ( \15637 , \15626 , \15635 );
or \U$15295 ( \15638 , \15631 , \15636 , \15637 );
and \U$15296 ( \15639 , \15622 , \15638 );
xor \U$15297 ( \15640 , \15309 , \15313 );
xor \U$15298 ( \15641 , \15640 , \15318 );
and \U$15299 ( \15642 , \15638 , \15641 );
and \U$15300 ( \15643 , \15622 , \15641 );
or \U$15301 ( \15644 , \15639 , \15642 , \15643 );
and \U$15302 ( \15645 , \15605 , \15644 );
and \U$15303 ( \15646 , \15557 , \15644 );
or \U$15304 ( \15647 , \15606 , \15645 , \15646 );
xor \U$15305 ( \15648 , \15293 , \15297 );
xor \U$15306 ( \15649 , \15648 , \15302 );
xor \U$15307 ( \15650 , \15386 , \15390 );
xor \U$15308 ( \15651 , \15650 , \15395 );
and \U$15309 ( \15652 , \15649 , \15651 );
xor \U$15310 ( \15653 , \15402 , \15406 );
xor \U$15311 ( \15654 , \15653 , \15411 );
and \U$15312 ( \15655 , \15651 , \15654 );
and \U$15313 ( \15656 , \15649 , \15654 );
or \U$15314 ( \15657 , \15652 , \15655 , \15656 );
xor \U$15315 ( \15658 , \15349 , \15353 );
xor \U$15316 ( \15659 , \15658 , \15358 );
xor \U$15317 ( \15660 , \15419 , \15423 );
xor \U$15318 ( \15661 , \15660 , \15428 );
and \U$15319 ( \15662 , \15659 , \15661 );
xor \U$15320 ( \15663 , \15366 , \15370 );
xor \U$15321 ( \15664 , \15663 , \15375 );
and \U$15322 ( \15665 , \15661 , \15664 );
and \U$15323 ( \15666 , \15659 , \15664 );
or \U$15324 ( \15667 , \15662 , \15665 , \15666 );
and \U$15325 ( \15668 , \15657 , \15667 );
xor \U$15326 ( \15669 , \15257 , \15259 );
xor \U$15327 ( \15670 , \15669 , \15262 );
and \U$15328 ( \15671 , \15667 , \15670 );
and \U$15329 ( \15672 , \15657 , \15670 );
or \U$15330 ( \15673 , \15668 , \15671 , \15672 );
and \U$15331 ( \15674 , \15647 , \15673 );
xor \U$15332 ( \15675 , \15305 , \15321 );
xor \U$15333 ( \15676 , \15675 , \15326 );
xor \U$15334 ( \15677 , \15267 , \15269 );
xor \U$15335 ( \15678 , \15677 , \15272 );
and \U$15336 ( \15679 , \15676 , \15678 );
xor \U$15337 ( \15680 , \15278 , \15280 );
xor \U$15338 ( \15681 , \15680 , \15283 );
and \U$15339 ( \15682 , \15678 , \15681 );
and \U$15340 ( \15683 , \15676 , \15681 );
or \U$15341 ( \15684 , \15679 , \15682 , \15683 );
and \U$15342 ( \15685 , \15673 , \15684 );
and \U$15343 ( \15686 , \15647 , \15684 );
or \U$15344 ( \15687 , \15674 , \15685 , \15686 );
xor \U$15345 ( \15688 , \15265 , \15275 );
xor \U$15346 ( \15689 , \15688 , \15286 );
xor \U$15347 ( \15690 , \15452 , \15454 );
xor \U$15348 ( \15691 , \15690 , \15457 );
and \U$15349 ( \15692 , \15689 , \15691 );
xor \U$15350 ( \15693 , \15440 , \15442 );
xor \U$15351 ( \15694 , \15693 , \15444 );
and \U$15352 ( \15695 , \15691 , \15694 );
and \U$15353 ( \15696 , \15689 , \15694 );
or \U$15354 ( \15697 , \15692 , \15695 , \15696 );
and \U$15355 ( \15698 , \15687 , \15697 );
xor \U$15356 ( \15699 , \15179 , \15189 );
xor \U$15357 ( \15700 , \15699 , \15195 );
and \U$15358 ( \15701 , \15697 , \15700 );
and \U$15359 ( \15702 , \15687 , \15700 );
or \U$15360 ( \15703 , \15698 , \15701 , \15702 );
xor \U$15361 ( \15704 , \15073 , \15113 );
xor \U$15362 ( \15705 , \15704 , \15166 );
xor \U$15363 ( \15706 , \15289 , \15437 );
xor \U$15364 ( \15707 , \15706 , \15447 );
and \U$15365 ( \15708 , \15705 , \15707 );
xor \U$15366 ( \15709 , \15460 , \15462 );
xor \U$15367 ( \15710 , \15709 , \15465 );
and \U$15368 ( \15711 , \15707 , \15710 );
and \U$15369 ( \15712 , \15705 , \15710 );
or \U$15370 ( \15713 , \15708 , \15711 , \15712 );
and \U$15371 ( \15714 , \15703 , \15713 );
xor \U$15372 ( \15715 , \15476 , \15478 );
xor \U$15373 ( \15716 , \15715 , \15481 );
and \U$15374 ( \15717 , \15713 , \15716 );
and \U$15375 ( \15718 , \15703 , \15716 );
or \U$15376 ( \15719 , \15714 , \15717 , \15718 );
xor \U$15377 ( \15720 , \15474 , \15484 );
xor \U$15378 ( \15721 , \15720 , \15487 );
and \U$15379 ( \15722 , \15719 , \15721 );
xor \U$15380 ( \15723 , \15492 , \15494 );
and \U$15381 ( \15724 , \15721 , \15723 );
and \U$15382 ( \15725 , \15719 , \15723 );
or \U$15383 ( \15726 , \15722 , \15724 , \15725 );
and \U$15384 ( \15727 , \15505 , \15726 );
xor \U$15385 ( \15728 , \15505 , \15726 );
xor \U$15386 ( \15729 , \15719 , \15721 );
xor \U$15387 ( \15730 , \15729 , \15723 );
and \U$15388 ( \15731 , \3813 , \5443 );
and \U$15389 ( \15732 , \3808 , \5441 );
nor \U$15390 ( \15733 , \15731 , \15732 );
xnor \U$15391 ( \15734 , \15733 , \5202 );
and \U$15392 ( \15735 , \4266 , \4977 );
and \U$15393 ( \15736 , \4069 , \4975 );
nor \U$15394 ( \15737 , \15735 , \15736 );
xnor \U$15395 ( \15738 , \15737 , \4789 );
and \U$15396 ( \15739 , \15734 , \15738 );
and \U$15397 ( \15740 , \4576 , \4603 );
and \U$15398 ( \15741 , \4568 , \4601 );
nor \U$15399 ( \15742 , \15740 , \15741 );
xnor \U$15400 ( \15743 , \15742 , \4371 );
and \U$15401 ( \15744 , \15738 , \15743 );
and \U$15402 ( \15745 , \15734 , \15743 );
or \U$15403 ( \15746 , \15739 , \15744 , \15745 );
and \U$15404 ( \15747 , \5050 , \4152 );
and \U$15405 ( \15748 , \5045 , \4150 );
nor \U$15406 ( \15749 , \15747 , \15748 );
xnor \U$15407 ( \15750 , \15749 , \4009 );
and \U$15408 ( \15751 , \5573 , \3829 );
and \U$15409 ( \15752 , \5314 , \3827 );
nor \U$15410 ( \15753 , \15751 , \15752 );
xnor \U$15411 ( \15754 , \15753 , \3583 );
and \U$15412 ( \15755 , \15750 , \15754 );
and \U$15413 ( \15756 , \5954 , \3434 );
and \U$15414 ( \15757 , \5945 , \3432 );
nor \U$15415 ( \15758 , \15756 , \15757 );
xnor \U$15416 ( \15759 , \15758 , \3247 );
and \U$15417 ( \15760 , \15754 , \15759 );
and \U$15418 ( \15761 , \15750 , \15759 );
or \U$15419 ( \15762 , \15755 , \15760 , \15761 );
and \U$15420 ( \15763 , \15746 , \15762 );
and \U$15421 ( \15764 , \6499 , \3121 );
and \U$15422 ( \15765 , \6297 , \3119 );
nor \U$15423 ( \15766 , \15764 , \15765 );
xnor \U$15424 ( \15767 , \15766 , \2916 );
and \U$15425 ( \15768 , \6974 , \2715 );
and \U$15426 ( \15769 , \6802 , \2713 );
nor \U$15427 ( \15770 , \15768 , \15769 );
xnor \U$15428 ( \15771 , \15770 , \2566 );
and \U$15429 ( \15772 , \15767 , \15771 );
and \U$15430 ( \15773 , \7924 , \2393 );
and \U$15431 ( \15774 , \7500 , \2391 );
nor \U$15432 ( \15775 , \15773 , \15774 );
xnor \U$15433 ( \15776 , \15775 , \2251 );
and \U$15434 ( \15777 , \15771 , \15776 );
and \U$15435 ( \15778 , \15767 , \15776 );
or \U$15436 ( \15779 , \15772 , \15777 , \15778 );
and \U$15437 ( \15780 , \15762 , \15779 );
and \U$15438 ( \15781 , \15746 , \15779 );
or \U$15439 ( \15782 , \15763 , \15780 , \15781 );
and \U$15440 ( \15783 , \1844 , \8693 );
and \U$15441 ( \15784 , \1839 , \8691 );
nor \U$15442 ( \15785 , \15783 , \15784 );
xnor \U$15443 ( \15786 , \15785 , \8322 );
and \U$15444 ( \15787 , \2174 , \8131 );
and \U$15445 ( \15788 , \2030 , \8129 );
nor \U$15446 ( \15789 , \15787 , \15788 );
xnor \U$15447 ( \15790 , \15789 , \7813 );
and \U$15448 ( \15791 , \15786 , \15790 );
and \U$15449 ( \15792 , \2463 , \7564 );
and \U$15450 ( \15793 , \2438 , \7562 );
nor \U$15451 ( \15794 , \15792 , \15793 );
xnor \U$15452 ( \15795 , \15794 , \7315 );
and \U$15453 ( \15796 , \15790 , \15795 );
and \U$15454 ( \15797 , \15786 , \15795 );
or \U$15455 ( \15798 , \15791 , \15796 , \15797 );
and \U$15456 ( \15799 , \2804 , \7035 );
and \U$15457 ( \15800 , \2637 , \7033 );
nor \U$15458 ( \15801 , \15799 , \15800 );
xnor \U$15459 ( \15802 , \15801 , \6775 );
and \U$15460 ( \15803 , \3061 , \6541 );
and \U$15461 ( \15804 , \2942 , \6539 );
nor \U$15462 ( \15805 , \15803 , \15804 );
xnor \U$15463 ( \15806 , \15805 , \6226 );
and \U$15464 ( \15807 , \15802 , \15806 );
and \U$15465 ( \15808 , \3686 , \6032 );
and \U$15466 ( \15809 , \3478 , \6030 );
nor \U$15467 ( \15810 , \15808 , \15809 );
xnor \U$15468 ( \15811 , \15810 , \5692 );
and \U$15469 ( \15812 , \15806 , \15811 );
and \U$15470 ( \15813 , \15802 , \15811 );
or \U$15471 ( \15814 , \15807 , \15812 , \15813 );
and \U$15472 ( \15815 , \15798 , \15814 );
and \U$15473 ( \15816 , \1181 , \10611 );
and \U$15474 ( \15817 , \1176 , \10608 );
nor \U$15475 ( \15818 , \15816 , \15817 );
xnor \U$15476 ( \15819 , \15818 , \9556 );
and \U$15477 ( \15820 , \1412 , \9798 );
and \U$15478 ( \15821 , \1297 , \9796 );
nor \U$15479 ( \15822 , \15820 , \15821 );
xnor \U$15480 ( \15823 , \15822 , \9559 );
and \U$15481 ( \15824 , \15819 , \15823 );
and \U$15482 ( \15825 , \1596 , \9230 );
and \U$15483 ( \15826 , \1588 , \9228 );
nor \U$15484 ( \15827 , \15825 , \15826 );
xnor \U$15485 ( \15828 , \15827 , \8920 );
and \U$15486 ( \15829 , \15823 , \15828 );
and \U$15487 ( \15830 , \15819 , \15828 );
or \U$15488 ( \15831 , \15824 , \15829 , \15830 );
and \U$15489 ( \15832 , \15814 , \15831 );
and \U$15490 ( \15833 , \15798 , \15831 );
or \U$15491 ( \15834 , \15815 , \15832 , \15833 );
and \U$15492 ( \15835 , \15782 , \15834 );
and \U$15493 ( \15836 , \8175 , \2097 );
and \U$15494 ( \15837 , \8170 , \2095 );
nor \U$15495 ( \15838 , \15836 , \15837 );
xnor \U$15496 ( \15839 , \15838 , \1960 );
and \U$15497 ( \15840 , \8778 , \1891 );
and \U$15498 ( \15841 , \8494 , \1889 );
nor \U$15499 ( \15842 , \15840 , \15841 );
xnor \U$15500 ( \15843 , \15842 , \1739 );
and \U$15501 ( \15844 , \15839 , \15843 );
and \U$15502 ( \15845 , \9355 , \1623 );
and \U$15503 ( \15846 , \9347 , \1621 );
nor \U$15504 ( \15847 , \15845 , \15846 );
xnor \U$15505 ( \15848 , \15847 , \1467 );
and \U$15506 ( \15849 , \15843 , \15848 );
and \U$15507 ( \15850 , \15839 , \15848 );
or \U$15508 ( \15851 , \15844 , \15849 , \15850 );
nand \U$15509 ( \15852 , \10764 , \955 );
xnor \U$15510 ( \15853 , \15852 , \879 );
and \U$15511 ( \15854 , \15851 , \15853 );
xor \U$15512 ( \15855 , \15626 , \15630 );
xor \U$15513 ( \15856 , \15855 , \15635 );
and \U$15514 ( \15857 , \15853 , \15856 );
and \U$15515 ( \15858 , \15851 , \15856 );
or \U$15516 ( \15859 , \15854 , \15857 , \15858 );
and \U$15517 ( \15860 , \15834 , \15859 );
and \U$15518 ( \15861 , \15782 , \15859 );
or \U$15519 ( \15862 , \15835 , \15860 , \15861 );
xor \U$15520 ( \15863 , \15509 , \15513 );
xor \U$15521 ( \15864 , \15863 , \15518 );
xor \U$15522 ( \15865 , \15610 , \15614 );
xor \U$15523 ( \15866 , \15865 , \15619 );
and \U$15524 ( \15867 , \15864 , \15866 );
xor \U$15525 ( \15868 , \15525 , \15529 );
xor \U$15526 ( \15869 , \15868 , \15534 );
and \U$15527 ( \15870 , \15866 , \15869 );
and \U$15528 ( \15871 , \15864 , \15869 );
or \U$15529 ( \15872 , \15867 , \15870 , \15871 );
xor \U$15530 ( \15873 , \15561 , \15565 );
xor \U$15531 ( \15874 , \15873 , \15570 );
xor \U$15532 ( \15875 , \15542 , \15546 );
xor \U$15533 ( \15876 , \15875 , \15551 );
and \U$15534 ( \15877 , \15874 , \15876 );
xor \U$15535 ( \15878 , \15590 , \15594 );
xor \U$15536 ( \15879 , \15878 , \15599 );
and \U$15537 ( \15880 , \15876 , \15879 );
and \U$15538 ( \15881 , \15874 , \15879 );
or \U$15539 ( \15882 , \15877 , \15880 , \15881 );
and \U$15540 ( \15883 , \15872 , \15882 );
xor \U$15541 ( \15884 , \15333 , \15337 );
xor \U$15542 ( \15885 , \15884 , \15342 );
and \U$15543 ( \15886 , \15882 , \15885 );
and \U$15544 ( \15887 , \15872 , \15885 );
or \U$15545 ( \15888 , \15883 , \15886 , \15887 );
and \U$15546 ( \15889 , \15862 , \15888 );
xor \U$15547 ( \15890 , \15649 , \15651 );
xor \U$15548 ( \15891 , \15890 , \15654 );
xor \U$15549 ( \15892 , \15659 , \15661 );
xor \U$15550 ( \15893 , \15892 , \15664 );
and \U$15551 ( \15894 , \15891 , \15893 );
xor \U$15552 ( \15895 , \15622 , \15638 );
xor \U$15553 ( \15896 , \15895 , \15641 );
and \U$15554 ( \15897 , \15893 , \15896 );
and \U$15555 ( \15898 , \15891 , \15896 );
or \U$15556 ( \15899 , \15894 , \15897 , \15898 );
and \U$15557 ( \15900 , \15888 , \15899 );
and \U$15558 ( \15901 , \15862 , \15899 );
or \U$15559 ( \15902 , \15889 , \15900 , \15901 );
xor \U$15560 ( \15903 , \15345 , \15361 );
xor \U$15561 ( \15904 , \15903 , \15378 );
xor \U$15562 ( \15905 , \15398 , \15414 );
xor \U$15563 ( \15906 , \15905 , \15431 );
and \U$15564 ( \15907 , \15904 , \15906 );
xor \U$15565 ( \15908 , \15676 , \15678 );
xor \U$15566 ( \15909 , \15908 , \15681 );
and \U$15567 ( \15910 , \15906 , \15909 );
and \U$15568 ( \15911 , \15904 , \15909 );
or \U$15569 ( \15912 , \15907 , \15910 , \15911 );
and \U$15570 ( \15913 , \15902 , \15912 );
xor \U$15571 ( \15914 , \15557 , \15605 );
xor \U$15572 ( \15915 , \15914 , \15644 );
xor \U$15573 ( \15916 , \15657 , \15667 );
xor \U$15574 ( \15917 , \15916 , \15670 );
and \U$15575 ( \15918 , \15915 , \15917 );
and \U$15576 ( \15919 , \15912 , \15918 );
and \U$15577 ( \15920 , \15902 , \15918 );
or \U$15578 ( \15921 , \15913 , \15919 , \15920 );
xor \U$15579 ( \15922 , \15329 , \15381 );
xor \U$15580 ( \15923 , \15922 , \15434 );
xor \U$15581 ( \15924 , \15647 , \15673 );
xor \U$15582 ( \15925 , \15924 , \15684 );
and \U$15583 ( \15926 , \15923 , \15925 );
xor \U$15584 ( \15927 , \15689 , \15691 );
xor \U$15585 ( \15928 , \15927 , \15694 );
and \U$15586 ( \15929 , \15925 , \15928 );
and \U$15587 ( \15930 , \15923 , \15928 );
or \U$15588 ( \15931 , \15926 , \15929 , \15930 );
and \U$15589 ( \15932 , \15921 , \15931 );
xor \U$15590 ( \15933 , \15705 , \15707 );
xor \U$15591 ( \15934 , \15933 , \15710 );
and \U$15592 ( \15935 , \15931 , \15934 );
and \U$15593 ( \15936 , \15921 , \15934 );
or \U$15594 ( \15937 , \15932 , \15935 , \15936 );
xor \U$15595 ( \15938 , \15450 , \15468 );
xor \U$15596 ( \15939 , \15938 , \15471 );
and \U$15597 ( \15940 , \15937 , \15939 );
xor \U$15598 ( \15941 , \15703 , \15713 );
xor \U$15599 ( \15942 , \15941 , \15716 );
and \U$15600 ( \15943 , \15939 , \15942 );
and \U$15601 ( \15944 , \15937 , \15942 );
or \U$15602 ( \15945 , \15940 , \15943 , \15944 );
and \U$15603 ( \15946 , \15730 , \15945 );
xor \U$15604 ( \15947 , \15730 , \15945 );
xor \U$15605 ( \15948 , \15937 , \15939 );
xor \U$15606 ( \15949 , \15948 , \15942 );
and \U$15607 ( \15950 , \1297 , \10611 );
and \U$15608 ( \15951 , \1181 , \10608 );
nor \U$15609 ( \15952 , \15950 , \15951 );
xnor \U$15610 ( \15953 , \15952 , \9556 );
and \U$15611 ( \15954 , \1588 , \9798 );
and \U$15612 ( \15955 , \1412 , \9796 );
nor \U$15613 ( \15956 , \15954 , \15955 );
xnor \U$15614 ( \15957 , \15956 , \9559 );
and \U$15615 ( \15958 , \15953 , \15957 );
and \U$15616 ( \15959 , \15957 , \1021 );
and \U$15617 ( \15960 , \15953 , \1021 );
or \U$15618 ( \15961 , \15958 , \15959 , \15960 );
and \U$15619 ( \15962 , \2637 , \7564 );
and \U$15620 ( \15963 , \2463 , \7562 );
nor \U$15621 ( \15964 , \15962 , \15963 );
xnor \U$15622 ( \15965 , \15964 , \7315 );
and \U$15623 ( \15966 , \2942 , \7035 );
and \U$15624 ( \15967 , \2804 , \7033 );
nor \U$15625 ( \15968 , \15966 , \15967 );
xnor \U$15626 ( \15969 , \15968 , \6775 );
and \U$15627 ( \15970 , \15965 , \15969 );
and \U$15628 ( \15971 , \3478 , \6541 );
and \U$15629 ( \15972 , \3061 , \6539 );
nor \U$15630 ( \15973 , \15971 , \15972 );
xnor \U$15631 ( \15974 , \15973 , \6226 );
and \U$15632 ( \15975 , \15969 , \15974 );
and \U$15633 ( \15976 , \15965 , \15974 );
or \U$15634 ( \15977 , \15970 , \15975 , \15976 );
and \U$15635 ( \15978 , \15961 , \15977 );
and \U$15636 ( \15979 , \1839 , \9230 );
and \U$15637 ( \15980 , \1596 , \9228 );
nor \U$15638 ( \15981 , \15979 , \15980 );
xnor \U$15639 ( \15982 , \15981 , \8920 );
and \U$15640 ( \15983 , \2030 , \8693 );
and \U$15641 ( \15984 , \1844 , \8691 );
nor \U$15642 ( \15985 , \15983 , \15984 );
xnor \U$15643 ( \15986 , \15985 , \8322 );
and \U$15644 ( \15987 , \15982 , \15986 );
and \U$15645 ( \15988 , \2438 , \8131 );
and \U$15646 ( \15989 , \2174 , \8129 );
nor \U$15647 ( \15990 , \15988 , \15989 );
xnor \U$15648 ( \15991 , \15990 , \7813 );
and \U$15649 ( \15992 , \15986 , \15991 );
and \U$15650 ( \15993 , \15982 , \15991 );
or \U$15651 ( \15994 , \15987 , \15992 , \15993 );
and \U$15652 ( \15995 , \15977 , \15994 );
and \U$15653 ( \15996 , \15961 , \15994 );
or \U$15654 ( \15997 , \15978 , \15995 , \15996 );
and \U$15655 ( \15998 , \3808 , \6032 );
and \U$15656 ( \15999 , \3686 , \6030 );
nor \U$15657 ( \16000 , \15998 , \15999 );
xnor \U$15658 ( \16001 , \16000 , \5692 );
and \U$15659 ( \16002 , \4069 , \5443 );
and \U$15660 ( \16003 , \3813 , \5441 );
nor \U$15661 ( \16004 , \16002 , \16003 );
xnor \U$15662 ( \16005 , \16004 , \5202 );
and \U$15663 ( \16006 , \16001 , \16005 );
and \U$15664 ( \16007 , \4568 , \4977 );
and \U$15665 ( \16008 , \4266 , \4975 );
nor \U$15666 ( \16009 , \16007 , \16008 );
xnor \U$15667 ( \16010 , \16009 , \4789 );
and \U$15668 ( \16011 , \16005 , \16010 );
and \U$15669 ( \16012 , \16001 , \16010 );
or \U$15670 ( \16013 , \16006 , \16011 , \16012 );
and \U$15671 ( \16014 , \5045 , \4603 );
and \U$15672 ( \16015 , \4576 , \4601 );
nor \U$15673 ( \16016 , \16014 , \16015 );
xnor \U$15674 ( \16017 , \16016 , \4371 );
and \U$15675 ( \16018 , \5314 , \4152 );
and \U$15676 ( \16019 , \5050 , \4150 );
nor \U$15677 ( \16020 , \16018 , \16019 );
xnor \U$15678 ( \16021 , \16020 , \4009 );
and \U$15679 ( \16022 , \16017 , \16021 );
and \U$15680 ( \16023 , \5945 , \3829 );
and \U$15681 ( \16024 , \5573 , \3827 );
nor \U$15682 ( \16025 , \16023 , \16024 );
xnor \U$15683 ( \16026 , \16025 , \3583 );
and \U$15684 ( \16027 , \16021 , \16026 );
and \U$15685 ( \16028 , \16017 , \16026 );
or \U$15686 ( \16029 , \16022 , \16027 , \16028 );
and \U$15687 ( \16030 , \16013 , \16029 );
and \U$15688 ( \16031 , \6297 , \3434 );
and \U$15689 ( \16032 , \5954 , \3432 );
nor \U$15690 ( \16033 , \16031 , \16032 );
xnor \U$15691 ( \16034 , \16033 , \3247 );
and \U$15692 ( \16035 , \6802 , \3121 );
and \U$15693 ( \16036 , \6499 , \3119 );
nor \U$15694 ( \16037 , \16035 , \16036 );
xnor \U$15695 ( \16038 , \16037 , \2916 );
and \U$15696 ( \16039 , \16034 , \16038 );
and \U$15697 ( \16040 , \7500 , \2715 );
and \U$15698 ( \16041 , \6974 , \2713 );
nor \U$15699 ( \16042 , \16040 , \16041 );
xnor \U$15700 ( \16043 , \16042 , \2566 );
and \U$15701 ( \16044 , \16038 , \16043 );
and \U$15702 ( \16045 , \16034 , \16043 );
or \U$15703 ( \16046 , \16039 , \16044 , \16045 );
and \U$15704 ( \16047 , \16029 , \16046 );
and \U$15705 ( \16048 , \16013 , \16046 );
or \U$15706 ( \16049 , \16030 , \16047 , \16048 );
and \U$15707 ( \16050 , \15997 , \16049 );
and \U$15708 ( \16051 , \9958 , \1623 );
and \U$15709 ( \16052 , \9355 , \1621 );
nor \U$15710 ( \16053 , \16051 , \16052 );
xnor \U$15711 ( \16054 , \16053 , \1467 );
and \U$15712 ( \16055 , \10144 , \1351 );
and \U$15713 ( \16056 , \9963 , \1349 );
nor \U$15714 ( \16057 , \16055 , \16056 );
xnor \U$15715 ( \16058 , \16057 , \1238 );
and \U$15716 ( \16059 , \16054 , \16058 );
nand \U$15717 ( \16060 , \10764 , \1155 );
xnor \U$15718 ( \16061 , \16060 , \1021 );
and \U$15719 ( \16062 , \16058 , \16061 );
and \U$15720 ( \16063 , \16054 , \16061 );
or \U$15721 ( \16064 , \16059 , \16062 , \16063 );
and \U$15722 ( \16065 , \8170 , \2393 );
and \U$15723 ( \16066 , \7924 , \2391 );
nor \U$15724 ( \16067 , \16065 , \16066 );
xnor \U$15725 ( \16068 , \16067 , \2251 );
and \U$15726 ( \16069 , \8494 , \2097 );
and \U$15727 ( \16070 , \8175 , \2095 );
nor \U$15728 ( \16071 , \16069 , \16070 );
xnor \U$15729 ( \16072 , \16071 , \1960 );
and \U$15730 ( \16073 , \16068 , \16072 );
and \U$15731 ( \16074 , \9347 , \1891 );
and \U$15732 ( \16075 , \8778 , \1889 );
nor \U$15733 ( \16076 , \16074 , \16075 );
xnor \U$15734 ( \16077 , \16076 , \1739 );
and \U$15735 ( \16078 , \16072 , \16077 );
and \U$15736 ( \16079 , \16068 , \16077 );
or \U$15737 ( \16080 , \16073 , \16078 , \16079 );
and \U$15738 ( \16081 , \16064 , \16080 );
and \U$15739 ( \16082 , \9963 , \1351 );
and \U$15740 ( \16083 , \9958 , \1349 );
nor \U$15741 ( \16084 , \16082 , \16083 );
xnor \U$15742 ( \16085 , \16084 , \1238 );
and \U$15743 ( \16086 , \16080 , \16085 );
and \U$15744 ( \16087 , \16064 , \16085 );
or \U$15745 ( \16088 , \16081 , \16086 , \16087 );
and \U$15746 ( \16089 , \16049 , \16088 );
and \U$15747 ( \16090 , \15997 , \16088 );
or \U$15748 ( \16091 , \16050 , \16089 , \16090 );
and \U$15749 ( \16092 , \10764 , \1157 );
and \U$15750 ( \16093 , \10144 , \1155 );
nor \U$15751 ( \16094 , \16092 , \16093 );
xnor \U$15752 ( \16095 , \16094 , \1021 );
xor \U$15753 ( \16096 , \15767 , \15771 );
xor \U$15754 ( \16097 , \16096 , \15776 );
and \U$15755 ( \16098 , \16095 , \16097 );
xor \U$15756 ( \16099 , \15839 , \15843 );
xor \U$15757 ( \16100 , \16099 , \15848 );
and \U$15758 ( \16101 , \16097 , \16100 );
and \U$15759 ( \16102 , \16095 , \16100 );
or \U$15760 ( \16103 , \16098 , \16101 , \16102 );
xor \U$15761 ( \16104 , \15734 , \15738 );
xor \U$15762 ( \16105 , \16104 , \15743 );
xor \U$15763 ( \16106 , \15750 , \15754 );
xor \U$15764 ( \16107 , \16106 , \15759 );
and \U$15765 ( \16108 , \16105 , \16107 );
xor \U$15766 ( \16109 , \15802 , \15806 );
xor \U$15767 ( \16110 , \16109 , \15811 );
and \U$15768 ( \16111 , \16107 , \16110 );
and \U$15769 ( \16112 , \16105 , \16110 );
or \U$15770 ( \16113 , \16108 , \16111 , \16112 );
and \U$15771 ( \16114 , \16103 , \16113 );
xor \U$15772 ( \16115 , \15577 , \15581 );
xor \U$15773 ( \16116 , \16115 , \879 );
and \U$15774 ( \16117 , \16113 , \16116 );
and \U$15775 ( \16118 , \16103 , \16116 );
or \U$15776 ( \16119 , \16114 , \16117 , \16118 );
and \U$15777 ( \16120 , \16091 , \16119 );
xor \U$15778 ( \16121 , \15851 , \15853 );
xor \U$15779 ( \16122 , \16121 , \15856 );
xor \U$15780 ( \16123 , \15864 , \15866 );
xor \U$15781 ( \16124 , \16123 , \15869 );
and \U$15782 ( \16125 , \16122 , \16124 );
xor \U$15783 ( \16126 , \15874 , \15876 );
xor \U$15784 ( \16127 , \16126 , \15879 );
and \U$15785 ( \16128 , \16124 , \16127 );
and \U$15786 ( \16129 , \16122 , \16127 );
or \U$15787 ( \16130 , \16125 , \16128 , \16129 );
and \U$15788 ( \16131 , \16119 , \16130 );
and \U$15789 ( \16132 , \16091 , \16130 );
or \U$15790 ( \16133 , \16120 , \16131 , \16132 );
xor \U$15791 ( \16134 , \15521 , \15537 );
xor \U$15792 ( \16135 , \16134 , \15554 );
xor \U$15793 ( \16136 , \15573 , \15585 );
xor \U$15794 ( \16137 , \16136 , \15602 );
and \U$15795 ( \16138 , \16135 , \16137 );
xor \U$15796 ( \16139 , \15891 , \15893 );
xor \U$15797 ( \16140 , \16139 , \15896 );
and \U$15798 ( \16141 , \16137 , \16140 );
and \U$15799 ( \16142 , \16135 , \16140 );
or \U$15800 ( \16143 , \16138 , \16141 , \16142 );
and \U$15801 ( \16144 , \16133 , \16143 );
xor \U$15802 ( \16145 , \15782 , \15834 );
xor \U$15803 ( \16146 , \16145 , \15859 );
xor \U$15804 ( \16147 , \15872 , \15882 );
xor \U$15805 ( \16148 , \16147 , \15885 );
and \U$15806 ( \16149 , \16146 , \16148 );
and \U$15807 ( \16150 , \16143 , \16149 );
and \U$15808 ( \16151 , \16133 , \16149 );
or \U$15809 ( \16152 , \16144 , \16150 , \16151 );
xor \U$15810 ( \16153 , \15862 , \15888 );
xor \U$15811 ( \16154 , \16153 , \15899 );
xor \U$15812 ( \16155 , \15904 , \15906 );
xor \U$15813 ( \16156 , \16155 , \15909 );
and \U$15814 ( \16157 , \16154 , \16156 );
xor \U$15815 ( \16158 , \15915 , \15917 );
and \U$15816 ( \16159 , \16156 , \16158 );
and \U$15817 ( \16160 , \16154 , \16158 );
or \U$15818 ( \16161 , \16157 , \16159 , \16160 );
and \U$15819 ( \16162 , \16152 , \16161 );
xor \U$15820 ( \16163 , \15923 , \15925 );
xor \U$15821 ( \16164 , \16163 , \15928 );
and \U$15822 ( \16165 , \16161 , \16164 );
and \U$15823 ( \16166 , \16152 , \16164 );
or \U$15824 ( \16167 , \16162 , \16165 , \16166 );
xor \U$15825 ( \16168 , \15687 , \15697 );
xor \U$15826 ( \16169 , \16168 , \15700 );
and \U$15827 ( \16170 , \16167 , \16169 );
xor \U$15828 ( \16171 , \15921 , \15931 );
xor \U$15829 ( \16172 , \16171 , \15934 );
and \U$15830 ( \16173 , \16169 , \16172 );
and \U$15831 ( \16174 , \16167 , \16172 );
or \U$15832 ( \16175 , \16170 , \16173 , \16174 );
and \U$15833 ( \16176 , \15949 , \16175 );
xor \U$15834 ( \16177 , \15949 , \16175 );
xor \U$15835 ( \16178 , \16167 , \16169 );
xor \U$15836 ( \16179 , \16178 , \16172 );
and \U$15837 ( \16180 , \1412 , \10611 );
and \U$15838 ( \16181 , \1297 , \10608 );
nor \U$15839 ( \16182 , \16180 , \16181 );
xnor \U$15840 ( \16183 , \16182 , \9556 );
and \U$15841 ( \16184 , \1596 , \9798 );
and \U$15842 ( \16185 , \1588 , \9796 );
nor \U$15843 ( \16186 , \16184 , \16185 );
xnor \U$15844 ( \16187 , \16186 , \9559 );
and \U$15845 ( \16188 , \16183 , \16187 );
and \U$15846 ( \16189 , \1844 , \9230 );
and \U$15847 ( \16190 , \1839 , \9228 );
nor \U$15848 ( \16191 , \16189 , \16190 );
xnor \U$15849 ( \16192 , \16191 , \8920 );
and \U$15850 ( \16193 , \16187 , \16192 );
and \U$15851 ( \16194 , \16183 , \16192 );
or \U$15852 ( \16195 , \16188 , \16193 , \16194 );
and \U$15853 ( \16196 , \2174 , \8693 );
and \U$15854 ( \16197 , \2030 , \8691 );
nor \U$15855 ( \16198 , \16196 , \16197 );
xnor \U$15856 ( \16199 , \16198 , \8322 );
and \U$15857 ( \16200 , \2463 , \8131 );
and \U$15858 ( \16201 , \2438 , \8129 );
nor \U$15859 ( \16202 , \16200 , \16201 );
xnor \U$15860 ( \16203 , \16202 , \7813 );
and \U$15861 ( \16204 , \16199 , \16203 );
and \U$15862 ( \16205 , \2804 , \7564 );
and \U$15863 ( \16206 , \2637 , \7562 );
nor \U$15864 ( \16207 , \16205 , \16206 );
xnor \U$15865 ( \16208 , \16207 , \7315 );
and \U$15866 ( \16209 , \16203 , \16208 );
and \U$15867 ( \16210 , \16199 , \16208 );
or \U$15868 ( \16211 , \16204 , \16209 , \16210 );
and \U$15869 ( \16212 , \16195 , \16211 );
and \U$15870 ( \16213 , \3061 , \7035 );
and \U$15871 ( \16214 , \2942 , \7033 );
nor \U$15872 ( \16215 , \16213 , \16214 );
xnor \U$15873 ( \16216 , \16215 , \6775 );
and \U$15874 ( \16217 , \3686 , \6541 );
and \U$15875 ( \16218 , \3478 , \6539 );
nor \U$15876 ( \16219 , \16217 , \16218 );
xnor \U$15877 ( \16220 , \16219 , \6226 );
and \U$15878 ( \16221 , \16216 , \16220 );
and \U$15879 ( \16222 , \3813 , \6032 );
and \U$15880 ( \16223 , \3808 , \6030 );
nor \U$15881 ( \16224 , \16222 , \16223 );
xnor \U$15882 ( \16225 , \16224 , \5692 );
and \U$15883 ( \16226 , \16220 , \16225 );
and \U$15884 ( \16227 , \16216 , \16225 );
or \U$15885 ( \16228 , \16221 , \16226 , \16227 );
and \U$15886 ( \16229 , \16211 , \16228 );
and \U$15887 ( \16230 , \16195 , \16228 );
or \U$15888 ( \16231 , \16212 , \16229 , \16230 );
and \U$15889 ( \16232 , \5573 , \4152 );
and \U$15890 ( \16233 , \5314 , \4150 );
nor \U$15891 ( \16234 , \16232 , \16233 );
xnor \U$15892 ( \16235 , \16234 , \4009 );
and \U$15893 ( \16236 , \5954 , \3829 );
and \U$15894 ( \16237 , \5945 , \3827 );
nor \U$15895 ( \16238 , \16236 , \16237 );
xnor \U$15896 ( \16239 , \16238 , \3583 );
and \U$15897 ( \16240 , \16235 , \16239 );
and \U$15898 ( \16241 , \6499 , \3434 );
and \U$15899 ( \16242 , \6297 , \3432 );
nor \U$15900 ( \16243 , \16241 , \16242 );
xnor \U$15901 ( \16244 , \16243 , \3247 );
and \U$15902 ( \16245 , \16239 , \16244 );
and \U$15903 ( \16246 , \16235 , \16244 );
or \U$15904 ( \16247 , \16240 , \16245 , \16246 );
and \U$15905 ( \16248 , \6974 , \3121 );
and \U$15906 ( \16249 , \6802 , \3119 );
nor \U$15907 ( \16250 , \16248 , \16249 );
xnor \U$15908 ( \16251 , \16250 , \2916 );
and \U$15909 ( \16252 , \7924 , \2715 );
and \U$15910 ( \16253 , \7500 , \2713 );
nor \U$15911 ( \16254 , \16252 , \16253 );
xnor \U$15912 ( \16255 , \16254 , \2566 );
and \U$15913 ( \16256 , \16251 , \16255 );
and \U$15914 ( \16257 , \8175 , \2393 );
and \U$15915 ( \16258 , \8170 , \2391 );
nor \U$15916 ( \16259 , \16257 , \16258 );
xnor \U$15917 ( \16260 , \16259 , \2251 );
and \U$15918 ( \16261 , \16255 , \16260 );
and \U$15919 ( \16262 , \16251 , \16260 );
or \U$15920 ( \16263 , \16256 , \16261 , \16262 );
and \U$15921 ( \16264 , \16247 , \16263 );
and \U$15922 ( \16265 , \4266 , \5443 );
and \U$15923 ( \16266 , \4069 , \5441 );
nor \U$15924 ( \16267 , \16265 , \16266 );
xnor \U$15925 ( \16268 , \16267 , \5202 );
and \U$15926 ( \16269 , \4576 , \4977 );
and \U$15927 ( \16270 , \4568 , \4975 );
nor \U$15928 ( \16271 , \16269 , \16270 );
xnor \U$15929 ( \16272 , \16271 , \4789 );
and \U$15930 ( \16273 , \16268 , \16272 );
and \U$15931 ( \16274 , \5050 , \4603 );
and \U$15932 ( \16275 , \5045 , \4601 );
nor \U$15933 ( \16276 , \16274 , \16275 );
xnor \U$15934 ( \16277 , \16276 , \4371 );
and \U$15935 ( \16278 , \16272 , \16277 );
and \U$15936 ( \16279 , \16268 , \16277 );
or \U$15937 ( \16280 , \16273 , \16278 , \16279 );
and \U$15938 ( \16281 , \16263 , \16280 );
and \U$15939 ( \16282 , \16247 , \16280 );
or \U$15940 ( \16283 , \16264 , \16281 , \16282 );
and \U$15941 ( \16284 , \16231 , \16283 );
and \U$15942 ( \16285 , \8778 , \2097 );
and \U$15943 ( \16286 , \8494 , \2095 );
nor \U$15944 ( \16287 , \16285 , \16286 );
xnor \U$15945 ( \16288 , \16287 , \1960 );
and \U$15946 ( \16289 , \9355 , \1891 );
and \U$15947 ( \16290 , \9347 , \1889 );
nor \U$15948 ( \16291 , \16289 , \16290 );
xnor \U$15949 ( \16292 , \16291 , \1739 );
and \U$15950 ( \16293 , \16288 , \16292 );
and \U$15951 ( \16294 , \9963 , \1623 );
and \U$15952 ( \16295 , \9958 , \1621 );
nor \U$15953 ( \16296 , \16294 , \16295 );
xnor \U$15954 ( \16297 , \16296 , \1467 );
and \U$15955 ( \16298 , \16292 , \16297 );
and \U$15956 ( \16299 , \16288 , \16297 );
or \U$15957 ( \16300 , \16293 , \16298 , \16299 );
xor \U$15958 ( \16301 , \16054 , \16058 );
xor \U$15959 ( \16302 , \16301 , \16061 );
and \U$15960 ( \16303 , \16300 , \16302 );
xor \U$15961 ( \16304 , \16068 , \16072 );
xor \U$15962 ( \16305 , \16304 , \16077 );
and \U$15963 ( \16306 , \16302 , \16305 );
and \U$15964 ( \16307 , \16300 , \16305 );
or \U$15965 ( \16308 , \16303 , \16306 , \16307 );
and \U$15966 ( \16309 , \16283 , \16308 );
and \U$15967 ( \16310 , \16231 , \16308 );
or \U$15968 ( \16311 , \16284 , \16309 , \16310 );
xor \U$15969 ( \16312 , \16001 , \16005 );
xor \U$15970 ( \16313 , \16312 , \16010 );
xor \U$15971 ( \16314 , \16017 , \16021 );
xor \U$15972 ( \16315 , \16314 , \16026 );
and \U$15973 ( \16316 , \16313 , \16315 );
xor \U$15974 ( \16317 , \16034 , \16038 );
xor \U$15975 ( \16318 , \16317 , \16043 );
and \U$15976 ( \16319 , \16315 , \16318 );
and \U$15977 ( \16320 , \16313 , \16318 );
or \U$15978 ( \16321 , \16316 , \16319 , \16320 );
xor \U$15979 ( \16322 , \15953 , \15957 );
xor \U$15980 ( \16323 , \16322 , \1021 );
xor \U$15981 ( \16324 , \15965 , \15969 );
xor \U$15982 ( \16325 , \16324 , \15974 );
and \U$15983 ( \16326 , \16323 , \16325 );
xor \U$15984 ( \16327 , \15982 , \15986 );
xor \U$15985 ( \16328 , \16327 , \15991 );
and \U$15986 ( \16329 , \16325 , \16328 );
and \U$15987 ( \16330 , \16323 , \16328 );
or \U$15988 ( \16331 , \16326 , \16329 , \16330 );
and \U$15989 ( \16332 , \16321 , \16331 );
xor \U$15990 ( \16333 , \15786 , \15790 );
xor \U$15991 ( \16334 , \16333 , \15795 );
and \U$15992 ( \16335 , \16331 , \16334 );
and \U$15993 ( \16336 , \16321 , \16334 );
or \U$15994 ( \16337 , \16332 , \16335 , \16336 );
and \U$15995 ( \16338 , \16311 , \16337 );
xor \U$15996 ( \16339 , \15819 , \15823 );
xor \U$15997 ( \16340 , \16339 , \15828 );
xor \U$15998 ( \16341 , \16095 , \16097 );
xor \U$15999 ( \16342 , \16341 , \16100 );
and \U$16000 ( \16343 , \16340 , \16342 );
xor \U$16001 ( \16344 , \16105 , \16107 );
xor \U$16002 ( \16345 , \16344 , \16110 );
and \U$16003 ( \16346 , \16342 , \16345 );
and \U$16004 ( \16347 , \16340 , \16345 );
or \U$16005 ( \16348 , \16343 , \16346 , \16347 );
and \U$16006 ( \16349 , \16337 , \16348 );
and \U$16007 ( \16350 , \16311 , \16348 );
or \U$16008 ( \16351 , \16338 , \16349 , \16350 );
xor \U$16009 ( \16352 , \15961 , \15977 );
xor \U$16010 ( \16353 , \16352 , \15994 );
xor \U$16011 ( \16354 , \16013 , \16029 );
xor \U$16012 ( \16355 , \16354 , \16046 );
and \U$16013 ( \16356 , \16353 , \16355 );
xor \U$16014 ( \16357 , \16064 , \16080 );
xor \U$16015 ( \16358 , \16357 , \16085 );
and \U$16016 ( \16359 , \16355 , \16358 );
and \U$16017 ( \16360 , \16353 , \16358 );
or \U$16018 ( \16361 , \16356 , \16359 , \16360 );
xor \U$16019 ( \16362 , \15746 , \15762 );
xor \U$16020 ( \16363 , \16362 , \15779 );
and \U$16021 ( \16364 , \16361 , \16363 );
xor \U$16022 ( \16365 , \15798 , \15814 );
xor \U$16023 ( \16366 , \16365 , \15831 );
and \U$16024 ( \16367 , \16363 , \16366 );
and \U$16025 ( \16368 , \16361 , \16366 );
or \U$16026 ( \16369 , \16364 , \16367 , \16368 );
and \U$16027 ( \16370 , \16351 , \16369 );
xor \U$16028 ( \16371 , \15997 , \16049 );
xor \U$16029 ( \16372 , \16371 , \16088 );
xor \U$16030 ( \16373 , \16103 , \16113 );
xor \U$16031 ( \16374 , \16373 , \16116 );
and \U$16032 ( \16375 , \16372 , \16374 );
xor \U$16033 ( \16376 , \16122 , \16124 );
xor \U$16034 ( \16377 , \16376 , \16127 );
and \U$16035 ( \16378 , \16374 , \16377 );
and \U$16036 ( \16379 , \16372 , \16377 );
or \U$16037 ( \16380 , \16375 , \16378 , \16379 );
and \U$16038 ( \16381 , \16369 , \16380 );
and \U$16039 ( \16382 , \16351 , \16380 );
or \U$16040 ( \16383 , \16370 , \16381 , \16382 );
xor \U$16041 ( \16384 , \16091 , \16119 );
xor \U$16042 ( \16385 , \16384 , \16130 );
xor \U$16043 ( \16386 , \16135 , \16137 );
xor \U$16044 ( \16387 , \16386 , \16140 );
and \U$16045 ( \16388 , \16385 , \16387 );
xor \U$16046 ( \16389 , \16146 , \16148 );
and \U$16047 ( \16390 , \16387 , \16389 );
and \U$16048 ( \16391 , \16385 , \16389 );
or \U$16049 ( \16392 , \16388 , \16390 , \16391 );
and \U$16050 ( \16393 , \16383 , \16392 );
xor \U$16051 ( \16394 , \16154 , \16156 );
xor \U$16052 ( \16395 , \16394 , \16158 );
and \U$16053 ( \16396 , \16392 , \16395 );
and \U$16054 ( \16397 , \16383 , \16395 );
or \U$16055 ( \16398 , \16393 , \16396 , \16397 );
xor \U$16056 ( \16399 , \15902 , \15912 );
xor \U$16057 ( \16400 , \16399 , \15918 );
and \U$16058 ( \16401 , \16398 , \16400 );
xor \U$16059 ( \16402 , \16152 , \16161 );
xor \U$16060 ( \16403 , \16402 , \16164 );
and \U$16061 ( \16404 , \16400 , \16403 );
and \U$16062 ( \16405 , \16398 , \16403 );
or \U$16063 ( \16406 , \16401 , \16404 , \16405 );
and \U$16064 ( \16407 , \16179 , \16406 );
xor \U$16065 ( \16408 , \16179 , \16406 );
xor \U$16066 ( \16409 , \16398 , \16400 );
xor \U$16067 ( \16410 , \16409 , \16403 );
and \U$16068 ( \16411 , \6802 , \3434 );
and \U$16069 ( \16412 , \6499 , \3432 );
nor \U$16070 ( \16413 , \16411 , \16412 );
xnor \U$16071 ( \16414 , \16413 , \3247 );
and \U$16072 ( \16415 , \7500 , \3121 );
and \U$16073 ( \16416 , \6974 , \3119 );
nor \U$16074 ( \16417 , \16415 , \16416 );
xnor \U$16075 ( \16418 , \16417 , \2916 );
and \U$16076 ( \16419 , \16414 , \16418 );
and \U$16077 ( \16420 , \8170 , \2715 );
and \U$16078 ( \16421 , \7924 , \2713 );
nor \U$16079 ( \16422 , \16420 , \16421 );
xnor \U$16080 ( \16423 , \16422 , \2566 );
and \U$16081 ( \16424 , \16418 , \16423 );
and \U$16082 ( \16425 , \16414 , \16423 );
or \U$16083 ( \16426 , \16419 , \16424 , \16425 );
and \U$16084 ( \16427 , \4069 , \6032 );
and \U$16085 ( \16428 , \3813 , \6030 );
nor \U$16086 ( \16429 , \16427 , \16428 );
xnor \U$16087 ( \16430 , \16429 , \5692 );
and \U$16088 ( \16431 , \4568 , \5443 );
and \U$16089 ( \16432 , \4266 , \5441 );
nor \U$16090 ( \16433 , \16431 , \16432 );
xnor \U$16091 ( \16434 , \16433 , \5202 );
and \U$16092 ( \16435 , \16430 , \16434 );
and \U$16093 ( \16436 , \5045 , \4977 );
and \U$16094 ( \16437 , \4576 , \4975 );
nor \U$16095 ( \16438 , \16436 , \16437 );
xnor \U$16096 ( \16439 , \16438 , \4789 );
and \U$16097 ( \16440 , \16434 , \16439 );
and \U$16098 ( \16441 , \16430 , \16439 );
or \U$16099 ( \16442 , \16435 , \16440 , \16441 );
and \U$16100 ( \16443 , \16426 , \16442 );
and \U$16101 ( \16444 , \5314 , \4603 );
and \U$16102 ( \16445 , \5050 , \4601 );
nor \U$16103 ( \16446 , \16444 , \16445 );
xnor \U$16104 ( \16447 , \16446 , \4371 );
and \U$16105 ( \16448 , \5945 , \4152 );
and \U$16106 ( \16449 , \5573 , \4150 );
nor \U$16107 ( \16450 , \16448 , \16449 );
xnor \U$16108 ( \16451 , \16450 , \4009 );
and \U$16109 ( \16452 , \16447 , \16451 );
and \U$16110 ( \16453 , \6297 , \3829 );
and \U$16111 ( \16454 , \5954 , \3827 );
nor \U$16112 ( \16455 , \16453 , \16454 );
xnor \U$16113 ( \16456 , \16455 , \3583 );
and \U$16114 ( \16457 , \16451 , \16456 );
and \U$16115 ( \16458 , \16447 , \16456 );
or \U$16116 ( \16459 , \16452 , \16457 , \16458 );
and \U$16117 ( \16460 , \16442 , \16459 );
and \U$16118 ( \16461 , \16426 , \16459 );
or \U$16119 ( \16462 , \16443 , \16460 , \16461 );
and \U$16120 ( \16463 , \1588 , \10611 );
and \U$16121 ( \16464 , \1412 , \10608 );
nor \U$16122 ( \16465 , \16463 , \16464 );
xnor \U$16123 ( \16466 , \16465 , \9556 );
and \U$16124 ( \16467 , \1839 , \9798 );
and \U$16125 ( \16468 , \1596 , \9796 );
nor \U$16126 ( \16469 , \16467 , \16468 );
xnor \U$16127 ( \16470 , \16469 , \9559 );
and \U$16128 ( \16471 , \16466 , \16470 );
and \U$16129 ( \16472 , \16470 , \1238 );
and \U$16130 ( \16473 , \16466 , \1238 );
or \U$16131 ( \16474 , \16471 , \16472 , \16473 );
and \U$16132 ( \16475 , \2942 , \7564 );
and \U$16133 ( \16476 , \2804 , \7562 );
nor \U$16134 ( \16477 , \16475 , \16476 );
xnor \U$16135 ( \16478 , \16477 , \7315 );
and \U$16136 ( \16479 , \3478 , \7035 );
and \U$16137 ( \16480 , \3061 , \7033 );
nor \U$16138 ( \16481 , \16479 , \16480 );
xnor \U$16139 ( \16482 , \16481 , \6775 );
and \U$16140 ( \16483 , \16478 , \16482 );
and \U$16141 ( \16484 , \3808 , \6541 );
and \U$16142 ( \16485 , \3686 , \6539 );
nor \U$16143 ( \16486 , \16484 , \16485 );
xnor \U$16144 ( \16487 , \16486 , \6226 );
and \U$16145 ( \16488 , \16482 , \16487 );
and \U$16146 ( \16489 , \16478 , \16487 );
or \U$16147 ( \16490 , \16483 , \16488 , \16489 );
and \U$16148 ( \16491 , \16474 , \16490 );
and \U$16149 ( \16492 , \2030 , \9230 );
and \U$16150 ( \16493 , \1844 , \9228 );
nor \U$16151 ( \16494 , \16492 , \16493 );
xnor \U$16152 ( \16495 , \16494 , \8920 );
and \U$16153 ( \16496 , \2438 , \8693 );
and \U$16154 ( \16497 , \2174 , \8691 );
nor \U$16155 ( \16498 , \16496 , \16497 );
xnor \U$16156 ( \16499 , \16498 , \8322 );
and \U$16157 ( \16500 , \16495 , \16499 );
and \U$16158 ( \16501 , \2637 , \8131 );
and \U$16159 ( \16502 , \2463 , \8129 );
nor \U$16160 ( \16503 , \16501 , \16502 );
xnor \U$16161 ( \16504 , \16503 , \7813 );
and \U$16162 ( \16505 , \16499 , \16504 );
and \U$16163 ( \16506 , \16495 , \16504 );
or \U$16164 ( \16507 , \16500 , \16505 , \16506 );
and \U$16165 ( \16508 , \16490 , \16507 );
and \U$16166 ( \16509 , \16474 , \16507 );
or \U$16167 ( \16510 , \16491 , \16508 , \16509 );
and \U$16168 ( \16511 , \16462 , \16510 );
and \U$16169 ( \16512 , \8494 , \2393 );
and \U$16170 ( \16513 , \8175 , \2391 );
nor \U$16171 ( \16514 , \16512 , \16513 );
xnor \U$16172 ( \16515 , \16514 , \2251 );
and \U$16173 ( \16516 , \9347 , \2097 );
and \U$16174 ( \16517 , \8778 , \2095 );
nor \U$16175 ( \16518 , \16516 , \16517 );
xnor \U$16176 ( \16519 , \16518 , \1960 );
and \U$16177 ( \16520 , \16515 , \16519 );
and \U$16178 ( \16521 , \9958 , \1891 );
and \U$16179 ( \16522 , \9355 , \1889 );
nor \U$16180 ( \16523 , \16521 , \16522 );
xnor \U$16181 ( \16524 , \16523 , \1739 );
and \U$16182 ( \16525 , \16519 , \16524 );
and \U$16183 ( \16526 , \16515 , \16524 );
or \U$16184 ( \16527 , \16520 , \16525 , \16526 );
and \U$16185 ( \16528 , \10144 , \1623 );
and \U$16186 ( \16529 , \9963 , \1621 );
nor \U$16187 ( \16530 , \16528 , \16529 );
xnor \U$16188 ( \16531 , \16530 , \1467 );
nand \U$16189 ( \16532 , \10764 , \1349 );
xnor \U$16190 ( \16533 , \16532 , \1238 );
and \U$16191 ( \16534 , \16531 , \16533 );
and \U$16192 ( \16535 , \16527 , \16534 );
and \U$16193 ( \16536 , \10764 , \1351 );
and \U$16194 ( \16537 , \10144 , \1349 );
nor \U$16195 ( \16538 , \16536 , \16537 );
xnor \U$16196 ( \16539 , \16538 , \1238 );
and \U$16197 ( \16540 , \16534 , \16539 );
and \U$16198 ( \16541 , \16527 , \16539 );
or \U$16199 ( \16542 , \16535 , \16540 , \16541 );
and \U$16200 ( \16543 , \16510 , \16542 );
and \U$16201 ( \16544 , \16462 , \16542 );
or \U$16202 ( \16545 , \16511 , \16543 , \16544 );
xor \U$16203 ( \16546 , \16199 , \16203 );
xor \U$16204 ( \16547 , \16546 , \16208 );
xor \U$16205 ( \16548 , \16268 , \16272 );
xor \U$16206 ( \16549 , \16548 , \16277 );
and \U$16207 ( \16550 , \16547 , \16549 );
xor \U$16208 ( \16551 , \16216 , \16220 );
xor \U$16209 ( \16552 , \16551 , \16225 );
and \U$16210 ( \16553 , \16549 , \16552 );
and \U$16211 ( \16554 , \16547 , \16552 );
or \U$16212 ( \16555 , \16550 , \16553 , \16554 );
xor \U$16213 ( \16556 , \16235 , \16239 );
xor \U$16214 ( \16557 , \16556 , \16244 );
xor \U$16215 ( \16558 , \16288 , \16292 );
xor \U$16216 ( \16559 , \16558 , \16297 );
and \U$16217 ( \16560 , \16557 , \16559 );
xor \U$16218 ( \16561 , \16251 , \16255 );
xor \U$16219 ( \16562 , \16561 , \16260 );
and \U$16220 ( \16563 , \16559 , \16562 );
and \U$16221 ( \16564 , \16557 , \16562 );
or \U$16222 ( \16565 , \16560 , \16563 , \16564 );
and \U$16223 ( \16566 , \16555 , \16565 );
xor \U$16224 ( \16567 , \16323 , \16325 );
xor \U$16225 ( \16568 , \16567 , \16328 );
and \U$16226 ( \16569 , \16565 , \16568 );
and \U$16227 ( \16570 , \16555 , \16568 );
or \U$16228 ( \16571 , \16566 , \16569 , \16570 );
and \U$16229 ( \16572 , \16545 , \16571 );
xor \U$16230 ( \16573 , \16247 , \16263 );
xor \U$16231 ( \16574 , \16573 , \16280 );
xor \U$16232 ( \16575 , \16313 , \16315 );
xor \U$16233 ( \16576 , \16575 , \16318 );
and \U$16234 ( \16577 , \16574 , \16576 );
xor \U$16235 ( \16578 , \16300 , \16302 );
xor \U$16236 ( \16579 , \16578 , \16305 );
and \U$16237 ( \16580 , \16576 , \16579 );
and \U$16238 ( \16581 , \16574 , \16579 );
or \U$16239 ( \16582 , \16577 , \16580 , \16581 );
and \U$16240 ( \16583 , \16571 , \16582 );
and \U$16241 ( \16584 , \16545 , \16582 );
or \U$16242 ( \16585 , \16572 , \16583 , \16584 );
xor \U$16243 ( \16586 , \16353 , \16355 );
xor \U$16244 ( \16587 , \16586 , \16358 );
xor \U$16245 ( \16588 , \16321 , \16331 );
xor \U$16246 ( \16589 , \16588 , \16334 );
and \U$16247 ( \16590 , \16587 , \16589 );
xor \U$16248 ( \16591 , \16340 , \16342 );
xor \U$16249 ( \16592 , \16591 , \16345 );
and \U$16250 ( \16593 , \16589 , \16592 );
and \U$16251 ( \16594 , \16587 , \16592 );
or \U$16252 ( \16595 , \16590 , \16593 , \16594 );
and \U$16253 ( \16596 , \16585 , \16595 );
xor \U$16254 ( \16597 , \16372 , \16374 );
xor \U$16255 ( \16598 , \16597 , \16377 );
and \U$16256 ( \16599 , \16595 , \16598 );
and \U$16257 ( \16600 , \16585 , \16598 );
or \U$16258 ( \16601 , \16596 , \16599 , \16600 );
xor \U$16259 ( \16602 , \16351 , \16369 );
xor \U$16260 ( \16603 , \16602 , \16380 );
and \U$16261 ( \16604 , \16601 , \16603 );
xor \U$16262 ( \16605 , \16385 , \16387 );
xor \U$16263 ( \16606 , \16605 , \16389 );
and \U$16264 ( \16607 , \16603 , \16606 );
and \U$16265 ( \16608 , \16601 , \16606 );
or \U$16266 ( \16609 , \16604 , \16607 , \16608 );
xor \U$16267 ( \16610 , \16133 , \16143 );
xor \U$16268 ( \16611 , \16610 , \16149 );
and \U$16269 ( \16612 , \16609 , \16611 );
xor \U$16270 ( \16613 , \16383 , \16392 );
xor \U$16271 ( \16614 , \16613 , \16395 );
and \U$16272 ( \16615 , \16611 , \16614 );
and \U$16273 ( \16616 , \16609 , \16614 );
or \U$16274 ( \16617 , \16612 , \16615 , \16616 );
and \U$16275 ( \16618 , \16410 , \16617 );
xor \U$16276 ( \16619 , \16410 , \16617 );
xor \U$16277 ( \16620 , \16609 , \16611 );
xor \U$16278 ( \16621 , \16620 , \16614 );
and \U$16279 ( \16622 , \5954 , \4152 );
and \U$16280 ( \16623 , \5945 , \4150 );
nor \U$16281 ( \16624 , \16622 , \16623 );
xnor \U$16282 ( \16625 , \16624 , \4009 );
and \U$16283 ( \16626 , \6499 , \3829 );
and \U$16284 ( \16627 , \6297 , \3827 );
nor \U$16285 ( \16628 , \16626 , \16627 );
xnor \U$16286 ( \16629 , \16628 , \3583 );
and \U$16287 ( \16630 , \16625 , \16629 );
and \U$16288 ( \16631 , \6974 , \3434 );
and \U$16289 ( \16632 , \6802 , \3432 );
nor \U$16290 ( \16633 , \16631 , \16632 );
xnor \U$16291 ( \16634 , \16633 , \3247 );
and \U$16292 ( \16635 , \16629 , \16634 );
and \U$16293 ( \16636 , \16625 , \16634 );
or \U$16294 ( \16637 , \16630 , \16635 , \16636 );
and \U$16295 ( \16638 , \7924 , \3121 );
and \U$16296 ( \16639 , \7500 , \3119 );
nor \U$16297 ( \16640 , \16638 , \16639 );
xnor \U$16298 ( \16641 , \16640 , \2916 );
and \U$16299 ( \16642 , \8175 , \2715 );
and \U$16300 ( \16643 , \8170 , \2713 );
nor \U$16301 ( \16644 , \16642 , \16643 );
xnor \U$16302 ( \16645 , \16644 , \2566 );
and \U$16303 ( \16646 , \16641 , \16645 );
and \U$16304 ( \16647 , \8778 , \2393 );
and \U$16305 ( \16648 , \8494 , \2391 );
nor \U$16306 ( \16649 , \16647 , \16648 );
xnor \U$16307 ( \16650 , \16649 , \2251 );
and \U$16308 ( \16651 , \16645 , \16650 );
and \U$16309 ( \16652 , \16641 , \16650 );
or \U$16310 ( \16653 , \16646 , \16651 , \16652 );
and \U$16311 ( \16654 , \16637 , \16653 );
and \U$16312 ( \16655 , \4576 , \5443 );
and \U$16313 ( \16656 , \4568 , \5441 );
nor \U$16314 ( \16657 , \16655 , \16656 );
xnor \U$16315 ( \16658 , \16657 , \5202 );
and \U$16316 ( \16659 , \5050 , \4977 );
and \U$16317 ( \16660 , \5045 , \4975 );
nor \U$16318 ( \16661 , \16659 , \16660 );
xnor \U$16319 ( \16662 , \16661 , \4789 );
and \U$16320 ( \16663 , \16658 , \16662 );
and \U$16321 ( \16664 , \5573 , \4603 );
and \U$16322 ( \16665 , \5314 , \4601 );
nor \U$16323 ( \16666 , \16664 , \16665 );
xnor \U$16324 ( \16667 , \16666 , \4371 );
and \U$16325 ( \16668 , \16662 , \16667 );
and \U$16326 ( \16669 , \16658 , \16667 );
or \U$16327 ( \16670 , \16663 , \16668 , \16669 );
and \U$16328 ( \16671 , \16653 , \16670 );
and \U$16329 ( \16672 , \16637 , \16670 );
or \U$16330 ( \16673 , \16654 , \16671 , \16672 );
and \U$16331 ( \16674 , \3686 , \7035 );
and \U$16332 ( \16675 , \3478 , \7033 );
nor \U$16333 ( \16676 , \16674 , \16675 );
xnor \U$16334 ( \16677 , \16676 , \6775 );
and \U$16335 ( \16678 , \3813 , \6541 );
and \U$16336 ( \16679 , \3808 , \6539 );
nor \U$16337 ( \16680 , \16678 , \16679 );
xnor \U$16338 ( \16681 , \16680 , \6226 );
and \U$16339 ( \16682 , \16677 , \16681 );
and \U$16340 ( \16683 , \4266 , \6032 );
and \U$16341 ( \16684 , \4069 , \6030 );
nor \U$16342 ( \16685 , \16683 , \16684 );
xnor \U$16343 ( \16686 , \16685 , \5692 );
and \U$16344 ( \16687 , \16681 , \16686 );
and \U$16345 ( \16688 , \16677 , \16686 );
or \U$16346 ( \16689 , \16682 , \16687 , \16688 );
and \U$16347 ( \16690 , \2463 , \8693 );
and \U$16348 ( \16691 , \2438 , \8691 );
nor \U$16349 ( \16692 , \16690 , \16691 );
xnor \U$16350 ( \16693 , \16692 , \8322 );
and \U$16351 ( \16694 , \2804 , \8131 );
and \U$16352 ( \16695 , \2637 , \8129 );
nor \U$16353 ( \16696 , \16694 , \16695 );
xnor \U$16354 ( \16697 , \16696 , \7813 );
and \U$16355 ( \16698 , \16693 , \16697 );
and \U$16356 ( \16699 , \3061 , \7564 );
and \U$16357 ( \16700 , \2942 , \7562 );
nor \U$16358 ( \16701 , \16699 , \16700 );
xnor \U$16359 ( \16702 , \16701 , \7315 );
and \U$16360 ( \16703 , \16697 , \16702 );
and \U$16361 ( \16704 , \16693 , \16702 );
or \U$16362 ( \16705 , \16698 , \16703 , \16704 );
and \U$16363 ( \16706 , \16689 , \16705 );
and \U$16364 ( \16707 , \1596 , \10611 );
and \U$16365 ( \16708 , \1588 , \10608 );
nor \U$16366 ( \16709 , \16707 , \16708 );
xnor \U$16367 ( \16710 , \16709 , \9556 );
and \U$16368 ( \16711 , \1844 , \9798 );
and \U$16369 ( \16712 , \1839 , \9796 );
nor \U$16370 ( \16713 , \16711 , \16712 );
xnor \U$16371 ( \16714 , \16713 , \9559 );
and \U$16372 ( \16715 , \16710 , \16714 );
and \U$16373 ( \16716 , \2174 , \9230 );
and \U$16374 ( \16717 , \2030 , \9228 );
nor \U$16375 ( \16718 , \16716 , \16717 );
xnor \U$16376 ( \16719 , \16718 , \8920 );
and \U$16377 ( \16720 , \16714 , \16719 );
and \U$16378 ( \16721 , \16710 , \16719 );
or \U$16379 ( \16722 , \16715 , \16720 , \16721 );
and \U$16380 ( \16723 , \16705 , \16722 );
and \U$16381 ( \16724 , \16689 , \16722 );
or \U$16382 ( \16725 , \16706 , \16723 , \16724 );
and \U$16383 ( \16726 , \16673 , \16725 );
and \U$16384 ( \16727 , \9355 , \2097 );
and \U$16385 ( \16728 , \9347 , \2095 );
nor \U$16386 ( \16729 , \16727 , \16728 );
xnor \U$16387 ( \16730 , \16729 , \1960 );
and \U$16388 ( \16731 , \9963 , \1891 );
and \U$16389 ( \16732 , \9958 , \1889 );
nor \U$16390 ( \16733 , \16731 , \16732 );
xnor \U$16391 ( \16734 , \16733 , \1739 );
and \U$16392 ( \16735 , \16730 , \16734 );
and \U$16393 ( \16736 , \10764 , \1623 );
and \U$16394 ( \16737 , \10144 , \1621 );
nor \U$16395 ( \16738 , \16736 , \16737 );
xnor \U$16396 ( \16739 , \16738 , \1467 );
and \U$16397 ( \16740 , \16734 , \16739 );
and \U$16398 ( \16741 , \16730 , \16739 );
or \U$16399 ( \16742 , \16735 , \16740 , \16741 );
xor \U$16400 ( \16743 , \16515 , \16519 );
xor \U$16401 ( \16744 , \16743 , \16524 );
and \U$16402 ( \16745 , \16742 , \16744 );
xor \U$16403 ( \16746 , \16531 , \16533 );
and \U$16404 ( \16747 , \16744 , \16746 );
and \U$16405 ( \16748 , \16742 , \16746 );
or \U$16406 ( \16749 , \16745 , \16747 , \16748 );
and \U$16407 ( \16750 , \16725 , \16749 );
and \U$16408 ( \16751 , \16673 , \16749 );
or \U$16409 ( \16752 , \16726 , \16750 , \16751 );
xor \U$16410 ( \16753 , \16466 , \16470 );
xor \U$16411 ( \16754 , \16753 , \1238 );
xor \U$16412 ( \16755 , \16478 , \16482 );
xor \U$16413 ( \16756 , \16755 , \16487 );
and \U$16414 ( \16757 , \16754 , \16756 );
xor \U$16415 ( \16758 , \16495 , \16499 );
xor \U$16416 ( \16759 , \16758 , \16504 );
and \U$16417 ( \16760 , \16756 , \16759 );
and \U$16418 ( \16761 , \16754 , \16759 );
or \U$16419 ( \16762 , \16757 , \16760 , \16761 );
xor \U$16420 ( \16763 , \16414 , \16418 );
xor \U$16421 ( \16764 , \16763 , \16423 );
xor \U$16422 ( \16765 , \16430 , \16434 );
xor \U$16423 ( \16766 , \16765 , \16439 );
and \U$16424 ( \16767 , \16764 , \16766 );
xor \U$16425 ( \16768 , \16447 , \16451 );
xor \U$16426 ( \16769 , \16768 , \16456 );
and \U$16427 ( \16770 , \16766 , \16769 );
and \U$16428 ( \16771 , \16764 , \16769 );
or \U$16429 ( \16772 , \16767 , \16770 , \16771 );
and \U$16430 ( \16773 , \16762 , \16772 );
xor \U$16431 ( \16774 , \16183 , \16187 );
xor \U$16432 ( \16775 , \16774 , \16192 );
and \U$16433 ( \16776 , \16772 , \16775 );
and \U$16434 ( \16777 , \16762 , \16775 );
or \U$16435 ( \16778 , \16773 , \16776 , \16777 );
and \U$16436 ( \16779 , \16752 , \16778 );
xor \U$16437 ( \16780 , \16527 , \16534 );
xor \U$16438 ( \16781 , \16780 , \16539 );
xor \U$16439 ( \16782 , \16547 , \16549 );
xor \U$16440 ( \16783 , \16782 , \16552 );
and \U$16441 ( \16784 , \16781 , \16783 );
xor \U$16442 ( \16785 , \16557 , \16559 );
xor \U$16443 ( \16786 , \16785 , \16562 );
and \U$16444 ( \16787 , \16783 , \16786 );
and \U$16445 ( \16788 , \16781 , \16786 );
or \U$16446 ( \16789 , \16784 , \16787 , \16788 );
and \U$16447 ( \16790 , \16778 , \16789 );
and \U$16448 ( \16791 , \16752 , \16789 );
or \U$16449 ( \16792 , \16779 , \16790 , \16791 );
xor \U$16450 ( \16793 , \16195 , \16211 );
xor \U$16451 ( \16794 , \16793 , \16228 );
xor \U$16452 ( \16795 , \16555 , \16565 );
xor \U$16453 ( \16796 , \16795 , \16568 );
and \U$16454 ( \16797 , \16794 , \16796 );
xor \U$16455 ( \16798 , \16574 , \16576 );
xor \U$16456 ( \16799 , \16798 , \16579 );
and \U$16457 ( \16800 , \16796 , \16799 );
and \U$16458 ( \16801 , \16794 , \16799 );
or \U$16459 ( \16802 , \16797 , \16800 , \16801 );
and \U$16460 ( \16803 , \16792 , \16802 );
xor \U$16461 ( \16804 , \16231 , \16283 );
xor \U$16462 ( \16805 , \16804 , \16308 );
and \U$16463 ( \16806 , \16802 , \16805 );
and \U$16464 ( \16807 , \16792 , \16805 );
or \U$16465 ( \16808 , \16803 , \16806 , \16807 );
xor \U$16466 ( \16809 , \16545 , \16571 );
xor \U$16467 ( \16810 , \16809 , \16582 );
xor \U$16468 ( \16811 , \16587 , \16589 );
xor \U$16469 ( \16812 , \16811 , \16592 );
and \U$16470 ( \16813 , \16810 , \16812 );
and \U$16471 ( \16814 , \16808 , \16813 );
xor \U$16472 ( \16815 , \16361 , \16363 );
xor \U$16473 ( \16816 , \16815 , \16366 );
and \U$16474 ( \16817 , \16813 , \16816 );
and \U$16475 ( \16818 , \16808 , \16816 );
or \U$16476 ( \16819 , \16814 , \16817 , \16818 );
xor \U$16477 ( \16820 , \16311 , \16337 );
xor \U$16478 ( \16821 , \16820 , \16348 );
xor \U$16479 ( \16822 , \16585 , \16595 );
xor \U$16480 ( \16823 , \16822 , \16598 );
and \U$16481 ( \16824 , \16821 , \16823 );
and \U$16482 ( \16825 , \16819 , \16824 );
xor \U$16483 ( \16826 , \16601 , \16603 );
xor \U$16484 ( \16827 , \16826 , \16606 );
and \U$16485 ( \16828 , \16824 , \16827 );
and \U$16486 ( \16829 , \16819 , \16827 );
or \U$16487 ( \16830 , \16825 , \16828 , \16829 );
and \U$16488 ( \16831 , \16621 , \16830 );
xor \U$16489 ( \16832 , \16621 , \16830 );
xor \U$16490 ( \16833 , \16819 , \16824 );
xor \U$16491 ( \16834 , \16833 , \16827 );
and \U$16492 ( \16835 , \3478 , \7564 );
and \U$16493 ( \16836 , \3061 , \7562 );
nor \U$16494 ( \16837 , \16835 , \16836 );
xnor \U$16495 ( \16838 , \16837 , \7315 );
and \U$16496 ( \16839 , \3808 , \7035 );
and \U$16497 ( \16840 , \3686 , \7033 );
nor \U$16498 ( \16841 , \16839 , \16840 );
xnor \U$16499 ( \16842 , \16841 , \6775 );
and \U$16500 ( \16843 , \16838 , \16842 );
and \U$16501 ( \16844 , \4069 , \6541 );
and \U$16502 ( \16845 , \3813 , \6539 );
nor \U$16503 ( \16846 , \16844 , \16845 );
xnor \U$16504 ( \16847 , \16846 , \6226 );
and \U$16505 ( \16848 , \16842 , \16847 );
and \U$16506 ( \16849 , \16838 , \16847 );
or \U$16507 ( \16850 , \16843 , \16848 , \16849 );
and \U$16508 ( \16851 , \2438 , \9230 );
and \U$16509 ( \16852 , \2174 , \9228 );
nor \U$16510 ( \16853 , \16851 , \16852 );
xnor \U$16511 ( \16854 , \16853 , \8920 );
and \U$16512 ( \16855 , \2637 , \8693 );
and \U$16513 ( \16856 , \2463 , \8691 );
nor \U$16514 ( \16857 , \16855 , \16856 );
xnor \U$16515 ( \16858 , \16857 , \8322 );
and \U$16516 ( \16859 , \16854 , \16858 );
and \U$16517 ( \16860 , \2942 , \8131 );
and \U$16518 ( \16861 , \2804 , \8129 );
nor \U$16519 ( \16862 , \16860 , \16861 );
xnor \U$16520 ( \16863 , \16862 , \7813 );
and \U$16521 ( \16864 , \16858 , \16863 );
and \U$16522 ( \16865 , \16854 , \16863 );
or \U$16523 ( \16866 , \16859 , \16864 , \16865 );
and \U$16524 ( \16867 , \16850 , \16866 );
and \U$16525 ( \16868 , \1839 , \10611 );
and \U$16526 ( \16869 , \1596 , \10608 );
nor \U$16527 ( \16870 , \16868 , \16869 );
xnor \U$16528 ( \16871 , \16870 , \9556 );
and \U$16529 ( \16872 , \2030 , \9798 );
and \U$16530 ( \16873 , \1844 , \9796 );
nor \U$16531 ( \16874 , \16872 , \16873 );
xnor \U$16532 ( \16875 , \16874 , \9559 );
and \U$16533 ( \16876 , \16871 , \16875 );
and \U$16534 ( \16877 , \16875 , \1467 );
and \U$16535 ( \16878 , \16871 , \1467 );
or \U$16536 ( \16879 , \16876 , \16877 , \16878 );
and \U$16537 ( \16880 , \16866 , \16879 );
and \U$16538 ( \16881 , \16850 , \16879 );
or \U$16539 ( \16882 , \16867 , \16880 , \16881 );
and \U$16540 ( \16883 , \7500 , \3434 );
and \U$16541 ( \16884 , \6974 , \3432 );
nor \U$16542 ( \16885 , \16883 , \16884 );
xnor \U$16543 ( \16886 , \16885 , \3247 );
and \U$16544 ( \16887 , \8170 , \3121 );
and \U$16545 ( \16888 , \7924 , \3119 );
nor \U$16546 ( \16889 , \16887 , \16888 );
xnor \U$16547 ( \16890 , \16889 , \2916 );
and \U$16548 ( \16891 , \16886 , \16890 );
and \U$16549 ( \16892 , \8494 , \2715 );
and \U$16550 ( \16893 , \8175 , \2713 );
nor \U$16551 ( \16894 , \16892 , \16893 );
xnor \U$16552 ( \16895 , \16894 , \2566 );
and \U$16553 ( \16896 , \16890 , \16895 );
and \U$16554 ( \16897 , \16886 , \16895 );
or \U$16555 ( \16898 , \16891 , \16896 , \16897 );
and \U$16556 ( \16899 , \4568 , \6032 );
and \U$16557 ( \16900 , \4266 , \6030 );
nor \U$16558 ( \16901 , \16899 , \16900 );
xnor \U$16559 ( \16902 , \16901 , \5692 );
and \U$16560 ( \16903 , \5045 , \5443 );
and \U$16561 ( \16904 , \4576 , \5441 );
nor \U$16562 ( \16905 , \16903 , \16904 );
xnor \U$16563 ( \16906 , \16905 , \5202 );
and \U$16564 ( \16907 , \16902 , \16906 );
and \U$16565 ( \16908 , \5314 , \4977 );
and \U$16566 ( \16909 , \5050 , \4975 );
nor \U$16567 ( \16910 , \16908 , \16909 );
xnor \U$16568 ( \16911 , \16910 , \4789 );
and \U$16569 ( \16912 , \16906 , \16911 );
and \U$16570 ( \16913 , \16902 , \16911 );
or \U$16571 ( \16914 , \16907 , \16912 , \16913 );
and \U$16572 ( \16915 , \16898 , \16914 );
and \U$16573 ( \16916 , \5945 , \4603 );
and \U$16574 ( \16917 , \5573 , \4601 );
nor \U$16575 ( \16918 , \16916 , \16917 );
xnor \U$16576 ( \16919 , \16918 , \4371 );
and \U$16577 ( \16920 , \6297 , \4152 );
and \U$16578 ( \16921 , \5954 , \4150 );
nor \U$16579 ( \16922 , \16920 , \16921 );
xnor \U$16580 ( \16923 , \16922 , \4009 );
and \U$16581 ( \16924 , \16919 , \16923 );
and \U$16582 ( \16925 , \6802 , \3829 );
and \U$16583 ( \16926 , \6499 , \3827 );
nor \U$16584 ( \16927 , \16925 , \16926 );
xnor \U$16585 ( \16928 , \16927 , \3583 );
and \U$16586 ( \16929 , \16923 , \16928 );
and \U$16587 ( \16930 , \16919 , \16928 );
or \U$16588 ( \16931 , \16924 , \16929 , \16930 );
and \U$16589 ( \16932 , \16914 , \16931 );
and \U$16590 ( \16933 , \16898 , \16931 );
or \U$16591 ( \16934 , \16915 , \16932 , \16933 );
and \U$16592 ( \16935 , \16882 , \16934 );
and \U$16593 ( \16936 , \9347 , \2393 );
and \U$16594 ( \16937 , \8778 , \2391 );
nor \U$16595 ( \16938 , \16936 , \16937 );
xnor \U$16596 ( \16939 , \16938 , \2251 );
and \U$16597 ( \16940 , \9958 , \2097 );
and \U$16598 ( \16941 , \9355 , \2095 );
nor \U$16599 ( \16942 , \16940 , \16941 );
xnor \U$16600 ( \16943 , \16942 , \1960 );
and \U$16601 ( \16944 , \16939 , \16943 );
and \U$16602 ( \16945 , \10144 , \1891 );
and \U$16603 ( \16946 , \9963 , \1889 );
nor \U$16604 ( \16947 , \16945 , \16946 );
xnor \U$16605 ( \16948 , \16947 , \1739 );
and \U$16606 ( \16949 , \16943 , \16948 );
and \U$16607 ( \16950 , \16939 , \16948 );
or \U$16608 ( \16951 , \16944 , \16949 , \16950 );
xor \U$16609 ( \16952 , \16641 , \16645 );
xor \U$16610 ( \16953 , \16952 , \16650 );
and \U$16611 ( \16954 , \16951 , \16953 );
xor \U$16612 ( \16955 , \16730 , \16734 );
xor \U$16613 ( \16956 , \16955 , \16739 );
and \U$16614 ( \16957 , \16953 , \16956 );
and \U$16615 ( \16958 , \16951 , \16956 );
or \U$16616 ( \16959 , \16954 , \16957 , \16958 );
and \U$16617 ( \16960 , \16934 , \16959 );
and \U$16618 ( \16961 , \16882 , \16959 );
or \U$16619 ( \16962 , \16935 , \16960 , \16961 );
xor \U$16620 ( \16963 , \16625 , \16629 );
xor \U$16621 ( \16964 , \16963 , \16634 );
xor \U$16622 ( \16965 , \16677 , \16681 );
xor \U$16623 ( \16966 , \16965 , \16686 );
and \U$16624 ( \16967 , \16964 , \16966 );
xor \U$16625 ( \16968 , \16658 , \16662 );
xor \U$16626 ( \16969 , \16968 , \16667 );
and \U$16627 ( \16970 , \16966 , \16969 );
and \U$16628 ( \16971 , \16964 , \16969 );
or \U$16629 ( \16972 , \16967 , \16970 , \16971 );
xor \U$16630 ( \16973 , \16693 , \16697 );
xor \U$16631 ( \16974 , \16973 , \16702 );
xor \U$16632 ( \16975 , \16710 , \16714 );
xor \U$16633 ( \16976 , \16975 , \16719 );
and \U$16634 ( \16977 , \16974 , \16976 );
and \U$16635 ( \16978 , \16972 , \16977 );
xor \U$16636 ( \16979 , \16754 , \16756 );
xor \U$16637 ( \16980 , \16979 , \16759 );
and \U$16638 ( \16981 , \16977 , \16980 );
and \U$16639 ( \16982 , \16972 , \16980 );
or \U$16640 ( \16983 , \16978 , \16981 , \16982 );
and \U$16641 ( \16984 , \16962 , \16983 );
xor \U$16642 ( \16985 , \16637 , \16653 );
xor \U$16643 ( \16986 , \16985 , \16670 );
xor \U$16644 ( \16987 , \16764 , \16766 );
xor \U$16645 ( \16988 , \16987 , \16769 );
and \U$16646 ( \16989 , \16986 , \16988 );
xor \U$16647 ( \16990 , \16742 , \16744 );
xor \U$16648 ( \16991 , \16990 , \16746 );
and \U$16649 ( \16992 , \16988 , \16991 );
and \U$16650 ( \16993 , \16986 , \16991 );
or \U$16651 ( \16994 , \16989 , \16992 , \16993 );
and \U$16652 ( \16995 , \16983 , \16994 );
and \U$16653 ( \16996 , \16962 , \16994 );
or \U$16654 ( \16997 , \16984 , \16995 , \16996 );
xor \U$16655 ( \16998 , \16426 , \16442 );
xor \U$16656 ( \16999 , \16998 , \16459 );
xor \U$16657 ( \17000 , \16474 , \16490 );
xor \U$16658 ( \17001 , \17000 , \16507 );
and \U$16659 ( \17002 , \16999 , \17001 );
xor \U$16660 ( \17003 , \16781 , \16783 );
xor \U$16661 ( \17004 , \17003 , \16786 );
and \U$16662 ( \17005 , \17001 , \17004 );
and \U$16663 ( \17006 , \16999 , \17004 );
or \U$16664 ( \17007 , \17002 , \17005 , \17006 );
and \U$16665 ( \17008 , \16997 , \17007 );
xor \U$16666 ( \17009 , \16462 , \16510 );
xor \U$16667 ( \17010 , \17009 , \16542 );
and \U$16668 ( \17011 , \17007 , \17010 );
and \U$16669 ( \17012 , \16997 , \17010 );
or \U$16670 ( \17013 , \17008 , \17011 , \17012 );
xor \U$16671 ( \17014 , \16792 , \16802 );
xor \U$16672 ( \17015 , \17014 , \16805 );
and \U$16673 ( \17016 , \17013 , \17015 );
xor \U$16674 ( \17017 , \16810 , \16812 );
and \U$16675 ( \17018 , \17015 , \17017 );
and \U$16676 ( \17019 , \17013 , \17017 );
or \U$16677 ( \17020 , \17016 , \17018 , \17019 );
xor \U$16678 ( \17021 , \16808 , \16813 );
xor \U$16679 ( \17022 , \17021 , \16816 );
and \U$16680 ( \17023 , \17020 , \17022 );
xor \U$16681 ( \17024 , \16821 , \16823 );
and \U$16682 ( \17025 , \17022 , \17024 );
and \U$16683 ( \17026 , \17020 , \17024 );
or \U$16684 ( \17027 , \17023 , \17025 , \17026 );
and \U$16685 ( \17028 , \16834 , \17027 );
xor \U$16686 ( \17029 , \16834 , \17027 );
xor \U$16687 ( \17030 , \17020 , \17022 );
xor \U$16688 ( \17031 , \17030 , \17024 );
and \U$16689 ( \17032 , \1844 , \10611 );
and \U$16690 ( \17033 , \1839 , \10608 );
nor \U$16691 ( \17034 , \17032 , \17033 );
xnor \U$16692 ( \17035 , \17034 , \9556 );
and \U$16693 ( \17036 , \2174 , \9798 );
and \U$16694 ( \17037 , \2030 , \9796 );
nor \U$16695 ( \17038 , \17036 , \17037 );
xnor \U$16696 ( \17039 , \17038 , \9559 );
and \U$16697 ( \17040 , \17035 , \17039 );
and \U$16698 ( \17041 , \2463 , \9230 );
and \U$16699 ( \17042 , \2438 , \9228 );
nor \U$16700 ( \17043 , \17041 , \17042 );
xnor \U$16701 ( \17044 , \17043 , \8920 );
and \U$16702 ( \17045 , \17039 , \17044 );
and \U$16703 ( \17046 , \17035 , \17044 );
or \U$16704 ( \17047 , \17040 , \17045 , \17046 );
and \U$16705 ( \17048 , \2804 , \8693 );
and \U$16706 ( \17049 , \2637 , \8691 );
nor \U$16707 ( \17050 , \17048 , \17049 );
xnor \U$16708 ( \17051 , \17050 , \8322 );
and \U$16709 ( \17052 , \3061 , \8131 );
and \U$16710 ( \17053 , \2942 , \8129 );
nor \U$16711 ( \17054 , \17052 , \17053 );
xnor \U$16712 ( \17055 , \17054 , \7813 );
and \U$16713 ( \17056 , \17051 , \17055 );
and \U$16714 ( \17057 , \3686 , \7564 );
and \U$16715 ( \17058 , \3478 , \7562 );
nor \U$16716 ( \17059 , \17057 , \17058 );
xnor \U$16717 ( \17060 , \17059 , \7315 );
and \U$16718 ( \17061 , \17055 , \17060 );
and \U$16719 ( \17062 , \17051 , \17060 );
or \U$16720 ( \17063 , \17056 , \17061 , \17062 );
and \U$16721 ( \17064 , \17047 , \17063 );
and \U$16722 ( \17065 , \3813 , \7035 );
and \U$16723 ( \17066 , \3808 , \7033 );
nor \U$16724 ( \17067 , \17065 , \17066 );
xnor \U$16725 ( \17068 , \17067 , \6775 );
and \U$16726 ( \17069 , \4266 , \6541 );
and \U$16727 ( \17070 , \4069 , \6539 );
nor \U$16728 ( \17071 , \17069 , \17070 );
xnor \U$16729 ( \17072 , \17071 , \6226 );
and \U$16730 ( \17073 , \17068 , \17072 );
and \U$16731 ( \17074 , \4576 , \6032 );
and \U$16732 ( \17075 , \4568 , \6030 );
nor \U$16733 ( \17076 , \17074 , \17075 );
xnor \U$16734 ( \17077 , \17076 , \5692 );
and \U$16735 ( \17078 , \17072 , \17077 );
and \U$16736 ( \17079 , \17068 , \17077 );
or \U$16737 ( \17080 , \17073 , \17078 , \17079 );
and \U$16738 ( \17081 , \17063 , \17080 );
and \U$16739 ( \17082 , \17047 , \17080 );
or \U$16740 ( \17083 , \17064 , \17081 , \17082 );
and \U$16741 ( \17084 , \6499 , \4152 );
and \U$16742 ( \17085 , \6297 , \4150 );
nor \U$16743 ( \17086 , \17084 , \17085 );
xnor \U$16744 ( \17087 , \17086 , \4009 );
and \U$16745 ( \17088 , \6974 , \3829 );
and \U$16746 ( \17089 , \6802 , \3827 );
nor \U$16747 ( \17090 , \17088 , \17089 );
xnor \U$16748 ( \17091 , \17090 , \3583 );
and \U$16749 ( \17092 , \17087 , \17091 );
and \U$16750 ( \17093 , \7924 , \3434 );
and \U$16751 ( \17094 , \7500 , \3432 );
nor \U$16752 ( \17095 , \17093 , \17094 );
xnor \U$16753 ( \17096 , \17095 , \3247 );
and \U$16754 ( \17097 , \17091 , \17096 );
and \U$16755 ( \17098 , \17087 , \17096 );
or \U$16756 ( \17099 , \17092 , \17097 , \17098 );
and \U$16757 ( \17100 , \5050 , \5443 );
and \U$16758 ( \17101 , \5045 , \5441 );
nor \U$16759 ( \17102 , \17100 , \17101 );
xnor \U$16760 ( \17103 , \17102 , \5202 );
and \U$16761 ( \17104 , \5573 , \4977 );
and \U$16762 ( \17105 , \5314 , \4975 );
nor \U$16763 ( \17106 , \17104 , \17105 );
xnor \U$16764 ( \17107 , \17106 , \4789 );
and \U$16765 ( \17108 , \17103 , \17107 );
and \U$16766 ( \17109 , \5954 , \4603 );
and \U$16767 ( \17110 , \5945 , \4601 );
nor \U$16768 ( \17111 , \17109 , \17110 );
xnor \U$16769 ( \17112 , \17111 , \4371 );
and \U$16770 ( \17113 , \17107 , \17112 );
and \U$16771 ( \17114 , \17103 , \17112 );
or \U$16772 ( \17115 , \17108 , \17113 , \17114 );
and \U$16773 ( \17116 , \17099 , \17115 );
and \U$16774 ( \17117 , \8175 , \3121 );
and \U$16775 ( \17118 , \8170 , \3119 );
nor \U$16776 ( \17119 , \17117 , \17118 );
xnor \U$16777 ( \17120 , \17119 , \2916 );
and \U$16778 ( \17121 , \8778 , \2715 );
and \U$16779 ( \17122 , \8494 , \2713 );
nor \U$16780 ( \17123 , \17121 , \17122 );
xnor \U$16781 ( \17124 , \17123 , \2566 );
and \U$16782 ( \17125 , \17120 , \17124 );
and \U$16783 ( \17126 , \9355 , \2393 );
and \U$16784 ( \17127 , \9347 , \2391 );
nor \U$16785 ( \17128 , \17126 , \17127 );
xnor \U$16786 ( \17129 , \17128 , \2251 );
and \U$16787 ( \17130 , \17124 , \17129 );
and \U$16788 ( \17131 , \17120 , \17129 );
or \U$16789 ( \17132 , \17125 , \17130 , \17131 );
and \U$16790 ( \17133 , \17115 , \17132 );
and \U$16791 ( \17134 , \17099 , \17132 );
or \U$16792 ( \17135 , \17116 , \17133 , \17134 );
and \U$16793 ( \17136 , \17083 , \17135 );
nand \U$16794 ( \17137 , \10764 , \1621 );
xnor \U$16795 ( \17138 , \17137 , \1467 );
xor \U$16796 ( \17139 , \16886 , \16890 );
xor \U$16797 ( \17140 , \17139 , \16895 );
and \U$16798 ( \17141 , \17138 , \17140 );
xor \U$16799 ( \17142 , \16939 , \16943 );
xor \U$16800 ( \17143 , \17142 , \16948 );
and \U$16801 ( \17144 , \17140 , \17143 );
and \U$16802 ( \17145 , \17138 , \17143 );
or \U$16803 ( \17146 , \17141 , \17144 , \17145 );
and \U$16804 ( \17147 , \17135 , \17146 );
and \U$16805 ( \17148 , \17083 , \17146 );
or \U$16806 ( \17149 , \17136 , \17147 , \17148 );
xor \U$16807 ( \17150 , \16850 , \16866 );
xor \U$16808 ( \17151 , \17150 , \16879 );
xor \U$16809 ( \17152 , \16898 , \16914 );
xor \U$16810 ( \17153 , \17152 , \16931 );
and \U$16811 ( \17154 , \17151 , \17153 );
xor \U$16812 ( \17155 , \16951 , \16953 );
xor \U$16813 ( \17156 , \17155 , \16956 );
and \U$16814 ( \17157 , \17153 , \17156 );
and \U$16815 ( \17158 , \17151 , \17156 );
or \U$16816 ( \17159 , \17154 , \17157 , \17158 );
and \U$16817 ( \17160 , \17149 , \17159 );
xor \U$16818 ( \17161 , \16838 , \16842 );
xor \U$16819 ( \17162 , \17161 , \16847 );
xor \U$16820 ( \17163 , \16902 , \16906 );
xor \U$16821 ( \17164 , \17163 , \16911 );
and \U$16822 ( \17165 , \17162 , \17164 );
xor \U$16823 ( \17166 , \16919 , \16923 );
xor \U$16824 ( \17167 , \17166 , \16928 );
and \U$16825 ( \17168 , \17164 , \17167 );
and \U$16826 ( \17169 , \17162 , \17167 );
or \U$16827 ( \17170 , \17165 , \17168 , \17169 );
xor \U$16828 ( \17171 , \16964 , \16966 );
xor \U$16829 ( \17172 , \17171 , \16969 );
and \U$16830 ( \17173 , \17170 , \17172 );
xor \U$16831 ( \17174 , \16974 , \16976 );
and \U$16832 ( \17175 , \17172 , \17174 );
and \U$16833 ( \17176 , \17170 , \17174 );
or \U$16834 ( \17177 , \17173 , \17175 , \17176 );
and \U$16835 ( \17178 , \17159 , \17177 );
and \U$16836 ( \17179 , \17149 , \17177 );
or \U$16837 ( \17180 , \17160 , \17178 , \17179 );
xor \U$16838 ( \17181 , \16689 , \16705 );
xor \U$16839 ( \17182 , \17181 , \16722 );
xor \U$16840 ( \17183 , \16972 , \16977 );
xor \U$16841 ( \17184 , \17183 , \16980 );
and \U$16842 ( \17185 , \17182 , \17184 );
xor \U$16843 ( \17186 , \16986 , \16988 );
xor \U$16844 ( \17187 , \17186 , \16991 );
and \U$16845 ( \17188 , \17184 , \17187 );
and \U$16846 ( \17189 , \17182 , \17187 );
or \U$16847 ( \17190 , \17185 , \17188 , \17189 );
and \U$16848 ( \17191 , \17180 , \17190 );
xor \U$16849 ( \17192 , \16762 , \16772 );
xor \U$16850 ( \17193 , \17192 , \16775 );
and \U$16851 ( \17194 , \17190 , \17193 );
and \U$16852 ( \17195 , \17180 , \17193 );
or \U$16853 ( \17196 , \17191 , \17194 , \17195 );
xor \U$16854 ( \17197 , \16673 , \16725 );
xor \U$16855 ( \17198 , \17197 , \16749 );
xor \U$16856 ( \17199 , \16962 , \16983 );
xor \U$16857 ( \17200 , \17199 , \16994 );
and \U$16858 ( \17201 , \17198 , \17200 );
xor \U$16859 ( \17202 , \16999 , \17001 );
xor \U$16860 ( \17203 , \17202 , \17004 );
and \U$16861 ( \17204 , \17200 , \17203 );
and \U$16862 ( \17205 , \17198 , \17203 );
or \U$16863 ( \17206 , \17201 , \17204 , \17205 );
and \U$16864 ( \17207 , \17196 , \17206 );
xor \U$16865 ( \17208 , \16794 , \16796 );
xor \U$16866 ( \17209 , \17208 , \16799 );
and \U$16867 ( \17210 , \17206 , \17209 );
and \U$16868 ( \17211 , \17196 , \17209 );
or \U$16869 ( \17212 , \17207 , \17210 , \17211 );
xor \U$16870 ( \17213 , \16752 , \16778 );
xor \U$16871 ( \17214 , \17213 , \16789 );
xor \U$16872 ( \17215 , \16997 , \17007 );
xor \U$16873 ( \17216 , \17215 , \17010 );
and \U$16874 ( \17217 , \17214 , \17216 );
and \U$16875 ( \17218 , \17212 , \17217 );
xor \U$16876 ( \17219 , \17013 , \17015 );
xor \U$16877 ( \17220 , \17219 , \17017 );
and \U$16878 ( \17221 , \17217 , \17220 );
and \U$16879 ( \17222 , \17212 , \17220 );
or \U$16880 ( \17223 , \17218 , \17221 , \17222 );
and \U$16881 ( \17224 , \17031 , \17223 );
xor \U$16882 ( \17225 , \17031 , \17223 );
xor \U$16883 ( \17226 , \17212 , \17217 );
xor \U$16884 ( \17227 , \17226 , \17220 );
and \U$16885 ( \17228 , \2030 , \10611 );
and \U$16886 ( \17229 , \1844 , \10608 );
nor \U$16887 ( \17230 , \17228 , \17229 );
xnor \U$16888 ( \17231 , \17230 , \9556 );
and \U$16889 ( \17232 , \2438 , \9798 );
and \U$16890 ( \17233 , \2174 , \9796 );
nor \U$16891 ( \17234 , \17232 , \17233 );
xnor \U$16892 ( \17235 , \17234 , \9559 );
and \U$16893 ( \17236 , \17231 , \17235 );
and \U$16894 ( \17237 , \17235 , \1739 );
and \U$16895 ( \17238 , \17231 , \1739 );
or \U$16896 ( \17239 , \17236 , \17237 , \17238 );
and \U$16897 ( \17240 , \3808 , \7564 );
and \U$16898 ( \17241 , \3686 , \7562 );
nor \U$16899 ( \17242 , \17240 , \17241 );
xnor \U$16900 ( \17243 , \17242 , \7315 );
and \U$16901 ( \17244 , \4069 , \7035 );
and \U$16902 ( \17245 , \3813 , \7033 );
nor \U$16903 ( \17246 , \17244 , \17245 );
xnor \U$16904 ( \17247 , \17246 , \6775 );
and \U$16905 ( \17248 , \17243 , \17247 );
and \U$16906 ( \17249 , \4568 , \6541 );
and \U$16907 ( \17250 , \4266 , \6539 );
nor \U$16908 ( \17251 , \17249 , \17250 );
xnor \U$16909 ( \17252 , \17251 , \6226 );
and \U$16910 ( \17253 , \17247 , \17252 );
and \U$16911 ( \17254 , \17243 , \17252 );
or \U$16912 ( \17255 , \17248 , \17253 , \17254 );
and \U$16913 ( \17256 , \17239 , \17255 );
and \U$16914 ( \17257 , \2637 , \9230 );
and \U$16915 ( \17258 , \2463 , \9228 );
nor \U$16916 ( \17259 , \17257 , \17258 );
xnor \U$16917 ( \17260 , \17259 , \8920 );
and \U$16918 ( \17261 , \2942 , \8693 );
and \U$16919 ( \17262 , \2804 , \8691 );
nor \U$16920 ( \17263 , \17261 , \17262 );
xnor \U$16921 ( \17264 , \17263 , \8322 );
and \U$16922 ( \17265 , \17260 , \17264 );
and \U$16923 ( \17266 , \3478 , \8131 );
and \U$16924 ( \17267 , \3061 , \8129 );
nor \U$16925 ( \17268 , \17266 , \17267 );
xnor \U$16926 ( \17269 , \17268 , \7813 );
and \U$16927 ( \17270 , \17264 , \17269 );
and \U$16928 ( \17271 , \17260 , \17269 );
or \U$16929 ( \17272 , \17265 , \17270 , \17271 );
and \U$16930 ( \17273 , \17255 , \17272 );
and \U$16931 ( \17274 , \17239 , \17272 );
or \U$16932 ( \17275 , \17256 , \17273 , \17274 );
and \U$16933 ( \17276 , \9958 , \2393 );
and \U$16934 ( \17277 , \9355 , \2391 );
nor \U$16935 ( \17278 , \17276 , \17277 );
xnor \U$16936 ( \17279 , \17278 , \2251 );
and \U$16937 ( \17280 , \10144 , \2097 );
and \U$16938 ( \17281 , \9963 , \2095 );
nor \U$16939 ( \17282 , \17280 , \17281 );
xnor \U$16940 ( \17283 , \17282 , \1960 );
and \U$16941 ( \17284 , \17279 , \17283 );
nand \U$16942 ( \17285 , \10764 , \1889 );
xnor \U$16943 ( \17286 , \17285 , \1739 );
and \U$16944 ( \17287 , \17283 , \17286 );
and \U$16945 ( \17288 , \17279 , \17286 );
or \U$16946 ( \17289 , \17284 , \17287 , \17288 );
and \U$16947 ( \17290 , \9963 , \2097 );
and \U$16948 ( \17291 , \9958 , \2095 );
nor \U$16949 ( \17292 , \17290 , \17291 );
xnor \U$16950 ( \17293 , \17292 , \1960 );
and \U$16951 ( \17294 , \17289 , \17293 );
and \U$16952 ( \17295 , \10764 , \1891 );
and \U$16953 ( \17296 , \10144 , \1889 );
nor \U$16954 ( \17297 , \17295 , \17296 );
xnor \U$16955 ( \17298 , \17297 , \1739 );
and \U$16956 ( \17299 , \17293 , \17298 );
and \U$16957 ( \17300 , \17289 , \17298 );
or \U$16958 ( \17301 , \17294 , \17299 , \17300 );
and \U$16959 ( \17302 , \17275 , \17301 );
and \U$16960 ( \17303 , \5045 , \6032 );
and \U$16961 ( \17304 , \4576 , \6030 );
nor \U$16962 ( \17305 , \17303 , \17304 );
xnor \U$16963 ( \17306 , \17305 , \5692 );
and \U$16964 ( \17307 , \5314 , \5443 );
and \U$16965 ( \17308 , \5050 , \5441 );
nor \U$16966 ( \17309 , \17307 , \17308 );
xnor \U$16967 ( \17310 , \17309 , \5202 );
and \U$16968 ( \17311 , \17306 , \17310 );
and \U$16969 ( \17312 , \5945 , \4977 );
and \U$16970 ( \17313 , \5573 , \4975 );
nor \U$16971 ( \17314 , \17312 , \17313 );
xnor \U$16972 ( \17315 , \17314 , \4789 );
and \U$16973 ( \17316 , \17310 , \17315 );
and \U$16974 ( \17317 , \17306 , \17315 );
or \U$16975 ( \17318 , \17311 , \17316 , \17317 );
and \U$16976 ( \17319 , \8170 , \3434 );
and \U$16977 ( \17320 , \7924 , \3432 );
nor \U$16978 ( \17321 , \17319 , \17320 );
xnor \U$16979 ( \17322 , \17321 , \3247 );
and \U$16980 ( \17323 , \8494 , \3121 );
and \U$16981 ( \17324 , \8175 , \3119 );
nor \U$16982 ( \17325 , \17323 , \17324 );
xnor \U$16983 ( \17326 , \17325 , \2916 );
and \U$16984 ( \17327 , \17322 , \17326 );
and \U$16985 ( \17328 , \9347 , \2715 );
and \U$16986 ( \17329 , \8778 , \2713 );
nor \U$16987 ( \17330 , \17328 , \17329 );
xnor \U$16988 ( \17331 , \17330 , \2566 );
and \U$16989 ( \17332 , \17326 , \17331 );
and \U$16990 ( \17333 , \17322 , \17331 );
or \U$16991 ( \17334 , \17327 , \17332 , \17333 );
and \U$16992 ( \17335 , \17318 , \17334 );
and \U$16993 ( \17336 , \6297 , \4603 );
and \U$16994 ( \17337 , \5954 , \4601 );
nor \U$16995 ( \17338 , \17336 , \17337 );
xnor \U$16996 ( \17339 , \17338 , \4371 );
and \U$16997 ( \17340 , \6802 , \4152 );
and \U$16998 ( \17341 , \6499 , \4150 );
nor \U$16999 ( \17342 , \17340 , \17341 );
xnor \U$17000 ( \17343 , \17342 , \4009 );
and \U$17001 ( \17344 , \17339 , \17343 );
and \U$17002 ( \17345 , \7500 , \3829 );
and \U$17003 ( \17346 , \6974 , \3827 );
nor \U$17004 ( \17347 , \17345 , \17346 );
xnor \U$17005 ( \17348 , \17347 , \3583 );
and \U$17006 ( \17349 , \17343 , \17348 );
and \U$17007 ( \17350 , \17339 , \17348 );
or \U$17008 ( \17351 , \17344 , \17349 , \17350 );
and \U$17009 ( \17352 , \17334 , \17351 );
and \U$17010 ( \17353 , \17318 , \17351 );
or \U$17011 ( \17354 , \17335 , \17352 , \17353 );
and \U$17012 ( \17355 , \17301 , \17354 );
and \U$17013 ( \17356 , \17275 , \17354 );
or \U$17014 ( \17357 , \17302 , \17355 , \17356 );
xor \U$17015 ( \17358 , \17035 , \17039 );
xor \U$17016 ( \17359 , \17358 , \17044 );
xor \U$17017 ( \17360 , \17051 , \17055 );
xor \U$17018 ( \17361 , \17360 , \17060 );
and \U$17019 ( \17362 , \17359 , \17361 );
xor \U$17020 ( \17363 , \17068 , \17072 );
xor \U$17021 ( \17364 , \17363 , \17077 );
and \U$17022 ( \17365 , \17361 , \17364 );
and \U$17023 ( \17366 , \17359 , \17364 );
or \U$17024 ( \17367 , \17362 , \17365 , \17366 );
xor \U$17025 ( \17368 , \17087 , \17091 );
xor \U$17026 ( \17369 , \17368 , \17096 );
xor \U$17027 ( \17370 , \17103 , \17107 );
xor \U$17028 ( \17371 , \17370 , \17112 );
and \U$17029 ( \17372 , \17369 , \17371 );
xor \U$17030 ( \17373 , \17120 , \17124 );
xor \U$17031 ( \17374 , \17373 , \17129 );
and \U$17032 ( \17375 , \17371 , \17374 );
and \U$17033 ( \17376 , \17369 , \17374 );
or \U$17034 ( \17377 , \17372 , \17375 , \17376 );
and \U$17035 ( \17378 , \17367 , \17377 );
xor \U$17036 ( \17379 , \16854 , \16858 );
xor \U$17037 ( \17380 , \17379 , \16863 );
and \U$17038 ( \17381 , \17377 , \17380 );
and \U$17039 ( \17382 , \17367 , \17380 );
or \U$17040 ( \17383 , \17378 , \17381 , \17382 );
and \U$17041 ( \17384 , \17357 , \17383 );
xor \U$17042 ( \17385 , \16871 , \16875 );
xor \U$17043 ( \17386 , \17385 , \1467 );
xor \U$17044 ( \17387 , \17162 , \17164 );
xor \U$17045 ( \17388 , \17387 , \17167 );
and \U$17046 ( \17389 , \17386 , \17388 );
xor \U$17047 ( \17390 , \17138 , \17140 );
xor \U$17048 ( \17391 , \17390 , \17143 );
and \U$17049 ( \17392 , \17388 , \17391 );
and \U$17050 ( \17393 , \17386 , \17391 );
or \U$17051 ( \17394 , \17389 , \17392 , \17393 );
and \U$17052 ( \17395 , \17383 , \17394 );
and \U$17053 ( \17396 , \17357 , \17394 );
or \U$17054 ( \17397 , \17384 , \17395 , \17396 );
xor \U$17055 ( \17398 , \17083 , \17135 );
xor \U$17056 ( \17399 , \17398 , \17146 );
xor \U$17057 ( \17400 , \17151 , \17153 );
xor \U$17058 ( \17401 , \17400 , \17156 );
and \U$17059 ( \17402 , \17399 , \17401 );
xor \U$17060 ( \17403 , \17170 , \17172 );
xor \U$17061 ( \17404 , \17403 , \17174 );
and \U$17062 ( \17405 , \17401 , \17404 );
and \U$17063 ( \17406 , \17399 , \17404 );
or \U$17064 ( \17407 , \17402 , \17405 , \17406 );
and \U$17065 ( \17408 , \17397 , \17407 );
xor \U$17066 ( \17409 , \16882 , \16934 );
xor \U$17067 ( \17410 , \17409 , \16959 );
and \U$17068 ( \17411 , \17407 , \17410 );
and \U$17069 ( \17412 , \17397 , \17410 );
or \U$17070 ( \17413 , \17408 , \17411 , \17412 );
xor \U$17071 ( \17414 , \17149 , \17159 );
xor \U$17072 ( \17415 , \17414 , \17177 );
xor \U$17073 ( \17416 , \17182 , \17184 );
xor \U$17074 ( \17417 , \17416 , \17187 );
and \U$17075 ( \17418 , \17415 , \17417 );
and \U$17076 ( \17419 , \17413 , \17418 );
xor \U$17077 ( \17420 , \17198 , \17200 );
xor \U$17078 ( \17421 , \17420 , \17203 );
and \U$17079 ( \17422 , \17418 , \17421 );
and \U$17080 ( \17423 , \17413 , \17421 );
or \U$17081 ( \17424 , \17419 , \17422 , \17423 );
xor \U$17082 ( \17425 , \17196 , \17206 );
xor \U$17083 ( \17426 , \17425 , \17209 );
and \U$17084 ( \17427 , \17424 , \17426 );
xor \U$17085 ( \17428 , \17214 , \17216 );
and \U$17086 ( \17429 , \17426 , \17428 );
and \U$17087 ( \17430 , \17424 , \17428 );
or \U$17088 ( \17431 , \17427 , \17429 , \17430 );
and \U$17089 ( \17432 , \17227 , \17431 );
xor \U$17090 ( \17433 , \17227 , \17431 );
xor \U$17091 ( \17434 , \17424 , \17426 );
xor \U$17092 ( \17435 , \17434 , \17428 );
and \U$17093 ( \17436 , \8778 , \3121 );
and \U$17094 ( \17437 , \8494 , \3119 );
nor \U$17095 ( \17438 , \17436 , \17437 );
xnor \U$17096 ( \17439 , \17438 , \2916 );
and \U$17097 ( \17440 , \9355 , \2715 );
and \U$17098 ( \17441 , \9347 , \2713 );
nor \U$17099 ( \17442 , \17440 , \17441 );
xnor \U$17100 ( \17443 , \17442 , \2566 );
and \U$17101 ( \17444 , \17439 , \17443 );
and \U$17102 ( \17445 , \9963 , \2393 );
and \U$17103 ( \17446 , \9958 , \2391 );
nor \U$17104 ( \17447 , \17445 , \17446 );
xnor \U$17105 ( \17448 , \17447 , \2251 );
and \U$17106 ( \17449 , \17443 , \17448 );
and \U$17107 ( \17450 , \17439 , \17448 );
or \U$17108 ( \17451 , \17444 , \17449 , \17450 );
and \U$17109 ( \17452 , \5573 , \5443 );
and \U$17110 ( \17453 , \5314 , \5441 );
nor \U$17111 ( \17454 , \17452 , \17453 );
xnor \U$17112 ( \17455 , \17454 , \5202 );
and \U$17113 ( \17456 , \5954 , \4977 );
and \U$17114 ( \17457 , \5945 , \4975 );
nor \U$17115 ( \17458 , \17456 , \17457 );
xnor \U$17116 ( \17459 , \17458 , \4789 );
and \U$17117 ( \17460 , \17455 , \17459 );
and \U$17118 ( \17461 , \6499 , \4603 );
and \U$17119 ( \17462 , \6297 , \4601 );
nor \U$17120 ( \17463 , \17461 , \17462 );
xnor \U$17121 ( \17464 , \17463 , \4371 );
and \U$17122 ( \17465 , \17459 , \17464 );
and \U$17123 ( \17466 , \17455 , \17464 );
or \U$17124 ( \17467 , \17460 , \17465 , \17466 );
and \U$17125 ( \17468 , \17451 , \17467 );
and \U$17126 ( \17469 , \6974 , \4152 );
and \U$17127 ( \17470 , \6802 , \4150 );
nor \U$17128 ( \17471 , \17469 , \17470 );
xnor \U$17129 ( \17472 , \17471 , \4009 );
and \U$17130 ( \17473 , \7924 , \3829 );
and \U$17131 ( \17474 , \7500 , \3827 );
nor \U$17132 ( \17475 , \17473 , \17474 );
xnor \U$17133 ( \17476 , \17475 , \3583 );
and \U$17134 ( \17477 , \17472 , \17476 );
and \U$17135 ( \17478 , \8175 , \3434 );
and \U$17136 ( \17479 , \8170 , \3432 );
nor \U$17137 ( \17480 , \17478 , \17479 );
xnor \U$17138 ( \17481 , \17480 , \3247 );
and \U$17139 ( \17482 , \17476 , \17481 );
and \U$17140 ( \17483 , \17472 , \17481 );
or \U$17141 ( \17484 , \17477 , \17482 , \17483 );
and \U$17142 ( \17485 , \17467 , \17484 );
and \U$17143 ( \17486 , \17451 , \17484 );
or \U$17144 ( \17487 , \17468 , \17485 , \17486 );
and \U$17145 ( \17488 , \4266 , \7035 );
and \U$17146 ( \17489 , \4069 , \7033 );
nor \U$17147 ( \17490 , \17488 , \17489 );
xnor \U$17148 ( \17491 , \17490 , \6775 );
and \U$17149 ( \17492 , \4576 , \6541 );
and \U$17150 ( \17493 , \4568 , \6539 );
nor \U$17151 ( \17494 , \17492 , \17493 );
xnor \U$17152 ( \17495 , \17494 , \6226 );
and \U$17153 ( \17496 , \17491 , \17495 );
and \U$17154 ( \17497 , \5050 , \6032 );
and \U$17155 ( \17498 , \5045 , \6030 );
nor \U$17156 ( \17499 , \17497 , \17498 );
xnor \U$17157 ( \17500 , \17499 , \5692 );
and \U$17158 ( \17501 , \17495 , \17500 );
and \U$17159 ( \17502 , \17491 , \17500 );
or \U$17160 ( \17503 , \17496 , \17501 , \17502 );
and \U$17161 ( \17504 , \3061 , \8693 );
and \U$17162 ( \17505 , \2942 , \8691 );
nor \U$17163 ( \17506 , \17504 , \17505 );
xnor \U$17164 ( \17507 , \17506 , \8322 );
and \U$17165 ( \17508 , \3686 , \8131 );
and \U$17166 ( \17509 , \3478 , \8129 );
nor \U$17167 ( \17510 , \17508 , \17509 );
xnor \U$17168 ( \17511 , \17510 , \7813 );
and \U$17169 ( \17512 , \17507 , \17511 );
and \U$17170 ( \17513 , \3813 , \7564 );
and \U$17171 ( \17514 , \3808 , \7562 );
nor \U$17172 ( \17515 , \17513 , \17514 );
xnor \U$17173 ( \17516 , \17515 , \7315 );
and \U$17174 ( \17517 , \17511 , \17516 );
and \U$17175 ( \17518 , \17507 , \17516 );
or \U$17176 ( \17519 , \17512 , \17517 , \17518 );
and \U$17177 ( \17520 , \17503 , \17519 );
and \U$17178 ( \17521 , \2174 , \10611 );
and \U$17179 ( \17522 , \2030 , \10608 );
nor \U$17180 ( \17523 , \17521 , \17522 );
xnor \U$17181 ( \17524 , \17523 , \9556 );
and \U$17182 ( \17525 , \2463 , \9798 );
and \U$17183 ( \17526 , \2438 , \9796 );
nor \U$17184 ( \17527 , \17525 , \17526 );
xnor \U$17185 ( \17528 , \17527 , \9559 );
and \U$17186 ( \17529 , \17524 , \17528 );
and \U$17187 ( \17530 , \2804 , \9230 );
and \U$17188 ( \17531 , \2637 , \9228 );
nor \U$17189 ( \17532 , \17530 , \17531 );
xnor \U$17190 ( \17533 , \17532 , \8920 );
and \U$17191 ( \17534 , \17528 , \17533 );
and \U$17192 ( \17535 , \17524 , \17533 );
or \U$17193 ( \17536 , \17529 , \17534 , \17535 );
and \U$17194 ( \17537 , \17519 , \17536 );
and \U$17195 ( \17538 , \17503 , \17536 );
or \U$17196 ( \17539 , \17520 , \17537 , \17538 );
and \U$17197 ( \17540 , \17487 , \17539 );
xor \U$17198 ( \17541 , \17279 , \17283 );
xor \U$17199 ( \17542 , \17541 , \17286 );
xor \U$17200 ( \17543 , \17322 , \17326 );
xor \U$17201 ( \17544 , \17543 , \17331 );
and \U$17202 ( \17545 , \17542 , \17544 );
xor \U$17203 ( \17546 , \17339 , \17343 );
xor \U$17204 ( \17547 , \17546 , \17348 );
and \U$17205 ( \17548 , \17544 , \17547 );
and \U$17206 ( \17549 , \17542 , \17547 );
or \U$17207 ( \17550 , \17545 , \17548 , \17549 );
and \U$17208 ( \17551 , \17539 , \17550 );
and \U$17209 ( \17552 , \17487 , \17550 );
or \U$17210 ( \17553 , \17540 , \17551 , \17552 );
xor \U$17211 ( \17554 , \17239 , \17255 );
xor \U$17212 ( \17555 , \17554 , \17272 );
xor \U$17213 ( \17556 , \17289 , \17293 );
xor \U$17214 ( \17557 , \17556 , \17298 );
and \U$17215 ( \17558 , \17555 , \17557 );
xor \U$17216 ( \17559 , \17318 , \17334 );
xor \U$17217 ( \17560 , \17559 , \17351 );
and \U$17218 ( \17561 , \17557 , \17560 );
and \U$17219 ( \17562 , \17555 , \17560 );
or \U$17220 ( \17563 , \17558 , \17561 , \17562 );
and \U$17221 ( \17564 , \17553 , \17563 );
xor \U$17222 ( \17565 , \17306 , \17310 );
xor \U$17223 ( \17566 , \17565 , \17315 );
xor \U$17224 ( \17567 , \17243 , \17247 );
xor \U$17225 ( \17568 , \17567 , \17252 );
and \U$17226 ( \17569 , \17566 , \17568 );
xor \U$17227 ( \17570 , \17260 , \17264 );
xor \U$17228 ( \17571 , \17570 , \17269 );
and \U$17229 ( \17572 , \17568 , \17571 );
and \U$17230 ( \17573 , \17566 , \17571 );
or \U$17231 ( \17574 , \17569 , \17572 , \17573 );
xor \U$17232 ( \17575 , \17359 , \17361 );
xor \U$17233 ( \17576 , \17575 , \17364 );
and \U$17234 ( \17577 , \17574 , \17576 );
xor \U$17235 ( \17578 , \17369 , \17371 );
xor \U$17236 ( \17579 , \17578 , \17374 );
and \U$17237 ( \17580 , \17576 , \17579 );
and \U$17238 ( \17581 , \17574 , \17579 );
or \U$17239 ( \17582 , \17577 , \17580 , \17581 );
and \U$17240 ( \17583 , \17563 , \17582 );
and \U$17241 ( \17584 , \17553 , \17582 );
or \U$17242 ( \17585 , \17564 , \17583 , \17584 );
xor \U$17243 ( \17586 , \17047 , \17063 );
xor \U$17244 ( \17587 , \17586 , \17080 );
xor \U$17245 ( \17588 , \17099 , \17115 );
xor \U$17246 ( \17589 , \17588 , \17132 );
and \U$17247 ( \17590 , \17587 , \17589 );
xor \U$17248 ( \17591 , \17386 , \17388 );
xor \U$17249 ( \17592 , \17591 , \17391 );
and \U$17250 ( \17593 , \17589 , \17592 );
and \U$17251 ( \17594 , \17587 , \17592 );
or \U$17252 ( \17595 , \17590 , \17593 , \17594 );
and \U$17253 ( \17596 , \17585 , \17595 );
xor \U$17254 ( \17597 , \17399 , \17401 );
xor \U$17255 ( \17598 , \17597 , \17404 );
and \U$17256 ( \17599 , \17595 , \17598 );
and \U$17257 ( \17600 , \17585 , \17598 );
or \U$17258 ( \17601 , \17596 , \17599 , \17600 );
xor \U$17259 ( \17602 , \17397 , \17407 );
xor \U$17260 ( \17603 , \17602 , \17410 );
and \U$17261 ( \17604 , \17601 , \17603 );
xor \U$17262 ( \17605 , \17415 , \17417 );
and \U$17263 ( \17606 , \17603 , \17605 );
and \U$17264 ( \17607 , \17601 , \17605 );
or \U$17265 ( \17608 , \17604 , \17606 , \17607 );
xor \U$17266 ( \17609 , \17180 , \17190 );
xor \U$17267 ( \17610 , \17609 , \17193 );
and \U$17268 ( \17611 , \17608 , \17610 );
xor \U$17269 ( \17612 , \17413 , \17418 );
xor \U$17270 ( \17613 , \17612 , \17421 );
and \U$17271 ( \17614 , \17610 , \17613 );
and \U$17272 ( \17615 , \17608 , \17613 );
or \U$17273 ( \17616 , \17611 , \17614 , \17615 );
and \U$17274 ( \17617 , \17435 , \17616 );
xor \U$17275 ( \17618 , \17435 , \17616 );
xor \U$17276 ( \17619 , \17608 , \17610 );
xor \U$17277 ( \17620 , \17619 , \17613 );
and \U$17278 ( \17621 , \4069 , \7564 );
and \U$17279 ( \17622 , \3813 , \7562 );
nor \U$17280 ( \17623 , \17621 , \17622 );
xnor \U$17281 ( \17624 , \17623 , \7315 );
and \U$17282 ( \17625 , \4568 , \7035 );
and \U$17283 ( \17626 , \4266 , \7033 );
nor \U$17284 ( \17627 , \17625 , \17626 );
xnor \U$17285 ( \17628 , \17627 , \6775 );
and \U$17286 ( \17629 , \17624 , \17628 );
and \U$17287 ( \17630 , \5045 , \6541 );
and \U$17288 ( \17631 , \4576 , \6539 );
nor \U$17289 ( \17632 , \17630 , \17631 );
xnor \U$17290 ( \17633 , \17632 , \6226 );
and \U$17291 ( \17634 , \17628 , \17633 );
and \U$17292 ( \17635 , \17624 , \17633 );
or \U$17293 ( \17636 , \17629 , \17634 , \17635 );
and \U$17294 ( \17637 , \2942 , \9230 );
and \U$17295 ( \17638 , \2804 , \9228 );
nor \U$17296 ( \17639 , \17637 , \17638 );
xnor \U$17297 ( \17640 , \17639 , \8920 );
and \U$17298 ( \17641 , \3478 , \8693 );
and \U$17299 ( \17642 , \3061 , \8691 );
nor \U$17300 ( \17643 , \17641 , \17642 );
xnor \U$17301 ( \17644 , \17643 , \8322 );
and \U$17302 ( \17645 , \17640 , \17644 );
and \U$17303 ( \17646 , \3808 , \8131 );
and \U$17304 ( \17647 , \3686 , \8129 );
nor \U$17305 ( \17648 , \17646 , \17647 );
xnor \U$17306 ( \17649 , \17648 , \7813 );
and \U$17307 ( \17650 , \17644 , \17649 );
and \U$17308 ( \17651 , \17640 , \17649 );
or \U$17309 ( \17652 , \17645 , \17650 , \17651 );
and \U$17310 ( \17653 , \17636 , \17652 );
and \U$17311 ( \17654 , \2438 , \10611 );
and \U$17312 ( \17655 , \2174 , \10608 );
nor \U$17313 ( \17656 , \17654 , \17655 );
xnor \U$17314 ( \17657 , \17656 , \9556 );
and \U$17315 ( \17658 , \2637 , \9798 );
and \U$17316 ( \17659 , \2463 , \9796 );
nor \U$17317 ( \17660 , \17658 , \17659 );
xnor \U$17318 ( \17661 , \17660 , \9559 );
and \U$17319 ( \17662 , \17657 , \17661 );
and \U$17320 ( \17663 , \17661 , \1960 );
and \U$17321 ( \17664 , \17657 , \1960 );
or \U$17322 ( \17665 , \17662 , \17663 , \17664 );
and \U$17323 ( \17666 , \17652 , \17665 );
and \U$17324 ( \17667 , \17636 , \17665 );
or \U$17325 ( \17668 , \17653 , \17666 , \17667 );
and \U$17326 ( \17669 , \8494 , \3434 );
and \U$17327 ( \17670 , \8175 , \3432 );
nor \U$17328 ( \17671 , \17669 , \17670 );
xnor \U$17329 ( \17672 , \17671 , \3247 );
and \U$17330 ( \17673 , \9347 , \3121 );
and \U$17331 ( \17674 , \8778 , \3119 );
nor \U$17332 ( \17675 , \17673 , \17674 );
xnor \U$17333 ( \17676 , \17675 , \2916 );
and \U$17334 ( \17677 , \17672 , \17676 );
and \U$17335 ( \17678 , \9958 , \2715 );
and \U$17336 ( \17679 , \9355 , \2713 );
nor \U$17337 ( \17680 , \17678 , \17679 );
xnor \U$17338 ( \17681 , \17680 , \2566 );
and \U$17339 ( \17682 , \17676 , \17681 );
and \U$17340 ( \17683 , \17672 , \17681 );
or \U$17341 ( \17684 , \17677 , \17682 , \17683 );
and \U$17342 ( \17685 , \5314 , \6032 );
and \U$17343 ( \17686 , \5050 , \6030 );
nor \U$17344 ( \17687 , \17685 , \17686 );
xnor \U$17345 ( \17688 , \17687 , \5692 );
and \U$17346 ( \17689 , \5945 , \5443 );
and \U$17347 ( \17690 , \5573 , \5441 );
nor \U$17348 ( \17691 , \17689 , \17690 );
xnor \U$17349 ( \17692 , \17691 , \5202 );
and \U$17350 ( \17693 , \17688 , \17692 );
and \U$17351 ( \17694 , \6297 , \4977 );
and \U$17352 ( \17695 , \5954 , \4975 );
nor \U$17353 ( \17696 , \17694 , \17695 );
xnor \U$17354 ( \17697 , \17696 , \4789 );
and \U$17355 ( \17698 , \17692 , \17697 );
and \U$17356 ( \17699 , \17688 , \17697 );
or \U$17357 ( \17700 , \17693 , \17698 , \17699 );
and \U$17358 ( \17701 , \17684 , \17700 );
and \U$17359 ( \17702 , \6802 , \4603 );
and \U$17360 ( \17703 , \6499 , \4601 );
nor \U$17361 ( \17704 , \17702 , \17703 );
xnor \U$17362 ( \17705 , \17704 , \4371 );
and \U$17363 ( \17706 , \7500 , \4152 );
and \U$17364 ( \17707 , \6974 , \4150 );
nor \U$17365 ( \17708 , \17706 , \17707 );
xnor \U$17366 ( \17709 , \17708 , \4009 );
and \U$17367 ( \17710 , \17705 , \17709 );
and \U$17368 ( \17711 , \8170 , \3829 );
and \U$17369 ( \17712 , \7924 , \3827 );
nor \U$17370 ( \17713 , \17711 , \17712 );
xnor \U$17371 ( \17714 , \17713 , \3583 );
and \U$17372 ( \17715 , \17709 , \17714 );
and \U$17373 ( \17716 , \17705 , \17714 );
or \U$17374 ( \17717 , \17710 , \17715 , \17716 );
and \U$17375 ( \17718 , \17700 , \17717 );
and \U$17376 ( \17719 , \17684 , \17717 );
or \U$17377 ( \17720 , \17701 , \17718 , \17719 );
and \U$17378 ( \17721 , \17668 , \17720 );
and \U$17379 ( \17722 , \10764 , \2097 );
and \U$17380 ( \17723 , \10144 , \2095 );
nor \U$17381 ( \17724 , \17722 , \17723 );
xnor \U$17382 ( \17725 , \17724 , \1960 );
xor \U$17383 ( \17726 , \17439 , \17443 );
xor \U$17384 ( \17727 , \17726 , \17448 );
and \U$17385 ( \17728 , \17725 , \17727 );
xor \U$17386 ( \17729 , \17472 , \17476 );
xor \U$17387 ( \17730 , \17729 , \17481 );
and \U$17388 ( \17731 , \17727 , \17730 );
and \U$17389 ( \17732 , \17725 , \17730 );
or \U$17390 ( \17733 , \17728 , \17731 , \17732 );
and \U$17391 ( \17734 , \17720 , \17733 );
and \U$17392 ( \17735 , \17668 , \17733 );
or \U$17393 ( \17736 , \17721 , \17734 , \17735 );
xor \U$17394 ( \17737 , \17491 , \17495 );
xor \U$17395 ( \17738 , \17737 , \17500 );
xor \U$17396 ( \17739 , \17455 , \17459 );
xor \U$17397 ( \17740 , \17739 , \17464 );
and \U$17398 ( \17741 , \17738 , \17740 );
xor \U$17399 ( \17742 , \17507 , \17511 );
xor \U$17400 ( \17743 , \17742 , \17516 );
and \U$17401 ( \17744 , \17740 , \17743 );
and \U$17402 ( \17745 , \17738 , \17743 );
or \U$17403 ( \17746 , \17741 , \17744 , \17745 );
xor \U$17404 ( \17747 , \17231 , \17235 );
xor \U$17405 ( \17748 , \17747 , \1739 );
and \U$17406 ( \17749 , \17746 , \17748 );
xor \U$17407 ( \17750 , \17566 , \17568 );
xor \U$17408 ( \17751 , \17750 , \17571 );
and \U$17409 ( \17752 , \17748 , \17751 );
and \U$17410 ( \17753 , \17746 , \17751 );
or \U$17411 ( \17754 , \17749 , \17752 , \17753 );
and \U$17412 ( \17755 , \17736 , \17754 );
xor \U$17413 ( \17756 , \17451 , \17467 );
xor \U$17414 ( \17757 , \17756 , \17484 );
xor \U$17415 ( \17758 , \17503 , \17519 );
xor \U$17416 ( \17759 , \17758 , \17536 );
and \U$17417 ( \17760 , \17757 , \17759 );
xor \U$17418 ( \17761 , \17542 , \17544 );
xor \U$17419 ( \17762 , \17761 , \17547 );
and \U$17420 ( \17763 , \17759 , \17762 );
and \U$17421 ( \17764 , \17757 , \17762 );
or \U$17422 ( \17765 , \17760 , \17763 , \17764 );
and \U$17423 ( \17766 , \17754 , \17765 );
and \U$17424 ( \17767 , \17736 , \17765 );
or \U$17425 ( \17768 , \17755 , \17766 , \17767 );
xor \U$17426 ( \17769 , \17487 , \17539 );
xor \U$17427 ( \17770 , \17769 , \17550 );
xor \U$17428 ( \17771 , \17555 , \17557 );
xor \U$17429 ( \17772 , \17771 , \17560 );
and \U$17430 ( \17773 , \17770 , \17772 );
xor \U$17431 ( \17774 , \17574 , \17576 );
xor \U$17432 ( \17775 , \17774 , \17579 );
and \U$17433 ( \17776 , \17772 , \17775 );
and \U$17434 ( \17777 , \17770 , \17775 );
or \U$17435 ( \17778 , \17773 , \17776 , \17777 );
and \U$17436 ( \17779 , \17768 , \17778 );
xor \U$17437 ( \17780 , \17367 , \17377 );
xor \U$17438 ( \17781 , \17780 , \17380 );
and \U$17439 ( \17782 , \17778 , \17781 );
and \U$17440 ( \17783 , \17768 , \17781 );
or \U$17441 ( \17784 , \17779 , \17782 , \17783 );
xor \U$17442 ( \17785 , \17275 , \17301 );
xor \U$17443 ( \17786 , \17785 , \17354 );
xor \U$17444 ( \17787 , \17553 , \17563 );
xor \U$17445 ( \17788 , \17787 , \17582 );
and \U$17446 ( \17789 , \17786 , \17788 );
xor \U$17447 ( \17790 , \17587 , \17589 );
xor \U$17448 ( \17791 , \17790 , \17592 );
and \U$17449 ( \17792 , \17788 , \17791 );
and \U$17450 ( \17793 , \17786 , \17791 );
or \U$17451 ( \17794 , \17789 , \17792 , \17793 );
and \U$17452 ( \17795 , \17784 , \17794 );
xor \U$17453 ( \17796 , \17357 , \17383 );
xor \U$17454 ( \17797 , \17796 , \17394 );
and \U$17455 ( \17798 , \17794 , \17797 );
and \U$17456 ( \17799 , \17784 , \17797 );
or \U$17457 ( \17800 , \17795 , \17798 , \17799 );
xor \U$17458 ( \17801 , \17601 , \17603 );
xor \U$17459 ( \17802 , \17801 , \17605 );
and \U$17460 ( \17803 , \17800 , \17802 );
and \U$17461 ( \17804 , \17620 , \17803 );
xor \U$17462 ( \17805 , \17620 , \17803 );
xor \U$17463 ( \17806 , \17800 , \17802 );
and \U$17464 ( \17807 , \2463 , \10611 );
and \U$17465 ( \17808 , \2438 , \10608 );
nor \U$17466 ( \17809 , \17807 , \17808 );
xnor \U$17467 ( \17810 , \17809 , \9556 );
and \U$17468 ( \17811 , \2804 , \9798 );
and \U$17469 ( \17812 , \2637 , \9796 );
nor \U$17470 ( \17813 , \17811 , \17812 );
xnor \U$17471 ( \17814 , \17813 , \9559 );
and \U$17472 ( \17815 , \17810 , \17814 );
and \U$17473 ( \17816 , \3061 , \9230 );
and \U$17474 ( \17817 , \2942 , \9228 );
nor \U$17475 ( \17818 , \17816 , \17817 );
xnor \U$17476 ( \17819 , \17818 , \8920 );
and \U$17477 ( \17820 , \17814 , \17819 );
and \U$17478 ( \17821 , \17810 , \17819 );
or \U$17479 ( \17822 , \17815 , \17820 , \17821 );
and \U$17480 ( \17823 , \3686 , \8693 );
and \U$17481 ( \17824 , \3478 , \8691 );
nor \U$17482 ( \17825 , \17823 , \17824 );
xnor \U$17483 ( \17826 , \17825 , \8322 );
and \U$17484 ( \17827 , \3813 , \8131 );
and \U$17485 ( \17828 , \3808 , \8129 );
nor \U$17486 ( \17829 , \17827 , \17828 );
xnor \U$17487 ( \17830 , \17829 , \7813 );
and \U$17488 ( \17831 , \17826 , \17830 );
and \U$17489 ( \17832 , \4266 , \7564 );
and \U$17490 ( \17833 , \4069 , \7562 );
nor \U$17491 ( \17834 , \17832 , \17833 );
xnor \U$17492 ( \17835 , \17834 , \7315 );
and \U$17493 ( \17836 , \17830 , \17835 );
and \U$17494 ( \17837 , \17826 , \17835 );
or \U$17495 ( \17838 , \17831 , \17836 , \17837 );
and \U$17496 ( \17839 , \17822 , \17838 );
and \U$17497 ( \17840 , \4576 , \7035 );
and \U$17498 ( \17841 , \4568 , \7033 );
nor \U$17499 ( \17842 , \17840 , \17841 );
xnor \U$17500 ( \17843 , \17842 , \6775 );
and \U$17501 ( \17844 , \5050 , \6541 );
and \U$17502 ( \17845 , \5045 , \6539 );
nor \U$17503 ( \17846 , \17844 , \17845 );
xnor \U$17504 ( \17847 , \17846 , \6226 );
and \U$17505 ( \17848 , \17843 , \17847 );
and \U$17506 ( \17849 , \5573 , \6032 );
and \U$17507 ( \17850 , \5314 , \6030 );
nor \U$17508 ( \17851 , \17849 , \17850 );
xnor \U$17509 ( \17852 , \17851 , \5692 );
and \U$17510 ( \17853 , \17847 , \17852 );
and \U$17511 ( \17854 , \17843 , \17852 );
or \U$17512 ( \17855 , \17848 , \17853 , \17854 );
and \U$17513 ( \17856 , \17838 , \17855 );
and \U$17514 ( \17857 , \17822 , \17855 );
or \U$17515 ( \17858 , \17839 , \17856 , \17857 );
and \U$17516 ( \17859 , \9355 , \3121 );
and \U$17517 ( \17860 , \9347 , \3119 );
nor \U$17518 ( \17861 , \17859 , \17860 );
xnor \U$17519 ( \17862 , \17861 , \2916 );
and \U$17520 ( \17863 , \9963 , \2715 );
and \U$17521 ( \17864 , \9958 , \2713 );
nor \U$17522 ( \17865 , \17863 , \17864 );
xnor \U$17523 ( \17866 , \17865 , \2566 );
and \U$17524 ( \17867 , \17862 , \17866 );
and \U$17525 ( \17868 , \10764 , \2393 );
and \U$17526 ( \17869 , \10144 , \2391 );
nor \U$17527 ( \17870 , \17868 , \17869 );
xnor \U$17528 ( \17871 , \17870 , \2251 );
and \U$17529 ( \17872 , \17866 , \17871 );
and \U$17530 ( \17873 , \17862 , \17871 );
or \U$17531 ( \17874 , \17867 , \17872 , \17873 );
and \U$17532 ( \17875 , \7924 , \4152 );
and \U$17533 ( \17876 , \7500 , \4150 );
nor \U$17534 ( \17877 , \17875 , \17876 );
xnor \U$17535 ( \17878 , \17877 , \4009 );
and \U$17536 ( \17879 , \8175 , \3829 );
and \U$17537 ( \17880 , \8170 , \3827 );
nor \U$17538 ( \17881 , \17879 , \17880 );
xnor \U$17539 ( \17882 , \17881 , \3583 );
and \U$17540 ( \17883 , \17878 , \17882 );
and \U$17541 ( \17884 , \8778 , \3434 );
and \U$17542 ( \17885 , \8494 , \3432 );
nor \U$17543 ( \17886 , \17884 , \17885 );
xnor \U$17544 ( \17887 , \17886 , \3247 );
and \U$17545 ( \17888 , \17882 , \17887 );
and \U$17546 ( \17889 , \17878 , \17887 );
or \U$17547 ( \17890 , \17883 , \17888 , \17889 );
and \U$17548 ( \17891 , \17874 , \17890 );
and \U$17549 ( \17892 , \5954 , \5443 );
and \U$17550 ( \17893 , \5945 , \5441 );
nor \U$17551 ( \17894 , \17892 , \17893 );
xnor \U$17552 ( \17895 , \17894 , \5202 );
and \U$17553 ( \17896 , \6499 , \4977 );
and \U$17554 ( \17897 , \6297 , \4975 );
nor \U$17555 ( \17898 , \17896 , \17897 );
xnor \U$17556 ( \17899 , \17898 , \4789 );
and \U$17557 ( \17900 , \17895 , \17899 );
and \U$17558 ( \17901 , \6974 , \4603 );
and \U$17559 ( \17902 , \6802 , \4601 );
nor \U$17560 ( \17903 , \17901 , \17902 );
xnor \U$17561 ( \17904 , \17903 , \4371 );
and \U$17562 ( \17905 , \17899 , \17904 );
and \U$17563 ( \17906 , \17895 , \17904 );
or \U$17564 ( \17907 , \17900 , \17905 , \17906 );
and \U$17565 ( \17908 , \17890 , \17907 );
and \U$17566 ( \17909 , \17874 , \17907 );
or \U$17567 ( \17910 , \17891 , \17908 , \17909 );
and \U$17568 ( \17911 , \17858 , \17910 );
and \U$17569 ( \17912 , \10144 , \2393 );
and \U$17570 ( \17913 , \9963 , \2391 );
nor \U$17571 ( \17914 , \17912 , \17913 );
xnor \U$17572 ( \17915 , \17914 , \2251 );
nand \U$17573 ( \17916 , \10764 , \2095 );
xnor \U$17574 ( \17917 , \17916 , \1960 );
and \U$17575 ( \17918 , \17915 , \17917 );
xor \U$17576 ( \17919 , \17672 , \17676 );
xor \U$17577 ( \17920 , \17919 , \17681 );
and \U$17578 ( \17921 , \17917 , \17920 );
and \U$17579 ( \17922 , \17915 , \17920 );
or \U$17580 ( \17923 , \17918 , \17921 , \17922 );
and \U$17581 ( \17924 , \17910 , \17923 );
and \U$17582 ( \17925 , \17858 , \17923 );
or \U$17583 ( \17926 , \17911 , \17924 , \17925 );
xor \U$17584 ( \17927 , \17624 , \17628 );
xor \U$17585 ( \17928 , \17927 , \17633 );
xor \U$17586 ( \17929 , \17688 , \17692 );
xor \U$17587 ( \17930 , \17929 , \17697 );
and \U$17588 ( \17931 , \17928 , \17930 );
xor \U$17589 ( \17932 , \17705 , \17709 );
xor \U$17590 ( \17933 , \17932 , \17714 );
and \U$17591 ( \17934 , \17930 , \17933 );
and \U$17592 ( \17935 , \17928 , \17933 );
or \U$17593 ( \17936 , \17931 , \17934 , \17935 );
xor \U$17594 ( \17937 , \17640 , \17644 );
xor \U$17595 ( \17938 , \17937 , \17649 );
xor \U$17596 ( \17939 , \17657 , \17661 );
xor \U$17597 ( \17940 , \17939 , \1960 );
and \U$17598 ( \17941 , \17938 , \17940 );
and \U$17599 ( \17942 , \17936 , \17941 );
xor \U$17600 ( \17943 , \17524 , \17528 );
xor \U$17601 ( \17944 , \17943 , \17533 );
and \U$17602 ( \17945 , \17941 , \17944 );
and \U$17603 ( \17946 , \17936 , \17944 );
or \U$17604 ( \17947 , \17942 , \17945 , \17946 );
and \U$17605 ( \17948 , \17926 , \17947 );
xor \U$17606 ( \17949 , \17684 , \17700 );
xor \U$17607 ( \17950 , \17949 , \17717 );
xor \U$17608 ( \17951 , \17738 , \17740 );
xor \U$17609 ( \17952 , \17951 , \17743 );
and \U$17610 ( \17953 , \17950 , \17952 );
xor \U$17611 ( \17954 , \17725 , \17727 );
xor \U$17612 ( \17955 , \17954 , \17730 );
and \U$17613 ( \17956 , \17952 , \17955 );
and \U$17614 ( \17957 , \17950 , \17955 );
or \U$17615 ( \17958 , \17953 , \17956 , \17957 );
and \U$17616 ( \17959 , \17947 , \17958 );
and \U$17617 ( \17960 , \17926 , \17958 );
or \U$17618 ( \17961 , \17948 , \17959 , \17960 );
xor \U$17619 ( \17962 , \17668 , \17720 );
xor \U$17620 ( \17963 , \17962 , \17733 );
xor \U$17621 ( \17964 , \17746 , \17748 );
xor \U$17622 ( \17965 , \17964 , \17751 );
and \U$17623 ( \17966 , \17963 , \17965 );
xor \U$17624 ( \17967 , \17757 , \17759 );
xor \U$17625 ( \17968 , \17967 , \17762 );
and \U$17626 ( \17969 , \17965 , \17968 );
and \U$17627 ( \17970 , \17963 , \17968 );
or \U$17628 ( \17971 , \17966 , \17969 , \17970 );
and \U$17629 ( \17972 , \17961 , \17971 );
xor \U$17630 ( \17973 , \17770 , \17772 );
xor \U$17631 ( \17974 , \17973 , \17775 );
and \U$17632 ( \17975 , \17971 , \17974 );
and \U$17633 ( \17976 , \17961 , \17974 );
or \U$17634 ( \17977 , \17972 , \17975 , \17976 );
xor \U$17635 ( \17978 , \17768 , \17778 );
xor \U$17636 ( \17979 , \17978 , \17781 );
and \U$17637 ( \17980 , \17977 , \17979 );
xor \U$17638 ( \17981 , \17786 , \17788 );
xor \U$17639 ( \17982 , \17981 , \17791 );
and \U$17640 ( \17983 , \17979 , \17982 );
and \U$17641 ( \17984 , \17977 , \17982 );
or \U$17642 ( \17985 , \17980 , \17983 , \17984 );
xor \U$17643 ( \17986 , \17784 , \17794 );
xor \U$17644 ( \17987 , \17986 , \17797 );
and \U$17645 ( \17988 , \17985 , \17987 );
xor \U$17646 ( \17989 , \17585 , \17595 );
xor \U$17647 ( \17990 , \17989 , \17598 );
and \U$17648 ( \17991 , \17987 , \17990 );
and \U$17649 ( \17992 , \17985 , \17990 );
or \U$17650 ( \17993 , \17988 , \17991 , \17992 );
and \U$17651 ( \17994 , \17806 , \17993 );
xor \U$17652 ( \17995 , \17806 , \17993 );
xor \U$17653 ( \17996 , \17985 , \17987 );
xor \U$17654 ( \17997 , \17996 , \17990 );
and \U$17655 ( \17998 , \2637 , \10611 );
and \U$17656 ( \17999 , \2463 , \10608 );
nor \U$17657 ( \18000 , \17998 , \17999 );
xnor \U$17658 ( \18001 , \18000 , \9556 );
and \U$17659 ( \18002 , \2942 , \9798 );
and \U$17660 ( \18003 , \2804 , \9796 );
nor \U$17661 ( \18004 , \18002 , \18003 );
xnor \U$17662 ( \18005 , \18004 , \9559 );
and \U$17663 ( \18006 , \18001 , \18005 );
and \U$17664 ( \18007 , \18005 , \2251 );
and \U$17665 ( \18008 , \18001 , \2251 );
or \U$17666 ( \18009 , \18006 , \18007 , \18008 );
and \U$17667 ( \18010 , \3478 , \9230 );
and \U$17668 ( \18011 , \3061 , \9228 );
nor \U$17669 ( \18012 , \18010 , \18011 );
xnor \U$17670 ( \18013 , \18012 , \8920 );
and \U$17671 ( \18014 , \3808 , \8693 );
and \U$17672 ( \18015 , \3686 , \8691 );
nor \U$17673 ( \18016 , \18014 , \18015 );
xnor \U$17674 ( \18017 , \18016 , \8322 );
and \U$17675 ( \18018 , \18013 , \18017 );
and \U$17676 ( \18019 , \4069 , \8131 );
and \U$17677 ( \18020 , \3813 , \8129 );
nor \U$17678 ( \18021 , \18019 , \18020 );
xnor \U$17679 ( \18022 , \18021 , \7813 );
and \U$17680 ( \18023 , \18017 , \18022 );
and \U$17681 ( \18024 , \18013 , \18022 );
or \U$17682 ( \18025 , \18018 , \18023 , \18024 );
and \U$17683 ( \18026 , \18009 , \18025 );
and \U$17684 ( \18027 , \4568 , \7564 );
and \U$17685 ( \18028 , \4266 , \7562 );
nor \U$17686 ( \18029 , \18027 , \18028 );
xnor \U$17687 ( \18030 , \18029 , \7315 );
and \U$17688 ( \18031 , \5045 , \7035 );
and \U$17689 ( \18032 , \4576 , \7033 );
nor \U$17690 ( \18033 , \18031 , \18032 );
xnor \U$17691 ( \18034 , \18033 , \6775 );
and \U$17692 ( \18035 , \18030 , \18034 );
and \U$17693 ( \18036 , \5314 , \6541 );
and \U$17694 ( \18037 , \5050 , \6539 );
nor \U$17695 ( \18038 , \18036 , \18037 );
xnor \U$17696 ( \18039 , \18038 , \6226 );
and \U$17697 ( \18040 , \18034 , \18039 );
and \U$17698 ( \18041 , \18030 , \18039 );
or \U$17699 ( \18042 , \18035 , \18040 , \18041 );
and \U$17700 ( \18043 , \18025 , \18042 );
and \U$17701 ( \18044 , \18009 , \18042 );
or \U$17702 ( \18045 , \18026 , \18043 , \18044 );
and \U$17703 ( \18046 , \5945 , \6032 );
and \U$17704 ( \18047 , \5573 , \6030 );
nor \U$17705 ( \18048 , \18046 , \18047 );
xnor \U$17706 ( \18049 , \18048 , \5692 );
and \U$17707 ( \18050 , \6297 , \5443 );
and \U$17708 ( \18051 , \5954 , \5441 );
nor \U$17709 ( \18052 , \18050 , \18051 );
xnor \U$17710 ( \18053 , \18052 , \5202 );
and \U$17711 ( \18054 , \18049 , \18053 );
and \U$17712 ( \18055 , \6802 , \4977 );
and \U$17713 ( \18056 , \6499 , \4975 );
nor \U$17714 ( \18057 , \18055 , \18056 );
xnor \U$17715 ( \18058 , \18057 , \4789 );
and \U$17716 ( \18059 , \18053 , \18058 );
and \U$17717 ( \18060 , \18049 , \18058 );
or \U$17718 ( \18061 , \18054 , \18059 , \18060 );
and \U$17719 ( \18062 , \7500 , \4603 );
and \U$17720 ( \18063 , \6974 , \4601 );
nor \U$17721 ( \18064 , \18062 , \18063 );
xnor \U$17722 ( \18065 , \18064 , \4371 );
and \U$17723 ( \18066 , \8170 , \4152 );
and \U$17724 ( \18067 , \7924 , \4150 );
nor \U$17725 ( \18068 , \18066 , \18067 );
xnor \U$17726 ( \18069 , \18068 , \4009 );
and \U$17727 ( \18070 , \18065 , \18069 );
and \U$17728 ( \18071 , \8494 , \3829 );
and \U$17729 ( \18072 , \8175 , \3827 );
nor \U$17730 ( \18073 , \18071 , \18072 );
xnor \U$17731 ( \18074 , \18073 , \3583 );
and \U$17732 ( \18075 , \18069 , \18074 );
and \U$17733 ( \18076 , \18065 , \18074 );
or \U$17734 ( \18077 , \18070 , \18075 , \18076 );
and \U$17735 ( \18078 , \18061 , \18077 );
and \U$17736 ( \18079 , \9347 , \3434 );
and \U$17737 ( \18080 , \8778 , \3432 );
nor \U$17738 ( \18081 , \18079 , \18080 );
xnor \U$17739 ( \18082 , \18081 , \3247 );
and \U$17740 ( \18083 , \9958 , \3121 );
and \U$17741 ( \18084 , \9355 , \3119 );
nor \U$17742 ( \18085 , \18083 , \18084 );
xnor \U$17743 ( \18086 , \18085 , \2916 );
and \U$17744 ( \18087 , \18082 , \18086 );
and \U$17745 ( \18088 , \10144 , \2715 );
and \U$17746 ( \18089 , \9963 , \2713 );
nor \U$17747 ( \18090 , \18088 , \18089 );
xnor \U$17748 ( \18091 , \18090 , \2566 );
and \U$17749 ( \18092 , \18086 , \18091 );
and \U$17750 ( \18093 , \18082 , \18091 );
or \U$17751 ( \18094 , \18087 , \18092 , \18093 );
and \U$17752 ( \18095 , \18077 , \18094 );
and \U$17753 ( \18096 , \18061 , \18094 );
or \U$17754 ( \18097 , \18078 , \18095 , \18096 );
and \U$17755 ( \18098 , \18045 , \18097 );
xor \U$17756 ( \18099 , \17862 , \17866 );
xor \U$17757 ( \18100 , \18099 , \17871 );
xor \U$17758 ( \18101 , \17878 , \17882 );
xor \U$17759 ( \18102 , \18101 , \17887 );
and \U$17760 ( \18103 , \18100 , \18102 );
xor \U$17761 ( \18104 , \17895 , \17899 );
xor \U$17762 ( \18105 , \18104 , \17904 );
and \U$17763 ( \18106 , \18102 , \18105 );
and \U$17764 ( \18107 , \18100 , \18105 );
or \U$17765 ( \18108 , \18103 , \18106 , \18107 );
and \U$17766 ( \18109 , \18097 , \18108 );
and \U$17767 ( \18110 , \18045 , \18108 );
or \U$17768 ( \18111 , \18098 , \18109 , \18110 );
xor \U$17769 ( \18112 , \17822 , \17838 );
xor \U$17770 ( \18113 , \18112 , \17855 );
xor \U$17771 ( \18114 , \17874 , \17890 );
xor \U$17772 ( \18115 , \18114 , \17907 );
and \U$17773 ( \18116 , \18113 , \18115 );
xor \U$17774 ( \18117 , \17915 , \17917 );
xor \U$17775 ( \18118 , \18117 , \17920 );
and \U$17776 ( \18119 , \18115 , \18118 );
and \U$17777 ( \18120 , \18113 , \18118 );
or \U$17778 ( \18121 , \18116 , \18119 , \18120 );
and \U$17779 ( \18122 , \18111 , \18121 );
xor \U$17780 ( \18123 , \17810 , \17814 );
xor \U$17781 ( \18124 , \18123 , \17819 );
xor \U$17782 ( \18125 , \17826 , \17830 );
xor \U$17783 ( \18126 , \18125 , \17835 );
and \U$17784 ( \18127 , \18124 , \18126 );
xor \U$17785 ( \18128 , \17843 , \17847 );
xor \U$17786 ( \18129 , \18128 , \17852 );
and \U$17787 ( \18130 , \18126 , \18129 );
and \U$17788 ( \18131 , \18124 , \18129 );
or \U$17789 ( \18132 , \18127 , \18130 , \18131 );
xor \U$17790 ( \18133 , \17928 , \17930 );
xor \U$17791 ( \18134 , \18133 , \17933 );
and \U$17792 ( \18135 , \18132 , \18134 );
xor \U$17793 ( \18136 , \17938 , \17940 );
and \U$17794 ( \18137 , \18134 , \18136 );
and \U$17795 ( \18138 , \18132 , \18136 );
or \U$17796 ( \18139 , \18135 , \18137 , \18138 );
and \U$17797 ( \18140 , \18121 , \18139 );
and \U$17798 ( \18141 , \18111 , \18139 );
or \U$17799 ( \18142 , \18122 , \18140 , \18141 );
xor \U$17800 ( \18143 , \17636 , \17652 );
xor \U$17801 ( \18144 , \18143 , \17665 );
xor \U$17802 ( \18145 , \17936 , \17941 );
xor \U$17803 ( \18146 , \18145 , \17944 );
and \U$17804 ( \18147 , \18144 , \18146 );
xor \U$17805 ( \18148 , \17950 , \17952 );
xor \U$17806 ( \18149 , \18148 , \17955 );
and \U$17807 ( \18150 , \18146 , \18149 );
and \U$17808 ( \18151 , \18144 , \18149 );
or \U$17809 ( \18152 , \18147 , \18150 , \18151 );
and \U$17810 ( \18153 , \18142 , \18152 );
xor \U$17811 ( \18154 , \17963 , \17965 );
xor \U$17812 ( \18155 , \18154 , \17968 );
and \U$17813 ( \18156 , \18152 , \18155 );
and \U$17814 ( \18157 , \18142 , \18155 );
or \U$17815 ( \18158 , \18153 , \18156 , \18157 );
xor \U$17816 ( \18159 , \17736 , \17754 );
xor \U$17817 ( \18160 , \18159 , \17765 );
and \U$17818 ( \18161 , \18158 , \18160 );
xor \U$17819 ( \18162 , \17961 , \17971 );
xor \U$17820 ( \18163 , \18162 , \17974 );
and \U$17821 ( \18164 , \18160 , \18163 );
and \U$17822 ( \18165 , \18158 , \18163 );
or \U$17823 ( \18166 , \18161 , \18164 , \18165 );
xor \U$17824 ( \18167 , \17977 , \17979 );
xor \U$17825 ( \18168 , \18167 , \17982 );
and \U$17826 ( \18169 , \18166 , \18168 );
and \U$17827 ( \18170 , \17997 , \18169 );
xor \U$17828 ( \18171 , \17997 , \18169 );
xor \U$17829 ( \18172 , \18166 , \18168 );
and \U$17830 ( \18173 , \5050 , \7035 );
and \U$17831 ( \18174 , \5045 , \7033 );
nor \U$17832 ( \18175 , \18173 , \18174 );
xnor \U$17833 ( \18176 , \18175 , \6775 );
and \U$17834 ( \18177 , \5573 , \6541 );
and \U$17835 ( \18178 , \5314 , \6539 );
nor \U$17836 ( \18179 , \18177 , \18178 );
xnor \U$17837 ( \18180 , \18179 , \6226 );
and \U$17838 ( \18181 , \18176 , \18180 );
and \U$17839 ( \18182 , \5954 , \6032 );
and \U$17840 ( \18183 , \5945 , \6030 );
nor \U$17841 ( \18184 , \18182 , \18183 );
xnor \U$17842 ( \18185 , \18184 , \5692 );
and \U$17843 ( \18186 , \18180 , \18185 );
and \U$17844 ( \18187 , \18176 , \18185 );
or \U$17845 ( \18188 , \18181 , \18186 , \18187 );
and \U$17846 ( \18189 , \2804 , \10611 );
and \U$17847 ( \18190 , \2637 , \10608 );
nor \U$17848 ( \18191 , \18189 , \18190 );
xnor \U$17849 ( \18192 , \18191 , \9556 );
and \U$17850 ( \18193 , \3061 , \9798 );
and \U$17851 ( \18194 , \2942 , \9796 );
nor \U$17852 ( \18195 , \18193 , \18194 );
xnor \U$17853 ( \18196 , \18195 , \9559 );
and \U$17854 ( \18197 , \18192 , \18196 );
and \U$17855 ( \18198 , \3686 , \9230 );
and \U$17856 ( \18199 , \3478 , \9228 );
nor \U$17857 ( \18200 , \18198 , \18199 );
xnor \U$17858 ( \18201 , \18200 , \8920 );
and \U$17859 ( \18202 , \18196 , \18201 );
and \U$17860 ( \18203 , \18192 , \18201 );
or \U$17861 ( \18204 , \18197 , \18202 , \18203 );
and \U$17862 ( \18205 , \18188 , \18204 );
and \U$17863 ( \18206 , \3813 , \8693 );
and \U$17864 ( \18207 , \3808 , \8691 );
nor \U$17865 ( \18208 , \18206 , \18207 );
xnor \U$17866 ( \18209 , \18208 , \8322 );
and \U$17867 ( \18210 , \4266 , \8131 );
and \U$17868 ( \18211 , \4069 , \8129 );
nor \U$17869 ( \18212 , \18210 , \18211 );
xnor \U$17870 ( \18213 , \18212 , \7813 );
and \U$17871 ( \18214 , \18209 , \18213 );
and \U$17872 ( \18215 , \4576 , \7564 );
and \U$17873 ( \18216 , \4568 , \7562 );
nor \U$17874 ( \18217 , \18215 , \18216 );
xnor \U$17875 ( \18218 , \18217 , \7315 );
and \U$17876 ( \18219 , \18213 , \18218 );
and \U$17877 ( \18220 , \18209 , \18218 );
or \U$17878 ( \18221 , \18214 , \18219 , \18220 );
and \U$17879 ( \18222 , \18204 , \18221 );
and \U$17880 ( \18223 , \18188 , \18221 );
or \U$17881 ( \18224 , \18205 , \18222 , \18223 );
and \U$17882 ( \18225 , \8175 , \4152 );
and \U$17883 ( \18226 , \8170 , \4150 );
nor \U$17884 ( \18227 , \18225 , \18226 );
xnor \U$17885 ( \18228 , \18227 , \4009 );
and \U$17886 ( \18229 , \8778 , \3829 );
and \U$17887 ( \18230 , \8494 , \3827 );
nor \U$17888 ( \18231 , \18229 , \18230 );
xnor \U$17889 ( \18232 , \18231 , \3583 );
and \U$17890 ( \18233 , \18228 , \18232 );
and \U$17891 ( \18234 , \9355 , \3434 );
and \U$17892 ( \18235 , \9347 , \3432 );
nor \U$17893 ( \18236 , \18234 , \18235 );
xnor \U$17894 ( \18237 , \18236 , \3247 );
and \U$17895 ( \18238 , \18232 , \18237 );
and \U$17896 ( \18239 , \18228 , \18237 );
or \U$17897 ( \18240 , \18233 , \18238 , \18239 );
and \U$17898 ( \18241 , \6499 , \5443 );
and \U$17899 ( \18242 , \6297 , \5441 );
nor \U$17900 ( \18243 , \18241 , \18242 );
xnor \U$17901 ( \18244 , \18243 , \5202 );
and \U$17902 ( \18245 , \6974 , \4977 );
and \U$17903 ( \18246 , \6802 , \4975 );
nor \U$17904 ( \18247 , \18245 , \18246 );
xnor \U$17905 ( \18248 , \18247 , \4789 );
and \U$17906 ( \18249 , \18244 , \18248 );
and \U$17907 ( \18250 , \7924 , \4603 );
and \U$17908 ( \18251 , \7500 , \4601 );
nor \U$17909 ( \18252 , \18250 , \18251 );
xnor \U$17910 ( \18253 , \18252 , \4371 );
and \U$17911 ( \18254 , \18248 , \18253 );
and \U$17912 ( \18255 , \18244 , \18253 );
or \U$17913 ( \18256 , \18249 , \18254 , \18255 );
and \U$17914 ( \18257 , \18240 , \18256 );
and \U$17915 ( \18258 , \9963 , \3121 );
and \U$17916 ( \18259 , \9958 , \3119 );
nor \U$17917 ( \18260 , \18258 , \18259 );
xnor \U$17918 ( \18261 , \18260 , \2916 );
and \U$17919 ( \18262 , \10764 , \2715 );
and \U$17920 ( \18263 , \10144 , \2713 );
nor \U$17921 ( \18264 , \18262 , \18263 );
xnor \U$17922 ( \18265 , \18264 , \2566 );
and \U$17923 ( \18266 , \18261 , \18265 );
and \U$17924 ( \18267 , \18256 , \18266 );
and \U$17925 ( \18268 , \18240 , \18266 );
or \U$17926 ( \18269 , \18257 , \18267 , \18268 );
and \U$17927 ( \18270 , \18224 , \18269 );
nand \U$17928 ( \18271 , \10764 , \2391 );
xnor \U$17929 ( \18272 , \18271 , \2251 );
xor \U$17930 ( \18273 , \18065 , \18069 );
xor \U$17931 ( \18274 , \18273 , \18074 );
and \U$17932 ( \18275 , \18272 , \18274 );
xor \U$17933 ( \18276 , \18082 , \18086 );
xor \U$17934 ( \18277 , \18276 , \18091 );
and \U$17935 ( \18278 , \18274 , \18277 );
and \U$17936 ( \18279 , \18272 , \18277 );
or \U$17937 ( \18280 , \18275 , \18278 , \18279 );
and \U$17938 ( \18281 , \18269 , \18280 );
and \U$17939 ( \18282 , \18224 , \18280 );
or \U$17940 ( \18283 , \18270 , \18281 , \18282 );
xor \U$17941 ( \18284 , \18013 , \18017 );
xor \U$17942 ( \18285 , \18284 , \18022 );
xor \U$17943 ( \18286 , \18049 , \18053 );
xor \U$17944 ( \18287 , \18286 , \18058 );
and \U$17945 ( \18288 , \18285 , \18287 );
xor \U$17946 ( \18289 , \18030 , \18034 );
xor \U$17947 ( \18290 , \18289 , \18039 );
and \U$17948 ( \18291 , \18287 , \18290 );
and \U$17949 ( \18292 , \18285 , \18290 );
or \U$17950 ( \18293 , \18288 , \18291 , \18292 );
xor \U$17951 ( \18294 , \18100 , \18102 );
xor \U$17952 ( \18295 , \18294 , \18105 );
and \U$17953 ( \18296 , \18293 , \18295 );
xor \U$17954 ( \18297 , \18124 , \18126 );
xor \U$17955 ( \18298 , \18297 , \18129 );
and \U$17956 ( \18299 , \18295 , \18298 );
and \U$17957 ( \18300 , \18293 , \18298 );
or \U$17958 ( \18301 , \18296 , \18299 , \18300 );
and \U$17959 ( \18302 , \18283 , \18301 );
xor \U$17960 ( \18303 , \18009 , \18025 );
xor \U$17961 ( \18304 , \18303 , \18042 );
xor \U$17962 ( \18305 , \18061 , \18077 );
xor \U$17963 ( \18306 , \18305 , \18094 );
and \U$17964 ( \18307 , \18304 , \18306 );
and \U$17965 ( \18308 , \18301 , \18307 );
and \U$17966 ( \18309 , \18283 , \18307 );
or \U$17967 ( \18310 , \18302 , \18308 , \18309 );
xor \U$17968 ( \18311 , \18045 , \18097 );
xor \U$17969 ( \18312 , \18311 , \18108 );
xor \U$17970 ( \18313 , \18113 , \18115 );
xor \U$17971 ( \18314 , \18313 , \18118 );
and \U$17972 ( \18315 , \18312 , \18314 );
xor \U$17973 ( \18316 , \18132 , \18134 );
xor \U$17974 ( \18317 , \18316 , \18136 );
and \U$17975 ( \18318 , \18314 , \18317 );
and \U$17976 ( \18319 , \18312 , \18317 );
or \U$17977 ( \18320 , \18315 , \18318 , \18319 );
and \U$17978 ( \18321 , \18310 , \18320 );
xor \U$17979 ( \18322 , \17858 , \17910 );
xor \U$17980 ( \18323 , \18322 , \17923 );
and \U$17981 ( \18324 , \18320 , \18323 );
and \U$17982 ( \18325 , \18310 , \18323 );
or \U$17983 ( \18326 , \18321 , \18324 , \18325 );
xor \U$17984 ( \18327 , \18111 , \18121 );
xor \U$17985 ( \18328 , \18327 , \18139 );
xor \U$17986 ( \18329 , \18144 , \18146 );
xor \U$17987 ( \18330 , \18329 , \18149 );
and \U$17988 ( \18331 , \18328 , \18330 );
and \U$17989 ( \18332 , \18326 , \18331 );
xor \U$17990 ( \18333 , \17926 , \17947 );
xor \U$17991 ( \18334 , \18333 , \17958 );
and \U$17992 ( \18335 , \18331 , \18334 );
and \U$17993 ( \18336 , \18326 , \18334 );
or \U$17994 ( \18337 , \18332 , \18335 , \18336 );
xor \U$17995 ( \18338 , \18158 , \18160 );
xor \U$17996 ( \18339 , \18338 , \18163 );
and \U$17997 ( \18340 , \18337 , \18339 );
and \U$17998 ( \18341 , \18172 , \18340 );
xor \U$17999 ( \18342 , \18172 , \18340 );
xor \U$18000 ( \18343 , \18337 , \18339 );
xor \U$18001 ( \18344 , \18326 , \18331 );
xor \U$18002 ( \18345 , \18344 , \18334 );
xor \U$18003 ( \18346 , \18142 , \18152 );
xor \U$18004 ( \18347 , \18346 , \18155 );
and \U$18005 ( \18348 , \18345 , \18347 );
and \U$18006 ( \18349 , \18343 , \18348 );
xor \U$18007 ( \18350 , \18343 , \18348 );
xor \U$18008 ( \18351 , \18345 , \18347 );
and \U$18009 ( \18352 , \8170 , \4603 );
and \U$18010 ( \18353 , \7924 , \4601 );
nor \U$18011 ( \18354 , \18352 , \18353 );
xnor \U$18012 ( \18355 , \18354 , \4371 );
and \U$18013 ( \18356 , \8494 , \4152 );
and \U$18014 ( \18357 , \8175 , \4150 );
nor \U$18015 ( \18358 , \18356 , \18357 );
xnor \U$18016 ( \18359 , \18358 , \4009 );
and \U$18017 ( \18360 , \18355 , \18359 );
and \U$18018 ( \18361 , \9347 , \3829 );
and \U$18019 ( \18362 , \8778 , \3827 );
nor \U$18020 ( \18363 , \18361 , \18362 );
xnor \U$18021 ( \18364 , \18363 , \3583 );
and \U$18022 ( \18365 , \18359 , \18364 );
and \U$18023 ( \18366 , \18355 , \18364 );
or \U$18024 ( \18367 , \18360 , \18365 , \18366 );
and \U$18025 ( \18368 , \9958 , \3434 );
and \U$18026 ( \18369 , \9355 , \3432 );
nor \U$18027 ( \18370 , \18368 , \18369 );
xnor \U$18028 ( \18371 , \18370 , \3247 );
and \U$18029 ( \18372 , \10144 , \3121 );
and \U$18030 ( \18373 , \9963 , \3119 );
nor \U$18031 ( \18374 , \18372 , \18373 );
xnor \U$18032 ( \18375 , \18374 , \2916 );
and \U$18033 ( \18376 , \18371 , \18375 );
nand \U$18034 ( \18377 , \10764 , \2713 );
xnor \U$18035 ( \18378 , \18377 , \2566 );
and \U$18036 ( \18379 , \18375 , \18378 );
and \U$18037 ( \18380 , \18371 , \18378 );
or \U$18038 ( \18381 , \18376 , \18379 , \18380 );
and \U$18039 ( \18382 , \18367 , \18381 );
and \U$18040 ( \18383 , \6297 , \6032 );
and \U$18041 ( \18384 , \5954 , \6030 );
nor \U$18042 ( \18385 , \18383 , \18384 );
xnor \U$18043 ( \18386 , \18385 , \5692 );
and \U$18044 ( \18387 , \6802 , \5443 );
and \U$18045 ( \18388 , \6499 , \5441 );
nor \U$18046 ( \18389 , \18387 , \18388 );
xnor \U$18047 ( \18390 , \18389 , \5202 );
and \U$18048 ( \18391 , \18386 , \18390 );
and \U$18049 ( \18392 , \7500 , \4977 );
and \U$18050 ( \18393 , \6974 , \4975 );
nor \U$18051 ( \18394 , \18392 , \18393 );
xnor \U$18052 ( \18395 , \18394 , \4789 );
and \U$18053 ( \18396 , \18390 , \18395 );
and \U$18054 ( \18397 , \18386 , \18395 );
or \U$18055 ( \18398 , \18391 , \18396 , \18397 );
and \U$18056 ( \18399 , \18381 , \18398 );
and \U$18057 ( \18400 , \18367 , \18398 );
or \U$18058 ( \18401 , \18382 , \18399 , \18400 );
and \U$18059 ( \18402 , \5045 , \7564 );
and \U$18060 ( \18403 , \4576 , \7562 );
nor \U$18061 ( \18404 , \18402 , \18403 );
xnor \U$18062 ( \18405 , \18404 , \7315 );
and \U$18063 ( \18406 , \5314 , \7035 );
and \U$18064 ( \18407 , \5050 , \7033 );
nor \U$18065 ( \18408 , \18406 , \18407 );
xnor \U$18066 ( \18409 , \18408 , \6775 );
and \U$18067 ( \18410 , \18405 , \18409 );
and \U$18068 ( \18411 , \5945 , \6541 );
and \U$18069 ( \18412 , \5573 , \6539 );
nor \U$18070 ( \18413 , \18411 , \18412 );
xnor \U$18071 ( \18414 , \18413 , \6226 );
and \U$18072 ( \18415 , \18409 , \18414 );
and \U$18073 ( \18416 , \18405 , \18414 );
or \U$18074 ( \18417 , \18410 , \18415 , \18416 );
and \U$18075 ( \18418 , \2942 , \10611 );
and \U$18076 ( \18419 , \2804 , \10608 );
nor \U$18077 ( \18420 , \18418 , \18419 );
xnor \U$18078 ( \18421 , \18420 , \9556 );
and \U$18079 ( \18422 , \3478 , \9798 );
and \U$18080 ( \18423 , \3061 , \9796 );
nor \U$18081 ( \18424 , \18422 , \18423 );
xnor \U$18082 ( \18425 , \18424 , \9559 );
and \U$18083 ( \18426 , \18421 , \18425 );
and \U$18084 ( \18427 , \18425 , \2566 );
and \U$18085 ( \18428 , \18421 , \2566 );
or \U$18086 ( \18429 , \18426 , \18427 , \18428 );
and \U$18087 ( \18430 , \18417 , \18429 );
and \U$18088 ( \18431 , \3808 , \9230 );
and \U$18089 ( \18432 , \3686 , \9228 );
nor \U$18090 ( \18433 , \18431 , \18432 );
xnor \U$18091 ( \18434 , \18433 , \8920 );
and \U$18092 ( \18435 , \4069 , \8693 );
and \U$18093 ( \18436 , \3813 , \8691 );
nor \U$18094 ( \18437 , \18435 , \18436 );
xnor \U$18095 ( \18438 , \18437 , \8322 );
and \U$18096 ( \18439 , \18434 , \18438 );
and \U$18097 ( \18440 , \4568 , \8131 );
and \U$18098 ( \18441 , \4266 , \8129 );
nor \U$18099 ( \18442 , \18440 , \18441 );
xnor \U$18100 ( \18443 , \18442 , \7813 );
and \U$18101 ( \18444 , \18438 , \18443 );
and \U$18102 ( \18445 , \18434 , \18443 );
or \U$18103 ( \18446 , \18439 , \18444 , \18445 );
and \U$18104 ( \18447 , \18429 , \18446 );
and \U$18105 ( \18448 , \18417 , \18446 );
or \U$18106 ( \18449 , \18430 , \18447 , \18448 );
and \U$18107 ( \18450 , \18401 , \18449 );
xor \U$18108 ( \18451 , \18228 , \18232 );
xor \U$18109 ( \18452 , \18451 , \18237 );
xor \U$18110 ( \18453 , \18244 , \18248 );
xor \U$18111 ( \18454 , \18453 , \18253 );
and \U$18112 ( \18455 , \18452 , \18454 );
xor \U$18113 ( \18456 , \18261 , \18265 );
and \U$18114 ( \18457 , \18454 , \18456 );
and \U$18115 ( \18458 , \18452 , \18456 );
or \U$18116 ( \18459 , \18455 , \18457 , \18458 );
and \U$18117 ( \18460 , \18449 , \18459 );
and \U$18118 ( \18461 , \18401 , \18459 );
or \U$18119 ( \18462 , \18450 , \18460 , \18461 );
xor \U$18120 ( \18463 , \18176 , \18180 );
xor \U$18121 ( \18464 , \18463 , \18185 );
xor \U$18122 ( \18465 , \18192 , \18196 );
xor \U$18123 ( \18466 , \18465 , \18201 );
and \U$18124 ( \18467 , \18464 , \18466 );
xor \U$18125 ( \18468 , \18209 , \18213 );
xor \U$18126 ( \18469 , \18468 , \18218 );
and \U$18127 ( \18470 , \18466 , \18469 );
and \U$18128 ( \18471 , \18464 , \18469 );
or \U$18129 ( \18472 , \18467 , \18470 , \18471 );
xor \U$18130 ( \18473 , \18001 , \18005 );
xor \U$18131 ( \18474 , \18473 , \2251 );
and \U$18132 ( \18475 , \18472 , \18474 );
xor \U$18133 ( \18476 , \18285 , \18287 );
xor \U$18134 ( \18477 , \18476 , \18290 );
and \U$18135 ( \18478 , \18474 , \18477 );
and \U$18136 ( \18479 , \18472 , \18477 );
or \U$18137 ( \18480 , \18475 , \18478 , \18479 );
and \U$18138 ( \18481 , \18462 , \18480 );
xor \U$18139 ( \18482 , \18188 , \18204 );
xor \U$18140 ( \18483 , \18482 , \18221 );
xor \U$18141 ( \18484 , \18240 , \18256 );
xor \U$18142 ( \18485 , \18484 , \18266 );
and \U$18143 ( \18486 , \18483 , \18485 );
xor \U$18144 ( \18487 , \18272 , \18274 );
xor \U$18145 ( \18488 , \18487 , \18277 );
and \U$18146 ( \18489 , \18485 , \18488 );
and \U$18147 ( \18490 , \18483 , \18488 );
or \U$18148 ( \18491 , \18486 , \18489 , \18490 );
and \U$18149 ( \18492 , \18480 , \18491 );
and \U$18150 ( \18493 , \18462 , \18491 );
or \U$18151 ( \18494 , \18481 , \18492 , \18493 );
xor \U$18152 ( \18495 , \18224 , \18269 );
xor \U$18153 ( \18496 , \18495 , \18280 );
xor \U$18154 ( \18497 , \18293 , \18295 );
xor \U$18155 ( \18498 , \18497 , \18298 );
and \U$18156 ( \18499 , \18496 , \18498 );
xor \U$18157 ( \18500 , \18304 , \18306 );
and \U$18158 ( \18501 , \18498 , \18500 );
and \U$18159 ( \18502 , \18496 , \18500 );
or \U$18160 ( \18503 , \18499 , \18501 , \18502 );
and \U$18161 ( \18504 , \18494 , \18503 );
xor \U$18162 ( \18505 , \18312 , \18314 );
xor \U$18163 ( \18506 , \18505 , \18317 );
and \U$18164 ( \18507 , \18503 , \18506 );
and \U$18165 ( \18508 , \18494 , \18506 );
or \U$18166 ( \18509 , \18504 , \18507 , \18508 );
xor \U$18167 ( \18510 , \18310 , \18320 );
xor \U$18168 ( \18511 , \18510 , \18323 );
and \U$18169 ( \18512 , \18509 , \18511 );
xor \U$18170 ( \18513 , \18328 , \18330 );
and \U$18171 ( \18514 , \18511 , \18513 );
and \U$18172 ( \18515 , \18509 , \18513 );
or \U$18173 ( \18516 , \18512 , \18514 , \18515 );
and \U$18174 ( \18517 , \18351 , \18516 );
xor \U$18175 ( \18518 , \18351 , \18516 );
xor \U$18176 ( \18519 , \18509 , \18511 );
xor \U$18177 ( \18520 , \18519 , \18513 );
and \U$18178 ( \18521 , \4266 , \8693 );
and \U$18179 ( \18522 , \4069 , \8691 );
nor \U$18180 ( \18523 , \18521 , \18522 );
xnor \U$18181 ( \18524 , \18523 , \8322 );
and \U$18182 ( \18525 , \4576 , \8131 );
and \U$18183 ( \18526 , \4568 , \8129 );
nor \U$18184 ( \18527 , \18525 , \18526 );
xnor \U$18185 ( \18528 , \18527 , \7813 );
and \U$18186 ( \18529 , \18524 , \18528 );
and \U$18187 ( \18530 , \5050 , \7564 );
and \U$18188 ( \18531 , \5045 , \7562 );
nor \U$18189 ( \18532 , \18530 , \18531 );
xnor \U$18190 ( \18533 , \18532 , \7315 );
and \U$18191 ( \18534 , \18528 , \18533 );
and \U$18192 ( \18535 , \18524 , \18533 );
or \U$18193 ( \18536 , \18529 , \18534 , \18535 );
and \U$18194 ( \18537 , \3061 , \10611 );
and \U$18195 ( \18538 , \2942 , \10608 );
nor \U$18196 ( \18539 , \18537 , \18538 );
xnor \U$18197 ( \18540 , \18539 , \9556 );
and \U$18198 ( \18541 , \3686 , \9798 );
and \U$18199 ( \18542 , \3478 , \9796 );
nor \U$18200 ( \18543 , \18541 , \18542 );
xnor \U$18201 ( \18544 , \18543 , \9559 );
and \U$18202 ( \18545 , \18540 , \18544 );
and \U$18203 ( \18546 , \3813 , \9230 );
and \U$18204 ( \18547 , \3808 , \9228 );
nor \U$18205 ( \18548 , \18546 , \18547 );
xnor \U$18206 ( \18549 , \18548 , \8920 );
and \U$18207 ( \18550 , \18544 , \18549 );
and \U$18208 ( \18551 , \18540 , \18549 );
or \U$18209 ( \18552 , \18545 , \18550 , \18551 );
and \U$18210 ( \18553 , \18536 , \18552 );
and \U$18211 ( \18554 , \5573 , \7035 );
and \U$18212 ( \18555 , \5314 , \7033 );
nor \U$18213 ( \18556 , \18554 , \18555 );
xnor \U$18214 ( \18557 , \18556 , \6775 );
and \U$18215 ( \18558 , \5954 , \6541 );
and \U$18216 ( \18559 , \5945 , \6539 );
nor \U$18217 ( \18560 , \18558 , \18559 );
xnor \U$18218 ( \18561 , \18560 , \6226 );
and \U$18219 ( \18562 , \18557 , \18561 );
and \U$18220 ( \18563 , \6499 , \6032 );
and \U$18221 ( \18564 , \6297 , \6030 );
nor \U$18222 ( \18565 , \18563 , \18564 );
xnor \U$18223 ( \18566 , \18565 , \5692 );
and \U$18224 ( \18567 , \18561 , \18566 );
and \U$18225 ( \18568 , \18557 , \18566 );
or \U$18226 ( \18569 , \18562 , \18567 , \18568 );
and \U$18227 ( \18570 , \18552 , \18569 );
and \U$18228 ( \18571 , \18536 , \18569 );
or \U$18229 ( \18572 , \18553 , \18570 , \18571 );
xor \U$18230 ( \18573 , \18355 , \18359 );
xor \U$18231 ( \18574 , \18573 , \18364 );
xor \U$18232 ( \18575 , \18405 , \18409 );
xor \U$18233 ( \18576 , \18575 , \18414 );
and \U$18234 ( \18577 , \18574 , \18576 );
xor \U$18235 ( \18578 , \18386 , \18390 );
xor \U$18236 ( \18579 , \18578 , \18395 );
and \U$18237 ( \18580 , \18576 , \18579 );
and \U$18238 ( \18581 , \18574 , \18579 );
or \U$18239 ( \18582 , \18577 , \18580 , \18581 );
and \U$18240 ( \18583 , \18572 , \18582 );
and \U$18241 ( \18584 , \6974 , \5443 );
and \U$18242 ( \18585 , \6802 , \5441 );
nor \U$18243 ( \18586 , \18584 , \18585 );
xnor \U$18244 ( \18587 , \18586 , \5202 );
and \U$18245 ( \18588 , \7924 , \4977 );
and \U$18246 ( \18589 , \7500 , \4975 );
nor \U$18247 ( \18590 , \18588 , \18589 );
xnor \U$18248 ( \18591 , \18590 , \4789 );
and \U$18249 ( \18592 , \18587 , \18591 );
and \U$18250 ( \18593 , \8175 , \4603 );
and \U$18251 ( \18594 , \8170 , \4601 );
nor \U$18252 ( \18595 , \18593 , \18594 );
xnor \U$18253 ( \18596 , \18595 , \4371 );
and \U$18254 ( \18597 , \18591 , \18596 );
and \U$18255 ( \18598 , \18587 , \18596 );
or \U$18256 ( \18599 , \18592 , \18597 , \18598 );
and \U$18257 ( \18600 , \8778 , \4152 );
and \U$18258 ( \18601 , \8494 , \4150 );
nor \U$18259 ( \18602 , \18600 , \18601 );
xnor \U$18260 ( \18603 , \18602 , \4009 );
and \U$18261 ( \18604 , \9355 , \3829 );
and \U$18262 ( \18605 , \9347 , \3827 );
nor \U$18263 ( \18606 , \18604 , \18605 );
xnor \U$18264 ( \18607 , \18606 , \3583 );
and \U$18265 ( \18608 , \18603 , \18607 );
and \U$18266 ( \18609 , \9963 , \3434 );
and \U$18267 ( \18610 , \9958 , \3432 );
nor \U$18268 ( \18611 , \18609 , \18610 );
xnor \U$18269 ( \18612 , \18611 , \3247 );
and \U$18270 ( \18613 , \18607 , \18612 );
and \U$18271 ( \18614 , \18603 , \18612 );
or \U$18272 ( \18615 , \18608 , \18613 , \18614 );
and \U$18273 ( \18616 , \18599 , \18615 );
xor \U$18274 ( \18617 , \18371 , \18375 );
xor \U$18275 ( \18618 , \18617 , \18378 );
and \U$18276 ( \18619 , \18615 , \18618 );
and \U$18277 ( \18620 , \18599 , \18618 );
or \U$18278 ( \18621 , \18616 , \18619 , \18620 );
and \U$18279 ( \18622 , \18582 , \18621 );
and \U$18280 ( \18623 , \18572 , \18621 );
or \U$18281 ( \18624 , \18583 , \18622 , \18623 );
xor \U$18282 ( \18625 , \18367 , \18381 );
xor \U$18283 ( \18626 , \18625 , \18398 );
xor \U$18284 ( \18627 , \18464 , \18466 );
xor \U$18285 ( \18628 , \18627 , \18469 );
and \U$18286 ( \18629 , \18626 , \18628 );
xor \U$18287 ( \18630 , \18452 , \18454 );
xor \U$18288 ( \18631 , \18630 , \18456 );
and \U$18289 ( \18632 , \18628 , \18631 );
and \U$18290 ( \18633 , \18626 , \18631 );
or \U$18291 ( \18634 , \18629 , \18632 , \18633 );
and \U$18292 ( \18635 , \18624 , \18634 );
xor \U$18293 ( \18636 , \18483 , \18485 );
xor \U$18294 ( \18637 , \18636 , \18488 );
and \U$18295 ( \18638 , \18634 , \18637 );
and \U$18296 ( \18639 , \18624 , \18637 );
or \U$18297 ( \18640 , \18635 , \18638 , \18639 );
xor \U$18298 ( \18641 , \18462 , \18480 );
xor \U$18299 ( \18642 , \18641 , \18491 );
and \U$18300 ( \18643 , \18640 , \18642 );
xor \U$18301 ( \18644 , \18496 , \18498 );
xor \U$18302 ( \18645 , \18644 , \18500 );
and \U$18303 ( \18646 , \18642 , \18645 );
and \U$18304 ( \18647 , \18640 , \18645 );
or \U$18305 ( \18648 , \18643 , \18646 , \18647 );
xor \U$18306 ( \18649 , \18283 , \18301 );
xor \U$18307 ( \18650 , \18649 , \18307 );
and \U$18308 ( \18651 , \18648 , \18650 );
xor \U$18309 ( \18652 , \18494 , \18503 );
xor \U$18310 ( \18653 , \18652 , \18506 );
and \U$18311 ( \18654 , \18650 , \18653 );
and \U$18312 ( \18655 , \18648 , \18653 );
or \U$18313 ( \18656 , \18651 , \18654 , \18655 );
and \U$18314 ( \18657 , \18520 , \18656 );
xor \U$18315 ( \18658 , \18520 , \18656 );
xor \U$18316 ( \18659 , \18648 , \18650 );
xor \U$18317 ( \18660 , \18659 , \18653 );
and \U$18318 ( \18661 , \4069 , \9230 );
and \U$18319 ( \18662 , \3813 , \9228 );
nor \U$18320 ( \18663 , \18661 , \18662 );
xnor \U$18321 ( \18664 , \18663 , \8920 );
and \U$18322 ( \18665 , \4568 , \8693 );
and \U$18323 ( \18666 , \4266 , \8691 );
nor \U$18324 ( \18667 , \18665 , \18666 );
xnor \U$18325 ( \18668 , \18667 , \8322 );
and \U$18326 ( \18669 , \18664 , \18668 );
and \U$18327 ( \18670 , \5045 , \8131 );
and \U$18328 ( \18671 , \4576 , \8129 );
nor \U$18329 ( \18672 , \18670 , \18671 );
xnor \U$18330 ( \18673 , \18672 , \7813 );
and \U$18331 ( \18674 , \18668 , \18673 );
and \U$18332 ( \18675 , \18664 , \18673 );
or \U$18333 ( \18676 , \18669 , \18674 , \18675 );
and \U$18334 ( \18677 , \5314 , \7564 );
and \U$18335 ( \18678 , \5050 , \7562 );
nor \U$18336 ( \18679 , \18677 , \18678 );
xnor \U$18337 ( \18680 , \18679 , \7315 );
and \U$18338 ( \18681 , \5945 , \7035 );
and \U$18339 ( \18682 , \5573 , \7033 );
nor \U$18340 ( \18683 , \18681 , \18682 );
xnor \U$18341 ( \18684 , \18683 , \6775 );
and \U$18342 ( \18685 , \18680 , \18684 );
and \U$18343 ( \18686 , \6297 , \6541 );
and \U$18344 ( \18687 , \5954 , \6539 );
nor \U$18345 ( \18688 , \18686 , \18687 );
xnor \U$18346 ( \18689 , \18688 , \6226 );
and \U$18347 ( \18690 , \18684 , \18689 );
and \U$18348 ( \18691 , \18680 , \18689 );
or \U$18349 ( \18692 , \18685 , \18690 , \18691 );
and \U$18350 ( \18693 , \18676 , \18692 );
and \U$18351 ( \18694 , \3478 , \10611 );
and \U$18352 ( \18695 , \3061 , \10608 );
nor \U$18353 ( \18696 , \18694 , \18695 );
xnor \U$18354 ( \18697 , \18696 , \9556 );
and \U$18355 ( \18698 , \3808 , \9798 );
and \U$18356 ( \18699 , \3686 , \9796 );
nor \U$18357 ( \18700 , \18698 , \18699 );
xnor \U$18358 ( \18701 , \18700 , \9559 );
and \U$18359 ( \18702 , \18697 , \18701 );
and \U$18360 ( \18703 , \18701 , \2916 );
and \U$18361 ( \18704 , \18697 , \2916 );
or \U$18362 ( \18705 , \18702 , \18703 , \18704 );
and \U$18363 ( \18706 , \18692 , \18705 );
and \U$18364 ( \18707 , \18676 , \18705 );
or \U$18365 ( \18708 , \18693 , \18706 , \18707 );
and \U$18366 ( \18709 , \8494 , \4603 );
and \U$18367 ( \18710 , \8175 , \4601 );
nor \U$18368 ( \18711 , \18709 , \18710 );
xnor \U$18369 ( \18712 , \18711 , \4371 );
and \U$18370 ( \18713 , \9347 , \4152 );
and \U$18371 ( \18714 , \8778 , \4150 );
nor \U$18372 ( \18715 , \18713 , \18714 );
xnor \U$18373 ( \18716 , \18715 , \4009 );
and \U$18374 ( \18717 , \18712 , \18716 );
and \U$18375 ( \18718 , \9958 , \3829 );
and \U$18376 ( \18719 , \9355 , \3827 );
nor \U$18377 ( \18720 , \18718 , \18719 );
xnor \U$18378 ( \18721 , \18720 , \3583 );
and \U$18379 ( \18722 , \18716 , \18721 );
and \U$18380 ( \18723 , \18712 , \18721 );
or \U$18381 ( \18724 , \18717 , \18722 , \18723 );
and \U$18382 ( \18725 , \6802 , \6032 );
and \U$18383 ( \18726 , \6499 , \6030 );
nor \U$18384 ( \18727 , \18725 , \18726 );
xnor \U$18385 ( \18728 , \18727 , \5692 );
and \U$18386 ( \18729 , \7500 , \5443 );
and \U$18387 ( \18730 , \6974 , \5441 );
nor \U$18388 ( \18731 , \18729 , \18730 );
xnor \U$18389 ( \18732 , \18731 , \5202 );
and \U$18390 ( \18733 , \18728 , \18732 );
and \U$18391 ( \18734 , \8170 , \4977 );
and \U$18392 ( \18735 , \7924 , \4975 );
nor \U$18393 ( \18736 , \18734 , \18735 );
xnor \U$18394 ( \18737 , \18736 , \4789 );
and \U$18395 ( \18738 , \18732 , \18737 );
and \U$18396 ( \18739 , \18728 , \18737 );
or \U$18397 ( \18740 , \18733 , \18738 , \18739 );
and \U$18398 ( \18741 , \18724 , \18740 );
and \U$18399 ( \18742 , \10764 , \3121 );
and \U$18400 ( \18743 , \10144 , \3119 );
nor \U$18401 ( \18744 , \18742 , \18743 );
xnor \U$18402 ( \18745 , \18744 , \2916 );
and \U$18403 ( \18746 , \18740 , \18745 );
and \U$18404 ( \18747 , \18724 , \18745 );
or \U$18405 ( \18748 , \18741 , \18746 , \18747 );
and \U$18406 ( \18749 , \18708 , \18748 );
xor \U$18407 ( \18750 , \18587 , \18591 );
xor \U$18408 ( \18751 , \18750 , \18596 );
xor \U$18409 ( \18752 , \18603 , \18607 );
xor \U$18410 ( \18753 , \18752 , \18612 );
and \U$18411 ( \18754 , \18751 , \18753 );
xor \U$18412 ( \18755 , \18557 , \18561 );
xor \U$18413 ( \18756 , \18755 , \18566 );
and \U$18414 ( \18757 , \18753 , \18756 );
and \U$18415 ( \18758 , \18751 , \18756 );
or \U$18416 ( \18759 , \18754 , \18757 , \18758 );
and \U$18417 ( \18760 , \18748 , \18759 );
and \U$18418 ( \18761 , \18708 , \18759 );
or \U$18419 ( \18762 , \18749 , \18760 , \18761 );
xor \U$18420 ( \18763 , \18421 , \18425 );
xor \U$18421 ( \18764 , \18763 , \2566 );
xor \U$18422 ( \18765 , \18434 , \18438 );
xor \U$18423 ( \18766 , \18765 , \18443 );
and \U$18424 ( \18767 , \18764 , \18766 );
xor \U$18425 ( \18768 , \18574 , \18576 );
xor \U$18426 ( \18769 , \18768 , \18579 );
and \U$18427 ( \18770 , \18766 , \18769 );
and \U$18428 ( \18771 , \18764 , \18769 );
or \U$18429 ( \18772 , \18767 , \18770 , \18771 );
and \U$18430 ( \18773 , \18762 , \18772 );
xor \U$18431 ( \18774 , \18536 , \18552 );
xor \U$18432 ( \18775 , \18774 , \18569 );
xor \U$18433 ( \18776 , \18599 , \18615 );
xor \U$18434 ( \18777 , \18776 , \18618 );
and \U$18435 ( \18778 , \18775 , \18777 );
and \U$18436 ( \18779 , \18772 , \18778 );
and \U$18437 ( \18780 , \18762 , \18778 );
or \U$18438 ( \18781 , \18773 , \18779 , \18780 );
xor \U$18439 ( \18782 , \18417 , \18429 );
xor \U$18440 ( \18783 , \18782 , \18446 );
xor \U$18441 ( \18784 , \18572 , \18582 );
xor \U$18442 ( \18785 , \18784 , \18621 );
and \U$18443 ( \18786 , \18783 , \18785 );
xor \U$18444 ( \18787 , \18626 , \18628 );
xor \U$18445 ( \18788 , \18787 , \18631 );
and \U$18446 ( \18789 , \18785 , \18788 );
and \U$18447 ( \18790 , \18783 , \18788 );
or \U$18448 ( \18791 , \18786 , \18789 , \18790 );
and \U$18449 ( \18792 , \18781 , \18791 );
xor \U$18450 ( \18793 , \18472 , \18474 );
xor \U$18451 ( \18794 , \18793 , \18477 );
and \U$18452 ( \18795 , \18791 , \18794 );
and \U$18453 ( \18796 , \18781 , \18794 );
or \U$18454 ( \18797 , \18792 , \18795 , \18796 );
xor \U$18455 ( \18798 , \18401 , \18449 );
xor \U$18456 ( \18799 , \18798 , \18459 );
xor \U$18457 ( \18800 , \18624 , \18634 );
xor \U$18458 ( \18801 , \18800 , \18637 );
and \U$18459 ( \18802 , \18799 , \18801 );
and \U$18460 ( \18803 , \18797 , \18802 );
xor \U$18461 ( \18804 , \18640 , \18642 );
xor \U$18462 ( \18805 , \18804 , \18645 );
and \U$18463 ( \18806 , \18802 , \18805 );
and \U$18464 ( \18807 , \18797 , \18805 );
or \U$18465 ( \18808 , \18803 , \18806 , \18807 );
and \U$18466 ( \18809 , \18660 , \18808 );
xor \U$18467 ( \18810 , \18660 , \18808 );
xor \U$18468 ( \18811 , \18797 , \18802 );
xor \U$18469 ( \18812 , \18811 , \18805 );
and \U$18470 ( \18813 , \5954 , \7035 );
and \U$18471 ( \18814 , \5945 , \7033 );
nor \U$18472 ( \18815 , \18813 , \18814 );
xnor \U$18473 ( \18816 , \18815 , \6775 );
and \U$18474 ( \18817 , \6499 , \6541 );
and \U$18475 ( \18818 , \6297 , \6539 );
nor \U$18476 ( \18819 , \18817 , \18818 );
xnor \U$18477 ( \18820 , \18819 , \6226 );
and \U$18478 ( \18821 , \18816 , \18820 );
and \U$18479 ( \18822 , \6974 , \6032 );
and \U$18480 ( \18823 , \6802 , \6030 );
nor \U$18481 ( \18824 , \18822 , \18823 );
xnor \U$18482 ( \18825 , \18824 , \5692 );
and \U$18483 ( \18826 , \18820 , \18825 );
and \U$18484 ( \18827 , \18816 , \18825 );
or \U$18485 ( \18828 , \18821 , \18826 , \18827 );
and \U$18486 ( \18829 , \4576 , \8693 );
and \U$18487 ( \18830 , \4568 , \8691 );
nor \U$18488 ( \18831 , \18829 , \18830 );
xnor \U$18489 ( \18832 , \18831 , \8322 );
and \U$18490 ( \18833 , \5050 , \8131 );
and \U$18491 ( \18834 , \5045 , \8129 );
nor \U$18492 ( \18835 , \18833 , \18834 );
xnor \U$18493 ( \18836 , \18835 , \7813 );
and \U$18494 ( \18837 , \18832 , \18836 );
and \U$18495 ( \18838 , \5573 , \7564 );
and \U$18496 ( \18839 , \5314 , \7562 );
nor \U$18497 ( \18840 , \18838 , \18839 );
xnor \U$18498 ( \18841 , \18840 , \7315 );
and \U$18499 ( \18842 , \18836 , \18841 );
and \U$18500 ( \18843 , \18832 , \18841 );
or \U$18501 ( \18844 , \18837 , \18842 , \18843 );
and \U$18502 ( \18845 , \18828 , \18844 );
and \U$18503 ( \18846 , \3686 , \10611 );
and \U$18504 ( \18847 , \3478 , \10608 );
nor \U$18505 ( \18848 , \18846 , \18847 );
xnor \U$18506 ( \18849 , \18848 , \9556 );
and \U$18507 ( \18850 , \3813 , \9798 );
and \U$18508 ( \18851 , \3808 , \9796 );
nor \U$18509 ( \18852 , \18850 , \18851 );
xnor \U$18510 ( \18853 , \18852 , \9559 );
and \U$18511 ( \18854 , \18849 , \18853 );
and \U$18512 ( \18855 , \4266 , \9230 );
and \U$18513 ( \18856 , \4069 , \9228 );
nor \U$18514 ( \18857 , \18855 , \18856 );
xnor \U$18515 ( \18858 , \18857 , \8920 );
and \U$18516 ( \18859 , \18853 , \18858 );
and \U$18517 ( \18860 , \18849 , \18858 );
or \U$18518 ( \18861 , \18854 , \18859 , \18860 );
and \U$18519 ( \18862 , \18844 , \18861 );
and \U$18520 ( \18863 , \18828 , \18861 );
or \U$18521 ( \18864 , \18845 , \18862 , \18863 );
and \U$18522 ( \18865 , \9355 , \4152 );
and \U$18523 ( \18866 , \9347 , \4150 );
nor \U$18524 ( \18867 , \18865 , \18866 );
xnor \U$18525 ( \18868 , \18867 , \4009 );
and \U$18526 ( \18869 , \9963 , \3829 );
and \U$18527 ( \18870 , \9958 , \3827 );
nor \U$18528 ( \18871 , \18869 , \18870 );
xnor \U$18529 ( \18872 , \18871 , \3583 );
and \U$18530 ( \18873 , \18868 , \18872 );
and \U$18531 ( \18874 , \10764 , \3434 );
and \U$18532 ( \18875 , \10144 , \3432 );
nor \U$18533 ( \18876 , \18874 , \18875 );
xnor \U$18534 ( \18877 , \18876 , \3247 );
and \U$18535 ( \18878 , \18872 , \18877 );
and \U$18536 ( \18879 , \18868 , \18877 );
or \U$18537 ( \18880 , \18873 , \18878 , \18879 );
and \U$18538 ( \18881 , \7924 , \5443 );
and \U$18539 ( \18882 , \7500 , \5441 );
nor \U$18540 ( \18883 , \18881 , \18882 );
xnor \U$18541 ( \18884 , \18883 , \5202 );
and \U$18542 ( \18885 , \8175 , \4977 );
and \U$18543 ( \18886 , \8170 , \4975 );
nor \U$18544 ( \18887 , \18885 , \18886 );
xnor \U$18545 ( \18888 , \18887 , \4789 );
and \U$18546 ( \18889 , \18884 , \18888 );
and \U$18547 ( \18890 , \8778 , \4603 );
and \U$18548 ( \18891 , \8494 , \4601 );
nor \U$18549 ( \18892 , \18890 , \18891 );
xnor \U$18550 ( \18893 , \18892 , \4371 );
and \U$18551 ( \18894 , \18888 , \18893 );
and \U$18552 ( \18895 , \18884 , \18893 );
or \U$18553 ( \18896 , \18889 , \18894 , \18895 );
and \U$18554 ( \18897 , \18880 , \18896 );
and \U$18555 ( \18898 , \10144 , \3434 );
and \U$18556 ( \18899 , \9963 , \3432 );
nor \U$18557 ( \18900 , \18898 , \18899 );
xnor \U$18558 ( \18901 , \18900 , \3247 );
and \U$18559 ( \18902 , \18896 , \18901 );
and \U$18560 ( \18903 , \18880 , \18901 );
or \U$18561 ( \18904 , \18897 , \18902 , \18903 );
and \U$18562 ( \18905 , \18864 , \18904 );
nand \U$18563 ( \18906 , \10764 , \3119 );
xnor \U$18564 ( \18907 , \18906 , \2916 );
xor \U$18565 ( \18908 , \18712 , \18716 );
xor \U$18566 ( \18909 , \18908 , \18721 );
and \U$18567 ( \18910 , \18907 , \18909 );
xor \U$18568 ( \18911 , \18728 , \18732 );
xor \U$18569 ( \18912 , \18911 , \18737 );
and \U$18570 ( \18913 , \18909 , \18912 );
and \U$18571 ( \18914 , \18907 , \18912 );
or \U$18572 ( \18915 , \18910 , \18913 , \18914 );
and \U$18573 ( \18916 , \18904 , \18915 );
and \U$18574 ( \18917 , \18864 , \18915 );
or \U$18575 ( \18918 , \18905 , \18916 , \18917 );
xor \U$18576 ( \18919 , \18664 , \18668 );
xor \U$18577 ( \18920 , \18919 , \18673 );
xor \U$18578 ( \18921 , \18680 , \18684 );
xor \U$18579 ( \18922 , \18921 , \18689 );
and \U$18580 ( \18923 , \18920 , \18922 );
xor \U$18581 ( \18924 , \18697 , \18701 );
xor \U$18582 ( \18925 , \18924 , \2916 );
and \U$18583 ( \18926 , \18922 , \18925 );
and \U$18584 ( \18927 , \18920 , \18925 );
or \U$18585 ( \18928 , \18923 , \18926 , \18927 );
xor \U$18586 ( \18929 , \18524 , \18528 );
xor \U$18587 ( \18930 , \18929 , \18533 );
and \U$18588 ( \18931 , \18928 , \18930 );
xor \U$18589 ( \18932 , \18540 , \18544 );
xor \U$18590 ( \18933 , \18932 , \18549 );
and \U$18591 ( \18934 , \18930 , \18933 );
and \U$18592 ( \18935 , \18928 , \18933 );
or \U$18593 ( \18936 , \18931 , \18934 , \18935 );
and \U$18594 ( \18937 , \18918 , \18936 );
xor \U$18595 ( \18938 , \18676 , \18692 );
xor \U$18596 ( \18939 , \18938 , \18705 );
xor \U$18597 ( \18940 , \18724 , \18740 );
xor \U$18598 ( \18941 , \18940 , \18745 );
and \U$18599 ( \18942 , \18939 , \18941 );
xor \U$18600 ( \18943 , \18751 , \18753 );
xor \U$18601 ( \18944 , \18943 , \18756 );
and \U$18602 ( \18945 , \18941 , \18944 );
and \U$18603 ( \18946 , \18939 , \18944 );
or \U$18604 ( \18947 , \18942 , \18945 , \18946 );
and \U$18605 ( \18948 , \18936 , \18947 );
and \U$18606 ( \18949 , \18918 , \18947 );
or \U$18607 ( \18950 , \18937 , \18948 , \18949 );
xor \U$18608 ( \18951 , \18708 , \18748 );
xor \U$18609 ( \18952 , \18951 , \18759 );
xor \U$18610 ( \18953 , \18764 , \18766 );
xor \U$18611 ( \18954 , \18953 , \18769 );
and \U$18612 ( \18955 , \18952 , \18954 );
xor \U$18613 ( \18956 , \18775 , \18777 );
and \U$18614 ( \18957 , \18954 , \18956 );
and \U$18615 ( \18958 , \18952 , \18956 );
or \U$18616 ( \18959 , \18955 , \18957 , \18958 );
and \U$18617 ( \18960 , \18950 , \18959 );
xor \U$18618 ( \18961 , \18783 , \18785 );
xor \U$18619 ( \18962 , \18961 , \18788 );
and \U$18620 ( \18963 , \18959 , \18962 );
and \U$18621 ( \18964 , \18950 , \18962 );
or \U$18622 ( \18965 , \18960 , \18963 , \18964 );
xor \U$18623 ( \18966 , \18781 , \18791 );
xor \U$18624 ( \18967 , \18966 , \18794 );
and \U$18625 ( \18968 , \18965 , \18967 );
xor \U$18626 ( \18969 , \18799 , \18801 );
and \U$18627 ( \18970 , \18967 , \18969 );
and \U$18628 ( \18971 , \18965 , \18969 );
or \U$18629 ( \18972 , \18968 , \18970 , \18971 );
and \U$18630 ( \18973 , \18812 , \18972 );
xor \U$18631 ( \18974 , \18812 , \18972 );
xor \U$18632 ( \18975 , \18965 , \18967 );
xor \U$18633 ( \18976 , \18975 , \18969 );
and \U$18634 ( \18977 , \5945 , \7564 );
and \U$18635 ( \18978 , \5573 , \7562 );
nor \U$18636 ( \18979 , \18977 , \18978 );
xnor \U$18637 ( \18980 , \18979 , \7315 );
and \U$18638 ( \18981 , \6297 , \7035 );
and \U$18639 ( \18982 , \5954 , \7033 );
nor \U$18640 ( \18983 , \18981 , \18982 );
xnor \U$18641 ( \18984 , \18983 , \6775 );
and \U$18642 ( \18985 , \18980 , \18984 );
and \U$18643 ( \18986 , \6802 , \6541 );
and \U$18644 ( \18987 , \6499 , \6539 );
nor \U$18645 ( \18988 , \18986 , \18987 );
xnor \U$18646 ( \18989 , \18988 , \6226 );
and \U$18647 ( \18990 , \18984 , \18989 );
and \U$18648 ( \18991 , \18980 , \18989 );
or \U$18649 ( \18992 , \18985 , \18990 , \18991 );
and \U$18650 ( \18993 , \4568 , \9230 );
and \U$18651 ( \18994 , \4266 , \9228 );
nor \U$18652 ( \18995 , \18993 , \18994 );
xnor \U$18653 ( \18996 , \18995 , \8920 );
and \U$18654 ( \18997 , \5045 , \8693 );
and \U$18655 ( \18998 , \4576 , \8691 );
nor \U$18656 ( \18999 , \18997 , \18998 );
xnor \U$18657 ( \19000 , \18999 , \8322 );
and \U$18658 ( \19001 , \18996 , \19000 );
and \U$18659 ( \19002 , \5314 , \8131 );
and \U$18660 ( \19003 , \5050 , \8129 );
nor \U$18661 ( \19004 , \19002 , \19003 );
xnor \U$18662 ( \19005 , \19004 , \7813 );
and \U$18663 ( \19006 , \19000 , \19005 );
and \U$18664 ( \19007 , \18996 , \19005 );
or \U$18665 ( \19008 , \19001 , \19006 , \19007 );
and \U$18666 ( \19009 , \18992 , \19008 );
and \U$18667 ( \19010 , \3808 , \10611 );
and \U$18668 ( \19011 , \3686 , \10608 );
nor \U$18669 ( \19012 , \19010 , \19011 );
xnor \U$18670 ( \19013 , \19012 , \9556 );
and \U$18671 ( \19014 , \4069 , \9798 );
and \U$18672 ( \19015 , \3813 , \9796 );
nor \U$18673 ( \19016 , \19014 , \19015 );
xnor \U$18674 ( \19017 , \19016 , \9559 );
and \U$18675 ( \19018 , \19013 , \19017 );
and \U$18676 ( \19019 , \19017 , \3247 );
and \U$18677 ( \19020 , \19013 , \3247 );
or \U$18678 ( \19021 , \19018 , \19019 , \19020 );
and \U$18679 ( \19022 , \19008 , \19021 );
and \U$18680 ( \19023 , \18992 , \19021 );
or \U$18681 ( \19024 , \19009 , \19022 , \19023 );
and \U$18682 ( \19025 , \7500 , \6032 );
and \U$18683 ( \19026 , \6974 , \6030 );
nor \U$18684 ( \19027 , \19025 , \19026 );
xnor \U$18685 ( \19028 , \19027 , \5692 );
and \U$18686 ( \19029 , \8170 , \5443 );
and \U$18687 ( \19030 , \7924 , \5441 );
nor \U$18688 ( \19031 , \19029 , \19030 );
xnor \U$18689 ( \19032 , \19031 , \5202 );
and \U$18690 ( \19033 , \19028 , \19032 );
and \U$18691 ( \19034 , \8494 , \4977 );
and \U$18692 ( \19035 , \8175 , \4975 );
nor \U$18693 ( \19036 , \19034 , \19035 );
xnor \U$18694 ( \19037 , \19036 , \4789 );
and \U$18695 ( \19038 , \19032 , \19037 );
and \U$18696 ( \19039 , \19028 , \19037 );
or \U$18697 ( \19040 , \19033 , \19038 , \19039 );
and \U$18698 ( \19041 , \9347 , \4603 );
and \U$18699 ( \19042 , \8778 , \4601 );
nor \U$18700 ( \19043 , \19041 , \19042 );
xnor \U$18701 ( \19044 , \19043 , \4371 );
and \U$18702 ( \19045 , \9958 , \4152 );
and \U$18703 ( \19046 , \9355 , \4150 );
nor \U$18704 ( \19047 , \19045 , \19046 );
xnor \U$18705 ( \19048 , \19047 , \4009 );
and \U$18706 ( \19049 , \19044 , \19048 );
and \U$18707 ( \19050 , \10144 , \3829 );
and \U$18708 ( \19051 , \9963 , \3827 );
nor \U$18709 ( \19052 , \19050 , \19051 );
xnor \U$18710 ( \19053 , \19052 , \3583 );
and \U$18711 ( \19054 , \19048 , \19053 );
and \U$18712 ( \19055 , \19044 , \19053 );
or \U$18713 ( \19056 , \19049 , \19054 , \19055 );
and \U$18714 ( \19057 , \19040 , \19056 );
xor \U$18715 ( \19058 , \18868 , \18872 );
xor \U$18716 ( \19059 , \19058 , \18877 );
and \U$18717 ( \19060 , \19056 , \19059 );
and \U$18718 ( \19061 , \19040 , \19059 );
or \U$18719 ( \19062 , \19057 , \19060 , \19061 );
and \U$18720 ( \19063 , \19024 , \19062 );
xor \U$18721 ( \19064 , \18816 , \18820 );
xor \U$18722 ( \19065 , \19064 , \18825 );
xor \U$18723 ( \19066 , \18832 , \18836 );
xor \U$18724 ( \19067 , \19066 , \18841 );
and \U$18725 ( \19068 , \19065 , \19067 );
xor \U$18726 ( \19069 , \18884 , \18888 );
xor \U$18727 ( \19070 , \19069 , \18893 );
and \U$18728 ( \19071 , \19067 , \19070 );
and \U$18729 ( \19072 , \19065 , \19070 );
or \U$18730 ( \19073 , \19068 , \19071 , \19072 );
and \U$18731 ( \19074 , \19062 , \19073 );
and \U$18732 ( \19075 , \19024 , \19073 );
or \U$18733 ( \19076 , \19063 , \19074 , \19075 );
xor \U$18734 ( \19077 , \18880 , \18896 );
xor \U$18735 ( \19078 , \19077 , \18901 );
xor \U$18736 ( \19079 , \18920 , \18922 );
xor \U$18737 ( \19080 , \19079 , \18925 );
and \U$18738 ( \19081 , \19078 , \19080 );
xor \U$18739 ( \19082 , \18907 , \18909 );
xor \U$18740 ( \19083 , \19082 , \18912 );
and \U$18741 ( \19084 , \19080 , \19083 );
and \U$18742 ( \19085 , \19078 , \19083 );
or \U$18743 ( \19086 , \19081 , \19084 , \19085 );
and \U$18744 ( \19087 , \19076 , \19086 );
xor \U$18745 ( \19088 , \18939 , \18941 );
xor \U$18746 ( \19089 , \19088 , \18944 );
and \U$18747 ( \19090 , \19086 , \19089 );
and \U$18748 ( \19091 , \19076 , \19089 );
or \U$18749 ( \19092 , \19087 , \19090 , \19091 );
xor \U$18750 ( \19093 , \18864 , \18904 );
xor \U$18751 ( \19094 , \19093 , \18915 );
xor \U$18752 ( \19095 , \18928 , \18930 );
xor \U$18753 ( \19096 , \19095 , \18933 );
and \U$18754 ( \19097 , \19094 , \19096 );
and \U$18755 ( \19098 , \19092 , \19097 );
xor \U$18756 ( \19099 , \18952 , \18954 );
xor \U$18757 ( \19100 , \19099 , \18956 );
and \U$18758 ( \19101 , \19097 , \19100 );
and \U$18759 ( \19102 , \19092 , \19100 );
or \U$18760 ( \19103 , \19098 , \19101 , \19102 );
xor \U$18761 ( \19104 , \18762 , \18772 );
xor \U$18762 ( \19105 , \19104 , \18778 );
and \U$18763 ( \19106 , \19103 , \19105 );
xor \U$18764 ( \19107 , \18950 , \18959 );
xor \U$18765 ( \19108 , \19107 , \18962 );
and \U$18766 ( \19109 , \19105 , \19108 );
and \U$18767 ( \19110 , \19103 , \19108 );
or \U$18768 ( \19111 , \19106 , \19109 , \19110 );
and \U$18769 ( \19112 , \18976 , \19111 );
xor \U$18770 ( \19113 , \18976 , \19111 );
xor \U$18771 ( \19114 , \19103 , \19105 );
xor \U$18772 ( \19115 , \19114 , \19108 );
and \U$18773 ( \19116 , \3813 , \10611 );
and \U$18774 ( \19117 , \3808 , \10608 );
nor \U$18775 ( \19118 , \19116 , \19117 );
xnor \U$18776 ( \19119 , \19118 , \9556 );
and \U$18777 ( \19120 , \4266 , \9798 );
and \U$18778 ( \19121 , \4069 , \9796 );
nor \U$18779 ( \19122 , \19120 , \19121 );
xnor \U$18780 ( \19123 , \19122 , \9559 );
and \U$18781 ( \19124 , \19119 , \19123 );
and \U$18782 ( \19125 , \4576 , \9230 );
and \U$18783 ( \19126 , \4568 , \9228 );
nor \U$18784 ( \19127 , \19125 , \19126 );
xnor \U$18785 ( \19128 , \19127 , \8920 );
and \U$18786 ( \19129 , \19123 , \19128 );
and \U$18787 ( \19130 , \19119 , \19128 );
or \U$18788 ( \19131 , \19124 , \19129 , \19130 );
and \U$18789 ( \19132 , \6499 , \7035 );
and \U$18790 ( \19133 , \6297 , \7033 );
nor \U$18791 ( \19134 , \19132 , \19133 );
xnor \U$18792 ( \19135 , \19134 , \6775 );
and \U$18793 ( \19136 , \6974 , \6541 );
and \U$18794 ( \19137 , \6802 , \6539 );
nor \U$18795 ( \19138 , \19136 , \19137 );
xnor \U$18796 ( \19139 , \19138 , \6226 );
and \U$18797 ( \19140 , \19135 , \19139 );
and \U$18798 ( \19141 , \7924 , \6032 );
and \U$18799 ( \19142 , \7500 , \6030 );
nor \U$18800 ( \19143 , \19141 , \19142 );
xnor \U$18801 ( \19144 , \19143 , \5692 );
and \U$18802 ( \19145 , \19139 , \19144 );
and \U$18803 ( \19146 , \19135 , \19144 );
or \U$18804 ( \19147 , \19140 , \19145 , \19146 );
and \U$18805 ( \19148 , \19131 , \19147 );
and \U$18806 ( \19149 , \5050 , \8693 );
and \U$18807 ( \19150 , \5045 , \8691 );
nor \U$18808 ( \19151 , \19149 , \19150 );
xnor \U$18809 ( \19152 , \19151 , \8322 );
and \U$18810 ( \19153 , \5573 , \8131 );
and \U$18811 ( \19154 , \5314 , \8129 );
nor \U$18812 ( \19155 , \19153 , \19154 );
xnor \U$18813 ( \19156 , \19155 , \7813 );
and \U$18814 ( \19157 , \19152 , \19156 );
and \U$18815 ( \19158 , \5954 , \7564 );
and \U$18816 ( \19159 , \5945 , \7562 );
nor \U$18817 ( \19160 , \19158 , \19159 );
xnor \U$18818 ( \19161 , \19160 , \7315 );
and \U$18819 ( \19162 , \19156 , \19161 );
and \U$18820 ( \19163 , \19152 , \19161 );
or \U$18821 ( \19164 , \19157 , \19162 , \19163 );
and \U$18822 ( \19165 , \19147 , \19164 );
and \U$18823 ( \19166 , \19131 , \19164 );
or \U$18824 ( \19167 , \19148 , \19165 , \19166 );
xor \U$18825 ( \19168 , \18980 , \18984 );
xor \U$18826 ( \19169 , \19168 , \18989 );
xor \U$18827 ( \19170 , \18996 , \19000 );
xor \U$18828 ( \19171 , \19170 , \19005 );
and \U$18829 ( \19172 , \19169 , \19171 );
xor \U$18830 ( \19173 , \19028 , \19032 );
xor \U$18831 ( \19174 , \19173 , \19037 );
and \U$18832 ( \19175 , \19171 , \19174 );
and \U$18833 ( \19176 , \19169 , \19174 );
or \U$18834 ( \19177 , \19172 , \19175 , \19176 );
and \U$18835 ( \19178 , \19167 , \19177 );
and \U$18836 ( \19179 , \8175 , \5443 );
and \U$18837 ( \19180 , \8170 , \5441 );
nor \U$18838 ( \19181 , \19179 , \19180 );
xnor \U$18839 ( \19182 , \19181 , \5202 );
and \U$18840 ( \19183 , \8778 , \4977 );
and \U$18841 ( \19184 , \8494 , \4975 );
nor \U$18842 ( \19185 , \19183 , \19184 );
xnor \U$18843 ( \19186 , \19185 , \4789 );
and \U$18844 ( \19187 , \19182 , \19186 );
and \U$18845 ( \19188 , \9355 , \4603 );
and \U$18846 ( \19189 , \9347 , \4601 );
nor \U$18847 ( \19190 , \19188 , \19189 );
xnor \U$18848 ( \19191 , \19190 , \4371 );
and \U$18849 ( \19192 , \19186 , \19191 );
and \U$18850 ( \19193 , \19182 , \19191 );
or \U$18851 ( \19194 , \19187 , \19192 , \19193 );
nand \U$18852 ( \19195 , \10764 , \3432 );
xnor \U$18853 ( \19196 , \19195 , \3247 );
and \U$18854 ( \19197 , \19194 , \19196 );
xor \U$18855 ( \19198 , \19044 , \19048 );
xor \U$18856 ( \19199 , \19198 , \19053 );
and \U$18857 ( \19200 , \19196 , \19199 );
and \U$18858 ( \19201 , \19194 , \19199 );
or \U$18859 ( \19202 , \19197 , \19200 , \19201 );
and \U$18860 ( \19203 , \19177 , \19202 );
and \U$18861 ( \19204 , \19167 , \19202 );
or \U$18862 ( \19205 , \19178 , \19203 , \19204 );
xor \U$18863 ( \19206 , \18849 , \18853 );
xor \U$18864 ( \19207 , \19206 , \18858 );
xor \U$18865 ( \19208 , \19040 , \19056 );
xor \U$18866 ( \19209 , \19208 , \19059 );
and \U$18867 ( \19210 , \19207 , \19209 );
xor \U$18868 ( \19211 , \19065 , \19067 );
xor \U$18869 ( \19212 , \19211 , \19070 );
and \U$18870 ( \19213 , \19209 , \19212 );
and \U$18871 ( \19214 , \19207 , \19212 );
or \U$18872 ( \19215 , \19210 , \19213 , \19214 );
and \U$18873 ( \19216 , \19205 , \19215 );
xor \U$18874 ( \19217 , \18828 , \18844 );
xor \U$18875 ( \19218 , \19217 , \18861 );
and \U$18876 ( \19219 , \19215 , \19218 );
and \U$18877 ( \19220 , \19205 , \19218 );
or \U$18878 ( \19221 , \19216 , \19219 , \19220 );
xor \U$18879 ( \19222 , \19076 , \19086 );
xor \U$18880 ( \19223 , \19222 , \19089 );
and \U$18881 ( \19224 , \19221 , \19223 );
xor \U$18882 ( \19225 , \19094 , \19096 );
and \U$18883 ( \19226 , \19223 , \19225 );
and \U$18884 ( \19227 , \19221 , \19225 );
or \U$18885 ( \19228 , \19224 , \19226 , \19227 );
xor \U$18886 ( \19229 , \18918 , \18936 );
xor \U$18887 ( \19230 , \19229 , \18947 );
and \U$18888 ( \19231 , \19228 , \19230 );
xor \U$18889 ( \19232 , \19092 , \19097 );
xor \U$18890 ( \19233 , \19232 , \19100 );
and \U$18891 ( \19234 , \19230 , \19233 );
and \U$18892 ( \19235 , \19228 , \19233 );
or \U$18893 ( \19236 , \19231 , \19234 , \19235 );
and \U$18894 ( \19237 , \19115 , \19236 );
xor \U$18895 ( \19238 , \19115 , \19236 );
xor \U$18896 ( \19239 , \19228 , \19230 );
xor \U$18897 ( \19240 , \19239 , \19233 );
and \U$18898 ( \19241 , \8170 , \6032 );
and \U$18899 ( \19242 , \7924 , \6030 );
nor \U$18900 ( \19243 , \19241 , \19242 );
xnor \U$18901 ( \19244 , \19243 , \5692 );
and \U$18902 ( \19245 , \8494 , \5443 );
and \U$18903 ( \19246 , \8175 , \5441 );
nor \U$18904 ( \19247 , \19245 , \19246 );
xnor \U$18905 ( \19248 , \19247 , \5202 );
and \U$18906 ( \19249 , \19244 , \19248 );
and \U$18907 ( \19250 , \9347 , \4977 );
and \U$18908 ( \19251 , \8778 , \4975 );
nor \U$18909 ( \19252 , \19250 , \19251 );
xnor \U$18910 ( \19253 , \19252 , \4789 );
and \U$18911 ( \19254 , \19248 , \19253 );
and \U$18912 ( \19255 , \19244 , \19253 );
or \U$18913 ( \19256 , \19249 , \19254 , \19255 );
and \U$18914 ( \19257 , \9958 , \4603 );
and \U$18915 ( \19258 , \9355 , \4601 );
nor \U$18916 ( \19259 , \19257 , \19258 );
xnor \U$18917 ( \19260 , \19259 , \4371 );
and \U$18918 ( \19261 , \10144 , \4152 );
and \U$18919 ( \19262 , \9963 , \4150 );
nor \U$18920 ( \19263 , \19261 , \19262 );
xnor \U$18921 ( \19264 , \19263 , \4009 );
and \U$18922 ( \19265 , \19260 , \19264 );
nand \U$18923 ( \19266 , \10764 , \3827 );
xnor \U$18924 ( \19267 , \19266 , \3583 );
and \U$18925 ( \19268 , \19264 , \19267 );
and \U$18926 ( \19269 , \19260 , \19267 );
or \U$18927 ( \19270 , \19265 , \19268 , \19269 );
and \U$18928 ( \19271 , \19256 , \19270 );
and \U$18929 ( \19272 , \9963 , \4152 );
and \U$18930 ( \19273 , \9958 , \4150 );
nor \U$18931 ( \19274 , \19272 , \19273 );
xnor \U$18932 ( \19275 , \19274 , \4009 );
and \U$18933 ( \19276 , \19270 , \19275 );
and \U$18934 ( \19277 , \19256 , \19275 );
or \U$18935 ( \19278 , \19271 , \19276 , \19277 );
and \U$18936 ( \19279 , \6297 , \7564 );
and \U$18937 ( \19280 , \5954 , \7562 );
nor \U$18938 ( \19281 , \19279 , \19280 );
xnor \U$18939 ( \19282 , \19281 , \7315 );
and \U$18940 ( \19283 , \6802 , \7035 );
and \U$18941 ( \19284 , \6499 , \7033 );
nor \U$18942 ( \19285 , \19283 , \19284 );
xnor \U$18943 ( \19286 , \19285 , \6775 );
and \U$18944 ( \19287 , \19282 , \19286 );
and \U$18945 ( \19288 , \7500 , \6541 );
and \U$18946 ( \19289 , \6974 , \6539 );
nor \U$18947 ( \19290 , \19288 , \19289 );
xnor \U$18948 ( \19291 , \19290 , \6226 );
and \U$18949 ( \19292 , \19286 , \19291 );
and \U$18950 ( \19293 , \19282 , \19291 );
or \U$18951 ( \19294 , \19287 , \19292 , \19293 );
and \U$18952 ( \19295 , \4069 , \10611 );
and \U$18953 ( \19296 , \3813 , \10608 );
nor \U$18954 ( \19297 , \19295 , \19296 );
xnor \U$18955 ( \19298 , \19297 , \9556 );
and \U$18956 ( \19299 , \4568 , \9798 );
and \U$18957 ( \19300 , \4266 , \9796 );
nor \U$18958 ( \19301 , \19299 , \19300 );
xnor \U$18959 ( \19302 , \19301 , \9559 );
and \U$18960 ( \19303 , \19298 , \19302 );
and \U$18961 ( \19304 , \19302 , \3583 );
and \U$18962 ( \19305 , \19298 , \3583 );
or \U$18963 ( \19306 , \19303 , \19304 , \19305 );
and \U$18964 ( \19307 , \19294 , \19306 );
and \U$18965 ( \19308 , \5045 , \9230 );
and \U$18966 ( \19309 , \4576 , \9228 );
nor \U$18967 ( \19310 , \19308 , \19309 );
xnor \U$18968 ( \19311 , \19310 , \8920 );
and \U$18969 ( \19312 , \5314 , \8693 );
and \U$18970 ( \19313 , \5050 , \8691 );
nor \U$18971 ( \19314 , \19312 , \19313 );
xnor \U$18972 ( \19315 , \19314 , \8322 );
and \U$18973 ( \19316 , \19311 , \19315 );
and \U$18974 ( \19317 , \5945 , \8131 );
and \U$18975 ( \19318 , \5573 , \8129 );
nor \U$18976 ( \19319 , \19317 , \19318 );
xnor \U$18977 ( \19320 , \19319 , \7813 );
and \U$18978 ( \19321 , \19315 , \19320 );
and \U$18979 ( \19322 , \19311 , \19320 );
or \U$18980 ( \19323 , \19316 , \19321 , \19322 );
and \U$18981 ( \19324 , \19306 , \19323 );
and \U$18982 ( \19325 , \19294 , \19323 );
or \U$18983 ( \19326 , \19307 , \19324 , \19325 );
and \U$18984 ( \19327 , \19278 , \19326 );
and \U$18985 ( \19328 , \10764 , \3829 );
and \U$18986 ( \19329 , \10144 , \3827 );
nor \U$18987 ( \19330 , \19328 , \19329 );
xnor \U$18988 ( \19331 , \19330 , \3583 );
xor \U$18989 ( \19332 , \19182 , \19186 );
xor \U$18990 ( \19333 , \19332 , \19191 );
and \U$18991 ( \19334 , \19331 , \19333 );
xor \U$18992 ( \19335 , \19135 , \19139 );
xor \U$18993 ( \19336 , \19335 , \19144 );
and \U$18994 ( \19337 , \19333 , \19336 );
and \U$18995 ( \19338 , \19331 , \19336 );
or \U$18996 ( \19339 , \19334 , \19337 , \19338 );
and \U$18997 ( \19340 , \19326 , \19339 );
and \U$18998 ( \19341 , \19278 , \19339 );
or \U$18999 ( \19342 , \19327 , \19340 , \19341 );
xor \U$19000 ( \19343 , \19013 , \19017 );
xor \U$19001 ( \19344 , \19343 , \3247 );
xor \U$19002 ( \19345 , \19169 , \19171 );
xor \U$19003 ( \19346 , \19345 , \19174 );
and \U$19004 ( \19347 , \19344 , \19346 );
xor \U$19005 ( \19348 , \19194 , \19196 );
xor \U$19006 ( \19349 , \19348 , \19199 );
and \U$19007 ( \19350 , \19346 , \19349 );
and \U$19008 ( \19351 , \19344 , \19349 );
or \U$19009 ( \19352 , \19347 , \19350 , \19351 );
and \U$19010 ( \19353 , \19342 , \19352 );
xor \U$19011 ( \19354 , \18992 , \19008 );
xor \U$19012 ( \19355 , \19354 , \19021 );
and \U$19013 ( \19356 , \19352 , \19355 );
and \U$19014 ( \19357 , \19342 , \19355 );
or \U$19015 ( \19358 , \19353 , \19356 , \19357 );
xor \U$19016 ( \19359 , \19167 , \19177 );
xor \U$19017 ( \19360 , \19359 , \19202 );
xor \U$19018 ( \19361 , \19207 , \19209 );
xor \U$19019 ( \19362 , \19361 , \19212 );
and \U$19020 ( \19363 , \19360 , \19362 );
and \U$19021 ( \19364 , \19358 , \19363 );
xor \U$19022 ( \19365 , \19078 , \19080 );
xor \U$19023 ( \19366 , \19365 , \19083 );
and \U$19024 ( \19367 , \19363 , \19366 );
and \U$19025 ( \19368 , \19358 , \19366 );
or \U$19026 ( \19369 , \19364 , \19367 , \19368 );
xor \U$19027 ( \19370 , \19024 , \19062 );
xor \U$19028 ( \19371 , \19370 , \19073 );
xor \U$19029 ( \19372 , \19205 , \19215 );
xor \U$19030 ( \19373 , \19372 , \19218 );
and \U$19031 ( \19374 , \19371 , \19373 );
and \U$19032 ( \19375 , \19369 , \19374 );
xor \U$19033 ( \19376 , \19221 , \19223 );
xor \U$19034 ( \19377 , \19376 , \19225 );
and \U$19035 ( \19378 , \19374 , \19377 );
and \U$19036 ( \19379 , \19369 , \19377 );
or \U$19037 ( \19380 , \19375 , \19378 , \19379 );
and \U$19038 ( \19381 , \19240 , \19380 );
xor \U$19039 ( \19382 , \19240 , \19380 );
xor \U$19040 ( \19383 , \19369 , \19374 );
xor \U$19041 ( \19384 , \19383 , \19377 );
and \U$19042 ( \19385 , \5573 , \8693 );
and \U$19043 ( \19386 , \5314 , \8691 );
nor \U$19044 ( \19387 , \19385 , \19386 );
xnor \U$19045 ( \19388 , \19387 , \8322 );
and \U$19046 ( \19389 , \5954 , \8131 );
and \U$19047 ( \19390 , \5945 , \8129 );
nor \U$19048 ( \19391 , \19389 , \19390 );
xnor \U$19049 ( \19392 , \19391 , \7813 );
and \U$19050 ( \19393 , \19388 , \19392 );
and \U$19051 ( \19394 , \6499 , \7564 );
and \U$19052 ( \19395 , \6297 , \7562 );
nor \U$19053 ( \19396 , \19394 , \19395 );
xnor \U$19054 ( \19397 , \19396 , \7315 );
and \U$19055 ( \19398 , \19392 , \19397 );
and \U$19056 ( \19399 , \19388 , \19397 );
or \U$19057 ( \19400 , \19393 , \19398 , \19399 );
and \U$19058 ( \19401 , \4266 , \10611 );
and \U$19059 ( \19402 , \4069 , \10608 );
nor \U$19060 ( \19403 , \19401 , \19402 );
xnor \U$19061 ( \19404 , \19403 , \9556 );
and \U$19062 ( \19405 , \4576 , \9798 );
and \U$19063 ( \19406 , \4568 , \9796 );
nor \U$19064 ( \19407 , \19405 , \19406 );
xnor \U$19065 ( \19408 , \19407 , \9559 );
and \U$19066 ( \19409 , \19404 , \19408 );
and \U$19067 ( \19410 , \5050 , \9230 );
and \U$19068 ( \19411 , \5045 , \9228 );
nor \U$19069 ( \19412 , \19410 , \19411 );
xnor \U$19070 ( \19413 , \19412 , \8920 );
and \U$19071 ( \19414 , \19408 , \19413 );
and \U$19072 ( \19415 , \19404 , \19413 );
or \U$19073 ( \19416 , \19409 , \19414 , \19415 );
and \U$19074 ( \19417 , \19400 , \19416 );
and \U$19075 ( \19418 , \6974 , \7035 );
and \U$19076 ( \19419 , \6802 , \7033 );
nor \U$19077 ( \19420 , \19418 , \19419 );
xnor \U$19078 ( \19421 , \19420 , \6775 );
and \U$19079 ( \19422 , \7924 , \6541 );
and \U$19080 ( \19423 , \7500 , \6539 );
nor \U$19081 ( \19424 , \19422 , \19423 );
xnor \U$19082 ( \19425 , \19424 , \6226 );
and \U$19083 ( \19426 , \19421 , \19425 );
and \U$19084 ( \19427 , \8175 , \6032 );
and \U$19085 ( \19428 , \8170 , \6030 );
nor \U$19086 ( \19429 , \19427 , \19428 );
xnor \U$19087 ( \19430 , \19429 , \5692 );
and \U$19088 ( \19431 , \19425 , \19430 );
and \U$19089 ( \19432 , \19421 , \19430 );
or \U$19090 ( \19433 , \19426 , \19431 , \19432 );
and \U$19091 ( \19434 , \19416 , \19433 );
and \U$19092 ( \19435 , \19400 , \19433 );
or \U$19093 ( \19436 , \19417 , \19434 , \19435 );
xor \U$19094 ( \19437 , \19282 , \19286 );
xor \U$19095 ( \19438 , \19437 , \19291 );
xor \U$19096 ( \19439 , \19298 , \19302 );
xor \U$19097 ( \19440 , \19439 , \3583 );
and \U$19098 ( \19441 , \19438 , \19440 );
xor \U$19099 ( \19442 , \19311 , \19315 );
xor \U$19100 ( \19443 , \19442 , \19320 );
and \U$19101 ( \19444 , \19440 , \19443 );
and \U$19102 ( \19445 , \19438 , \19443 );
or \U$19103 ( \19446 , \19441 , \19444 , \19445 );
and \U$19104 ( \19447 , \19436 , \19446 );
and \U$19105 ( \19448 , \8778 , \5443 );
and \U$19106 ( \19449 , \8494 , \5441 );
nor \U$19107 ( \19450 , \19448 , \19449 );
xnor \U$19108 ( \19451 , \19450 , \5202 );
and \U$19109 ( \19452 , \9355 , \4977 );
and \U$19110 ( \19453 , \9347 , \4975 );
nor \U$19111 ( \19454 , \19452 , \19453 );
xnor \U$19112 ( \19455 , \19454 , \4789 );
and \U$19113 ( \19456 , \19451 , \19455 );
and \U$19114 ( \19457 , \9963 , \4603 );
and \U$19115 ( \19458 , \9958 , \4601 );
nor \U$19116 ( \19459 , \19457 , \19458 );
xnor \U$19117 ( \19460 , \19459 , \4371 );
and \U$19118 ( \19461 , \19455 , \19460 );
and \U$19119 ( \19462 , \19451 , \19460 );
or \U$19120 ( \19463 , \19456 , \19461 , \19462 );
xor \U$19121 ( \19464 , \19244 , \19248 );
xor \U$19122 ( \19465 , \19464 , \19253 );
and \U$19123 ( \19466 , \19463 , \19465 );
xor \U$19124 ( \19467 , \19260 , \19264 );
xor \U$19125 ( \19468 , \19467 , \19267 );
and \U$19126 ( \19469 , \19465 , \19468 );
and \U$19127 ( \19470 , \19463 , \19468 );
or \U$19128 ( \19471 , \19466 , \19469 , \19470 );
and \U$19129 ( \19472 , \19446 , \19471 );
and \U$19130 ( \19473 , \19436 , \19471 );
or \U$19131 ( \19474 , \19447 , \19472 , \19473 );
xor \U$19132 ( \19475 , \19119 , \19123 );
xor \U$19133 ( \19476 , \19475 , \19128 );
xor \U$19134 ( \19477 , \19152 , \19156 );
xor \U$19135 ( \19478 , \19477 , \19161 );
and \U$19136 ( \19479 , \19476 , \19478 );
xor \U$19137 ( \19480 , \19331 , \19333 );
xor \U$19138 ( \19481 , \19480 , \19336 );
and \U$19139 ( \19482 , \19478 , \19481 );
and \U$19140 ( \19483 , \19476 , \19481 );
or \U$19141 ( \19484 , \19479 , \19482 , \19483 );
and \U$19142 ( \19485 , \19474 , \19484 );
xor \U$19143 ( \19486 , \19131 , \19147 );
xor \U$19144 ( \19487 , \19486 , \19164 );
and \U$19145 ( \19488 , \19484 , \19487 );
and \U$19146 ( \19489 , \19474 , \19487 );
or \U$19147 ( \19490 , \19485 , \19488 , \19489 );
xor \U$19148 ( \19491 , \19342 , \19352 );
xor \U$19149 ( \19492 , \19491 , \19355 );
and \U$19150 ( \19493 , \19490 , \19492 );
xor \U$19151 ( \19494 , \19360 , \19362 );
and \U$19152 ( \19495 , \19492 , \19494 );
and \U$19153 ( \19496 , \19490 , \19494 );
or \U$19154 ( \19497 , \19493 , \19495 , \19496 );
xor \U$19155 ( \19498 , \19358 , \19363 );
xor \U$19156 ( \19499 , \19498 , \19366 );
and \U$19157 ( \19500 , \19497 , \19499 );
xor \U$19158 ( \19501 , \19371 , \19373 );
and \U$19159 ( \19502 , \19499 , \19501 );
and \U$19160 ( \19503 , \19497 , \19501 );
or \U$19161 ( \19504 , \19500 , \19502 , \19503 );
and \U$19162 ( \19505 , \19384 , \19504 );
xor \U$19163 ( \19506 , \19384 , \19504 );
xor \U$19164 ( \19507 , \19497 , \19499 );
xor \U$19165 ( \19508 , \19507 , \19501 );
and \U$19166 ( \19509 , \5314 , \9230 );
and \U$19167 ( \19510 , \5050 , \9228 );
nor \U$19168 ( \19511 , \19509 , \19510 );
xnor \U$19169 ( \19512 , \19511 , \8920 );
and \U$19170 ( \19513 , \5945 , \8693 );
and \U$19171 ( \19514 , \5573 , \8691 );
nor \U$19172 ( \19515 , \19513 , \19514 );
xnor \U$19173 ( \19516 , \19515 , \8322 );
and \U$19174 ( \19517 , \19512 , \19516 );
and \U$19175 ( \19518 , \6297 , \8131 );
and \U$19176 ( \19519 , \5954 , \8129 );
nor \U$19177 ( \19520 , \19518 , \19519 );
xnor \U$19178 ( \19521 , \19520 , \7813 );
and \U$19179 ( \19522 , \19516 , \19521 );
and \U$19180 ( \19523 , \19512 , \19521 );
or \U$19181 ( \19524 , \19517 , \19522 , \19523 );
and \U$19182 ( \19525 , \4568 , \10611 );
and \U$19183 ( \19526 , \4266 , \10608 );
nor \U$19184 ( \19527 , \19525 , \19526 );
xnor \U$19185 ( \19528 , \19527 , \9556 );
and \U$19186 ( \19529 , \5045 , \9798 );
and \U$19187 ( \19530 , \4576 , \9796 );
nor \U$19188 ( \19531 , \19529 , \19530 );
xnor \U$19189 ( \19532 , \19531 , \9559 );
and \U$19190 ( \19533 , \19528 , \19532 );
and \U$19191 ( \19534 , \19532 , \4009 );
and \U$19192 ( \19535 , \19528 , \4009 );
or \U$19193 ( \19536 , \19533 , \19534 , \19535 );
and \U$19194 ( \19537 , \19524 , \19536 );
and \U$19195 ( \19538 , \6802 , \7564 );
and \U$19196 ( \19539 , \6499 , \7562 );
nor \U$19197 ( \19540 , \19538 , \19539 );
xnor \U$19198 ( \19541 , \19540 , \7315 );
and \U$19199 ( \19542 , \7500 , \7035 );
and \U$19200 ( \19543 , \6974 , \7033 );
nor \U$19201 ( \19544 , \19542 , \19543 );
xnor \U$19202 ( \19545 , \19544 , \6775 );
and \U$19203 ( \19546 , \19541 , \19545 );
and \U$19204 ( \19547 , \8170 , \6541 );
and \U$19205 ( \19548 , \7924 , \6539 );
nor \U$19206 ( \19549 , \19547 , \19548 );
xnor \U$19207 ( \19550 , \19549 , \6226 );
and \U$19208 ( \19551 , \19545 , \19550 );
and \U$19209 ( \19552 , \19541 , \19550 );
or \U$19210 ( \19553 , \19546 , \19551 , \19552 );
and \U$19211 ( \19554 , \19536 , \19553 );
and \U$19212 ( \19555 , \19524 , \19553 );
or \U$19213 ( \19556 , \19537 , \19554 , \19555 );
and \U$19214 ( \19557 , \8494 , \6032 );
and \U$19215 ( \19558 , \8175 , \6030 );
nor \U$19216 ( \19559 , \19557 , \19558 );
xnor \U$19217 ( \19560 , \19559 , \5692 );
and \U$19218 ( \19561 , \9347 , \5443 );
and \U$19219 ( \19562 , \8778 , \5441 );
nor \U$19220 ( \19563 , \19561 , \19562 );
xnor \U$19221 ( \19564 , \19563 , \5202 );
and \U$19222 ( \19565 , \19560 , \19564 );
and \U$19223 ( \19566 , \9958 , \4977 );
and \U$19224 ( \19567 , \9355 , \4975 );
nor \U$19225 ( \19568 , \19566 , \19567 );
xnor \U$19226 ( \19569 , \19568 , \4789 );
and \U$19227 ( \19570 , \19564 , \19569 );
and \U$19228 ( \19571 , \19560 , \19569 );
or \U$19229 ( \19572 , \19565 , \19570 , \19571 );
and \U$19230 ( \19573 , \10144 , \4603 );
and \U$19231 ( \19574 , \9963 , \4601 );
nor \U$19232 ( \19575 , \19573 , \19574 );
xnor \U$19233 ( \19576 , \19575 , \4371 );
nand \U$19234 ( \19577 , \10764 , \4150 );
xnor \U$19235 ( \19578 , \19577 , \4009 );
and \U$19236 ( \19579 , \19576 , \19578 );
and \U$19237 ( \19580 , \19572 , \19579 );
and \U$19238 ( \19581 , \10764 , \4152 );
and \U$19239 ( \19582 , \10144 , \4150 );
nor \U$19240 ( \19583 , \19581 , \19582 );
xnor \U$19241 ( \19584 , \19583 , \4009 );
and \U$19242 ( \19585 , \19579 , \19584 );
and \U$19243 ( \19586 , \19572 , \19584 );
or \U$19244 ( \19587 , \19580 , \19585 , \19586 );
and \U$19245 ( \19588 , \19556 , \19587 );
xor \U$19246 ( \19589 , \19388 , \19392 );
xor \U$19247 ( \19590 , \19589 , \19397 );
xor \U$19248 ( \19591 , \19451 , \19455 );
xor \U$19249 ( \19592 , \19591 , \19460 );
and \U$19250 ( \19593 , \19590 , \19592 );
xor \U$19251 ( \19594 , \19421 , \19425 );
xor \U$19252 ( \19595 , \19594 , \19430 );
and \U$19253 ( \19596 , \19592 , \19595 );
and \U$19254 ( \19597 , \19590 , \19595 );
or \U$19255 ( \19598 , \19593 , \19596 , \19597 );
and \U$19256 ( \19599 , \19587 , \19598 );
and \U$19257 ( \19600 , \19556 , \19598 );
or \U$19258 ( \19601 , \19588 , \19599 , \19600 );
xor \U$19259 ( \19602 , \19400 , \19416 );
xor \U$19260 ( \19603 , \19602 , \19433 );
xor \U$19261 ( \19604 , \19438 , \19440 );
xor \U$19262 ( \19605 , \19604 , \19443 );
and \U$19263 ( \19606 , \19603 , \19605 );
xor \U$19264 ( \19607 , \19463 , \19465 );
xor \U$19265 ( \19608 , \19607 , \19468 );
and \U$19266 ( \19609 , \19605 , \19608 );
and \U$19267 ( \19610 , \19603 , \19608 );
or \U$19268 ( \19611 , \19606 , \19609 , \19610 );
and \U$19269 ( \19612 , \19601 , \19611 );
xor \U$19270 ( \19613 , \19256 , \19270 );
xor \U$19271 ( \19614 , \19613 , \19275 );
and \U$19272 ( \19615 , \19611 , \19614 );
and \U$19273 ( \19616 , \19601 , \19614 );
or \U$19274 ( \19617 , \19612 , \19615 , \19616 );
xor \U$19275 ( \19618 , \19294 , \19306 );
xor \U$19276 ( \19619 , \19618 , \19323 );
xor \U$19277 ( \19620 , \19436 , \19446 );
xor \U$19278 ( \19621 , \19620 , \19471 );
and \U$19279 ( \19622 , \19619 , \19621 );
xor \U$19280 ( \19623 , \19476 , \19478 );
xor \U$19281 ( \19624 , \19623 , \19481 );
and \U$19282 ( \19625 , \19621 , \19624 );
and \U$19283 ( \19626 , \19619 , \19624 );
or \U$19284 ( \19627 , \19622 , \19625 , \19626 );
and \U$19285 ( \19628 , \19617 , \19627 );
xor \U$19286 ( \19629 , \19344 , \19346 );
xor \U$19287 ( \19630 , \19629 , \19349 );
and \U$19288 ( \19631 , \19627 , \19630 );
and \U$19289 ( \19632 , \19617 , \19630 );
or \U$19290 ( \19633 , \19628 , \19631 , \19632 );
xor \U$19291 ( \19634 , \19278 , \19326 );
xor \U$19292 ( \19635 , \19634 , \19339 );
xor \U$19293 ( \19636 , \19474 , \19484 );
xor \U$19294 ( \19637 , \19636 , \19487 );
and \U$19295 ( \19638 , \19635 , \19637 );
and \U$19296 ( \19639 , \19633 , \19638 );
xor \U$19297 ( \19640 , \19490 , \19492 );
xor \U$19298 ( \19641 , \19640 , \19494 );
and \U$19299 ( \19642 , \19638 , \19641 );
and \U$19300 ( \19643 , \19633 , \19641 );
or \U$19301 ( \19644 , \19639 , \19642 , \19643 );
and \U$19302 ( \19645 , \19508 , \19644 );
xor \U$19303 ( \19646 , \19508 , \19644 );
xor \U$19304 ( \19647 , \19633 , \19638 );
xor \U$19305 ( \19648 , \19647 , \19641 );
and \U$19306 ( \19649 , \5954 , \8693 );
and \U$19307 ( \19650 , \5945 , \8691 );
nor \U$19308 ( \19651 , \19649 , \19650 );
xnor \U$19309 ( \19652 , \19651 , \8322 );
and \U$19310 ( \19653 , \6499 , \8131 );
and \U$19311 ( \19654 , \6297 , \8129 );
nor \U$19312 ( \19655 , \19653 , \19654 );
xnor \U$19313 ( \19656 , \19655 , \7813 );
and \U$19314 ( \19657 , \19652 , \19656 );
and \U$19315 ( \19658 , \6974 , \7564 );
and \U$19316 ( \19659 , \6802 , \7562 );
nor \U$19317 ( \19660 , \19658 , \19659 );
xnor \U$19318 ( \19661 , \19660 , \7315 );
and \U$19319 ( \19662 , \19656 , \19661 );
and \U$19320 ( \19663 , \19652 , \19661 );
or \U$19321 ( \19664 , \19657 , \19662 , \19663 );
and \U$19322 ( \19665 , \7924 , \7035 );
and \U$19323 ( \19666 , \7500 , \7033 );
nor \U$19324 ( \19667 , \19665 , \19666 );
xnor \U$19325 ( \19668 , \19667 , \6775 );
and \U$19326 ( \19669 , \8175 , \6541 );
and \U$19327 ( \19670 , \8170 , \6539 );
nor \U$19328 ( \19671 , \19669 , \19670 );
xnor \U$19329 ( \19672 , \19671 , \6226 );
and \U$19330 ( \19673 , \19668 , \19672 );
and \U$19331 ( \19674 , \8778 , \6032 );
and \U$19332 ( \19675 , \8494 , \6030 );
nor \U$19333 ( \19676 , \19674 , \19675 );
xnor \U$19334 ( \19677 , \19676 , \5692 );
and \U$19335 ( \19678 , \19672 , \19677 );
and \U$19336 ( \19679 , \19668 , \19677 );
or \U$19337 ( \19680 , \19673 , \19678 , \19679 );
and \U$19338 ( \19681 , \19664 , \19680 );
and \U$19339 ( \19682 , \4576 , \10611 );
and \U$19340 ( \19683 , \4568 , \10608 );
nor \U$19341 ( \19684 , \19682 , \19683 );
xnor \U$19342 ( \19685 , \19684 , \9556 );
and \U$19343 ( \19686 , \5050 , \9798 );
and \U$19344 ( \19687 , \5045 , \9796 );
nor \U$19345 ( \19688 , \19686 , \19687 );
xnor \U$19346 ( \19689 , \19688 , \9559 );
and \U$19347 ( \19690 , \19685 , \19689 );
and \U$19348 ( \19691 , \5573 , \9230 );
and \U$19349 ( \19692 , \5314 , \9228 );
nor \U$19350 ( \19693 , \19691 , \19692 );
xnor \U$19351 ( \19694 , \19693 , \8920 );
and \U$19352 ( \19695 , \19689 , \19694 );
and \U$19353 ( \19696 , \19685 , \19694 );
or \U$19354 ( \19697 , \19690 , \19695 , \19696 );
and \U$19355 ( \19698 , \19680 , \19697 );
and \U$19356 ( \19699 , \19664 , \19697 );
or \U$19357 ( \19700 , \19681 , \19698 , \19699 );
xor \U$19358 ( \19701 , \19512 , \19516 );
xor \U$19359 ( \19702 , \19701 , \19521 );
xor \U$19360 ( \19703 , \19528 , \19532 );
xor \U$19361 ( \19704 , \19703 , \4009 );
and \U$19362 ( \19705 , \19702 , \19704 );
xor \U$19363 ( \19706 , \19541 , \19545 );
xor \U$19364 ( \19707 , \19706 , \19550 );
and \U$19365 ( \19708 , \19704 , \19707 );
and \U$19366 ( \19709 , \19702 , \19707 );
or \U$19367 ( \19710 , \19705 , \19708 , \19709 );
and \U$19368 ( \19711 , \19700 , \19710 );
and \U$19369 ( \19712 , \9355 , \5443 );
and \U$19370 ( \19713 , \9347 , \5441 );
nor \U$19371 ( \19714 , \19712 , \19713 );
xnor \U$19372 ( \19715 , \19714 , \5202 );
and \U$19373 ( \19716 , \9963 , \4977 );
and \U$19374 ( \19717 , \9958 , \4975 );
nor \U$19375 ( \19718 , \19716 , \19717 );
xnor \U$19376 ( \19719 , \19718 , \4789 );
and \U$19377 ( \19720 , \19715 , \19719 );
and \U$19378 ( \19721 , \10764 , \4603 );
and \U$19379 ( \19722 , \10144 , \4601 );
nor \U$19380 ( \19723 , \19721 , \19722 );
xnor \U$19381 ( \19724 , \19723 , \4371 );
and \U$19382 ( \19725 , \19719 , \19724 );
and \U$19383 ( \19726 , \19715 , \19724 );
or \U$19384 ( \19727 , \19720 , \19725 , \19726 );
xor \U$19385 ( \19728 , \19560 , \19564 );
xor \U$19386 ( \19729 , \19728 , \19569 );
and \U$19387 ( \19730 , \19727 , \19729 );
xor \U$19388 ( \19731 , \19576 , \19578 );
and \U$19389 ( \19732 , \19729 , \19731 );
and \U$19390 ( \19733 , \19727 , \19731 );
or \U$19391 ( \19734 , \19730 , \19732 , \19733 );
and \U$19392 ( \19735 , \19710 , \19734 );
and \U$19393 ( \19736 , \19700 , \19734 );
or \U$19394 ( \19737 , \19711 , \19735 , \19736 );
xor \U$19395 ( \19738 , \19404 , \19408 );
xor \U$19396 ( \19739 , \19738 , \19413 );
xor \U$19397 ( \19740 , \19572 , \19579 );
xor \U$19398 ( \19741 , \19740 , \19584 );
and \U$19399 ( \19742 , \19739 , \19741 );
xor \U$19400 ( \19743 , \19590 , \19592 );
xor \U$19401 ( \19744 , \19743 , \19595 );
and \U$19402 ( \19745 , \19741 , \19744 );
and \U$19403 ( \19746 , \19739 , \19744 );
or \U$19404 ( \19747 , \19742 , \19745 , \19746 );
and \U$19405 ( \19748 , \19737 , \19747 );
xor \U$19406 ( \19749 , \19603 , \19605 );
xor \U$19407 ( \19750 , \19749 , \19608 );
and \U$19408 ( \19751 , \19747 , \19750 );
and \U$19409 ( \19752 , \19737 , \19750 );
or \U$19410 ( \19753 , \19748 , \19751 , \19752 );
xor \U$19411 ( \19754 , \19601 , \19611 );
xor \U$19412 ( \19755 , \19754 , \19614 );
and \U$19413 ( \19756 , \19753 , \19755 );
xor \U$19414 ( \19757 , \19619 , \19621 );
xor \U$19415 ( \19758 , \19757 , \19624 );
and \U$19416 ( \19759 , \19755 , \19758 );
and \U$19417 ( \19760 , \19753 , \19758 );
or \U$19418 ( \19761 , \19756 , \19759 , \19760 );
xor \U$19419 ( \19762 , \19617 , \19627 );
xor \U$19420 ( \19763 , \19762 , \19630 );
and \U$19421 ( \19764 , \19761 , \19763 );
xor \U$19422 ( \19765 , \19635 , \19637 );
and \U$19423 ( \19766 , \19763 , \19765 );
and \U$19424 ( \19767 , \19761 , \19765 );
or \U$19425 ( \19768 , \19764 , \19766 , \19767 );
and \U$19426 ( \19769 , \19648 , \19768 );
xor \U$19427 ( \19770 , \19648 , \19768 );
xor \U$19428 ( \19771 , \19761 , \19763 );
xor \U$19429 ( \19772 , \19771 , \19765 );
and \U$19430 ( \19773 , \5945 , \9230 );
and \U$19431 ( \19774 , \5573 , \9228 );
nor \U$19432 ( \19775 , \19773 , \19774 );
xnor \U$19433 ( \19776 , \19775 , \8920 );
and \U$19434 ( \19777 , \6297 , \8693 );
and \U$19435 ( \19778 , \5954 , \8691 );
nor \U$19436 ( \19779 , \19777 , \19778 );
xnor \U$19437 ( \19780 , \19779 , \8322 );
and \U$19438 ( \19781 , \19776 , \19780 );
and \U$19439 ( \19782 , \6802 , \8131 );
and \U$19440 ( \19783 , \6499 , \8129 );
nor \U$19441 ( \19784 , \19782 , \19783 );
xnor \U$19442 ( \19785 , \19784 , \7813 );
and \U$19443 ( \19786 , \19780 , \19785 );
and \U$19444 ( \19787 , \19776 , \19785 );
or \U$19445 ( \19788 , \19781 , \19786 , \19787 );
and \U$19446 ( \19789 , \7500 , \7564 );
and \U$19447 ( \19790 , \6974 , \7562 );
nor \U$19448 ( \19791 , \19789 , \19790 );
xnor \U$19449 ( \19792 , \19791 , \7315 );
and \U$19450 ( \19793 , \8170 , \7035 );
and \U$19451 ( \19794 , \7924 , \7033 );
nor \U$19452 ( \19795 , \19793 , \19794 );
xnor \U$19453 ( \19796 , \19795 , \6775 );
and \U$19454 ( \19797 , \19792 , \19796 );
and \U$19455 ( \19798 , \8494 , \6541 );
and \U$19456 ( \19799 , \8175 , \6539 );
nor \U$19457 ( \19800 , \19798 , \19799 );
xnor \U$19458 ( \19801 , \19800 , \6226 );
and \U$19459 ( \19802 , \19796 , \19801 );
and \U$19460 ( \19803 , \19792 , \19801 );
or \U$19461 ( \19804 , \19797 , \19802 , \19803 );
and \U$19462 ( \19805 , \19788 , \19804 );
and \U$19463 ( \19806 , \5045 , \10611 );
and \U$19464 ( \19807 , \4576 , \10608 );
nor \U$19465 ( \19808 , \19806 , \19807 );
xnor \U$19466 ( \19809 , \19808 , \9556 );
and \U$19467 ( \19810 , \5314 , \9798 );
and \U$19468 ( \19811 , \5050 , \9796 );
nor \U$19469 ( \19812 , \19810 , \19811 );
xnor \U$19470 ( \19813 , \19812 , \9559 );
and \U$19471 ( \19814 , \19809 , \19813 );
and \U$19472 ( \19815 , \19813 , \4371 );
and \U$19473 ( \19816 , \19809 , \4371 );
or \U$19474 ( \19817 , \19814 , \19815 , \19816 );
and \U$19475 ( \19818 , \19804 , \19817 );
and \U$19476 ( \19819 , \19788 , \19817 );
or \U$19477 ( \19820 , \19805 , \19818 , \19819 );
and \U$19478 ( \19821 , \9347 , \6032 );
and \U$19479 ( \19822 , \8778 , \6030 );
nor \U$19480 ( \19823 , \19821 , \19822 );
xnor \U$19481 ( \19824 , \19823 , \5692 );
and \U$19482 ( \19825 , \9958 , \5443 );
and \U$19483 ( \19826 , \9355 , \5441 );
nor \U$19484 ( \19827 , \19825 , \19826 );
xnor \U$19485 ( \19828 , \19827 , \5202 );
and \U$19486 ( \19829 , \19824 , \19828 );
and \U$19487 ( \19830 , \10144 , \4977 );
and \U$19488 ( \19831 , \9963 , \4975 );
nor \U$19489 ( \19832 , \19830 , \19831 );
xnor \U$19490 ( \19833 , \19832 , \4789 );
and \U$19491 ( \19834 , \19828 , \19833 );
and \U$19492 ( \19835 , \19824 , \19833 );
or \U$19493 ( \19836 , \19829 , \19834 , \19835 );
xor \U$19494 ( \19837 , \19668 , \19672 );
xor \U$19495 ( \19838 , \19837 , \19677 );
and \U$19496 ( \19839 , \19836 , \19838 );
xor \U$19497 ( \19840 , \19715 , \19719 );
xor \U$19498 ( \19841 , \19840 , \19724 );
and \U$19499 ( \19842 , \19838 , \19841 );
and \U$19500 ( \19843 , \19836 , \19841 );
or \U$19501 ( \19844 , \19839 , \19842 , \19843 );
and \U$19502 ( \19845 , \19820 , \19844 );
xor \U$19503 ( \19846 , \19652 , \19656 );
xor \U$19504 ( \19847 , \19846 , \19661 );
xor \U$19505 ( \19848 , \19685 , \19689 );
xor \U$19506 ( \19849 , \19848 , \19694 );
and \U$19507 ( \19850 , \19847 , \19849 );
and \U$19508 ( \19851 , \19844 , \19850 );
and \U$19509 ( \19852 , \19820 , \19850 );
or \U$19510 ( \19853 , \19845 , \19851 , \19852 );
xor \U$19511 ( \19854 , \19664 , \19680 );
xor \U$19512 ( \19855 , \19854 , \19697 );
xor \U$19513 ( \19856 , \19702 , \19704 );
xor \U$19514 ( \19857 , \19856 , \19707 );
and \U$19515 ( \19858 , \19855 , \19857 );
xor \U$19516 ( \19859 , \19727 , \19729 );
xor \U$19517 ( \19860 , \19859 , \19731 );
and \U$19518 ( \19861 , \19857 , \19860 );
and \U$19519 ( \19862 , \19855 , \19860 );
or \U$19520 ( \19863 , \19858 , \19861 , \19862 );
and \U$19521 ( \19864 , \19853 , \19863 );
xor \U$19522 ( \19865 , \19524 , \19536 );
xor \U$19523 ( \19866 , \19865 , \19553 );
and \U$19524 ( \19867 , \19863 , \19866 );
and \U$19525 ( \19868 , \19853 , \19866 );
or \U$19526 ( \19869 , \19864 , \19867 , \19868 );
xor \U$19527 ( \19870 , \19700 , \19710 );
xor \U$19528 ( \19871 , \19870 , \19734 );
xor \U$19529 ( \19872 , \19739 , \19741 );
xor \U$19530 ( \19873 , \19872 , \19744 );
and \U$19531 ( \19874 , \19871 , \19873 );
and \U$19532 ( \19875 , \19869 , \19874 );
xor \U$19533 ( \19876 , \19556 , \19587 );
xor \U$19534 ( \19877 , \19876 , \19598 );
and \U$19535 ( \19878 , \19874 , \19877 );
and \U$19536 ( \19879 , \19869 , \19877 );
or \U$19537 ( \19880 , \19875 , \19878 , \19879 );
xor \U$19538 ( \19881 , \19753 , \19755 );
xor \U$19539 ( \19882 , \19881 , \19758 );
and \U$19540 ( \19883 , \19880 , \19882 );
and \U$19541 ( \19884 , \19772 , \19883 );
xor \U$19542 ( \19885 , \19772 , \19883 );
xor \U$19543 ( \19886 , \19880 , \19882 );
xor \U$19544 ( \19887 , \19869 , \19874 );
xor \U$19545 ( \19888 , \19887 , \19877 );
xor \U$19546 ( \19889 , \19737 , \19747 );
xor \U$19547 ( \19890 , \19889 , \19750 );
and \U$19548 ( \19891 , \19888 , \19890 );
and \U$19549 ( \19892 , \19886 , \19891 );
xor \U$19550 ( \19893 , \19886 , \19891 );
xor \U$19551 ( \19894 , \19888 , \19890 );
and \U$19552 ( \19895 , \5050 , \10611 );
and \U$19553 ( \19896 , \5045 , \10608 );
nor \U$19554 ( \19897 , \19895 , \19896 );
xnor \U$19555 ( \19898 , \19897 , \9556 );
and \U$19556 ( \19899 , \5573 , \9798 );
and \U$19557 ( \19900 , \5314 , \9796 );
nor \U$19558 ( \19901 , \19899 , \19900 );
xnor \U$19559 ( \19902 , \19901 , \9559 );
and \U$19560 ( \19903 , \19898 , \19902 );
and \U$19561 ( \19904 , \5954 , \9230 );
and \U$19562 ( \19905 , \5945 , \9228 );
nor \U$19563 ( \19906 , \19904 , \19905 );
xnor \U$19564 ( \19907 , \19906 , \8920 );
and \U$19565 ( \19908 , \19902 , \19907 );
and \U$19566 ( \19909 , \19898 , \19907 );
or \U$19567 ( \19910 , \19903 , \19908 , \19909 );
and \U$19568 ( \19911 , \8175 , \7035 );
and \U$19569 ( \19912 , \8170 , \7033 );
nor \U$19570 ( \19913 , \19911 , \19912 );
xnor \U$19571 ( \19914 , \19913 , \6775 );
and \U$19572 ( \19915 , \8778 , \6541 );
and \U$19573 ( \19916 , \8494 , \6539 );
nor \U$19574 ( \19917 , \19915 , \19916 );
xnor \U$19575 ( \19918 , \19917 , \6226 );
and \U$19576 ( \19919 , \19914 , \19918 );
and \U$19577 ( \19920 , \9355 , \6032 );
and \U$19578 ( \19921 , \9347 , \6030 );
nor \U$19579 ( \19922 , \19920 , \19921 );
xnor \U$19580 ( \19923 , \19922 , \5692 );
and \U$19581 ( \19924 , \19918 , \19923 );
and \U$19582 ( \19925 , \19914 , \19923 );
or \U$19583 ( \19926 , \19919 , \19924 , \19925 );
and \U$19584 ( \19927 , \19910 , \19926 );
and \U$19585 ( \19928 , \6499 , \8693 );
and \U$19586 ( \19929 , \6297 , \8691 );
nor \U$19587 ( \19930 , \19928 , \19929 );
xnor \U$19588 ( \19931 , \19930 , \8322 );
and \U$19589 ( \19932 , \6974 , \8131 );
and \U$19590 ( \19933 , \6802 , \8129 );
nor \U$19591 ( \19934 , \19932 , \19933 );
xnor \U$19592 ( \19935 , \19934 , \7813 );
and \U$19593 ( \19936 , \19931 , \19935 );
and \U$19594 ( \19937 , \7924 , \7564 );
and \U$19595 ( \19938 , \7500 , \7562 );
nor \U$19596 ( \19939 , \19937 , \19938 );
xnor \U$19597 ( \19940 , \19939 , \7315 );
and \U$19598 ( \19941 , \19935 , \19940 );
and \U$19599 ( \19942 , \19931 , \19940 );
or \U$19600 ( \19943 , \19936 , \19941 , \19942 );
and \U$19601 ( \19944 , \19926 , \19943 );
and \U$19602 ( \19945 , \19910 , \19943 );
or \U$19603 ( \19946 , \19927 , \19944 , \19945 );
nand \U$19604 ( \19947 , \10764 , \4601 );
xnor \U$19605 ( \19948 , \19947 , \4371 );
xor \U$19606 ( \19949 , \19792 , \19796 );
xor \U$19607 ( \19950 , \19949 , \19801 );
and \U$19608 ( \19951 , \19948 , \19950 );
xor \U$19609 ( \19952 , \19824 , \19828 );
xor \U$19610 ( \19953 , \19952 , \19833 );
and \U$19611 ( \19954 , \19950 , \19953 );
and \U$19612 ( \19955 , \19948 , \19953 );
or \U$19613 ( \19956 , \19951 , \19954 , \19955 );
and \U$19614 ( \19957 , \19946 , \19956 );
xor \U$19615 ( \19958 , \19776 , \19780 );
xor \U$19616 ( \19959 , \19958 , \19785 );
xor \U$19617 ( \19960 , \19809 , \19813 );
xor \U$19618 ( \19961 , \19960 , \4371 );
and \U$19619 ( \19962 , \19959 , \19961 );
and \U$19620 ( \19963 , \19956 , \19962 );
and \U$19621 ( \19964 , \19946 , \19962 );
or \U$19622 ( \19965 , \19957 , \19963 , \19964 );
xor \U$19623 ( \19966 , \19788 , \19804 );
xor \U$19624 ( \19967 , \19966 , \19817 );
xor \U$19625 ( \19968 , \19836 , \19838 );
xor \U$19626 ( \19969 , \19968 , \19841 );
and \U$19627 ( \19970 , \19967 , \19969 );
xor \U$19628 ( \19971 , \19847 , \19849 );
and \U$19629 ( \19972 , \19969 , \19971 );
and \U$19630 ( \19973 , \19967 , \19971 );
or \U$19631 ( \19974 , \19970 , \19972 , \19973 );
and \U$19632 ( \19975 , \19965 , \19974 );
xor \U$19633 ( \19976 , \19855 , \19857 );
xor \U$19634 ( \19977 , \19976 , \19860 );
and \U$19635 ( \19978 , \19974 , \19977 );
and \U$19636 ( \19979 , \19965 , \19977 );
or \U$19637 ( \19980 , \19975 , \19978 , \19979 );
xor \U$19638 ( \19981 , \19853 , \19863 );
xor \U$19639 ( \19982 , \19981 , \19866 );
and \U$19640 ( \19983 , \19980 , \19982 );
xor \U$19641 ( \19984 , \19871 , \19873 );
and \U$19642 ( \19985 , \19982 , \19984 );
and \U$19643 ( \19986 , \19980 , \19984 );
or \U$19644 ( \19987 , \19983 , \19985 , \19986 );
and \U$19645 ( \19988 , \19894 , \19987 );
xor \U$19646 ( \19989 , \19894 , \19987 );
xor \U$19647 ( \19990 , \19980 , \19982 );
xor \U$19648 ( \19991 , \19990 , \19984 );
and \U$19649 ( \19992 , \9958 , \6032 );
and \U$19650 ( \19993 , \9355 , \6030 );
nor \U$19651 ( \19994 , \19992 , \19993 );
xnor \U$19652 ( \19995 , \19994 , \5692 );
and \U$19653 ( \19996 , \10144 , \5443 );
and \U$19654 ( \19997 , \9963 , \5441 );
nor \U$19655 ( \19998 , \19996 , \19997 );
xnor \U$19656 ( \19999 , \19998 , \5202 );
and \U$19657 ( \20000 , \19995 , \19999 );
nand \U$19658 ( \20001 , \10764 , \4975 );
xnor \U$19659 ( \20002 , \20001 , \4789 );
and \U$19660 ( \20003 , \19999 , \20002 );
and \U$19661 ( \20004 , \19995 , \20002 );
or \U$19662 ( \20005 , \20000 , \20003 , \20004 );
and \U$19663 ( \20006 , \9963 , \5443 );
and \U$19664 ( \20007 , \9958 , \5441 );
nor \U$19665 ( \20008 , \20006 , \20007 );
xnor \U$19666 ( \20009 , \20008 , \5202 );
and \U$19667 ( \20010 , \20005 , \20009 );
and \U$19668 ( \20011 , \10764 , \4977 );
and \U$19669 ( \20012 , \10144 , \4975 );
nor \U$19670 ( \20013 , \20011 , \20012 );
xnor \U$19671 ( \20014 , \20013 , \4789 );
and \U$19672 ( \20015 , \20009 , \20014 );
and \U$19673 ( \20016 , \20005 , \20014 );
or \U$19674 ( \20017 , \20010 , \20015 , \20016 );
and \U$19675 ( \20018 , \5314 , \10611 );
and \U$19676 ( \20019 , \5050 , \10608 );
nor \U$19677 ( \20020 , \20018 , \20019 );
xnor \U$19678 ( \20021 , \20020 , \9556 );
and \U$19679 ( \20022 , \5945 , \9798 );
and \U$19680 ( \20023 , \5573 , \9796 );
nor \U$19681 ( \20024 , \20022 , \20023 );
xnor \U$19682 ( \20025 , \20024 , \9559 );
and \U$19683 ( \20026 , \20021 , \20025 );
and \U$19684 ( \20027 , \20025 , \4789 );
and \U$19685 ( \20028 , \20021 , \4789 );
or \U$19686 ( \20029 , \20026 , \20027 , \20028 );
and \U$19687 ( \20030 , \6297 , \9230 );
and \U$19688 ( \20031 , \5954 , \9228 );
nor \U$19689 ( \20032 , \20030 , \20031 );
xnor \U$19690 ( \20033 , \20032 , \8920 );
and \U$19691 ( \20034 , \6802 , \8693 );
and \U$19692 ( \20035 , \6499 , \8691 );
nor \U$19693 ( \20036 , \20034 , \20035 );
xnor \U$19694 ( \20037 , \20036 , \8322 );
and \U$19695 ( \20038 , \20033 , \20037 );
and \U$19696 ( \20039 , \7500 , \8131 );
and \U$19697 ( \20040 , \6974 , \8129 );
nor \U$19698 ( \20041 , \20039 , \20040 );
xnor \U$19699 ( \20042 , \20041 , \7813 );
and \U$19700 ( \20043 , \20037 , \20042 );
and \U$19701 ( \20044 , \20033 , \20042 );
or \U$19702 ( \20045 , \20038 , \20043 , \20044 );
and \U$19703 ( \20046 , \20029 , \20045 );
and \U$19704 ( \20047 , \8170 , \7564 );
and \U$19705 ( \20048 , \7924 , \7562 );
nor \U$19706 ( \20049 , \20047 , \20048 );
xnor \U$19707 ( \20050 , \20049 , \7315 );
and \U$19708 ( \20051 , \8494 , \7035 );
and \U$19709 ( \20052 , \8175 , \7033 );
nor \U$19710 ( \20053 , \20051 , \20052 );
xnor \U$19711 ( \20054 , \20053 , \6775 );
and \U$19712 ( \20055 , \20050 , \20054 );
and \U$19713 ( \20056 , \9347 , \6541 );
and \U$19714 ( \20057 , \8778 , \6539 );
nor \U$19715 ( \20058 , \20056 , \20057 );
xnor \U$19716 ( \20059 , \20058 , \6226 );
and \U$19717 ( \20060 , \20054 , \20059 );
and \U$19718 ( \20061 , \20050 , \20059 );
or \U$19719 ( \20062 , \20055 , \20060 , \20061 );
and \U$19720 ( \20063 , \20045 , \20062 );
and \U$19721 ( \20064 , \20029 , \20062 );
or \U$19722 ( \20065 , \20046 , \20063 , \20064 );
and \U$19723 ( \20066 , \20017 , \20065 );
xor \U$19724 ( \20067 , \19898 , \19902 );
xor \U$19725 ( \20068 , \20067 , \19907 );
xor \U$19726 ( \20069 , \19914 , \19918 );
xor \U$19727 ( \20070 , \20069 , \19923 );
and \U$19728 ( \20071 , \20068 , \20070 );
xor \U$19729 ( \20072 , \19931 , \19935 );
xor \U$19730 ( \20073 , \20072 , \19940 );
and \U$19731 ( \20074 , \20070 , \20073 );
and \U$19732 ( \20075 , \20068 , \20073 );
or \U$19733 ( \20076 , \20071 , \20074 , \20075 );
and \U$19734 ( \20077 , \20065 , \20076 );
and \U$19735 ( \20078 , \20017 , \20076 );
or \U$19736 ( \20079 , \20066 , \20077 , \20078 );
xor \U$19737 ( \20080 , \19910 , \19926 );
xor \U$19738 ( \20081 , \20080 , \19943 );
xor \U$19739 ( \20082 , \19948 , \19950 );
xor \U$19740 ( \20083 , \20082 , \19953 );
and \U$19741 ( \20084 , \20081 , \20083 );
xor \U$19742 ( \20085 , \19959 , \19961 );
and \U$19743 ( \20086 , \20083 , \20085 );
and \U$19744 ( \20087 , \20081 , \20085 );
or \U$19745 ( \20088 , \20084 , \20086 , \20087 );
and \U$19746 ( \20089 , \20079 , \20088 );
xor \U$19747 ( \20090 , \19967 , \19969 );
xor \U$19748 ( \20091 , \20090 , \19971 );
and \U$19749 ( \20092 , \20088 , \20091 );
and \U$19750 ( \20093 , \20079 , \20091 );
or \U$19751 ( \20094 , \20089 , \20092 , \20093 );
xor \U$19752 ( \20095 , \19820 , \19844 );
xor \U$19753 ( \20096 , \20095 , \19850 );
and \U$19754 ( \20097 , \20094 , \20096 );
xor \U$19755 ( \20098 , \19965 , \19974 );
xor \U$19756 ( \20099 , \20098 , \19977 );
and \U$19757 ( \20100 , \20096 , \20099 );
and \U$19758 ( \20101 , \20094 , \20099 );
or \U$19759 ( \20102 , \20097 , \20100 , \20101 );
and \U$19760 ( \20103 , \19991 , \20102 );
xor \U$19761 ( \20104 , \19991 , \20102 );
xor \U$19762 ( \20105 , \20094 , \20096 );
xor \U$19763 ( \20106 , \20105 , \20099 );
and \U$19764 ( \20107 , \8778 , \7035 );
and \U$19765 ( \20108 , \8494 , \7033 );
nor \U$19766 ( \20109 , \20107 , \20108 );
xnor \U$19767 ( \20110 , \20109 , \6775 );
and \U$19768 ( \20111 , \9355 , \6541 );
and \U$19769 ( \20112 , \9347 , \6539 );
nor \U$19770 ( \20113 , \20111 , \20112 );
xnor \U$19771 ( \20114 , \20113 , \6226 );
and \U$19772 ( \20115 , \20110 , \20114 );
and \U$19773 ( \20116 , \9963 , \6032 );
and \U$19774 ( \20117 , \9958 , \6030 );
nor \U$19775 ( \20118 , \20116 , \20117 );
xnor \U$19776 ( \20119 , \20118 , \5692 );
and \U$19777 ( \20120 , \20114 , \20119 );
and \U$19778 ( \20121 , \20110 , \20119 );
or \U$19779 ( \20122 , \20115 , \20120 , \20121 );
and \U$19780 ( \20123 , \5573 , \10611 );
and \U$19781 ( \20124 , \5314 , \10608 );
nor \U$19782 ( \20125 , \20123 , \20124 );
xnor \U$19783 ( \20126 , \20125 , \9556 );
and \U$19784 ( \20127 , \5954 , \9798 );
and \U$19785 ( \20128 , \5945 , \9796 );
nor \U$19786 ( \20129 , \20127 , \20128 );
xnor \U$19787 ( \20130 , \20129 , \9559 );
and \U$19788 ( \20131 , \20126 , \20130 );
and \U$19789 ( \20132 , \6499 , \9230 );
and \U$19790 ( \20133 , \6297 , \9228 );
nor \U$19791 ( \20134 , \20132 , \20133 );
xnor \U$19792 ( \20135 , \20134 , \8920 );
and \U$19793 ( \20136 , \20130 , \20135 );
and \U$19794 ( \20137 , \20126 , \20135 );
or \U$19795 ( \20138 , \20131 , \20136 , \20137 );
and \U$19796 ( \20139 , \20122 , \20138 );
and \U$19797 ( \20140 , \6974 , \8693 );
and \U$19798 ( \20141 , \6802 , \8691 );
nor \U$19799 ( \20142 , \20140 , \20141 );
xnor \U$19800 ( \20143 , \20142 , \8322 );
and \U$19801 ( \20144 , \7924 , \8131 );
and \U$19802 ( \20145 , \7500 , \8129 );
nor \U$19803 ( \20146 , \20144 , \20145 );
xnor \U$19804 ( \20147 , \20146 , \7813 );
and \U$19805 ( \20148 , \20143 , \20147 );
and \U$19806 ( \20149 , \8175 , \7564 );
and \U$19807 ( \20150 , \8170 , \7562 );
nor \U$19808 ( \20151 , \20149 , \20150 );
xnor \U$19809 ( \20152 , \20151 , \7315 );
and \U$19810 ( \20153 , \20147 , \20152 );
and \U$19811 ( \20154 , \20143 , \20152 );
or \U$19812 ( \20155 , \20148 , \20153 , \20154 );
and \U$19813 ( \20156 , \20138 , \20155 );
and \U$19814 ( \20157 , \20122 , \20155 );
or \U$19815 ( \20158 , \20139 , \20156 , \20157 );
xor \U$19816 ( \20159 , \20033 , \20037 );
xor \U$19817 ( \20160 , \20159 , \20042 );
xor \U$19818 ( \20161 , \19995 , \19999 );
xor \U$19819 ( \20162 , \20161 , \20002 );
and \U$19820 ( \20163 , \20160 , \20162 );
xor \U$19821 ( \20164 , \20050 , \20054 );
xor \U$19822 ( \20165 , \20164 , \20059 );
and \U$19823 ( \20166 , \20162 , \20165 );
and \U$19824 ( \20167 , \20160 , \20165 );
or \U$19825 ( \20168 , \20163 , \20166 , \20167 );
and \U$19826 ( \20169 , \20158 , \20168 );
xor \U$19827 ( \20170 , \20068 , \20070 );
xor \U$19828 ( \20171 , \20170 , \20073 );
and \U$19829 ( \20172 , \20168 , \20171 );
and \U$19830 ( \20173 , \20158 , \20171 );
or \U$19831 ( \20174 , \20169 , \20172 , \20173 );
xor \U$19832 ( \20175 , \20017 , \20065 );
xor \U$19833 ( \20176 , \20175 , \20076 );
and \U$19834 ( \20177 , \20174 , \20176 );
xor \U$19835 ( \20178 , \20081 , \20083 );
xor \U$19836 ( \20179 , \20178 , \20085 );
and \U$19837 ( \20180 , \20176 , \20179 );
and \U$19838 ( \20181 , \20174 , \20179 );
or \U$19839 ( \20182 , \20177 , \20180 , \20181 );
xor \U$19840 ( \20183 , \19946 , \19956 );
xor \U$19841 ( \20184 , \20183 , \19962 );
and \U$19842 ( \20185 , \20182 , \20184 );
xor \U$19843 ( \20186 , \20079 , \20088 );
xor \U$19844 ( \20187 , \20186 , \20091 );
and \U$19845 ( \20188 , \20184 , \20187 );
and \U$19846 ( \20189 , \20182 , \20187 );
or \U$19847 ( \20190 , \20185 , \20188 , \20189 );
and \U$19848 ( \20191 , \20106 , \20190 );
xor \U$19849 ( \20192 , \20106 , \20190 );
xor \U$19850 ( \20193 , \20182 , \20184 );
xor \U$19851 ( \20194 , \20193 , \20187 );
and \U$19852 ( \20195 , \5945 , \10611 );
and \U$19853 ( \20196 , \5573 , \10608 );
nor \U$19854 ( \20197 , \20195 , \20196 );
xnor \U$19855 ( \20198 , \20197 , \9556 );
and \U$19856 ( \20199 , \6297 , \9798 );
and \U$19857 ( \20200 , \5954 , \9796 );
nor \U$19858 ( \20201 , \20199 , \20200 );
xnor \U$19859 ( \20202 , \20201 , \9559 );
and \U$19860 ( \20203 , \20198 , \20202 );
and \U$19861 ( \20204 , \20202 , \5202 );
and \U$19862 ( \20205 , \20198 , \5202 );
or \U$19863 ( \20206 , \20203 , \20204 , \20205 );
and \U$19864 ( \20207 , \8494 , \7564 );
and \U$19865 ( \20208 , \8175 , \7562 );
nor \U$19866 ( \20209 , \20207 , \20208 );
xnor \U$19867 ( \20210 , \20209 , \7315 );
and \U$19868 ( \20211 , \9347 , \7035 );
and \U$19869 ( \20212 , \8778 , \7033 );
nor \U$19870 ( \20213 , \20211 , \20212 );
xnor \U$19871 ( \20214 , \20213 , \6775 );
and \U$19872 ( \20215 , \20210 , \20214 );
and \U$19873 ( \20216 , \9958 , \6541 );
and \U$19874 ( \20217 , \9355 , \6539 );
nor \U$19875 ( \20218 , \20216 , \20217 );
xnor \U$19876 ( \20219 , \20218 , \6226 );
and \U$19877 ( \20220 , \20214 , \20219 );
and \U$19878 ( \20221 , \20210 , \20219 );
or \U$19879 ( \20222 , \20215 , \20220 , \20221 );
and \U$19880 ( \20223 , \20206 , \20222 );
and \U$19881 ( \20224 , \6802 , \9230 );
and \U$19882 ( \20225 , \6499 , \9228 );
nor \U$19883 ( \20226 , \20224 , \20225 );
xnor \U$19884 ( \20227 , \20226 , \8920 );
and \U$19885 ( \20228 , \7500 , \8693 );
and \U$19886 ( \20229 , \6974 , \8691 );
nor \U$19887 ( \20230 , \20228 , \20229 );
xnor \U$19888 ( \20231 , \20230 , \8322 );
and \U$19889 ( \20232 , \20227 , \20231 );
and \U$19890 ( \20233 , \8170 , \8131 );
and \U$19891 ( \20234 , \7924 , \8129 );
nor \U$19892 ( \20235 , \20233 , \20234 );
xnor \U$19893 ( \20236 , \20235 , \7813 );
and \U$19894 ( \20237 , \20231 , \20236 );
and \U$19895 ( \20238 , \20227 , \20236 );
or \U$19896 ( \20239 , \20232 , \20237 , \20238 );
and \U$19897 ( \20240 , \20222 , \20239 );
and \U$19898 ( \20241 , \20206 , \20239 );
or \U$19899 ( \20242 , \20223 , \20240 , \20241 );
and \U$19900 ( \20243 , \10764 , \5443 );
and \U$19901 ( \20244 , \10144 , \5441 );
nor \U$19902 ( \20245 , \20243 , \20244 );
xnor \U$19903 ( \20246 , \20245 , \5202 );
xor \U$19904 ( \20247 , \20110 , \20114 );
xor \U$19905 ( \20248 , \20247 , \20119 );
and \U$19906 ( \20249 , \20246 , \20248 );
xor \U$19907 ( \20250 , \20143 , \20147 );
xor \U$19908 ( \20251 , \20250 , \20152 );
and \U$19909 ( \20252 , \20248 , \20251 );
and \U$19910 ( \20253 , \20246 , \20251 );
or \U$19911 ( \20254 , \20249 , \20252 , \20253 );
and \U$19912 ( \20255 , \20242 , \20254 );
xor \U$19913 ( \20256 , \20021 , \20025 );
xor \U$19914 ( \20257 , \20256 , \4789 );
and \U$19915 ( \20258 , \20254 , \20257 );
and \U$19916 ( \20259 , \20242 , \20257 );
or \U$19917 ( \20260 , \20255 , \20258 , \20259 );
xor \U$19918 ( \20261 , \20122 , \20138 );
xor \U$19919 ( \20262 , \20261 , \20155 );
xor \U$19920 ( \20263 , \20160 , \20162 );
xor \U$19921 ( \20264 , \20263 , \20165 );
and \U$19922 ( \20265 , \20262 , \20264 );
and \U$19923 ( \20266 , \20260 , \20265 );
xor \U$19924 ( \20267 , \20005 , \20009 );
xor \U$19925 ( \20268 , \20267 , \20014 );
and \U$19926 ( \20269 , \20265 , \20268 );
and \U$19927 ( \20270 , \20260 , \20268 );
or \U$19928 ( \20271 , \20266 , \20269 , \20270 );
xor \U$19929 ( \20272 , \20029 , \20045 );
xor \U$19930 ( \20273 , \20272 , \20062 );
xor \U$19931 ( \20274 , \20158 , \20168 );
xor \U$19932 ( \20275 , \20274 , \20171 );
and \U$19933 ( \20276 , \20273 , \20275 );
and \U$19934 ( \20277 , \20271 , \20276 );
xor \U$19935 ( \20278 , \20174 , \20176 );
xor \U$19936 ( \20279 , \20278 , \20179 );
and \U$19937 ( \20280 , \20276 , \20279 );
and \U$19938 ( \20281 , \20271 , \20279 );
or \U$19939 ( \20282 , \20277 , \20280 , \20281 );
and \U$19940 ( \20283 , \20194 , \20282 );
xor \U$19941 ( \20284 , \20194 , \20282 );
xor \U$19942 ( \20285 , \20271 , \20276 );
xor \U$19943 ( \20286 , \20285 , \20279 );
and \U$19944 ( \20287 , \7924 , \8693 );
and \U$19945 ( \20288 , \7500 , \8691 );
nor \U$19946 ( \20289 , \20287 , \20288 );
xnor \U$19947 ( \20290 , \20289 , \8322 );
and \U$19948 ( \20291 , \8175 , \8131 );
and \U$19949 ( \20292 , \8170 , \8129 );
nor \U$19950 ( \20293 , \20291 , \20292 );
xnor \U$19951 ( \20294 , \20293 , \7813 );
and \U$19952 ( \20295 , \20290 , \20294 );
and \U$19953 ( \20296 , \8778 , \7564 );
and \U$19954 ( \20297 , \8494 , \7562 );
nor \U$19955 ( \20298 , \20296 , \20297 );
xnor \U$19956 ( \20299 , \20298 , \7315 );
and \U$19957 ( \20300 , \20294 , \20299 );
and \U$19958 ( \20301 , \20290 , \20299 );
or \U$19959 ( \20302 , \20295 , \20300 , \20301 );
and \U$19960 ( \20303 , \5954 , \10611 );
and \U$19961 ( \20304 , \5945 , \10608 );
nor \U$19962 ( \20305 , \20303 , \20304 );
xnor \U$19963 ( \20306 , \20305 , \9556 );
and \U$19964 ( \20307 , \6499 , \9798 );
and \U$19965 ( \20308 , \6297 , \9796 );
nor \U$19966 ( \20309 , \20307 , \20308 );
xnor \U$19967 ( \20310 , \20309 , \9559 );
and \U$19968 ( \20311 , \20306 , \20310 );
and \U$19969 ( \20312 , \6974 , \9230 );
and \U$19970 ( \20313 , \6802 , \9228 );
nor \U$19971 ( \20314 , \20312 , \20313 );
xnor \U$19972 ( \20315 , \20314 , \8920 );
and \U$19973 ( \20316 , \20310 , \20315 );
and \U$19974 ( \20317 , \20306 , \20315 );
or \U$19975 ( \20318 , \20311 , \20316 , \20317 );
and \U$19976 ( \20319 , \20302 , \20318 );
and \U$19977 ( \20320 , \9355 , \7035 );
and \U$19978 ( \20321 , \9347 , \7033 );
nor \U$19979 ( \20322 , \20320 , \20321 );
xnor \U$19980 ( \20323 , \20322 , \6775 );
and \U$19981 ( \20324 , \9963 , \6541 );
and \U$19982 ( \20325 , \9958 , \6539 );
nor \U$19983 ( \20326 , \20324 , \20325 );
xnor \U$19984 ( \20327 , \20326 , \6226 );
and \U$19985 ( \20328 , \20323 , \20327 );
and \U$19986 ( \20329 , \10764 , \6032 );
and \U$19987 ( \20330 , \10144 , \6030 );
nor \U$19988 ( \20331 , \20329 , \20330 );
xnor \U$19989 ( \20332 , \20331 , \5692 );
and \U$19990 ( \20333 , \20327 , \20332 );
and \U$19991 ( \20334 , \20323 , \20332 );
or \U$19992 ( \20335 , \20328 , \20333 , \20334 );
and \U$19993 ( \20336 , \20318 , \20335 );
and \U$19994 ( \20337 , \20302 , \20335 );
or \U$19995 ( \20338 , \20319 , \20336 , \20337 );
and \U$19996 ( \20339 , \10144 , \6032 );
and \U$19997 ( \20340 , \9963 , \6030 );
nor \U$19998 ( \20341 , \20339 , \20340 );
xnor \U$19999 ( \20342 , \20341 , \5692 );
nand \U$20000 ( \20343 , \10764 , \5441 );
xnor \U$20001 ( \20344 , \20343 , \5202 );
and \U$20002 ( \20345 , \20342 , \20344 );
xor \U$20003 ( \20346 , \20210 , \20214 );
xor \U$20004 ( \20347 , \20346 , \20219 );
and \U$20005 ( \20348 , \20344 , \20347 );
and \U$20006 ( \20349 , \20342 , \20347 );
or \U$20007 ( \20350 , \20345 , \20348 , \20349 );
and \U$20008 ( \20351 , \20338 , \20350 );
xor \U$20009 ( \20352 , \20126 , \20130 );
xor \U$20010 ( \20353 , \20352 , \20135 );
and \U$20011 ( \20354 , \20350 , \20353 );
and \U$20012 ( \20355 , \20338 , \20353 );
or \U$20013 ( \20356 , \20351 , \20354 , \20355 );
xor \U$20014 ( \20357 , \20242 , \20254 );
xor \U$20015 ( \20358 , \20357 , \20257 );
and \U$20016 ( \20359 , \20356 , \20358 );
xor \U$20017 ( \20360 , \20262 , \20264 );
and \U$20018 ( \20361 , \20358 , \20360 );
and \U$20019 ( \20362 , \20356 , \20360 );
or \U$20020 ( \20363 , \20359 , \20361 , \20362 );
xor \U$20021 ( \20364 , \20260 , \20265 );
xor \U$20022 ( \20365 , \20364 , \20268 );
and \U$20023 ( \20366 , \20363 , \20365 );
xor \U$20024 ( \20367 , \20273 , \20275 );
and \U$20025 ( \20368 , \20365 , \20367 );
and \U$20026 ( \20369 , \20363 , \20367 );
or \U$20027 ( \20370 , \20366 , \20368 , \20369 );
and \U$20028 ( \20371 , \20286 , \20370 );
xor \U$20029 ( \20372 , \20286 , \20370 );
xor \U$20030 ( \20373 , \20363 , \20365 );
xor \U$20031 ( \20374 , \20373 , \20367 );
and \U$20032 ( \20375 , \7500 , \9230 );
and \U$20033 ( \20376 , \6974 , \9228 );
nor \U$20034 ( \20377 , \20375 , \20376 );
xnor \U$20035 ( \20378 , \20377 , \8920 );
and \U$20036 ( \20379 , \8170 , \8693 );
and \U$20037 ( \20380 , \7924 , \8691 );
nor \U$20038 ( \20381 , \20379 , \20380 );
xnor \U$20039 ( \20382 , \20381 , \8322 );
and \U$20040 ( \20383 , \20378 , \20382 );
and \U$20041 ( \20384 , \8494 , \8131 );
and \U$20042 ( \20385 , \8175 , \8129 );
nor \U$20043 ( \20386 , \20384 , \20385 );
xnor \U$20044 ( \20387 , \20386 , \7813 );
and \U$20045 ( \20388 , \20382 , \20387 );
and \U$20046 ( \20389 , \20378 , \20387 );
or \U$20047 ( \20390 , \20383 , \20388 , \20389 );
and \U$20048 ( \20391 , \6297 , \10611 );
and \U$20049 ( \20392 , \5954 , \10608 );
nor \U$20050 ( \20393 , \20391 , \20392 );
xnor \U$20051 ( \20394 , \20393 , \9556 );
and \U$20052 ( \20395 , \6802 , \9798 );
and \U$20053 ( \20396 , \6499 , \9796 );
nor \U$20054 ( \20397 , \20395 , \20396 );
xnor \U$20055 ( \20398 , \20397 , \9559 );
and \U$20056 ( \20399 , \20394 , \20398 );
and \U$20057 ( \20400 , \20398 , \5692 );
and \U$20058 ( \20401 , \20394 , \5692 );
or \U$20059 ( \20402 , \20399 , \20400 , \20401 );
and \U$20060 ( \20403 , \20390 , \20402 );
and \U$20061 ( \20404 , \9347 , \7564 );
and \U$20062 ( \20405 , \8778 , \7562 );
nor \U$20063 ( \20406 , \20404 , \20405 );
xnor \U$20064 ( \20407 , \20406 , \7315 );
and \U$20065 ( \20408 , \9958 , \7035 );
and \U$20066 ( \20409 , \9355 , \7033 );
nor \U$20067 ( \20410 , \20408 , \20409 );
xnor \U$20068 ( \20411 , \20410 , \6775 );
and \U$20069 ( \20412 , \20407 , \20411 );
and \U$20070 ( \20413 , \10144 , \6541 );
and \U$20071 ( \20414 , \9963 , \6539 );
nor \U$20072 ( \20415 , \20413 , \20414 );
xnor \U$20073 ( \20416 , \20415 , \6226 );
and \U$20074 ( \20417 , \20411 , \20416 );
and \U$20075 ( \20418 , \20407 , \20416 );
or \U$20076 ( \20419 , \20412 , \20417 , \20418 );
and \U$20077 ( \20420 , \20402 , \20419 );
and \U$20078 ( \20421 , \20390 , \20419 );
or \U$20079 ( \20422 , \20403 , \20420 , \20421 );
xor \U$20080 ( \20423 , \20290 , \20294 );
xor \U$20081 ( \20424 , \20423 , \20299 );
xor \U$20082 ( \20425 , \20306 , \20310 );
xor \U$20083 ( \20426 , \20425 , \20315 );
and \U$20084 ( \20427 , \20424 , \20426 );
xor \U$20085 ( \20428 , \20323 , \20327 );
xor \U$20086 ( \20429 , \20428 , \20332 );
and \U$20087 ( \20430 , \20426 , \20429 );
and \U$20088 ( \20431 , \20424 , \20429 );
or \U$20089 ( \20432 , \20427 , \20430 , \20431 );
and \U$20090 ( \20433 , \20422 , \20432 );
xor \U$20091 ( \20434 , \20227 , \20231 );
xor \U$20092 ( \20435 , \20434 , \20236 );
and \U$20093 ( \20436 , \20432 , \20435 );
and \U$20094 ( \20437 , \20422 , \20435 );
or \U$20095 ( \20438 , \20433 , \20436 , \20437 );
xor \U$20096 ( \20439 , \20198 , \20202 );
xor \U$20097 ( \20440 , \20439 , \5202 );
xor \U$20098 ( \20441 , \20302 , \20318 );
xor \U$20099 ( \20442 , \20441 , \20335 );
and \U$20100 ( \20443 , \20440 , \20442 );
xor \U$20101 ( \20444 , \20342 , \20344 );
xor \U$20102 ( \20445 , \20444 , \20347 );
and \U$20103 ( \20446 , \20442 , \20445 );
and \U$20104 ( \20447 , \20440 , \20445 );
or \U$20105 ( \20448 , \20443 , \20446 , \20447 );
and \U$20106 ( \20449 , \20438 , \20448 );
xor \U$20107 ( \20450 , \20246 , \20248 );
xor \U$20108 ( \20451 , \20450 , \20251 );
and \U$20109 ( \20452 , \20448 , \20451 );
and \U$20110 ( \20453 , \20438 , \20451 );
or \U$20111 ( \20454 , \20449 , \20452 , \20453 );
xor \U$20112 ( \20455 , \20206 , \20222 );
xor \U$20113 ( \20456 , \20455 , \20239 );
xor \U$20114 ( \20457 , \20338 , \20350 );
xor \U$20115 ( \20458 , \20457 , \20353 );
and \U$20116 ( \20459 , \20456 , \20458 );
and \U$20117 ( \20460 , \20454 , \20459 );
xor \U$20118 ( \20461 , \20356 , \20358 );
xor \U$20119 ( \20462 , \20461 , \20360 );
and \U$20120 ( \20463 , \20459 , \20462 );
and \U$20121 ( \20464 , \20454 , \20462 );
or \U$20122 ( \20465 , \20460 , \20463 , \20464 );
and \U$20123 ( \20466 , \20374 , \20465 );
xor \U$20124 ( \20467 , \20374 , \20465 );
xor \U$20125 ( \20468 , \20454 , \20459 );
xor \U$20126 ( \20469 , \20468 , \20462 );
and \U$20127 ( \20470 , \6499 , \10611 );
and \U$20128 ( \20471 , \6297 , \10608 );
nor \U$20129 ( \20472 , \20470 , \20471 );
xnor \U$20130 ( \20473 , \20472 , \9556 );
and \U$20131 ( \20474 , \6974 , \9798 );
and \U$20132 ( \20475 , \6802 , \9796 );
nor \U$20133 ( \20476 , \20474 , \20475 );
xnor \U$20134 ( \20477 , \20476 , \9559 );
and \U$20135 ( \20478 , \20473 , \20477 );
and \U$20136 ( \20479 , \7924 , \9230 );
and \U$20137 ( \20480 , \7500 , \9228 );
nor \U$20138 ( \20481 , \20479 , \20480 );
xnor \U$20139 ( \20482 , \20481 , \8920 );
and \U$20140 ( \20483 , \20477 , \20482 );
and \U$20141 ( \20484 , \20473 , \20482 );
or \U$20142 ( \20485 , \20478 , \20483 , \20484 );
and \U$20143 ( \20486 , \8175 , \8693 );
and \U$20144 ( \20487 , \8170 , \8691 );
nor \U$20145 ( \20488 , \20486 , \20487 );
xnor \U$20146 ( \20489 , \20488 , \8322 );
and \U$20147 ( \20490 , \8778 , \8131 );
and \U$20148 ( \20491 , \8494 , \8129 );
nor \U$20149 ( \20492 , \20490 , \20491 );
xnor \U$20150 ( \20493 , \20492 , \7813 );
and \U$20151 ( \20494 , \20489 , \20493 );
and \U$20152 ( \20495 , \9355 , \7564 );
and \U$20153 ( \20496 , \9347 , \7562 );
nor \U$20154 ( \20497 , \20495 , \20496 );
xnor \U$20155 ( \20498 , \20497 , \7315 );
and \U$20156 ( \20499 , \20493 , \20498 );
and \U$20157 ( \20500 , \20489 , \20498 );
or \U$20158 ( \20501 , \20494 , \20499 , \20500 );
and \U$20159 ( \20502 , \20485 , \20501 );
and \U$20160 ( \20503 , \9963 , \7035 );
and \U$20161 ( \20504 , \9958 , \7033 );
nor \U$20162 ( \20505 , \20503 , \20504 );
xnor \U$20163 ( \20506 , \20505 , \6775 );
and \U$20164 ( \20507 , \10764 , \6541 );
and \U$20165 ( \20508 , \10144 , \6539 );
nor \U$20166 ( \20509 , \20507 , \20508 );
xnor \U$20167 ( \20510 , \20509 , \6226 );
and \U$20168 ( \20511 , \20506 , \20510 );
and \U$20169 ( \20512 , \20501 , \20511 );
and \U$20170 ( \20513 , \20485 , \20511 );
or \U$20171 ( \20514 , \20502 , \20512 , \20513 );
nand \U$20172 ( \20515 , \10764 , \6030 );
xnor \U$20173 ( \20516 , \20515 , \5692 );
xor \U$20174 ( \20517 , \20378 , \20382 );
xor \U$20175 ( \20518 , \20517 , \20387 );
and \U$20176 ( \20519 , \20516 , \20518 );
xor \U$20177 ( \20520 , \20407 , \20411 );
xor \U$20178 ( \20521 , \20520 , \20416 );
and \U$20179 ( \20522 , \20518 , \20521 );
and \U$20180 ( \20523 , \20516 , \20521 );
or \U$20181 ( \20524 , \20519 , \20522 , \20523 );
and \U$20182 ( \20525 , \20514 , \20524 );
xor \U$20183 ( \20526 , \20424 , \20426 );
xor \U$20184 ( \20527 , \20526 , \20429 );
and \U$20185 ( \20528 , \20524 , \20527 );
and \U$20186 ( \20529 , \20514 , \20527 );
or \U$20187 ( \20530 , \20525 , \20528 , \20529 );
xor \U$20188 ( \20531 , \20422 , \20432 );
xor \U$20189 ( \20532 , \20531 , \20435 );
and \U$20190 ( \20533 , \20530 , \20532 );
xor \U$20191 ( \20534 , \20440 , \20442 );
xor \U$20192 ( \20535 , \20534 , \20445 );
and \U$20193 ( \20536 , \20532 , \20535 );
and \U$20194 ( \20537 , \20530 , \20535 );
or \U$20195 ( \20538 , \20533 , \20536 , \20537 );
xor \U$20196 ( \20539 , \20438 , \20448 );
xor \U$20197 ( \20540 , \20539 , \20451 );
and \U$20198 ( \20541 , \20538 , \20540 );
xor \U$20199 ( \20542 , \20456 , \20458 );
and \U$20200 ( \20543 , \20540 , \20542 );
and \U$20201 ( \20544 , \20538 , \20542 );
or \U$20202 ( \20545 , \20541 , \20543 , \20544 );
and \U$20203 ( \20546 , \20469 , \20545 );
xor \U$20204 ( \20547 , \20469 , \20545 );
xor \U$20205 ( \20548 , \20538 , \20540 );
xor \U$20206 ( \20549 , \20548 , \20542 );
and \U$20207 ( \20550 , \9958 , \7564 );
and \U$20208 ( \20551 , \9355 , \7562 );
nor \U$20209 ( \20552 , \20550 , \20551 );
xnor \U$20210 ( \20553 , \20552 , \7315 );
and \U$20211 ( \20554 , \10144 , \7035 );
and \U$20212 ( \20555 , \9963 , \7033 );
nor \U$20213 ( \20556 , \20554 , \20555 );
xnor \U$20214 ( \20557 , \20556 , \6775 );
and \U$20215 ( \20558 , \20553 , \20557 );
nand \U$20216 ( \20559 , \10764 , \6539 );
xnor \U$20217 ( \20560 , \20559 , \6226 );
and \U$20218 ( \20561 , \20557 , \20560 );
and \U$20219 ( \20562 , \20553 , \20560 );
or \U$20220 ( \20563 , \20558 , \20561 , \20562 );
and \U$20221 ( \20564 , \6802 , \10611 );
and \U$20222 ( \20565 , \6499 , \10608 );
nor \U$20223 ( \20566 , \20564 , \20565 );
xnor \U$20224 ( \20567 , \20566 , \9556 );
and \U$20225 ( \20568 , \7500 , \9798 );
and \U$20226 ( \20569 , \6974 , \9796 );
nor \U$20227 ( \20570 , \20568 , \20569 );
xnor \U$20228 ( \20571 , \20570 , \9559 );
and \U$20229 ( \20572 , \20567 , \20571 );
and \U$20230 ( \20573 , \20571 , \6226 );
and \U$20231 ( \20574 , \20567 , \6226 );
or \U$20232 ( \20575 , \20572 , \20573 , \20574 );
and \U$20233 ( \20576 , \20563 , \20575 );
and \U$20234 ( \20577 , \8170 , \9230 );
and \U$20235 ( \20578 , \7924 , \9228 );
nor \U$20236 ( \20579 , \20577 , \20578 );
xnor \U$20237 ( \20580 , \20579 , \8920 );
and \U$20238 ( \20581 , \8494 , \8693 );
and \U$20239 ( \20582 , \8175 , \8691 );
nor \U$20240 ( \20583 , \20581 , \20582 );
xnor \U$20241 ( \20584 , \20583 , \8322 );
and \U$20242 ( \20585 , \20580 , \20584 );
and \U$20243 ( \20586 , \9347 , \8131 );
and \U$20244 ( \20587 , \8778 , \8129 );
nor \U$20245 ( \20588 , \20586 , \20587 );
xnor \U$20246 ( \20589 , \20588 , \7813 );
and \U$20247 ( \20590 , \20584 , \20589 );
and \U$20248 ( \20591 , \20580 , \20589 );
or \U$20249 ( \20592 , \20585 , \20590 , \20591 );
and \U$20250 ( \20593 , \20575 , \20592 );
and \U$20251 ( \20594 , \20563 , \20592 );
or \U$20252 ( \20595 , \20576 , \20593 , \20594 );
xor \U$20253 ( \20596 , \20473 , \20477 );
xor \U$20254 ( \20597 , \20596 , \20482 );
xor \U$20255 ( \20598 , \20489 , \20493 );
xor \U$20256 ( \20599 , \20598 , \20498 );
and \U$20257 ( \20600 , \20597 , \20599 );
xor \U$20258 ( \20601 , \20506 , \20510 );
and \U$20259 ( \20602 , \20599 , \20601 );
and \U$20260 ( \20603 , \20597 , \20601 );
or \U$20261 ( \20604 , \20600 , \20602 , \20603 );
and \U$20262 ( \20605 , \20595 , \20604 );
xor \U$20263 ( \20606 , \20394 , \20398 );
xor \U$20264 ( \20607 , \20606 , \5692 );
and \U$20265 ( \20608 , \20604 , \20607 );
and \U$20266 ( \20609 , \20595 , \20607 );
or \U$20267 ( \20610 , \20605 , \20608 , \20609 );
xor \U$20268 ( \20611 , \20485 , \20501 );
xor \U$20269 ( \20612 , \20611 , \20511 );
xor \U$20270 ( \20613 , \20516 , \20518 );
xor \U$20271 ( \20614 , \20613 , \20521 );
and \U$20272 ( \20615 , \20612 , \20614 );
and \U$20273 ( \20616 , \20610 , \20615 );
xor \U$20274 ( \20617 , \20390 , \20402 );
xor \U$20275 ( \20618 , \20617 , \20419 );
and \U$20276 ( \20619 , \20615 , \20618 );
and \U$20277 ( \20620 , \20610 , \20618 );
or \U$20278 ( \20621 , \20616 , \20619 , \20620 );
xor \U$20279 ( \20622 , \20530 , \20532 );
xor \U$20280 ( \20623 , \20622 , \20535 );
and \U$20281 ( \20624 , \20621 , \20623 );
and \U$20282 ( \20625 , \20549 , \20624 );
xor \U$20283 ( \20626 , \20549 , \20624 );
xor \U$20284 ( \20627 , \20621 , \20623 );
xor \U$20285 ( \20628 , \20610 , \20615 );
xor \U$20286 ( \20629 , \20628 , \20618 );
xor \U$20287 ( \20630 , \20514 , \20524 );
xor \U$20288 ( \20631 , \20630 , \20527 );
and \U$20289 ( \20632 , \20629 , \20631 );
and \U$20290 ( \20633 , \20627 , \20632 );
xor \U$20291 ( \20634 , \20627 , \20632 );
xor \U$20292 ( \20635 , \20629 , \20631 );
and \U$20293 ( \20636 , \6974 , \10611 );
and \U$20294 ( \20637 , \6802 , \10608 );
nor \U$20295 ( \20638 , \20636 , \20637 );
xnor \U$20296 ( \20639 , \20638 , \9556 );
and \U$20297 ( \20640 , \7924 , \9798 );
and \U$20298 ( \20641 , \7500 , \9796 );
nor \U$20299 ( \20642 , \20640 , \20641 );
xnor \U$20300 ( \20643 , \20642 , \9559 );
and \U$20301 ( \20644 , \20639 , \20643 );
and \U$20302 ( \20645 , \8175 , \9230 );
and \U$20303 ( \20646 , \8170 , \9228 );
nor \U$20304 ( \20647 , \20645 , \20646 );
xnor \U$20305 ( \20648 , \20647 , \8920 );
and \U$20306 ( \20649 , \20643 , \20648 );
and \U$20307 ( \20650 , \20639 , \20648 );
or \U$20308 ( \20651 , \20644 , \20649 , \20650 );
and \U$20309 ( \20652 , \8778 , \8693 );
and \U$20310 ( \20653 , \8494 , \8691 );
nor \U$20311 ( \20654 , \20652 , \20653 );
xnor \U$20312 ( \20655 , \20654 , \8322 );
and \U$20313 ( \20656 , \9355 , \8131 );
and \U$20314 ( \20657 , \9347 , \8129 );
nor \U$20315 ( \20658 , \20656 , \20657 );
xnor \U$20316 ( \20659 , \20658 , \7813 );
and \U$20317 ( \20660 , \20655 , \20659 );
and \U$20318 ( \20661 , \9963 , \7564 );
and \U$20319 ( \20662 , \9958 , \7562 );
nor \U$20320 ( \20663 , \20661 , \20662 );
xnor \U$20321 ( \20664 , \20663 , \7315 );
and \U$20322 ( \20665 , \20659 , \20664 );
and \U$20323 ( \20666 , \20655 , \20664 );
or \U$20324 ( \20667 , \20660 , \20665 , \20666 );
and \U$20325 ( \20668 , \20651 , \20667 );
xor \U$20326 ( \20669 , \20553 , \20557 );
xor \U$20327 ( \20670 , \20669 , \20560 );
and \U$20328 ( \20671 , \20667 , \20670 );
and \U$20329 ( \20672 , \20651 , \20670 );
or \U$20330 ( \20673 , \20668 , \20671 , \20672 );
xor \U$20331 ( \20674 , \20567 , \20571 );
xor \U$20332 ( \20675 , \20674 , \6226 );
xor \U$20333 ( \20676 , \20580 , \20584 );
xor \U$20334 ( \20677 , \20676 , \20589 );
and \U$20335 ( \20678 , \20675 , \20677 );
and \U$20336 ( \20679 , \20673 , \20678 );
xor \U$20337 ( \20680 , \20597 , \20599 );
xor \U$20338 ( \20681 , \20680 , \20601 );
and \U$20339 ( \20682 , \20678 , \20681 );
and \U$20340 ( \20683 , \20673 , \20681 );
or \U$20341 ( \20684 , \20679 , \20682 , \20683 );
xor \U$20342 ( \20685 , \20595 , \20604 );
xor \U$20343 ( \20686 , \20685 , \20607 );
and \U$20344 ( \20687 , \20684 , \20686 );
xor \U$20345 ( \20688 , \20612 , \20614 );
and \U$20346 ( \20689 , \20686 , \20688 );
and \U$20347 ( \20690 , \20684 , \20688 );
or \U$20348 ( \20691 , \20687 , \20689 , \20690 );
and \U$20349 ( \20692 , \20635 , \20691 );
xor \U$20350 ( \20693 , \20635 , \20691 );
xor \U$20351 ( \20694 , \20684 , \20686 );
xor \U$20352 ( \20695 , \20694 , \20688 );
and \U$20353 ( \20696 , \7500 , \10611 );
and \U$20354 ( \20697 , \6974 , \10608 );
nor \U$20355 ( \20698 , \20696 , \20697 );
xnor \U$20356 ( \20699 , \20698 , \9556 );
and \U$20357 ( \20700 , \8170 , \9798 );
and \U$20358 ( \20701 , \7924 , \9796 );
nor \U$20359 ( \20702 , \20700 , \20701 );
xnor \U$20360 ( \20703 , \20702 , \9559 );
and \U$20361 ( \20704 , \20699 , \20703 );
and \U$20362 ( \20705 , \20703 , \6775 );
and \U$20363 ( \20706 , \20699 , \6775 );
or \U$20364 ( \20707 , \20704 , \20705 , \20706 );
and \U$20365 ( \20708 , \8494 , \9230 );
and \U$20366 ( \20709 , \8175 , \9228 );
nor \U$20367 ( \20710 , \20708 , \20709 );
xnor \U$20368 ( \20711 , \20710 , \8920 );
and \U$20369 ( \20712 , \9347 , \8693 );
and \U$20370 ( \20713 , \8778 , \8691 );
nor \U$20371 ( \20714 , \20712 , \20713 );
xnor \U$20372 ( \20715 , \20714 , \8322 );
and \U$20373 ( \20716 , \20711 , \20715 );
and \U$20374 ( \20717 , \9958 , \8131 );
and \U$20375 ( \20718 , \9355 , \8129 );
nor \U$20376 ( \20719 , \20717 , \20718 );
xnor \U$20377 ( \20720 , \20719 , \7813 );
and \U$20378 ( \20721 , \20715 , \20720 );
and \U$20379 ( \20722 , \20711 , \20720 );
or \U$20380 ( \20723 , \20716 , \20721 , \20722 );
and \U$20381 ( \20724 , \20707 , \20723 );
and \U$20382 ( \20725 , \10764 , \7035 );
and \U$20383 ( \20726 , \10144 , \7033 );
nor \U$20384 ( \20727 , \20725 , \20726 );
xnor \U$20385 ( \20728 , \20727 , \6775 );
and \U$20386 ( \20729 , \20723 , \20728 );
and \U$20387 ( \20730 , \20707 , \20728 );
or \U$20388 ( \20731 , \20724 , \20729 , \20730 );
xor \U$20389 ( \20732 , \20651 , \20667 );
xor \U$20390 ( \20733 , \20732 , \20670 );
and \U$20391 ( \20734 , \20731 , \20733 );
xor \U$20392 ( \20735 , \20675 , \20677 );
and \U$20393 ( \20736 , \20733 , \20735 );
and \U$20394 ( \20737 , \20731 , \20735 );
or \U$20395 ( \20738 , \20734 , \20736 , \20737 );
xor \U$20396 ( \20739 , \20563 , \20575 );
xor \U$20397 ( \20740 , \20739 , \20592 );
and \U$20398 ( \20741 , \20738 , \20740 );
xor \U$20399 ( \20742 , \20673 , \20678 );
xor \U$20400 ( \20743 , \20742 , \20681 );
and \U$20401 ( \20744 , \20740 , \20743 );
and \U$20402 ( \20745 , \20738 , \20743 );
or \U$20403 ( \20746 , \20741 , \20744 , \20745 );
and \U$20404 ( \20747 , \20695 , \20746 );
xor \U$20405 ( \20748 , \20695 , \20746 );
xor \U$20406 ( \20749 , \20738 , \20740 );
xor \U$20407 ( \20750 , \20749 , \20743 );
and \U$20408 ( \20751 , \9355 , \8693 );
and \U$20409 ( \20752 , \9347 , \8691 );
nor \U$20410 ( \20753 , \20751 , \20752 );
xnor \U$20411 ( \20754 , \20753 , \8322 );
and \U$20412 ( \20755 , \9963 , \8131 );
and \U$20413 ( \20756 , \9958 , \8129 );
nor \U$20414 ( \20757 , \20755 , \20756 );
xnor \U$20415 ( \20758 , \20757 , \7813 );
and \U$20416 ( \20759 , \20754 , \20758 );
and \U$20417 ( \20760 , \10764 , \7564 );
and \U$20418 ( \20761 , \10144 , \7562 );
nor \U$20419 ( \20762 , \20760 , \20761 );
xnor \U$20420 ( \20763 , \20762 , \7315 );
and \U$20421 ( \20764 , \20758 , \20763 );
and \U$20422 ( \20765 , \20754 , \20763 );
or \U$20423 ( \20766 , \20759 , \20764 , \20765 );
and \U$20424 ( \20767 , \7924 , \10611 );
and \U$20425 ( \20768 , \7500 , \10608 );
nor \U$20426 ( \20769 , \20767 , \20768 );
xnor \U$20427 ( \20770 , \20769 , \9556 );
and \U$20428 ( \20771 , \8175 , \9798 );
and \U$20429 ( \20772 , \8170 , \9796 );
nor \U$20430 ( \20773 , \20771 , \20772 );
xnor \U$20431 ( \20774 , \20773 , \9559 );
and \U$20432 ( \20775 , \20770 , \20774 );
and \U$20433 ( \20776 , \8778 , \9230 );
and \U$20434 ( \20777 , \8494 , \9228 );
nor \U$20435 ( \20778 , \20776 , \20777 );
xnor \U$20436 ( \20779 , \20778 , \8920 );
and \U$20437 ( \20780 , \20774 , \20779 );
and \U$20438 ( \20781 , \20770 , \20779 );
or \U$20439 ( \20782 , \20775 , \20780 , \20781 );
and \U$20440 ( \20783 , \20766 , \20782 );
and \U$20441 ( \20784 , \10144 , \7564 );
and \U$20442 ( \20785 , \9963 , \7562 );
nor \U$20443 ( \20786 , \20784 , \20785 );
xnor \U$20444 ( \20787 , \20786 , \7315 );
and \U$20445 ( \20788 , \20782 , \20787 );
and \U$20446 ( \20789 , \20766 , \20787 );
or \U$20447 ( \20790 , \20783 , \20788 , \20789 );
nand \U$20448 ( \20791 , \10764 , \7033 );
xnor \U$20449 ( \20792 , \20791 , \6775 );
xor \U$20450 ( \20793 , \20699 , \20703 );
xor \U$20451 ( \20794 , \20793 , \6775 );
and \U$20452 ( \20795 , \20792 , \20794 );
xor \U$20453 ( \20796 , \20711 , \20715 );
xor \U$20454 ( \20797 , \20796 , \20720 );
and \U$20455 ( \20798 , \20794 , \20797 );
and \U$20456 ( \20799 , \20792 , \20797 );
or \U$20457 ( \20800 , \20795 , \20798 , \20799 );
and \U$20458 ( \20801 , \20790 , \20800 );
xor \U$20459 ( \20802 , \20655 , \20659 );
xor \U$20460 ( \20803 , \20802 , \20664 );
and \U$20461 ( \20804 , \20800 , \20803 );
and \U$20462 ( \20805 , \20790 , \20803 );
or \U$20463 ( \20806 , \20801 , \20804 , \20805 );
xor \U$20464 ( \20807 , \20639 , \20643 );
xor \U$20465 ( \20808 , \20807 , \20648 );
xor \U$20466 ( \20809 , \20707 , \20723 );
xor \U$20467 ( \20810 , \20809 , \20728 );
and \U$20468 ( \20811 , \20808 , \20810 );
and \U$20469 ( \20812 , \20806 , \20811 );
xor \U$20470 ( \20813 , \20731 , \20733 );
xor \U$20471 ( \20814 , \20813 , \20735 );
and \U$20472 ( \20815 , \20811 , \20814 );
and \U$20473 ( \20816 , \20806 , \20814 );
or \U$20474 ( \20817 , \20812 , \20815 , \20816 );
and \U$20475 ( \20818 , \20750 , \20817 );
xor \U$20476 ( \20819 , \20750 , \20817 );
xor \U$20477 ( \20820 , \20806 , \20811 );
xor \U$20478 ( \20821 , \20820 , \20814 );
and \U$20479 ( \20822 , \9347 , \9230 );
and \U$20480 ( \20823 , \8778 , \9228 );
nor \U$20481 ( \20824 , \20822 , \20823 );
xnor \U$20482 ( \20825 , \20824 , \8920 );
and \U$20483 ( \20826 , \9958 , \8693 );
and \U$20484 ( \20827 , \9355 , \8691 );
nor \U$20485 ( \20828 , \20826 , \20827 );
xnor \U$20486 ( \20829 , \20828 , \8322 );
and \U$20487 ( \20830 , \20825 , \20829 );
and \U$20488 ( \20831 , \10144 , \8131 );
and \U$20489 ( \20832 , \9963 , \8129 );
nor \U$20490 ( \20833 , \20831 , \20832 );
xnor \U$20491 ( \20834 , \20833 , \7813 );
and \U$20492 ( \20835 , \20829 , \20834 );
and \U$20493 ( \20836 , \20825 , \20834 );
or \U$20494 ( \20837 , \20830 , \20835 , \20836 );
and \U$20495 ( \20838 , \8170 , \10611 );
and \U$20496 ( \20839 , \7924 , \10608 );
nor \U$20497 ( \20840 , \20838 , \20839 );
xnor \U$20498 ( \20841 , \20840 , \9556 );
and \U$20499 ( \20842 , \8494 , \9798 );
and \U$20500 ( \20843 , \8175 , \9796 );
nor \U$20501 ( \20844 , \20842 , \20843 );
xnor \U$20502 ( \20845 , \20844 , \9559 );
and \U$20503 ( \20846 , \20841 , \20845 );
and \U$20504 ( \20847 , \20845 , \7315 );
and \U$20505 ( \20848 , \20841 , \7315 );
or \U$20506 ( \20849 , \20846 , \20847 , \20848 );
and \U$20507 ( \20850 , \20837 , \20849 );
xor \U$20508 ( \20851 , \20754 , \20758 );
xor \U$20509 ( \20852 , \20851 , \20763 );
and \U$20510 ( \20853 , \20849 , \20852 );
and \U$20511 ( \20854 , \20837 , \20852 );
or \U$20512 ( \20855 , \20850 , \20853 , \20854 );
xor \U$20513 ( \20856 , \20766 , \20782 );
xor \U$20514 ( \20857 , \20856 , \20787 );
and \U$20515 ( \20858 , \20855 , \20857 );
xor \U$20516 ( \20859 , \20792 , \20794 );
xor \U$20517 ( \20860 , \20859 , \20797 );
and \U$20518 ( \20861 , \20857 , \20860 );
and \U$20519 ( \20862 , \20855 , \20860 );
or \U$20520 ( \20863 , \20858 , \20861 , \20862 );
xor \U$20521 ( \20864 , \20790 , \20800 );
xor \U$20522 ( \20865 , \20864 , \20803 );
and \U$20523 ( \20866 , \20863 , \20865 );
xor \U$20524 ( \20867 , \20808 , \20810 );
and \U$20525 ( \20868 , \20865 , \20867 );
and \U$20526 ( \20869 , \20863 , \20867 );
or \U$20527 ( \20870 , \20866 , \20868 , \20869 );
and \U$20528 ( \20871 , \20821 , \20870 );
xor \U$20529 ( \20872 , \20821 , \20870 );
xor \U$20530 ( \20873 , \20863 , \20865 );
xor \U$20531 ( \20874 , \20873 , \20867 );
and \U$20532 ( \20875 , \8175 , \10611 );
and \U$20533 ( \20876 , \8170 , \10608 );
nor \U$20534 ( \20877 , \20875 , \20876 );
xnor \U$20535 ( \20878 , \20877 , \9556 );
and \U$20536 ( \20879 , \8778 , \9798 );
and \U$20537 ( \20880 , \8494 , \9796 );
nor \U$20538 ( \20881 , \20879 , \20880 );
xnor \U$20539 ( \20882 , \20881 , \9559 );
and \U$20540 ( \20883 , \20878 , \20882 );
and \U$20541 ( \20884 , \9355 , \9230 );
and \U$20542 ( \20885 , \9347 , \9228 );
nor \U$20543 ( \20886 , \20884 , \20885 );
xnor \U$20544 ( \20887 , \20886 , \8920 );
and \U$20545 ( \20888 , \20882 , \20887 );
and \U$20546 ( \20889 , \20878 , \20887 );
or \U$20547 ( \20890 , \20883 , \20888 , \20889 );
nand \U$20548 ( \20891 , \10764 , \7562 );
xnor \U$20549 ( \20892 , \20891 , \7315 );
and \U$20550 ( \20893 , \20890 , \20892 );
xor \U$20551 ( \20894 , \20825 , \20829 );
xor \U$20552 ( \20895 , \20894 , \20834 );
and \U$20553 ( \20896 , \20892 , \20895 );
and \U$20554 ( \20897 , \20890 , \20895 );
or \U$20555 ( \20898 , \20893 , \20896 , \20897 );
xor \U$20556 ( \20899 , \20770 , \20774 );
xor \U$20557 ( \20900 , \20899 , \20779 );
and \U$20558 ( \20901 , \20898 , \20900 );
xor \U$20559 ( \20902 , \20837 , \20849 );
xor \U$20560 ( \20903 , \20902 , \20852 );
and \U$20561 ( \20904 , \20900 , \20903 );
and \U$20562 ( \20905 , \20898 , \20903 );
or \U$20563 ( \20906 , \20901 , \20904 , \20905 );
xor \U$20564 ( \20907 , \20855 , \20857 );
xor \U$20565 ( \20908 , \20907 , \20860 );
and \U$20566 ( \20909 , \20906 , \20908 );
and \U$20567 ( \20910 , \20874 , \20909 );
xor \U$20568 ( \20911 , \20874 , \20909 );
xor \U$20569 ( \20912 , \20906 , \20908 );
and \U$20570 ( \20913 , \9958 , \9230 );
and \U$20571 ( \20914 , \9355 , \9228 );
nor \U$20572 ( \20915 , \20913 , \20914 );
xnor \U$20573 ( \20916 , \20915 , \8920 );
and \U$20574 ( \20917 , \10144 , \8693 );
and \U$20575 ( \20918 , \9963 , \8691 );
nor \U$20576 ( \20919 , \20917 , \20918 );
xnor \U$20577 ( \20920 , \20919 , \8322 );
and \U$20578 ( \20921 , \20916 , \20920 );
nand \U$20579 ( \20922 , \10764 , \8129 );
xnor \U$20580 ( \20923 , \20922 , \7813 );
and \U$20581 ( \20924 , \20920 , \20923 );
and \U$20582 ( \20925 , \20916 , \20923 );
or \U$20583 ( \20926 , \20921 , \20924 , \20925 );
and \U$20584 ( \20927 , \8494 , \10611 );
and \U$20585 ( \20928 , \8175 , \10608 );
nor \U$20586 ( \20929 , \20927 , \20928 );
xnor \U$20587 ( \20930 , \20929 , \9556 );
and \U$20588 ( \20931 , \9347 , \9798 );
and \U$20589 ( \20932 , \8778 , \9796 );
nor \U$20590 ( \20933 , \20931 , \20932 );
xnor \U$20591 ( \20934 , \20933 , \9559 );
and \U$20592 ( \20935 , \20930 , \20934 );
and \U$20593 ( \20936 , \20934 , \7813 );
and \U$20594 ( \20937 , \20930 , \7813 );
or \U$20595 ( \20938 , \20935 , \20936 , \20937 );
and \U$20596 ( \20939 , \20926 , \20938 );
and \U$20597 ( \20940 , \9963 , \8693 );
and \U$20598 ( \20941 , \9958 , \8691 );
nor \U$20599 ( \20942 , \20940 , \20941 );
xnor \U$20600 ( \20943 , \20942 , \8322 );
and \U$20601 ( \20944 , \20938 , \20943 );
and \U$20602 ( \20945 , \20926 , \20943 );
or \U$20603 ( \20946 , \20939 , \20944 , \20945 );
and \U$20604 ( \20947 , \10764 , \8131 );
and \U$20605 ( \20948 , \10144 , \8129 );
nor \U$20606 ( \20949 , \20947 , \20948 );
xnor \U$20607 ( \20950 , \20949 , \7813 );
xor \U$20608 ( \20951 , \20878 , \20882 );
xor \U$20609 ( \20952 , \20951 , \20887 );
and \U$20610 ( \20953 , \20950 , \20952 );
and \U$20611 ( \20954 , \20946 , \20953 );
xor \U$20612 ( \20955 , \20841 , \20845 );
xor \U$20613 ( \20956 , \20955 , \7315 );
and \U$20614 ( \20957 , \20953 , \20956 );
and \U$20615 ( \20958 , \20946 , \20956 );
or \U$20616 ( \20959 , \20954 , \20957 , \20958 );
xor \U$20617 ( \20960 , \20898 , \20900 );
xor \U$20618 ( \20961 , \20960 , \20903 );
and \U$20619 ( \20962 , \20959 , \20961 );
and \U$20620 ( \20963 , \20912 , \20962 );
xor \U$20621 ( \20964 , \20912 , \20962 );
xor \U$20622 ( \20965 , \20959 , \20961 );
xor \U$20623 ( \20966 , \20890 , \20892 );
xor \U$20624 ( \20967 , \20966 , \20895 );
xor \U$20625 ( \20968 , \20946 , \20953 );
xor \U$20626 ( \20969 , \20968 , \20956 );
and \U$20627 ( \20970 , \20967 , \20969 );
and \U$20628 ( \20971 , \20965 , \20970 );
xor \U$20629 ( \20972 , \20965 , \20970 );
xor \U$20630 ( \20973 , \20967 , \20969 );
and \U$20631 ( \20974 , \8778 , \10611 );
and \U$20632 ( \20975 , \8494 , \10608 );
nor \U$20633 ( \20976 , \20974 , \20975 );
xnor \U$20634 ( \20977 , \20976 , \9556 );
and \U$20635 ( \20978 , \9355 , \9798 );
and \U$20636 ( \20979 , \9347 , \9796 );
nor \U$20637 ( \20980 , \20978 , \20979 );
xnor \U$20638 ( \20981 , \20980 , \9559 );
and \U$20639 ( \20982 , \20977 , \20981 );
and \U$20640 ( \20983 , \9963 , \9230 );
and \U$20641 ( \20984 , \9958 , \9228 );
nor \U$20642 ( \20985 , \20983 , \20984 );
xnor \U$20643 ( \20986 , \20985 , \8920 );
and \U$20644 ( \20987 , \20981 , \20986 );
and \U$20645 ( \20988 , \20977 , \20986 );
or \U$20646 ( \20989 , \20982 , \20987 , \20988 );
xor \U$20647 ( \20990 , \20916 , \20920 );
xor \U$20648 ( \20991 , \20990 , \20923 );
and \U$20649 ( \20992 , \20989 , \20991 );
xor \U$20650 ( \20993 , \20930 , \20934 );
xor \U$20651 ( \20994 , \20993 , \7813 );
and \U$20652 ( \20995 , \20991 , \20994 );
and \U$20653 ( \20996 , \20989 , \20994 );
or \U$20654 ( \20997 , \20992 , \20995 , \20996 );
xor \U$20655 ( \20998 , \20926 , \20938 );
xor \U$20656 ( \20999 , \20998 , \20943 );
and \U$20657 ( \21000 , \20997 , \20999 );
xor \U$20658 ( \21001 , \20950 , \20952 );
and \U$20659 ( \21002 , \20999 , \21001 );
and \U$20660 ( \21003 , \20997 , \21001 );
or \U$20661 ( \21004 , \21000 , \21002 , \21003 );
and \U$20662 ( \21005 , \20973 , \21004 );
xor \U$20663 ( \21006 , \20973 , \21004 );
xor \U$20664 ( \21007 , \20997 , \20999 );
xor \U$20665 ( \21008 , \21007 , \21001 );
and \U$20666 ( \21009 , \9347 , \10611 );
and \U$20667 ( \21010 , \8778 , \10608 );
nor \U$20668 ( \21011 , \21009 , \21010 );
xnor \U$20669 ( \21012 , \21011 , \9556 );
and \U$20670 ( \21013 , \9958 , \9798 );
and \U$20671 ( \21014 , \9355 , \9796 );
nor \U$20672 ( \21015 , \21013 , \21014 );
xnor \U$20673 ( \21016 , \21015 , \9559 );
and \U$20674 ( \21017 , \21012 , \21016 );
and \U$20675 ( \21018 , \21016 , \8322 );
and \U$20676 ( \21019 , \21012 , \8322 );
or \U$20677 ( \21020 , \21017 , \21018 , \21019 );
and \U$20678 ( \21021 , \10144 , \9230 );
and \U$20679 ( \21022 , \9963 , \9228 );
nor \U$20680 ( \21023 , \21021 , \21022 );
xnor \U$20681 ( \21024 , \21023 , \8920 );
nand \U$20682 ( \21025 , \10764 , \8691 );
xnor \U$20683 ( \21026 , \21025 , \8322 );
and \U$20684 ( \21027 , \21024 , \21026 );
and \U$20685 ( \21028 , \21020 , \21027 );
and \U$20686 ( \21029 , \10764 , \8693 );
and \U$20687 ( \21030 , \10144 , \8691 );
nor \U$20688 ( \21031 , \21029 , \21030 );
xnor \U$20689 ( \21032 , \21031 , \8322 );
and \U$20690 ( \21033 , \21027 , \21032 );
and \U$20691 ( \21034 , \21020 , \21032 );
or \U$20692 ( \21035 , \21028 , \21033 , \21034 );
xor \U$20693 ( \21036 , \20989 , \20991 );
xor \U$20694 ( \21037 , \21036 , \20994 );
and \U$20695 ( \21038 , \21035 , \21037 );
and \U$20696 ( \21039 , \21008 , \21038 );
xor \U$20697 ( \21040 , \21008 , \21038 );
xor \U$20698 ( \21041 , \21035 , \21037 );
xor \U$20699 ( \21042 , \20977 , \20981 );
xor \U$20700 ( \21043 , \21042 , \20986 );
xor \U$20701 ( \21044 , \21020 , \21027 );
xor \U$20702 ( \21045 , \21044 , \21032 );
and \U$20703 ( \21046 , \21043 , \21045 );
and \U$20704 ( \21047 , \21041 , \21046 );
xor \U$20705 ( \21048 , \21041 , \21046 );
xor \U$20706 ( \21049 , \21043 , \21045 );
and \U$20707 ( \21050 , \9355 , \10611 );
and \U$20708 ( \21051 , \9347 , \10608 );
nor \U$20709 ( \21052 , \21050 , \21051 );
xnor \U$20710 ( \21053 , \21052 , \9556 );
and \U$20711 ( \21054 , \9963 , \9798 );
and \U$20712 ( \21055 , \9958 , \9796 );
nor \U$20713 ( \21056 , \21054 , \21055 );
xnor \U$20714 ( \21057 , \21056 , \9559 );
and \U$20715 ( \21058 , \21053 , \21057 );
and \U$20716 ( \21059 , \10764 , \9230 );
and \U$20717 ( \21060 , \10144 , \9228 );
nor \U$20718 ( \21061 , \21059 , \21060 );
xnor \U$20719 ( \21062 , \21061 , \8920 );
and \U$20720 ( \21063 , \21057 , \21062 );
and \U$20721 ( \21064 , \21053 , \21062 );
or \U$20722 ( \21065 , \21058 , \21063 , \21064 );
xor \U$20723 ( \21066 , \21012 , \21016 );
xor \U$20724 ( \21067 , \21066 , \8322 );
and \U$20725 ( \21068 , \21065 , \21067 );
xor \U$20726 ( \21069 , \21024 , \21026 );
and \U$20727 ( \21070 , \21067 , \21069 );
and \U$20728 ( \21071 , \21065 , \21069 );
or \U$20729 ( \21072 , \21068 , \21070 , \21071 );
and \U$20730 ( \21073 , \21049 , \21072 );
xor \U$20731 ( \21074 , \21049 , \21072 );
xor \U$20732 ( \21075 , \21065 , \21067 );
xor \U$20733 ( \21076 , \21075 , \21069 );
and \U$20734 ( \21077 , \9958 , \10611 );
and \U$20735 ( \21078 , \9355 , \10608 );
nor \U$20736 ( \21079 , \21077 , \21078 );
xnor \U$20737 ( \21080 , \21079 , \9556 );
and \U$20738 ( \21081 , \10144 , \9798 );
and \U$20739 ( \21082 , \9963 , \9796 );
nor \U$20740 ( \21083 , \21081 , \21082 );
xnor \U$20741 ( \21084 , \21083 , \9559 );
and \U$20742 ( \21085 , \21080 , \21084 );
and \U$20743 ( \21086 , \21084 , \8920 );
and \U$20744 ( \21087 , \21080 , \8920 );
or \U$20745 ( \21088 , \21085 , \21086 , \21087 );
xor \U$20746 ( \21089 , \21053 , \21057 );
xor \U$20747 ( \21090 , \21089 , \21062 );
and \U$20748 ( \21091 , \21088 , \21090 );
and \U$20749 ( \21092 , \21076 , \21091 );
xor \U$20750 ( \21093 , \21076 , \21091 );
xor \U$20751 ( \21094 , \21088 , \21090 );
nand \U$20752 ( \21095 , \10764 , \9228 );
xnor \U$20753 ( \21096 , \21095 , \8920 );
xor \U$20754 ( \21097 , \21080 , \21084 );
xor \U$20755 ( \21098 , \21097 , \8920 );
and \U$20756 ( \21099 , \21096 , \21098 );
and \U$20757 ( \21100 , \21094 , \21099 );
xor \U$20758 ( \21101 , \21094 , \21099 );
xor \U$20759 ( \21102 , \21096 , \21098 );
and \U$20760 ( \21103 , \9963 , \10611 );
and \U$20761 ( \21104 , \9958 , \10608 );
nor \U$20762 ( \21105 , \21103 , \21104 );
xnor \U$20763 ( \21106 , \21105 , \9556 );
and \U$20764 ( \21107 , \10764 , \9798 );
and \U$20765 ( \21108 , \10144 , \9796 );
nor \U$20766 ( \21109 , \21107 , \21108 );
xnor \U$20767 ( \21110 , \21109 , \9559 );
and \U$20768 ( \21111 , \21106 , \21110 );
and \U$20769 ( \21112 , \21102 , \21111 );
xor \U$20770 ( \21113 , \21102 , \21111 );
xor \U$20771 ( \21114 , \21106 , \21110 );
and \U$20772 ( \21115 , \10144 , \10611 );
and \U$20773 ( \21116 , \9963 , \10608 );
nor \U$20774 ( \21117 , \21115 , \21116 );
xnor \U$20775 ( \21118 , \21117 , \9556 );
and \U$20776 ( \21119 , \21118 , \9559 );
and \U$20777 ( \21120 , \21114 , \21119 );
xor \U$20778 ( \21121 , \21114 , \21119 );
nand \U$20779 ( \21122 , \10764 , \9796 );
xnor \U$20780 ( \21123 , \21122 , \9559 );
xor \U$20781 ( \21124 , \21118 , \9559 );
and \U$20782 ( \21125 , \21123 , \21124 );
xor \U$20783 ( \21126 , \21123 , \21124 );
and \U$20784 ( \21127 , \10764 , \10611 );
and \U$20785 ( \21128 , \10144 , \10608 );
nor \U$20786 ( \21129 , \21127 , \21128 );
xnor \U$20787 ( \21130 , \21129 , \9556 );
nand \U$20788 ( \21131 , \10764 , \10608 );
xnor \U$20789 ( \21132 , \21131 , \9556 );
and \U$20790 ( \21133 , \21132 , \9556 );
and \U$20791 ( \21134 , \21130 , \21133 );
and \U$20792 ( \21135 , \21126 , \21134 );
or \U$20793 ( \21136 , \21125 , \21135 );
and \U$20794 ( \21137 , \21121 , \21136 );
or \U$20795 ( \21138 , \21120 , \21137 );
and \U$20796 ( \21139 , \21113 , \21138 );
or \U$20797 ( \21140 , \21112 , \21139 );
and \U$20798 ( \21141 , \21101 , \21140 );
or \U$20799 ( \21142 , \21100 , \21141 );
and \U$20800 ( \21143 , \21093 , \21142 );
or \U$20801 ( \21144 , \21092 , \21143 );
and \U$20802 ( \21145 , \21074 , \21144 );
or \U$20803 ( \21146 , \21073 , \21145 );
and \U$20804 ( \21147 , \21048 , \21146 );
or \U$20805 ( \21148 , \21047 , \21147 );
and \U$20806 ( \21149 , \21040 , \21148 );
or \U$20807 ( \21150 , \21039 , \21149 );
and \U$20808 ( \21151 , \21006 , \21150 );
or \U$20809 ( \21152 , \21005 , \21151 );
and \U$20810 ( \21153 , \20972 , \21152 );
or \U$20811 ( \21154 , \20971 , \21153 );
and \U$20812 ( \21155 , \20964 , \21154 );
or \U$20813 ( \21156 , \20963 , \21155 );
and \U$20814 ( \21157 , \20911 , \21156 );
or \U$20815 ( \21158 , \20910 , \21157 );
and \U$20816 ( \21159 , \20872 , \21158 );
or \U$20817 ( \21160 , \20871 , \21159 );
and \U$20818 ( \21161 , \20819 , \21160 );
or \U$20819 ( \21162 , \20818 , \21161 );
and \U$20820 ( \21163 , \20748 , \21162 );
or \U$20821 ( \21164 , \20747 , \21163 );
and \U$20822 ( \21165 , \20693 , \21164 );
or \U$20823 ( \21166 , \20692 , \21165 );
and \U$20824 ( \21167 , \20634 , \21166 );
or \U$20825 ( \21168 , \20633 , \21167 );
and \U$20826 ( \21169 , \20626 , \21168 );
or \U$20827 ( \21170 , \20625 , \21169 );
and \U$20828 ( \21171 , \20547 , \21170 );
or \U$20829 ( \21172 , \20546 , \21171 );
and \U$20830 ( \21173 , \20467 , \21172 );
or \U$20831 ( \21174 , \20466 , \21173 );
and \U$20832 ( \21175 , \20372 , \21174 );
or \U$20833 ( \21176 , \20371 , \21175 );
and \U$20834 ( \21177 , \20284 , \21176 );
or \U$20835 ( \21178 , \20283 , \21177 );
and \U$20836 ( \21179 , \20192 , \21178 );
or \U$20837 ( \21180 , \20191 , \21179 );
and \U$20838 ( \21181 , \20104 , \21180 );
or \U$20839 ( \21182 , \20103 , \21181 );
and \U$20840 ( \21183 , \19989 , \21182 );
or \U$20841 ( \21184 , \19988 , \21183 );
and \U$20842 ( \21185 , \19893 , \21184 );
or \U$20843 ( \21186 , \19892 , \21185 );
and \U$20844 ( \21187 , \19885 , \21186 );
or \U$20845 ( \21188 , \19884 , \21187 );
and \U$20846 ( \21189 , \19770 , \21188 );
or \U$20847 ( \21190 , \19769 , \21189 );
and \U$20848 ( \21191 , \19646 , \21190 );
or \U$20849 ( \21192 , \19645 , \21191 );
and \U$20850 ( \21193 , \19506 , \21192 );
or \U$20851 ( \21194 , \19505 , \21193 );
and \U$20852 ( \21195 , \19382 , \21194 );
or \U$20853 ( \21196 , \19381 , \21195 );
and \U$20854 ( \21197 , \19238 , \21196 );
or \U$20855 ( \21198 , \19237 , \21197 );
and \U$20856 ( \21199 , \19113 , \21198 );
or \U$20857 ( \21200 , \19112 , \21199 );
and \U$20858 ( \21201 , \18974 , \21200 );
or \U$20859 ( \21202 , \18973 , \21201 );
and \U$20860 ( \21203 , \18810 , \21202 );
or \U$20861 ( \21204 , \18809 , \21203 );
and \U$20862 ( \21205 , \18658 , \21204 );
or \U$20863 ( \21206 , \18657 , \21205 );
and \U$20864 ( \21207 , \18518 , \21206 );
or \U$20865 ( \21208 , \18517 , \21207 );
and \U$20866 ( \21209 , \18350 , \21208 );
or \U$20867 ( \21210 , \18349 , \21209 );
and \U$20868 ( \21211 , \18342 , \21210 );
or \U$20869 ( \21212 , \18341 , \21211 );
and \U$20870 ( \21213 , \18171 , \21212 );
or \U$20871 ( \21214 , \18170 , \21213 );
and \U$20872 ( \21215 , \17995 , \21214 );
or \U$20873 ( \21216 , \17994 , \21215 );
and \U$20874 ( \21217 , \17805 , \21216 );
or \U$20875 ( \21218 , \17804 , \21217 );
and \U$20876 ( \21219 , \17618 , \21218 );
or \U$20877 ( \21220 , \17617 , \21219 );
and \U$20878 ( \21221 , \17433 , \21220 );
or \U$20879 ( \21222 , \17432 , \21221 );
and \U$20880 ( \21223 , \17225 , \21222 );
or \U$20881 ( \21224 , \17224 , \21223 );
and \U$20882 ( \21225 , \17029 , \21224 );
or \U$20883 ( \21226 , \17028 , \21225 );
and \U$20884 ( \21227 , \16832 , \21226 );
or \U$20885 ( \21228 , \16831 , \21227 );
and \U$20886 ( \21229 , \16619 , \21228 );
or \U$20887 ( \21230 , \16618 , \21229 );
and \U$20888 ( \21231 , \16408 , \21230 );
or \U$20889 ( \21232 , \16407 , \21231 );
and \U$20890 ( \21233 , \16177 , \21232 );
or \U$20891 ( \21234 , \16176 , \21233 );
and \U$20892 ( \21235 , \15947 , \21234 );
or \U$20893 ( \21236 , \15946 , \21235 );
and \U$20894 ( \21237 , \15728 , \21236 );
or \U$20895 ( \21238 , \15727 , \21237 );
and \U$20896 ( \21239 , \15503 , \21238 );
or \U$20897 ( \21240 , \15502 , \21239 );
and \U$20898 ( \21241 , \15253 , \21240 );
or \U$20899 ( \21242 , \15252 , \21241 );
and \U$20900 ( \21243 , \15023 , \21242 );
or \U$20901 ( \21244 , \15022 , \21243 );
and \U$20902 ( \21245 , \14777 , \21244 );
or \U$20903 ( \21246 , \14776 , \21245 );
and \U$20904 ( \21247 , \14769 , \21246 );
or \U$20905 ( \21248 , \14768 , \21247 );
and \U$20906 ( \21249 , \14508 , \21248 );
or \U$20907 ( \21250 , \14507 , \21249 );
and \U$20908 ( \21251 , \14246 , \21250 );
or \U$20909 ( \21252 , \14245 , \21251 );
and \U$20910 ( \21253 , \13976 , \21252 );
or \U$20911 ( \21254 , \13975 , \21253 );
and \U$20912 ( \21255 , \13699 , \21254 );
or \U$20913 ( \21256 , \13698 , \21255 );
and \U$20914 ( \21257 , \13423 , \21256 );
or \U$20915 ( \21258 , \13422 , \21257 );
and \U$20916 ( \21259 , \13152 , \21258 );
or \U$20917 ( \21260 , \13151 , \21259 );
and \U$20918 ( \21261 , \12849 , \21260 );
or \U$20919 ( \21262 , \12848 , \21261 );
and \U$20920 ( \21263 , \12570 , \21262 );
or \U$20921 ( \21264 , \12569 , \21263 );
and \U$20922 ( \21265 , \12285 , \21264 );
or \U$20923 ( \21266 , \12284 , \21265 );
and \U$20924 ( \21267 , \11969 , \21266 );
or \U$20925 ( \21268 , \11968 , \21267 );
and \U$20926 ( \21269 , \11669 , \21268 );
or \U$20927 ( \21270 , \11668 , \21269 );
and \U$20928 ( \21271 , \11353 , \21270 );
or \U$20929 ( \21272 , \11352 , \21271 );
and \U$20930 ( \21273 , \11035 , \21272 );
or \U$20931 ( \21274 , \11034 , \21273 );
and \U$20932 ( \21275 , \10724 , \21274 );
or \U$20933 ( \21276 , \10723 , \21275 );
and \U$20934 ( \21277 , \10411 , \21276 );
or \U$20935 ( \21278 , \10410 , \21277 );
and \U$20936 ( \21279 , \10095 , \21278 );
or \U$20937 ( \21280 , \10094 , \21279 );
and \U$20938 ( \21281 , \9777 , \21280 );
or \U$20939 ( \21282 , \9776 , \21281 );
and \U$20940 ( \21283 , \9468 , \21282 );
or \U$20941 ( \21284 , \9467 , \21283 );
and \U$20942 ( \21285 , \9172 , \21284 );
or \U$20943 ( \21286 , \9171 , \21285 );
and \U$20944 ( \21287 , \8871 , \21286 );
or \U$20945 ( \21288 , \8870 , \21287 );
and \U$20946 ( \21289 , \8583 , \21288 );
or \U$20947 ( \21290 , \8582 , \21289 );
and \U$20948 ( \21291 , \8300 , \21290 );
or \U$20949 ( \21292 , \8299 , \21291 );
and \U$20950 ( \21293 , \8005 , \21292 );
or \U$20951 ( \21294 , \8004 , \21293 );
and \U$20952 ( \21295 , \7739 , \21294 );
or \U$20953 ( \21296 , \7738 , \21295 );
and \U$20954 ( \21297 , \7473 , \21296 );
or \U$20955 ( \21298 , \7472 , \21297 );
and \U$20956 ( \21299 , \7212 , \21298 );
or \U$20957 ( \21300 , \7211 , \21299 );
and \U$20958 ( \21301 , \6947 , \21300 );
or \U$20959 ( \21302 , \6946 , \21301 );
and \U$20960 ( \21303 , \6684 , \21302 );
or \U$20961 ( \21304 , \6683 , \21303 );
and \U$20962 ( \21305 , \6427 , \21304 );
or \U$20963 ( \21306 , \6426 , \21305 );
and \U$20964 ( \21307 , \6171 , \21306 );
or \U$20965 ( \21308 , \6170 , \21307 );
and \U$20966 ( \21309 , \5918 , \21308 );
or \U$20967 ( \21310 , \5917 , \21309 );
and \U$20968 ( \21311 , \5670 , \21310 );
or \U$20969 ( \21312 , \5669 , \21311 );
and \U$20970 ( \21313 , \5438 , \21312 );
or \U$20971 ( \21314 , \5437 , \21313 );
and \U$20972 ( \21315 , \5195 , \21314 );
or \U$20973 ( \21316 , \5194 , \21315 );
and \U$20974 ( \21317 , \4766 , \21316 );
or \U$20975 ( \21318 , \4765 , \21317 );
and \U$20976 ( \21319 , \4556 , \21318 );
or \U$20977 ( \21320 , \4555 , \21319 );
and \U$20978 ( \21321 , \4349 , \21320 );
or \U$20979 ( \21322 , \4348 , \21321 );
and \U$20980 ( \21323 , \4147 , \21322 );
or \U$20981 ( \21324 , \4146 , \21323 );
and \U$20982 ( \21325 , \3951 , \21324 );
or \U$20983 ( \21326 , \3950 , \21325 );
and \U$20984 ( \21327 , \3754 , \21326 );
or \U$20985 ( \21328 , \3753 , \21327 );
and \U$20986 ( \21329 , \3577 , \21328 );
or \U$20987 ( \21330 , \3576 , \21329 );
and \U$20988 ( \21331 , \3396 , \21330 );
or \U$20989 ( \21332 , \3395 , \21331 );
and \U$20990 ( \21333 , \3225 , \21332 );
or \U$20991 ( \21334 , \3224 , \21333 );
and \U$20992 ( \21335 , \3050 , \21334 );
or \U$20993 ( \21336 , \3049 , \21335 );
and \U$20994 ( \21337 , \2877 , \21336 );
or \U$20995 ( \21338 , \2876 , \21337 );
and \U$20996 ( \21339 , \2710 , \21338 );
or \U$20997 ( \21340 , \2709 , \21339 );
and \U$20998 ( \21341 , \2544 , \21340 );
or \U$20999 ( \21342 , \2543 , \21341 );
and \U$21000 ( \21343 , \2371 , \21342 );
or \U$21001 ( \21344 , \2370 , \21343 );
and \U$21002 ( \21345 , \2091 , \21344 );
or \U$21003 ( \21346 , \2090 , \21345 );
and \U$21004 ( \21347 , \1954 , \21346 );
or \U$21005 ( \21348 , \1953 , \21347 );
and \U$21006 ( \21349 , \1821 , \21348 );
or \U$21007 ( \21350 , \1820 , \21349 );
and \U$21008 ( \21351 , \1700 , \21350 );
or \U$21009 ( \21352 , \1699 , \21351 );
and \U$21010 ( \21353 , \1577 , \21352 );
or \U$21011 ( \21354 , \1576 , \21353 );
and \U$21012 ( \21355 , \1461 , \21354 );
or \U$21013 ( \21356 , \1460 , \21355 );
and \U$21014 ( \21357 , \1346 , \21356 );
or \U$21015 ( \21358 , \1345 , \21357 );
and \U$21016 ( \21359 , \1232 , \21358 );
or \U$21017 ( \21360 , \1231 , \21359 );
and \U$21018 ( \21361 , \1118 , \21360 );
or \U$21019 ( \21362 , \1117 , \21361 );
and \U$21020 ( \21363 , \936 , \21362 );
or \U$21021 ( \21364 , \935 , \21363 );
and \U$21022 ( \21365 , \857 , \21364 );
or \U$21023 ( \21366 , \856 , \21365 );
and \U$21024 ( \21367 , \774 , \21366 );
or \U$21025 ( \21368 , \773 , \21367 );
xor \U$21026 ( \21369 , \693 , \21368 );
buf gac4c_GF_PartitionCandidate( \21370_nGac4c , \21369 );
buf \U$21027 ( \21371 , \21370_nGac4c );
buf \U$21028 ( \21372 , RIbb2f070_13);
buf \U$21029 ( \21373 , RIbb2eff8_14);
buf \U$21030 ( \21374 , RIbb2ef80_15);
and \U$21031 ( \21375 , \21373 , \21374 );
not \U$21032 ( \21376 , \21375 );
and \U$21033 ( \21377 , \21372 , \21376 );
not \U$21034 ( \21378 , \21377 );
buf \U$21035 ( \21379 , RIbb31668_130);
buf \U$21036 ( \21380 , RIbb2f160_11);
buf \U$21037 ( \21381 , RIbb2f0e8_12);
xor \U$21038 ( \21382 , \21380 , \21381 );
xor \U$21039 ( \21383 , \21381 , \21372 );
not \U$21040 ( \21384 , \21383 );
and \U$21041 ( \21385 , \21382 , \21384 );
and \U$21042 ( \21386 , \21379 , \21385 );
buf \U$21043 ( \21387 , RIbb315f0_129);
and \U$21044 ( \21388 , \21387 , \21383 );
nor \U$21045 ( \21389 , \21386 , \21388 );
and \U$21046 ( \21390 , \21381 , \21372 );
not \U$21047 ( \21391 , \21390 );
and \U$21048 ( \21392 , \21380 , \21391 );
xnor \U$21049 ( \21393 , \21389 , \21392 );
and \U$21050 ( \21394 , \21378 , \21393 );
buf \U$21051 ( \21395 , RIbb31758_132);
buf \U$21052 ( \21396 , RIbb2f250_9);
buf \U$21053 ( \21397 , RIbb2f1d8_10);
xor \U$21054 ( \21398 , \21396 , \21397 );
xor \U$21055 ( \21399 , \21397 , \21380 );
not \U$21056 ( \21400 , \21399 );
and \U$21057 ( \21401 , \21398 , \21400 );
and \U$21058 ( \21402 , \21395 , \21401 );
buf \U$21059 ( \21403 , RIbb316e0_131);
and \U$21060 ( \21404 , \21403 , \21399 );
nor \U$21061 ( \21405 , \21402 , \21404 );
and \U$21062 ( \21406 , \21397 , \21380 );
not \U$21063 ( \21407 , \21406 );
and \U$21064 ( \21408 , \21396 , \21407 );
xnor \U$21065 ( \21409 , \21405 , \21408 );
and \U$21066 ( \21410 , \21393 , \21409 );
and \U$21067 ( \21411 , \21378 , \21409 );
or \U$21068 ( \21412 , \21394 , \21410 , \21411 );
buf \U$21069 ( \21413 , RIbb31848_134);
buf \U$21070 ( \21414 , RIbb2f340_7);
buf \U$21071 ( \21415 , RIbb2f2c8_8);
xor \U$21072 ( \21416 , \21414 , \21415 );
xor \U$21073 ( \21417 , \21415 , \21396 );
not \U$21074 ( \21418 , \21417 );
and \U$21075 ( \21419 , \21416 , \21418 );
and \U$21076 ( \21420 , \21413 , \21419 );
buf \U$21077 ( \21421 , RIbb317d0_133);
and \U$21078 ( \21422 , \21421 , \21417 );
nor \U$21079 ( \21423 , \21420 , \21422 );
and \U$21080 ( \21424 , \21415 , \21396 );
not \U$21081 ( \21425 , \21424 );
and \U$21082 ( \21426 , \21414 , \21425 );
xnor \U$21083 ( \21427 , \21423 , \21426 );
buf \U$21084 ( \21428 , RIbb31938_136);
buf \U$21085 ( \21429 , RIbb2f430_5);
buf \U$21086 ( \21430 , RIbb2f3b8_6);
xor \U$21087 ( \21431 , \21429 , \21430 );
xor \U$21088 ( \21432 , \21430 , \21414 );
not \U$21089 ( \21433 , \21432 );
and \U$21090 ( \21434 , \21431 , \21433 );
and \U$21091 ( \21435 , \21428 , \21434 );
buf \U$21092 ( \21436 , RIbb318c0_135);
and \U$21093 ( \21437 , \21436 , \21432 );
nor \U$21094 ( \21438 , \21435 , \21437 );
and \U$21095 ( \21439 , \21430 , \21414 );
not \U$21096 ( \21440 , \21439 );
and \U$21097 ( \21441 , \21429 , \21440 );
xnor \U$21098 ( \21442 , \21438 , \21441 );
and \U$21099 ( \21443 , \21427 , \21442 );
buf \U$21100 ( \21444 , RIbb31a28_138);
buf \U$21101 ( \21445 , RIbb2f520_3);
buf \U$21102 ( \21446 , RIbb2f4a8_4);
xor \U$21103 ( \21447 , \21445 , \21446 );
xor \U$21104 ( \21448 , \21446 , \21429 );
not \U$21105 ( \21449 , \21448 );
and \U$21106 ( \21450 , \21447 , \21449 );
and \U$21107 ( \21451 , \21444 , \21450 );
buf \U$21108 ( \21452 , RIbb319b0_137);
and \U$21109 ( \21453 , \21452 , \21448 );
nor \U$21110 ( \21454 , \21451 , \21453 );
and \U$21111 ( \21455 , \21446 , \21429 );
not \U$21112 ( \21456 , \21455 );
and \U$21113 ( \21457 , \21445 , \21456 );
xnor \U$21114 ( \21458 , \21454 , \21457 );
and \U$21115 ( \21459 , \21442 , \21458 );
and \U$21116 ( \21460 , \21427 , \21458 );
or \U$21117 ( \21461 , \21443 , \21459 , \21460 );
and \U$21118 ( \21462 , \21412 , \21461 );
buf \U$21119 ( \21463 , RIbb31b18_140);
buf \U$21120 ( \21464 , RIbb2f610_1);
buf \U$21121 ( \21465 , RIbb2f598_2);
xor \U$21122 ( \21466 , \21464 , \21465 );
xor \U$21123 ( \21467 , \21465 , \21445 );
not \U$21124 ( \21468 , \21467 );
and \U$21125 ( \21469 , \21466 , \21468 );
and \U$21126 ( \21470 , \21463 , \21469 );
buf \U$21127 ( \21471 , RIbb31aa0_139);
and \U$21128 ( \21472 , \21471 , \21467 );
nor \U$21129 ( \21473 , \21470 , \21472 );
and \U$21130 ( \21474 , \21465 , \21445 );
not \U$21131 ( \21475 , \21474 );
and \U$21132 ( \21476 , \21464 , \21475 );
xnor \U$21133 ( \21477 , \21473 , \21476 );
buf \U$21134 ( \21478 , RIbb31b90_141);
and \U$21135 ( \21479 , \21478 , \21464 );
and \U$21136 ( \21480 , \21477 , \21479 );
and \U$21137 ( \21481 , \21461 , \21480 );
and \U$21138 ( \21482 , \21412 , \21480 );
or \U$21139 ( \21483 , \21462 , \21481 , \21482 );
and \U$21140 ( \21484 , \21436 , \21434 );
and \U$21141 ( \21485 , \21413 , \21432 );
nor \U$21142 ( \21486 , \21484 , \21485 );
xnor \U$21143 ( \21487 , \21486 , \21441 );
and \U$21144 ( \21488 , \21452 , \21450 );
and \U$21145 ( \21489 , \21428 , \21448 );
nor \U$21146 ( \21490 , \21488 , \21489 );
xnor \U$21147 ( \21491 , \21490 , \21457 );
xor \U$21148 ( \21492 , \21487 , \21491 );
and \U$21149 ( \21493 , \21471 , \21469 );
and \U$21150 ( \21494 , \21444 , \21467 );
nor \U$21151 ( \21495 , \21493 , \21494 );
xnor \U$21152 ( \21496 , \21495 , \21476 );
xor \U$21153 ( \21497 , \21492 , \21496 );
and \U$21154 ( \21498 , \21387 , \21385 );
not \U$21155 ( \21499 , \21498 );
xnor \U$21156 ( \21500 , \21499 , \21392 );
and \U$21157 ( \21501 , \21403 , \21401 );
and \U$21158 ( \21502 , \21379 , \21399 );
nor \U$21159 ( \21503 , \21501 , \21502 );
xnor \U$21160 ( \21504 , \21503 , \21408 );
xor \U$21161 ( \21505 , \21500 , \21504 );
and \U$21162 ( \21506 , \21421 , \21419 );
and \U$21163 ( \21507 , \21395 , \21417 );
nor \U$21164 ( \21508 , \21506 , \21507 );
xnor \U$21165 ( \21509 , \21508 , \21426 );
xor \U$21166 ( \21510 , \21505 , \21509 );
and \U$21167 ( \21511 , \21497 , \21510 );
and \U$21168 ( \21512 , \21463 , \21464 );
not \U$21169 ( \21513 , \21512 );
and \U$21170 ( \21514 , \21510 , \21513 );
and \U$21171 ( \21515 , \21497 , \21513 );
or \U$21172 ( \21516 , \21511 , \21514 , \21515 );
and \U$21173 ( \21517 , \21483 , \21516 );
and \U$21174 ( \21518 , \21471 , \21464 );
and \U$21175 ( \21519 , \21413 , \21434 );
and \U$21176 ( \21520 , \21421 , \21432 );
nor \U$21177 ( \21521 , \21519 , \21520 );
xnor \U$21178 ( \21522 , \21521 , \21441 );
and \U$21179 ( \21523 , \21428 , \21450 );
and \U$21180 ( \21524 , \21436 , \21448 );
nor \U$21181 ( \21525 , \21523 , \21524 );
xnor \U$21182 ( \21526 , \21525 , \21457 );
xor \U$21183 ( \21527 , \21522 , \21526 );
and \U$21184 ( \21528 , \21444 , \21469 );
and \U$21185 ( \21529 , \21452 , \21467 );
nor \U$21186 ( \21530 , \21528 , \21529 );
xnor \U$21187 ( \21531 , \21530 , \21476 );
xor \U$21188 ( \21532 , \21527 , \21531 );
xor \U$21189 ( \21533 , \21518 , \21532 );
not \U$21190 ( \21534 , \21392 );
and \U$21191 ( \21535 , \21379 , \21401 );
and \U$21192 ( \21536 , \21387 , \21399 );
nor \U$21193 ( \21537 , \21535 , \21536 );
xnor \U$21194 ( \21538 , \21537 , \21408 );
xor \U$21195 ( \21539 , \21534 , \21538 );
and \U$21196 ( \21540 , \21395 , \21419 );
and \U$21197 ( \21541 , \21403 , \21417 );
nor \U$21198 ( \21542 , \21540 , \21541 );
xnor \U$21199 ( \21543 , \21542 , \21426 );
xor \U$21200 ( \21544 , \21539 , \21543 );
xor \U$21201 ( \21545 , \21533 , \21544 );
and \U$21202 ( \21546 , \21516 , \21545 );
and \U$21203 ( \21547 , \21483 , \21545 );
or \U$21204 ( \21548 , \21517 , \21546 , \21547 );
and \U$21205 ( \21549 , \21487 , \21491 );
and \U$21206 ( \21550 , \21491 , \21496 );
and \U$21207 ( \21551 , \21487 , \21496 );
or \U$21208 ( \21552 , \21549 , \21550 , \21551 );
and \U$21209 ( \21553 , \21500 , \21504 );
and \U$21210 ( \21554 , \21504 , \21509 );
and \U$21211 ( \21555 , \21500 , \21509 );
or \U$21212 ( \21556 , \21553 , \21554 , \21555 );
and \U$21213 ( \21557 , \21552 , \21556 );
buf \U$21214 ( \21558 , \21512 );
and \U$21215 ( \21559 , \21556 , \21558 );
and \U$21216 ( \21560 , \21552 , \21558 );
or \U$21217 ( \21561 , \21557 , \21559 , \21560 );
and \U$21218 ( \21562 , \21518 , \21532 );
and \U$21219 ( \21563 , \21532 , \21544 );
and \U$21220 ( \21564 , \21518 , \21544 );
or \U$21221 ( \21565 , \21562 , \21563 , \21564 );
xor \U$21222 ( \21566 , \21561 , \21565 );
and \U$21223 ( \21567 , \21436 , \21450 );
and \U$21224 ( \21568 , \21413 , \21448 );
nor \U$21225 ( \21569 , \21567 , \21568 );
xnor \U$21226 ( \21570 , \21569 , \21457 );
and \U$21227 ( \21571 , \21452 , \21469 );
and \U$21228 ( \21572 , \21428 , \21467 );
nor \U$21229 ( \21573 , \21571 , \21572 );
xnor \U$21230 ( \21574 , \21573 , \21476 );
xor \U$21231 ( \21575 , \21570 , \21574 );
and \U$21232 ( \21576 , \21444 , \21464 );
xor \U$21233 ( \21577 , \21575 , \21576 );
xor \U$21234 ( \21578 , \21566 , \21577 );
and \U$21235 ( \21579 , \21548 , \21578 );
and \U$21236 ( \21580 , \21387 , \21401 );
not \U$21237 ( \21581 , \21580 );
xnor \U$21238 ( \21582 , \21581 , \21408 );
and \U$21239 ( \21583 , \21403 , \21419 );
and \U$21240 ( \21584 , \21379 , \21417 );
nor \U$21241 ( \21585 , \21583 , \21584 );
xnor \U$21242 ( \21586 , \21585 , \21426 );
xor \U$21243 ( \21587 , \21582 , \21586 );
and \U$21244 ( \21588 , \21421 , \21434 );
and \U$21245 ( \21589 , \21395 , \21432 );
nor \U$21246 ( \21590 , \21588 , \21589 );
xnor \U$21247 ( \21591 , \21590 , \21441 );
xor \U$21248 ( \21592 , \21587 , \21591 );
and \U$21249 ( \21593 , \21522 , \21526 );
and \U$21250 ( \21594 , \21526 , \21531 );
and \U$21251 ( \21595 , \21522 , \21531 );
or \U$21252 ( \21596 , \21593 , \21594 , \21595 );
and \U$21253 ( \21597 , \21534 , \21538 );
and \U$21254 ( \21598 , \21538 , \21543 );
and \U$21255 ( \21599 , \21534 , \21543 );
or \U$21256 ( \21600 , \21597 , \21598 , \21599 );
xnor \U$21257 ( \21601 , \21596 , \21600 );
xor \U$21258 ( \21602 , \21592 , \21601 );
and \U$21259 ( \21603 , \21578 , \21602 );
and \U$21260 ( \21604 , \21548 , \21602 );
or \U$21261 ( \21605 , \21579 , \21603 , \21604 );
and \U$21262 ( \21606 , \21561 , \21565 );
and \U$21263 ( \21607 , \21565 , \21577 );
and \U$21264 ( \21608 , \21561 , \21577 );
or \U$21265 ( \21609 , \21606 , \21607 , \21608 );
and \U$21266 ( \21610 , \21592 , \21601 );
xor \U$21267 ( \21611 , \21609 , \21610 );
or \U$21268 ( \21612 , \21596 , \21600 );
not \U$21269 ( \21613 , \21408 );
and \U$21270 ( \21614 , \21379 , \21419 );
and \U$21271 ( \21615 , \21387 , \21417 );
nor \U$21272 ( \21616 , \21614 , \21615 );
xnor \U$21273 ( \21617 , \21616 , \21426 );
xor \U$21274 ( \21618 , \21613 , \21617 );
and \U$21275 ( \21619 , \21395 , \21434 );
and \U$21276 ( \21620 , \21403 , \21432 );
nor \U$21277 ( \21621 , \21619 , \21620 );
xnor \U$21278 ( \21622 , \21621 , \21441 );
xor \U$21279 ( \21623 , \21618 , \21622 );
xor \U$21280 ( \21624 , \21612 , \21623 );
and \U$21281 ( \21625 , \21582 , \21586 );
and \U$21282 ( \21626 , \21586 , \21591 );
and \U$21283 ( \21627 , \21582 , \21591 );
or \U$21284 ( \21628 , \21625 , \21626 , \21627 );
and \U$21285 ( \21629 , \21570 , \21574 );
and \U$21286 ( \21630 , \21574 , \21576 );
and \U$21287 ( \21631 , \21570 , \21576 );
or \U$21288 ( \21632 , \21629 , \21630 , \21631 );
xor \U$21289 ( \21633 , \21628 , \21632 );
and \U$21290 ( \21634 , \21413 , \21450 );
and \U$21291 ( \21635 , \21421 , \21448 );
nor \U$21292 ( \21636 , \21634 , \21635 );
xnor \U$21293 ( \21637 , \21636 , \21457 );
and \U$21294 ( \21638 , \21428 , \21469 );
and \U$21295 ( \21639 , \21436 , \21467 );
nor \U$21296 ( \21640 , \21638 , \21639 );
xnor \U$21297 ( \21641 , \21640 , \21476 );
xor \U$21298 ( \21642 , \21637 , \21641 );
and \U$21299 ( \21643 , \21452 , \21464 );
xor \U$21300 ( \21644 , \21642 , \21643 );
xor \U$21301 ( \21645 , \21633 , \21644 );
xor \U$21302 ( \21646 , \21624 , \21645 );
xor \U$21303 ( \21647 , \21611 , \21646 );
xor \U$21304 ( \21648 , \21605 , \21647 );
xor \U$21305 ( \21649 , \21372 , \21373 );
xor \U$21306 ( \21650 , \21373 , \21374 );
not \U$21307 ( \21651 , \21650 );
and \U$21308 ( \21652 , \21649 , \21651 );
and \U$21309 ( \21653 , \21387 , \21652 );
not \U$21310 ( \21654 , \21653 );
xnor \U$21311 ( \21655 , \21654 , \21377 );
and \U$21312 ( \21656 , \21403 , \21385 );
and \U$21313 ( \21657 , \21379 , \21383 );
nor \U$21314 ( \21658 , \21656 , \21657 );
xnor \U$21315 ( \21659 , \21658 , \21392 );
and \U$21316 ( \21660 , \21655 , \21659 );
and \U$21317 ( \21661 , \21421 , \21401 );
and \U$21318 ( \21662 , \21395 , \21399 );
nor \U$21319 ( \21663 , \21661 , \21662 );
xnor \U$21320 ( \21664 , \21663 , \21408 );
and \U$21321 ( \21665 , \21659 , \21664 );
and \U$21322 ( \21666 , \21655 , \21664 );
or \U$21323 ( \21667 , \21660 , \21665 , \21666 );
and \U$21324 ( \21668 , \21436 , \21419 );
and \U$21325 ( \21669 , \21413 , \21417 );
nor \U$21326 ( \21670 , \21668 , \21669 );
xnor \U$21327 ( \21671 , \21670 , \21426 );
and \U$21328 ( \21672 , \21452 , \21434 );
and \U$21329 ( \21673 , \21428 , \21432 );
nor \U$21330 ( \21674 , \21672 , \21673 );
xnor \U$21331 ( \21675 , \21674 , \21441 );
and \U$21332 ( \21676 , \21671 , \21675 );
and \U$21333 ( \21677 , \21471 , \21450 );
and \U$21334 ( \21678 , \21444 , \21448 );
nor \U$21335 ( \21679 , \21677 , \21678 );
xnor \U$21336 ( \21680 , \21679 , \21457 );
and \U$21337 ( \21681 , \21675 , \21680 );
and \U$21338 ( \21682 , \21671 , \21680 );
or \U$21339 ( \21683 , \21676 , \21681 , \21682 );
and \U$21340 ( \21684 , \21667 , \21683 );
and \U$21341 ( \21685 , \21478 , \21469 );
and \U$21342 ( \21686 , \21463 , \21467 );
nor \U$21343 ( \21687 , \21685 , \21686 );
xnor \U$21344 ( \21688 , \21687 , \21476 );
buf \U$21345 ( \21689 , RIbb31c08_142);
and \U$21346 ( \21690 , \21689 , \21464 );
or \U$21347 ( \21691 , \21688 , \21690 );
and \U$21348 ( \21692 , \21683 , \21691 );
and \U$21349 ( \21693 , \21667 , \21691 );
or \U$21350 ( \21694 , \21684 , \21692 , \21693 );
xor \U$21351 ( \21695 , \21378 , \21393 );
xor \U$21352 ( \21696 , \21695 , \21409 );
xor \U$21353 ( \21697 , \21427 , \21442 );
xor \U$21354 ( \21698 , \21697 , \21458 );
and \U$21355 ( \21699 , \21696 , \21698 );
xor \U$21356 ( \21700 , \21477 , \21479 );
and \U$21357 ( \21701 , \21698 , \21700 );
and \U$21358 ( \21702 , \21696 , \21700 );
or \U$21359 ( \21703 , \21699 , \21701 , \21702 );
and \U$21360 ( \21704 , \21694 , \21703 );
xor \U$21361 ( \21705 , \21497 , \21510 );
xor \U$21362 ( \21706 , \21705 , \21513 );
and \U$21363 ( \21707 , \21703 , \21706 );
and \U$21364 ( \21708 , \21694 , \21706 );
or \U$21365 ( \21709 , \21704 , \21707 , \21708 );
xor \U$21366 ( \21710 , \21552 , \21556 );
xor \U$21367 ( \21711 , \21710 , \21558 );
and \U$21368 ( \21712 , \21709 , \21711 );
xor \U$21369 ( \21713 , \21483 , \21516 );
xor \U$21370 ( \21714 , \21713 , \21545 );
and \U$21371 ( \21715 , \21711 , \21714 );
and \U$21372 ( \21716 , \21709 , \21714 );
or \U$21373 ( \21717 , \21712 , \21715 , \21716 );
xor \U$21374 ( \21718 , \21548 , \21578 );
xor \U$21375 ( \21719 , \21718 , \21602 );
and \U$21376 ( \21720 , \21717 , \21719 );
xor \U$21377 ( \21721 , \21648 , \21720 );
xor \U$21378 ( \21722 , \21717 , \21719 );
buf \U$21379 ( \21723 , RIbb2ef08_16);
buf \U$21380 ( \21724 , RIbb2ee90_17);
and \U$21381 ( \21725 , \21723 , \21724 );
not \U$21382 ( \21726 , \21725 );
and \U$21383 ( \21727 , \21374 , \21726 );
not \U$21384 ( \21728 , \21727 );
and \U$21385 ( \21729 , \21379 , \21652 );
and \U$21386 ( \21730 , \21387 , \21650 );
nor \U$21387 ( \21731 , \21729 , \21730 );
xnor \U$21388 ( \21732 , \21731 , \21377 );
and \U$21389 ( \21733 , \21728 , \21732 );
and \U$21390 ( \21734 , \21395 , \21385 );
and \U$21391 ( \21735 , \21403 , \21383 );
nor \U$21392 ( \21736 , \21734 , \21735 );
xnor \U$21393 ( \21737 , \21736 , \21392 );
and \U$21394 ( \21738 , \21732 , \21737 );
and \U$21395 ( \21739 , \21728 , \21737 );
or \U$21396 ( \21740 , \21733 , \21738 , \21739 );
and \U$21397 ( \21741 , \21463 , \21450 );
and \U$21398 ( \21742 , \21471 , \21448 );
nor \U$21399 ( \21743 , \21741 , \21742 );
xnor \U$21400 ( \21744 , \21743 , \21457 );
and \U$21401 ( \21745 , \21689 , \21469 );
and \U$21402 ( \21746 , \21478 , \21467 );
nor \U$21403 ( \21747 , \21745 , \21746 );
xnor \U$21404 ( \21748 , \21747 , \21476 );
and \U$21405 ( \21749 , \21744 , \21748 );
buf \U$21406 ( \21750 , RIbb31c80_143);
and \U$21407 ( \21751 , \21750 , \21464 );
and \U$21408 ( \21752 , \21748 , \21751 );
and \U$21409 ( \21753 , \21744 , \21751 );
or \U$21410 ( \21754 , \21749 , \21752 , \21753 );
and \U$21411 ( \21755 , \21740 , \21754 );
and \U$21412 ( \21756 , \21413 , \21401 );
and \U$21413 ( \21757 , \21421 , \21399 );
nor \U$21414 ( \21758 , \21756 , \21757 );
xnor \U$21415 ( \21759 , \21758 , \21408 );
and \U$21416 ( \21760 , \21428 , \21419 );
and \U$21417 ( \21761 , \21436 , \21417 );
nor \U$21418 ( \21762 , \21760 , \21761 );
xnor \U$21419 ( \21763 , \21762 , \21426 );
and \U$21420 ( \21764 , \21759 , \21763 );
and \U$21421 ( \21765 , \21444 , \21434 );
and \U$21422 ( \21766 , \21452 , \21432 );
nor \U$21423 ( \21767 , \21765 , \21766 );
xnor \U$21424 ( \21768 , \21767 , \21441 );
and \U$21425 ( \21769 , \21763 , \21768 );
and \U$21426 ( \21770 , \21759 , \21768 );
or \U$21427 ( \21771 , \21764 , \21769 , \21770 );
and \U$21428 ( \21772 , \21754 , \21771 );
and \U$21429 ( \21773 , \21740 , \21771 );
or \U$21430 ( \21774 , \21755 , \21772 , \21773 );
xor \U$21431 ( \21775 , \21655 , \21659 );
xor \U$21432 ( \21776 , \21775 , \21664 );
xor \U$21433 ( \21777 , \21671 , \21675 );
xor \U$21434 ( \21778 , \21777 , \21680 );
and \U$21435 ( \21779 , \21776 , \21778 );
xnor \U$21436 ( \21780 , \21688 , \21690 );
and \U$21437 ( \21781 , \21778 , \21780 );
and \U$21438 ( \21782 , \21776 , \21780 );
or \U$21439 ( \21783 , \21779 , \21781 , \21782 );
and \U$21440 ( \21784 , \21774 , \21783 );
xor \U$21441 ( \21785 , \21696 , \21698 );
xor \U$21442 ( \21786 , \21785 , \21700 );
and \U$21443 ( \21787 , \21783 , \21786 );
and \U$21444 ( \21788 , \21774 , \21786 );
or \U$21445 ( \21789 , \21784 , \21787 , \21788 );
xor \U$21446 ( \21790 , \21412 , \21461 );
xor \U$21447 ( \21791 , \21790 , \21480 );
and \U$21448 ( \21792 , \21789 , \21791 );
xor \U$21449 ( \21793 , \21694 , \21703 );
xor \U$21450 ( \21794 , \21793 , \21706 );
and \U$21451 ( \21795 , \21791 , \21794 );
and \U$21452 ( \21796 , \21789 , \21794 );
or \U$21453 ( \21797 , \21792 , \21795 , \21796 );
xor \U$21454 ( \21798 , \21709 , \21711 );
xor \U$21455 ( \21799 , \21798 , \21714 );
and \U$21456 ( \21800 , \21797 , \21799 );
and \U$21457 ( \21801 , \21722 , \21800 );
xor \U$21458 ( \21802 , \21722 , \21800 );
xor \U$21459 ( \21803 , \21797 , \21799 );
and \U$21460 ( \21804 , \21478 , \21450 );
and \U$21461 ( \21805 , \21463 , \21448 );
nor \U$21462 ( \21806 , \21804 , \21805 );
xnor \U$21463 ( \21807 , \21806 , \21457 );
and \U$21464 ( \21808 , \21750 , \21469 );
and \U$21465 ( \21809 , \21689 , \21467 );
nor \U$21466 ( \21810 , \21808 , \21809 );
xnor \U$21467 ( \21811 , \21810 , \21476 );
and \U$21468 ( \21812 , \21807 , \21811 );
buf \U$21469 ( \21813 , RIbb31cf8_144);
and \U$21470 ( \21814 , \21813 , \21464 );
and \U$21471 ( \21815 , \21811 , \21814 );
and \U$21472 ( \21816 , \21807 , \21814 );
or \U$21473 ( \21817 , \21812 , \21815 , \21816 );
xor \U$21474 ( \21818 , \21374 , \21723 );
xor \U$21475 ( \21819 , \21723 , \21724 );
not \U$21476 ( \21820 , \21819 );
and \U$21477 ( \21821 , \21818 , \21820 );
and \U$21478 ( \21822 , \21387 , \21821 );
not \U$21479 ( \21823 , \21822 );
xnor \U$21480 ( \21824 , \21823 , \21727 );
and \U$21481 ( \21825 , \21403 , \21652 );
and \U$21482 ( \21826 , \21379 , \21650 );
nor \U$21483 ( \21827 , \21825 , \21826 );
xnor \U$21484 ( \21828 , \21827 , \21377 );
and \U$21485 ( \21829 , \21824 , \21828 );
and \U$21486 ( \21830 , \21421 , \21385 );
and \U$21487 ( \21831 , \21395 , \21383 );
nor \U$21488 ( \21832 , \21830 , \21831 );
xnor \U$21489 ( \21833 , \21832 , \21392 );
and \U$21490 ( \21834 , \21828 , \21833 );
and \U$21491 ( \21835 , \21824 , \21833 );
or \U$21492 ( \21836 , \21829 , \21834 , \21835 );
and \U$21493 ( \21837 , \21817 , \21836 );
and \U$21494 ( \21838 , \21436 , \21401 );
and \U$21495 ( \21839 , \21413 , \21399 );
nor \U$21496 ( \21840 , \21838 , \21839 );
xnor \U$21497 ( \21841 , \21840 , \21408 );
and \U$21498 ( \21842 , \21452 , \21419 );
and \U$21499 ( \21843 , \21428 , \21417 );
nor \U$21500 ( \21844 , \21842 , \21843 );
xnor \U$21501 ( \21845 , \21844 , \21426 );
and \U$21502 ( \21846 , \21841 , \21845 );
and \U$21503 ( \21847 , \21471 , \21434 );
and \U$21504 ( \21848 , \21444 , \21432 );
nor \U$21505 ( \21849 , \21847 , \21848 );
xnor \U$21506 ( \21850 , \21849 , \21441 );
and \U$21507 ( \21851 , \21845 , \21850 );
and \U$21508 ( \21852 , \21841 , \21850 );
or \U$21509 ( \21853 , \21846 , \21851 , \21852 );
and \U$21510 ( \21854 , \21836 , \21853 );
and \U$21511 ( \21855 , \21817 , \21853 );
or \U$21512 ( \21856 , \21837 , \21854 , \21855 );
xor \U$21513 ( \21857 , \21728 , \21732 );
xor \U$21514 ( \21858 , \21857 , \21737 );
xor \U$21515 ( \21859 , \21744 , \21748 );
xor \U$21516 ( \21860 , \21859 , \21751 );
and \U$21517 ( \21861 , \21858 , \21860 );
xor \U$21518 ( \21862 , \21759 , \21763 );
xor \U$21519 ( \21863 , \21862 , \21768 );
and \U$21520 ( \21864 , \21860 , \21863 );
and \U$21521 ( \21865 , \21858 , \21863 );
or \U$21522 ( \21866 , \21861 , \21864 , \21865 );
and \U$21523 ( \21867 , \21856 , \21866 );
xor \U$21524 ( \21868 , \21776 , \21778 );
xor \U$21525 ( \21869 , \21868 , \21780 );
and \U$21526 ( \21870 , \21866 , \21869 );
and \U$21527 ( \21871 , \21856 , \21869 );
or \U$21528 ( \21872 , \21867 , \21870 , \21871 );
xor \U$21529 ( \21873 , \21667 , \21683 );
xor \U$21530 ( \21874 , \21873 , \21691 );
and \U$21531 ( \21875 , \21872 , \21874 );
xor \U$21532 ( \21876 , \21774 , \21783 );
xor \U$21533 ( \21877 , \21876 , \21786 );
and \U$21534 ( \21878 , \21874 , \21877 );
and \U$21535 ( \21879 , \21872 , \21877 );
or \U$21536 ( \21880 , \21875 , \21878 , \21879 );
xor \U$21537 ( \21881 , \21789 , \21791 );
xor \U$21538 ( \21882 , \21881 , \21794 );
and \U$21539 ( \21883 , \21880 , \21882 );
and \U$21540 ( \21884 , \21803 , \21883 );
xor \U$21541 ( \21885 , \21803 , \21883 );
xor \U$21542 ( \21886 , \21880 , \21882 );
and \U$21543 ( \21887 , \21413 , \21385 );
and \U$21544 ( \21888 , \21421 , \21383 );
nor \U$21545 ( \21889 , \21887 , \21888 );
xnor \U$21546 ( \21890 , \21889 , \21392 );
and \U$21547 ( \21891 , \21428 , \21401 );
and \U$21548 ( \21892 , \21436 , \21399 );
nor \U$21549 ( \21893 , \21891 , \21892 );
xnor \U$21550 ( \21894 , \21893 , \21408 );
and \U$21551 ( \21895 , \21890 , \21894 );
and \U$21552 ( \21896 , \21444 , \21419 );
and \U$21553 ( \21897 , \21452 , \21417 );
nor \U$21554 ( \21898 , \21896 , \21897 );
xnor \U$21555 ( \21899 , \21898 , \21426 );
and \U$21556 ( \21900 , \21894 , \21899 );
and \U$21557 ( \21901 , \21890 , \21899 );
or \U$21558 ( \21902 , \21895 , \21900 , \21901 );
buf \U$21559 ( \21903 , RIbb2ee18_18);
buf \U$21560 ( \21904 , RIbb2eda0_19);
and \U$21561 ( \21905 , \21903 , \21904 );
not \U$21562 ( \21906 , \21905 );
and \U$21563 ( \21907 , \21724 , \21906 );
not \U$21564 ( \21908 , \21907 );
and \U$21565 ( \21909 , \21379 , \21821 );
and \U$21566 ( \21910 , \21387 , \21819 );
nor \U$21567 ( \21911 , \21909 , \21910 );
xnor \U$21568 ( \21912 , \21911 , \21727 );
and \U$21569 ( \21913 , \21908 , \21912 );
and \U$21570 ( \21914 , \21395 , \21652 );
and \U$21571 ( \21915 , \21403 , \21650 );
nor \U$21572 ( \21916 , \21914 , \21915 );
xnor \U$21573 ( \21917 , \21916 , \21377 );
and \U$21574 ( \21918 , \21912 , \21917 );
and \U$21575 ( \21919 , \21908 , \21917 );
or \U$21576 ( \21920 , \21913 , \21918 , \21919 );
and \U$21577 ( \21921 , \21902 , \21920 );
and \U$21578 ( \21922 , \21463 , \21434 );
and \U$21579 ( \21923 , \21471 , \21432 );
nor \U$21580 ( \21924 , \21922 , \21923 );
xnor \U$21581 ( \21925 , \21924 , \21441 );
and \U$21582 ( \21926 , \21689 , \21450 );
and \U$21583 ( \21927 , \21478 , \21448 );
nor \U$21584 ( \21928 , \21926 , \21927 );
xnor \U$21585 ( \21929 , \21928 , \21457 );
and \U$21586 ( \21930 , \21925 , \21929 );
and \U$21587 ( \21931 , \21813 , \21469 );
and \U$21588 ( \21932 , \21750 , \21467 );
nor \U$21589 ( \21933 , \21931 , \21932 );
xnor \U$21590 ( \21934 , \21933 , \21476 );
and \U$21591 ( \21935 , \21929 , \21934 );
and \U$21592 ( \21936 , \21925 , \21934 );
or \U$21593 ( \21937 , \21930 , \21935 , \21936 );
and \U$21594 ( \21938 , \21920 , \21937 );
and \U$21595 ( \21939 , \21902 , \21937 );
or \U$21596 ( \21940 , \21921 , \21938 , \21939 );
xor \U$21597 ( \21941 , \21807 , \21811 );
xor \U$21598 ( \21942 , \21941 , \21814 );
xor \U$21599 ( \21943 , \21841 , \21845 );
xor \U$21600 ( \21944 , \21943 , \21850 );
or \U$21601 ( \21945 , \21942 , \21944 );
and \U$21602 ( \21946 , \21940 , \21945 );
xor \U$21603 ( \21947 , \21858 , \21860 );
xor \U$21604 ( \21948 , \21947 , \21863 );
and \U$21605 ( \21949 , \21945 , \21948 );
and \U$21606 ( \21950 , \21940 , \21948 );
or \U$21607 ( \21951 , \21946 , \21949 , \21950 );
xor \U$21608 ( \21952 , \21740 , \21754 );
xor \U$21609 ( \21953 , \21952 , \21771 );
and \U$21610 ( \21954 , \21951 , \21953 );
xor \U$21611 ( \21955 , \21856 , \21866 );
xor \U$21612 ( \21956 , \21955 , \21869 );
and \U$21613 ( \21957 , \21953 , \21956 );
and \U$21614 ( \21958 , \21951 , \21956 );
or \U$21615 ( \21959 , \21954 , \21957 , \21958 );
xor \U$21616 ( \21960 , \21872 , \21874 );
xor \U$21617 ( \21961 , \21960 , \21877 );
and \U$21618 ( \21962 , \21959 , \21961 );
and \U$21619 ( \21963 , \21886 , \21962 );
xor \U$21620 ( \21964 , \21886 , \21962 );
xor \U$21621 ( \21965 , \21959 , \21961 );
and \U$21622 ( \21966 , \21436 , \21385 );
and \U$21623 ( \21967 , \21413 , \21383 );
nor \U$21624 ( \21968 , \21966 , \21967 );
xnor \U$21625 ( \21969 , \21968 , \21392 );
and \U$21626 ( \21970 , \21452 , \21401 );
and \U$21627 ( \21971 , \21428 , \21399 );
nor \U$21628 ( \21972 , \21970 , \21971 );
xnor \U$21629 ( \21973 , \21972 , \21408 );
and \U$21630 ( \21974 , \21969 , \21973 );
and \U$21631 ( \21975 , \21471 , \21419 );
and \U$21632 ( \21976 , \21444 , \21417 );
nor \U$21633 ( \21977 , \21975 , \21976 );
xnor \U$21634 ( \21978 , \21977 , \21426 );
and \U$21635 ( \21979 , \21973 , \21978 );
and \U$21636 ( \21980 , \21969 , \21978 );
or \U$21637 ( \21981 , \21974 , \21979 , \21980 );
xor \U$21638 ( \21982 , \21724 , \21903 );
xor \U$21639 ( \21983 , \21903 , \21904 );
not \U$21640 ( \21984 , \21983 );
and \U$21641 ( \21985 , \21982 , \21984 );
and \U$21642 ( \21986 , \21387 , \21985 );
not \U$21643 ( \21987 , \21986 );
xnor \U$21644 ( \21988 , \21987 , \21907 );
and \U$21645 ( \21989 , \21403 , \21821 );
and \U$21646 ( \21990 , \21379 , \21819 );
nor \U$21647 ( \21991 , \21989 , \21990 );
xnor \U$21648 ( \21992 , \21991 , \21727 );
and \U$21649 ( \21993 , \21988 , \21992 );
and \U$21650 ( \21994 , \21421 , \21652 );
and \U$21651 ( \21995 , \21395 , \21650 );
nor \U$21652 ( \21996 , \21994 , \21995 );
xnor \U$21653 ( \21997 , \21996 , \21377 );
and \U$21654 ( \21998 , \21992 , \21997 );
and \U$21655 ( \21999 , \21988 , \21997 );
or \U$21656 ( \22000 , \21993 , \21998 , \21999 );
and \U$21657 ( \22001 , \21981 , \22000 );
and \U$21658 ( \22002 , \21478 , \21434 );
and \U$21659 ( \22003 , \21463 , \21432 );
nor \U$21660 ( \22004 , \22002 , \22003 );
xnor \U$21661 ( \22005 , \22004 , \21441 );
and \U$21662 ( \22006 , \21750 , \21450 );
and \U$21663 ( \22007 , \21689 , \21448 );
nor \U$21664 ( \22008 , \22006 , \22007 );
xnor \U$21665 ( \22009 , \22008 , \21457 );
and \U$21666 ( \22010 , \22005 , \22009 );
buf \U$21667 ( \22011 , RIbb31d70_145);
and \U$21668 ( \22012 , \22011 , \21469 );
and \U$21669 ( \22013 , \21813 , \21467 );
nor \U$21670 ( \22014 , \22012 , \22013 );
xnor \U$21671 ( \22015 , \22014 , \21476 );
and \U$21672 ( \22016 , \22009 , \22015 );
and \U$21673 ( \22017 , \22005 , \22015 );
or \U$21674 ( \22018 , \22010 , \22016 , \22017 );
and \U$21675 ( \22019 , \22000 , \22018 );
and \U$21676 ( \22020 , \21981 , \22018 );
or \U$21677 ( \22021 , \22001 , \22019 , \22020 );
and \U$21678 ( \22022 , \22011 , \21464 );
xor \U$21679 ( \22023 , \21890 , \21894 );
xor \U$21680 ( \22024 , \22023 , \21899 );
and \U$21681 ( \22025 , \22022 , \22024 );
xor \U$21682 ( \22026 , \21925 , \21929 );
xor \U$21683 ( \22027 , \22026 , \21934 );
and \U$21684 ( \22028 , \22024 , \22027 );
and \U$21685 ( \22029 , \22022 , \22027 );
or \U$21686 ( \22030 , \22025 , \22028 , \22029 );
and \U$21687 ( \22031 , \22021 , \22030 );
xor \U$21688 ( \22032 , \21824 , \21828 );
xor \U$21689 ( \22033 , \22032 , \21833 );
and \U$21690 ( \22034 , \22030 , \22033 );
and \U$21691 ( \22035 , \22021 , \22033 );
or \U$21692 ( \22036 , \22031 , \22034 , \22035 );
xor \U$21693 ( \22037 , \21817 , \21836 );
xor \U$21694 ( \22038 , \22037 , \21853 );
and \U$21695 ( \22039 , \22036 , \22038 );
xor \U$21696 ( \22040 , \21940 , \21945 );
xor \U$21697 ( \22041 , \22040 , \21948 );
and \U$21698 ( \22042 , \22038 , \22041 );
and \U$21699 ( \22043 , \22036 , \22041 );
or \U$21700 ( \22044 , \22039 , \22042 , \22043 );
buf \U$21701 ( \22045 , RIbb2ed28_20);
buf \U$21702 ( \22046 , RIbb2ecb0_21);
and \U$21703 ( \22047 , \22045 , \22046 );
not \U$21704 ( \22048 , \22047 );
and \U$21705 ( \22049 , \21904 , \22048 );
not \U$21706 ( \22050 , \22049 );
and \U$21707 ( \22051 , \21379 , \21985 );
and \U$21708 ( \22052 , \21387 , \21983 );
nor \U$21709 ( \22053 , \22051 , \22052 );
xnor \U$21710 ( \22054 , \22053 , \21907 );
and \U$21711 ( \22055 , \22050 , \22054 );
and \U$21712 ( \22056 , \21395 , \21821 );
and \U$21713 ( \22057 , \21403 , \21819 );
nor \U$21714 ( \22058 , \22056 , \22057 );
xnor \U$21715 ( \22059 , \22058 , \21727 );
and \U$21716 ( \22060 , \22054 , \22059 );
and \U$21717 ( \22061 , \22050 , \22059 );
or \U$21718 ( \22062 , \22055 , \22060 , \22061 );
and \U$21719 ( \22063 , \21413 , \21652 );
and \U$21720 ( \22064 , \21421 , \21650 );
nor \U$21721 ( \22065 , \22063 , \22064 );
xnor \U$21722 ( \22066 , \22065 , \21377 );
and \U$21723 ( \22067 , \21428 , \21385 );
and \U$21724 ( \22068 , \21436 , \21383 );
nor \U$21725 ( \22069 , \22067 , \22068 );
xnor \U$21726 ( \22070 , \22069 , \21392 );
and \U$21727 ( \22071 , \22066 , \22070 );
and \U$21728 ( \22072 , \21444 , \21401 );
and \U$21729 ( \22073 , \21452 , \21399 );
nor \U$21730 ( \22074 , \22072 , \22073 );
xnor \U$21731 ( \22075 , \22074 , \21408 );
and \U$21732 ( \22076 , \22070 , \22075 );
and \U$21733 ( \22077 , \22066 , \22075 );
or \U$21734 ( \22078 , \22071 , \22076 , \22077 );
and \U$21735 ( \22079 , \22062 , \22078 );
and \U$21736 ( \22080 , \21463 , \21419 );
and \U$21737 ( \22081 , \21471 , \21417 );
nor \U$21738 ( \22082 , \22080 , \22081 );
xnor \U$21739 ( \22083 , \22082 , \21426 );
and \U$21740 ( \22084 , \21689 , \21434 );
and \U$21741 ( \22085 , \21478 , \21432 );
nor \U$21742 ( \22086 , \22084 , \22085 );
xnor \U$21743 ( \22087 , \22086 , \21441 );
and \U$21744 ( \22088 , \22083 , \22087 );
and \U$21745 ( \22089 , \21813 , \21450 );
and \U$21746 ( \22090 , \21750 , \21448 );
nor \U$21747 ( \22091 , \22089 , \22090 );
xnor \U$21748 ( \22092 , \22091 , \21457 );
and \U$21749 ( \22093 , \22087 , \22092 );
and \U$21750 ( \22094 , \22083 , \22092 );
or \U$21751 ( \22095 , \22088 , \22093 , \22094 );
and \U$21752 ( \22096 , \22078 , \22095 );
and \U$21753 ( \22097 , \22062 , \22095 );
or \U$21754 ( \22098 , \22079 , \22096 , \22097 );
buf \U$21755 ( \22099 , RIbb31de8_146);
and \U$21756 ( \22100 , \22099 , \21464 );
xor \U$21757 ( \22101 , \22005 , \22009 );
xor \U$21758 ( \22102 , \22101 , \22015 );
or \U$21759 ( \22103 , \22100 , \22102 );
and \U$21760 ( \22104 , \22098 , \22103 );
xor \U$21761 ( \22105 , \21969 , \21973 );
xor \U$21762 ( \22106 , \22105 , \21978 );
xor \U$21763 ( \22107 , \21988 , \21992 );
xor \U$21764 ( \22108 , \22107 , \21997 );
and \U$21765 ( \22109 , \22106 , \22108 );
and \U$21766 ( \22110 , \22103 , \22109 );
and \U$21767 ( \22111 , \22098 , \22109 );
or \U$21768 ( \22112 , \22104 , \22110 , \22111 );
xor \U$21769 ( \22113 , \21908 , \21912 );
xor \U$21770 ( \22114 , \22113 , \21917 );
xor \U$21771 ( \22115 , \21981 , \22000 );
xor \U$21772 ( \22116 , \22115 , \22018 );
and \U$21773 ( \22117 , \22114 , \22116 );
xor \U$21774 ( \22118 , \22022 , \22024 );
xor \U$21775 ( \22119 , \22118 , \22027 );
and \U$21776 ( \22120 , \22116 , \22119 );
and \U$21777 ( \22121 , \22114 , \22119 );
or \U$21778 ( \22122 , \22117 , \22120 , \22121 );
and \U$21779 ( \22123 , \22112 , \22122 );
xnor \U$21780 ( \22124 , \21942 , \21944 );
and \U$21781 ( \22125 , \22122 , \22124 );
and \U$21782 ( \22126 , \22112 , \22124 );
or \U$21783 ( \22127 , \22123 , \22125 , \22126 );
xor \U$21784 ( \22128 , \21902 , \21920 );
xor \U$21785 ( \22129 , \22128 , \21937 );
xor \U$21786 ( \22130 , \22021 , \22030 );
xor \U$21787 ( \22131 , \22130 , \22033 );
and \U$21788 ( \22132 , \22129 , \22131 );
and \U$21789 ( \22133 , \22127 , \22132 );
xor \U$21790 ( \22134 , \22036 , \22038 );
xor \U$21791 ( \22135 , \22134 , \22041 );
and \U$21792 ( \22136 , \22132 , \22135 );
and \U$21793 ( \22137 , \22127 , \22135 );
or \U$21794 ( \22138 , \22133 , \22136 , \22137 );
and \U$21795 ( \22139 , \22044 , \22138 );
xor \U$21796 ( \22140 , \21951 , \21953 );
xor \U$21797 ( \22141 , \22140 , \21956 );
and \U$21798 ( \22142 , \22138 , \22141 );
and \U$21799 ( \22143 , \22044 , \22141 );
or \U$21800 ( \22144 , \22139 , \22142 , \22143 );
and \U$21801 ( \22145 , \21965 , \22144 );
xor \U$21802 ( \22146 , \21965 , \22144 );
xor \U$21803 ( \22147 , \22044 , \22138 );
xor \U$21804 ( \22148 , \22147 , \22141 );
and \U$21805 ( \22149 , \21478 , \21419 );
and \U$21806 ( \22150 , \21463 , \21417 );
nor \U$21807 ( \22151 , \22149 , \22150 );
xnor \U$21808 ( \22152 , \22151 , \21426 );
and \U$21809 ( \22153 , \21750 , \21434 );
and \U$21810 ( \22154 , \21689 , \21432 );
nor \U$21811 ( \22155 , \22153 , \22154 );
xnor \U$21812 ( \22156 , \22155 , \21441 );
and \U$21813 ( \22157 , \22152 , \22156 );
and \U$21814 ( \22158 , \22011 , \21450 );
and \U$21815 ( \22159 , \21813 , \21448 );
nor \U$21816 ( \22160 , \22158 , \22159 );
xnor \U$21817 ( \22161 , \22160 , \21457 );
and \U$21818 ( \22162 , \22156 , \22161 );
and \U$21819 ( \22163 , \22152 , \22161 );
or \U$21820 ( \22164 , \22157 , \22162 , \22163 );
and \U$21821 ( \22165 , \21436 , \21652 );
and \U$21822 ( \22166 , \21413 , \21650 );
nor \U$21823 ( \22167 , \22165 , \22166 );
xnor \U$21824 ( \22168 , \22167 , \21377 );
and \U$21825 ( \22169 , \21452 , \21385 );
and \U$21826 ( \22170 , \21428 , \21383 );
nor \U$21827 ( \22171 , \22169 , \22170 );
xnor \U$21828 ( \22172 , \22171 , \21392 );
and \U$21829 ( \22173 , \22168 , \22172 );
and \U$21830 ( \22174 , \21471 , \21401 );
and \U$21831 ( \22175 , \21444 , \21399 );
nor \U$21832 ( \22176 , \22174 , \22175 );
xnor \U$21833 ( \22177 , \22176 , \21408 );
and \U$21834 ( \22178 , \22172 , \22177 );
and \U$21835 ( \22179 , \22168 , \22177 );
or \U$21836 ( \22180 , \22173 , \22178 , \22179 );
and \U$21837 ( \22181 , \22164 , \22180 );
xor \U$21838 ( \22182 , \21904 , \22045 );
xor \U$21839 ( \22183 , \22045 , \22046 );
not \U$21840 ( \22184 , \22183 );
and \U$21841 ( \22185 , \22182 , \22184 );
and \U$21842 ( \22186 , \21387 , \22185 );
not \U$21843 ( \22187 , \22186 );
xnor \U$21844 ( \22188 , \22187 , \22049 );
and \U$21845 ( \22189 , \21403 , \21985 );
and \U$21846 ( \22190 , \21379 , \21983 );
nor \U$21847 ( \22191 , \22189 , \22190 );
xnor \U$21848 ( \22192 , \22191 , \21907 );
and \U$21849 ( \22193 , \22188 , \22192 );
and \U$21850 ( \22194 , \21421 , \21821 );
and \U$21851 ( \22195 , \21395 , \21819 );
nor \U$21852 ( \22196 , \22194 , \22195 );
xnor \U$21853 ( \22197 , \22196 , \21727 );
and \U$21854 ( \22198 , \22192 , \22197 );
and \U$21855 ( \22199 , \22188 , \22197 );
or \U$21856 ( \22200 , \22193 , \22198 , \22199 );
and \U$21857 ( \22201 , \22180 , \22200 );
and \U$21858 ( \22202 , \22164 , \22200 );
or \U$21859 ( \22203 , \22181 , \22201 , \22202 );
buf \U$21860 ( \22204 , RIbb31e60_147);
and \U$21861 ( \22205 , \22204 , \21469 );
and \U$21862 ( \22206 , \22099 , \21467 );
nor \U$21863 ( \22207 , \22205 , \22206 );
xnor \U$21864 ( \22208 , \22207 , \21476 );
buf \U$21865 ( \22209 , RIbb31ed8_148);
and \U$21866 ( \22210 , \22209 , \21464 );
or \U$21867 ( \22211 , \22208 , \22210 );
and \U$21868 ( \22212 , \22099 , \21469 );
and \U$21869 ( \22213 , \22011 , \21467 );
nor \U$21870 ( \22214 , \22212 , \22213 );
xnor \U$21871 ( \22215 , \22214 , \21476 );
and \U$21872 ( \22216 , \22211 , \22215 );
and \U$21873 ( \22217 , \22204 , \21464 );
and \U$21874 ( \22218 , \22215 , \22217 );
and \U$21875 ( \22219 , \22211 , \22217 );
or \U$21876 ( \22220 , \22216 , \22218 , \22219 );
and \U$21877 ( \22221 , \22203 , \22220 );
xor \U$21878 ( \22222 , \22050 , \22054 );
xor \U$21879 ( \22223 , \22222 , \22059 );
xor \U$21880 ( \22224 , \22066 , \22070 );
xor \U$21881 ( \22225 , \22224 , \22075 );
and \U$21882 ( \22226 , \22223 , \22225 );
xor \U$21883 ( \22227 , \22083 , \22087 );
xor \U$21884 ( \22228 , \22227 , \22092 );
and \U$21885 ( \22229 , \22225 , \22228 );
and \U$21886 ( \22230 , \22223 , \22228 );
or \U$21887 ( \22231 , \22226 , \22229 , \22230 );
and \U$21888 ( \22232 , \22220 , \22231 );
and \U$21889 ( \22233 , \22203 , \22231 );
or \U$21890 ( \22234 , \22221 , \22232 , \22233 );
xor \U$21891 ( \22235 , \22062 , \22078 );
xor \U$21892 ( \22236 , \22235 , \22095 );
xnor \U$21893 ( \22237 , \22100 , \22102 );
and \U$21894 ( \22238 , \22236 , \22237 );
xor \U$21895 ( \22239 , \22106 , \22108 );
and \U$21896 ( \22240 , \22237 , \22239 );
and \U$21897 ( \22241 , \22236 , \22239 );
or \U$21898 ( \22242 , \22238 , \22240 , \22241 );
and \U$21899 ( \22243 , \22234 , \22242 );
xor \U$21900 ( \22244 , \22114 , \22116 );
xor \U$21901 ( \22245 , \22244 , \22119 );
and \U$21902 ( \22246 , \22242 , \22245 );
and \U$21903 ( \22247 , \22234 , \22245 );
or \U$21904 ( \22248 , \22243 , \22246 , \22247 );
xor \U$21905 ( \22249 , \22112 , \22122 );
xor \U$21906 ( \22250 , \22249 , \22124 );
and \U$21907 ( \22251 , \22248 , \22250 );
xor \U$21908 ( \22252 , \22129 , \22131 );
and \U$21909 ( \22253 , \22250 , \22252 );
and \U$21910 ( \22254 , \22248 , \22252 );
or \U$21911 ( \22255 , \22251 , \22253 , \22254 );
xor \U$21912 ( \22256 , \22127 , \22132 );
xor \U$21913 ( \22257 , \22256 , \22135 );
and \U$21914 ( \22258 , \22255 , \22257 );
and \U$21915 ( \22259 , \22148 , \22258 );
xor \U$21916 ( \22260 , \22148 , \22258 );
xor \U$21917 ( \22261 , \22255 , \22257 );
buf \U$21918 ( \22262 , RIbb2ec38_22);
buf \U$21919 ( \22263 , RIbb2ebc0_23);
and \U$21920 ( \22264 , \22262 , \22263 );
not \U$21921 ( \22265 , \22264 );
and \U$21922 ( \22266 , \22046 , \22265 );
not \U$21923 ( \22267 , \22266 );
and \U$21924 ( \22268 , \21379 , \22185 );
and \U$21925 ( \22269 , \21387 , \22183 );
nor \U$21926 ( \22270 , \22268 , \22269 );
xnor \U$21927 ( \22271 , \22270 , \22049 );
and \U$21928 ( \22272 , \22267 , \22271 );
and \U$21929 ( \22273 , \21395 , \21985 );
and \U$21930 ( \22274 , \21403 , \21983 );
nor \U$21931 ( \22275 , \22273 , \22274 );
xnor \U$21932 ( \22276 , \22275 , \21907 );
and \U$21933 ( \22277 , \22271 , \22276 );
and \U$21934 ( \22278 , \22267 , \22276 );
or \U$21935 ( \22279 , \22272 , \22277 , \22278 );
and \U$21936 ( \22280 , \21463 , \21401 );
and \U$21937 ( \22281 , \21471 , \21399 );
nor \U$21938 ( \22282 , \22280 , \22281 );
xnor \U$21939 ( \22283 , \22282 , \21408 );
and \U$21940 ( \22284 , \21689 , \21419 );
and \U$21941 ( \22285 , \21478 , \21417 );
nor \U$21942 ( \22286 , \22284 , \22285 );
xnor \U$21943 ( \22287 , \22286 , \21426 );
and \U$21944 ( \22288 , \22283 , \22287 );
and \U$21945 ( \22289 , \21813 , \21434 );
and \U$21946 ( \22290 , \21750 , \21432 );
nor \U$21947 ( \22291 , \22289 , \22290 );
xnor \U$21948 ( \22292 , \22291 , \21441 );
and \U$21949 ( \22293 , \22287 , \22292 );
and \U$21950 ( \22294 , \22283 , \22292 );
or \U$21951 ( \22295 , \22288 , \22293 , \22294 );
and \U$21952 ( \22296 , \22279 , \22295 );
and \U$21953 ( \22297 , \21413 , \21821 );
and \U$21954 ( \22298 , \21421 , \21819 );
nor \U$21955 ( \22299 , \22297 , \22298 );
xnor \U$21956 ( \22300 , \22299 , \21727 );
and \U$21957 ( \22301 , \21428 , \21652 );
and \U$21958 ( \22302 , \21436 , \21650 );
nor \U$21959 ( \22303 , \22301 , \22302 );
xnor \U$21960 ( \22304 , \22303 , \21377 );
and \U$21961 ( \22305 , \22300 , \22304 );
and \U$21962 ( \22306 , \21444 , \21385 );
and \U$21963 ( \22307 , \21452 , \21383 );
nor \U$21964 ( \22308 , \22306 , \22307 );
xnor \U$21965 ( \22309 , \22308 , \21392 );
and \U$21966 ( \22310 , \22304 , \22309 );
and \U$21967 ( \22311 , \22300 , \22309 );
or \U$21968 ( \22312 , \22305 , \22310 , \22311 );
and \U$21969 ( \22313 , \22295 , \22312 );
and \U$21970 ( \22314 , \22279 , \22312 );
or \U$21971 ( \22315 , \22296 , \22313 , \22314 );
and \U$21972 ( \22316 , \22099 , \21450 );
and \U$21973 ( \22317 , \22011 , \21448 );
nor \U$21974 ( \22318 , \22316 , \22317 );
xnor \U$21975 ( \22319 , \22318 , \21457 );
and \U$21976 ( \22320 , \22209 , \21469 );
and \U$21977 ( \22321 , \22204 , \21467 );
nor \U$21978 ( \22322 , \22320 , \22321 );
xnor \U$21979 ( \22323 , \22322 , \21476 );
and \U$21980 ( \22324 , \22319 , \22323 );
buf \U$21981 ( \22325 , RIbb31f50_149);
and \U$21982 ( \22326 , \22325 , \21464 );
and \U$21983 ( \22327 , \22323 , \22326 );
and \U$21984 ( \22328 , \22319 , \22326 );
or \U$21985 ( \22329 , \22324 , \22327 , \22328 );
xor \U$21986 ( \22330 , \22152 , \22156 );
xor \U$21987 ( \22331 , \22330 , \22161 );
and \U$21988 ( \22332 , \22329 , \22331 );
xnor \U$21989 ( \22333 , \22208 , \22210 );
and \U$21990 ( \22334 , \22331 , \22333 );
and \U$21991 ( \22335 , \22329 , \22333 );
or \U$21992 ( \22336 , \22332 , \22334 , \22335 );
and \U$21993 ( \22337 , \22315 , \22336 );
xor \U$21994 ( \22338 , \22168 , \22172 );
xor \U$21995 ( \22339 , \22338 , \22177 );
xor \U$21996 ( \22340 , \22188 , \22192 );
xor \U$21997 ( \22341 , \22340 , \22197 );
and \U$21998 ( \22342 , \22339 , \22341 );
and \U$21999 ( \22343 , \22336 , \22342 );
and \U$22000 ( \22344 , \22315 , \22342 );
or \U$22001 ( \22345 , \22337 , \22343 , \22344 );
xor \U$22002 ( \22346 , \22164 , \22180 );
xor \U$22003 ( \22347 , \22346 , \22200 );
xor \U$22004 ( \22348 , \22211 , \22215 );
xor \U$22005 ( \22349 , \22348 , \22217 );
and \U$22006 ( \22350 , \22347 , \22349 );
xor \U$22007 ( \22351 , \22223 , \22225 );
xor \U$22008 ( \22352 , \22351 , \22228 );
and \U$22009 ( \22353 , \22349 , \22352 );
and \U$22010 ( \22354 , \22347 , \22352 );
or \U$22011 ( \22355 , \22350 , \22353 , \22354 );
and \U$22012 ( \22356 , \22345 , \22355 );
xor \U$22013 ( \22357 , \22236 , \22237 );
xor \U$22014 ( \22358 , \22357 , \22239 );
and \U$22015 ( \22359 , \22355 , \22358 );
and \U$22016 ( \22360 , \22345 , \22358 );
or \U$22017 ( \22361 , \22356 , \22359 , \22360 );
xor \U$22018 ( \22362 , \22098 , \22103 );
xor \U$22019 ( \22363 , \22362 , \22109 );
and \U$22020 ( \22364 , \22361 , \22363 );
xor \U$22021 ( \22365 , \22234 , \22242 );
xor \U$22022 ( \22366 , \22365 , \22245 );
and \U$22023 ( \22367 , \22363 , \22366 );
and \U$22024 ( \22368 , \22361 , \22366 );
or \U$22025 ( \22369 , \22364 , \22367 , \22368 );
xor \U$22026 ( \22370 , \22248 , \22250 );
xor \U$22027 ( \22371 , \22370 , \22252 );
and \U$22028 ( \22372 , \22369 , \22371 );
and \U$22029 ( \22373 , \22261 , \22372 );
xor \U$22030 ( \22374 , \22261 , \22372 );
xor \U$22031 ( \22375 , \22369 , \22371 );
xor \U$22032 ( \22376 , \22046 , \22262 );
xor \U$22033 ( \22377 , \22262 , \22263 );
not \U$22034 ( \22378 , \22377 );
and \U$22035 ( \22379 , \22376 , \22378 );
and \U$22036 ( \22380 , \21387 , \22379 );
not \U$22037 ( \22381 , \22380 );
xnor \U$22038 ( \22382 , \22381 , \22266 );
and \U$22039 ( \22383 , \21403 , \22185 );
and \U$22040 ( \22384 , \21379 , \22183 );
nor \U$22041 ( \22385 , \22383 , \22384 );
xnor \U$22042 ( \22386 , \22385 , \22049 );
and \U$22043 ( \22387 , \22382 , \22386 );
and \U$22044 ( \22388 , \21421 , \21985 );
and \U$22045 ( \22389 , \21395 , \21983 );
nor \U$22046 ( \22390 , \22388 , \22389 );
xnor \U$22047 ( \22391 , \22390 , \21907 );
and \U$22048 ( \22392 , \22386 , \22391 );
and \U$22049 ( \22393 , \22382 , \22391 );
or \U$22050 ( \22394 , \22387 , \22392 , \22393 );
and \U$22051 ( \22395 , \21478 , \21401 );
and \U$22052 ( \22396 , \21463 , \21399 );
nor \U$22053 ( \22397 , \22395 , \22396 );
xnor \U$22054 ( \22398 , \22397 , \21408 );
and \U$22055 ( \22399 , \21750 , \21419 );
and \U$22056 ( \22400 , \21689 , \21417 );
nor \U$22057 ( \22401 , \22399 , \22400 );
xnor \U$22058 ( \22402 , \22401 , \21426 );
and \U$22059 ( \22403 , \22398 , \22402 );
and \U$22060 ( \22404 , \22011 , \21434 );
and \U$22061 ( \22405 , \21813 , \21432 );
nor \U$22062 ( \22406 , \22404 , \22405 );
xnor \U$22063 ( \22407 , \22406 , \21441 );
and \U$22064 ( \22408 , \22402 , \22407 );
and \U$22065 ( \22409 , \22398 , \22407 );
or \U$22066 ( \22410 , \22403 , \22408 , \22409 );
and \U$22067 ( \22411 , \22394 , \22410 );
and \U$22068 ( \22412 , \21436 , \21821 );
and \U$22069 ( \22413 , \21413 , \21819 );
nor \U$22070 ( \22414 , \22412 , \22413 );
xnor \U$22071 ( \22415 , \22414 , \21727 );
and \U$22072 ( \22416 , \21452 , \21652 );
and \U$22073 ( \22417 , \21428 , \21650 );
nor \U$22074 ( \22418 , \22416 , \22417 );
xnor \U$22075 ( \22419 , \22418 , \21377 );
and \U$22076 ( \22420 , \22415 , \22419 );
and \U$22077 ( \22421 , \21471 , \21385 );
and \U$22078 ( \22422 , \21444 , \21383 );
nor \U$22079 ( \22423 , \22421 , \22422 );
xnor \U$22080 ( \22424 , \22423 , \21392 );
and \U$22081 ( \22425 , \22419 , \22424 );
and \U$22082 ( \22426 , \22415 , \22424 );
or \U$22083 ( \22427 , \22420 , \22425 , \22426 );
and \U$22084 ( \22428 , \22410 , \22427 );
and \U$22085 ( \22429 , \22394 , \22427 );
or \U$22086 ( \22430 , \22411 , \22428 , \22429 );
and \U$22087 ( \22431 , \22204 , \21450 );
and \U$22088 ( \22432 , \22099 , \21448 );
nor \U$22089 ( \22433 , \22431 , \22432 );
xnor \U$22090 ( \22434 , \22433 , \21457 );
and \U$22091 ( \22435 , \22325 , \21469 );
and \U$22092 ( \22436 , \22209 , \21467 );
nor \U$22093 ( \22437 , \22435 , \22436 );
xnor \U$22094 ( \22438 , \22437 , \21476 );
and \U$22095 ( \22439 , \22434 , \22438 );
buf \U$22096 ( \22440 , RIbb31fc8_150);
and \U$22097 ( \22441 , \22440 , \21464 );
and \U$22098 ( \22442 , \22438 , \22441 );
and \U$22099 ( \22443 , \22434 , \22441 );
or \U$22100 ( \22444 , \22439 , \22442 , \22443 );
xor \U$22101 ( \22445 , \22319 , \22323 );
xor \U$22102 ( \22446 , \22445 , \22326 );
and \U$22103 ( \22447 , \22444 , \22446 );
xor \U$22104 ( \22448 , \22283 , \22287 );
xor \U$22105 ( \22449 , \22448 , \22292 );
and \U$22106 ( \22450 , \22446 , \22449 );
and \U$22107 ( \22451 , \22444 , \22449 );
or \U$22108 ( \22452 , \22447 , \22450 , \22451 );
and \U$22109 ( \22453 , \22430 , \22452 );
xor \U$22110 ( \22454 , \22267 , \22271 );
xor \U$22111 ( \22455 , \22454 , \22276 );
xor \U$22112 ( \22456 , \22300 , \22304 );
xor \U$22113 ( \22457 , \22456 , \22309 );
and \U$22114 ( \22458 , \22455 , \22457 );
and \U$22115 ( \22459 , \22452 , \22458 );
and \U$22116 ( \22460 , \22430 , \22458 );
or \U$22117 ( \22461 , \22453 , \22459 , \22460 );
xor \U$22118 ( \22462 , \22279 , \22295 );
xor \U$22119 ( \22463 , \22462 , \22312 );
xor \U$22120 ( \22464 , \22329 , \22331 );
xor \U$22121 ( \22465 , \22464 , \22333 );
and \U$22122 ( \22466 , \22463 , \22465 );
xor \U$22123 ( \22467 , \22339 , \22341 );
and \U$22124 ( \22468 , \22465 , \22467 );
and \U$22125 ( \22469 , \22463 , \22467 );
or \U$22126 ( \22470 , \22466 , \22468 , \22469 );
and \U$22127 ( \22471 , \22461 , \22470 );
xor \U$22128 ( \22472 , \22347 , \22349 );
xor \U$22129 ( \22473 , \22472 , \22352 );
and \U$22130 ( \22474 , \22470 , \22473 );
and \U$22131 ( \22475 , \22461 , \22473 );
or \U$22132 ( \22476 , \22471 , \22474 , \22475 );
xor \U$22133 ( \22477 , \22203 , \22220 );
xor \U$22134 ( \22478 , \22477 , \22231 );
and \U$22135 ( \22479 , \22476 , \22478 );
xor \U$22136 ( \22480 , \22345 , \22355 );
xor \U$22137 ( \22481 , \22480 , \22358 );
and \U$22138 ( \22482 , \22478 , \22481 );
and \U$22139 ( \22483 , \22476 , \22481 );
or \U$22140 ( \22484 , \22479 , \22482 , \22483 );
xor \U$22141 ( \22485 , \22361 , \22363 );
xor \U$22142 ( \22486 , \22485 , \22366 );
and \U$22143 ( \22487 , \22484 , \22486 );
and \U$22144 ( \22488 , \22375 , \22487 );
xor \U$22145 ( \22489 , \22375 , \22487 );
xor \U$22146 ( \22490 , \22484 , \22486 );
buf \U$22147 ( \22491 , RIbb2eb48_24);
buf \U$22148 ( \22492 , RIbb2ead0_25);
and \U$22149 ( \22493 , \22491 , \22492 );
not \U$22150 ( \22494 , \22493 );
and \U$22151 ( \22495 , \22263 , \22494 );
not \U$22152 ( \22496 , \22495 );
and \U$22153 ( \22497 , \21379 , \22379 );
and \U$22154 ( \22498 , \21387 , \22377 );
nor \U$22155 ( \22499 , \22497 , \22498 );
xnor \U$22156 ( \22500 , \22499 , \22266 );
and \U$22157 ( \22501 , \22496 , \22500 );
and \U$22158 ( \22502 , \21395 , \22185 );
and \U$22159 ( \22503 , \21403 , \22183 );
nor \U$22160 ( \22504 , \22502 , \22503 );
xnor \U$22161 ( \22505 , \22504 , \22049 );
and \U$22162 ( \22506 , \22500 , \22505 );
and \U$22163 ( \22507 , \22496 , \22505 );
or \U$22164 ( \22508 , \22501 , \22506 , \22507 );
and \U$22165 ( \22509 , \21413 , \21985 );
and \U$22166 ( \22510 , \21421 , \21983 );
nor \U$22167 ( \22511 , \22509 , \22510 );
xnor \U$22168 ( \22512 , \22511 , \21907 );
and \U$22169 ( \22513 , \21428 , \21821 );
and \U$22170 ( \22514 , \21436 , \21819 );
nor \U$22171 ( \22515 , \22513 , \22514 );
xnor \U$22172 ( \22516 , \22515 , \21727 );
and \U$22173 ( \22517 , \22512 , \22516 );
and \U$22174 ( \22518 , \21444 , \21652 );
and \U$22175 ( \22519 , \21452 , \21650 );
nor \U$22176 ( \22520 , \22518 , \22519 );
xnor \U$22177 ( \22521 , \22520 , \21377 );
and \U$22178 ( \22522 , \22516 , \22521 );
and \U$22179 ( \22523 , \22512 , \22521 );
or \U$22180 ( \22524 , \22517 , \22522 , \22523 );
and \U$22181 ( \22525 , \22508 , \22524 );
and \U$22182 ( \22526 , \21463 , \21385 );
and \U$22183 ( \22527 , \21471 , \21383 );
nor \U$22184 ( \22528 , \22526 , \22527 );
xnor \U$22185 ( \22529 , \22528 , \21392 );
and \U$22186 ( \22530 , \21689 , \21401 );
and \U$22187 ( \22531 , \21478 , \21399 );
nor \U$22188 ( \22532 , \22530 , \22531 );
xnor \U$22189 ( \22533 , \22532 , \21408 );
and \U$22190 ( \22534 , \22529 , \22533 );
and \U$22191 ( \22535 , \21813 , \21419 );
and \U$22192 ( \22536 , \21750 , \21417 );
nor \U$22193 ( \22537 , \22535 , \22536 );
xnor \U$22194 ( \22538 , \22537 , \21426 );
and \U$22195 ( \22539 , \22533 , \22538 );
and \U$22196 ( \22540 , \22529 , \22538 );
or \U$22197 ( \22541 , \22534 , \22539 , \22540 );
and \U$22198 ( \22542 , \22524 , \22541 );
and \U$22199 ( \22543 , \22508 , \22541 );
or \U$22200 ( \22544 , \22525 , \22542 , \22543 );
xor \U$22201 ( \22545 , \22382 , \22386 );
xor \U$22202 ( \22546 , \22545 , \22391 );
xor \U$22203 ( \22547 , \22398 , \22402 );
xor \U$22204 ( \22548 , \22547 , \22407 );
and \U$22205 ( \22549 , \22546 , \22548 );
xor \U$22206 ( \22550 , \22415 , \22419 );
xor \U$22207 ( \22551 , \22550 , \22424 );
and \U$22208 ( \22552 , \22548 , \22551 );
and \U$22209 ( \22553 , \22546 , \22551 );
or \U$22210 ( \22554 , \22549 , \22552 , \22553 );
and \U$22211 ( \22555 , \22544 , \22554 );
and \U$22212 ( \22556 , \22099 , \21434 );
and \U$22213 ( \22557 , \22011 , \21432 );
nor \U$22214 ( \22558 , \22556 , \22557 );
xnor \U$22215 ( \22559 , \22558 , \21441 );
and \U$22216 ( \22560 , \22209 , \21450 );
and \U$22217 ( \22561 , \22204 , \21448 );
nor \U$22218 ( \22562 , \22560 , \22561 );
xnor \U$22219 ( \22563 , \22562 , \21457 );
and \U$22220 ( \22564 , \22559 , \22563 );
and \U$22221 ( \22565 , \22440 , \21469 );
and \U$22222 ( \22566 , \22325 , \21467 );
nor \U$22223 ( \22567 , \22565 , \22566 );
xnor \U$22224 ( \22568 , \22567 , \21476 );
and \U$22225 ( \22569 , \22563 , \22568 );
and \U$22226 ( \22570 , \22559 , \22568 );
or \U$22227 ( \22571 , \22564 , \22569 , \22570 );
xor \U$22228 ( \22572 , \22434 , \22438 );
xor \U$22229 ( \22573 , \22572 , \22441 );
or \U$22230 ( \22574 , \22571 , \22573 );
and \U$22231 ( \22575 , \22554 , \22574 );
and \U$22232 ( \22576 , \22544 , \22574 );
or \U$22233 ( \22577 , \22555 , \22575 , \22576 );
xor \U$22234 ( \22578 , \22394 , \22410 );
xor \U$22235 ( \22579 , \22578 , \22427 );
xor \U$22236 ( \22580 , \22444 , \22446 );
xor \U$22237 ( \22581 , \22580 , \22449 );
and \U$22238 ( \22582 , \22579 , \22581 );
xor \U$22239 ( \22583 , \22455 , \22457 );
and \U$22240 ( \22584 , \22581 , \22583 );
and \U$22241 ( \22585 , \22579 , \22583 );
or \U$22242 ( \22586 , \22582 , \22584 , \22585 );
and \U$22243 ( \22587 , \22577 , \22586 );
xor \U$22244 ( \22588 , \22463 , \22465 );
xor \U$22245 ( \22589 , \22588 , \22467 );
and \U$22246 ( \22590 , \22586 , \22589 );
and \U$22247 ( \22591 , \22577 , \22589 );
or \U$22248 ( \22592 , \22587 , \22590 , \22591 );
xor \U$22249 ( \22593 , \22315 , \22336 );
xor \U$22250 ( \22594 , \22593 , \22342 );
and \U$22251 ( \22595 , \22592 , \22594 );
xor \U$22252 ( \22596 , \22461 , \22470 );
xor \U$22253 ( \22597 , \22596 , \22473 );
and \U$22254 ( \22598 , \22594 , \22597 );
and \U$22255 ( \22599 , \22592 , \22597 );
or \U$22256 ( \22600 , \22595 , \22598 , \22599 );
xor \U$22257 ( \22601 , \22476 , \22478 );
xor \U$22258 ( \22602 , \22601 , \22481 );
and \U$22259 ( \22603 , \22600 , \22602 );
and \U$22260 ( \22604 , \22490 , \22603 );
xor \U$22261 ( \22605 , \22490 , \22603 );
xor \U$22262 ( \22606 , \22600 , \22602 );
and \U$22263 ( \22607 , \22204 , \21434 );
and \U$22264 ( \22608 , \22099 , \21432 );
nor \U$22265 ( \22609 , \22607 , \22608 );
xnor \U$22266 ( \22610 , \22609 , \21441 );
and \U$22267 ( \22611 , \22325 , \21450 );
and \U$22268 ( \22612 , \22209 , \21448 );
nor \U$22269 ( \22613 , \22611 , \22612 );
xnor \U$22270 ( \22614 , \22613 , \21457 );
and \U$22271 ( \22615 , \22610 , \22614 );
buf \U$22272 ( \22616 , RIbb32040_151);
and \U$22273 ( \22617 , \22616 , \21469 );
and \U$22274 ( \22618 , \22440 , \21467 );
nor \U$22275 ( \22619 , \22617 , \22618 );
xnor \U$22276 ( \22620 , \22619 , \21476 );
and \U$22277 ( \22621 , \22614 , \22620 );
and \U$22278 ( \22622 , \22610 , \22620 );
or \U$22279 ( \22623 , \22615 , \22621 , \22622 );
buf \U$22280 ( \22624 , RIbb320b8_152);
and \U$22281 ( \22625 , \22624 , \21464 );
buf \U$22282 ( \22626 , \22625 );
and \U$22283 ( \22627 , \22623 , \22626 );
and \U$22284 ( \22628 , \22616 , \21464 );
and \U$22285 ( \22629 , \22626 , \22628 );
and \U$22286 ( \22630 , \22623 , \22628 );
or \U$22287 ( \22631 , \22627 , \22629 , \22630 );
and \U$22288 ( \22632 , \21436 , \21985 );
and \U$22289 ( \22633 , \21413 , \21983 );
nor \U$22290 ( \22634 , \22632 , \22633 );
xnor \U$22291 ( \22635 , \22634 , \21907 );
and \U$22292 ( \22636 , \21452 , \21821 );
and \U$22293 ( \22637 , \21428 , \21819 );
nor \U$22294 ( \22638 , \22636 , \22637 );
xnor \U$22295 ( \22639 , \22638 , \21727 );
and \U$22296 ( \22640 , \22635 , \22639 );
and \U$22297 ( \22641 , \21471 , \21652 );
and \U$22298 ( \22642 , \21444 , \21650 );
nor \U$22299 ( \22643 , \22641 , \22642 );
xnor \U$22300 ( \22644 , \22643 , \21377 );
and \U$22301 ( \22645 , \22639 , \22644 );
and \U$22302 ( \22646 , \22635 , \22644 );
or \U$22303 ( \22647 , \22640 , \22645 , \22646 );
xor \U$22304 ( \22648 , \22263 , \22491 );
xor \U$22305 ( \22649 , \22491 , \22492 );
not \U$22306 ( \22650 , \22649 );
and \U$22307 ( \22651 , \22648 , \22650 );
and \U$22308 ( \22652 , \21387 , \22651 );
not \U$22309 ( \22653 , \22652 );
xnor \U$22310 ( \22654 , \22653 , \22495 );
and \U$22311 ( \22655 , \21403 , \22379 );
and \U$22312 ( \22656 , \21379 , \22377 );
nor \U$22313 ( \22657 , \22655 , \22656 );
xnor \U$22314 ( \22658 , \22657 , \22266 );
and \U$22315 ( \22659 , \22654 , \22658 );
and \U$22316 ( \22660 , \21421 , \22185 );
and \U$22317 ( \22661 , \21395 , \22183 );
nor \U$22318 ( \22662 , \22660 , \22661 );
xnor \U$22319 ( \22663 , \22662 , \22049 );
and \U$22320 ( \22664 , \22658 , \22663 );
and \U$22321 ( \22665 , \22654 , \22663 );
or \U$22322 ( \22666 , \22659 , \22664 , \22665 );
and \U$22323 ( \22667 , \22647 , \22666 );
and \U$22324 ( \22668 , \21478 , \21385 );
and \U$22325 ( \22669 , \21463 , \21383 );
nor \U$22326 ( \22670 , \22668 , \22669 );
xnor \U$22327 ( \22671 , \22670 , \21392 );
and \U$22328 ( \22672 , \21750 , \21401 );
and \U$22329 ( \22673 , \21689 , \21399 );
nor \U$22330 ( \22674 , \22672 , \22673 );
xnor \U$22331 ( \22675 , \22674 , \21408 );
and \U$22332 ( \22676 , \22671 , \22675 );
and \U$22333 ( \22677 , \22011 , \21419 );
and \U$22334 ( \22678 , \21813 , \21417 );
nor \U$22335 ( \22679 , \22677 , \22678 );
xnor \U$22336 ( \22680 , \22679 , \21426 );
and \U$22337 ( \22681 , \22675 , \22680 );
and \U$22338 ( \22682 , \22671 , \22680 );
or \U$22339 ( \22683 , \22676 , \22681 , \22682 );
and \U$22340 ( \22684 , \22666 , \22683 );
and \U$22341 ( \22685 , \22647 , \22683 );
or \U$22342 ( \22686 , \22667 , \22684 , \22685 );
and \U$22343 ( \22687 , \22631 , \22686 );
xor \U$22344 ( \22688 , \22512 , \22516 );
xor \U$22345 ( \22689 , \22688 , \22521 );
xor \U$22346 ( \22690 , \22559 , \22563 );
xor \U$22347 ( \22691 , \22690 , \22568 );
and \U$22348 ( \22692 , \22689 , \22691 );
xor \U$22349 ( \22693 , \22529 , \22533 );
xor \U$22350 ( \22694 , \22693 , \22538 );
and \U$22351 ( \22695 , \22691 , \22694 );
and \U$22352 ( \22696 , \22689 , \22694 );
or \U$22353 ( \22697 , \22692 , \22695 , \22696 );
and \U$22354 ( \22698 , \22686 , \22697 );
and \U$22355 ( \22699 , \22631 , \22697 );
or \U$22356 ( \22700 , \22687 , \22698 , \22699 );
xor \U$22357 ( \22701 , \22508 , \22524 );
xor \U$22358 ( \22702 , \22701 , \22541 );
xor \U$22359 ( \22703 , \22546 , \22548 );
xor \U$22360 ( \22704 , \22703 , \22551 );
and \U$22361 ( \22705 , \22702 , \22704 );
xnor \U$22362 ( \22706 , \22571 , \22573 );
and \U$22363 ( \22707 , \22704 , \22706 );
and \U$22364 ( \22708 , \22702 , \22706 );
or \U$22365 ( \22709 , \22705 , \22707 , \22708 );
and \U$22366 ( \22710 , \22700 , \22709 );
xor \U$22367 ( \22711 , \22579 , \22581 );
xor \U$22368 ( \22712 , \22711 , \22583 );
and \U$22369 ( \22713 , \22709 , \22712 );
and \U$22370 ( \22714 , \22700 , \22712 );
or \U$22371 ( \22715 , \22710 , \22713 , \22714 );
xor \U$22372 ( \22716 , \22430 , \22452 );
xor \U$22373 ( \22717 , \22716 , \22458 );
and \U$22374 ( \22718 , \22715 , \22717 );
xor \U$22375 ( \22719 , \22577 , \22586 );
xor \U$22376 ( \22720 , \22719 , \22589 );
and \U$22377 ( \22721 , \22717 , \22720 );
and \U$22378 ( \22722 , \22715 , \22720 );
or \U$22379 ( \22723 , \22718 , \22721 , \22722 );
xor \U$22380 ( \22724 , \22592 , \22594 );
xor \U$22381 ( \22725 , \22724 , \22597 );
and \U$22382 ( \22726 , \22723 , \22725 );
and \U$22383 ( \22727 , \22606 , \22726 );
xor \U$22384 ( \22728 , \22606 , \22726 );
xor \U$22385 ( \22729 , \22723 , \22725 );
and \U$22386 ( \22730 , \21463 , \21652 );
and \U$22387 ( \22731 , \21471 , \21650 );
nor \U$22388 ( \22732 , \22730 , \22731 );
xnor \U$22389 ( \22733 , \22732 , \21377 );
and \U$22390 ( \22734 , \21689 , \21385 );
and \U$22391 ( \22735 , \21478 , \21383 );
nor \U$22392 ( \22736 , \22734 , \22735 );
xnor \U$22393 ( \22737 , \22736 , \21392 );
and \U$22394 ( \22738 , \22733 , \22737 );
and \U$22395 ( \22739 , \21813 , \21401 );
and \U$22396 ( \22740 , \21750 , \21399 );
nor \U$22397 ( \22741 , \22739 , \22740 );
xnor \U$22398 ( \22742 , \22741 , \21408 );
and \U$22399 ( \22743 , \22737 , \22742 );
and \U$22400 ( \22744 , \22733 , \22742 );
or \U$22401 ( \22745 , \22738 , \22743 , \22744 );
and \U$22402 ( \22746 , \21413 , \22185 );
and \U$22403 ( \22747 , \21421 , \22183 );
nor \U$22404 ( \22748 , \22746 , \22747 );
xnor \U$22405 ( \22749 , \22748 , \22049 );
and \U$22406 ( \22750 , \21428 , \21985 );
and \U$22407 ( \22751 , \21436 , \21983 );
nor \U$22408 ( \22752 , \22750 , \22751 );
xnor \U$22409 ( \22753 , \22752 , \21907 );
and \U$22410 ( \22754 , \22749 , \22753 );
and \U$22411 ( \22755 , \21444 , \21821 );
and \U$22412 ( \22756 , \21452 , \21819 );
nor \U$22413 ( \22757 , \22755 , \22756 );
xnor \U$22414 ( \22758 , \22757 , \21727 );
and \U$22415 ( \22759 , \22753 , \22758 );
and \U$22416 ( \22760 , \22749 , \22758 );
or \U$22417 ( \22761 , \22754 , \22759 , \22760 );
and \U$22418 ( \22762 , \22745 , \22761 );
buf \U$22419 ( \22763 , RIbb2ea58_26);
buf \U$22420 ( \22764 , RIbb2e9e0_27);
and \U$22421 ( \22765 , \22763 , \22764 );
not \U$22422 ( \22766 , \22765 );
and \U$22423 ( \22767 , \22492 , \22766 );
not \U$22424 ( \22768 , \22767 );
and \U$22425 ( \22769 , \21379 , \22651 );
and \U$22426 ( \22770 , \21387 , \22649 );
nor \U$22427 ( \22771 , \22769 , \22770 );
xnor \U$22428 ( \22772 , \22771 , \22495 );
and \U$22429 ( \22773 , \22768 , \22772 );
and \U$22430 ( \22774 , \21395 , \22379 );
and \U$22431 ( \22775 , \21403 , \22377 );
nor \U$22432 ( \22776 , \22774 , \22775 );
xnor \U$22433 ( \22777 , \22776 , \22266 );
and \U$22434 ( \22778 , \22772 , \22777 );
and \U$22435 ( \22779 , \22768 , \22777 );
or \U$22436 ( \22780 , \22773 , \22778 , \22779 );
and \U$22437 ( \22781 , \22761 , \22780 );
and \U$22438 ( \22782 , \22745 , \22780 );
or \U$22439 ( \22783 , \22762 , \22781 , \22782 );
xor \U$22440 ( \22784 , \22635 , \22639 );
xor \U$22441 ( \22785 , \22784 , \22644 );
xor \U$22442 ( \22786 , \22654 , \22658 );
xor \U$22443 ( \22787 , \22786 , \22663 );
and \U$22444 ( \22788 , \22785 , \22787 );
xor \U$22445 ( \22789 , \22671 , \22675 );
xor \U$22446 ( \22790 , \22789 , \22680 );
and \U$22447 ( \22791 , \22787 , \22790 );
and \U$22448 ( \22792 , \22785 , \22790 );
or \U$22449 ( \22793 , \22788 , \22791 , \22792 );
and \U$22450 ( \22794 , \22783 , \22793 );
and \U$22451 ( \22795 , \22099 , \21419 );
and \U$22452 ( \22796 , \22011 , \21417 );
nor \U$22453 ( \22797 , \22795 , \22796 );
xnor \U$22454 ( \22798 , \22797 , \21426 );
and \U$22455 ( \22799 , \22209 , \21434 );
and \U$22456 ( \22800 , \22204 , \21432 );
nor \U$22457 ( \22801 , \22799 , \22800 );
xnor \U$22458 ( \22802 , \22801 , \21441 );
and \U$22459 ( \22803 , \22798 , \22802 );
and \U$22460 ( \22804 , \22440 , \21450 );
and \U$22461 ( \22805 , \22325 , \21448 );
nor \U$22462 ( \22806 , \22804 , \22805 );
xnor \U$22463 ( \22807 , \22806 , \21457 );
and \U$22464 ( \22808 , \22802 , \22807 );
and \U$22465 ( \22809 , \22798 , \22807 );
or \U$22466 ( \22810 , \22803 , \22808 , \22809 );
xor \U$22467 ( \22811 , \22610 , \22614 );
xor \U$22468 ( \22812 , \22811 , \22620 );
and \U$22469 ( \22813 , \22810 , \22812 );
not \U$22470 ( \22814 , \22625 );
and \U$22471 ( \22815 , \22812 , \22814 );
and \U$22472 ( \22816 , \22810 , \22814 );
or \U$22473 ( \22817 , \22813 , \22815 , \22816 );
and \U$22474 ( \22818 , \22793 , \22817 );
and \U$22475 ( \22819 , \22783 , \22817 );
or \U$22476 ( \22820 , \22794 , \22818 , \22819 );
xor \U$22477 ( \22821 , \22496 , \22500 );
xor \U$22478 ( \22822 , \22821 , \22505 );
xor \U$22479 ( \22823 , \22623 , \22626 );
xor \U$22480 ( \22824 , \22823 , \22628 );
and \U$22481 ( \22825 , \22822 , \22824 );
xor \U$22482 ( \22826 , \22689 , \22691 );
xor \U$22483 ( \22827 , \22826 , \22694 );
and \U$22484 ( \22828 , \22824 , \22827 );
and \U$22485 ( \22829 , \22822 , \22827 );
or \U$22486 ( \22830 , \22825 , \22828 , \22829 );
and \U$22487 ( \22831 , \22820 , \22830 );
xor \U$22488 ( \22832 , \22702 , \22704 );
xor \U$22489 ( \22833 , \22832 , \22706 );
and \U$22490 ( \22834 , \22830 , \22833 );
and \U$22491 ( \22835 , \22820 , \22833 );
or \U$22492 ( \22836 , \22831 , \22834 , \22835 );
xor \U$22493 ( \22837 , \22544 , \22554 );
xor \U$22494 ( \22838 , \22837 , \22574 );
and \U$22495 ( \22839 , \22836 , \22838 );
xor \U$22496 ( \22840 , \22700 , \22709 );
xor \U$22497 ( \22841 , \22840 , \22712 );
and \U$22498 ( \22842 , \22838 , \22841 );
and \U$22499 ( \22843 , \22836 , \22841 );
or \U$22500 ( \22844 , \22839 , \22842 , \22843 );
xor \U$22501 ( \22845 , \22715 , \22717 );
xor \U$22502 ( \22846 , \22845 , \22720 );
and \U$22503 ( \22847 , \22844 , \22846 );
and \U$22504 ( \22848 , \22729 , \22847 );
xor \U$22505 ( \22849 , \22729 , \22847 );
xor \U$22506 ( \22850 , \22844 , \22846 );
and \U$22507 ( \22851 , \22204 , \21419 );
and \U$22508 ( \22852 , \22099 , \21417 );
nor \U$22509 ( \22853 , \22851 , \22852 );
xnor \U$22510 ( \22854 , \22853 , \21426 );
and \U$22511 ( \22855 , \22325 , \21434 );
and \U$22512 ( \22856 , \22209 , \21432 );
nor \U$22513 ( \22857 , \22855 , \22856 );
xnor \U$22514 ( \22858 , \22857 , \21441 );
and \U$22515 ( \22859 , \22854 , \22858 );
and \U$22516 ( \22860 , \22616 , \21450 );
and \U$22517 ( \22861 , \22440 , \21448 );
nor \U$22518 ( \22862 , \22860 , \22861 );
xnor \U$22519 ( \22863 , \22862 , \21457 );
and \U$22520 ( \22864 , \22858 , \22863 );
and \U$22521 ( \22865 , \22854 , \22863 );
or \U$22522 ( \22866 , \22859 , \22864 , \22865 );
buf \U$22523 ( \22867 , RIbb32130_153);
and \U$22524 ( \22868 , \22867 , \21469 );
and \U$22525 ( \22869 , \22624 , \21467 );
nor \U$22526 ( \22870 , \22868 , \22869 );
xnor \U$22527 ( \22871 , \22870 , \21476 );
buf \U$22528 ( \22872 , RIbb321a8_154);
and \U$22529 ( \22873 , \22872 , \21464 );
or \U$22530 ( \22874 , \22871 , \22873 );
and \U$22531 ( \22875 , \22866 , \22874 );
and \U$22532 ( \22876 , \22624 , \21469 );
and \U$22533 ( \22877 , \22616 , \21467 );
nor \U$22534 ( \22878 , \22876 , \22877 );
xnor \U$22535 ( \22879 , \22878 , \21476 );
and \U$22536 ( \22880 , \22874 , \22879 );
and \U$22537 ( \22881 , \22866 , \22879 );
or \U$22538 ( \22882 , \22875 , \22880 , \22881 );
and \U$22539 ( \22883 , \21478 , \21652 );
and \U$22540 ( \22884 , \21463 , \21650 );
nor \U$22541 ( \22885 , \22883 , \22884 );
xnor \U$22542 ( \22886 , \22885 , \21377 );
and \U$22543 ( \22887 , \21750 , \21385 );
and \U$22544 ( \22888 , \21689 , \21383 );
nor \U$22545 ( \22889 , \22887 , \22888 );
xnor \U$22546 ( \22890 , \22889 , \21392 );
and \U$22547 ( \22891 , \22886 , \22890 );
and \U$22548 ( \22892 , \22011 , \21401 );
and \U$22549 ( \22893 , \21813 , \21399 );
nor \U$22550 ( \22894 , \22892 , \22893 );
xnor \U$22551 ( \22895 , \22894 , \21408 );
and \U$22552 ( \22896 , \22890 , \22895 );
and \U$22553 ( \22897 , \22886 , \22895 );
or \U$22554 ( \22898 , \22891 , \22896 , \22897 );
and \U$22555 ( \22899 , \21436 , \22185 );
and \U$22556 ( \22900 , \21413 , \22183 );
nor \U$22557 ( \22901 , \22899 , \22900 );
xnor \U$22558 ( \22902 , \22901 , \22049 );
and \U$22559 ( \22903 , \21452 , \21985 );
and \U$22560 ( \22904 , \21428 , \21983 );
nor \U$22561 ( \22905 , \22903 , \22904 );
xnor \U$22562 ( \22906 , \22905 , \21907 );
and \U$22563 ( \22907 , \22902 , \22906 );
and \U$22564 ( \22908 , \21471 , \21821 );
and \U$22565 ( \22909 , \21444 , \21819 );
nor \U$22566 ( \22910 , \22908 , \22909 );
xnor \U$22567 ( \22911 , \22910 , \21727 );
and \U$22568 ( \22912 , \22906 , \22911 );
and \U$22569 ( \22913 , \22902 , \22911 );
or \U$22570 ( \22914 , \22907 , \22912 , \22913 );
and \U$22571 ( \22915 , \22898 , \22914 );
xor \U$22572 ( \22916 , \22492 , \22763 );
xor \U$22573 ( \22917 , \22763 , \22764 );
not \U$22574 ( \22918 , \22917 );
and \U$22575 ( \22919 , \22916 , \22918 );
and \U$22576 ( \22920 , \21387 , \22919 );
not \U$22577 ( \22921 , \22920 );
xnor \U$22578 ( \22922 , \22921 , \22767 );
and \U$22579 ( \22923 , \21403 , \22651 );
and \U$22580 ( \22924 , \21379 , \22649 );
nor \U$22581 ( \22925 , \22923 , \22924 );
xnor \U$22582 ( \22926 , \22925 , \22495 );
and \U$22583 ( \22927 , \22922 , \22926 );
and \U$22584 ( \22928 , \21421 , \22379 );
and \U$22585 ( \22929 , \21395 , \22377 );
nor \U$22586 ( \22930 , \22928 , \22929 );
xnor \U$22587 ( \22931 , \22930 , \22266 );
and \U$22588 ( \22932 , \22926 , \22931 );
and \U$22589 ( \22933 , \22922 , \22931 );
or \U$22590 ( \22934 , \22927 , \22932 , \22933 );
and \U$22591 ( \22935 , \22914 , \22934 );
and \U$22592 ( \22936 , \22898 , \22934 );
or \U$22593 ( \22937 , \22915 , \22935 , \22936 );
and \U$22594 ( \22938 , \22882 , \22937 );
and \U$22595 ( \22939 , \22867 , \21464 );
xor \U$22596 ( \22940 , \22733 , \22737 );
xor \U$22597 ( \22941 , \22940 , \22742 );
and \U$22598 ( \22942 , \22939 , \22941 );
xor \U$22599 ( \22943 , \22798 , \22802 );
xor \U$22600 ( \22944 , \22943 , \22807 );
and \U$22601 ( \22945 , \22941 , \22944 );
and \U$22602 ( \22946 , \22939 , \22944 );
or \U$22603 ( \22947 , \22942 , \22945 , \22946 );
and \U$22604 ( \22948 , \22937 , \22947 );
and \U$22605 ( \22949 , \22882 , \22947 );
or \U$22606 ( \22950 , \22938 , \22948 , \22949 );
xor \U$22607 ( \22951 , \22745 , \22761 );
xor \U$22608 ( \22952 , \22951 , \22780 );
xor \U$22609 ( \22953 , \22785 , \22787 );
xor \U$22610 ( \22954 , \22953 , \22790 );
and \U$22611 ( \22955 , \22952 , \22954 );
xor \U$22612 ( \22956 , \22810 , \22812 );
xor \U$22613 ( \22957 , \22956 , \22814 );
and \U$22614 ( \22958 , \22954 , \22957 );
and \U$22615 ( \22959 , \22952 , \22957 );
or \U$22616 ( \22960 , \22955 , \22958 , \22959 );
and \U$22617 ( \22961 , \22950 , \22960 );
xor \U$22618 ( \22962 , \22647 , \22666 );
xor \U$22619 ( \22963 , \22962 , \22683 );
and \U$22620 ( \22964 , \22960 , \22963 );
and \U$22621 ( \22965 , \22950 , \22963 );
or \U$22622 ( \22966 , \22961 , \22964 , \22965 );
xor \U$22623 ( \22967 , \22783 , \22793 );
xor \U$22624 ( \22968 , \22967 , \22817 );
xor \U$22625 ( \22969 , \22822 , \22824 );
xor \U$22626 ( \22970 , \22969 , \22827 );
and \U$22627 ( \22971 , \22968 , \22970 );
and \U$22628 ( \22972 , \22966 , \22971 );
xor \U$22629 ( \22973 , \22631 , \22686 );
xor \U$22630 ( \22974 , \22973 , \22697 );
and \U$22631 ( \22975 , \22971 , \22974 );
and \U$22632 ( \22976 , \22966 , \22974 );
or \U$22633 ( \22977 , \22972 , \22975 , \22976 );
xor \U$22634 ( \22978 , \22836 , \22838 );
xor \U$22635 ( \22979 , \22978 , \22841 );
and \U$22636 ( \22980 , \22977 , \22979 );
and \U$22637 ( \22981 , \22850 , \22980 );
xor \U$22638 ( \22982 , \22850 , \22980 );
xor \U$22639 ( \22983 , \22977 , \22979 );
buf \U$22640 ( \22984 , RIbb2e968_28);
buf \U$22641 ( \22985 , RIbb2e8f0_29);
and \U$22642 ( \22986 , \22984 , \22985 );
not \U$22643 ( \22987 , \22986 );
and \U$22644 ( \22988 , \22764 , \22987 );
not \U$22645 ( \22989 , \22988 );
and \U$22646 ( \22990 , \21379 , \22919 );
and \U$22647 ( \22991 , \21387 , \22917 );
nor \U$22648 ( \22992 , \22990 , \22991 );
xnor \U$22649 ( \22993 , \22992 , \22767 );
and \U$22650 ( \22994 , \22989 , \22993 );
and \U$22651 ( \22995 , \21395 , \22651 );
and \U$22652 ( \22996 , \21403 , \22649 );
nor \U$22653 ( \22997 , \22995 , \22996 );
xnor \U$22654 ( \22998 , \22997 , \22495 );
and \U$22655 ( \22999 , \22993 , \22998 );
and \U$22656 ( \23000 , \22989 , \22998 );
or \U$22657 ( \23001 , \22994 , \22999 , \23000 );
and \U$22658 ( \23002 , \21413 , \22379 );
and \U$22659 ( \23003 , \21421 , \22377 );
nor \U$22660 ( \23004 , \23002 , \23003 );
xnor \U$22661 ( \23005 , \23004 , \22266 );
and \U$22662 ( \23006 , \21428 , \22185 );
and \U$22663 ( \23007 , \21436 , \22183 );
nor \U$22664 ( \23008 , \23006 , \23007 );
xnor \U$22665 ( \23009 , \23008 , \22049 );
and \U$22666 ( \23010 , \23005 , \23009 );
and \U$22667 ( \23011 , \21444 , \21985 );
and \U$22668 ( \23012 , \21452 , \21983 );
nor \U$22669 ( \23013 , \23011 , \23012 );
xnor \U$22670 ( \23014 , \23013 , \21907 );
and \U$22671 ( \23015 , \23009 , \23014 );
and \U$22672 ( \23016 , \23005 , \23014 );
or \U$22673 ( \23017 , \23010 , \23015 , \23016 );
and \U$22674 ( \23018 , \23001 , \23017 );
and \U$22675 ( \23019 , \21463 , \21821 );
and \U$22676 ( \23020 , \21471 , \21819 );
nor \U$22677 ( \23021 , \23019 , \23020 );
xnor \U$22678 ( \23022 , \23021 , \21727 );
and \U$22679 ( \23023 , \21689 , \21652 );
and \U$22680 ( \23024 , \21478 , \21650 );
nor \U$22681 ( \23025 , \23023 , \23024 );
xnor \U$22682 ( \23026 , \23025 , \21377 );
and \U$22683 ( \23027 , \23022 , \23026 );
and \U$22684 ( \23028 , \21813 , \21385 );
and \U$22685 ( \23029 , \21750 , \21383 );
nor \U$22686 ( \23030 , \23028 , \23029 );
xnor \U$22687 ( \23031 , \23030 , \21392 );
and \U$22688 ( \23032 , \23026 , \23031 );
and \U$22689 ( \23033 , \23022 , \23031 );
or \U$22690 ( \23034 , \23027 , \23032 , \23033 );
and \U$22691 ( \23035 , \23017 , \23034 );
and \U$22692 ( \23036 , \23001 , \23034 );
or \U$22693 ( \23037 , \23018 , \23035 , \23036 );
xor \U$22694 ( \23038 , \22886 , \22890 );
xor \U$22695 ( \23039 , \23038 , \22895 );
xor \U$22696 ( \23040 , \22902 , \22906 );
xor \U$22697 ( \23041 , \23040 , \22911 );
and \U$22698 ( \23042 , \23039 , \23041 );
xor \U$22699 ( \23043 , \22854 , \22858 );
xor \U$22700 ( \23044 , \23043 , \22863 );
and \U$22701 ( \23045 , \23041 , \23044 );
and \U$22702 ( \23046 , \23039 , \23044 );
or \U$22703 ( \23047 , \23042 , \23045 , \23046 );
and \U$22704 ( \23048 , \23037 , \23047 );
and \U$22705 ( \23049 , \22624 , \21450 );
and \U$22706 ( \23050 , \22616 , \21448 );
nor \U$22707 ( \23051 , \23049 , \23050 );
xnor \U$22708 ( \23052 , \23051 , \21457 );
and \U$22709 ( \23053 , \22872 , \21469 );
and \U$22710 ( \23054 , \22867 , \21467 );
nor \U$22711 ( \23055 , \23053 , \23054 );
xnor \U$22712 ( \23056 , \23055 , \21476 );
and \U$22713 ( \23057 , \23052 , \23056 );
buf \U$22714 ( \23058 , RIbb32220_155);
and \U$22715 ( \23059 , \23058 , \21464 );
and \U$22716 ( \23060 , \23056 , \23059 );
and \U$22717 ( \23061 , \23052 , \23059 );
or \U$22718 ( \23062 , \23057 , \23060 , \23061 );
and \U$22719 ( \23063 , \22099 , \21401 );
and \U$22720 ( \23064 , \22011 , \21399 );
nor \U$22721 ( \23065 , \23063 , \23064 );
xnor \U$22722 ( \23066 , \23065 , \21408 );
and \U$22723 ( \23067 , \22209 , \21419 );
and \U$22724 ( \23068 , \22204 , \21417 );
nor \U$22725 ( \23069 , \23067 , \23068 );
xnor \U$22726 ( \23070 , \23069 , \21426 );
and \U$22727 ( \23071 , \23066 , \23070 );
and \U$22728 ( \23072 , \22440 , \21434 );
and \U$22729 ( \23073 , \22325 , \21432 );
nor \U$22730 ( \23074 , \23072 , \23073 );
xnor \U$22731 ( \23075 , \23074 , \21441 );
and \U$22732 ( \23076 , \23070 , \23075 );
and \U$22733 ( \23077 , \23066 , \23075 );
or \U$22734 ( \23078 , \23071 , \23076 , \23077 );
and \U$22735 ( \23079 , \23062 , \23078 );
xnor \U$22736 ( \23080 , \22871 , \22873 );
and \U$22737 ( \23081 , \23078 , \23080 );
and \U$22738 ( \23082 , \23062 , \23080 );
or \U$22739 ( \23083 , \23079 , \23081 , \23082 );
and \U$22740 ( \23084 , \23047 , \23083 );
and \U$22741 ( \23085 , \23037 , \23083 );
or \U$22742 ( \23086 , \23048 , \23084 , \23085 );
xor \U$22743 ( \23087 , \22749 , \22753 );
xor \U$22744 ( \23088 , \23087 , \22758 );
xor \U$22745 ( \23089 , \22768 , \22772 );
xor \U$22746 ( \23090 , \23089 , \22777 );
and \U$22747 ( \23091 , \23088 , \23090 );
xor \U$22748 ( \23092 , \22939 , \22941 );
xor \U$22749 ( \23093 , \23092 , \22944 );
and \U$22750 ( \23094 , \23090 , \23093 );
and \U$22751 ( \23095 , \23088 , \23093 );
or \U$22752 ( \23096 , \23091 , \23094 , \23095 );
and \U$22753 ( \23097 , \23086 , \23096 );
xor \U$22754 ( \23098 , \22952 , \22954 );
xor \U$22755 ( \23099 , \23098 , \22957 );
and \U$22756 ( \23100 , \23096 , \23099 );
and \U$22757 ( \23101 , \23086 , \23099 );
or \U$22758 ( \23102 , \23097 , \23100 , \23101 );
xor \U$22759 ( \23103 , \22950 , \22960 );
xor \U$22760 ( \23104 , \23103 , \22963 );
and \U$22761 ( \23105 , \23102 , \23104 );
xor \U$22762 ( \23106 , \22968 , \22970 );
and \U$22763 ( \23107 , \23104 , \23106 );
and \U$22764 ( \23108 , \23102 , \23106 );
or \U$22765 ( \23109 , \23105 , \23107 , \23108 );
xor \U$22766 ( \23110 , \22966 , \22971 );
xor \U$22767 ( \23111 , \23110 , \22974 );
and \U$22768 ( \23112 , \23109 , \23111 );
xor \U$22769 ( \23113 , \22820 , \22830 );
xor \U$22770 ( \23114 , \23113 , \22833 );
and \U$22771 ( \23115 , \23111 , \23114 );
and \U$22772 ( \23116 , \23109 , \23114 );
or \U$22773 ( \23117 , \23112 , \23115 , \23116 );
and \U$22774 ( \23118 , \22983 , \23117 );
xor \U$22775 ( \23119 , \22983 , \23117 );
xor \U$22776 ( \23120 , \23109 , \23111 );
xor \U$22777 ( \23121 , \23120 , \23114 );
xor \U$22778 ( \23122 , \22764 , \22984 );
xor \U$22779 ( \23123 , \22984 , \22985 );
not \U$22780 ( \23124 , \23123 );
and \U$22781 ( \23125 , \23122 , \23124 );
and \U$22782 ( \23126 , \21387 , \23125 );
not \U$22783 ( \23127 , \23126 );
xnor \U$22784 ( \23128 , \23127 , \22988 );
and \U$22785 ( \23129 , \21403 , \22919 );
and \U$22786 ( \23130 , \21379 , \22917 );
nor \U$22787 ( \23131 , \23129 , \23130 );
xnor \U$22788 ( \23132 , \23131 , \22767 );
and \U$22789 ( \23133 , \23128 , \23132 );
and \U$22790 ( \23134 , \21421 , \22651 );
and \U$22791 ( \23135 , \21395 , \22649 );
nor \U$22792 ( \23136 , \23134 , \23135 );
xnor \U$22793 ( \23137 , \23136 , \22495 );
and \U$22794 ( \23138 , \23132 , \23137 );
and \U$22795 ( \23139 , \23128 , \23137 );
or \U$22796 ( \23140 , \23133 , \23138 , \23139 );
and \U$22797 ( \23141 , \21436 , \22379 );
and \U$22798 ( \23142 , \21413 , \22377 );
nor \U$22799 ( \23143 , \23141 , \23142 );
xnor \U$22800 ( \23144 , \23143 , \22266 );
and \U$22801 ( \23145 , \21452 , \22185 );
and \U$22802 ( \23146 , \21428 , \22183 );
nor \U$22803 ( \23147 , \23145 , \23146 );
xnor \U$22804 ( \23148 , \23147 , \22049 );
and \U$22805 ( \23149 , \23144 , \23148 );
and \U$22806 ( \23150 , \21471 , \21985 );
and \U$22807 ( \23151 , \21444 , \21983 );
nor \U$22808 ( \23152 , \23150 , \23151 );
xnor \U$22809 ( \23153 , \23152 , \21907 );
and \U$22810 ( \23154 , \23148 , \23153 );
and \U$22811 ( \23155 , \23144 , \23153 );
or \U$22812 ( \23156 , \23149 , \23154 , \23155 );
and \U$22813 ( \23157 , \23140 , \23156 );
and \U$22814 ( \23158 , \21478 , \21821 );
and \U$22815 ( \23159 , \21463 , \21819 );
nor \U$22816 ( \23160 , \23158 , \23159 );
xnor \U$22817 ( \23161 , \23160 , \21727 );
and \U$22818 ( \23162 , \21750 , \21652 );
and \U$22819 ( \23163 , \21689 , \21650 );
nor \U$22820 ( \23164 , \23162 , \23163 );
xnor \U$22821 ( \23165 , \23164 , \21377 );
and \U$22822 ( \23166 , \23161 , \23165 );
and \U$22823 ( \23167 , \22011 , \21385 );
and \U$22824 ( \23168 , \21813 , \21383 );
nor \U$22825 ( \23169 , \23167 , \23168 );
xnor \U$22826 ( \23170 , \23169 , \21392 );
and \U$22827 ( \23171 , \23165 , \23170 );
and \U$22828 ( \23172 , \23161 , \23170 );
or \U$22829 ( \23173 , \23166 , \23171 , \23172 );
and \U$22830 ( \23174 , \23156 , \23173 );
and \U$22831 ( \23175 , \23140 , \23173 );
or \U$22832 ( \23176 , \23157 , \23174 , \23175 );
and \U$22833 ( \23177 , \22204 , \21401 );
and \U$22834 ( \23178 , \22099 , \21399 );
nor \U$22835 ( \23179 , \23177 , \23178 );
xnor \U$22836 ( \23180 , \23179 , \21408 );
and \U$22837 ( \23181 , \22325 , \21419 );
and \U$22838 ( \23182 , \22209 , \21417 );
nor \U$22839 ( \23183 , \23181 , \23182 );
xnor \U$22840 ( \23184 , \23183 , \21426 );
and \U$22841 ( \23185 , \23180 , \23184 );
and \U$22842 ( \23186 , \22616 , \21434 );
and \U$22843 ( \23187 , \22440 , \21432 );
nor \U$22844 ( \23188 , \23186 , \23187 );
xnor \U$22845 ( \23189 , \23188 , \21441 );
and \U$22846 ( \23190 , \23184 , \23189 );
and \U$22847 ( \23191 , \23180 , \23189 );
or \U$22848 ( \23192 , \23185 , \23190 , \23191 );
and \U$22849 ( \23193 , \22867 , \21450 );
and \U$22850 ( \23194 , \22624 , \21448 );
nor \U$22851 ( \23195 , \23193 , \23194 );
xnor \U$22852 ( \23196 , \23195 , \21457 );
and \U$22853 ( \23197 , \23058 , \21469 );
and \U$22854 ( \23198 , \22872 , \21467 );
nor \U$22855 ( \23199 , \23197 , \23198 );
xnor \U$22856 ( \23200 , \23199 , \21476 );
and \U$22857 ( \23201 , \23196 , \23200 );
buf \U$22858 ( \23202 , RIbb32298_156);
and \U$22859 ( \23203 , \23202 , \21464 );
and \U$22860 ( \23204 , \23200 , \23203 );
and \U$22861 ( \23205 , \23196 , \23203 );
or \U$22862 ( \23206 , \23201 , \23204 , \23205 );
and \U$22863 ( \23207 , \23192 , \23206 );
xor \U$22864 ( \23208 , \23052 , \23056 );
xor \U$22865 ( \23209 , \23208 , \23059 );
and \U$22866 ( \23210 , \23206 , \23209 );
and \U$22867 ( \23211 , \23192 , \23209 );
or \U$22868 ( \23212 , \23207 , \23210 , \23211 );
and \U$22869 ( \23213 , \23176 , \23212 );
xor \U$22870 ( \23214 , \23005 , \23009 );
xor \U$22871 ( \23215 , \23214 , \23014 );
xor \U$22872 ( \23216 , \23066 , \23070 );
xor \U$22873 ( \23217 , \23216 , \23075 );
and \U$22874 ( \23218 , \23215 , \23217 );
xor \U$22875 ( \23219 , \23022 , \23026 );
xor \U$22876 ( \23220 , \23219 , \23031 );
and \U$22877 ( \23221 , \23217 , \23220 );
and \U$22878 ( \23222 , \23215 , \23220 );
or \U$22879 ( \23223 , \23218 , \23221 , \23222 );
and \U$22880 ( \23224 , \23212 , \23223 );
and \U$22881 ( \23225 , \23176 , \23223 );
or \U$22882 ( \23226 , \23213 , \23224 , \23225 );
xor \U$22883 ( \23227 , \22922 , \22926 );
xor \U$22884 ( \23228 , \23227 , \22931 );
xor \U$22885 ( \23229 , \23039 , \23041 );
xor \U$22886 ( \23230 , \23229 , \23044 );
and \U$22887 ( \23231 , \23228 , \23230 );
xor \U$22888 ( \23232 , \23062 , \23078 );
xor \U$22889 ( \23233 , \23232 , \23080 );
and \U$22890 ( \23234 , \23230 , \23233 );
and \U$22891 ( \23235 , \23228 , \23233 );
or \U$22892 ( \23236 , \23231 , \23234 , \23235 );
and \U$22893 ( \23237 , \23226 , \23236 );
xor \U$22894 ( \23238 , \22866 , \22874 );
xor \U$22895 ( \23239 , \23238 , \22879 );
and \U$22896 ( \23240 , \23236 , \23239 );
and \U$22897 ( \23241 , \23226 , \23239 );
or \U$22898 ( \23242 , \23237 , \23240 , \23241 );
xor \U$22899 ( \23243 , \22898 , \22914 );
xor \U$22900 ( \23244 , \23243 , \22934 );
xor \U$22901 ( \23245 , \23037 , \23047 );
xor \U$22902 ( \23246 , \23245 , \23083 );
and \U$22903 ( \23247 , \23244 , \23246 );
xor \U$22904 ( \23248 , \23088 , \23090 );
xor \U$22905 ( \23249 , \23248 , \23093 );
and \U$22906 ( \23250 , \23246 , \23249 );
and \U$22907 ( \23251 , \23244 , \23249 );
or \U$22908 ( \23252 , \23247 , \23250 , \23251 );
and \U$22909 ( \23253 , \23242 , \23252 );
xor \U$22910 ( \23254 , \22882 , \22937 );
xor \U$22911 ( \23255 , \23254 , \22947 );
and \U$22912 ( \23256 , \23252 , \23255 );
and \U$22913 ( \23257 , \23242 , \23255 );
or \U$22914 ( \23258 , \23253 , \23256 , \23257 );
and \U$22915 ( \23259 , \21413 , \22651 );
and \U$22916 ( \23260 , \21421 , \22649 );
nor \U$22917 ( \23261 , \23259 , \23260 );
xnor \U$22918 ( \23262 , \23261 , \22495 );
and \U$22919 ( \23263 , \21428 , \22379 );
and \U$22920 ( \23264 , \21436 , \22377 );
nor \U$22921 ( \23265 , \23263 , \23264 );
xnor \U$22922 ( \23266 , \23265 , \22266 );
and \U$22923 ( \23267 , \23262 , \23266 );
and \U$22924 ( \23268 , \21444 , \22185 );
and \U$22925 ( \23269 , \21452 , \22183 );
nor \U$22926 ( \23270 , \23268 , \23269 );
xnor \U$22927 ( \23271 , \23270 , \22049 );
and \U$22928 ( \23272 , \23266 , \23271 );
and \U$22929 ( \23273 , \23262 , \23271 );
or \U$22930 ( \23274 , \23267 , \23272 , \23273 );
buf \U$22931 ( \23275 , RIbb2e878_30);
buf \U$22932 ( \23276 , RIbb2e800_31);
and \U$22933 ( \23277 , \23275 , \23276 );
not \U$22934 ( \23278 , \23277 );
and \U$22935 ( \23279 , \22985 , \23278 );
not \U$22936 ( \23280 , \23279 );
and \U$22937 ( \23281 , \21379 , \23125 );
and \U$22938 ( \23282 , \21387 , \23123 );
nor \U$22939 ( \23283 , \23281 , \23282 );
xnor \U$22940 ( \23284 , \23283 , \22988 );
and \U$22941 ( \23285 , \23280 , \23284 );
and \U$22942 ( \23286 , \21395 , \22919 );
and \U$22943 ( \23287 , \21403 , \22917 );
nor \U$22944 ( \23288 , \23286 , \23287 );
xnor \U$22945 ( \23289 , \23288 , \22767 );
and \U$22946 ( \23290 , \23284 , \23289 );
and \U$22947 ( \23291 , \23280 , \23289 );
or \U$22948 ( \23292 , \23285 , \23290 , \23291 );
and \U$22949 ( \23293 , \23274 , \23292 );
and \U$22950 ( \23294 , \21463 , \21985 );
and \U$22951 ( \23295 , \21471 , \21983 );
nor \U$22952 ( \23296 , \23294 , \23295 );
xnor \U$22953 ( \23297 , \23296 , \21907 );
and \U$22954 ( \23298 , \21689 , \21821 );
and \U$22955 ( \23299 , \21478 , \21819 );
nor \U$22956 ( \23300 , \23298 , \23299 );
xnor \U$22957 ( \23301 , \23300 , \21727 );
and \U$22958 ( \23302 , \23297 , \23301 );
and \U$22959 ( \23303 , \21813 , \21652 );
and \U$22960 ( \23304 , \21750 , \21650 );
nor \U$22961 ( \23305 , \23303 , \23304 );
xnor \U$22962 ( \23306 , \23305 , \21377 );
and \U$22963 ( \23307 , \23301 , \23306 );
and \U$22964 ( \23308 , \23297 , \23306 );
or \U$22965 ( \23309 , \23302 , \23307 , \23308 );
and \U$22966 ( \23310 , \23292 , \23309 );
and \U$22967 ( \23311 , \23274 , \23309 );
or \U$22968 ( \23312 , \23293 , \23310 , \23311 );
xor \U$22969 ( \23313 , \23180 , \23184 );
xor \U$22970 ( \23314 , \23313 , \23189 );
xor \U$22971 ( \23315 , \23196 , \23200 );
xor \U$22972 ( \23316 , \23315 , \23203 );
and \U$22973 ( \23317 , \23314 , \23316 );
xor \U$22974 ( \23318 , \23161 , \23165 );
xor \U$22975 ( \23319 , \23318 , \23170 );
and \U$22976 ( \23320 , \23316 , \23319 );
and \U$22977 ( \23321 , \23314 , \23319 );
or \U$22978 ( \23322 , \23317 , \23320 , \23321 );
and \U$22979 ( \23323 , \23312 , \23322 );
and \U$22980 ( \23324 , \22624 , \21434 );
and \U$22981 ( \23325 , \22616 , \21432 );
nor \U$22982 ( \23326 , \23324 , \23325 );
xnor \U$22983 ( \23327 , \23326 , \21441 );
and \U$22984 ( \23328 , \22872 , \21450 );
and \U$22985 ( \23329 , \22867 , \21448 );
nor \U$22986 ( \23330 , \23328 , \23329 );
xnor \U$22987 ( \23331 , \23330 , \21457 );
and \U$22988 ( \23332 , \23327 , \23331 );
and \U$22989 ( \23333 , \23202 , \21469 );
and \U$22990 ( \23334 , \23058 , \21467 );
nor \U$22991 ( \23335 , \23333 , \23334 );
xnor \U$22992 ( \23336 , \23335 , \21476 );
and \U$22993 ( \23337 , \23331 , \23336 );
and \U$22994 ( \23338 , \23327 , \23336 );
or \U$22995 ( \23339 , \23332 , \23337 , \23338 );
and \U$22996 ( \23340 , \22099 , \21385 );
and \U$22997 ( \23341 , \22011 , \21383 );
nor \U$22998 ( \23342 , \23340 , \23341 );
xnor \U$22999 ( \23343 , \23342 , \21392 );
and \U$23000 ( \23344 , \22209 , \21401 );
and \U$23001 ( \23345 , \22204 , \21399 );
nor \U$23002 ( \23346 , \23344 , \23345 );
xnor \U$23003 ( \23347 , \23346 , \21408 );
and \U$23004 ( \23348 , \23343 , \23347 );
and \U$23005 ( \23349 , \22440 , \21419 );
and \U$23006 ( \23350 , \22325 , \21417 );
nor \U$23007 ( \23351 , \23349 , \23350 );
xnor \U$23008 ( \23352 , \23351 , \21426 );
and \U$23009 ( \23353 , \23347 , \23352 );
and \U$23010 ( \23354 , \23343 , \23352 );
or \U$23011 ( \23355 , \23348 , \23353 , \23354 );
or \U$23012 ( \23356 , \23339 , \23355 );
and \U$23013 ( \23357 , \23322 , \23356 );
and \U$23014 ( \23358 , \23312 , \23356 );
or \U$23015 ( \23359 , \23323 , \23357 , \23358 );
xor \U$23016 ( \23360 , \22989 , \22993 );
xor \U$23017 ( \23361 , \23360 , \22998 );
xor \U$23018 ( \23362 , \23192 , \23206 );
xor \U$23019 ( \23363 , \23362 , \23209 );
and \U$23020 ( \23364 , \23361 , \23363 );
xor \U$23021 ( \23365 , \23215 , \23217 );
xor \U$23022 ( \23366 , \23365 , \23220 );
and \U$23023 ( \23367 , \23363 , \23366 );
and \U$23024 ( \23368 , \23361 , \23366 );
or \U$23025 ( \23369 , \23364 , \23367 , \23368 );
and \U$23026 ( \23370 , \23359 , \23369 );
xor \U$23027 ( \23371 , \23001 , \23017 );
xor \U$23028 ( \23372 , \23371 , \23034 );
and \U$23029 ( \23373 , \23369 , \23372 );
and \U$23030 ( \23374 , \23359 , \23372 );
or \U$23031 ( \23375 , \23370 , \23373 , \23374 );
xor \U$23032 ( \23376 , \23226 , \23236 );
xor \U$23033 ( \23377 , \23376 , \23239 );
and \U$23034 ( \23378 , \23375 , \23377 );
xor \U$23035 ( \23379 , \23244 , \23246 );
xor \U$23036 ( \23380 , \23379 , \23249 );
and \U$23037 ( \23381 , \23377 , \23380 );
and \U$23038 ( \23382 , \23375 , \23380 );
or \U$23039 ( \23383 , \23378 , \23381 , \23382 );
xor \U$23040 ( \23384 , \23242 , \23252 );
xor \U$23041 ( \23385 , \23384 , \23255 );
and \U$23042 ( \23386 , \23383 , \23385 );
xor \U$23043 ( \23387 , \23086 , \23096 );
xor \U$23044 ( \23388 , \23387 , \23099 );
and \U$23045 ( \23389 , \23385 , \23388 );
and \U$23046 ( \23390 , \23383 , \23388 );
or \U$23047 ( \23391 , \23386 , \23389 , \23390 );
and \U$23048 ( \23392 , \23258 , \23391 );
xor \U$23049 ( \23393 , \23102 , \23104 );
xor \U$23050 ( \23394 , \23393 , \23106 );
and \U$23051 ( \23395 , \23391 , \23394 );
and \U$23052 ( \23396 , \23258 , \23394 );
or \U$23053 ( \23397 , \23392 , \23395 , \23396 );
and \U$23054 ( \23398 , \23121 , \23397 );
xor \U$23055 ( \23399 , \23121 , \23397 );
xor \U$23056 ( \23400 , \23258 , \23391 );
xor \U$23057 ( \23401 , \23400 , \23394 );
and \U$23058 ( \23402 , \21436 , \22651 );
and \U$23059 ( \23403 , \21413 , \22649 );
nor \U$23060 ( \23404 , \23402 , \23403 );
xnor \U$23061 ( \23405 , \23404 , \22495 );
and \U$23062 ( \23406 , \21452 , \22379 );
and \U$23063 ( \23407 , \21428 , \22377 );
nor \U$23064 ( \23408 , \23406 , \23407 );
xnor \U$23065 ( \23409 , \23408 , \22266 );
and \U$23066 ( \23410 , \23405 , \23409 );
and \U$23067 ( \23411 , \21471 , \22185 );
and \U$23068 ( \23412 , \21444 , \22183 );
nor \U$23069 ( \23413 , \23411 , \23412 );
xnor \U$23070 ( \23414 , \23413 , \22049 );
and \U$23071 ( \23415 , \23409 , \23414 );
and \U$23072 ( \23416 , \23405 , \23414 );
or \U$23073 ( \23417 , \23410 , \23415 , \23416 );
xor \U$23074 ( \23418 , \22985 , \23275 );
xor \U$23075 ( \23419 , \23275 , \23276 );
not \U$23076 ( \23420 , \23419 );
and \U$23077 ( \23421 , \23418 , \23420 );
and \U$23078 ( \23422 , \21387 , \23421 );
not \U$23079 ( \23423 , \23422 );
xnor \U$23080 ( \23424 , \23423 , \23279 );
and \U$23081 ( \23425 , \21403 , \23125 );
and \U$23082 ( \23426 , \21379 , \23123 );
nor \U$23083 ( \23427 , \23425 , \23426 );
xnor \U$23084 ( \23428 , \23427 , \22988 );
and \U$23085 ( \23429 , \23424 , \23428 );
and \U$23086 ( \23430 , \21421 , \22919 );
and \U$23087 ( \23431 , \21395 , \22917 );
nor \U$23088 ( \23432 , \23430 , \23431 );
xnor \U$23089 ( \23433 , \23432 , \22767 );
and \U$23090 ( \23434 , \23428 , \23433 );
and \U$23091 ( \23435 , \23424 , \23433 );
or \U$23092 ( \23436 , \23429 , \23434 , \23435 );
and \U$23093 ( \23437 , \23417 , \23436 );
and \U$23094 ( \23438 , \21478 , \21985 );
and \U$23095 ( \23439 , \21463 , \21983 );
nor \U$23096 ( \23440 , \23438 , \23439 );
xnor \U$23097 ( \23441 , \23440 , \21907 );
and \U$23098 ( \23442 , \21750 , \21821 );
and \U$23099 ( \23443 , \21689 , \21819 );
nor \U$23100 ( \23444 , \23442 , \23443 );
xnor \U$23101 ( \23445 , \23444 , \21727 );
and \U$23102 ( \23446 , \23441 , \23445 );
and \U$23103 ( \23447 , \22011 , \21652 );
and \U$23104 ( \23448 , \21813 , \21650 );
nor \U$23105 ( \23449 , \23447 , \23448 );
xnor \U$23106 ( \23450 , \23449 , \21377 );
and \U$23107 ( \23451 , \23445 , \23450 );
and \U$23108 ( \23452 , \23441 , \23450 );
or \U$23109 ( \23453 , \23446 , \23451 , \23452 );
and \U$23110 ( \23454 , \23436 , \23453 );
and \U$23111 ( \23455 , \23417 , \23453 );
or \U$23112 ( \23456 , \23437 , \23454 , \23455 );
and \U$23113 ( \23457 , \22867 , \21434 );
and \U$23114 ( \23458 , \22624 , \21432 );
nor \U$23115 ( \23459 , \23457 , \23458 );
xnor \U$23116 ( \23460 , \23459 , \21441 );
and \U$23117 ( \23461 , \23058 , \21450 );
and \U$23118 ( \23462 , \22872 , \21448 );
nor \U$23119 ( \23463 , \23461 , \23462 );
xnor \U$23120 ( \23464 , \23463 , \21457 );
and \U$23121 ( \23465 , \23460 , \23464 );
buf \U$23122 ( \23466 , RIbb32310_157);
and \U$23123 ( \23467 , \23466 , \21469 );
and \U$23124 ( \23468 , \23202 , \21467 );
nor \U$23125 ( \23469 , \23467 , \23468 );
xnor \U$23126 ( \23470 , \23469 , \21476 );
and \U$23127 ( \23471 , \23464 , \23470 );
and \U$23128 ( \23472 , \23460 , \23470 );
or \U$23129 ( \23473 , \23465 , \23471 , \23472 );
and \U$23130 ( \23474 , \22204 , \21385 );
and \U$23131 ( \23475 , \22099 , \21383 );
nor \U$23132 ( \23476 , \23474 , \23475 );
xnor \U$23133 ( \23477 , \23476 , \21392 );
and \U$23134 ( \23478 , \22325 , \21401 );
and \U$23135 ( \23479 , \22209 , \21399 );
nor \U$23136 ( \23480 , \23478 , \23479 );
xnor \U$23137 ( \23481 , \23480 , \21408 );
and \U$23138 ( \23482 , \23477 , \23481 );
and \U$23139 ( \23483 , \22616 , \21419 );
and \U$23140 ( \23484 , \22440 , \21417 );
nor \U$23141 ( \23485 , \23483 , \23484 );
xnor \U$23142 ( \23486 , \23485 , \21426 );
and \U$23143 ( \23487 , \23481 , \23486 );
and \U$23144 ( \23488 , \23477 , \23486 );
or \U$23145 ( \23489 , \23482 , \23487 , \23488 );
and \U$23146 ( \23490 , \23473 , \23489 );
buf \U$23147 ( \23491 , RIbb32388_158);
and \U$23148 ( \23492 , \23491 , \21464 );
buf \U$23149 ( \23493 , \23492 );
and \U$23150 ( \23494 , \23489 , \23493 );
and \U$23151 ( \23495 , \23473 , \23493 );
or \U$23152 ( \23496 , \23490 , \23494 , \23495 );
and \U$23153 ( \23497 , \23456 , \23496 );
and \U$23154 ( \23498 , \23466 , \21464 );
xor \U$23155 ( \23499 , \23327 , \23331 );
xor \U$23156 ( \23500 , \23499 , \23336 );
and \U$23157 ( \23501 , \23498 , \23500 );
xor \U$23158 ( \23502 , \23343 , \23347 );
xor \U$23159 ( \23503 , \23502 , \23352 );
and \U$23160 ( \23504 , \23500 , \23503 );
and \U$23161 ( \23505 , \23498 , \23503 );
or \U$23162 ( \23506 , \23501 , \23504 , \23505 );
and \U$23163 ( \23507 , \23496 , \23506 );
and \U$23164 ( \23508 , \23456 , \23506 );
or \U$23165 ( \23509 , \23497 , \23507 , \23508 );
xor \U$23166 ( \23510 , \23262 , \23266 );
xor \U$23167 ( \23511 , \23510 , \23271 );
xor \U$23168 ( \23512 , \23280 , \23284 );
xor \U$23169 ( \23513 , \23512 , \23289 );
and \U$23170 ( \23514 , \23511 , \23513 );
xor \U$23171 ( \23515 , \23297 , \23301 );
xor \U$23172 ( \23516 , \23515 , \23306 );
and \U$23173 ( \23517 , \23513 , \23516 );
and \U$23174 ( \23518 , \23511 , \23516 );
or \U$23175 ( \23519 , \23514 , \23517 , \23518 );
xor \U$23176 ( \23520 , \23128 , \23132 );
xor \U$23177 ( \23521 , \23520 , \23137 );
and \U$23178 ( \23522 , \23519 , \23521 );
xor \U$23179 ( \23523 , \23144 , \23148 );
xor \U$23180 ( \23524 , \23523 , \23153 );
and \U$23181 ( \23525 , \23521 , \23524 );
and \U$23182 ( \23526 , \23519 , \23524 );
or \U$23183 ( \23527 , \23522 , \23525 , \23526 );
and \U$23184 ( \23528 , \23509 , \23527 );
xor \U$23185 ( \23529 , \23274 , \23292 );
xor \U$23186 ( \23530 , \23529 , \23309 );
xor \U$23187 ( \23531 , \23314 , \23316 );
xor \U$23188 ( \23532 , \23531 , \23319 );
and \U$23189 ( \23533 , \23530 , \23532 );
xnor \U$23190 ( \23534 , \23339 , \23355 );
and \U$23191 ( \23535 , \23532 , \23534 );
and \U$23192 ( \23536 , \23530 , \23534 );
or \U$23193 ( \23537 , \23533 , \23535 , \23536 );
and \U$23194 ( \23538 , \23527 , \23537 );
and \U$23195 ( \23539 , \23509 , \23537 );
or \U$23196 ( \23540 , \23528 , \23538 , \23539 );
xor \U$23197 ( \23541 , \23140 , \23156 );
xor \U$23198 ( \23542 , \23541 , \23173 );
xor \U$23199 ( \23543 , \23312 , \23322 );
xor \U$23200 ( \23544 , \23543 , \23356 );
and \U$23201 ( \23545 , \23542 , \23544 );
xor \U$23202 ( \23546 , \23361 , \23363 );
xor \U$23203 ( \23547 , \23546 , \23366 );
and \U$23204 ( \23548 , \23544 , \23547 );
and \U$23205 ( \23549 , \23542 , \23547 );
or \U$23206 ( \23550 , \23545 , \23548 , \23549 );
and \U$23207 ( \23551 , \23540 , \23550 );
xor \U$23208 ( \23552 , \23228 , \23230 );
xor \U$23209 ( \23553 , \23552 , \23233 );
and \U$23210 ( \23554 , \23550 , \23553 );
and \U$23211 ( \23555 , \23540 , \23553 );
or \U$23212 ( \23556 , \23551 , \23554 , \23555 );
xor \U$23213 ( \23557 , \23176 , \23212 );
xor \U$23214 ( \23558 , \23557 , \23223 );
xor \U$23215 ( \23559 , \23359 , \23369 );
xor \U$23216 ( \23560 , \23559 , \23372 );
and \U$23217 ( \23561 , \23558 , \23560 );
and \U$23218 ( \23562 , \23556 , \23561 );
xor \U$23219 ( \23563 , \23375 , \23377 );
xor \U$23220 ( \23564 , \23563 , \23380 );
and \U$23221 ( \23565 , \23561 , \23564 );
and \U$23222 ( \23566 , \23556 , \23564 );
or \U$23223 ( \23567 , \23562 , \23565 , \23566 );
xor \U$23224 ( \23568 , \23383 , \23385 );
xor \U$23225 ( \23569 , \23568 , \23388 );
and \U$23226 ( \23570 , \23567 , \23569 );
and \U$23227 ( \23571 , \23401 , \23570 );
xor \U$23228 ( \23572 , \23401 , \23570 );
xor \U$23229 ( \23573 , \23567 , \23569 );
and \U$23230 ( \23574 , \21463 , \22185 );
and \U$23231 ( \23575 , \21471 , \22183 );
nor \U$23232 ( \23576 , \23574 , \23575 );
xnor \U$23233 ( \23577 , \23576 , \22049 );
and \U$23234 ( \23578 , \21689 , \21985 );
and \U$23235 ( \23579 , \21478 , \21983 );
nor \U$23236 ( \23580 , \23578 , \23579 );
xnor \U$23237 ( \23581 , \23580 , \21907 );
and \U$23238 ( \23582 , \23577 , \23581 );
and \U$23239 ( \23583 , \21813 , \21821 );
and \U$23240 ( \23584 , \21750 , \21819 );
nor \U$23241 ( \23585 , \23583 , \23584 );
xnor \U$23242 ( \23586 , \23585 , \21727 );
and \U$23243 ( \23587 , \23581 , \23586 );
and \U$23244 ( \23588 , \23577 , \23586 );
or \U$23245 ( \23589 , \23582 , \23587 , \23588 );
buf \U$23246 ( \23590 , RIbb2e788_32);
buf \U$23247 ( \23591 , RIbb2e710_33);
and \U$23248 ( \23592 , \23590 , \23591 );
not \U$23249 ( \23593 , \23592 );
and \U$23250 ( \23594 , \23276 , \23593 );
not \U$23251 ( \23595 , \23594 );
and \U$23252 ( \23596 , \21379 , \23421 );
and \U$23253 ( \23597 , \21387 , \23419 );
nor \U$23254 ( \23598 , \23596 , \23597 );
xnor \U$23255 ( \23599 , \23598 , \23279 );
and \U$23256 ( \23600 , \23595 , \23599 );
and \U$23257 ( \23601 , \21395 , \23125 );
and \U$23258 ( \23602 , \21403 , \23123 );
nor \U$23259 ( \23603 , \23601 , \23602 );
xnor \U$23260 ( \23604 , \23603 , \22988 );
and \U$23261 ( \23605 , \23599 , \23604 );
and \U$23262 ( \23606 , \23595 , \23604 );
or \U$23263 ( \23607 , \23600 , \23605 , \23606 );
and \U$23264 ( \23608 , \23589 , \23607 );
and \U$23265 ( \23609 , \21413 , \22919 );
and \U$23266 ( \23610 , \21421 , \22917 );
nor \U$23267 ( \23611 , \23609 , \23610 );
xnor \U$23268 ( \23612 , \23611 , \22767 );
and \U$23269 ( \23613 , \21428 , \22651 );
and \U$23270 ( \23614 , \21436 , \22649 );
nor \U$23271 ( \23615 , \23613 , \23614 );
xnor \U$23272 ( \23616 , \23615 , \22495 );
and \U$23273 ( \23617 , \23612 , \23616 );
and \U$23274 ( \23618 , \21444 , \22379 );
and \U$23275 ( \23619 , \21452 , \22377 );
nor \U$23276 ( \23620 , \23618 , \23619 );
xnor \U$23277 ( \23621 , \23620 , \22266 );
and \U$23278 ( \23622 , \23616 , \23621 );
and \U$23279 ( \23623 , \23612 , \23621 );
or \U$23280 ( \23624 , \23617 , \23622 , \23623 );
and \U$23281 ( \23625 , \23607 , \23624 );
and \U$23282 ( \23626 , \23589 , \23624 );
or \U$23283 ( \23627 , \23608 , \23625 , \23626 );
and \U$23284 ( \23628 , \22624 , \21419 );
and \U$23285 ( \23629 , \22616 , \21417 );
nor \U$23286 ( \23630 , \23628 , \23629 );
xnor \U$23287 ( \23631 , \23630 , \21426 );
and \U$23288 ( \23632 , \22872 , \21434 );
and \U$23289 ( \23633 , \22867 , \21432 );
nor \U$23290 ( \23634 , \23632 , \23633 );
xnor \U$23291 ( \23635 , \23634 , \21441 );
and \U$23292 ( \23636 , \23631 , \23635 );
and \U$23293 ( \23637 , \23202 , \21450 );
and \U$23294 ( \23638 , \23058 , \21448 );
nor \U$23295 ( \23639 , \23637 , \23638 );
xnor \U$23296 ( \23640 , \23639 , \21457 );
and \U$23297 ( \23641 , \23635 , \23640 );
and \U$23298 ( \23642 , \23631 , \23640 );
or \U$23299 ( \23643 , \23636 , \23641 , \23642 );
and \U$23300 ( \23644 , \22099 , \21652 );
and \U$23301 ( \23645 , \22011 , \21650 );
nor \U$23302 ( \23646 , \23644 , \23645 );
xnor \U$23303 ( \23647 , \23646 , \21377 );
and \U$23304 ( \23648 , \22209 , \21385 );
and \U$23305 ( \23649 , \22204 , \21383 );
nor \U$23306 ( \23650 , \23648 , \23649 );
xnor \U$23307 ( \23651 , \23650 , \21392 );
and \U$23308 ( \23652 , \23647 , \23651 );
and \U$23309 ( \23653 , \22440 , \21401 );
and \U$23310 ( \23654 , \22325 , \21399 );
nor \U$23311 ( \23655 , \23653 , \23654 );
xnor \U$23312 ( \23656 , \23655 , \21408 );
and \U$23313 ( \23657 , \23651 , \23656 );
and \U$23314 ( \23658 , \23647 , \23656 );
or \U$23315 ( \23659 , \23652 , \23657 , \23658 );
and \U$23316 ( \23660 , \23643 , \23659 );
and \U$23317 ( \23661 , \23491 , \21469 );
and \U$23318 ( \23662 , \23466 , \21467 );
nor \U$23319 ( \23663 , \23661 , \23662 );
xnor \U$23320 ( \23664 , \23663 , \21476 );
buf \U$23321 ( \23665 , RIbb32400_159);
and \U$23322 ( \23666 , \23665 , \21464 );
and \U$23323 ( \23667 , \23664 , \23666 );
and \U$23324 ( \23668 , \23659 , \23667 );
and \U$23325 ( \23669 , \23643 , \23667 );
or \U$23326 ( \23670 , \23660 , \23668 , \23669 );
and \U$23327 ( \23671 , \23627 , \23670 );
xor \U$23328 ( \23672 , \23460 , \23464 );
xor \U$23329 ( \23673 , \23672 , \23470 );
xor \U$23330 ( \23674 , \23477 , \23481 );
xor \U$23331 ( \23675 , \23674 , \23486 );
and \U$23332 ( \23676 , \23673 , \23675 );
not \U$23333 ( \23677 , \23492 );
and \U$23334 ( \23678 , \23675 , \23677 );
and \U$23335 ( \23679 , \23673 , \23677 );
or \U$23336 ( \23680 , \23676 , \23678 , \23679 );
and \U$23337 ( \23681 , \23670 , \23680 );
and \U$23338 ( \23682 , \23627 , \23680 );
or \U$23339 ( \23683 , \23671 , \23681 , \23682 );
xor \U$23340 ( \23684 , \23405 , \23409 );
xor \U$23341 ( \23685 , \23684 , \23414 );
xor \U$23342 ( \23686 , \23424 , \23428 );
xor \U$23343 ( \23687 , \23686 , \23433 );
and \U$23344 ( \23688 , \23685 , \23687 );
xor \U$23345 ( \23689 , \23441 , \23445 );
xor \U$23346 ( \23690 , \23689 , \23450 );
and \U$23347 ( \23691 , \23687 , \23690 );
and \U$23348 ( \23692 , \23685 , \23690 );
or \U$23349 ( \23693 , \23688 , \23691 , \23692 );
xor \U$23350 ( \23694 , \23511 , \23513 );
xor \U$23351 ( \23695 , \23694 , \23516 );
and \U$23352 ( \23696 , \23693 , \23695 );
xor \U$23353 ( \23697 , \23498 , \23500 );
xor \U$23354 ( \23698 , \23697 , \23503 );
and \U$23355 ( \23699 , \23695 , \23698 );
and \U$23356 ( \23700 , \23693 , \23698 );
or \U$23357 ( \23701 , \23696 , \23699 , \23700 );
and \U$23358 ( \23702 , \23683 , \23701 );
xor \U$23359 ( \23703 , \23417 , \23436 );
xor \U$23360 ( \23704 , \23703 , \23453 );
xor \U$23361 ( \23705 , \23473 , \23489 );
xor \U$23362 ( \23706 , \23705 , \23493 );
and \U$23363 ( \23707 , \23704 , \23706 );
and \U$23364 ( \23708 , \23701 , \23707 );
and \U$23365 ( \23709 , \23683 , \23707 );
or \U$23366 ( \23710 , \23702 , \23708 , \23709 );
xor \U$23367 ( \23711 , \23456 , \23496 );
xor \U$23368 ( \23712 , \23711 , \23506 );
xor \U$23369 ( \23713 , \23519 , \23521 );
xor \U$23370 ( \23714 , \23713 , \23524 );
and \U$23371 ( \23715 , \23712 , \23714 );
xor \U$23372 ( \23716 , \23530 , \23532 );
xor \U$23373 ( \23717 , \23716 , \23534 );
and \U$23374 ( \23718 , \23714 , \23717 );
and \U$23375 ( \23719 , \23712 , \23717 );
or \U$23376 ( \23720 , \23715 , \23718 , \23719 );
and \U$23377 ( \23721 , \23710 , \23720 );
xor \U$23378 ( \23722 , \23542 , \23544 );
xor \U$23379 ( \23723 , \23722 , \23547 );
and \U$23380 ( \23724 , \23720 , \23723 );
and \U$23381 ( \23725 , \23710 , \23723 );
or \U$23382 ( \23726 , \23721 , \23724 , \23725 );
xor \U$23383 ( \23727 , \23540 , \23550 );
xor \U$23384 ( \23728 , \23727 , \23553 );
and \U$23385 ( \23729 , \23726 , \23728 );
xor \U$23386 ( \23730 , \23558 , \23560 );
and \U$23387 ( \23731 , \23728 , \23730 );
and \U$23388 ( \23732 , \23726 , \23730 );
or \U$23389 ( \23733 , \23729 , \23731 , \23732 );
xor \U$23390 ( \23734 , \23556 , \23561 );
xor \U$23391 ( \23735 , \23734 , \23564 );
and \U$23392 ( \23736 , \23733 , \23735 );
and \U$23393 ( \23737 , \23573 , \23736 );
xor \U$23394 ( \23738 , \23573 , \23736 );
xor \U$23395 ( \23739 , \23733 , \23735 );
xor \U$23396 ( \23740 , \23276 , \23590 );
xor \U$23397 ( \23741 , \23590 , \23591 );
not \U$23398 ( \23742 , \23741 );
and \U$23399 ( \23743 , \23740 , \23742 );
and \U$23400 ( \23744 , \21387 , \23743 );
not \U$23401 ( \23745 , \23744 );
xnor \U$23402 ( \23746 , \23745 , \23594 );
and \U$23403 ( \23747 , \21403 , \23421 );
and \U$23404 ( \23748 , \21379 , \23419 );
nor \U$23405 ( \23749 , \23747 , \23748 );
xnor \U$23406 ( \23750 , \23749 , \23279 );
and \U$23407 ( \23751 , \23746 , \23750 );
and \U$23408 ( \23752 , \21421 , \23125 );
and \U$23409 ( \23753 , \21395 , \23123 );
nor \U$23410 ( \23754 , \23752 , \23753 );
xnor \U$23411 ( \23755 , \23754 , \22988 );
and \U$23412 ( \23756 , \23750 , \23755 );
and \U$23413 ( \23757 , \23746 , \23755 );
or \U$23414 ( \23758 , \23751 , \23756 , \23757 );
and \U$23415 ( \23759 , \21478 , \22185 );
and \U$23416 ( \23760 , \21463 , \22183 );
nor \U$23417 ( \23761 , \23759 , \23760 );
xnor \U$23418 ( \23762 , \23761 , \22049 );
and \U$23419 ( \23763 , \21750 , \21985 );
and \U$23420 ( \23764 , \21689 , \21983 );
nor \U$23421 ( \23765 , \23763 , \23764 );
xnor \U$23422 ( \23766 , \23765 , \21907 );
and \U$23423 ( \23767 , \23762 , \23766 );
and \U$23424 ( \23768 , \22011 , \21821 );
and \U$23425 ( \23769 , \21813 , \21819 );
nor \U$23426 ( \23770 , \23768 , \23769 );
xnor \U$23427 ( \23771 , \23770 , \21727 );
and \U$23428 ( \23772 , \23766 , \23771 );
and \U$23429 ( \23773 , \23762 , \23771 );
or \U$23430 ( \23774 , \23767 , \23772 , \23773 );
and \U$23431 ( \23775 , \23758 , \23774 );
and \U$23432 ( \23776 , \21436 , \22919 );
and \U$23433 ( \23777 , \21413 , \22917 );
nor \U$23434 ( \23778 , \23776 , \23777 );
xnor \U$23435 ( \23779 , \23778 , \22767 );
and \U$23436 ( \23780 , \21452 , \22651 );
and \U$23437 ( \23781 , \21428 , \22649 );
nor \U$23438 ( \23782 , \23780 , \23781 );
xnor \U$23439 ( \23783 , \23782 , \22495 );
and \U$23440 ( \23784 , \23779 , \23783 );
and \U$23441 ( \23785 , \21471 , \22379 );
and \U$23442 ( \23786 , \21444 , \22377 );
nor \U$23443 ( \23787 , \23785 , \23786 );
xnor \U$23444 ( \23788 , \23787 , \22266 );
and \U$23445 ( \23789 , \23783 , \23788 );
and \U$23446 ( \23790 , \23779 , \23788 );
or \U$23447 ( \23791 , \23784 , \23789 , \23790 );
and \U$23448 ( \23792 , \23774 , \23791 );
and \U$23449 ( \23793 , \23758 , \23791 );
or \U$23450 ( \23794 , \23775 , \23792 , \23793 );
and \U$23451 ( \23795 , \22867 , \21419 );
and \U$23452 ( \23796 , \22624 , \21417 );
nor \U$23453 ( \23797 , \23795 , \23796 );
xnor \U$23454 ( \23798 , \23797 , \21426 );
and \U$23455 ( \23799 , \23058 , \21434 );
and \U$23456 ( \23800 , \22872 , \21432 );
nor \U$23457 ( \23801 , \23799 , \23800 );
xnor \U$23458 ( \23802 , \23801 , \21441 );
and \U$23459 ( \23803 , \23798 , \23802 );
and \U$23460 ( \23804 , \23466 , \21450 );
and \U$23461 ( \23805 , \23202 , \21448 );
nor \U$23462 ( \23806 , \23804 , \23805 );
xnor \U$23463 ( \23807 , \23806 , \21457 );
and \U$23464 ( \23808 , \23802 , \23807 );
and \U$23465 ( \23809 , \23798 , \23807 );
or \U$23466 ( \23810 , \23803 , \23808 , \23809 );
and \U$23467 ( \23811 , \22204 , \21652 );
and \U$23468 ( \23812 , \22099 , \21650 );
nor \U$23469 ( \23813 , \23811 , \23812 );
xnor \U$23470 ( \23814 , \23813 , \21377 );
and \U$23471 ( \23815 , \22325 , \21385 );
and \U$23472 ( \23816 , \22209 , \21383 );
nor \U$23473 ( \23817 , \23815 , \23816 );
xnor \U$23474 ( \23818 , \23817 , \21392 );
and \U$23475 ( \23819 , \23814 , \23818 );
and \U$23476 ( \23820 , \22616 , \21401 );
and \U$23477 ( \23821 , \22440 , \21399 );
nor \U$23478 ( \23822 , \23820 , \23821 );
xnor \U$23479 ( \23823 , \23822 , \21408 );
and \U$23480 ( \23824 , \23818 , \23823 );
and \U$23481 ( \23825 , \23814 , \23823 );
or \U$23482 ( \23826 , \23819 , \23824 , \23825 );
and \U$23483 ( \23827 , \23810 , \23826 );
and \U$23484 ( \23828 , \23665 , \21469 );
and \U$23485 ( \23829 , \23491 , \21467 );
nor \U$23486 ( \23830 , \23828 , \23829 );
xnor \U$23487 ( \23831 , \23830 , \21476 );
buf \U$23488 ( \23832 , RIbb32478_160);
and \U$23489 ( \23833 , \23832 , \21464 );
or \U$23490 ( \23834 , \23831 , \23833 );
and \U$23491 ( \23835 , \23826 , \23834 );
and \U$23492 ( \23836 , \23810 , \23834 );
or \U$23493 ( \23837 , \23827 , \23835 , \23836 );
and \U$23494 ( \23838 , \23794 , \23837 );
xor \U$23495 ( \23839 , \23631 , \23635 );
xor \U$23496 ( \23840 , \23839 , \23640 );
xor \U$23497 ( \23841 , \23647 , \23651 );
xor \U$23498 ( \23842 , \23841 , \23656 );
and \U$23499 ( \23843 , \23840 , \23842 );
xor \U$23500 ( \23844 , \23664 , \23666 );
and \U$23501 ( \23845 , \23842 , \23844 );
and \U$23502 ( \23846 , \23840 , \23844 );
or \U$23503 ( \23847 , \23843 , \23845 , \23846 );
and \U$23504 ( \23848 , \23837 , \23847 );
and \U$23505 ( \23849 , \23794 , \23847 );
or \U$23506 ( \23850 , \23838 , \23848 , \23849 );
xor \U$23507 ( \23851 , \23577 , \23581 );
xor \U$23508 ( \23852 , \23851 , \23586 );
xor \U$23509 ( \23853 , \23595 , \23599 );
xor \U$23510 ( \23854 , \23853 , \23604 );
and \U$23511 ( \23855 , \23852 , \23854 );
xor \U$23512 ( \23856 , \23612 , \23616 );
xor \U$23513 ( \23857 , \23856 , \23621 );
and \U$23514 ( \23858 , \23854 , \23857 );
and \U$23515 ( \23859 , \23852 , \23857 );
or \U$23516 ( \23860 , \23855 , \23858 , \23859 );
xor \U$23517 ( \23861 , \23685 , \23687 );
xor \U$23518 ( \23862 , \23861 , \23690 );
and \U$23519 ( \23863 , \23860 , \23862 );
xor \U$23520 ( \23864 , \23673 , \23675 );
xor \U$23521 ( \23865 , \23864 , \23677 );
and \U$23522 ( \23866 , \23862 , \23865 );
and \U$23523 ( \23867 , \23860 , \23865 );
or \U$23524 ( \23868 , \23863 , \23866 , \23867 );
and \U$23525 ( \23869 , \23850 , \23868 );
xor \U$23526 ( \23870 , \23589 , \23607 );
xor \U$23527 ( \23871 , \23870 , \23624 );
xor \U$23528 ( \23872 , \23643 , \23659 );
xor \U$23529 ( \23873 , \23872 , \23667 );
and \U$23530 ( \23874 , \23871 , \23873 );
and \U$23531 ( \23875 , \23868 , \23874 );
and \U$23532 ( \23876 , \23850 , \23874 );
or \U$23533 ( \23877 , \23869 , \23875 , \23876 );
xor \U$23534 ( \23878 , \23627 , \23670 );
xor \U$23535 ( \23879 , \23878 , \23680 );
xor \U$23536 ( \23880 , \23693 , \23695 );
xor \U$23537 ( \23881 , \23880 , \23698 );
and \U$23538 ( \23882 , \23879 , \23881 );
xor \U$23539 ( \23883 , \23704 , \23706 );
and \U$23540 ( \23884 , \23881 , \23883 );
and \U$23541 ( \23885 , \23879 , \23883 );
or \U$23542 ( \23886 , \23882 , \23884 , \23885 );
and \U$23543 ( \23887 , \23877 , \23886 );
xor \U$23544 ( \23888 , \23712 , \23714 );
xor \U$23545 ( \23889 , \23888 , \23717 );
and \U$23546 ( \23890 , \23886 , \23889 );
and \U$23547 ( \23891 , \23877 , \23889 );
or \U$23548 ( \23892 , \23887 , \23890 , \23891 );
xor \U$23549 ( \23893 , \23509 , \23527 );
xor \U$23550 ( \23894 , \23893 , \23537 );
and \U$23551 ( \23895 , \23892 , \23894 );
xor \U$23552 ( \23896 , \23710 , \23720 );
xor \U$23553 ( \23897 , \23896 , \23723 );
and \U$23554 ( \23898 , \23894 , \23897 );
and \U$23555 ( \23899 , \23892 , \23897 );
or \U$23556 ( \23900 , \23895 , \23898 , \23899 );
xor \U$23557 ( \23901 , \23726 , \23728 );
xor \U$23558 ( \23902 , \23901 , \23730 );
and \U$23559 ( \23903 , \23900 , \23902 );
and \U$23560 ( \23904 , \23739 , \23903 );
xor \U$23561 ( \23905 , \23739 , \23903 );
xor \U$23562 ( \23906 , \23900 , \23902 );
and \U$23563 ( \23907 , \21413 , \23125 );
and \U$23564 ( \23908 , \21421 , \23123 );
nor \U$23565 ( \23909 , \23907 , \23908 );
xnor \U$23566 ( \23910 , \23909 , \22988 );
and \U$23567 ( \23911 , \21428 , \22919 );
and \U$23568 ( \23912 , \21436 , \22917 );
nor \U$23569 ( \23913 , \23911 , \23912 );
xnor \U$23570 ( \23914 , \23913 , \22767 );
and \U$23571 ( \23915 , \23910 , \23914 );
and \U$23572 ( \23916 , \21444 , \22651 );
and \U$23573 ( \23917 , \21452 , \22649 );
nor \U$23574 ( \23918 , \23916 , \23917 );
xnor \U$23575 ( \23919 , \23918 , \22495 );
and \U$23576 ( \23920 , \23914 , \23919 );
and \U$23577 ( \23921 , \23910 , \23919 );
or \U$23578 ( \23922 , \23915 , \23920 , \23921 );
and \U$23579 ( \23923 , \21463 , \22379 );
and \U$23580 ( \23924 , \21471 , \22377 );
nor \U$23581 ( \23925 , \23923 , \23924 );
xnor \U$23582 ( \23926 , \23925 , \22266 );
and \U$23583 ( \23927 , \21689 , \22185 );
and \U$23584 ( \23928 , \21478 , \22183 );
nor \U$23585 ( \23929 , \23927 , \23928 );
xnor \U$23586 ( \23930 , \23929 , \22049 );
and \U$23587 ( \23931 , \23926 , \23930 );
and \U$23588 ( \23932 , \21813 , \21985 );
and \U$23589 ( \23933 , \21750 , \21983 );
nor \U$23590 ( \23934 , \23932 , \23933 );
xnor \U$23591 ( \23935 , \23934 , \21907 );
and \U$23592 ( \23936 , \23930 , \23935 );
and \U$23593 ( \23937 , \23926 , \23935 );
or \U$23594 ( \23938 , \23931 , \23936 , \23937 );
and \U$23595 ( \23939 , \23922 , \23938 );
buf \U$23596 ( \23940 , RIbb2e698_34);
buf \U$23597 ( \23941 , RIbb2e620_35);
and \U$23598 ( \23942 , \23940 , \23941 );
not \U$23599 ( \23943 , \23942 );
and \U$23600 ( \23944 , \23591 , \23943 );
not \U$23601 ( \23945 , \23944 );
and \U$23602 ( \23946 , \21379 , \23743 );
and \U$23603 ( \23947 , \21387 , \23741 );
nor \U$23604 ( \23948 , \23946 , \23947 );
xnor \U$23605 ( \23949 , \23948 , \23594 );
and \U$23606 ( \23950 , \23945 , \23949 );
and \U$23607 ( \23951 , \21395 , \23421 );
and \U$23608 ( \23952 , \21403 , \23419 );
nor \U$23609 ( \23953 , \23951 , \23952 );
xnor \U$23610 ( \23954 , \23953 , \23279 );
and \U$23611 ( \23955 , \23949 , \23954 );
and \U$23612 ( \23956 , \23945 , \23954 );
or \U$23613 ( \23957 , \23950 , \23955 , \23956 );
and \U$23614 ( \23958 , \23938 , \23957 );
and \U$23615 ( \23959 , \23922 , \23957 );
or \U$23616 ( \23960 , \23939 , \23958 , \23959 );
and \U$23617 ( \23961 , \23491 , \21450 );
and \U$23618 ( \23962 , \23466 , \21448 );
nor \U$23619 ( \23963 , \23961 , \23962 );
xnor \U$23620 ( \23964 , \23963 , \21457 );
and \U$23621 ( \23965 , \23832 , \21469 );
and \U$23622 ( \23966 , \23665 , \21467 );
nor \U$23623 ( \23967 , \23965 , \23966 );
xnor \U$23624 ( \23968 , \23967 , \21476 );
and \U$23625 ( \23969 , \23964 , \23968 );
buf \U$23626 ( \23970 , RIbb324f0_161);
and \U$23627 ( \23971 , \23970 , \21464 );
and \U$23628 ( \23972 , \23968 , \23971 );
and \U$23629 ( \23973 , \23964 , \23971 );
or \U$23630 ( \23974 , \23969 , \23972 , \23973 );
and \U$23631 ( \23975 , \22624 , \21401 );
and \U$23632 ( \23976 , \22616 , \21399 );
nor \U$23633 ( \23977 , \23975 , \23976 );
xnor \U$23634 ( \23978 , \23977 , \21408 );
and \U$23635 ( \23979 , \22872 , \21419 );
and \U$23636 ( \23980 , \22867 , \21417 );
nor \U$23637 ( \23981 , \23979 , \23980 );
xnor \U$23638 ( \23982 , \23981 , \21426 );
and \U$23639 ( \23983 , \23978 , \23982 );
and \U$23640 ( \23984 , \23202 , \21434 );
and \U$23641 ( \23985 , \23058 , \21432 );
nor \U$23642 ( \23986 , \23984 , \23985 );
xnor \U$23643 ( \23987 , \23986 , \21441 );
and \U$23644 ( \23988 , \23982 , \23987 );
and \U$23645 ( \23989 , \23978 , \23987 );
or \U$23646 ( \23990 , \23983 , \23988 , \23989 );
and \U$23647 ( \23991 , \23974 , \23990 );
and \U$23648 ( \23992 , \22099 , \21821 );
and \U$23649 ( \23993 , \22011 , \21819 );
nor \U$23650 ( \23994 , \23992 , \23993 );
xnor \U$23651 ( \23995 , \23994 , \21727 );
and \U$23652 ( \23996 , \22209 , \21652 );
and \U$23653 ( \23997 , \22204 , \21650 );
nor \U$23654 ( \23998 , \23996 , \23997 );
xnor \U$23655 ( \23999 , \23998 , \21377 );
and \U$23656 ( \24000 , \23995 , \23999 );
and \U$23657 ( \24001 , \22440 , \21385 );
and \U$23658 ( \24002 , \22325 , \21383 );
nor \U$23659 ( \24003 , \24001 , \24002 );
xnor \U$23660 ( \24004 , \24003 , \21392 );
and \U$23661 ( \24005 , \23999 , \24004 );
and \U$23662 ( \24006 , \23995 , \24004 );
or \U$23663 ( \24007 , \24000 , \24005 , \24006 );
and \U$23664 ( \24008 , \23990 , \24007 );
and \U$23665 ( \24009 , \23974 , \24007 );
or \U$23666 ( \24010 , \23991 , \24008 , \24009 );
and \U$23667 ( \24011 , \23960 , \24010 );
xor \U$23668 ( \24012 , \23798 , \23802 );
xor \U$23669 ( \24013 , \24012 , \23807 );
xor \U$23670 ( \24014 , \23814 , \23818 );
xor \U$23671 ( \24015 , \24014 , \23823 );
and \U$23672 ( \24016 , \24013 , \24015 );
xnor \U$23673 ( \24017 , \23831 , \23833 );
and \U$23674 ( \24018 , \24015 , \24017 );
and \U$23675 ( \24019 , \24013 , \24017 );
or \U$23676 ( \24020 , \24016 , \24018 , \24019 );
and \U$23677 ( \24021 , \24010 , \24020 );
and \U$23678 ( \24022 , \23960 , \24020 );
or \U$23679 ( \24023 , \24011 , \24021 , \24022 );
xor \U$23680 ( \24024 , \23746 , \23750 );
xor \U$23681 ( \24025 , \24024 , \23755 );
xor \U$23682 ( \24026 , \23762 , \23766 );
xor \U$23683 ( \24027 , \24026 , \23771 );
and \U$23684 ( \24028 , \24025 , \24027 );
xor \U$23685 ( \24029 , \23779 , \23783 );
xor \U$23686 ( \24030 , \24029 , \23788 );
and \U$23687 ( \24031 , \24027 , \24030 );
and \U$23688 ( \24032 , \24025 , \24030 );
or \U$23689 ( \24033 , \24028 , \24031 , \24032 );
xor \U$23690 ( \24034 , \23852 , \23854 );
xor \U$23691 ( \24035 , \24034 , \23857 );
and \U$23692 ( \24036 , \24033 , \24035 );
xor \U$23693 ( \24037 , \23840 , \23842 );
xor \U$23694 ( \24038 , \24037 , \23844 );
and \U$23695 ( \24039 , \24035 , \24038 );
and \U$23696 ( \24040 , \24033 , \24038 );
or \U$23697 ( \24041 , \24036 , \24039 , \24040 );
and \U$23698 ( \24042 , \24023 , \24041 );
xor \U$23699 ( \24043 , \23758 , \23774 );
xor \U$23700 ( \24044 , \24043 , \23791 );
xor \U$23701 ( \24045 , \23810 , \23826 );
xor \U$23702 ( \24046 , \24045 , \23834 );
and \U$23703 ( \24047 , \24044 , \24046 );
and \U$23704 ( \24048 , \24041 , \24047 );
and \U$23705 ( \24049 , \24023 , \24047 );
or \U$23706 ( \24050 , \24042 , \24048 , \24049 );
xor \U$23707 ( \24051 , \23794 , \23837 );
xor \U$23708 ( \24052 , \24051 , \23847 );
xor \U$23709 ( \24053 , \23860 , \23862 );
xor \U$23710 ( \24054 , \24053 , \23865 );
and \U$23711 ( \24055 , \24052 , \24054 );
xor \U$23712 ( \24056 , \23871 , \23873 );
and \U$23713 ( \24057 , \24054 , \24056 );
and \U$23714 ( \24058 , \24052 , \24056 );
or \U$23715 ( \24059 , \24055 , \24057 , \24058 );
and \U$23716 ( \24060 , \24050 , \24059 );
xor \U$23717 ( \24061 , \23879 , \23881 );
xor \U$23718 ( \24062 , \24061 , \23883 );
and \U$23719 ( \24063 , \24059 , \24062 );
and \U$23720 ( \24064 , \24050 , \24062 );
or \U$23721 ( \24065 , \24060 , \24063 , \24064 );
xor \U$23722 ( \24066 , \23683 , \23701 );
xor \U$23723 ( \24067 , \24066 , \23707 );
and \U$23724 ( \24068 , \24065 , \24067 );
xor \U$23725 ( \24069 , \23877 , \23886 );
xor \U$23726 ( \24070 , \24069 , \23889 );
and \U$23727 ( \24071 , \24067 , \24070 );
and \U$23728 ( \24072 , \24065 , \24070 );
or \U$23729 ( \24073 , \24068 , \24071 , \24072 );
xor \U$23730 ( \24074 , \23892 , \23894 );
xor \U$23731 ( \24075 , \24074 , \23897 );
and \U$23732 ( \24076 , \24073 , \24075 );
and \U$23733 ( \24077 , \23906 , \24076 );
xor \U$23734 ( \24078 , \23906 , \24076 );
xor \U$23735 ( \24079 , \24073 , \24075 );
and \U$23736 ( \24080 , \23665 , \21450 );
and \U$23737 ( \24081 , \23491 , \21448 );
nor \U$23738 ( \24082 , \24080 , \24081 );
xnor \U$23739 ( \24083 , \24082 , \21457 );
and \U$23740 ( \24084 , \23970 , \21469 );
and \U$23741 ( \24085 , \23832 , \21467 );
nor \U$23742 ( \24086 , \24084 , \24085 );
xnor \U$23743 ( \24087 , \24086 , \21476 );
and \U$23744 ( \24088 , \24083 , \24087 );
buf \U$23745 ( \24089 , RIbb32568_162);
and \U$23746 ( \24090 , \24089 , \21464 );
and \U$23747 ( \24091 , \24087 , \24090 );
and \U$23748 ( \24092 , \24083 , \24090 );
or \U$23749 ( \24093 , \24088 , \24091 , \24092 );
and \U$23750 ( \24094 , \22867 , \21401 );
and \U$23751 ( \24095 , \22624 , \21399 );
nor \U$23752 ( \24096 , \24094 , \24095 );
xnor \U$23753 ( \24097 , \24096 , \21408 );
and \U$23754 ( \24098 , \23058 , \21419 );
and \U$23755 ( \24099 , \22872 , \21417 );
nor \U$23756 ( \24100 , \24098 , \24099 );
xnor \U$23757 ( \24101 , \24100 , \21426 );
and \U$23758 ( \24102 , \24097 , \24101 );
and \U$23759 ( \24103 , \23466 , \21434 );
and \U$23760 ( \24104 , \23202 , \21432 );
nor \U$23761 ( \24105 , \24103 , \24104 );
xnor \U$23762 ( \24106 , \24105 , \21441 );
and \U$23763 ( \24107 , \24101 , \24106 );
and \U$23764 ( \24108 , \24097 , \24106 );
or \U$23765 ( \24109 , \24102 , \24107 , \24108 );
and \U$23766 ( \24110 , \24093 , \24109 );
and \U$23767 ( \24111 , \22204 , \21821 );
and \U$23768 ( \24112 , \22099 , \21819 );
nor \U$23769 ( \24113 , \24111 , \24112 );
xnor \U$23770 ( \24114 , \24113 , \21727 );
and \U$23771 ( \24115 , \22325 , \21652 );
and \U$23772 ( \24116 , \22209 , \21650 );
nor \U$23773 ( \24117 , \24115 , \24116 );
xnor \U$23774 ( \24118 , \24117 , \21377 );
and \U$23775 ( \24119 , \24114 , \24118 );
and \U$23776 ( \24120 , \22616 , \21385 );
and \U$23777 ( \24121 , \22440 , \21383 );
nor \U$23778 ( \24122 , \24120 , \24121 );
xnor \U$23779 ( \24123 , \24122 , \21392 );
and \U$23780 ( \24124 , \24118 , \24123 );
and \U$23781 ( \24125 , \24114 , \24123 );
or \U$23782 ( \24126 , \24119 , \24124 , \24125 );
and \U$23783 ( \24127 , \24109 , \24126 );
and \U$23784 ( \24128 , \24093 , \24126 );
or \U$23785 ( \24129 , \24110 , \24127 , \24128 );
and \U$23786 ( \24130 , \21436 , \23125 );
and \U$23787 ( \24131 , \21413 , \23123 );
nor \U$23788 ( \24132 , \24130 , \24131 );
xnor \U$23789 ( \24133 , \24132 , \22988 );
and \U$23790 ( \24134 , \21452 , \22919 );
and \U$23791 ( \24135 , \21428 , \22917 );
nor \U$23792 ( \24136 , \24134 , \24135 );
xnor \U$23793 ( \24137 , \24136 , \22767 );
and \U$23794 ( \24138 , \24133 , \24137 );
and \U$23795 ( \24139 , \21471 , \22651 );
and \U$23796 ( \24140 , \21444 , \22649 );
nor \U$23797 ( \24141 , \24139 , \24140 );
xnor \U$23798 ( \24142 , \24141 , \22495 );
and \U$23799 ( \24143 , \24137 , \24142 );
and \U$23800 ( \24144 , \24133 , \24142 );
or \U$23801 ( \24145 , \24138 , \24143 , \24144 );
xor \U$23802 ( \24146 , \23591 , \23940 );
xor \U$23803 ( \24147 , \23940 , \23941 );
not \U$23804 ( \24148 , \24147 );
and \U$23805 ( \24149 , \24146 , \24148 );
and \U$23806 ( \24150 , \21387 , \24149 );
not \U$23807 ( \24151 , \24150 );
xnor \U$23808 ( \24152 , \24151 , \23944 );
and \U$23809 ( \24153 , \21403 , \23743 );
and \U$23810 ( \24154 , \21379 , \23741 );
nor \U$23811 ( \24155 , \24153 , \24154 );
xnor \U$23812 ( \24156 , \24155 , \23594 );
and \U$23813 ( \24157 , \24152 , \24156 );
and \U$23814 ( \24158 , \21421 , \23421 );
and \U$23815 ( \24159 , \21395 , \23419 );
nor \U$23816 ( \24160 , \24158 , \24159 );
xnor \U$23817 ( \24161 , \24160 , \23279 );
and \U$23818 ( \24162 , \24156 , \24161 );
and \U$23819 ( \24163 , \24152 , \24161 );
or \U$23820 ( \24164 , \24157 , \24162 , \24163 );
and \U$23821 ( \24165 , \24145 , \24164 );
and \U$23822 ( \24166 , \21478 , \22379 );
and \U$23823 ( \24167 , \21463 , \22377 );
nor \U$23824 ( \24168 , \24166 , \24167 );
xnor \U$23825 ( \24169 , \24168 , \22266 );
and \U$23826 ( \24170 , \21750 , \22185 );
and \U$23827 ( \24171 , \21689 , \22183 );
nor \U$23828 ( \24172 , \24170 , \24171 );
xnor \U$23829 ( \24173 , \24172 , \22049 );
and \U$23830 ( \24174 , \24169 , \24173 );
and \U$23831 ( \24175 , \22011 , \21985 );
and \U$23832 ( \24176 , \21813 , \21983 );
nor \U$23833 ( \24177 , \24175 , \24176 );
xnor \U$23834 ( \24178 , \24177 , \21907 );
and \U$23835 ( \24179 , \24173 , \24178 );
and \U$23836 ( \24180 , \24169 , \24178 );
or \U$23837 ( \24181 , \24174 , \24179 , \24180 );
and \U$23838 ( \24182 , \24164 , \24181 );
and \U$23839 ( \24183 , \24145 , \24181 );
or \U$23840 ( \24184 , \24165 , \24182 , \24183 );
and \U$23841 ( \24185 , \24129 , \24184 );
xor \U$23842 ( \24186 , \23964 , \23968 );
xor \U$23843 ( \24187 , \24186 , \23971 );
xor \U$23844 ( \24188 , \23978 , \23982 );
xor \U$23845 ( \24189 , \24188 , \23987 );
and \U$23846 ( \24190 , \24187 , \24189 );
xor \U$23847 ( \24191 , \23995 , \23999 );
xor \U$23848 ( \24192 , \24191 , \24004 );
and \U$23849 ( \24193 , \24189 , \24192 );
and \U$23850 ( \24194 , \24187 , \24192 );
or \U$23851 ( \24195 , \24190 , \24193 , \24194 );
and \U$23852 ( \24196 , \24184 , \24195 );
and \U$23853 ( \24197 , \24129 , \24195 );
or \U$23854 ( \24198 , \24185 , \24196 , \24197 );
xor \U$23855 ( \24199 , \23910 , \23914 );
xor \U$23856 ( \24200 , \24199 , \23919 );
xor \U$23857 ( \24201 , \23926 , \23930 );
xor \U$23858 ( \24202 , \24201 , \23935 );
and \U$23859 ( \24203 , \24200 , \24202 );
xor \U$23860 ( \24204 , \23945 , \23949 );
xor \U$23861 ( \24205 , \24204 , \23954 );
and \U$23862 ( \24206 , \24202 , \24205 );
and \U$23863 ( \24207 , \24200 , \24205 );
or \U$23864 ( \24208 , \24203 , \24206 , \24207 );
xor \U$23865 ( \24209 , \24025 , \24027 );
xor \U$23866 ( \24210 , \24209 , \24030 );
and \U$23867 ( \24211 , \24208 , \24210 );
xor \U$23868 ( \24212 , \24013 , \24015 );
xor \U$23869 ( \24213 , \24212 , \24017 );
and \U$23870 ( \24214 , \24210 , \24213 );
and \U$23871 ( \24215 , \24208 , \24213 );
or \U$23872 ( \24216 , \24211 , \24214 , \24215 );
and \U$23873 ( \24217 , \24198 , \24216 );
xor \U$23874 ( \24218 , \23922 , \23938 );
xor \U$23875 ( \24219 , \24218 , \23957 );
xor \U$23876 ( \24220 , \23974 , \23990 );
xor \U$23877 ( \24221 , \24220 , \24007 );
and \U$23878 ( \24222 , \24219 , \24221 );
and \U$23879 ( \24223 , \24216 , \24222 );
and \U$23880 ( \24224 , \24198 , \24222 );
or \U$23881 ( \24225 , \24217 , \24223 , \24224 );
xor \U$23882 ( \24226 , \23960 , \24010 );
xor \U$23883 ( \24227 , \24226 , \24020 );
xor \U$23884 ( \24228 , \24033 , \24035 );
xor \U$23885 ( \24229 , \24228 , \24038 );
and \U$23886 ( \24230 , \24227 , \24229 );
xor \U$23887 ( \24231 , \24044 , \24046 );
and \U$23888 ( \24232 , \24229 , \24231 );
and \U$23889 ( \24233 , \24227 , \24231 );
or \U$23890 ( \24234 , \24230 , \24232 , \24233 );
and \U$23891 ( \24235 , \24225 , \24234 );
xor \U$23892 ( \24236 , \24052 , \24054 );
xor \U$23893 ( \24237 , \24236 , \24056 );
and \U$23894 ( \24238 , \24234 , \24237 );
and \U$23895 ( \24239 , \24225 , \24237 );
or \U$23896 ( \24240 , \24235 , \24238 , \24239 );
xor \U$23897 ( \24241 , \23850 , \23868 );
xor \U$23898 ( \24242 , \24241 , \23874 );
and \U$23899 ( \24243 , \24240 , \24242 );
xor \U$23900 ( \24244 , \24050 , \24059 );
xor \U$23901 ( \24245 , \24244 , \24062 );
and \U$23902 ( \24246 , \24242 , \24245 );
and \U$23903 ( \24247 , \24240 , \24245 );
or \U$23904 ( \24248 , \24243 , \24246 , \24247 );
xor \U$23905 ( \24249 , \24065 , \24067 );
xor \U$23906 ( \24250 , \24249 , \24070 );
and \U$23907 ( \24251 , \24248 , \24250 );
and \U$23908 ( \24252 , \24079 , \24251 );
xor \U$23909 ( \24253 , \24079 , \24251 );
xor \U$23910 ( \24254 , \24248 , \24250 );
and \U$23911 ( \24255 , \21463 , \22651 );
and \U$23912 ( \24256 , \21471 , \22649 );
nor \U$23913 ( \24257 , \24255 , \24256 );
xnor \U$23914 ( \24258 , \24257 , \22495 );
and \U$23915 ( \24259 , \21689 , \22379 );
and \U$23916 ( \24260 , \21478 , \22377 );
nor \U$23917 ( \24261 , \24259 , \24260 );
xnor \U$23918 ( \24262 , \24261 , \22266 );
and \U$23919 ( \24263 , \24258 , \24262 );
and \U$23920 ( \24264 , \21813 , \22185 );
and \U$23921 ( \24265 , \21750 , \22183 );
nor \U$23922 ( \24266 , \24264 , \24265 );
xnor \U$23923 ( \24267 , \24266 , \22049 );
and \U$23924 ( \24268 , \24262 , \24267 );
and \U$23925 ( \24269 , \24258 , \24267 );
or \U$23926 ( \24270 , \24263 , \24268 , \24269 );
buf \U$23927 ( \24271 , RIbb2e5a8_36);
buf \U$23928 ( \24272 , RIbb2e530_37);
and \U$23929 ( \24273 , \24271 , \24272 );
not \U$23930 ( \24274 , \24273 );
and \U$23931 ( \24275 , \23941 , \24274 );
not \U$23932 ( \24276 , \24275 );
and \U$23933 ( \24277 , \21379 , \24149 );
and \U$23934 ( \24278 , \21387 , \24147 );
nor \U$23935 ( \24279 , \24277 , \24278 );
xnor \U$23936 ( \24280 , \24279 , \23944 );
and \U$23937 ( \24281 , \24276 , \24280 );
and \U$23938 ( \24282 , \21395 , \23743 );
and \U$23939 ( \24283 , \21403 , \23741 );
nor \U$23940 ( \24284 , \24282 , \24283 );
xnor \U$23941 ( \24285 , \24284 , \23594 );
and \U$23942 ( \24286 , \24280 , \24285 );
and \U$23943 ( \24287 , \24276 , \24285 );
or \U$23944 ( \24288 , \24281 , \24286 , \24287 );
and \U$23945 ( \24289 , \24270 , \24288 );
and \U$23946 ( \24290 , \21413 , \23421 );
and \U$23947 ( \24291 , \21421 , \23419 );
nor \U$23948 ( \24292 , \24290 , \24291 );
xnor \U$23949 ( \24293 , \24292 , \23279 );
and \U$23950 ( \24294 , \21428 , \23125 );
and \U$23951 ( \24295 , \21436 , \23123 );
nor \U$23952 ( \24296 , \24294 , \24295 );
xnor \U$23953 ( \24297 , \24296 , \22988 );
and \U$23954 ( \24298 , \24293 , \24297 );
and \U$23955 ( \24299 , \21444 , \22919 );
and \U$23956 ( \24300 , \21452 , \22917 );
nor \U$23957 ( \24301 , \24299 , \24300 );
xnor \U$23958 ( \24302 , \24301 , \22767 );
and \U$23959 ( \24303 , \24297 , \24302 );
and \U$23960 ( \24304 , \24293 , \24302 );
or \U$23961 ( \24305 , \24298 , \24303 , \24304 );
and \U$23962 ( \24306 , \24288 , \24305 );
and \U$23963 ( \24307 , \24270 , \24305 );
or \U$23964 ( \24308 , \24289 , \24306 , \24307 );
and \U$23965 ( \24309 , \23491 , \21434 );
and \U$23966 ( \24310 , \23466 , \21432 );
nor \U$23967 ( \24311 , \24309 , \24310 );
xnor \U$23968 ( \24312 , \24311 , \21441 );
and \U$23969 ( \24313 , \23832 , \21450 );
and \U$23970 ( \24314 , \23665 , \21448 );
nor \U$23971 ( \24315 , \24313 , \24314 );
xnor \U$23972 ( \24316 , \24315 , \21457 );
and \U$23973 ( \24317 , \24312 , \24316 );
and \U$23974 ( \24318 , \24089 , \21469 );
and \U$23975 ( \24319 , \23970 , \21467 );
nor \U$23976 ( \24320 , \24318 , \24319 );
xnor \U$23977 ( \24321 , \24320 , \21476 );
and \U$23978 ( \24322 , \24316 , \24321 );
and \U$23979 ( \24323 , \24312 , \24321 );
or \U$23980 ( \24324 , \24317 , \24322 , \24323 );
and \U$23981 ( \24325 , \22099 , \21985 );
and \U$23982 ( \24326 , \22011 , \21983 );
nor \U$23983 ( \24327 , \24325 , \24326 );
xnor \U$23984 ( \24328 , \24327 , \21907 );
and \U$23985 ( \24329 , \22209 , \21821 );
and \U$23986 ( \24330 , \22204 , \21819 );
nor \U$23987 ( \24331 , \24329 , \24330 );
xnor \U$23988 ( \24332 , \24331 , \21727 );
and \U$23989 ( \24333 , \24328 , \24332 );
and \U$23990 ( \24334 , \22440 , \21652 );
and \U$23991 ( \24335 , \22325 , \21650 );
nor \U$23992 ( \24336 , \24334 , \24335 );
xnor \U$23993 ( \24337 , \24336 , \21377 );
and \U$23994 ( \24338 , \24332 , \24337 );
and \U$23995 ( \24339 , \24328 , \24337 );
or \U$23996 ( \24340 , \24333 , \24338 , \24339 );
and \U$23997 ( \24341 , \24324 , \24340 );
and \U$23998 ( \24342 , \22624 , \21385 );
and \U$23999 ( \24343 , \22616 , \21383 );
nor \U$24000 ( \24344 , \24342 , \24343 );
xnor \U$24001 ( \24345 , \24344 , \21392 );
and \U$24002 ( \24346 , \22872 , \21401 );
and \U$24003 ( \24347 , \22867 , \21399 );
nor \U$24004 ( \24348 , \24346 , \24347 );
xnor \U$24005 ( \24349 , \24348 , \21408 );
and \U$24006 ( \24350 , \24345 , \24349 );
and \U$24007 ( \24351 , \23202 , \21419 );
and \U$24008 ( \24352 , \23058 , \21417 );
nor \U$24009 ( \24353 , \24351 , \24352 );
xnor \U$24010 ( \24354 , \24353 , \21426 );
and \U$24011 ( \24355 , \24349 , \24354 );
and \U$24012 ( \24356 , \24345 , \24354 );
or \U$24013 ( \24357 , \24350 , \24355 , \24356 );
and \U$24014 ( \24358 , \24340 , \24357 );
and \U$24015 ( \24359 , \24324 , \24357 );
or \U$24016 ( \24360 , \24341 , \24358 , \24359 );
and \U$24017 ( \24361 , \24308 , \24360 );
xor \U$24018 ( \24362 , \24083 , \24087 );
xor \U$24019 ( \24363 , \24362 , \24090 );
xor \U$24020 ( \24364 , \24097 , \24101 );
xor \U$24021 ( \24365 , \24364 , \24106 );
or \U$24022 ( \24366 , \24363 , \24365 );
and \U$24023 ( \24367 , \24360 , \24366 );
and \U$24024 ( \24368 , \24308 , \24366 );
or \U$24025 ( \24369 , \24361 , \24367 , \24368 );
xor \U$24026 ( \24370 , \24133 , \24137 );
xor \U$24027 ( \24371 , \24370 , \24142 );
xor \U$24028 ( \24372 , \24169 , \24173 );
xor \U$24029 ( \24373 , \24372 , \24178 );
and \U$24030 ( \24374 , \24371 , \24373 );
xor \U$24031 ( \24375 , \24114 , \24118 );
xor \U$24032 ( \24376 , \24375 , \24123 );
and \U$24033 ( \24377 , \24373 , \24376 );
and \U$24034 ( \24378 , \24371 , \24376 );
or \U$24035 ( \24379 , \24374 , \24377 , \24378 );
xor \U$24036 ( \24380 , \24187 , \24189 );
xor \U$24037 ( \24381 , \24380 , \24192 );
and \U$24038 ( \24382 , \24379 , \24381 );
xor \U$24039 ( \24383 , \24200 , \24202 );
xor \U$24040 ( \24384 , \24383 , \24205 );
and \U$24041 ( \24385 , \24381 , \24384 );
and \U$24042 ( \24386 , \24379 , \24384 );
or \U$24043 ( \24387 , \24382 , \24385 , \24386 );
and \U$24044 ( \24388 , \24369 , \24387 );
xor \U$24045 ( \24389 , \24093 , \24109 );
xor \U$24046 ( \24390 , \24389 , \24126 );
xor \U$24047 ( \24391 , \24145 , \24164 );
xor \U$24048 ( \24392 , \24391 , \24181 );
and \U$24049 ( \24393 , \24390 , \24392 );
and \U$24050 ( \24394 , \24387 , \24393 );
and \U$24051 ( \24395 , \24369 , \24393 );
or \U$24052 ( \24396 , \24388 , \24394 , \24395 );
xor \U$24053 ( \24397 , \24129 , \24184 );
xor \U$24054 ( \24398 , \24397 , \24195 );
xor \U$24055 ( \24399 , \24208 , \24210 );
xor \U$24056 ( \24400 , \24399 , \24213 );
and \U$24057 ( \24401 , \24398 , \24400 );
xor \U$24058 ( \24402 , \24219 , \24221 );
and \U$24059 ( \24403 , \24400 , \24402 );
and \U$24060 ( \24404 , \24398 , \24402 );
or \U$24061 ( \24405 , \24401 , \24403 , \24404 );
and \U$24062 ( \24406 , \24396 , \24405 );
xor \U$24063 ( \24407 , \24227 , \24229 );
xor \U$24064 ( \24408 , \24407 , \24231 );
and \U$24065 ( \24409 , \24405 , \24408 );
and \U$24066 ( \24410 , \24396 , \24408 );
or \U$24067 ( \24411 , \24406 , \24409 , \24410 );
xor \U$24068 ( \24412 , \24023 , \24041 );
xor \U$24069 ( \24413 , \24412 , \24047 );
and \U$24070 ( \24414 , \24411 , \24413 );
xor \U$24071 ( \24415 , \24225 , \24234 );
xor \U$24072 ( \24416 , \24415 , \24237 );
and \U$24073 ( \24417 , \24413 , \24416 );
and \U$24074 ( \24418 , \24411 , \24416 );
or \U$24075 ( \24419 , \24414 , \24417 , \24418 );
xor \U$24076 ( \24420 , \24240 , \24242 );
xor \U$24077 ( \24421 , \24420 , \24245 );
and \U$24078 ( \24422 , \24419 , \24421 );
and \U$24079 ( \24423 , \24254 , \24422 );
xor \U$24080 ( \24424 , \24254 , \24422 );
xor \U$24081 ( \24425 , \24419 , \24421 );
and \U$24082 ( \24426 , \21478 , \22651 );
and \U$24083 ( \24427 , \21463 , \22649 );
nor \U$24084 ( \24428 , \24426 , \24427 );
xnor \U$24085 ( \24429 , \24428 , \22495 );
and \U$24086 ( \24430 , \21750 , \22379 );
and \U$24087 ( \24431 , \21689 , \22377 );
nor \U$24088 ( \24432 , \24430 , \24431 );
xnor \U$24089 ( \24433 , \24432 , \22266 );
and \U$24090 ( \24434 , \24429 , \24433 );
and \U$24091 ( \24435 , \22011 , \22185 );
and \U$24092 ( \24436 , \21813 , \22183 );
nor \U$24093 ( \24437 , \24435 , \24436 );
xnor \U$24094 ( \24438 , \24437 , \22049 );
and \U$24095 ( \24439 , \24433 , \24438 );
and \U$24096 ( \24440 , \24429 , \24438 );
or \U$24097 ( \24441 , \24434 , \24439 , \24440 );
and \U$24098 ( \24442 , \21436 , \23421 );
and \U$24099 ( \24443 , \21413 , \23419 );
nor \U$24100 ( \24444 , \24442 , \24443 );
xnor \U$24101 ( \24445 , \24444 , \23279 );
and \U$24102 ( \24446 , \21452 , \23125 );
and \U$24103 ( \24447 , \21428 , \23123 );
nor \U$24104 ( \24448 , \24446 , \24447 );
xnor \U$24105 ( \24449 , \24448 , \22988 );
and \U$24106 ( \24450 , \24445 , \24449 );
and \U$24107 ( \24451 , \21471 , \22919 );
and \U$24108 ( \24452 , \21444 , \22917 );
nor \U$24109 ( \24453 , \24451 , \24452 );
xnor \U$24110 ( \24454 , \24453 , \22767 );
and \U$24111 ( \24455 , \24449 , \24454 );
and \U$24112 ( \24456 , \24445 , \24454 );
or \U$24113 ( \24457 , \24450 , \24455 , \24456 );
and \U$24114 ( \24458 , \24441 , \24457 );
xor \U$24115 ( \24459 , \23941 , \24271 );
xor \U$24116 ( \24460 , \24271 , \24272 );
not \U$24117 ( \24461 , \24460 );
and \U$24118 ( \24462 , \24459 , \24461 );
and \U$24119 ( \24463 , \21387 , \24462 );
not \U$24120 ( \24464 , \24463 );
xnor \U$24121 ( \24465 , \24464 , \24275 );
and \U$24122 ( \24466 , \21403 , \24149 );
and \U$24123 ( \24467 , \21379 , \24147 );
nor \U$24124 ( \24468 , \24466 , \24467 );
xnor \U$24125 ( \24469 , \24468 , \23944 );
and \U$24126 ( \24470 , \24465 , \24469 );
and \U$24127 ( \24471 , \21421 , \23743 );
and \U$24128 ( \24472 , \21395 , \23741 );
nor \U$24129 ( \24473 , \24471 , \24472 );
xnor \U$24130 ( \24474 , \24473 , \23594 );
and \U$24131 ( \24475 , \24469 , \24474 );
and \U$24132 ( \24476 , \24465 , \24474 );
or \U$24133 ( \24477 , \24470 , \24475 , \24476 );
and \U$24134 ( \24478 , \24457 , \24477 );
and \U$24135 ( \24479 , \24441 , \24477 );
or \U$24136 ( \24480 , \24458 , \24478 , \24479 );
and \U$24137 ( \24481 , \22204 , \21985 );
and \U$24138 ( \24482 , \22099 , \21983 );
nor \U$24139 ( \24483 , \24481 , \24482 );
xnor \U$24140 ( \24484 , \24483 , \21907 );
and \U$24141 ( \24485 , \22325 , \21821 );
and \U$24142 ( \24486 , \22209 , \21819 );
nor \U$24143 ( \24487 , \24485 , \24486 );
xnor \U$24144 ( \24488 , \24487 , \21727 );
and \U$24145 ( \24489 , \24484 , \24488 );
and \U$24146 ( \24490 , \22616 , \21652 );
and \U$24147 ( \24491 , \22440 , \21650 );
nor \U$24148 ( \24492 , \24490 , \24491 );
xnor \U$24149 ( \24493 , \24492 , \21377 );
and \U$24150 ( \24494 , \24488 , \24493 );
and \U$24151 ( \24495 , \24484 , \24493 );
or \U$24152 ( \24496 , \24489 , \24494 , \24495 );
and \U$24153 ( \24497 , \23665 , \21434 );
and \U$24154 ( \24498 , \23491 , \21432 );
nor \U$24155 ( \24499 , \24497 , \24498 );
xnor \U$24156 ( \24500 , \24499 , \21441 );
and \U$24157 ( \24501 , \23970 , \21450 );
and \U$24158 ( \24502 , \23832 , \21448 );
nor \U$24159 ( \24503 , \24501 , \24502 );
xnor \U$24160 ( \24504 , \24503 , \21457 );
and \U$24161 ( \24505 , \24500 , \24504 );
buf \U$24162 ( \24506 , RIbb325e0_163);
and \U$24163 ( \24507 , \24506 , \21469 );
and \U$24164 ( \24508 , \24089 , \21467 );
nor \U$24165 ( \24509 , \24507 , \24508 );
xnor \U$24166 ( \24510 , \24509 , \21476 );
and \U$24167 ( \24511 , \24504 , \24510 );
and \U$24168 ( \24512 , \24500 , \24510 );
or \U$24169 ( \24513 , \24505 , \24511 , \24512 );
and \U$24170 ( \24514 , \24496 , \24513 );
and \U$24171 ( \24515 , \22867 , \21385 );
and \U$24172 ( \24516 , \22624 , \21383 );
nor \U$24173 ( \24517 , \24515 , \24516 );
xnor \U$24174 ( \24518 , \24517 , \21392 );
and \U$24175 ( \24519 , \23058 , \21401 );
and \U$24176 ( \24520 , \22872 , \21399 );
nor \U$24177 ( \24521 , \24519 , \24520 );
xnor \U$24178 ( \24522 , \24521 , \21408 );
and \U$24179 ( \24523 , \24518 , \24522 );
and \U$24180 ( \24524 , \23466 , \21419 );
and \U$24181 ( \24525 , \23202 , \21417 );
nor \U$24182 ( \24526 , \24524 , \24525 );
xnor \U$24183 ( \24527 , \24526 , \21426 );
and \U$24184 ( \24528 , \24522 , \24527 );
and \U$24185 ( \24529 , \24518 , \24527 );
or \U$24186 ( \24530 , \24523 , \24528 , \24529 );
and \U$24187 ( \24531 , \24513 , \24530 );
and \U$24188 ( \24532 , \24496 , \24530 );
or \U$24189 ( \24533 , \24514 , \24531 , \24532 );
and \U$24190 ( \24534 , \24480 , \24533 );
and \U$24191 ( \24535 , \24506 , \21464 );
xor \U$24192 ( \24536 , \24312 , \24316 );
xor \U$24193 ( \24537 , \24536 , \24321 );
and \U$24194 ( \24538 , \24535 , \24537 );
xor \U$24195 ( \24539 , \24345 , \24349 );
xor \U$24196 ( \24540 , \24539 , \24354 );
and \U$24197 ( \24541 , \24537 , \24540 );
and \U$24198 ( \24542 , \24535 , \24540 );
or \U$24199 ( \24543 , \24538 , \24541 , \24542 );
and \U$24200 ( \24544 , \24533 , \24543 );
and \U$24201 ( \24545 , \24480 , \24543 );
or \U$24202 ( \24546 , \24534 , \24544 , \24545 );
xor \U$24203 ( \24547 , \24258 , \24262 );
xor \U$24204 ( \24548 , \24547 , \24267 );
xor \U$24205 ( \24549 , \24328 , \24332 );
xor \U$24206 ( \24550 , \24549 , \24337 );
and \U$24207 ( \24551 , \24548 , \24550 );
xor \U$24208 ( \24552 , \24293 , \24297 );
xor \U$24209 ( \24553 , \24552 , \24302 );
and \U$24210 ( \24554 , \24550 , \24553 );
and \U$24211 ( \24555 , \24548 , \24553 );
or \U$24212 ( \24556 , \24551 , \24554 , \24555 );
xor \U$24213 ( \24557 , \24152 , \24156 );
xor \U$24214 ( \24558 , \24557 , \24161 );
and \U$24215 ( \24559 , \24556 , \24558 );
xor \U$24216 ( \24560 , \24371 , \24373 );
xor \U$24217 ( \24561 , \24560 , \24376 );
and \U$24218 ( \24562 , \24558 , \24561 );
and \U$24219 ( \24563 , \24556 , \24561 );
or \U$24220 ( \24564 , \24559 , \24562 , \24563 );
and \U$24221 ( \24565 , \24546 , \24564 );
xor \U$24222 ( \24566 , \24270 , \24288 );
xor \U$24223 ( \24567 , \24566 , \24305 );
xor \U$24224 ( \24568 , \24324 , \24340 );
xor \U$24225 ( \24569 , \24568 , \24357 );
and \U$24226 ( \24570 , \24567 , \24569 );
xnor \U$24227 ( \24571 , \24363 , \24365 );
and \U$24228 ( \24572 , \24569 , \24571 );
and \U$24229 ( \24573 , \24567 , \24571 );
or \U$24230 ( \24574 , \24570 , \24572 , \24573 );
and \U$24231 ( \24575 , \24564 , \24574 );
and \U$24232 ( \24576 , \24546 , \24574 );
or \U$24233 ( \24577 , \24565 , \24575 , \24576 );
xor \U$24234 ( \24578 , \24308 , \24360 );
xor \U$24235 ( \24579 , \24578 , \24366 );
xor \U$24236 ( \24580 , \24379 , \24381 );
xor \U$24237 ( \24581 , \24580 , \24384 );
and \U$24238 ( \24582 , \24579 , \24581 );
xor \U$24239 ( \24583 , \24390 , \24392 );
and \U$24240 ( \24584 , \24581 , \24583 );
and \U$24241 ( \24585 , \24579 , \24583 );
or \U$24242 ( \24586 , \24582 , \24584 , \24585 );
and \U$24243 ( \24587 , \24577 , \24586 );
xor \U$24244 ( \24588 , \24398 , \24400 );
xor \U$24245 ( \24589 , \24588 , \24402 );
and \U$24246 ( \24590 , \24586 , \24589 );
and \U$24247 ( \24591 , \24577 , \24589 );
or \U$24248 ( \24592 , \24587 , \24590 , \24591 );
xor \U$24249 ( \24593 , \24198 , \24216 );
xor \U$24250 ( \24594 , \24593 , \24222 );
and \U$24251 ( \24595 , \24592 , \24594 );
xor \U$24252 ( \24596 , \24396 , \24405 );
xor \U$24253 ( \24597 , \24596 , \24408 );
and \U$24254 ( \24598 , \24594 , \24597 );
and \U$24255 ( \24599 , \24592 , \24597 );
or \U$24256 ( \24600 , \24595 , \24598 , \24599 );
xor \U$24257 ( \24601 , \24411 , \24413 );
xor \U$24258 ( \24602 , \24601 , \24416 );
and \U$24259 ( \24603 , \24600 , \24602 );
and \U$24260 ( \24604 , \24425 , \24603 );
xor \U$24261 ( \24605 , \24425 , \24603 );
xor \U$24262 ( \24606 , \24600 , \24602 );
buf \U$24263 ( \24607 , RIbb2e4b8_38);
buf \U$24264 ( \24608 , RIbb2e440_39);
and \U$24265 ( \24609 , \24607 , \24608 );
not \U$24266 ( \24610 , \24609 );
and \U$24267 ( \24611 , \24272 , \24610 );
not \U$24268 ( \24612 , \24611 );
and \U$24269 ( \24613 , \21379 , \24462 );
and \U$24270 ( \24614 , \21387 , \24460 );
nor \U$24271 ( \24615 , \24613 , \24614 );
xnor \U$24272 ( \24616 , \24615 , \24275 );
and \U$24273 ( \24617 , \24612 , \24616 );
and \U$24274 ( \24618 , \21395 , \24149 );
and \U$24275 ( \24619 , \21403 , \24147 );
nor \U$24276 ( \24620 , \24618 , \24619 );
xnor \U$24277 ( \24621 , \24620 , \23944 );
and \U$24278 ( \24622 , \24616 , \24621 );
and \U$24279 ( \24623 , \24612 , \24621 );
or \U$24280 ( \24624 , \24617 , \24622 , \24623 );
and \U$24281 ( \24625 , \21413 , \23743 );
and \U$24282 ( \24626 , \21421 , \23741 );
nor \U$24283 ( \24627 , \24625 , \24626 );
xnor \U$24284 ( \24628 , \24627 , \23594 );
and \U$24285 ( \24629 , \21428 , \23421 );
and \U$24286 ( \24630 , \21436 , \23419 );
nor \U$24287 ( \24631 , \24629 , \24630 );
xnor \U$24288 ( \24632 , \24631 , \23279 );
and \U$24289 ( \24633 , \24628 , \24632 );
and \U$24290 ( \24634 , \21444 , \23125 );
and \U$24291 ( \24635 , \21452 , \23123 );
nor \U$24292 ( \24636 , \24634 , \24635 );
xnor \U$24293 ( \24637 , \24636 , \22988 );
and \U$24294 ( \24638 , \24632 , \24637 );
and \U$24295 ( \24639 , \24628 , \24637 );
or \U$24296 ( \24640 , \24633 , \24638 , \24639 );
and \U$24297 ( \24641 , \24624 , \24640 );
and \U$24298 ( \24642 , \21463 , \22919 );
and \U$24299 ( \24643 , \21471 , \22917 );
nor \U$24300 ( \24644 , \24642 , \24643 );
xnor \U$24301 ( \24645 , \24644 , \22767 );
and \U$24302 ( \24646 , \21689 , \22651 );
and \U$24303 ( \24647 , \21478 , \22649 );
nor \U$24304 ( \24648 , \24646 , \24647 );
xnor \U$24305 ( \24649 , \24648 , \22495 );
and \U$24306 ( \24650 , \24645 , \24649 );
and \U$24307 ( \24651 , \21813 , \22379 );
and \U$24308 ( \24652 , \21750 , \22377 );
nor \U$24309 ( \24653 , \24651 , \24652 );
xnor \U$24310 ( \24654 , \24653 , \22266 );
and \U$24311 ( \24655 , \24649 , \24654 );
and \U$24312 ( \24656 , \24645 , \24654 );
or \U$24313 ( \24657 , \24650 , \24655 , \24656 );
and \U$24314 ( \24658 , \24640 , \24657 );
and \U$24315 ( \24659 , \24624 , \24657 );
or \U$24316 ( \24660 , \24641 , \24658 , \24659 );
and \U$24317 ( \24661 , \22624 , \21652 );
and \U$24318 ( \24662 , \22616 , \21650 );
nor \U$24319 ( \24663 , \24661 , \24662 );
xnor \U$24320 ( \24664 , \24663 , \21377 );
and \U$24321 ( \24665 , \22872 , \21385 );
and \U$24322 ( \24666 , \22867 , \21383 );
nor \U$24323 ( \24667 , \24665 , \24666 );
xnor \U$24324 ( \24668 , \24667 , \21392 );
and \U$24325 ( \24669 , \24664 , \24668 );
and \U$24326 ( \24670 , \23202 , \21401 );
and \U$24327 ( \24671 , \23058 , \21399 );
nor \U$24328 ( \24672 , \24670 , \24671 );
xnor \U$24329 ( \24673 , \24672 , \21408 );
and \U$24330 ( \24674 , \24668 , \24673 );
and \U$24331 ( \24675 , \24664 , \24673 );
or \U$24332 ( \24676 , \24669 , \24674 , \24675 );
and \U$24333 ( \24677 , \22099 , \22185 );
and \U$24334 ( \24678 , \22011 , \22183 );
nor \U$24335 ( \24679 , \24677 , \24678 );
xnor \U$24336 ( \24680 , \24679 , \22049 );
and \U$24337 ( \24681 , \22209 , \21985 );
and \U$24338 ( \24682 , \22204 , \21983 );
nor \U$24339 ( \24683 , \24681 , \24682 );
xnor \U$24340 ( \24684 , \24683 , \21907 );
and \U$24341 ( \24685 , \24680 , \24684 );
and \U$24342 ( \24686 , \22440 , \21821 );
and \U$24343 ( \24687 , \22325 , \21819 );
nor \U$24344 ( \24688 , \24686 , \24687 );
xnor \U$24345 ( \24689 , \24688 , \21727 );
and \U$24346 ( \24690 , \24684 , \24689 );
and \U$24347 ( \24691 , \24680 , \24689 );
or \U$24348 ( \24692 , \24685 , \24690 , \24691 );
and \U$24349 ( \24693 , \24676 , \24692 );
and \U$24350 ( \24694 , \23491 , \21419 );
and \U$24351 ( \24695 , \23466 , \21417 );
nor \U$24352 ( \24696 , \24694 , \24695 );
xnor \U$24353 ( \24697 , \24696 , \21426 );
and \U$24354 ( \24698 , \23832 , \21434 );
and \U$24355 ( \24699 , \23665 , \21432 );
nor \U$24356 ( \24700 , \24698 , \24699 );
xnor \U$24357 ( \24701 , \24700 , \21441 );
and \U$24358 ( \24702 , \24697 , \24701 );
and \U$24359 ( \24703 , \24089 , \21450 );
and \U$24360 ( \24704 , \23970 , \21448 );
nor \U$24361 ( \24705 , \24703 , \24704 );
xnor \U$24362 ( \24706 , \24705 , \21457 );
and \U$24363 ( \24707 , \24701 , \24706 );
and \U$24364 ( \24708 , \24697 , \24706 );
or \U$24365 ( \24709 , \24702 , \24707 , \24708 );
and \U$24366 ( \24710 , \24692 , \24709 );
and \U$24367 ( \24711 , \24676 , \24709 );
or \U$24368 ( \24712 , \24693 , \24710 , \24711 );
and \U$24369 ( \24713 , \24660 , \24712 );
buf \U$24370 ( \24714 , RIbb32658_164);
and \U$24371 ( \24715 , \24714 , \21464 );
xor \U$24372 ( \24716 , \24500 , \24504 );
xor \U$24373 ( \24717 , \24716 , \24510 );
or \U$24374 ( \24718 , \24715 , \24717 );
and \U$24375 ( \24719 , \24712 , \24718 );
and \U$24376 ( \24720 , \24660 , \24718 );
or \U$24377 ( \24721 , \24713 , \24719 , \24720 );
xor \U$24378 ( \24722 , \24429 , \24433 );
xor \U$24379 ( \24723 , \24722 , \24438 );
xor \U$24380 ( \24724 , \24484 , \24488 );
xor \U$24381 ( \24725 , \24724 , \24493 );
and \U$24382 ( \24726 , \24723 , \24725 );
xor \U$24383 ( \24727 , \24518 , \24522 );
xor \U$24384 ( \24728 , \24727 , \24527 );
and \U$24385 ( \24729 , \24725 , \24728 );
and \U$24386 ( \24730 , \24723 , \24728 );
or \U$24387 ( \24731 , \24726 , \24729 , \24730 );
xor \U$24388 ( \24732 , \24276 , \24280 );
xor \U$24389 ( \24733 , \24732 , \24285 );
and \U$24390 ( \24734 , \24731 , \24733 );
xor \U$24391 ( \24735 , \24548 , \24550 );
xor \U$24392 ( \24736 , \24735 , \24553 );
and \U$24393 ( \24737 , \24733 , \24736 );
and \U$24394 ( \24738 , \24731 , \24736 );
or \U$24395 ( \24739 , \24734 , \24737 , \24738 );
and \U$24396 ( \24740 , \24721 , \24739 );
xor \U$24397 ( \24741 , \24441 , \24457 );
xor \U$24398 ( \24742 , \24741 , \24477 );
xor \U$24399 ( \24743 , \24496 , \24513 );
xor \U$24400 ( \24744 , \24743 , \24530 );
and \U$24401 ( \24745 , \24742 , \24744 );
xor \U$24402 ( \24746 , \24535 , \24537 );
xor \U$24403 ( \24747 , \24746 , \24540 );
and \U$24404 ( \24748 , \24744 , \24747 );
and \U$24405 ( \24749 , \24742 , \24747 );
or \U$24406 ( \24750 , \24745 , \24748 , \24749 );
and \U$24407 ( \24751 , \24739 , \24750 );
and \U$24408 ( \24752 , \24721 , \24750 );
or \U$24409 ( \24753 , \24740 , \24751 , \24752 );
xor \U$24410 ( \24754 , \24480 , \24533 );
xor \U$24411 ( \24755 , \24754 , \24543 );
xor \U$24412 ( \24756 , \24556 , \24558 );
xor \U$24413 ( \24757 , \24756 , \24561 );
and \U$24414 ( \24758 , \24755 , \24757 );
xor \U$24415 ( \24759 , \24567 , \24569 );
xor \U$24416 ( \24760 , \24759 , \24571 );
and \U$24417 ( \24761 , \24757 , \24760 );
and \U$24418 ( \24762 , \24755 , \24760 );
or \U$24419 ( \24763 , \24758 , \24761 , \24762 );
and \U$24420 ( \24764 , \24753 , \24763 );
xor \U$24421 ( \24765 , \24579 , \24581 );
xor \U$24422 ( \24766 , \24765 , \24583 );
and \U$24423 ( \24767 , \24763 , \24766 );
and \U$24424 ( \24768 , \24753 , \24766 );
or \U$24425 ( \24769 , \24764 , \24767 , \24768 );
xor \U$24426 ( \24770 , \24369 , \24387 );
xor \U$24427 ( \24771 , \24770 , \24393 );
and \U$24428 ( \24772 , \24769 , \24771 );
xor \U$24429 ( \24773 , \24577 , \24586 );
xor \U$24430 ( \24774 , \24773 , \24589 );
and \U$24431 ( \24775 , \24771 , \24774 );
and \U$24432 ( \24776 , \24769 , \24774 );
or \U$24433 ( \24777 , \24772 , \24775 , \24776 );
xor \U$24434 ( \24778 , \24592 , \24594 );
xor \U$24435 ( \24779 , \24778 , \24597 );
and \U$24436 ( \24780 , \24777 , \24779 );
and \U$24437 ( \24781 , \24606 , \24780 );
xor \U$24438 ( \24782 , \24606 , \24780 );
xor \U$24439 ( \24783 , \24777 , \24779 );
and \U$24440 ( \24784 , \22204 , \22185 );
and \U$24441 ( \24785 , \22099 , \22183 );
nor \U$24442 ( \24786 , \24784 , \24785 );
xnor \U$24443 ( \24787 , \24786 , \22049 );
and \U$24444 ( \24788 , \22325 , \21985 );
and \U$24445 ( \24789 , \22209 , \21983 );
nor \U$24446 ( \24790 , \24788 , \24789 );
xnor \U$24447 ( \24791 , \24790 , \21907 );
and \U$24448 ( \24792 , \24787 , \24791 );
and \U$24449 ( \24793 , \22616 , \21821 );
and \U$24450 ( \24794 , \22440 , \21819 );
nor \U$24451 ( \24795 , \24793 , \24794 );
xnor \U$24452 ( \24796 , \24795 , \21727 );
and \U$24453 ( \24797 , \24791 , \24796 );
and \U$24454 ( \24798 , \24787 , \24796 );
or \U$24455 ( \24799 , \24792 , \24797 , \24798 );
and \U$24456 ( \24800 , \22867 , \21652 );
and \U$24457 ( \24801 , \22624 , \21650 );
nor \U$24458 ( \24802 , \24800 , \24801 );
xnor \U$24459 ( \24803 , \24802 , \21377 );
and \U$24460 ( \24804 , \23058 , \21385 );
and \U$24461 ( \24805 , \22872 , \21383 );
nor \U$24462 ( \24806 , \24804 , \24805 );
xnor \U$24463 ( \24807 , \24806 , \21392 );
and \U$24464 ( \24808 , \24803 , \24807 );
and \U$24465 ( \24809 , \23466 , \21401 );
and \U$24466 ( \24810 , \23202 , \21399 );
nor \U$24467 ( \24811 , \24809 , \24810 );
xnor \U$24468 ( \24812 , \24811 , \21408 );
and \U$24469 ( \24813 , \24807 , \24812 );
and \U$24470 ( \24814 , \24803 , \24812 );
or \U$24471 ( \24815 , \24808 , \24813 , \24814 );
and \U$24472 ( \24816 , \24799 , \24815 );
and \U$24473 ( \24817 , \23665 , \21419 );
and \U$24474 ( \24818 , \23491 , \21417 );
nor \U$24475 ( \24819 , \24817 , \24818 );
xnor \U$24476 ( \24820 , \24819 , \21426 );
and \U$24477 ( \24821 , \23970 , \21434 );
and \U$24478 ( \24822 , \23832 , \21432 );
nor \U$24479 ( \24823 , \24821 , \24822 );
xnor \U$24480 ( \24824 , \24823 , \21441 );
and \U$24481 ( \24825 , \24820 , \24824 );
and \U$24482 ( \24826 , \24506 , \21450 );
and \U$24483 ( \24827 , \24089 , \21448 );
nor \U$24484 ( \24828 , \24826 , \24827 );
xnor \U$24485 ( \24829 , \24828 , \21457 );
and \U$24486 ( \24830 , \24824 , \24829 );
and \U$24487 ( \24831 , \24820 , \24829 );
or \U$24488 ( \24832 , \24825 , \24830 , \24831 );
and \U$24489 ( \24833 , \24815 , \24832 );
and \U$24490 ( \24834 , \24799 , \24832 );
or \U$24491 ( \24835 , \24816 , \24833 , \24834 );
buf \U$24492 ( \24836 , RIbb326d0_165);
and \U$24493 ( \24837 , \24836 , \21469 );
and \U$24494 ( \24838 , \24714 , \21467 );
nor \U$24495 ( \24839 , \24837 , \24838 );
xnor \U$24496 ( \24840 , \24839 , \21476 );
buf \U$24497 ( \24841 , RIbb32748_166);
and \U$24498 ( \24842 , \24841 , \21464 );
or \U$24499 ( \24843 , \24840 , \24842 );
and \U$24500 ( \24844 , \24714 , \21469 );
and \U$24501 ( \24845 , \24506 , \21467 );
nor \U$24502 ( \24846 , \24844 , \24845 );
xnor \U$24503 ( \24847 , \24846 , \21476 );
and \U$24504 ( \24848 , \24843 , \24847 );
and \U$24505 ( \24849 , \24836 , \21464 );
and \U$24506 ( \24850 , \24847 , \24849 );
and \U$24507 ( \24851 , \24843 , \24849 );
or \U$24508 ( \24852 , \24848 , \24850 , \24851 );
and \U$24509 ( \24853 , \24835 , \24852 );
xor \U$24510 ( \24854 , \24272 , \24607 );
xor \U$24511 ( \24855 , \24607 , \24608 );
not \U$24512 ( \24856 , \24855 );
and \U$24513 ( \24857 , \24854 , \24856 );
and \U$24514 ( \24858 , \21387 , \24857 );
not \U$24515 ( \24859 , \24858 );
xnor \U$24516 ( \24860 , \24859 , \24611 );
and \U$24517 ( \24861 , \21403 , \24462 );
and \U$24518 ( \24862 , \21379 , \24460 );
nor \U$24519 ( \24863 , \24861 , \24862 );
xnor \U$24520 ( \24864 , \24863 , \24275 );
and \U$24521 ( \24865 , \24860 , \24864 );
and \U$24522 ( \24866 , \21421 , \24149 );
and \U$24523 ( \24867 , \21395 , \24147 );
nor \U$24524 ( \24868 , \24866 , \24867 );
xnor \U$24525 ( \24869 , \24868 , \23944 );
and \U$24526 ( \24870 , \24864 , \24869 );
and \U$24527 ( \24871 , \24860 , \24869 );
or \U$24528 ( \24872 , \24865 , \24870 , \24871 );
and \U$24529 ( \24873 , \21436 , \23743 );
and \U$24530 ( \24874 , \21413 , \23741 );
nor \U$24531 ( \24875 , \24873 , \24874 );
xnor \U$24532 ( \24876 , \24875 , \23594 );
and \U$24533 ( \24877 , \21452 , \23421 );
and \U$24534 ( \24878 , \21428 , \23419 );
nor \U$24535 ( \24879 , \24877 , \24878 );
xnor \U$24536 ( \24880 , \24879 , \23279 );
and \U$24537 ( \24881 , \24876 , \24880 );
and \U$24538 ( \24882 , \21471 , \23125 );
and \U$24539 ( \24883 , \21444 , \23123 );
nor \U$24540 ( \24884 , \24882 , \24883 );
xnor \U$24541 ( \24885 , \24884 , \22988 );
and \U$24542 ( \24886 , \24880 , \24885 );
and \U$24543 ( \24887 , \24876 , \24885 );
or \U$24544 ( \24888 , \24881 , \24886 , \24887 );
and \U$24545 ( \24889 , \24872 , \24888 );
and \U$24546 ( \24890 , \21478 , \22919 );
and \U$24547 ( \24891 , \21463 , \22917 );
nor \U$24548 ( \24892 , \24890 , \24891 );
xnor \U$24549 ( \24893 , \24892 , \22767 );
and \U$24550 ( \24894 , \21750 , \22651 );
and \U$24551 ( \24895 , \21689 , \22649 );
nor \U$24552 ( \24896 , \24894 , \24895 );
xnor \U$24553 ( \24897 , \24896 , \22495 );
and \U$24554 ( \24898 , \24893 , \24897 );
and \U$24555 ( \24899 , \22011 , \22379 );
and \U$24556 ( \24900 , \21813 , \22377 );
nor \U$24557 ( \24901 , \24899 , \24900 );
xnor \U$24558 ( \24902 , \24901 , \22266 );
and \U$24559 ( \24903 , \24897 , \24902 );
and \U$24560 ( \24904 , \24893 , \24902 );
or \U$24561 ( \24905 , \24898 , \24903 , \24904 );
and \U$24562 ( \24906 , \24888 , \24905 );
and \U$24563 ( \24907 , \24872 , \24905 );
or \U$24564 ( \24908 , \24889 , \24906 , \24907 );
and \U$24565 ( \24909 , \24852 , \24908 );
and \U$24566 ( \24910 , \24835 , \24908 );
or \U$24567 ( \24911 , \24853 , \24909 , \24910 );
xor \U$24568 ( \24912 , \24664 , \24668 );
xor \U$24569 ( \24913 , \24912 , \24673 );
xor \U$24570 ( \24914 , \24680 , \24684 );
xor \U$24571 ( \24915 , \24914 , \24689 );
and \U$24572 ( \24916 , \24913 , \24915 );
xor \U$24573 ( \24917 , \24697 , \24701 );
xor \U$24574 ( \24918 , \24917 , \24706 );
and \U$24575 ( \24919 , \24915 , \24918 );
and \U$24576 ( \24920 , \24913 , \24918 );
or \U$24577 ( \24921 , \24916 , \24919 , \24920 );
xor \U$24578 ( \24922 , \24612 , \24616 );
xor \U$24579 ( \24923 , \24922 , \24621 );
xor \U$24580 ( \24924 , \24628 , \24632 );
xor \U$24581 ( \24925 , \24924 , \24637 );
and \U$24582 ( \24926 , \24923 , \24925 );
xor \U$24583 ( \24927 , \24645 , \24649 );
xor \U$24584 ( \24928 , \24927 , \24654 );
and \U$24585 ( \24929 , \24925 , \24928 );
and \U$24586 ( \24930 , \24923 , \24928 );
or \U$24587 ( \24931 , \24926 , \24929 , \24930 );
and \U$24588 ( \24932 , \24921 , \24931 );
xor \U$24589 ( \24933 , \24445 , \24449 );
xor \U$24590 ( \24934 , \24933 , \24454 );
and \U$24591 ( \24935 , \24931 , \24934 );
and \U$24592 ( \24936 , \24921 , \24934 );
or \U$24593 ( \24937 , \24932 , \24935 , \24936 );
and \U$24594 ( \24938 , \24911 , \24937 );
xor \U$24595 ( \24939 , \24465 , \24469 );
xor \U$24596 ( \24940 , \24939 , \24474 );
xor \U$24597 ( \24941 , \24723 , \24725 );
xor \U$24598 ( \24942 , \24941 , \24728 );
and \U$24599 ( \24943 , \24940 , \24942 );
xnor \U$24600 ( \24944 , \24715 , \24717 );
and \U$24601 ( \24945 , \24942 , \24944 );
and \U$24602 ( \24946 , \24940 , \24944 );
or \U$24603 ( \24947 , \24943 , \24945 , \24946 );
and \U$24604 ( \24948 , \24937 , \24947 );
and \U$24605 ( \24949 , \24911 , \24947 );
or \U$24606 ( \24950 , \24938 , \24948 , \24949 );
xor \U$24607 ( \24951 , \24660 , \24712 );
xor \U$24608 ( \24952 , \24951 , \24718 );
xor \U$24609 ( \24953 , \24731 , \24733 );
xor \U$24610 ( \24954 , \24953 , \24736 );
and \U$24611 ( \24955 , \24952 , \24954 );
xor \U$24612 ( \24956 , \24742 , \24744 );
xor \U$24613 ( \24957 , \24956 , \24747 );
and \U$24614 ( \24958 , \24954 , \24957 );
and \U$24615 ( \24959 , \24952 , \24957 );
or \U$24616 ( \24960 , \24955 , \24958 , \24959 );
and \U$24617 ( \24961 , \24950 , \24960 );
xor \U$24618 ( \24962 , \24755 , \24757 );
xor \U$24619 ( \24963 , \24962 , \24760 );
and \U$24620 ( \24964 , \24960 , \24963 );
and \U$24621 ( \24965 , \24950 , \24963 );
or \U$24622 ( \24966 , \24961 , \24964 , \24965 );
xor \U$24623 ( \24967 , \24546 , \24564 );
xor \U$24624 ( \24968 , \24967 , \24574 );
and \U$24625 ( \24969 , \24966 , \24968 );
xor \U$24626 ( \24970 , \24753 , \24763 );
xor \U$24627 ( \24971 , \24970 , \24766 );
and \U$24628 ( \24972 , \24968 , \24971 );
and \U$24629 ( \24973 , \24966 , \24971 );
or \U$24630 ( \24974 , \24969 , \24972 , \24973 );
xor \U$24631 ( \24975 , \24769 , \24771 );
xor \U$24632 ( \24976 , \24975 , \24774 );
and \U$24633 ( \24977 , \24974 , \24976 );
and \U$24634 ( \24978 , \24783 , \24977 );
xor \U$24635 ( \24979 , \24783 , \24977 );
xor \U$24636 ( \24980 , \24974 , \24976 );
and \U$24637 ( \24981 , \22624 , \21821 );
and \U$24638 ( \24982 , \22616 , \21819 );
nor \U$24639 ( \24983 , \24981 , \24982 );
xnor \U$24640 ( \24984 , \24983 , \21727 );
and \U$24641 ( \24985 , \22872 , \21652 );
and \U$24642 ( \24986 , \22867 , \21650 );
nor \U$24643 ( \24987 , \24985 , \24986 );
xnor \U$24644 ( \24988 , \24987 , \21377 );
and \U$24645 ( \24989 , \24984 , \24988 );
and \U$24646 ( \24990 , \23202 , \21385 );
and \U$24647 ( \24991 , \23058 , \21383 );
nor \U$24648 ( \24992 , \24990 , \24991 );
xnor \U$24649 ( \24993 , \24992 , \21392 );
and \U$24650 ( \24994 , \24988 , \24993 );
and \U$24651 ( \24995 , \24984 , \24993 );
or \U$24652 ( \24996 , \24989 , \24994 , \24995 );
and \U$24653 ( \24997 , \22099 , \22379 );
and \U$24654 ( \24998 , \22011 , \22377 );
nor \U$24655 ( \24999 , \24997 , \24998 );
xnor \U$24656 ( \25000 , \24999 , \22266 );
and \U$24657 ( \25001 , \22209 , \22185 );
and \U$24658 ( \25002 , \22204 , \22183 );
nor \U$24659 ( \25003 , \25001 , \25002 );
xnor \U$24660 ( \25004 , \25003 , \22049 );
and \U$24661 ( \25005 , \25000 , \25004 );
and \U$24662 ( \25006 , \22440 , \21985 );
and \U$24663 ( \25007 , \22325 , \21983 );
nor \U$24664 ( \25008 , \25006 , \25007 );
xnor \U$24665 ( \25009 , \25008 , \21907 );
and \U$24666 ( \25010 , \25004 , \25009 );
and \U$24667 ( \25011 , \25000 , \25009 );
or \U$24668 ( \25012 , \25005 , \25010 , \25011 );
and \U$24669 ( \25013 , \24996 , \25012 );
and \U$24670 ( \25014 , \23491 , \21401 );
and \U$24671 ( \25015 , \23466 , \21399 );
nor \U$24672 ( \25016 , \25014 , \25015 );
xnor \U$24673 ( \25017 , \25016 , \21408 );
and \U$24674 ( \25018 , \23832 , \21419 );
and \U$24675 ( \25019 , \23665 , \21417 );
nor \U$24676 ( \25020 , \25018 , \25019 );
xnor \U$24677 ( \25021 , \25020 , \21426 );
and \U$24678 ( \25022 , \25017 , \25021 );
and \U$24679 ( \25023 , \24089 , \21434 );
and \U$24680 ( \25024 , \23970 , \21432 );
nor \U$24681 ( \25025 , \25023 , \25024 );
xnor \U$24682 ( \25026 , \25025 , \21441 );
and \U$24683 ( \25027 , \25021 , \25026 );
and \U$24684 ( \25028 , \25017 , \25026 );
or \U$24685 ( \25029 , \25022 , \25027 , \25028 );
and \U$24686 ( \25030 , \25012 , \25029 );
and \U$24687 ( \25031 , \24996 , \25029 );
or \U$24688 ( \25032 , \25013 , \25030 , \25031 );
buf \U$24689 ( \25033 , RIbb2e3c8_40);
buf \U$24690 ( \25034 , RIbb2e350_41);
and \U$24691 ( \25035 , \25033 , \25034 );
not \U$24692 ( \25036 , \25035 );
and \U$24693 ( \25037 , \24608 , \25036 );
not \U$24694 ( \25038 , \25037 );
and \U$24695 ( \25039 , \21379 , \24857 );
and \U$24696 ( \25040 , \21387 , \24855 );
nor \U$24697 ( \25041 , \25039 , \25040 );
xnor \U$24698 ( \25042 , \25041 , \24611 );
and \U$24699 ( \25043 , \25038 , \25042 );
and \U$24700 ( \25044 , \21395 , \24462 );
and \U$24701 ( \25045 , \21403 , \24460 );
nor \U$24702 ( \25046 , \25044 , \25045 );
xnor \U$24703 ( \25047 , \25046 , \24275 );
and \U$24704 ( \25048 , \25042 , \25047 );
and \U$24705 ( \25049 , \25038 , \25047 );
or \U$24706 ( \25050 , \25043 , \25048 , \25049 );
and \U$24707 ( \25051 , \21413 , \24149 );
and \U$24708 ( \25052 , \21421 , \24147 );
nor \U$24709 ( \25053 , \25051 , \25052 );
xnor \U$24710 ( \25054 , \25053 , \23944 );
and \U$24711 ( \25055 , \21428 , \23743 );
and \U$24712 ( \25056 , \21436 , \23741 );
nor \U$24713 ( \25057 , \25055 , \25056 );
xnor \U$24714 ( \25058 , \25057 , \23594 );
and \U$24715 ( \25059 , \25054 , \25058 );
and \U$24716 ( \25060 , \21444 , \23421 );
and \U$24717 ( \25061 , \21452 , \23419 );
nor \U$24718 ( \25062 , \25060 , \25061 );
xnor \U$24719 ( \25063 , \25062 , \23279 );
and \U$24720 ( \25064 , \25058 , \25063 );
and \U$24721 ( \25065 , \25054 , \25063 );
or \U$24722 ( \25066 , \25059 , \25064 , \25065 );
and \U$24723 ( \25067 , \25050 , \25066 );
and \U$24724 ( \25068 , \21463 , \23125 );
and \U$24725 ( \25069 , \21471 , \23123 );
nor \U$24726 ( \25070 , \25068 , \25069 );
xnor \U$24727 ( \25071 , \25070 , \22988 );
and \U$24728 ( \25072 , \21689 , \22919 );
and \U$24729 ( \25073 , \21478 , \22917 );
nor \U$24730 ( \25074 , \25072 , \25073 );
xnor \U$24731 ( \25075 , \25074 , \22767 );
and \U$24732 ( \25076 , \25071 , \25075 );
and \U$24733 ( \25077 , \21813 , \22651 );
and \U$24734 ( \25078 , \21750 , \22649 );
nor \U$24735 ( \25079 , \25077 , \25078 );
xnor \U$24736 ( \25080 , \25079 , \22495 );
and \U$24737 ( \25081 , \25075 , \25080 );
and \U$24738 ( \25082 , \25071 , \25080 );
or \U$24739 ( \25083 , \25076 , \25081 , \25082 );
and \U$24740 ( \25084 , \25066 , \25083 );
and \U$24741 ( \25085 , \25050 , \25083 );
or \U$24742 ( \25086 , \25067 , \25084 , \25085 );
and \U$24743 ( \25087 , \25032 , \25086 );
and \U$24744 ( \25088 , \24714 , \21450 );
and \U$24745 ( \25089 , \24506 , \21448 );
nor \U$24746 ( \25090 , \25088 , \25089 );
xnor \U$24747 ( \25091 , \25090 , \21457 );
and \U$24748 ( \25092 , \24841 , \21469 );
and \U$24749 ( \25093 , \24836 , \21467 );
nor \U$24750 ( \25094 , \25092 , \25093 );
xnor \U$24751 ( \25095 , \25094 , \21476 );
and \U$24752 ( \25096 , \25091 , \25095 );
buf \U$24753 ( \25097 , RIbb327c0_167);
and \U$24754 ( \25098 , \25097 , \21464 );
and \U$24755 ( \25099 , \25095 , \25098 );
and \U$24756 ( \25100 , \25091 , \25098 );
or \U$24757 ( \25101 , \25096 , \25099 , \25100 );
xor \U$24758 ( \25102 , \24820 , \24824 );
xor \U$24759 ( \25103 , \25102 , \24829 );
and \U$24760 ( \25104 , \25101 , \25103 );
xnor \U$24761 ( \25105 , \24840 , \24842 );
and \U$24762 ( \25106 , \25103 , \25105 );
and \U$24763 ( \25107 , \25101 , \25105 );
or \U$24764 ( \25108 , \25104 , \25106 , \25107 );
and \U$24765 ( \25109 , \25086 , \25108 );
and \U$24766 ( \25110 , \25032 , \25108 );
or \U$24767 ( \25111 , \25087 , \25109 , \25110 );
xor \U$24768 ( \25112 , \24787 , \24791 );
xor \U$24769 ( \25113 , \25112 , \24796 );
xor \U$24770 ( \25114 , \24803 , \24807 );
xor \U$24771 ( \25115 , \25114 , \24812 );
and \U$24772 ( \25116 , \25113 , \25115 );
xor \U$24773 ( \25117 , \24893 , \24897 );
xor \U$24774 ( \25118 , \25117 , \24902 );
and \U$24775 ( \25119 , \25115 , \25118 );
and \U$24776 ( \25120 , \25113 , \25118 );
or \U$24777 ( \25121 , \25116 , \25119 , \25120 );
xor \U$24778 ( \25122 , \24860 , \24864 );
xor \U$24779 ( \25123 , \25122 , \24869 );
xor \U$24780 ( \25124 , \24876 , \24880 );
xor \U$24781 ( \25125 , \25124 , \24885 );
and \U$24782 ( \25126 , \25123 , \25125 );
and \U$24783 ( \25127 , \25121 , \25126 );
xor \U$24784 ( \25128 , \24923 , \24925 );
xor \U$24785 ( \25129 , \25128 , \24928 );
and \U$24786 ( \25130 , \25126 , \25129 );
and \U$24787 ( \25131 , \25121 , \25129 );
or \U$24788 ( \25132 , \25127 , \25130 , \25131 );
and \U$24789 ( \25133 , \25111 , \25132 );
xor \U$24790 ( \25134 , \24799 , \24815 );
xor \U$24791 ( \25135 , \25134 , \24832 );
xor \U$24792 ( \25136 , \24843 , \24847 );
xor \U$24793 ( \25137 , \25136 , \24849 );
and \U$24794 ( \25138 , \25135 , \25137 );
xor \U$24795 ( \25139 , \24913 , \24915 );
xor \U$24796 ( \25140 , \25139 , \24918 );
and \U$24797 ( \25141 , \25137 , \25140 );
and \U$24798 ( \25142 , \25135 , \25140 );
or \U$24799 ( \25143 , \25138 , \25141 , \25142 );
and \U$24800 ( \25144 , \25132 , \25143 );
and \U$24801 ( \25145 , \25111 , \25143 );
or \U$24802 ( \25146 , \25133 , \25144 , \25145 );
xor \U$24803 ( \25147 , \24624 , \24640 );
xor \U$24804 ( \25148 , \25147 , \24657 );
xor \U$24805 ( \25149 , \24676 , \24692 );
xor \U$24806 ( \25150 , \25149 , \24709 );
and \U$24807 ( \25151 , \25148 , \25150 );
xor \U$24808 ( \25152 , \24940 , \24942 );
xor \U$24809 ( \25153 , \25152 , \24944 );
and \U$24810 ( \25154 , \25150 , \25153 );
and \U$24811 ( \25155 , \25148 , \25153 );
or \U$24812 ( \25156 , \25151 , \25154 , \25155 );
and \U$24813 ( \25157 , \25146 , \25156 );
xor \U$24814 ( \25158 , \24952 , \24954 );
xor \U$24815 ( \25159 , \25158 , \24957 );
and \U$24816 ( \25160 , \25156 , \25159 );
and \U$24817 ( \25161 , \25146 , \25159 );
or \U$24818 ( \25162 , \25157 , \25160 , \25161 );
xor \U$24819 ( \25163 , \24721 , \24739 );
xor \U$24820 ( \25164 , \25163 , \24750 );
and \U$24821 ( \25165 , \25162 , \25164 );
xor \U$24822 ( \25166 , \24950 , \24960 );
xor \U$24823 ( \25167 , \25166 , \24963 );
and \U$24824 ( \25168 , \25164 , \25167 );
and \U$24825 ( \25169 , \25162 , \25167 );
or \U$24826 ( \25170 , \25165 , \25168 , \25169 );
xor \U$24827 ( \25171 , \24966 , \24968 );
xor \U$24828 ( \25172 , \25171 , \24971 );
and \U$24829 ( \25173 , \25170 , \25172 );
and \U$24830 ( \25174 , \24980 , \25173 );
xor \U$24831 ( \25175 , \24980 , \25173 );
xor \U$24832 ( \25176 , \25170 , \25172 );
xor \U$24833 ( \25177 , \24608 , \25033 );
xor \U$24834 ( \25178 , \25033 , \25034 );
not \U$24835 ( \25179 , \25178 );
and \U$24836 ( \25180 , \25177 , \25179 );
and \U$24837 ( \25181 , \21387 , \25180 );
not \U$24838 ( \25182 , \25181 );
xnor \U$24839 ( \25183 , \25182 , \25037 );
and \U$24840 ( \25184 , \21403 , \24857 );
and \U$24841 ( \25185 , \21379 , \24855 );
nor \U$24842 ( \25186 , \25184 , \25185 );
xnor \U$24843 ( \25187 , \25186 , \24611 );
and \U$24844 ( \25188 , \25183 , \25187 );
and \U$24845 ( \25189 , \21421 , \24462 );
and \U$24846 ( \25190 , \21395 , \24460 );
nor \U$24847 ( \25191 , \25189 , \25190 );
xnor \U$24848 ( \25192 , \25191 , \24275 );
and \U$24849 ( \25193 , \25187 , \25192 );
and \U$24850 ( \25194 , \25183 , \25192 );
or \U$24851 ( \25195 , \25188 , \25193 , \25194 );
and \U$24852 ( \25196 , \21436 , \24149 );
and \U$24853 ( \25197 , \21413 , \24147 );
nor \U$24854 ( \25198 , \25196 , \25197 );
xnor \U$24855 ( \25199 , \25198 , \23944 );
and \U$24856 ( \25200 , \21452 , \23743 );
and \U$24857 ( \25201 , \21428 , \23741 );
nor \U$24858 ( \25202 , \25200 , \25201 );
xnor \U$24859 ( \25203 , \25202 , \23594 );
and \U$24860 ( \25204 , \25199 , \25203 );
and \U$24861 ( \25205 , \21471 , \23421 );
and \U$24862 ( \25206 , \21444 , \23419 );
nor \U$24863 ( \25207 , \25205 , \25206 );
xnor \U$24864 ( \25208 , \25207 , \23279 );
and \U$24865 ( \25209 , \25203 , \25208 );
and \U$24866 ( \25210 , \25199 , \25208 );
or \U$24867 ( \25211 , \25204 , \25209 , \25210 );
and \U$24868 ( \25212 , \25195 , \25211 );
and \U$24869 ( \25213 , \21478 , \23125 );
and \U$24870 ( \25214 , \21463 , \23123 );
nor \U$24871 ( \25215 , \25213 , \25214 );
xnor \U$24872 ( \25216 , \25215 , \22988 );
and \U$24873 ( \25217 , \21750 , \22919 );
and \U$24874 ( \25218 , \21689 , \22917 );
nor \U$24875 ( \25219 , \25217 , \25218 );
xnor \U$24876 ( \25220 , \25219 , \22767 );
and \U$24877 ( \25221 , \25216 , \25220 );
and \U$24878 ( \25222 , \22011 , \22651 );
and \U$24879 ( \25223 , \21813 , \22649 );
nor \U$24880 ( \25224 , \25222 , \25223 );
xnor \U$24881 ( \25225 , \25224 , \22495 );
and \U$24882 ( \25226 , \25220 , \25225 );
and \U$24883 ( \25227 , \25216 , \25225 );
or \U$24884 ( \25228 , \25221 , \25226 , \25227 );
and \U$24885 ( \25229 , \25211 , \25228 );
and \U$24886 ( \25230 , \25195 , \25228 );
or \U$24887 ( \25231 , \25212 , \25229 , \25230 );
and \U$24888 ( \25232 , \23665 , \21401 );
and \U$24889 ( \25233 , \23491 , \21399 );
nor \U$24890 ( \25234 , \25232 , \25233 );
xnor \U$24891 ( \25235 , \25234 , \21408 );
and \U$24892 ( \25236 , \23970 , \21419 );
and \U$24893 ( \25237 , \23832 , \21417 );
nor \U$24894 ( \25238 , \25236 , \25237 );
xnor \U$24895 ( \25239 , \25238 , \21426 );
and \U$24896 ( \25240 , \25235 , \25239 );
and \U$24897 ( \25241 , \24506 , \21434 );
and \U$24898 ( \25242 , \24089 , \21432 );
nor \U$24899 ( \25243 , \25241 , \25242 );
xnor \U$24900 ( \25244 , \25243 , \21441 );
and \U$24901 ( \25245 , \25239 , \25244 );
and \U$24902 ( \25246 , \25235 , \25244 );
or \U$24903 ( \25247 , \25240 , \25245 , \25246 );
and \U$24904 ( \25248 , \22204 , \22379 );
and \U$24905 ( \25249 , \22099 , \22377 );
nor \U$24906 ( \25250 , \25248 , \25249 );
xnor \U$24907 ( \25251 , \25250 , \22266 );
and \U$24908 ( \25252 , \22325 , \22185 );
and \U$24909 ( \25253 , \22209 , \22183 );
nor \U$24910 ( \25254 , \25252 , \25253 );
xnor \U$24911 ( \25255 , \25254 , \22049 );
and \U$24912 ( \25256 , \25251 , \25255 );
and \U$24913 ( \25257 , \22616 , \21985 );
and \U$24914 ( \25258 , \22440 , \21983 );
nor \U$24915 ( \25259 , \25257 , \25258 );
xnor \U$24916 ( \25260 , \25259 , \21907 );
and \U$24917 ( \25261 , \25255 , \25260 );
and \U$24918 ( \25262 , \25251 , \25260 );
or \U$24919 ( \25263 , \25256 , \25261 , \25262 );
and \U$24920 ( \25264 , \25247 , \25263 );
and \U$24921 ( \25265 , \22867 , \21821 );
and \U$24922 ( \25266 , \22624 , \21819 );
nor \U$24923 ( \25267 , \25265 , \25266 );
xnor \U$24924 ( \25268 , \25267 , \21727 );
and \U$24925 ( \25269 , \23058 , \21652 );
and \U$24926 ( \25270 , \22872 , \21650 );
nor \U$24927 ( \25271 , \25269 , \25270 );
xnor \U$24928 ( \25272 , \25271 , \21377 );
and \U$24929 ( \25273 , \25268 , \25272 );
and \U$24930 ( \25274 , \23466 , \21385 );
and \U$24931 ( \25275 , \23202 , \21383 );
nor \U$24932 ( \25276 , \25274 , \25275 );
xnor \U$24933 ( \25277 , \25276 , \21392 );
and \U$24934 ( \25278 , \25272 , \25277 );
and \U$24935 ( \25279 , \25268 , \25277 );
or \U$24936 ( \25280 , \25273 , \25278 , \25279 );
and \U$24937 ( \25281 , \25263 , \25280 );
and \U$24938 ( \25282 , \25247 , \25280 );
or \U$24939 ( \25283 , \25264 , \25281 , \25282 );
and \U$24940 ( \25284 , \25231 , \25283 );
and \U$24941 ( \25285 , \24836 , \21450 );
and \U$24942 ( \25286 , \24714 , \21448 );
nor \U$24943 ( \25287 , \25285 , \25286 );
xnor \U$24944 ( \25288 , \25287 , \21457 );
and \U$24945 ( \25289 , \25097 , \21469 );
and \U$24946 ( \25290 , \24841 , \21467 );
nor \U$24947 ( \25291 , \25289 , \25290 );
xnor \U$24948 ( \25292 , \25291 , \21476 );
and \U$24949 ( \25293 , \25288 , \25292 );
buf \U$24950 ( \25294 , RIbb32838_168);
and \U$24951 ( \25295 , \25294 , \21464 );
and \U$24952 ( \25296 , \25292 , \25295 );
and \U$24953 ( \25297 , \25288 , \25295 );
or \U$24954 ( \25298 , \25293 , \25296 , \25297 );
xor \U$24955 ( \25299 , \25091 , \25095 );
xor \U$24956 ( \25300 , \25299 , \25098 );
and \U$24957 ( \25301 , \25298 , \25300 );
xor \U$24958 ( \25302 , \25017 , \25021 );
xor \U$24959 ( \25303 , \25302 , \25026 );
and \U$24960 ( \25304 , \25300 , \25303 );
and \U$24961 ( \25305 , \25298 , \25303 );
or \U$24962 ( \25306 , \25301 , \25304 , \25305 );
and \U$24963 ( \25307 , \25283 , \25306 );
and \U$24964 ( \25308 , \25231 , \25306 );
or \U$24965 ( \25309 , \25284 , \25307 , \25308 );
xor \U$24966 ( \25310 , \24996 , \25012 );
xor \U$24967 ( \25311 , \25310 , \25029 );
xor \U$24968 ( \25312 , \25050 , \25066 );
xor \U$24969 ( \25313 , \25312 , \25083 );
and \U$24970 ( \25314 , \25311 , \25313 );
xor \U$24971 ( \25315 , \25101 , \25103 );
xor \U$24972 ( \25316 , \25315 , \25105 );
and \U$24973 ( \25317 , \25313 , \25316 );
and \U$24974 ( \25318 , \25311 , \25316 );
or \U$24975 ( \25319 , \25314 , \25317 , \25318 );
and \U$24976 ( \25320 , \25309 , \25319 );
xor \U$24977 ( \25321 , \24984 , \24988 );
xor \U$24978 ( \25322 , \25321 , \24993 );
xor \U$24979 ( \25323 , \25000 , \25004 );
xor \U$24980 ( \25324 , \25323 , \25009 );
and \U$24981 ( \25325 , \25322 , \25324 );
xor \U$24982 ( \25326 , \25071 , \25075 );
xor \U$24983 ( \25327 , \25326 , \25080 );
and \U$24984 ( \25328 , \25324 , \25327 );
and \U$24985 ( \25329 , \25322 , \25327 );
or \U$24986 ( \25330 , \25325 , \25328 , \25329 );
xor \U$24987 ( \25331 , \25113 , \25115 );
xor \U$24988 ( \25332 , \25331 , \25118 );
and \U$24989 ( \25333 , \25330 , \25332 );
xor \U$24990 ( \25334 , \25123 , \25125 );
and \U$24991 ( \25335 , \25332 , \25334 );
and \U$24992 ( \25336 , \25330 , \25334 );
or \U$24993 ( \25337 , \25333 , \25335 , \25336 );
and \U$24994 ( \25338 , \25319 , \25337 );
and \U$24995 ( \25339 , \25309 , \25337 );
or \U$24996 ( \25340 , \25320 , \25338 , \25339 );
xor \U$24997 ( \25341 , \24872 , \24888 );
xor \U$24998 ( \25342 , \25341 , \24905 );
xor \U$24999 ( \25343 , \25121 , \25126 );
xor \U$25000 ( \25344 , \25343 , \25129 );
and \U$25001 ( \25345 , \25342 , \25344 );
xor \U$25002 ( \25346 , \25135 , \25137 );
xor \U$25003 ( \25347 , \25346 , \25140 );
and \U$25004 ( \25348 , \25344 , \25347 );
and \U$25005 ( \25349 , \25342 , \25347 );
or \U$25006 ( \25350 , \25345 , \25348 , \25349 );
and \U$25007 ( \25351 , \25340 , \25350 );
xor \U$25008 ( \25352 , \24921 , \24931 );
xor \U$25009 ( \25353 , \25352 , \24934 );
and \U$25010 ( \25354 , \25350 , \25353 );
and \U$25011 ( \25355 , \25340 , \25353 );
or \U$25012 ( \25356 , \25351 , \25354 , \25355 );
xor \U$25013 ( \25357 , \24835 , \24852 );
xor \U$25014 ( \25358 , \25357 , \24908 );
xor \U$25015 ( \25359 , \25111 , \25132 );
xor \U$25016 ( \25360 , \25359 , \25143 );
and \U$25017 ( \25361 , \25358 , \25360 );
xor \U$25018 ( \25362 , \25148 , \25150 );
xor \U$25019 ( \25363 , \25362 , \25153 );
and \U$25020 ( \25364 , \25360 , \25363 );
and \U$25021 ( \25365 , \25358 , \25363 );
or \U$25022 ( \25366 , \25361 , \25364 , \25365 );
and \U$25023 ( \25367 , \25356 , \25366 );
xor \U$25024 ( \25368 , \24911 , \24937 );
xor \U$25025 ( \25369 , \25368 , \24947 );
and \U$25026 ( \25370 , \25366 , \25369 );
and \U$25027 ( \25371 , \25356 , \25369 );
or \U$25028 ( \25372 , \25367 , \25370 , \25371 );
xor \U$25029 ( \25373 , \25162 , \25164 );
xor \U$25030 ( \25374 , \25373 , \25167 );
and \U$25031 ( \25375 , \25372 , \25374 );
and \U$25032 ( \25376 , \25176 , \25375 );
xor \U$25033 ( \25377 , \25176 , \25375 );
xor \U$25034 ( \25378 , \25372 , \25374 );
and \U$25035 ( \25379 , \21463 , \23421 );
and \U$25036 ( \25380 , \21471 , \23419 );
nor \U$25037 ( \25381 , \25379 , \25380 );
xnor \U$25038 ( \25382 , \25381 , \23279 );
and \U$25039 ( \25383 , \21689 , \23125 );
and \U$25040 ( \25384 , \21478 , \23123 );
nor \U$25041 ( \25385 , \25383 , \25384 );
xnor \U$25042 ( \25386 , \25385 , \22988 );
and \U$25043 ( \25387 , \25382 , \25386 );
and \U$25044 ( \25388 , \21813 , \22919 );
and \U$25045 ( \25389 , \21750 , \22917 );
nor \U$25046 ( \25390 , \25388 , \25389 );
xnor \U$25047 ( \25391 , \25390 , \22767 );
and \U$25048 ( \25392 , \25386 , \25391 );
and \U$25049 ( \25393 , \25382 , \25391 );
or \U$25050 ( \25394 , \25387 , \25392 , \25393 );
buf \U$25051 ( \25395 , RIbb2e2d8_42);
buf \U$25052 ( \25396 , RIbb2e260_43);
and \U$25053 ( \25397 , \25395 , \25396 );
not \U$25054 ( \25398 , \25397 );
and \U$25055 ( \25399 , \25034 , \25398 );
not \U$25056 ( \25400 , \25399 );
and \U$25057 ( \25401 , \21379 , \25180 );
and \U$25058 ( \25402 , \21387 , \25178 );
nor \U$25059 ( \25403 , \25401 , \25402 );
xnor \U$25060 ( \25404 , \25403 , \25037 );
and \U$25061 ( \25405 , \25400 , \25404 );
and \U$25062 ( \25406 , \21395 , \24857 );
and \U$25063 ( \25407 , \21403 , \24855 );
nor \U$25064 ( \25408 , \25406 , \25407 );
xnor \U$25065 ( \25409 , \25408 , \24611 );
and \U$25066 ( \25410 , \25404 , \25409 );
and \U$25067 ( \25411 , \25400 , \25409 );
or \U$25068 ( \25412 , \25405 , \25410 , \25411 );
and \U$25069 ( \25413 , \25394 , \25412 );
and \U$25070 ( \25414 , \21413 , \24462 );
and \U$25071 ( \25415 , \21421 , \24460 );
nor \U$25072 ( \25416 , \25414 , \25415 );
xnor \U$25073 ( \25417 , \25416 , \24275 );
and \U$25074 ( \25418 , \21428 , \24149 );
and \U$25075 ( \25419 , \21436 , \24147 );
nor \U$25076 ( \25420 , \25418 , \25419 );
xnor \U$25077 ( \25421 , \25420 , \23944 );
and \U$25078 ( \25422 , \25417 , \25421 );
and \U$25079 ( \25423 , \21444 , \23743 );
and \U$25080 ( \25424 , \21452 , \23741 );
nor \U$25081 ( \25425 , \25423 , \25424 );
xnor \U$25082 ( \25426 , \25425 , \23594 );
and \U$25083 ( \25427 , \25421 , \25426 );
and \U$25084 ( \25428 , \25417 , \25426 );
or \U$25085 ( \25429 , \25422 , \25427 , \25428 );
and \U$25086 ( \25430 , \25412 , \25429 );
and \U$25087 ( \25431 , \25394 , \25429 );
or \U$25088 ( \25432 , \25413 , \25430 , \25431 );
and \U$25089 ( \25433 , \23491 , \21385 );
and \U$25090 ( \25434 , \23466 , \21383 );
nor \U$25091 ( \25435 , \25433 , \25434 );
xnor \U$25092 ( \25436 , \25435 , \21392 );
and \U$25093 ( \25437 , \23832 , \21401 );
and \U$25094 ( \25438 , \23665 , \21399 );
nor \U$25095 ( \25439 , \25437 , \25438 );
xnor \U$25096 ( \25440 , \25439 , \21408 );
and \U$25097 ( \25441 , \25436 , \25440 );
and \U$25098 ( \25442 , \24089 , \21419 );
and \U$25099 ( \25443 , \23970 , \21417 );
nor \U$25100 ( \25444 , \25442 , \25443 );
xnor \U$25101 ( \25445 , \25444 , \21426 );
and \U$25102 ( \25446 , \25440 , \25445 );
and \U$25103 ( \25447 , \25436 , \25445 );
or \U$25104 ( \25448 , \25441 , \25446 , \25447 );
and \U$25105 ( \25449 , \22099 , \22651 );
and \U$25106 ( \25450 , \22011 , \22649 );
nor \U$25107 ( \25451 , \25449 , \25450 );
xnor \U$25108 ( \25452 , \25451 , \22495 );
and \U$25109 ( \25453 , \22209 , \22379 );
and \U$25110 ( \25454 , \22204 , \22377 );
nor \U$25111 ( \25455 , \25453 , \25454 );
xnor \U$25112 ( \25456 , \25455 , \22266 );
and \U$25113 ( \25457 , \25452 , \25456 );
and \U$25114 ( \25458 , \22440 , \22185 );
and \U$25115 ( \25459 , \22325 , \22183 );
nor \U$25116 ( \25460 , \25458 , \25459 );
xnor \U$25117 ( \25461 , \25460 , \22049 );
and \U$25118 ( \25462 , \25456 , \25461 );
and \U$25119 ( \25463 , \25452 , \25461 );
or \U$25120 ( \25464 , \25457 , \25462 , \25463 );
and \U$25121 ( \25465 , \25448 , \25464 );
and \U$25122 ( \25466 , \22624 , \21985 );
and \U$25123 ( \25467 , \22616 , \21983 );
nor \U$25124 ( \25468 , \25466 , \25467 );
xnor \U$25125 ( \25469 , \25468 , \21907 );
and \U$25126 ( \25470 , \22872 , \21821 );
and \U$25127 ( \25471 , \22867 , \21819 );
nor \U$25128 ( \25472 , \25470 , \25471 );
xnor \U$25129 ( \25473 , \25472 , \21727 );
and \U$25130 ( \25474 , \25469 , \25473 );
and \U$25131 ( \25475 , \23202 , \21652 );
and \U$25132 ( \25476 , \23058 , \21650 );
nor \U$25133 ( \25477 , \25475 , \25476 );
xnor \U$25134 ( \25478 , \25477 , \21377 );
and \U$25135 ( \25479 , \25473 , \25478 );
and \U$25136 ( \25480 , \25469 , \25478 );
or \U$25137 ( \25481 , \25474 , \25479 , \25480 );
and \U$25138 ( \25482 , \25464 , \25481 );
and \U$25139 ( \25483 , \25448 , \25481 );
or \U$25140 ( \25484 , \25465 , \25482 , \25483 );
and \U$25141 ( \25485 , \25432 , \25484 );
and \U$25142 ( \25486 , \24714 , \21434 );
and \U$25143 ( \25487 , \24506 , \21432 );
nor \U$25144 ( \25488 , \25486 , \25487 );
xnor \U$25145 ( \25489 , \25488 , \21441 );
and \U$25146 ( \25490 , \24841 , \21450 );
and \U$25147 ( \25491 , \24836 , \21448 );
nor \U$25148 ( \25492 , \25490 , \25491 );
xnor \U$25149 ( \25493 , \25492 , \21457 );
and \U$25150 ( \25494 , \25489 , \25493 );
and \U$25151 ( \25495 , \25294 , \21469 );
and \U$25152 ( \25496 , \25097 , \21467 );
nor \U$25153 ( \25497 , \25495 , \25496 );
xnor \U$25154 ( \25498 , \25497 , \21476 );
and \U$25155 ( \25499 , \25493 , \25498 );
and \U$25156 ( \25500 , \25489 , \25498 );
or \U$25157 ( \25501 , \25494 , \25499 , \25500 );
xor \U$25158 ( \25502 , \25288 , \25292 );
xor \U$25159 ( \25503 , \25502 , \25295 );
or \U$25160 ( \25504 , \25501 , \25503 );
and \U$25161 ( \25505 , \25484 , \25504 );
and \U$25162 ( \25506 , \25432 , \25504 );
or \U$25163 ( \25507 , \25485 , \25505 , \25506 );
xor \U$25164 ( \25508 , \25235 , \25239 );
xor \U$25165 ( \25509 , \25508 , \25244 );
xor \U$25166 ( \25510 , \25251 , \25255 );
xor \U$25167 ( \25511 , \25510 , \25260 );
and \U$25168 ( \25512 , \25509 , \25511 );
xor \U$25169 ( \25513 , \25268 , \25272 );
xor \U$25170 ( \25514 , \25513 , \25277 );
and \U$25171 ( \25515 , \25511 , \25514 );
and \U$25172 ( \25516 , \25509 , \25514 );
or \U$25173 ( \25517 , \25512 , \25515 , \25516 );
xor \U$25174 ( \25518 , \25183 , \25187 );
xor \U$25175 ( \25519 , \25518 , \25192 );
xor \U$25176 ( \25520 , \25199 , \25203 );
xor \U$25177 ( \25521 , \25520 , \25208 );
and \U$25178 ( \25522 , \25519 , \25521 );
xor \U$25179 ( \25523 , \25216 , \25220 );
xor \U$25180 ( \25524 , \25523 , \25225 );
and \U$25181 ( \25525 , \25521 , \25524 );
and \U$25182 ( \25526 , \25519 , \25524 );
or \U$25183 ( \25527 , \25522 , \25525 , \25526 );
and \U$25184 ( \25528 , \25517 , \25527 );
xor \U$25185 ( \25529 , \25054 , \25058 );
xor \U$25186 ( \25530 , \25529 , \25063 );
and \U$25187 ( \25531 , \25527 , \25530 );
and \U$25188 ( \25532 , \25517 , \25530 );
or \U$25189 ( \25533 , \25528 , \25531 , \25532 );
and \U$25190 ( \25534 , \25507 , \25533 );
xor \U$25191 ( \25535 , \25038 , \25042 );
xor \U$25192 ( \25536 , \25535 , \25047 );
xor \U$25193 ( \25537 , \25322 , \25324 );
xor \U$25194 ( \25538 , \25537 , \25327 );
and \U$25195 ( \25539 , \25536 , \25538 );
xor \U$25196 ( \25540 , \25298 , \25300 );
xor \U$25197 ( \25541 , \25540 , \25303 );
and \U$25198 ( \25542 , \25538 , \25541 );
and \U$25199 ( \25543 , \25536 , \25541 );
or \U$25200 ( \25544 , \25539 , \25542 , \25543 );
and \U$25201 ( \25545 , \25533 , \25544 );
and \U$25202 ( \25546 , \25507 , \25544 );
or \U$25203 ( \25547 , \25534 , \25545 , \25546 );
xor \U$25204 ( \25548 , \25231 , \25283 );
xor \U$25205 ( \25549 , \25548 , \25306 );
xor \U$25206 ( \25550 , \25311 , \25313 );
xor \U$25207 ( \25551 , \25550 , \25316 );
and \U$25208 ( \25552 , \25549 , \25551 );
xor \U$25209 ( \25553 , \25330 , \25332 );
xor \U$25210 ( \25554 , \25553 , \25334 );
and \U$25211 ( \25555 , \25551 , \25554 );
and \U$25212 ( \25556 , \25549 , \25554 );
or \U$25213 ( \25557 , \25552 , \25555 , \25556 );
and \U$25214 ( \25558 , \25547 , \25557 );
xor \U$25215 ( \25559 , \25032 , \25086 );
xor \U$25216 ( \25560 , \25559 , \25108 );
and \U$25217 ( \25561 , \25557 , \25560 );
and \U$25218 ( \25562 , \25547 , \25560 );
or \U$25219 ( \25563 , \25558 , \25561 , \25562 );
xor \U$25220 ( \25564 , \25309 , \25319 );
xor \U$25221 ( \25565 , \25564 , \25337 );
xor \U$25222 ( \25566 , \25342 , \25344 );
xor \U$25223 ( \25567 , \25566 , \25347 );
and \U$25224 ( \25568 , \25565 , \25567 );
and \U$25225 ( \25569 , \25563 , \25568 );
xor \U$25226 ( \25570 , \25358 , \25360 );
xor \U$25227 ( \25571 , \25570 , \25363 );
and \U$25228 ( \25572 , \25568 , \25571 );
and \U$25229 ( \25573 , \25563 , \25571 );
or \U$25230 ( \25574 , \25569 , \25572 , \25573 );
xor \U$25231 ( \25575 , \25356 , \25366 );
xor \U$25232 ( \25576 , \25575 , \25369 );
and \U$25233 ( \25577 , \25574 , \25576 );
xor \U$25234 ( \25578 , \25146 , \25156 );
xor \U$25235 ( \25579 , \25578 , \25159 );
and \U$25236 ( \25580 , \25576 , \25579 );
and \U$25237 ( \25581 , \25574 , \25579 );
or \U$25238 ( \25582 , \25577 , \25580 , \25581 );
and \U$25239 ( \25583 , \25378 , \25582 );
xor \U$25240 ( \25584 , \25378 , \25582 );
xor \U$25241 ( \25585 , \25574 , \25576 );
xor \U$25242 ( \25586 , \25585 , \25579 );
and \U$25243 ( \25587 , \24836 , \21434 );
and \U$25244 ( \25588 , \24714 , \21432 );
nor \U$25245 ( \25589 , \25587 , \25588 );
xnor \U$25246 ( \25590 , \25589 , \21441 );
and \U$25247 ( \25591 , \25097 , \21450 );
and \U$25248 ( \25592 , \24841 , \21448 );
nor \U$25249 ( \25593 , \25591 , \25592 );
xnor \U$25250 ( \25594 , \25593 , \21457 );
and \U$25251 ( \25595 , \25590 , \25594 );
buf \U$25252 ( \25596 , RIbb328b0_169);
and \U$25253 ( \25597 , \25596 , \21469 );
and \U$25254 ( \25598 , \25294 , \21467 );
nor \U$25255 ( \25599 , \25597 , \25598 );
xnor \U$25256 ( \25600 , \25599 , \21476 );
and \U$25257 ( \25601 , \25594 , \25600 );
and \U$25258 ( \25602 , \25590 , \25600 );
or \U$25259 ( \25603 , \25595 , \25601 , \25602 );
buf \U$25260 ( \25604 , RIbb32928_170);
and \U$25261 ( \25605 , \25604 , \21464 );
buf \U$25262 ( \25606 , \25605 );
and \U$25263 ( \25607 , \25603 , \25606 );
and \U$25264 ( \25608 , \25596 , \21464 );
and \U$25265 ( \25609 , \25606 , \25608 );
and \U$25266 ( \25610 , \25603 , \25608 );
or \U$25267 ( \25611 , \25607 , \25609 , \25610 );
and \U$25268 ( \25612 , \21478 , \23421 );
and \U$25269 ( \25613 , \21463 , \23419 );
nor \U$25270 ( \25614 , \25612 , \25613 );
xnor \U$25271 ( \25615 , \25614 , \23279 );
and \U$25272 ( \25616 , \21750 , \23125 );
and \U$25273 ( \25617 , \21689 , \23123 );
nor \U$25274 ( \25618 , \25616 , \25617 );
xnor \U$25275 ( \25619 , \25618 , \22988 );
and \U$25276 ( \25620 , \25615 , \25619 );
and \U$25277 ( \25621 , \22011 , \22919 );
and \U$25278 ( \25622 , \21813 , \22917 );
nor \U$25279 ( \25623 , \25621 , \25622 );
xnor \U$25280 ( \25624 , \25623 , \22767 );
and \U$25281 ( \25625 , \25619 , \25624 );
and \U$25282 ( \25626 , \25615 , \25624 );
or \U$25283 ( \25627 , \25620 , \25625 , \25626 );
xor \U$25284 ( \25628 , \25034 , \25395 );
xor \U$25285 ( \25629 , \25395 , \25396 );
not \U$25286 ( \25630 , \25629 );
and \U$25287 ( \25631 , \25628 , \25630 );
and \U$25288 ( \25632 , \21387 , \25631 );
not \U$25289 ( \25633 , \25632 );
xnor \U$25290 ( \25634 , \25633 , \25399 );
and \U$25291 ( \25635 , \21403 , \25180 );
and \U$25292 ( \25636 , \21379 , \25178 );
nor \U$25293 ( \25637 , \25635 , \25636 );
xnor \U$25294 ( \25638 , \25637 , \25037 );
and \U$25295 ( \25639 , \25634 , \25638 );
and \U$25296 ( \25640 , \21421 , \24857 );
and \U$25297 ( \25641 , \21395 , \24855 );
nor \U$25298 ( \25642 , \25640 , \25641 );
xnor \U$25299 ( \25643 , \25642 , \24611 );
and \U$25300 ( \25644 , \25638 , \25643 );
and \U$25301 ( \25645 , \25634 , \25643 );
or \U$25302 ( \25646 , \25639 , \25644 , \25645 );
and \U$25303 ( \25647 , \25627 , \25646 );
and \U$25304 ( \25648 , \21436 , \24462 );
and \U$25305 ( \25649 , \21413 , \24460 );
nor \U$25306 ( \25650 , \25648 , \25649 );
xnor \U$25307 ( \25651 , \25650 , \24275 );
and \U$25308 ( \25652 , \21452 , \24149 );
and \U$25309 ( \25653 , \21428 , \24147 );
nor \U$25310 ( \25654 , \25652 , \25653 );
xnor \U$25311 ( \25655 , \25654 , \23944 );
and \U$25312 ( \25656 , \25651 , \25655 );
and \U$25313 ( \25657 , \21471 , \23743 );
and \U$25314 ( \25658 , \21444 , \23741 );
nor \U$25315 ( \25659 , \25657 , \25658 );
xnor \U$25316 ( \25660 , \25659 , \23594 );
and \U$25317 ( \25661 , \25655 , \25660 );
and \U$25318 ( \25662 , \25651 , \25660 );
or \U$25319 ( \25663 , \25656 , \25661 , \25662 );
and \U$25320 ( \25664 , \25646 , \25663 );
and \U$25321 ( \25665 , \25627 , \25663 );
or \U$25322 ( \25666 , \25647 , \25664 , \25665 );
and \U$25323 ( \25667 , \25611 , \25666 );
and \U$25324 ( \25668 , \23665 , \21385 );
and \U$25325 ( \25669 , \23491 , \21383 );
nor \U$25326 ( \25670 , \25668 , \25669 );
xnor \U$25327 ( \25671 , \25670 , \21392 );
and \U$25328 ( \25672 , \23970 , \21401 );
and \U$25329 ( \25673 , \23832 , \21399 );
nor \U$25330 ( \25674 , \25672 , \25673 );
xnor \U$25331 ( \25675 , \25674 , \21408 );
and \U$25332 ( \25676 , \25671 , \25675 );
and \U$25333 ( \25677 , \24506 , \21419 );
and \U$25334 ( \25678 , \24089 , \21417 );
nor \U$25335 ( \25679 , \25677 , \25678 );
xnor \U$25336 ( \25680 , \25679 , \21426 );
and \U$25337 ( \25681 , \25675 , \25680 );
and \U$25338 ( \25682 , \25671 , \25680 );
or \U$25339 ( \25683 , \25676 , \25681 , \25682 );
and \U$25340 ( \25684 , \22867 , \21985 );
and \U$25341 ( \25685 , \22624 , \21983 );
nor \U$25342 ( \25686 , \25684 , \25685 );
xnor \U$25343 ( \25687 , \25686 , \21907 );
and \U$25344 ( \25688 , \23058 , \21821 );
and \U$25345 ( \25689 , \22872 , \21819 );
nor \U$25346 ( \25690 , \25688 , \25689 );
xnor \U$25347 ( \25691 , \25690 , \21727 );
and \U$25348 ( \25692 , \25687 , \25691 );
and \U$25349 ( \25693 , \23466 , \21652 );
and \U$25350 ( \25694 , \23202 , \21650 );
nor \U$25351 ( \25695 , \25693 , \25694 );
xnor \U$25352 ( \25696 , \25695 , \21377 );
and \U$25353 ( \25697 , \25691 , \25696 );
and \U$25354 ( \25698 , \25687 , \25696 );
or \U$25355 ( \25699 , \25692 , \25697 , \25698 );
and \U$25356 ( \25700 , \25683 , \25699 );
and \U$25357 ( \25701 , \22204 , \22651 );
and \U$25358 ( \25702 , \22099 , \22649 );
nor \U$25359 ( \25703 , \25701 , \25702 );
xnor \U$25360 ( \25704 , \25703 , \22495 );
and \U$25361 ( \25705 , \22325 , \22379 );
and \U$25362 ( \25706 , \22209 , \22377 );
nor \U$25363 ( \25707 , \25705 , \25706 );
xnor \U$25364 ( \25708 , \25707 , \22266 );
and \U$25365 ( \25709 , \25704 , \25708 );
and \U$25366 ( \25710 , \22616 , \22185 );
and \U$25367 ( \25711 , \22440 , \22183 );
nor \U$25368 ( \25712 , \25710 , \25711 );
xnor \U$25369 ( \25713 , \25712 , \22049 );
and \U$25370 ( \25714 , \25708 , \25713 );
and \U$25371 ( \25715 , \25704 , \25713 );
or \U$25372 ( \25716 , \25709 , \25714 , \25715 );
and \U$25373 ( \25717 , \25699 , \25716 );
and \U$25374 ( \25718 , \25683 , \25716 );
or \U$25375 ( \25719 , \25700 , \25717 , \25718 );
and \U$25376 ( \25720 , \25666 , \25719 );
and \U$25377 ( \25721 , \25611 , \25719 );
or \U$25378 ( \25722 , \25667 , \25720 , \25721 );
xor \U$25379 ( \25723 , \25436 , \25440 );
xor \U$25380 ( \25724 , \25723 , \25445 );
xor \U$25381 ( \25725 , \25469 , \25473 );
xor \U$25382 ( \25726 , \25725 , \25478 );
and \U$25383 ( \25727 , \25724 , \25726 );
xor \U$25384 ( \25728 , \25489 , \25493 );
xor \U$25385 ( \25729 , \25728 , \25498 );
and \U$25386 ( \25730 , \25726 , \25729 );
and \U$25387 ( \25731 , \25724 , \25729 );
or \U$25388 ( \25732 , \25727 , \25730 , \25731 );
xor \U$25389 ( \25733 , \25382 , \25386 );
xor \U$25390 ( \25734 , \25733 , \25391 );
xor \U$25391 ( \25735 , \25452 , \25456 );
xor \U$25392 ( \25736 , \25735 , \25461 );
and \U$25393 ( \25737 , \25734 , \25736 );
xor \U$25394 ( \25738 , \25417 , \25421 );
xor \U$25395 ( \25739 , \25738 , \25426 );
and \U$25396 ( \25740 , \25736 , \25739 );
and \U$25397 ( \25741 , \25734 , \25739 );
or \U$25398 ( \25742 , \25737 , \25740 , \25741 );
and \U$25399 ( \25743 , \25732 , \25742 );
xor \U$25400 ( \25744 , \25519 , \25521 );
xor \U$25401 ( \25745 , \25744 , \25524 );
and \U$25402 ( \25746 , \25742 , \25745 );
and \U$25403 ( \25747 , \25732 , \25745 );
or \U$25404 ( \25748 , \25743 , \25746 , \25747 );
and \U$25405 ( \25749 , \25722 , \25748 );
xor \U$25406 ( \25750 , \25448 , \25464 );
xor \U$25407 ( \25751 , \25750 , \25481 );
xor \U$25408 ( \25752 , \25509 , \25511 );
xor \U$25409 ( \25753 , \25752 , \25514 );
and \U$25410 ( \25754 , \25751 , \25753 );
xnor \U$25411 ( \25755 , \25501 , \25503 );
and \U$25412 ( \25756 , \25753 , \25755 );
and \U$25413 ( \25757 , \25751 , \25755 );
or \U$25414 ( \25758 , \25754 , \25756 , \25757 );
and \U$25415 ( \25759 , \25748 , \25758 );
and \U$25416 ( \25760 , \25722 , \25758 );
or \U$25417 ( \25761 , \25749 , \25759 , \25760 );
xor \U$25418 ( \25762 , \25195 , \25211 );
xor \U$25419 ( \25763 , \25762 , \25228 );
xor \U$25420 ( \25764 , \25247 , \25263 );
xor \U$25421 ( \25765 , \25764 , \25280 );
and \U$25422 ( \25766 , \25763 , \25765 );
xor \U$25423 ( \25767 , \25536 , \25538 );
xor \U$25424 ( \25768 , \25767 , \25541 );
and \U$25425 ( \25769 , \25765 , \25768 );
and \U$25426 ( \25770 , \25763 , \25768 );
or \U$25427 ( \25771 , \25766 , \25769 , \25770 );
and \U$25428 ( \25772 , \25761 , \25771 );
xor \U$25429 ( \25773 , \25549 , \25551 );
xor \U$25430 ( \25774 , \25773 , \25554 );
and \U$25431 ( \25775 , \25771 , \25774 );
and \U$25432 ( \25776 , \25761 , \25774 );
or \U$25433 ( \25777 , \25772 , \25775 , \25776 );
xor \U$25434 ( \25778 , \25547 , \25557 );
xor \U$25435 ( \25779 , \25778 , \25560 );
and \U$25436 ( \25780 , \25777 , \25779 );
xor \U$25437 ( \25781 , \25565 , \25567 );
and \U$25438 ( \25782 , \25779 , \25781 );
and \U$25439 ( \25783 , \25777 , \25781 );
or \U$25440 ( \25784 , \25780 , \25782 , \25783 );
xor \U$25441 ( \25785 , \25340 , \25350 );
xor \U$25442 ( \25786 , \25785 , \25353 );
and \U$25443 ( \25787 , \25784 , \25786 );
xor \U$25444 ( \25788 , \25563 , \25568 );
xor \U$25445 ( \25789 , \25788 , \25571 );
and \U$25446 ( \25790 , \25786 , \25789 );
and \U$25447 ( \25791 , \25784 , \25789 );
or \U$25448 ( \25792 , \25787 , \25790 , \25791 );
and \U$25449 ( \25793 , \25586 , \25792 );
xor \U$25450 ( \25794 , \25586 , \25792 );
xor \U$25451 ( \25795 , \25784 , \25786 );
xor \U$25452 ( \25796 , \25795 , \25789 );
and \U$25453 ( \25797 , \21463 , \23743 );
and \U$25454 ( \25798 , \21471 , \23741 );
nor \U$25455 ( \25799 , \25797 , \25798 );
xnor \U$25456 ( \25800 , \25799 , \23594 );
and \U$25457 ( \25801 , \21689 , \23421 );
and \U$25458 ( \25802 , \21478 , \23419 );
nor \U$25459 ( \25803 , \25801 , \25802 );
xnor \U$25460 ( \25804 , \25803 , \23279 );
and \U$25461 ( \25805 , \25800 , \25804 );
and \U$25462 ( \25806 , \21813 , \23125 );
and \U$25463 ( \25807 , \21750 , \23123 );
nor \U$25464 ( \25808 , \25806 , \25807 );
xnor \U$25465 ( \25809 , \25808 , \22988 );
and \U$25466 ( \25810 , \25804 , \25809 );
and \U$25467 ( \25811 , \25800 , \25809 );
or \U$25468 ( \25812 , \25805 , \25810 , \25811 );
buf \U$25469 ( \25813 , RIbb2e1e8_44);
buf \U$25470 ( \25814 , RIbb2e170_45);
and \U$25471 ( \25815 , \25813 , \25814 );
not \U$25472 ( \25816 , \25815 );
and \U$25473 ( \25817 , \25396 , \25816 );
not \U$25474 ( \25818 , \25817 );
and \U$25475 ( \25819 , \21379 , \25631 );
and \U$25476 ( \25820 , \21387 , \25629 );
nor \U$25477 ( \25821 , \25819 , \25820 );
xnor \U$25478 ( \25822 , \25821 , \25399 );
and \U$25479 ( \25823 , \25818 , \25822 );
and \U$25480 ( \25824 , \21395 , \25180 );
and \U$25481 ( \25825 , \21403 , \25178 );
nor \U$25482 ( \25826 , \25824 , \25825 );
xnor \U$25483 ( \25827 , \25826 , \25037 );
and \U$25484 ( \25828 , \25822 , \25827 );
and \U$25485 ( \25829 , \25818 , \25827 );
or \U$25486 ( \25830 , \25823 , \25828 , \25829 );
and \U$25487 ( \25831 , \25812 , \25830 );
and \U$25488 ( \25832 , \21413 , \24857 );
and \U$25489 ( \25833 , \21421 , \24855 );
nor \U$25490 ( \25834 , \25832 , \25833 );
xnor \U$25491 ( \25835 , \25834 , \24611 );
and \U$25492 ( \25836 , \21428 , \24462 );
and \U$25493 ( \25837 , \21436 , \24460 );
nor \U$25494 ( \25838 , \25836 , \25837 );
xnor \U$25495 ( \25839 , \25838 , \24275 );
and \U$25496 ( \25840 , \25835 , \25839 );
and \U$25497 ( \25841 , \21444 , \24149 );
and \U$25498 ( \25842 , \21452 , \24147 );
nor \U$25499 ( \25843 , \25841 , \25842 );
xnor \U$25500 ( \25844 , \25843 , \23944 );
and \U$25501 ( \25845 , \25839 , \25844 );
and \U$25502 ( \25846 , \25835 , \25844 );
or \U$25503 ( \25847 , \25840 , \25845 , \25846 );
and \U$25504 ( \25848 , \25830 , \25847 );
and \U$25505 ( \25849 , \25812 , \25847 );
or \U$25506 ( \25850 , \25831 , \25848 , \25849 );
and \U$25507 ( \25851 , \22099 , \22919 );
and \U$25508 ( \25852 , \22011 , \22917 );
nor \U$25509 ( \25853 , \25851 , \25852 );
xnor \U$25510 ( \25854 , \25853 , \22767 );
and \U$25511 ( \25855 , \22209 , \22651 );
and \U$25512 ( \25856 , \22204 , \22649 );
nor \U$25513 ( \25857 , \25855 , \25856 );
xnor \U$25514 ( \25858 , \25857 , \22495 );
and \U$25515 ( \25859 , \25854 , \25858 );
and \U$25516 ( \25860 , \22440 , \22379 );
and \U$25517 ( \25861 , \22325 , \22377 );
nor \U$25518 ( \25862 , \25860 , \25861 );
xnor \U$25519 ( \25863 , \25862 , \22266 );
and \U$25520 ( \25864 , \25858 , \25863 );
and \U$25521 ( \25865 , \25854 , \25863 );
or \U$25522 ( \25866 , \25859 , \25864 , \25865 );
and \U$25523 ( \25867 , \23491 , \21652 );
and \U$25524 ( \25868 , \23466 , \21650 );
nor \U$25525 ( \25869 , \25867 , \25868 );
xnor \U$25526 ( \25870 , \25869 , \21377 );
and \U$25527 ( \25871 , \23832 , \21385 );
and \U$25528 ( \25872 , \23665 , \21383 );
nor \U$25529 ( \25873 , \25871 , \25872 );
xnor \U$25530 ( \25874 , \25873 , \21392 );
and \U$25531 ( \25875 , \25870 , \25874 );
and \U$25532 ( \25876 , \24089 , \21401 );
and \U$25533 ( \25877 , \23970 , \21399 );
nor \U$25534 ( \25878 , \25876 , \25877 );
xnor \U$25535 ( \25879 , \25878 , \21408 );
and \U$25536 ( \25880 , \25874 , \25879 );
and \U$25537 ( \25881 , \25870 , \25879 );
or \U$25538 ( \25882 , \25875 , \25880 , \25881 );
and \U$25539 ( \25883 , \25866 , \25882 );
and \U$25540 ( \25884 , \22624 , \22185 );
and \U$25541 ( \25885 , \22616 , \22183 );
nor \U$25542 ( \25886 , \25884 , \25885 );
xnor \U$25543 ( \25887 , \25886 , \22049 );
and \U$25544 ( \25888 , \22872 , \21985 );
and \U$25545 ( \25889 , \22867 , \21983 );
nor \U$25546 ( \25890 , \25888 , \25889 );
xnor \U$25547 ( \25891 , \25890 , \21907 );
and \U$25548 ( \25892 , \25887 , \25891 );
and \U$25549 ( \25893 , \23202 , \21821 );
and \U$25550 ( \25894 , \23058 , \21819 );
nor \U$25551 ( \25895 , \25893 , \25894 );
xnor \U$25552 ( \25896 , \25895 , \21727 );
and \U$25553 ( \25897 , \25891 , \25896 );
and \U$25554 ( \25898 , \25887 , \25896 );
or \U$25555 ( \25899 , \25892 , \25897 , \25898 );
and \U$25556 ( \25900 , \25882 , \25899 );
and \U$25557 ( \25901 , \25866 , \25899 );
or \U$25558 ( \25902 , \25883 , \25900 , \25901 );
and \U$25559 ( \25903 , \25850 , \25902 );
and \U$25560 ( \25904 , \24714 , \21419 );
and \U$25561 ( \25905 , \24506 , \21417 );
nor \U$25562 ( \25906 , \25904 , \25905 );
xnor \U$25563 ( \25907 , \25906 , \21426 );
and \U$25564 ( \25908 , \24841 , \21434 );
and \U$25565 ( \25909 , \24836 , \21432 );
nor \U$25566 ( \25910 , \25908 , \25909 );
xnor \U$25567 ( \25911 , \25910 , \21441 );
and \U$25568 ( \25912 , \25907 , \25911 );
and \U$25569 ( \25913 , \25294 , \21450 );
and \U$25570 ( \25914 , \25097 , \21448 );
nor \U$25571 ( \25915 , \25913 , \25914 );
xnor \U$25572 ( \25916 , \25915 , \21457 );
and \U$25573 ( \25917 , \25911 , \25916 );
and \U$25574 ( \25918 , \25907 , \25916 );
or \U$25575 ( \25919 , \25912 , \25917 , \25918 );
xor \U$25576 ( \25920 , \25590 , \25594 );
xor \U$25577 ( \25921 , \25920 , \25600 );
and \U$25578 ( \25922 , \25919 , \25921 );
not \U$25579 ( \25923 , \25605 );
and \U$25580 ( \25924 , \25921 , \25923 );
and \U$25581 ( \25925 , \25919 , \25923 );
or \U$25582 ( \25926 , \25922 , \25924 , \25925 );
and \U$25583 ( \25927 , \25902 , \25926 );
and \U$25584 ( \25928 , \25850 , \25926 );
or \U$25585 ( \25929 , \25903 , \25927 , \25928 );
xor \U$25586 ( \25930 , \25671 , \25675 );
xor \U$25587 ( \25931 , \25930 , \25680 );
xor \U$25588 ( \25932 , \25687 , \25691 );
xor \U$25589 ( \25933 , \25932 , \25696 );
and \U$25590 ( \25934 , \25931 , \25933 );
xor \U$25591 ( \25935 , \25704 , \25708 );
xor \U$25592 ( \25936 , \25935 , \25713 );
and \U$25593 ( \25937 , \25933 , \25936 );
and \U$25594 ( \25938 , \25931 , \25936 );
or \U$25595 ( \25939 , \25934 , \25937 , \25938 );
xor \U$25596 ( \25940 , \25615 , \25619 );
xor \U$25597 ( \25941 , \25940 , \25624 );
xor \U$25598 ( \25942 , \25634 , \25638 );
xor \U$25599 ( \25943 , \25942 , \25643 );
and \U$25600 ( \25944 , \25941 , \25943 );
xor \U$25601 ( \25945 , \25651 , \25655 );
xor \U$25602 ( \25946 , \25945 , \25660 );
and \U$25603 ( \25947 , \25943 , \25946 );
and \U$25604 ( \25948 , \25941 , \25946 );
or \U$25605 ( \25949 , \25944 , \25947 , \25948 );
and \U$25606 ( \25950 , \25939 , \25949 );
xor \U$25607 ( \25951 , \25400 , \25404 );
xor \U$25608 ( \25952 , \25951 , \25409 );
and \U$25609 ( \25953 , \25949 , \25952 );
and \U$25610 ( \25954 , \25939 , \25952 );
or \U$25611 ( \25955 , \25950 , \25953 , \25954 );
and \U$25612 ( \25956 , \25929 , \25955 );
xor \U$25613 ( \25957 , \25603 , \25606 );
xor \U$25614 ( \25958 , \25957 , \25608 );
xor \U$25615 ( \25959 , \25724 , \25726 );
xor \U$25616 ( \25960 , \25959 , \25729 );
and \U$25617 ( \25961 , \25958 , \25960 );
xor \U$25618 ( \25962 , \25734 , \25736 );
xor \U$25619 ( \25963 , \25962 , \25739 );
and \U$25620 ( \25964 , \25960 , \25963 );
and \U$25621 ( \25965 , \25958 , \25963 );
or \U$25622 ( \25966 , \25961 , \25964 , \25965 );
and \U$25623 ( \25967 , \25955 , \25966 );
and \U$25624 ( \25968 , \25929 , \25966 );
or \U$25625 ( \25969 , \25956 , \25967 , \25968 );
xor \U$25626 ( \25970 , \25394 , \25412 );
xor \U$25627 ( \25971 , \25970 , \25429 );
xor \U$25628 ( \25972 , \25732 , \25742 );
xor \U$25629 ( \25973 , \25972 , \25745 );
and \U$25630 ( \25974 , \25971 , \25973 );
xor \U$25631 ( \25975 , \25751 , \25753 );
xor \U$25632 ( \25976 , \25975 , \25755 );
and \U$25633 ( \25977 , \25973 , \25976 );
and \U$25634 ( \25978 , \25971 , \25976 );
or \U$25635 ( \25979 , \25974 , \25977 , \25978 );
and \U$25636 ( \25980 , \25969 , \25979 );
xor \U$25637 ( \25981 , \25517 , \25527 );
xor \U$25638 ( \25982 , \25981 , \25530 );
and \U$25639 ( \25983 , \25979 , \25982 );
and \U$25640 ( \25984 , \25969 , \25982 );
or \U$25641 ( \25985 , \25980 , \25983 , \25984 );
xor \U$25642 ( \25986 , \25432 , \25484 );
xor \U$25643 ( \25987 , \25986 , \25504 );
xor \U$25644 ( \25988 , \25722 , \25748 );
xor \U$25645 ( \25989 , \25988 , \25758 );
and \U$25646 ( \25990 , \25987 , \25989 );
xor \U$25647 ( \25991 , \25763 , \25765 );
xor \U$25648 ( \25992 , \25991 , \25768 );
and \U$25649 ( \25993 , \25989 , \25992 );
and \U$25650 ( \25994 , \25987 , \25992 );
or \U$25651 ( \25995 , \25990 , \25993 , \25994 );
and \U$25652 ( \25996 , \25985 , \25995 );
xor \U$25653 ( \25997 , \25507 , \25533 );
xor \U$25654 ( \25998 , \25997 , \25544 );
and \U$25655 ( \25999 , \25995 , \25998 );
and \U$25656 ( \26000 , \25985 , \25998 );
or \U$25657 ( \26001 , \25996 , \25999 , \26000 );
xor \U$25658 ( \26002 , \25396 , \25813 );
xor \U$25659 ( \26003 , \25813 , \25814 );
not \U$25660 ( \26004 , \26003 );
and \U$25661 ( \26005 , \26002 , \26004 );
and \U$25662 ( \26006 , \21387 , \26005 );
not \U$25663 ( \26007 , \26006 );
xnor \U$25664 ( \26008 , \26007 , \25817 );
and \U$25665 ( \26009 , \21403 , \25631 );
and \U$25666 ( \26010 , \21379 , \25629 );
nor \U$25667 ( \26011 , \26009 , \26010 );
xnor \U$25668 ( \26012 , \26011 , \25399 );
and \U$25669 ( \26013 , \26008 , \26012 );
and \U$25670 ( \26014 , \21421 , \25180 );
and \U$25671 ( \26015 , \21395 , \25178 );
nor \U$25672 ( \26016 , \26014 , \26015 );
xnor \U$25673 ( \26017 , \26016 , \25037 );
and \U$25674 ( \26018 , \26012 , \26017 );
and \U$25675 ( \26019 , \26008 , \26017 );
or \U$25676 ( \26020 , \26013 , \26018 , \26019 );
and \U$25677 ( \26021 , \21478 , \23743 );
and \U$25678 ( \26022 , \21463 , \23741 );
nor \U$25679 ( \26023 , \26021 , \26022 );
xnor \U$25680 ( \26024 , \26023 , \23594 );
and \U$25681 ( \26025 , \21750 , \23421 );
and \U$25682 ( \26026 , \21689 , \23419 );
nor \U$25683 ( \26027 , \26025 , \26026 );
xnor \U$25684 ( \26028 , \26027 , \23279 );
and \U$25685 ( \26029 , \26024 , \26028 );
and \U$25686 ( \26030 , \22011 , \23125 );
and \U$25687 ( \26031 , \21813 , \23123 );
nor \U$25688 ( \26032 , \26030 , \26031 );
xnor \U$25689 ( \26033 , \26032 , \22988 );
and \U$25690 ( \26034 , \26028 , \26033 );
and \U$25691 ( \26035 , \26024 , \26033 );
or \U$25692 ( \26036 , \26029 , \26034 , \26035 );
and \U$25693 ( \26037 , \26020 , \26036 );
and \U$25694 ( \26038 , \21436 , \24857 );
and \U$25695 ( \26039 , \21413 , \24855 );
nor \U$25696 ( \26040 , \26038 , \26039 );
xnor \U$25697 ( \26041 , \26040 , \24611 );
and \U$25698 ( \26042 , \21452 , \24462 );
and \U$25699 ( \26043 , \21428 , \24460 );
nor \U$25700 ( \26044 , \26042 , \26043 );
xnor \U$25701 ( \26045 , \26044 , \24275 );
and \U$25702 ( \26046 , \26041 , \26045 );
and \U$25703 ( \26047 , \21471 , \24149 );
and \U$25704 ( \26048 , \21444 , \24147 );
nor \U$25705 ( \26049 , \26047 , \26048 );
xnor \U$25706 ( \26050 , \26049 , \23944 );
and \U$25707 ( \26051 , \26045 , \26050 );
and \U$25708 ( \26052 , \26041 , \26050 );
or \U$25709 ( \26053 , \26046 , \26051 , \26052 );
and \U$25710 ( \26054 , \26036 , \26053 );
and \U$25711 ( \26055 , \26020 , \26053 );
or \U$25712 ( \26056 , \26037 , \26054 , \26055 );
and \U$25713 ( \26057 , \24836 , \21419 );
and \U$25714 ( \26058 , \24714 , \21417 );
nor \U$25715 ( \26059 , \26057 , \26058 );
xnor \U$25716 ( \26060 , \26059 , \21426 );
and \U$25717 ( \26061 , \25097 , \21434 );
and \U$25718 ( \26062 , \24841 , \21432 );
nor \U$25719 ( \26063 , \26061 , \26062 );
xnor \U$25720 ( \26064 , \26063 , \21441 );
and \U$25721 ( \26065 , \26060 , \26064 );
and \U$25722 ( \26066 , \25596 , \21450 );
and \U$25723 ( \26067 , \25294 , \21448 );
nor \U$25724 ( \26068 , \26066 , \26067 );
xnor \U$25725 ( \26069 , \26068 , \21457 );
and \U$25726 ( \26070 , \26064 , \26069 );
and \U$25727 ( \26071 , \26060 , \26069 );
or \U$25728 ( \26072 , \26065 , \26070 , \26071 );
buf \U$25729 ( \26073 , RIbb329a0_171);
and \U$25730 ( \26074 , \26073 , \21469 );
and \U$25731 ( \26075 , \25604 , \21467 );
nor \U$25732 ( \26076 , \26074 , \26075 );
xnor \U$25733 ( \26077 , \26076 , \21476 );
buf \U$25734 ( \26078 , RIbb32a18_172);
and \U$25735 ( \26079 , \26078 , \21464 );
or \U$25736 ( \26080 , \26077 , \26079 );
and \U$25737 ( \26081 , \26072 , \26080 );
and \U$25738 ( \26082 , \25604 , \21469 );
and \U$25739 ( \26083 , \25596 , \21467 );
nor \U$25740 ( \26084 , \26082 , \26083 );
xnor \U$25741 ( \26085 , \26084 , \21476 );
and \U$25742 ( \26086 , \26080 , \26085 );
and \U$25743 ( \26087 , \26072 , \26085 );
or \U$25744 ( \26088 , \26081 , \26086 , \26087 );
and \U$25745 ( \26089 , \26056 , \26088 );
and \U$25746 ( \26090 , \22204 , \22919 );
and \U$25747 ( \26091 , \22099 , \22917 );
nor \U$25748 ( \26092 , \26090 , \26091 );
xnor \U$25749 ( \26093 , \26092 , \22767 );
and \U$25750 ( \26094 , \22325 , \22651 );
and \U$25751 ( \26095 , \22209 , \22649 );
nor \U$25752 ( \26096 , \26094 , \26095 );
xnor \U$25753 ( \26097 , \26096 , \22495 );
and \U$25754 ( \26098 , \26093 , \26097 );
and \U$25755 ( \26099 , \22616 , \22379 );
and \U$25756 ( \26100 , \22440 , \22377 );
nor \U$25757 ( \26101 , \26099 , \26100 );
xnor \U$25758 ( \26102 , \26101 , \22266 );
and \U$25759 ( \26103 , \26097 , \26102 );
and \U$25760 ( \26104 , \26093 , \26102 );
or \U$25761 ( \26105 , \26098 , \26103 , \26104 );
and \U$25762 ( \26106 , \22867 , \22185 );
and \U$25763 ( \26107 , \22624 , \22183 );
nor \U$25764 ( \26108 , \26106 , \26107 );
xnor \U$25765 ( \26109 , \26108 , \22049 );
and \U$25766 ( \26110 , \23058 , \21985 );
and \U$25767 ( \26111 , \22872 , \21983 );
nor \U$25768 ( \26112 , \26110 , \26111 );
xnor \U$25769 ( \26113 , \26112 , \21907 );
and \U$25770 ( \26114 , \26109 , \26113 );
and \U$25771 ( \26115 , \23466 , \21821 );
and \U$25772 ( \26116 , \23202 , \21819 );
nor \U$25773 ( \26117 , \26115 , \26116 );
xnor \U$25774 ( \26118 , \26117 , \21727 );
and \U$25775 ( \26119 , \26113 , \26118 );
and \U$25776 ( \26120 , \26109 , \26118 );
or \U$25777 ( \26121 , \26114 , \26119 , \26120 );
and \U$25778 ( \26122 , \26105 , \26121 );
and \U$25779 ( \26123 , \23665 , \21652 );
and \U$25780 ( \26124 , \23491 , \21650 );
nor \U$25781 ( \26125 , \26123 , \26124 );
xnor \U$25782 ( \26126 , \26125 , \21377 );
and \U$25783 ( \26127 , \23970 , \21385 );
and \U$25784 ( \26128 , \23832 , \21383 );
nor \U$25785 ( \26129 , \26127 , \26128 );
xnor \U$25786 ( \26130 , \26129 , \21392 );
and \U$25787 ( \26131 , \26126 , \26130 );
and \U$25788 ( \26132 , \24506 , \21401 );
and \U$25789 ( \26133 , \24089 , \21399 );
nor \U$25790 ( \26134 , \26132 , \26133 );
xnor \U$25791 ( \26135 , \26134 , \21408 );
and \U$25792 ( \26136 , \26130 , \26135 );
and \U$25793 ( \26137 , \26126 , \26135 );
or \U$25794 ( \26138 , \26131 , \26136 , \26137 );
and \U$25795 ( \26139 , \26121 , \26138 );
and \U$25796 ( \26140 , \26105 , \26138 );
or \U$25797 ( \26141 , \26122 , \26139 , \26140 );
and \U$25798 ( \26142 , \26088 , \26141 );
and \U$25799 ( \26143 , \26056 , \26141 );
or \U$25800 ( \26144 , \26089 , \26142 , \26143 );
and \U$25801 ( \26145 , \26073 , \21464 );
xor \U$25802 ( \26146 , \25907 , \25911 );
xor \U$25803 ( \26147 , \26146 , \25916 );
and \U$25804 ( \26148 , \26145 , \26147 );
xor \U$25805 ( \26149 , \25870 , \25874 );
xor \U$25806 ( \26150 , \26149 , \25879 );
and \U$25807 ( \26151 , \26147 , \26150 );
and \U$25808 ( \26152 , \26145 , \26150 );
or \U$25809 ( \26153 , \26148 , \26151 , \26152 );
xor \U$25810 ( \26154 , \25854 , \25858 );
xor \U$25811 ( \26155 , \26154 , \25863 );
xor \U$25812 ( \26156 , \25800 , \25804 );
xor \U$25813 ( \26157 , \26156 , \25809 );
and \U$25814 ( \26158 , \26155 , \26157 );
xor \U$25815 ( \26159 , \25887 , \25891 );
xor \U$25816 ( \26160 , \26159 , \25896 );
and \U$25817 ( \26161 , \26157 , \26160 );
and \U$25818 ( \26162 , \26155 , \26160 );
or \U$25819 ( \26163 , \26158 , \26161 , \26162 );
and \U$25820 ( \26164 , \26153 , \26163 );
xor \U$25821 ( \26165 , \25941 , \25943 );
xor \U$25822 ( \26166 , \26165 , \25946 );
and \U$25823 ( \26167 , \26163 , \26166 );
and \U$25824 ( \26168 , \26153 , \26166 );
or \U$25825 ( \26169 , \26164 , \26167 , \26168 );
and \U$25826 ( \26170 , \26144 , \26169 );
xor \U$25827 ( \26171 , \25866 , \25882 );
xor \U$25828 ( \26172 , \26171 , \25899 );
xor \U$25829 ( \26173 , \25931 , \25933 );
xor \U$25830 ( \26174 , \26173 , \25936 );
and \U$25831 ( \26175 , \26172 , \26174 );
xor \U$25832 ( \26176 , \25919 , \25921 );
xor \U$25833 ( \26177 , \26176 , \25923 );
and \U$25834 ( \26178 , \26174 , \26177 );
and \U$25835 ( \26179 , \26172 , \26177 );
or \U$25836 ( \26180 , \26175 , \26178 , \26179 );
and \U$25837 ( \26181 , \26169 , \26180 );
and \U$25838 ( \26182 , \26144 , \26180 );
or \U$25839 ( \26183 , \26170 , \26181 , \26182 );
xor \U$25840 ( \26184 , \25627 , \25646 );
xor \U$25841 ( \26185 , \26184 , \25663 );
xor \U$25842 ( \26186 , \25683 , \25699 );
xor \U$25843 ( \26187 , \26186 , \25716 );
and \U$25844 ( \26188 , \26185 , \26187 );
xor \U$25845 ( \26189 , \25958 , \25960 );
xor \U$25846 ( \26190 , \26189 , \25963 );
and \U$25847 ( \26191 , \26187 , \26190 );
and \U$25848 ( \26192 , \26185 , \26190 );
or \U$25849 ( \26193 , \26188 , \26191 , \26192 );
and \U$25850 ( \26194 , \26183 , \26193 );
xor \U$25851 ( \26195 , \25611 , \25666 );
xor \U$25852 ( \26196 , \26195 , \25719 );
and \U$25853 ( \26197 , \26193 , \26196 );
and \U$25854 ( \26198 , \26183 , \26196 );
or \U$25855 ( \26199 , \26194 , \26197 , \26198 );
xor \U$25856 ( \26200 , \25969 , \25979 );
xor \U$25857 ( \26201 , \26200 , \25982 );
and \U$25858 ( \26202 , \26199 , \26201 );
xor \U$25859 ( \26203 , \25987 , \25989 );
xor \U$25860 ( \26204 , \26203 , \25992 );
and \U$25861 ( \26205 , \26201 , \26204 );
and \U$25862 ( \26206 , \26199 , \26204 );
or \U$25863 ( \26207 , \26202 , \26205 , \26206 );
xor \U$25864 ( \26208 , \25985 , \25995 );
xor \U$25865 ( \26209 , \26208 , \25998 );
and \U$25866 ( \26210 , \26207 , \26209 );
xor \U$25867 ( \26211 , \25761 , \25771 );
xor \U$25868 ( \26212 , \26211 , \25774 );
and \U$25869 ( \26213 , \26209 , \26212 );
and \U$25870 ( \26214 , \26207 , \26212 );
or \U$25871 ( \26215 , \26210 , \26213 , \26214 );
and \U$25872 ( \26216 , \26001 , \26215 );
xor \U$25873 ( \26217 , \25777 , \25779 );
xor \U$25874 ( \26218 , \26217 , \25781 );
and \U$25875 ( \26219 , \26215 , \26218 );
and \U$25876 ( \26220 , \26001 , \26218 );
or \U$25877 ( \26221 , \26216 , \26219 , \26220 );
and \U$25878 ( \26222 , \25796 , \26221 );
xor \U$25879 ( \26223 , \25796 , \26221 );
xor \U$25880 ( \26224 , \26001 , \26215 );
xor \U$25881 ( \26225 , \26224 , \26218 );
buf \U$25882 ( \26226 , RIbb2e0f8_46);
buf \U$25883 ( \26227 , RIbb2e080_47);
and \U$25884 ( \26228 , \26226 , \26227 );
not \U$25885 ( \26229 , \26228 );
and \U$25886 ( \26230 , \25814 , \26229 );
not \U$25887 ( \26231 , \26230 );
and \U$25888 ( \26232 , \21379 , \26005 );
and \U$25889 ( \26233 , \21387 , \26003 );
nor \U$25890 ( \26234 , \26232 , \26233 );
xnor \U$25891 ( \26235 , \26234 , \25817 );
and \U$25892 ( \26236 , \26231 , \26235 );
and \U$25893 ( \26237 , \21395 , \25631 );
and \U$25894 ( \26238 , \21403 , \25629 );
nor \U$25895 ( \26239 , \26237 , \26238 );
xnor \U$25896 ( \26240 , \26239 , \25399 );
and \U$25897 ( \26241 , \26235 , \26240 );
and \U$25898 ( \26242 , \26231 , \26240 );
or \U$25899 ( \26243 , \26236 , \26241 , \26242 );
and \U$25900 ( \26244 , \21413 , \25180 );
and \U$25901 ( \26245 , \21421 , \25178 );
nor \U$25902 ( \26246 , \26244 , \26245 );
xnor \U$25903 ( \26247 , \26246 , \25037 );
and \U$25904 ( \26248 , \21428 , \24857 );
and \U$25905 ( \26249 , \21436 , \24855 );
nor \U$25906 ( \26250 , \26248 , \26249 );
xnor \U$25907 ( \26251 , \26250 , \24611 );
and \U$25908 ( \26252 , \26247 , \26251 );
and \U$25909 ( \26253 , \21444 , \24462 );
and \U$25910 ( \26254 , \21452 , \24460 );
nor \U$25911 ( \26255 , \26253 , \26254 );
xnor \U$25912 ( \26256 , \26255 , \24275 );
and \U$25913 ( \26257 , \26251 , \26256 );
and \U$25914 ( \26258 , \26247 , \26256 );
or \U$25915 ( \26259 , \26252 , \26257 , \26258 );
and \U$25916 ( \26260 , \26243 , \26259 );
and \U$25917 ( \26261 , \21463 , \24149 );
and \U$25918 ( \26262 , \21471 , \24147 );
nor \U$25919 ( \26263 , \26261 , \26262 );
xnor \U$25920 ( \26264 , \26263 , \23944 );
and \U$25921 ( \26265 , \21689 , \23743 );
and \U$25922 ( \26266 , \21478 , \23741 );
nor \U$25923 ( \26267 , \26265 , \26266 );
xnor \U$25924 ( \26268 , \26267 , \23594 );
and \U$25925 ( \26269 , \26264 , \26268 );
and \U$25926 ( \26270 , \21813 , \23421 );
and \U$25927 ( \26271 , \21750 , \23419 );
nor \U$25928 ( \26272 , \26270 , \26271 );
xnor \U$25929 ( \26273 , \26272 , \23279 );
and \U$25930 ( \26274 , \26268 , \26273 );
and \U$25931 ( \26275 , \26264 , \26273 );
or \U$25932 ( \26276 , \26269 , \26274 , \26275 );
and \U$25933 ( \26277 , \26259 , \26276 );
and \U$25934 ( \26278 , \26243 , \26276 );
or \U$25935 ( \26279 , \26260 , \26277 , \26278 );
and \U$25936 ( \26280 , \22099 , \23125 );
and \U$25937 ( \26281 , \22011 , \23123 );
nor \U$25938 ( \26282 , \26280 , \26281 );
xnor \U$25939 ( \26283 , \26282 , \22988 );
and \U$25940 ( \26284 , \22209 , \22919 );
and \U$25941 ( \26285 , \22204 , \22917 );
nor \U$25942 ( \26286 , \26284 , \26285 );
xnor \U$25943 ( \26287 , \26286 , \22767 );
and \U$25944 ( \26288 , \26283 , \26287 );
and \U$25945 ( \26289 , \22440 , \22651 );
and \U$25946 ( \26290 , \22325 , \22649 );
nor \U$25947 ( \26291 , \26289 , \26290 );
xnor \U$25948 ( \26292 , \26291 , \22495 );
and \U$25949 ( \26293 , \26287 , \26292 );
and \U$25950 ( \26294 , \26283 , \26292 );
or \U$25951 ( \26295 , \26288 , \26293 , \26294 );
and \U$25952 ( \26296 , \22624 , \22379 );
and \U$25953 ( \26297 , \22616 , \22377 );
nor \U$25954 ( \26298 , \26296 , \26297 );
xnor \U$25955 ( \26299 , \26298 , \22266 );
and \U$25956 ( \26300 , \22872 , \22185 );
and \U$25957 ( \26301 , \22867 , \22183 );
nor \U$25958 ( \26302 , \26300 , \26301 );
xnor \U$25959 ( \26303 , \26302 , \22049 );
and \U$25960 ( \26304 , \26299 , \26303 );
and \U$25961 ( \26305 , \23202 , \21985 );
and \U$25962 ( \26306 , \23058 , \21983 );
nor \U$25963 ( \26307 , \26305 , \26306 );
xnor \U$25964 ( \26308 , \26307 , \21907 );
and \U$25965 ( \26309 , \26303 , \26308 );
and \U$25966 ( \26310 , \26299 , \26308 );
or \U$25967 ( \26311 , \26304 , \26309 , \26310 );
and \U$25968 ( \26312 , \26295 , \26311 );
and \U$25969 ( \26313 , \23491 , \21821 );
and \U$25970 ( \26314 , \23466 , \21819 );
nor \U$25971 ( \26315 , \26313 , \26314 );
xnor \U$25972 ( \26316 , \26315 , \21727 );
and \U$25973 ( \26317 , \23832 , \21652 );
and \U$25974 ( \26318 , \23665 , \21650 );
nor \U$25975 ( \26319 , \26317 , \26318 );
xnor \U$25976 ( \26320 , \26319 , \21377 );
and \U$25977 ( \26321 , \26316 , \26320 );
and \U$25978 ( \26322 , \24089 , \21385 );
and \U$25979 ( \26323 , \23970 , \21383 );
nor \U$25980 ( \26324 , \26322 , \26323 );
xnor \U$25981 ( \26325 , \26324 , \21392 );
and \U$25982 ( \26326 , \26320 , \26325 );
and \U$25983 ( \26327 , \26316 , \26325 );
or \U$25984 ( \26328 , \26321 , \26326 , \26327 );
and \U$25985 ( \26329 , \26311 , \26328 );
and \U$25986 ( \26330 , \26295 , \26328 );
or \U$25987 ( \26331 , \26312 , \26329 , \26330 );
and \U$25988 ( \26332 , \26279 , \26331 );
and \U$25989 ( \26333 , \25604 , \21450 );
and \U$25990 ( \26334 , \25596 , \21448 );
nor \U$25991 ( \26335 , \26333 , \26334 );
xnor \U$25992 ( \26336 , \26335 , \21457 );
and \U$25993 ( \26337 , \26078 , \21469 );
and \U$25994 ( \26338 , \26073 , \21467 );
nor \U$25995 ( \26339 , \26337 , \26338 );
xnor \U$25996 ( \26340 , \26339 , \21476 );
and \U$25997 ( \26341 , \26336 , \26340 );
buf \U$25998 ( \26342 , RIbb32a90_173);
and \U$25999 ( \26343 , \26342 , \21464 );
and \U$26000 ( \26344 , \26340 , \26343 );
and \U$26001 ( \26345 , \26336 , \26343 );
or \U$26002 ( \26346 , \26341 , \26344 , \26345 );
and \U$26003 ( \26347 , \24714 , \21401 );
and \U$26004 ( \26348 , \24506 , \21399 );
nor \U$26005 ( \26349 , \26347 , \26348 );
xnor \U$26006 ( \26350 , \26349 , \21408 );
and \U$26007 ( \26351 , \24841 , \21419 );
and \U$26008 ( \26352 , \24836 , \21417 );
nor \U$26009 ( \26353 , \26351 , \26352 );
xnor \U$26010 ( \26354 , \26353 , \21426 );
and \U$26011 ( \26355 , \26350 , \26354 );
and \U$26012 ( \26356 , \25294 , \21434 );
and \U$26013 ( \26357 , \25097 , \21432 );
nor \U$26014 ( \26358 , \26356 , \26357 );
xnor \U$26015 ( \26359 , \26358 , \21441 );
and \U$26016 ( \26360 , \26354 , \26359 );
and \U$26017 ( \26361 , \26350 , \26359 );
or \U$26018 ( \26362 , \26355 , \26360 , \26361 );
and \U$26019 ( \26363 , \26346 , \26362 );
xnor \U$26020 ( \26364 , \26077 , \26079 );
and \U$26021 ( \26365 , \26362 , \26364 );
and \U$26022 ( \26366 , \26346 , \26364 );
or \U$26023 ( \26367 , \26363 , \26365 , \26366 );
and \U$26024 ( \26368 , \26331 , \26367 );
and \U$26025 ( \26369 , \26279 , \26367 );
or \U$26026 ( \26370 , \26332 , \26368 , \26369 );
xor \U$26027 ( \26371 , \26060 , \26064 );
xor \U$26028 ( \26372 , \26371 , \26069 );
xor \U$26029 ( \26373 , \26109 , \26113 );
xor \U$26030 ( \26374 , \26373 , \26118 );
and \U$26031 ( \26375 , \26372 , \26374 );
xor \U$26032 ( \26376 , \26126 , \26130 );
xor \U$26033 ( \26377 , \26376 , \26135 );
and \U$26034 ( \26378 , \26374 , \26377 );
and \U$26035 ( \26379 , \26372 , \26377 );
or \U$26036 ( \26380 , \26375 , \26378 , \26379 );
xor \U$26037 ( \26381 , \26093 , \26097 );
xor \U$26038 ( \26382 , \26381 , \26102 );
xor \U$26039 ( \26383 , \26024 , \26028 );
xor \U$26040 ( \26384 , \26383 , \26033 );
and \U$26041 ( \26385 , \26382 , \26384 );
xor \U$26042 ( \26386 , \26041 , \26045 );
xor \U$26043 ( \26387 , \26386 , \26050 );
and \U$26044 ( \26388 , \26384 , \26387 );
and \U$26045 ( \26389 , \26382 , \26387 );
or \U$26046 ( \26390 , \26385 , \26388 , \26389 );
and \U$26047 ( \26391 , \26380 , \26390 );
xor \U$26048 ( \26392 , \25835 , \25839 );
xor \U$26049 ( \26393 , \26392 , \25844 );
and \U$26050 ( \26394 , \26390 , \26393 );
and \U$26051 ( \26395 , \26380 , \26393 );
or \U$26052 ( \26396 , \26391 , \26394 , \26395 );
and \U$26053 ( \26397 , \26370 , \26396 );
xor \U$26054 ( \26398 , \25818 , \25822 );
xor \U$26055 ( \26399 , \26398 , \25827 );
xor \U$26056 ( \26400 , \26145 , \26147 );
xor \U$26057 ( \26401 , \26400 , \26150 );
and \U$26058 ( \26402 , \26399 , \26401 );
xor \U$26059 ( \26403 , \26155 , \26157 );
xor \U$26060 ( \26404 , \26403 , \26160 );
and \U$26061 ( \26405 , \26401 , \26404 );
and \U$26062 ( \26406 , \26399 , \26404 );
or \U$26063 ( \26407 , \26402 , \26405 , \26406 );
and \U$26064 ( \26408 , \26396 , \26407 );
and \U$26065 ( \26409 , \26370 , \26407 );
or \U$26066 ( \26410 , \26397 , \26408 , \26409 );
xor \U$26067 ( \26411 , \26020 , \26036 );
xor \U$26068 ( \26412 , \26411 , \26053 );
xor \U$26069 ( \26413 , \26072 , \26080 );
xor \U$26070 ( \26414 , \26413 , \26085 );
and \U$26071 ( \26415 , \26412 , \26414 );
xor \U$26072 ( \26416 , \26105 , \26121 );
xor \U$26073 ( \26417 , \26416 , \26138 );
and \U$26074 ( \26418 , \26414 , \26417 );
and \U$26075 ( \26419 , \26412 , \26417 );
or \U$26076 ( \26420 , \26415 , \26418 , \26419 );
xor \U$26077 ( \26421 , \25812 , \25830 );
xor \U$26078 ( \26422 , \26421 , \25847 );
and \U$26079 ( \26423 , \26420 , \26422 );
xor \U$26080 ( \26424 , \26172 , \26174 );
xor \U$26081 ( \26425 , \26424 , \26177 );
and \U$26082 ( \26426 , \26422 , \26425 );
and \U$26083 ( \26427 , \26420 , \26425 );
or \U$26084 ( \26428 , \26423 , \26426 , \26427 );
and \U$26085 ( \26429 , \26410 , \26428 );
xor \U$26086 ( \26430 , \25939 , \25949 );
xor \U$26087 ( \26431 , \26430 , \25952 );
and \U$26088 ( \26432 , \26428 , \26431 );
and \U$26089 ( \26433 , \26410 , \26431 );
or \U$26090 ( \26434 , \26429 , \26432 , \26433 );
xor \U$26091 ( \26435 , \25850 , \25902 );
xor \U$26092 ( \26436 , \26435 , \25926 );
xor \U$26093 ( \26437 , \26144 , \26169 );
xor \U$26094 ( \26438 , \26437 , \26180 );
and \U$26095 ( \26439 , \26436 , \26438 );
xor \U$26096 ( \26440 , \26185 , \26187 );
xor \U$26097 ( \26441 , \26440 , \26190 );
and \U$26098 ( \26442 , \26438 , \26441 );
and \U$26099 ( \26443 , \26436 , \26441 );
or \U$26100 ( \26444 , \26439 , \26442 , \26443 );
and \U$26101 ( \26445 , \26434 , \26444 );
xor \U$26102 ( \26446 , \25971 , \25973 );
xor \U$26103 ( \26447 , \26446 , \25976 );
and \U$26104 ( \26448 , \26444 , \26447 );
and \U$26105 ( \26449 , \26434 , \26447 );
or \U$26106 ( \26450 , \26445 , \26448 , \26449 );
xor \U$26107 ( \26451 , \25929 , \25955 );
xor \U$26108 ( \26452 , \26451 , \25966 );
xor \U$26109 ( \26453 , \26183 , \26193 );
xor \U$26110 ( \26454 , \26453 , \26196 );
and \U$26111 ( \26455 , \26452 , \26454 );
and \U$26112 ( \26456 , \26450 , \26455 );
xor \U$26113 ( \26457 , \26199 , \26201 );
xor \U$26114 ( \26458 , \26457 , \26204 );
and \U$26115 ( \26459 , \26455 , \26458 );
and \U$26116 ( \26460 , \26450 , \26458 );
or \U$26117 ( \26461 , \26456 , \26459 , \26460 );
xor \U$26118 ( \26462 , \26207 , \26209 );
xor \U$26119 ( \26463 , \26462 , \26212 );
and \U$26120 ( \26464 , \26461 , \26463 );
and \U$26121 ( \26465 , \26225 , \26464 );
xor \U$26122 ( \26466 , \26225 , \26464 );
xor \U$26123 ( \26467 , \26461 , \26463 );
xor \U$26124 ( \26468 , \25814 , \26226 );
xor \U$26125 ( \26469 , \26226 , \26227 );
not \U$26126 ( \26470 , \26469 );
and \U$26127 ( \26471 , \26468 , \26470 );
and \U$26128 ( \26472 , \21387 , \26471 );
not \U$26129 ( \26473 , \26472 );
xnor \U$26130 ( \26474 , \26473 , \26230 );
and \U$26131 ( \26475 , \21403 , \26005 );
and \U$26132 ( \26476 , \21379 , \26003 );
nor \U$26133 ( \26477 , \26475 , \26476 );
xnor \U$26134 ( \26478 , \26477 , \25817 );
and \U$26135 ( \26479 , \26474 , \26478 );
and \U$26136 ( \26480 , \21421 , \25631 );
and \U$26137 ( \26481 , \21395 , \25629 );
nor \U$26138 ( \26482 , \26480 , \26481 );
xnor \U$26139 ( \26483 , \26482 , \25399 );
and \U$26140 ( \26484 , \26478 , \26483 );
and \U$26141 ( \26485 , \26474 , \26483 );
or \U$26142 ( \26486 , \26479 , \26484 , \26485 );
and \U$26143 ( \26487 , \21436 , \25180 );
and \U$26144 ( \26488 , \21413 , \25178 );
nor \U$26145 ( \26489 , \26487 , \26488 );
xnor \U$26146 ( \26490 , \26489 , \25037 );
and \U$26147 ( \26491 , \21452 , \24857 );
and \U$26148 ( \26492 , \21428 , \24855 );
nor \U$26149 ( \26493 , \26491 , \26492 );
xnor \U$26150 ( \26494 , \26493 , \24611 );
and \U$26151 ( \26495 , \26490 , \26494 );
and \U$26152 ( \26496 , \21471 , \24462 );
and \U$26153 ( \26497 , \21444 , \24460 );
nor \U$26154 ( \26498 , \26496 , \26497 );
xnor \U$26155 ( \26499 , \26498 , \24275 );
and \U$26156 ( \26500 , \26494 , \26499 );
and \U$26157 ( \26501 , \26490 , \26499 );
or \U$26158 ( \26502 , \26495 , \26500 , \26501 );
and \U$26159 ( \26503 , \26486 , \26502 );
and \U$26160 ( \26504 , \21478 , \24149 );
and \U$26161 ( \26505 , \21463 , \24147 );
nor \U$26162 ( \26506 , \26504 , \26505 );
xnor \U$26163 ( \26507 , \26506 , \23944 );
and \U$26164 ( \26508 , \21750 , \23743 );
and \U$26165 ( \26509 , \21689 , \23741 );
nor \U$26166 ( \26510 , \26508 , \26509 );
xnor \U$26167 ( \26511 , \26510 , \23594 );
and \U$26168 ( \26512 , \26507 , \26511 );
and \U$26169 ( \26513 , \22011 , \23421 );
and \U$26170 ( \26514 , \21813 , \23419 );
nor \U$26171 ( \26515 , \26513 , \26514 );
xnor \U$26172 ( \26516 , \26515 , \23279 );
and \U$26173 ( \26517 , \26511 , \26516 );
and \U$26174 ( \26518 , \26507 , \26516 );
or \U$26175 ( \26519 , \26512 , \26517 , \26518 );
and \U$26176 ( \26520 , \26502 , \26519 );
and \U$26177 ( \26521 , \26486 , \26519 );
or \U$26178 ( \26522 , \26503 , \26520 , \26521 );
and \U$26179 ( \26523 , \22204 , \23125 );
and \U$26180 ( \26524 , \22099 , \23123 );
nor \U$26181 ( \26525 , \26523 , \26524 );
xnor \U$26182 ( \26526 , \26525 , \22988 );
and \U$26183 ( \26527 , \22325 , \22919 );
and \U$26184 ( \26528 , \22209 , \22917 );
nor \U$26185 ( \26529 , \26527 , \26528 );
xnor \U$26186 ( \26530 , \26529 , \22767 );
and \U$26187 ( \26531 , \26526 , \26530 );
and \U$26188 ( \26532 , \22616 , \22651 );
and \U$26189 ( \26533 , \22440 , \22649 );
nor \U$26190 ( \26534 , \26532 , \26533 );
xnor \U$26191 ( \26535 , \26534 , \22495 );
and \U$26192 ( \26536 , \26530 , \26535 );
and \U$26193 ( \26537 , \26526 , \26535 );
or \U$26194 ( \26538 , \26531 , \26536 , \26537 );
and \U$26195 ( \26539 , \22867 , \22379 );
and \U$26196 ( \26540 , \22624 , \22377 );
nor \U$26197 ( \26541 , \26539 , \26540 );
xnor \U$26198 ( \26542 , \26541 , \22266 );
and \U$26199 ( \26543 , \23058 , \22185 );
and \U$26200 ( \26544 , \22872 , \22183 );
nor \U$26201 ( \26545 , \26543 , \26544 );
xnor \U$26202 ( \26546 , \26545 , \22049 );
and \U$26203 ( \26547 , \26542 , \26546 );
and \U$26204 ( \26548 , \23466 , \21985 );
and \U$26205 ( \26549 , \23202 , \21983 );
nor \U$26206 ( \26550 , \26548 , \26549 );
xnor \U$26207 ( \26551 , \26550 , \21907 );
and \U$26208 ( \26552 , \26546 , \26551 );
and \U$26209 ( \26553 , \26542 , \26551 );
or \U$26210 ( \26554 , \26547 , \26552 , \26553 );
and \U$26211 ( \26555 , \26538 , \26554 );
and \U$26212 ( \26556 , \23665 , \21821 );
and \U$26213 ( \26557 , \23491 , \21819 );
nor \U$26214 ( \26558 , \26556 , \26557 );
xnor \U$26215 ( \26559 , \26558 , \21727 );
and \U$26216 ( \26560 , \23970 , \21652 );
and \U$26217 ( \26561 , \23832 , \21650 );
nor \U$26218 ( \26562 , \26560 , \26561 );
xnor \U$26219 ( \26563 , \26562 , \21377 );
and \U$26220 ( \26564 , \26559 , \26563 );
and \U$26221 ( \26565 , \24506 , \21385 );
and \U$26222 ( \26566 , \24089 , \21383 );
nor \U$26223 ( \26567 , \26565 , \26566 );
xnor \U$26224 ( \26568 , \26567 , \21392 );
and \U$26225 ( \26569 , \26563 , \26568 );
and \U$26226 ( \26570 , \26559 , \26568 );
or \U$26227 ( \26571 , \26564 , \26569 , \26570 );
and \U$26228 ( \26572 , \26554 , \26571 );
and \U$26229 ( \26573 , \26538 , \26571 );
or \U$26230 ( \26574 , \26555 , \26572 , \26573 );
and \U$26231 ( \26575 , \26522 , \26574 );
and \U$26232 ( \26576 , \24836 , \21401 );
and \U$26233 ( \26577 , \24714 , \21399 );
nor \U$26234 ( \26578 , \26576 , \26577 );
xnor \U$26235 ( \26579 , \26578 , \21408 );
and \U$26236 ( \26580 , \25097 , \21419 );
and \U$26237 ( \26581 , \24841 , \21417 );
nor \U$26238 ( \26582 , \26580 , \26581 );
xnor \U$26239 ( \26583 , \26582 , \21426 );
and \U$26240 ( \26584 , \26579 , \26583 );
and \U$26241 ( \26585 , \25596 , \21434 );
and \U$26242 ( \26586 , \25294 , \21432 );
nor \U$26243 ( \26587 , \26585 , \26586 );
xnor \U$26244 ( \26588 , \26587 , \21441 );
and \U$26245 ( \26589 , \26583 , \26588 );
and \U$26246 ( \26590 , \26579 , \26588 );
or \U$26247 ( \26591 , \26584 , \26589 , \26590 );
and \U$26248 ( \26592 , \26073 , \21450 );
and \U$26249 ( \26593 , \25604 , \21448 );
nor \U$26250 ( \26594 , \26592 , \26593 );
xnor \U$26251 ( \26595 , \26594 , \21457 );
and \U$26252 ( \26596 , \26342 , \21469 );
and \U$26253 ( \26597 , \26078 , \21467 );
nor \U$26254 ( \26598 , \26596 , \26597 );
xnor \U$26255 ( \26599 , \26598 , \21476 );
and \U$26256 ( \26600 , \26595 , \26599 );
buf \U$26257 ( \26601 , RIbb32b08_174);
and \U$26258 ( \26602 , \26601 , \21464 );
and \U$26259 ( \26603 , \26599 , \26602 );
and \U$26260 ( \26604 , \26595 , \26602 );
or \U$26261 ( \26605 , \26600 , \26603 , \26604 );
and \U$26262 ( \26606 , \26591 , \26605 );
xor \U$26263 ( \26607 , \26336 , \26340 );
xor \U$26264 ( \26608 , \26607 , \26343 );
and \U$26265 ( \26609 , \26605 , \26608 );
and \U$26266 ( \26610 , \26591 , \26608 );
or \U$26267 ( \26611 , \26606 , \26609 , \26610 );
and \U$26268 ( \26612 , \26574 , \26611 );
and \U$26269 ( \26613 , \26522 , \26611 );
or \U$26270 ( \26614 , \26575 , \26612 , \26613 );
xor \U$26271 ( \26615 , \26283 , \26287 );
xor \U$26272 ( \26616 , \26615 , \26292 );
xor \U$26273 ( \26617 , \26247 , \26251 );
xor \U$26274 ( \26618 , \26617 , \26256 );
and \U$26275 ( \26619 , \26616 , \26618 );
xor \U$26276 ( \26620 , \26264 , \26268 );
xor \U$26277 ( \26621 , \26620 , \26273 );
and \U$26278 ( \26622 , \26618 , \26621 );
and \U$26279 ( \26623 , \26616 , \26621 );
or \U$26280 ( \26624 , \26619 , \26622 , \26623 );
xor \U$26281 ( \26625 , \26299 , \26303 );
xor \U$26282 ( \26626 , \26625 , \26308 );
xor \U$26283 ( \26627 , \26316 , \26320 );
xor \U$26284 ( \26628 , \26627 , \26325 );
and \U$26285 ( \26629 , \26626 , \26628 );
xor \U$26286 ( \26630 , \26350 , \26354 );
xor \U$26287 ( \26631 , \26630 , \26359 );
and \U$26288 ( \26632 , \26628 , \26631 );
and \U$26289 ( \26633 , \26626 , \26631 );
or \U$26290 ( \26634 , \26629 , \26632 , \26633 );
and \U$26291 ( \26635 , \26624 , \26634 );
xor \U$26292 ( \26636 , \26008 , \26012 );
xor \U$26293 ( \26637 , \26636 , \26017 );
and \U$26294 ( \26638 , \26634 , \26637 );
and \U$26295 ( \26639 , \26624 , \26637 );
or \U$26296 ( \26640 , \26635 , \26638 , \26639 );
and \U$26297 ( \26641 , \26614 , \26640 );
xor \U$26298 ( \26642 , \26372 , \26374 );
xor \U$26299 ( \26643 , \26642 , \26377 );
xor \U$26300 ( \26644 , \26382 , \26384 );
xor \U$26301 ( \26645 , \26644 , \26387 );
and \U$26302 ( \26646 , \26643 , \26645 );
xor \U$26303 ( \26647 , \26346 , \26362 );
xor \U$26304 ( \26648 , \26647 , \26364 );
and \U$26305 ( \26649 , \26645 , \26648 );
and \U$26306 ( \26650 , \26643 , \26648 );
or \U$26307 ( \26651 , \26646 , \26649 , \26650 );
and \U$26308 ( \26652 , \26640 , \26651 );
and \U$26309 ( \26653 , \26614 , \26651 );
or \U$26310 ( \26654 , \26641 , \26652 , \26653 );
xor \U$26311 ( \26655 , \26380 , \26390 );
xor \U$26312 ( \26656 , \26655 , \26393 );
xor \U$26313 ( \26657 , \26412 , \26414 );
xor \U$26314 ( \26658 , \26657 , \26417 );
and \U$26315 ( \26659 , \26656 , \26658 );
xor \U$26316 ( \26660 , \26399 , \26401 );
xor \U$26317 ( \26661 , \26660 , \26404 );
and \U$26318 ( \26662 , \26658 , \26661 );
and \U$26319 ( \26663 , \26656 , \26661 );
or \U$26320 ( \26664 , \26659 , \26662 , \26663 );
and \U$26321 ( \26665 , \26654 , \26664 );
xor \U$26322 ( \26666 , \26153 , \26163 );
xor \U$26323 ( \26667 , \26666 , \26166 );
and \U$26324 ( \26668 , \26664 , \26667 );
and \U$26325 ( \26669 , \26654 , \26667 );
or \U$26326 ( \26670 , \26665 , \26668 , \26669 );
xor \U$26327 ( \26671 , \26056 , \26088 );
xor \U$26328 ( \26672 , \26671 , \26141 );
xor \U$26329 ( \26673 , \26370 , \26396 );
xor \U$26330 ( \26674 , \26673 , \26407 );
and \U$26331 ( \26675 , \26672 , \26674 );
xor \U$26332 ( \26676 , \26420 , \26422 );
xor \U$26333 ( \26677 , \26676 , \26425 );
and \U$26334 ( \26678 , \26674 , \26677 );
and \U$26335 ( \26679 , \26672 , \26677 );
or \U$26336 ( \26680 , \26675 , \26678 , \26679 );
and \U$26337 ( \26681 , \26670 , \26680 );
xor \U$26338 ( \26682 , \26436 , \26438 );
xor \U$26339 ( \26683 , \26682 , \26441 );
and \U$26340 ( \26684 , \26680 , \26683 );
and \U$26341 ( \26685 , \26670 , \26683 );
or \U$26342 ( \26686 , \26681 , \26684 , \26685 );
xor \U$26343 ( \26687 , \26434 , \26444 );
xor \U$26344 ( \26688 , \26687 , \26447 );
and \U$26345 ( \26689 , \26686 , \26688 );
xor \U$26346 ( \26690 , \26452 , \26454 );
and \U$26347 ( \26691 , \26688 , \26690 );
and \U$26348 ( \26692 , \26686 , \26690 );
or \U$26349 ( \26693 , \26689 , \26691 , \26692 );
xor \U$26350 ( \26694 , \26450 , \26455 );
xor \U$26351 ( \26695 , \26694 , \26458 );
and \U$26352 ( \26696 , \26693 , \26695 );
and \U$26353 ( \26697 , \26467 , \26696 );
xor \U$26354 ( \26698 , \26467 , \26696 );
xor \U$26355 ( \26699 , \26693 , \26695 );
and \U$26356 ( \26700 , \21413 , \25631 );
and \U$26357 ( \26701 , \21421 , \25629 );
nor \U$26358 ( \26702 , \26700 , \26701 );
xnor \U$26359 ( \26703 , \26702 , \25399 );
and \U$26360 ( \26704 , \21428 , \25180 );
and \U$26361 ( \26705 , \21436 , \25178 );
nor \U$26362 ( \26706 , \26704 , \26705 );
xnor \U$26363 ( \26707 , \26706 , \25037 );
and \U$26364 ( \26708 , \26703 , \26707 );
and \U$26365 ( \26709 , \21444 , \24857 );
and \U$26366 ( \26710 , \21452 , \24855 );
nor \U$26367 ( \26711 , \26709 , \26710 );
xnor \U$26368 ( \26712 , \26711 , \24611 );
and \U$26369 ( \26713 , \26707 , \26712 );
and \U$26370 ( \26714 , \26703 , \26712 );
or \U$26371 ( \26715 , \26708 , \26713 , \26714 );
buf \U$26372 ( \26716 , RIbb2e008_48);
buf \U$26373 ( \26717 , RIbb2df90_49);
and \U$26374 ( \26718 , \26716 , \26717 );
not \U$26375 ( \26719 , \26718 );
and \U$26376 ( \26720 , \26227 , \26719 );
not \U$26377 ( \26721 , \26720 );
and \U$26378 ( \26722 , \21379 , \26471 );
and \U$26379 ( \26723 , \21387 , \26469 );
nor \U$26380 ( \26724 , \26722 , \26723 );
xnor \U$26381 ( \26725 , \26724 , \26230 );
and \U$26382 ( \26726 , \26721 , \26725 );
and \U$26383 ( \26727 , \21395 , \26005 );
and \U$26384 ( \26728 , \21403 , \26003 );
nor \U$26385 ( \26729 , \26727 , \26728 );
xnor \U$26386 ( \26730 , \26729 , \25817 );
and \U$26387 ( \26731 , \26725 , \26730 );
and \U$26388 ( \26732 , \26721 , \26730 );
or \U$26389 ( \26733 , \26726 , \26731 , \26732 );
and \U$26390 ( \26734 , \26715 , \26733 );
and \U$26391 ( \26735 , \21463 , \24462 );
and \U$26392 ( \26736 , \21471 , \24460 );
nor \U$26393 ( \26737 , \26735 , \26736 );
xnor \U$26394 ( \26738 , \26737 , \24275 );
and \U$26395 ( \26739 , \21689 , \24149 );
and \U$26396 ( \26740 , \21478 , \24147 );
nor \U$26397 ( \26741 , \26739 , \26740 );
xnor \U$26398 ( \26742 , \26741 , \23944 );
and \U$26399 ( \26743 , \26738 , \26742 );
and \U$26400 ( \26744 , \21813 , \23743 );
and \U$26401 ( \26745 , \21750 , \23741 );
nor \U$26402 ( \26746 , \26744 , \26745 );
xnor \U$26403 ( \26747 , \26746 , \23594 );
and \U$26404 ( \26748 , \26742 , \26747 );
and \U$26405 ( \26749 , \26738 , \26747 );
or \U$26406 ( \26750 , \26743 , \26748 , \26749 );
and \U$26407 ( \26751 , \26733 , \26750 );
and \U$26408 ( \26752 , \26715 , \26750 );
or \U$26409 ( \26753 , \26734 , \26751 , \26752 );
and \U$26410 ( \26754 , \23491 , \21985 );
and \U$26411 ( \26755 , \23466 , \21983 );
nor \U$26412 ( \26756 , \26754 , \26755 );
xnor \U$26413 ( \26757 , \26756 , \21907 );
and \U$26414 ( \26758 , \23832 , \21821 );
and \U$26415 ( \26759 , \23665 , \21819 );
nor \U$26416 ( \26760 , \26758 , \26759 );
xnor \U$26417 ( \26761 , \26760 , \21727 );
and \U$26418 ( \26762 , \26757 , \26761 );
and \U$26419 ( \26763 , \24089 , \21652 );
and \U$26420 ( \26764 , \23970 , \21650 );
nor \U$26421 ( \26765 , \26763 , \26764 );
xnor \U$26422 ( \26766 , \26765 , \21377 );
and \U$26423 ( \26767 , \26761 , \26766 );
and \U$26424 ( \26768 , \26757 , \26766 );
or \U$26425 ( \26769 , \26762 , \26767 , \26768 );
and \U$26426 ( \26770 , \22624 , \22651 );
and \U$26427 ( \26771 , \22616 , \22649 );
nor \U$26428 ( \26772 , \26770 , \26771 );
xnor \U$26429 ( \26773 , \26772 , \22495 );
and \U$26430 ( \26774 , \22872 , \22379 );
and \U$26431 ( \26775 , \22867 , \22377 );
nor \U$26432 ( \26776 , \26774 , \26775 );
xnor \U$26433 ( \26777 , \26776 , \22266 );
and \U$26434 ( \26778 , \26773 , \26777 );
and \U$26435 ( \26779 , \23202 , \22185 );
and \U$26436 ( \26780 , \23058 , \22183 );
nor \U$26437 ( \26781 , \26779 , \26780 );
xnor \U$26438 ( \26782 , \26781 , \22049 );
and \U$26439 ( \26783 , \26777 , \26782 );
and \U$26440 ( \26784 , \26773 , \26782 );
or \U$26441 ( \26785 , \26778 , \26783 , \26784 );
and \U$26442 ( \26786 , \26769 , \26785 );
and \U$26443 ( \26787 , \22099 , \23421 );
and \U$26444 ( \26788 , \22011 , \23419 );
nor \U$26445 ( \26789 , \26787 , \26788 );
xnor \U$26446 ( \26790 , \26789 , \23279 );
and \U$26447 ( \26791 , \22209 , \23125 );
and \U$26448 ( \26792 , \22204 , \23123 );
nor \U$26449 ( \26793 , \26791 , \26792 );
xnor \U$26450 ( \26794 , \26793 , \22988 );
and \U$26451 ( \26795 , \26790 , \26794 );
and \U$26452 ( \26796 , \22440 , \22919 );
and \U$26453 ( \26797 , \22325 , \22917 );
nor \U$26454 ( \26798 , \26796 , \26797 );
xnor \U$26455 ( \26799 , \26798 , \22767 );
and \U$26456 ( \26800 , \26794 , \26799 );
and \U$26457 ( \26801 , \26790 , \26799 );
or \U$26458 ( \26802 , \26795 , \26800 , \26801 );
and \U$26459 ( \26803 , \26785 , \26802 );
and \U$26460 ( \26804 , \26769 , \26802 );
or \U$26461 ( \26805 , \26786 , \26803 , \26804 );
and \U$26462 ( \26806 , \26753 , \26805 );
and \U$26463 ( \26807 , \24714 , \21385 );
and \U$26464 ( \26808 , \24506 , \21383 );
nor \U$26465 ( \26809 , \26807 , \26808 );
xnor \U$26466 ( \26810 , \26809 , \21392 );
and \U$26467 ( \26811 , \24841 , \21401 );
and \U$26468 ( \26812 , \24836 , \21399 );
nor \U$26469 ( \26813 , \26811 , \26812 );
xnor \U$26470 ( \26814 , \26813 , \21408 );
and \U$26471 ( \26815 , \26810 , \26814 );
and \U$26472 ( \26816 , \25294 , \21419 );
and \U$26473 ( \26817 , \25097 , \21417 );
nor \U$26474 ( \26818 , \26816 , \26817 );
xnor \U$26475 ( \26819 , \26818 , \21426 );
and \U$26476 ( \26820 , \26814 , \26819 );
and \U$26477 ( \26821 , \26810 , \26819 );
or \U$26478 ( \26822 , \26815 , \26820 , \26821 );
and \U$26479 ( \26823 , \25604 , \21434 );
and \U$26480 ( \26824 , \25596 , \21432 );
nor \U$26481 ( \26825 , \26823 , \26824 );
xnor \U$26482 ( \26826 , \26825 , \21441 );
and \U$26483 ( \26827 , \26078 , \21450 );
and \U$26484 ( \26828 , \26073 , \21448 );
nor \U$26485 ( \26829 , \26827 , \26828 );
xnor \U$26486 ( \26830 , \26829 , \21457 );
and \U$26487 ( \26831 , \26826 , \26830 );
and \U$26488 ( \26832 , \26601 , \21469 );
and \U$26489 ( \26833 , \26342 , \21467 );
nor \U$26490 ( \26834 , \26832 , \26833 );
xnor \U$26491 ( \26835 , \26834 , \21476 );
and \U$26492 ( \26836 , \26830 , \26835 );
and \U$26493 ( \26837 , \26826 , \26835 );
or \U$26494 ( \26838 , \26831 , \26836 , \26837 );
or \U$26495 ( \26839 , \26822 , \26838 );
and \U$26496 ( \26840 , \26805 , \26839 );
and \U$26497 ( \26841 , \26753 , \26839 );
or \U$26498 ( \26842 , \26806 , \26840 , \26841 );
xor \U$26499 ( \26843 , \26526 , \26530 );
xor \U$26500 ( \26844 , \26843 , \26535 );
xor \U$26501 ( \26845 , \26542 , \26546 );
xor \U$26502 ( \26846 , \26845 , \26551 );
and \U$26503 ( \26847 , \26844 , \26846 );
xor \U$26504 ( \26848 , \26507 , \26511 );
xor \U$26505 ( \26849 , \26848 , \26516 );
and \U$26506 ( \26850 , \26846 , \26849 );
and \U$26507 ( \26851 , \26844 , \26849 );
or \U$26508 ( \26852 , \26847 , \26850 , \26851 );
xor \U$26509 ( \26853 , \26559 , \26563 );
xor \U$26510 ( \26854 , \26853 , \26568 );
xor \U$26511 ( \26855 , \26579 , \26583 );
xor \U$26512 ( \26856 , \26855 , \26588 );
and \U$26513 ( \26857 , \26854 , \26856 );
xor \U$26514 ( \26858 , \26595 , \26599 );
xor \U$26515 ( \26859 , \26858 , \26602 );
and \U$26516 ( \26860 , \26856 , \26859 );
and \U$26517 ( \26861 , \26854 , \26859 );
or \U$26518 ( \26862 , \26857 , \26860 , \26861 );
and \U$26519 ( \26863 , \26852 , \26862 );
xor \U$26520 ( \26864 , \26474 , \26478 );
xor \U$26521 ( \26865 , \26864 , \26483 );
xor \U$26522 ( \26866 , \26490 , \26494 );
xor \U$26523 ( \26867 , \26866 , \26499 );
and \U$26524 ( \26868 , \26865 , \26867 );
and \U$26525 ( \26869 , \26862 , \26868 );
and \U$26526 ( \26870 , \26852 , \26868 );
or \U$26527 ( \26871 , \26863 , \26869 , \26870 );
and \U$26528 ( \26872 , \26842 , \26871 );
xor \U$26529 ( \26873 , \26231 , \26235 );
xor \U$26530 ( \26874 , \26873 , \26240 );
xor \U$26531 ( \26875 , \26616 , \26618 );
xor \U$26532 ( \26876 , \26875 , \26621 );
and \U$26533 ( \26877 , \26874 , \26876 );
xor \U$26534 ( \26878 , \26626 , \26628 );
xor \U$26535 ( \26879 , \26878 , \26631 );
and \U$26536 ( \26880 , \26876 , \26879 );
and \U$26537 ( \26881 , \26874 , \26879 );
or \U$26538 ( \26882 , \26877 , \26880 , \26881 );
and \U$26539 ( \26883 , \26871 , \26882 );
and \U$26540 ( \26884 , \26842 , \26882 );
or \U$26541 ( \26885 , \26872 , \26883 , \26884 );
xor \U$26542 ( \26886 , \26486 , \26502 );
xor \U$26543 ( \26887 , \26886 , \26519 );
xor \U$26544 ( \26888 , \26538 , \26554 );
xor \U$26545 ( \26889 , \26888 , \26571 );
and \U$26546 ( \26890 , \26887 , \26889 );
xor \U$26547 ( \26891 , \26591 , \26605 );
xor \U$26548 ( \26892 , \26891 , \26608 );
and \U$26549 ( \26893 , \26889 , \26892 );
and \U$26550 ( \26894 , \26887 , \26892 );
or \U$26551 ( \26895 , \26890 , \26893 , \26894 );
xor \U$26552 ( \26896 , \26243 , \26259 );
xor \U$26553 ( \26897 , \26896 , \26276 );
and \U$26554 ( \26898 , \26895 , \26897 );
xor \U$26555 ( \26899 , \26295 , \26311 );
xor \U$26556 ( \26900 , \26899 , \26328 );
and \U$26557 ( \26901 , \26897 , \26900 );
and \U$26558 ( \26902 , \26895 , \26900 );
or \U$26559 ( \26903 , \26898 , \26901 , \26902 );
and \U$26560 ( \26904 , \26885 , \26903 );
xor \U$26561 ( \26905 , \26522 , \26574 );
xor \U$26562 ( \26906 , \26905 , \26611 );
xor \U$26563 ( \26907 , \26624 , \26634 );
xor \U$26564 ( \26908 , \26907 , \26637 );
and \U$26565 ( \26909 , \26906 , \26908 );
xor \U$26566 ( \26910 , \26643 , \26645 );
xor \U$26567 ( \26911 , \26910 , \26648 );
and \U$26568 ( \26912 , \26908 , \26911 );
and \U$26569 ( \26913 , \26906 , \26911 );
or \U$26570 ( \26914 , \26909 , \26912 , \26913 );
and \U$26571 ( \26915 , \26903 , \26914 );
and \U$26572 ( \26916 , \26885 , \26914 );
or \U$26573 ( \26917 , \26904 , \26915 , \26916 );
xor \U$26574 ( \26918 , \26279 , \26331 );
xor \U$26575 ( \26919 , \26918 , \26367 );
xor \U$26576 ( \26920 , \26614 , \26640 );
xor \U$26577 ( \26921 , \26920 , \26651 );
and \U$26578 ( \26922 , \26919 , \26921 );
xor \U$26579 ( \26923 , \26656 , \26658 );
xor \U$26580 ( \26924 , \26923 , \26661 );
and \U$26581 ( \26925 , \26921 , \26924 );
and \U$26582 ( \26926 , \26919 , \26924 );
or \U$26583 ( \26927 , \26922 , \26925 , \26926 );
and \U$26584 ( \26928 , \26917 , \26927 );
xor \U$26585 ( \26929 , \26672 , \26674 );
xor \U$26586 ( \26930 , \26929 , \26677 );
and \U$26587 ( \26931 , \26927 , \26930 );
and \U$26588 ( \26932 , \26917 , \26930 );
or \U$26589 ( \26933 , \26928 , \26931 , \26932 );
xor \U$26590 ( \26934 , \26410 , \26428 );
xor \U$26591 ( \26935 , \26934 , \26431 );
and \U$26592 ( \26936 , \26933 , \26935 );
xor \U$26593 ( \26937 , \26670 , \26680 );
xor \U$26594 ( \26938 , \26937 , \26683 );
and \U$26595 ( \26939 , \26935 , \26938 );
and \U$26596 ( \26940 , \26933 , \26938 );
or \U$26597 ( \26941 , \26936 , \26939 , \26940 );
xor \U$26598 ( \26942 , \26686 , \26688 );
xor \U$26599 ( \26943 , \26942 , \26690 );
and \U$26600 ( \26944 , \26941 , \26943 );
and \U$26601 ( \26945 , \26699 , \26944 );
xor \U$26602 ( \26946 , \26699 , \26944 );
xor \U$26603 ( \26947 , \26941 , \26943 );
and \U$26604 ( \26948 , \24836 , \21385 );
and \U$26605 ( \26949 , \24714 , \21383 );
nor \U$26606 ( \26950 , \26948 , \26949 );
xnor \U$26607 ( \26951 , \26950 , \21392 );
and \U$26608 ( \26952 , \25097 , \21401 );
and \U$26609 ( \26953 , \24841 , \21399 );
nor \U$26610 ( \26954 , \26952 , \26953 );
xnor \U$26611 ( \26955 , \26954 , \21408 );
and \U$26612 ( \26956 , \26951 , \26955 );
and \U$26613 ( \26957 , \25596 , \21419 );
and \U$26614 ( \26958 , \25294 , \21417 );
nor \U$26615 ( \26959 , \26957 , \26958 );
xnor \U$26616 ( \26960 , \26959 , \21426 );
and \U$26617 ( \26961 , \26955 , \26960 );
and \U$26618 ( \26962 , \26951 , \26960 );
or \U$26619 ( \26963 , \26956 , \26961 , \26962 );
and \U$26620 ( \26964 , \26073 , \21434 );
and \U$26621 ( \26965 , \25604 , \21432 );
nor \U$26622 ( \26966 , \26964 , \26965 );
xnor \U$26623 ( \26967 , \26966 , \21441 );
and \U$26624 ( \26968 , \26342 , \21450 );
and \U$26625 ( \26969 , \26078 , \21448 );
nor \U$26626 ( \26970 , \26968 , \26969 );
xnor \U$26627 ( \26971 , \26970 , \21457 );
and \U$26628 ( \26972 , \26967 , \26971 );
buf \U$26629 ( \26973 , RIbb32b80_175);
and \U$26630 ( \26974 , \26973 , \21469 );
and \U$26631 ( \26975 , \26601 , \21467 );
nor \U$26632 ( \26976 , \26974 , \26975 );
xnor \U$26633 ( \26977 , \26976 , \21476 );
and \U$26634 ( \26978 , \26971 , \26977 );
and \U$26635 ( \26979 , \26967 , \26977 );
or \U$26636 ( \26980 , \26972 , \26978 , \26979 );
and \U$26637 ( \26981 , \26963 , \26980 );
buf \U$26638 ( \26982 , RIbb32bf8_176);
and \U$26639 ( \26983 , \26982 , \21464 );
buf \U$26640 ( \26984 , \26983 );
and \U$26641 ( \26985 , \26980 , \26984 );
and \U$26642 ( \26986 , \26963 , \26984 );
or \U$26643 ( \26987 , \26981 , \26985 , \26986 );
and \U$26644 ( \26988 , \22867 , \22651 );
and \U$26645 ( \26989 , \22624 , \22649 );
nor \U$26646 ( \26990 , \26988 , \26989 );
xnor \U$26647 ( \26991 , \26990 , \22495 );
and \U$26648 ( \26992 , \23058 , \22379 );
and \U$26649 ( \26993 , \22872 , \22377 );
nor \U$26650 ( \26994 , \26992 , \26993 );
xnor \U$26651 ( \26995 , \26994 , \22266 );
and \U$26652 ( \26996 , \26991 , \26995 );
and \U$26653 ( \26997 , \23466 , \22185 );
and \U$26654 ( \26998 , \23202 , \22183 );
nor \U$26655 ( \26999 , \26997 , \26998 );
xnor \U$26656 ( \27000 , \26999 , \22049 );
and \U$26657 ( \27001 , \26995 , \27000 );
and \U$26658 ( \27002 , \26991 , \27000 );
or \U$26659 ( \27003 , \26996 , \27001 , \27002 );
and \U$26660 ( \27004 , \22204 , \23421 );
and \U$26661 ( \27005 , \22099 , \23419 );
nor \U$26662 ( \27006 , \27004 , \27005 );
xnor \U$26663 ( \27007 , \27006 , \23279 );
and \U$26664 ( \27008 , \22325 , \23125 );
and \U$26665 ( \27009 , \22209 , \23123 );
nor \U$26666 ( \27010 , \27008 , \27009 );
xnor \U$26667 ( \27011 , \27010 , \22988 );
and \U$26668 ( \27012 , \27007 , \27011 );
and \U$26669 ( \27013 , \22616 , \22919 );
and \U$26670 ( \27014 , \22440 , \22917 );
nor \U$26671 ( \27015 , \27013 , \27014 );
xnor \U$26672 ( \27016 , \27015 , \22767 );
and \U$26673 ( \27017 , \27011 , \27016 );
and \U$26674 ( \27018 , \27007 , \27016 );
or \U$26675 ( \27019 , \27012 , \27017 , \27018 );
and \U$26676 ( \27020 , \27003 , \27019 );
and \U$26677 ( \27021 , \23665 , \21985 );
and \U$26678 ( \27022 , \23491 , \21983 );
nor \U$26679 ( \27023 , \27021 , \27022 );
xnor \U$26680 ( \27024 , \27023 , \21907 );
and \U$26681 ( \27025 , \23970 , \21821 );
and \U$26682 ( \27026 , \23832 , \21819 );
nor \U$26683 ( \27027 , \27025 , \27026 );
xnor \U$26684 ( \27028 , \27027 , \21727 );
and \U$26685 ( \27029 , \27024 , \27028 );
and \U$26686 ( \27030 , \24506 , \21652 );
and \U$26687 ( \27031 , \24089 , \21650 );
nor \U$26688 ( \27032 , \27030 , \27031 );
xnor \U$26689 ( \27033 , \27032 , \21377 );
and \U$26690 ( \27034 , \27028 , \27033 );
and \U$26691 ( \27035 , \27024 , \27033 );
or \U$26692 ( \27036 , \27029 , \27034 , \27035 );
and \U$26693 ( \27037 , \27019 , \27036 );
and \U$26694 ( \27038 , \27003 , \27036 );
or \U$26695 ( \27039 , \27020 , \27037 , \27038 );
and \U$26696 ( \27040 , \26987 , \27039 );
and \U$26697 ( \27041 , \21436 , \25631 );
and \U$26698 ( \27042 , \21413 , \25629 );
nor \U$26699 ( \27043 , \27041 , \27042 );
xnor \U$26700 ( \27044 , \27043 , \25399 );
and \U$26701 ( \27045 , \21452 , \25180 );
and \U$26702 ( \27046 , \21428 , \25178 );
nor \U$26703 ( \27047 , \27045 , \27046 );
xnor \U$26704 ( \27048 , \27047 , \25037 );
and \U$26705 ( \27049 , \27044 , \27048 );
and \U$26706 ( \27050 , \21471 , \24857 );
and \U$26707 ( \27051 , \21444 , \24855 );
nor \U$26708 ( \27052 , \27050 , \27051 );
xnor \U$26709 ( \27053 , \27052 , \24611 );
and \U$26710 ( \27054 , \27048 , \27053 );
and \U$26711 ( \27055 , \27044 , \27053 );
or \U$26712 ( \27056 , \27049 , \27054 , \27055 );
xor \U$26713 ( \27057 , \26227 , \26716 );
xor \U$26714 ( \27058 , \26716 , \26717 );
not \U$26715 ( \27059 , \27058 );
and \U$26716 ( \27060 , \27057 , \27059 );
and \U$26717 ( \27061 , \21387 , \27060 );
not \U$26718 ( \27062 , \27061 );
xnor \U$26719 ( \27063 , \27062 , \26720 );
and \U$26720 ( \27064 , \21403 , \26471 );
and \U$26721 ( \27065 , \21379 , \26469 );
nor \U$26722 ( \27066 , \27064 , \27065 );
xnor \U$26723 ( \27067 , \27066 , \26230 );
and \U$26724 ( \27068 , \27063 , \27067 );
and \U$26725 ( \27069 , \21421 , \26005 );
and \U$26726 ( \27070 , \21395 , \26003 );
nor \U$26727 ( \27071 , \27069 , \27070 );
xnor \U$26728 ( \27072 , \27071 , \25817 );
and \U$26729 ( \27073 , \27067 , \27072 );
and \U$26730 ( \27074 , \27063 , \27072 );
or \U$26731 ( \27075 , \27068 , \27073 , \27074 );
and \U$26732 ( \27076 , \27056 , \27075 );
and \U$26733 ( \27077 , \21478 , \24462 );
and \U$26734 ( \27078 , \21463 , \24460 );
nor \U$26735 ( \27079 , \27077 , \27078 );
xnor \U$26736 ( \27080 , \27079 , \24275 );
and \U$26737 ( \27081 , \21750 , \24149 );
and \U$26738 ( \27082 , \21689 , \24147 );
nor \U$26739 ( \27083 , \27081 , \27082 );
xnor \U$26740 ( \27084 , \27083 , \23944 );
and \U$26741 ( \27085 , \27080 , \27084 );
and \U$26742 ( \27086 , \22011 , \23743 );
and \U$26743 ( \27087 , \21813 , \23741 );
nor \U$26744 ( \27088 , \27086 , \27087 );
xnor \U$26745 ( \27089 , \27088 , \23594 );
and \U$26746 ( \27090 , \27084 , \27089 );
and \U$26747 ( \27091 , \27080 , \27089 );
or \U$26748 ( \27092 , \27085 , \27090 , \27091 );
and \U$26749 ( \27093 , \27075 , \27092 );
and \U$26750 ( \27094 , \27056 , \27092 );
or \U$26751 ( \27095 , \27076 , \27093 , \27094 );
and \U$26752 ( \27096 , \27039 , \27095 );
and \U$26753 ( \27097 , \26987 , \27095 );
or \U$26754 ( \27098 , \27040 , \27096 , \27097 );
xor \U$26755 ( \27099 , \26703 , \26707 );
xor \U$26756 ( \27100 , \27099 , \26712 );
xor \U$26757 ( \27101 , \26721 , \26725 );
xor \U$26758 ( \27102 , \27101 , \26730 );
and \U$26759 ( \27103 , \27100 , \27102 );
xor \U$26760 ( \27104 , \26738 , \26742 );
xor \U$26761 ( \27105 , \27104 , \26747 );
and \U$26762 ( \27106 , \27102 , \27105 );
and \U$26763 ( \27107 , \27100 , \27105 );
or \U$26764 ( \27108 , \27103 , \27106 , \27107 );
xor \U$26765 ( \27109 , \26757 , \26761 );
xor \U$26766 ( \27110 , \27109 , \26766 );
xor \U$26767 ( \27111 , \26773 , \26777 );
xor \U$26768 ( \27112 , \27111 , \26782 );
and \U$26769 ( \27113 , \27110 , \27112 );
xor \U$26770 ( \27114 , \26790 , \26794 );
xor \U$26771 ( \27115 , \27114 , \26799 );
and \U$26772 ( \27116 , \27112 , \27115 );
and \U$26773 ( \27117 , \27110 , \27115 );
or \U$26774 ( \27118 , \27113 , \27116 , \27117 );
and \U$26775 ( \27119 , \27108 , \27118 );
and \U$26776 ( \27120 , \26973 , \21464 );
xor \U$26777 ( \27121 , \26810 , \26814 );
xor \U$26778 ( \27122 , \27121 , \26819 );
and \U$26779 ( \27123 , \27120 , \27122 );
xor \U$26780 ( \27124 , \26826 , \26830 );
xor \U$26781 ( \27125 , \27124 , \26835 );
and \U$26782 ( \27126 , \27122 , \27125 );
and \U$26783 ( \27127 , \27120 , \27125 );
or \U$26784 ( \27128 , \27123 , \27126 , \27127 );
and \U$26785 ( \27129 , \27118 , \27128 );
and \U$26786 ( \27130 , \27108 , \27128 );
or \U$26787 ( \27131 , \27119 , \27129 , \27130 );
and \U$26788 ( \27132 , \27098 , \27131 );
xor \U$26789 ( \27133 , \26844 , \26846 );
xor \U$26790 ( \27134 , \27133 , \26849 );
xor \U$26791 ( \27135 , \26854 , \26856 );
xor \U$26792 ( \27136 , \27135 , \26859 );
and \U$26793 ( \27137 , \27134 , \27136 );
xor \U$26794 ( \27138 , \26865 , \26867 );
and \U$26795 ( \27139 , \27136 , \27138 );
and \U$26796 ( \27140 , \27134 , \27138 );
or \U$26797 ( \27141 , \27137 , \27139 , \27140 );
and \U$26798 ( \27142 , \27131 , \27141 );
and \U$26799 ( \27143 , \27098 , \27141 );
or \U$26800 ( \27144 , \27132 , \27142 , \27143 );
xor \U$26801 ( \27145 , \26715 , \26733 );
xor \U$26802 ( \27146 , \27145 , \26750 );
xor \U$26803 ( \27147 , \26769 , \26785 );
xor \U$26804 ( \27148 , \27147 , \26802 );
and \U$26805 ( \27149 , \27146 , \27148 );
xnor \U$26806 ( \27150 , \26822 , \26838 );
and \U$26807 ( \27151 , \27148 , \27150 );
and \U$26808 ( \27152 , \27146 , \27150 );
or \U$26809 ( \27153 , \27149 , \27151 , \27152 );
xor \U$26810 ( \27154 , \26874 , \26876 );
xor \U$26811 ( \27155 , \27154 , \26879 );
and \U$26812 ( \27156 , \27153 , \27155 );
xor \U$26813 ( \27157 , \26887 , \26889 );
xor \U$26814 ( \27158 , \27157 , \26892 );
and \U$26815 ( \27159 , \27155 , \27158 );
and \U$26816 ( \27160 , \27153 , \27158 );
or \U$26817 ( \27161 , \27156 , \27159 , \27160 );
and \U$26818 ( \27162 , \27144 , \27161 );
xor \U$26819 ( \27163 , \26753 , \26805 );
xor \U$26820 ( \27164 , \27163 , \26839 );
xor \U$26821 ( \27165 , \26852 , \26862 );
xor \U$26822 ( \27166 , \27165 , \26868 );
and \U$26823 ( \27167 , \27164 , \27166 );
and \U$26824 ( \27168 , \27161 , \27167 );
and \U$26825 ( \27169 , \27144 , \27167 );
or \U$26826 ( \27170 , \27162 , \27168 , \27169 );
xor \U$26827 ( \27171 , \26842 , \26871 );
xor \U$26828 ( \27172 , \27171 , \26882 );
xor \U$26829 ( \27173 , \26895 , \26897 );
xor \U$26830 ( \27174 , \27173 , \26900 );
and \U$26831 ( \27175 , \27172 , \27174 );
xor \U$26832 ( \27176 , \26906 , \26908 );
xor \U$26833 ( \27177 , \27176 , \26911 );
and \U$26834 ( \27178 , \27174 , \27177 );
and \U$26835 ( \27179 , \27172 , \27177 );
or \U$26836 ( \27180 , \27175 , \27178 , \27179 );
and \U$26837 ( \27181 , \27170 , \27180 );
xor \U$26838 ( \27182 , \26919 , \26921 );
xor \U$26839 ( \27183 , \27182 , \26924 );
and \U$26840 ( \27184 , \27180 , \27183 );
and \U$26841 ( \27185 , \27170 , \27183 );
or \U$26842 ( \27186 , \27181 , \27184 , \27185 );
xor \U$26843 ( \27187 , \26654 , \26664 );
xor \U$26844 ( \27188 , \27187 , \26667 );
and \U$26845 ( \27189 , \27186 , \27188 );
xor \U$26846 ( \27190 , \26917 , \26927 );
xor \U$26847 ( \27191 , \27190 , \26930 );
and \U$26848 ( \27192 , \27188 , \27191 );
and \U$26849 ( \27193 , \27186 , \27191 );
or \U$26850 ( \27194 , \27189 , \27192 , \27193 );
xor \U$26851 ( \27195 , \26933 , \26935 );
xor \U$26852 ( \27196 , \27195 , \26938 );
and \U$26853 ( \27197 , \27194 , \27196 );
and \U$26854 ( \27198 , \26947 , \27197 );
xor \U$26855 ( \27199 , \26947 , \27197 );
xor \U$26856 ( \27200 , \27194 , \27196 );
xor \U$26857 ( \27201 , \26991 , \26995 );
xor \U$26858 ( \27202 , \27201 , \27000 );
xor \U$26859 ( \27203 , \27007 , \27011 );
xor \U$26860 ( \27204 , \27203 , \27016 );
and \U$26861 ( \27205 , \27202 , \27204 );
xor \U$26862 ( \27206 , \27024 , \27028 );
xor \U$26863 ( \27207 , \27206 , \27033 );
and \U$26864 ( \27208 , \27204 , \27207 );
and \U$26865 ( \27209 , \27202 , \27207 );
or \U$26866 ( \27210 , \27205 , \27208 , \27209 );
xor \U$26867 ( \27211 , \27044 , \27048 );
xor \U$26868 ( \27212 , \27211 , \27053 );
xor \U$26869 ( \27213 , \27063 , \27067 );
xor \U$26870 ( \27214 , \27213 , \27072 );
and \U$26871 ( \27215 , \27212 , \27214 );
xor \U$26872 ( \27216 , \27080 , \27084 );
xor \U$26873 ( \27217 , \27216 , \27089 );
and \U$26874 ( \27218 , \27214 , \27217 );
and \U$26875 ( \27219 , \27212 , \27217 );
or \U$26876 ( \27220 , \27215 , \27218 , \27219 );
and \U$26877 ( \27221 , \27210 , \27220 );
xor \U$26878 ( \27222 , \26951 , \26955 );
xor \U$26879 ( \27223 , \27222 , \26960 );
xor \U$26880 ( \27224 , \26967 , \26971 );
xor \U$26881 ( \27225 , \27224 , \26977 );
and \U$26882 ( \27226 , \27223 , \27225 );
not \U$26883 ( \27227 , \26983 );
and \U$26884 ( \27228 , \27225 , \27227 );
and \U$26885 ( \27229 , \27223 , \27227 );
or \U$26886 ( \27230 , \27226 , \27228 , \27229 );
and \U$26887 ( \27231 , \27220 , \27230 );
and \U$26888 ( \27232 , \27210 , \27230 );
or \U$26889 ( \27233 , \27221 , \27231 , \27232 );
and \U$26890 ( \27234 , \21413 , \26005 );
and \U$26891 ( \27235 , \21421 , \26003 );
nor \U$26892 ( \27236 , \27234 , \27235 );
xnor \U$26893 ( \27237 , \27236 , \25817 );
and \U$26894 ( \27238 , \21428 , \25631 );
and \U$26895 ( \27239 , \21436 , \25629 );
nor \U$26896 ( \27240 , \27238 , \27239 );
xnor \U$26897 ( \27241 , \27240 , \25399 );
and \U$26898 ( \27242 , \27237 , \27241 );
and \U$26899 ( \27243 , \21444 , \25180 );
and \U$26900 ( \27244 , \21452 , \25178 );
nor \U$26901 ( \27245 , \27243 , \27244 );
xnor \U$26902 ( \27246 , \27245 , \25037 );
and \U$26903 ( \27247 , \27241 , \27246 );
and \U$26904 ( \27248 , \27237 , \27246 );
or \U$26905 ( \27249 , \27242 , \27247 , \27248 );
buf \U$26906 ( \27250 , RIbb2df18_50);
buf \U$26907 ( \27251 , RIbb2dea0_51);
and \U$26908 ( \27252 , \27250 , \27251 );
not \U$26909 ( \27253 , \27252 );
and \U$26910 ( \27254 , \26717 , \27253 );
not \U$26911 ( \27255 , \27254 );
and \U$26912 ( \27256 , \21379 , \27060 );
and \U$26913 ( \27257 , \21387 , \27058 );
nor \U$26914 ( \27258 , \27256 , \27257 );
xnor \U$26915 ( \27259 , \27258 , \26720 );
and \U$26916 ( \27260 , \27255 , \27259 );
and \U$26917 ( \27261 , \21395 , \26471 );
and \U$26918 ( \27262 , \21403 , \26469 );
nor \U$26919 ( \27263 , \27261 , \27262 );
xnor \U$26920 ( \27264 , \27263 , \26230 );
and \U$26921 ( \27265 , \27259 , \27264 );
and \U$26922 ( \27266 , \27255 , \27264 );
or \U$26923 ( \27267 , \27260 , \27265 , \27266 );
and \U$26924 ( \27268 , \27249 , \27267 );
and \U$26925 ( \27269 , \21463 , \24857 );
and \U$26926 ( \27270 , \21471 , \24855 );
nor \U$26927 ( \27271 , \27269 , \27270 );
xnor \U$26928 ( \27272 , \27271 , \24611 );
and \U$26929 ( \27273 , \21689 , \24462 );
and \U$26930 ( \27274 , \21478 , \24460 );
nor \U$26931 ( \27275 , \27273 , \27274 );
xnor \U$26932 ( \27276 , \27275 , \24275 );
and \U$26933 ( \27277 , \27272 , \27276 );
and \U$26934 ( \27278 , \21813 , \24149 );
and \U$26935 ( \27279 , \21750 , \24147 );
nor \U$26936 ( \27280 , \27278 , \27279 );
xnor \U$26937 ( \27281 , \27280 , \23944 );
and \U$26938 ( \27282 , \27276 , \27281 );
and \U$26939 ( \27283 , \27272 , \27281 );
or \U$26940 ( \27284 , \27277 , \27282 , \27283 );
and \U$26941 ( \27285 , \27267 , \27284 );
and \U$26942 ( \27286 , \27249 , \27284 );
or \U$26943 ( \27287 , \27268 , \27285 , \27286 );
and \U$26944 ( \27288 , \24714 , \21652 );
and \U$26945 ( \27289 , \24506 , \21650 );
nor \U$26946 ( \27290 , \27288 , \27289 );
xnor \U$26947 ( \27291 , \27290 , \21377 );
and \U$26948 ( \27292 , \24841 , \21385 );
and \U$26949 ( \27293 , \24836 , \21383 );
nor \U$26950 ( \27294 , \27292 , \27293 );
xnor \U$26951 ( \27295 , \27294 , \21392 );
and \U$26952 ( \27296 , \27291 , \27295 );
and \U$26953 ( \27297 , \25294 , \21401 );
and \U$26954 ( \27298 , \25097 , \21399 );
nor \U$26955 ( \27299 , \27297 , \27298 );
xnor \U$26956 ( \27300 , \27299 , \21408 );
and \U$26957 ( \27301 , \27295 , \27300 );
and \U$26958 ( \27302 , \27291 , \27300 );
or \U$26959 ( \27303 , \27296 , \27301 , \27302 );
and \U$26960 ( \27304 , \25604 , \21419 );
and \U$26961 ( \27305 , \25596 , \21417 );
nor \U$26962 ( \27306 , \27304 , \27305 );
xnor \U$26963 ( \27307 , \27306 , \21426 );
and \U$26964 ( \27308 , \26078 , \21434 );
and \U$26965 ( \27309 , \26073 , \21432 );
nor \U$26966 ( \27310 , \27308 , \27309 );
xnor \U$26967 ( \27311 , \27310 , \21441 );
and \U$26968 ( \27312 , \27307 , \27311 );
and \U$26969 ( \27313 , \26601 , \21450 );
and \U$26970 ( \27314 , \26342 , \21448 );
nor \U$26971 ( \27315 , \27313 , \27314 );
xnor \U$26972 ( \27316 , \27315 , \21457 );
and \U$26973 ( \27317 , \27311 , \27316 );
and \U$26974 ( \27318 , \27307 , \27316 );
or \U$26975 ( \27319 , \27312 , \27317 , \27318 );
and \U$26976 ( \27320 , \27303 , \27319 );
and \U$26977 ( \27321 , \26982 , \21469 );
and \U$26978 ( \27322 , \26973 , \21467 );
nor \U$26979 ( \27323 , \27321 , \27322 );
xnor \U$26980 ( \27324 , \27323 , \21476 );
buf \U$26981 ( \27325 , RIbb32c70_177);
and \U$26982 ( \27326 , \27325 , \21464 );
and \U$26983 ( \27327 , \27324 , \27326 );
and \U$26984 ( \27328 , \27319 , \27327 );
and \U$26985 ( \27329 , \27303 , \27327 );
or \U$26986 ( \27330 , \27320 , \27328 , \27329 );
and \U$26987 ( \27331 , \27287 , \27330 );
and \U$26988 ( \27332 , \22099 , \23743 );
and \U$26989 ( \27333 , \22011 , \23741 );
nor \U$26990 ( \27334 , \27332 , \27333 );
xnor \U$26991 ( \27335 , \27334 , \23594 );
and \U$26992 ( \27336 , \22209 , \23421 );
and \U$26993 ( \27337 , \22204 , \23419 );
nor \U$26994 ( \27338 , \27336 , \27337 );
xnor \U$26995 ( \27339 , \27338 , \23279 );
and \U$26996 ( \27340 , \27335 , \27339 );
and \U$26997 ( \27341 , \22440 , \23125 );
and \U$26998 ( \27342 , \22325 , \23123 );
nor \U$26999 ( \27343 , \27341 , \27342 );
xnor \U$27000 ( \27344 , \27343 , \22988 );
and \U$27001 ( \27345 , \27339 , \27344 );
and \U$27002 ( \27346 , \27335 , \27344 );
or \U$27003 ( \27347 , \27340 , \27345 , \27346 );
and \U$27004 ( \27348 , \22624 , \22919 );
and \U$27005 ( \27349 , \22616 , \22917 );
nor \U$27006 ( \27350 , \27348 , \27349 );
xnor \U$27007 ( \27351 , \27350 , \22767 );
and \U$27008 ( \27352 , \22872 , \22651 );
and \U$27009 ( \27353 , \22867 , \22649 );
nor \U$27010 ( \27354 , \27352 , \27353 );
xnor \U$27011 ( \27355 , \27354 , \22495 );
and \U$27012 ( \27356 , \27351 , \27355 );
and \U$27013 ( \27357 , \23202 , \22379 );
and \U$27014 ( \27358 , \23058 , \22377 );
nor \U$27015 ( \27359 , \27357 , \27358 );
xnor \U$27016 ( \27360 , \27359 , \22266 );
and \U$27017 ( \27361 , \27355 , \27360 );
and \U$27018 ( \27362 , \27351 , \27360 );
or \U$27019 ( \27363 , \27356 , \27361 , \27362 );
and \U$27020 ( \27364 , \27347 , \27363 );
and \U$27021 ( \27365 , \23491 , \22185 );
and \U$27022 ( \27366 , \23466 , \22183 );
nor \U$27023 ( \27367 , \27365 , \27366 );
xnor \U$27024 ( \27368 , \27367 , \22049 );
and \U$27025 ( \27369 , \23832 , \21985 );
and \U$27026 ( \27370 , \23665 , \21983 );
nor \U$27027 ( \27371 , \27369 , \27370 );
xnor \U$27028 ( \27372 , \27371 , \21907 );
and \U$27029 ( \27373 , \27368 , \27372 );
and \U$27030 ( \27374 , \24089 , \21821 );
and \U$27031 ( \27375 , \23970 , \21819 );
nor \U$27032 ( \27376 , \27374 , \27375 );
xnor \U$27033 ( \27377 , \27376 , \21727 );
and \U$27034 ( \27378 , \27372 , \27377 );
and \U$27035 ( \27379 , \27368 , \27377 );
or \U$27036 ( \27380 , \27373 , \27378 , \27379 );
and \U$27037 ( \27381 , \27363 , \27380 );
and \U$27038 ( \27382 , \27347 , \27380 );
or \U$27039 ( \27383 , \27364 , \27381 , \27382 );
and \U$27040 ( \27384 , \27330 , \27383 );
and \U$27041 ( \27385 , \27287 , \27383 );
or \U$27042 ( \27386 , \27331 , \27384 , \27385 );
and \U$27043 ( \27387 , \27233 , \27386 );
xor \U$27044 ( \27388 , \27100 , \27102 );
xor \U$27045 ( \27389 , \27388 , \27105 );
xor \U$27046 ( \27390 , \27110 , \27112 );
xor \U$27047 ( \27391 , \27390 , \27115 );
and \U$27048 ( \27392 , \27389 , \27391 );
xor \U$27049 ( \27393 , \27120 , \27122 );
xor \U$27050 ( \27394 , \27393 , \27125 );
and \U$27051 ( \27395 , \27391 , \27394 );
and \U$27052 ( \27396 , \27389 , \27394 );
or \U$27053 ( \27397 , \27392 , \27395 , \27396 );
and \U$27054 ( \27398 , \27386 , \27397 );
and \U$27055 ( \27399 , \27233 , \27397 );
or \U$27056 ( \27400 , \27387 , \27398 , \27399 );
xor \U$27057 ( \27401 , \26963 , \26980 );
xor \U$27058 ( \27402 , \27401 , \26984 );
xor \U$27059 ( \27403 , \27003 , \27019 );
xor \U$27060 ( \27404 , \27403 , \27036 );
and \U$27061 ( \27405 , \27402 , \27404 );
xor \U$27062 ( \27406 , \27056 , \27075 );
xor \U$27063 ( \27407 , \27406 , \27092 );
and \U$27064 ( \27408 , \27404 , \27407 );
and \U$27065 ( \27409 , \27402 , \27407 );
or \U$27066 ( \27410 , \27405 , \27408 , \27409 );
xor \U$27067 ( \27411 , \27146 , \27148 );
xor \U$27068 ( \27412 , \27411 , \27150 );
and \U$27069 ( \27413 , \27410 , \27412 );
xor \U$27070 ( \27414 , \27134 , \27136 );
xor \U$27071 ( \27415 , \27414 , \27138 );
and \U$27072 ( \27416 , \27412 , \27415 );
and \U$27073 ( \27417 , \27410 , \27415 );
or \U$27074 ( \27418 , \27413 , \27416 , \27417 );
and \U$27075 ( \27419 , \27400 , \27418 );
xor \U$27076 ( \27420 , \26987 , \27039 );
xor \U$27077 ( \27421 , \27420 , \27095 );
xor \U$27078 ( \27422 , \27108 , \27118 );
xor \U$27079 ( \27423 , \27422 , \27128 );
and \U$27080 ( \27424 , \27421 , \27423 );
and \U$27081 ( \27425 , \27418 , \27424 );
and \U$27082 ( \27426 , \27400 , \27424 );
or \U$27083 ( \27427 , \27419 , \27425 , \27426 );
xor \U$27084 ( \27428 , \27098 , \27131 );
xor \U$27085 ( \27429 , \27428 , \27141 );
xor \U$27086 ( \27430 , \27153 , \27155 );
xor \U$27087 ( \27431 , \27430 , \27158 );
and \U$27088 ( \27432 , \27429 , \27431 );
xor \U$27089 ( \27433 , \27164 , \27166 );
and \U$27090 ( \27434 , \27431 , \27433 );
and \U$27091 ( \27435 , \27429 , \27433 );
or \U$27092 ( \27436 , \27432 , \27434 , \27435 );
and \U$27093 ( \27437 , \27427 , \27436 );
xor \U$27094 ( \27438 , \27172 , \27174 );
xor \U$27095 ( \27439 , \27438 , \27177 );
and \U$27096 ( \27440 , \27436 , \27439 );
and \U$27097 ( \27441 , \27427 , \27439 );
or \U$27098 ( \27442 , \27437 , \27440 , \27441 );
xor \U$27099 ( \27443 , \26885 , \26903 );
xor \U$27100 ( \27444 , \27443 , \26914 );
and \U$27101 ( \27445 , \27442 , \27444 );
xor \U$27102 ( \27446 , \27170 , \27180 );
xor \U$27103 ( \27447 , \27446 , \27183 );
and \U$27104 ( \27448 , \27444 , \27447 );
and \U$27105 ( \27449 , \27442 , \27447 );
or \U$27106 ( \27450 , \27445 , \27448 , \27449 );
xor \U$27107 ( \27451 , \27186 , \27188 );
xor \U$27108 ( \27452 , \27451 , \27191 );
and \U$27109 ( \27453 , \27450 , \27452 );
and \U$27110 ( \27454 , \27200 , \27453 );
xor \U$27111 ( \27455 , \27200 , \27453 );
xor \U$27112 ( \27456 , \27450 , \27452 );
xor \U$27113 ( \27457 , \27335 , \27339 );
xor \U$27114 ( \27458 , \27457 , \27344 );
xor \U$27115 ( \27459 , \27351 , \27355 );
xor \U$27116 ( \27460 , \27459 , \27360 );
and \U$27117 ( \27461 , \27458 , \27460 );
xor \U$27118 ( \27462 , \27368 , \27372 );
xor \U$27119 ( \27463 , \27462 , \27377 );
and \U$27120 ( \27464 , \27460 , \27463 );
and \U$27121 ( \27465 , \27458 , \27463 );
or \U$27122 ( \27466 , \27461 , \27464 , \27465 );
xor \U$27123 ( \27467 , \27237 , \27241 );
xor \U$27124 ( \27468 , \27467 , \27246 );
xor \U$27125 ( \27469 , \27255 , \27259 );
xor \U$27126 ( \27470 , \27469 , \27264 );
and \U$27127 ( \27471 , \27468 , \27470 );
xor \U$27128 ( \27472 , \27272 , \27276 );
xor \U$27129 ( \27473 , \27472 , \27281 );
and \U$27130 ( \27474 , \27470 , \27473 );
and \U$27131 ( \27475 , \27468 , \27473 );
or \U$27132 ( \27476 , \27471 , \27474 , \27475 );
and \U$27133 ( \27477 , \27466 , \27476 );
xor \U$27134 ( \27478 , \27291 , \27295 );
xor \U$27135 ( \27479 , \27478 , \27300 );
xor \U$27136 ( \27480 , \27307 , \27311 );
xor \U$27137 ( \27481 , \27480 , \27316 );
and \U$27138 ( \27482 , \27479 , \27481 );
xor \U$27139 ( \27483 , \27324 , \27326 );
and \U$27140 ( \27484 , \27481 , \27483 );
and \U$27141 ( \27485 , \27479 , \27483 );
or \U$27142 ( \27486 , \27482 , \27484 , \27485 );
and \U$27143 ( \27487 , \27476 , \27486 );
and \U$27144 ( \27488 , \27466 , \27486 );
or \U$27145 ( \27489 , \27477 , \27487 , \27488 );
and \U$27146 ( \27490 , \24836 , \21652 );
and \U$27147 ( \27491 , \24714 , \21650 );
nor \U$27148 ( \27492 , \27490 , \27491 );
xnor \U$27149 ( \27493 , \27492 , \21377 );
and \U$27150 ( \27494 , \25097 , \21385 );
and \U$27151 ( \27495 , \24841 , \21383 );
nor \U$27152 ( \27496 , \27494 , \27495 );
xnor \U$27153 ( \27497 , \27496 , \21392 );
and \U$27154 ( \27498 , \27493 , \27497 );
and \U$27155 ( \27499 , \25596 , \21401 );
and \U$27156 ( \27500 , \25294 , \21399 );
nor \U$27157 ( \27501 , \27499 , \27500 );
xnor \U$27158 ( \27502 , \27501 , \21408 );
and \U$27159 ( \27503 , \27497 , \27502 );
and \U$27160 ( \27504 , \27493 , \27502 );
or \U$27161 ( \27505 , \27498 , \27503 , \27504 );
and \U$27162 ( \27506 , \26073 , \21419 );
and \U$27163 ( \27507 , \25604 , \21417 );
nor \U$27164 ( \27508 , \27506 , \27507 );
xnor \U$27165 ( \27509 , \27508 , \21426 );
and \U$27166 ( \27510 , \26342 , \21434 );
and \U$27167 ( \27511 , \26078 , \21432 );
nor \U$27168 ( \27512 , \27510 , \27511 );
xnor \U$27169 ( \27513 , \27512 , \21441 );
and \U$27170 ( \27514 , \27509 , \27513 );
and \U$27171 ( \27515 , \26973 , \21450 );
and \U$27172 ( \27516 , \26601 , \21448 );
nor \U$27173 ( \27517 , \27515 , \27516 );
xnor \U$27174 ( \27518 , \27517 , \21457 );
and \U$27175 ( \27519 , \27513 , \27518 );
and \U$27176 ( \27520 , \27509 , \27518 );
or \U$27177 ( \27521 , \27514 , \27519 , \27520 );
and \U$27178 ( \27522 , \27505 , \27521 );
and \U$27179 ( \27523 , \27325 , \21469 );
and \U$27180 ( \27524 , \26982 , \21467 );
nor \U$27181 ( \27525 , \27523 , \27524 );
xnor \U$27182 ( \27526 , \27525 , \21476 );
buf \U$27183 ( \27527 , RIbb32ce8_178);
and \U$27184 ( \27528 , \27527 , \21464 );
or \U$27185 ( \27529 , \27526 , \27528 );
and \U$27186 ( \27530 , \27521 , \27529 );
and \U$27187 ( \27531 , \27505 , \27529 );
or \U$27188 ( \27532 , \27522 , \27530 , \27531 );
and \U$27189 ( \27533 , \21478 , \24857 );
and \U$27190 ( \27534 , \21463 , \24855 );
nor \U$27191 ( \27535 , \27533 , \27534 );
xnor \U$27192 ( \27536 , \27535 , \24611 );
and \U$27193 ( \27537 , \21750 , \24462 );
and \U$27194 ( \27538 , \21689 , \24460 );
nor \U$27195 ( \27539 , \27537 , \27538 );
xnor \U$27196 ( \27540 , \27539 , \24275 );
and \U$27197 ( \27541 , \27536 , \27540 );
and \U$27198 ( \27542 , \22011 , \24149 );
and \U$27199 ( \27543 , \21813 , \24147 );
nor \U$27200 ( \27544 , \27542 , \27543 );
xnor \U$27201 ( \27545 , \27544 , \23944 );
and \U$27202 ( \27546 , \27540 , \27545 );
and \U$27203 ( \27547 , \27536 , \27545 );
or \U$27204 ( \27548 , \27541 , \27546 , \27547 );
and \U$27205 ( \27549 , \21436 , \26005 );
and \U$27206 ( \27550 , \21413 , \26003 );
nor \U$27207 ( \27551 , \27549 , \27550 );
xnor \U$27208 ( \27552 , \27551 , \25817 );
and \U$27209 ( \27553 , \21452 , \25631 );
and \U$27210 ( \27554 , \21428 , \25629 );
nor \U$27211 ( \27555 , \27553 , \27554 );
xnor \U$27212 ( \27556 , \27555 , \25399 );
and \U$27213 ( \27557 , \27552 , \27556 );
and \U$27214 ( \27558 , \21471 , \25180 );
and \U$27215 ( \27559 , \21444 , \25178 );
nor \U$27216 ( \27560 , \27558 , \27559 );
xnor \U$27217 ( \27561 , \27560 , \25037 );
and \U$27218 ( \27562 , \27556 , \27561 );
and \U$27219 ( \27563 , \27552 , \27561 );
or \U$27220 ( \27564 , \27557 , \27562 , \27563 );
and \U$27221 ( \27565 , \27548 , \27564 );
xor \U$27222 ( \27566 , \26717 , \27250 );
xor \U$27223 ( \27567 , \27250 , \27251 );
not \U$27224 ( \27568 , \27567 );
and \U$27225 ( \27569 , \27566 , \27568 );
and \U$27226 ( \27570 , \21387 , \27569 );
not \U$27227 ( \27571 , \27570 );
xnor \U$27228 ( \27572 , \27571 , \27254 );
and \U$27229 ( \27573 , \21403 , \27060 );
and \U$27230 ( \27574 , \21379 , \27058 );
nor \U$27231 ( \27575 , \27573 , \27574 );
xnor \U$27232 ( \27576 , \27575 , \26720 );
and \U$27233 ( \27577 , \27572 , \27576 );
and \U$27234 ( \27578 , \21421 , \26471 );
and \U$27235 ( \27579 , \21395 , \26469 );
nor \U$27236 ( \27580 , \27578 , \27579 );
xnor \U$27237 ( \27581 , \27580 , \26230 );
and \U$27238 ( \27582 , \27576 , \27581 );
and \U$27239 ( \27583 , \27572 , \27581 );
or \U$27240 ( \27584 , \27577 , \27582 , \27583 );
and \U$27241 ( \27585 , \27564 , \27584 );
and \U$27242 ( \27586 , \27548 , \27584 );
or \U$27243 ( \27587 , \27565 , \27585 , \27586 );
and \U$27244 ( \27588 , \27532 , \27587 );
and \U$27245 ( \27589 , \22867 , \22919 );
and \U$27246 ( \27590 , \22624 , \22917 );
nor \U$27247 ( \27591 , \27589 , \27590 );
xnor \U$27248 ( \27592 , \27591 , \22767 );
and \U$27249 ( \27593 , \23058 , \22651 );
and \U$27250 ( \27594 , \22872 , \22649 );
nor \U$27251 ( \27595 , \27593 , \27594 );
xnor \U$27252 ( \27596 , \27595 , \22495 );
and \U$27253 ( \27597 , \27592 , \27596 );
and \U$27254 ( \27598 , \23466 , \22379 );
and \U$27255 ( \27599 , \23202 , \22377 );
nor \U$27256 ( \27600 , \27598 , \27599 );
xnor \U$27257 ( \27601 , \27600 , \22266 );
and \U$27258 ( \27602 , \27596 , \27601 );
and \U$27259 ( \27603 , \27592 , \27601 );
or \U$27260 ( \27604 , \27597 , \27602 , \27603 );
and \U$27261 ( \27605 , \23665 , \22185 );
and \U$27262 ( \27606 , \23491 , \22183 );
nor \U$27263 ( \27607 , \27605 , \27606 );
xnor \U$27264 ( \27608 , \27607 , \22049 );
and \U$27265 ( \27609 , \23970 , \21985 );
and \U$27266 ( \27610 , \23832 , \21983 );
nor \U$27267 ( \27611 , \27609 , \27610 );
xnor \U$27268 ( \27612 , \27611 , \21907 );
and \U$27269 ( \27613 , \27608 , \27612 );
and \U$27270 ( \27614 , \24506 , \21821 );
and \U$27271 ( \27615 , \24089 , \21819 );
nor \U$27272 ( \27616 , \27614 , \27615 );
xnor \U$27273 ( \27617 , \27616 , \21727 );
and \U$27274 ( \27618 , \27612 , \27617 );
and \U$27275 ( \27619 , \27608 , \27617 );
or \U$27276 ( \27620 , \27613 , \27618 , \27619 );
and \U$27277 ( \27621 , \27604 , \27620 );
and \U$27278 ( \27622 , \22204 , \23743 );
and \U$27279 ( \27623 , \22099 , \23741 );
nor \U$27280 ( \27624 , \27622 , \27623 );
xnor \U$27281 ( \27625 , \27624 , \23594 );
and \U$27282 ( \27626 , \22325 , \23421 );
and \U$27283 ( \27627 , \22209 , \23419 );
nor \U$27284 ( \27628 , \27626 , \27627 );
xnor \U$27285 ( \27629 , \27628 , \23279 );
and \U$27286 ( \27630 , \27625 , \27629 );
and \U$27287 ( \27631 , \22616 , \23125 );
and \U$27288 ( \27632 , \22440 , \23123 );
nor \U$27289 ( \27633 , \27631 , \27632 );
xnor \U$27290 ( \27634 , \27633 , \22988 );
and \U$27291 ( \27635 , \27629 , \27634 );
and \U$27292 ( \27636 , \27625 , \27634 );
or \U$27293 ( \27637 , \27630 , \27635 , \27636 );
and \U$27294 ( \27638 , \27620 , \27637 );
and \U$27295 ( \27639 , \27604 , \27637 );
or \U$27296 ( \27640 , \27621 , \27638 , \27639 );
and \U$27297 ( \27641 , \27587 , \27640 );
and \U$27298 ( \27642 , \27532 , \27640 );
or \U$27299 ( \27643 , \27588 , \27641 , \27642 );
and \U$27300 ( \27644 , \27489 , \27643 );
xor \U$27301 ( \27645 , \27202 , \27204 );
xor \U$27302 ( \27646 , \27645 , \27207 );
xor \U$27303 ( \27647 , \27212 , \27214 );
xor \U$27304 ( \27648 , \27647 , \27217 );
and \U$27305 ( \27649 , \27646 , \27648 );
xor \U$27306 ( \27650 , \27223 , \27225 );
xor \U$27307 ( \27651 , \27650 , \27227 );
and \U$27308 ( \27652 , \27648 , \27651 );
and \U$27309 ( \27653 , \27646 , \27651 );
or \U$27310 ( \27654 , \27649 , \27652 , \27653 );
and \U$27311 ( \27655 , \27643 , \27654 );
and \U$27312 ( \27656 , \27489 , \27654 );
or \U$27313 ( \27657 , \27644 , \27655 , \27656 );
xor \U$27314 ( \27658 , \27249 , \27267 );
xor \U$27315 ( \27659 , \27658 , \27284 );
xor \U$27316 ( \27660 , \27303 , \27319 );
xor \U$27317 ( \27661 , \27660 , \27327 );
and \U$27318 ( \27662 , \27659 , \27661 );
xor \U$27319 ( \27663 , \27347 , \27363 );
xor \U$27320 ( \27664 , \27663 , \27380 );
and \U$27321 ( \27665 , \27661 , \27664 );
and \U$27322 ( \27666 , \27659 , \27664 );
or \U$27323 ( \27667 , \27662 , \27665 , \27666 );
xor \U$27324 ( \27668 , \27402 , \27404 );
xor \U$27325 ( \27669 , \27668 , \27407 );
and \U$27326 ( \27670 , \27667 , \27669 );
xor \U$27327 ( \27671 , \27389 , \27391 );
xor \U$27328 ( \27672 , \27671 , \27394 );
and \U$27329 ( \27673 , \27669 , \27672 );
and \U$27330 ( \27674 , \27667 , \27672 );
or \U$27331 ( \27675 , \27670 , \27673 , \27674 );
and \U$27332 ( \27676 , \27657 , \27675 );
xor \U$27333 ( \27677 , \27210 , \27220 );
xor \U$27334 ( \27678 , \27677 , \27230 );
xor \U$27335 ( \27679 , \27287 , \27330 );
xor \U$27336 ( \27680 , \27679 , \27383 );
and \U$27337 ( \27681 , \27678 , \27680 );
and \U$27338 ( \27682 , \27675 , \27681 );
and \U$27339 ( \27683 , \27657 , \27681 );
or \U$27340 ( \27684 , \27676 , \27682 , \27683 );
xor \U$27341 ( \27685 , \27233 , \27386 );
xor \U$27342 ( \27686 , \27685 , \27397 );
xor \U$27343 ( \27687 , \27410 , \27412 );
xor \U$27344 ( \27688 , \27687 , \27415 );
and \U$27345 ( \27689 , \27686 , \27688 );
xor \U$27346 ( \27690 , \27421 , \27423 );
and \U$27347 ( \27691 , \27688 , \27690 );
and \U$27348 ( \27692 , \27686 , \27690 );
or \U$27349 ( \27693 , \27689 , \27691 , \27692 );
and \U$27350 ( \27694 , \27684 , \27693 );
xor \U$27351 ( \27695 , \27429 , \27431 );
xor \U$27352 ( \27696 , \27695 , \27433 );
and \U$27353 ( \27697 , \27693 , \27696 );
and \U$27354 ( \27698 , \27684 , \27696 );
or \U$27355 ( \27699 , \27694 , \27697 , \27698 );
xor \U$27356 ( \27700 , \27144 , \27161 );
xor \U$27357 ( \27701 , \27700 , \27167 );
and \U$27358 ( \27702 , \27699 , \27701 );
xor \U$27359 ( \27703 , \27427 , \27436 );
xor \U$27360 ( \27704 , \27703 , \27439 );
and \U$27361 ( \27705 , \27701 , \27704 );
and \U$27362 ( \27706 , \27699 , \27704 );
or \U$27363 ( \27707 , \27702 , \27705 , \27706 );
xor \U$27364 ( \27708 , \27442 , \27444 );
xor \U$27365 ( \27709 , \27708 , \27447 );
and \U$27366 ( \27710 , \27707 , \27709 );
and \U$27367 ( \27711 , \27456 , \27710 );
xor \U$27368 ( \27712 , \27456 , \27710 );
xor \U$27369 ( \27713 , \27707 , \27709 );
and \U$27370 ( \27714 , \22099 , \24149 );
and \U$27371 ( \27715 , \22011 , \24147 );
nor \U$27372 ( \27716 , \27714 , \27715 );
xnor \U$27373 ( \27717 , \27716 , \23944 );
and \U$27374 ( \27718 , \22209 , \23743 );
and \U$27375 ( \27719 , \22204 , \23741 );
nor \U$27376 ( \27720 , \27718 , \27719 );
xnor \U$27377 ( \27721 , \27720 , \23594 );
and \U$27378 ( \27722 , \27717 , \27721 );
and \U$27379 ( \27723 , \22440 , \23421 );
and \U$27380 ( \27724 , \22325 , \23419 );
nor \U$27381 ( \27725 , \27723 , \27724 );
xnor \U$27382 ( \27726 , \27725 , \23279 );
and \U$27383 ( \27727 , \27721 , \27726 );
and \U$27384 ( \27728 , \27717 , \27726 );
or \U$27385 ( \27729 , \27722 , \27727 , \27728 );
and \U$27386 ( \27730 , \22624 , \23125 );
and \U$27387 ( \27731 , \22616 , \23123 );
nor \U$27388 ( \27732 , \27730 , \27731 );
xnor \U$27389 ( \27733 , \27732 , \22988 );
and \U$27390 ( \27734 , \22872 , \22919 );
and \U$27391 ( \27735 , \22867 , \22917 );
nor \U$27392 ( \27736 , \27734 , \27735 );
xnor \U$27393 ( \27737 , \27736 , \22767 );
and \U$27394 ( \27738 , \27733 , \27737 );
and \U$27395 ( \27739 , \23202 , \22651 );
and \U$27396 ( \27740 , \23058 , \22649 );
nor \U$27397 ( \27741 , \27739 , \27740 );
xnor \U$27398 ( \27742 , \27741 , \22495 );
and \U$27399 ( \27743 , \27737 , \27742 );
and \U$27400 ( \27744 , \27733 , \27742 );
or \U$27401 ( \27745 , \27738 , \27743 , \27744 );
and \U$27402 ( \27746 , \27729 , \27745 );
and \U$27403 ( \27747 , \23491 , \22379 );
and \U$27404 ( \27748 , \23466 , \22377 );
nor \U$27405 ( \27749 , \27747 , \27748 );
xnor \U$27406 ( \27750 , \27749 , \22266 );
and \U$27407 ( \27751 , \23832 , \22185 );
and \U$27408 ( \27752 , \23665 , \22183 );
nor \U$27409 ( \27753 , \27751 , \27752 );
xnor \U$27410 ( \27754 , \27753 , \22049 );
and \U$27411 ( \27755 , \27750 , \27754 );
and \U$27412 ( \27756 , \24089 , \21985 );
and \U$27413 ( \27757 , \23970 , \21983 );
nor \U$27414 ( \27758 , \27756 , \27757 );
xnor \U$27415 ( \27759 , \27758 , \21907 );
and \U$27416 ( \27760 , \27754 , \27759 );
and \U$27417 ( \27761 , \27750 , \27759 );
or \U$27418 ( \27762 , \27755 , \27760 , \27761 );
and \U$27419 ( \27763 , \27745 , \27762 );
and \U$27420 ( \27764 , \27729 , \27762 );
or \U$27421 ( \27765 , \27746 , \27763 , \27764 );
and \U$27422 ( \27766 , \21413 , \26471 );
and \U$27423 ( \27767 , \21421 , \26469 );
nor \U$27424 ( \27768 , \27766 , \27767 );
xnor \U$27425 ( \27769 , \27768 , \26230 );
and \U$27426 ( \27770 , \21428 , \26005 );
and \U$27427 ( \27771 , \21436 , \26003 );
nor \U$27428 ( \27772 , \27770 , \27771 );
xnor \U$27429 ( \27773 , \27772 , \25817 );
and \U$27430 ( \27774 , \27769 , \27773 );
and \U$27431 ( \27775 , \21444 , \25631 );
and \U$27432 ( \27776 , \21452 , \25629 );
nor \U$27433 ( \27777 , \27775 , \27776 );
xnor \U$27434 ( \27778 , \27777 , \25399 );
and \U$27435 ( \27779 , \27773 , \27778 );
and \U$27436 ( \27780 , \27769 , \27778 );
or \U$27437 ( \27781 , \27774 , \27779 , \27780 );
and \U$27438 ( \27782 , \21463 , \25180 );
and \U$27439 ( \27783 , \21471 , \25178 );
nor \U$27440 ( \27784 , \27782 , \27783 );
xnor \U$27441 ( \27785 , \27784 , \25037 );
and \U$27442 ( \27786 , \21689 , \24857 );
and \U$27443 ( \27787 , \21478 , \24855 );
nor \U$27444 ( \27788 , \27786 , \27787 );
xnor \U$27445 ( \27789 , \27788 , \24611 );
and \U$27446 ( \27790 , \27785 , \27789 );
and \U$27447 ( \27791 , \21813 , \24462 );
and \U$27448 ( \27792 , \21750 , \24460 );
nor \U$27449 ( \27793 , \27791 , \27792 );
xnor \U$27450 ( \27794 , \27793 , \24275 );
and \U$27451 ( \27795 , \27789 , \27794 );
and \U$27452 ( \27796 , \27785 , \27794 );
or \U$27453 ( \27797 , \27790 , \27795 , \27796 );
and \U$27454 ( \27798 , \27781 , \27797 );
buf \U$27455 ( \27799 , RIbb2de28_52);
buf \U$27456 ( \27800 , RIbb2ddb0_53);
and \U$27457 ( \27801 , \27799 , \27800 );
not \U$27458 ( \27802 , \27801 );
and \U$27459 ( \27803 , \27251 , \27802 );
not \U$27460 ( \27804 , \27803 );
and \U$27461 ( \27805 , \21379 , \27569 );
and \U$27462 ( \27806 , \21387 , \27567 );
nor \U$27463 ( \27807 , \27805 , \27806 );
xnor \U$27464 ( \27808 , \27807 , \27254 );
and \U$27465 ( \27809 , \27804 , \27808 );
and \U$27466 ( \27810 , \21395 , \27060 );
and \U$27467 ( \27811 , \21403 , \27058 );
nor \U$27468 ( \27812 , \27810 , \27811 );
xnor \U$27469 ( \27813 , \27812 , \26720 );
and \U$27470 ( \27814 , \27808 , \27813 );
and \U$27471 ( \27815 , \27804 , \27813 );
or \U$27472 ( \27816 , \27809 , \27814 , \27815 );
and \U$27473 ( \27817 , \27797 , \27816 );
and \U$27474 ( \27818 , \27781 , \27816 );
or \U$27475 ( \27819 , \27798 , \27817 , \27818 );
and \U$27476 ( \27820 , \27765 , \27819 );
and \U$27477 ( \27821 , \26982 , \21450 );
and \U$27478 ( \27822 , \26973 , \21448 );
nor \U$27479 ( \27823 , \27821 , \27822 );
xnor \U$27480 ( \27824 , \27823 , \21457 );
and \U$27481 ( \27825 , \27527 , \21469 );
and \U$27482 ( \27826 , \27325 , \21467 );
nor \U$27483 ( \27827 , \27825 , \27826 );
xnor \U$27484 ( \27828 , \27827 , \21476 );
and \U$27485 ( \27829 , \27824 , \27828 );
buf \U$27486 ( \27830 , RIbb32d60_179);
and \U$27487 ( \27831 , \27830 , \21464 );
and \U$27488 ( \27832 , \27828 , \27831 );
and \U$27489 ( \27833 , \27824 , \27831 );
or \U$27490 ( \27834 , \27829 , \27832 , \27833 );
and \U$27491 ( \27835 , \24714 , \21821 );
and \U$27492 ( \27836 , \24506 , \21819 );
nor \U$27493 ( \27837 , \27835 , \27836 );
xnor \U$27494 ( \27838 , \27837 , \21727 );
and \U$27495 ( \27839 , \24841 , \21652 );
and \U$27496 ( \27840 , \24836 , \21650 );
nor \U$27497 ( \27841 , \27839 , \27840 );
xnor \U$27498 ( \27842 , \27841 , \21377 );
and \U$27499 ( \27843 , \27838 , \27842 );
and \U$27500 ( \27844 , \25294 , \21385 );
and \U$27501 ( \27845 , \25097 , \21383 );
nor \U$27502 ( \27846 , \27844 , \27845 );
xnor \U$27503 ( \27847 , \27846 , \21392 );
and \U$27504 ( \27848 , \27842 , \27847 );
and \U$27505 ( \27849 , \27838 , \27847 );
or \U$27506 ( \27850 , \27843 , \27848 , \27849 );
and \U$27507 ( \27851 , \27834 , \27850 );
and \U$27508 ( \27852 , \25604 , \21401 );
and \U$27509 ( \27853 , \25596 , \21399 );
nor \U$27510 ( \27854 , \27852 , \27853 );
xnor \U$27511 ( \27855 , \27854 , \21408 );
and \U$27512 ( \27856 , \26078 , \21419 );
and \U$27513 ( \27857 , \26073 , \21417 );
nor \U$27514 ( \27858 , \27856 , \27857 );
xnor \U$27515 ( \27859 , \27858 , \21426 );
and \U$27516 ( \27860 , \27855 , \27859 );
and \U$27517 ( \27861 , \26601 , \21434 );
and \U$27518 ( \27862 , \26342 , \21432 );
nor \U$27519 ( \27863 , \27861 , \27862 );
xnor \U$27520 ( \27864 , \27863 , \21441 );
and \U$27521 ( \27865 , \27859 , \27864 );
and \U$27522 ( \27866 , \27855 , \27864 );
or \U$27523 ( \27867 , \27860 , \27865 , \27866 );
and \U$27524 ( \27868 , \27850 , \27867 );
and \U$27525 ( \27869 , \27834 , \27867 );
or \U$27526 ( \27870 , \27851 , \27868 , \27869 );
and \U$27527 ( \27871 , \27819 , \27870 );
and \U$27528 ( \27872 , \27765 , \27870 );
or \U$27529 ( \27873 , \27820 , \27871 , \27872 );
xor \U$27530 ( \27874 , \27592 , \27596 );
xor \U$27531 ( \27875 , \27874 , \27601 );
xor \U$27532 ( \27876 , \27608 , \27612 );
xor \U$27533 ( \27877 , \27876 , \27617 );
and \U$27534 ( \27878 , \27875 , \27877 );
xor \U$27535 ( \27879 , \27625 , \27629 );
xor \U$27536 ( \27880 , \27879 , \27634 );
and \U$27537 ( \27881 , \27877 , \27880 );
and \U$27538 ( \27882 , \27875 , \27880 );
or \U$27539 ( \27883 , \27878 , \27881 , \27882 );
xor \U$27540 ( \27884 , \27536 , \27540 );
xor \U$27541 ( \27885 , \27884 , \27545 );
xor \U$27542 ( \27886 , \27552 , \27556 );
xor \U$27543 ( \27887 , \27886 , \27561 );
and \U$27544 ( \27888 , \27885 , \27887 );
xor \U$27545 ( \27889 , \27572 , \27576 );
xor \U$27546 ( \27890 , \27889 , \27581 );
and \U$27547 ( \27891 , \27887 , \27890 );
and \U$27548 ( \27892 , \27885 , \27890 );
or \U$27549 ( \27893 , \27888 , \27891 , \27892 );
and \U$27550 ( \27894 , \27883 , \27893 );
xor \U$27551 ( \27895 , \27493 , \27497 );
xor \U$27552 ( \27896 , \27895 , \27502 );
xor \U$27553 ( \27897 , \27509 , \27513 );
xor \U$27554 ( \27898 , \27897 , \27518 );
and \U$27555 ( \27899 , \27896 , \27898 );
xnor \U$27556 ( \27900 , \27526 , \27528 );
and \U$27557 ( \27901 , \27898 , \27900 );
and \U$27558 ( \27902 , \27896 , \27900 );
or \U$27559 ( \27903 , \27899 , \27901 , \27902 );
and \U$27560 ( \27904 , \27893 , \27903 );
and \U$27561 ( \27905 , \27883 , \27903 );
or \U$27562 ( \27906 , \27894 , \27904 , \27905 );
and \U$27563 ( \27907 , \27873 , \27906 );
xor \U$27564 ( \27908 , \27458 , \27460 );
xor \U$27565 ( \27909 , \27908 , \27463 );
xor \U$27566 ( \27910 , \27468 , \27470 );
xor \U$27567 ( \27911 , \27910 , \27473 );
and \U$27568 ( \27912 , \27909 , \27911 );
xor \U$27569 ( \27913 , \27479 , \27481 );
xor \U$27570 ( \27914 , \27913 , \27483 );
and \U$27571 ( \27915 , \27911 , \27914 );
and \U$27572 ( \27916 , \27909 , \27914 );
or \U$27573 ( \27917 , \27912 , \27915 , \27916 );
and \U$27574 ( \27918 , \27906 , \27917 );
and \U$27575 ( \27919 , \27873 , \27917 );
or \U$27576 ( \27920 , \27907 , \27918 , \27919 );
xor \U$27577 ( \27921 , \27505 , \27521 );
xor \U$27578 ( \27922 , \27921 , \27529 );
xor \U$27579 ( \27923 , \27548 , \27564 );
xor \U$27580 ( \27924 , \27923 , \27584 );
and \U$27581 ( \27925 , \27922 , \27924 );
xor \U$27582 ( \27926 , \27604 , \27620 );
xor \U$27583 ( \27927 , \27926 , \27637 );
and \U$27584 ( \27928 , \27924 , \27927 );
and \U$27585 ( \27929 , \27922 , \27927 );
or \U$27586 ( \27930 , \27925 , \27928 , \27929 );
xor \U$27587 ( \27931 , \27659 , \27661 );
xor \U$27588 ( \27932 , \27931 , \27664 );
and \U$27589 ( \27933 , \27930 , \27932 );
xor \U$27590 ( \27934 , \27646 , \27648 );
xor \U$27591 ( \27935 , \27934 , \27651 );
and \U$27592 ( \27936 , \27932 , \27935 );
and \U$27593 ( \27937 , \27930 , \27935 );
or \U$27594 ( \27938 , \27933 , \27936 , \27937 );
and \U$27595 ( \27939 , \27920 , \27938 );
xor \U$27596 ( \27940 , \27466 , \27476 );
xor \U$27597 ( \27941 , \27940 , \27486 );
xor \U$27598 ( \27942 , \27532 , \27587 );
xor \U$27599 ( \27943 , \27942 , \27640 );
and \U$27600 ( \27944 , \27941 , \27943 );
and \U$27601 ( \27945 , \27938 , \27944 );
and \U$27602 ( \27946 , \27920 , \27944 );
or \U$27603 ( \27947 , \27939 , \27945 , \27946 );
xor \U$27604 ( \27948 , \27489 , \27643 );
xor \U$27605 ( \27949 , \27948 , \27654 );
xor \U$27606 ( \27950 , \27667 , \27669 );
xor \U$27607 ( \27951 , \27950 , \27672 );
and \U$27608 ( \27952 , \27949 , \27951 );
xor \U$27609 ( \27953 , \27678 , \27680 );
and \U$27610 ( \27954 , \27951 , \27953 );
and \U$27611 ( \27955 , \27949 , \27953 );
or \U$27612 ( \27956 , \27952 , \27954 , \27955 );
and \U$27613 ( \27957 , \27947 , \27956 );
xor \U$27614 ( \27958 , \27686 , \27688 );
xor \U$27615 ( \27959 , \27958 , \27690 );
and \U$27616 ( \27960 , \27956 , \27959 );
and \U$27617 ( \27961 , \27947 , \27959 );
or \U$27618 ( \27962 , \27957 , \27960 , \27961 );
xor \U$27619 ( \27963 , \27400 , \27418 );
xor \U$27620 ( \27964 , \27963 , \27424 );
and \U$27621 ( \27965 , \27962 , \27964 );
xor \U$27622 ( \27966 , \27684 , \27693 );
xor \U$27623 ( \27967 , \27966 , \27696 );
and \U$27624 ( \27968 , \27964 , \27967 );
and \U$27625 ( \27969 , \27962 , \27967 );
or \U$27626 ( \27970 , \27965 , \27968 , \27969 );
xor \U$27627 ( \27971 , \27699 , \27701 );
xor \U$27628 ( \27972 , \27971 , \27704 );
and \U$27629 ( \27973 , \27970 , \27972 );
and \U$27630 ( \27974 , \27713 , \27973 );
xor \U$27631 ( \27975 , \27713 , \27973 );
xor \U$27632 ( \27976 , \27970 , \27972 );
and \U$27633 ( \27977 , \24836 , \21821 );
and \U$27634 ( \27978 , \24714 , \21819 );
nor \U$27635 ( \27979 , \27977 , \27978 );
xnor \U$27636 ( \27980 , \27979 , \21727 );
and \U$27637 ( \27981 , \25097 , \21652 );
and \U$27638 ( \27982 , \24841 , \21650 );
nor \U$27639 ( \27983 , \27981 , \27982 );
xnor \U$27640 ( \27984 , \27983 , \21377 );
and \U$27641 ( \27985 , \27980 , \27984 );
and \U$27642 ( \27986 , \25596 , \21385 );
and \U$27643 ( \27987 , \25294 , \21383 );
nor \U$27644 ( \27988 , \27986 , \27987 );
xnor \U$27645 ( \27989 , \27988 , \21392 );
and \U$27646 ( \27990 , \27984 , \27989 );
and \U$27647 ( \27991 , \27980 , \27989 );
or \U$27648 ( \27992 , \27985 , \27990 , \27991 );
and \U$27649 ( \27993 , \27325 , \21450 );
and \U$27650 ( \27994 , \26982 , \21448 );
nor \U$27651 ( \27995 , \27993 , \27994 );
xnor \U$27652 ( \27996 , \27995 , \21457 );
and \U$27653 ( \27997 , \27830 , \21469 );
and \U$27654 ( \27998 , \27527 , \21467 );
nor \U$27655 ( \27999 , \27997 , \27998 );
xnor \U$27656 ( \28000 , \27999 , \21476 );
and \U$27657 ( \28001 , \27996 , \28000 );
buf \U$27658 ( \28002 , RIbb32dd8_180);
and \U$27659 ( \28003 , \28002 , \21464 );
and \U$27660 ( \28004 , \28000 , \28003 );
and \U$27661 ( \28005 , \27996 , \28003 );
or \U$27662 ( \28006 , \28001 , \28004 , \28005 );
and \U$27663 ( \28007 , \27992 , \28006 );
and \U$27664 ( \28008 , \26073 , \21401 );
and \U$27665 ( \28009 , \25604 , \21399 );
nor \U$27666 ( \28010 , \28008 , \28009 );
xnor \U$27667 ( \28011 , \28010 , \21408 );
and \U$27668 ( \28012 , \26342 , \21419 );
and \U$27669 ( \28013 , \26078 , \21417 );
nor \U$27670 ( \28014 , \28012 , \28013 );
xnor \U$27671 ( \28015 , \28014 , \21426 );
and \U$27672 ( \28016 , \28011 , \28015 );
and \U$27673 ( \28017 , \26973 , \21434 );
and \U$27674 ( \28018 , \26601 , \21432 );
nor \U$27675 ( \28019 , \28017 , \28018 );
xnor \U$27676 ( \28020 , \28019 , \21441 );
and \U$27677 ( \28021 , \28015 , \28020 );
and \U$27678 ( \28022 , \28011 , \28020 );
or \U$27679 ( \28023 , \28016 , \28021 , \28022 );
and \U$27680 ( \28024 , \28006 , \28023 );
and \U$27681 ( \28025 , \27992 , \28023 );
or \U$27682 ( \28026 , \28007 , \28024 , \28025 );
and \U$27683 ( \28027 , \21436 , \26471 );
and \U$27684 ( \28028 , \21413 , \26469 );
nor \U$27685 ( \28029 , \28027 , \28028 );
xnor \U$27686 ( \28030 , \28029 , \26230 );
and \U$27687 ( \28031 , \21452 , \26005 );
and \U$27688 ( \28032 , \21428 , \26003 );
nor \U$27689 ( \28033 , \28031 , \28032 );
xnor \U$27690 ( \28034 , \28033 , \25817 );
and \U$27691 ( \28035 , \28030 , \28034 );
and \U$27692 ( \28036 , \21471 , \25631 );
and \U$27693 ( \28037 , \21444 , \25629 );
nor \U$27694 ( \28038 , \28036 , \28037 );
xnor \U$27695 ( \28039 , \28038 , \25399 );
and \U$27696 ( \28040 , \28034 , \28039 );
and \U$27697 ( \28041 , \28030 , \28039 );
or \U$27698 ( \28042 , \28035 , \28040 , \28041 );
and \U$27699 ( \28043 , \21478 , \25180 );
and \U$27700 ( \28044 , \21463 , \25178 );
nor \U$27701 ( \28045 , \28043 , \28044 );
xnor \U$27702 ( \28046 , \28045 , \25037 );
and \U$27703 ( \28047 , \21750 , \24857 );
and \U$27704 ( \28048 , \21689 , \24855 );
nor \U$27705 ( \28049 , \28047 , \28048 );
xnor \U$27706 ( \28050 , \28049 , \24611 );
and \U$27707 ( \28051 , \28046 , \28050 );
and \U$27708 ( \28052 , \22011 , \24462 );
and \U$27709 ( \28053 , \21813 , \24460 );
nor \U$27710 ( \28054 , \28052 , \28053 );
xnor \U$27711 ( \28055 , \28054 , \24275 );
and \U$27712 ( \28056 , \28050 , \28055 );
and \U$27713 ( \28057 , \28046 , \28055 );
or \U$27714 ( \28058 , \28051 , \28056 , \28057 );
and \U$27715 ( \28059 , \28042 , \28058 );
xor \U$27716 ( \28060 , \27251 , \27799 );
xor \U$27717 ( \28061 , \27799 , \27800 );
not \U$27718 ( \28062 , \28061 );
and \U$27719 ( \28063 , \28060 , \28062 );
and \U$27720 ( \28064 , \21387 , \28063 );
not \U$27721 ( \28065 , \28064 );
xnor \U$27722 ( \28066 , \28065 , \27803 );
and \U$27723 ( \28067 , \21403 , \27569 );
and \U$27724 ( \28068 , \21379 , \27567 );
nor \U$27725 ( \28069 , \28067 , \28068 );
xnor \U$27726 ( \28070 , \28069 , \27254 );
and \U$27727 ( \28071 , \28066 , \28070 );
and \U$27728 ( \28072 , \21421 , \27060 );
and \U$27729 ( \28073 , \21395 , \27058 );
nor \U$27730 ( \28074 , \28072 , \28073 );
xnor \U$27731 ( \28075 , \28074 , \26720 );
and \U$27732 ( \28076 , \28070 , \28075 );
and \U$27733 ( \28077 , \28066 , \28075 );
or \U$27734 ( \28078 , \28071 , \28076 , \28077 );
and \U$27735 ( \28079 , \28058 , \28078 );
and \U$27736 ( \28080 , \28042 , \28078 );
or \U$27737 ( \28081 , \28059 , \28079 , \28080 );
and \U$27738 ( \28082 , \28026 , \28081 );
and \U$27739 ( \28083 , \22204 , \24149 );
and \U$27740 ( \28084 , \22099 , \24147 );
nor \U$27741 ( \28085 , \28083 , \28084 );
xnor \U$27742 ( \28086 , \28085 , \23944 );
and \U$27743 ( \28087 , \22325 , \23743 );
and \U$27744 ( \28088 , \22209 , \23741 );
nor \U$27745 ( \28089 , \28087 , \28088 );
xnor \U$27746 ( \28090 , \28089 , \23594 );
and \U$27747 ( \28091 , \28086 , \28090 );
and \U$27748 ( \28092 , \22616 , \23421 );
and \U$27749 ( \28093 , \22440 , \23419 );
nor \U$27750 ( \28094 , \28092 , \28093 );
xnor \U$27751 ( \28095 , \28094 , \23279 );
and \U$27752 ( \28096 , \28090 , \28095 );
and \U$27753 ( \28097 , \28086 , \28095 );
or \U$27754 ( \28098 , \28091 , \28096 , \28097 );
and \U$27755 ( \28099 , \22867 , \23125 );
and \U$27756 ( \28100 , \22624 , \23123 );
nor \U$27757 ( \28101 , \28099 , \28100 );
xnor \U$27758 ( \28102 , \28101 , \22988 );
and \U$27759 ( \28103 , \23058 , \22919 );
and \U$27760 ( \28104 , \22872 , \22917 );
nor \U$27761 ( \28105 , \28103 , \28104 );
xnor \U$27762 ( \28106 , \28105 , \22767 );
and \U$27763 ( \28107 , \28102 , \28106 );
and \U$27764 ( \28108 , \23466 , \22651 );
and \U$27765 ( \28109 , \23202 , \22649 );
nor \U$27766 ( \28110 , \28108 , \28109 );
xnor \U$27767 ( \28111 , \28110 , \22495 );
and \U$27768 ( \28112 , \28106 , \28111 );
and \U$27769 ( \28113 , \28102 , \28111 );
or \U$27770 ( \28114 , \28107 , \28112 , \28113 );
and \U$27771 ( \28115 , \28098 , \28114 );
and \U$27772 ( \28116 , \23665 , \22379 );
and \U$27773 ( \28117 , \23491 , \22377 );
nor \U$27774 ( \28118 , \28116 , \28117 );
xnor \U$27775 ( \28119 , \28118 , \22266 );
and \U$27776 ( \28120 , \23970 , \22185 );
and \U$27777 ( \28121 , \23832 , \22183 );
nor \U$27778 ( \28122 , \28120 , \28121 );
xnor \U$27779 ( \28123 , \28122 , \22049 );
and \U$27780 ( \28124 , \28119 , \28123 );
and \U$27781 ( \28125 , \24506 , \21985 );
and \U$27782 ( \28126 , \24089 , \21983 );
nor \U$27783 ( \28127 , \28125 , \28126 );
xnor \U$27784 ( \28128 , \28127 , \21907 );
and \U$27785 ( \28129 , \28123 , \28128 );
and \U$27786 ( \28130 , \28119 , \28128 );
or \U$27787 ( \28131 , \28124 , \28129 , \28130 );
and \U$27788 ( \28132 , \28114 , \28131 );
and \U$27789 ( \28133 , \28098 , \28131 );
or \U$27790 ( \28134 , \28115 , \28132 , \28133 );
and \U$27791 ( \28135 , \28081 , \28134 );
and \U$27792 ( \28136 , \28026 , \28134 );
or \U$27793 ( \28137 , \28082 , \28135 , \28136 );
xor \U$27794 ( \28138 , \27824 , \27828 );
xor \U$27795 ( \28139 , \28138 , \27831 );
xor \U$27796 ( \28140 , \27838 , \27842 );
xor \U$27797 ( \28141 , \28140 , \27847 );
and \U$27798 ( \28142 , \28139 , \28141 );
xor \U$27799 ( \28143 , \27855 , \27859 );
xor \U$27800 ( \28144 , \28143 , \27864 );
and \U$27801 ( \28145 , \28141 , \28144 );
and \U$27802 ( \28146 , \28139 , \28144 );
or \U$27803 ( \28147 , \28142 , \28145 , \28146 );
xor \U$27804 ( \28148 , \27717 , \27721 );
xor \U$27805 ( \28149 , \28148 , \27726 );
xor \U$27806 ( \28150 , \27733 , \27737 );
xor \U$27807 ( \28151 , \28150 , \27742 );
and \U$27808 ( \28152 , \28149 , \28151 );
xor \U$27809 ( \28153 , \27750 , \27754 );
xor \U$27810 ( \28154 , \28153 , \27759 );
and \U$27811 ( \28155 , \28151 , \28154 );
and \U$27812 ( \28156 , \28149 , \28154 );
or \U$27813 ( \28157 , \28152 , \28155 , \28156 );
and \U$27814 ( \28158 , \28147 , \28157 );
xor \U$27815 ( \28159 , \27769 , \27773 );
xor \U$27816 ( \28160 , \28159 , \27778 );
xor \U$27817 ( \28161 , \27785 , \27789 );
xor \U$27818 ( \28162 , \28161 , \27794 );
and \U$27819 ( \28163 , \28160 , \28162 );
xor \U$27820 ( \28164 , \27804 , \27808 );
xor \U$27821 ( \28165 , \28164 , \27813 );
and \U$27822 ( \28166 , \28162 , \28165 );
and \U$27823 ( \28167 , \28160 , \28165 );
or \U$27824 ( \28168 , \28163 , \28166 , \28167 );
and \U$27825 ( \28169 , \28157 , \28168 );
and \U$27826 ( \28170 , \28147 , \28168 );
or \U$27827 ( \28171 , \28158 , \28169 , \28170 );
and \U$27828 ( \28172 , \28137 , \28171 );
xor \U$27829 ( \28173 , \27875 , \27877 );
xor \U$27830 ( \28174 , \28173 , \27880 );
xor \U$27831 ( \28175 , \27885 , \27887 );
xor \U$27832 ( \28176 , \28175 , \27890 );
and \U$27833 ( \28177 , \28174 , \28176 );
xor \U$27834 ( \28178 , \27896 , \27898 );
xor \U$27835 ( \28179 , \28178 , \27900 );
and \U$27836 ( \28180 , \28176 , \28179 );
and \U$27837 ( \28181 , \28174 , \28179 );
or \U$27838 ( \28182 , \28177 , \28180 , \28181 );
and \U$27839 ( \28183 , \28171 , \28182 );
and \U$27840 ( \28184 , \28137 , \28182 );
or \U$27841 ( \28185 , \28172 , \28183 , \28184 );
xor \U$27842 ( \28186 , \27729 , \27745 );
xor \U$27843 ( \28187 , \28186 , \27762 );
xor \U$27844 ( \28188 , \27781 , \27797 );
xor \U$27845 ( \28189 , \28188 , \27816 );
and \U$27846 ( \28190 , \28187 , \28189 );
xor \U$27847 ( \28191 , \27834 , \27850 );
xor \U$27848 ( \28192 , \28191 , \27867 );
and \U$27849 ( \28193 , \28189 , \28192 );
and \U$27850 ( \28194 , \28187 , \28192 );
or \U$27851 ( \28195 , \28190 , \28193 , \28194 );
xor \U$27852 ( \28196 , \27922 , \27924 );
xor \U$27853 ( \28197 , \28196 , \27927 );
and \U$27854 ( \28198 , \28195 , \28197 );
xor \U$27855 ( \28199 , \27909 , \27911 );
xor \U$27856 ( \28200 , \28199 , \27914 );
and \U$27857 ( \28201 , \28197 , \28200 );
and \U$27858 ( \28202 , \28195 , \28200 );
or \U$27859 ( \28203 , \28198 , \28201 , \28202 );
and \U$27860 ( \28204 , \28185 , \28203 );
xor \U$27861 ( \28205 , \27765 , \27819 );
xor \U$27862 ( \28206 , \28205 , \27870 );
xor \U$27863 ( \28207 , \27883 , \27893 );
xor \U$27864 ( \28208 , \28207 , \27903 );
and \U$27865 ( \28209 , \28206 , \28208 );
and \U$27866 ( \28210 , \28203 , \28209 );
and \U$27867 ( \28211 , \28185 , \28209 );
or \U$27868 ( \28212 , \28204 , \28210 , \28211 );
xor \U$27869 ( \28213 , \27873 , \27906 );
xor \U$27870 ( \28214 , \28213 , \27917 );
xor \U$27871 ( \28215 , \27930 , \27932 );
xor \U$27872 ( \28216 , \28215 , \27935 );
and \U$27873 ( \28217 , \28214 , \28216 );
xor \U$27874 ( \28218 , \27941 , \27943 );
and \U$27875 ( \28219 , \28216 , \28218 );
and \U$27876 ( \28220 , \28214 , \28218 );
or \U$27877 ( \28221 , \28217 , \28219 , \28220 );
and \U$27878 ( \28222 , \28212 , \28221 );
xor \U$27879 ( \28223 , \27949 , \27951 );
xor \U$27880 ( \28224 , \28223 , \27953 );
and \U$27881 ( \28225 , \28221 , \28224 );
and \U$27882 ( \28226 , \28212 , \28224 );
or \U$27883 ( \28227 , \28222 , \28225 , \28226 );
xor \U$27884 ( \28228 , \27657 , \27675 );
xor \U$27885 ( \28229 , \28228 , \27681 );
and \U$27886 ( \28230 , \28227 , \28229 );
xor \U$27887 ( \28231 , \27947 , \27956 );
xor \U$27888 ( \28232 , \28231 , \27959 );
and \U$27889 ( \28233 , \28229 , \28232 );
and \U$27890 ( \28234 , \28227 , \28232 );
or \U$27891 ( \28235 , \28230 , \28233 , \28234 );
xor \U$27892 ( \28236 , \27962 , \27964 );
xor \U$27893 ( \28237 , \28236 , \27967 );
and \U$27894 ( \28238 , \28235 , \28237 );
and \U$27895 ( \28239 , \27976 , \28238 );
xor \U$27896 ( \28240 , \27976 , \28238 );
xor \U$27897 ( \28241 , \28235 , \28237 );
xor \U$27898 ( \28242 , \28030 , \28034 );
xor \U$27899 ( \28243 , \28242 , \28039 );
xor \U$27900 ( \28244 , \28086 , \28090 );
xor \U$27901 ( \28245 , \28244 , \28095 );
and \U$27902 ( \28246 , \28243 , \28245 );
xor \U$27903 ( \28247 , \28046 , \28050 );
xor \U$27904 ( \28248 , \28247 , \28055 );
and \U$27905 ( \28249 , \28245 , \28248 );
and \U$27906 ( \28250 , \28243 , \28248 );
or \U$27907 ( \28251 , \28246 , \28249 , \28250 );
xor \U$27908 ( \28252 , \28102 , \28106 );
xor \U$27909 ( \28253 , \28252 , \28111 );
xor \U$27910 ( \28254 , \27980 , \27984 );
xor \U$27911 ( \28255 , \28254 , \27989 );
and \U$27912 ( \28256 , \28253 , \28255 );
xor \U$27913 ( \28257 , \28119 , \28123 );
xor \U$27914 ( \28258 , \28257 , \28128 );
and \U$27915 ( \28259 , \28255 , \28258 );
and \U$27916 ( \28260 , \28253 , \28258 );
or \U$27917 ( \28261 , \28256 , \28259 , \28260 );
and \U$27918 ( \28262 , \28251 , \28261 );
xor \U$27919 ( \28263 , \27996 , \28000 );
xor \U$27920 ( \28264 , \28263 , \28003 );
xor \U$27921 ( \28265 , \28011 , \28015 );
xor \U$27922 ( \28266 , \28265 , \28020 );
or \U$27923 ( \28267 , \28264 , \28266 );
and \U$27924 ( \28268 , \28261 , \28267 );
and \U$27925 ( \28269 , \28251 , \28267 );
or \U$27926 ( \28270 , \28262 , \28268 , \28269 );
and \U$27927 ( \28271 , \22624 , \23421 );
and \U$27928 ( \28272 , \22616 , \23419 );
nor \U$27929 ( \28273 , \28271 , \28272 );
xnor \U$27930 ( \28274 , \28273 , \23279 );
and \U$27931 ( \28275 , \22872 , \23125 );
and \U$27932 ( \28276 , \22867 , \23123 );
nor \U$27933 ( \28277 , \28275 , \28276 );
xnor \U$27934 ( \28278 , \28277 , \22988 );
and \U$27935 ( \28279 , \28274 , \28278 );
and \U$27936 ( \28280 , \23202 , \22919 );
and \U$27937 ( \28281 , \23058 , \22917 );
nor \U$27938 ( \28282 , \28280 , \28281 );
xnor \U$27939 ( \28283 , \28282 , \22767 );
and \U$27940 ( \28284 , \28278 , \28283 );
and \U$27941 ( \28285 , \28274 , \28283 );
or \U$27942 ( \28286 , \28279 , \28284 , \28285 );
and \U$27943 ( \28287 , \22099 , \24462 );
and \U$27944 ( \28288 , \22011 , \24460 );
nor \U$27945 ( \28289 , \28287 , \28288 );
xnor \U$27946 ( \28290 , \28289 , \24275 );
and \U$27947 ( \28291 , \22209 , \24149 );
and \U$27948 ( \28292 , \22204 , \24147 );
nor \U$27949 ( \28293 , \28291 , \28292 );
xnor \U$27950 ( \28294 , \28293 , \23944 );
and \U$27951 ( \28295 , \28290 , \28294 );
and \U$27952 ( \28296 , \22440 , \23743 );
and \U$27953 ( \28297 , \22325 , \23741 );
nor \U$27954 ( \28298 , \28296 , \28297 );
xnor \U$27955 ( \28299 , \28298 , \23594 );
and \U$27956 ( \28300 , \28294 , \28299 );
and \U$27957 ( \28301 , \28290 , \28299 );
or \U$27958 ( \28302 , \28295 , \28300 , \28301 );
and \U$27959 ( \28303 , \28286 , \28302 );
and \U$27960 ( \28304 , \23491 , \22651 );
and \U$27961 ( \28305 , \23466 , \22649 );
nor \U$27962 ( \28306 , \28304 , \28305 );
xnor \U$27963 ( \28307 , \28306 , \22495 );
and \U$27964 ( \28308 , \23832 , \22379 );
and \U$27965 ( \28309 , \23665 , \22377 );
nor \U$27966 ( \28310 , \28308 , \28309 );
xnor \U$27967 ( \28311 , \28310 , \22266 );
and \U$27968 ( \28312 , \28307 , \28311 );
and \U$27969 ( \28313 , \24089 , \22185 );
and \U$27970 ( \28314 , \23970 , \22183 );
nor \U$27971 ( \28315 , \28313 , \28314 );
xnor \U$27972 ( \28316 , \28315 , \22049 );
and \U$27973 ( \28317 , \28311 , \28316 );
and \U$27974 ( \28318 , \28307 , \28316 );
or \U$27975 ( \28319 , \28312 , \28317 , \28318 );
and \U$27976 ( \28320 , \28302 , \28319 );
and \U$27977 ( \28321 , \28286 , \28319 );
or \U$27978 ( \28322 , \28303 , \28320 , \28321 );
and \U$27979 ( \28323 , \21413 , \27060 );
and \U$27980 ( \28324 , \21421 , \27058 );
nor \U$27981 ( \28325 , \28323 , \28324 );
xnor \U$27982 ( \28326 , \28325 , \26720 );
and \U$27983 ( \28327 , \21428 , \26471 );
and \U$27984 ( \28328 , \21436 , \26469 );
nor \U$27985 ( \28329 , \28327 , \28328 );
xnor \U$27986 ( \28330 , \28329 , \26230 );
and \U$27987 ( \28331 , \28326 , \28330 );
and \U$27988 ( \28332 , \21444 , \26005 );
and \U$27989 ( \28333 , \21452 , \26003 );
nor \U$27990 ( \28334 , \28332 , \28333 );
xnor \U$27991 ( \28335 , \28334 , \25817 );
and \U$27992 ( \28336 , \28330 , \28335 );
and \U$27993 ( \28337 , \28326 , \28335 );
or \U$27994 ( \28338 , \28331 , \28336 , \28337 );
buf \U$27995 ( \28339 , RIbb2dd38_54);
buf \U$27996 ( \28340 , RIbb2dcc0_55);
and \U$27997 ( \28341 , \28339 , \28340 );
not \U$27998 ( \28342 , \28341 );
and \U$27999 ( \28343 , \27800 , \28342 );
not \U$28000 ( \28344 , \28343 );
and \U$28001 ( \28345 , \21379 , \28063 );
and \U$28002 ( \28346 , \21387 , \28061 );
nor \U$28003 ( \28347 , \28345 , \28346 );
xnor \U$28004 ( \28348 , \28347 , \27803 );
and \U$28005 ( \28349 , \28344 , \28348 );
and \U$28006 ( \28350 , \21395 , \27569 );
and \U$28007 ( \28351 , \21403 , \27567 );
nor \U$28008 ( \28352 , \28350 , \28351 );
xnor \U$28009 ( \28353 , \28352 , \27254 );
and \U$28010 ( \28354 , \28348 , \28353 );
and \U$28011 ( \28355 , \28344 , \28353 );
or \U$28012 ( \28356 , \28349 , \28354 , \28355 );
and \U$28013 ( \28357 , \28338 , \28356 );
and \U$28014 ( \28358 , \21463 , \25631 );
and \U$28015 ( \28359 , \21471 , \25629 );
nor \U$28016 ( \28360 , \28358 , \28359 );
xnor \U$28017 ( \28361 , \28360 , \25399 );
and \U$28018 ( \28362 , \21689 , \25180 );
and \U$28019 ( \28363 , \21478 , \25178 );
nor \U$28020 ( \28364 , \28362 , \28363 );
xnor \U$28021 ( \28365 , \28364 , \25037 );
and \U$28022 ( \28366 , \28361 , \28365 );
and \U$28023 ( \28367 , \21813 , \24857 );
and \U$28024 ( \28368 , \21750 , \24855 );
nor \U$28025 ( \28369 , \28367 , \28368 );
xnor \U$28026 ( \28370 , \28369 , \24611 );
and \U$28027 ( \28371 , \28365 , \28370 );
and \U$28028 ( \28372 , \28361 , \28370 );
or \U$28029 ( \28373 , \28366 , \28371 , \28372 );
and \U$28030 ( \28374 , \28356 , \28373 );
and \U$28031 ( \28375 , \28338 , \28373 );
or \U$28032 ( \28376 , \28357 , \28374 , \28375 );
and \U$28033 ( \28377 , \28322 , \28376 );
and \U$28034 ( \28378 , \24714 , \21985 );
and \U$28035 ( \28379 , \24506 , \21983 );
nor \U$28036 ( \28380 , \28378 , \28379 );
xnor \U$28037 ( \28381 , \28380 , \21907 );
and \U$28038 ( \28382 , \24841 , \21821 );
and \U$28039 ( \28383 , \24836 , \21819 );
nor \U$28040 ( \28384 , \28382 , \28383 );
xnor \U$28041 ( \28385 , \28384 , \21727 );
and \U$28042 ( \28386 , \28381 , \28385 );
and \U$28043 ( \28387 , \25294 , \21652 );
and \U$28044 ( \28388 , \25097 , \21650 );
nor \U$28045 ( \28389 , \28387 , \28388 );
xnor \U$28046 ( \28390 , \28389 , \21377 );
and \U$28047 ( \28391 , \28385 , \28390 );
and \U$28048 ( \28392 , \28381 , \28390 );
or \U$28049 ( \28393 , \28386 , \28391 , \28392 );
and \U$28050 ( \28394 , \25604 , \21385 );
and \U$28051 ( \28395 , \25596 , \21383 );
nor \U$28052 ( \28396 , \28394 , \28395 );
xnor \U$28053 ( \28397 , \28396 , \21392 );
and \U$28054 ( \28398 , \26078 , \21401 );
and \U$28055 ( \28399 , \26073 , \21399 );
nor \U$28056 ( \28400 , \28398 , \28399 );
xnor \U$28057 ( \28401 , \28400 , \21408 );
and \U$28058 ( \28402 , \28397 , \28401 );
and \U$28059 ( \28403 , \26601 , \21419 );
and \U$28060 ( \28404 , \26342 , \21417 );
nor \U$28061 ( \28405 , \28403 , \28404 );
xnor \U$28062 ( \28406 , \28405 , \21426 );
and \U$28063 ( \28407 , \28401 , \28406 );
and \U$28064 ( \28408 , \28397 , \28406 );
or \U$28065 ( \28409 , \28402 , \28407 , \28408 );
and \U$28066 ( \28410 , \28393 , \28409 );
and \U$28067 ( \28411 , \26982 , \21434 );
and \U$28068 ( \28412 , \26973 , \21432 );
nor \U$28069 ( \28413 , \28411 , \28412 );
xnor \U$28070 ( \28414 , \28413 , \21441 );
and \U$28071 ( \28415 , \27527 , \21450 );
and \U$28072 ( \28416 , \27325 , \21448 );
nor \U$28073 ( \28417 , \28415 , \28416 );
xnor \U$28074 ( \28418 , \28417 , \21457 );
and \U$28075 ( \28419 , \28414 , \28418 );
and \U$28076 ( \28420 , \28002 , \21469 );
and \U$28077 ( \28421 , \27830 , \21467 );
nor \U$28078 ( \28422 , \28420 , \28421 );
xnor \U$28079 ( \28423 , \28422 , \21476 );
and \U$28080 ( \28424 , \28418 , \28423 );
and \U$28081 ( \28425 , \28414 , \28423 );
or \U$28082 ( \28426 , \28419 , \28424 , \28425 );
and \U$28083 ( \28427 , \28409 , \28426 );
and \U$28084 ( \28428 , \28393 , \28426 );
or \U$28085 ( \28429 , \28410 , \28427 , \28428 );
and \U$28086 ( \28430 , \28376 , \28429 );
and \U$28087 ( \28431 , \28322 , \28429 );
or \U$28088 ( \28432 , \28377 , \28430 , \28431 );
and \U$28089 ( \28433 , \28270 , \28432 );
xor \U$28090 ( \28434 , \28139 , \28141 );
xor \U$28091 ( \28435 , \28434 , \28144 );
xor \U$28092 ( \28436 , \28149 , \28151 );
xor \U$28093 ( \28437 , \28436 , \28154 );
and \U$28094 ( \28438 , \28435 , \28437 );
xor \U$28095 ( \28439 , \28160 , \28162 );
xor \U$28096 ( \28440 , \28439 , \28165 );
and \U$28097 ( \28441 , \28437 , \28440 );
and \U$28098 ( \28442 , \28435 , \28440 );
or \U$28099 ( \28443 , \28438 , \28441 , \28442 );
and \U$28100 ( \28444 , \28432 , \28443 );
and \U$28101 ( \28445 , \28270 , \28443 );
or \U$28102 ( \28446 , \28433 , \28444 , \28445 );
xor \U$28103 ( \28447 , \27992 , \28006 );
xor \U$28104 ( \28448 , \28447 , \28023 );
xor \U$28105 ( \28449 , \28042 , \28058 );
xor \U$28106 ( \28450 , \28449 , \28078 );
and \U$28107 ( \28451 , \28448 , \28450 );
xor \U$28108 ( \28452 , \28098 , \28114 );
xor \U$28109 ( \28453 , \28452 , \28131 );
and \U$28110 ( \28454 , \28450 , \28453 );
and \U$28111 ( \28455 , \28448 , \28453 );
or \U$28112 ( \28456 , \28451 , \28454 , \28455 );
xor \U$28113 ( \28457 , \28187 , \28189 );
xor \U$28114 ( \28458 , \28457 , \28192 );
and \U$28115 ( \28459 , \28456 , \28458 );
xor \U$28116 ( \28460 , \28174 , \28176 );
xor \U$28117 ( \28461 , \28460 , \28179 );
and \U$28118 ( \28462 , \28458 , \28461 );
and \U$28119 ( \28463 , \28456 , \28461 );
or \U$28120 ( \28464 , \28459 , \28462 , \28463 );
and \U$28121 ( \28465 , \28446 , \28464 );
xor \U$28122 ( \28466 , \28026 , \28081 );
xor \U$28123 ( \28467 , \28466 , \28134 );
xor \U$28124 ( \28468 , \28147 , \28157 );
xor \U$28125 ( \28469 , \28468 , \28168 );
and \U$28126 ( \28470 , \28467 , \28469 );
and \U$28127 ( \28471 , \28464 , \28470 );
and \U$28128 ( \28472 , \28446 , \28470 );
or \U$28129 ( \28473 , \28465 , \28471 , \28472 );
xor \U$28130 ( \28474 , \28137 , \28171 );
xor \U$28131 ( \28475 , \28474 , \28182 );
xor \U$28132 ( \28476 , \28195 , \28197 );
xor \U$28133 ( \28477 , \28476 , \28200 );
and \U$28134 ( \28478 , \28475 , \28477 );
xor \U$28135 ( \28479 , \28206 , \28208 );
and \U$28136 ( \28480 , \28477 , \28479 );
and \U$28137 ( \28481 , \28475 , \28479 );
or \U$28138 ( \28482 , \28478 , \28480 , \28481 );
and \U$28139 ( \28483 , \28473 , \28482 );
xor \U$28140 ( \28484 , \28214 , \28216 );
xor \U$28141 ( \28485 , \28484 , \28218 );
and \U$28142 ( \28486 , \28482 , \28485 );
and \U$28143 ( \28487 , \28473 , \28485 );
or \U$28144 ( \28488 , \28483 , \28486 , \28487 );
xor \U$28145 ( \28489 , \27920 , \27938 );
xor \U$28146 ( \28490 , \28489 , \27944 );
and \U$28147 ( \28491 , \28488 , \28490 );
xor \U$28148 ( \28492 , \28212 , \28221 );
xor \U$28149 ( \28493 , \28492 , \28224 );
and \U$28150 ( \28494 , \28490 , \28493 );
and \U$28151 ( \28495 , \28488 , \28493 );
or \U$28152 ( \28496 , \28491 , \28494 , \28495 );
xor \U$28153 ( \28497 , \28227 , \28229 );
xor \U$28154 ( \28498 , \28497 , \28232 );
and \U$28155 ( \28499 , \28496 , \28498 );
and \U$28156 ( \28500 , \28241 , \28499 );
xor \U$28157 ( \28501 , \28241 , \28499 );
xor \U$28158 ( \28502 , \28496 , \28498 );
and \U$28159 ( \28503 , \24836 , \21985 );
and \U$28160 ( \28504 , \24714 , \21983 );
nor \U$28161 ( \28505 , \28503 , \28504 );
xnor \U$28162 ( \28506 , \28505 , \21907 );
and \U$28163 ( \28507 , \25097 , \21821 );
and \U$28164 ( \28508 , \24841 , \21819 );
nor \U$28165 ( \28509 , \28507 , \28508 );
xnor \U$28166 ( \28510 , \28509 , \21727 );
and \U$28167 ( \28511 , \28506 , \28510 );
and \U$28168 ( \28512 , \25596 , \21652 );
and \U$28169 ( \28513 , \25294 , \21650 );
nor \U$28170 ( \28514 , \28512 , \28513 );
xnor \U$28171 ( \28515 , \28514 , \21377 );
and \U$28172 ( \28516 , \28510 , \28515 );
and \U$28173 ( \28517 , \28506 , \28515 );
or \U$28174 ( \28518 , \28511 , \28516 , \28517 );
and \U$28175 ( \28519 , \27325 , \21434 );
and \U$28176 ( \28520 , \26982 , \21432 );
nor \U$28177 ( \28521 , \28519 , \28520 );
xnor \U$28178 ( \28522 , \28521 , \21441 );
and \U$28179 ( \28523 , \27830 , \21450 );
and \U$28180 ( \28524 , \27527 , \21448 );
nor \U$28181 ( \28525 , \28523 , \28524 );
xnor \U$28182 ( \28526 , \28525 , \21457 );
and \U$28183 ( \28527 , \28522 , \28526 );
buf \U$28184 ( \28528 , RIbb32e50_181);
and \U$28185 ( \28529 , \28528 , \21469 );
and \U$28186 ( \28530 , \28002 , \21467 );
nor \U$28187 ( \28531 , \28529 , \28530 );
xnor \U$28188 ( \28532 , \28531 , \21476 );
and \U$28189 ( \28533 , \28526 , \28532 );
and \U$28190 ( \28534 , \28522 , \28532 );
or \U$28191 ( \28535 , \28527 , \28533 , \28534 );
and \U$28192 ( \28536 , \28518 , \28535 );
and \U$28193 ( \28537 , \26073 , \21385 );
and \U$28194 ( \28538 , \25604 , \21383 );
nor \U$28195 ( \28539 , \28537 , \28538 );
xnor \U$28196 ( \28540 , \28539 , \21392 );
and \U$28197 ( \28541 , \26342 , \21401 );
and \U$28198 ( \28542 , \26078 , \21399 );
nor \U$28199 ( \28543 , \28541 , \28542 );
xnor \U$28200 ( \28544 , \28543 , \21408 );
and \U$28201 ( \28545 , \28540 , \28544 );
and \U$28202 ( \28546 , \26973 , \21419 );
and \U$28203 ( \28547 , \26601 , \21417 );
nor \U$28204 ( \28548 , \28546 , \28547 );
xnor \U$28205 ( \28549 , \28548 , \21426 );
and \U$28206 ( \28550 , \28544 , \28549 );
and \U$28207 ( \28551 , \28540 , \28549 );
or \U$28208 ( \28552 , \28545 , \28550 , \28551 );
and \U$28209 ( \28553 , \28535 , \28552 );
and \U$28210 ( \28554 , \28518 , \28552 );
or \U$28211 ( \28555 , \28536 , \28553 , \28554 );
and \U$28212 ( \28556 , \21436 , \27060 );
and \U$28213 ( \28557 , \21413 , \27058 );
nor \U$28214 ( \28558 , \28556 , \28557 );
xnor \U$28215 ( \28559 , \28558 , \26720 );
and \U$28216 ( \28560 , \21452 , \26471 );
and \U$28217 ( \28561 , \21428 , \26469 );
nor \U$28218 ( \28562 , \28560 , \28561 );
xnor \U$28219 ( \28563 , \28562 , \26230 );
and \U$28220 ( \28564 , \28559 , \28563 );
and \U$28221 ( \28565 , \21471 , \26005 );
and \U$28222 ( \28566 , \21444 , \26003 );
nor \U$28223 ( \28567 , \28565 , \28566 );
xnor \U$28224 ( \28568 , \28567 , \25817 );
and \U$28225 ( \28569 , \28563 , \28568 );
and \U$28226 ( \28570 , \28559 , \28568 );
or \U$28227 ( \28571 , \28564 , \28569 , \28570 );
and \U$28228 ( \28572 , \21478 , \25631 );
and \U$28229 ( \28573 , \21463 , \25629 );
nor \U$28230 ( \28574 , \28572 , \28573 );
xnor \U$28231 ( \28575 , \28574 , \25399 );
and \U$28232 ( \28576 , \21750 , \25180 );
and \U$28233 ( \28577 , \21689 , \25178 );
nor \U$28234 ( \28578 , \28576 , \28577 );
xnor \U$28235 ( \28579 , \28578 , \25037 );
and \U$28236 ( \28580 , \28575 , \28579 );
and \U$28237 ( \28581 , \22011 , \24857 );
and \U$28238 ( \28582 , \21813 , \24855 );
nor \U$28239 ( \28583 , \28581 , \28582 );
xnor \U$28240 ( \28584 , \28583 , \24611 );
and \U$28241 ( \28585 , \28579 , \28584 );
and \U$28242 ( \28586 , \28575 , \28584 );
or \U$28243 ( \28587 , \28580 , \28585 , \28586 );
and \U$28244 ( \28588 , \28571 , \28587 );
xor \U$28245 ( \28589 , \27800 , \28339 );
xor \U$28246 ( \28590 , \28339 , \28340 );
not \U$28247 ( \28591 , \28590 );
and \U$28248 ( \28592 , \28589 , \28591 );
and \U$28249 ( \28593 , \21387 , \28592 );
not \U$28250 ( \28594 , \28593 );
xnor \U$28251 ( \28595 , \28594 , \28343 );
and \U$28252 ( \28596 , \21403 , \28063 );
and \U$28253 ( \28597 , \21379 , \28061 );
nor \U$28254 ( \28598 , \28596 , \28597 );
xnor \U$28255 ( \28599 , \28598 , \27803 );
and \U$28256 ( \28600 , \28595 , \28599 );
and \U$28257 ( \28601 , \21421 , \27569 );
and \U$28258 ( \28602 , \21395 , \27567 );
nor \U$28259 ( \28603 , \28601 , \28602 );
xnor \U$28260 ( \28604 , \28603 , \27254 );
and \U$28261 ( \28605 , \28599 , \28604 );
and \U$28262 ( \28606 , \28595 , \28604 );
or \U$28263 ( \28607 , \28600 , \28605 , \28606 );
and \U$28264 ( \28608 , \28587 , \28607 );
and \U$28265 ( \28609 , \28571 , \28607 );
or \U$28266 ( \28610 , \28588 , \28608 , \28609 );
and \U$28267 ( \28611 , \28555 , \28610 );
and \U$28268 ( \28612 , \23665 , \22651 );
and \U$28269 ( \28613 , \23491 , \22649 );
nor \U$28270 ( \28614 , \28612 , \28613 );
xnor \U$28271 ( \28615 , \28614 , \22495 );
and \U$28272 ( \28616 , \23970 , \22379 );
and \U$28273 ( \28617 , \23832 , \22377 );
nor \U$28274 ( \28618 , \28616 , \28617 );
xnor \U$28275 ( \28619 , \28618 , \22266 );
and \U$28276 ( \28620 , \28615 , \28619 );
and \U$28277 ( \28621 , \24506 , \22185 );
and \U$28278 ( \28622 , \24089 , \22183 );
nor \U$28279 ( \28623 , \28621 , \28622 );
xnor \U$28280 ( \28624 , \28623 , \22049 );
and \U$28281 ( \28625 , \28619 , \28624 );
and \U$28282 ( \28626 , \28615 , \28624 );
or \U$28283 ( \28627 , \28620 , \28625 , \28626 );
and \U$28284 ( \28628 , \22204 , \24462 );
and \U$28285 ( \28629 , \22099 , \24460 );
nor \U$28286 ( \28630 , \28628 , \28629 );
xnor \U$28287 ( \28631 , \28630 , \24275 );
and \U$28288 ( \28632 , \22325 , \24149 );
and \U$28289 ( \28633 , \22209 , \24147 );
nor \U$28290 ( \28634 , \28632 , \28633 );
xnor \U$28291 ( \28635 , \28634 , \23944 );
and \U$28292 ( \28636 , \28631 , \28635 );
and \U$28293 ( \28637 , \22616 , \23743 );
and \U$28294 ( \28638 , \22440 , \23741 );
nor \U$28295 ( \28639 , \28637 , \28638 );
xnor \U$28296 ( \28640 , \28639 , \23594 );
and \U$28297 ( \28641 , \28635 , \28640 );
and \U$28298 ( \28642 , \28631 , \28640 );
or \U$28299 ( \28643 , \28636 , \28641 , \28642 );
and \U$28300 ( \28644 , \28627 , \28643 );
and \U$28301 ( \28645 , \22867 , \23421 );
and \U$28302 ( \28646 , \22624 , \23419 );
nor \U$28303 ( \28647 , \28645 , \28646 );
xnor \U$28304 ( \28648 , \28647 , \23279 );
and \U$28305 ( \28649 , \23058 , \23125 );
and \U$28306 ( \28650 , \22872 , \23123 );
nor \U$28307 ( \28651 , \28649 , \28650 );
xnor \U$28308 ( \28652 , \28651 , \22988 );
and \U$28309 ( \28653 , \28648 , \28652 );
and \U$28310 ( \28654 , \23466 , \22919 );
and \U$28311 ( \28655 , \23202 , \22917 );
nor \U$28312 ( \28656 , \28654 , \28655 );
xnor \U$28313 ( \28657 , \28656 , \22767 );
and \U$28314 ( \28658 , \28652 , \28657 );
and \U$28315 ( \28659 , \28648 , \28657 );
or \U$28316 ( \28660 , \28653 , \28658 , \28659 );
and \U$28317 ( \28661 , \28643 , \28660 );
and \U$28318 ( \28662 , \28627 , \28660 );
or \U$28319 ( \28663 , \28644 , \28661 , \28662 );
and \U$28320 ( \28664 , \28610 , \28663 );
and \U$28321 ( \28665 , \28555 , \28663 );
or \U$28322 ( \28666 , \28611 , \28664 , \28665 );
xor \U$28323 ( \28667 , \28326 , \28330 );
xor \U$28324 ( \28668 , \28667 , \28335 );
xor \U$28325 ( \28669 , \28290 , \28294 );
xor \U$28326 ( \28670 , \28669 , \28299 );
and \U$28327 ( \28671 , \28668 , \28670 );
xor \U$28328 ( \28672 , \28361 , \28365 );
xor \U$28329 ( \28673 , \28672 , \28370 );
and \U$28330 ( \28674 , \28670 , \28673 );
and \U$28331 ( \28675 , \28668 , \28673 );
or \U$28332 ( \28676 , \28671 , \28674 , \28675 );
and \U$28333 ( \28677 , \28528 , \21464 );
xor \U$28334 ( \28678 , \28397 , \28401 );
xor \U$28335 ( \28679 , \28678 , \28406 );
and \U$28336 ( \28680 , \28677 , \28679 );
xor \U$28337 ( \28681 , \28414 , \28418 );
xor \U$28338 ( \28682 , \28681 , \28423 );
and \U$28339 ( \28683 , \28679 , \28682 );
and \U$28340 ( \28684 , \28677 , \28682 );
or \U$28341 ( \28685 , \28680 , \28683 , \28684 );
and \U$28342 ( \28686 , \28676 , \28685 );
xor \U$28343 ( \28687 , \28381 , \28385 );
xor \U$28344 ( \28688 , \28687 , \28390 );
xor \U$28345 ( \28689 , \28274 , \28278 );
xor \U$28346 ( \28690 , \28689 , \28283 );
and \U$28347 ( \28691 , \28688 , \28690 );
xor \U$28348 ( \28692 , \28307 , \28311 );
xor \U$28349 ( \28693 , \28692 , \28316 );
and \U$28350 ( \28694 , \28690 , \28693 );
and \U$28351 ( \28695 , \28688 , \28693 );
or \U$28352 ( \28696 , \28691 , \28694 , \28695 );
and \U$28353 ( \28697 , \28685 , \28696 );
and \U$28354 ( \28698 , \28676 , \28696 );
or \U$28355 ( \28699 , \28686 , \28697 , \28698 );
and \U$28356 ( \28700 , \28666 , \28699 );
xor \U$28357 ( \28701 , \28066 , \28070 );
xor \U$28358 ( \28702 , \28701 , \28075 );
xor \U$28359 ( \28703 , \28243 , \28245 );
xor \U$28360 ( \28704 , \28703 , \28248 );
and \U$28361 ( \28705 , \28702 , \28704 );
xor \U$28362 ( \28706 , \28253 , \28255 );
xor \U$28363 ( \28707 , \28706 , \28258 );
and \U$28364 ( \28708 , \28704 , \28707 );
and \U$28365 ( \28709 , \28702 , \28707 );
or \U$28366 ( \28710 , \28705 , \28708 , \28709 );
and \U$28367 ( \28711 , \28699 , \28710 );
and \U$28368 ( \28712 , \28666 , \28710 );
or \U$28369 ( \28713 , \28700 , \28711 , \28712 );
xor \U$28370 ( \28714 , \28286 , \28302 );
xor \U$28371 ( \28715 , \28714 , \28319 );
xor \U$28372 ( \28716 , \28393 , \28409 );
xor \U$28373 ( \28717 , \28716 , \28426 );
and \U$28374 ( \28718 , \28715 , \28717 );
xnor \U$28375 ( \28719 , \28264 , \28266 );
and \U$28376 ( \28720 , \28717 , \28719 );
and \U$28377 ( \28721 , \28715 , \28719 );
or \U$28378 ( \28722 , \28718 , \28720 , \28721 );
xor \U$28379 ( \28723 , \28448 , \28450 );
xor \U$28380 ( \28724 , \28723 , \28453 );
and \U$28381 ( \28725 , \28722 , \28724 );
xor \U$28382 ( \28726 , \28435 , \28437 );
xor \U$28383 ( \28727 , \28726 , \28440 );
and \U$28384 ( \28728 , \28724 , \28727 );
and \U$28385 ( \28729 , \28722 , \28727 );
or \U$28386 ( \28730 , \28725 , \28728 , \28729 );
and \U$28387 ( \28731 , \28713 , \28730 );
xor \U$28388 ( \28732 , \28251 , \28261 );
xor \U$28389 ( \28733 , \28732 , \28267 );
xor \U$28390 ( \28734 , \28322 , \28376 );
xor \U$28391 ( \28735 , \28734 , \28429 );
and \U$28392 ( \28736 , \28733 , \28735 );
and \U$28393 ( \28737 , \28730 , \28736 );
and \U$28394 ( \28738 , \28713 , \28736 );
or \U$28395 ( \28739 , \28731 , \28737 , \28738 );
xor \U$28396 ( \28740 , \28270 , \28432 );
xor \U$28397 ( \28741 , \28740 , \28443 );
xor \U$28398 ( \28742 , \28456 , \28458 );
xor \U$28399 ( \28743 , \28742 , \28461 );
and \U$28400 ( \28744 , \28741 , \28743 );
xor \U$28401 ( \28745 , \28467 , \28469 );
and \U$28402 ( \28746 , \28743 , \28745 );
and \U$28403 ( \28747 , \28741 , \28745 );
or \U$28404 ( \28748 , \28744 , \28746 , \28747 );
and \U$28405 ( \28749 , \28739 , \28748 );
xor \U$28406 ( \28750 , \28475 , \28477 );
xor \U$28407 ( \28751 , \28750 , \28479 );
and \U$28408 ( \28752 , \28748 , \28751 );
and \U$28409 ( \28753 , \28739 , \28751 );
or \U$28410 ( \28754 , \28749 , \28752 , \28753 );
xor \U$28411 ( \28755 , \28185 , \28203 );
xor \U$28412 ( \28756 , \28755 , \28209 );
and \U$28413 ( \28757 , \28754 , \28756 );
xor \U$28414 ( \28758 , \28473 , \28482 );
xor \U$28415 ( \28759 , \28758 , \28485 );
and \U$28416 ( \28760 , \28756 , \28759 );
and \U$28417 ( \28761 , \28754 , \28759 );
or \U$28418 ( \28762 , \28757 , \28760 , \28761 );
xor \U$28419 ( \28763 , \28488 , \28490 );
xor \U$28420 ( \28764 , \28763 , \28493 );
and \U$28421 ( \28765 , \28762 , \28764 );
and \U$28422 ( \28766 , \28502 , \28765 );
xor \U$28423 ( \28767 , \28502 , \28765 );
xor \U$28424 ( \28768 , \28762 , \28764 );
and \U$28425 ( \28769 , \23491 , \22919 );
and \U$28426 ( \28770 , \23466 , \22917 );
nor \U$28427 ( \28771 , \28769 , \28770 );
xnor \U$28428 ( \28772 , \28771 , \22767 );
and \U$28429 ( \28773 , \23832 , \22651 );
and \U$28430 ( \28774 , \23665 , \22649 );
nor \U$28431 ( \28775 , \28773 , \28774 );
xnor \U$28432 ( \28776 , \28775 , \22495 );
and \U$28433 ( \28777 , \28772 , \28776 );
and \U$28434 ( \28778 , \24089 , \22379 );
and \U$28435 ( \28779 , \23970 , \22377 );
nor \U$28436 ( \28780 , \28778 , \28779 );
xnor \U$28437 ( \28781 , \28780 , \22266 );
and \U$28438 ( \28782 , \28776 , \28781 );
and \U$28439 ( \28783 , \28772 , \28781 );
or \U$28440 ( \28784 , \28777 , \28782 , \28783 );
and \U$28441 ( \28785 , \22099 , \24857 );
and \U$28442 ( \28786 , \22011 , \24855 );
nor \U$28443 ( \28787 , \28785 , \28786 );
xnor \U$28444 ( \28788 , \28787 , \24611 );
and \U$28445 ( \28789 , \22209 , \24462 );
and \U$28446 ( \28790 , \22204 , \24460 );
nor \U$28447 ( \28791 , \28789 , \28790 );
xnor \U$28448 ( \28792 , \28791 , \24275 );
and \U$28449 ( \28793 , \28788 , \28792 );
and \U$28450 ( \28794 , \22440 , \24149 );
and \U$28451 ( \28795 , \22325 , \24147 );
nor \U$28452 ( \28796 , \28794 , \28795 );
xnor \U$28453 ( \28797 , \28796 , \23944 );
and \U$28454 ( \28798 , \28792 , \28797 );
and \U$28455 ( \28799 , \28788 , \28797 );
or \U$28456 ( \28800 , \28793 , \28798 , \28799 );
and \U$28457 ( \28801 , \28784 , \28800 );
and \U$28458 ( \28802 , \22624 , \23743 );
and \U$28459 ( \28803 , \22616 , \23741 );
nor \U$28460 ( \28804 , \28802 , \28803 );
xnor \U$28461 ( \28805 , \28804 , \23594 );
and \U$28462 ( \28806 , \22872 , \23421 );
and \U$28463 ( \28807 , \22867 , \23419 );
nor \U$28464 ( \28808 , \28806 , \28807 );
xnor \U$28465 ( \28809 , \28808 , \23279 );
and \U$28466 ( \28810 , \28805 , \28809 );
and \U$28467 ( \28811 , \23202 , \23125 );
and \U$28468 ( \28812 , \23058 , \23123 );
nor \U$28469 ( \28813 , \28811 , \28812 );
xnor \U$28470 ( \28814 , \28813 , \22988 );
and \U$28471 ( \28815 , \28809 , \28814 );
and \U$28472 ( \28816 , \28805 , \28814 );
or \U$28473 ( \28817 , \28810 , \28815 , \28816 );
and \U$28474 ( \28818 , \28800 , \28817 );
and \U$28475 ( \28819 , \28784 , \28817 );
or \U$28476 ( \28820 , \28801 , \28818 , \28819 );
and \U$28477 ( \28821 , \21463 , \26005 );
and \U$28478 ( \28822 , \21471 , \26003 );
nor \U$28479 ( \28823 , \28821 , \28822 );
xnor \U$28480 ( \28824 , \28823 , \25817 );
and \U$28481 ( \28825 , \21689 , \25631 );
and \U$28482 ( \28826 , \21478 , \25629 );
nor \U$28483 ( \28827 , \28825 , \28826 );
xnor \U$28484 ( \28828 , \28827 , \25399 );
and \U$28485 ( \28829 , \28824 , \28828 );
and \U$28486 ( \28830 , \21813 , \25180 );
and \U$28487 ( \28831 , \21750 , \25178 );
nor \U$28488 ( \28832 , \28830 , \28831 );
xnor \U$28489 ( \28833 , \28832 , \25037 );
and \U$28490 ( \28834 , \28828 , \28833 );
and \U$28491 ( \28835 , \28824 , \28833 );
or \U$28492 ( \28836 , \28829 , \28834 , \28835 );
buf \U$28493 ( \28837 , RIbb2dc48_56);
buf \U$28494 ( \28838 , RIbb2dbd0_57);
and \U$28495 ( \28839 , \28837 , \28838 );
not \U$28496 ( \28840 , \28839 );
and \U$28497 ( \28841 , \28340 , \28840 );
not \U$28498 ( \28842 , \28841 );
and \U$28499 ( \28843 , \21379 , \28592 );
and \U$28500 ( \28844 , \21387 , \28590 );
nor \U$28501 ( \28845 , \28843 , \28844 );
xnor \U$28502 ( \28846 , \28845 , \28343 );
and \U$28503 ( \28847 , \28842 , \28846 );
and \U$28504 ( \28848 , \21395 , \28063 );
and \U$28505 ( \28849 , \21403 , \28061 );
nor \U$28506 ( \28850 , \28848 , \28849 );
xnor \U$28507 ( \28851 , \28850 , \27803 );
and \U$28508 ( \28852 , \28846 , \28851 );
and \U$28509 ( \28853 , \28842 , \28851 );
or \U$28510 ( \28854 , \28847 , \28852 , \28853 );
and \U$28511 ( \28855 , \28836 , \28854 );
and \U$28512 ( \28856 , \21413 , \27569 );
and \U$28513 ( \28857 , \21421 , \27567 );
nor \U$28514 ( \28858 , \28856 , \28857 );
xnor \U$28515 ( \28859 , \28858 , \27254 );
and \U$28516 ( \28860 , \21428 , \27060 );
and \U$28517 ( \28861 , \21436 , \27058 );
nor \U$28518 ( \28862 , \28860 , \28861 );
xnor \U$28519 ( \28863 , \28862 , \26720 );
and \U$28520 ( \28864 , \28859 , \28863 );
and \U$28521 ( \28865 , \21444 , \26471 );
and \U$28522 ( \28866 , \21452 , \26469 );
nor \U$28523 ( \28867 , \28865 , \28866 );
xnor \U$28524 ( \28868 , \28867 , \26230 );
and \U$28525 ( \28869 , \28863 , \28868 );
and \U$28526 ( \28870 , \28859 , \28868 );
or \U$28527 ( \28871 , \28864 , \28869 , \28870 );
and \U$28528 ( \28872 , \28854 , \28871 );
and \U$28529 ( \28873 , \28836 , \28871 );
or \U$28530 ( \28874 , \28855 , \28872 , \28873 );
and \U$28531 ( \28875 , \28820 , \28874 );
and \U$28532 ( \28876 , \25604 , \21652 );
and \U$28533 ( \28877 , \25596 , \21650 );
nor \U$28534 ( \28878 , \28876 , \28877 );
xnor \U$28535 ( \28879 , \28878 , \21377 );
and \U$28536 ( \28880 , \26078 , \21385 );
and \U$28537 ( \28881 , \26073 , \21383 );
nor \U$28538 ( \28882 , \28880 , \28881 );
xnor \U$28539 ( \28883 , \28882 , \21392 );
and \U$28540 ( \28884 , \28879 , \28883 );
and \U$28541 ( \28885 , \26601 , \21401 );
and \U$28542 ( \28886 , \26342 , \21399 );
nor \U$28543 ( \28887 , \28885 , \28886 );
xnor \U$28544 ( \28888 , \28887 , \21408 );
and \U$28545 ( \28889 , \28883 , \28888 );
and \U$28546 ( \28890 , \28879 , \28888 );
or \U$28547 ( \28891 , \28884 , \28889 , \28890 );
and \U$28548 ( \28892 , \26982 , \21419 );
and \U$28549 ( \28893 , \26973 , \21417 );
nor \U$28550 ( \28894 , \28892 , \28893 );
xnor \U$28551 ( \28895 , \28894 , \21426 );
and \U$28552 ( \28896 , \27527 , \21434 );
and \U$28553 ( \28897 , \27325 , \21432 );
nor \U$28554 ( \28898 , \28896 , \28897 );
xnor \U$28555 ( \28899 , \28898 , \21441 );
and \U$28556 ( \28900 , \28895 , \28899 );
and \U$28557 ( \28901 , \28002 , \21450 );
and \U$28558 ( \28902 , \27830 , \21448 );
nor \U$28559 ( \28903 , \28901 , \28902 );
xnor \U$28560 ( \28904 , \28903 , \21457 );
and \U$28561 ( \28905 , \28899 , \28904 );
and \U$28562 ( \28906 , \28895 , \28904 );
or \U$28563 ( \28907 , \28900 , \28905 , \28906 );
and \U$28564 ( \28908 , \28891 , \28907 );
and \U$28565 ( \28909 , \24714 , \22185 );
and \U$28566 ( \28910 , \24506 , \22183 );
nor \U$28567 ( \28911 , \28909 , \28910 );
xnor \U$28568 ( \28912 , \28911 , \22049 );
and \U$28569 ( \28913 , \24841 , \21985 );
and \U$28570 ( \28914 , \24836 , \21983 );
nor \U$28571 ( \28915 , \28913 , \28914 );
xnor \U$28572 ( \28916 , \28915 , \21907 );
and \U$28573 ( \28917 , \28912 , \28916 );
and \U$28574 ( \28918 , \25294 , \21821 );
and \U$28575 ( \28919 , \25097 , \21819 );
nor \U$28576 ( \28920 , \28918 , \28919 );
xnor \U$28577 ( \28921 , \28920 , \21727 );
and \U$28578 ( \28922 , \28916 , \28921 );
and \U$28579 ( \28923 , \28912 , \28921 );
or \U$28580 ( \28924 , \28917 , \28922 , \28923 );
and \U$28581 ( \28925 , \28907 , \28924 );
and \U$28582 ( \28926 , \28891 , \28924 );
or \U$28583 ( \28927 , \28908 , \28925 , \28926 );
and \U$28584 ( \28928 , \28874 , \28927 );
and \U$28585 ( \28929 , \28820 , \28927 );
or \U$28586 ( \28930 , \28875 , \28928 , \28929 );
xor \U$28587 ( \28931 , \28506 , \28510 );
xor \U$28588 ( \28932 , \28931 , \28515 );
xor \U$28589 ( \28933 , \28615 , \28619 );
xor \U$28590 ( \28934 , \28933 , \28624 );
and \U$28591 ( \28935 , \28932 , \28934 );
xor \U$28592 ( \28936 , \28540 , \28544 );
xor \U$28593 ( \28937 , \28936 , \28549 );
and \U$28594 ( \28938 , \28934 , \28937 );
and \U$28595 ( \28939 , \28932 , \28937 );
or \U$28596 ( \28940 , \28935 , \28938 , \28939 );
xor \U$28597 ( \28941 , \28575 , \28579 );
xor \U$28598 ( \28942 , \28941 , \28584 );
xor \U$28599 ( \28943 , \28631 , \28635 );
xor \U$28600 ( \28944 , \28943 , \28640 );
and \U$28601 ( \28945 , \28942 , \28944 );
xor \U$28602 ( \28946 , \28648 , \28652 );
xor \U$28603 ( \28947 , \28946 , \28657 );
and \U$28604 ( \28948 , \28944 , \28947 );
and \U$28605 ( \28949 , \28942 , \28947 );
or \U$28606 ( \28950 , \28945 , \28948 , \28949 );
and \U$28607 ( \28951 , \28940 , \28950 );
buf \U$28608 ( \28952 , RIbb32ec8_182);
and \U$28609 ( \28953 , \28952 , \21464 );
xor \U$28610 ( \28954 , \28522 , \28526 );
xor \U$28611 ( \28955 , \28954 , \28532 );
or \U$28612 ( \28956 , \28953 , \28955 );
and \U$28613 ( \28957 , \28950 , \28956 );
and \U$28614 ( \28958 , \28940 , \28956 );
or \U$28615 ( \28959 , \28951 , \28957 , \28958 );
and \U$28616 ( \28960 , \28930 , \28959 );
xor \U$28617 ( \28961 , \28344 , \28348 );
xor \U$28618 ( \28962 , \28961 , \28353 );
xor \U$28619 ( \28963 , \28668 , \28670 );
xor \U$28620 ( \28964 , \28963 , \28673 );
and \U$28621 ( \28965 , \28962 , \28964 );
xor \U$28622 ( \28966 , \28688 , \28690 );
xor \U$28623 ( \28967 , \28966 , \28693 );
and \U$28624 ( \28968 , \28964 , \28967 );
and \U$28625 ( \28969 , \28962 , \28967 );
or \U$28626 ( \28970 , \28965 , \28968 , \28969 );
and \U$28627 ( \28971 , \28959 , \28970 );
and \U$28628 ( \28972 , \28930 , \28970 );
or \U$28629 ( \28973 , \28960 , \28971 , \28972 );
xor \U$28630 ( \28974 , \28555 , \28610 );
xor \U$28631 ( \28975 , \28974 , \28663 );
xor \U$28632 ( \28976 , \28676 , \28685 );
xor \U$28633 ( \28977 , \28976 , \28696 );
and \U$28634 ( \28978 , \28975 , \28977 );
xor \U$28635 ( \28979 , \28702 , \28704 );
xor \U$28636 ( \28980 , \28979 , \28707 );
and \U$28637 ( \28981 , \28977 , \28980 );
and \U$28638 ( \28982 , \28975 , \28980 );
or \U$28639 ( \28983 , \28978 , \28981 , \28982 );
and \U$28640 ( \28984 , \28973 , \28983 );
xor \U$28641 ( \28985 , \28518 , \28535 );
xor \U$28642 ( \28986 , \28985 , \28552 );
xor \U$28643 ( \28987 , \28627 , \28643 );
xor \U$28644 ( \28988 , \28987 , \28660 );
and \U$28645 ( \28989 , \28986 , \28988 );
xor \U$28646 ( \28990 , \28677 , \28679 );
xor \U$28647 ( \28991 , \28990 , \28682 );
and \U$28648 ( \28992 , \28988 , \28991 );
and \U$28649 ( \28993 , \28986 , \28991 );
or \U$28650 ( \28994 , \28989 , \28992 , \28993 );
xor \U$28651 ( \28995 , \28338 , \28356 );
xor \U$28652 ( \28996 , \28995 , \28373 );
and \U$28653 ( \28997 , \28994 , \28996 );
xor \U$28654 ( \28998 , \28715 , \28717 );
xor \U$28655 ( \28999 , \28998 , \28719 );
and \U$28656 ( \29000 , \28996 , \28999 );
and \U$28657 ( \29001 , \28994 , \28999 );
or \U$28658 ( \29002 , \28997 , \29000 , \29001 );
and \U$28659 ( \29003 , \28983 , \29002 );
and \U$28660 ( \29004 , \28973 , \29002 );
or \U$28661 ( \29005 , \28984 , \29003 , \29004 );
xor \U$28662 ( \29006 , \28666 , \28699 );
xor \U$28663 ( \29007 , \29006 , \28710 );
xor \U$28664 ( \29008 , \28722 , \28724 );
xor \U$28665 ( \29009 , \29008 , \28727 );
and \U$28666 ( \29010 , \29007 , \29009 );
xor \U$28667 ( \29011 , \28733 , \28735 );
and \U$28668 ( \29012 , \29009 , \29011 );
and \U$28669 ( \29013 , \29007 , \29011 );
or \U$28670 ( \29014 , \29010 , \29012 , \29013 );
and \U$28671 ( \29015 , \29005 , \29014 );
xor \U$28672 ( \29016 , \28741 , \28743 );
xor \U$28673 ( \29017 , \29016 , \28745 );
and \U$28674 ( \29018 , \29014 , \29017 );
and \U$28675 ( \29019 , \29005 , \29017 );
or \U$28676 ( \29020 , \29015 , \29018 , \29019 );
xor \U$28677 ( \29021 , \28446 , \28464 );
xor \U$28678 ( \29022 , \29021 , \28470 );
and \U$28679 ( \29023 , \29020 , \29022 );
xor \U$28680 ( \29024 , \28739 , \28748 );
xor \U$28681 ( \29025 , \29024 , \28751 );
and \U$28682 ( \29026 , \29022 , \29025 );
and \U$28683 ( \29027 , \29020 , \29025 );
or \U$28684 ( \29028 , \29023 , \29026 , \29027 );
xor \U$28685 ( \29029 , \28754 , \28756 );
xor \U$28686 ( \29030 , \29029 , \28759 );
and \U$28687 ( \29031 , \29028 , \29030 );
and \U$28688 ( \29032 , \28768 , \29031 );
xor \U$28689 ( \29033 , \28768 , \29031 );
xor \U$28690 ( \29034 , \29028 , \29030 );
and \U$28691 ( \29035 , \22867 , \23743 );
and \U$28692 ( \29036 , \22624 , \23741 );
nor \U$28693 ( \29037 , \29035 , \29036 );
xnor \U$28694 ( \29038 , \29037 , \23594 );
and \U$28695 ( \29039 , \23058 , \23421 );
and \U$28696 ( \29040 , \22872 , \23419 );
nor \U$28697 ( \29041 , \29039 , \29040 );
xnor \U$28698 ( \29042 , \29041 , \23279 );
and \U$28699 ( \29043 , \29038 , \29042 );
and \U$28700 ( \29044 , \23466 , \23125 );
and \U$28701 ( \29045 , \23202 , \23123 );
nor \U$28702 ( \29046 , \29044 , \29045 );
xnor \U$28703 ( \29047 , \29046 , \22988 );
and \U$28704 ( \29048 , \29042 , \29047 );
and \U$28705 ( \29049 , \29038 , \29047 );
or \U$28706 ( \29050 , \29043 , \29048 , \29049 );
and \U$28707 ( \29051 , \23665 , \22919 );
and \U$28708 ( \29052 , \23491 , \22917 );
nor \U$28709 ( \29053 , \29051 , \29052 );
xnor \U$28710 ( \29054 , \29053 , \22767 );
and \U$28711 ( \29055 , \23970 , \22651 );
and \U$28712 ( \29056 , \23832 , \22649 );
nor \U$28713 ( \29057 , \29055 , \29056 );
xnor \U$28714 ( \29058 , \29057 , \22495 );
and \U$28715 ( \29059 , \29054 , \29058 );
and \U$28716 ( \29060 , \24506 , \22379 );
and \U$28717 ( \29061 , \24089 , \22377 );
nor \U$28718 ( \29062 , \29060 , \29061 );
xnor \U$28719 ( \29063 , \29062 , \22266 );
and \U$28720 ( \29064 , \29058 , \29063 );
and \U$28721 ( \29065 , \29054 , \29063 );
or \U$28722 ( \29066 , \29059 , \29064 , \29065 );
and \U$28723 ( \29067 , \29050 , \29066 );
and \U$28724 ( \29068 , \22204 , \24857 );
and \U$28725 ( \29069 , \22099 , \24855 );
nor \U$28726 ( \29070 , \29068 , \29069 );
xnor \U$28727 ( \29071 , \29070 , \24611 );
and \U$28728 ( \29072 , \22325 , \24462 );
and \U$28729 ( \29073 , \22209 , \24460 );
nor \U$28730 ( \29074 , \29072 , \29073 );
xnor \U$28731 ( \29075 , \29074 , \24275 );
and \U$28732 ( \29076 , \29071 , \29075 );
and \U$28733 ( \29077 , \22616 , \24149 );
and \U$28734 ( \29078 , \22440 , \24147 );
nor \U$28735 ( \29079 , \29077 , \29078 );
xnor \U$28736 ( \29080 , \29079 , \23944 );
and \U$28737 ( \29081 , \29075 , \29080 );
and \U$28738 ( \29082 , \29071 , \29080 );
or \U$28739 ( \29083 , \29076 , \29081 , \29082 );
and \U$28740 ( \29084 , \29066 , \29083 );
and \U$28741 ( \29085 , \29050 , \29083 );
or \U$28742 ( \29086 , \29067 , \29084 , \29085 );
and \U$28743 ( \29087 , \26073 , \21652 );
and \U$28744 ( \29088 , \25604 , \21650 );
nor \U$28745 ( \29089 , \29087 , \29088 );
xnor \U$28746 ( \29090 , \29089 , \21377 );
and \U$28747 ( \29091 , \26342 , \21385 );
and \U$28748 ( \29092 , \26078 , \21383 );
nor \U$28749 ( \29093 , \29091 , \29092 );
xnor \U$28750 ( \29094 , \29093 , \21392 );
and \U$28751 ( \29095 , \29090 , \29094 );
and \U$28752 ( \29096 , \26973 , \21401 );
and \U$28753 ( \29097 , \26601 , \21399 );
nor \U$28754 ( \29098 , \29096 , \29097 );
xnor \U$28755 ( \29099 , \29098 , \21408 );
and \U$28756 ( \29100 , \29094 , \29099 );
and \U$28757 ( \29101 , \29090 , \29099 );
or \U$28758 ( \29102 , \29095 , \29100 , \29101 );
and \U$28759 ( \29103 , \24836 , \22185 );
and \U$28760 ( \29104 , \24714 , \22183 );
nor \U$28761 ( \29105 , \29103 , \29104 );
xnor \U$28762 ( \29106 , \29105 , \22049 );
and \U$28763 ( \29107 , \25097 , \21985 );
and \U$28764 ( \29108 , \24841 , \21983 );
nor \U$28765 ( \29109 , \29107 , \29108 );
xnor \U$28766 ( \29110 , \29109 , \21907 );
and \U$28767 ( \29111 , \29106 , \29110 );
and \U$28768 ( \29112 , \25596 , \21821 );
and \U$28769 ( \29113 , \25294 , \21819 );
nor \U$28770 ( \29114 , \29112 , \29113 );
xnor \U$28771 ( \29115 , \29114 , \21727 );
and \U$28772 ( \29116 , \29110 , \29115 );
and \U$28773 ( \29117 , \29106 , \29115 );
or \U$28774 ( \29118 , \29111 , \29116 , \29117 );
and \U$28775 ( \29119 , \29102 , \29118 );
and \U$28776 ( \29120 , \27325 , \21419 );
and \U$28777 ( \29121 , \26982 , \21417 );
nor \U$28778 ( \29122 , \29120 , \29121 );
xnor \U$28779 ( \29123 , \29122 , \21426 );
and \U$28780 ( \29124 , \27830 , \21434 );
and \U$28781 ( \29125 , \27527 , \21432 );
nor \U$28782 ( \29126 , \29124 , \29125 );
xnor \U$28783 ( \29127 , \29126 , \21441 );
and \U$28784 ( \29128 , \29123 , \29127 );
and \U$28785 ( \29129 , \28528 , \21450 );
and \U$28786 ( \29130 , \28002 , \21448 );
nor \U$28787 ( \29131 , \29129 , \29130 );
xnor \U$28788 ( \29132 , \29131 , \21457 );
and \U$28789 ( \29133 , \29127 , \29132 );
and \U$28790 ( \29134 , \29123 , \29132 );
or \U$28791 ( \29135 , \29128 , \29133 , \29134 );
and \U$28792 ( \29136 , \29118 , \29135 );
and \U$28793 ( \29137 , \29102 , \29135 );
or \U$28794 ( \29138 , \29119 , \29136 , \29137 );
and \U$28795 ( \29139 , \29086 , \29138 );
and \U$28796 ( \29140 , \21478 , \26005 );
and \U$28797 ( \29141 , \21463 , \26003 );
nor \U$28798 ( \29142 , \29140 , \29141 );
xnor \U$28799 ( \29143 , \29142 , \25817 );
and \U$28800 ( \29144 , \21750 , \25631 );
and \U$28801 ( \29145 , \21689 , \25629 );
nor \U$28802 ( \29146 , \29144 , \29145 );
xnor \U$28803 ( \29147 , \29146 , \25399 );
and \U$28804 ( \29148 , \29143 , \29147 );
and \U$28805 ( \29149 , \22011 , \25180 );
and \U$28806 ( \29150 , \21813 , \25178 );
nor \U$28807 ( \29151 , \29149 , \29150 );
xnor \U$28808 ( \29152 , \29151 , \25037 );
and \U$28809 ( \29153 , \29147 , \29152 );
and \U$28810 ( \29154 , \29143 , \29152 );
or \U$28811 ( \29155 , \29148 , \29153 , \29154 );
xor \U$28812 ( \29156 , \28340 , \28837 );
xor \U$28813 ( \29157 , \28837 , \28838 );
not \U$28814 ( \29158 , \29157 );
and \U$28815 ( \29159 , \29156 , \29158 );
and \U$28816 ( \29160 , \21387 , \29159 );
not \U$28817 ( \29161 , \29160 );
xnor \U$28818 ( \29162 , \29161 , \28841 );
and \U$28819 ( \29163 , \21403 , \28592 );
and \U$28820 ( \29164 , \21379 , \28590 );
nor \U$28821 ( \29165 , \29163 , \29164 );
xnor \U$28822 ( \29166 , \29165 , \28343 );
and \U$28823 ( \29167 , \29162 , \29166 );
and \U$28824 ( \29168 , \21421 , \28063 );
and \U$28825 ( \29169 , \21395 , \28061 );
nor \U$28826 ( \29170 , \29168 , \29169 );
xnor \U$28827 ( \29171 , \29170 , \27803 );
and \U$28828 ( \29172 , \29166 , \29171 );
and \U$28829 ( \29173 , \29162 , \29171 );
or \U$28830 ( \29174 , \29167 , \29172 , \29173 );
and \U$28831 ( \29175 , \29155 , \29174 );
and \U$28832 ( \29176 , \21436 , \27569 );
and \U$28833 ( \29177 , \21413 , \27567 );
nor \U$28834 ( \29178 , \29176 , \29177 );
xnor \U$28835 ( \29179 , \29178 , \27254 );
and \U$28836 ( \29180 , \21452 , \27060 );
and \U$28837 ( \29181 , \21428 , \27058 );
nor \U$28838 ( \29182 , \29180 , \29181 );
xnor \U$28839 ( \29183 , \29182 , \26720 );
and \U$28840 ( \29184 , \29179 , \29183 );
and \U$28841 ( \29185 , \21471 , \26471 );
and \U$28842 ( \29186 , \21444 , \26469 );
nor \U$28843 ( \29187 , \29185 , \29186 );
xnor \U$28844 ( \29188 , \29187 , \26230 );
and \U$28845 ( \29189 , \29183 , \29188 );
and \U$28846 ( \29190 , \29179 , \29188 );
or \U$28847 ( \29191 , \29184 , \29189 , \29190 );
and \U$28848 ( \29192 , \29174 , \29191 );
and \U$28849 ( \29193 , \29155 , \29191 );
or \U$28850 ( \29194 , \29175 , \29192 , \29193 );
and \U$28851 ( \29195 , \29138 , \29194 );
and \U$28852 ( \29196 , \29086 , \29194 );
or \U$28853 ( \29197 , \29139 , \29195 , \29196 );
buf \U$28854 ( \29198 , RIbb32f40_183);
and \U$28855 ( \29199 , \29198 , \21469 );
and \U$28856 ( \29200 , \28952 , \21467 );
nor \U$28857 ( \29201 , \29199 , \29200 );
xnor \U$28858 ( \29202 , \29201 , \21476 );
buf \U$28859 ( \29203 , RIbb32fb8_184);
and \U$28860 ( \29204 , \29203 , \21464 );
or \U$28861 ( \29205 , \29202 , \29204 );
and \U$28862 ( \29206 , \28952 , \21469 );
and \U$28863 ( \29207 , \28528 , \21467 );
nor \U$28864 ( \29208 , \29206 , \29207 );
xnor \U$28865 ( \29209 , \29208 , \21476 );
and \U$28866 ( \29210 , \29205 , \29209 );
and \U$28867 ( \29211 , \29198 , \21464 );
and \U$28868 ( \29212 , \29209 , \29211 );
and \U$28869 ( \29213 , \29205 , \29211 );
or \U$28870 ( \29214 , \29210 , \29212 , \29213 );
xor \U$28871 ( \29215 , \28879 , \28883 );
xor \U$28872 ( \29216 , \29215 , \28888 );
xor \U$28873 ( \29217 , \28895 , \28899 );
xor \U$28874 ( \29218 , \29217 , \28904 );
and \U$28875 ( \29219 , \29216 , \29218 );
xor \U$28876 ( \29220 , \28912 , \28916 );
xor \U$28877 ( \29221 , \29220 , \28921 );
and \U$28878 ( \29222 , \29218 , \29221 );
and \U$28879 ( \29223 , \29216 , \29221 );
or \U$28880 ( \29224 , \29219 , \29222 , \29223 );
and \U$28881 ( \29225 , \29214 , \29224 );
xor \U$28882 ( \29226 , \28772 , \28776 );
xor \U$28883 ( \29227 , \29226 , \28781 );
xor \U$28884 ( \29228 , \28788 , \28792 );
xor \U$28885 ( \29229 , \29228 , \28797 );
and \U$28886 ( \29230 , \29227 , \29229 );
xor \U$28887 ( \29231 , \28805 , \28809 );
xor \U$28888 ( \29232 , \29231 , \28814 );
and \U$28889 ( \29233 , \29229 , \29232 );
and \U$28890 ( \29234 , \29227 , \29232 );
or \U$28891 ( \29235 , \29230 , \29233 , \29234 );
and \U$28892 ( \29236 , \29224 , \29235 );
and \U$28893 ( \29237 , \29214 , \29235 );
or \U$28894 ( \29238 , \29225 , \29236 , \29237 );
and \U$28895 ( \29239 , \29197 , \29238 );
xor \U$28896 ( \29240 , \28824 , \28828 );
xor \U$28897 ( \29241 , \29240 , \28833 );
xor \U$28898 ( \29242 , \28842 , \28846 );
xor \U$28899 ( \29243 , \29242 , \28851 );
and \U$28900 ( \29244 , \29241 , \29243 );
xor \U$28901 ( \29245 , \28859 , \28863 );
xor \U$28902 ( \29246 , \29245 , \28868 );
and \U$28903 ( \29247 , \29243 , \29246 );
and \U$28904 ( \29248 , \29241 , \29246 );
or \U$28905 ( \29249 , \29244 , \29247 , \29248 );
xor \U$28906 ( \29250 , \28559 , \28563 );
xor \U$28907 ( \29251 , \29250 , \28568 );
and \U$28908 ( \29252 , \29249 , \29251 );
xor \U$28909 ( \29253 , \28595 , \28599 );
xor \U$28910 ( \29254 , \29253 , \28604 );
and \U$28911 ( \29255 , \29251 , \29254 );
and \U$28912 ( \29256 , \29249 , \29254 );
or \U$28913 ( \29257 , \29252 , \29255 , \29256 );
and \U$28914 ( \29258 , \29238 , \29257 );
and \U$28915 ( \29259 , \29197 , \29257 );
or \U$28916 ( \29260 , \29239 , \29258 , \29259 );
xor \U$28917 ( \29261 , \28784 , \28800 );
xor \U$28918 ( \29262 , \29261 , \28817 );
xor \U$28919 ( \29263 , \28836 , \28854 );
xor \U$28920 ( \29264 , \29263 , \28871 );
and \U$28921 ( \29265 , \29262 , \29264 );
xor \U$28922 ( \29266 , \28891 , \28907 );
xor \U$28923 ( \29267 , \29266 , \28924 );
and \U$28924 ( \29268 , \29264 , \29267 );
and \U$28925 ( \29269 , \29262 , \29267 );
or \U$28926 ( \29270 , \29265 , \29268 , \29269 );
xor \U$28927 ( \29271 , \28932 , \28934 );
xor \U$28928 ( \29272 , \29271 , \28937 );
xor \U$28929 ( \29273 , \28942 , \28944 );
xor \U$28930 ( \29274 , \29273 , \28947 );
and \U$28931 ( \29275 , \29272 , \29274 );
xnor \U$28932 ( \29276 , \28953 , \28955 );
and \U$28933 ( \29277 , \29274 , \29276 );
and \U$28934 ( \29278 , \29272 , \29276 );
or \U$28935 ( \29279 , \29275 , \29277 , \29278 );
and \U$28936 ( \29280 , \29270 , \29279 );
xor \U$28937 ( \29281 , \28571 , \28587 );
xor \U$28938 ( \29282 , \29281 , \28607 );
and \U$28939 ( \29283 , \29279 , \29282 );
and \U$28940 ( \29284 , \29270 , \29282 );
or \U$28941 ( \29285 , \29280 , \29283 , \29284 );
and \U$28942 ( \29286 , \29260 , \29285 );
xor \U$28943 ( \29287 , \28940 , \28950 );
xor \U$28944 ( \29288 , \29287 , \28956 );
xor \U$28945 ( \29289 , \28986 , \28988 );
xor \U$28946 ( \29290 , \29289 , \28991 );
and \U$28947 ( \29291 , \29288 , \29290 );
xor \U$28948 ( \29292 , \28962 , \28964 );
xor \U$28949 ( \29293 , \29292 , \28967 );
and \U$28950 ( \29294 , \29290 , \29293 );
and \U$28951 ( \29295 , \29288 , \29293 );
or \U$28952 ( \29296 , \29291 , \29294 , \29295 );
and \U$28953 ( \29297 , \29285 , \29296 );
and \U$28954 ( \29298 , \29260 , \29296 );
or \U$28955 ( \29299 , \29286 , \29297 , \29298 );
xor \U$28956 ( \29300 , \28930 , \28959 );
xor \U$28957 ( \29301 , \29300 , \28970 );
xor \U$28958 ( \29302 , \28975 , \28977 );
xor \U$28959 ( \29303 , \29302 , \28980 );
and \U$28960 ( \29304 , \29301 , \29303 );
xor \U$28961 ( \29305 , \28994 , \28996 );
xor \U$28962 ( \29306 , \29305 , \28999 );
and \U$28963 ( \29307 , \29303 , \29306 );
and \U$28964 ( \29308 , \29301 , \29306 );
or \U$28965 ( \29309 , \29304 , \29307 , \29308 );
and \U$28966 ( \29310 , \29299 , \29309 );
xor \U$28967 ( \29311 , \29007 , \29009 );
xor \U$28968 ( \29312 , \29311 , \29011 );
and \U$28969 ( \29313 , \29309 , \29312 );
and \U$28970 ( \29314 , \29299 , \29312 );
or \U$28971 ( \29315 , \29310 , \29313 , \29314 );
xor \U$28972 ( \29316 , \28713 , \28730 );
xor \U$28973 ( \29317 , \29316 , \28736 );
and \U$28974 ( \29318 , \29315 , \29317 );
xor \U$28975 ( \29319 , \29005 , \29014 );
xor \U$28976 ( \29320 , \29319 , \29017 );
and \U$28977 ( \29321 , \29317 , \29320 );
and \U$28978 ( \29322 , \29315 , \29320 );
or \U$28979 ( \29323 , \29318 , \29321 , \29322 );
xor \U$28980 ( \29324 , \29020 , \29022 );
xor \U$28981 ( \29325 , \29324 , \29025 );
and \U$28982 ( \29326 , \29323 , \29325 );
and \U$28983 ( \29327 , \29034 , \29326 );
xor \U$28984 ( \29328 , \29034 , \29326 );
xor \U$28985 ( \29329 , \29323 , \29325 );
and \U$28986 ( \29330 , \21413 , \28063 );
and \U$28987 ( \29331 , \21421 , \28061 );
nor \U$28988 ( \29332 , \29330 , \29331 );
xnor \U$28989 ( \29333 , \29332 , \27803 );
and \U$28990 ( \29334 , \21428 , \27569 );
and \U$28991 ( \29335 , \21436 , \27567 );
nor \U$28992 ( \29336 , \29334 , \29335 );
xnor \U$28993 ( \29337 , \29336 , \27254 );
and \U$28994 ( \29338 , \29333 , \29337 );
and \U$28995 ( \29339 , \21444 , \27060 );
and \U$28996 ( \29340 , \21452 , \27058 );
nor \U$28997 ( \29341 , \29339 , \29340 );
xnor \U$28998 ( \29342 , \29341 , \26720 );
and \U$28999 ( \29343 , \29337 , \29342 );
and \U$29000 ( \29344 , \29333 , \29342 );
or \U$29001 ( \29345 , \29338 , \29343 , \29344 );
buf \U$29002 ( \29346 , RIbb2db58_58);
buf \U$29003 ( \29347 , RIbb2dae0_59);
and \U$29004 ( \29348 , \29346 , \29347 );
not \U$29005 ( \29349 , \29348 );
and \U$29006 ( \29350 , \28838 , \29349 );
not \U$29007 ( \29351 , \29350 );
and \U$29008 ( \29352 , \21379 , \29159 );
and \U$29009 ( \29353 , \21387 , \29157 );
nor \U$29010 ( \29354 , \29352 , \29353 );
xnor \U$29011 ( \29355 , \29354 , \28841 );
and \U$29012 ( \29356 , \29351 , \29355 );
and \U$29013 ( \29357 , \21395 , \28592 );
and \U$29014 ( \29358 , \21403 , \28590 );
nor \U$29015 ( \29359 , \29357 , \29358 );
xnor \U$29016 ( \29360 , \29359 , \28343 );
and \U$29017 ( \29361 , \29355 , \29360 );
and \U$29018 ( \29362 , \29351 , \29360 );
or \U$29019 ( \29363 , \29356 , \29361 , \29362 );
and \U$29020 ( \29364 , \29345 , \29363 );
and \U$29021 ( \29365 , \21463 , \26471 );
and \U$29022 ( \29366 , \21471 , \26469 );
nor \U$29023 ( \29367 , \29365 , \29366 );
xnor \U$29024 ( \29368 , \29367 , \26230 );
and \U$29025 ( \29369 , \21689 , \26005 );
and \U$29026 ( \29370 , \21478 , \26003 );
nor \U$29027 ( \29371 , \29369 , \29370 );
xnor \U$29028 ( \29372 , \29371 , \25817 );
and \U$29029 ( \29373 , \29368 , \29372 );
and \U$29030 ( \29374 , \21813 , \25631 );
and \U$29031 ( \29375 , \21750 , \25629 );
nor \U$29032 ( \29376 , \29374 , \29375 );
xnor \U$29033 ( \29377 , \29376 , \25399 );
and \U$29034 ( \29378 , \29372 , \29377 );
and \U$29035 ( \29379 , \29368 , \29377 );
or \U$29036 ( \29380 , \29373 , \29378 , \29379 );
and \U$29037 ( \29381 , \29363 , \29380 );
and \U$29038 ( \29382 , \29345 , \29380 );
or \U$29039 ( \29383 , \29364 , \29381 , \29382 );
and \U$29040 ( \29384 , \23491 , \23125 );
and \U$29041 ( \29385 , \23466 , \23123 );
nor \U$29042 ( \29386 , \29384 , \29385 );
xnor \U$29043 ( \29387 , \29386 , \22988 );
and \U$29044 ( \29388 , \23832 , \22919 );
and \U$29045 ( \29389 , \23665 , \22917 );
nor \U$29046 ( \29390 , \29388 , \29389 );
xnor \U$29047 ( \29391 , \29390 , \22767 );
and \U$29048 ( \29392 , \29387 , \29391 );
and \U$29049 ( \29393 , \24089 , \22651 );
and \U$29050 ( \29394 , \23970 , \22649 );
nor \U$29051 ( \29395 , \29393 , \29394 );
xnor \U$29052 ( \29396 , \29395 , \22495 );
and \U$29053 ( \29397 , \29391 , \29396 );
and \U$29054 ( \29398 , \29387 , \29396 );
or \U$29055 ( \29399 , \29392 , \29397 , \29398 );
and \U$29056 ( \29400 , \22624 , \24149 );
and \U$29057 ( \29401 , \22616 , \24147 );
nor \U$29058 ( \29402 , \29400 , \29401 );
xnor \U$29059 ( \29403 , \29402 , \23944 );
and \U$29060 ( \29404 , \22872 , \23743 );
and \U$29061 ( \29405 , \22867 , \23741 );
nor \U$29062 ( \29406 , \29404 , \29405 );
xnor \U$29063 ( \29407 , \29406 , \23594 );
and \U$29064 ( \29408 , \29403 , \29407 );
and \U$29065 ( \29409 , \23202 , \23421 );
and \U$29066 ( \29410 , \23058 , \23419 );
nor \U$29067 ( \29411 , \29409 , \29410 );
xnor \U$29068 ( \29412 , \29411 , \23279 );
and \U$29069 ( \29413 , \29407 , \29412 );
and \U$29070 ( \29414 , \29403 , \29412 );
or \U$29071 ( \29415 , \29408 , \29413 , \29414 );
and \U$29072 ( \29416 , \29399 , \29415 );
and \U$29073 ( \29417 , \22099 , \25180 );
and \U$29074 ( \29418 , \22011 , \25178 );
nor \U$29075 ( \29419 , \29417 , \29418 );
xnor \U$29076 ( \29420 , \29419 , \25037 );
and \U$29077 ( \29421 , \22209 , \24857 );
and \U$29078 ( \29422 , \22204 , \24855 );
nor \U$29079 ( \29423 , \29421 , \29422 );
xnor \U$29080 ( \29424 , \29423 , \24611 );
and \U$29081 ( \29425 , \29420 , \29424 );
and \U$29082 ( \29426 , \22440 , \24462 );
and \U$29083 ( \29427 , \22325 , \24460 );
nor \U$29084 ( \29428 , \29426 , \29427 );
xnor \U$29085 ( \29429 , \29428 , \24275 );
and \U$29086 ( \29430 , \29424 , \29429 );
and \U$29087 ( \29431 , \29420 , \29429 );
or \U$29088 ( \29432 , \29425 , \29430 , \29431 );
and \U$29089 ( \29433 , \29415 , \29432 );
and \U$29090 ( \29434 , \29399 , \29432 );
or \U$29091 ( \29435 , \29416 , \29433 , \29434 );
and \U$29092 ( \29436 , \29383 , \29435 );
and \U$29093 ( \29437 , \25604 , \21821 );
and \U$29094 ( \29438 , \25596 , \21819 );
nor \U$29095 ( \29439 , \29437 , \29438 );
xnor \U$29096 ( \29440 , \29439 , \21727 );
and \U$29097 ( \29441 , \26078 , \21652 );
and \U$29098 ( \29442 , \26073 , \21650 );
nor \U$29099 ( \29443 , \29441 , \29442 );
xnor \U$29100 ( \29444 , \29443 , \21377 );
and \U$29101 ( \29445 , \29440 , \29444 );
and \U$29102 ( \29446 , \26601 , \21385 );
and \U$29103 ( \29447 , \26342 , \21383 );
nor \U$29104 ( \29448 , \29446 , \29447 );
xnor \U$29105 ( \29449 , \29448 , \21392 );
and \U$29106 ( \29450 , \29444 , \29449 );
and \U$29107 ( \29451 , \29440 , \29449 );
or \U$29108 ( \29452 , \29445 , \29450 , \29451 );
and \U$29109 ( \29453 , \24714 , \22379 );
and \U$29110 ( \29454 , \24506 , \22377 );
nor \U$29111 ( \29455 , \29453 , \29454 );
xnor \U$29112 ( \29456 , \29455 , \22266 );
and \U$29113 ( \29457 , \24841 , \22185 );
and \U$29114 ( \29458 , \24836 , \22183 );
nor \U$29115 ( \29459 , \29457 , \29458 );
xnor \U$29116 ( \29460 , \29459 , \22049 );
and \U$29117 ( \29461 , \29456 , \29460 );
and \U$29118 ( \29462 , \25294 , \21985 );
and \U$29119 ( \29463 , \25097 , \21983 );
nor \U$29120 ( \29464 , \29462 , \29463 );
xnor \U$29121 ( \29465 , \29464 , \21907 );
and \U$29122 ( \29466 , \29460 , \29465 );
and \U$29123 ( \29467 , \29456 , \29465 );
or \U$29124 ( \29468 , \29461 , \29466 , \29467 );
and \U$29125 ( \29469 , \29452 , \29468 );
and \U$29126 ( \29470 , \26982 , \21401 );
and \U$29127 ( \29471 , \26973 , \21399 );
nor \U$29128 ( \29472 , \29470 , \29471 );
xnor \U$29129 ( \29473 , \29472 , \21408 );
and \U$29130 ( \29474 , \27527 , \21419 );
and \U$29131 ( \29475 , \27325 , \21417 );
nor \U$29132 ( \29476 , \29474 , \29475 );
xnor \U$29133 ( \29477 , \29476 , \21426 );
and \U$29134 ( \29478 , \29473 , \29477 );
and \U$29135 ( \29479 , \28002 , \21434 );
and \U$29136 ( \29480 , \27830 , \21432 );
nor \U$29137 ( \29481 , \29479 , \29480 );
xnor \U$29138 ( \29482 , \29481 , \21441 );
and \U$29139 ( \29483 , \29477 , \29482 );
and \U$29140 ( \29484 , \29473 , \29482 );
or \U$29141 ( \29485 , \29478 , \29483 , \29484 );
and \U$29142 ( \29486 , \29468 , \29485 );
and \U$29143 ( \29487 , \29452 , \29485 );
or \U$29144 ( \29488 , \29469 , \29486 , \29487 );
and \U$29145 ( \29489 , \29435 , \29488 );
and \U$29146 ( \29490 , \29383 , \29488 );
or \U$29147 ( \29491 , \29436 , \29489 , \29490 );
xor \U$29148 ( \29492 , \29038 , \29042 );
xor \U$29149 ( \29493 , \29492 , \29047 );
xor \U$29150 ( \29494 , \29143 , \29147 );
xor \U$29151 ( \29495 , \29494 , \29152 );
and \U$29152 ( \29496 , \29493 , \29495 );
xor \U$29153 ( \29497 , \29071 , \29075 );
xor \U$29154 ( \29498 , \29497 , \29080 );
and \U$29155 ( \29499 , \29495 , \29498 );
and \U$29156 ( \29500 , \29493 , \29498 );
or \U$29157 ( \29501 , \29496 , \29499 , \29500 );
xor \U$29158 ( \29502 , \29054 , \29058 );
xor \U$29159 ( \29503 , \29502 , \29063 );
xor \U$29160 ( \29504 , \29090 , \29094 );
xor \U$29161 ( \29505 , \29504 , \29099 );
and \U$29162 ( \29506 , \29503 , \29505 );
xor \U$29163 ( \29507 , \29106 , \29110 );
xor \U$29164 ( \29508 , \29507 , \29115 );
and \U$29165 ( \29509 , \29505 , \29508 );
and \U$29166 ( \29510 , \29503 , \29508 );
or \U$29167 ( \29511 , \29506 , \29509 , \29510 );
and \U$29168 ( \29512 , \29501 , \29511 );
and \U$29169 ( \29513 , \28952 , \21450 );
and \U$29170 ( \29514 , \28528 , \21448 );
nor \U$29171 ( \29515 , \29513 , \29514 );
xnor \U$29172 ( \29516 , \29515 , \21457 );
and \U$29173 ( \29517 , \29203 , \21469 );
and \U$29174 ( \29518 , \29198 , \21467 );
nor \U$29175 ( \29519 , \29517 , \29518 );
xnor \U$29176 ( \29520 , \29519 , \21476 );
and \U$29177 ( \29521 , \29516 , \29520 );
buf \U$29178 ( \29522 , RIbb33030_185);
and \U$29179 ( \29523 , \29522 , \21464 );
and \U$29180 ( \29524 , \29520 , \29523 );
and \U$29181 ( \29525 , \29516 , \29523 );
or \U$29182 ( \29526 , \29521 , \29524 , \29525 );
xor \U$29183 ( \29527 , \29123 , \29127 );
xor \U$29184 ( \29528 , \29527 , \29132 );
and \U$29185 ( \29529 , \29526 , \29528 );
xnor \U$29186 ( \29530 , \29202 , \29204 );
and \U$29187 ( \29531 , \29528 , \29530 );
and \U$29188 ( \29532 , \29526 , \29530 );
or \U$29189 ( \29533 , \29529 , \29531 , \29532 );
and \U$29190 ( \29534 , \29511 , \29533 );
and \U$29191 ( \29535 , \29501 , \29533 );
or \U$29192 ( \29536 , \29512 , \29534 , \29535 );
and \U$29193 ( \29537 , \29491 , \29536 );
xor \U$29194 ( \29538 , \29216 , \29218 );
xor \U$29195 ( \29539 , \29538 , \29221 );
xor \U$29196 ( \29540 , \29227 , \29229 );
xor \U$29197 ( \29541 , \29540 , \29232 );
and \U$29198 ( \29542 , \29539 , \29541 );
xor \U$29199 ( \29543 , \29241 , \29243 );
xor \U$29200 ( \29544 , \29543 , \29246 );
and \U$29201 ( \29545 , \29541 , \29544 );
and \U$29202 ( \29546 , \29539 , \29544 );
or \U$29203 ( \29547 , \29542 , \29545 , \29546 );
and \U$29204 ( \29548 , \29536 , \29547 );
and \U$29205 ( \29549 , \29491 , \29547 );
or \U$29206 ( \29550 , \29537 , \29548 , \29549 );
xor \U$29207 ( \29551 , \29086 , \29138 );
xor \U$29208 ( \29552 , \29551 , \29194 );
xor \U$29209 ( \29553 , \29214 , \29224 );
xor \U$29210 ( \29554 , \29553 , \29235 );
and \U$29211 ( \29555 , \29552 , \29554 );
xor \U$29212 ( \29556 , \29249 , \29251 );
xor \U$29213 ( \29557 , \29556 , \29254 );
and \U$29214 ( \29558 , \29554 , \29557 );
and \U$29215 ( \29559 , \29552 , \29557 );
or \U$29216 ( \29560 , \29555 , \29558 , \29559 );
and \U$29217 ( \29561 , \29550 , \29560 );
xor \U$29218 ( \29562 , \29050 , \29066 );
xor \U$29219 ( \29563 , \29562 , \29083 );
xor \U$29220 ( \29564 , \29102 , \29118 );
xor \U$29221 ( \29565 , \29564 , \29135 );
and \U$29222 ( \29566 , \29563 , \29565 );
xor \U$29223 ( \29567 , \29205 , \29209 );
xor \U$29224 ( \29568 , \29567 , \29211 );
and \U$29225 ( \29569 , \29565 , \29568 );
and \U$29226 ( \29570 , \29563 , \29568 );
or \U$29227 ( \29571 , \29566 , \29569 , \29570 );
xor \U$29228 ( \29572 , \29262 , \29264 );
xor \U$29229 ( \29573 , \29572 , \29267 );
and \U$29230 ( \29574 , \29571 , \29573 );
xor \U$29231 ( \29575 , \29272 , \29274 );
xor \U$29232 ( \29576 , \29575 , \29276 );
and \U$29233 ( \29577 , \29573 , \29576 );
and \U$29234 ( \29578 , \29571 , \29576 );
or \U$29235 ( \29579 , \29574 , \29577 , \29578 );
and \U$29236 ( \29580 , \29560 , \29579 );
and \U$29237 ( \29581 , \29550 , \29579 );
or \U$29238 ( \29582 , \29561 , \29580 , \29581 );
xor \U$29239 ( \29583 , \28820 , \28874 );
xor \U$29240 ( \29584 , \29583 , \28927 );
xor \U$29241 ( \29585 , \29270 , \29279 );
xor \U$29242 ( \29586 , \29585 , \29282 );
and \U$29243 ( \29587 , \29584 , \29586 );
xor \U$29244 ( \29588 , \29288 , \29290 );
xor \U$29245 ( \29589 , \29588 , \29293 );
and \U$29246 ( \29590 , \29586 , \29589 );
and \U$29247 ( \29591 , \29584 , \29589 );
or \U$29248 ( \29592 , \29587 , \29590 , \29591 );
and \U$29249 ( \29593 , \29582 , \29592 );
xor \U$29250 ( \29594 , \29301 , \29303 );
xor \U$29251 ( \29595 , \29594 , \29306 );
and \U$29252 ( \29596 , \29592 , \29595 );
and \U$29253 ( \29597 , \29582 , \29595 );
or \U$29254 ( \29598 , \29593 , \29596 , \29597 );
xor \U$29255 ( \29599 , \28973 , \28983 );
xor \U$29256 ( \29600 , \29599 , \29002 );
and \U$29257 ( \29601 , \29598 , \29600 );
xor \U$29258 ( \29602 , \29299 , \29309 );
xor \U$29259 ( \29603 , \29602 , \29312 );
and \U$29260 ( \29604 , \29600 , \29603 );
and \U$29261 ( \29605 , \29598 , \29603 );
or \U$29262 ( \29606 , \29601 , \29604 , \29605 );
xor \U$29263 ( \29607 , \29315 , \29317 );
xor \U$29264 ( \29608 , \29607 , \29320 );
and \U$29265 ( \29609 , \29606 , \29608 );
and \U$29266 ( \29610 , \29329 , \29609 );
xor \U$29267 ( \29611 , \29329 , \29609 );
xor \U$29268 ( \29612 , \29606 , \29608 );
and \U$29269 ( \29613 , \23665 , \23125 );
and \U$29270 ( \29614 , \23491 , \23123 );
nor \U$29271 ( \29615 , \29613 , \29614 );
xnor \U$29272 ( \29616 , \29615 , \22988 );
and \U$29273 ( \29617 , \23970 , \22919 );
and \U$29274 ( \29618 , \23832 , \22917 );
nor \U$29275 ( \29619 , \29617 , \29618 );
xnor \U$29276 ( \29620 , \29619 , \22767 );
and \U$29277 ( \29621 , \29616 , \29620 );
and \U$29278 ( \29622 , \24506 , \22651 );
and \U$29279 ( \29623 , \24089 , \22649 );
nor \U$29280 ( \29624 , \29622 , \29623 );
xnor \U$29281 ( \29625 , \29624 , \22495 );
and \U$29282 ( \29626 , \29620 , \29625 );
and \U$29283 ( \29627 , \29616 , \29625 );
or \U$29284 ( \29628 , \29621 , \29626 , \29627 );
and \U$29285 ( \29629 , \22204 , \25180 );
and \U$29286 ( \29630 , \22099 , \25178 );
nor \U$29287 ( \29631 , \29629 , \29630 );
xnor \U$29288 ( \29632 , \29631 , \25037 );
and \U$29289 ( \29633 , \22325 , \24857 );
and \U$29290 ( \29634 , \22209 , \24855 );
nor \U$29291 ( \29635 , \29633 , \29634 );
xnor \U$29292 ( \29636 , \29635 , \24611 );
and \U$29293 ( \29637 , \29632 , \29636 );
and \U$29294 ( \29638 , \22616 , \24462 );
and \U$29295 ( \29639 , \22440 , \24460 );
nor \U$29296 ( \29640 , \29638 , \29639 );
xnor \U$29297 ( \29641 , \29640 , \24275 );
and \U$29298 ( \29642 , \29636 , \29641 );
and \U$29299 ( \29643 , \29632 , \29641 );
or \U$29300 ( \29644 , \29637 , \29642 , \29643 );
and \U$29301 ( \29645 , \29628 , \29644 );
and \U$29302 ( \29646 , \22867 , \24149 );
and \U$29303 ( \29647 , \22624 , \24147 );
nor \U$29304 ( \29648 , \29646 , \29647 );
xnor \U$29305 ( \29649 , \29648 , \23944 );
and \U$29306 ( \29650 , \23058 , \23743 );
and \U$29307 ( \29651 , \22872 , \23741 );
nor \U$29308 ( \29652 , \29650 , \29651 );
xnor \U$29309 ( \29653 , \29652 , \23594 );
and \U$29310 ( \29654 , \29649 , \29653 );
and \U$29311 ( \29655 , \23466 , \23421 );
and \U$29312 ( \29656 , \23202 , \23419 );
nor \U$29313 ( \29657 , \29655 , \29656 );
xnor \U$29314 ( \29658 , \29657 , \23279 );
and \U$29315 ( \29659 , \29653 , \29658 );
and \U$29316 ( \29660 , \29649 , \29658 );
or \U$29317 ( \29661 , \29654 , \29659 , \29660 );
and \U$29318 ( \29662 , \29644 , \29661 );
and \U$29319 ( \29663 , \29628 , \29661 );
or \U$29320 ( \29664 , \29645 , \29662 , \29663 );
and \U$29321 ( \29665 , \27325 , \21401 );
and \U$29322 ( \29666 , \26982 , \21399 );
nor \U$29323 ( \29667 , \29665 , \29666 );
xnor \U$29324 ( \29668 , \29667 , \21408 );
and \U$29325 ( \29669 , \27830 , \21419 );
and \U$29326 ( \29670 , \27527 , \21417 );
nor \U$29327 ( \29671 , \29669 , \29670 );
xnor \U$29328 ( \29672 , \29671 , \21426 );
and \U$29329 ( \29673 , \29668 , \29672 );
and \U$29330 ( \29674 , \28528 , \21434 );
and \U$29331 ( \29675 , \28002 , \21432 );
nor \U$29332 ( \29676 , \29674 , \29675 );
xnor \U$29333 ( \29677 , \29676 , \21441 );
and \U$29334 ( \29678 , \29672 , \29677 );
and \U$29335 ( \29679 , \29668 , \29677 );
or \U$29336 ( \29680 , \29673 , \29678 , \29679 );
and \U$29337 ( \29681 , \26073 , \21821 );
and \U$29338 ( \29682 , \25604 , \21819 );
nor \U$29339 ( \29683 , \29681 , \29682 );
xnor \U$29340 ( \29684 , \29683 , \21727 );
and \U$29341 ( \29685 , \26342 , \21652 );
and \U$29342 ( \29686 , \26078 , \21650 );
nor \U$29343 ( \29687 , \29685 , \29686 );
xnor \U$29344 ( \29688 , \29687 , \21377 );
and \U$29345 ( \29689 , \29684 , \29688 );
and \U$29346 ( \29690 , \26973 , \21385 );
and \U$29347 ( \29691 , \26601 , \21383 );
nor \U$29348 ( \29692 , \29690 , \29691 );
xnor \U$29349 ( \29693 , \29692 , \21392 );
and \U$29350 ( \29694 , \29688 , \29693 );
and \U$29351 ( \29695 , \29684 , \29693 );
or \U$29352 ( \29696 , \29689 , \29694 , \29695 );
and \U$29353 ( \29697 , \29680 , \29696 );
and \U$29354 ( \29698 , \24836 , \22379 );
and \U$29355 ( \29699 , \24714 , \22377 );
nor \U$29356 ( \29700 , \29698 , \29699 );
xnor \U$29357 ( \29701 , \29700 , \22266 );
and \U$29358 ( \29702 , \25097 , \22185 );
and \U$29359 ( \29703 , \24841 , \22183 );
nor \U$29360 ( \29704 , \29702 , \29703 );
xnor \U$29361 ( \29705 , \29704 , \22049 );
and \U$29362 ( \29706 , \29701 , \29705 );
and \U$29363 ( \29707 , \25596 , \21985 );
and \U$29364 ( \29708 , \25294 , \21983 );
nor \U$29365 ( \29709 , \29707 , \29708 );
xnor \U$29366 ( \29710 , \29709 , \21907 );
and \U$29367 ( \29711 , \29705 , \29710 );
and \U$29368 ( \29712 , \29701 , \29710 );
or \U$29369 ( \29713 , \29706 , \29711 , \29712 );
and \U$29370 ( \29714 , \29696 , \29713 );
and \U$29371 ( \29715 , \29680 , \29713 );
or \U$29372 ( \29716 , \29697 , \29714 , \29715 );
and \U$29373 ( \29717 , \29664 , \29716 );
xor \U$29374 ( \29718 , \28838 , \29346 );
xor \U$29375 ( \29719 , \29346 , \29347 );
not \U$29376 ( \29720 , \29719 );
and \U$29377 ( \29721 , \29718 , \29720 );
and \U$29378 ( \29722 , \21387 , \29721 );
not \U$29379 ( \29723 , \29722 );
xnor \U$29380 ( \29724 , \29723 , \29350 );
and \U$29381 ( \29725 , \21403 , \29159 );
and \U$29382 ( \29726 , \21379 , \29157 );
nor \U$29383 ( \29727 , \29725 , \29726 );
xnor \U$29384 ( \29728 , \29727 , \28841 );
and \U$29385 ( \29729 , \29724 , \29728 );
and \U$29386 ( \29730 , \21421 , \28592 );
and \U$29387 ( \29731 , \21395 , \28590 );
nor \U$29388 ( \29732 , \29730 , \29731 );
xnor \U$29389 ( \29733 , \29732 , \28343 );
and \U$29390 ( \29734 , \29728 , \29733 );
and \U$29391 ( \29735 , \29724 , \29733 );
or \U$29392 ( \29736 , \29729 , \29734 , \29735 );
and \U$29393 ( \29737 , \21478 , \26471 );
and \U$29394 ( \29738 , \21463 , \26469 );
nor \U$29395 ( \29739 , \29737 , \29738 );
xnor \U$29396 ( \29740 , \29739 , \26230 );
and \U$29397 ( \29741 , \21750 , \26005 );
and \U$29398 ( \29742 , \21689 , \26003 );
nor \U$29399 ( \29743 , \29741 , \29742 );
xnor \U$29400 ( \29744 , \29743 , \25817 );
and \U$29401 ( \29745 , \29740 , \29744 );
and \U$29402 ( \29746 , \22011 , \25631 );
and \U$29403 ( \29747 , \21813 , \25629 );
nor \U$29404 ( \29748 , \29746 , \29747 );
xnor \U$29405 ( \29749 , \29748 , \25399 );
and \U$29406 ( \29750 , \29744 , \29749 );
and \U$29407 ( \29751 , \29740 , \29749 );
or \U$29408 ( \29752 , \29745 , \29750 , \29751 );
and \U$29409 ( \29753 , \29736 , \29752 );
and \U$29410 ( \29754 , \21436 , \28063 );
and \U$29411 ( \29755 , \21413 , \28061 );
nor \U$29412 ( \29756 , \29754 , \29755 );
xnor \U$29413 ( \29757 , \29756 , \27803 );
and \U$29414 ( \29758 , \21452 , \27569 );
and \U$29415 ( \29759 , \21428 , \27567 );
nor \U$29416 ( \29760 , \29758 , \29759 );
xnor \U$29417 ( \29761 , \29760 , \27254 );
and \U$29418 ( \29762 , \29757 , \29761 );
and \U$29419 ( \29763 , \21471 , \27060 );
and \U$29420 ( \29764 , \21444 , \27058 );
nor \U$29421 ( \29765 , \29763 , \29764 );
xnor \U$29422 ( \29766 , \29765 , \26720 );
and \U$29423 ( \29767 , \29761 , \29766 );
and \U$29424 ( \29768 , \29757 , \29766 );
or \U$29425 ( \29769 , \29762 , \29767 , \29768 );
and \U$29426 ( \29770 , \29752 , \29769 );
and \U$29427 ( \29771 , \29736 , \29769 );
or \U$29428 ( \29772 , \29753 , \29770 , \29771 );
and \U$29429 ( \29773 , \29716 , \29772 );
and \U$29430 ( \29774 , \29664 , \29772 );
or \U$29431 ( \29775 , \29717 , \29773 , \29774 );
xor \U$29432 ( \29776 , \29368 , \29372 );
xor \U$29433 ( \29777 , \29776 , \29377 );
xor \U$29434 ( \29778 , \29403 , \29407 );
xor \U$29435 ( \29779 , \29778 , \29412 );
and \U$29436 ( \29780 , \29777 , \29779 );
xor \U$29437 ( \29781 , \29420 , \29424 );
xor \U$29438 ( \29782 , \29781 , \29429 );
and \U$29439 ( \29783 , \29779 , \29782 );
and \U$29440 ( \29784 , \29777 , \29782 );
or \U$29441 ( \29785 , \29780 , \29783 , \29784 );
xor \U$29442 ( \29786 , \29387 , \29391 );
xor \U$29443 ( \29787 , \29786 , \29396 );
xor \U$29444 ( \29788 , \29440 , \29444 );
xor \U$29445 ( \29789 , \29788 , \29449 );
and \U$29446 ( \29790 , \29787 , \29789 );
xor \U$29447 ( \29791 , \29456 , \29460 );
xor \U$29448 ( \29792 , \29791 , \29465 );
and \U$29449 ( \29793 , \29789 , \29792 );
and \U$29450 ( \29794 , \29787 , \29792 );
or \U$29451 ( \29795 , \29790 , \29793 , \29794 );
and \U$29452 ( \29796 , \29785 , \29795 );
and \U$29453 ( \29797 , \29198 , \21450 );
and \U$29454 ( \29798 , \28952 , \21448 );
nor \U$29455 ( \29799 , \29797 , \29798 );
xnor \U$29456 ( \29800 , \29799 , \21457 );
and \U$29457 ( \29801 , \29522 , \21469 );
and \U$29458 ( \29802 , \29203 , \21467 );
nor \U$29459 ( \29803 , \29801 , \29802 );
xnor \U$29460 ( \29804 , \29803 , \21476 );
and \U$29461 ( \29805 , \29800 , \29804 );
buf \U$29462 ( \29806 , RIbb330a8_186);
and \U$29463 ( \29807 , \29806 , \21464 );
and \U$29464 ( \29808 , \29804 , \29807 );
and \U$29465 ( \29809 , \29800 , \29807 );
or \U$29466 ( \29810 , \29805 , \29808 , \29809 );
xor \U$29467 ( \29811 , \29516 , \29520 );
xor \U$29468 ( \29812 , \29811 , \29523 );
and \U$29469 ( \29813 , \29810 , \29812 );
xor \U$29470 ( \29814 , \29473 , \29477 );
xor \U$29471 ( \29815 , \29814 , \29482 );
and \U$29472 ( \29816 , \29812 , \29815 );
and \U$29473 ( \29817 , \29810 , \29815 );
or \U$29474 ( \29818 , \29813 , \29816 , \29817 );
and \U$29475 ( \29819 , \29795 , \29818 );
and \U$29476 ( \29820 , \29785 , \29818 );
or \U$29477 ( \29821 , \29796 , \29819 , \29820 );
and \U$29478 ( \29822 , \29775 , \29821 );
xor \U$29479 ( \29823 , \29162 , \29166 );
xor \U$29480 ( \29824 , \29823 , \29171 );
xor \U$29481 ( \29825 , \29179 , \29183 );
xor \U$29482 ( \29826 , \29825 , \29188 );
and \U$29483 ( \29827 , \29824 , \29826 );
xor \U$29484 ( \29828 , \29493 , \29495 );
xor \U$29485 ( \29829 , \29828 , \29498 );
and \U$29486 ( \29830 , \29826 , \29829 );
and \U$29487 ( \29831 , \29824 , \29829 );
or \U$29488 ( \29832 , \29827 , \29830 , \29831 );
and \U$29489 ( \29833 , \29821 , \29832 );
and \U$29490 ( \29834 , \29775 , \29832 );
or \U$29491 ( \29835 , \29822 , \29833 , \29834 );
xor \U$29492 ( \29836 , \29452 , \29468 );
xor \U$29493 ( \29837 , \29836 , \29485 );
xor \U$29494 ( \29838 , \29503 , \29505 );
xor \U$29495 ( \29839 , \29838 , \29508 );
and \U$29496 ( \29840 , \29837 , \29839 );
xor \U$29497 ( \29841 , \29526 , \29528 );
xor \U$29498 ( \29842 , \29841 , \29530 );
and \U$29499 ( \29843 , \29839 , \29842 );
and \U$29500 ( \29844 , \29837 , \29842 );
or \U$29501 ( \29845 , \29840 , \29843 , \29844 );
xor \U$29502 ( \29846 , \29155 , \29174 );
xor \U$29503 ( \29847 , \29846 , \29191 );
and \U$29504 ( \29848 , \29845 , \29847 );
xor \U$29505 ( \29849 , \29563 , \29565 );
xor \U$29506 ( \29850 , \29849 , \29568 );
and \U$29507 ( \29851 , \29847 , \29850 );
and \U$29508 ( \29852 , \29845 , \29850 );
or \U$29509 ( \29853 , \29848 , \29851 , \29852 );
and \U$29510 ( \29854 , \29835 , \29853 );
xor \U$29511 ( \29855 , \29383 , \29435 );
xor \U$29512 ( \29856 , \29855 , \29488 );
xor \U$29513 ( \29857 , \29501 , \29511 );
xor \U$29514 ( \29858 , \29857 , \29533 );
and \U$29515 ( \29859 , \29856 , \29858 );
xor \U$29516 ( \29860 , \29539 , \29541 );
xor \U$29517 ( \29861 , \29860 , \29544 );
and \U$29518 ( \29862 , \29858 , \29861 );
and \U$29519 ( \29863 , \29856 , \29861 );
or \U$29520 ( \29864 , \29859 , \29862 , \29863 );
and \U$29521 ( \29865 , \29853 , \29864 );
and \U$29522 ( \29866 , \29835 , \29864 );
or \U$29523 ( \29867 , \29854 , \29865 , \29866 );
xor \U$29524 ( \29868 , \29491 , \29536 );
xor \U$29525 ( \29869 , \29868 , \29547 );
xor \U$29526 ( \29870 , \29552 , \29554 );
xor \U$29527 ( \29871 , \29870 , \29557 );
and \U$29528 ( \29872 , \29869 , \29871 );
xor \U$29529 ( \29873 , \29571 , \29573 );
xor \U$29530 ( \29874 , \29873 , \29576 );
and \U$29531 ( \29875 , \29871 , \29874 );
and \U$29532 ( \29876 , \29869 , \29874 );
or \U$29533 ( \29877 , \29872 , \29875 , \29876 );
and \U$29534 ( \29878 , \29867 , \29877 );
xor \U$29535 ( \29879 , \29197 , \29238 );
xor \U$29536 ( \29880 , \29879 , \29257 );
and \U$29537 ( \29881 , \29877 , \29880 );
and \U$29538 ( \29882 , \29867 , \29880 );
or \U$29539 ( \29883 , \29878 , \29881 , \29882 );
xor \U$29540 ( \29884 , \29550 , \29560 );
xor \U$29541 ( \29885 , \29884 , \29579 );
xor \U$29542 ( \29886 , \29584 , \29586 );
xor \U$29543 ( \29887 , \29886 , \29589 );
and \U$29544 ( \29888 , \29885 , \29887 );
and \U$29545 ( \29889 , \29883 , \29888 );
xor \U$29546 ( \29890 , \29260 , \29285 );
xor \U$29547 ( \29891 , \29890 , \29296 );
and \U$29548 ( \29892 , \29888 , \29891 );
and \U$29549 ( \29893 , \29883 , \29891 );
or \U$29550 ( \29894 , \29889 , \29892 , \29893 );
xor \U$29551 ( \29895 , \29598 , \29600 );
xor \U$29552 ( \29896 , \29895 , \29603 );
and \U$29553 ( \29897 , \29894 , \29896 );
and \U$29554 ( \29898 , \29612 , \29897 );
xor \U$29555 ( \29899 , \29612 , \29897 );
xor \U$29556 ( \29900 , \29894 , \29896 );
xor \U$29557 ( \29901 , \29668 , \29672 );
xor \U$29558 ( \29902 , \29901 , \29677 );
xor \U$29559 ( \29903 , \29684 , \29688 );
xor \U$29560 ( \29904 , \29903 , \29693 );
and \U$29561 ( \29905 , \29902 , \29904 );
xor \U$29562 ( \29906 , \29701 , \29705 );
xor \U$29563 ( \29907 , \29906 , \29710 );
and \U$29564 ( \29908 , \29904 , \29907 );
and \U$29565 ( \29909 , \29902 , \29907 );
or \U$29566 ( \29910 , \29905 , \29908 , \29909 );
xor \U$29567 ( \29911 , \29616 , \29620 );
xor \U$29568 ( \29912 , \29911 , \29625 );
xor \U$29569 ( \29913 , \29632 , \29636 );
xor \U$29570 ( \29914 , \29913 , \29641 );
and \U$29571 ( \29915 , \29912 , \29914 );
xor \U$29572 ( \29916 , \29649 , \29653 );
xor \U$29573 ( \29917 , \29916 , \29658 );
and \U$29574 ( \29918 , \29914 , \29917 );
and \U$29575 ( \29919 , \29912 , \29917 );
or \U$29576 ( \29920 , \29915 , \29918 , \29919 );
and \U$29577 ( \29921 , \29910 , \29920 );
and \U$29578 ( \29922 , \28952 , \21434 );
and \U$29579 ( \29923 , \28528 , \21432 );
nor \U$29580 ( \29924 , \29922 , \29923 );
xnor \U$29581 ( \29925 , \29924 , \21441 );
and \U$29582 ( \29926 , \29203 , \21450 );
and \U$29583 ( \29927 , \29198 , \21448 );
nor \U$29584 ( \29928 , \29926 , \29927 );
xnor \U$29585 ( \29929 , \29928 , \21457 );
and \U$29586 ( \29930 , \29925 , \29929 );
and \U$29587 ( \29931 , \29806 , \21469 );
and \U$29588 ( \29932 , \29522 , \21467 );
nor \U$29589 ( \29933 , \29931 , \29932 );
xnor \U$29590 ( \29934 , \29933 , \21476 );
and \U$29591 ( \29935 , \29929 , \29934 );
and \U$29592 ( \29936 , \29925 , \29934 );
or \U$29593 ( \29937 , \29930 , \29935 , \29936 );
xor \U$29594 ( \29938 , \29800 , \29804 );
xor \U$29595 ( \29939 , \29938 , \29807 );
or \U$29596 ( \29940 , \29937 , \29939 );
and \U$29597 ( \29941 , \29920 , \29940 );
and \U$29598 ( \29942 , \29910 , \29940 );
or \U$29599 ( \29943 , \29921 , \29941 , \29942 );
buf \U$29600 ( \29944 , RIbb2da68_60);
buf \U$29601 ( \29945 , RIbb2d9f0_61);
and \U$29602 ( \29946 , \29944 , \29945 );
not \U$29603 ( \29947 , \29946 );
and \U$29604 ( \29948 , \29347 , \29947 );
not \U$29605 ( \29949 , \29948 );
and \U$29606 ( \29950 , \21379 , \29721 );
and \U$29607 ( \29951 , \21387 , \29719 );
nor \U$29608 ( \29952 , \29950 , \29951 );
xnor \U$29609 ( \29953 , \29952 , \29350 );
and \U$29610 ( \29954 , \29949 , \29953 );
and \U$29611 ( \29955 , \21395 , \29159 );
and \U$29612 ( \29956 , \21403 , \29157 );
nor \U$29613 ( \29957 , \29955 , \29956 );
xnor \U$29614 ( \29958 , \29957 , \28841 );
and \U$29615 ( \29959 , \29953 , \29958 );
and \U$29616 ( \29960 , \29949 , \29958 );
or \U$29617 ( \29961 , \29954 , \29959 , \29960 );
and \U$29618 ( \29962 , \21463 , \27060 );
and \U$29619 ( \29963 , \21471 , \27058 );
nor \U$29620 ( \29964 , \29962 , \29963 );
xnor \U$29621 ( \29965 , \29964 , \26720 );
and \U$29622 ( \29966 , \21689 , \26471 );
and \U$29623 ( \29967 , \21478 , \26469 );
nor \U$29624 ( \29968 , \29966 , \29967 );
xnor \U$29625 ( \29969 , \29968 , \26230 );
and \U$29626 ( \29970 , \29965 , \29969 );
and \U$29627 ( \29971 , \21813 , \26005 );
and \U$29628 ( \29972 , \21750 , \26003 );
nor \U$29629 ( \29973 , \29971 , \29972 );
xnor \U$29630 ( \29974 , \29973 , \25817 );
and \U$29631 ( \29975 , \29969 , \29974 );
and \U$29632 ( \29976 , \29965 , \29974 );
or \U$29633 ( \29977 , \29970 , \29975 , \29976 );
and \U$29634 ( \29978 , \29961 , \29977 );
and \U$29635 ( \29979 , \21413 , \28592 );
and \U$29636 ( \29980 , \21421 , \28590 );
nor \U$29637 ( \29981 , \29979 , \29980 );
xnor \U$29638 ( \29982 , \29981 , \28343 );
and \U$29639 ( \29983 , \21428 , \28063 );
and \U$29640 ( \29984 , \21436 , \28061 );
nor \U$29641 ( \29985 , \29983 , \29984 );
xnor \U$29642 ( \29986 , \29985 , \27803 );
and \U$29643 ( \29987 , \29982 , \29986 );
and \U$29644 ( \29988 , \21444 , \27569 );
and \U$29645 ( \29989 , \21452 , \27567 );
nor \U$29646 ( \29990 , \29988 , \29989 );
xnor \U$29647 ( \29991 , \29990 , \27254 );
and \U$29648 ( \29992 , \29986 , \29991 );
and \U$29649 ( \29993 , \29982 , \29991 );
or \U$29650 ( \29994 , \29987 , \29992 , \29993 );
and \U$29651 ( \29995 , \29977 , \29994 );
and \U$29652 ( \29996 , \29961 , \29994 );
or \U$29653 ( \29997 , \29978 , \29995 , \29996 );
and \U$29654 ( \29998 , \22624 , \24462 );
and \U$29655 ( \29999 , \22616 , \24460 );
nor \U$29656 ( \30000 , \29998 , \29999 );
xnor \U$29657 ( \30001 , \30000 , \24275 );
and \U$29658 ( \30002 , \22872 , \24149 );
and \U$29659 ( \30003 , \22867 , \24147 );
nor \U$29660 ( \30004 , \30002 , \30003 );
xnor \U$29661 ( \30005 , \30004 , \23944 );
and \U$29662 ( \30006 , \30001 , \30005 );
and \U$29663 ( \30007 , \23202 , \23743 );
and \U$29664 ( \30008 , \23058 , \23741 );
nor \U$29665 ( \30009 , \30007 , \30008 );
xnor \U$29666 ( \30010 , \30009 , \23594 );
and \U$29667 ( \30011 , \30005 , \30010 );
and \U$29668 ( \30012 , \30001 , \30010 );
or \U$29669 ( \30013 , \30006 , \30011 , \30012 );
and \U$29670 ( \30014 , \23491 , \23421 );
and \U$29671 ( \30015 , \23466 , \23419 );
nor \U$29672 ( \30016 , \30014 , \30015 );
xnor \U$29673 ( \30017 , \30016 , \23279 );
and \U$29674 ( \30018 , \23832 , \23125 );
and \U$29675 ( \30019 , \23665 , \23123 );
nor \U$29676 ( \30020 , \30018 , \30019 );
xnor \U$29677 ( \30021 , \30020 , \22988 );
and \U$29678 ( \30022 , \30017 , \30021 );
and \U$29679 ( \30023 , \24089 , \22919 );
and \U$29680 ( \30024 , \23970 , \22917 );
nor \U$29681 ( \30025 , \30023 , \30024 );
xnor \U$29682 ( \30026 , \30025 , \22767 );
and \U$29683 ( \30027 , \30021 , \30026 );
and \U$29684 ( \30028 , \30017 , \30026 );
or \U$29685 ( \30029 , \30022 , \30027 , \30028 );
and \U$29686 ( \30030 , \30013 , \30029 );
and \U$29687 ( \30031 , \22099 , \25631 );
and \U$29688 ( \30032 , \22011 , \25629 );
nor \U$29689 ( \30033 , \30031 , \30032 );
xnor \U$29690 ( \30034 , \30033 , \25399 );
and \U$29691 ( \30035 , \22209 , \25180 );
and \U$29692 ( \30036 , \22204 , \25178 );
nor \U$29693 ( \30037 , \30035 , \30036 );
xnor \U$29694 ( \30038 , \30037 , \25037 );
and \U$29695 ( \30039 , \30034 , \30038 );
and \U$29696 ( \30040 , \22440 , \24857 );
and \U$29697 ( \30041 , \22325 , \24855 );
nor \U$29698 ( \30042 , \30040 , \30041 );
xnor \U$29699 ( \30043 , \30042 , \24611 );
and \U$29700 ( \30044 , \30038 , \30043 );
and \U$29701 ( \30045 , \30034 , \30043 );
or \U$29702 ( \30046 , \30039 , \30044 , \30045 );
and \U$29703 ( \30047 , \30029 , \30046 );
and \U$29704 ( \30048 , \30013 , \30046 );
or \U$29705 ( \30049 , \30030 , \30047 , \30048 );
and \U$29706 ( \30050 , \29997 , \30049 );
and \U$29707 ( \30051 , \26982 , \21385 );
and \U$29708 ( \30052 , \26973 , \21383 );
nor \U$29709 ( \30053 , \30051 , \30052 );
xnor \U$29710 ( \30054 , \30053 , \21392 );
and \U$29711 ( \30055 , \27527 , \21401 );
and \U$29712 ( \30056 , \27325 , \21399 );
nor \U$29713 ( \30057 , \30055 , \30056 );
xnor \U$29714 ( \30058 , \30057 , \21408 );
and \U$29715 ( \30059 , \30054 , \30058 );
and \U$29716 ( \30060 , \28002 , \21419 );
and \U$29717 ( \30061 , \27830 , \21417 );
nor \U$29718 ( \30062 , \30060 , \30061 );
xnor \U$29719 ( \30063 , \30062 , \21426 );
and \U$29720 ( \30064 , \30058 , \30063 );
and \U$29721 ( \30065 , \30054 , \30063 );
or \U$29722 ( \30066 , \30059 , \30064 , \30065 );
and \U$29723 ( \30067 , \25604 , \21985 );
and \U$29724 ( \30068 , \25596 , \21983 );
nor \U$29725 ( \30069 , \30067 , \30068 );
xnor \U$29726 ( \30070 , \30069 , \21907 );
and \U$29727 ( \30071 , \26078 , \21821 );
and \U$29728 ( \30072 , \26073 , \21819 );
nor \U$29729 ( \30073 , \30071 , \30072 );
xnor \U$29730 ( \30074 , \30073 , \21727 );
and \U$29731 ( \30075 , \30070 , \30074 );
and \U$29732 ( \30076 , \26601 , \21652 );
and \U$29733 ( \30077 , \26342 , \21650 );
nor \U$29734 ( \30078 , \30076 , \30077 );
xnor \U$29735 ( \30079 , \30078 , \21377 );
and \U$29736 ( \30080 , \30074 , \30079 );
and \U$29737 ( \30081 , \30070 , \30079 );
or \U$29738 ( \30082 , \30075 , \30080 , \30081 );
and \U$29739 ( \30083 , \30066 , \30082 );
and \U$29740 ( \30084 , \24714 , \22651 );
and \U$29741 ( \30085 , \24506 , \22649 );
nor \U$29742 ( \30086 , \30084 , \30085 );
xnor \U$29743 ( \30087 , \30086 , \22495 );
and \U$29744 ( \30088 , \24841 , \22379 );
and \U$29745 ( \30089 , \24836 , \22377 );
nor \U$29746 ( \30090 , \30088 , \30089 );
xnor \U$29747 ( \30091 , \30090 , \22266 );
and \U$29748 ( \30092 , \30087 , \30091 );
and \U$29749 ( \30093 , \25294 , \22185 );
and \U$29750 ( \30094 , \25097 , \22183 );
nor \U$29751 ( \30095 , \30093 , \30094 );
xnor \U$29752 ( \30096 , \30095 , \22049 );
and \U$29753 ( \30097 , \30091 , \30096 );
and \U$29754 ( \30098 , \30087 , \30096 );
or \U$29755 ( \30099 , \30092 , \30097 , \30098 );
and \U$29756 ( \30100 , \30082 , \30099 );
and \U$29757 ( \30101 , \30066 , \30099 );
or \U$29758 ( \30102 , \30083 , \30100 , \30101 );
and \U$29759 ( \30103 , \30049 , \30102 );
and \U$29760 ( \30104 , \29997 , \30102 );
or \U$29761 ( \30105 , \30050 , \30103 , \30104 );
and \U$29762 ( \30106 , \29943 , \30105 );
xor \U$29763 ( \30107 , \29724 , \29728 );
xor \U$29764 ( \30108 , \30107 , \29733 );
xor \U$29765 ( \30109 , \29740 , \29744 );
xor \U$29766 ( \30110 , \30109 , \29749 );
and \U$29767 ( \30111 , \30108 , \30110 );
xor \U$29768 ( \30112 , \29757 , \29761 );
xor \U$29769 ( \30113 , \30112 , \29766 );
and \U$29770 ( \30114 , \30110 , \30113 );
and \U$29771 ( \30115 , \30108 , \30113 );
or \U$29772 ( \30116 , \30111 , \30114 , \30115 );
xor \U$29773 ( \30117 , \29333 , \29337 );
xor \U$29774 ( \30118 , \30117 , \29342 );
and \U$29775 ( \30119 , \30116 , \30118 );
xor \U$29776 ( \30120 , \29351 , \29355 );
xor \U$29777 ( \30121 , \30120 , \29360 );
and \U$29778 ( \30122 , \30118 , \30121 );
and \U$29779 ( \30123 , \30116 , \30121 );
or \U$29780 ( \30124 , \30119 , \30122 , \30123 );
and \U$29781 ( \30125 , \30105 , \30124 );
and \U$29782 ( \30126 , \29943 , \30124 );
or \U$29783 ( \30127 , \30106 , \30125 , \30126 );
xor \U$29784 ( \30128 , \29628 , \29644 );
xor \U$29785 ( \30129 , \30128 , \29661 );
xor \U$29786 ( \30130 , \29680 , \29696 );
xor \U$29787 ( \30131 , \30130 , \29713 );
and \U$29788 ( \30132 , \30129 , \30131 );
xor \U$29789 ( \30133 , \29736 , \29752 );
xor \U$29790 ( \30134 , \30133 , \29769 );
and \U$29791 ( \30135 , \30131 , \30134 );
and \U$29792 ( \30136 , \30129 , \30134 );
or \U$29793 ( \30137 , \30132 , \30135 , \30136 );
xor \U$29794 ( \30138 , \29777 , \29779 );
xor \U$29795 ( \30139 , \30138 , \29782 );
xor \U$29796 ( \30140 , \29787 , \29789 );
xor \U$29797 ( \30141 , \30140 , \29792 );
and \U$29798 ( \30142 , \30139 , \30141 );
xor \U$29799 ( \30143 , \29810 , \29812 );
xor \U$29800 ( \30144 , \30143 , \29815 );
and \U$29801 ( \30145 , \30141 , \30144 );
and \U$29802 ( \30146 , \30139 , \30144 );
or \U$29803 ( \30147 , \30142 , \30145 , \30146 );
and \U$29804 ( \30148 , \30137 , \30147 );
xor \U$29805 ( \30149 , \29399 , \29415 );
xor \U$29806 ( \30150 , \30149 , \29432 );
and \U$29807 ( \30151 , \30147 , \30150 );
and \U$29808 ( \30152 , \30137 , \30150 );
or \U$29809 ( \30153 , \30148 , \30151 , \30152 );
and \U$29810 ( \30154 , \30127 , \30153 );
xor \U$29811 ( \30155 , \29345 , \29363 );
xor \U$29812 ( \30156 , \30155 , \29380 );
xor \U$29813 ( \30157 , \29824 , \29826 );
xor \U$29814 ( \30158 , \30157 , \29829 );
and \U$29815 ( \30159 , \30156 , \30158 );
xor \U$29816 ( \30160 , \29837 , \29839 );
xor \U$29817 ( \30161 , \30160 , \29842 );
and \U$29818 ( \30162 , \30158 , \30161 );
and \U$29819 ( \30163 , \30156 , \30161 );
or \U$29820 ( \30164 , \30159 , \30162 , \30163 );
and \U$29821 ( \30165 , \30153 , \30164 );
and \U$29822 ( \30166 , \30127 , \30164 );
or \U$29823 ( \30167 , \30154 , \30165 , \30166 );
xor \U$29824 ( \30168 , \29775 , \29821 );
xor \U$29825 ( \30169 , \30168 , \29832 );
xor \U$29826 ( \30170 , \29845 , \29847 );
xor \U$29827 ( \30171 , \30170 , \29850 );
and \U$29828 ( \30172 , \30169 , \30171 );
xor \U$29829 ( \30173 , \29856 , \29858 );
xor \U$29830 ( \30174 , \30173 , \29861 );
and \U$29831 ( \30175 , \30171 , \30174 );
and \U$29832 ( \30176 , \30169 , \30174 );
or \U$29833 ( \30177 , \30172 , \30175 , \30176 );
and \U$29834 ( \30178 , \30167 , \30177 );
xor \U$29835 ( \30179 , \29869 , \29871 );
xor \U$29836 ( \30180 , \30179 , \29874 );
and \U$29837 ( \30181 , \30177 , \30180 );
and \U$29838 ( \30182 , \30167 , \30180 );
or \U$29839 ( \30183 , \30178 , \30181 , \30182 );
xor \U$29840 ( \30184 , \29867 , \29877 );
xor \U$29841 ( \30185 , \30184 , \29880 );
and \U$29842 ( \30186 , \30183 , \30185 );
xor \U$29843 ( \30187 , \29885 , \29887 );
and \U$29844 ( \30188 , \30185 , \30187 );
and \U$29845 ( \30189 , \30183 , \30187 );
or \U$29846 ( \30190 , \30186 , \30188 , \30189 );
xor \U$29847 ( \30191 , \29883 , \29888 );
xor \U$29848 ( \30192 , \30191 , \29891 );
and \U$29849 ( \30193 , \30190 , \30192 );
xor \U$29850 ( \30194 , \29582 , \29592 );
xor \U$29851 ( \30195 , \30194 , \29595 );
and \U$29852 ( \30196 , \30192 , \30195 );
and \U$29853 ( \30197 , \30190 , \30195 );
or \U$29854 ( \30198 , \30193 , \30196 , \30197 );
and \U$29855 ( \30199 , \29900 , \30198 );
xor \U$29856 ( \30200 , \29900 , \30198 );
xor \U$29857 ( \30201 , \30190 , \30192 );
xor \U$29858 ( \30202 , \30201 , \30195 );
and \U$29859 ( \30203 , \26073 , \21985 );
and \U$29860 ( \30204 , \25604 , \21983 );
nor \U$29861 ( \30205 , \30203 , \30204 );
xnor \U$29862 ( \30206 , \30205 , \21907 );
and \U$29863 ( \30207 , \26342 , \21821 );
and \U$29864 ( \30208 , \26078 , \21819 );
nor \U$29865 ( \30209 , \30207 , \30208 );
xnor \U$29866 ( \30210 , \30209 , \21727 );
and \U$29867 ( \30211 , \30206 , \30210 );
and \U$29868 ( \30212 , \26973 , \21652 );
and \U$29869 ( \30213 , \26601 , \21650 );
nor \U$29870 ( \30214 , \30212 , \30213 );
xnor \U$29871 ( \30215 , \30214 , \21377 );
and \U$29872 ( \30216 , \30210 , \30215 );
and \U$29873 ( \30217 , \30206 , \30215 );
or \U$29874 ( \30218 , \30211 , \30216 , \30217 );
and \U$29875 ( \30219 , \24836 , \22651 );
and \U$29876 ( \30220 , \24714 , \22649 );
nor \U$29877 ( \30221 , \30219 , \30220 );
xnor \U$29878 ( \30222 , \30221 , \22495 );
and \U$29879 ( \30223 , \25097 , \22379 );
and \U$29880 ( \30224 , \24841 , \22377 );
nor \U$29881 ( \30225 , \30223 , \30224 );
xnor \U$29882 ( \30226 , \30225 , \22266 );
and \U$29883 ( \30227 , \30222 , \30226 );
and \U$29884 ( \30228 , \25596 , \22185 );
and \U$29885 ( \30229 , \25294 , \22183 );
nor \U$29886 ( \30230 , \30228 , \30229 );
xnor \U$29887 ( \30231 , \30230 , \22049 );
and \U$29888 ( \30232 , \30226 , \30231 );
and \U$29889 ( \30233 , \30222 , \30231 );
or \U$29890 ( \30234 , \30227 , \30232 , \30233 );
and \U$29891 ( \30235 , \30218 , \30234 );
and \U$29892 ( \30236 , \27325 , \21385 );
and \U$29893 ( \30237 , \26982 , \21383 );
nor \U$29894 ( \30238 , \30236 , \30237 );
xnor \U$29895 ( \30239 , \30238 , \21392 );
and \U$29896 ( \30240 , \27830 , \21401 );
and \U$29897 ( \30241 , \27527 , \21399 );
nor \U$29898 ( \30242 , \30240 , \30241 );
xnor \U$29899 ( \30243 , \30242 , \21408 );
and \U$29900 ( \30244 , \30239 , \30243 );
and \U$29901 ( \30245 , \28528 , \21419 );
and \U$29902 ( \30246 , \28002 , \21417 );
nor \U$29903 ( \30247 , \30245 , \30246 );
xnor \U$29904 ( \30248 , \30247 , \21426 );
and \U$29905 ( \30249 , \30243 , \30248 );
and \U$29906 ( \30250 , \30239 , \30248 );
or \U$29907 ( \30251 , \30244 , \30249 , \30250 );
and \U$29908 ( \30252 , \30234 , \30251 );
and \U$29909 ( \30253 , \30218 , \30251 );
or \U$29910 ( \30254 , \30235 , \30252 , \30253 );
xor \U$29911 ( \30255 , \29347 , \29944 );
xor \U$29912 ( \30256 , \29944 , \29945 );
not \U$29913 ( \30257 , \30256 );
and \U$29914 ( \30258 , \30255 , \30257 );
and \U$29915 ( \30259 , \21387 , \30258 );
not \U$29916 ( \30260 , \30259 );
xnor \U$29917 ( \30261 , \30260 , \29948 );
and \U$29918 ( \30262 , \21403 , \29721 );
and \U$29919 ( \30263 , \21379 , \29719 );
nor \U$29920 ( \30264 , \30262 , \30263 );
xnor \U$29921 ( \30265 , \30264 , \29350 );
and \U$29922 ( \30266 , \30261 , \30265 );
and \U$29923 ( \30267 , \21421 , \29159 );
and \U$29924 ( \30268 , \21395 , \29157 );
nor \U$29925 ( \30269 , \30267 , \30268 );
xnor \U$29926 ( \30270 , \30269 , \28841 );
and \U$29927 ( \30271 , \30265 , \30270 );
and \U$29928 ( \30272 , \30261 , \30270 );
or \U$29929 ( \30273 , \30266 , \30271 , \30272 );
and \U$29930 ( \30274 , \21478 , \27060 );
and \U$29931 ( \30275 , \21463 , \27058 );
nor \U$29932 ( \30276 , \30274 , \30275 );
xnor \U$29933 ( \30277 , \30276 , \26720 );
and \U$29934 ( \30278 , \21750 , \26471 );
and \U$29935 ( \30279 , \21689 , \26469 );
nor \U$29936 ( \30280 , \30278 , \30279 );
xnor \U$29937 ( \30281 , \30280 , \26230 );
and \U$29938 ( \30282 , \30277 , \30281 );
and \U$29939 ( \30283 , \22011 , \26005 );
and \U$29940 ( \30284 , \21813 , \26003 );
nor \U$29941 ( \30285 , \30283 , \30284 );
xnor \U$29942 ( \30286 , \30285 , \25817 );
and \U$29943 ( \30287 , \30281 , \30286 );
and \U$29944 ( \30288 , \30277 , \30286 );
or \U$29945 ( \30289 , \30282 , \30287 , \30288 );
and \U$29946 ( \30290 , \30273 , \30289 );
and \U$29947 ( \30291 , \21436 , \28592 );
and \U$29948 ( \30292 , \21413 , \28590 );
nor \U$29949 ( \30293 , \30291 , \30292 );
xnor \U$29950 ( \30294 , \30293 , \28343 );
and \U$29951 ( \30295 , \21452 , \28063 );
and \U$29952 ( \30296 , \21428 , \28061 );
nor \U$29953 ( \30297 , \30295 , \30296 );
xnor \U$29954 ( \30298 , \30297 , \27803 );
and \U$29955 ( \30299 , \30294 , \30298 );
and \U$29956 ( \30300 , \21471 , \27569 );
and \U$29957 ( \30301 , \21444 , \27567 );
nor \U$29958 ( \30302 , \30300 , \30301 );
xnor \U$29959 ( \30303 , \30302 , \27254 );
and \U$29960 ( \30304 , \30298 , \30303 );
and \U$29961 ( \30305 , \30294 , \30303 );
or \U$29962 ( \30306 , \30299 , \30304 , \30305 );
and \U$29963 ( \30307 , \30289 , \30306 );
and \U$29964 ( \30308 , \30273 , \30306 );
or \U$29965 ( \30309 , \30290 , \30307 , \30308 );
and \U$29966 ( \30310 , \30254 , \30309 );
and \U$29967 ( \30311 , \22204 , \25631 );
and \U$29968 ( \30312 , \22099 , \25629 );
nor \U$29969 ( \30313 , \30311 , \30312 );
xnor \U$29970 ( \30314 , \30313 , \25399 );
and \U$29971 ( \30315 , \22325 , \25180 );
and \U$29972 ( \30316 , \22209 , \25178 );
nor \U$29973 ( \30317 , \30315 , \30316 );
xnor \U$29974 ( \30318 , \30317 , \25037 );
and \U$29975 ( \30319 , \30314 , \30318 );
and \U$29976 ( \30320 , \22616 , \24857 );
and \U$29977 ( \30321 , \22440 , \24855 );
nor \U$29978 ( \30322 , \30320 , \30321 );
xnor \U$29979 ( \30323 , \30322 , \24611 );
and \U$29980 ( \30324 , \30318 , \30323 );
and \U$29981 ( \30325 , \30314 , \30323 );
or \U$29982 ( \30326 , \30319 , \30324 , \30325 );
and \U$29983 ( \30327 , \23665 , \23421 );
and \U$29984 ( \30328 , \23491 , \23419 );
nor \U$29985 ( \30329 , \30327 , \30328 );
xnor \U$29986 ( \30330 , \30329 , \23279 );
and \U$29987 ( \30331 , \23970 , \23125 );
and \U$29988 ( \30332 , \23832 , \23123 );
nor \U$29989 ( \30333 , \30331 , \30332 );
xnor \U$29990 ( \30334 , \30333 , \22988 );
and \U$29991 ( \30335 , \30330 , \30334 );
and \U$29992 ( \30336 , \24506 , \22919 );
and \U$29993 ( \30337 , \24089 , \22917 );
nor \U$29994 ( \30338 , \30336 , \30337 );
xnor \U$29995 ( \30339 , \30338 , \22767 );
and \U$29996 ( \30340 , \30334 , \30339 );
and \U$29997 ( \30341 , \30330 , \30339 );
or \U$29998 ( \30342 , \30335 , \30340 , \30341 );
and \U$29999 ( \30343 , \30326 , \30342 );
and \U$30000 ( \30344 , \22867 , \24462 );
and \U$30001 ( \30345 , \22624 , \24460 );
nor \U$30002 ( \30346 , \30344 , \30345 );
xnor \U$30003 ( \30347 , \30346 , \24275 );
and \U$30004 ( \30348 , \23058 , \24149 );
and \U$30005 ( \30349 , \22872 , \24147 );
nor \U$30006 ( \30350 , \30348 , \30349 );
xnor \U$30007 ( \30351 , \30350 , \23944 );
and \U$30008 ( \30352 , \30347 , \30351 );
and \U$30009 ( \30353 , \23466 , \23743 );
and \U$30010 ( \30354 , \23202 , \23741 );
nor \U$30011 ( \30355 , \30353 , \30354 );
xnor \U$30012 ( \30356 , \30355 , \23594 );
and \U$30013 ( \30357 , \30351 , \30356 );
and \U$30014 ( \30358 , \30347 , \30356 );
or \U$30015 ( \30359 , \30352 , \30357 , \30358 );
and \U$30016 ( \30360 , \30342 , \30359 );
and \U$30017 ( \30361 , \30326 , \30359 );
or \U$30018 ( \30362 , \30343 , \30360 , \30361 );
and \U$30019 ( \30363 , \30309 , \30362 );
and \U$30020 ( \30364 , \30254 , \30362 );
or \U$30021 ( \30365 , \30310 , \30363 , \30364 );
and \U$30022 ( \30366 , \29198 , \21434 );
and \U$30023 ( \30367 , \28952 , \21432 );
nor \U$30024 ( \30368 , \30366 , \30367 );
xnor \U$30025 ( \30369 , \30368 , \21441 );
and \U$30026 ( \30370 , \29522 , \21450 );
and \U$30027 ( \30371 , \29203 , \21448 );
nor \U$30028 ( \30372 , \30370 , \30371 );
xnor \U$30029 ( \30373 , \30372 , \21457 );
and \U$30030 ( \30374 , \30369 , \30373 );
buf \U$30031 ( \30375 , RIbb33120_187);
and \U$30032 ( \30376 , \30375 , \21469 );
and \U$30033 ( \30377 , \29806 , \21467 );
nor \U$30034 ( \30378 , \30376 , \30377 );
xnor \U$30035 ( \30379 , \30378 , \21476 );
and \U$30036 ( \30380 , \30373 , \30379 );
and \U$30037 ( \30381 , \30369 , \30379 );
or \U$30038 ( \30382 , \30374 , \30380 , \30381 );
buf \U$30039 ( \30383 , RIbb33198_188);
and \U$30040 ( \30384 , \30383 , \21464 );
buf \U$30041 ( \30385 , \30384 );
and \U$30042 ( \30386 , \30382 , \30385 );
and \U$30043 ( \30387 , \30375 , \21464 );
and \U$30044 ( \30388 , \30385 , \30387 );
and \U$30045 ( \30389 , \30382 , \30387 );
or \U$30046 ( \30390 , \30386 , \30388 , \30389 );
xor \U$30047 ( \30391 , \29925 , \29929 );
xor \U$30048 ( \30392 , \30391 , \29934 );
xor \U$30049 ( \30393 , \30054 , \30058 );
xor \U$30050 ( \30394 , \30393 , \30063 );
and \U$30051 ( \30395 , \30392 , \30394 );
xor \U$30052 ( \30396 , \30070 , \30074 );
xor \U$30053 ( \30397 , \30396 , \30079 );
and \U$30054 ( \30398 , \30394 , \30397 );
and \U$30055 ( \30399 , \30392 , \30397 );
or \U$30056 ( \30400 , \30395 , \30398 , \30399 );
and \U$30057 ( \30401 , \30390 , \30400 );
xor \U$30058 ( \30402 , \30087 , \30091 );
xor \U$30059 ( \30403 , \30402 , \30096 );
xor \U$30060 ( \30404 , \30001 , \30005 );
xor \U$30061 ( \30405 , \30404 , \30010 );
and \U$30062 ( \30406 , \30403 , \30405 );
xor \U$30063 ( \30407 , \30017 , \30021 );
xor \U$30064 ( \30408 , \30407 , \30026 );
and \U$30065 ( \30409 , \30405 , \30408 );
and \U$30066 ( \30410 , \30403 , \30408 );
or \U$30067 ( \30411 , \30406 , \30409 , \30410 );
and \U$30068 ( \30412 , \30400 , \30411 );
and \U$30069 ( \30413 , \30390 , \30411 );
or \U$30070 ( \30414 , \30401 , \30412 , \30413 );
and \U$30071 ( \30415 , \30365 , \30414 );
xor \U$30072 ( \30416 , \29965 , \29969 );
xor \U$30073 ( \30417 , \30416 , \29974 );
xor \U$30074 ( \30418 , \29982 , \29986 );
xor \U$30075 ( \30419 , \30418 , \29991 );
and \U$30076 ( \30420 , \30417 , \30419 );
xor \U$30077 ( \30421 , \30034 , \30038 );
xor \U$30078 ( \30422 , \30421 , \30043 );
and \U$30079 ( \30423 , \30419 , \30422 );
and \U$30080 ( \30424 , \30417 , \30422 );
or \U$30081 ( \30425 , \30420 , \30423 , \30424 );
xor \U$30082 ( \30426 , \30108 , \30110 );
xor \U$30083 ( \30427 , \30426 , \30113 );
and \U$30084 ( \30428 , \30425 , \30427 );
xor \U$30085 ( \30429 , \29912 , \29914 );
xor \U$30086 ( \30430 , \30429 , \29917 );
and \U$30087 ( \30431 , \30427 , \30430 );
and \U$30088 ( \30432 , \30425 , \30430 );
or \U$30089 ( \30433 , \30428 , \30431 , \30432 );
and \U$30090 ( \30434 , \30414 , \30433 );
and \U$30091 ( \30435 , \30365 , \30433 );
or \U$30092 ( \30436 , \30415 , \30434 , \30435 );
xor \U$30093 ( \30437 , \29910 , \29920 );
xor \U$30094 ( \30438 , \30437 , \29940 );
xor \U$30095 ( \30439 , \29997 , \30049 );
xor \U$30096 ( \30440 , \30439 , \30102 );
and \U$30097 ( \30441 , \30438 , \30440 );
xor \U$30098 ( \30442 , \30116 , \30118 );
xor \U$30099 ( \30443 , \30442 , \30121 );
and \U$30100 ( \30444 , \30440 , \30443 );
and \U$30101 ( \30445 , \30438 , \30443 );
or \U$30102 ( \30446 , \30441 , \30444 , \30445 );
and \U$30103 ( \30447 , \30436 , \30446 );
xor \U$30104 ( \30448 , \30066 , \30082 );
xor \U$30105 ( \30449 , \30448 , \30099 );
xor \U$30106 ( \30450 , \29902 , \29904 );
xor \U$30107 ( \30451 , \30450 , \29907 );
and \U$30108 ( \30452 , \30449 , \30451 );
xnor \U$30109 ( \30453 , \29937 , \29939 );
and \U$30110 ( \30454 , \30451 , \30453 );
and \U$30111 ( \30455 , \30449 , \30453 );
or \U$30112 ( \30456 , \30452 , \30454 , \30455 );
xor \U$30113 ( \30457 , \30129 , \30131 );
xor \U$30114 ( \30458 , \30457 , \30134 );
and \U$30115 ( \30459 , \30456 , \30458 );
xor \U$30116 ( \30460 , \30139 , \30141 );
xor \U$30117 ( \30461 , \30460 , \30144 );
and \U$30118 ( \30462 , \30458 , \30461 );
and \U$30119 ( \30463 , \30456 , \30461 );
or \U$30120 ( \30464 , \30459 , \30462 , \30463 );
and \U$30121 ( \30465 , \30446 , \30464 );
and \U$30122 ( \30466 , \30436 , \30464 );
or \U$30123 ( \30467 , \30447 , \30465 , \30466 );
xor \U$30124 ( \30468 , \29664 , \29716 );
xor \U$30125 ( \30469 , \30468 , \29772 );
xor \U$30126 ( \30470 , \29785 , \29795 );
xor \U$30127 ( \30471 , \30470 , \29818 );
and \U$30128 ( \30472 , \30469 , \30471 );
xor \U$30129 ( \30473 , \30156 , \30158 );
xor \U$30130 ( \30474 , \30473 , \30161 );
and \U$30131 ( \30475 , \30471 , \30474 );
and \U$30132 ( \30476 , \30469 , \30474 );
or \U$30133 ( \30477 , \30472 , \30475 , \30476 );
and \U$30134 ( \30478 , \30467 , \30477 );
xor \U$30135 ( \30479 , \30169 , \30171 );
xor \U$30136 ( \30480 , \30479 , \30174 );
and \U$30137 ( \30481 , \30477 , \30480 );
and \U$30138 ( \30482 , \30467 , \30480 );
or \U$30139 ( \30483 , \30478 , \30481 , \30482 );
xor \U$30140 ( \30484 , \29835 , \29853 );
xor \U$30141 ( \30485 , \30484 , \29864 );
and \U$30142 ( \30486 , \30483 , \30485 );
xor \U$30143 ( \30487 , \30167 , \30177 );
xor \U$30144 ( \30488 , \30487 , \30180 );
and \U$30145 ( \30489 , \30485 , \30488 );
and \U$30146 ( \30490 , \30483 , \30488 );
or \U$30147 ( \30491 , \30486 , \30489 , \30490 );
xor \U$30148 ( \30492 , \30183 , \30185 );
xor \U$30149 ( \30493 , \30492 , \30187 );
and \U$30150 ( \30494 , \30491 , \30493 );
and \U$30151 ( \30495 , \30202 , \30494 );
xor \U$30152 ( \30496 , \30202 , \30494 );
xor \U$30153 ( \30497 , \30491 , \30493 );
and \U$30154 ( \30498 , \23491 , \23743 );
and \U$30155 ( \30499 , \23466 , \23741 );
nor \U$30156 ( \30500 , \30498 , \30499 );
xnor \U$30157 ( \30501 , \30500 , \23594 );
and \U$30158 ( \30502 , \23832 , \23421 );
and \U$30159 ( \30503 , \23665 , \23419 );
nor \U$30160 ( \30504 , \30502 , \30503 );
xnor \U$30161 ( \30505 , \30504 , \23279 );
and \U$30162 ( \30506 , \30501 , \30505 );
and \U$30163 ( \30507 , \24089 , \23125 );
and \U$30164 ( \30508 , \23970 , \23123 );
nor \U$30165 ( \30509 , \30507 , \30508 );
xnor \U$30166 ( \30510 , \30509 , \22988 );
and \U$30167 ( \30511 , \30505 , \30510 );
and \U$30168 ( \30512 , \30501 , \30510 );
or \U$30169 ( \30513 , \30506 , \30511 , \30512 );
and \U$30170 ( \30514 , \22624 , \24857 );
and \U$30171 ( \30515 , \22616 , \24855 );
nor \U$30172 ( \30516 , \30514 , \30515 );
xnor \U$30173 ( \30517 , \30516 , \24611 );
and \U$30174 ( \30518 , \22872 , \24462 );
and \U$30175 ( \30519 , \22867 , \24460 );
nor \U$30176 ( \30520 , \30518 , \30519 );
xnor \U$30177 ( \30521 , \30520 , \24275 );
and \U$30178 ( \30522 , \30517 , \30521 );
and \U$30179 ( \30523 , \23202 , \24149 );
and \U$30180 ( \30524 , \23058 , \24147 );
nor \U$30181 ( \30525 , \30523 , \30524 );
xnor \U$30182 ( \30526 , \30525 , \23944 );
and \U$30183 ( \30527 , \30521 , \30526 );
and \U$30184 ( \30528 , \30517 , \30526 );
or \U$30185 ( \30529 , \30522 , \30527 , \30528 );
and \U$30186 ( \30530 , \30513 , \30529 );
and \U$30187 ( \30531 , \22099 , \26005 );
and \U$30188 ( \30532 , \22011 , \26003 );
nor \U$30189 ( \30533 , \30531 , \30532 );
xnor \U$30190 ( \30534 , \30533 , \25817 );
and \U$30191 ( \30535 , \22209 , \25631 );
and \U$30192 ( \30536 , \22204 , \25629 );
nor \U$30193 ( \30537 , \30535 , \30536 );
xnor \U$30194 ( \30538 , \30537 , \25399 );
and \U$30195 ( \30539 , \30534 , \30538 );
and \U$30196 ( \30540 , \22440 , \25180 );
and \U$30197 ( \30541 , \22325 , \25178 );
nor \U$30198 ( \30542 , \30540 , \30541 );
xnor \U$30199 ( \30543 , \30542 , \25037 );
and \U$30200 ( \30544 , \30538 , \30543 );
and \U$30201 ( \30545 , \30534 , \30543 );
or \U$30202 ( \30546 , \30539 , \30544 , \30545 );
and \U$30203 ( \30547 , \30529 , \30546 );
and \U$30204 ( \30548 , \30513 , \30546 );
or \U$30205 ( \30549 , \30530 , \30547 , \30548 );
and \U$30206 ( \30550 , \21463 , \27569 );
and \U$30207 ( \30551 , \21471 , \27567 );
nor \U$30208 ( \30552 , \30550 , \30551 );
xnor \U$30209 ( \30553 , \30552 , \27254 );
and \U$30210 ( \30554 , \21689 , \27060 );
and \U$30211 ( \30555 , \21478 , \27058 );
nor \U$30212 ( \30556 , \30554 , \30555 );
xnor \U$30213 ( \30557 , \30556 , \26720 );
and \U$30214 ( \30558 , \30553 , \30557 );
and \U$30215 ( \30559 , \21813 , \26471 );
and \U$30216 ( \30560 , \21750 , \26469 );
nor \U$30217 ( \30561 , \30559 , \30560 );
xnor \U$30218 ( \30562 , \30561 , \26230 );
and \U$30219 ( \30563 , \30557 , \30562 );
and \U$30220 ( \30564 , \30553 , \30562 );
or \U$30221 ( \30565 , \30558 , \30563 , \30564 );
and \U$30222 ( \30566 , \21413 , \29159 );
and \U$30223 ( \30567 , \21421 , \29157 );
nor \U$30224 ( \30568 , \30566 , \30567 );
xnor \U$30225 ( \30569 , \30568 , \28841 );
and \U$30226 ( \30570 , \21428 , \28592 );
and \U$30227 ( \30571 , \21436 , \28590 );
nor \U$30228 ( \30572 , \30570 , \30571 );
xnor \U$30229 ( \30573 , \30572 , \28343 );
and \U$30230 ( \30574 , \30569 , \30573 );
and \U$30231 ( \30575 , \21444 , \28063 );
and \U$30232 ( \30576 , \21452 , \28061 );
nor \U$30233 ( \30577 , \30575 , \30576 );
xnor \U$30234 ( \30578 , \30577 , \27803 );
and \U$30235 ( \30579 , \30573 , \30578 );
and \U$30236 ( \30580 , \30569 , \30578 );
or \U$30237 ( \30581 , \30574 , \30579 , \30580 );
and \U$30238 ( \30582 , \30565 , \30581 );
buf \U$30239 ( \30583 , RIbb2d978_62);
buf \U$30240 ( \30584 , RIbb2d900_63);
and \U$30241 ( \30585 , \30583 , \30584 );
not \U$30242 ( \30586 , \30585 );
and \U$30243 ( \30587 , \29945 , \30586 );
not \U$30244 ( \30588 , \30587 );
and \U$30245 ( \30589 , \21379 , \30258 );
and \U$30246 ( \30590 , \21387 , \30256 );
nor \U$30247 ( \30591 , \30589 , \30590 );
xnor \U$30248 ( \30592 , \30591 , \29948 );
and \U$30249 ( \30593 , \30588 , \30592 );
and \U$30250 ( \30594 , \21395 , \29721 );
and \U$30251 ( \30595 , \21403 , \29719 );
nor \U$30252 ( \30596 , \30594 , \30595 );
xnor \U$30253 ( \30597 , \30596 , \29350 );
and \U$30254 ( \30598 , \30592 , \30597 );
and \U$30255 ( \30599 , \30588 , \30597 );
or \U$30256 ( \30600 , \30593 , \30598 , \30599 );
and \U$30257 ( \30601 , \30581 , \30600 );
and \U$30258 ( \30602 , \30565 , \30600 );
or \U$30259 ( \30603 , \30582 , \30601 , \30602 );
and \U$30260 ( \30604 , \30549 , \30603 );
and \U$30261 ( \30605 , \26982 , \21652 );
and \U$30262 ( \30606 , \26973 , \21650 );
nor \U$30263 ( \30607 , \30605 , \30606 );
xnor \U$30264 ( \30608 , \30607 , \21377 );
and \U$30265 ( \30609 , \27527 , \21385 );
and \U$30266 ( \30610 , \27325 , \21383 );
nor \U$30267 ( \30611 , \30609 , \30610 );
xnor \U$30268 ( \30612 , \30611 , \21392 );
and \U$30269 ( \30613 , \30608 , \30612 );
and \U$30270 ( \30614 , \28002 , \21401 );
and \U$30271 ( \30615 , \27830 , \21399 );
nor \U$30272 ( \30616 , \30614 , \30615 );
xnor \U$30273 ( \30617 , \30616 , \21408 );
and \U$30274 ( \30618 , \30612 , \30617 );
and \U$30275 ( \30619 , \30608 , \30617 );
or \U$30276 ( \30620 , \30613 , \30618 , \30619 );
and \U$30277 ( \30621 , \25604 , \22185 );
and \U$30278 ( \30622 , \25596 , \22183 );
nor \U$30279 ( \30623 , \30621 , \30622 );
xnor \U$30280 ( \30624 , \30623 , \22049 );
and \U$30281 ( \30625 , \26078 , \21985 );
and \U$30282 ( \30626 , \26073 , \21983 );
nor \U$30283 ( \30627 , \30625 , \30626 );
xnor \U$30284 ( \30628 , \30627 , \21907 );
and \U$30285 ( \30629 , \30624 , \30628 );
and \U$30286 ( \30630 , \26601 , \21821 );
and \U$30287 ( \30631 , \26342 , \21819 );
nor \U$30288 ( \30632 , \30630 , \30631 );
xnor \U$30289 ( \30633 , \30632 , \21727 );
and \U$30290 ( \30634 , \30628 , \30633 );
and \U$30291 ( \30635 , \30624 , \30633 );
or \U$30292 ( \30636 , \30629 , \30634 , \30635 );
and \U$30293 ( \30637 , \30620 , \30636 );
and \U$30294 ( \30638 , \24714 , \22919 );
and \U$30295 ( \30639 , \24506 , \22917 );
nor \U$30296 ( \30640 , \30638 , \30639 );
xnor \U$30297 ( \30641 , \30640 , \22767 );
and \U$30298 ( \30642 , \24841 , \22651 );
and \U$30299 ( \30643 , \24836 , \22649 );
nor \U$30300 ( \30644 , \30642 , \30643 );
xnor \U$30301 ( \30645 , \30644 , \22495 );
and \U$30302 ( \30646 , \30641 , \30645 );
and \U$30303 ( \30647 , \25294 , \22379 );
and \U$30304 ( \30648 , \25097 , \22377 );
nor \U$30305 ( \30649 , \30647 , \30648 );
xnor \U$30306 ( \30650 , \30649 , \22266 );
and \U$30307 ( \30651 , \30645 , \30650 );
and \U$30308 ( \30652 , \30641 , \30650 );
or \U$30309 ( \30653 , \30646 , \30651 , \30652 );
and \U$30310 ( \30654 , \30636 , \30653 );
and \U$30311 ( \30655 , \30620 , \30653 );
or \U$30312 ( \30656 , \30637 , \30654 , \30655 );
and \U$30313 ( \30657 , \30603 , \30656 );
and \U$30314 ( \30658 , \30549 , \30656 );
or \U$30315 ( \30659 , \30604 , \30657 , \30658 );
xor \U$30316 ( \30660 , \30314 , \30318 );
xor \U$30317 ( \30661 , \30660 , \30323 );
xor \U$30318 ( \30662 , \30330 , \30334 );
xor \U$30319 ( \30663 , \30662 , \30339 );
and \U$30320 ( \30664 , \30661 , \30663 );
xor \U$30321 ( \30665 , \30347 , \30351 );
xor \U$30322 ( \30666 , \30665 , \30356 );
and \U$30323 ( \30667 , \30663 , \30666 );
and \U$30324 ( \30668 , \30661 , \30666 );
or \U$30325 ( \30669 , \30664 , \30667 , \30668 );
xor \U$30326 ( \30670 , \30206 , \30210 );
xor \U$30327 ( \30671 , \30670 , \30215 );
xor \U$30328 ( \30672 , \30222 , \30226 );
xor \U$30329 ( \30673 , \30672 , \30231 );
and \U$30330 ( \30674 , \30671 , \30673 );
xor \U$30331 ( \30675 , \30239 , \30243 );
xor \U$30332 ( \30676 , \30675 , \30248 );
and \U$30333 ( \30677 , \30673 , \30676 );
and \U$30334 ( \30678 , \30671 , \30676 );
or \U$30335 ( \30679 , \30674 , \30677 , \30678 );
and \U$30336 ( \30680 , \30669 , \30679 );
and \U$30337 ( \30681 , \28952 , \21419 );
and \U$30338 ( \30682 , \28528 , \21417 );
nor \U$30339 ( \30683 , \30681 , \30682 );
xnor \U$30340 ( \30684 , \30683 , \21426 );
and \U$30341 ( \30685 , \29203 , \21434 );
and \U$30342 ( \30686 , \29198 , \21432 );
nor \U$30343 ( \30687 , \30685 , \30686 );
xnor \U$30344 ( \30688 , \30687 , \21441 );
and \U$30345 ( \30689 , \30684 , \30688 );
and \U$30346 ( \30690 , \29806 , \21450 );
and \U$30347 ( \30691 , \29522 , \21448 );
nor \U$30348 ( \30692 , \30690 , \30691 );
xnor \U$30349 ( \30693 , \30692 , \21457 );
and \U$30350 ( \30694 , \30688 , \30693 );
and \U$30351 ( \30695 , \30684 , \30693 );
or \U$30352 ( \30696 , \30689 , \30694 , \30695 );
xor \U$30353 ( \30697 , \30369 , \30373 );
xor \U$30354 ( \30698 , \30697 , \30379 );
and \U$30355 ( \30699 , \30696 , \30698 );
not \U$30356 ( \30700 , \30384 );
and \U$30357 ( \30701 , \30698 , \30700 );
and \U$30358 ( \30702 , \30696 , \30700 );
or \U$30359 ( \30703 , \30699 , \30701 , \30702 );
and \U$30360 ( \30704 , \30679 , \30703 );
and \U$30361 ( \30705 , \30669 , \30703 );
or \U$30362 ( \30706 , \30680 , \30704 , \30705 );
and \U$30363 ( \30707 , \30659 , \30706 );
xor \U$30364 ( \30708 , \30261 , \30265 );
xor \U$30365 ( \30709 , \30708 , \30270 );
xor \U$30366 ( \30710 , \30277 , \30281 );
xor \U$30367 ( \30711 , \30710 , \30286 );
and \U$30368 ( \30712 , \30709 , \30711 );
xor \U$30369 ( \30713 , \30294 , \30298 );
xor \U$30370 ( \30714 , \30713 , \30303 );
and \U$30371 ( \30715 , \30711 , \30714 );
and \U$30372 ( \30716 , \30709 , \30714 );
or \U$30373 ( \30717 , \30712 , \30715 , \30716 );
xor \U$30374 ( \30718 , \29949 , \29953 );
xor \U$30375 ( \30719 , \30718 , \29958 );
and \U$30376 ( \30720 , \30717 , \30719 );
xor \U$30377 ( \30721 , \30417 , \30419 );
xor \U$30378 ( \30722 , \30721 , \30422 );
and \U$30379 ( \30723 , \30719 , \30722 );
and \U$30380 ( \30724 , \30717 , \30722 );
or \U$30381 ( \30725 , \30720 , \30723 , \30724 );
and \U$30382 ( \30726 , \30706 , \30725 );
and \U$30383 ( \30727 , \30659 , \30725 );
or \U$30384 ( \30728 , \30707 , \30726 , \30727 );
xor \U$30385 ( \30729 , \30218 , \30234 );
xor \U$30386 ( \30730 , \30729 , \30251 );
xor \U$30387 ( \30731 , \30273 , \30289 );
xor \U$30388 ( \30732 , \30731 , \30306 );
and \U$30389 ( \30733 , \30730 , \30732 );
xor \U$30390 ( \30734 , \30326 , \30342 );
xor \U$30391 ( \30735 , \30734 , \30359 );
and \U$30392 ( \30736 , \30732 , \30735 );
and \U$30393 ( \30737 , \30730 , \30735 );
or \U$30394 ( \30738 , \30733 , \30736 , \30737 );
xor \U$30395 ( \30739 , \30382 , \30385 );
xor \U$30396 ( \30740 , \30739 , \30387 );
xor \U$30397 ( \30741 , \30392 , \30394 );
xor \U$30398 ( \30742 , \30741 , \30397 );
and \U$30399 ( \30743 , \30740 , \30742 );
xor \U$30400 ( \30744 , \30403 , \30405 );
xor \U$30401 ( \30745 , \30744 , \30408 );
and \U$30402 ( \30746 , \30742 , \30745 );
and \U$30403 ( \30747 , \30740 , \30745 );
or \U$30404 ( \30748 , \30743 , \30746 , \30747 );
and \U$30405 ( \30749 , \30738 , \30748 );
xor \U$30406 ( \30750 , \30013 , \30029 );
xor \U$30407 ( \30751 , \30750 , \30046 );
and \U$30408 ( \30752 , \30748 , \30751 );
and \U$30409 ( \30753 , \30738 , \30751 );
or \U$30410 ( \30754 , \30749 , \30752 , \30753 );
and \U$30411 ( \30755 , \30728 , \30754 );
xor \U$30412 ( \30756 , \29961 , \29977 );
xor \U$30413 ( \30757 , \30756 , \29994 );
xor \U$30414 ( \30758 , \30425 , \30427 );
xor \U$30415 ( \30759 , \30758 , \30430 );
and \U$30416 ( \30760 , \30757 , \30759 );
xor \U$30417 ( \30761 , \30449 , \30451 );
xor \U$30418 ( \30762 , \30761 , \30453 );
and \U$30419 ( \30763 , \30759 , \30762 );
and \U$30420 ( \30764 , \30757 , \30762 );
or \U$30421 ( \30765 , \30760 , \30763 , \30764 );
and \U$30422 ( \30766 , \30754 , \30765 );
and \U$30423 ( \30767 , \30728 , \30765 );
or \U$30424 ( \30768 , \30755 , \30766 , \30767 );
xor \U$30425 ( \30769 , \30365 , \30414 );
xor \U$30426 ( \30770 , \30769 , \30433 );
xor \U$30427 ( \30771 , \30438 , \30440 );
xor \U$30428 ( \30772 , \30771 , \30443 );
and \U$30429 ( \30773 , \30770 , \30772 );
xor \U$30430 ( \30774 , \30456 , \30458 );
xor \U$30431 ( \30775 , \30774 , \30461 );
and \U$30432 ( \30776 , \30772 , \30775 );
and \U$30433 ( \30777 , \30770 , \30775 );
or \U$30434 ( \30778 , \30773 , \30776 , \30777 );
and \U$30435 ( \30779 , \30768 , \30778 );
xor \U$30436 ( \30780 , \30137 , \30147 );
xor \U$30437 ( \30781 , \30780 , \30150 );
and \U$30438 ( \30782 , \30778 , \30781 );
and \U$30439 ( \30783 , \30768 , \30781 );
or \U$30440 ( \30784 , \30779 , \30782 , \30783 );
xor \U$30441 ( \30785 , \29943 , \30105 );
xor \U$30442 ( \30786 , \30785 , \30124 );
xor \U$30443 ( \30787 , \30436 , \30446 );
xor \U$30444 ( \30788 , \30787 , \30464 );
and \U$30445 ( \30789 , \30786 , \30788 );
xor \U$30446 ( \30790 , \30469 , \30471 );
xor \U$30447 ( \30791 , \30790 , \30474 );
and \U$30448 ( \30792 , \30788 , \30791 );
and \U$30449 ( \30793 , \30786 , \30791 );
or \U$30450 ( \30794 , \30789 , \30792 , \30793 );
and \U$30451 ( \30795 , \30784 , \30794 );
xor \U$30452 ( \30796 , \30127 , \30153 );
xor \U$30453 ( \30797 , \30796 , \30164 );
and \U$30454 ( \30798 , \30794 , \30797 );
and \U$30455 ( \30799 , \30784 , \30797 );
or \U$30456 ( \30800 , \30795 , \30798 , \30799 );
xor \U$30457 ( \30801 , \30483 , \30485 );
xor \U$30458 ( \30802 , \30801 , \30488 );
and \U$30459 ( \30803 , \30800 , \30802 );
and \U$30460 ( \30804 , \30497 , \30803 );
xor \U$30461 ( \30805 , \30497 , \30803 );
xor \U$30462 ( \30806 , \30800 , \30802 );
and \U$30463 ( \30807 , \21478 , \27569 );
and \U$30464 ( \30808 , \21463 , \27567 );
nor \U$30465 ( \30809 , \30807 , \30808 );
xnor \U$30466 ( \30810 , \30809 , \27254 );
and \U$30467 ( \30811 , \21750 , \27060 );
and \U$30468 ( \30812 , \21689 , \27058 );
nor \U$30469 ( \30813 , \30811 , \30812 );
xnor \U$30470 ( \30814 , \30813 , \26720 );
and \U$30471 ( \30815 , \30810 , \30814 );
and \U$30472 ( \30816 , \22011 , \26471 );
and \U$30473 ( \30817 , \21813 , \26469 );
nor \U$30474 ( \30818 , \30816 , \30817 );
xnor \U$30475 ( \30819 , \30818 , \26230 );
and \U$30476 ( \30820 , \30814 , \30819 );
and \U$30477 ( \30821 , \30810 , \30819 );
or \U$30478 ( \30822 , \30815 , \30820 , \30821 );
xor \U$30479 ( \30823 , \29945 , \30583 );
xor \U$30480 ( \30824 , \30583 , \30584 );
not \U$30481 ( \30825 , \30824 );
and \U$30482 ( \30826 , \30823 , \30825 );
and \U$30483 ( \30827 , \21387 , \30826 );
not \U$30484 ( \30828 , \30827 );
xnor \U$30485 ( \30829 , \30828 , \30587 );
and \U$30486 ( \30830 , \21403 , \30258 );
and \U$30487 ( \30831 , \21379 , \30256 );
nor \U$30488 ( \30832 , \30830 , \30831 );
xnor \U$30489 ( \30833 , \30832 , \29948 );
and \U$30490 ( \30834 , \30829 , \30833 );
and \U$30491 ( \30835 , \21421 , \29721 );
and \U$30492 ( \30836 , \21395 , \29719 );
nor \U$30493 ( \30837 , \30835 , \30836 );
xnor \U$30494 ( \30838 , \30837 , \29350 );
and \U$30495 ( \30839 , \30833 , \30838 );
and \U$30496 ( \30840 , \30829 , \30838 );
or \U$30497 ( \30841 , \30834 , \30839 , \30840 );
and \U$30498 ( \30842 , \30822 , \30841 );
and \U$30499 ( \30843 , \21436 , \29159 );
and \U$30500 ( \30844 , \21413 , \29157 );
nor \U$30501 ( \30845 , \30843 , \30844 );
xnor \U$30502 ( \30846 , \30845 , \28841 );
and \U$30503 ( \30847 , \21452 , \28592 );
and \U$30504 ( \30848 , \21428 , \28590 );
nor \U$30505 ( \30849 , \30847 , \30848 );
xnor \U$30506 ( \30850 , \30849 , \28343 );
and \U$30507 ( \30851 , \30846 , \30850 );
and \U$30508 ( \30852 , \21471 , \28063 );
and \U$30509 ( \30853 , \21444 , \28061 );
nor \U$30510 ( \30854 , \30852 , \30853 );
xnor \U$30511 ( \30855 , \30854 , \27803 );
and \U$30512 ( \30856 , \30850 , \30855 );
and \U$30513 ( \30857 , \30846 , \30855 );
or \U$30514 ( \30858 , \30851 , \30856 , \30857 );
and \U$30515 ( \30859 , \30841 , \30858 );
and \U$30516 ( \30860 , \30822 , \30858 );
or \U$30517 ( \30861 , \30842 , \30859 , \30860 );
and \U$30518 ( \30862 , \27325 , \21652 );
and \U$30519 ( \30863 , \26982 , \21650 );
nor \U$30520 ( \30864 , \30862 , \30863 );
xnor \U$30521 ( \30865 , \30864 , \21377 );
and \U$30522 ( \30866 , \27830 , \21385 );
and \U$30523 ( \30867 , \27527 , \21383 );
nor \U$30524 ( \30868 , \30866 , \30867 );
xnor \U$30525 ( \30869 , \30868 , \21392 );
and \U$30526 ( \30870 , \30865 , \30869 );
and \U$30527 ( \30871 , \28528 , \21401 );
and \U$30528 ( \30872 , \28002 , \21399 );
nor \U$30529 ( \30873 , \30871 , \30872 );
xnor \U$30530 ( \30874 , \30873 , \21408 );
and \U$30531 ( \30875 , \30869 , \30874 );
and \U$30532 ( \30876 , \30865 , \30874 );
or \U$30533 ( \30877 , \30870 , \30875 , \30876 );
and \U$30534 ( \30878 , \24836 , \22919 );
and \U$30535 ( \30879 , \24714 , \22917 );
nor \U$30536 ( \30880 , \30878 , \30879 );
xnor \U$30537 ( \30881 , \30880 , \22767 );
and \U$30538 ( \30882 , \25097 , \22651 );
and \U$30539 ( \30883 , \24841 , \22649 );
nor \U$30540 ( \30884 , \30882 , \30883 );
xnor \U$30541 ( \30885 , \30884 , \22495 );
and \U$30542 ( \30886 , \30881 , \30885 );
and \U$30543 ( \30887 , \25596 , \22379 );
and \U$30544 ( \30888 , \25294 , \22377 );
nor \U$30545 ( \30889 , \30887 , \30888 );
xnor \U$30546 ( \30890 , \30889 , \22266 );
and \U$30547 ( \30891 , \30885 , \30890 );
and \U$30548 ( \30892 , \30881 , \30890 );
or \U$30549 ( \30893 , \30886 , \30891 , \30892 );
and \U$30550 ( \30894 , \30877 , \30893 );
and \U$30551 ( \30895 , \26073 , \22185 );
and \U$30552 ( \30896 , \25604 , \22183 );
nor \U$30553 ( \30897 , \30895 , \30896 );
xnor \U$30554 ( \30898 , \30897 , \22049 );
and \U$30555 ( \30899 , \26342 , \21985 );
and \U$30556 ( \30900 , \26078 , \21983 );
nor \U$30557 ( \30901 , \30899 , \30900 );
xnor \U$30558 ( \30902 , \30901 , \21907 );
and \U$30559 ( \30903 , \30898 , \30902 );
and \U$30560 ( \30904 , \26973 , \21821 );
and \U$30561 ( \30905 , \26601 , \21819 );
nor \U$30562 ( \30906 , \30904 , \30905 );
xnor \U$30563 ( \30907 , \30906 , \21727 );
and \U$30564 ( \30908 , \30902 , \30907 );
and \U$30565 ( \30909 , \30898 , \30907 );
or \U$30566 ( \30910 , \30903 , \30908 , \30909 );
and \U$30567 ( \30911 , \30893 , \30910 );
and \U$30568 ( \30912 , \30877 , \30910 );
or \U$30569 ( \30913 , \30894 , \30911 , \30912 );
and \U$30570 ( \30914 , \30861 , \30913 );
and \U$30571 ( \30915 , \22204 , \26005 );
and \U$30572 ( \30916 , \22099 , \26003 );
nor \U$30573 ( \30917 , \30915 , \30916 );
xnor \U$30574 ( \30918 , \30917 , \25817 );
and \U$30575 ( \30919 , \22325 , \25631 );
and \U$30576 ( \30920 , \22209 , \25629 );
nor \U$30577 ( \30921 , \30919 , \30920 );
xnor \U$30578 ( \30922 , \30921 , \25399 );
and \U$30579 ( \30923 , \30918 , \30922 );
and \U$30580 ( \30924 , \22616 , \25180 );
and \U$30581 ( \30925 , \22440 , \25178 );
nor \U$30582 ( \30926 , \30924 , \30925 );
xnor \U$30583 ( \30927 , \30926 , \25037 );
and \U$30584 ( \30928 , \30922 , \30927 );
and \U$30585 ( \30929 , \30918 , \30927 );
or \U$30586 ( \30930 , \30923 , \30928 , \30929 );
and \U$30587 ( \30931 , \23665 , \23743 );
and \U$30588 ( \30932 , \23491 , \23741 );
nor \U$30589 ( \30933 , \30931 , \30932 );
xnor \U$30590 ( \30934 , \30933 , \23594 );
and \U$30591 ( \30935 , \23970 , \23421 );
and \U$30592 ( \30936 , \23832 , \23419 );
nor \U$30593 ( \30937 , \30935 , \30936 );
xnor \U$30594 ( \30938 , \30937 , \23279 );
and \U$30595 ( \30939 , \30934 , \30938 );
and \U$30596 ( \30940 , \24506 , \23125 );
and \U$30597 ( \30941 , \24089 , \23123 );
nor \U$30598 ( \30942 , \30940 , \30941 );
xnor \U$30599 ( \30943 , \30942 , \22988 );
and \U$30600 ( \30944 , \30938 , \30943 );
and \U$30601 ( \30945 , \30934 , \30943 );
or \U$30602 ( \30946 , \30939 , \30944 , \30945 );
and \U$30603 ( \30947 , \30930 , \30946 );
and \U$30604 ( \30948 , \22867 , \24857 );
and \U$30605 ( \30949 , \22624 , \24855 );
nor \U$30606 ( \30950 , \30948 , \30949 );
xnor \U$30607 ( \30951 , \30950 , \24611 );
and \U$30608 ( \30952 , \23058 , \24462 );
and \U$30609 ( \30953 , \22872 , \24460 );
nor \U$30610 ( \30954 , \30952 , \30953 );
xnor \U$30611 ( \30955 , \30954 , \24275 );
and \U$30612 ( \30956 , \30951 , \30955 );
and \U$30613 ( \30957 , \23466 , \24149 );
and \U$30614 ( \30958 , \23202 , \24147 );
nor \U$30615 ( \30959 , \30957 , \30958 );
xnor \U$30616 ( \30960 , \30959 , \23944 );
and \U$30617 ( \30961 , \30955 , \30960 );
and \U$30618 ( \30962 , \30951 , \30960 );
or \U$30619 ( \30963 , \30956 , \30961 , \30962 );
and \U$30620 ( \30964 , \30946 , \30963 );
and \U$30621 ( \30965 , \30930 , \30963 );
or \U$30622 ( \30966 , \30947 , \30964 , \30965 );
and \U$30623 ( \30967 , \30913 , \30966 );
and \U$30624 ( \30968 , \30861 , \30966 );
or \U$30625 ( \30969 , \30914 , \30967 , \30968 );
and \U$30626 ( \30970 , \29198 , \21419 );
and \U$30627 ( \30971 , \28952 , \21417 );
nor \U$30628 ( \30972 , \30970 , \30971 );
xnor \U$30629 ( \30973 , \30972 , \21426 );
and \U$30630 ( \30974 , \29522 , \21434 );
and \U$30631 ( \30975 , \29203 , \21432 );
nor \U$30632 ( \30976 , \30974 , \30975 );
xnor \U$30633 ( \30977 , \30976 , \21441 );
and \U$30634 ( \30978 , \30973 , \30977 );
and \U$30635 ( \30979 , \30375 , \21450 );
and \U$30636 ( \30980 , \29806 , \21448 );
nor \U$30637 ( \30981 , \30979 , \30980 );
xnor \U$30638 ( \30982 , \30981 , \21457 );
and \U$30639 ( \30983 , \30977 , \30982 );
and \U$30640 ( \30984 , \30973 , \30982 );
or \U$30641 ( \30985 , \30978 , \30983 , \30984 );
buf \U$30642 ( \30986 , RIbb33210_189);
and \U$30643 ( \30987 , \30986 , \21469 );
and \U$30644 ( \30988 , \30383 , \21467 );
nor \U$30645 ( \30989 , \30987 , \30988 );
xnor \U$30646 ( \30990 , \30989 , \21476 );
buf \U$30647 ( \30991 , RIbb33288_190);
and \U$30648 ( \30992 , \30991 , \21464 );
or \U$30649 ( \30993 , \30990 , \30992 );
and \U$30650 ( \30994 , \30985 , \30993 );
and \U$30651 ( \30995 , \30383 , \21469 );
and \U$30652 ( \30996 , \30375 , \21467 );
nor \U$30653 ( \30997 , \30995 , \30996 );
xnor \U$30654 ( \30998 , \30997 , \21476 );
and \U$30655 ( \30999 , \30993 , \30998 );
and \U$30656 ( \31000 , \30985 , \30998 );
or \U$30657 ( \31001 , \30994 , \30999 , \31000 );
and \U$30658 ( \31002 , \30986 , \21464 );
xor \U$30659 ( \31003 , \30608 , \30612 );
xor \U$30660 ( \31004 , \31003 , \30617 );
and \U$30661 ( \31005 , \31002 , \31004 );
xor \U$30662 ( \31006 , \30684 , \30688 );
xor \U$30663 ( \31007 , \31006 , \30693 );
and \U$30664 ( \31008 , \31004 , \31007 );
and \U$30665 ( \31009 , \31002 , \31007 );
or \U$30666 ( \31010 , \31005 , \31008 , \31009 );
and \U$30667 ( \31011 , \31001 , \31010 );
xor \U$30668 ( \31012 , \30501 , \30505 );
xor \U$30669 ( \31013 , \31012 , \30510 );
xor \U$30670 ( \31014 , \30624 , \30628 );
xor \U$30671 ( \31015 , \31014 , \30633 );
and \U$30672 ( \31016 , \31013 , \31015 );
xor \U$30673 ( \31017 , \30641 , \30645 );
xor \U$30674 ( \31018 , \31017 , \30650 );
and \U$30675 ( \31019 , \31015 , \31018 );
and \U$30676 ( \31020 , \31013 , \31018 );
or \U$30677 ( \31021 , \31016 , \31019 , \31020 );
and \U$30678 ( \31022 , \31010 , \31021 );
and \U$30679 ( \31023 , \31001 , \31021 );
or \U$30680 ( \31024 , \31011 , \31022 , \31023 );
and \U$30681 ( \31025 , \30969 , \31024 );
xor \U$30682 ( \31026 , \30553 , \30557 );
xor \U$30683 ( \31027 , \31026 , \30562 );
xor \U$30684 ( \31028 , \30517 , \30521 );
xor \U$30685 ( \31029 , \31028 , \30526 );
and \U$30686 ( \31030 , \31027 , \31029 );
xor \U$30687 ( \31031 , \30534 , \30538 );
xor \U$30688 ( \31032 , \31031 , \30543 );
and \U$30689 ( \31033 , \31029 , \31032 );
and \U$30690 ( \31034 , \31027 , \31032 );
or \U$30691 ( \31035 , \31030 , \31033 , \31034 );
xor \U$30692 ( \31036 , \30569 , \30573 );
xor \U$30693 ( \31037 , \31036 , \30578 );
xor \U$30694 ( \31038 , \30588 , \30592 );
xor \U$30695 ( \31039 , \31038 , \30597 );
and \U$30696 ( \31040 , \31037 , \31039 );
and \U$30697 ( \31041 , \31035 , \31040 );
xor \U$30698 ( \31042 , \30709 , \30711 );
xor \U$30699 ( \31043 , \31042 , \30714 );
and \U$30700 ( \31044 , \31040 , \31043 );
and \U$30701 ( \31045 , \31035 , \31043 );
or \U$30702 ( \31046 , \31041 , \31044 , \31045 );
and \U$30703 ( \31047 , \31024 , \31046 );
and \U$30704 ( \31048 , \30969 , \31046 );
or \U$30705 ( \31049 , \31025 , \31047 , \31048 );
xor \U$30706 ( \31050 , \30513 , \30529 );
xor \U$30707 ( \31051 , \31050 , \30546 );
xor \U$30708 ( \31052 , \30565 , \30581 );
xor \U$30709 ( \31053 , \31052 , \30600 );
and \U$30710 ( \31054 , \31051 , \31053 );
xor \U$30711 ( \31055 , \30620 , \30636 );
xor \U$30712 ( \31056 , \31055 , \30653 );
and \U$30713 ( \31057 , \31053 , \31056 );
and \U$30714 ( \31058 , \31051 , \31056 );
or \U$30715 ( \31059 , \31054 , \31057 , \31058 );
xor \U$30716 ( \31060 , \30661 , \30663 );
xor \U$30717 ( \31061 , \31060 , \30666 );
xor \U$30718 ( \31062 , \30671 , \30673 );
xor \U$30719 ( \31063 , \31062 , \30676 );
and \U$30720 ( \31064 , \31061 , \31063 );
xor \U$30721 ( \31065 , \30696 , \30698 );
xor \U$30722 ( \31066 , \31065 , \30700 );
and \U$30723 ( \31067 , \31063 , \31066 );
and \U$30724 ( \31068 , \31061 , \31066 );
or \U$30725 ( \31069 , \31064 , \31067 , \31068 );
and \U$30726 ( \31070 , \31059 , \31069 );
xor \U$30727 ( \31071 , \30730 , \30732 );
xor \U$30728 ( \31072 , \31071 , \30735 );
and \U$30729 ( \31073 , \31069 , \31072 );
and \U$30730 ( \31074 , \31059 , \31072 );
or \U$30731 ( \31075 , \31070 , \31073 , \31074 );
and \U$30732 ( \31076 , \31049 , \31075 );
xor \U$30733 ( \31077 , \30669 , \30679 );
xor \U$30734 ( \31078 , \31077 , \30703 );
xor \U$30735 ( \31079 , \30740 , \30742 );
xor \U$30736 ( \31080 , \31079 , \30745 );
and \U$30737 ( \31081 , \31078 , \31080 );
xor \U$30738 ( \31082 , \30717 , \30719 );
xor \U$30739 ( \31083 , \31082 , \30722 );
and \U$30740 ( \31084 , \31080 , \31083 );
and \U$30741 ( \31085 , \31078 , \31083 );
or \U$30742 ( \31086 , \31081 , \31084 , \31085 );
and \U$30743 ( \31087 , \31075 , \31086 );
and \U$30744 ( \31088 , \31049 , \31086 );
or \U$30745 ( \31089 , \31076 , \31087 , \31088 );
xor \U$30746 ( \31090 , \30254 , \30309 );
xor \U$30747 ( \31091 , \31090 , \30362 );
xor \U$30748 ( \31092 , \30390 , \30400 );
xor \U$30749 ( \31093 , \31092 , \30411 );
and \U$30750 ( \31094 , \31091 , \31093 );
xor \U$30751 ( \31095 , \30757 , \30759 );
xor \U$30752 ( \31096 , \31095 , \30762 );
and \U$30753 ( \31097 , \31093 , \31096 );
and \U$30754 ( \31098 , \31091 , \31096 );
or \U$30755 ( \31099 , \31094 , \31097 , \31098 );
and \U$30756 ( \31100 , \31089 , \31099 );
xor \U$30757 ( \31101 , \30770 , \30772 );
xor \U$30758 ( \31102 , \31101 , \30775 );
and \U$30759 ( \31103 , \31099 , \31102 );
and \U$30760 ( \31104 , \31089 , \31102 );
or \U$30761 ( \31105 , \31100 , \31103 , \31104 );
xor \U$30762 ( \31106 , \30768 , \30778 );
xor \U$30763 ( \31107 , \31106 , \30781 );
and \U$30764 ( \31108 , \31105 , \31107 );
xor \U$30765 ( \31109 , \30786 , \30788 );
xor \U$30766 ( \31110 , \31109 , \30791 );
and \U$30767 ( \31111 , \31107 , \31110 );
and \U$30768 ( \31112 , \31105 , \31110 );
or \U$30769 ( \31113 , \31108 , \31111 , \31112 );
xor \U$30770 ( \31114 , \30784 , \30794 );
xor \U$30771 ( \31115 , \31114 , \30797 );
and \U$30772 ( \31116 , \31113 , \31115 );
xor \U$30773 ( \31117 , \30467 , \30477 );
xor \U$30774 ( \31118 , \31117 , \30480 );
and \U$30775 ( \31119 , \31115 , \31118 );
and \U$30776 ( \31120 , \31113 , \31118 );
or \U$30777 ( \31121 , \31116 , \31119 , \31120 );
and \U$30778 ( \31122 , \30806 , \31121 );
xor \U$30779 ( \31123 , \30806 , \31121 );
xor \U$30780 ( \31124 , \31113 , \31115 );
xor \U$30781 ( \31125 , \31124 , \31118 );
xor \U$30782 ( \31126 , \30934 , \30938 );
xor \U$30783 ( \31127 , \31126 , \30943 );
xor \U$30784 ( \31128 , \30951 , \30955 );
xor \U$30785 ( \31129 , \31128 , \30960 );
and \U$30786 ( \31130 , \31127 , \31129 );
xor \U$30787 ( \31131 , \30881 , \30885 );
xor \U$30788 ( \31132 , \31131 , \30890 );
and \U$30789 ( \31133 , \31129 , \31132 );
and \U$30790 ( \31134 , \31127 , \31132 );
or \U$30791 ( \31135 , \31130 , \31133 , \31134 );
xor \U$30792 ( \31136 , \30865 , \30869 );
xor \U$30793 ( \31137 , \31136 , \30874 );
xor \U$30794 ( \31138 , \30973 , \30977 );
xor \U$30795 ( \31139 , \31138 , \30982 );
and \U$30796 ( \31140 , \31137 , \31139 );
xor \U$30797 ( \31141 , \30898 , \30902 );
xor \U$30798 ( \31142 , \31141 , \30907 );
and \U$30799 ( \31143 , \31139 , \31142 );
and \U$30800 ( \31144 , \31137 , \31142 );
or \U$30801 ( \31145 , \31140 , \31143 , \31144 );
and \U$30802 ( \31146 , \31135 , \31145 );
and \U$30803 ( \31147 , \28952 , \21401 );
and \U$30804 ( \31148 , \28528 , \21399 );
nor \U$30805 ( \31149 , \31147 , \31148 );
xnor \U$30806 ( \31150 , \31149 , \21408 );
and \U$30807 ( \31151 , \29203 , \21419 );
and \U$30808 ( \31152 , \29198 , \21417 );
nor \U$30809 ( \31153 , \31151 , \31152 );
xnor \U$30810 ( \31154 , \31153 , \21426 );
and \U$30811 ( \31155 , \31150 , \31154 );
and \U$30812 ( \31156 , \29806 , \21434 );
and \U$30813 ( \31157 , \29522 , \21432 );
nor \U$30814 ( \31158 , \31156 , \31157 );
xnor \U$30815 ( \31159 , \31158 , \21441 );
and \U$30816 ( \31160 , \31154 , \31159 );
and \U$30817 ( \31161 , \31150 , \31159 );
or \U$30818 ( \31162 , \31155 , \31160 , \31161 );
and \U$30819 ( \31163 , \30383 , \21450 );
and \U$30820 ( \31164 , \30375 , \21448 );
nor \U$30821 ( \31165 , \31163 , \31164 );
xnor \U$30822 ( \31166 , \31165 , \21457 );
and \U$30823 ( \31167 , \30991 , \21469 );
and \U$30824 ( \31168 , \30986 , \21467 );
nor \U$30825 ( \31169 , \31167 , \31168 );
xnor \U$30826 ( \31170 , \31169 , \21476 );
and \U$30827 ( \31171 , \31166 , \31170 );
buf \U$30828 ( \31172 , RIbb33300_191);
and \U$30829 ( \31173 , \31172 , \21464 );
and \U$30830 ( \31174 , \31170 , \31173 );
and \U$30831 ( \31175 , \31166 , \31173 );
or \U$30832 ( \31176 , \31171 , \31174 , \31175 );
and \U$30833 ( \31177 , \31162 , \31176 );
xnor \U$30834 ( \31178 , \30990 , \30992 );
and \U$30835 ( \31179 , \31176 , \31178 );
and \U$30836 ( \31180 , \31162 , \31178 );
or \U$30837 ( \31181 , \31177 , \31179 , \31180 );
and \U$30838 ( \31182 , \31145 , \31181 );
and \U$30839 ( \31183 , \31135 , \31181 );
or \U$30840 ( \31184 , \31146 , \31182 , \31183 );
not \U$30841 ( \31185 , \30584 );
and \U$30842 ( \31186 , \21379 , \30826 );
and \U$30843 ( \31187 , \21387 , \30824 );
nor \U$30844 ( \31188 , \31186 , \31187 );
xnor \U$30845 ( \31189 , \31188 , \30587 );
and \U$30846 ( \31190 , \31185 , \31189 );
and \U$30847 ( \31191 , \21395 , \30258 );
and \U$30848 ( \31192 , \21403 , \30256 );
nor \U$30849 ( \31193 , \31191 , \31192 );
xnor \U$30850 ( \31194 , \31193 , \29948 );
and \U$30851 ( \31195 , \31189 , \31194 );
and \U$30852 ( \31196 , \31185 , \31194 );
or \U$30853 ( \31197 , \31190 , \31195 , \31196 );
and \U$30854 ( \31198 , \21413 , \29721 );
and \U$30855 ( \31199 , \21421 , \29719 );
nor \U$30856 ( \31200 , \31198 , \31199 );
xnor \U$30857 ( \31201 , \31200 , \29350 );
and \U$30858 ( \31202 , \21428 , \29159 );
and \U$30859 ( \31203 , \21436 , \29157 );
nor \U$30860 ( \31204 , \31202 , \31203 );
xnor \U$30861 ( \31205 , \31204 , \28841 );
and \U$30862 ( \31206 , \31201 , \31205 );
and \U$30863 ( \31207 , \21444 , \28592 );
and \U$30864 ( \31208 , \21452 , \28590 );
nor \U$30865 ( \31209 , \31207 , \31208 );
xnor \U$30866 ( \31210 , \31209 , \28343 );
and \U$30867 ( \31211 , \31205 , \31210 );
and \U$30868 ( \31212 , \31201 , \31210 );
or \U$30869 ( \31213 , \31206 , \31211 , \31212 );
and \U$30870 ( \31214 , \31197 , \31213 );
and \U$30871 ( \31215 , \21463 , \28063 );
and \U$30872 ( \31216 , \21471 , \28061 );
nor \U$30873 ( \31217 , \31215 , \31216 );
xnor \U$30874 ( \31218 , \31217 , \27803 );
and \U$30875 ( \31219 , \21689 , \27569 );
and \U$30876 ( \31220 , \21478 , \27567 );
nor \U$30877 ( \31221 , \31219 , \31220 );
xnor \U$30878 ( \31222 , \31221 , \27254 );
and \U$30879 ( \31223 , \31218 , \31222 );
and \U$30880 ( \31224 , \21813 , \27060 );
and \U$30881 ( \31225 , \21750 , \27058 );
nor \U$30882 ( \31226 , \31224 , \31225 );
xnor \U$30883 ( \31227 , \31226 , \26720 );
and \U$30884 ( \31228 , \31222 , \31227 );
and \U$30885 ( \31229 , \31218 , \31227 );
or \U$30886 ( \31230 , \31223 , \31228 , \31229 );
and \U$30887 ( \31231 , \31213 , \31230 );
and \U$30888 ( \31232 , \31197 , \31230 );
or \U$30889 ( \31233 , \31214 , \31231 , \31232 );
and \U$30890 ( \31234 , \25604 , \22379 );
and \U$30891 ( \31235 , \25596 , \22377 );
nor \U$30892 ( \31236 , \31234 , \31235 );
xnor \U$30893 ( \31237 , \31236 , \22266 );
and \U$30894 ( \31238 , \26078 , \22185 );
and \U$30895 ( \31239 , \26073 , \22183 );
nor \U$30896 ( \31240 , \31238 , \31239 );
xnor \U$30897 ( \31241 , \31240 , \22049 );
and \U$30898 ( \31242 , \31237 , \31241 );
and \U$30899 ( \31243 , \26601 , \21985 );
and \U$30900 ( \31244 , \26342 , \21983 );
nor \U$30901 ( \31245 , \31243 , \31244 );
xnor \U$30902 ( \31246 , \31245 , \21907 );
and \U$30903 ( \31247 , \31241 , \31246 );
and \U$30904 ( \31248 , \31237 , \31246 );
or \U$30905 ( \31249 , \31242 , \31247 , \31248 );
and \U$30906 ( \31250 , \24714 , \23125 );
and \U$30907 ( \31251 , \24506 , \23123 );
nor \U$30908 ( \31252 , \31250 , \31251 );
xnor \U$30909 ( \31253 , \31252 , \22988 );
and \U$30910 ( \31254 , \24841 , \22919 );
and \U$30911 ( \31255 , \24836 , \22917 );
nor \U$30912 ( \31256 , \31254 , \31255 );
xnor \U$30913 ( \31257 , \31256 , \22767 );
and \U$30914 ( \31258 , \31253 , \31257 );
and \U$30915 ( \31259 , \25294 , \22651 );
and \U$30916 ( \31260 , \25097 , \22649 );
nor \U$30917 ( \31261 , \31259 , \31260 );
xnor \U$30918 ( \31262 , \31261 , \22495 );
and \U$30919 ( \31263 , \31257 , \31262 );
and \U$30920 ( \31264 , \31253 , \31262 );
or \U$30921 ( \31265 , \31258 , \31263 , \31264 );
and \U$30922 ( \31266 , \31249 , \31265 );
and \U$30923 ( \31267 , \26982 , \21821 );
and \U$30924 ( \31268 , \26973 , \21819 );
nor \U$30925 ( \31269 , \31267 , \31268 );
xnor \U$30926 ( \31270 , \31269 , \21727 );
and \U$30927 ( \31271 , \27527 , \21652 );
and \U$30928 ( \31272 , \27325 , \21650 );
nor \U$30929 ( \31273 , \31271 , \31272 );
xnor \U$30930 ( \31274 , \31273 , \21377 );
and \U$30931 ( \31275 , \31270 , \31274 );
and \U$30932 ( \31276 , \28002 , \21385 );
and \U$30933 ( \31277 , \27830 , \21383 );
nor \U$30934 ( \31278 , \31276 , \31277 );
xnor \U$30935 ( \31279 , \31278 , \21392 );
and \U$30936 ( \31280 , \31274 , \31279 );
and \U$30937 ( \31281 , \31270 , \31279 );
or \U$30938 ( \31282 , \31275 , \31280 , \31281 );
and \U$30939 ( \31283 , \31265 , \31282 );
and \U$30940 ( \31284 , \31249 , \31282 );
or \U$30941 ( \31285 , \31266 , \31283 , \31284 );
and \U$30942 ( \31286 , \31233 , \31285 );
and \U$30943 ( \31287 , \22624 , \25180 );
and \U$30944 ( \31288 , \22616 , \25178 );
nor \U$30945 ( \31289 , \31287 , \31288 );
xnor \U$30946 ( \31290 , \31289 , \25037 );
and \U$30947 ( \31291 , \22872 , \24857 );
and \U$30948 ( \31292 , \22867 , \24855 );
nor \U$30949 ( \31293 , \31291 , \31292 );
xnor \U$30950 ( \31294 , \31293 , \24611 );
and \U$30951 ( \31295 , \31290 , \31294 );
and \U$30952 ( \31296 , \23202 , \24462 );
and \U$30953 ( \31297 , \23058 , \24460 );
nor \U$30954 ( \31298 , \31296 , \31297 );
xnor \U$30955 ( \31299 , \31298 , \24275 );
and \U$30956 ( \31300 , \31294 , \31299 );
and \U$30957 ( \31301 , \31290 , \31299 );
or \U$30958 ( \31302 , \31295 , \31300 , \31301 );
and \U$30959 ( \31303 , \23491 , \24149 );
and \U$30960 ( \31304 , \23466 , \24147 );
nor \U$30961 ( \31305 , \31303 , \31304 );
xnor \U$30962 ( \31306 , \31305 , \23944 );
and \U$30963 ( \31307 , \23832 , \23743 );
and \U$30964 ( \31308 , \23665 , \23741 );
nor \U$30965 ( \31309 , \31307 , \31308 );
xnor \U$30966 ( \31310 , \31309 , \23594 );
and \U$30967 ( \31311 , \31306 , \31310 );
and \U$30968 ( \31312 , \24089 , \23421 );
and \U$30969 ( \31313 , \23970 , \23419 );
nor \U$30970 ( \31314 , \31312 , \31313 );
xnor \U$30971 ( \31315 , \31314 , \23279 );
and \U$30972 ( \31316 , \31310 , \31315 );
and \U$30973 ( \31317 , \31306 , \31315 );
or \U$30974 ( \31318 , \31311 , \31316 , \31317 );
and \U$30975 ( \31319 , \31302 , \31318 );
and \U$30976 ( \31320 , \22099 , \26471 );
and \U$30977 ( \31321 , \22011 , \26469 );
nor \U$30978 ( \31322 , \31320 , \31321 );
xnor \U$30979 ( \31323 , \31322 , \26230 );
and \U$30980 ( \31324 , \22209 , \26005 );
and \U$30981 ( \31325 , \22204 , \26003 );
nor \U$30982 ( \31326 , \31324 , \31325 );
xnor \U$30983 ( \31327 , \31326 , \25817 );
and \U$30984 ( \31328 , \31323 , \31327 );
and \U$30985 ( \31329 , \22440 , \25631 );
and \U$30986 ( \31330 , \22325 , \25629 );
nor \U$30987 ( \31331 , \31329 , \31330 );
xnor \U$30988 ( \31332 , \31331 , \25399 );
and \U$30989 ( \31333 , \31327 , \31332 );
and \U$30990 ( \31334 , \31323 , \31332 );
or \U$30991 ( \31335 , \31328 , \31333 , \31334 );
and \U$30992 ( \31336 , \31318 , \31335 );
and \U$30993 ( \31337 , \31302 , \31335 );
or \U$30994 ( \31338 , \31319 , \31336 , \31337 );
and \U$30995 ( \31339 , \31285 , \31338 );
and \U$30996 ( \31340 , \31233 , \31338 );
or \U$30997 ( \31341 , \31286 , \31339 , \31340 );
and \U$30998 ( \31342 , \31184 , \31341 );
xor \U$30999 ( \31343 , \30918 , \30922 );
xor \U$31000 ( \31344 , \31343 , \30927 );
xor \U$31001 ( \31345 , \30810 , \30814 );
xor \U$31002 ( \31346 , \31345 , \30819 );
and \U$31003 ( \31347 , \31344 , \31346 );
xor \U$31004 ( \31348 , \30846 , \30850 );
xor \U$31005 ( \31349 , \31348 , \30855 );
and \U$31006 ( \31350 , \31346 , \31349 );
and \U$31007 ( \31351 , \31344 , \31349 );
or \U$31008 ( \31352 , \31347 , \31350 , \31351 );
xor \U$31009 ( \31353 , \31027 , \31029 );
xor \U$31010 ( \31354 , \31353 , \31032 );
and \U$31011 ( \31355 , \31352 , \31354 );
xor \U$31012 ( \31356 , \31037 , \31039 );
and \U$31013 ( \31357 , \31354 , \31356 );
and \U$31014 ( \31358 , \31352 , \31356 );
or \U$31015 ( \31359 , \31355 , \31357 , \31358 );
and \U$31016 ( \31360 , \31341 , \31359 );
and \U$31017 ( \31361 , \31184 , \31359 );
or \U$31018 ( \31362 , \31342 , \31360 , \31361 );
xor \U$31019 ( \31363 , \30822 , \30841 );
xor \U$31020 ( \31364 , \31363 , \30858 );
xor \U$31021 ( \31365 , \30877 , \30893 );
xor \U$31022 ( \31366 , \31365 , \30910 );
and \U$31023 ( \31367 , \31364 , \31366 );
xor \U$31024 ( \31368 , \30930 , \30946 );
xor \U$31025 ( \31369 , \31368 , \30963 );
and \U$31026 ( \31370 , \31366 , \31369 );
and \U$31027 ( \31371 , \31364 , \31369 );
or \U$31028 ( \31372 , \31367 , \31370 , \31371 );
xor \U$31029 ( \31373 , \30985 , \30993 );
xor \U$31030 ( \31374 , \31373 , \30998 );
xor \U$31031 ( \31375 , \31002 , \31004 );
xor \U$31032 ( \31376 , \31375 , \31007 );
and \U$31033 ( \31377 , \31374 , \31376 );
xor \U$31034 ( \31378 , \31013 , \31015 );
xor \U$31035 ( \31379 , \31378 , \31018 );
and \U$31036 ( \31380 , \31376 , \31379 );
and \U$31037 ( \31381 , \31374 , \31379 );
or \U$31038 ( \31382 , \31377 , \31380 , \31381 );
and \U$31039 ( \31383 , \31372 , \31382 );
xor \U$31040 ( \31384 , \31051 , \31053 );
xor \U$31041 ( \31385 , \31384 , \31056 );
and \U$31042 ( \31386 , \31382 , \31385 );
and \U$31043 ( \31387 , \31372 , \31385 );
or \U$31044 ( \31388 , \31383 , \31386 , \31387 );
and \U$31045 ( \31389 , \31362 , \31388 );
xor \U$31046 ( \31390 , \31001 , \31010 );
xor \U$31047 ( \31391 , \31390 , \31021 );
xor \U$31048 ( \31392 , \31035 , \31040 );
xor \U$31049 ( \31393 , \31392 , \31043 );
and \U$31050 ( \31394 , \31391 , \31393 );
xor \U$31051 ( \31395 , \31061 , \31063 );
xor \U$31052 ( \31396 , \31395 , \31066 );
and \U$31053 ( \31397 , \31393 , \31396 );
and \U$31054 ( \31398 , \31391 , \31396 );
or \U$31055 ( \31399 , \31394 , \31397 , \31398 );
and \U$31056 ( \31400 , \31388 , \31399 );
and \U$31057 ( \31401 , \31362 , \31399 );
or \U$31058 ( \31402 , \31389 , \31400 , \31401 );
xor \U$31059 ( \31403 , \30549 , \30603 );
xor \U$31060 ( \31404 , \31403 , \30656 );
xor \U$31061 ( \31405 , \31059 , \31069 );
xor \U$31062 ( \31406 , \31405 , \31072 );
and \U$31063 ( \31407 , \31404 , \31406 );
xor \U$31064 ( \31408 , \31078 , \31080 );
xor \U$31065 ( \31409 , \31408 , \31083 );
and \U$31066 ( \31410 , \31406 , \31409 );
and \U$31067 ( \31411 , \31404 , \31409 );
or \U$31068 ( \31412 , \31407 , \31410 , \31411 );
and \U$31069 ( \31413 , \31402 , \31412 );
xor \U$31070 ( \31414 , \30738 , \30748 );
xor \U$31071 ( \31415 , \31414 , \30751 );
and \U$31072 ( \31416 , \31412 , \31415 );
and \U$31073 ( \31417 , \31402 , \31415 );
or \U$31074 ( \31418 , \31413 , \31416 , \31417 );
xor \U$31075 ( \31419 , \30659 , \30706 );
xor \U$31076 ( \31420 , \31419 , \30725 );
xor \U$31077 ( \31421 , \31049 , \31075 );
xor \U$31078 ( \31422 , \31421 , \31086 );
and \U$31079 ( \31423 , \31420 , \31422 );
xor \U$31080 ( \31424 , \31091 , \31093 );
xor \U$31081 ( \31425 , \31424 , \31096 );
and \U$31082 ( \31426 , \31422 , \31425 );
and \U$31083 ( \31427 , \31420 , \31425 );
or \U$31084 ( \31428 , \31423 , \31426 , \31427 );
and \U$31085 ( \31429 , \31418 , \31428 );
xor \U$31086 ( \31430 , \30728 , \30754 );
xor \U$31087 ( \31431 , \31430 , \30765 );
and \U$31088 ( \31432 , \31428 , \31431 );
and \U$31089 ( \31433 , \31418 , \31431 );
or \U$31090 ( \31434 , \31429 , \31432 , \31433 );
xor \U$31091 ( \31435 , \31105 , \31107 );
xor \U$31092 ( \31436 , \31435 , \31110 );
and \U$31093 ( \31437 , \31434 , \31436 );
and \U$31094 ( \31438 , \31125 , \31437 );
xor \U$31095 ( \31439 , \31125 , \31437 );
xor \U$31096 ( \31440 , \31434 , \31436 );
xor \U$31097 ( \31441 , \31237 , \31241 );
xor \U$31098 ( \31442 , \31441 , \31246 );
xor \U$31099 ( \31443 , \31253 , \31257 );
xor \U$31100 ( \31444 , \31443 , \31262 );
and \U$31101 ( \31445 , \31442 , \31444 );
xor \U$31102 ( \31446 , \31306 , \31310 );
xor \U$31103 ( \31447 , \31446 , \31315 );
and \U$31104 ( \31448 , \31444 , \31447 );
and \U$31105 ( \31449 , \31442 , \31447 );
or \U$31106 ( \31450 , \31445 , \31448 , \31449 );
xor \U$31107 ( \31451 , \31150 , \31154 );
xor \U$31108 ( \31452 , \31451 , \31159 );
xor \U$31109 ( \31453 , \31166 , \31170 );
xor \U$31110 ( \31454 , \31453 , \31173 );
and \U$31111 ( \31455 , \31452 , \31454 );
xor \U$31112 ( \31456 , \31270 , \31274 );
xor \U$31113 ( \31457 , \31456 , \31279 );
and \U$31114 ( \31458 , \31454 , \31457 );
and \U$31115 ( \31459 , \31452 , \31457 );
or \U$31116 ( \31460 , \31455 , \31458 , \31459 );
and \U$31117 ( \31461 , \31450 , \31460 );
and \U$31118 ( \31462 , \28528 , \21385 );
and \U$31119 ( \31463 , \28002 , \21383 );
nor \U$31120 ( \31464 , \31462 , \31463 );
xnor \U$31121 ( \31465 , \31464 , \21392 );
and \U$31122 ( \31466 , \29198 , \21401 );
and \U$31123 ( \31467 , \28952 , \21399 );
nor \U$31124 ( \31468 , \31466 , \31467 );
xnor \U$31125 ( \31469 , \31468 , \21408 );
and \U$31126 ( \31470 , \31465 , \31469 );
and \U$31127 ( \31471 , \29522 , \21419 );
and \U$31128 ( \31472 , \29203 , \21417 );
nor \U$31129 ( \31473 , \31471 , \31472 );
xnor \U$31130 ( \31474 , \31473 , \21426 );
and \U$31131 ( \31475 , \31469 , \31474 );
and \U$31132 ( \31476 , \31465 , \31474 );
or \U$31133 ( \31477 , \31470 , \31475 , \31476 );
and \U$31134 ( \31478 , \30375 , \21434 );
and \U$31135 ( \31479 , \29806 , \21432 );
nor \U$31136 ( \31480 , \31478 , \31479 );
xnor \U$31137 ( \31481 , \31480 , \21441 );
and \U$31138 ( \31482 , \30986 , \21450 );
and \U$31139 ( \31483 , \30383 , \21448 );
nor \U$31140 ( \31484 , \31482 , \31483 );
xnor \U$31141 ( \31485 , \31484 , \21457 );
and \U$31142 ( \31486 , \31481 , \31485 );
and \U$31143 ( \31487 , \31172 , \21469 );
and \U$31144 ( \31488 , \30991 , \21467 );
nor \U$31145 ( \31489 , \31487 , \31488 );
xnor \U$31146 ( \31490 , \31489 , \21476 );
and \U$31147 ( \31491 , \31485 , \31490 );
and \U$31148 ( \31492 , \31481 , \31490 );
or \U$31149 ( \31493 , \31486 , \31491 , \31492 );
or \U$31150 ( \31494 , \31477 , \31493 );
and \U$31151 ( \31495 , \31460 , \31494 );
and \U$31152 ( \31496 , \31450 , \31494 );
or \U$31153 ( \31497 , \31461 , \31495 , \31496 );
and \U$31154 ( \31498 , \25596 , \22651 );
and \U$31155 ( \31499 , \25294 , \22649 );
nor \U$31156 ( \31500 , \31498 , \31499 );
xnor \U$31157 ( \31501 , \31500 , \22495 );
and \U$31158 ( \31502 , \26073 , \22379 );
and \U$31159 ( \31503 , \25604 , \22377 );
nor \U$31160 ( \31504 , \31502 , \31503 );
xnor \U$31161 ( \31505 , \31504 , \22266 );
and \U$31162 ( \31506 , \31501 , \31505 );
and \U$31163 ( \31507 , \26342 , \22185 );
and \U$31164 ( \31508 , \26078 , \22183 );
nor \U$31165 ( \31509 , \31507 , \31508 );
xnor \U$31166 ( \31510 , \31509 , \22049 );
and \U$31167 ( \31511 , \31505 , \31510 );
and \U$31168 ( \31512 , \31501 , \31510 );
or \U$31169 ( \31513 , \31506 , \31511 , \31512 );
and \U$31170 ( \31514 , \26973 , \21985 );
and \U$31171 ( \31515 , \26601 , \21983 );
nor \U$31172 ( \31516 , \31514 , \31515 );
xnor \U$31173 ( \31517 , \31516 , \21907 );
and \U$31174 ( \31518 , \27325 , \21821 );
and \U$31175 ( \31519 , \26982 , \21819 );
nor \U$31176 ( \31520 , \31518 , \31519 );
xnor \U$31177 ( \31521 , \31520 , \21727 );
and \U$31178 ( \31522 , \31517 , \31521 );
and \U$31179 ( \31523 , \27830 , \21652 );
and \U$31180 ( \31524 , \27527 , \21650 );
nor \U$31181 ( \31525 , \31523 , \31524 );
xnor \U$31182 ( \31526 , \31525 , \21377 );
and \U$31183 ( \31527 , \31521 , \31526 );
and \U$31184 ( \31528 , \31517 , \31526 );
or \U$31185 ( \31529 , \31522 , \31527 , \31528 );
and \U$31186 ( \31530 , \31513 , \31529 );
and \U$31187 ( \31531 , \24506 , \23421 );
and \U$31188 ( \31532 , \24089 , \23419 );
nor \U$31189 ( \31533 , \31531 , \31532 );
xnor \U$31190 ( \31534 , \31533 , \23279 );
and \U$31191 ( \31535 , \24836 , \23125 );
and \U$31192 ( \31536 , \24714 , \23123 );
nor \U$31193 ( \31537 , \31535 , \31536 );
xnor \U$31194 ( \31538 , \31537 , \22988 );
and \U$31195 ( \31539 , \31534 , \31538 );
and \U$31196 ( \31540 , \25097 , \22919 );
and \U$31197 ( \31541 , \24841 , \22917 );
nor \U$31198 ( \31542 , \31540 , \31541 );
xnor \U$31199 ( \31543 , \31542 , \22767 );
and \U$31200 ( \31544 , \31538 , \31543 );
and \U$31201 ( \31545 , \31534 , \31543 );
or \U$31202 ( \31546 , \31539 , \31544 , \31545 );
and \U$31203 ( \31547 , \31529 , \31546 );
and \U$31204 ( \31548 , \31513 , \31546 );
or \U$31205 ( \31549 , \31530 , \31547 , \31548 );
and \U$31206 ( \31550 , \22616 , \25631 );
and \U$31207 ( \31551 , \22440 , \25629 );
nor \U$31208 ( \31552 , \31550 , \31551 );
xnor \U$31209 ( \31553 , \31552 , \25399 );
and \U$31210 ( \31554 , \22867 , \25180 );
and \U$31211 ( \31555 , \22624 , \25178 );
nor \U$31212 ( \31556 , \31554 , \31555 );
xnor \U$31213 ( \31557 , \31556 , \25037 );
and \U$31214 ( \31558 , \31553 , \31557 );
and \U$31215 ( \31559 , \23058 , \24857 );
and \U$31216 ( \31560 , \22872 , \24855 );
nor \U$31217 ( \31561 , \31559 , \31560 );
xnor \U$31218 ( \31562 , \31561 , \24611 );
and \U$31219 ( \31563 , \31557 , \31562 );
and \U$31220 ( \31564 , \31553 , \31562 );
or \U$31221 ( \31565 , \31558 , \31563 , \31564 );
and \U$31222 ( \31566 , \23466 , \24462 );
and \U$31223 ( \31567 , \23202 , \24460 );
nor \U$31224 ( \31568 , \31566 , \31567 );
xnor \U$31225 ( \31569 , \31568 , \24275 );
and \U$31226 ( \31570 , \23665 , \24149 );
and \U$31227 ( \31571 , \23491 , \24147 );
nor \U$31228 ( \31572 , \31570 , \31571 );
xnor \U$31229 ( \31573 , \31572 , \23944 );
and \U$31230 ( \31574 , \31569 , \31573 );
and \U$31231 ( \31575 , \23970 , \23743 );
and \U$31232 ( \31576 , \23832 , \23741 );
nor \U$31233 ( \31577 , \31575 , \31576 );
xnor \U$31234 ( \31578 , \31577 , \23594 );
and \U$31235 ( \31579 , \31573 , \31578 );
and \U$31236 ( \31580 , \31569 , \31578 );
or \U$31237 ( \31581 , \31574 , \31579 , \31580 );
and \U$31238 ( \31582 , \31565 , \31581 );
and \U$31239 ( \31583 , \22011 , \27060 );
and \U$31240 ( \31584 , \21813 , \27058 );
nor \U$31241 ( \31585 , \31583 , \31584 );
xnor \U$31242 ( \31586 , \31585 , \26720 );
and \U$31243 ( \31587 , \22204 , \26471 );
and \U$31244 ( \31588 , \22099 , \26469 );
nor \U$31245 ( \31589 , \31587 , \31588 );
xnor \U$31246 ( \31590 , \31589 , \26230 );
and \U$31247 ( \31591 , \31586 , \31590 );
and \U$31248 ( \31592 , \22325 , \26005 );
and \U$31249 ( \31593 , \22209 , \26003 );
nor \U$31250 ( \31594 , \31592 , \31593 );
xnor \U$31251 ( \31595 , \31594 , \25817 );
and \U$31252 ( \31596 , \31590 , \31595 );
and \U$31253 ( \31597 , \31586 , \31595 );
or \U$31254 ( \31598 , \31591 , \31596 , \31597 );
and \U$31255 ( \31599 , \31581 , \31598 );
and \U$31256 ( \31600 , \31565 , \31598 );
or \U$31257 ( \31601 , \31582 , \31599 , \31600 );
and \U$31258 ( \31602 , \31549 , \31601 );
and \U$31259 ( \31603 , \21421 , \30258 );
and \U$31260 ( \31604 , \21395 , \30256 );
nor \U$31261 ( \31605 , \31603 , \31604 );
xnor \U$31262 ( \31606 , \31605 , \29948 );
and \U$31263 ( \31607 , \21436 , \29721 );
and \U$31264 ( \31608 , \21413 , \29719 );
nor \U$31265 ( \31609 , \31607 , \31608 );
xnor \U$31266 ( \31610 , \31609 , \29350 );
and \U$31267 ( \31611 , \31606 , \31610 );
and \U$31268 ( \31612 , \21452 , \29159 );
and \U$31269 ( \31613 , \21428 , \29157 );
nor \U$31270 ( \31614 , \31612 , \31613 );
xnor \U$31271 ( \31615 , \31614 , \28841 );
and \U$31272 ( \31616 , \31610 , \31615 );
and \U$31273 ( \31617 , \31606 , \31615 );
or \U$31274 ( \31618 , \31611 , \31616 , \31617 );
and \U$31275 ( \31619 , \21471 , \28592 );
and \U$31276 ( \31620 , \21444 , \28590 );
nor \U$31277 ( \31621 , \31619 , \31620 );
xnor \U$31278 ( \31622 , \31621 , \28343 );
and \U$31279 ( \31623 , \21478 , \28063 );
and \U$31280 ( \31624 , \21463 , \28061 );
nor \U$31281 ( \31625 , \31623 , \31624 );
xnor \U$31282 ( \31626 , \31625 , \27803 );
and \U$31283 ( \31627 , \31622 , \31626 );
and \U$31284 ( \31628 , \21750 , \27569 );
and \U$31285 ( \31629 , \21689 , \27567 );
nor \U$31286 ( \31630 , \31628 , \31629 );
xnor \U$31287 ( \31631 , \31630 , \27254 );
and \U$31288 ( \31632 , \31626 , \31631 );
and \U$31289 ( \31633 , \31622 , \31631 );
or \U$31290 ( \31634 , \31627 , \31632 , \31633 );
and \U$31291 ( \31635 , \31618 , \31634 );
buf \U$31292 ( \31636 , RIbb2d888_64);
xor \U$31293 ( \31637 , \30584 , \31636 );
not \U$31294 ( \31638 , \31636 );
and \U$31295 ( \31639 , \31637 , \31638 );
and \U$31296 ( \31640 , \21387 , \31639 );
not \U$31297 ( \31641 , \31640 );
xnor \U$31298 ( \31642 , \31641 , \30584 );
and \U$31299 ( \31643 , \21403 , \30826 );
and \U$31300 ( \31644 , \21379 , \30824 );
nor \U$31301 ( \31645 , \31643 , \31644 );
xnor \U$31302 ( \31646 , \31645 , \30587 );
and \U$31303 ( \31647 , \31642 , \31646 );
and \U$31304 ( \31648 , \31634 , \31647 );
and \U$31305 ( \31649 , \31618 , \31647 );
or \U$31306 ( \31650 , \31635 , \31648 , \31649 );
and \U$31307 ( \31651 , \31601 , \31650 );
and \U$31308 ( \31652 , \31549 , \31650 );
or \U$31309 ( \31653 , \31602 , \31651 , \31652 );
and \U$31310 ( \31654 , \31497 , \31653 );
xor \U$31311 ( \31655 , \31290 , \31294 );
xor \U$31312 ( \31656 , \31655 , \31299 );
xor \U$31313 ( \31657 , \31218 , \31222 );
xor \U$31314 ( \31658 , \31657 , \31227 );
and \U$31315 ( \31659 , \31656 , \31658 );
xor \U$31316 ( \31660 , \31323 , \31327 );
xor \U$31317 ( \31661 , \31660 , \31332 );
and \U$31318 ( \31662 , \31658 , \31661 );
and \U$31319 ( \31663 , \31656 , \31661 );
or \U$31320 ( \31664 , \31659 , \31662 , \31663 );
xor \U$31321 ( \31665 , \31185 , \31189 );
xor \U$31322 ( \31666 , \31665 , \31194 );
xor \U$31323 ( \31667 , \31201 , \31205 );
xor \U$31324 ( \31668 , \31667 , \31210 );
and \U$31325 ( \31669 , \31666 , \31668 );
and \U$31326 ( \31670 , \31664 , \31669 );
xor \U$31327 ( \31671 , \30829 , \30833 );
xor \U$31328 ( \31672 , \31671 , \30838 );
and \U$31329 ( \31673 , \31669 , \31672 );
and \U$31330 ( \31674 , \31664 , \31672 );
or \U$31331 ( \31675 , \31670 , \31673 , \31674 );
and \U$31332 ( \31676 , \31653 , \31675 );
and \U$31333 ( \31677 , \31497 , \31675 );
or \U$31334 ( \31678 , \31654 , \31676 , \31677 );
xor \U$31335 ( \31679 , \31344 , \31346 );
xor \U$31336 ( \31680 , \31679 , \31349 );
xor \U$31337 ( \31681 , \31127 , \31129 );
xor \U$31338 ( \31682 , \31681 , \31132 );
and \U$31339 ( \31683 , \31680 , \31682 );
xor \U$31340 ( \31684 , \31137 , \31139 );
xor \U$31341 ( \31685 , \31684 , \31142 );
and \U$31342 ( \31686 , \31682 , \31685 );
and \U$31343 ( \31687 , \31680 , \31685 );
or \U$31344 ( \31688 , \31683 , \31686 , \31687 );
xor \U$31345 ( \31689 , \31249 , \31265 );
xor \U$31346 ( \31690 , \31689 , \31282 );
xor \U$31347 ( \31691 , \31302 , \31318 );
xor \U$31348 ( \31692 , \31691 , \31335 );
and \U$31349 ( \31693 , \31690 , \31692 );
xor \U$31350 ( \31694 , \31162 , \31176 );
xor \U$31351 ( \31695 , \31694 , \31178 );
and \U$31352 ( \31696 , \31692 , \31695 );
and \U$31353 ( \31697 , \31690 , \31695 );
or \U$31354 ( \31698 , \31693 , \31696 , \31697 );
and \U$31355 ( \31699 , \31688 , \31698 );
xor \U$31356 ( \31700 , \31364 , \31366 );
xor \U$31357 ( \31701 , \31700 , \31369 );
and \U$31358 ( \31702 , \31698 , \31701 );
and \U$31359 ( \31703 , \31688 , \31701 );
or \U$31360 ( \31704 , \31699 , \31702 , \31703 );
and \U$31361 ( \31705 , \31678 , \31704 );
xor \U$31362 ( \31706 , \31135 , \31145 );
xor \U$31363 ( \31707 , \31706 , \31181 );
xor \U$31364 ( \31708 , \31374 , \31376 );
xor \U$31365 ( \31709 , \31708 , \31379 );
and \U$31366 ( \31710 , \31707 , \31709 );
xor \U$31367 ( \31711 , \31352 , \31354 );
xor \U$31368 ( \31712 , \31711 , \31356 );
and \U$31369 ( \31713 , \31709 , \31712 );
and \U$31370 ( \31714 , \31707 , \31712 );
or \U$31371 ( \31715 , \31710 , \31713 , \31714 );
and \U$31372 ( \31716 , \31704 , \31715 );
and \U$31373 ( \31717 , \31678 , \31715 );
or \U$31374 ( \31718 , \31705 , \31716 , \31717 );
xor \U$31375 ( \31719 , \30861 , \30913 );
xor \U$31376 ( \31720 , \31719 , \30966 );
xor \U$31377 ( \31721 , \31372 , \31382 );
xor \U$31378 ( \31722 , \31721 , \31385 );
and \U$31379 ( \31723 , \31720 , \31722 );
xor \U$31380 ( \31724 , \31391 , \31393 );
xor \U$31381 ( \31725 , \31724 , \31396 );
and \U$31382 ( \31726 , \31722 , \31725 );
and \U$31383 ( \31727 , \31720 , \31725 );
or \U$31384 ( \31728 , \31723 , \31726 , \31727 );
and \U$31385 ( \31729 , \31718 , \31728 );
xor \U$31386 ( \31730 , \30969 , \31024 );
xor \U$31387 ( \31731 , \31730 , \31046 );
and \U$31388 ( \31732 , \31728 , \31731 );
and \U$31389 ( \31733 , \31718 , \31731 );
or \U$31390 ( \31734 , \31729 , \31732 , \31733 );
xor \U$31391 ( \31735 , \31402 , \31412 );
xor \U$31392 ( \31736 , \31735 , \31415 );
and \U$31393 ( \31737 , \31734 , \31736 );
xor \U$31394 ( \31738 , \31420 , \31422 );
xor \U$31395 ( \31739 , \31738 , \31425 );
and \U$31396 ( \31740 , \31736 , \31739 );
and \U$31397 ( \31741 , \31734 , \31739 );
or \U$31398 ( \31742 , \31737 , \31740 , \31741 );
xor \U$31399 ( \31743 , \31418 , \31428 );
xor \U$31400 ( \31744 , \31743 , \31431 );
and \U$31401 ( \31745 , \31742 , \31744 );
xor \U$31402 ( \31746 , \31089 , \31099 );
xor \U$31403 ( \31747 , \31746 , \31102 );
and \U$31404 ( \31748 , \31744 , \31747 );
and \U$31405 ( \31749 , \31742 , \31747 );
or \U$31406 ( \31750 , \31745 , \31748 , \31749 );
and \U$31407 ( \31751 , \31440 , \31750 );
xor \U$31408 ( \31752 , \31440 , \31750 );
xor \U$31409 ( \31753 , \31742 , \31744 );
xor \U$31410 ( \31754 , \31753 , \31747 );
xor \U$31411 ( \31755 , \31501 , \31505 );
xor \U$31412 ( \31756 , \31755 , \31510 );
xor \U$31413 ( \31757 , \31465 , \31469 );
xor \U$31414 ( \31758 , \31757 , \31474 );
and \U$31415 ( \31759 , \31756 , \31758 );
xor \U$31416 ( \31760 , \31517 , \31521 );
xor \U$31417 ( \31761 , \31760 , \31526 );
and \U$31418 ( \31762 , \31758 , \31761 );
and \U$31419 ( \31763 , \31756 , \31761 );
or \U$31420 ( \31764 , \31759 , \31762 , \31763 );
xor \U$31421 ( \31765 , \31553 , \31557 );
xor \U$31422 ( \31766 , \31765 , \31562 );
xor \U$31423 ( \31767 , \31569 , \31573 );
xor \U$31424 ( \31768 , \31767 , \31578 );
and \U$31425 ( \31769 , \31766 , \31768 );
xor \U$31426 ( \31770 , \31534 , \31538 );
xor \U$31427 ( \31771 , \31770 , \31543 );
and \U$31428 ( \31772 , \31768 , \31771 );
and \U$31429 ( \31773 , \31766 , \31771 );
or \U$31430 ( \31774 , \31769 , \31772 , \31773 );
and \U$31431 ( \31775 , \31764 , \31774 );
and \U$31432 ( \31776 , \29203 , \21401 );
and \U$31433 ( \31777 , \29198 , \21399 );
nor \U$31434 ( \31778 , \31776 , \31777 );
xnor \U$31435 ( \31779 , \31778 , \21408 );
and \U$31436 ( \31780 , \29806 , \21419 );
and \U$31437 ( \31781 , \29522 , \21417 );
nor \U$31438 ( \31782 , \31780 , \31781 );
xnor \U$31439 ( \31783 , \31782 , \21426 );
and \U$31440 ( \31784 , \31779 , \31783 );
and \U$31441 ( \31785 , \30383 , \21434 );
and \U$31442 ( \31786 , \30375 , \21432 );
nor \U$31443 ( \31787 , \31785 , \31786 );
xnor \U$31444 ( \31788 , \31787 , \21441 );
and \U$31445 ( \31789 , \31783 , \31788 );
and \U$31446 ( \31790 , \31779 , \31788 );
or \U$31447 ( \31791 , \31784 , \31789 , \31790 );
buf \U$31448 ( \31792 , RIbb33378_192);
nand \U$31449 ( \31793 , \31792 , \21464 );
not \U$31450 ( \31794 , \31793 );
and \U$31451 ( \31795 , \31791 , \31794 );
xor \U$31452 ( \31796 , \31481 , \31485 );
xor \U$31453 ( \31797 , \31796 , \31490 );
and \U$31454 ( \31798 , \31794 , \31797 );
and \U$31455 ( \31799 , \31791 , \31797 );
or \U$31456 ( \31800 , \31795 , \31798 , \31799 );
and \U$31457 ( \31801 , \31774 , \31800 );
and \U$31458 ( \31802 , \31764 , \31800 );
or \U$31459 ( \31803 , \31775 , \31801 , \31802 );
and \U$31460 ( \31804 , \22872 , \25180 );
and \U$31461 ( \31805 , \22867 , \25178 );
nor \U$31462 ( \31806 , \31804 , \31805 );
xnor \U$31463 ( \31807 , \31806 , \25037 );
and \U$31464 ( \31808 , \23202 , \24857 );
and \U$31465 ( \31809 , \23058 , \24855 );
nor \U$31466 ( \31810 , \31808 , \31809 );
xnor \U$31467 ( \31811 , \31810 , \24611 );
and \U$31468 ( \31812 , \31807 , \31811 );
and \U$31469 ( \31813 , \23491 , \24462 );
and \U$31470 ( \31814 , \23466 , \24460 );
nor \U$31471 ( \31815 , \31813 , \31814 );
xnor \U$31472 ( \31816 , \31815 , \24275 );
and \U$31473 ( \31817 , \31811 , \31816 );
and \U$31474 ( \31818 , \31807 , \31816 );
or \U$31475 ( \31819 , \31812 , \31817 , \31818 );
and \U$31476 ( \31820 , \22209 , \26471 );
and \U$31477 ( \31821 , \22204 , \26469 );
nor \U$31478 ( \31822 , \31820 , \31821 );
xnor \U$31479 ( \31823 , \31822 , \26230 );
and \U$31480 ( \31824 , \22440 , \26005 );
and \U$31481 ( \31825 , \22325 , \26003 );
nor \U$31482 ( \31826 , \31824 , \31825 );
xnor \U$31483 ( \31827 , \31826 , \25817 );
and \U$31484 ( \31828 , \31823 , \31827 );
and \U$31485 ( \31829 , \22624 , \25631 );
and \U$31486 ( \31830 , \22616 , \25629 );
nor \U$31487 ( \31831 , \31829 , \31830 );
xnor \U$31488 ( \31832 , \31831 , \25399 );
and \U$31489 ( \31833 , \31827 , \31832 );
and \U$31490 ( \31834 , \31823 , \31832 );
or \U$31491 ( \31835 , \31828 , \31833 , \31834 );
and \U$31492 ( \31836 , \31819 , \31835 );
and \U$31493 ( \31837 , \23832 , \24149 );
and \U$31494 ( \31838 , \23665 , \24147 );
nor \U$31495 ( \31839 , \31837 , \31838 );
xnor \U$31496 ( \31840 , \31839 , \23944 );
and \U$31497 ( \31841 , \24089 , \23743 );
and \U$31498 ( \31842 , \23970 , \23741 );
nor \U$31499 ( \31843 , \31841 , \31842 );
xnor \U$31500 ( \31844 , \31843 , \23594 );
and \U$31501 ( \31845 , \31840 , \31844 );
and \U$31502 ( \31846 , \24714 , \23421 );
and \U$31503 ( \31847 , \24506 , \23419 );
nor \U$31504 ( \31848 , \31846 , \31847 );
xnor \U$31505 ( \31849 , \31848 , \23279 );
and \U$31506 ( \31850 , \31844 , \31849 );
and \U$31507 ( \31851 , \31840 , \31849 );
or \U$31508 ( \31852 , \31845 , \31850 , \31851 );
and \U$31509 ( \31853 , \31835 , \31852 );
and \U$31510 ( \31854 , \31819 , \31852 );
or \U$31511 ( \31855 , \31836 , \31853 , \31854 );
and \U$31512 ( \31856 , \21689 , \28063 );
and \U$31513 ( \31857 , \21478 , \28061 );
nor \U$31514 ( \31858 , \31856 , \31857 );
xnor \U$31515 ( \31859 , \31858 , \27803 );
and \U$31516 ( \31860 , \21813 , \27569 );
and \U$31517 ( \31861 , \21750 , \27567 );
nor \U$31518 ( \31862 , \31860 , \31861 );
xnor \U$31519 ( \31863 , \31862 , \27254 );
and \U$31520 ( \31864 , \31859 , \31863 );
and \U$31521 ( \31865 , \22099 , \27060 );
and \U$31522 ( \31866 , \22011 , \27058 );
nor \U$31523 ( \31867 , \31865 , \31866 );
xnor \U$31524 ( \31868 , \31867 , \26720 );
and \U$31525 ( \31869 , \31863 , \31868 );
and \U$31526 ( \31870 , \31859 , \31868 );
or \U$31527 ( \31871 , \31864 , \31869 , \31870 );
and \U$31528 ( \31872 , \21428 , \29721 );
and \U$31529 ( \31873 , \21436 , \29719 );
nor \U$31530 ( \31874 , \31872 , \31873 );
xnor \U$31531 ( \31875 , \31874 , \29350 );
and \U$31532 ( \31876 , \21444 , \29159 );
and \U$31533 ( \31877 , \21452 , \29157 );
nor \U$31534 ( \31878 , \31876 , \31877 );
xnor \U$31535 ( \31879 , \31878 , \28841 );
and \U$31536 ( \31880 , \31875 , \31879 );
and \U$31537 ( \31881 , \21463 , \28592 );
and \U$31538 ( \31882 , \21471 , \28590 );
nor \U$31539 ( \31883 , \31881 , \31882 );
xnor \U$31540 ( \31884 , \31883 , \28343 );
and \U$31541 ( \31885 , \31879 , \31884 );
and \U$31542 ( \31886 , \31875 , \31884 );
or \U$31543 ( \31887 , \31880 , \31885 , \31886 );
and \U$31544 ( \31888 , \31871 , \31887 );
and \U$31545 ( \31889 , \21379 , \31639 );
and \U$31546 ( \31890 , \21387 , \31636 );
nor \U$31547 ( \31891 , \31889 , \31890 );
xnor \U$31548 ( \31892 , \31891 , \30584 );
and \U$31549 ( \31893 , \21395 , \30826 );
and \U$31550 ( \31894 , \21403 , \30824 );
nor \U$31551 ( \31895 , \31893 , \31894 );
xnor \U$31552 ( \31896 , \31895 , \30587 );
and \U$31553 ( \31897 , \31892 , \31896 );
and \U$31554 ( \31898 , \21413 , \30258 );
and \U$31555 ( \31899 , \21421 , \30256 );
nor \U$31556 ( \31900 , \31898 , \31899 );
xnor \U$31557 ( \31901 , \31900 , \29948 );
and \U$31558 ( \31902 , \31896 , \31901 );
and \U$31559 ( \31903 , \31892 , \31901 );
or \U$31560 ( \31904 , \31897 , \31902 , \31903 );
and \U$31561 ( \31905 , \31887 , \31904 );
and \U$31562 ( \31906 , \31871 , \31904 );
or \U$31563 ( \31907 , \31888 , \31905 , \31906 );
and \U$31564 ( \31908 , \31855 , \31907 );
and \U$31565 ( \31909 , \26078 , \22379 );
and \U$31566 ( \31910 , \26073 , \22377 );
nor \U$31567 ( \31911 , \31909 , \31910 );
xnor \U$31568 ( \31912 , \31911 , \22266 );
and \U$31569 ( \31913 , \26601 , \22185 );
and \U$31570 ( \31914 , \26342 , \22183 );
nor \U$31571 ( \31915 , \31913 , \31914 );
xnor \U$31572 ( \31916 , \31915 , \22049 );
and \U$31573 ( \31917 , \31912 , \31916 );
and \U$31574 ( \31918 , \26982 , \21985 );
and \U$31575 ( \31919 , \26973 , \21983 );
nor \U$31576 ( \31920 , \31918 , \31919 );
xnor \U$31577 ( \31921 , \31920 , \21907 );
and \U$31578 ( \31922 , \31916 , \31921 );
and \U$31579 ( \31923 , \31912 , \31921 );
or \U$31580 ( \31924 , \31917 , \31922 , \31923 );
and \U$31581 ( \31925 , \24841 , \23125 );
and \U$31582 ( \31926 , \24836 , \23123 );
nor \U$31583 ( \31927 , \31925 , \31926 );
xnor \U$31584 ( \31928 , \31927 , \22988 );
and \U$31585 ( \31929 , \25294 , \22919 );
and \U$31586 ( \31930 , \25097 , \22917 );
nor \U$31587 ( \31931 , \31929 , \31930 );
xnor \U$31588 ( \31932 , \31931 , \22767 );
and \U$31589 ( \31933 , \31928 , \31932 );
and \U$31590 ( \31934 , \25604 , \22651 );
and \U$31591 ( \31935 , \25596 , \22649 );
nor \U$31592 ( \31936 , \31934 , \31935 );
xnor \U$31593 ( \31937 , \31936 , \22495 );
and \U$31594 ( \31938 , \31932 , \31937 );
and \U$31595 ( \31939 , \31928 , \31937 );
or \U$31596 ( \31940 , \31933 , \31938 , \31939 );
and \U$31597 ( \31941 , \31924 , \31940 );
and \U$31598 ( \31942 , \27527 , \21821 );
and \U$31599 ( \31943 , \27325 , \21819 );
nor \U$31600 ( \31944 , \31942 , \31943 );
xnor \U$31601 ( \31945 , \31944 , \21727 );
and \U$31602 ( \31946 , \28002 , \21652 );
and \U$31603 ( \31947 , \27830 , \21650 );
nor \U$31604 ( \31948 , \31946 , \31947 );
xnor \U$31605 ( \31949 , \31948 , \21377 );
and \U$31606 ( \31950 , \31945 , \31949 );
and \U$31607 ( \31951 , \28952 , \21385 );
and \U$31608 ( \31952 , \28528 , \21383 );
nor \U$31609 ( \31953 , \31951 , \31952 );
xnor \U$31610 ( \31954 , \31953 , \21392 );
and \U$31611 ( \31955 , \31949 , \31954 );
and \U$31612 ( \31956 , \31945 , \31954 );
or \U$31613 ( \31957 , \31950 , \31955 , \31956 );
and \U$31614 ( \31958 , \31940 , \31957 );
and \U$31615 ( \31959 , \31924 , \31957 );
or \U$31616 ( \31960 , \31941 , \31958 , \31959 );
and \U$31617 ( \31961 , \31907 , \31960 );
and \U$31618 ( \31962 , \31855 , \31960 );
or \U$31619 ( \31963 , \31908 , \31961 , \31962 );
and \U$31620 ( \31964 , \31803 , \31963 );
xor \U$31621 ( \31965 , \31606 , \31610 );
xor \U$31622 ( \31966 , \31965 , \31615 );
xor \U$31623 ( \31967 , \31622 , \31626 );
xor \U$31624 ( \31968 , \31967 , \31631 );
and \U$31625 ( \31969 , \31966 , \31968 );
xor \U$31626 ( \31970 , \31586 , \31590 );
xor \U$31627 ( \31971 , \31970 , \31595 );
and \U$31628 ( \31972 , \31968 , \31971 );
and \U$31629 ( \31973 , \31966 , \31971 );
or \U$31630 ( \31974 , \31969 , \31972 , \31973 );
xor \U$31631 ( \31975 , \31656 , \31658 );
xor \U$31632 ( \31976 , \31975 , \31661 );
and \U$31633 ( \31977 , \31974 , \31976 );
xor \U$31634 ( \31978 , \31666 , \31668 );
and \U$31635 ( \31979 , \31976 , \31978 );
and \U$31636 ( \31980 , \31974 , \31978 );
or \U$31637 ( \31981 , \31977 , \31979 , \31980 );
and \U$31638 ( \31982 , \31963 , \31981 );
and \U$31639 ( \31983 , \31803 , \31981 );
or \U$31640 ( \31984 , \31964 , \31982 , \31983 );
xor \U$31641 ( \31985 , \31513 , \31529 );
xor \U$31642 ( \31986 , \31985 , \31546 );
xor \U$31643 ( \31987 , \31565 , \31581 );
xor \U$31644 ( \31988 , \31987 , \31598 );
and \U$31645 ( \31989 , \31986 , \31988 );
xor \U$31646 ( \31990 , \31618 , \31634 );
xor \U$31647 ( \31991 , \31990 , \31647 );
and \U$31648 ( \31992 , \31988 , \31991 );
and \U$31649 ( \31993 , \31986 , \31991 );
or \U$31650 ( \31994 , \31989 , \31992 , \31993 );
xor \U$31651 ( \31995 , \31442 , \31444 );
xor \U$31652 ( \31996 , \31995 , \31447 );
xor \U$31653 ( \31997 , \31452 , \31454 );
xor \U$31654 ( \31998 , \31997 , \31457 );
and \U$31655 ( \31999 , \31996 , \31998 );
xnor \U$31656 ( \32000 , \31477 , \31493 );
and \U$31657 ( \32001 , \31998 , \32000 );
and \U$31658 ( \32002 , \31996 , \32000 );
or \U$31659 ( \32003 , \31999 , \32001 , \32002 );
and \U$31660 ( \32004 , \31994 , \32003 );
xor \U$31661 ( \32005 , \31197 , \31213 );
xor \U$31662 ( \32006 , \32005 , \31230 );
and \U$31663 ( \32007 , \32003 , \32006 );
and \U$31664 ( \32008 , \31994 , \32006 );
or \U$31665 ( \32009 , \32004 , \32007 , \32008 );
and \U$31666 ( \32010 , \31984 , \32009 );
xor \U$31667 ( \32011 , \31664 , \31669 );
xor \U$31668 ( \32012 , \32011 , \31672 );
xor \U$31669 ( \32013 , \31680 , \31682 );
xor \U$31670 ( \32014 , \32013 , \31685 );
and \U$31671 ( \32015 , \32012 , \32014 );
xor \U$31672 ( \32016 , \31690 , \31692 );
xor \U$31673 ( \32017 , \32016 , \31695 );
and \U$31674 ( \32018 , \32014 , \32017 );
and \U$31675 ( \32019 , \32012 , \32017 );
or \U$31676 ( \32020 , \32015 , \32018 , \32019 );
and \U$31677 ( \32021 , \32009 , \32020 );
and \U$31678 ( \32022 , \31984 , \32020 );
or \U$31679 ( \32023 , \32010 , \32021 , \32022 );
xor \U$31680 ( \32024 , \31233 , \31285 );
xor \U$31681 ( \32025 , \32024 , \31338 );
xor \U$31682 ( \32026 , \31688 , \31698 );
xor \U$31683 ( \32027 , \32026 , \31701 );
and \U$31684 ( \32028 , \32025 , \32027 );
xor \U$31685 ( \32029 , \31707 , \31709 );
xor \U$31686 ( \32030 , \32029 , \31712 );
and \U$31687 ( \32031 , \32027 , \32030 );
and \U$31688 ( \32032 , \32025 , \32030 );
or \U$31689 ( \32033 , \32028 , \32031 , \32032 );
and \U$31690 ( \32034 , \32023 , \32033 );
xor \U$31691 ( \32035 , \31184 , \31341 );
xor \U$31692 ( \32036 , \32035 , \31359 );
and \U$31693 ( \32037 , \32033 , \32036 );
and \U$31694 ( \32038 , \32023 , \32036 );
or \U$31695 ( \32039 , \32034 , \32037 , \32038 );
xor \U$31696 ( \32040 , \31678 , \31704 );
xor \U$31697 ( \32041 , \32040 , \31715 );
xor \U$31698 ( \32042 , \31720 , \31722 );
xor \U$31699 ( \32043 , \32042 , \31725 );
and \U$31700 ( \32044 , \32041 , \32043 );
and \U$31701 ( \32045 , \32039 , \32044 );
xor \U$31702 ( \32046 , \31404 , \31406 );
xor \U$31703 ( \32047 , \32046 , \31409 );
and \U$31704 ( \32048 , \32044 , \32047 );
and \U$31705 ( \32049 , \32039 , \32047 );
or \U$31706 ( \32050 , \32045 , \32048 , \32049 );
xor \U$31707 ( \32051 , \31362 , \31388 );
xor \U$31708 ( \32052 , \32051 , \31399 );
xor \U$31709 ( \32053 , \31718 , \31728 );
xor \U$31710 ( \32054 , \32053 , \31731 );
and \U$31711 ( \32055 , \32052 , \32054 );
and \U$31712 ( \32056 , \32050 , \32055 );
xor \U$31713 ( \32057 , \31734 , \31736 );
xor \U$31714 ( \32058 , \32057 , \31739 );
and \U$31715 ( \32059 , \32055 , \32058 );
and \U$31716 ( \32060 , \32050 , \32058 );
or \U$31717 ( \32061 , \32056 , \32059 , \32060 );
and \U$31718 ( \32062 , \31754 , \32061 );
xor \U$31719 ( \32063 , \31754 , \32061 );
xor \U$31720 ( \32064 , \32050 , \32055 );
xor \U$31721 ( \32065 , \32064 , \32058 );
and \U$31722 ( \32066 , \30986 , \21434 );
and \U$31723 ( \32067 , \30383 , \21432 );
nor \U$31724 ( \32068 , \32066 , \32067 );
xnor \U$31725 ( \32069 , \32068 , \21441 );
and \U$31726 ( \32070 , \31172 , \21450 );
and \U$31727 ( \32071 , \30991 , \21448 );
nor \U$31728 ( \32072 , \32070 , \32071 );
xnor \U$31729 ( \32073 , \32072 , \21457 );
and \U$31730 ( \32074 , \32069 , \32073 );
nand \U$31731 ( \32075 , \31792 , \21467 );
xnor \U$31732 ( \32076 , \32075 , \21476 );
and \U$31733 ( \32077 , \32073 , \32076 );
and \U$31734 ( \32078 , \32069 , \32076 );
or \U$31735 ( \32079 , \32074 , \32077 , \32078 );
and \U$31736 ( \32080 , \29198 , \21385 );
and \U$31737 ( \32081 , \28952 , \21383 );
nor \U$31738 ( \32082 , \32080 , \32081 );
xnor \U$31739 ( \32083 , \32082 , \21392 );
and \U$31740 ( \32084 , \29522 , \21401 );
and \U$31741 ( \32085 , \29203 , \21399 );
nor \U$31742 ( \32086 , \32084 , \32085 );
xnor \U$31743 ( \32087 , \32086 , \21408 );
and \U$31744 ( \32088 , \32083 , \32087 );
and \U$31745 ( \32089 , \30375 , \21419 );
and \U$31746 ( \32090 , \29806 , \21417 );
nor \U$31747 ( \32091 , \32089 , \32090 );
xnor \U$31748 ( \32092 , \32091 , \21426 );
and \U$31749 ( \32093 , \32087 , \32092 );
and \U$31750 ( \32094 , \32083 , \32092 );
or \U$31751 ( \32095 , \32088 , \32093 , \32094 );
and \U$31752 ( \32096 , \32079 , \32095 );
and \U$31753 ( \32097 , \30991 , \21450 );
and \U$31754 ( \32098 , \30986 , \21448 );
nor \U$31755 ( \32099 , \32097 , \32098 );
xnor \U$31756 ( \32100 , \32099 , \21457 );
and \U$31757 ( \32101 , \32095 , \32100 );
and \U$31758 ( \32102 , \32079 , \32100 );
or \U$31759 ( \32103 , \32096 , \32101 , \32102 );
and \U$31760 ( \32104 , \31792 , \21469 );
and \U$31761 ( \32105 , \31172 , \21467 );
nor \U$31762 ( \32106 , \32104 , \32105 );
xnor \U$31763 ( \32107 , \32106 , \21476 );
xor \U$31764 ( \32108 , \31945 , \31949 );
xor \U$31765 ( \32109 , \32108 , \31954 );
and \U$31766 ( \32110 , \32107 , \32109 );
xor \U$31767 ( \32111 , \31779 , \31783 );
xor \U$31768 ( \32112 , \32111 , \31788 );
and \U$31769 ( \32113 , \32109 , \32112 );
and \U$31770 ( \32114 , \32107 , \32112 );
or \U$31771 ( \32115 , \32110 , \32113 , \32114 );
and \U$31772 ( \32116 , \32103 , \32115 );
xor \U$31773 ( \32117 , \31912 , \31916 );
xor \U$31774 ( \32118 , \32117 , \31921 );
xor \U$31775 ( \32119 , \31928 , \31932 );
xor \U$31776 ( \32120 , \32119 , \31937 );
and \U$31777 ( \32121 , \32118 , \32120 );
xor \U$31778 ( \32122 , \31840 , \31844 );
xor \U$31779 ( \32123 , \32122 , \31849 );
and \U$31780 ( \32124 , \32120 , \32123 );
and \U$31781 ( \32125 , \32118 , \32123 );
or \U$31782 ( \32126 , \32121 , \32124 , \32125 );
and \U$31783 ( \32127 , \32115 , \32126 );
and \U$31784 ( \32128 , \32103 , \32126 );
or \U$31785 ( \32129 , \32116 , \32127 , \32128 );
and \U$31786 ( \32130 , \26073 , \22651 );
and \U$31787 ( \32131 , \25604 , \22649 );
nor \U$31788 ( \32132 , \32130 , \32131 );
xnor \U$31789 ( \32133 , \32132 , \22495 );
and \U$31790 ( \32134 , \26342 , \22379 );
and \U$31791 ( \32135 , \26078 , \22377 );
nor \U$31792 ( \32136 , \32134 , \32135 );
xnor \U$31793 ( \32137 , \32136 , \22266 );
and \U$31794 ( \32138 , \32133 , \32137 );
and \U$31795 ( \32139 , \26973 , \22185 );
and \U$31796 ( \32140 , \26601 , \22183 );
nor \U$31797 ( \32141 , \32139 , \32140 );
xnor \U$31798 ( \32142 , \32141 , \22049 );
and \U$31799 ( \32143 , \32137 , \32142 );
and \U$31800 ( \32144 , \32133 , \32142 );
or \U$31801 ( \32145 , \32138 , \32143 , \32144 );
and \U$31802 ( \32146 , \24836 , \23421 );
and \U$31803 ( \32147 , \24714 , \23419 );
nor \U$31804 ( \32148 , \32146 , \32147 );
xnor \U$31805 ( \32149 , \32148 , \23279 );
and \U$31806 ( \32150 , \25097 , \23125 );
and \U$31807 ( \32151 , \24841 , \23123 );
nor \U$31808 ( \32152 , \32150 , \32151 );
xnor \U$31809 ( \32153 , \32152 , \22988 );
and \U$31810 ( \32154 , \32149 , \32153 );
and \U$31811 ( \32155 , \25596 , \22919 );
and \U$31812 ( \32156 , \25294 , \22917 );
nor \U$31813 ( \32157 , \32155 , \32156 );
xnor \U$31814 ( \32158 , \32157 , \22767 );
and \U$31815 ( \32159 , \32153 , \32158 );
and \U$31816 ( \32160 , \32149 , \32158 );
or \U$31817 ( \32161 , \32154 , \32159 , \32160 );
and \U$31818 ( \32162 , \32145 , \32161 );
and \U$31819 ( \32163 , \27325 , \21985 );
and \U$31820 ( \32164 , \26982 , \21983 );
nor \U$31821 ( \32165 , \32163 , \32164 );
xnor \U$31822 ( \32166 , \32165 , \21907 );
and \U$31823 ( \32167 , \27830 , \21821 );
and \U$31824 ( \32168 , \27527 , \21819 );
nor \U$31825 ( \32169 , \32167 , \32168 );
xnor \U$31826 ( \32170 , \32169 , \21727 );
and \U$31827 ( \32171 , \32166 , \32170 );
and \U$31828 ( \32172 , \28528 , \21652 );
and \U$31829 ( \32173 , \28002 , \21650 );
nor \U$31830 ( \32174 , \32172 , \32173 );
xnor \U$31831 ( \32175 , \32174 , \21377 );
and \U$31832 ( \32176 , \32170 , \32175 );
and \U$31833 ( \32177 , \32166 , \32175 );
or \U$31834 ( \32178 , \32171 , \32176 , \32177 );
and \U$31835 ( \32179 , \32161 , \32178 );
and \U$31836 ( \32180 , \32145 , \32178 );
or \U$31837 ( \32181 , \32162 , \32179 , \32180 );
and \U$31838 ( \32182 , \21478 , \28592 );
and \U$31839 ( \32183 , \21463 , \28590 );
nor \U$31840 ( \32184 , \32182 , \32183 );
xnor \U$31841 ( \32185 , \32184 , \28343 );
and \U$31842 ( \32186 , \21750 , \28063 );
and \U$31843 ( \32187 , \21689 , \28061 );
nor \U$31844 ( \32188 , \32186 , \32187 );
xnor \U$31845 ( \32189 , \32188 , \27803 );
and \U$31846 ( \32190 , \32185 , \32189 );
and \U$31847 ( \32191 , \22011 , \27569 );
and \U$31848 ( \32192 , \21813 , \27567 );
nor \U$31849 ( \32193 , \32191 , \32192 );
xnor \U$31850 ( \32194 , \32193 , \27254 );
and \U$31851 ( \32195 , \32189 , \32194 );
and \U$31852 ( \32196 , \32185 , \32194 );
or \U$31853 ( \32197 , \32190 , \32195 , \32196 );
and \U$31854 ( \32198 , \21403 , \31639 );
and \U$31855 ( \32199 , \21379 , \31636 );
nor \U$31856 ( \32200 , \32198 , \32199 );
xnor \U$31857 ( \32201 , \32200 , \30584 );
and \U$31858 ( \32202 , \21421 , \30826 );
and \U$31859 ( \32203 , \21395 , \30824 );
nor \U$31860 ( \32204 , \32202 , \32203 );
xnor \U$31861 ( \32205 , \32204 , \30587 );
and \U$31862 ( \32206 , \32201 , \32205 );
and \U$31863 ( \32207 , \32205 , \21476 );
and \U$31864 ( \32208 , \32201 , \21476 );
or \U$31865 ( \32209 , \32206 , \32207 , \32208 );
and \U$31866 ( \32210 , \32197 , \32209 );
and \U$31867 ( \32211 , \21436 , \30258 );
and \U$31868 ( \32212 , \21413 , \30256 );
nor \U$31869 ( \32213 , \32211 , \32212 );
xnor \U$31870 ( \32214 , \32213 , \29948 );
and \U$31871 ( \32215 , \21452 , \29721 );
and \U$31872 ( \32216 , \21428 , \29719 );
nor \U$31873 ( \32217 , \32215 , \32216 );
xnor \U$31874 ( \32218 , \32217 , \29350 );
and \U$31875 ( \32219 , \32214 , \32218 );
and \U$31876 ( \32220 , \21471 , \29159 );
and \U$31877 ( \32221 , \21444 , \29157 );
nor \U$31878 ( \32222 , \32220 , \32221 );
xnor \U$31879 ( \32223 , \32222 , \28841 );
and \U$31880 ( \32224 , \32218 , \32223 );
and \U$31881 ( \32225 , \32214 , \32223 );
or \U$31882 ( \32226 , \32219 , \32224 , \32225 );
and \U$31883 ( \32227 , \32209 , \32226 );
and \U$31884 ( \32228 , \32197 , \32226 );
or \U$31885 ( \32229 , \32210 , \32227 , \32228 );
and \U$31886 ( \32230 , \32181 , \32229 );
and \U$31887 ( \32231 , \22867 , \25631 );
and \U$31888 ( \32232 , \22624 , \25629 );
nor \U$31889 ( \32233 , \32231 , \32232 );
xnor \U$31890 ( \32234 , \32233 , \25399 );
and \U$31891 ( \32235 , \23058 , \25180 );
and \U$31892 ( \32236 , \22872 , \25178 );
nor \U$31893 ( \32237 , \32235 , \32236 );
xnor \U$31894 ( \32238 , \32237 , \25037 );
and \U$31895 ( \32239 , \32234 , \32238 );
and \U$31896 ( \32240 , \23466 , \24857 );
and \U$31897 ( \32241 , \23202 , \24855 );
nor \U$31898 ( \32242 , \32240 , \32241 );
xnor \U$31899 ( \32243 , \32242 , \24611 );
and \U$31900 ( \32244 , \32238 , \32243 );
and \U$31901 ( \32245 , \32234 , \32243 );
or \U$31902 ( \32246 , \32239 , \32244 , \32245 );
and \U$31903 ( \32247 , \22204 , \27060 );
and \U$31904 ( \32248 , \22099 , \27058 );
nor \U$31905 ( \32249 , \32247 , \32248 );
xnor \U$31906 ( \32250 , \32249 , \26720 );
and \U$31907 ( \32251 , \22325 , \26471 );
and \U$31908 ( \32252 , \22209 , \26469 );
nor \U$31909 ( \32253 , \32251 , \32252 );
xnor \U$31910 ( \32254 , \32253 , \26230 );
and \U$31911 ( \32255 , \32250 , \32254 );
and \U$31912 ( \32256 , \22616 , \26005 );
and \U$31913 ( \32257 , \22440 , \26003 );
nor \U$31914 ( \32258 , \32256 , \32257 );
xnor \U$31915 ( \32259 , \32258 , \25817 );
and \U$31916 ( \32260 , \32254 , \32259 );
and \U$31917 ( \32261 , \32250 , \32259 );
or \U$31918 ( \32262 , \32255 , \32260 , \32261 );
and \U$31919 ( \32263 , \32246 , \32262 );
and \U$31920 ( \32264 , \23665 , \24462 );
and \U$31921 ( \32265 , \23491 , \24460 );
nor \U$31922 ( \32266 , \32264 , \32265 );
xnor \U$31923 ( \32267 , \32266 , \24275 );
and \U$31924 ( \32268 , \23970 , \24149 );
and \U$31925 ( \32269 , \23832 , \24147 );
nor \U$31926 ( \32270 , \32268 , \32269 );
xnor \U$31927 ( \32271 , \32270 , \23944 );
and \U$31928 ( \32272 , \32267 , \32271 );
and \U$31929 ( \32273 , \24506 , \23743 );
and \U$31930 ( \32274 , \24089 , \23741 );
nor \U$31931 ( \32275 , \32273 , \32274 );
xnor \U$31932 ( \32276 , \32275 , \23594 );
and \U$31933 ( \32277 , \32271 , \32276 );
and \U$31934 ( \32278 , \32267 , \32276 );
or \U$31935 ( \32279 , \32272 , \32277 , \32278 );
and \U$31936 ( \32280 , \32262 , \32279 );
and \U$31937 ( \32281 , \32246 , \32279 );
or \U$31938 ( \32282 , \32263 , \32280 , \32281 );
and \U$31939 ( \32283 , \32229 , \32282 );
and \U$31940 ( \32284 , \32181 , \32282 );
or \U$31941 ( \32285 , \32230 , \32283 , \32284 );
and \U$31942 ( \32286 , \32129 , \32285 );
xor \U$31943 ( \32287 , \31807 , \31811 );
xor \U$31944 ( \32288 , \32287 , \31816 );
xor \U$31945 ( \32289 , \31823 , \31827 );
xor \U$31946 ( \32290 , \32289 , \31832 );
and \U$31947 ( \32291 , \32288 , \32290 );
xor \U$31948 ( \32292 , \31859 , \31863 );
xor \U$31949 ( \32293 , \32292 , \31868 );
and \U$31950 ( \32294 , \32290 , \32293 );
and \U$31951 ( \32295 , \32288 , \32293 );
or \U$31952 ( \32296 , \32291 , \32294 , \32295 );
xor \U$31953 ( \32297 , \31875 , \31879 );
xor \U$31954 ( \32298 , \32297 , \31884 );
xor \U$31955 ( \32299 , \31892 , \31896 );
xor \U$31956 ( \32300 , \32299 , \31901 );
and \U$31957 ( \32301 , \32298 , \32300 );
and \U$31958 ( \32302 , \32296 , \32301 );
xor \U$31959 ( \32303 , \31642 , \31646 );
and \U$31960 ( \32304 , \32301 , \32303 );
and \U$31961 ( \32305 , \32296 , \32303 );
or \U$31962 ( \32306 , \32302 , \32304 , \32305 );
and \U$31963 ( \32307 , \32285 , \32306 );
and \U$31964 ( \32308 , \32129 , \32306 );
or \U$31965 ( \32309 , \32286 , \32307 , \32308 );
xor \U$31966 ( \32310 , \31819 , \31835 );
xor \U$31967 ( \32311 , \32310 , \31852 );
xor \U$31968 ( \32312 , \31924 , \31940 );
xor \U$31969 ( \32313 , \32312 , \31957 );
and \U$31970 ( \32314 , \32311 , \32313 );
xor \U$31971 ( \32315 , \31791 , \31794 );
xor \U$31972 ( \32316 , \32315 , \31797 );
and \U$31973 ( \32317 , \32313 , \32316 );
and \U$31974 ( \32318 , \32311 , \32316 );
or \U$31975 ( \32319 , \32314 , \32317 , \32318 );
xor \U$31976 ( \32320 , \31966 , \31968 );
xor \U$31977 ( \32321 , \32320 , \31971 );
xor \U$31978 ( \32322 , \31756 , \31758 );
xor \U$31979 ( \32323 , \32322 , \31761 );
and \U$31980 ( \32324 , \32321 , \32323 );
xor \U$31981 ( \32325 , \31766 , \31768 );
xor \U$31982 ( \32326 , \32325 , \31771 );
and \U$31983 ( \32327 , \32323 , \32326 );
and \U$31984 ( \32328 , \32321 , \32326 );
or \U$31985 ( \32329 , \32324 , \32327 , \32328 );
and \U$31986 ( \32330 , \32319 , \32329 );
xor \U$31987 ( \32331 , \31986 , \31988 );
xor \U$31988 ( \32332 , \32331 , \31991 );
and \U$31989 ( \32333 , \32329 , \32332 );
and \U$31990 ( \32334 , \32319 , \32332 );
or \U$31991 ( \32335 , \32330 , \32333 , \32334 );
and \U$31992 ( \32336 , \32309 , \32335 );
xor \U$31993 ( \32337 , \31764 , \31774 );
xor \U$31994 ( \32338 , \32337 , \31800 );
xor \U$31995 ( \32339 , \31996 , \31998 );
xor \U$31996 ( \32340 , \32339 , \32000 );
and \U$31997 ( \32341 , \32338 , \32340 );
xor \U$31998 ( \32342 , \31974 , \31976 );
xor \U$31999 ( \32343 , \32342 , \31978 );
and \U$32000 ( \32344 , \32340 , \32343 );
and \U$32001 ( \32345 , \32338 , \32343 );
or \U$32002 ( \32346 , \32341 , \32344 , \32345 );
and \U$32003 ( \32347 , \32335 , \32346 );
and \U$32004 ( \32348 , \32309 , \32346 );
or \U$32005 ( \32349 , \32336 , \32347 , \32348 );
xor \U$32006 ( \32350 , \31450 , \31460 );
xor \U$32007 ( \32351 , \32350 , \31494 );
xor \U$32008 ( \32352 , \31549 , \31601 );
xor \U$32009 ( \32353 , \32352 , \31650 );
and \U$32010 ( \32354 , \32351 , \32353 );
xor \U$32011 ( \32355 , \32012 , \32014 );
xor \U$32012 ( \32356 , \32355 , \32017 );
and \U$32013 ( \32357 , \32353 , \32356 );
and \U$32014 ( \32358 , \32351 , \32356 );
or \U$32015 ( \32359 , \32354 , \32357 , \32358 );
and \U$32016 ( \32360 , \32349 , \32359 );
xor \U$32017 ( \32361 , \31497 , \31653 );
xor \U$32018 ( \32362 , \32361 , \31675 );
and \U$32019 ( \32363 , \32359 , \32362 );
and \U$32020 ( \32364 , \32349 , \32362 );
or \U$32021 ( \32365 , \32360 , \32363 , \32364 );
xor \U$32022 ( \32366 , \32023 , \32033 );
xor \U$32023 ( \32367 , \32366 , \32036 );
and \U$32024 ( \32368 , \32365 , \32367 );
xor \U$32025 ( \32369 , \32041 , \32043 );
and \U$32026 ( \32370 , \32367 , \32369 );
and \U$32027 ( \32371 , \32365 , \32369 );
or \U$32028 ( \32372 , \32368 , \32370 , \32371 );
xor \U$32029 ( \32373 , \32039 , \32044 );
xor \U$32030 ( \32374 , \32373 , \32047 );
and \U$32031 ( \32375 , \32372 , \32374 );
xor \U$32032 ( \32376 , \32052 , \32054 );
and \U$32033 ( \32377 , \32374 , \32376 );
and \U$32034 ( \32378 , \32372 , \32376 );
or \U$32035 ( \32379 , \32375 , \32377 , \32378 );
and \U$32036 ( \32380 , \32065 , \32379 );
xor \U$32037 ( \32381 , \32065 , \32379 );
xor \U$32038 ( \32382 , \32372 , \32374 );
xor \U$32039 ( \32383 , \32382 , \32376 );
and \U$32040 ( \32384 , \21444 , \29721 );
and \U$32041 ( \32385 , \21452 , \29719 );
nor \U$32042 ( \32386 , \32384 , \32385 );
xnor \U$32043 ( \32387 , \32386 , \29350 );
and \U$32044 ( \32388 , \21463 , \29159 );
and \U$32045 ( \32389 , \21471 , \29157 );
nor \U$32046 ( \32390 , \32388 , \32389 );
xnor \U$32047 ( \32391 , \32390 , \28841 );
and \U$32048 ( \32392 , \32387 , \32391 );
and \U$32049 ( \32393 , \21689 , \28592 );
and \U$32050 ( \32394 , \21478 , \28590 );
nor \U$32051 ( \32395 , \32393 , \32394 );
xnor \U$32052 ( \32396 , \32395 , \28343 );
and \U$32053 ( \32397 , \32391 , \32396 );
and \U$32054 ( \32398 , \32387 , \32396 );
or \U$32055 ( \32399 , \32392 , \32397 , \32398 );
and \U$32056 ( \32400 , \21395 , \31639 );
and \U$32057 ( \32401 , \21403 , \31636 );
nor \U$32058 ( \32402 , \32400 , \32401 );
xnor \U$32059 ( \32403 , \32402 , \30584 );
and \U$32060 ( \32404 , \21413 , \30826 );
and \U$32061 ( \32405 , \21421 , \30824 );
nor \U$32062 ( \32406 , \32404 , \32405 );
xnor \U$32063 ( \32407 , \32406 , \30587 );
and \U$32064 ( \32408 , \32403 , \32407 );
and \U$32065 ( \32409 , \21428 , \30258 );
and \U$32066 ( \32410 , \21436 , \30256 );
nor \U$32067 ( \32411 , \32409 , \32410 );
xnor \U$32068 ( \32412 , \32411 , \29948 );
and \U$32069 ( \32413 , \32407 , \32412 );
and \U$32070 ( \32414 , \32403 , \32412 );
or \U$32071 ( \32415 , \32408 , \32413 , \32414 );
and \U$32072 ( \32416 , \32399 , \32415 );
and \U$32073 ( \32417 , \21813 , \28063 );
and \U$32074 ( \32418 , \21750 , \28061 );
nor \U$32075 ( \32419 , \32417 , \32418 );
xnor \U$32076 ( \32420 , \32419 , \27803 );
and \U$32077 ( \32421 , \22099 , \27569 );
and \U$32078 ( \32422 , \22011 , \27567 );
nor \U$32079 ( \32423 , \32421 , \32422 );
xnor \U$32080 ( \32424 , \32423 , \27254 );
and \U$32081 ( \32425 , \32420 , \32424 );
and \U$32082 ( \32426 , \22209 , \27060 );
and \U$32083 ( \32427 , \22204 , \27058 );
nor \U$32084 ( \32428 , \32426 , \32427 );
xnor \U$32085 ( \32429 , \32428 , \26720 );
and \U$32086 ( \32430 , \32424 , \32429 );
and \U$32087 ( \32431 , \32420 , \32429 );
or \U$32088 ( \32432 , \32425 , \32430 , \32431 );
and \U$32089 ( \32433 , \32415 , \32432 );
and \U$32090 ( \32434 , \32399 , \32432 );
or \U$32091 ( \32435 , \32416 , \32433 , \32434 );
and \U$32092 ( \32436 , \26601 , \22379 );
and \U$32093 ( \32437 , \26342 , \22377 );
nor \U$32094 ( \32438 , \32436 , \32437 );
xnor \U$32095 ( \32439 , \32438 , \22266 );
and \U$32096 ( \32440 , \26982 , \22185 );
and \U$32097 ( \32441 , \26973 , \22183 );
nor \U$32098 ( \32442 , \32440 , \32441 );
xnor \U$32099 ( \32443 , \32442 , \22049 );
and \U$32100 ( \32444 , \32439 , \32443 );
and \U$32101 ( \32445 , \27527 , \21985 );
and \U$32102 ( \32446 , \27325 , \21983 );
nor \U$32103 ( \32447 , \32445 , \32446 );
xnor \U$32104 ( \32448 , \32447 , \21907 );
and \U$32105 ( \32449 , \32443 , \32448 );
and \U$32106 ( \32450 , \32439 , \32448 );
or \U$32107 ( \32451 , \32444 , \32449 , \32450 );
and \U$32108 ( \32452 , \28002 , \21821 );
and \U$32109 ( \32453 , \27830 , \21819 );
nor \U$32110 ( \32454 , \32452 , \32453 );
xnor \U$32111 ( \32455 , \32454 , \21727 );
and \U$32112 ( \32456 , \28952 , \21652 );
and \U$32113 ( \32457 , \28528 , \21650 );
nor \U$32114 ( \32458 , \32456 , \32457 );
xnor \U$32115 ( \32459 , \32458 , \21377 );
and \U$32116 ( \32460 , \32455 , \32459 );
and \U$32117 ( \32461 , \29203 , \21385 );
and \U$32118 ( \32462 , \29198 , \21383 );
nor \U$32119 ( \32463 , \32461 , \32462 );
xnor \U$32120 ( \32464 , \32463 , \21392 );
and \U$32121 ( \32465 , \32459 , \32464 );
and \U$32122 ( \32466 , \32455 , \32464 );
or \U$32123 ( \32467 , \32460 , \32465 , \32466 );
and \U$32124 ( \32468 , \32451 , \32467 );
and \U$32125 ( \32469 , \25294 , \23125 );
and \U$32126 ( \32470 , \25097 , \23123 );
nor \U$32127 ( \32471 , \32469 , \32470 );
xnor \U$32128 ( \32472 , \32471 , \22988 );
and \U$32129 ( \32473 , \25604 , \22919 );
and \U$32130 ( \32474 , \25596 , \22917 );
nor \U$32131 ( \32475 , \32473 , \32474 );
xnor \U$32132 ( \32476 , \32475 , \22767 );
and \U$32133 ( \32477 , \32472 , \32476 );
and \U$32134 ( \32478 , \26078 , \22651 );
and \U$32135 ( \32479 , \26073 , \22649 );
nor \U$32136 ( \32480 , \32478 , \32479 );
xnor \U$32137 ( \32481 , \32480 , \22495 );
and \U$32138 ( \32482 , \32476 , \32481 );
and \U$32139 ( \32483 , \32472 , \32481 );
or \U$32140 ( \32484 , \32477 , \32482 , \32483 );
and \U$32141 ( \32485 , \32467 , \32484 );
and \U$32142 ( \32486 , \32451 , \32484 );
or \U$32143 ( \32487 , \32468 , \32485 , \32486 );
and \U$32144 ( \32488 , \32435 , \32487 );
and \U$32145 ( \32489 , \22440 , \26471 );
and \U$32146 ( \32490 , \22325 , \26469 );
nor \U$32147 ( \32491 , \32489 , \32490 );
xnor \U$32148 ( \32492 , \32491 , \26230 );
and \U$32149 ( \32493 , \22624 , \26005 );
and \U$32150 ( \32494 , \22616 , \26003 );
nor \U$32151 ( \32495 , \32493 , \32494 );
xnor \U$32152 ( \32496 , \32495 , \25817 );
and \U$32153 ( \32497 , \32492 , \32496 );
and \U$32154 ( \32498 , \22872 , \25631 );
and \U$32155 ( \32499 , \22867 , \25629 );
nor \U$32156 ( \32500 , \32498 , \32499 );
xnor \U$32157 ( \32501 , \32500 , \25399 );
and \U$32158 ( \32502 , \32496 , \32501 );
and \U$32159 ( \32503 , \32492 , \32501 );
or \U$32160 ( \32504 , \32497 , \32502 , \32503 );
and \U$32161 ( \32505 , \24089 , \24149 );
and \U$32162 ( \32506 , \23970 , \24147 );
nor \U$32163 ( \32507 , \32505 , \32506 );
xnor \U$32164 ( \32508 , \32507 , \23944 );
and \U$32165 ( \32509 , \24714 , \23743 );
and \U$32166 ( \32510 , \24506 , \23741 );
nor \U$32167 ( \32511 , \32509 , \32510 );
xnor \U$32168 ( \32512 , \32511 , \23594 );
and \U$32169 ( \32513 , \32508 , \32512 );
and \U$32170 ( \32514 , \24841 , \23421 );
and \U$32171 ( \32515 , \24836 , \23419 );
nor \U$32172 ( \32516 , \32514 , \32515 );
xnor \U$32173 ( \32517 , \32516 , \23279 );
and \U$32174 ( \32518 , \32512 , \32517 );
and \U$32175 ( \32519 , \32508 , \32517 );
or \U$32176 ( \32520 , \32513 , \32518 , \32519 );
and \U$32177 ( \32521 , \32504 , \32520 );
and \U$32178 ( \32522 , \23202 , \25180 );
and \U$32179 ( \32523 , \23058 , \25178 );
nor \U$32180 ( \32524 , \32522 , \32523 );
xnor \U$32181 ( \32525 , \32524 , \25037 );
and \U$32182 ( \32526 , \23491 , \24857 );
and \U$32183 ( \32527 , \23466 , \24855 );
nor \U$32184 ( \32528 , \32526 , \32527 );
xnor \U$32185 ( \32529 , \32528 , \24611 );
and \U$32186 ( \32530 , \32525 , \32529 );
and \U$32187 ( \32531 , \23832 , \24462 );
and \U$32188 ( \32532 , \23665 , \24460 );
nor \U$32189 ( \32533 , \32531 , \32532 );
xnor \U$32190 ( \32534 , \32533 , \24275 );
and \U$32191 ( \32535 , \32529 , \32534 );
and \U$32192 ( \32536 , \32525 , \32534 );
or \U$32193 ( \32537 , \32530 , \32535 , \32536 );
and \U$32194 ( \32538 , \32520 , \32537 );
and \U$32195 ( \32539 , \32504 , \32537 );
or \U$32196 ( \32540 , \32521 , \32538 , \32539 );
and \U$32197 ( \32541 , \32487 , \32540 );
and \U$32198 ( \32542 , \32435 , \32540 );
or \U$32199 ( \32543 , \32488 , \32541 , \32542 );
xor \U$32200 ( \32544 , \32234 , \32238 );
xor \U$32201 ( \32545 , \32544 , \32243 );
xor \U$32202 ( \32546 , \32250 , \32254 );
xor \U$32203 ( \32547 , \32546 , \32259 );
and \U$32204 ( \32548 , \32545 , \32547 );
xor \U$32205 ( \32549 , \32267 , \32271 );
xor \U$32206 ( \32550 , \32549 , \32276 );
and \U$32207 ( \32551 , \32547 , \32550 );
and \U$32208 ( \32552 , \32545 , \32550 );
or \U$32209 ( \32553 , \32548 , \32551 , \32552 );
and \U$32210 ( \32554 , \29806 , \21401 );
and \U$32211 ( \32555 , \29522 , \21399 );
nor \U$32212 ( \32556 , \32554 , \32555 );
xnor \U$32213 ( \32557 , \32556 , \21408 );
and \U$32214 ( \32558 , \30383 , \21419 );
and \U$32215 ( \32559 , \30375 , \21417 );
nor \U$32216 ( \32560 , \32558 , \32559 );
xnor \U$32217 ( \32561 , \32560 , \21426 );
and \U$32218 ( \32562 , \32557 , \32561 );
and \U$32219 ( \32563 , \30991 , \21434 );
and \U$32220 ( \32564 , \30986 , \21432 );
nor \U$32221 ( \32565 , \32563 , \32564 );
xnor \U$32222 ( \32566 , \32565 , \21441 );
and \U$32223 ( \32567 , \32561 , \32566 );
and \U$32224 ( \32568 , \32557 , \32566 );
or \U$32225 ( \32569 , \32562 , \32567 , \32568 );
xor \U$32226 ( \32570 , \32069 , \32073 );
xor \U$32227 ( \32571 , \32570 , \32076 );
and \U$32228 ( \32572 , \32569 , \32571 );
xor \U$32229 ( \32573 , \32083 , \32087 );
xor \U$32230 ( \32574 , \32573 , \32092 );
and \U$32231 ( \32575 , \32571 , \32574 );
and \U$32232 ( \32576 , \32569 , \32574 );
or \U$32233 ( \32577 , \32572 , \32575 , \32576 );
and \U$32234 ( \32578 , \32553 , \32577 );
xor \U$32235 ( \32579 , \32133 , \32137 );
xor \U$32236 ( \32580 , \32579 , \32142 );
xor \U$32237 ( \32581 , \32149 , \32153 );
xor \U$32238 ( \32582 , \32581 , \32158 );
and \U$32239 ( \32583 , \32580 , \32582 );
xor \U$32240 ( \32584 , \32166 , \32170 );
xor \U$32241 ( \32585 , \32584 , \32175 );
and \U$32242 ( \32586 , \32582 , \32585 );
and \U$32243 ( \32587 , \32580 , \32585 );
or \U$32244 ( \32588 , \32583 , \32586 , \32587 );
and \U$32245 ( \32589 , \32577 , \32588 );
and \U$32246 ( \32590 , \32553 , \32588 );
or \U$32247 ( \32591 , \32578 , \32589 , \32590 );
and \U$32248 ( \32592 , \32543 , \32591 );
xor \U$32249 ( \32593 , \32185 , \32189 );
xor \U$32250 ( \32594 , \32593 , \32194 );
xor \U$32251 ( \32595 , \32201 , \32205 );
xor \U$32252 ( \32596 , \32595 , \21476 );
and \U$32253 ( \32597 , \32594 , \32596 );
xor \U$32254 ( \32598 , \32214 , \32218 );
xor \U$32255 ( \32599 , \32598 , \32223 );
and \U$32256 ( \32600 , \32596 , \32599 );
and \U$32257 ( \32601 , \32594 , \32599 );
or \U$32258 ( \32602 , \32597 , \32600 , \32601 );
xor \U$32259 ( \32603 , \32288 , \32290 );
xor \U$32260 ( \32604 , \32603 , \32293 );
and \U$32261 ( \32605 , \32602 , \32604 );
xor \U$32262 ( \32606 , \32298 , \32300 );
and \U$32263 ( \32607 , \32604 , \32606 );
and \U$32264 ( \32608 , \32602 , \32606 );
or \U$32265 ( \32609 , \32605 , \32607 , \32608 );
and \U$32266 ( \32610 , \32591 , \32609 );
and \U$32267 ( \32611 , \32543 , \32609 );
or \U$32268 ( \32612 , \32592 , \32610 , \32611 );
xor \U$32269 ( \32613 , \32145 , \32161 );
xor \U$32270 ( \32614 , \32613 , \32178 );
xor \U$32271 ( \32615 , \32197 , \32209 );
xor \U$32272 ( \32616 , \32615 , \32226 );
and \U$32273 ( \32617 , \32614 , \32616 );
xor \U$32274 ( \32618 , \32246 , \32262 );
xor \U$32275 ( \32619 , \32618 , \32279 );
and \U$32276 ( \32620 , \32616 , \32619 );
and \U$32277 ( \32621 , \32614 , \32619 );
or \U$32278 ( \32622 , \32617 , \32620 , \32621 );
xor \U$32279 ( \32623 , \32079 , \32095 );
xor \U$32280 ( \32624 , \32623 , \32100 );
xor \U$32281 ( \32625 , \32107 , \32109 );
xor \U$32282 ( \32626 , \32625 , \32112 );
and \U$32283 ( \32627 , \32624 , \32626 );
xor \U$32284 ( \32628 , \32118 , \32120 );
xor \U$32285 ( \32629 , \32628 , \32123 );
and \U$32286 ( \32630 , \32626 , \32629 );
and \U$32287 ( \32631 , \32624 , \32629 );
or \U$32288 ( \32632 , \32627 , \32630 , \32631 );
and \U$32289 ( \32633 , \32622 , \32632 );
xor \U$32290 ( \32634 , \31871 , \31887 );
xor \U$32291 ( \32635 , \32634 , \31904 );
and \U$32292 ( \32636 , \32632 , \32635 );
and \U$32293 ( \32637 , \32622 , \32635 );
or \U$32294 ( \32638 , \32633 , \32636 , \32637 );
and \U$32295 ( \32639 , \32612 , \32638 );
xor \U$32296 ( \32640 , \32311 , \32313 );
xor \U$32297 ( \32641 , \32640 , \32316 );
xor \U$32298 ( \32642 , \32321 , \32323 );
xor \U$32299 ( \32643 , \32642 , \32326 );
and \U$32300 ( \32644 , \32641 , \32643 );
xor \U$32301 ( \32645 , \32296 , \32301 );
xor \U$32302 ( \32646 , \32645 , \32303 );
and \U$32303 ( \32647 , \32643 , \32646 );
and \U$32304 ( \32648 , \32641 , \32646 );
or \U$32305 ( \32649 , \32644 , \32647 , \32648 );
and \U$32306 ( \32650 , \32638 , \32649 );
and \U$32307 ( \32651 , \32612 , \32649 );
or \U$32308 ( \32652 , \32639 , \32650 , \32651 );
xor \U$32309 ( \32653 , \31855 , \31907 );
xor \U$32310 ( \32654 , \32653 , \31960 );
xor \U$32311 ( \32655 , \32319 , \32329 );
xor \U$32312 ( \32656 , \32655 , \32332 );
and \U$32313 ( \32657 , \32654 , \32656 );
xor \U$32314 ( \32658 , \32338 , \32340 );
xor \U$32315 ( \32659 , \32658 , \32343 );
and \U$32316 ( \32660 , \32656 , \32659 );
and \U$32317 ( \32661 , \32654 , \32659 );
or \U$32318 ( \32662 , \32657 , \32660 , \32661 );
and \U$32319 ( \32663 , \32652 , \32662 );
xor \U$32320 ( \32664 , \31994 , \32003 );
xor \U$32321 ( \32665 , \32664 , \32006 );
and \U$32322 ( \32666 , \32662 , \32665 );
and \U$32323 ( \32667 , \32652 , \32665 );
or \U$32324 ( \32668 , \32663 , \32666 , \32667 );
xor \U$32325 ( \32669 , \31803 , \31963 );
xor \U$32326 ( \32670 , \32669 , \31981 );
xor \U$32327 ( \32671 , \32309 , \32335 );
xor \U$32328 ( \32672 , \32671 , \32346 );
and \U$32329 ( \32673 , \32670 , \32672 );
xor \U$32330 ( \32674 , \32351 , \32353 );
xor \U$32331 ( \32675 , \32674 , \32356 );
and \U$32332 ( \32676 , \32672 , \32675 );
and \U$32333 ( \32677 , \32670 , \32675 );
or \U$32334 ( \32678 , \32673 , \32676 , \32677 );
and \U$32335 ( \32679 , \32668 , \32678 );
xor \U$32336 ( \32680 , \32025 , \32027 );
xor \U$32337 ( \32681 , \32680 , \32030 );
and \U$32338 ( \32682 , \32678 , \32681 );
and \U$32339 ( \32683 , \32668 , \32681 );
or \U$32340 ( \32684 , \32679 , \32682 , \32683 );
xor \U$32341 ( \32685 , \31984 , \32009 );
xor \U$32342 ( \32686 , \32685 , \32020 );
xor \U$32343 ( \32687 , \32349 , \32359 );
xor \U$32344 ( \32688 , \32687 , \32362 );
and \U$32345 ( \32689 , \32686 , \32688 );
and \U$32346 ( \32690 , \32684 , \32689 );
xor \U$32347 ( \32691 , \32365 , \32367 );
xor \U$32348 ( \32692 , \32691 , \32369 );
and \U$32349 ( \32693 , \32689 , \32692 );
and \U$32350 ( \32694 , \32684 , \32692 );
or \U$32351 ( \32695 , \32690 , \32693 , \32694 );
and \U$32352 ( \32696 , \32383 , \32695 );
xor \U$32353 ( \32697 , \32383 , \32695 );
xor \U$32354 ( \32698 , \32684 , \32689 );
xor \U$32355 ( \32699 , \32698 , \32692 );
and \U$32356 ( \32700 , \27830 , \21985 );
and \U$32357 ( \32701 , \27527 , \21983 );
nor \U$32358 ( \32702 , \32700 , \32701 );
xnor \U$32359 ( \32703 , \32702 , \21907 );
and \U$32360 ( \32704 , \28528 , \21821 );
and \U$32361 ( \32705 , \28002 , \21819 );
nor \U$32362 ( \32706 , \32704 , \32705 );
xnor \U$32363 ( \32707 , \32706 , \21727 );
and \U$32364 ( \32708 , \32703 , \32707 );
and \U$32365 ( \32709 , \29198 , \21652 );
and \U$32366 ( \32710 , \28952 , \21650 );
nor \U$32367 ( \32711 , \32709 , \32710 );
xnor \U$32368 ( \32712 , \32711 , \21377 );
and \U$32369 ( \32713 , \32707 , \32712 );
and \U$32370 ( \32714 , \32703 , \32712 );
or \U$32371 ( \32715 , \32708 , \32713 , \32714 );
and \U$32372 ( \32716 , \25097 , \23421 );
and \U$32373 ( \32717 , \24841 , \23419 );
nor \U$32374 ( \32718 , \32716 , \32717 );
xnor \U$32375 ( \32719 , \32718 , \23279 );
and \U$32376 ( \32720 , \25596 , \23125 );
and \U$32377 ( \32721 , \25294 , \23123 );
nor \U$32378 ( \32722 , \32720 , \32721 );
xnor \U$32379 ( \32723 , \32722 , \22988 );
and \U$32380 ( \32724 , \32719 , \32723 );
and \U$32381 ( \32725 , \26073 , \22919 );
and \U$32382 ( \32726 , \25604 , \22917 );
nor \U$32383 ( \32727 , \32725 , \32726 );
xnor \U$32384 ( \32728 , \32727 , \22767 );
and \U$32385 ( \32729 , \32723 , \32728 );
and \U$32386 ( \32730 , \32719 , \32728 );
or \U$32387 ( \32731 , \32724 , \32729 , \32730 );
and \U$32388 ( \32732 , \32715 , \32731 );
and \U$32389 ( \32733 , \26342 , \22651 );
and \U$32390 ( \32734 , \26078 , \22649 );
nor \U$32391 ( \32735 , \32733 , \32734 );
xnor \U$32392 ( \32736 , \32735 , \22495 );
and \U$32393 ( \32737 , \26973 , \22379 );
and \U$32394 ( \32738 , \26601 , \22377 );
nor \U$32395 ( \32739 , \32737 , \32738 );
xnor \U$32396 ( \32740 , \32739 , \22266 );
and \U$32397 ( \32741 , \32736 , \32740 );
and \U$32398 ( \32742 , \27325 , \22185 );
and \U$32399 ( \32743 , \26982 , \22183 );
nor \U$32400 ( \32744 , \32742 , \32743 );
xnor \U$32401 ( \32745 , \32744 , \22049 );
and \U$32402 ( \32746 , \32740 , \32745 );
and \U$32403 ( \32747 , \32736 , \32745 );
or \U$32404 ( \32748 , \32741 , \32746 , \32747 );
and \U$32405 ( \32749 , \32731 , \32748 );
and \U$32406 ( \32750 , \32715 , \32748 );
or \U$32407 ( \32751 , \32732 , \32749 , \32750 );
and \U$32408 ( \32752 , \21750 , \28592 );
and \U$32409 ( \32753 , \21689 , \28590 );
nor \U$32410 ( \32754 , \32752 , \32753 );
xnor \U$32411 ( \32755 , \32754 , \28343 );
and \U$32412 ( \32756 , \22011 , \28063 );
and \U$32413 ( \32757 , \21813 , \28061 );
nor \U$32414 ( \32758 , \32756 , \32757 );
xnor \U$32415 ( \32759 , \32758 , \27803 );
and \U$32416 ( \32760 , \32755 , \32759 );
and \U$32417 ( \32761 , \22204 , \27569 );
and \U$32418 ( \32762 , \22099 , \27567 );
nor \U$32419 ( \32763 , \32761 , \32762 );
xnor \U$32420 ( \32764 , \32763 , \27254 );
and \U$32421 ( \32765 , \32759 , \32764 );
and \U$32422 ( \32766 , \32755 , \32764 );
or \U$32423 ( \32767 , \32760 , \32765 , \32766 );
and \U$32424 ( \32768 , \21452 , \30258 );
and \U$32425 ( \32769 , \21428 , \30256 );
nor \U$32426 ( \32770 , \32768 , \32769 );
xnor \U$32427 ( \32771 , \32770 , \29948 );
and \U$32428 ( \32772 , \21471 , \29721 );
and \U$32429 ( \32773 , \21444 , \29719 );
nor \U$32430 ( \32774 , \32772 , \32773 );
xnor \U$32431 ( \32775 , \32774 , \29350 );
and \U$32432 ( \32776 , \32771 , \32775 );
and \U$32433 ( \32777 , \21478 , \29159 );
and \U$32434 ( \32778 , \21463 , \29157 );
nor \U$32435 ( \32779 , \32777 , \32778 );
xnor \U$32436 ( \32780 , \32779 , \28841 );
and \U$32437 ( \32781 , \32775 , \32780 );
and \U$32438 ( \32782 , \32771 , \32780 );
or \U$32439 ( \32783 , \32776 , \32781 , \32782 );
and \U$32440 ( \32784 , \32767 , \32783 );
and \U$32441 ( \32785 , \21421 , \31639 );
and \U$32442 ( \32786 , \21395 , \31636 );
nor \U$32443 ( \32787 , \32785 , \32786 );
xnor \U$32444 ( \32788 , \32787 , \30584 );
and \U$32445 ( \32789 , \21436 , \30826 );
and \U$32446 ( \32790 , \21413 , \30824 );
nor \U$32447 ( \32791 , \32789 , \32790 );
xnor \U$32448 ( \32792 , \32791 , \30587 );
and \U$32449 ( \32793 , \32788 , \32792 );
and \U$32450 ( \32794 , \32792 , \21457 );
and \U$32451 ( \32795 , \32788 , \21457 );
or \U$32452 ( \32796 , \32793 , \32794 , \32795 );
and \U$32453 ( \32797 , \32783 , \32796 );
and \U$32454 ( \32798 , \32767 , \32796 );
or \U$32455 ( \32799 , \32784 , \32797 , \32798 );
and \U$32456 ( \32800 , \32751 , \32799 );
and \U$32457 ( \32801 , \22325 , \27060 );
and \U$32458 ( \32802 , \22209 , \27058 );
nor \U$32459 ( \32803 , \32801 , \32802 );
xnor \U$32460 ( \32804 , \32803 , \26720 );
and \U$32461 ( \32805 , \22616 , \26471 );
and \U$32462 ( \32806 , \22440 , \26469 );
nor \U$32463 ( \32807 , \32805 , \32806 );
xnor \U$32464 ( \32808 , \32807 , \26230 );
and \U$32465 ( \32809 , \32804 , \32808 );
and \U$32466 ( \32810 , \22867 , \26005 );
and \U$32467 ( \32811 , \22624 , \26003 );
nor \U$32468 ( \32812 , \32810 , \32811 );
xnor \U$32469 ( \32813 , \32812 , \25817 );
and \U$32470 ( \32814 , \32808 , \32813 );
and \U$32471 ( \32815 , \32804 , \32813 );
or \U$32472 ( \32816 , \32809 , \32814 , \32815 );
and \U$32473 ( \32817 , \23058 , \25631 );
and \U$32474 ( \32818 , \22872 , \25629 );
nor \U$32475 ( \32819 , \32817 , \32818 );
xnor \U$32476 ( \32820 , \32819 , \25399 );
and \U$32477 ( \32821 , \23466 , \25180 );
and \U$32478 ( \32822 , \23202 , \25178 );
nor \U$32479 ( \32823 , \32821 , \32822 );
xnor \U$32480 ( \32824 , \32823 , \25037 );
and \U$32481 ( \32825 , \32820 , \32824 );
and \U$32482 ( \32826 , \23665 , \24857 );
and \U$32483 ( \32827 , \23491 , \24855 );
nor \U$32484 ( \32828 , \32826 , \32827 );
xnor \U$32485 ( \32829 , \32828 , \24611 );
and \U$32486 ( \32830 , \32824 , \32829 );
and \U$32487 ( \32831 , \32820 , \32829 );
or \U$32488 ( \32832 , \32825 , \32830 , \32831 );
and \U$32489 ( \32833 , \32816 , \32832 );
and \U$32490 ( \32834 , \23970 , \24462 );
and \U$32491 ( \32835 , \23832 , \24460 );
nor \U$32492 ( \32836 , \32834 , \32835 );
xnor \U$32493 ( \32837 , \32836 , \24275 );
and \U$32494 ( \32838 , \24506 , \24149 );
and \U$32495 ( \32839 , \24089 , \24147 );
nor \U$32496 ( \32840 , \32838 , \32839 );
xnor \U$32497 ( \32841 , \32840 , \23944 );
and \U$32498 ( \32842 , \32837 , \32841 );
and \U$32499 ( \32843 , \24836 , \23743 );
and \U$32500 ( \32844 , \24714 , \23741 );
nor \U$32501 ( \32845 , \32843 , \32844 );
xnor \U$32502 ( \32846 , \32845 , \23594 );
and \U$32503 ( \32847 , \32841 , \32846 );
and \U$32504 ( \32848 , \32837 , \32846 );
or \U$32505 ( \32849 , \32842 , \32847 , \32848 );
and \U$32506 ( \32850 , \32832 , \32849 );
and \U$32507 ( \32851 , \32816 , \32849 );
or \U$32508 ( \32852 , \32833 , \32850 , \32851 );
and \U$32509 ( \32853 , \32799 , \32852 );
and \U$32510 ( \32854 , \32751 , \32852 );
or \U$32511 ( \32855 , \32800 , \32853 , \32854 );
and \U$32512 ( \32856 , \29522 , \21385 );
and \U$32513 ( \32857 , \29203 , \21383 );
nor \U$32514 ( \32858 , \32856 , \32857 );
xnor \U$32515 ( \32859 , \32858 , \21392 );
and \U$32516 ( \32860 , \30375 , \21401 );
and \U$32517 ( \32861 , \29806 , \21399 );
nor \U$32518 ( \32862 , \32860 , \32861 );
xnor \U$32519 ( \32863 , \32862 , \21408 );
and \U$32520 ( \32864 , \32859 , \32863 );
and \U$32521 ( \32865 , \30986 , \21419 );
and \U$32522 ( \32866 , \30383 , \21417 );
nor \U$32523 ( \32867 , \32865 , \32866 );
xnor \U$32524 ( \32868 , \32867 , \21426 );
and \U$32525 ( \32869 , \32863 , \32868 );
and \U$32526 ( \32870 , \32859 , \32868 );
or \U$32527 ( \32871 , \32864 , \32869 , \32870 );
and \U$32528 ( \32872 , \31172 , \21434 );
and \U$32529 ( \32873 , \30991 , \21432 );
nor \U$32530 ( \32874 , \32872 , \32873 );
xnor \U$32531 ( \32875 , \32874 , \21441 );
nand \U$32532 ( \32876 , \31792 , \21448 );
xnor \U$32533 ( \32877 , \32876 , \21457 );
and \U$32534 ( \32878 , \32875 , \32877 );
and \U$32535 ( \32879 , \32871 , \32878 );
and \U$32536 ( \32880 , \31792 , \21450 );
and \U$32537 ( \32881 , \31172 , \21448 );
nor \U$32538 ( \32882 , \32880 , \32881 );
xnor \U$32539 ( \32883 , \32882 , \21457 );
and \U$32540 ( \32884 , \32878 , \32883 );
and \U$32541 ( \32885 , \32871 , \32883 );
or \U$32542 ( \32886 , \32879 , \32884 , \32885 );
xor \U$32543 ( \32887 , \32472 , \32476 );
xor \U$32544 ( \32888 , \32887 , \32481 );
xor \U$32545 ( \32889 , \32508 , \32512 );
xor \U$32546 ( \32890 , \32889 , \32517 );
and \U$32547 ( \32891 , \32888 , \32890 );
xor \U$32548 ( \32892 , \32525 , \32529 );
xor \U$32549 ( \32893 , \32892 , \32534 );
and \U$32550 ( \32894 , \32890 , \32893 );
and \U$32551 ( \32895 , \32888 , \32893 );
or \U$32552 ( \32896 , \32891 , \32894 , \32895 );
and \U$32553 ( \32897 , \32886 , \32896 );
xor \U$32554 ( \32898 , \32439 , \32443 );
xor \U$32555 ( \32899 , \32898 , \32448 );
xor \U$32556 ( \32900 , \32455 , \32459 );
xor \U$32557 ( \32901 , \32900 , \32464 );
and \U$32558 ( \32902 , \32899 , \32901 );
xor \U$32559 ( \32903 , \32557 , \32561 );
xor \U$32560 ( \32904 , \32903 , \32566 );
and \U$32561 ( \32905 , \32901 , \32904 );
and \U$32562 ( \32906 , \32899 , \32904 );
or \U$32563 ( \32907 , \32902 , \32905 , \32906 );
and \U$32564 ( \32908 , \32896 , \32907 );
and \U$32565 ( \32909 , \32886 , \32907 );
or \U$32566 ( \32910 , \32897 , \32908 , \32909 );
and \U$32567 ( \32911 , \32855 , \32910 );
xor \U$32568 ( \32912 , \32387 , \32391 );
xor \U$32569 ( \32913 , \32912 , \32396 );
xor \U$32570 ( \32914 , \32492 , \32496 );
xor \U$32571 ( \32915 , \32914 , \32501 );
and \U$32572 ( \32916 , \32913 , \32915 );
xor \U$32573 ( \32917 , \32420 , \32424 );
xor \U$32574 ( \32918 , \32917 , \32429 );
and \U$32575 ( \32919 , \32915 , \32918 );
and \U$32576 ( \32920 , \32913 , \32918 );
or \U$32577 ( \32921 , \32916 , \32919 , \32920 );
xor \U$32578 ( \32922 , \32594 , \32596 );
xor \U$32579 ( \32923 , \32922 , \32599 );
and \U$32580 ( \32924 , \32921 , \32923 );
xor \U$32581 ( \32925 , \32545 , \32547 );
xor \U$32582 ( \32926 , \32925 , \32550 );
and \U$32583 ( \32927 , \32923 , \32926 );
and \U$32584 ( \32928 , \32921 , \32926 );
or \U$32585 ( \32929 , \32924 , \32927 , \32928 );
and \U$32586 ( \32930 , \32910 , \32929 );
and \U$32587 ( \32931 , \32855 , \32929 );
or \U$32588 ( \32932 , \32911 , \32930 , \32931 );
xor \U$32589 ( \32933 , \32451 , \32467 );
xor \U$32590 ( \32934 , \32933 , \32484 );
xor \U$32591 ( \32935 , \32569 , \32571 );
xor \U$32592 ( \32936 , \32935 , \32574 );
and \U$32593 ( \32937 , \32934 , \32936 );
xor \U$32594 ( \32938 , \32580 , \32582 );
xor \U$32595 ( \32939 , \32938 , \32585 );
and \U$32596 ( \32940 , \32936 , \32939 );
and \U$32597 ( \32941 , \32934 , \32939 );
or \U$32598 ( \32942 , \32937 , \32940 , \32941 );
xor \U$32599 ( \32943 , \32614 , \32616 );
xor \U$32600 ( \32944 , \32943 , \32619 );
and \U$32601 ( \32945 , \32942 , \32944 );
xor \U$32602 ( \32946 , \32624 , \32626 );
xor \U$32603 ( \32947 , \32946 , \32629 );
and \U$32604 ( \32948 , \32944 , \32947 );
and \U$32605 ( \32949 , \32942 , \32947 );
or \U$32606 ( \32950 , \32945 , \32948 , \32949 );
and \U$32607 ( \32951 , \32932 , \32950 );
xor \U$32608 ( \32952 , \32435 , \32487 );
xor \U$32609 ( \32953 , \32952 , \32540 );
xor \U$32610 ( \32954 , \32553 , \32577 );
xor \U$32611 ( \32955 , \32954 , \32588 );
and \U$32612 ( \32956 , \32953 , \32955 );
xor \U$32613 ( \32957 , \32602 , \32604 );
xor \U$32614 ( \32958 , \32957 , \32606 );
and \U$32615 ( \32959 , \32955 , \32958 );
and \U$32616 ( \32960 , \32953 , \32958 );
or \U$32617 ( \32961 , \32956 , \32959 , \32960 );
and \U$32618 ( \32962 , \32950 , \32961 );
and \U$32619 ( \32963 , \32932 , \32961 );
or \U$32620 ( \32964 , \32951 , \32962 , \32963 );
xor \U$32621 ( \32965 , \32103 , \32115 );
xor \U$32622 ( \32966 , \32965 , \32126 );
xor \U$32623 ( \32967 , \32181 , \32229 );
xor \U$32624 ( \32968 , \32967 , \32282 );
and \U$32625 ( \32969 , \32966 , \32968 );
xor \U$32626 ( \32970 , \32641 , \32643 );
xor \U$32627 ( \32971 , \32970 , \32646 );
and \U$32628 ( \32972 , \32968 , \32971 );
and \U$32629 ( \32973 , \32966 , \32971 );
or \U$32630 ( \32974 , \32969 , \32972 , \32973 );
and \U$32631 ( \32975 , \32964 , \32974 );
xor \U$32632 ( \32976 , \32129 , \32285 );
xor \U$32633 ( \32977 , \32976 , \32306 );
and \U$32634 ( \32978 , \32974 , \32977 );
and \U$32635 ( \32979 , \32964 , \32977 );
or \U$32636 ( \32980 , \32975 , \32978 , \32979 );
xor \U$32637 ( \32981 , \32652 , \32662 );
xor \U$32638 ( \32982 , \32981 , \32665 );
and \U$32639 ( \32983 , \32980 , \32982 );
xor \U$32640 ( \32984 , \32670 , \32672 );
xor \U$32641 ( \32985 , \32984 , \32675 );
and \U$32642 ( \32986 , \32982 , \32985 );
and \U$32643 ( \32987 , \32980 , \32985 );
or \U$32644 ( \32988 , \32983 , \32986 , \32987 );
xor \U$32645 ( \32989 , \32668 , \32678 );
xor \U$32646 ( \32990 , \32989 , \32681 );
and \U$32647 ( \32991 , \32988 , \32990 );
xor \U$32648 ( \32992 , \32686 , \32688 );
and \U$32649 ( \32993 , \32990 , \32992 );
and \U$32650 ( \32994 , \32988 , \32992 );
or \U$32651 ( \32995 , \32991 , \32993 , \32994 );
and \U$32652 ( \32996 , \32699 , \32995 );
xor \U$32653 ( \32997 , \32699 , \32995 );
xor \U$32654 ( \32998 , \32988 , \32990 );
xor \U$32655 ( \32999 , \32998 , \32992 );
xor \U$32656 ( \33000 , \32703 , \32707 );
xor \U$32657 ( \33001 , \33000 , \32712 );
xor \U$32658 ( \33002 , \32719 , \32723 );
xor \U$32659 ( \33003 , \33002 , \32728 );
and \U$32660 ( \33004 , \33001 , \33003 );
xor \U$32661 ( \33005 , \32736 , \32740 );
xor \U$32662 ( \33006 , \33005 , \32745 );
and \U$32663 ( \33007 , \33003 , \33006 );
and \U$32664 ( \33008 , \33001 , \33006 );
or \U$32665 ( \33009 , \33004 , \33007 , \33008 );
xor \U$32666 ( \33010 , \32804 , \32808 );
xor \U$32667 ( \33011 , \33010 , \32813 );
xor \U$32668 ( \33012 , \32820 , \32824 );
xor \U$32669 ( \33013 , \33012 , \32829 );
and \U$32670 ( \33014 , \33011 , \33013 );
xor \U$32671 ( \33015 , \32837 , \32841 );
xor \U$32672 ( \33016 , \33015 , \32846 );
and \U$32673 ( \33017 , \33013 , \33016 );
and \U$32674 ( \33018 , \33011 , \33016 );
or \U$32675 ( \33019 , \33014 , \33017 , \33018 );
and \U$32676 ( \33020 , \33009 , \33019 );
and \U$32677 ( \33021 , \30383 , \21401 );
and \U$32678 ( \33022 , \30375 , \21399 );
nor \U$32679 ( \33023 , \33021 , \33022 );
xnor \U$32680 ( \33024 , \33023 , \21408 );
and \U$32681 ( \33025 , \30991 , \21419 );
and \U$32682 ( \33026 , \30986 , \21417 );
nor \U$32683 ( \33027 , \33025 , \33026 );
xnor \U$32684 ( \33028 , \33027 , \21426 );
and \U$32685 ( \33029 , \33024 , \33028 );
and \U$32686 ( \33030 , \31792 , \21434 );
and \U$32687 ( \33031 , \31172 , \21432 );
nor \U$32688 ( \33032 , \33030 , \33031 );
xnor \U$32689 ( \33033 , \33032 , \21441 );
and \U$32690 ( \33034 , \33028 , \33033 );
and \U$32691 ( \33035 , \33024 , \33033 );
or \U$32692 ( \33036 , \33029 , \33034 , \33035 );
xor \U$32693 ( \33037 , \32859 , \32863 );
xor \U$32694 ( \33038 , \33037 , \32868 );
and \U$32695 ( \33039 , \33036 , \33038 );
xor \U$32696 ( \33040 , \32875 , \32877 );
and \U$32697 ( \33041 , \33038 , \33040 );
and \U$32698 ( \33042 , \33036 , \33040 );
or \U$32699 ( \33043 , \33039 , \33041 , \33042 );
and \U$32700 ( \33044 , \33019 , \33043 );
and \U$32701 ( \33045 , \33009 , \33043 );
or \U$32702 ( \33046 , \33020 , \33044 , \33045 );
and \U$32703 ( \33047 , \24714 , \24149 );
and \U$32704 ( \33048 , \24506 , \24147 );
nor \U$32705 ( \33049 , \33047 , \33048 );
xnor \U$32706 ( \33050 , \33049 , \23944 );
and \U$32707 ( \33051 , \24841 , \23743 );
and \U$32708 ( \33052 , \24836 , \23741 );
nor \U$32709 ( \33053 , \33051 , \33052 );
xnor \U$32710 ( \33054 , \33053 , \23594 );
and \U$32711 ( \33055 , \33050 , \33054 );
and \U$32712 ( \33056 , \25294 , \23421 );
and \U$32713 ( \33057 , \25097 , \23419 );
nor \U$32714 ( \33058 , \33056 , \33057 );
xnor \U$32715 ( \33059 , \33058 , \23279 );
and \U$32716 ( \33060 , \33054 , \33059 );
and \U$32717 ( \33061 , \33050 , \33059 );
or \U$32718 ( \33062 , \33055 , \33060 , \33061 );
and \U$32719 ( \33063 , \22624 , \26471 );
and \U$32720 ( \33064 , \22616 , \26469 );
nor \U$32721 ( \33065 , \33063 , \33064 );
xnor \U$32722 ( \33066 , \33065 , \26230 );
and \U$32723 ( \33067 , \22872 , \26005 );
and \U$32724 ( \33068 , \22867 , \26003 );
nor \U$32725 ( \33069 , \33067 , \33068 );
xnor \U$32726 ( \33070 , \33069 , \25817 );
and \U$32727 ( \33071 , \33066 , \33070 );
and \U$32728 ( \33072 , \23202 , \25631 );
and \U$32729 ( \33073 , \23058 , \25629 );
nor \U$32730 ( \33074 , \33072 , \33073 );
xnor \U$32731 ( \33075 , \33074 , \25399 );
and \U$32732 ( \33076 , \33070 , \33075 );
and \U$32733 ( \33077 , \33066 , \33075 );
or \U$32734 ( \33078 , \33071 , \33076 , \33077 );
and \U$32735 ( \33079 , \33062 , \33078 );
and \U$32736 ( \33080 , \23491 , \25180 );
and \U$32737 ( \33081 , \23466 , \25178 );
nor \U$32738 ( \33082 , \33080 , \33081 );
xnor \U$32739 ( \33083 , \33082 , \25037 );
and \U$32740 ( \33084 , \23832 , \24857 );
and \U$32741 ( \33085 , \23665 , \24855 );
nor \U$32742 ( \33086 , \33084 , \33085 );
xnor \U$32743 ( \33087 , \33086 , \24611 );
and \U$32744 ( \33088 , \33083 , \33087 );
and \U$32745 ( \33089 , \24089 , \24462 );
and \U$32746 ( \33090 , \23970 , \24460 );
nor \U$32747 ( \33091 , \33089 , \33090 );
xnor \U$32748 ( \33092 , \33091 , \24275 );
and \U$32749 ( \33093 , \33087 , \33092 );
and \U$32750 ( \33094 , \33083 , \33092 );
or \U$32751 ( \33095 , \33088 , \33093 , \33094 );
and \U$32752 ( \33096 , \33078 , \33095 );
and \U$32753 ( \33097 , \33062 , \33095 );
or \U$32754 ( \33098 , \33079 , \33096 , \33097 );
and \U$32755 ( \33099 , \22099 , \28063 );
and \U$32756 ( \33100 , \22011 , \28061 );
nor \U$32757 ( \33101 , \33099 , \33100 );
xnor \U$32758 ( \33102 , \33101 , \27803 );
and \U$32759 ( \33103 , \22209 , \27569 );
and \U$32760 ( \33104 , \22204 , \27567 );
nor \U$32761 ( \33105 , \33103 , \33104 );
xnor \U$32762 ( \33106 , \33105 , \27254 );
and \U$32763 ( \33107 , \33102 , \33106 );
and \U$32764 ( \33108 , \22440 , \27060 );
and \U$32765 ( \33109 , \22325 , \27058 );
nor \U$32766 ( \33110 , \33108 , \33109 );
xnor \U$32767 ( \33111 , \33110 , \26720 );
and \U$32768 ( \33112 , \33106 , \33111 );
and \U$32769 ( \33113 , \33102 , \33111 );
or \U$32770 ( \33114 , \33107 , \33112 , \33113 );
and \U$32771 ( \33115 , \21413 , \31639 );
and \U$32772 ( \33116 , \21421 , \31636 );
nor \U$32773 ( \33117 , \33115 , \33116 );
xnor \U$32774 ( \33118 , \33117 , \30584 );
and \U$32775 ( \33119 , \21428 , \30826 );
and \U$32776 ( \33120 , \21436 , \30824 );
nor \U$32777 ( \33121 , \33119 , \33120 );
xnor \U$32778 ( \33122 , \33121 , \30587 );
and \U$32779 ( \33123 , \33118 , \33122 );
and \U$32780 ( \33124 , \21444 , \30258 );
and \U$32781 ( \33125 , \21452 , \30256 );
nor \U$32782 ( \33126 , \33124 , \33125 );
xnor \U$32783 ( \33127 , \33126 , \29948 );
and \U$32784 ( \33128 , \33122 , \33127 );
and \U$32785 ( \33129 , \33118 , \33127 );
or \U$32786 ( \33130 , \33123 , \33128 , \33129 );
and \U$32787 ( \33131 , \33114 , \33130 );
and \U$32788 ( \33132 , \21463 , \29721 );
and \U$32789 ( \33133 , \21471 , \29719 );
nor \U$32790 ( \33134 , \33132 , \33133 );
xnor \U$32791 ( \33135 , \33134 , \29350 );
and \U$32792 ( \33136 , \21689 , \29159 );
and \U$32793 ( \33137 , \21478 , \29157 );
nor \U$32794 ( \33138 , \33136 , \33137 );
xnor \U$32795 ( \33139 , \33138 , \28841 );
and \U$32796 ( \33140 , \33135 , \33139 );
and \U$32797 ( \33141 , \21813 , \28592 );
and \U$32798 ( \33142 , \21750 , \28590 );
nor \U$32799 ( \33143 , \33141 , \33142 );
xnor \U$32800 ( \33144 , \33143 , \28343 );
and \U$32801 ( \33145 , \33139 , \33144 );
and \U$32802 ( \33146 , \33135 , \33144 );
or \U$32803 ( \33147 , \33140 , \33145 , \33146 );
and \U$32804 ( \33148 , \33130 , \33147 );
and \U$32805 ( \33149 , \33114 , \33147 );
or \U$32806 ( \33150 , \33131 , \33148 , \33149 );
and \U$32807 ( \33151 , \33098 , \33150 );
and \U$32808 ( \33152 , \25604 , \23125 );
and \U$32809 ( \33153 , \25596 , \23123 );
nor \U$32810 ( \33154 , \33152 , \33153 );
xnor \U$32811 ( \33155 , \33154 , \22988 );
and \U$32812 ( \33156 , \26078 , \22919 );
and \U$32813 ( \33157 , \26073 , \22917 );
nor \U$32814 ( \33158 , \33156 , \33157 );
xnor \U$32815 ( \33159 , \33158 , \22767 );
and \U$32816 ( \33160 , \33155 , \33159 );
and \U$32817 ( \33161 , \26601 , \22651 );
and \U$32818 ( \33162 , \26342 , \22649 );
nor \U$32819 ( \33163 , \33161 , \33162 );
xnor \U$32820 ( \33164 , \33163 , \22495 );
and \U$32821 ( \33165 , \33159 , \33164 );
and \U$32822 ( \33166 , \33155 , \33164 );
or \U$32823 ( \33167 , \33160 , \33165 , \33166 );
and \U$32824 ( \33168 , \28952 , \21821 );
and \U$32825 ( \33169 , \28528 , \21819 );
nor \U$32826 ( \33170 , \33168 , \33169 );
xnor \U$32827 ( \33171 , \33170 , \21727 );
and \U$32828 ( \33172 , \29203 , \21652 );
and \U$32829 ( \33173 , \29198 , \21650 );
nor \U$32830 ( \33174 , \33172 , \33173 );
xnor \U$32831 ( \33175 , \33174 , \21377 );
and \U$32832 ( \33176 , \33171 , \33175 );
and \U$32833 ( \33177 , \29806 , \21385 );
and \U$32834 ( \33178 , \29522 , \21383 );
nor \U$32835 ( \33179 , \33177 , \33178 );
xnor \U$32836 ( \33180 , \33179 , \21392 );
and \U$32837 ( \33181 , \33175 , \33180 );
and \U$32838 ( \33182 , \33171 , \33180 );
or \U$32839 ( \33183 , \33176 , \33181 , \33182 );
and \U$32840 ( \33184 , \33167 , \33183 );
and \U$32841 ( \33185 , \26982 , \22379 );
and \U$32842 ( \33186 , \26973 , \22377 );
nor \U$32843 ( \33187 , \33185 , \33186 );
xnor \U$32844 ( \33188 , \33187 , \22266 );
and \U$32845 ( \33189 , \27527 , \22185 );
and \U$32846 ( \33190 , \27325 , \22183 );
nor \U$32847 ( \33191 , \33189 , \33190 );
xnor \U$32848 ( \33192 , \33191 , \22049 );
and \U$32849 ( \33193 , \33188 , \33192 );
and \U$32850 ( \33194 , \28002 , \21985 );
and \U$32851 ( \33195 , \27830 , \21983 );
nor \U$32852 ( \33196 , \33194 , \33195 );
xnor \U$32853 ( \33197 , \33196 , \21907 );
and \U$32854 ( \33198 , \33192 , \33197 );
and \U$32855 ( \33199 , \33188 , \33197 );
or \U$32856 ( \33200 , \33193 , \33198 , \33199 );
and \U$32857 ( \33201 , \33183 , \33200 );
and \U$32858 ( \33202 , \33167 , \33200 );
or \U$32859 ( \33203 , \33184 , \33201 , \33202 );
and \U$32860 ( \33204 , \33150 , \33203 );
and \U$32861 ( \33205 , \33098 , \33203 );
or \U$32862 ( \33206 , \33151 , \33204 , \33205 );
and \U$32863 ( \33207 , \33046 , \33206 );
xor \U$32864 ( \33208 , \32755 , \32759 );
xor \U$32865 ( \33209 , \33208 , \32764 );
xor \U$32866 ( \33210 , \32771 , \32775 );
xor \U$32867 ( \33211 , \33210 , \32780 );
and \U$32868 ( \33212 , \33209 , \33211 );
xor \U$32869 ( \33213 , \32788 , \32792 );
xor \U$32870 ( \33214 , \33213 , \21457 );
and \U$32871 ( \33215 , \33211 , \33214 );
and \U$32872 ( \33216 , \33209 , \33214 );
or \U$32873 ( \33217 , \33212 , \33215 , \33216 );
xor \U$32874 ( \33218 , \32403 , \32407 );
xor \U$32875 ( \33219 , \33218 , \32412 );
and \U$32876 ( \33220 , \33217 , \33219 );
xor \U$32877 ( \33221 , \32913 , \32915 );
xor \U$32878 ( \33222 , \33221 , \32918 );
and \U$32879 ( \33223 , \33219 , \33222 );
and \U$32880 ( \33224 , \33217 , \33222 );
or \U$32881 ( \33225 , \33220 , \33223 , \33224 );
and \U$32882 ( \33226 , \33206 , \33225 );
and \U$32883 ( \33227 , \33046 , \33225 );
or \U$32884 ( \33228 , \33207 , \33226 , \33227 );
xor \U$32885 ( \33229 , \32715 , \32731 );
xor \U$32886 ( \33230 , \33229 , \32748 );
xor \U$32887 ( \33231 , \32767 , \32783 );
xor \U$32888 ( \33232 , \33231 , \32796 );
and \U$32889 ( \33233 , \33230 , \33232 );
xor \U$32890 ( \33234 , \32816 , \32832 );
xor \U$32891 ( \33235 , \33234 , \32849 );
and \U$32892 ( \33236 , \33232 , \33235 );
and \U$32893 ( \33237 , \33230 , \33235 );
or \U$32894 ( \33238 , \33233 , \33236 , \33237 );
xor \U$32895 ( \33239 , \32871 , \32878 );
xor \U$32896 ( \33240 , \33239 , \32883 );
xor \U$32897 ( \33241 , \32888 , \32890 );
xor \U$32898 ( \33242 , \33241 , \32893 );
and \U$32899 ( \33243 , \33240 , \33242 );
xor \U$32900 ( \33244 , \32899 , \32901 );
xor \U$32901 ( \33245 , \33244 , \32904 );
and \U$32902 ( \33246 , \33242 , \33245 );
and \U$32903 ( \33247 , \33240 , \33245 );
or \U$32904 ( \33248 , \33243 , \33246 , \33247 );
and \U$32905 ( \33249 , \33238 , \33248 );
xor \U$32906 ( \33250 , \32504 , \32520 );
xor \U$32907 ( \33251 , \33250 , \32537 );
and \U$32908 ( \33252 , \33248 , \33251 );
and \U$32909 ( \33253 , \33238 , \33251 );
or \U$32910 ( \33254 , \33249 , \33252 , \33253 );
and \U$32911 ( \33255 , \33228 , \33254 );
xor \U$32912 ( \33256 , \32399 , \32415 );
xor \U$32913 ( \33257 , \33256 , \32432 );
xor \U$32914 ( \33258 , \32934 , \32936 );
xor \U$32915 ( \33259 , \33258 , \32939 );
and \U$32916 ( \33260 , \33257 , \33259 );
xor \U$32917 ( \33261 , \32921 , \32923 );
xor \U$32918 ( \33262 , \33261 , \32926 );
and \U$32919 ( \33263 , \33259 , \33262 );
and \U$32920 ( \33264 , \33257 , \33262 );
or \U$32921 ( \33265 , \33260 , \33263 , \33264 );
and \U$32922 ( \33266 , \33254 , \33265 );
and \U$32923 ( \33267 , \33228 , \33265 );
or \U$32924 ( \33268 , \33255 , \33266 , \33267 );
xor \U$32925 ( \33269 , \32855 , \32910 );
xor \U$32926 ( \33270 , \33269 , \32929 );
xor \U$32927 ( \33271 , \32942 , \32944 );
xor \U$32928 ( \33272 , \33271 , \32947 );
and \U$32929 ( \33273 , \33270 , \33272 );
xor \U$32930 ( \33274 , \32953 , \32955 );
xor \U$32931 ( \33275 , \33274 , \32958 );
and \U$32932 ( \33276 , \33272 , \33275 );
and \U$32933 ( \33277 , \33270 , \33275 );
or \U$32934 ( \33278 , \33273 , \33276 , \33277 );
and \U$32935 ( \33279 , \33268 , \33278 );
xor \U$32936 ( \33280 , \32622 , \32632 );
xor \U$32937 ( \33281 , \33280 , \32635 );
and \U$32938 ( \33282 , \33278 , \33281 );
and \U$32939 ( \33283 , \33268 , \33281 );
or \U$32940 ( \33284 , \33279 , \33282 , \33283 );
xor \U$32941 ( \33285 , \32543 , \32591 );
xor \U$32942 ( \33286 , \33285 , \32609 );
xor \U$32943 ( \33287 , \32932 , \32950 );
xor \U$32944 ( \33288 , \33287 , \32961 );
and \U$32945 ( \33289 , \33286 , \33288 );
xor \U$32946 ( \33290 , \32966 , \32968 );
xor \U$32947 ( \33291 , \33290 , \32971 );
and \U$32948 ( \33292 , \33288 , \33291 );
and \U$32949 ( \33293 , \33286 , \33291 );
or \U$32950 ( \33294 , \33289 , \33292 , \33293 );
and \U$32951 ( \33295 , \33284 , \33294 );
xor \U$32952 ( \33296 , \32654 , \32656 );
xor \U$32953 ( \33297 , \33296 , \32659 );
and \U$32954 ( \33298 , \33294 , \33297 );
and \U$32955 ( \33299 , \33284 , \33297 );
or \U$32956 ( \33300 , \33295 , \33298 , \33299 );
xor \U$32957 ( \33301 , \32612 , \32638 );
xor \U$32958 ( \33302 , \33301 , \32649 );
xor \U$32959 ( \33303 , \32964 , \32974 );
xor \U$32960 ( \33304 , \33303 , \32977 );
and \U$32961 ( \33305 , \33302 , \33304 );
and \U$32962 ( \33306 , \33300 , \33305 );
xor \U$32963 ( \33307 , \32980 , \32982 );
xor \U$32964 ( \33308 , \33307 , \32985 );
and \U$32965 ( \33309 , \33305 , \33308 );
and \U$32966 ( \33310 , \33300 , \33308 );
or \U$32967 ( \33311 , \33306 , \33309 , \33310 );
and \U$32968 ( \33312 , \32999 , \33311 );
xor \U$32969 ( \33313 , \32999 , \33311 );
xor \U$32970 ( \33314 , \33300 , \33305 );
xor \U$32971 ( \33315 , \33314 , \33308 );
xor \U$32972 ( \33316 , \33050 , \33054 );
xor \U$32973 ( \33317 , \33316 , \33059 );
xor \U$32974 ( \33318 , \33155 , \33159 );
xor \U$32975 ( \33319 , \33318 , \33164 );
and \U$32976 ( \33320 , \33317 , \33319 );
xor \U$32977 ( \33321 , \33188 , \33192 );
xor \U$32978 ( \33322 , \33321 , \33197 );
and \U$32979 ( \33323 , \33319 , \33322 );
and \U$32980 ( \33324 , \33317 , \33322 );
or \U$32981 ( \33325 , \33320 , \33323 , \33324 );
and \U$32982 ( \33326 , \30375 , \21385 );
and \U$32983 ( \33327 , \29806 , \21383 );
nor \U$32984 ( \33328 , \33326 , \33327 );
xnor \U$32985 ( \33329 , \33328 , \21392 );
and \U$32986 ( \33330 , \30986 , \21401 );
and \U$32987 ( \33331 , \30383 , \21399 );
nor \U$32988 ( \33332 , \33330 , \33331 );
xnor \U$32989 ( \33333 , \33332 , \21408 );
and \U$32990 ( \33334 , \33329 , \33333 );
and \U$32991 ( \33335 , \31172 , \21419 );
and \U$32992 ( \33336 , \30991 , \21417 );
nor \U$32993 ( \33337 , \33335 , \33336 );
xnor \U$32994 ( \33338 , \33337 , \21426 );
and \U$32995 ( \33339 , \33333 , \33338 );
and \U$32996 ( \33340 , \33329 , \33338 );
or \U$32997 ( \33341 , \33334 , \33339 , \33340 );
xor \U$32998 ( \33342 , \33171 , \33175 );
xor \U$32999 ( \33343 , \33342 , \33180 );
and \U$33000 ( \33344 , \33341 , \33343 );
xor \U$33001 ( \33345 , \33024 , \33028 );
xor \U$33002 ( \33346 , \33345 , \33033 );
and \U$33003 ( \33347 , \33343 , \33346 );
and \U$33004 ( \33348 , \33341 , \33346 );
or \U$33005 ( \33349 , \33344 , \33347 , \33348 );
and \U$33006 ( \33350 , \33325 , \33349 );
xor \U$33007 ( \33351 , \33102 , \33106 );
xor \U$33008 ( \33352 , \33351 , \33111 );
xor \U$33009 ( \33353 , \33066 , \33070 );
xor \U$33010 ( \33354 , \33353 , \33075 );
and \U$33011 ( \33355 , \33352 , \33354 );
xor \U$33012 ( \33356 , \33083 , \33087 );
xor \U$33013 ( \33357 , \33356 , \33092 );
and \U$33014 ( \33358 , \33354 , \33357 );
and \U$33015 ( \33359 , \33352 , \33357 );
or \U$33016 ( \33360 , \33355 , \33358 , \33359 );
and \U$33017 ( \33361 , \33349 , \33360 );
and \U$33018 ( \33362 , \33325 , \33360 );
or \U$33019 ( \33363 , \33350 , \33361 , \33362 );
and \U$33020 ( \33364 , \22011 , \28592 );
and \U$33021 ( \33365 , \21813 , \28590 );
nor \U$33022 ( \33366 , \33364 , \33365 );
xnor \U$33023 ( \33367 , \33366 , \28343 );
and \U$33024 ( \33368 , \22204 , \28063 );
and \U$33025 ( \33369 , \22099 , \28061 );
nor \U$33026 ( \33370 , \33368 , \33369 );
xnor \U$33027 ( \33371 , \33370 , \27803 );
and \U$33028 ( \33372 , \33367 , \33371 );
and \U$33029 ( \33373 , \22325 , \27569 );
and \U$33030 ( \33374 , \22209 , \27567 );
nor \U$33031 ( \33375 , \33373 , \33374 );
xnor \U$33032 ( \33376 , \33375 , \27254 );
and \U$33033 ( \33377 , \33371 , \33376 );
and \U$33034 ( \33378 , \33367 , \33376 );
or \U$33035 ( \33379 , \33372 , \33377 , \33378 );
and \U$33036 ( \33380 , \21436 , \31639 );
and \U$33037 ( \33381 , \21413 , \31636 );
nor \U$33038 ( \33382 , \33380 , \33381 );
xnor \U$33039 ( \33383 , \33382 , \30584 );
and \U$33040 ( \33384 , \21452 , \30826 );
and \U$33041 ( \33385 , \21428 , \30824 );
nor \U$33042 ( \33386 , \33384 , \33385 );
xnor \U$33043 ( \33387 , \33386 , \30587 );
and \U$33044 ( \33388 , \33383 , \33387 );
and \U$33045 ( \33389 , \33387 , \21441 );
and \U$33046 ( \33390 , \33383 , \21441 );
or \U$33047 ( \33391 , \33388 , \33389 , \33390 );
and \U$33048 ( \33392 , \33379 , \33391 );
and \U$33049 ( \33393 , \21471 , \30258 );
and \U$33050 ( \33394 , \21444 , \30256 );
nor \U$33051 ( \33395 , \33393 , \33394 );
xnor \U$33052 ( \33396 , \33395 , \29948 );
and \U$33053 ( \33397 , \21478 , \29721 );
and \U$33054 ( \33398 , \21463 , \29719 );
nor \U$33055 ( \33399 , \33397 , \33398 );
xnor \U$33056 ( \33400 , \33399 , \29350 );
and \U$33057 ( \33401 , \33396 , \33400 );
and \U$33058 ( \33402 , \21750 , \29159 );
and \U$33059 ( \33403 , \21689 , \29157 );
nor \U$33060 ( \33404 , \33402 , \33403 );
xnor \U$33061 ( \33405 , \33404 , \28841 );
and \U$33062 ( \33406 , \33400 , \33405 );
and \U$33063 ( \33407 , \33396 , \33405 );
or \U$33064 ( \33408 , \33401 , \33406 , \33407 );
and \U$33065 ( \33409 , \33391 , \33408 );
and \U$33066 ( \33410 , \33379 , \33408 );
or \U$33067 ( \33411 , \33392 , \33409 , \33410 );
and \U$33068 ( \33412 , \24506 , \24462 );
and \U$33069 ( \33413 , \24089 , \24460 );
nor \U$33070 ( \33414 , \33412 , \33413 );
xnor \U$33071 ( \33415 , \33414 , \24275 );
and \U$33072 ( \33416 , \24836 , \24149 );
and \U$33073 ( \33417 , \24714 , \24147 );
nor \U$33074 ( \33418 , \33416 , \33417 );
xnor \U$33075 ( \33419 , \33418 , \23944 );
and \U$33076 ( \33420 , \33415 , \33419 );
and \U$33077 ( \33421 , \25097 , \23743 );
and \U$33078 ( \33422 , \24841 , \23741 );
nor \U$33079 ( \33423 , \33421 , \33422 );
xnor \U$33080 ( \33424 , \33423 , \23594 );
and \U$33081 ( \33425 , \33419 , \33424 );
and \U$33082 ( \33426 , \33415 , \33424 );
or \U$33083 ( \33427 , \33420 , \33425 , \33426 );
and \U$33084 ( \33428 , \23466 , \25631 );
and \U$33085 ( \33429 , \23202 , \25629 );
nor \U$33086 ( \33430 , \33428 , \33429 );
xnor \U$33087 ( \33431 , \33430 , \25399 );
and \U$33088 ( \33432 , \23665 , \25180 );
and \U$33089 ( \33433 , \23491 , \25178 );
nor \U$33090 ( \33434 , \33432 , \33433 );
xnor \U$33091 ( \33435 , \33434 , \25037 );
and \U$33092 ( \33436 , \33431 , \33435 );
and \U$33093 ( \33437 , \23970 , \24857 );
and \U$33094 ( \33438 , \23832 , \24855 );
nor \U$33095 ( \33439 , \33437 , \33438 );
xnor \U$33096 ( \33440 , \33439 , \24611 );
and \U$33097 ( \33441 , \33435 , \33440 );
and \U$33098 ( \33442 , \33431 , \33440 );
or \U$33099 ( \33443 , \33436 , \33441 , \33442 );
and \U$33100 ( \33444 , \33427 , \33443 );
and \U$33101 ( \33445 , \22616 , \27060 );
and \U$33102 ( \33446 , \22440 , \27058 );
nor \U$33103 ( \33447 , \33445 , \33446 );
xnor \U$33104 ( \33448 , \33447 , \26720 );
and \U$33105 ( \33449 , \22867 , \26471 );
and \U$33106 ( \33450 , \22624 , \26469 );
nor \U$33107 ( \33451 , \33449 , \33450 );
xnor \U$33108 ( \33452 , \33451 , \26230 );
and \U$33109 ( \33453 , \33448 , \33452 );
and \U$33110 ( \33454 , \23058 , \26005 );
and \U$33111 ( \33455 , \22872 , \26003 );
nor \U$33112 ( \33456 , \33454 , \33455 );
xnor \U$33113 ( \33457 , \33456 , \25817 );
and \U$33114 ( \33458 , \33452 , \33457 );
and \U$33115 ( \33459 , \33448 , \33457 );
or \U$33116 ( \33460 , \33453 , \33458 , \33459 );
and \U$33117 ( \33461 , \33443 , \33460 );
and \U$33118 ( \33462 , \33427 , \33460 );
or \U$33119 ( \33463 , \33444 , \33461 , \33462 );
and \U$33120 ( \33464 , \33411 , \33463 );
and \U$33121 ( \33465 , \25596 , \23421 );
and \U$33122 ( \33466 , \25294 , \23419 );
nor \U$33123 ( \33467 , \33465 , \33466 );
xnor \U$33124 ( \33468 , \33467 , \23279 );
and \U$33125 ( \33469 , \26073 , \23125 );
and \U$33126 ( \33470 , \25604 , \23123 );
nor \U$33127 ( \33471 , \33469 , \33470 );
xnor \U$33128 ( \33472 , \33471 , \22988 );
and \U$33129 ( \33473 , \33468 , \33472 );
and \U$33130 ( \33474 , \26342 , \22919 );
and \U$33131 ( \33475 , \26078 , \22917 );
nor \U$33132 ( \33476 , \33474 , \33475 );
xnor \U$33133 ( \33477 , \33476 , \22767 );
and \U$33134 ( \33478 , \33472 , \33477 );
and \U$33135 ( \33479 , \33468 , \33477 );
or \U$33136 ( \33480 , \33473 , \33478 , \33479 );
and \U$33137 ( \33481 , \26973 , \22651 );
and \U$33138 ( \33482 , \26601 , \22649 );
nor \U$33139 ( \33483 , \33481 , \33482 );
xnor \U$33140 ( \33484 , \33483 , \22495 );
and \U$33141 ( \33485 , \27325 , \22379 );
and \U$33142 ( \33486 , \26982 , \22377 );
nor \U$33143 ( \33487 , \33485 , \33486 );
xnor \U$33144 ( \33488 , \33487 , \22266 );
and \U$33145 ( \33489 , \33484 , \33488 );
and \U$33146 ( \33490 , \27830 , \22185 );
and \U$33147 ( \33491 , \27527 , \22183 );
nor \U$33148 ( \33492 , \33490 , \33491 );
xnor \U$33149 ( \33493 , \33492 , \22049 );
and \U$33150 ( \33494 , \33488 , \33493 );
and \U$33151 ( \33495 , \33484 , \33493 );
or \U$33152 ( \33496 , \33489 , \33494 , \33495 );
and \U$33153 ( \33497 , \33480 , \33496 );
and \U$33154 ( \33498 , \28528 , \21985 );
and \U$33155 ( \33499 , \28002 , \21983 );
nor \U$33156 ( \33500 , \33498 , \33499 );
xnor \U$33157 ( \33501 , \33500 , \21907 );
and \U$33158 ( \33502 , \29198 , \21821 );
and \U$33159 ( \33503 , \28952 , \21819 );
nor \U$33160 ( \33504 , \33502 , \33503 );
xnor \U$33161 ( \33505 , \33504 , \21727 );
and \U$33162 ( \33506 , \33501 , \33505 );
and \U$33163 ( \33507 , \29522 , \21652 );
and \U$33164 ( \33508 , \29203 , \21650 );
nor \U$33165 ( \33509 , \33507 , \33508 );
xnor \U$33166 ( \33510 , \33509 , \21377 );
and \U$33167 ( \33511 , \33505 , \33510 );
and \U$33168 ( \33512 , \33501 , \33510 );
or \U$33169 ( \33513 , \33506 , \33511 , \33512 );
and \U$33170 ( \33514 , \33496 , \33513 );
and \U$33171 ( \33515 , \33480 , \33513 );
or \U$33172 ( \33516 , \33497 , \33514 , \33515 );
and \U$33173 ( \33517 , \33463 , \33516 );
and \U$33174 ( \33518 , \33411 , \33516 );
or \U$33175 ( \33519 , \33464 , \33517 , \33518 );
and \U$33176 ( \33520 , \33363 , \33519 );
xor \U$33177 ( \33521 , \33209 , \33211 );
xor \U$33178 ( \33522 , \33521 , \33214 );
xor \U$33179 ( \33523 , \33001 , \33003 );
xor \U$33180 ( \33524 , \33523 , \33006 );
and \U$33181 ( \33525 , \33522 , \33524 );
xor \U$33182 ( \33526 , \33011 , \33013 );
xor \U$33183 ( \33527 , \33526 , \33016 );
and \U$33184 ( \33528 , \33524 , \33527 );
and \U$33185 ( \33529 , \33522 , \33527 );
or \U$33186 ( \33530 , \33525 , \33528 , \33529 );
and \U$33187 ( \33531 , \33519 , \33530 );
and \U$33188 ( \33532 , \33363 , \33530 );
or \U$33189 ( \33533 , \33520 , \33531 , \33532 );
xor \U$33190 ( \33534 , \33062 , \33078 );
xor \U$33191 ( \33535 , \33534 , \33095 );
xor \U$33192 ( \33536 , \33167 , \33183 );
xor \U$33193 ( \33537 , \33536 , \33200 );
and \U$33194 ( \33538 , \33535 , \33537 );
xor \U$33195 ( \33539 , \33036 , \33038 );
xor \U$33196 ( \33540 , \33539 , \33040 );
and \U$33197 ( \33541 , \33537 , \33540 );
and \U$33198 ( \33542 , \33535 , \33540 );
or \U$33199 ( \33543 , \33538 , \33541 , \33542 );
xor \U$33200 ( \33544 , \33230 , \33232 );
xor \U$33201 ( \33545 , \33544 , \33235 );
and \U$33202 ( \33546 , \33543 , \33545 );
xor \U$33203 ( \33547 , \33240 , \33242 );
xor \U$33204 ( \33548 , \33547 , \33245 );
and \U$33205 ( \33549 , \33545 , \33548 );
and \U$33206 ( \33550 , \33543 , \33548 );
or \U$33207 ( \33551 , \33546 , \33549 , \33550 );
and \U$33208 ( \33552 , \33533 , \33551 );
xor \U$33209 ( \33553 , \33009 , \33019 );
xor \U$33210 ( \33554 , \33553 , \33043 );
xor \U$33211 ( \33555 , \33098 , \33150 );
xor \U$33212 ( \33556 , \33555 , \33203 );
and \U$33213 ( \33557 , \33554 , \33556 );
xor \U$33214 ( \33558 , \33217 , \33219 );
xor \U$33215 ( \33559 , \33558 , \33222 );
and \U$33216 ( \33560 , \33556 , \33559 );
and \U$33217 ( \33561 , \33554 , \33559 );
or \U$33218 ( \33562 , \33557 , \33560 , \33561 );
and \U$33219 ( \33563 , \33551 , \33562 );
and \U$33220 ( \33564 , \33533 , \33562 );
or \U$33221 ( \33565 , \33552 , \33563 , \33564 );
xor \U$33222 ( \33566 , \32751 , \32799 );
xor \U$33223 ( \33567 , \33566 , \32852 );
xor \U$33224 ( \33568 , \32886 , \32896 );
xor \U$33225 ( \33569 , \33568 , \32907 );
and \U$33226 ( \33570 , \33567 , \33569 );
xor \U$33227 ( \33571 , \33257 , \33259 );
xor \U$33228 ( \33572 , \33571 , \33262 );
and \U$33229 ( \33573 , \33569 , \33572 );
and \U$33230 ( \33574 , \33567 , \33572 );
or \U$33231 ( \33575 , \33570 , \33573 , \33574 );
and \U$33232 ( \33576 , \33565 , \33575 );
xor \U$33233 ( \33577 , \33270 , \33272 );
xor \U$33234 ( \33578 , \33577 , \33275 );
and \U$33235 ( \33579 , \33575 , \33578 );
and \U$33236 ( \33580 , \33565 , \33578 );
or \U$33237 ( \33581 , \33576 , \33579 , \33580 );
xor \U$33238 ( \33582 , \33268 , \33278 );
xor \U$33239 ( \33583 , \33582 , \33281 );
and \U$33240 ( \33584 , \33581 , \33583 );
xor \U$33241 ( \33585 , \33286 , \33288 );
xor \U$33242 ( \33586 , \33585 , \33291 );
and \U$33243 ( \33587 , \33583 , \33586 );
and \U$33244 ( \33588 , \33581 , \33586 );
or \U$33245 ( \33589 , \33584 , \33587 , \33588 );
xor \U$33246 ( \33590 , \33284 , \33294 );
xor \U$33247 ( \33591 , \33590 , \33297 );
and \U$33248 ( \33592 , \33589 , \33591 );
xor \U$33249 ( \33593 , \33302 , \33304 );
and \U$33250 ( \33594 , \33591 , \33593 );
and \U$33251 ( \33595 , \33589 , \33593 );
or \U$33252 ( \33596 , \33592 , \33594 , \33595 );
and \U$33253 ( \33597 , \33315 , \33596 );
xor \U$33254 ( \33598 , \33315 , \33596 );
xor \U$33255 ( \33599 , \33589 , \33591 );
xor \U$33256 ( \33600 , \33599 , \33593 );
and \U$33257 ( \33601 , \23832 , \25180 );
and \U$33258 ( \33602 , \23665 , \25178 );
nor \U$33259 ( \33603 , \33601 , \33602 );
xnor \U$33260 ( \33604 , \33603 , \25037 );
and \U$33261 ( \33605 , \24089 , \24857 );
and \U$33262 ( \33606 , \23970 , \24855 );
nor \U$33263 ( \33607 , \33605 , \33606 );
xnor \U$33264 ( \33608 , \33607 , \24611 );
and \U$33265 ( \33609 , \33604 , \33608 );
and \U$33266 ( \33610 , \24714 , \24462 );
and \U$33267 ( \33611 , \24506 , \24460 );
nor \U$33268 ( \33612 , \33610 , \33611 );
xnor \U$33269 ( \33613 , \33612 , \24275 );
and \U$33270 ( \33614 , \33608 , \33613 );
and \U$33271 ( \33615 , \33604 , \33613 );
or \U$33272 ( \33616 , \33609 , \33614 , \33615 );
and \U$33273 ( \33617 , \24841 , \24149 );
and \U$33274 ( \33618 , \24836 , \24147 );
nor \U$33275 ( \33619 , \33617 , \33618 );
xnor \U$33276 ( \33620 , \33619 , \23944 );
and \U$33277 ( \33621 , \25294 , \23743 );
and \U$33278 ( \33622 , \25097 , \23741 );
nor \U$33279 ( \33623 , \33621 , \33622 );
xnor \U$33280 ( \33624 , \33623 , \23594 );
and \U$33281 ( \33625 , \33620 , \33624 );
and \U$33282 ( \33626 , \25604 , \23421 );
and \U$33283 ( \33627 , \25596 , \23419 );
nor \U$33284 ( \33628 , \33626 , \33627 );
xnor \U$33285 ( \33629 , \33628 , \23279 );
and \U$33286 ( \33630 , \33624 , \33629 );
and \U$33287 ( \33631 , \33620 , \33629 );
or \U$33288 ( \33632 , \33625 , \33630 , \33631 );
and \U$33289 ( \33633 , \33616 , \33632 );
and \U$33290 ( \33634 , \22872 , \26471 );
and \U$33291 ( \33635 , \22867 , \26469 );
nor \U$33292 ( \33636 , \33634 , \33635 );
xnor \U$33293 ( \33637 , \33636 , \26230 );
and \U$33294 ( \33638 , \23202 , \26005 );
and \U$33295 ( \33639 , \23058 , \26003 );
nor \U$33296 ( \33640 , \33638 , \33639 );
xnor \U$33297 ( \33641 , \33640 , \25817 );
and \U$33298 ( \33642 , \33637 , \33641 );
and \U$33299 ( \33643 , \23491 , \25631 );
and \U$33300 ( \33644 , \23466 , \25629 );
nor \U$33301 ( \33645 , \33643 , \33644 );
xnor \U$33302 ( \33646 , \33645 , \25399 );
and \U$33303 ( \33647 , \33641 , \33646 );
and \U$33304 ( \33648 , \33637 , \33646 );
or \U$33305 ( \33649 , \33642 , \33647 , \33648 );
and \U$33306 ( \33650 , \33632 , \33649 );
and \U$33307 ( \33651 , \33616 , \33649 );
or \U$33308 ( \33652 , \33633 , \33650 , \33651 );
and \U$33309 ( \33653 , \27527 , \22379 );
and \U$33310 ( \33654 , \27325 , \22377 );
nor \U$33311 ( \33655 , \33653 , \33654 );
xnor \U$33312 ( \33656 , \33655 , \22266 );
and \U$33313 ( \33657 , \28002 , \22185 );
and \U$33314 ( \33658 , \27830 , \22183 );
nor \U$33315 ( \33659 , \33657 , \33658 );
xnor \U$33316 ( \33660 , \33659 , \22049 );
and \U$33317 ( \33661 , \33656 , \33660 );
and \U$33318 ( \33662 , \28952 , \21985 );
and \U$33319 ( \33663 , \28528 , \21983 );
nor \U$33320 ( \33664 , \33662 , \33663 );
xnor \U$33321 ( \33665 , \33664 , \21907 );
and \U$33322 ( \33666 , \33660 , \33665 );
and \U$33323 ( \33667 , \33656 , \33665 );
or \U$33324 ( \33668 , \33661 , \33666 , \33667 );
and \U$33325 ( \33669 , \29203 , \21821 );
and \U$33326 ( \33670 , \29198 , \21819 );
nor \U$33327 ( \33671 , \33669 , \33670 );
xnor \U$33328 ( \33672 , \33671 , \21727 );
and \U$33329 ( \33673 , \29806 , \21652 );
and \U$33330 ( \33674 , \29522 , \21650 );
nor \U$33331 ( \33675 , \33673 , \33674 );
xnor \U$33332 ( \33676 , \33675 , \21377 );
and \U$33333 ( \33677 , \33672 , \33676 );
and \U$33334 ( \33678 , \30383 , \21385 );
and \U$33335 ( \33679 , \30375 , \21383 );
nor \U$33336 ( \33680 , \33678 , \33679 );
xnor \U$33337 ( \33681 , \33680 , \21392 );
and \U$33338 ( \33682 , \33676 , \33681 );
and \U$33339 ( \33683 , \33672 , \33681 );
or \U$33340 ( \33684 , \33677 , \33682 , \33683 );
and \U$33341 ( \33685 , \33668 , \33684 );
and \U$33342 ( \33686 , \26078 , \23125 );
and \U$33343 ( \33687 , \26073 , \23123 );
nor \U$33344 ( \33688 , \33686 , \33687 );
xnor \U$33345 ( \33689 , \33688 , \22988 );
and \U$33346 ( \33690 , \26601 , \22919 );
and \U$33347 ( \33691 , \26342 , \22917 );
nor \U$33348 ( \33692 , \33690 , \33691 );
xnor \U$33349 ( \33693 , \33692 , \22767 );
and \U$33350 ( \33694 , \33689 , \33693 );
and \U$33351 ( \33695 , \26982 , \22651 );
and \U$33352 ( \33696 , \26973 , \22649 );
nor \U$33353 ( \33697 , \33695 , \33696 );
xnor \U$33354 ( \33698 , \33697 , \22495 );
and \U$33355 ( \33699 , \33693 , \33698 );
and \U$33356 ( \33700 , \33689 , \33698 );
or \U$33357 ( \33701 , \33694 , \33699 , \33700 );
and \U$33358 ( \33702 , \33684 , \33701 );
and \U$33359 ( \33703 , \33668 , \33701 );
or \U$33360 ( \33704 , \33685 , \33702 , \33703 );
and \U$33361 ( \33705 , \33652 , \33704 );
and \U$33362 ( \33706 , \21428 , \31639 );
and \U$33363 ( \33707 , \21436 , \31636 );
nor \U$33364 ( \33708 , \33706 , \33707 );
xnor \U$33365 ( \33709 , \33708 , \30584 );
and \U$33366 ( \33710 , \21444 , \30826 );
and \U$33367 ( \33711 , \21452 , \30824 );
nor \U$33368 ( \33712 , \33710 , \33711 );
xnor \U$33369 ( \33713 , \33712 , \30587 );
and \U$33370 ( \33714 , \33709 , \33713 );
and \U$33371 ( \33715 , \21463 , \30258 );
and \U$33372 ( \33716 , \21471 , \30256 );
nor \U$33373 ( \33717 , \33715 , \33716 );
xnor \U$33374 ( \33718 , \33717 , \29948 );
and \U$33375 ( \33719 , \33713 , \33718 );
and \U$33376 ( \33720 , \33709 , \33718 );
or \U$33377 ( \33721 , \33714 , \33719 , \33720 );
and \U$33378 ( \33722 , \21689 , \29721 );
and \U$33379 ( \33723 , \21478 , \29719 );
nor \U$33380 ( \33724 , \33722 , \33723 );
xnor \U$33381 ( \33725 , \33724 , \29350 );
and \U$33382 ( \33726 , \21813 , \29159 );
and \U$33383 ( \33727 , \21750 , \29157 );
nor \U$33384 ( \33728 , \33726 , \33727 );
xnor \U$33385 ( \33729 , \33728 , \28841 );
and \U$33386 ( \33730 , \33725 , \33729 );
and \U$33387 ( \33731 , \22099 , \28592 );
and \U$33388 ( \33732 , \22011 , \28590 );
nor \U$33389 ( \33733 , \33731 , \33732 );
xnor \U$33390 ( \33734 , \33733 , \28343 );
and \U$33391 ( \33735 , \33729 , \33734 );
and \U$33392 ( \33736 , \33725 , \33734 );
or \U$33393 ( \33737 , \33730 , \33735 , \33736 );
and \U$33394 ( \33738 , \33721 , \33737 );
and \U$33395 ( \33739 , \22209 , \28063 );
and \U$33396 ( \33740 , \22204 , \28061 );
nor \U$33397 ( \33741 , \33739 , \33740 );
xnor \U$33398 ( \33742 , \33741 , \27803 );
and \U$33399 ( \33743 , \22440 , \27569 );
and \U$33400 ( \33744 , \22325 , \27567 );
nor \U$33401 ( \33745 , \33743 , \33744 );
xnor \U$33402 ( \33746 , \33745 , \27254 );
and \U$33403 ( \33747 , \33742 , \33746 );
and \U$33404 ( \33748 , \22624 , \27060 );
and \U$33405 ( \33749 , \22616 , \27058 );
nor \U$33406 ( \33750 , \33748 , \33749 );
xnor \U$33407 ( \33751 , \33750 , \26720 );
and \U$33408 ( \33752 , \33746 , \33751 );
and \U$33409 ( \33753 , \33742 , \33751 );
or \U$33410 ( \33754 , \33747 , \33752 , \33753 );
and \U$33411 ( \33755 , \33737 , \33754 );
and \U$33412 ( \33756 , \33721 , \33754 );
or \U$33413 ( \33757 , \33738 , \33755 , \33756 );
and \U$33414 ( \33758 , \33704 , \33757 );
and \U$33415 ( \33759 , \33652 , \33757 );
or \U$33416 ( \33760 , \33705 , \33758 , \33759 );
xor \U$33417 ( \33761 , \33367 , \33371 );
xor \U$33418 ( \33762 , \33761 , \33376 );
xor \U$33419 ( \33763 , \33431 , \33435 );
xor \U$33420 ( \33764 , \33763 , \33440 );
and \U$33421 ( \33765 , \33762 , \33764 );
xor \U$33422 ( \33766 , \33448 , \33452 );
xor \U$33423 ( \33767 , \33766 , \33457 );
and \U$33424 ( \33768 , \33764 , \33767 );
and \U$33425 ( \33769 , \33762 , \33767 );
or \U$33426 ( \33770 , \33765 , \33768 , \33769 );
xor \U$33427 ( \33771 , \33415 , \33419 );
xor \U$33428 ( \33772 , \33771 , \33424 );
xor \U$33429 ( \33773 , \33468 , \33472 );
xor \U$33430 ( \33774 , \33773 , \33477 );
and \U$33431 ( \33775 , \33772 , \33774 );
xor \U$33432 ( \33776 , \33484 , \33488 );
xor \U$33433 ( \33777 , \33776 , \33493 );
and \U$33434 ( \33778 , \33774 , \33777 );
and \U$33435 ( \33779 , \33772 , \33777 );
or \U$33436 ( \33780 , \33775 , \33778 , \33779 );
and \U$33437 ( \33781 , \33770 , \33780 );
nand \U$33438 ( \33782 , \31792 , \21432 );
xnor \U$33439 ( \33783 , \33782 , \21441 );
xor \U$33440 ( \33784 , \33501 , \33505 );
xor \U$33441 ( \33785 , \33784 , \33510 );
and \U$33442 ( \33786 , \33783 , \33785 );
xor \U$33443 ( \33787 , \33329 , \33333 );
xor \U$33444 ( \33788 , \33787 , \33338 );
and \U$33445 ( \33789 , \33785 , \33788 );
and \U$33446 ( \33790 , \33783 , \33788 );
or \U$33447 ( \33791 , \33786 , \33789 , \33790 );
and \U$33448 ( \33792 , \33780 , \33791 );
and \U$33449 ( \33793 , \33770 , \33791 );
or \U$33450 ( \33794 , \33781 , \33792 , \33793 );
and \U$33451 ( \33795 , \33760 , \33794 );
xor \U$33452 ( \33796 , \33118 , \33122 );
xor \U$33453 ( \33797 , \33796 , \33127 );
xor \U$33454 ( \33798 , \33135 , \33139 );
xor \U$33455 ( \33799 , \33798 , \33144 );
and \U$33456 ( \33800 , \33797 , \33799 );
xor \U$33457 ( \33801 , \33352 , \33354 );
xor \U$33458 ( \33802 , \33801 , \33357 );
and \U$33459 ( \33803 , \33799 , \33802 );
and \U$33460 ( \33804 , \33797 , \33802 );
or \U$33461 ( \33805 , \33800 , \33803 , \33804 );
and \U$33462 ( \33806 , \33794 , \33805 );
and \U$33463 ( \33807 , \33760 , \33805 );
or \U$33464 ( \33808 , \33795 , \33806 , \33807 );
xor \U$33465 ( \33809 , \33325 , \33349 );
xor \U$33466 ( \33810 , \33809 , \33360 );
xor \U$33467 ( \33811 , \33411 , \33463 );
xor \U$33468 ( \33812 , \33811 , \33516 );
and \U$33469 ( \33813 , \33810 , \33812 );
xor \U$33470 ( \33814 , \33522 , \33524 );
xor \U$33471 ( \33815 , \33814 , \33527 );
and \U$33472 ( \33816 , \33812 , \33815 );
and \U$33473 ( \33817 , \33810 , \33815 );
or \U$33474 ( \33818 , \33813 , \33816 , \33817 );
and \U$33475 ( \33819 , \33808 , \33818 );
xor \U$33476 ( \33820 , \33480 , \33496 );
xor \U$33477 ( \33821 , \33820 , \33513 );
xor \U$33478 ( \33822 , \33317 , \33319 );
xor \U$33479 ( \33823 , \33822 , \33322 );
and \U$33480 ( \33824 , \33821 , \33823 );
xor \U$33481 ( \33825 , \33341 , \33343 );
xor \U$33482 ( \33826 , \33825 , \33346 );
and \U$33483 ( \33827 , \33823 , \33826 );
and \U$33484 ( \33828 , \33821 , \33826 );
or \U$33485 ( \33829 , \33824 , \33827 , \33828 );
xor \U$33486 ( \33830 , \33114 , \33130 );
xor \U$33487 ( \33831 , \33830 , \33147 );
and \U$33488 ( \33832 , \33829 , \33831 );
xor \U$33489 ( \33833 , \33535 , \33537 );
xor \U$33490 ( \33834 , \33833 , \33540 );
and \U$33491 ( \33835 , \33831 , \33834 );
and \U$33492 ( \33836 , \33829 , \33834 );
or \U$33493 ( \33837 , \33832 , \33835 , \33836 );
and \U$33494 ( \33838 , \33818 , \33837 );
and \U$33495 ( \33839 , \33808 , \33837 );
or \U$33496 ( \33840 , \33819 , \33838 , \33839 );
xor \U$33497 ( \33841 , \33363 , \33519 );
xor \U$33498 ( \33842 , \33841 , \33530 );
xor \U$33499 ( \33843 , \33543 , \33545 );
xor \U$33500 ( \33844 , \33843 , \33548 );
and \U$33501 ( \33845 , \33842 , \33844 );
xor \U$33502 ( \33846 , \33554 , \33556 );
xor \U$33503 ( \33847 , \33846 , \33559 );
and \U$33504 ( \33848 , \33844 , \33847 );
and \U$33505 ( \33849 , \33842 , \33847 );
or \U$33506 ( \33850 , \33845 , \33848 , \33849 );
and \U$33507 ( \33851 , \33840 , \33850 );
xor \U$33508 ( \33852 , \33238 , \33248 );
xor \U$33509 ( \33853 , \33852 , \33251 );
and \U$33510 ( \33854 , \33850 , \33853 );
and \U$33511 ( \33855 , \33840 , \33853 );
or \U$33512 ( \33856 , \33851 , \33854 , \33855 );
xor \U$33513 ( \33857 , \33046 , \33206 );
xor \U$33514 ( \33858 , \33857 , \33225 );
xor \U$33515 ( \33859 , \33533 , \33551 );
xor \U$33516 ( \33860 , \33859 , \33562 );
and \U$33517 ( \33861 , \33858 , \33860 );
xor \U$33518 ( \33862 , \33567 , \33569 );
xor \U$33519 ( \33863 , \33862 , \33572 );
and \U$33520 ( \33864 , \33860 , \33863 );
and \U$33521 ( \33865 , \33858 , \33863 );
or \U$33522 ( \33866 , \33861 , \33864 , \33865 );
and \U$33523 ( \33867 , \33856 , \33866 );
xor \U$33524 ( \33868 , \33228 , \33254 );
xor \U$33525 ( \33869 , \33868 , \33265 );
and \U$33526 ( \33870 , \33866 , \33869 );
and \U$33527 ( \33871 , \33856 , \33869 );
or \U$33528 ( \33872 , \33867 , \33870 , \33871 );
xor \U$33529 ( \33873 , \33581 , \33583 );
xor \U$33530 ( \33874 , \33873 , \33586 );
and \U$33531 ( \33875 , \33872 , \33874 );
and \U$33532 ( \33876 , \33600 , \33875 );
xor \U$33533 ( \33877 , \33600 , \33875 );
xor \U$33534 ( \33878 , \33872 , \33874 );
and \U$33535 ( \33879 , \30986 , \21385 );
and \U$33536 ( \33880 , \30383 , \21383 );
nor \U$33537 ( \33881 , \33879 , \33880 );
xnor \U$33538 ( \33882 , \33881 , \21392 );
and \U$33539 ( \33883 , \31172 , \21401 );
and \U$33540 ( \33884 , \30991 , \21399 );
nor \U$33541 ( \33885 , \33883 , \33884 );
xnor \U$33542 ( \33886 , \33885 , \21408 );
and \U$33543 ( \33887 , \33882 , \33886 );
nand \U$33544 ( \33888 , \31792 , \21417 );
xnor \U$33545 ( \33889 , \33888 , \21426 );
and \U$33546 ( \33890 , \33886 , \33889 );
and \U$33547 ( \33891 , \33882 , \33889 );
or \U$33548 ( \33892 , \33887 , \33890 , \33891 );
and \U$33549 ( \33893 , \30991 , \21401 );
and \U$33550 ( \33894 , \30986 , \21399 );
nor \U$33551 ( \33895 , \33893 , \33894 );
xnor \U$33552 ( \33896 , \33895 , \21408 );
and \U$33553 ( \33897 , \33892 , \33896 );
and \U$33554 ( \33898 , \31792 , \21419 );
and \U$33555 ( \33899 , \31172 , \21417 );
nor \U$33556 ( \33900 , \33898 , \33899 );
xnor \U$33557 ( \33901 , \33900 , \21426 );
and \U$33558 ( \33902 , \33896 , \33901 );
and \U$33559 ( \33903 , \33892 , \33901 );
or \U$33560 ( \33904 , \33897 , \33902 , \33903 );
xor \U$33561 ( \33905 , \33656 , \33660 );
xor \U$33562 ( \33906 , \33905 , \33665 );
xor \U$33563 ( \33907 , \33672 , \33676 );
xor \U$33564 ( \33908 , \33907 , \33681 );
and \U$33565 ( \33909 , \33906 , \33908 );
xor \U$33566 ( \33910 , \33689 , \33693 );
xor \U$33567 ( \33911 , \33910 , \33698 );
and \U$33568 ( \33912 , \33908 , \33911 );
and \U$33569 ( \33913 , \33906 , \33911 );
or \U$33570 ( \33914 , \33909 , \33912 , \33913 );
and \U$33571 ( \33915 , \33904 , \33914 );
xor \U$33572 ( \33916 , \33604 , \33608 );
xor \U$33573 ( \33917 , \33916 , \33613 );
xor \U$33574 ( \33918 , \33620 , \33624 );
xor \U$33575 ( \33919 , \33918 , \33629 );
and \U$33576 ( \33920 , \33917 , \33919 );
xor \U$33577 ( \33921 , \33637 , \33641 );
xor \U$33578 ( \33922 , \33921 , \33646 );
and \U$33579 ( \33923 , \33919 , \33922 );
and \U$33580 ( \33924 , \33917 , \33922 );
or \U$33581 ( \33925 , \33920 , \33923 , \33924 );
and \U$33582 ( \33926 , \33914 , \33925 );
and \U$33583 ( \33927 , \33904 , \33925 );
or \U$33584 ( \33928 , \33915 , \33926 , \33927 );
and \U$33585 ( \33929 , \21478 , \30258 );
and \U$33586 ( \33930 , \21463 , \30256 );
nor \U$33587 ( \33931 , \33929 , \33930 );
xnor \U$33588 ( \33932 , \33931 , \29948 );
and \U$33589 ( \33933 , \21750 , \29721 );
and \U$33590 ( \33934 , \21689 , \29719 );
nor \U$33591 ( \33935 , \33933 , \33934 );
xnor \U$33592 ( \33936 , \33935 , \29350 );
and \U$33593 ( \33937 , \33932 , \33936 );
and \U$33594 ( \33938 , \22011 , \29159 );
and \U$33595 ( \33939 , \21813 , \29157 );
nor \U$33596 ( \33940 , \33938 , \33939 );
xnor \U$33597 ( \33941 , \33940 , \28841 );
and \U$33598 ( \33942 , \33936 , \33941 );
and \U$33599 ( \33943 , \33932 , \33941 );
or \U$33600 ( \33944 , \33937 , \33942 , \33943 );
and \U$33601 ( \33945 , \22204 , \28592 );
and \U$33602 ( \33946 , \22099 , \28590 );
nor \U$33603 ( \33947 , \33945 , \33946 );
xnor \U$33604 ( \33948 , \33947 , \28343 );
and \U$33605 ( \33949 , \22325 , \28063 );
and \U$33606 ( \33950 , \22209 , \28061 );
nor \U$33607 ( \33951 , \33949 , \33950 );
xnor \U$33608 ( \33952 , \33951 , \27803 );
and \U$33609 ( \33953 , \33948 , \33952 );
and \U$33610 ( \33954 , \22616 , \27569 );
and \U$33611 ( \33955 , \22440 , \27567 );
nor \U$33612 ( \33956 , \33954 , \33955 );
xnor \U$33613 ( \33957 , \33956 , \27254 );
and \U$33614 ( \33958 , \33952 , \33957 );
and \U$33615 ( \33959 , \33948 , \33957 );
or \U$33616 ( \33960 , \33953 , \33958 , \33959 );
and \U$33617 ( \33961 , \33944 , \33960 );
and \U$33618 ( \33962 , \21452 , \31639 );
and \U$33619 ( \33963 , \21428 , \31636 );
nor \U$33620 ( \33964 , \33962 , \33963 );
xnor \U$33621 ( \33965 , \33964 , \30584 );
and \U$33622 ( \33966 , \21471 , \30826 );
and \U$33623 ( \33967 , \21444 , \30824 );
nor \U$33624 ( \33968 , \33966 , \33967 );
xnor \U$33625 ( \33969 , \33968 , \30587 );
and \U$33626 ( \33970 , \33965 , \33969 );
and \U$33627 ( \33971 , \33969 , \21426 );
and \U$33628 ( \33972 , \33965 , \21426 );
or \U$33629 ( \33973 , \33970 , \33971 , \33972 );
and \U$33630 ( \33974 , \33960 , \33973 );
and \U$33631 ( \33975 , \33944 , \33973 );
or \U$33632 ( \33976 , \33961 , \33974 , \33975 );
and \U$33633 ( \33977 , \24836 , \24462 );
and \U$33634 ( \33978 , \24714 , \24460 );
nor \U$33635 ( \33979 , \33977 , \33978 );
xnor \U$33636 ( \33980 , \33979 , \24275 );
and \U$33637 ( \33981 , \25097 , \24149 );
and \U$33638 ( \33982 , \24841 , \24147 );
nor \U$33639 ( \33983 , \33981 , \33982 );
xnor \U$33640 ( \33984 , \33983 , \23944 );
and \U$33641 ( \33985 , \33980 , \33984 );
and \U$33642 ( \33986 , \25596 , \23743 );
and \U$33643 ( \33987 , \25294 , \23741 );
nor \U$33644 ( \33988 , \33986 , \33987 );
xnor \U$33645 ( \33989 , \33988 , \23594 );
and \U$33646 ( \33990 , \33984 , \33989 );
and \U$33647 ( \33991 , \33980 , \33989 );
or \U$33648 ( \33992 , \33985 , \33990 , \33991 );
and \U$33649 ( \33993 , \22867 , \27060 );
and \U$33650 ( \33994 , \22624 , \27058 );
nor \U$33651 ( \33995 , \33993 , \33994 );
xnor \U$33652 ( \33996 , \33995 , \26720 );
and \U$33653 ( \33997 , \23058 , \26471 );
and \U$33654 ( \33998 , \22872 , \26469 );
nor \U$33655 ( \33999 , \33997 , \33998 );
xnor \U$33656 ( \34000 , \33999 , \26230 );
and \U$33657 ( \34001 , \33996 , \34000 );
and \U$33658 ( \34002 , \23466 , \26005 );
and \U$33659 ( \34003 , \23202 , \26003 );
nor \U$33660 ( \34004 , \34002 , \34003 );
xnor \U$33661 ( \34005 , \34004 , \25817 );
and \U$33662 ( \34006 , \34000 , \34005 );
and \U$33663 ( \34007 , \33996 , \34005 );
or \U$33664 ( \34008 , \34001 , \34006 , \34007 );
and \U$33665 ( \34009 , \33992 , \34008 );
and \U$33666 ( \34010 , \23665 , \25631 );
and \U$33667 ( \34011 , \23491 , \25629 );
nor \U$33668 ( \34012 , \34010 , \34011 );
xnor \U$33669 ( \34013 , \34012 , \25399 );
and \U$33670 ( \34014 , \23970 , \25180 );
and \U$33671 ( \34015 , \23832 , \25178 );
nor \U$33672 ( \34016 , \34014 , \34015 );
xnor \U$33673 ( \34017 , \34016 , \25037 );
and \U$33674 ( \34018 , \34013 , \34017 );
and \U$33675 ( \34019 , \24506 , \24857 );
and \U$33676 ( \34020 , \24089 , \24855 );
nor \U$33677 ( \34021 , \34019 , \34020 );
xnor \U$33678 ( \34022 , \34021 , \24611 );
and \U$33679 ( \34023 , \34017 , \34022 );
and \U$33680 ( \34024 , \34013 , \34022 );
or \U$33681 ( \34025 , \34018 , \34023 , \34024 );
and \U$33682 ( \34026 , \34008 , \34025 );
and \U$33683 ( \34027 , \33992 , \34025 );
or \U$33684 ( \34028 , \34009 , \34026 , \34027 );
and \U$33685 ( \34029 , \33976 , \34028 );
and \U$33686 ( \34030 , \27325 , \22651 );
and \U$33687 ( \34031 , \26982 , \22649 );
nor \U$33688 ( \34032 , \34030 , \34031 );
xnor \U$33689 ( \34033 , \34032 , \22495 );
and \U$33690 ( \34034 , \27830 , \22379 );
and \U$33691 ( \34035 , \27527 , \22377 );
nor \U$33692 ( \34036 , \34034 , \34035 );
xnor \U$33693 ( \34037 , \34036 , \22266 );
and \U$33694 ( \34038 , \34033 , \34037 );
and \U$33695 ( \34039 , \28528 , \22185 );
and \U$33696 ( \34040 , \28002 , \22183 );
nor \U$33697 ( \34041 , \34039 , \34040 );
xnor \U$33698 ( \34042 , \34041 , \22049 );
and \U$33699 ( \34043 , \34037 , \34042 );
and \U$33700 ( \34044 , \34033 , \34042 );
or \U$33701 ( \34045 , \34038 , \34043 , \34044 );
and \U$33702 ( \34046 , \29198 , \21985 );
and \U$33703 ( \34047 , \28952 , \21983 );
nor \U$33704 ( \34048 , \34046 , \34047 );
xnor \U$33705 ( \34049 , \34048 , \21907 );
and \U$33706 ( \34050 , \29522 , \21821 );
and \U$33707 ( \34051 , \29203 , \21819 );
nor \U$33708 ( \34052 , \34050 , \34051 );
xnor \U$33709 ( \34053 , \34052 , \21727 );
and \U$33710 ( \34054 , \34049 , \34053 );
and \U$33711 ( \34055 , \30375 , \21652 );
and \U$33712 ( \34056 , \29806 , \21650 );
nor \U$33713 ( \34057 , \34055 , \34056 );
xnor \U$33714 ( \34058 , \34057 , \21377 );
and \U$33715 ( \34059 , \34053 , \34058 );
and \U$33716 ( \34060 , \34049 , \34058 );
or \U$33717 ( \34061 , \34054 , \34059 , \34060 );
and \U$33718 ( \34062 , \34045 , \34061 );
and \U$33719 ( \34063 , \26073 , \23421 );
and \U$33720 ( \34064 , \25604 , \23419 );
nor \U$33721 ( \34065 , \34063 , \34064 );
xnor \U$33722 ( \34066 , \34065 , \23279 );
and \U$33723 ( \34067 , \26342 , \23125 );
and \U$33724 ( \34068 , \26078 , \23123 );
nor \U$33725 ( \34069 , \34067 , \34068 );
xnor \U$33726 ( \34070 , \34069 , \22988 );
and \U$33727 ( \34071 , \34066 , \34070 );
and \U$33728 ( \34072 , \26973 , \22919 );
and \U$33729 ( \34073 , \26601 , \22917 );
nor \U$33730 ( \34074 , \34072 , \34073 );
xnor \U$33731 ( \34075 , \34074 , \22767 );
and \U$33732 ( \34076 , \34070 , \34075 );
and \U$33733 ( \34077 , \34066 , \34075 );
or \U$33734 ( \34078 , \34071 , \34076 , \34077 );
and \U$33735 ( \34079 , \34061 , \34078 );
and \U$33736 ( \34080 , \34045 , \34078 );
or \U$33737 ( \34081 , \34062 , \34079 , \34080 );
and \U$33738 ( \34082 , \34028 , \34081 );
and \U$33739 ( \34083 , \33976 , \34081 );
or \U$33740 ( \34084 , \34029 , \34082 , \34083 );
and \U$33741 ( \34085 , \33928 , \34084 );
xor \U$33742 ( \34086 , \33709 , \33713 );
xor \U$33743 ( \34087 , \34086 , \33718 );
xor \U$33744 ( \34088 , \33725 , \33729 );
xor \U$33745 ( \34089 , \34088 , \33734 );
and \U$33746 ( \34090 , \34087 , \34089 );
xor \U$33747 ( \34091 , \33742 , \33746 );
xor \U$33748 ( \34092 , \34091 , \33751 );
and \U$33749 ( \34093 , \34089 , \34092 );
and \U$33750 ( \34094 , \34087 , \34092 );
or \U$33751 ( \34095 , \34090 , \34093 , \34094 );
xor \U$33752 ( \34096 , \33383 , \33387 );
xor \U$33753 ( \34097 , \34096 , \21441 );
and \U$33754 ( \34098 , \34095 , \34097 );
xor \U$33755 ( \34099 , \33396 , \33400 );
xor \U$33756 ( \34100 , \34099 , \33405 );
and \U$33757 ( \34101 , \34097 , \34100 );
and \U$33758 ( \34102 , \34095 , \34100 );
or \U$33759 ( \34103 , \34098 , \34101 , \34102 );
and \U$33760 ( \34104 , \34084 , \34103 );
and \U$33761 ( \34105 , \33928 , \34103 );
or \U$33762 ( \34106 , \34085 , \34104 , \34105 );
xor \U$33763 ( \34107 , \33616 , \33632 );
xor \U$33764 ( \34108 , \34107 , \33649 );
xor \U$33765 ( \34109 , \33668 , \33684 );
xor \U$33766 ( \34110 , \34109 , \33701 );
and \U$33767 ( \34111 , \34108 , \34110 );
xor \U$33768 ( \34112 , \33721 , \33737 );
xor \U$33769 ( \34113 , \34112 , \33754 );
and \U$33770 ( \34114 , \34110 , \34113 );
and \U$33771 ( \34115 , \34108 , \34113 );
or \U$33772 ( \34116 , \34111 , \34114 , \34115 );
xor \U$33773 ( \34117 , \33762 , \33764 );
xor \U$33774 ( \34118 , \34117 , \33767 );
xor \U$33775 ( \34119 , \33772 , \33774 );
xor \U$33776 ( \34120 , \34119 , \33777 );
and \U$33777 ( \34121 , \34118 , \34120 );
xor \U$33778 ( \34122 , \33783 , \33785 );
xor \U$33779 ( \34123 , \34122 , \33788 );
and \U$33780 ( \34124 , \34120 , \34123 );
and \U$33781 ( \34125 , \34118 , \34123 );
or \U$33782 ( \34126 , \34121 , \34124 , \34125 );
and \U$33783 ( \34127 , \34116 , \34126 );
xor \U$33784 ( \34128 , \33427 , \33443 );
xor \U$33785 ( \34129 , \34128 , \33460 );
and \U$33786 ( \34130 , \34126 , \34129 );
and \U$33787 ( \34131 , \34116 , \34129 );
or \U$33788 ( \34132 , \34127 , \34130 , \34131 );
and \U$33789 ( \34133 , \34106 , \34132 );
xor \U$33790 ( \34134 , \33379 , \33391 );
xor \U$33791 ( \34135 , \34134 , \33408 );
xor \U$33792 ( \34136 , \33797 , \33799 );
xor \U$33793 ( \34137 , \34136 , \33802 );
and \U$33794 ( \34138 , \34135 , \34137 );
xor \U$33795 ( \34139 , \33821 , \33823 );
xor \U$33796 ( \34140 , \34139 , \33826 );
and \U$33797 ( \34141 , \34137 , \34140 );
and \U$33798 ( \34142 , \34135 , \34140 );
or \U$33799 ( \34143 , \34138 , \34141 , \34142 );
and \U$33800 ( \34144 , \34132 , \34143 );
and \U$33801 ( \34145 , \34106 , \34143 );
or \U$33802 ( \34146 , \34133 , \34144 , \34145 );
xor \U$33803 ( \34147 , \33760 , \33794 );
xor \U$33804 ( \34148 , \34147 , \33805 );
xor \U$33805 ( \34149 , \33810 , \33812 );
xor \U$33806 ( \34150 , \34149 , \33815 );
and \U$33807 ( \34151 , \34148 , \34150 );
xor \U$33808 ( \34152 , \33829 , \33831 );
xor \U$33809 ( \34153 , \34152 , \33834 );
and \U$33810 ( \34154 , \34150 , \34153 );
and \U$33811 ( \34155 , \34148 , \34153 );
or \U$33812 ( \34156 , \34151 , \34154 , \34155 );
and \U$33813 ( \34157 , \34146 , \34156 );
xor \U$33814 ( \34158 , \33842 , \33844 );
xor \U$33815 ( \34159 , \34158 , \33847 );
and \U$33816 ( \34160 , \34156 , \34159 );
and \U$33817 ( \34161 , \34146 , \34159 );
or \U$33818 ( \34162 , \34157 , \34160 , \34161 );
xor \U$33819 ( \34163 , \33840 , \33850 );
xor \U$33820 ( \34164 , \34163 , \33853 );
and \U$33821 ( \34165 , \34162 , \34164 );
xor \U$33822 ( \34166 , \33858 , \33860 );
xor \U$33823 ( \34167 , \34166 , \33863 );
and \U$33824 ( \34168 , \34164 , \34167 );
and \U$33825 ( \34169 , \34162 , \34167 );
or \U$33826 ( \34170 , \34165 , \34168 , \34169 );
xor \U$33827 ( \34171 , \33856 , \33866 );
xor \U$33828 ( \34172 , \34171 , \33869 );
and \U$33829 ( \34173 , \34170 , \34172 );
xor \U$33830 ( \34174 , \33565 , \33575 );
xor \U$33831 ( \34175 , \34174 , \33578 );
and \U$33832 ( \34176 , \34172 , \34175 );
and \U$33833 ( \34177 , \34170 , \34175 );
or \U$33834 ( \34178 , \34173 , \34176 , \34177 );
and \U$33835 ( \34179 , \33878 , \34178 );
xor \U$33836 ( \34180 , \33878 , \34178 );
xor \U$33837 ( \34181 , \34170 , \34172 );
xor \U$33838 ( \34182 , \34181 , \34175 );
xor \U$33839 ( \34183 , \33932 , \33936 );
xor \U$33840 ( \34184 , \34183 , \33941 );
xor \U$33841 ( \34185 , \33948 , \33952 );
xor \U$33842 ( \34186 , \34185 , \33957 );
and \U$33843 ( \34187 , \34184 , \34186 );
xor \U$33844 ( \34188 , \33996 , \34000 );
xor \U$33845 ( \34189 , \34188 , \34005 );
and \U$33846 ( \34190 , \34186 , \34189 );
and \U$33847 ( \34191 , \34184 , \34189 );
or \U$33848 ( \34192 , \34187 , \34190 , \34191 );
xor \U$33849 ( \34193 , \33980 , \33984 );
xor \U$33850 ( \34194 , \34193 , \33989 );
xor \U$33851 ( \34195 , \34013 , \34017 );
xor \U$33852 ( \34196 , \34195 , \34022 );
and \U$33853 ( \34197 , \34194 , \34196 );
xor \U$33854 ( \34198 , \34066 , \34070 );
xor \U$33855 ( \34199 , \34198 , \34075 );
and \U$33856 ( \34200 , \34196 , \34199 );
and \U$33857 ( \34201 , \34194 , \34199 );
or \U$33858 ( \34202 , \34197 , \34200 , \34201 );
and \U$33859 ( \34203 , \34192 , \34202 );
xor \U$33860 ( \34204 , \34033 , \34037 );
xor \U$33861 ( \34205 , \34204 , \34042 );
xor \U$33862 ( \34206 , \33882 , \33886 );
xor \U$33863 ( \34207 , \34206 , \33889 );
and \U$33864 ( \34208 , \34205 , \34207 );
xor \U$33865 ( \34209 , \34049 , \34053 );
xor \U$33866 ( \34210 , \34209 , \34058 );
and \U$33867 ( \34211 , \34207 , \34210 );
and \U$33868 ( \34212 , \34205 , \34210 );
or \U$33869 ( \34213 , \34208 , \34211 , \34212 );
and \U$33870 ( \34214 , \34202 , \34213 );
and \U$33871 ( \34215 , \34192 , \34213 );
or \U$33872 ( \34216 , \34203 , \34214 , \34215 );
and \U$33873 ( \34217 , \23202 , \26471 );
and \U$33874 ( \34218 , \23058 , \26469 );
nor \U$33875 ( \34219 , \34217 , \34218 );
xnor \U$33876 ( \34220 , \34219 , \26230 );
and \U$33877 ( \34221 , \23491 , \26005 );
and \U$33878 ( \34222 , \23466 , \26003 );
nor \U$33879 ( \34223 , \34221 , \34222 );
xnor \U$33880 ( \34224 , \34223 , \25817 );
and \U$33881 ( \34225 , \34220 , \34224 );
and \U$33882 ( \34226 , \23832 , \25631 );
and \U$33883 ( \34227 , \23665 , \25629 );
nor \U$33884 ( \34228 , \34226 , \34227 );
xnor \U$33885 ( \34229 , \34228 , \25399 );
and \U$33886 ( \34230 , \34224 , \34229 );
and \U$33887 ( \34231 , \34220 , \34229 );
or \U$33888 ( \34232 , \34225 , \34230 , \34231 );
and \U$33889 ( \34233 , \25294 , \24149 );
and \U$33890 ( \34234 , \25097 , \24147 );
nor \U$33891 ( \34235 , \34233 , \34234 );
xnor \U$33892 ( \34236 , \34235 , \23944 );
and \U$33893 ( \34237 , \25604 , \23743 );
and \U$33894 ( \34238 , \25596 , \23741 );
nor \U$33895 ( \34239 , \34237 , \34238 );
xnor \U$33896 ( \34240 , \34239 , \23594 );
and \U$33897 ( \34241 , \34236 , \34240 );
and \U$33898 ( \34242 , \26078 , \23421 );
and \U$33899 ( \34243 , \26073 , \23419 );
nor \U$33900 ( \34244 , \34242 , \34243 );
xnor \U$33901 ( \34245 , \34244 , \23279 );
and \U$33902 ( \34246 , \34240 , \34245 );
and \U$33903 ( \34247 , \34236 , \34245 );
or \U$33904 ( \34248 , \34241 , \34246 , \34247 );
and \U$33905 ( \34249 , \34232 , \34248 );
and \U$33906 ( \34250 , \24089 , \25180 );
and \U$33907 ( \34251 , \23970 , \25178 );
nor \U$33908 ( \34252 , \34250 , \34251 );
xnor \U$33909 ( \34253 , \34252 , \25037 );
and \U$33910 ( \34254 , \24714 , \24857 );
and \U$33911 ( \34255 , \24506 , \24855 );
nor \U$33912 ( \34256 , \34254 , \34255 );
xnor \U$33913 ( \34257 , \34256 , \24611 );
and \U$33914 ( \34258 , \34253 , \34257 );
and \U$33915 ( \34259 , \24841 , \24462 );
and \U$33916 ( \34260 , \24836 , \24460 );
nor \U$33917 ( \34261 , \34259 , \34260 );
xnor \U$33918 ( \34262 , \34261 , \24275 );
and \U$33919 ( \34263 , \34257 , \34262 );
and \U$33920 ( \34264 , \34253 , \34262 );
or \U$33921 ( \34265 , \34258 , \34263 , \34264 );
and \U$33922 ( \34266 , \34248 , \34265 );
and \U$33923 ( \34267 , \34232 , \34265 );
or \U$33924 ( \34268 , \34249 , \34266 , \34267 );
and \U$33925 ( \34269 , \29806 , \21821 );
and \U$33926 ( \34270 , \29522 , \21819 );
nor \U$33927 ( \34271 , \34269 , \34270 );
xnor \U$33928 ( \34272 , \34271 , \21727 );
and \U$33929 ( \34273 , \30383 , \21652 );
and \U$33930 ( \34274 , \30375 , \21650 );
nor \U$33931 ( \34275 , \34273 , \34274 );
xnor \U$33932 ( \34276 , \34275 , \21377 );
and \U$33933 ( \34277 , \34272 , \34276 );
and \U$33934 ( \34278 , \30991 , \21385 );
and \U$33935 ( \34279 , \30986 , \21383 );
nor \U$33936 ( \34280 , \34278 , \34279 );
xnor \U$33937 ( \34281 , \34280 , \21392 );
and \U$33938 ( \34282 , \34276 , \34281 );
and \U$33939 ( \34283 , \34272 , \34281 );
or \U$33940 ( \34284 , \34277 , \34282 , \34283 );
and \U$33941 ( \34285 , \28002 , \22379 );
and \U$33942 ( \34286 , \27830 , \22377 );
nor \U$33943 ( \34287 , \34285 , \34286 );
xnor \U$33944 ( \34288 , \34287 , \22266 );
and \U$33945 ( \34289 , \28952 , \22185 );
and \U$33946 ( \34290 , \28528 , \22183 );
nor \U$33947 ( \34291 , \34289 , \34290 );
xnor \U$33948 ( \34292 , \34291 , \22049 );
and \U$33949 ( \34293 , \34288 , \34292 );
and \U$33950 ( \34294 , \29203 , \21985 );
and \U$33951 ( \34295 , \29198 , \21983 );
nor \U$33952 ( \34296 , \34294 , \34295 );
xnor \U$33953 ( \34297 , \34296 , \21907 );
and \U$33954 ( \34298 , \34292 , \34297 );
and \U$33955 ( \34299 , \34288 , \34297 );
or \U$33956 ( \34300 , \34293 , \34298 , \34299 );
and \U$33957 ( \34301 , \34284 , \34300 );
and \U$33958 ( \34302 , \26601 , \23125 );
and \U$33959 ( \34303 , \26342 , \23123 );
nor \U$33960 ( \34304 , \34302 , \34303 );
xnor \U$33961 ( \34305 , \34304 , \22988 );
and \U$33962 ( \34306 , \26982 , \22919 );
and \U$33963 ( \34307 , \26973 , \22917 );
nor \U$33964 ( \34308 , \34306 , \34307 );
xnor \U$33965 ( \34309 , \34308 , \22767 );
and \U$33966 ( \34310 , \34305 , \34309 );
and \U$33967 ( \34311 , \27527 , \22651 );
and \U$33968 ( \34312 , \27325 , \22649 );
nor \U$33969 ( \34313 , \34311 , \34312 );
xnor \U$33970 ( \34314 , \34313 , \22495 );
and \U$33971 ( \34315 , \34309 , \34314 );
and \U$33972 ( \34316 , \34305 , \34314 );
or \U$33973 ( \34317 , \34310 , \34315 , \34316 );
and \U$33974 ( \34318 , \34300 , \34317 );
and \U$33975 ( \34319 , \34284 , \34317 );
or \U$33976 ( \34320 , \34301 , \34318 , \34319 );
and \U$33977 ( \34321 , \34268 , \34320 );
and \U$33978 ( \34322 , \22440 , \28063 );
and \U$33979 ( \34323 , \22325 , \28061 );
nor \U$33980 ( \34324 , \34322 , \34323 );
xnor \U$33981 ( \34325 , \34324 , \27803 );
and \U$33982 ( \34326 , \22624 , \27569 );
and \U$33983 ( \34327 , \22616 , \27567 );
nor \U$33984 ( \34328 , \34326 , \34327 );
xnor \U$33985 ( \34329 , \34328 , \27254 );
and \U$33986 ( \34330 , \34325 , \34329 );
and \U$33987 ( \34331 , \22872 , \27060 );
and \U$33988 ( \34332 , \22867 , \27058 );
nor \U$33989 ( \34333 , \34331 , \34332 );
xnor \U$33990 ( \34334 , \34333 , \26720 );
and \U$33991 ( \34335 , \34329 , \34334 );
and \U$33992 ( \34336 , \34325 , \34334 );
or \U$33993 ( \34337 , \34330 , \34335 , \34336 );
and \U$33994 ( \34338 , \21444 , \31639 );
and \U$33995 ( \34339 , \21452 , \31636 );
nor \U$33996 ( \34340 , \34338 , \34339 );
xnor \U$33997 ( \34341 , \34340 , \30584 );
and \U$33998 ( \34342 , \21463 , \30826 );
and \U$33999 ( \34343 , \21471 , \30824 );
nor \U$34000 ( \34344 , \34342 , \34343 );
xnor \U$34001 ( \34345 , \34344 , \30587 );
and \U$34002 ( \34346 , \34341 , \34345 );
and \U$34003 ( \34347 , \21689 , \30258 );
and \U$34004 ( \34348 , \21478 , \30256 );
nor \U$34005 ( \34349 , \34347 , \34348 );
xnor \U$34006 ( \34350 , \34349 , \29948 );
and \U$34007 ( \34351 , \34345 , \34350 );
and \U$34008 ( \34352 , \34341 , \34350 );
or \U$34009 ( \34353 , \34346 , \34351 , \34352 );
and \U$34010 ( \34354 , \34337 , \34353 );
and \U$34011 ( \34355 , \21813 , \29721 );
and \U$34012 ( \34356 , \21750 , \29719 );
nor \U$34013 ( \34357 , \34355 , \34356 );
xnor \U$34014 ( \34358 , \34357 , \29350 );
and \U$34015 ( \34359 , \22099 , \29159 );
and \U$34016 ( \34360 , \22011 , \29157 );
nor \U$34017 ( \34361 , \34359 , \34360 );
xnor \U$34018 ( \34362 , \34361 , \28841 );
and \U$34019 ( \34363 , \34358 , \34362 );
and \U$34020 ( \34364 , \22209 , \28592 );
and \U$34021 ( \34365 , \22204 , \28590 );
nor \U$34022 ( \34366 , \34364 , \34365 );
xnor \U$34023 ( \34367 , \34366 , \28343 );
and \U$34024 ( \34368 , \34362 , \34367 );
and \U$34025 ( \34369 , \34358 , \34367 );
or \U$34026 ( \34370 , \34363 , \34368 , \34369 );
and \U$34027 ( \34371 , \34353 , \34370 );
and \U$34028 ( \34372 , \34337 , \34370 );
or \U$34029 ( \34373 , \34354 , \34371 , \34372 );
and \U$34030 ( \34374 , \34320 , \34373 );
and \U$34031 ( \34375 , \34268 , \34373 );
or \U$34032 ( \34376 , \34321 , \34374 , \34375 );
and \U$34033 ( \34377 , \34216 , \34376 );
xor \U$34034 ( \34378 , \33906 , \33908 );
xor \U$34035 ( \34379 , \34378 , \33911 );
xor \U$34036 ( \34380 , \34087 , \34089 );
xor \U$34037 ( \34381 , \34380 , \34092 );
and \U$34038 ( \34382 , \34379 , \34381 );
xor \U$34039 ( \34383 , \33917 , \33919 );
xor \U$34040 ( \34384 , \34383 , \33922 );
and \U$34041 ( \34385 , \34381 , \34384 );
and \U$34042 ( \34386 , \34379 , \34384 );
or \U$34043 ( \34387 , \34382 , \34385 , \34386 );
and \U$34044 ( \34388 , \34376 , \34387 );
and \U$34045 ( \34389 , \34216 , \34387 );
or \U$34046 ( \34390 , \34377 , \34388 , \34389 );
xor \U$34047 ( \34391 , \33904 , \33914 );
xor \U$34048 ( \34392 , \34391 , \33925 );
xor \U$34049 ( \34393 , \33976 , \34028 );
xor \U$34050 ( \34394 , \34393 , \34081 );
and \U$34051 ( \34395 , \34392 , \34394 );
xor \U$34052 ( \34396 , \34095 , \34097 );
xor \U$34053 ( \34397 , \34396 , \34100 );
and \U$34054 ( \34398 , \34394 , \34397 );
and \U$34055 ( \34399 , \34392 , \34397 );
or \U$34056 ( \34400 , \34395 , \34398 , \34399 );
and \U$34057 ( \34401 , \34390 , \34400 );
xor \U$34058 ( \34402 , \33892 , \33896 );
xor \U$34059 ( \34403 , \34402 , \33901 );
xor \U$34060 ( \34404 , \33992 , \34008 );
xor \U$34061 ( \34405 , \34404 , \34025 );
and \U$34062 ( \34406 , \34403 , \34405 );
xor \U$34063 ( \34407 , \34045 , \34061 );
xor \U$34064 ( \34408 , \34407 , \34078 );
and \U$34065 ( \34409 , \34405 , \34408 );
and \U$34066 ( \34410 , \34403 , \34408 );
or \U$34067 ( \34411 , \34406 , \34409 , \34410 );
xor \U$34068 ( \34412 , \34108 , \34110 );
xor \U$34069 ( \34413 , \34412 , \34113 );
and \U$34070 ( \34414 , \34411 , \34413 );
xor \U$34071 ( \34415 , \34118 , \34120 );
xor \U$34072 ( \34416 , \34415 , \34123 );
and \U$34073 ( \34417 , \34413 , \34416 );
and \U$34074 ( \34418 , \34411 , \34416 );
or \U$34075 ( \34419 , \34414 , \34417 , \34418 );
and \U$34076 ( \34420 , \34400 , \34419 );
and \U$34077 ( \34421 , \34390 , \34419 );
or \U$34078 ( \34422 , \34401 , \34420 , \34421 );
xor \U$34079 ( \34423 , \33652 , \33704 );
xor \U$34080 ( \34424 , \34423 , \33757 );
xor \U$34081 ( \34425 , \33770 , \33780 );
xor \U$34082 ( \34426 , \34425 , \33791 );
and \U$34083 ( \34427 , \34424 , \34426 );
xor \U$34084 ( \34428 , \34135 , \34137 );
xor \U$34085 ( \34429 , \34428 , \34140 );
and \U$34086 ( \34430 , \34426 , \34429 );
and \U$34087 ( \34431 , \34424 , \34429 );
or \U$34088 ( \34432 , \34427 , \34430 , \34431 );
and \U$34089 ( \34433 , \34422 , \34432 );
xor \U$34090 ( \34434 , \34148 , \34150 );
xor \U$34091 ( \34435 , \34434 , \34153 );
and \U$34092 ( \34436 , \34432 , \34435 );
and \U$34093 ( \34437 , \34422 , \34435 );
or \U$34094 ( \34438 , \34433 , \34436 , \34437 );
xor \U$34095 ( \34439 , \33808 , \33818 );
xor \U$34096 ( \34440 , \34439 , \33837 );
and \U$34097 ( \34441 , \34438 , \34440 );
xor \U$34098 ( \34442 , \34146 , \34156 );
xor \U$34099 ( \34443 , \34442 , \34159 );
and \U$34100 ( \34444 , \34440 , \34443 );
and \U$34101 ( \34445 , \34438 , \34443 );
or \U$34102 ( \34446 , \34441 , \34444 , \34445 );
xor \U$34103 ( \34447 , \34162 , \34164 );
xor \U$34104 ( \34448 , \34447 , \34167 );
and \U$34105 ( \34449 , \34446 , \34448 );
and \U$34106 ( \34450 , \34182 , \34449 );
xor \U$34107 ( \34451 , \34182 , \34449 );
xor \U$34108 ( \34452 , \34446 , \34448 );
xor \U$34109 ( \34453 , \34236 , \34240 );
xor \U$34110 ( \34454 , \34453 , \34245 );
xor \U$34111 ( \34455 , \34253 , \34257 );
xor \U$34112 ( \34456 , \34455 , \34262 );
and \U$34113 ( \34457 , \34454 , \34456 );
xor \U$34114 ( \34458 , \34305 , \34309 );
xor \U$34115 ( \34459 , \34458 , \34314 );
and \U$34116 ( \34460 , \34456 , \34459 );
and \U$34117 ( \34461 , \34454 , \34459 );
or \U$34118 ( \34462 , \34457 , \34460 , \34461 );
xor \U$34119 ( \34463 , \34220 , \34224 );
xor \U$34120 ( \34464 , \34463 , \34229 );
xor \U$34121 ( \34465 , \34325 , \34329 );
xor \U$34122 ( \34466 , \34465 , \34334 );
and \U$34123 ( \34467 , \34464 , \34466 );
xor \U$34124 ( \34468 , \34358 , \34362 );
xor \U$34125 ( \34469 , \34468 , \34367 );
and \U$34126 ( \34470 , \34466 , \34469 );
and \U$34127 ( \34471 , \34464 , \34469 );
or \U$34128 ( \34472 , \34467 , \34470 , \34471 );
and \U$34129 ( \34473 , \34462 , \34472 );
and \U$34130 ( \34474 , \31792 , \21401 );
and \U$34131 ( \34475 , \31172 , \21399 );
nor \U$34132 ( \34476 , \34474 , \34475 );
xnor \U$34133 ( \34477 , \34476 , \21408 );
xor \U$34134 ( \34478 , \34272 , \34276 );
xor \U$34135 ( \34479 , \34478 , \34281 );
and \U$34136 ( \34480 , \34477 , \34479 );
xor \U$34137 ( \34481 , \34288 , \34292 );
xor \U$34138 ( \34482 , \34481 , \34297 );
and \U$34139 ( \34483 , \34479 , \34482 );
and \U$34140 ( \34484 , \34477 , \34482 );
or \U$34141 ( \34485 , \34480 , \34483 , \34484 );
and \U$34142 ( \34486 , \34472 , \34485 );
and \U$34143 ( \34487 , \34462 , \34485 );
or \U$34144 ( \34488 , \34473 , \34486 , \34487 );
and \U$34145 ( \34489 , \22325 , \28592 );
and \U$34146 ( \34490 , \22209 , \28590 );
nor \U$34147 ( \34491 , \34489 , \34490 );
xnor \U$34148 ( \34492 , \34491 , \28343 );
and \U$34149 ( \34493 , \22616 , \28063 );
and \U$34150 ( \34494 , \22440 , \28061 );
nor \U$34151 ( \34495 , \34493 , \34494 );
xnor \U$34152 ( \34496 , \34495 , \27803 );
and \U$34153 ( \34497 , \34492 , \34496 );
and \U$34154 ( \34498 , \22867 , \27569 );
and \U$34155 ( \34499 , \22624 , \27567 );
nor \U$34156 ( \34500 , \34498 , \34499 );
xnor \U$34157 ( \34501 , \34500 , \27254 );
and \U$34158 ( \34502 , \34496 , \34501 );
and \U$34159 ( \34503 , \34492 , \34501 );
or \U$34160 ( \34504 , \34497 , \34502 , \34503 );
and \U$34161 ( \34505 , \21750 , \30258 );
and \U$34162 ( \34506 , \21689 , \30256 );
nor \U$34163 ( \34507 , \34505 , \34506 );
xnor \U$34164 ( \34508 , \34507 , \29948 );
and \U$34165 ( \34509 , \22011 , \29721 );
and \U$34166 ( \34510 , \21813 , \29719 );
nor \U$34167 ( \34511 , \34509 , \34510 );
xnor \U$34168 ( \34512 , \34511 , \29350 );
and \U$34169 ( \34513 , \34508 , \34512 );
and \U$34170 ( \34514 , \22204 , \29159 );
and \U$34171 ( \34515 , \22099 , \29157 );
nor \U$34172 ( \34516 , \34514 , \34515 );
xnor \U$34173 ( \34517 , \34516 , \28841 );
and \U$34174 ( \34518 , \34512 , \34517 );
and \U$34175 ( \34519 , \34508 , \34517 );
or \U$34176 ( \34520 , \34513 , \34518 , \34519 );
and \U$34177 ( \34521 , \34504 , \34520 );
and \U$34178 ( \34522 , \21471 , \31639 );
and \U$34179 ( \34523 , \21444 , \31636 );
nor \U$34180 ( \34524 , \34522 , \34523 );
xnor \U$34181 ( \34525 , \34524 , \30584 );
and \U$34182 ( \34526 , \21478 , \30826 );
and \U$34183 ( \34527 , \21463 , \30824 );
nor \U$34184 ( \34528 , \34526 , \34527 );
xnor \U$34185 ( \34529 , \34528 , \30587 );
and \U$34186 ( \34530 , \34525 , \34529 );
and \U$34187 ( \34531 , \34529 , \21408 );
and \U$34188 ( \34532 , \34525 , \21408 );
or \U$34189 ( \34533 , \34530 , \34531 , \34532 );
and \U$34190 ( \34534 , \34520 , \34533 );
and \U$34191 ( \34535 , \34504 , \34533 );
or \U$34192 ( \34536 , \34521 , \34534 , \34535 );
and \U$34193 ( \34537 , \29522 , \21985 );
and \U$34194 ( \34538 , \29203 , \21983 );
nor \U$34195 ( \34539 , \34537 , \34538 );
xnor \U$34196 ( \34540 , \34539 , \21907 );
and \U$34197 ( \34541 , \30375 , \21821 );
and \U$34198 ( \34542 , \29806 , \21819 );
nor \U$34199 ( \34543 , \34541 , \34542 );
xnor \U$34200 ( \34544 , \34543 , \21727 );
and \U$34201 ( \34545 , \34540 , \34544 );
and \U$34202 ( \34546 , \30986 , \21652 );
and \U$34203 ( \34547 , \30383 , \21650 );
nor \U$34204 ( \34548 , \34546 , \34547 );
xnor \U$34205 ( \34549 , \34548 , \21377 );
and \U$34206 ( \34550 , \34544 , \34549 );
and \U$34207 ( \34551 , \34540 , \34549 );
or \U$34208 ( \34552 , \34545 , \34550 , \34551 );
and \U$34209 ( \34553 , \26342 , \23421 );
and \U$34210 ( \34554 , \26078 , \23419 );
nor \U$34211 ( \34555 , \34553 , \34554 );
xnor \U$34212 ( \34556 , \34555 , \23279 );
and \U$34213 ( \34557 , \26973 , \23125 );
and \U$34214 ( \34558 , \26601 , \23123 );
nor \U$34215 ( \34559 , \34557 , \34558 );
xnor \U$34216 ( \34560 , \34559 , \22988 );
and \U$34217 ( \34561 , \34556 , \34560 );
and \U$34218 ( \34562 , \27325 , \22919 );
and \U$34219 ( \34563 , \26982 , \22917 );
nor \U$34220 ( \34564 , \34562 , \34563 );
xnor \U$34221 ( \34565 , \34564 , \22767 );
and \U$34222 ( \34566 , \34560 , \34565 );
and \U$34223 ( \34567 , \34556 , \34565 );
or \U$34224 ( \34568 , \34561 , \34566 , \34567 );
and \U$34225 ( \34569 , \34552 , \34568 );
and \U$34226 ( \34570 , \27830 , \22651 );
and \U$34227 ( \34571 , \27527 , \22649 );
nor \U$34228 ( \34572 , \34570 , \34571 );
xnor \U$34229 ( \34573 , \34572 , \22495 );
and \U$34230 ( \34574 , \28528 , \22379 );
and \U$34231 ( \34575 , \28002 , \22377 );
nor \U$34232 ( \34576 , \34574 , \34575 );
xnor \U$34233 ( \34577 , \34576 , \22266 );
and \U$34234 ( \34578 , \34573 , \34577 );
and \U$34235 ( \34579 , \29198 , \22185 );
and \U$34236 ( \34580 , \28952 , \22183 );
nor \U$34237 ( \34581 , \34579 , \34580 );
xnor \U$34238 ( \34582 , \34581 , \22049 );
and \U$34239 ( \34583 , \34577 , \34582 );
and \U$34240 ( \34584 , \34573 , \34582 );
or \U$34241 ( \34585 , \34578 , \34583 , \34584 );
and \U$34242 ( \34586 , \34568 , \34585 );
and \U$34243 ( \34587 , \34552 , \34585 );
or \U$34244 ( \34588 , \34569 , \34586 , \34587 );
and \U$34245 ( \34589 , \34536 , \34588 );
and \U$34246 ( \34590 , \25097 , \24462 );
and \U$34247 ( \34591 , \24841 , \24460 );
nor \U$34248 ( \34592 , \34590 , \34591 );
xnor \U$34249 ( \34593 , \34592 , \24275 );
and \U$34250 ( \34594 , \25596 , \24149 );
and \U$34251 ( \34595 , \25294 , \24147 );
nor \U$34252 ( \34596 , \34594 , \34595 );
xnor \U$34253 ( \34597 , \34596 , \23944 );
and \U$34254 ( \34598 , \34593 , \34597 );
and \U$34255 ( \34599 , \26073 , \23743 );
and \U$34256 ( \34600 , \25604 , \23741 );
nor \U$34257 ( \34601 , \34599 , \34600 );
xnor \U$34258 ( \34602 , \34601 , \23594 );
and \U$34259 ( \34603 , \34597 , \34602 );
and \U$34260 ( \34604 , \34593 , \34602 );
or \U$34261 ( \34605 , \34598 , \34603 , \34604 );
and \U$34262 ( \34606 , \23970 , \25631 );
and \U$34263 ( \34607 , \23832 , \25629 );
nor \U$34264 ( \34608 , \34606 , \34607 );
xnor \U$34265 ( \34609 , \34608 , \25399 );
and \U$34266 ( \34610 , \24506 , \25180 );
and \U$34267 ( \34611 , \24089 , \25178 );
nor \U$34268 ( \34612 , \34610 , \34611 );
xnor \U$34269 ( \34613 , \34612 , \25037 );
and \U$34270 ( \34614 , \34609 , \34613 );
and \U$34271 ( \34615 , \24836 , \24857 );
and \U$34272 ( \34616 , \24714 , \24855 );
nor \U$34273 ( \34617 , \34615 , \34616 );
xnor \U$34274 ( \34618 , \34617 , \24611 );
and \U$34275 ( \34619 , \34613 , \34618 );
and \U$34276 ( \34620 , \34609 , \34618 );
or \U$34277 ( \34621 , \34614 , \34619 , \34620 );
and \U$34278 ( \34622 , \34605 , \34621 );
and \U$34279 ( \34623 , \23058 , \27060 );
and \U$34280 ( \34624 , \22872 , \27058 );
nor \U$34281 ( \34625 , \34623 , \34624 );
xnor \U$34282 ( \34626 , \34625 , \26720 );
and \U$34283 ( \34627 , \23466 , \26471 );
and \U$34284 ( \34628 , \23202 , \26469 );
nor \U$34285 ( \34629 , \34627 , \34628 );
xnor \U$34286 ( \34630 , \34629 , \26230 );
and \U$34287 ( \34631 , \34626 , \34630 );
and \U$34288 ( \34632 , \23665 , \26005 );
and \U$34289 ( \34633 , \23491 , \26003 );
nor \U$34290 ( \34634 , \34632 , \34633 );
xnor \U$34291 ( \34635 , \34634 , \25817 );
and \U$34292 ( \34636 , \34630 , \34635 );
and \U$34293 ( \34637 , \34626 , \34635 );
or \U$34294 ( \34638 , \34631 , \34636 , \34637 );
and \U$34295 ( \34639 , \34621 , \34638 );
and \U$34296 ( \34640 , \34605 , \34638 );
or \U$34297 ( \34641 , \34622 , \34639 , \34640 );
and \U$34298 ( \34642 , \34588 , \34641 );
and \U$34299 ( \34643 , \34536 , \34641 );
or \U$34300 ( \34644 , \34589 , \34642 , \34643 );
and \U$34301 ( \34645 , \34488 , \34644 );
xor \U$34302 ( \34646 , \33965 , \33969 );
xor \U$34303 ( \34647 , \34646 , \21426 );
xor \U$34304 ( \34648 , \34184 , \34186 );
xor \U$34305 ( \34649 , \34648 , \34189 );
and \U$34306 ( \34650 , \34647 , \34649 );
xor \U$34307 ( \34651 , \34194 , \34196 );
xor \U$34308 ( \34652 , \34651 , \34199 );
and \U$34309 ( \34653 , \34649 , \34652 );
and \U$34310 ( \34654 , \34647 , \34652 );
or \U$34311 ( \34655 , \34650 , \34653 , \34654 );
and \U$34312 ( \34656 , \34644 , \34655 );
and \U$34313 ( \34657 , \34488 , \34655 );
or \U$34314 ( \34658 , \34645 , \34656 , \34657 );
xor \U$34315 ( \34659 , \34232 , \34248 );
xor \U$34316 ( \34660 , \34659 , \34265 );
xor \U$34317 ( \34661 , \34284 , \34300 );
xor \U$34318 ( \34662 , \34661 , \34317 );
and \U$34319 ( \34663 , \34660 , \34662 );
xor \U$34320 ( \34664 , \34205 , \34207 );
xor \U$34321 ( \34665 , \34664 , \34210 );
and \U$34322 ( \34666 , \34662 , \34665 );
and \U$34323 ( \34667 , \34660 , \34665 );
or \U$34324 ( \34668 , \34663 , \34666 , \34667 );
xor \U$34325 ( \34669 , \33944 , \33960 );
xor \U$34326 ( \34670 , \34669 , \33973 );
and \U$34327 ( \34671 , \34668 , \34670 );
xor \U$34328 ( \34672 , \34403 , \34405 );
xor \U$34329 ( \34673 , \34672 , \34408 );
and \U$34330 ( \34674 , \34670 , \34673 );
and \U$34331 ( \34675 , \34668 , \34673 );
or \U$34332 ( \34676 , \34671 , \34674 , \34675 );
and \U$34333 ( \34677 , \34658 , \34676 );
xor \U$34334 ( \34678 , \34192 , \34202 );
xor \U$34335 ( \34679 , \34678 , \34213 );
xor \U$34336 ( \34680 , \34268 , \34320 );
xor \U$34337 ( \34681 , \34680 , \34373 );
and \U$34338 ( \34682 , \34679 , \34681 );
xor \U$34339 ( \34683 , \34379 , \34381 );
xor \U$34340 ( \34684 , \34683 , \34384 );
and \U$34341 ( \34685 , \34681 , \34684 );
and \U$34342 ( \34686 , \34679 , \34684 );
or \U$34343 ( \34687 , \34682 , \34685 , \34686 );
and \U$34344 ( \34688 , \34676 , \34687 );
and \U$34345 ( \34689 , \34658 , \34687 );
or \U$34346 ( \34690 , \34677 , \34688 , \34689 );
xor \U$34347 ( \34691 , \34216 , \34376 );
xor \U$34348 ( \34692 , \34691 , \34387 );
xor \U$34349 ( \34693 , \34392 , \34394 );
xor \U$34350 ( \34694 , \34693 , \34397 );
and \U$34351 ( \34695 , \34692 , \34694 );
xor \U$34352 ( \34696 , \34411 , \34413 );
xor \U$34353 ( \34697 , \34696 , \34416 );
and \U$34354 ( \34698 , \34694 , \34697 );
and \U$34355 ( \34699 , \34692 , \34697 );
or \U$34356 ( \34700 , \34695 , \34698 , \34699 );
and \U$34357 ( \34701 , \34690 , \34700 );
xor \U$34358 ( \34702 , \34116 , \34126 );
xor \U$34359 ( \34703 , \34702 , \34129 );
and \U$34360 ( \34704 , \34700 , \34703 );
and \U$34361 ( \34705 , \34690 , \34703 );
or \U$34362 ( \34706 , \34701 , \34704 , \34705 );
xor \U$34363 ( \34707 , \33928 , \34084 );
xor \U$34364 ( \34708 , \34707 , \34103 );
xor \U$34365 ( \34709 , \34390 , \34400 );
xor \U$34366 ( \34710 , \34709 , \34419 );
and \U$34367 ( \34711 , \34708 , \34710 );
xor \U$34368 ( \34712 , \34424 , \34426 );
xor \U$34369 ( \34713 , \34712 , \34429 );
and \U$34370 ( \34714 , \34710 , \34713 );
and \U$34371 ( \34715 , \34708 , \34713 );
or \U$34372 ( \34716 , \34711 , \34714 , \34715 );
and \U$34373 ( \34717 , \34706 , \34716 );
xor \U$34374 ( \34718 , \34106 , \34132 );
xor \U$34375 ( \34719 , \34718 , \34143 );
and \U$34376 ( \34720 , \34716 , \34719 );
and \U$34377 ( \34721 , \34706 , \34719 );
or \U$34378 ( \34722 , \34717 , \34720 , \34721 );
xor \U$34379 ( \34723 , \34438 , \34440 );
xor \U$34380 ( \34724 , \34723 , \34443 );
and \U$34381 ( \34725 , \34722 , \34724 );
and \U$34382 ( \34726 , \34452 , \34725 );
xor \U$34383 ( \34727 , \34452 , \34725 );
xor \U$34384 ( \34728 , \34722 , \34724 );
xor \U$34385 ( \34729 , \34593 , \34597 );
xor \U$34386 ( \34730 , \34729 , \34602 );
xor \U$34387 ( \34731 , \34556 , \34560 );
xor \U$34388 ( \34732 , \34731 , \34565 );
and \U$34389 ( \34733 , \34730 , \34732 );
xor \U$34390 ( \34734 , \34573 , \34577 );
xor \U$34391 ( \34735 , \34734 , \34582 );
and \U$34392 ( \34736 , \34732 , \34735 );
and \U$34393 ( \34737 , \34730 , \34735 );
or \U$34394 ( \34738 , \34733 , \34736 , \34737 );
and \U$34395 ( \34739 , \31172 , \21385 );
and \U$34396 ( \34740 , \30991 , \21383 );
nor \U$34397 ( \34741 , \34739 , \34740 );
xnor \U$34398 ( \34742 , \34741 , \21392 );
nand \U$34399 ( \34743 , \31792 , \21399 );
xnor \U$34400 ( \34744 , \34743 , \21408 );
and \U$34401 ( \34745 , \34742 , \34744 );
xor \U$34402 ( \34746 , \34540 , \34544 );
xor \U$34403 ( \34747 , \34746 , \34549 );
and \U$34404 ( \34748 , \34744 , \34747 );
and \U$34405 ( \34749 , \34742 , \34747 );
or \U$34406 ( \34750 , \34745 , \34748 , \34749 );
and \U$34407 ( \34751 , \34738 , \34750 );
xor \U$34408 ( \34752 , \34492 , \34496 );
xor \U$34409 ( \34753 , \34752 , \34501 );
xor \U$34410 ( \34754 , \34609 , \34613 );
xor \U$34411 ( \34755 , \34754 , \34618 );
and \U$34412 ( \34756 , \34753 , \34755 );
xor \U$34413 ( \34757 , \34626 , \34630 );
xor \U$34414 ( \34758 , \34757 , \34635 );
and \U$34415 ( \34759 , \34755 , \34758 );
and \U$34416 ( \34760 , \34753 , \34758 );
or \U$34417 ( \34761 , \34756 , \34759 , \34760 );
and \U$34418 ( \34762 , \34750 , \34761 );
and \U$34419 ( \34763 , \34738 , \34761 );
or \U$34420 ( \34764 , \34751 , \34762 , \34763 );
and \U$34421 ( \34765 , \30383 , \21821 );
and \U$34422 ( \34766 , \30375 , \21819 );
nor \U$34423 ( \34767 , \34765 , \34766 );
xnor \U$34424 ( \34768 , \34767 , \21727 );
and \U$34425 ( \34769 , \30991 , \21652 );
and \U$34426 ( \34770 , \30986 , \21650 );
nor \U$34427 ( \34771 , \34769 , \34770 );
xnor \U$34428 ( \34772 , \34771 , \21377 );
and \U$34429 ( \34773 , \34768 , \34772 );
and \U$34430 ( \34774 , \31792 , \21385 );
and \U$34431 ( \34775 , \31172 , \21383 );
nor \U$34432 ( \34776 , \34774 , \34775 );
xnor \U$34433 ( \34777 , \34776 , \21392 );
and \U$34434 ( \34778 , \34772 , \34777 );
and \U$34435 ( \34779 , \34768 , \34777 );
or \U$34436 ( \34780 , \34773 , \34778 , \34779 );
and \U$34437 ( \34781 , \26982 , \23125 );
and \U$34438 ( \34782 , \26973 , \23123 );
nor \U$34439 ( \34783 , \34781 , \34782 );
xnor \U$34440 ( \34784 , \34783 , \22988 );
and \U$34441 ( \34785 , \27527 , \22919 );
and \U$34442 ( \34786 , \27325 , \22917 );
nor \U$34443 ( \34787 , \34785 , \34786 );
xnor \U$34444 ( \34788 , \34787 , \22767 );
and \U$34445 ( \34789 , \34784 , \34788 );
and \U$34446 ( \34790 , \28002 , \22651 );
and \U$34447 ( \34791 , \27830 , \22649 );
nor \U$34448 ( \34792 , \34790 , \34791 );
xnor \U$34449 ( \34793 , \34792 , \22495 );
and \U$34450 ( \34794 , \34788 , \34793 );
and \U$34451 ( \34795 , \34784 , \34793 );
or \U$34452 ( \34796 , \34789 , \34794 , \34795 );
and \U$34453 ( \34797 , \34780 , \34796 );
and \U$34454 ( \34798 , \28952 , \22379 );
and \U$34455 ( \34799 , \28528 , \22377 );
nor \U$34456 ( \34800 , \34798 , \34799 );
xnor \U$34457 ( \34801 , \34800 , \22266 );
and \U$34458 ( \34802 , \29203 , \22185 );
and \U$34459 ( \34803 , \29198 , \22183 );
nor \U$34460 ( \34804 , \34802 , \34803 );
xnor \U$34461 ( \34805 , \34804 , \22049 );
and \U$34462 ( \34806 , \34801 , \34805 );
and \U$34463 ( \34807 , \29806 , \21985 );
and \U$34464 ( \34808 , \29522 , \21983 );
nor \U$34465 ( \34809 , \34807 , \34808 );
xnor \U$34466 ( \34810 , \34809 , \21907 );
and \U$34467 ( \34811 , \34805 , \34810 );
and \U$34468 ( \34812 , \34801 , \34810 );
or \U$34469 ( \34813 , \34806 , \34811 , \34812 );
and \U$34470 ( \34814 , \34796 , \34813 );
and \U$34471 ( \34815 , \34780 , \34813 );
or \U$34472 ( \34816 , \34797 , \34814 , \34815 );
and \U$34473 ( \34817 , \22099 , \29721 );
and \U$34474 ( \34818 , \22011 , \29719 );
nor \U$34475 ( \34819 , \34817 , \34818 );
xnor \U$34476 ( \34820 , \34819 , \29350 );
and \U$34477 ( \34821 , \22209 , \29159 );
and \U$34478 ( \34822 , \22204 , \29157 );
nor \U$34479 ( \34823 , \34821 , \34822 );
xnor \U$34480 ( \34824 , \34823 , \28841 );
and \U$34481 ( \34825 , \34820 , \34824 );
and \U$34482 ( \34826 , \22440 , \28592 );
and \U$34483 ( \34827 , \22325 , \28590 );
nor \U$34484 ( \34828 , \34826 , \34827 );
xnor \U$34485 ( \34829 , \34828 , \28343 );
and \U$34486 ( \34830 , \34824 , \34829 );
and \U$34487 ( \34831 , \34820 , \34829 );
or \U$34488 ( \34832 , \34825 , \34830 , \34831 );
and \U$34489 ( \34833 , \22624 , \28063 );
and \U$34490 ( \34834 , \22616 , \28061 );
nor \U$34491 ( \34835 , \34833 , \34834 );
xnor \U$34492 ( \34836 , \34835 , \27803 );
and \U$34493 ( \34837 , \22872 , \27569 );
and \U$34494 ( \34838 , \22867 , \27567 );
nor \U$34495 ( \34839 , \34837 , \34838 );
xnor \U$34496 ( \34840 , \34839 , \27254 );
and \U$34497 ( \34841 , \34836 , \34840 );
and \U$34498 ( \34842 , \23202 , \27060 );
and \U$34499 ( \34843 , \23058 , \27058 );
nor \U$34500 ( \34844 , \34842 , \34843 );
xnor \U$34501 ( \34845 , \34844 , \26720 );
and \U$34502 ( \34846 , \34840 , \34845 );
and \U$34503 ( \34847 , \34836 , \34845 );
or \U$34504 ( \34848 , \34841 , \34846 , \34847 );
and \U$34505 ( \34849 , \34832 , \34848 );
and \U$34506 ( \34850 , \21463 , \31639 );
and \U$34507 ( \34851 , \21471 , \31636 );
nor \U$34508 ( \34852 , \34850 , \34851 );
xnor \U$34509 ( \34853 , \34852 , \30584 );
and \U$34510 ( \34854 , \21689 , \30826 );
and \U$34511 ( \34855 , \21478 , \30824 );
nor \U$34512 ( \34856 , \34854 , \34855 );
xnor \U$34513 ( \34857 , \34856 , \30587 );
and \U$34514 ( \34858 , \34853 , \34857 );
and \U$34515 ( \34859 , \21813 , \30258 );
and \U$34516 ( \34860 , \21750 , \30256 );
nor \U$34517 ( \34861 , \34859 , \34860 );
xnor \U$34518 ( \34862 , \34861 , \29948 );
and \U$34519 ( \34863 , \34857 , \34862 );
and \U$34520 ( \34864 , \34853 , \34862 );
or \U$34521 ( \34865 , \34858 , \34863 , \34864 );
and \U$34522 ( \34866 , \34848 , \34865 );
and \U$34523 ( \34867 , \34832 , \34865 );
or \U$34524 ( \34868 , \34849 , \34866 , \34867 );
and \U$34525 ( \34869 , \34816 , \34868 );
and \U$34526 ( \34870 , \25604 , \24149 );
and \U$34527 ( \34871 , \25596 , \24147 );
nor \U$34528 ( \34872 , \34870 , \34871 );
xnor \U$34529 ( \34873 , \34872 , \23944 );
and \U$34530 ( \34874 , \26078 , \23743 );
and \U$34531 ( \34875 , \26073 , \23741 );
nor \U$34532 ( \34876 , \34874 , \34875 );
xnor \U$34533 ( \34877 , \34876 , \23594 );
and \U$34534 ( \34878 , \34873 , \34877 );
and \U$34535 ( \34879 , \26601 , \23421 );
and \U$34536 ( \34880 , \26342 , \23419 );
nor \U$34537 ( \34881 , \34879 , \34880 );
xnor \U$34538 ( \34882 , \34881 , \23279 );
and \U$34539 ( \34883 , \34877 , \34882 );
and \U$34540 ( \34884 , \34873 , \34882 );
or \U$34541 ( \34885 , \34878 , \34883 , \34884 );
and \U$34542 ( \34886 , \24714 , \25180 );
and \U$34543 ( \34887 , \24506 , \25178 );
nor \U$34544 ( \34888 , \34886 , \34887 );
xnor \U$34545 ( \34889 , \34888 , \25037 );
and \U$34546 ( \34890 , \24841 , \24857 );
and \U$34547 ( \34891 , \24836 , \24855 );
nor \U$34548 ( \34892 , \34890 , \34891 );
xnor \U$34549 ( \34893 , \34892 , \24611 );
and \U$34550 ( \34894 , \34889 , \34893 );
and \U$34551 ( \34895 , \25294 , \24462 );
and \U$34552 ( \34896 , \25097 , \24460 );
nor \U$34553 ( \34897 , \34895 , \34896 );
xnor \U$34554 ( \34898 , \34897 , \24275 );
and \U$34555 ( \34899 , \34893 , \34898 );
and \U$34556 ( \34900 , \34889 , \34898 );
or \U$34557 ( \34901 , \34894 , \34899 , \34900 );
and \U$34558 ( \34902 , \34885 , \34901 );
and \U$34559 ( \34903 , \23491 , \26471 );
and \U$34560 ( \34904 , \23466 , \26469 );
nor \U$34561 ( \34905 , \34903 , \34904 );
xnor \U$34562 ( \34906 , \34905 , \26230 );
and \U$34563 ( \34907 , \23832 , \26005 );
and \U$34564 ( \34908 , \23665 , \26003 );
nor \U$34565 ( \34909 , \34907 , \34908 );
xnor \U$34566 ( \34910 , \34909 , \25817 );
and \U$34567 ( \34911 , \34906 , \34910 );
and \U$34568 ( \34912 , \24089 , \25631 );
and \U$34569 ( \34913 , \23970 , \25629 );
nor \U$34570 ( \34914 , \34912 , \34913 );
xnor \U$34571 ( \34915 , \34914 , \25399 );
and \U$34572 ( \34916 , \34910 , \34915 );
and \U$34573 ( \34917 , \34906 , \34915 );
or \U$34574 ( \34918 , \34911 , \34916 , \34917 );
and \U$34575 ( \34919 , \34901 , \34918 );
and \U$34576 ( \34920 , \34885 , \34918 );
or \U$34577 ( \34921 , \34902 , \34919 , \34920 );
and \U$34578 ( \34922 , \34868 , \34921 );
and \U$34579 ( \34923 , \34816 , \34921 );
or \U$34580 ( \34924 , \34869 , \34922 , \34923 );
and \U$34581 ( \34925 , \34764 , \34924 );
xor \U$34582 ( \34926 , \34341 , \34345 );
xor \U$34583 ( \34927 , \34926 , \34350 );
xor \U$34584 ( \34928 , \34454 , \34456 );
xor \U$34585 ( \34929 , \34928 , \34459 );
and \U$34586 ( \34930 , \34927 , \34929 );
xor \U$34587 ( \34931 , \34464 , \34466 );
xor \U$34588 ( \34932 , \34931 , \34469 );
and \U$34589 ( \34933 , \34929 , \34932 );
and \U$34590 ( \34934 , \34927 , \34932 );
or \U$34591 ( \34935 , \34930 , \34933 , \34934 );
and \U$34592 ( \34936 , \34924 , \34935 );
and \U$34593 ( \34937 , \34764 , \34935 );
or \U$34594 ( \34938 , \34925 , \34936 , \34937 );
xor \U$34595 ( \34939 , \34552 , \34568 );
xor \U$34596 ( \34940 , \34939 , \34585 );
xor \U$34597 ( \34941 , \34605 , \34621 );
xor \U$34598 ( \34942 , \34941 , \34638 );
and \U$34599 ( \34943 , \34940 , \34942 );
xor \U$34600 ( \34944 , \34477 , \34479 );
xor \U$34601 ( \34945 , \34944 , \34482 );
and \U$34602 ( \34946 , \34942 , \34945 );
and \U$34603 ( \34947 , \34940 , \34945 );
or \U$34604 ( \34948 , \34943 , \34946 , \34947 );
xor \U$34605 ( \34949 , \34337 , \34353 );
xor \U$34606 ( \34950 , \34949 , \34370 );
and \U$34607 ( \34951 , \34948 , \34950 );
xor \U$34608 ( \34952 , \34660 , \34662 );
xor \U$34609 ( \34953 , \34952 , \34665 );
and \U$34610 ( \34954 , \34950 , \34953 );
and \U$34611 ( \34955 , \34948 , \34953 );
or \U$34612 ( \34956 , \34951 , \34954 , \34955 );
and \U$34613 ( \34957 , \34938 , \34956 );
xor \U$34614 ( \34958 , \34462 , \34472 );
xor \U$34615 ( \34959 , \34958 , \34485 );
xor \U$34616 ( \34960 , \34536 , \34588 );
xor \U$34617 ( \34961 , \34960 , \34641 );
and \U$34618 ( \34962 , \34959 , \34961 );
xor \U$34619 ( \34963 , \34647 , \34649 );
xor \U$34620 ( \34964 , \34963 , \34652 );
and \U$34621 ( \34965 , \34961 , \34964 );
and \U$34622 ( \34966 , \34959 , \34964 );
or \U$34623 ( \34967 , \34962 , \34965 , \34966 );
and \U$34624 ( \34968 , \34956 , \34967 );
and \U$34625 ( \34969 , \34938 , \34967 );
or \U$34626 ( \34970 , \34957 , \34968 , \34969 );
xor \U$34627 ( \34971 , \34488 , \34644 );
xor \U$34628 ( \34972 , \34971 , \34655 );
xor \U$34629 ( \34973 , \34668 , \34670 );
xor \U$34630 ( \34974 , \34973 , \34673 );
and \U$34631 ( \34975 , \34972 , \34974 );
xor \U$34632 ( \34976 , \34679 , \34681 );
xor \U$34633 ( \34977 , \34976 , \34684 );
and \U$34634 ( \34978 , \34974 , \34977 );
and \U$34635 ( \34979 , \34972 , \34977 );
or \U$34636 ( \34980 , \34975 , \34978 , \34979 );
and \U$34637 ( \34981 , \34970 , \34980 );
xor \U$34638 ( \34982 , \34692 , \34694 );
xor \U$34639 ( \34983 , \34982 , \34697 );
and \U$34640 ( \34984 , \34980 , \34983 );
and \U$34641 ( \34985 , \34970 , \34983 );
or \U$34642 ( \34986 , \34981 , \34984 , \34985 );
xor \U$34643 ( \34987 , \34690 , \34700 );
xor \U$34644 ( \34988 , \34987 , \34703 );
and \U$34645 ( \34989 , \34986 , \34988 );
xor \U$34646 ( \34990 , \34708 , \34710 );
xor \U$34647 ( \34991 , \34990 , \34713 );
and \U$34648 ( \34992 , \34988 , \34991 );
and \U$34649 ( \34993 , \34986 , \34991 );
or \U$34650 ( \34994 , \34989 , \34992 , \34993 );
xor \U$34651 ( \34995 , \34706 , \34716 );
xor \U$34652 ( \34996 , \34995 , \34719 );
and \U$34653 ( \34997 , \34994 , \34996 );
xor \U$34654 ( \34998 , \34422 , \34432 );
xor \U$34655 ( \34999 , \34998 , \34435 );
and \U$34656 ( \35000 , \34996 , \34999 );
and \U$34657 ( \35001 , \34994 , \34999 );
or \U$34658 ( \35002 , \34997 , \35000 , \35001 );
and \U$34659 ( \35003 , \34728 , \35002 );
xor \U$34660 ( \35004 , \34728 , \35002 );
xor \U$34661 ( \35005 , \34994 , \34996 );
xor \U$34662 ( \35006 , \35005 , \34999 );
xor \U$34663 ( \35007 , \34873 , \34877 );
xor \U$34664 ( \35008 , \35007 , \34882 );
xor \U$34665 ( \35009 , \34889 , \34893 );
xor \U$34666 ( \35010 , \35009 , \34898 );
and \U$34667 ( \35011 , \35008 , \35010 );
xor \U$34668 ( \35012 , \34906 , \34910 );
xor \U$34669 ( \35013 , \35012 , \34915 );
and \U$34670 ( \35014 , \35010 , \35013 );
and \U$34671 ( \35015 , \35008 , \35013 );
or \U$34672 ( \35016 , \35011 , \35014 , \35015 );
xor \U$34673 ( \35017 , \34768 , \34772 );
xor \U$34674 ( \35018 , \35017 , \34777 );
xor \U$34675 ( \35019 , \34784 , \34788 );
xor \U$34676 ( \35020 , \35019 , \34793 );
and \U$34677 ( \35021 , \35018 , \35020 );
xor \U$34678 ( \35022 , \34801 , \34805 );
xor \U$34679 ( \35023 , \35022 , \34810 );
and \U$34680 ( \35024 , \35020 , \35023 );
and \U$34681 ( \35025 , \35018 , \35023 );
or \U$34682 ( \35026 , \35021 , \35024 , \35025 );
and \U$34683 ( \35027 , \35016 , \35026 );
xor \U$34684 ( \35028 , \34820 , \34824 );
xor \U$34685 ( \35029 , \35028 , \34829 );
xor \U$34686 ( \35030 , \34836 , \34840 );
xor \U$34687 ( \35031 , \35030 , \34845 );
and \U$34688 ( \35032 , \35029 , \35031 );
xor \U$34689 ( \35033 , \34853 , \34857 );
xor \U$34690 ( \35034 , \35033 , \34862 );
and \U$34691 ( \35035 , \35031 , \35034 );
and \U$34692 ( \35036 , \35029 , \35034 );
or \U$34693 ( \35037 , \35032 , \35035 , \35036 );
and \U$34694 ( \35038 , \35026 , \35037 );
and \U$34695 ( \35039 , \35016 , \35037 );
or \U$34696 ( \35040 , \35027 , \35038 , \35039 );
and \U$34697 ( \35041 , \25596 , \24462 );
and \U$34698 ( \35042 , \25294 , \24460 );
nor \U$34699 ( \35043 , \35041 , \35042 );
xnor \U$34700 ( \35044 , \35043 , \24275 );
and \U$34701 ( \35045 , \26073 , \24149 );
and \U$34702 ( \35046 , \25604 , \24147 );
nor \U$34703 ( \35047 , \35045 , \35046 );
xnor \U$34704 ( \35048 , \35047 , \23944 );
and \U$34705 ( \35049 , \35044 , \35048 );
and \U$34706 ( \35050 , \26342 , \23743 );
and \U$34707 ( \35051 , \26078 , \23741 );
nor \U$34708 ( \35052 , \35050 , \35051 );
xnor \U$34709 ( \35053 , \35052 , \23594 );
and \U$34710 ( \35054 , \35048 , \35053 );
and \U$34711 ( \35055 , \35044 , \35053 );
or \U$34712 ( \35056 , \35049 , \35054 , \35055 );
and \U$34713 ( \35057 , \23466 , \27060 );
and \U$34714 ( \35058 , \23202 , \27058 );
nor \U$34715 ( \35059 , \35057 , \35058 );
xnor \U$34716 ( \35060 , \35059 , \26720 );
and \U$34717 ( \35061 , \23665 , \26471 );
and \U$34718 ( \35062 , \23491 , \26469 );
nor \U$34719 ( \35063 , \35061 , \35062 );
xnor \U$34720 ( \35064 , \35063 , \26230 );
and \U$34721 ( \35065 , \35060 , \35064 );
and \U$34722 ( \35066 , \23970 , \26005 );
and \U$34723 ( \35067 , \23832 , \26003 );
nor \U$34724 ( \35068 , \35066 , \35067 );
xnor \U$34725 ( \35069 , \35068 , \25817 );
and \U$34726 ( \35070 , \35064 , \35069 );
and \U$34727 ( \35071 , \35060 , \35069 );
or \U$34728 ( \35072 , \35065 , \35070 , \35071 );
and \U$34729 ( \35073 , \35056 , \35072 );
and \U$34730 ( \35074 , \24506 , \25631 );
and \U$34731 ( \35075 , \24089 , \25629 );
nor \U$34732 ( \35076 , \35074 , \35075 );
xnor \U$34733 ( \35077 , \35076 , \25399 );
and \U$34734 ( \35078 , \24836 , \25180 );
and \U$34735 ( \35079 , \24714 , \25178 );
nor \U$34736 ( \35080 , \35078 , \35079 );
xnor \U$34737 ( \35081 , \35080 , \25037 );
and \U$34738 ( \35082 , \35077 , \35081 );
and \U$34739 ( \35083 , \25097 , \24857 );
and \U$34740 ( \35084 , \24841 , \24855 );
nor \U$34741 ( \35085 , \35083 , \35084 );
xnor \U$34742 ( \35086 , \35085 , \24611 );
and \U$34743 ( \35087 , \35081 , \35086 );
and \U$34744 ( \35088 , \35077 , \35086 );
or \U$34745 ( \35089 , \35082 , \35087 , \35088 );
and \U$34746 ( \35090 , \35072 , \35089 );
and \U$34747 ( \35091 , \35056 , \35089 );
or \U$34748 ( \35092 , \35073 , \35090 , \35091 );
and \U$34749 ( \35093 , \22011 , \30258 );
and \U$34750 ( \35094 , \21813 , \30256 );
nor \U$34751 ( \35095 , \35093 , \35094 );
xnor \U$34752 ( \35096 , \35095 , \29948 );
and \U$34753 ( \35097 , \22204 , \29721 );
and \U$34754 ( \35098 , \22099 , \29719 );
nor \U$34755 ( \35099 , \35097 , \35098 );
xnor \U$34756 ( \35100 , \35099 , \29350 );
and \U$34757 ( \35101 , \35096 , \35100 );
and \U$34758 ( \35102 , \22325 , \29159 );
and \U$34759 ( \35103 , \22209 , \29157 );
nor \U$34760 ( \35104 , \35102 , \35103 );
xnor \U$34761 ( \35105 , \35104 , \28841 );
and \U$34762 ( \35106 , \35100 , \35105 );
and \U$34763 ( \35107 , \35096 , \35105 );
or \U$34764 ( \35108 , \35101 , \35106 , \35107 );
and \U$34765 ( \35109 , \21478 , \31639 );
and \U$34766 ( \35110 , \21463 , \31636 );
nor \U$34767 ( \35111 , \35109 , \35110 );
xnor \U$34768 ( \35112 , \35111 , \30584 );
and \U$34769 ( \35113 , \21750 , \30826 );
and \U$34770 ( \35114 , \21689 , \30824 );
nor \U$34771 ( \35115 , \35113 , \35114 );
xnor \U$34772 ( \35116 , \35115 , \30587 );
and \U$34773 ( \35117 , \35112 , \35116 );
and \U$34774 ( \35118 , \35116 , \21392 );
and \U$34775 ( \35119 , \35112 , \21392 );
or \U$34776 ( \35120 , \35117 , \35118 , \35119 );
and \U$34777 ( \35121 , \35108 , \35120 );
and \U$34778 ( \35122 , \22616 , \28592 );
and \U$34779 ( \35123 , \22440 , \28590 );
nor \U$34780 ( \35124 , \35122 , \35123 );
xnor \U$34781 ( \35125 , \35124 , \28343 );
and \U$34782 ( \35126 , \22867 , \28063 );
and \U$34783 ( \35127 , \22624 , \28061 );
nor \U$34784 ( \35128 , \35126 , \35127 );
xnor \U$34785 ( \35129 , \35128 , \27803 );
and \U$34786 ( \35130 , \35125 , \35129 );
and \U$34787 ( \35131 , \23058 , \27569 );
and \U$34788 ( \35132 , \22872 , \27567 );
nor \U$34789 ( \35133 , \35131 , \35132 );
xnor \U$34790 ( \35134 , \35133 , \27254 );
and \U$34791 ( \35135 , \35129 , \35134 );
and \U$34792 ( \35136 , \35125 , \35134 );
or \U$34793 ( \35137 , \35130 , \35135 , \35136 );
and \U$34794 ( \35138 , \35120 , \35137 );
and \U$34795 ( \35139 , \35108 , \35137 );
or \U$34796 ( \35140 , \35121 , \35138 , \35139 );
and \U$34797 ( \35141 , \35092 , \35140 );
and \U$34798 ( \35142 , \30375 , \21985 );
and \U$34799 ( \35143 , \29806 , \21983 );
nor \U$34800 ( \35144 , \35142 , \35143 );
xnor \U$34801 ( \35145 , \35144 , \21907 );
and \U$34802 ( \35146 , \30986 , \21821 );
and \U$34803 ( \35147 , \30383 , \21819 );
nor \U$34804 ( \35148 , \35146 , \35147 );
xnor \U$34805 ( \35149 , \35148 , \21727 );
and \U$34806 ( \35150 , \35145 , \35149 );
and \U$34807 ( \35151 , \31172 , \21652 );
and \U$34808 ( \35152 , \30991 , \21650 );
nor \U$34809 ( \35153 , \35151 , \35152 );
xnor \U$34810 ( \35154 , \35153 , \21377 );
and \U$34811 ( \35155 , \35149 , \35154 );
and \U$34812 ( \35156 , \35145 , \35154 );
or \U$34813 ( \35157 , \35150 , \35155 , \35156 );
and \U$34814 ( \35158 , \26973 , \23421 );
and \U$34815 ( \35159 , \26601 , \23419 );
nor \U$34816 ( \35160 , \35158 , \35159 );
xnor \U$34817 ( \35161 , \35160 , \23279 );
and \U$34818 ( \35162 , \27325 , \23125 );
and \U$34819 ( \35163 , \26982 , \23123 );
nor \U$34820 ( \35164 , \35162 , \35163 );
xnor \U$34821 ( \35165 , \35164 , \22988 );
and \U$34822 ( \35166 , \35161 , \35165 );
and \U$34823 ( \35167 , \27830 , \22919 );
and \U$34824 ( \35168 , \27527 , \22917 );
nor \U$34825 ( \35169 , \35167 , \35168 );
xnor \U$34826 ( \35170 , \35169 , \22767 );
and \U$34827 ( \35171 , \35165 , \35170 );
and \U$34828 ( \35172 , \35161 , \35170 );
or \U$34829 ( \35173 , \35166 , \35171 , \35172 );
and \U$34830 ( \35174 , \35157 , \35173 );
and \U$34831 ( \35175 , \28528 , \22651 );
and \U$34832 ( \35176 , \28002 , \22649 );
nor \U$34833 ( \35177 , \35175 , \35176 );
xnor \U$34834 ( \35178 , \35177 , \22495 );
and \U$34835 ( \35179 , \29198 , \22379 );
and \U$34836 ( \35180 , \28952 , \22377 );
nor \U$34837 ( \35181 , \35179 , \35180 );
xnor \U$34838 ( \35182 , \35181 , \22266 );
and \U$34839 ( \35183 , \35178 , \35182 );
and \U$34840 ( \35184 , \29522 , \22185 );
and \U$34841 ( \35185 , \29203 , \22183 );
nor \U$34842 ( \35186 , \35184 , \35185 );
xnor \U$34843 ( \35187 , \35186 , \22049 );
and \U$34844 ( \35188 , \35182 , \35187 );
and \U$34845 ( \35189 , \35178 , \35187 );
or \U$34846 ( \35190 , \35183 , \35188 , \35189 );
and \U$34847 ( \35191 , \35173 , \35190 );
and \U$34848 ( \35192 , \35157 , \35190 );
or \U$34849 ( \35193 , \35174 , \35191 , \35192 );
and \U$34850 ( \35194 , \35140 , \35193 );
and \U$34851 ( \35195 , \35092 , \35193 );
or \U$34852 ( \35196 , \35141 , \35194 , \35195 );
and \U$34853 ( \35197 , \35040 , \35196 );
xor \U$34854 ( \35198 , \34508 , \34512 );
xor \U$34855 ( \35199 , \35198 , \34517 );
xor \U$34856 ( \35200 , \34525 , \34529 );
xor \U$34857 ( \35201 , \35200 , \21408 );
and \U$34858 ( \35202 , \35199 , \35201 );
xor \U$34859 ( \35203 , \34753 , \34755 );
xor \U$34860 ( \35204 , \35203 , \34758 );
and \U$34861 ( \35205 , \35201 , \35204 );
and \U$34862 ( \35206 , \35199 , \35204 );
or \U$34863 ( \35207 , \35202 , \35205 , \35206 );
and \U$34864 ( \35208 , \35196 , \35207 );
and \U$34865 ( \35209 , \35040 , \35207 );
or \U$34866 ( \35210 , \35197 , \35208 , \35209 );
xor \U$34867 ( \35211 , \34780 , \34796 );
xor \U$34868 ( \35212 , \35211 , \34813 );
xor \U$34869 ( \35213 , \34730 , \34732 );
xor \U$34870 ( \35214 , \35213 , \34735 );
and \U$34871 ( \35215 , \35212 , \35214 );
xor \U$34872 ( \35216 , \34742 , \34744 );
xor \U$34873 ( \35217 , \35216 , \34747 );
and \U$34874 ( \35218 , \35214 , \35217 );
and \U$34875 ( \35219 , \35212 , \35217 );
or \U$34876 ( \35220 , \35215 , \35218 , \35219 );
xor \U$34877 ( \35221 , \34832 , \34848 );
xor \U$34878 ( \35222 , \35221 , \34865 );
xor \U$34879 ( \35223 , \34885 , \34901 );
xor \U$34880 ( \35224 , \35223 , \34918 );
and \U$34881 ( \35225 , \35222 , \35224 );
and \U$34882 ( \35226 , \35220 , \35225 );
xor \U$34883 ( \35227 , \34504 , \34520 );
xor \U$34884 ( \35228 , \35227 , \34533 );
and \U$34885 ( \35229 , \35225 , \35228 );
and \U$34886 ( \35230 , \35220 , \35228 );
or \U$34887 ( \35231 , \35226 , \35229 , \35230 );
and \U$34888 ( \35232 , \35210 , \35231 );
xor \U$34889 ( \35233 , \34738 , \34750 );
xor \U$34890 ( \35234 , \35233 , \34761 );
xor \U$34891 ( \35235 , \34940 , \34942 );
xor \U$34892 ( \35236 , \35235 , \34945 );
and \U$34893 ( \35237 , \35234 , \35236 );
xor \U$34894 ( \35238 , \34927 , \34929 );
xor \U$34895 ( \35239 , \35238 , \34932 );
and \U$34896 ( \35240 , \35236 , \35239 );
and \U$34897 ( \35241 , \35234 , \35239 );
or \U$34898 ( \35242 , \35237 , \35240 , \35241 );
and \U$34899 ( \35243 , \35231 , \35242 );
and \U$34900 ( \35244 , \35210 , \35242 );
or \U$34901 ( \35245 , \35232 , \35243 , \35244 );
xor \U$34902 ( \35246 , \34764 , \34924 );
xor \U$34903 ( \35247 , \35246 , \34935 );
xor \U$34904 ( \35248 , \34948 , \34950 );
xor \U$34905 ( \35249 , \35248 , \34953 );
and \U$34906 ( \35250 , \35247 , \35249 );
xor \U$34907 ( \35251 , \34959 , \34961 );
xor \U$34908 ( \35252 , \35251 , \34964 );
and \U$34909 ( \35253 , \35249 , \35252 );
and \U$34910 ( \35254 , \35247 , \35252 );
or \U$34911 ( \35255 , \35250 , \35253 , \35254 );
and \U$34912 ( \35256 , \35245 , \35255 );
xor \U$34913 ( \35257 , \34972 , \34974 );
xor \U$34914 ( \35258 , \35257 , \34977 );
and \U$34915 ( \35259 , \35255 , \35258 );
and \U$34916 ( \35260 , \35245 , \35258 );
or \U$34917 ( \35261 , \35256 , \35259 , \35260 );
xor \U$34918 ( \35262 , \34658 , \34676 );
xor \U$34919 ( \35263 , \35262 , \34687 );
and \U$34920 ( \35264 , \35261 , \35263 );
xor \U$34921 ( \35265 , \34970 , \34980 );
xor \U$34922 ( \35266 , \35265 , \34983 );
and \U$34923 ( \35267 , \35263 , \35266 );
and \U$34924 ( \35268 , \35261 , \35266 );
or \U$34925 ( \35269 , \35264 , \35267 , \35268 );
xor \U$34926 ( \35270 , \34986 , \34988 );
xor \U$34927 ( \35271 , \35270 , \34991 );
and \U$34928 ( \35272 , \35269 , \35271 );
and \U$34929 ( \35273 , \35006 , \35272 );
xor \U$34930 ( \35274 , \35006 , \35272 );
xor \U$34931 ( \35275 , \35269 , \35271 );
and \U$34932 ( \35276 , \24841 , \25180 );
and \U$34933 ( \35277 , \24836 , \25178 );
nor \U$34934 ( \35278 , \35276 , \35277 );
xnor \U$34935 ( \35279 , \35278 , \25037 );
and \U$34936 ( \35280 , \25294 , \24857 );
and \U$34937 ( \35281 , \25097 , \24855 );
nor \U$34938 ( \35282 , \35280 , \35281 );
xnor \U$34939 ( \35283 , \35282 , \24611 );
and \U$34940 ( \35284 , \35279 , \35283 );
and \U$34941 ( \35285 , \25604 , \24462 );
and \U$34942 ( \35286 , \25596 , \24460 );
nor \U$34943 ( \35287 , \35285 , \35286 );
xnor \U$34944 ( \35288 , \35287 , \24275 );
and \U$34945 ( \35289 , \35283 , \35288 );
and \U$34946 ( \35290 , \35279 , \35288 );
or \U$34947 ( \35291 , \35284 , \35289 , \35290 );
and \U$34948 ( \35292 , \23832 , \26471 );
and \U$34949 ( \35293 , \23665 , \26469 );
nor \U$34950 ( \35294 , \35292 , \35293 );
xnor \U$34951 ( \35295 , \35294 , \26230 );
and \U$34952 ( \35296 , \24089 , \26005 );
and \U$34953 ( \35297 , \23970 , \26003 );
nor \U$34954 ( \35298 , \35296 , \35297 );
xnor \U$34955 ( \35299 , \35298 , \25817 );
and \U$34956 ( \35300 , \35295 , \35299 );
and \U$34957 ( \35301 , \24714 , \25631 );
and \U$34958 ( \35302 , \24506 , \25629 );
nor \U$34959 ( \35303 , \35301 , \35302 );
xnor \U$34960 ( \35304 , \35303 , \25399 );
and \U$34961 ( \35305 , \35299 , \35304 );
and \U$34962 ( \35306 , \35295 , \35304 );
or \U$34963 ( \35307 , \35300 , \35305 , \35306 );
and \U$34964 ( \35308 , \35291 , \35307 );
and \U$34965 ( \35309 , \26078 , \24149 );
and \U$34966 ( \35310 , \26073 , \24147 );
nor \U$34967 ( \35311 , \35309 , \35310 );
xnor \U$34968 ( \35312 , \35311 , \23944 );
and \U$34969 ( \35313 , \26601 , \23743 );
and \U$34970 ( \35314 , \26342 , \23741 );
nor \U$34971 ( \35315 , \35313 , \35314 );
xnor \U$34972 ( \35316 , \35315 , \23594 );
and \U$34973 ( \35317 , \35312 , \35316 );
and \U$34974 ( \35318 , \26982 , \23421 );
and \U$34975 ( \35319 , \26973 , \23419 );
nor \U$34976 ( \35320 , \35318 , \35319 );
xnor \U$34977 ( \35321 , \35320 , \23279 );
and \U$34978 ( \35322 , \35316 , \35321 );
and \U$34979 ( \35323 , \35312 , \35321 );
or \U$34980 ( \35324 , \35317 , \35322 , \35323 );
and \U$34981 ( \35325 , \35307 , \35324 );
and \U$34982 ( \35326 , \35291 , \35324 );
or \U$34983 ( \35327 , \35308 , \35325 , \35326 );
and \U$34984 ( \35328 , \29203 , \22379 );
and \U$34985 ( \35329 , \29198 , \22377 );
nor \U$34986 ( \35330 , \35328 , \35329 );
xnor \U$34987 ( \35331 , \35330 , \22266 );
and \U$34988 ( \35332 , \29806 , \22185 );
and \U$34989 ( \35333 , \29522 , \22183 );
nor \U$34990 ( \35334 , \35332 , \35333 );
xnor \U$34991 ( \35335 , \35334 , \22049 );
and \U$34992 ( \35336 , \35331 , \35335 );
and \U$34993 ( \35337 , \30383 , \21985 );
and \U$34994 ( \35338 , \30375 , \21983 );
nor \U$34995 ( \35339 , \35337 , \35338 );
xnor \U$34996 ( \35340 , \35339 , \21907 );
and \U$34997 ( \35341 , \35335 , \35340 );
and \U$34998 ( \35342 , \35331 , \35340 );
or \U$34999 ( \35343 , \35336 , \35341 , \35342 );
and \U$35000 ( \35344 , \27527 , \23125 );
and \U$35001 ( \35345 , \27325 , \23123 );
nor \U$35002 ( \35346 , \35344 , \35345 );
xnor \U$35003 ( \35347 , \35346 , \22988 );
and \U$35004 ( \35348 , \28002 , \22919 );
and \U$35005 ( \35349 , \27830 , \22917 );
nor \U$35006 ( \35350 , \35348 , \35349 );
xnor \U$35007 ( \35351 , \35350 , \22767 );
and \U$35008 ( \35352 , \35347 , \35351 );
and \U$35009 ( \35353 , \28952 , \22651 );
and \U$35010 ( \35354 , \28528 , \22649 );
nor \U$35011 ( \35355 , \35353 , \35354 );
xnor \U$35012 ( \35356 , \35355 , \22495 );
and \U$35013 ( \35357 , \35351 , \35356 );
and \U$35014 ( \35358 , \35347 , \35356 );
or \U$35015 ( \35359 , \35352 , \35357 , \35358 );
and \U$35016 ( \35360 , \35343 , \35359 );
and \U$35017 ( \35361 , \30991 , \21821 );
and \U$35018 ( \35362 , \30986 , \21819 );
nor \U$35019 ( \35363 , \35361 , \35362 );
xnor \U$35020 ( \35364 , \35363 , \21727 );
and \U$35021 ( \35365 , \31792 , \21652 );
and \U$35022 ( \35366 , \31172 , \21650 );
nor \U$35023 ( \35367 , \35365 , \35366 );
xnor \U$35024 ( \35368 , \35367 , \21377 );
and \U$35025 ( \35369 , \35364 , \35368 );
and \U$35026 ( \35370 , \35359 , \35369 );
and \U$35027 ( \35371 , \35343 , \35369 );
or \U$35028 ( \35372 , \35360 , \35370 , \35371 );
and \U$35029 ( \35373 , \35327 , \35372 );
and \U$35030 ( \35374 , \22872 , \28063 );
and \U$35031 ( \35375 , \22867 , \28061 );
nor \U$35032 ( \35376 , \35374 , \35375 );
xnor \U$35033 ( \35377 , \35376 , \27803 );
and \U$35034 ( \35378 , \23202 , \27569 );
and \U$35035 ( \35379 , \23058 , \27567 );
nor \U$35036 ( \35380 , \35378 , \35379 );
xnor \U$35037 ( \35381 , \35380 , \27254 );
and \U$35038 ( \35382 , \35377 , \35381 );
and \U$35039 ( \35383 , \23491 , \27060 );
and \U$35040 ( \35384 , \23466 , \27058 );
nor \U$35041 ( \35385 , \35383 , \35384 );
xnor \U$35042 ( \35386 , \35385 , \26720 );
and \U$35043 ( \35387 , \35381 , \35386 );
and \U$35044 ( \35388 , \35377 , \35386 );
or \U$35045 ( \35389 , \35382 , \35387 , \35388 );
and \U$35046 ( \35390 , \21689 , \31639 );
and \U$35047 ( \35391 , \21478 , \31636 );
nor \U$35048 ( \35392 , \35390 , \35391 );
xnor \U$35049 ( \35393 , \35392 , \30584 );
and \U$35050 ( \35394 , \21813 , \30826 );
and \U$35051 ( \35395 , \21750 , \30824 );
nor \U$35052 ( \35396 , \35394 , \35395 );
xnor \U$35053 ( \35397 , \35396 , \30587 );
and \U$35054 ( \35398 , \35393 , \35397 );
and \U$35055 ( \35399 , \22099 , \30258 );
and \U$35056 ( \35400 , \22011 , \30256 );
nor \U$35057 ( \35401 , \35399 , \35400 );
xnor \U$35058 ( \35402 , \35401 , \29948 );
and \U$35059 ( \35403 , \35397 , \35402 );
and \U$35060 ( \35404 , \35393 , \35402 );
or \U$35061 ( \35405 , \35398 , \35403 , \35404 );
and \U$35062 ( \35406 , \35389 , \35405 );
and \U$35063 ( \35407 , \22209 , \29721 );
and \U$35064 ( \35408 , \22204 , \29719 );
nor \U$35065 ( \35409 , \35407 , \35408 );
xnor \U$35066 ( \35410 , \35409 , \29350 );
and \U$35067 ( \35411 , \22440 , \29159 );
and \U$35068 ( \35412 , \22325 , \29157 );
nor \U$35069 ( \35413 , \35411 , \35412 );
xnor \U$35070 ( \35414 , \35413 , \28841 );
and \U$35071 ( \35415 , \35410 , \35414 );
and \U$35072 ( \35416 , \22624 , \28592 );
and \U$35073 ( \35417 , \22616 , \28590 );
nor \U$35074 ( \35418 , \35416 , \35417 );
xnor \U$35075 ( \35419 , \35418 , \28343 );
and \U$35076 ( \35420 , \35414 , \35419 );
and \U$35077 ( \35421 , \35410 , \35419 );
or \U$35078 ( \35422 , \35415 , \35420 , \35421 );
and \U$35079 ( \35423 , \35405 , \35422 );
and \U$35080 ( \35424 , \35389 , \35422 );
or \U$35081 ( \35425 , \35406 , \35423 , \35424 );
and \U$35082 ( \35426 , \35372 , \35425 );
and \U$35083 ( \35427 , \35327 , \35425 );
or \U$35084 ( \35428 , \35373 , \35426 , \35427 );
xor \U$35085 ( \35429 , \35096 , \35100 );
xor \U$35086 ( \35430 , \35429 , \35105 );
xor \U$35087 ( \35431 , \35125 , \35129 );
xor \U$35088 ( \35432 , \35431 , \35134 );
and \U$35089 ( \35433 , \35430 , \35432 );
xor \U$35090 ( \35434 , \35060 , \35064 );
xor \U$35091 ( \35435 , \35434 , \35069 );
and \U$35092 ( \35436 , \35432 , \35435 );
and \U$35093 ( \35437 , \35430 , \35435 );
or \U$35094 ( \35438 , \35433 , \35436 , \35437 );
nand \U$35095 ( \35439 , \31792 , \21383 );
xnor \U$35096 ( \35440 , \35439 , \21392 );
xor \U$35097 ( \35441 , \35145 , \35149 );
xor \U$35098 ( \35442 , \35441 , \35154 );
and \U$35099 ( \35443 , \35440 , \35442 );
xor \U$35100 ( \35444 , \35178 , \35182 );
xor \U$35101 ( \35445 , \35444 , \35187 );
and \U$35102 ( \35446 , \35442 , \35445 );
and \U$35103 ( \35447 , \35440 , \35445 );
or \U$35104 ( \35448 , \35443 , \35446 , \35447 );
and \U$35105 ( \35449 , \35438 , \35448 );
xor \U$35106 ( \35450 , \35161 , \35165 );
xor \U$35107 ( \35451 , \35450 , \35170 );
xor \U$35108 ( \35452 , \35044 , \35048 );
xor \U$35109 ( \35453 , \35452 , \35053 );
and \U$35110 ( \35454 , \35451 , \35453 );
xor \U$35111 ( \35455 , \35077 , \35081 );
xor \U$35112 ( \35456 , \35455 , \35086 );
and \U$35113 ( \35457 , \35453 , \35456 );
and \U$35114 ( \35458 , \35451 , \35456 );
or \U$35115 ( \35459 , \35454 , \35457 , \35458 );
and \U$35116 ( \35460 , \35448 , \35459 );
and \U$35117 ( \35461 , \35438 , \35459 );
or \U$35118 ( \35462 , \35449 , \35460 , \35461 );
and \U$35119 ( \35463 , \35428 , \35462 );
xor \U$35120 ( \35464 , \35008 , \35010 );
xor \U$35121 ( \35465 , \35464 , \35013 );
xor \U$35122 ( \35466 , \35018 , \35020 );
xor \U$35123 ( \35467 , \35466 , \35023 );
and \U$35124 ( \35468 , \35465 , \35467 );
xor \U$35125 ( \35469 , \35029 , \35031 );
xor \U$35126 ( \35470 , \35469 , \35034 );
and \U$35127 ( \35471 , \35467 , \35470 );
and \U$35128 ( \35472 , \35465 , \35470 );
or \U$35129 ( \35473 , \35468 , \35471 , \35472 );
and \U$35130 ( \35474 , \35462 , \35473 );
and \U$35131 ( \35475 , \35428 , \35473 );
or \U$35132 ( \35476 , \35463 , \35474 , \35475 );
xor \U$35133 ( \35477 , \35016 , \35026 );
xor \U$35134 ( \35478 , \35477 , \35037 );
xor \U$35135 ( \35479 , \35092 , \35140 );
xor \U$35136 ( \35480 , \35479 , \35193 );
and \U$35137 ( \35481 , \35478 , \35480 );
xor \U$35138 ( \35482 , \35199 , \35201 );
xor \U$35139 ( \35483 , \35482 , \35204 );
and \U$35140 ( \35484 , \35480 , \35483 );
and \U$35141 ( \35485 , \35478 , \35483 );
or \U$35142 ( \35486 , \35481 , \35484 , \35485 );
and \U$35143 ( \35487 , \35476 , \35486 );
xor \U$35144 ( \35488 , \35056 , \35072 );
xor \U$35145 ( \35489 , \35488 , \35089 );
xor \U$35146 ( \35490 , \35108 , \35120 );
xor \U$35147 ( \35491 , \35490 , \35137 );
and \U$35148 ( \35492 , \35489 , \35491 );
xor \U$35149 ( \35493 , \35157 , \35173 );
xor \U$35150 ( \35494 , \35493 , \35190 );
and \U$35151 ( \35495 , \35491 , \35494 );
and \U$35152 ( \35496 , \35489 , \35494 );
or \U$35153 ( \35497 , \35492 , \35495 , \35496 );
xor \U$35154 ( \35498 , \35212 , \35214 );
xor \U$35155 ( \35499 , \35498 , \35217 );
and \U$35156 ( \35500 , \35497 , \35499 );
xor \U$35157 ( \35501 , \35222 , \35224 );
and \U$35158 ( \35502 , \35499 , \35501 );
and \U$35159 ( \35503 , \35497 , \35501 );
or \U$35160 ( \35504 , \35500 , \35502 , \35503 );
and \U$35161 ( \35505 , \35486 , \35504 );
and \U$35162 ( \35506 , \35476 , \35504 );
or \U$35163 ( \35507 , \35487 , \35505 , \35506 );
xor \U$35164 ( \35508 , \34816 , \34868 );
xor \U$35165 ( \35509 , \35508 , \34921 );
xor \U$35166 ( \35510 , \35220 , \35225 );
xor \U$35167 ( \35511 , \35510 , \35228 );
and \U$35168 ( \35512 , \35509 , \35511 );
xor \U$35169 ( \35513 , \35234 , \35236 );
xor \U$35170 ( \35514 , \35513 , \35239 );
and \U$35171 ( \35515 , \35511 , \35514 );
and \U$35172 ( \35516 , \35509 , \35514 );
or \U$35173 ( \35517 , \35512 , \35515 , \35516 );
and \U$35174 ( \35518 , \35507 , \35517 );
xor \U$35175 ( \35519 , \35247 , \35249 );
xor \U$35176 ( \35520 , \35519 , \35252 );
and \U$35177 ( \35521 , \35517 , \35520 );
and \U$35178 ( \35522 , \35507 , \35520 );
or \U$35179 ( \35523 , \35518 , \35521 , \35522 );
xor \U$35180 ( \35524 , \34938 , \34956 );
xor \U$35181 ( \35525 , \35524 , \34967 );
and \U$35182 ( \35526 , \35523 , \35525 );
xor \U$35183 ( \35527 , \35245 , \35255 );
xor \U$35184 ( \35528 , \35527 , \35258 );
and \U$35185 ( \35529 , \35525 , \35528 );
and \U$35186 ( \35530 , \35523 , \35528 );
or \U$35187 ( \35531 , \35526 , \35529 , \35530 );
xor \U$35188 ( \35532 , \35261 , \35263 );
xor \U$35189 ( \35533 , \35532 , \35266 );
and \U$35190 ( \35534 , \35531 , \35533 );
and \U$35191 ( \35535 , \35275 , \35534 );
xor \U$35192 ( \35536 , \35275 , \35534 );
xor \U$35193 ( \35537 , \35531 , \35533 );
and \U$35194 ( \35538 , \24836 , \25631 );
and \U$35195 ( \35539 , \24714 , \25629 );
nor \U$35196 ( \35540 , \35538 , \35539 );
xnor \U$35197 ( \35541 , \35540 , \25399 );
and \U$35198 ( \35542 , \25097 , \25180 );
and \U$35199 ( \35543 , \24841 , \25178 );
nor \U$35200 ( \35544 , \35542 , \35543 );
xnor \U$35201 ( \35545 , \35544 , \25037 );
and \U$35202 ( \35546 , \35541 , \35545 );
and \U$35203 ( \35547 , \25596 , \24857 );
and \U$35204 ( \35548 , \25294 , \24855 );
nor \U$35205 ( \35549 , \35547 , \35548 );
xnor \U$35206 ( \35550 , \35549 , \24611 );
and \U$35207 ( \35551 , \35545 , \35550 );
and \U$35208 ( \35552 , \35541 , \35550 );
or \U$35209 ( \35553 , \35546 , \35551 , \35552 );
and \U$35210 ( \35554 , \23665 , \27060 );
and \U$35211 ( \35555 , \23491 , \27058 );
nor \U$35212 ( \35556 , \35554 , \35555 );
xnor \U$35213 ( \35557 , \35556 , \26720 );
and \U$35214 ( \35558 , \23970 , \26471 );
and \U$35215 ( \35559 , \23832 , \26469 );
nor \U$35216 ( \35560 , \35558 , \35559 );
xnor \U$35217 ( \35561 , \35560 , \26230 );
and \U$35218 ( \35562 , \35557 , \35561 );
and \U$35219 ( \35563 , \24506 , \26005 );
and \U$35220 ( \35564 , \24089 , \26003 );
nor \U$35221 ( \35565 , \35563 , \35564 );
xnor \U$35222 ( \35566 , \35565 , \25817 );
and \U$35223 ( \35567 , \35561 , \35566 );
and \U$35224 ( \35568 , \35557 , \35566 );
or \U$35225 ( \35569 , \35562 , \35567 , \35568 );
and \U$35226 ( \35570 , \35553 , \35569 );
and \U$35227 ( \35571 , \26073 , \24462 );
and \U$35228 ( \35572 , \25604 , \24460 );
nor \U$35229 ( \35573 , \35571 , \35572 );
xnor \U$35230 ( \35574 , \35573 , \24275 );
and \U$35231 ( \35575 , \26342 , \24149 );
and \U$35232 ( \35576 , \26078 , \24147 );
nor \U$35233 ( \35577 , \35575 , \35576 );
xnor \U$35234 ( \35578 , \35577 , \23944 );
and \U$35235 ( \35579 , \35574 , \35578 );
and \U$35236 ( \35580 , \26973 , \23743 );
and \U$35237 ( \35581 , \26601 , \23741 );
nor \U$35238 ( \35582 , \35580 , \35581 );
xnor \U$35239 ( \35583 , \35582 , \23594 );
and \U$35240 ( \35584 , \35578 , \35583 );
and \U$35241 ( \35585 , \35574 , \35583 );
or \U$35242 ( \35586 , \35579 , \35584 , \35585 );
and \U$35243 ( \35587 , \35569 , \35586 );
and \U$35244 ( \35588 , \35553 , \35586 );
or \U$35245 ( \35589 , \35570 , \35587 , \35588 );
and \U$35246 ( \35590 , \22867 , \28592 );
and \U$35247 ( \35591 , \22624 , \28590 );
nor \U$35248 ( \35592 , \35590 , \35591 );
xnor \U$35249 ( \35593 , \35592 , \28343 );
and \U$35250 ( \35594 , \23058 , \28063 );
and \U$35251 ( \35595 , \22872 , \28061 );
nor \U$35252 ( \35596 , \35594 , \35595 );
xnor \U$35253 ( \35597 , \35596 , \27803 );
and \U$35254 ( \35598 , \35593 , \35597 );
and \U$35255 ( \35599 , \23466 , \27569 );
and \U$35256 ( \35600 , \23202 , \27567 );
nor \U$35257 ( \35601 , \35599 , \35600 );
xnor \U$35258 ( \35602 , \35601 , \27254 );
and \U$35259 ( \35603 , \35597 , \35602 );
and \U$35260 ( \35604 , \35593 , \35602 );
or \U$35261 ( \35605 , \35598 , \35603 , \35604 );
and \U$35262 ( \35606 , \22204 , \30258 );
and \U$35263 ( \35607 , \22099 , \30256 );
nor \U$35264 ( \35608 , \35606 , \35607 );
xnor \U$35265 ( \35609 , \35608 , \29948 );
and \U$35266 ( \35610 , \22325 , \29721 );
and \U$35267 ( \35611 , \22209 , \29719 );
nor \U$35268 ( \35612 , \35610 , \35611 );
xnor \U$35269 ( \35613 , \35612 , \29350 );
and \U$35270 ( \35614 , \35609 , \35613 );
and \U$35271 ( \35615 , \22616 , \29159 );
and \U$35272 ( \35616 , \22440 , \29157 );
nor \U$35273 ( \35617 , \35615 , \35616 );
xnor \U$35274 ( \35618 , \35617 , \28841 );
and \U$35275 ( \35619 , \35613 , \35618 );
and \U$35276 ( \35620 , \35609 , \35618 );
or \U$35277 ( \35621 , \35614 , \35619 , \35620 );
and \U$35278 ( \35622 , \35605 , \35621 );
and \U$35279 ( \35623 , \21750 , \31639 );
and \U$35280 ( \35624 , \21689 , \31636 );
nor \U$35281 ( \35625 , \35623 , \35624 );
xnor \U$35282 ( \35626 , \35625 , \30584 );
and \U$35283 ( \35627 , \22011 , \30826 );
and \U$35284 ( \35628 , \21813 , \30824 );
nor \U$35285 ( \35629 , \35627 , \35628 );
xnor \U$35286 ( \35630 , \35629 , \30587 );
and \U$35287 ( \35631 , \35626 , \35630 );
and \U$35288 ( \35632 , \35630 , \21377 );
and \U$35289 ( \35633 , \35626 , \21377 );
or \U$35290 ( \35634 , \35631 , \35632 , \35633 );
and \U$35291 ( \35635 , \35621 , \35634 );
and \U$35292 ( \35636 , \35605 , \35634 );
or \U$35293 ( \35637 , \35622 , \35635 , \35636 );
and \U$35294 ( \35638 , \35589 , \35637 );
and \U$35295 ( \35639 , \27325 , \23421 );
and \U$35296 ( \35640 , \26982 , \23419 );
nor \U$35297 ( \35641 , \35639 , \35640 );
xnor \U$35298 ( \35642 , \35641 , \23279 );
and \U$35299 ( \35643 , \27830 , \23125 );
and \U$35300 ( \35644 , \27527 , \23123 );
nor \U$35301 ( \35645 , \35643 , \35644 );
xnor \U$35302 ( \35646 , \35645 , \22988 );
and \U$35303 ( \35647 , \35642 , \35646 );
and \U$35304 ( \35648 , \28528 , \22919 );
and \U$35305 ( \35649 , \28002 , \22917 );
nor \U$35306 ( \35650 , \35648 , \35649 );
xnor \U$35307 ( \35651 , \35650 , \22767 );
and \U$35308 ( \35652 , \35646 , \35651 );
and \U$35309 ( \35653 , \35642 , \35651 );
or \U$35310 ( \35654 , \35647 , \35652 , \35653 );
and \U$35311 ( \35655 , \30986 , \21985 );
and \U$35312 ( \35656 , \30383 , \21983 );
nor \U$35313 ( \35657 , \35655 , \35656 );
xnor \U$35314 ( \35658 , \35657 , \21907 );
and \U$35315 ( \35659 , \31172 , \21821 );
and \U$35316 ( \35660 , \30991 , \21819 );
nor \U$35317 ( \35661 , \35659 , \35660 );
xnor \U$35318 ( \35662 , \35661 , \21727 );
and \U$35319 ( \35663 , \35658 , \35662 );
nand \U$35320 ( \35664 , \31792 , \21650 );
xnor \U$35321 ( \35665 , \35664 , \21377 );
and \U$35322 ( \35666 , \35662 , \35665 );
and \U$35323 ( \35667 , \35658 , \35665 );
or \U$35324 ( \35668 , \35663 , \35666 , \35667 );
and \U$35325 ( \35669 , \35654 , \35668 );
and \U$35326 ( \35670 , \29198 , \22651 );
and \U$35327 ( \35671 , \28952 , \22649 );
nor \U$35328 ( \35672 , \35670 , \35671 );
xnor \U$35329 ( \35673 , \35672 , \22495 );
and \U$35330 ( \35674 , \29522 , \22379 );
and \U$35331 ( \35675 , \29203 , \22377 );
nor \U$35332 ( \35676 , \35674 , \35675 );
xnor \U$35333 ( \35677 , \35676 , \22266 );
and \U$35334 ( \35678 , \35673 , \35677 );
and \U$35335 ( \35679 , \30375 , \22185 );
and \U$35336 ( \35680 , \29806 , \22183 );
nor \U$35337 ( \35681 , \35679 , \35680 );
xnor \U$35338 ( \35682 , \35681 , \22049 );
and \U$35339 ( \35683 , \35677 , \35682 );
and \U$35340 ( \35684 , \35673 , \35682 );
or \U$35341 ( \35685 , \35678 , \35683 , \35684 );
and \U$35342 ( \35686 , \35668 , \35685 );
and \U$35343 ( \35687 , \35654 , \35685 );
or \U$35344 ( \35688 , \35669 , \35686 , \35687 );
and \U$35345 ( \35689 , \35637 , \35688 );
and \U$35346 ( \35690 , \35589 , \35688 );
or \U$35347 ( \35691 , \35638 , \35689 , \35690 );
xor \U$35348 ( \35692 , \35377 , \35381 );
xor \U$35349 ( \35693 , \35692 , \35386 );
xor \U$35350 ( \35694 , \35393 , \35397 );
xor \U$35351 ( \35695 , \35694 , \35402 );
and \U$35352 ( \35696 , \35693 , \35695 );
xor \U$35353 ( \35697 , \35410 , \35414 );
xor \U$35354 ( \35698 , \35697 , \35419 );
and \U$35355 ( \35699 , \35695 , \35698 );
and \U$35356 ( \35700 , \35693 , \35698 );
or \U$35357 ( \35701 , \35696 , \35699 , \35700 );
xor \U$35358 ( \35702 , \35279 , \35283 );
xor \U$35359 ( \35703 , \35702 , \35288 );
xor \U$35360 ( \35704 , \35295 , \35299 );
xor \U$35361 ( \35705 , \35704 , \35304 );
and \U$35362 ( \35706 , \35703 , \35705 );
xor \U$35363 ( \35707 , \35312 , \35316 );
xor \U$35364 ( \35708 , \35707 , \35321 );
and \U$35365 ( \35709 , \35705 , \35708 );
and \U$35366 ( \35710 , \35703 , \35708 );
or \U$35367 ( \35711 , \35706 , \35709 , \35710 );
and \U$35368 ( \35712 , \35701 , \35711 );
xor \U$35369 ( \35713 , \35331 , \35335 );
xor \U$35370 ( \35714 , \35713 , \35340 );
xor \U$35371 ( \35715 , \35347 , \35351 );
xor \U$35372 ( \35716 , \35715 , \35356 );
and \U$35373 ( \35717 , \35714 , \35716 );
xor \U$35374 ( \35718 , \35364 , \35368 );
and \U$35375 ( \35719 , \35716 , \35718 );
and \U$35376 ( \35720 , \35714 , \35718 );
or \U$35377 ( \35721 , \35717 , \35719 , \35720 );
and \U$35378 ( \35722 , \35711 , \35721 );
and \U$35379 ( \35723 , \35701 , \35721 );
or \U$35380 ( \35724 , \35712 , \35722 , \35723 );
and \U$35381 ( \35725 , \35691 , \35724 );
xor \U$35382 ( \35726 , \35112 , \35116 );
xor \U$35383 ( \35727 , \35726 , \21392 );
xor \U$35384 ( \35728 , \35430 , \35432 );
xor \U$35385 ( \35729 , \35728 , \35435 );
and \U$35386 ( \35730 , \35727 , \35729 );
xor \U$35387 ( \35731 , \35451 , \35453 );
xor \U$35388 ( \35732 , \35731 , \35456 );
and \U$35389 ( \35733 , \35729 , \35732 );
and \U$35390 ( \35734 , \35727 , \35732 );
or \U$35391 ( \35735 , \35730 , \35733 , \35734 );
and \U$35392 ( \35736 , \35724 , \35735 );
and \U$35393 ( \35737 , \35691 , \35735 );
or \U$35394 ( \35738 , \35725 , \35736 , \35737 );
xor \U$35395 ( \35739 , \35291 , \35307 );
xor \U$35396 ( \35740 , \35739 , \35324 );
xor \U$35397 ( \35741 , \35343 , \35359 );
xor \U$35398 ( \35742 , \35741 , \35369 );
and \U$35399 ( \35743 , \35740 , \35742 );
xor \U$35400 ( \35744 , \35440 , \35442 );
xor \U$35401 ( \35745 , \35744 , \35445 );
and \U$35402 ( \35746 , \35742 , \35745 );
and \U$35403 ( \35747 , \35740 , \35745 );
or \U$35404 ( \35748 , \35743 , \35746 , \35747 );
xor \U$35405 ( \35749 , \35489 , \35491 );
xor \U$35406 ( \35750 , \35749 , \35494 );
and \U$35407 ( \35751 , \35748 , \35750 );
xor \U$35408 ( \35752 , \35465 , \35467 );
xor \U$35409 ( \35753 , \35752 , \35470 );
and \U$35410 ( \35754 , \35750 , \35753 );
and \U$35411 ( \35755 , \35748 , \35753 );
or \U$35412 ( \35756 , \35751 , \35754 , \35755 );
and \U$35413 ( \35757 , \35738 , \35756 );
xor \U$35414 ( \35758 , \35327 , \35372 );
xor \U$35415 ( \35759 , \35758 , \35425 );
xor \U$35416 ( \35760 , \35438 , \35448 );
xor \U$35417 ( \35761 , \35760 , \35459 );
and \U$35418 ( \35762 , \35759 , \35761 );
and \U$35419 ( \35763 , \35756 , \35762 );
and \U$35420 ( \35764 , \35738 , \35762 );
or \U$35421 ( \35765 , \35757 , \35763 , \35764 );
xor \U$35422 ( \35766 , \35428 , \35462 );
xor \U$35423 ( \35767 , \35766 , \35473 );
xor \U$35424 ( \35768 , \35478 , \35480 );
xor \U$35425 ( \35769 , \35768 , \35483 );
and \U$35426 ( \35770 , \35767 , \35769 );
xor \U$35427 ( \35771 , \35497 , \35499 );
xor \U$35428 ( \35772 , \35771 , \35501 );
and \U$35429 ( \35773 , \35769 , \35772 );
and \U$35430 ( \35774 , \35767 , \35772 );
or \U$35431 ( \35775 , \35770 , \35773 , \35774 );
and \U$35432 ( \35776 , \35765 , \35775 );
xor \U$35433 ( \35777 , \35040 , \35196 );
xor \U$35434 ( \35778 , \35777 , \35207 );
and \U$35435 ( \35779 , \35775 , \35778 );
and \U$35436 ( \35780 , \35765 , \35778 );
or \U$35437 ( \35781 , \35776 , \35779 , \35780 );
xor \U$35438 ( \35782 , \35476 , \35486 );
xor \U$35439 ( \35783 , \35782 , \35504 );
xor \U$35440 ( \35784 , \35509 , \35511 );
xor \U$35441 ( \35785 , \35784 , \35514 );
and \U$35442 ( \35786 , \35783 , \35785 );
and \U$35443 ( \35787 , \35781 , \35786 );
xor \U$35444 ( \35788 , \35210 , \35231 );
xor \U$35445 ( \35789 , \35788 , \35242 );
and \U$35446 ( \35790 , \35786 , \35789 );
and \U$35447 ( \35791 , \35781 , \35789 );
or \U$35448 ( \35792 , \35787 , \35790 , \35791 );
xor \U$35449 ( \35793 , \35523 , \35525 );
xor \U$35450 ( \35794 , \35793 , \35528 );
and \U$35451 ( \35795 , \35792 , \35794 );
and \U$35452 ( \35796 , \35537 , \35795 );
xor \U$35453 ( \35797 , \35537 , \35795 );
xor \U$35454 ( \35798 , \35792 , \35794 );
xor \U$35455 ( \35799 , \35781 , \35786 );
xor \U$35456 ( \35800 , \35799 , \35789 );
xor \U$35457 ( \35801 , \35507 , \35517 );
xor \U$35458 ( \35802 , \35801 , \35520 );
and \U$35459 ( \35803 , \35800 , \35802 );
and \U$35460 ( \35804 , \35798 , \35803 );
xor \U$35461 ( \35805 , \35798 , \35803 );
xor \U$35462 ( \35806 , \35800 , \35802 );
and \U$35463 ( \35807 , \23202 , \28063 );
and \U$35464 ( \35808 , \23058 , \28061 );
nor \U$35465 ( \35809 , \35807 , \35808 );
xnor \U$35466 ( \35810 , \35809 , \27803 );
and \U$35467 ( \35811 , \23491 , \27569 );
and \U$35468 ( \35812 , \23466 , \27567 );
nor \U$35469 ( \35813 , \35811 , \35812 );
xnor \U$35470 ( \35814 , \35813 , \27254 );
and \U$35471 ( \35815 , \35810 , \35814 );
and \U$35472 ( \35816 , \23832 , \27060 );
and \U$35473 ( \35817 , \23665 , \27058 );
nor \U$35474 ( \35818 , \35816 , \35817 );
xnor \U$35475 ( \35819 , \35818 , \26720 );
and \U$35476 ( \35820 , \35814 , \35819 );
and \U$35477 ( \35821 , \35810 , \35819 );
or \U$35478 ( \35822 , \35815 , \35820 , \35821 );
and \U$35479 ( \35823 , \21813 , \31639 );
and \U$35480 ( \35824 , \21750 , \31636 );
nor \U$35481 ( \35825 , \35823 , \35824 );
xnor \U$35482 ( \35826 , \35825 , \30584 );
and \U$35483 ( \35827 , \22099 , \30826 );
and \U$35484 ( \35828 , \22011 , \30824 );
nor \U$35485 ( \35829 , \35827 , \35828 );
xnor \U$35486 ( \35830 , \35829 , \30587 );
and \U$35487 ( \35831 , \35826 , \35830 );
and \U$35488 ( \35832 , \22209 , \30258 );
and \U$35489 ( \35833 , \22204 , \30256 );
nor \U$35490 ( \35834 , \35832 , \35833 );
xnor \U$35491 ( \35835 , \35834 , \29948 );
and \U$35492 ( \35836 , \35830 , \35835 );
and \U$35493 ( \35837 , \35826 , \35835 );
or \U$35494 ( \35838 , \35831 , \35836 , \35837 );
and \U$35495 ( \35839 , \35822 , \35838 );
and \U$35496 ( \35840 , \22440 , \29721 );
and \U$35497 ( \35841 , \22325 , \29719 );
nor \U$35498 ( \35842 , \35840 , \35841 );
xnor \U$35499 ( \35843 , \35842 , \29350 );
and \U$35500 ( \35844 , \22624 , \29159 );
and \U$35501 ( \35845 , \22616 , \29157 );
nor \U$35502 ( \35846 , \35844 , \35845 );
xnor \U$35503 ( \35847 , \35846 , \28841 );
and \U$35504 ( \35848 , \35843 , \35847 );
and \U$35505 ( \35849 , \22872 , \28592 );
and \U$35506 ( \35850 , \22867 , \28590 );
nor \U$35507 ( \35851 , \35849 , \35850 );
xnor \U$35508 ( \35852 , \35851 , \28343 );
and \U$35509 ( \35853 , \35847 , \35852 );
and \U$35510 ( \35854 , \35843 , \35852 );
or \U$35511 ( \35855 , \35848 , \35853 , \35854 );
and \U$35512 ( \35856 , \35838 , \35855 );
and \U$35513 ( \35857 , \35822 , \35855 );
or \U$35514 ( \35858 , \35839 , \35856 , \35857 );
and \U$35515 ( \35859 , \25294 , \25180 );
and \U$35516 ( \35860 , \25097 , \25178 );
nor \U$35517 ( \35861 , \35859 , \35860 );
xnor \U$35518 ( \35862 , \35861 , \25037 );
and \U$35519 ( \35863 , \25604 , \24857 );
and \U$35520 ( \35864 , \25596 , \24855 );
nor \U$35521 ( \35865 , \35863 , \35864 );
xnor \U$35522 ( \35866 , \35865 , \24611 );
and \U$35523 ( \35867 , \35862 , \35866 );
and \U$35524 ( \35868 , \26078 , \24462 );
and \U$35525 ( \35869 , \26073 , \24460 );
nor \U$35526 ( \35870 , \35868 , \35869 );
xnor \U$35527 ( \35871 , \35870 , \24275 );
and \U$35528 ( \35872 , \35866 , \35871 );
and \U$35529 ( \35873 , \35862 , \35871 );
or \U$35530 ( \35874 , \35867 , \35872 , \35873 );
and \U$35531 ( \35875 , \24089 , \26471 );
and \U$35532 ( \35876 , \23970 , \26469 );
nor \U$35533 ( \35877 , \35875 , \35876 );
xnor \U$35534 ( \35878 , \35877 , \26230 );
and \U$35535 ( \35879 , \24714 , \26005 );
and \U$35536 ( \35880 , \24506 , \26003 );
nor \U$35537 ( \35881 , \35879 , \35880 );
xnor \U$35538 ( \35882 , \35881 , \25817 );
and \U$35539 ( \35883 , \35878 , \35882 );
and \U$35540 ( \35884 , \24841 , \25631 );
and \U$35541 ( \35885 , \24836 , \25629 );
nor \U$35542 ( \35886 , \35884 , \35885 );
xnor \U$35543 ( \35887 , \35886 , \25399 );
and \U$35544 ( \35888 , \35882 , \35887 );
and \U$35545 ( \35889 , \35878 , \35887 );
or \U$35546 ( \35890 , \35883 , \35888 , \35889 );
and \U$35547 ( \35891 , \35874 , \35890 );
and \U$35548 ( \35892 , \26601 , \24149 );
and \U$35549 ( \35893 , \26342 , \24147 );
nor \U$35550 ( \35894 , \35892 , \35893 );
xnor \U$35551 ( \35895 , \35894 , \23944 );
and \U$35552 ( \35896 , \26982 , \23743 );
and \U$35553 ( \35897 , \26973 , \23741 );
nor \U$35554 ( \35898 , \35896 , \35897 );
xnor \U$35555 ( \35899 , \35898 , \23594 );
and \U$35556 ( \35900 , \35895 , \35899 );
and \U$35557 ( \35901 , \27527 , \23421 );
and \U$35558 ( \35902 , \27325 , \23419 );
nor \U$35559 ( \35903 , \35901 , \35902 );
xnor \U$35560 ( \35904 , \35903 , \23279 );
and \U$35561 ( \35905 , \35899 , \35904 );
and \U$35562 ( \35906 , \35895 , \35904 );
or \U$35563 ( \35907 , \35900 , \35905 , \35906 );
and \U$35564 ( \35908 , \35890 , \35907 );
and \U$35565 ( \35909 , \35874 , \35907 );
or \U$35566 ( \35910 , \35891 , \35908 , \35909 );
and \U$35567 ( \35911 , \35858 , \35910 );
and \U$35568 ( \35912 , \29806 , \22379 );
and \U$35569 ( \35913 , \29522 , \22377 );
nor \U$35570 ( \35914 , \35912 , \35913 );
xnor \U$35571 ( \35915 , \35914 , \22266 );
and \U$35572 ( \35916 , \30383 , \22185 );
and \U$35573 ( \35917 , \30375 , \22183 );
nor \U$35574 ( \35918 , \35916 , \35917 );
xnor \U$35575 ( \35919 , \35918 , \22049 );
and \U$35576 ( \35920 , \35915 , \35919 );
and \U$35577 ( \35921 , \30991 , \21985 );
and \U$35578 ( \35922 , \30986 , \21983 );
nor \U$35579 ( \35923 , \35921 , \35922 );
xnor \U$35580 ( \35924 , \35923 , \21907 );
and \U$35581 ( \35925 , \35919 , \35924 );
and \U$35582 ( \35926 , \35915 , \35924 );
or \U$35583 ( \35927 , \35920 , \35925 , \35926 );
and \U$35584 ( \35928 , \28002 , \23125 );
and \U$35585 ( \35929 , \27830 , \23123 );
nor \U$35586 ( \35930 , \35928 , \35929 );
xnor \U$35587 ( \35931 , \35930 , \22988 );
and \U$35588 ( \35932 , \28952 , \22919 );
and \U$35589 ( \35933 , \28528 , \22917 );
nor \U$35590 ( \35934 , \35932 , \35933 );
xnor \U$35591 ( \35935 , \35934 , \22767 );
and \U$35592 ( \35936 , \35931 , \35935 );
and \U$35593 ( \35937 , \29203 , \22651 );
and \U$35594 ( \35938 , \29198 , \22649 );
nor \U$35595 ( \35939 , \35937 , \35938 );
xnor \U$35596 ( \35940 , \35939 , \22495 );
and \U$35597 ( \35941 , \35935 , \35940 );
and \U$35598 ( \35942 , \35931 , \35940 );
or \U$35599 ( \35943 , \35936 , \35941 , \35942 );
and \U$35600 ( \35944 , \35927 , \35943 );
xor \U$35601 ( \35945 , \35658 , \35662 );
xor \U$35602 ( \35946 , \35945 , \35665 );
and \U$35603 ( \35947 , \35943 , \35946 );
and \U$35604 ( \35948 , \35927 , \35946 );
or \U$35605 ( \35949 , \35944 , \35947 , \35948 );
and \U$35606 ( \35950 , \35910 , \35949 );
and \U$35607 ( \35951 , \35858 , \35949 );
or \U$35608 ( \35952 , \35911 , \35950 , \35951 );
xor \U$35609 ( \35953 , \35642 , \35646 );
xor \U$35610 ( \35954 , \35953 , \35651 );
xor \U$35611 ( \35955 , \35574 , \35578 );
xor \U$35612 ( \35956 , \35955 , \35583 );
and \U$35613 ( \35957 , \35954 , \35956 );
xor \U$35614 ( \35958 , \35673 , \35677 );
xor \U$35615 ( \35959 , \35958 , \35682 );
and \U$35616 ( \35960 , \35956 , \35959 );
and \U$35617 ( \35961 , \35954 , \35959 );
or \U$35618 ( \35962 , \35957 , \35960 , \35961 );
xor \U$35619 ( \35963 , \35541 , \35545 );
xor \U$35620 ( \35964 , \35963 , \35550 );
xor \U$35621 ( \35965 , \35557 , \35561 );
xor \U$35622 ( \35966 , \35965 , \35566 );
and \U$35623 ( \35967 , \35964 , \35966 );
xor \U$35624 ( \35968 , \35593 , \35597 );
xor \U$35625 ( \35969 , \35968 , \35602 );
and \U$35626 ( \35970 , \35966 , \35969 );
and \U$35627 ( \35971 , \35964 , \35969 );
or \U$35628 ( \35972 , \35967 , \35970 , \35971 );
and \U$35629 ( \35973 , \35962 , \35972 );
xor \U$35630 ( \35974 , \35609 , \35613 );
xor \U$35631 ( \35975 , \35974 , \35618 );
xor \U$35632 ( \35976 , \35626 , \35630 );
xor \U$35633 ( \35977 , \35976 , \21377 );
and \U$35634 ( \35978 , \35975 , \35977 );
and \U$35635 ( \35979 , \35972 , \35978 );
and \U$35636 ( \35980 , \35962 , \35978 );
or \U$35637 ( \35981 , \35973 , \35979 , \35980 );
and \U$35638 ( \35982 , \35952 , \35981 );
xor \U$35639 ( \35983 , \35693 , \35695 );
xor \U$35640 ( \35984 , \35983 , \35698 );
xor \U$35641 ( \35985 , \35703 , \35705 );
xor \U$35642 ( \35986 , \35985 , \35708 );
and \U$35643 ( \35987 , \35984 , \35986 );
xor \U$35644 ( \35988 , \35714 , \35716 );
xor \U$35645 ( \35989 , \35988 , \35718 );
and \U$35646 ( \35990 , \35986 , \35989 );
and \U$35647 ( \35991 , \35984 , \35989 );
or \U$35648 ( \35992 , \35987 , \35990 , \35991 );
and \U$35649 ( \35993 , \35981 , \35992 );
and \U$35650 ( \35994 , \35952 , \35992 );
or \U$35651 ( \35995 , \35982 , \35993 , \35994 );
xor \U$35652 ( \35996 , \35553 , \35569 );
xor \U$35653 ( \35997 , \35996 , \35586 );
xor \U$35654 ( \35998 , \35605 , \35621 );
xor \U$35655 ( \35999 , \35998 , \35634 );
and \U$35656 ( \36000 , \35997 , \35999 );
xor \U$35657 ( \36001 , \35654 , \35668 );
xor \U$35658 ( \36002 , \36001 , \35685 );
and \U$35659 ( \36003 , \35999 , \36002 );
and \U$35660 ( \36004 , \35997 , \36002 );
or \U$35661 ( \36005 , \36000 , \36003 , \36004 );
xor \U$35662 ( \36006 , \35389 , \35405 );
xor \U$35663 ( \36007 , \36006 , \35422 );
and \U$35664 ( \36008 , \36005 , \36007 );
xor \U$35665 ( \36009 , \35740 , \35742 );
xor \U$35666 ( \36010 , \36009 , \35745 );
and \U$35667 ( \36011 , \36007 , \36010 );
and \U$35668 ( \36012 , \36005 , \36010 );
or \U$35669 ( \36013 , \36008 , \36011 , \36012 );
and \U$35670 ( \36014 , \35995 , \36013 );
xor \U$35671 ( \36015 , \35589 , \35637 );
xor \U$35672 ( \36016 , \36015 , \35688 );
xor \U$35673 ( \36017 , \35701 , \35711 );
xor \U$35674 ( \36018 , \36017 , \35721 );
and \U$35675 ( \36019 , \36016 , \36018 );
xor \U$35676 ( \36020 , \35727 , \35729 );
xor \U$35677 ( \36021 , \36020 , \35732 );
and \U$35678 ( \36022 , \36018 , \36021 );
and \U$35679 ( \36023 , \36016 , \36021 );
or \U$35680 ( \36024 , \36019 , \36022 , \36023 );
and \U$35681 ( \36025 , \36013 , \36024 );
and \U$35682 ( \36026 , \35995 , \36024 );
or \U$35683 ( \36027 , \36014 , \36025 , \36026 );
xor \U$35684 ( \36028 , \35691 , \35724 );
xor \U$35685 ( \36029 , \36028 , \35735 );
xor \U$35686 ( \36030 , \35748 , \35750 );
xor \U$35687 ( \36031 , \36030 , \35753 );
and \U$35688 ( \36032 , \36029 , \36031 );
xor \U$35689 ( \36033 , \35759 , \35761 );
and \U$35690 ( \36034 , \36031 , \36033 );
and \U$35691 ( \36035 , \36029 , \36033 );
or \U$35692 ( \36036 , \36032 , \36034 , \36035 );
and \U$35693 ( \36037 , \36027 , \36036 );
xor \U$35694 ( \36038 , \35767 , \35769 );
xor \U$35695 ( \36039 , \36038 , \35772 );
and \U$35696 ( \36040 , \36036 , \36039 );
and \U$35697 ( \36041 , \36027 , \36039 );
or \U$35698 ( \36042 , \36037 , \36040 , \36041 );
xor \U$35699 ( \36043 , \35765 , \35775 );
xor \U$35700 ( \36044 , \36043 , \35778 );
and \U$35701 ( \36045 , \36042 , \36044 );
xor \U$35702 ( \36046 , \35783 , \35785 );
and \U$35703 ( \36047 , \36044 , \36046 );
and \U$35704 ( \36048 , \36042 , \36046 );
or \U$35705 ( \36049 , \36045 , \36047 , \36048 );
and \U$35706 ( \36050 , \35806 , \36049 );
xor \U$35707 ( \36051 , \35806 , \36049 );
xor \U$35708 ( \36052 , \36042 , \36044 );
xor \U$35709 ( \36053 , \36052 , \36046 );
and \U$35710 ( \36054 , \23058 , \28592 );
and \U$35711 ( \36055 , \22872 , \28590 );
nor \U$35712 ( \36056 , \36054 , \36055 );
xnor \U$35713 ( \36057 , \36056 , \28343 );
and \U$35714 ( \36058 , \23466 , \28063 );
and \U$35715 ( \36059 , \23202 , \28061 );
nor \U$35716 ( \36060 , \36058 , \36059 );
xnor \U$35717 ( \36061 , \36060 , \27803 );
and \U$35718 ( \36062 , \36057 , \36061 );
and \U$35719 ( \36063 , \23665 , \27569 );
and \U$35720 ( \36064 , \23491 , \27567 );
nor \U$35721 ( \36065 , \36063 , \36064 );
xnor \U$35722 ( \36066 , \36065 , \27254 );
and \U$35723 ( \36067 , \36061 , \36066 );
and \U$35724 ( \36068 , \36057 , \36066 );
or \U$35725 ( \36069 , \36062 , \36067 , \36068 );
and \U$35726 ( \36070 , \22325 , \30258 );
and \U$35727 ( \36071 , \22209 , \30256 );
nor \U$35728 ( \36072 , \36070 , \36071 );
xnor \U$35729 ( \36073 , \36072 , \29948 );
and \U$35730 ( \36074 , \22616 , \29721 );
and \U$35731 ( \36075 , \22440 , \29719 );
nor \U$35732 ( \36076 , \36074 , \36075 );
xnor \U$35733 ( \36077 , \36076 , \29350 );
and \U$35734 ( \36078 , \36073 , \36077 );
and \U$35735 ( \36079 , \22867 , \29159 );
and \U$35736 ( \36080 , \22624 , \29157 );
nor \U$35737 ( \36081 , \36079 , \36080 );
xnor \U$35738 ( \36082 , \36081 , \28841 );
and \U$35739 ( \36083 , \36077 , \36082 );
and \U$35740 ( \36084 , \36073 , \36082 );
or \U$35741 ( \36085 , \36078 , \36083 , \36084 );
and \U$35742 ( \36086 , \36069 , \36085 );
and \U$35743 ( \36087 , \22011 , \31639 );
and \U$35744 ( \36088 , \21813 , \31636 );
nor \U$35745 ( \36089 , \36087 , \36088 );
xnor \U$35746 ( \36090 , \36089 , \30584 );
and \U$35747 ( \36091 , \22204 , \30826 );
and \U$35748 ( \36092 , \22099 , \30824 );
nor \U$35749 ( \36093 , \36091 , \36092 );
xnor \U$35750 ( \36094 , \36093 , \30587 );
and \U$35751 ( \36095 , \36090 , \36094 );
and \U$35752 ( \36096 , \36094 , \21727 );
and \U$35753 ( \36097 , \36090 , \21727 );
or \U$35754 ( \36098 , \36095 , \36096 , \36097 );
and \U$35755 ( \36099 , \36085 , \36098 );
and \U$35756 ( \36100 , \36069 , \36098 );
or \U$35757 ( \36101 , \36086 , \36099 , \36100 );
and \U$35758 ( \36102 , \27830 , \23421 );
and \U$35759 ( \36103 , \27527 , \23419 );
nor \U$35760 ( \36104 , \36102 , \36103 );
xnor \U$35761 ( \36105 , \36104 , \23279 );
and \U$35762 ( \36106 , \28528 , \23125 );
and \U$35763 ( \36107 , \28002 , \23123 );
nor \U$35764 ( \36108 , \36106 , \36107 );
xnor \U$35765 ( \36109 , \36108 , \22988 );
and \U$35766 ( \36110 , \36105 , \36109 );
and \U$35767 ( \36111 , \29198 , \22919 );
and \U$35768 ( \36112 , \28952 , \22917 );
nor \U$35769 ( \36113 , \36111 , \36112 );
xnor \U$35770 ( \36114 , \36113 , \22767 );
and \U$35771 ( \36115 , \36109 , \36114 );
and \U$35772 ( \36116 , \36105 , \36114 );
or \U$35773 ( \36117 , \36110 , \36115 , \36116 );
and \U$35774 ( \36118 , \29522 , \22651 );
and \U$35775 ( \36119 , \29203 , \22649 );
nor \U$35776 ( \36120 , \36118 , \36119 );
xnor \U$35777 ( \36121 , \36120 , \22495 );
and \U$35778 ( \36122 , \30375 , \22379 );
and \U$35779 ( \36123 , \29806 , \22377 );
nor \U$35780 ( \36124 , \36122 , \36123 );
xnor \U$35781 ( \36125 , \36124 , \22266 );
and \U$35782 ( \36126 , \36121 , \36125 );
and \U$35783 ( \36127 , \30986 , \22185 );
and \U$35784 ( \36128 , \30383 , \22183 );
nor \U$35785 ( \36129 , \36127 , \36128 );
xnor \U$35786 ( \36130 , \36129 , \22049 );
and \U$35787 ( \36131 , \36125 , \36130 );
and \U$35788 ( \36132 , \36121 , \36130 );
or \U$35789 ( \36133 , \36126 , \36131 , \36132 );
and \U$35790 ( \36134 , \36117 , \36133 );
and \U$35791 ( \36135 , \31792 , \21821 );
and \U$35792 ( \36136 , \31172 , \21819 );
nor \U$35793 ( \36137 , \36135 , \36136 );
xnor \U$35794 ( \36138 , \36137 , \21727 );
and \U$35795 ( \36139 , \36133 , \36138 );
and \U$35796 ( \36140 , \36117 , \36138 );
or \U$35797 ( \36141 , \36134 , \36139 , \36140 );
and \U$35798 ( \36142 , \36101 , \36141 );
and \U$35799 ( \36143 , \25097 , \25631 );
and \U$35800 ( \36144 , \24841 , \25629 );
nor \U$35801 ( \36145 , \36143 , \36144 );
xnor \U$35802 ( \36146 , \36145 , \25399 );
and \U$35803 ( \36147 , \25596 , \25180 );
and \U$35804 ( \36148 , \25294 , \25178 );
nor \U$35805 ( \36149 , \36147 , \36148 );
xnor \U$35806 ( \36150 , \36149 , \25037 );
and \U$35807 ( \36151 , \36146 , \36150 );
and \U$35808 ( \36152 , \26073 , \24857 );
and \U$35809 ( \36153 , \25604 , \24855 );
nor \U$35810 ( \36154 , \36152 , \36153 );
xnor \U$35811 ( \36155 , \36154 , \24611 );
and \U$35812 ( \36156 , \36150 , \36155 );
and \U$35813 ( \36157 , \36146 , \36155 );
or \U$35814 ( \36158 , \36151 , \36156 , \36157 );
and \U$35815 ( \36159 , \23970 , \27060 );
and \U$35816 ( \36160 , \23832 , \27058 );
nor \U$35817 ( \36161 , \36159 , \36160 );
xnor \U$35818 ( \36162 , \36161 , \26720 );
and \U$35819 ( \36163 , \24506 , \26471 );
and \U$35820 ( \36164 , \24089 , \26469 );
nor \U$35821 ( \36165 , \36163 , \36164 );
xnor \U$35822 ( \36166 , \36165 , \26230 );
and \U$35823 ( \36167 , \36162 , \36166 );
and \U$35824 ( \36168 , \24836 , \26005 );
and \U$35825 ( \36169 , \24714 , \26003 );
nor \U$35826 ( \36170 , \36168 , \36169 );
xnor \U$35827 ( \36171 , \36170 , \25817 );
and \U$35828 ( \36172 , \36166 , \36171 );
and \U$35829 ( \36173 , \36162 , \36171 );
or \U$35830 ( \36174 , \36167 , \36172 , \36173 );
and \U$35831 ( \36175 , \36158 , \36174 );
and \U$35832 ( \36176 , \26342 , \24462 );
and \U$35833 ( \36177 , \26078 , \24460 );
nor \U$35834 ( \36178 , \36176 , \36177 );
xnor \U$35835 ( \36179 , \36178 , \24275 );
and \U$35836 ( \36180 , \26973 , \24149 );
and \U$35837 ( \36181 , \26601 , \24147 );
nor \U$35838 ( \36182 , \36180 , \36181 );
xnor \U$35839 ( \36183 , \36182 , \23944 );
and \U$35840 ( \36184 , \36179 , \36183 );
and \U$35841 ( \36185 , \27325 , \23743 );
and \U$35842 ( \36186 , \26982 , \23741 );
nor \U$35843 ( \36187 , \36185 , \36186 );
xnor \U$35844 ( \36188 , \36187 , \23594 );
and \U$35845 ( \36189 , \36183 , \36188 );
and \U$35846 ( \36190 , \36179 , \36188 );
or \U$35847 ( \36191 , \36184 , \36189 , \36190 );
and \U$35848 ( \36192 , \36174 , \36191 );
and \U$35849 ( \36193 , \36158 , \36191 );
or \U$35850 ( \36194 , \36175 , \36192 , \36193 );
and \U$35851 ( \36195 , \36141 , \36194 );
and \U$35852 ( \36196 , \36101 , \36194 );
or \U$35853 ( \36197 , \36142 , \36195 , \36196 );
xor \U$35854 ( \36198 , \35915 , \35919 );
xor \U$35855 ( \36199 , \36198 , \35924 );
xor \U$35856 ( \36200 , \35895 , \35899 );
xor \U$35857 ( \36201 , \36200 , \35904 );
and \U$35858 ( \36202 , \36199 , \36201 );
xor \U$35859 ( \36203 , \35931 , \35935 );
xor \U$35860 ( \36204 , \36203 , \35940 );
and \U$35861 ( \36205 , \36201 , \36204 );
and \U$35862 ( \36206 , \36199 , \36204 );
or \U$35863 ( \36207 , \36202 , \36205 , \36206 );
xor \U$35864 ( \36208 , \35862 , \35866 );
xor \U$35865 ( \36209 , \36208 , \35871 );
xor \U$35866 ( \36210 , \35878 , \35882 );
xor \U$35867 ( \36211 , \36210 , \35887 );
and \U$35868 ( \36212 , \36209 , \36211 );
xor \U$35869 ( \36213 , \35810 , \35814 );
xor \U$35870 ( \36214 , \36213 , \35819 );
and \U$35871 ( \36215 , \36211 , \36214 );
and \U$35872 ( \36216 , \36209 , \36214 );
or \U$35873 ( \36217 , \36212 , \36215 , \36216 );
and \U$35874 ( \36218 , \36207 , \36217 );
xor \U$35875 ( \36219 , \35826 , \35830 );
xor \U$35876 ( \36220 , \36219 , \35835 );
xor \U$35877 ( \36221 , \35843 , \35847 );
xor \U$35878 ( \36222 , \36221 , \35852 );
and \U$35879 ( \36223 , \36220 , \36222 );
and \U$35880 ( \36224 , \36217 , \36223 );
and \U$35881 ( \36225 , \36207 , \36223 );
or \U$35882 ( \36226 , \36218 , \36224 , \36225 );
and \U$35883 ( \36227 , \36197 , \36226 );
xor \U$35884 ( \36228 , \35954 , \35956 );
xor \U$35885 ( \36229 , \36228 , \35959 );
xor \U$35886 ( \36230 , \35964 , \35966 );
xor \U$35887 ( \36231 , \36230 , \35969 );
and \U$35888 ( \36232 , \36229 , \36231 );
xor \U$35889 ( \36233 , \35975 , \35977 );
and \U$35890 ( \36234 , \36231 , \36233 );
and \U$35891 ( \36235 , \36229 , \36233 );
or \U$35892 ( \36236 , \36232 , \36234 , \36235 );
and \U$35893 ( \36237 , \36226 , \36236 );
and \U$35894 ( \36238 , \36197 , \36236 );
or \U$35895 ( \36239 , \36227 , \36237 , \36238 );
xor \U$35896 ( \36240 , \35822 , \35838 );
xor \U$35897 ( \36241 , \36240 , \35855 );
xor \U$35898 ( \36242 , \35874 , \35890 );
xor \U$35899 ( \36243 , \36242 , \35907 );
and \U$35900 ( \36244 , \36241 , \36243 );
xor \U$35901 ( \36245 , \35927 , \35943 );
xor \U$35902 ( \36246 , \36245 , \35946 );
and \U$35903 ( \36247 , \36243 , \36246 );
and \U$35904 ( \36248 , \36241 , \36246 );
or \U$35905 ( \36249 , \36244 , \36247 , \36248 );
xor \U$35906 ( \36250 , \35997 , \35999 );
xor \U$35907 ( \36251 , \36250 , \36002 );
and \U$35908 ( \36252 , \36249 , \36251 );
xor \U$35909 ( \36253 , \35984 , \35986 );
xor \U$35910 ( \36254 , \36253 , \35989 );
and \U$35911 ( \36255 , \36251 , \36254 );
and \U$35912 ( \36256 , \36249 , \36254 );
or \U$35913 ( \36257 , \36252 , \36255 , \36256 );
and \U$35914 ( \36258 , \36239 , \36257 );
xor \U$35915 ( \36259 , \36016 , \36018 );
xor \U$35916 ( \36260 , \36259 , \36021 );
and \U$35917 ( \36261 , \36257 , \36260 );
and \U$35918 ( \36262 , \36239 , \36260 );
or \U$35919 ( \36263 , \36258 , \36261 , \36262 );
xor \U$35920 ( \36264 , \35995 , \36013 );
xor \U$35921 ( \36265 , \36264 , \36024 );
and \U$35922 ( \36266 , \36263 , \36265 );
xor \U$35923 ( \36267 , \36029 , \36031 );
xor \U$35924 ( \36268 , \36267 , \36033 );
and \U$35925 ( \36269 , \36265 , \36268 );
and \U$35926 ( \36270 , \36263 , \36268 );
or \U$35927 ( \36271 , \36266 , \36269 , \36270 );
xor \U$35928 ( \36272 , \35738 , \35756 );
xor \U$35929 ( \36273 , \36272 , \35762 );
and \U$35930 ( \36274 , \36271 , \36273 );
xor \U$35931 ( \36275 , \36027 , \36036 );
xor \U$35932 ( \36276 , \36275 , \36039 );
and \U$35933 ( \36277 , \36273 , \36276 );
and \U$35934 ( \36278 , \36271 , \36276 );
or \U$35935 ( \36279 , \36274 , \36277 , \36278 );
and \U$35936 ( \36280 , \36053 , \36279 );
xor \U$35937 ( \36281 , \36053 , \36279 );
xor \U$35938 ( \36282 , \36271 , \36273 );
xor \U$35939 ( \36283 , \36282 , \36276 );
xor \U$35940 ( \36284 , \36057 , \36061 );
xor \U$35941 ( \36285 , \36284 , \36066 );
xor \U$35942 ( \36286 , \36073 , \36077 );
xor \U$35943 ( \36287 , \36286 , \36082 );
and \U$35944 ( \36288 , \36285 , \36287 );
xor \U$35945 ( \36289 , \36090 , \36094 );
xor \U$35946 ( \36290 , \36289 , \21727 );
and \U$35947 ( \36291 , \36287 , \36290 );
and \U$35948 ( \36292 , \36285 , \36290 );
or \U$35949 ( \36293 , \36288 , \36291 , \36292 );
nand \U$35950 ( \36294 , \31792 , \21819 );
xnor \U$35951 ( \36295 , \36294 , \21727 );
xor \U$35952 ( \36296 , \36105 , \36109 );
xor \U$35953 ( \36297 , \36296 , \36114 );
and \U$35954 ( \36298 , \36295 , \36297 );
xor \U$35955 ( \36299 , \36121 , \36125 );
xor \U$35956 ( \36300 , \36299 , \36130 );
and \U$35957 ( \36301 , \36297 , \36300 );
and \U$35958 ( \36302 , \36295 , \36300 );
or \U$35959 ( \36303 , \36298 , \36301 , \36302 );
and \U$35960 ( \36304 , \36293 , \36303 );
xor \U$35961 ( \36305 , \36146 , \36150 );
xor \U$35962 ( \36306 , \36305 , \36155 );
xor \U$35963 ( \36307 , \36162 , \36166 );
xor \U$35964 ( \36308 , \36307 , \36171 );
and \U$35965 ( \36309 , \36306 , \36308 );
xor \U$35966 ( \36310 , \36179 , \36183 );
xor \U$35967 ( \36311 , \36310 , \36188 );
and \U$35968 ( \36312 , \36308 , \36311 );
and \U$35969 ( \36313 , \36306 , \36311 );
or \U$35970 ( \36314 , \36309 , \36312 , \36313 );
and \U$35971 ( \36315 , \36303 , \36314 );
and \U$35972 ( \36316 , \36293 , \36314 );
or \U$35973 ( \36317 , \36304 , \36315 , \36316 );
and \U$35974 ( \36318 , \28952 , \23125 );
and \U$35975 ( \36319 , \28528 , \23123 );
nor \U$35976 ( \36320 , \36318 , \36319 );
xnor \U$35977 ( \36321 , \36320 , \22988 );
and \U$35978 ( \36322 , \29203 , \22919 );
and \U$35979 ( \36323 , \29198 , \22917 );
nor \U$35980 ( \36324 , \36322 , \36323 );
xnor \U$35981 ( \36325 , \36324 , \22767 );
and \U$35982 ( \36326 , \36321 , \36325 );
and \U$35983 ( \36327 , \29806 , \22651 );
and \U$35984 ( \36328 , \29522 , \22649 );
nor \U$35985 ( \36329 , \36327 , \36328 );
xnor \U$35986 ( \36330 , \36329 , \22495 );
and \U$35987 ( \36331 , \36325 , \36330 );
and \U$35988 ( \36332 , \36321 , \36330 );
or \U$35989 ( \36333 , \36326 , \36331 , \36332 );
and \U$35990 ( \36334 , \30383 , \22379 );
and \U$35991 ( \36335 , \30375 , \22377 );
nor \U$35992 ( \36336 , \36334 , \36335 );
xnor \U$35993 ( \36337 , \36336 , \22266 );
and \U$35994 ( \36338 , \30991 , \22185 );
and \U$35995 ( \36339 , \30986 , \22183 );
nor \U$35996 ( \36340 , \36338 , \36339 );
xnor \U$35997 ( \36341 , \36340 , \22049 );
and \U$35998 ( \36342 , \36337 , \36341 );
and \U$35999 ( \36343 , \31792 , \21985 );
and \U$36000 ( \36344 , \31172 , \21983 );
nor \U$36001 ( \36345 , \36343 , \36344 );
xnor \U$36002 ( \36346 , \36345 , \21907 );
and \U$36003 ( \36347 , \36341 , \36346 );
and \U$36004 ( \36348 , \36337 , \36346 );
or \U$36005 ( \36349 , \36342 , \36347 , \36348 );
and \U$36006 ( \36350 , \36333 , \36349 );
and \U$36007 ( \36351 , \31172 , \21985 );
and \U$36008 ( \36352 , \30991 , \21983 );
nor \U$36009 ( \36353 , \36351 , \36352 );
xnor \U$36010 ( \36354 , \36353 , \21907 );
and \U$36011 ( \36355 , \36349 , \36354 );
and \U$36012 ( \36356 , \36333 , \36354 );
or \U$36013 ( \36357 , \36350 , \36355 , \36356 );
and \U$36014 ( \36358 , \22099 , \31639 );
and \U$36015 ( \36359 , \22011 , \31636 );
nor \U$36016 ( \36360 , \36358 , \36359 );
xnor \U$36017 ( \36361 , \36360 , \30584 );
and \U$36018 ( \36362 , \22209 , \30826 );
and \U$36019 ( \36363 , \22204 , \30824 );
nor \U$36020 ( \36364 , \36362 , \36363 );
xnor \U$36021 ( \36365 , \36364 , \30587 );
and \U$36022 ( \36366 , \36361 , \36365 );
and \U$36023 ( \36367 , \22440 , \30258 );
and \U$36024 ( \36368 , \22325 , \30256 );
nor \U$36025 ( \36369 , \36367 , \36368 );
xnor \U$36026 ( \36370 , \36369 , \29948 );
and \U$36027 ( \36371 , \36365 , \36370 );
and \U$36028 ( \36372 , \36361 , \36370 );
or \U$36029 ( \36373 , \36366 , \36371 , \36372 );
and \U$36030 ( \36374 , \22624 , \29721 );
and \U$36031 ( \36375 , \22616 , \29719 );
nor \U$36032 ( \36376 , \36374 , \36375 );
xnor \U$36033 ( \36377 , \36376 , \29350 );
and \U$36034 ( \36378 , \22872 , \29159 );
and \U$36035 ( \36379 , \22867 , \29157 );
nor \U$36036 ( \36380 , \36378 , \36379 );
xnor \U$36037 ( \36381 , \36380 , \28841 );
and \U$36038 ( \36382 , \36377 , \36381 );
and \U$36039 ( \36383 , \23202 , \28592 );
and \U$36040 ( \36384 , \23058 , \28590 );
nor \U$36041 ( \36385 , \36383 , \36384 );
xnor \U$36042 ( \36386 , \36385 , \28343 );
and \U$36043 ( \36387 , \36381 , \36386 );
and \U$36044 ( \36388 , \36377 , \36386 );
or \U$36045 ( \36389 , \36382 , \36387 , \36388 );
and \U$36046 ( \36390 , \36373 , \36389 );
and \U$36047 ( \36391 , \23491 , \28063 );
and \U$36048 ( \36392 , \23466 , \28061 );
nor \U$36049 ( \36393 , \36391 , \36392 );
xnor \U$36050 ( \36394 , \36393 , \27803 );
and \U$36051 ( \36395 , \23832 , \27569 );
and \U$36052 ( \36396 , \23665 , \27567 );
nor \U$36053 ( \36397 , \36395 , \36396 );
xnor \U$36054 ( \36398 , \36397 , \27254 );
and \U$36055 ( \36399 , \36394 , \36398 );
and \U$36056 ( \36400 , \24089 , \27060 );
and \U$36057 ( \36401 , \23970 , \27058 );
nor \U$36058 ( \36402 , \36400 , \36401 );
xnor \U$36059 ( \36403 , \36402 , \26720 );
and \U$36060 ( \36404 , \36398 , \36403 );
and \U$36061 ( \36405 , \36394 , \36403 );
or \U$36062 ( \36406 , \36399 , \36404 , \36405 );
and \U$36063 ( \36407 , \36389 , \36406 );
and \U$36064 ( \36408 , \36373 , \36406 );
or \U$36065 ( \36409 , \36390 , \36407 , \36408 );
and \U$36066 ( \36410 , \36357 , \36409 );
and \U$36067 ( \36411 , \25604 , \25180 );
and \U$36068 ( \36412 , \25596 , \25178 );
nor \U$36069 ( \36413 , \36411 , \36412 );
xnor \U$36070 ( \36414 , \36413 , \25037 );
and \U$36071 ( \36415 , \26078 , \24857 );
and \U$36072 ( \36416 , \26073 , \24855 );
nor \U$36073 ( \36417 , \36415 , \36416 );
xnor \U$36074 ( \36418 , \36417 , \24611 );
and \U$36075 ( \36419 , \36414 , \36418 );
and \U$36076 ( \36420 , \26601 , \24462 );
and \U$36077 ( \36421 , \26342 , \24460 );
nor \U$36078 ( \36422 , \36420 , \36421 );
xnor \U$36079 ( \36423 , \36422 , \24275 );
and \U$36080 ( \36424 , \36418 , \36423 );
and \U$36081 ( \36425 , \36414 , \36423 );
or \U$36082 ( \36426 , \36419 , \36424 , \36425 );
and \U$36083 ( \36427 , \26982 , \24149 );
and \U$36084 ( \36428 , \26973 , \24147 );
nor \U$36085 ( \36429 , \36427 , \36428 );
xnor \U$36086 ( \36430 , \36429 , \23944 );
and \U$36087 ( \36431 , \27527 , \23743 );
and \U$36088 ( \36432 , \27325 , \23741 );
nor \U$36089 ( \36433 , \36431 , \36432 );
xnor \U$36090 ( \36434 , \36433 , \23594 );
and \U$36091 ( \36435 , \36430 , \36434 );
and \U$36092 ( \36436 , \28002 , \23421 );
and \U$36093 ( \36437 , \27830 , \23419 );
nor \U$36094 ( \36438 , \36436 , \36437 );
xnor \U$36095 ( \36439 , \36438 , \23279 );
and \U$36096 ( \36440 , \36434 , \36439 );
and \U$36097 ( \36441 , \36430 , \36439 );
or \U$36098 ( \36442 , \36435 , \36440 , \36441 );
and \U$36099 ( \36443 , \36426 , \36442 );
and \U$36100 ( \36444 , \24714 , \26471 );
and \U$36101 ( \36445 , \24506 , \26469 );
nor \U$36102 ( \36446 , \36444 , \36445 );
xnor \U$36103 ( \36447 , \36446 , \26230 );
and \U$36104 ( \36448 , \24841 , \26005 );
and \U$36105 ( \36449 , \24836 , \26003 );
nor \U$36106 ( \36450 , \36448 , \36449 );
xnor \U$36107 ( \36451 , \36450 , \25817 );
and \U$36108 ( \36452 , \36447 , \36451 );
and \U$36109 ( \36453 , \25294 , \25631 );
and \U$36110 ( \36454 , \25097 , \25629 );
nor \U$36111 ( \36455 , \36453 , \36454 );
xnor \U$36112 ( \36456 , \36455 , \25399 );
and \U$36113 ( \36457 , \36451 , \36456 );
and \U$36114 ( \36458 , \36447 , \36456 );
or \U$36115 ( \36459 , \36452 , \36457 , \36458 );
and \U$36116 ( \36460 , \36442 , \36459 );
and \U$36117 ( \36461 , \36426 , \36459 );
or \U$36118 ( \36462 , \36443 , \36460 , \36461 );
and \U$36119 ( \36463 , \36409 , \36462 );
and \U$36120 ( \36464 , \36357 , \36462 );
or \U$36121 ( \36465 , \36410 , \36463 , \36464 );
and \U$36122 ( \36466 , \36317 , \36465 );
xor \U$36123 ( \36467 , \36199 , \36201 );
xor \U$36124 ( \36468 , \36467 , \36204 );
xor \U$36125 ( \36469 , \36209 , \36211 );
xor \U$36126 ( \36470 , \36469 , \36214 );
and \U$36127 ( \36471 , \36468 , \36470 );
xor \U$36128 ( \36472 , \36220 , \36222 );
and \U$36129 ( \36473 , \36470 , \36472 );
and \U$36130 ( \36474 , \36468 , \36472 );
or \U$36131 ( \36475 , \36471 , \36473 , \36474 );
and \U$36132 ( \36476 , \36465 , \36475 );
and \U$36133 ( \36477 , \36317 , \36475 );
or \U$36134 ( \36478 , \36466 , \36476 , \36477 );
xor \U$36135 ( \36479 , \36069 , \36085 );
xor \U$36136 ( \36480 , \36479 , \36098 );
xor \U$36137 ( \36481 , \36117 , \36133 );
xor \U$36138 ( \36482 , \36481 , \36138 );
and \U$36139 ( \36483 , \36480 , \36482 );
xor \U$36140 ( \36484 , \36158 , \36174 );
xor \U$36141 ( \36485 , \36484 , \36191 );
and \U$36142 ( \36486 , \36482 , \36485 );
and \U$36143 ( \36487 , \36480 , \36485 );
or \U$36144 ( \36488 , \36483 , \36486 , \36487 );
xor \U$36145 ( \36489 , \36241 , \36243 );
xor \U$36146 ( \36490 , \36489 , \36246 );
and \U$36147 ( \36491 , \36488 , \36490 );
xor \U$36148 ( \36492 , \36229 , \36231 );
xor \U$36149 ( \36493 , \36492 , \36233 );
and \U$36150 ( \36494 , \36490 , \36493 );
and \U$36151 ( \36495 , \36488 , \36493 );
or \U$36152 ( \36496 , \36491 , \36494 , \36495 );
and \U$36153 ( \36497 , \36478 , \36496 );
xor \U$36154 ( \36498 , \35962 , \35972 );
xor \U$36155 ( \36499 , \36498 , \35978 );
and \U$36156 ( \36500 , \36496 , \36499 );
and \U$36157 ( \36501 , \36478 , \36499 );
or \U$36158 ( \36502 , \36497 , \36500 , \36501 );
xor \U$36159 ( \36503 , \35858 , \35910 );
xor \U$36160 ( \36504 , \36503 , \35949 );
xor \U$36161 ( \36505 , \36197 , \36226 );
xor \U$36162 ( \36506 , \36505 , \36236 );
and \U$36163 ( \36507 , \36504 , \36506 );
xor \U$36164 ( \36508 , \36249 , \36251 );
xor \U$36165 ( \36509 , \36508 , \36254 );
and \U$36166 ( \36510 , \36506 , \36509 );
and \U$36167 ( \36511 , \36504 , \36509 );
or \U$36168 ( \36512 , \36507 , \36510 , \36511 );
and \U$36169 ( \36513 , \36502 , \36512 );
xor \U$36170 ( \36514 , \36005 , \36007 );
xor \U$36171 ( \36515 , \36514 , \36010 );
and \U$36172 ( \36516 , \36512 , \36515 );
and \U$36173 ( \36517 , \36502 , \36515 );
or \U$36174 ( \36518 , \36513 , \36516 , \36517 );
xor \U$36175 ( \36519 , \35952 , \35981 );
xor \U$36176 ( \36520 , \36519 , \35992 );
xor \U$36177 ( \36521 , \36239 , \36257 );
xor \U$36178 ( \36522 , \36521 , \36260 );
and \U$36179 ( \36523 , \36520 , \36522 );
and \U$36180 ( \36524 , \36518 , \36523 );
xor \U$36181 ( \36525 , \36263 , \36265 );
xor \U$36182 ( \36526 , \36525 , \36268 );
and \U$36183 ( \36527 , \36523 , \36526 );
and \U$36184 ( \36528 , \36518 , \36526 );
or \U$36185 ( \36529 , \36524 , \36527 , \36528 );
and \U$36186 ( \36530 , \36283 , \36529 );
xor \U$36187 ( \36531 , \36283 , \36529 );
xor \U$36188 ( \36532 , \36518 , \36523 );
xor \U$36189 ( \36533 , \36532 , \36526 );
and \U$36190 ( \36534 , \26973 , \24462 );
and \U$36191 ( \36535 , \26601 , \24460 );
nor \U$36192 ( \36536 , \36534 , \36535 );
xnor \U$36193 ( \36537 , \36536 , \24275 );
and \U$36194 ( \36538 , \27325 , \24149 );
and \U$36195 ( \36539 , \26982 , \24147 );
nor \U$36196 ( \36540 , \36538 , \36539 );
xnor \U$36197 ( \36541 , \36540 , \23944 );
and \U$36198 ( \36542 , \36537 , \36541 );
and \U$36199 ( \36543 , \27830 , \23743 );
and \U$36200 ( \36544 , \27527 , \23741 );
nor \U$36201 ( \36545 , \36543 , \36544 );
xnor \U$36202 ( \36546 , \36545 , \23594 );
and \U$36203 ( \36547 , \36541 , \36546 );
and \U$36204 ( \36548 , \36537 , \36546 );
or \U$36205 ( \36549 , \36542 , \36547 , \36548 );
and \U$36206 ( \36550 , \25596 , \25631 );
and \U$36207 ( \36551 , \25294 , \25629 );
nor \U$36208 ( \36552 , \36550 , \36551 );
xnor \U$36209 ( \36553 , \36552 , \25399 );
and \U$36210 ( \36554 , \26073 , \25180 );
and \U$36211 ( \36555 , \25604 , \25178 );
nor \U$36212 ( \36556 , \36554 , \36555 );
xnor \U$36213 ( \36557 , \36556 , \25037 );
and \U$36214 ( \36558 , \36553 , \36557 );
and \U$36215 ( \36559 , \26342 , \24857 );
and \U$36216 ( \36560 , \26078 , \24855 );
nor \U$36217 ( \36561 , \36559 , \36560 );
xnor \U$36218 ( \36562 , \36561 , \24611 );
and \U$36219 ( \36563 , \36557 , \36562 );
and \U$36220 ( \36564 , \36553 , \36562 );
or \U$36221 ( \36565 , \36558 , \36563 , \36564 );
and \U$36222 ( \36566 , \36549 , \36565 );
and \U$36223 ( \36567 , \24506 , \27060 );
and \U$36224 ( \36568 , \24089 , \27058 );
nor \U$36225 ( \36569 , \36567 , \36568 );
xnor \U$36226 ( \36570 , \36569 , \26720 );
and \U$36227 ( \36571 , \24836 , \26471 );
and \U$36228 ( \36572 , \24714 , \26469 );
nor \U$36229 ( \36573 , \36571 , \36572 );
xnor \U$36230 ( \36574 , \36573 , \26230 );
and \U$36231 ( \36575 , \36570 , \36574 );
and \U$36232 ( \36576 , \25097 , \26005 );
and \U$36233 ( \36577 , \24841 , \26003 );
nor \U$36234 ( \36578 , \36576 , \36577 );
xnor \U$36235 ( \36579 , \36578 , \25817 );
and \U$36236 ( \36580 , \36574 , \36579 );
and \U$36237 ( \36581 , \36570 , \36579 );
or \U$36238 ( \36582 , \36575 , \36580 , \36581 );
and \U$36239 ( \36583 , \36565 , \36582 );
and \U$36240 ( \36584 , \36549 , \36582 );
or \U$36241 ( \36585 , \36566 , \36583 , \36584 );
and \U$36242 ( \36586 , \22616 , \30258 );
and \U$36243 ( \36587 , \22440 , \30256 );
nor \U$36244 ( \36588 , \36586 , \36587 );
xnor \U$36245 ( \36589 , \36588 , \29948 );
and \U$36246 ( \36590 , \22867 , \29721 );
and \U$36247 ( \36591 , \22624 , \29719 );
nor \U$36248 ( \36592 , \36590 , \36591 );
xnor \U$36249 ( \36593 , \36592 , \29350 );
and \U$36250 ( \36594 , \36589 , \36593 );
and \U$36251 ( \36595 , \23058 , \29159 );
and \U$36252 ( \36596 , \22872 , \29157 );
nor \U$36253 ( \36597 , \36595 , \36596 );
xnor \U$36254 ( \36598 , \36597 , \28841 );
and \U$36255 ( \36599 , \36593 , \36598 );
and \U$36256 ( \36600 , \36589 , \36598 );
or \U$36257 ( \36601 , \36594 , \36599 , \36600 );
and \U$36258 ( \36602 , \22204 , \31639 );
and \U$36259 ( \36603 , \22099 , \31636 );
nor \U$36260 ( \36604 , \36602 , \36603 );
xnor \U$36261 ( \36605 , \36604 , \30584 );
and \U$36262 ( \36606 , \22325 , \30826 );
and \U$36263 ( \36607 , \22209 , \30824 );
nor \U$36264 ( \36608 , \36606 , \36607 );
xnor \U$36265 ( \36609 , \36608 , \30587 );
and \U$36266 ( \36610 , \36605 , \36609 );
and \U$36267 ( \36611 , \36609 , \21907 );
and \U$36268 ( \36612 , \36605 , \21907 );
or \U$36269 ( \36613 , \36610 , \36611 , \36612 );
and \U$36270 ( \36614 , \36601 , \36613 );
and \U$36271 ( \36615 , \23466 , \28592 );
and \U$36272 ( \36616 , \23202 , \28590 );
nor \U$36273 ( \36617 , \36615 , \36616 );
xnor \U$36274 ( \36618 , \36617 , \28343 );
and \U$36275 ( \36619 , \23665 , \28063 );
and \U$36276 ( \36620 , \23491 , \28061 );
nor \U$36277 ( \36621 , \36619 , \36620 );
xnor \U$36278 ( \36622 , \36621 , \27803 );
and \U$36279 ( \36623 , \36618 , \36622 );
and \U$36280 ( \36624 , \23970 , \27569 );
and \U$36281 ( \36625 , \23832 , \27567 );
nor \U$36282 ( \36626 , \36624 , \36625 );
xnor \U$36283 ( \36627 , \36626 , \27254 );
and \U$36284 ( \36628 , \36622 , \36627 );
and \U$36285 ( \36629 , \36618 , \36627 );
or \U$36286 ( \36630 , \36623 , \36628 , \36629 );
and \U$36287 ( \36631 , \36613 , \36630 );
and \U$36288 ( \36632 , \36601 , \36630 );
or \U$36289 ( \36633 , \36614 , \36631 , \36632 );
and \U$36290 ( \36634 , \36585 , \36633 );
and \U$36291 ( \36635 , \28528 , \23421 );
and \U$36292 ( \36636 , \28002 , \23419 );
nor \U$36293 ( \36637 , \36635 , \36636 );
xnor \U$36294 ( \36638 , \36637 , \23279 );
and \U$36295 ( \36639 , \29198 , \23125 );
and \U$36296 ( \36640 , \28952 , \23123 );
nor \U$36297 ( \36641 , \36639 , \36640 );
xnor \U$36298 ( \36642 , \36641 , \22988 );
and \U$36299 ( \36643 , \36638 , \36642 );
and \U$36300 ( \36644 , \29522 , \22919 );
and \U$36301 ( \36645 , \29203 , \22917 );
nor \U$36302 ( \36646 , \36644 , \36645 );
xnor \U$36303 ( \36647 , \36646 , \22767 );
and \U$36304 ( \36648 , \36642 , \36647 );
and \U$36305 ( \36649 , \36638 , \36647 );
or \U$36306 ( \36650 , \36643 , \36648 , \36649 );
and \U$36307 ( \36651 , \30375 , \22651 );
and \U$36308 ( \36652 , \29806 , \22649 );
nor \U$36309 ( \36653 , \36651 , \36652 );
xnor \U$36310 ( \36654 , \36653 , \22495 );
and \U$36311 ( \36655 , \30986 , \22379 );
and \U$36312 ( \36656 , \30383 , \22377 );
nor \U$36313 ( \36657 , \36655 , \36656 );
xnor \U$36314 ( \36658 , \36657 , \22266 );
and \U$36315 ( \36659 , \36654 , \36658 );
and \U$36316 ( \36660 , \31172 , \22185 );
and \U$36317 ( \36661 , \30991 , \22183 );
nor \U$36318 ( \36662 , \36660 , \36661 );
xnor \U$36319 ( \36663 , \36662 , \22049 );
and \U$36320 ( \36664 , \36658 , \36663 );
and \U$36321 ( \36665 , \36654 , \36663 );
or \U$36322 ( \36666 , \36659 , \36664 , \36665 );
and \U$36323 ( \36667 , \36650 , \36666 );
xor \U$36324 ( \36668 , \36337 , \36341 );
xor \U$36325 ( \36669 , \36668 , \36346 );
and \U$36326 ( \36670 , \36666 , \36669 );
and \U$36327 ( \36671 , \36650 , \36669 );
or \U$36328 ( \36672 , \36667 , \36670 , \36671 );
and \U$36329 ( \36673 , \36633 , \36672 );
and \U$36330 ( \36674 , \36585 , \36672 );
or \U$36331 ( \36675 , \36634 , \36673 , \36674 );
xor \U$36332 ( \36676 , \36321 , \36325 );
xor \U$36333 ( \36677 , \36676 , \36330 );
xor \U$36334 ( \36678 , \36414 , \36418 );
xor \U$36335 ( \36679 , \36678 , \36423 );
and \U$36336 ( \36680 , \36677 , \36679 );
xor \U$36337 ( \36681 , \36430 , \36434 );
xor \U$36338 ( \36682 , \36681 , \36439 );
and \U$36339 ( \36683 , \36679 , \36682 );
and \U$36340 ( \36684 , \36677 , \36682 );
or \U$36341 ( \36685 , \36680 , \36683 , \36684 );
xor \U$36342 ( \36686 , \36377 , \36381 );
xor \U$36343 ( \36687 , \36686 , \36386 );
xor \U$36344 ( \36688 , \36447 , \36451 );
xor \U$36345 ( \36689 , \36688 , \36456 );
and \U$36346 ( \36690 , \36687 , \36689 );
xor \U$36347 ( \36691 , \36394 , \36398 );
xor \U$36348 ( \36692 , \36691 , \36403 );
and \U$36349 ( \36693 , \36689 , \36692 );
and \U$36350 ( \36694 , \36687 , \36692 );
or \U$36351 ( \36695 , \36690 , \36693 , \36694 );
and \U$36352 ( \36696 , \36685 , \36695 );
xor \U$36353 ( \36697 , \36285 , \36287 );
xor \U$36354 ( \36698 , \36697 , \36290 );
and \U$36355 ( \36699 , \36695 , \36698 );
and \U$36356 ( \36700 , \36685 , \36698 );
or \U$36357 ( \36701 , \36696 , \36699 , \36700 );
and \U$36358 ( \36702 , \36675 , \36701 );
xor \U$36359 ( \36703 , \36333 , \36349 );
xor \U$36360 ( \36704 , \36703 , \36354 );
xor \U$36361 ( \36705 , \36295 , \36297 );
xor \U$36362 ( \36706 , \36705 , \36300 );
and \U$36363 ( \36707 , \36704 , \36706 );
xor \U$36364 ( \36708 , \36306 , \36308 );
xor \U$36365 ( \36709 , \36708 , \36311 );
and \U$36366 ( \36710 , \36706 , \36709 );
and \U$36367 ( \36711 , \36704 , \36709 );
or \U$36368 ( \36712 , \36707 , \36710 , \36711 );
and \U$36369 ( \36713 , \36701 , \36712 );
and \U$36370 ( \36714 , \36675 , \36712 );
or \U$36371 ( \36715 , \36702 , \36713 , \36714 );
xor \U$36372 ( \36716 , \36293 , \36303 );
xor \U$36373 ( \36717 , \36716 , \36314 );
xor \U$36374 ( \36718 , \36480 , \36482 );
xor \U$36375 ( \36719 , \36718 , \36485 );
and \U$36376 ( \36720 , \36717 , \36719 );
xor \U$36377 ( \36721 , \36468 , \36470 );
xor \U$36378 ( \36722 , \36721 , \36472 );
and \U$36379 ( \36723 , \36719 , \36722 );
and \U$36380 ( \36724 , \36717 , \36722 );
or \U$36381 ( \36725 , \36720 , \36723 , \36724 );
and \U$36382 ( \36726 , \36715 , \36725 );
xor \U$36383 ( \36727 , \36207 , \36217 );
xor \U$36384 ( \36728 , \36727 , \36223 );
and \U$36385 ( \36729 , \36725 , \36728 );
and \U$36386 ( \36730 , \36715 , \36728 );
or \U$36387 ( \36731 , \36726 , \36729 , \36730 );
xor \U$36388 ( \36732 , \36101 , \36141 );
xor \U$36389 ( \36733 , \36732 , \36194 );
xor \U$36390 ( \36734 , \36317 , \36465 );
xor \U$36391 ( \36735 , \36734 , \36475 );
and \U$36392 ( \36736 , \36733 , \36735 );
xor \U$36393 ( \36737 , \36488 , \36490 );
xor \U$36394 ( \36738 , \36737 , \36493 );
and \U$36395 ( \36739 , \36735 , \36738 );
and \U$36396 ( \36740 , \36733 , \36738 );
or \U$36397 ( \36741 , \36736 , \36739 , \36740 );
and \U$36398 ( \36742 , \36731 , \36741 );
xor \U$36399 ( \36743 , \36504 , \36506 );
xor \U$36400 ( \36744 , \36743 , \36509 );
and \U$36401 ( \36745 , \36741 , \36744 );
and \U$36402 ( \36746 , \36731 , \36744 );
or \U$36403 ( \36747 , \36742 , \36745 , \36746 );
xor \U$36404 ( \36748 , \36502 , \36512 );
xor \U$36405 ( \36749 , \36748 , \36515 );
and \U$36406 ( \36750 , \36747 , \36749 );
xor \U$36407 ( \36751 , \36520 , \36522 );
and \U$36408 ( \36752 , \36749 , \36751 );
and \U$36409 ( \36753 , \36747 , \36751 );
or \U$36410 ( \36754 , \36750 , \36752 , \36753 );
and \U$36411 ( \36755 , \36533 , \36754 );
xor \U$36412 ( \36756 , \36533 , \36754 );
xor \U$36413 ( \36757 , \36747 , \36749 );
xor \U$36414 ( \36758 , \36757 , \36751 );
and \U$36415 ( \36759 , \24841 , \26471 );
and \U$36416 ( \36760 , \24836 , \26469 );
nor \U$36417 ( \36761 , \36759 , \36760 );
xnor \U$36418 ( \36762 , \36761 , \26230 );
and \U$36419 ( \36763 , \25294 , \26005 );
and \U$36420 ( \36764 , \25097 , \26003 );
nor \U$36421 ( \36765 , \36763 , \36764 );
xnor \U$36422 ( \36766 , \36765 , \25817 );
and \U$36423 ( \36767 , \36762 , \36766 );
and \U$36424 ( \36768 , \25604 , \25631 );
and \U$36425 ( \36769 , \25596 , \25629 );
nor \U$36426 ( \36770 , \36768 , \36769 );
xnor \U$36427 ( \36771 , \36770 , \25399 );
and \U$36428 ( \36772 , \36766 , \36771 );
and \U$36429 ( \36773 , \36762 , \36771 );
or \U$36430 ( \36774 , \36767 , \36772 , \36773 );
and \U$36431 ( \36775 , \26078 , \25180 );
and \U$36432 ( \36776 , \26073 , \25178 );
nor \U$36433 ( \36777 , \36775 , \36776 );
xnor \U$36434 ( \36778 , \36777 , \25037 );
and \U$36435 ( \36779 , \26601 , \24857 );
and \U$36436 ( \36780 , \26342 , \24855 );
nor \U$36437 ( \36781 , \36779 , \36780 );
xnor \U$36438 ( \36782 , \36781 , \24611 );
and \U$36439 ( \36783 , \36778 , \36782 );
and \U$36440 ( \36784 , \26982 , \24462 );
and \U$36441 ( \36785 , \26973 , \24460 );
nor \U$36442 ( \36786 , \36784 , \36785 );
xnor \U$36443 ( \36787 , \36786 , \24275 );
and \U$36444 ( \36788 , \36782 , \36787 );
and \U$36445 ( \36789 , \36778 , \36787 );
or \U$36446 ( \36790 , \36783 , \36788 , \36789 );
and \U$36447 ( \36791 , \36774 , \36790 );
and \U$36448 ( \36792 , \27527 , \24149 );
and \U$36449 ( \36793 , \27325 , \24147 );
nor \U$36450 ( \36794 , \36792 , \36793 );
xnor \U$36451 ( \36795 , \36794 , \23944 );
and \U$36452 ( \36796 , \28002 , \23743 );
and \U$36453 ( \36797 , \27830 , \23741 );
nor \U$36454 ( \36798 , \36796 , \36797 );
xnor \U$36455 ( \36799 , \36798 , \23594 );
and \U$36456 ( \36800 , \36795 , \36799 );
and \U$36457 ( \36801 , \28952 , \23421 );
and \U$36458 ( \36802 , \28528 , \23419 );
nor \U$36459 ( \36803 , \36801 , \36802 );
xnor \U$36460 ( \36804 , \36803 , \23279 );
and \U$36461 ( \36805 , \36799 , \36804 );
and \U$36462 ( \36806 , \36795 , \36804 );
or \U$36463 ( \36807 , \36800 , \36805 , \36806 );
and \U$36464 ( \36808 , \36790 , \36807 );
and \U$36465 ( \36809 , \36774 , \36807 );
or \U$36466 ( \36810 , \36791 , \36808 , \36809 );
and \U$36467 ( \36811 , \22872 , \29721 );
and \U$36468 ( \36812 , \22867 , \29719 );
nor \U$36469 ( \36813 , \36811 , \36812 );
xnor \U$36470 ( \36814 , \36813 , \29350 );
and \U$36471 ( \36815 , \23202 , \29159 );
and \U$36472 ( \36816 , \23058 , \29157 );
nor \U$36473 ( \36817 , \36815 , \36816 );
xnor \U$36474 ( \36818 , \36817 , \28841 );
and \U$36475 ( \36819 , \36814 , \36818 );
and \U$36476 ( \36820 , \23491 , \28592 );
and \U$36477 ( \36821 , \23466 , \28590 );
nor \U$36478 ( \36822 , \36820 , \36821 );
xnor \U$36479 ( \36823 , \36822 , \28343 );
and \U$36480 ( \36824 , \36818 , \36823 );
and \U$36481 ( \36825 , \36814 , \36823 );
or \U$36482 ( \36826 , \36819 , \36824 , \36825 );
and \U$36483 ( \36827 , \23832 , \28063 );
and \U$36484 ( \36828 , \23665 , \28061 );
nor \U$36485 ( \36829 , \36827 , \36828 );
xnor \U$36486 ( \36830 , \36829 , \27803 );
and \U$36487 ( \36831 , \24089 , \27569 );
and \U$36488 ( \36832 , \23970 , \27567 );
nor \U$36489 ( \36833 , \36831 , \36832 );
xnor \U$36490 ( \36834 , \36833 , \27254 );
and \U$36491 ( \36835 , \36830 , \36834 );
and \U$36492 ( \36836 , \24714 , \27060 );
and \U$36493 ( \36837 , \24506 , \27058 );
nor \U$36494 ( \36838 , \36836 , \36837 );
xnor \U$36495 ( \36839 , \36838 , \26720 );
and \U$36496 ( \36840 , \36834 , \36839 );
and \U$36497 ( \36841 , \36830 , \36839 );
or \U$36498 ( \36842 , \36835 , \36840 , \36841 );
and \U$36499 ( \36843 , \36826 , \36842 );
and \U$36500 ( \36844 , \22209 , \31639 );
and \U$36501 ( \36845 , \22204 , \31636 );
nor \U$36502 ( \36846 , \36844 , \36845 );
xnor \U$36503 ( \36847 , \36846 , \30584 );
and \U$36504 ( \36848 , \22440 , \30826 );
and \U$36505 ( \36849 , \22325 , \30824 );
nor \U$36506 ( \36850 , \36848 , \36849 );
xnor \U$36507 ( \36851 , \36850 , \30587 );
and \U$36508 ( \36852 , \36847 , \36851 );
and \U$36509 ( \36853 , \22624 , \30258 );
and \U$36510 ( \36854 , \22616 , \30256 );
nor \U$36511 ( \36855 , \36853 , \36854 );
xnor \U$36512 ( \36856 , \36855 , \29948 );
and \U$36513 ( \36857 , \36851 , \36856 );
and \U$36514 ( \36858 , \36847 , \36856 );
or \U$36515 ( \36859 , \36852 , \36857 , \36858 );
and \U$36516 ( \36860 , \36842 , \36859 );
and \U$36517 ( \36861 , \36826 , \36859 );
or \U$36518 ( \36862 , \36843 , \36860 , \36861 );
and \U$36519 ( \36863 , \36810 , \36862 );
and \U$36520 ( \36864 , \29203 , \23125 );
and \U$36521 ( \36865 , \29198 , \23123 );
nor \U$36522 ( \36866 , \36864 , \36865 );
xnor \U$36523 ( \36867 , \36866 , \22988 );
and \U$36524 ( \36868 , \29806 , \22919 );
and \U$36525 ( \36869 , \29522 , \22917 );
nor \U$36526 ( \36870 , \36868 , \36869 );
xnor \U$36527 ( \36871 , \36870 , \22767 );
and \U$36528 ( \36872 , \36867 , \36871 );
and \U$36529 ( \36873 , \30383 , \22651 );
and \U$36530 ( \36874 , \30375 , \22649 );
nor \U$36531 ( \36875 , \36873 , \36874 );
xnor \U$36532 ( \36876 , \36875 , \22495 );
and \U$36533 ( \36877 , \36871 , \36876 );
and \U$36534 ( \36878 , \36867 , \36876 );
or \U$36535 ( \36879 , \36872 , \36877 , \36878 );
nand \U$36536 ( \36880 , \31792 , \21983 );
xnor \U$36537 ( \36881 , \36880 , \21907 );
and \U$36538 ( \36882 , \36879 , \36881 );
xor \U$36539 ( \36883 , \36654 , \36658 );
xor \U$36540 ( \36884 , \36883 , \36663 );
and \U$36541 ( \36885 , \36881 , \36884 );
and \U$36542 ( \36886 , \36879 , \36884 );
or \U$36543 ( \36887 , \36882 , \36885 , \36886 );
and \U$36544 ( \36888 , \36862 , \36887 );
and \U$36545 ( \36889 , \36810 , \36887 );
or \U$36546 ( \36890 , \36863 , \36888 , \36889 );
xor \U$36547 ( \36891 , \36537 , \36541 );
xor \U$36548 ( \36892 , \36891 , \36546 );
xor \U$36549 ( \36893 , \36638 , \36642 );
xor \U$36550 ( \36894 , \36893 , \36647 );
and \U$36551 ( \36895 , \36892 , \36894 );
xor \U$36552 ( \36896 , \36553 , \36557 );
xor \U$36553 ( \36897 , \36896 , \36562 );
and \U$36554 ( \36898 , \36894 , \36897 );
and \U$36555 ( \36899 , \36892 , \36897 );
or \U$36556 ( \36900 , \36895 , \36898 , \36899 );
xor \U$36557 ( \36901 , \36589 , \36593 );
xor \U$36558 ( \36902 , \36901 , \36598 );
xor \U$36559 ( \36903 , \36570 , \36574 );
xor \U$36560 ( \36904 , \36903 , \36579 );
and \U$36561 ( \36905 , \36902 , \36904 );
xor \U$36562 ( \36906 , \36618 , \36622 );
xor \U$36563 ( \36907 , \36906 , \36627 );
and \U$36564 ( \36908 , \36904 , \36907 );
and \U$36565 ( \36909 , \36902 , \36907 );
or \U$36566 ( \36910 , \36905 , \36908 , \36909 );
and \U$36567 ( \36911 , \36900 , \36910 );
xor \U$36568 ( \36912 , \36361 , \36365 );
xor \U$36569 ( \36913 , \36912 , \36370 );
and \U$36570 ( \36914 , \36910 , \36913 );
and \U$36571 ( \36915 , \36900 , \36913 );
or \U$36572 ( \36916 , \36911 , \36914 , \36915 );
and \U$36573 ( \36917 , \36890 , \36916 );
xor \U$36574 ( \36918 , \36677 , \36679 );
xor \U$36575 ( \36919 , \36918 , \36682 );
xor \U$36576 ( \36920 , \36687 , \36689 );
xor \U$36577 ( \36921 , \36920 , \36692 );
and \U$36578 ( \36922 , \36919 , \36921 );
xor \U$36579 ( \36923 , \36650 , \36666 );
xor \U$36580 ( \36924 , \36923 , \36669 );
and \U$36581 ( \36925 , \36921 , \36924 );
and \U$36582 ( \36926 , \36919 , \36924 );
or \U$36583 ( \36927 , \36922 , \36925 , \36926 );
and \U$36584 ( \36928 , \36916 , \36927 );
and \U$36585 ( \36929 , \36890 , \36927 );
or \U$36586 ( \36930 , \36917 , \36928 , \36929 );
xor \U$36587 ( \36931 , \36373 , \36389 );
xor \U$36588 ( \36932 , \36931 , \36406 );
xor \U$36589 ( \36933 , \36426 , \36442 );
xor \U$36590 ( \36934 , \36933 , \36459 );
and \U$36591 ( \36935 , \36932 , \36934 );
xor \U$36592 ( \36936 , \36704 , \36706 );
xor \U$36593 ( \36937 , \36936 , \36709 );
and \U$36594 ( \36938 , \36934 , \36937 );
and \U$36595 ( \36939 , \36932 , \36937 );
or \U$36596 ( \36940 , \36935 , \36938 , \36939 );
and \U$36597 ( \36941 , \36930 , \36940 );
xor \U$36598 ( \36942 , \36585 , \36633 );
xor \U$36599 ( \36943 , \36942 , \36672 );
xor \U$36600 ( \36944 , \36685 , \36695 );
xor \U$36601 ( \36945 , \36944 , \36698 );
and \U$36602 ( \36946 , \36943 , \36945 );
and \U$36603 ( \36947 , \36940 , \36946 );
and \U$36604 ( \36948 , \36930 , \36946 );
or \U$36605 ( \36949 , \36941 , \36947 , \36948 );
xor \U$36606 ( \36950 , \36357 , \36409 );
xor \U$36607 ( \36951 , \36950 , \36462 );
xor \U$36608 ( \36952 , \36675 , \36701 );
xor \U$36609 ( \36953 , \36952 , \36712 );
and \U$36610 ( \36954 , \36951 , \36953 );
xor \U$36611 ( \36955 , \36717 , \36719 );
xor \U$36612 ( \36956 , \36955 , \36722 );
and \U$36613 ( \36957 , \36953 , \36956 );
and \U$36614 ( \36958 , \36951 , \36956 );
or \U$36615 ( \36959 , \36954 , \36957 , \36958 );
and \U$36616 ( \36960 , \36949 , \36959 );
xor \U$36617 ( \36961 , \36733 , \36735 );
xor \U$36618 ( \36962 , \36961 , \36738 );
and \U$36619 ( \36963 , \36959 , \36962 );
and \U$36620 ( \36964 , \36949 , \36962 );
or \U$36621 ( \36965 , \36960 , \36963 , \36964 );
xor \U$36622 ( \36966 , \36478 , \36496 );
xor \U$36623 ( \36967 , \36966 , \36499 );
and \U$36624 ( \36968 , \36965 , \36967 );
xor \U$36625 ( \36969 , \36731 , \36741 );
xor \U$36626 ( \36970 , \36969 , \36744 );
and \U$36627 ( \36971 , \36967 , \36970 );
and \U$36628 ( \36972 , \36965 , \36970 );
or \U$36629 ( \36973 , \36968 , \36971 , \36972 );
and \U$36630 ( \36974 , \36758 , \36973 );
xor \U$36631 ( \36975 , \36758 , \36973 );
xor \U$36632 ( \36976 , \36965 , \36967 );
xor \U$36633 ( \36977 , \36976 , \36970 );
and \U$36634 ( \36978 , \22325 , \31639 );
and \U$36635 ( \36979 , \22209 , \31636 );
nor \U$36636 ( \36980 , \36978 , \36979 );
xnor \U$36637 ( \36981 , \36980 , \30584 );
and \U$36638 ( \36982 , \22616 , \30826 );
and \U$36639 ( \36983 , \22440 , \30824 );
nor \U$36640 ( \36984 , \36982 , \36983 );
xnor \U$36641 ( \36985 , \36984 , \30587 );
and \U$36642 ( \36986 , \36981 , \36985 );
and \U$36643 ( \36987 , \36985 , \22049 );
and \U$36644 ( \36988 , \36981 , \22049 );
or \U$36645 ( \36989 , \36986 , \36987 , \36988 );
and \U$36646 ( \36990 , \23665 , \28592 );
and \U$36647 ( \36991 , \23491 , \28590 );
nor \U$36648 ( \36992 , \36990 , \36991 );
xnor \U$36649 ( \36993 , \36992 , \28343 );
and \U$36650 ( \36994 , \23970 , \28063 );
and \U$36651 ( \36995 , \23832 , \28061 );
nor \U$36652 ( \36996 , \36994 , \36995 );
xnor \U$36653 ( \36997 , \36996 , \27803 );
and \U$36654 ( \36998 , \36993 , \36997 );
and \U$36655 ( \36999 , \24506 , \27569 );
and \U$36656 ( \37000 , \24089 , \27567 );
nor \U$36657 ( \37001 , \36999 , \37000 );
xnor \U$36658 ( \37002 , \37001 , \27254 );
and \U$36659 ( \37003 , \36997 , \37002 );
and \U$36660 ( \37004 , \36993 , \37002 );
or \U$36661 ( \37005 , \36998 , \37003 , \37004 );
and \U$36662 ( \37006 , \36989 , \37005 );
and \U$36663 ( \37007 , \22867 , \30258 );
and \U$36664 ( \37008 , \22624 , \30256 );
nor \U$36665 ( \37009 , \37007 , \37008 );
xnor \U$36666 ( \37010 , \37009 , \29948 );
and \U$36667 ( \37011 , \23058 , \29721 );
and \U$36668 ( \37012 , \22872 , \29719 );
nor \U$36669 ( \37013 , \37011 , \37012 );
xnor \U$36670 ( \37014 , \37013 , \29350 );
and \U$36671 ( \37015 , \37010 , \37014 );
and \U$36672 ( \37016 , \23466 , \29159 );
and \U$36673 ( \37017 , \23202 , \29157 );
nor \U$36674 ( \37018 , \37016 , \37017 );
xnor \U$36675 ( \37019 , \37018 , \28841 );
and \U$36676 ( \37020 , \37014 , \37019 );
and \U$36677 ( \37021 , \37010 , \37019 );
or \U$36678 ( \37022 , \37015 , \37020 , \37021 );
and \U$36679 ( \37023 , \37005 , \37022 );
and \U$36680 ( \37024 , \36989 , \37022 );
or \U$36681 ( \37025 , \37006 , \37023 , \37024 );
and \U$36682 ( \37026 , \24836 , \27060 );
and \U$36683 ( \37027 , \24714 , \27058 );
nor \U$36684 ( \37028 , \37026 , \37027 );
xnor \U$36685 ( \37029 , \37028 , \26720 );
and \U$36686 ( \37030 , \25097 , \26471 );
and \U$36687 ( \37031 , \24841 , \26469 );
nor \U$36688 ( \37032 , \37030 , \37031 );
xnor \U$36689 ( \37033 , \37032 , \26230 );
and \U$36690 ( \37034 , \37029 , \37033 );
and \U$36691 ( \37035 , \25596 , \26005 );
and \U$36692 ( \37036 , \25294 , \26003 );
nor \U$36693 ( \37037 , \37035 , \37036 );
xnor \U$36694 ( \37038 , \37037 , \25817 );
and \U$36695 ( \37039 , \37033 , \37038 );
and \U$36696 ( \37040 , \37029 , \37038 );
or \U$36697 ( \37041 , \37034 , \37039 , \37040 );
and \U$36698 ( \37042 , \26073 , \25631 );
and \U$36699 ( \37043 , \25604 , \25629 );
nor \U$36700 ( \37044 , \37042 , \37043 );
xnor \U$36701 ( \37045 , \37044 , \25399 );
and \U$36702 ( \37046 , \26342 , \25180 );
and \U$36703 ( \37047 , \26078 , \25178 );
nor \U$36704 ( \37048 , \37046 , \37047 );
xnor \U$36705 ( \37049 , \37048 , \25037 );
and \U$36706 ( \37050 , \37045 , \37049 );
and \U$36707 ( \37051 , \26973 , \24857 );
and \U$36708 ( \37052 , \26601 , \24855 );
nor \U$36709 ( \37053 , \37051 , \37052 );
xnor \U$36710 ( \37054 , \37053 , \24611 );
and \U$36711 ( \37055 , \37049 , \37054 );
and \U$36712 ( \37056 , \37045 , \37054 );
or \U$36713 ( \37057 , \37050 , \37055 , \37056 );
and \U$36714 ( \37058 , \37041 , \37057 );
and \U$36715 ( \37059 , \27325 , \24462 );
and \U$36716 ( \37060 , \26982 , \24460 );
nor \U$36717 ( \37061 , \37059 , \37060 );
xnor \U$36718 ( \37062 , \37061 , \24275 );
and \U$36719 ( \37063 , \27830 , \24149 );
and \U$36720 ( \37064 , \27527 , \24147 );
nor \U$36721 ( \37065 , \37063 , \37064 );
xnor \U$36722 ( \37066 , \37065 , \23944 );
and \U$36723 ( \37067 , \37062 , \37066 );
and \U$36724 ( \37068 , \28528 , \23743 );
and \U$36725 ( \37069 , \28002 , \23741 );
nor \U$36726 ( \37070 , \37068 , \37069 );
xnor \U$36727 ( \37071 , \37070 , \23594 );
and \U$36728 ( \37072 , \37066 , \37071 );
and \U$36729 ( \37073 , \37062 , \37071 );
or \U$36730 ( \37074 , \37067 , \37072 , \37073 );
and \U$36731 ( \37075 , \37057 , \37074 );
and \U$36732 ( \37076 , \37041 , \37074 );
or \U$36733 ( \37077 , \37058 , \37075 , \37076 );
and \U$36734 ( \37078 , \37025 , \37077 );
and \U$36735 ( \37079 , \30986 , \22651 );
and \U$36736 ( \37080 , \30383 , \22649 );
nor \U$36737 ( \37081 , \37079 , \37080 );
xnor \U$36738 ( \37082 , \37081 , \22495 );
and \U$36739 ( \37083 , \31172 , \22379 );
and \U$36740 ( \37084 , \30991 , \22377 );
nor \U$36741 ( \37085 , \37083 , \37084 );
xnor \U$36742 ( \37086 , \37085 , \22266 );
and \U$36743 ( \37087 , \37082 , \37086 );
nand \U$36744 ( \37088 , \31792 , \22183 );
xnor \U$36745 ( \37089 , \37088 , \22049 );
and \U$36746 ( \37090 , \37086 , \37089 );
and \U$36747 ( \37091 , \37082 , \37089 );
or \U$36748 ( \37092 , \37087 , \37090 , \37091 );
and \U$36749 ( \37093 , \29198 , \23421 );
and \U$36750 ( \37094 , \28952 , \23419 );
nor \U$36751 ( \37095 , \37093 , \37094 );
xnor \U$36752 ( \37096 , \37095 , \23279 );
and \U$36753 ( \37097 , \29522 , \23125 );
and \U$36754 ( \37098 , \29203 , \23123 );
nor \U$36755 ( \37099 , \37097 , \37098 );
xnor \U$36756 ( \37100 , \37099 , \22988 );
and \U$36757 ( \37101 , \37096 , \37100 );
and \U$36758 ( \37102 , \30375 , \22919 );
and \U$36759 ( \37103 , \29806 , \22917 );
nor \U$36760 ( \37104 , \37102 , \37103 );
xnor \U$36761 ( \37105 , \37104 , \22767 );
and \U$36762 ( \37106 , \37100 , \37105 );
and \U$36763 ( \37107 , \37096 , \37105 );
or \U$36764 ( \37108 , \37101 , \37106 , \37107 );
and \U$36765 ( \37109 , \37092 , \37108 );
and \U$36766 ( \37110 , \30991 , \22379 );
and \U$36767 ( \37111 , \30986 , \22377 );
nor \U$36768 ( \37112 , \37110 , \37111 );
xnor \U$36769 ( \37113 , \37112 , \22266 );
and \U$36770 ( \37114 , \37108 , \37113 );
and \U$36771 ( \37115 , \37092 , \37113 );
or \U$36772 ( \37116 , \37109 , \37114 , \37115 );
and \U$36773 ( \37117 , \37077 , \37116 );
and \U$36774 ( \37118 , \37025 , \37116 );
or \U$36775 ( \37119 , \37078 , \37117 , \37118 );
and \U$36776 ( \37120 , \31792 , \22185 );
and \U$36777 ( \37121 , \31172 , \22183 );
nor \U$36778 ( \37122 , \37120 , \37121 );
xnor \U$36779 ( \37123 , \37122 , \22049 );
xor \U$36780 ( \37124 , \36795 , \36799 );
xor \U$36781 ( \37125 , \37124 , \36804 );
and \U$36782 ( \37126 , \37123 , \37125 );
xor \U$36783 ( \37127 , \36867 , \36871 );
xor \U$36784 ( \37128 , \37127 , \36876 );
and \U$36785 ( \37129 , \37125 , \37128 );
and \U$36786 ( \37130 , \37123 , \37128 );
or \U$36787 ( \37131 , \37126 , \37129 , \37130 );
xor \U$36788 ( \37132 , \36762 , \36766 );
xor \U$36789 ( \37133 , \37132 , \36771 );
xor \U$36790 ( \37134 , \36778 , \36782 );
xor \U$36791 ( \37135 , \37134 , \36787 );
and \U$36792 ( \37136 , \37133 , \37135 );
xor \U$36793 ( \37137 , \36830 , \36834 );
xor \U$36794 ( \37138 , \37137 , \36839 );
and \U$36795 ( \37139 , \37135 , \37138 );
and \U$36796 ( \37140 , \37133 , \37138 );
or \U$36797 ( \37141 , \37136 , \37139 , \37140 );
and \U$36798 ( \37142 , \37131 , \37141 );
xor \U$36799 ( \37143 , \36605 , \36609 );
xor \U$36800 ( \37144 , \37143 , \21907 );
and \U$36801 ( \37145 , \37141 , \37144 );
and \U$36802 ( \37146 , \37131 , \37144 );
or \U$36803 ( \37147 , \37142 , \37145 , \37146 );
and \U$36804 ( \37148 , \37119 , \37147 );
xor \U$36805 ( \37149 , \36879 , \36881 );
xor \U$36806 ( \37150 , \37149 , \36884 );
xor \U$36807 ( \37151 , \36892 , \36894 );
xor \U$36808 ( \37152 , \37151 , \36897 );
and \U$36809 ( \37153 , \37150 , \37152 );
xor \U$36810 ( \37154 , \36902 , \36904 );
xor \U$36811 ( \37155 , \37154 , \36907 );
and \U$36812 ( \37156 , \37152 , \37155 );
and \U$36813 ( \37157 , \37150 , \37155 );
or \U$36814 ( \37158 , \37153 , \37156 , \37157 );
and \U$36815 ( \37159 , \37147 , \37158 );
and \U$36816 ( \37160 , \37119 , \37158 );
or \U$36817 ( \37161 , \37148 , \37159 , \37160 );
xor \U$36818 ( \37162 , \36549 , \36565 );
xor \U$36819 ( \37163 , \37162 , \36582 );
xor \U$36820 ( \37164 , \36601 , \36613 );
xor \U$36821 ( \37165 , \37164 , \36630 );
and \U$36822 ( \37166 , \37163 , \37165 );
xor \U$36823 ( \37167 , \36919 , \36921 );
xor \U$36824 ( \37168 , \37167 , \36924 );
and \U$36825 ( \37169 , \37165 , \37168 );
and \U$36826 ( \37170 , \37163 , \37168 );
or \U$36827 ( \37171 , \37166 , \37169 , \37170 );
and \U$36828 ( \37172 , \37161 , \37171 );
xor \U$36829 ( \37173 , \36810 , \36862 );
xor \U$36830 ( \37174 , \37173 , \36887 );
xor \U$36831 ( \37175 , \36900 , \36910 );
xor \U$36832 ( \37176 , \37175 , \36913 );
and \U$36833 ( \37177 , \37174 , \37176 );
and \U$36834 ( \37178 , \37171 , \37177 );
and \U$36835 ( \37179 , \37161 , \37177 );
or \U$36836 ( \37180 , \37172 , \37178 , \37179 );
xor \U$36837 ( \37181 , \36890 , \36916 );
xor \U$36838 ( \37182 , \37181 , \36927 );
xor \U$36839 ( \37183 , \36932 , \36934 );
xor \U$36840 ( \37184 , \37183 , \36937 );
and \U$36841 ( \37185 , \37182 , \37184 );
xor \U$36842 ( \37186 , \36943 , \36945 );
and \U$36843 ( \37187 , \37184 , \37186 );
and \U$36844 ( \37188 , \37182 , \37186 );
or \U$36845 ( \37189 , \37185 , \37187 , \37188 );
and \U$36846 ( \37190 , \37180 , \37189 );
xor \U$36847 ( \37191 , \36951 , \36953 );
xor \U$36848 ( \37192 , \37191 , \36956 );
and \U$36849 ( \37193 , \37189 , \37192 );
and \U$36850 ( \37194 , \37180 , \37192 );
or \U$36851 ( \37195 , \37190 , \37193 , \37194 );
xor \U$36852 ( \37196 , \36715 , \36725 );
xor \U$36853 ( \37197 , \37196 , \36728 );
and \U$36854 ( \37198 , \37195 , \37197 );
xor \U$36855 ( \37199 , \36949 , \36959 );
xor \U$36856 ( \37200 , \37199 , \36962 );
and \U$36857 ( \37201 , \37197 , \37200 );
and \U$36858 ( \37202 , \37195 , \37200 );
or \U$36859 ( \37203 , \37198 , \37201 , \37202 );
and \U$36860 ( \37204 , \36977 , \37203 );
xor \U$36861 ( \37205 , \36977 , \37203 );
xor \U$36862 ( \37206 , \37195 , \37197 );
xor \U$36863 ( \37207 , \37206 , \37200 );
and \U$36864 ( \37208 , \22440 , \31639 );
and \U$36865 ( \37209 , \22325 , \31636 );
nor \U$36866 ( \37210 , \37208 , \37209 );
xnor \U$36867 ( \37211 , \37210 , \30584 );
and \U$36868 ( \37212 , \22624 , \30826 );
and \U$36869 ( \37213 , \22616 , \30824 );
nor \U$36870 ( \37214 , \37212 , \37213 );
xnor \U$36871 ( \37215 , \37214 , \30587 );
and \U$36872 ( \37216 , \37211 , \37215 );
and \U$36873 ( \37217 , \22872 , \30258 );
and \U$36874 ( \37218 , \22867 , \30256 );
nor \U$36875 ( \37219 , \37217 , \37218 );
xnor \U$36876 ( \37220 , \37219 , \29948 );
and \U$36877 ( \37221 , \37215 , \37220 );
and \U$36878 ( \37222 , \37211 , \37220 );
or \U$36879 ( \37223 , \37216 , \37221 , \37222 );
and \U$36880 ( \37224 , \23202 , \29721 );
and \U$36881 ( \37225 , \23058 , \29719 );
nor \U$36882 ( \37226 , \37224 , \37225 );
xnor \U$36883 ( \37227 , \37226 , \29350 );
and \U$36884 ( \37228 , \23491 , \29159 );
and \U$36885 ( \37229 , \23466 , \29157 );
nor \U$36886 ( \37230 , \37228 , \37229 );
xnor \U$36887 ( \37231 , \37230 , \28841 );
and \U$36888 ( \37232 , \37227 , \37231 );
and \U$36889 ( \37233 , \23832 , \28592 );
and \U$36890 ( \37234 , \23665 , \28590 );
nor \U$36891 ( \37235 , \37233 , \37234 );
xnor \U$36892 ( \37236 , \37235 , \28343 );
and \U$36893 ( \37237 , \37231 , \37236 );
and \U$36894 ( \37238 , \37227 , \37236 );
or \U$36895 ( \37239 , \37232 , \37237 , \37238 );
and \U$36896 ( \37240 , \37223 , \37239 );
and \U$36897 ( \37241 , \24089 , \28063 );
and \U$36898 ( \37242 , \23970 , \28061 );
nor \U$36899 ( \37243 , \37241 , \37242 );
xnor \U$36900 ( \37244 , \37243 , \27803 );
and \U$36901 ( \37245 , \24714 , \27569 );
and \U$36902 ( \37246 , \24506 , \27567 );
nor \U$36903 ( \37247 , \37245 , \37246 );
xnor \U$36904 ( \37248 , \37247 , \27254 );
and \U$36905 ( \37249 , \37244 , \37248 );
and \U$36906 ( \37250 , \24841 , \27060 );
and \U$36907 ( \37251 , \24836 , \27058 );
nor \U$36908 ( \37252 , \37250 , \37251 );
xnor \U$36909 ( \37253 , \37252 , \26720 );
and \U$36910 ( \37254 , \37248 , \37253 );
and \U$36911 ( \37255 , \37244 , \37253 );
or \U$36912 ( \37256 , \37249 , \37254 , \37255 );
and \U$36913 ( \37257 , \37239 , \37256 );
and \U$36914 ( \37258 , \37223 , \37256 );
or \U$36915 ( \37259 , \37240 , \37257 , \37258 );
and \U$36916 ( \37260 , \26601 , \25180 );
and \U$36917 ( \37261 , \26342 , \25178 );
nor \U$36918 ( \37262 , \37260 , \37261 );
xnor \U$36919 ( \37263 , \37262 , \25037 );
and \U$36920 ( \37264 , \26982 , \24857 );
and \U$36921 ( \37265 , \26973 , \24855 );
nor \U$36922 ( \37266 , \37264 , \37265 );
xnor \U$36923 ( \37267 , \37266 , \24611 );
and \U$36924 ( \37268 , \37263 , \37267 );
and \U$36925 ( \37269 , \27527 , \24462 );
and \U$36926 ( \37270 , \27325 , \24460 );
nor \U$36927 ( \37271 , \37269 , \37270 );
xnor \U$36928 ( \37272 , \37271 , \24275 );
and \U$36929 ( \37273 , \37267 , \37272 );
and \U$36930 ( \37274 , \37263 , \37272 );
or \U$36931 ( \37275 , \37268 , \37273 , \37274 );
and \U$36932 ( \37276 , \28002 , \24149 );
and \U$36933 ( \37277 , \27830 , \24147 );
nor \U$36934 ( \37278 , \37276 , \37277 );
xnor \U$36935 ( \37279 , \37278 , \23944 );
and \U$36936 ( \37280 , \28952 , \23743 );
and \U$36937 ( \37281 , \28528 , \23741 );
nor \U$36938 ( \37282 , \37280 , \37281 );
xnor \U$36939 ( \37283 , \37282 , \23594 );
and \U$36940 ( \37284 , \37279 , \37283 );
and \U$36941 ( \37285 , \29203 , \23421 );
and \U$36942 ( \37286 , \29198 , \23419 );
nor \U$36943 ( \37287 , \37285 , \37286 );
xnor \U$36944 ( \37288 , \37287 , \23279 );
and \U$36945 ( \37289 , \37283 , \37288 );
and \U$36946 ( \37290 , \37279 , \37288 );
or \U$36947 ( \37291 , \37284 , \37289 , \37290 );
and \U$36948 ( \37292 , \37275 , \37291 );
and \U$36949 ( \37293 , \25294 , \26471 );
and \U$36950 ( \37294 , \25097 , \26469 );
nor \U$36951 ( \37295 , \37293 , \37294 );
xnor \U$36952 ( \37296 , \37295 , \26230 );
and \U$36953 ( \37297 , \25604 , \26005 );
and \U$36954 ( \37298 , \25596 , \26003 );
nor \U$36955 ( \37299 , \37297 , \37298 );
xnor \U$36956 ( \37300 , \37299 , \25817 );
and \U$36957 ( \37301 , \37296 , \37300 );
and \U$36958 ( \37302 , \26078 , \25631 );
and \U$36959 ( \37303 , \26073 , \25629 );
nor \U$36960 ( \37304 , \37302 , \37303 );
xnor \U$36961 ( \37305 , \37304 , \25399 );
and \U$36962 ( \37306 , \37300 , \37305 );
and \U$36963 ( \37307 , \37296 , \37305 );
or \U$36964 ( \37308 , \37301 , \37306 , \37307 );
and \U$36965 ( \37309 , \37291 , \37308 );
and \U$36966 ( \37310 , \37275 , \37308 );
or \U$36967 ( \37311 , \37292 , \37309 , \37310 );
and \U$36968 ( \37312 , \37259 , \37311 );
and \U$36969 ( \37313 , \29806 , \23125 );
and \U$36970 ( \37314 , \29522 , \23123 );
nor \U$36971 ( \37315 , \37313 , \37314 );
xnor \U$36972 ( \37316 , \37315 , \22988 );
and \U$36973 ( \37317 , \30383 , \22919 );
and \U$36974 ( \37318 , \30375 , \22917 );
nor \U$36975 ( \37319 , \37317 , \37318 );
xnor \U$36976 ( \37320 , \37319 , \22767 );
and \U$36977 ( \37321 , \37316 , \37320 );
and \U$36978 ( \37322 , \30991 , \22651 );
and \U$36979 ( \37323 , \30986 , \22649 );
nor \U$36980 ( \37324 , \37322 , \37323 );
xnor \U$36981 ( \37325 , \37324 , \22495 );
and \U$36982 ( \37326 , \37320 , \37325 );
and \U$36983 ( \37327 , \37316 , \37325 );
or \U$36984 ( \37328 , \37321 , \37326 , \37327 );
xor \U$36985 ( \37329 , \37082 , \37086 );
xor \U$36986 ( \37330 , \37329 , \37089 );
and \U$36987 ( \37331 , \37328 , \37330 );
xor \U$36988 ( \37332 , \37096 , \37100 );
xor \U$36989 ( \37333 , \37332 , \37105 );
and \U$36990 ( \37334 , \37330 , \37333 );
and \U$36991 ( \37335 , \37328 , \37333 );
or \U$36992 ( \37336 , \37331 , \37334 , \37335 );
and \U$36993 ( \37337 , \37311 , \37336 );
and \U$36994 ( \37338 , \37259 , \37336 );
or \U$36995 ( \37339 , \37312 , \37337 , \37338 );
xor \U$36996 ( \37340 , \37029 , \37033 );
xor \U$36997 ( \37341 , \37340 , \37038 );
xor \U$36998 ( \37342 , \37045 , \37049 );
xor \U$36999 ( \37343 , \37342 , \37054 );
and \U$37000 ( \37344 , \37341 , \37343 );
xor \U$37001 ( \37345 , \37062 , \37066 );
xor \U$37002 ( \37346 , \37345 , \37071 );
and \U$37003 ( \37347 , \37343 , \37346 );
and \U$37004 ( \37348 , \37341 , \37346 );
or \U$37005 ( \37349 , \37344 , \37347 , \37348 );
xor \U$37006 ( \37350 , \36981 , \36985 );
xor \U$37007 ( \37351 , \37350 , \22049 );
xor \U$37008 ( \37352 , \36993 , \36997 );
xor \U$37009 ( \37353 , \37352 , \37002 );
and \U$37010 ( \37354 , \37351 , \37353 );
xor \U$37011 ( \37355 , \37010 , \37014 );
xor \U$37012 ( \37356 , \37355 , \37019 );
and \U$37013 ( \37357 , \37353 , \37356 );
and \U$37014 ( \37358 , \37351 , \37356 );
or \U$37015 ( \37359 , \37354 , \37357 , \37358 );
and \U$37016 ( \37360 , \37349 , \37359 );
xor \U$37017 ( \37361 , \36814 , \36818 );
xor \U$37018 ( \37362 , \37361 , \36823 );
and \U$37019 ( \37363 , \37359 , \37362 );
and \U$37020 ( \37364 , \37349 , \37362 );
or \U$37021 ( \37365 , \37360 , \37363 , \37364 );
and \U$37022 ( \37366 , \37339 , \37365 );
xor \U$37023 ( \37367 , \36847 , \36851 );
xor \U$37024 ( \37368 , \37367 , \36856 );
xor \U$37025 ( \37369 , \37123 , \37125 );
xor \U$37026 ( \37370 , \37369 , \37128 );
and \U$37027 ( \37371 , \37368 , \37370 );
xor \U$37028 ( \37372 , \37133 , \37135 );
xor \U$37029 ( \37373 , \37372 , \37138 );
and \U$37030 ( \37374 , \37370 , \37373 );
and \U$37031 ( \37375 , \37368 , \37373 );
or \U$37032 ( \37376 , \37371 , \37374 , \37375 );
and \U$37033 ( \37377 , \37365 , \37376 );
and \U$37034 ( \37378 , \37339 , \37376 );
or \U$37035 ( \37379 , \37366 , \37377 , \37378 );
xor \U$37036 ( \37380 , \36989 , \37005 );
xor \U$37037 ( \37381 , \37380 , \37022 );
xor \U$37038 ( \37382 , \37041 , \37057 );
xor \U$37039 ( \37383 , \37382 , \37074 );
and \U$37040 ( \37384 , \37381 , \37383 );
xor \U$37041 ( \37385 , \37092 , \37108 );
xor \U$37042 ( \37386 , \37385 , \37113 );
and \U$37043 ( \37387 , \37383 , \37386 );
and \U$37044 ( \37388 , \37381 , \37386 );
or \U$37045 ( \37389 , \37384 , \37387 , \37388 );
xor \U$37046 ( \37390 , \36774 , \36790 );
xor \U$37047 ( \37391 , \37390 , \36807 );
and \U$37048 ( \37392 , \37389 , \37391 );
xor \U$37049 ( \37393 , \36826 , \36842 );
xor \U$37050 ( \37394 , \37393 , \36859 );
and \U$37051 ( \37395 , \37391 , \37394 );
and \U$37052 ( \37396 , \37389 , \37394 );
or \U$37053 ( \37397 , \37392 , \37395 , \37396 );
and \U$37054 ( \37398 , \37379 , \37397 );
xor \U$37055 ( \37399 , \37025 , \37077 );
xor \U$37056 ( \37400 , \37399 , \37116 );
xor \U$37057 ( \37401 , \37131 , \37141 );
xor \U$37058 ( \37402 , \37401 , \37144 );
and \U$37059 ( \37403 , \37400 , \37402 );
xor \U$37060 ( \37404 , \37150 , \37152 );
xor \U$37061 ( \37405 , \37404 , \37155 );
and \U$37062 ( \37406 , \37402 , \37405 );
and \U$37063 ( \37407 , \37400 , \37405 );
or \U$37064 ( \37408 , \37403 , \37406 , \37407 );
and \U$37065 ( \37409 , \37397 , \37408 );
and \U$37066 ( \37410 , \37379 , \37408 );
or \U$37067 ( \37411 , \37398 , \37409 , \37410 );
xor \U$37068 ( \37412 , \37119 , \37147 );
xor \U$37069 ( \37413 , \37412 , \37158 );
xor \U$37070 ( \37414 , \37163 , \37165 );
xor \U$37071 ( \37415 , \37414 , \37168 );
and \U$37072 ( \37416 , \37413 , \37415 );
xor \U$37073 ( \37417 , \37174 , \37176 );
and \U$37074 ( \37418 , \37415 , \37417 );
and \U$37075 ( \37419 , \37413 , \37417 );
or \U$37076 ( \37420 , \37416 , \37418 , \37419 );
and \U$37077 ( \37421 , \37411 , \37420 );
xor \U$37078 ( \37422 , \37182 , \37184 );
xor \U$37079 ( \37423 , \37422 , \37186 );
and \U$37080 ( \37424 , \37420 , \37423 );
and \U$37081 ( \37425 , \37411 , \37423 );
or \U$37082 ( \37426 , \37421 , \37424 , \37425 );
xor \U$37083 ( \37427 , \36930 , \36940 );
xor \U$37084 ( \37428 , \37427 , \36946 );
and \U$37085 ( \37429 , \37426 , \37428 );
xor \U$37086 ( \37430 , \37180 , \37189 );
xor \U$37087 ( \37431 , \37430 , \37192 );
and \U$37088 ( \37432 , \37428 , \37431 );
and \U$37089 ( \37433 , \37426 , \37431 );
or \U$37090 ( \37434 , \37429 , \37432 , \37433 );
and \U$37091 ( \37435 , \37207 , \37434 );
xor \U$37092 ( \37436 , \37207 , \37434 );
xor \U$37093 ( \37437 , \37426 , \37428 );
xor \U$37094 ( \37438 , \37437 , \37431 );
and \U$37095 ( \37439 , \27830 , \24462 );
and \U$37096 ( \37440 , \27527 , \24460 );
nor \U$37097 ( \37441 , \37439 , \37440 );
xnor \U$37098 ( \37442 , \37441 , \24275 );
and \U$37099 ( \37443 , \28528 , \24149 );
and \U$37100 ( \37444 , \28002 , \24147 );
nor \U$37101 ( \37445 , \37443 , \37444 );
xnor \U$37102 ( \37446 , \37445 , \23944 );
and \U$37103 ( \37447 , \37442 , \37446 );
and \U$37104 ( \37448 , \29198 , \23743 );
and \U$37105 ( \37449 , \28952 , \23741 );
nor \U$37106 ( \37450 , \37448 , \37449 );
xnor \U$37107 ( \37451 , \37450 , \23594 );
and \U$37108 ( \37452 , \37446 , \37451 );
and \U$37109 ( \37453 , \37442 , \37451 );
or \U$37110 ( \37454 , \37447 , \37452 , \37453 );
and \U$37111 ( \37455 , \25097 , \27060 );
and \U$37112 ( \37456 , \24841 , \27058 );
nor \U$37113 ( \37457 , \37455 , \37456 );
xnor \U$37114 ( \37458 , \37457 , \26720 );
and \U$37115 ( \37459 , \25596 , \26471 );
and \U$37116 ( \37460 , \25294 , \26469 );
nor \U$37117 ( \37461 , \37459 , \37460 );
xnor \U$37118 ( \37462 , \37461 , \26230 );
and \U$37119 ( \37463 , \37458 , \37462 );
and \U$37120 ( \37464 , \26073 , \26005 );
and \U$37121 ( \37465 , \25604 , \26003 );
nor \U$37122 ( \37466 , \37464 , \37465 );
xnor \U$37123 ( \37467 , \37466 , \25817 );
and \U$37124 ( \37468 , \37462 , \37467 );
and \U$37125 ( \37469 , \37458 , \37467 );
or \U$37126 ( \37470 , \37463 , \37468 , \37469 );
and \U$37127 ( \37471 , \37454 , \37470 );
and \U$37128 ( \37472 , \26342 , \25631 );
and \U$37129 ( \37473 , \26078 , \25629 );
nor \U$37130 ( \37474 , \37472 , \37473 );
xnor \U$37131 ( \37475 , \37474 , \25399 );
and \U$37132 ( \37476 , \26973 , \25180 );
and \U$37133 ( \37477 , \26601 , \25178 );
nor \U$37134 ( \37478 , \37476 , \37477 );
xnor \U$37135 ( \37479 , \37478 , \25037 );
and \U$37136 ( \37480 , \37475 , \37479 );
and \U$37137 ( \37481 , \27325 , \24857 );
and \U$37138 ( \37482 , \26982 , \24855 );
nor \U$37139 ( \37483 , \37481 , \37482 );
xnor \U$37140 ( \37484 , \37483 , \24611 );
and \U$37141 ( \37485 , \37479 , \37484 );
and \U$37142 ( \37486 , \37475 , \37484 );
or \U$37143 ( \37487 , \37480 , \37485 , \37486 );
and \U$37144 ( \37488 , \37470 , \37487 );
and \U$37145 ( \37489 , \37454 , \37487 );
or \U$37146 ( \37490 , \37471 , \37488 , \37489 );
and \U$37147 ( \37491 , \22616 , \31639 );
and \U$37148 ( \37492 , \22440 , \31636 );
nor \U$37149 ( \37493 , \37491 , \37492 );
xnor \U$37150 ( \37494 , \37493 , \30584 );
and \U$37151 ( \37495 , \22867 , \30826 );
and \U$37152 ( \37496 , \22624 , \30824 );
nor \U$37153 ( \37497 , \37495 , \37496 );
xnor \U$37154 ( \37498 , \37497 , \30587 );
and \U$37155 ( \37499 , \37494 , \37498 );
and \U$37156 ( \37500 , \37498 , \22266 );
and \U$37157 ( \37501 , \37494 , \22266 );
or \U$37158 ( \37502 , \37499 , \37500 , \37501 );
and \U$37159 ( \37503 , \23970 , \28592 );
and \U$37160 ( \37504 , \23832 , \28590 );
nor \U$37161 ( \37505 , \37503 , \37504 );
xnor \U$37162 ( \37506 , \37505 , \28343 );
and \U$37163 ( \37507 , \24506 , \28063 );
and \U$37164 ( \37508 , \24089 , \28061 );
nor \U$37165 ( \37509 , \37507 , \37508 );
xnor \U$37166 ( \37510 , \37509 , \27803 );
and \U$37167 ( \37511 , \37506 , \37510 );
and \U$37168 ( \37512 , \24836 , \27569 );
and \U$37169 ( \37513 , \24714 , \27567 );
nor \U$37170 ( \37514 , \37512 , \37513 );
xnor \U$37171 ( \37515 , \37514 , \27254 );
and \U$37172 ( \37516 , \37510 , \37515 );
and \U$37173 ( \37517 , \37506 , \37515 );
or \U$37174 ( \37518 , \37511 , \37516 , \37517 );
and \U$37175 ( \37519 , \37502 , \37518 );
and \U$37176 ( \37520 , \23058 , \30258 );
and \U$37177 ( \37521 , \22872 , \30256 );
nor \U$37178 ( \37522 , \37520 , \37521 );
xnor \U$37179 ( \37523 , \37522 , \29948 );
and \U$37180 ( \37524 , \23466 , \29721 );
and \U$37181 ( \37525 , \23202 , \29719 );
nor \U$37182 ( \37526 , \37524 , \37525 );
xnor \U$37183 ( \37527 , \37526 , \29350 );
and \U$37184 ( \37528 , \37523 , \37527 );
and \U$37185 ( \37529 , \23665 , \29159 );
and \U$37186 ( \37530 , \23491 , \29157 );
nor \U$37187 ( \37531 , \37529 , \37530 );
xnor \U$37188 ( \37532 , \37531 , \28841 );
and \U$37189 ( \37533 , \37527 , \37532 );
and \U$37190 ( \37534 , \37523 , \37532 );
or \U$37191 ( \37535 , \37528 , \37533 , \37534 );
and \U$37192 ( \37536 , \37518 , \37535 );
and \U$37193 ( \37537 , \37502 , \37535 );
or \U$37194 ( \37538 , \37519 , \37536 , \37537 );
and \U$37195 ( \37539 , \37490 , \37538 );
and \U$37196 ( \37540 , \29522 , \23421 );
and \U$37197 ( \37541 , \29203 , \23419 );
nor \U$37198 ( \37542 , \37540 , \37541 );
xnor \U$37199 ( \37543 , \37542 , \23279 );
and \U$37200 ( \37544 , \30375 , \23125 );
and \U$37201 ( \37545 , \29806 , \23123 );
nor \U$37202 ( \37546 , \37544 , \37545 );
xnor \U$37203 ( \37547 , \37546 , \22988 );
and \U$37204 ( \37548 , \37543 , \37547 );
and \U$37205 ( \37549 , \30986 , \22919 );
and \U$37206 ( \37550 , \30383 , \22917 );
nor \U$37207 ( \37551 , \37549 , \37550 );
xnor \U$37208 ( \37552 , \37551 , \22767 );
and \U$37209 ( \37553 , \37547 , \37552 );
and \U$37210 ( \37554 , \37543 , \37552 );
or \U$37211 ( \37555 , \37548 , \37553 , \37554 );
and \U$37212 ( \37556 , \31172 , \22651 );
and \U$37213 ( \37557 , \30991 , \22649 );
nor \U$37214 ( \37558 , \37556 , \37557 );
xnor \U$37215 ( \37559 , \37558 , \22495 );
nand \U$37216 ( \37560 , \31792 , \22377 );
xnor \U$37217 ( \37561 , \37560 , \22266 );
and \U$37218 ( \37562 , \37559 , \37561 );
and \U$37219 ( \37563 , \37555 , \37562 );
and \U$37220 ( \37564 , \31792 , \22379 );
and \U$37221 ( \37565 , \31172 , \22377 );
nor \U$37222 ( \37566 , \37564 , \37565 );
xnor \U$37223 ( \37567 , \37566 , \22266 );
and \U$37224 ( \37568 , \37562 , \37567 );
and \U$37225 ( \37569 , \37555 , \37567 );
or \U$37226 ( \37570 , \37563 , \37568 , \37569 );
and \U$37227 ( \37571 , \37538 , \37570 );
and \U$37228 ( \37572 , \37490 , \37570 );
or \U$37229 ( \37573 , \37539 , \37571 , \37572 );
xor \U$37230 ( \37574 , \37227 , \37231 );
xor \U$37231 ( \37575 , \37574 , \37236 );
xor \U$37232 ( \37576 , \37296 , \37300 );
xor \U$37233 ( \37577 , \37576 , \37305 );
and \U$37234 ( \37578 , \37575 , \37577 );
xor \U$37235 ( \37579 , \37244 , \37248 );
xor \U$37236 ( \37580 , \37579 , \37253 );
and \U$37237 ( \37581 , \37577 , \37580 );
and \U$37238 ( \37582 , \37575 , \37580 );
or \U$37239 ( \37583 , \37578 , \37581 , \37582 );
xor \U$37240 ( \37584 , \37263 , \37267 );
xor \U$37241 ( \37585 , \37584 , \37272 );
xor \U$37242 ( \37586 , \37316 , \37320 );
xor \U$37243 ( \37587 , \37586 , \37325 );
and \U$37244 ( \37588 , \37585 , \37587 );
xor \U$37245 ( \37589 , \37279 , \37283 );
xor \U$37246 ( \37590 , \37589 , \37288 );
and \U$37247 ( \37591 , \37587 , \37590 );
and \U$37248 ( \37592 , \37585 , \37590 );
or \U$37249 ( \37593 , \37588 , \37591 , \37592 );
and \U$37250 ( \37594 , \37583 , \37593 );
xor \U$37251 ( \37595 , \37351 , \37353 );
xor \U$37252 ( \37596 , \37595 , \37356 );
and \U$37253 ( \37597 , \37593 , \37596 );
and \U$37254 ( \37598 , \37583 , \37596 );
or \U$37255 ( \37599 , \37594 , \37597 , \37598 );
and \U$37256 ( \37600 , \37573 , \37599 );
xor \U$37257 ( \37601 , \37275 , \37291 );
xor \U$37258 ( \37602 , \37601 , \37308 );
xor \U$37259 ( \37603 , \37341 , \37343 );
xor \U$37260 ( \37604 , \37603 , \37346 );
and \U$37261 ( \37605 , \37602 , \37604 );
xor \U$37262 ( \37606 , \37328 , \37330 );
xor \U$37263 ( \37607 , \37606 , \37333 );
and \U$37264 ( \37608 , \37604 , \37607 );
and \U$37265 ( \37609 , \37602 , \37607 );
or \U$37266 ( \37610 , \37605 , \37608 , \37609 );
and \U$37267 ( \37611 , \37599 , \37610 );
and \U$37268 ( \37612 , \37573 , \37610 );
or \U$37269 ( \37613 , \37600 , \37611 , \37612 );
xor \U$37270 ( \37614 , \37381 , \37383 );
xor \U$37271 ( \37615 , \37614 , \37386 );
xor \U$37272 ( \37616 , \37349 , \37359 );
xor \U$37273 ( \37617 , \37616 , \37362 );
and \U$37274 ( \37618 , \37615 , \37617 );
xor \U$37275 ( \37619 , \37368 , \37370 );
xor \U$37276 ( \37620 , \37619 , \37373 );
and \U$37277 ( \37621 , \37617 , \37620 );
and \U$37278 ( \37622 , \37615 , \37620 );
or \U$37279 ( \37623 , \37618 , \37621 , \37622 );
and \U$37280 ( \37624 , \37613 , \37623 );
xor \U$37281 ( \37625 , \37400 , \37402 );
xor \U$37282 ( \37626 , \37625 , \37405 );
and \U$37283 ( \37627 , \37623 , \37626 );
and \U$37284 ( \37628 , \37613 , \37626 );
or \U$37285 ( \37629 , \37624 , \37627 , \37628 );
xor \U$37286 ( \37630 , \37379 , \37397 );
xor \U$37287 ( \37631 , \37630 , \37408 );
and \U$37288 ( \37632 , \37629 , \37631 );
xor \U$37289 ( \37633 , \37413 , \37415 );
xor \U$37290 ( \37634 , \37633 , \37417 );
and \U$37291 ( \37635 , \37631 , \37634 );
and \U$37292 ( \37636 , \37629 , \37634 );
or \U$37293 ( \37637 , \37632 , \37635 , \37636 );
xor \U$37294 ( \37638 , \37161 , \37171 );
xor \U$37295 ( \37639 , \37638 , \37177 );
and \U$37296 ( \37640 , \37637 , \37639 );
xor \U$37297 ( \37641 , \37411 , \37420 );
xor \U$37298 ( \37642 , \37641 , \37423 );
and \U$37299 ( \37643 , \37639 , \37642 );
and \U$37300 ( \37644 , \37637 , \37642 );
or \U$37301 ( \37645 , \37640 , \37643 , \37644 );
and \U$37302 ( \37646 , \37438 , \37645 );
xor \U$37303 ( \37647 , \37438 , \37645 );
xor \U$37304 ( \37648 , \37637 , \37639 );
xor \U$37305 ( \37649 , \37648 , \37642 );
and \U$37306 ( \37650 , \26982 , \25180 );
and \U$37307 ( \37651 , \26973 , \25178 );
nor \U$37308 ( \37652 , \37650 , \37651 );
xnor \U$37309 ( \37653 , \37652 , \25037 );
and \U$37310 ( \37654 , \27527 , \24857 );
and \U$37311 ( \37655 , \27325 , \24855 );
nor \U$37312 ( \37656 , \37654 , \37655 );
xnor \U$37313 ( \37657 , \37656 , \24611 );
and \U$37314 ( \37658 , \37653 , \37657 );
and \U$37315 ( \37659 , \28002 , \24462 );
and \U$37316 ( \37660 , \27830 , \24460 );
nor \U$37317 ( \37661 , \37659 , \37660 );
xnor \U$37318 ( \37662 , \37661 , \24275 );
and \U$37319 ( \37663 , \37657 , \37662 );
and \U$37320 ( \37664 , \37653 , \37662 );
or \U$37321 ( \37665 , \37658 , \37663 , \37664 );
and \U$37322 ( \37666 , \28952 , \24149 );
and \U$37323 ( \37667 , \28528 , \24147 );
nor \U$37324 ( \37668 , \37666 , \37667 );
xnor \U$37325 ( \37669 , \37668 , \23944 );
and \U$37326 ( \37670 , \29203 , \23743 );
and \U$37327 ( \37671 , \29198 , \23741 );
nor \U$37328 ( \37672 , \37670 , \37671 );
xnor \U$37329 ( \37673 , \37672 , \23594 );
and \U$37330 ( \37674 , \37669 , \37673 );
and \U$37331 ( \37675 , \29806 , \23421 );
and \U$37332 ( \37676 , \29522 , \23419 );
nor \U$37333 ( \37677 , \37675 , \37676 );
xnor \U$37334 ( \37678 , \37677 , \23279 );
and \U$37335 ( \37679 , \37673 , \37678 );
and \U$37336 ( \37680 , \37669 , \37678 );
or \U$37337 ( \37681 , \37674 , \37679 , \37680 );
and \U$37338 ( \37682 , \37665 , \37681 );
and \U$37339 ( \37683 , \25604 , \26471 );
and \U$37340 ( \37684 , \25596 , \26469 );
nor \U$37341 ( \37685 , \37683 , \37684 );
xnor \U$37342 ( \37686 , \37685 , \26230 );
and \U$37343 ( \37687 , \26078 , \26005 );
and \U$37344 ( \37688 , \26073 , \26003 );
nor \U$37345 ( \37689 , \37687 , \37688 );
xnor \U$37346 ( \37690 , \37689 , \25817 );
and \U$37347 ( \37691 , \37686 , \37690 );
and \U$37348 ( \37692 , \26601 , \25631 );
and \U$37349 ( \37693 , \26342 , \25629 );
nor \U$37350 ( \37694 , \37692 , \37693 );
xnor \U$37351 ( \37695 , \37694 , \25399 );
and \U$37352 ( \37696 , \37690 , \37695 );
and \U$37353 ( \37697 , \37686 , \37695 );
or \U$37354 ( \37698 , \37691 , \37696 , \37697 );
and \U$37355 ( \37699 , \37681 , \37698 );
and \U$37356 ( \37700 , \37665 , \37698 );
or \U$37357 ( \37701 , \37682 , \37699 , \37700 );
and \U$37358 ( \37702 , \24714 , \28063 );
and \U$37359 ( \37703 , \24506 , \28061 );
nor \U$37360 ( \37704 , \37702 , \37703 );
xnor \U$37361 ( \37705 , \37704 , \27803 );
and \U$37362 ( \37706 , \24841 , \27569 );
and \U$37363 ( \37707 , \24836 , \27567 );
nor \U$37364 ( \37708 , \37706 , \37707 );
xnor \U$37365 ( \37709 , \37708 , \27254 );
and \U$37366 ( \37710 , \37705 , \37709 );
and \U$37367 ( \37711 , \25294 , \27060 );
and \U$37368 ( \37712 , \25097 , \27058 );
nor \U$37369 ( \37713 , \37711 , \37712 );
xnor \U$37370 ( \37714 , \37713 , \26720 );
and \U$37371 ( \37715 , \37709 , \37714 );
and \U$37372 ( \37716 , \37705 , \37714 );
or \U$37373 ( \37717 , \37710 , \37715 , \37716 );
and \U$37374 ( \37718 , \23491 , \29721 );
and \U$37375 ( \37719 , \23466 , \29719 );
nor \U$37376 ( \37720 , \37718 , \37719 );
xnor \U$37377 ( \37721 , \37720 , \29350 );
and \U$37378 ( \37722 , \23832 , \29159 );
and \U$37379 ( \37723 , \23665 , \29157 );
nor \U$37380 ( \37724 , \37722 , \37723 );
xnor \U$37381 ( \37725 , \37724 , \28841 );
and \U$37382 ( \37726 , \37721 , \37725 );
and \U$37383 ( \37727 , \24089 , \28592 );
and \U$37384 ( \37728 , \23970 , \28590 );
nor \U$37385 ( \37729 , \37727 , \37728 );
xnor \U$37386 ( \37730 , \37729 , \28343 );
and \U$37387 ( \37731 , \37725 , \37730 );
and \U$37388 ( \37732 , \37721 , \37730 );
or \U$37389 ( \37733 , \37726 , \37731 , \37732 );
and \U$37390 ( \37734 , \37717 , \37733 );
and \U$37391 ( \37735 , \22624 , \31639 );
and \U$37392 ( \37736 , \22616 , \31636 );
nor \U$37393 ( \37737 , \37735 , \37736 );
xnor \U$37394 ( \37738 , \37737 , \30584 );
and \U$37395 ( \37739 , \22872 , \30826 );
and \U$37396 ( \37740 , \22867 , \30824 );
nor \U$37397 ( \37741 , \37739 , \37740 );
xnor \U$37398 ( \37742 , \37741 , \30587 );
and \U$37399 ( \37743 , \37738 , \37742 );
and \U$37400 ( \37744 , \23202 , \30258 );
and \U$37401 ( \37745 , \23058 , \30256 );
nor \U$37402 ( \37746 , \37744 , \37745 );
xnor \U$37403 ( \37747 , \37746 , \29948 );
and \U$37404 ( \37748 , \37742 , \37747 );
and \U$37405 ( \37749 , \37738 , \37747 );
or \U$37406 ( \37750 , \37743 , \37748 , \37749 );
and \U$37407 ( \37751 , \37733 , \37750 );
and \U$37408 ( \37752 , \37717 , \37750 );
or \U$37409 ( \37753 , \37734 , \37751 , \37752 );
and \U$37410 ( \37754 , \37701 , \37753 );
and \U$37411 ( \37755 , \30383 , \23125 );
and \U$37412 ( \37756 , \30375 , \23123 );
nor \U$37413 ( \37757 , \37755 , \37756 );
xnor \U$37414 ( \37758 , \37757 , \22988 );
and \U$37415 ( \37759 , \30991 , \22919 );
and \U$37416 ( \37760 , \30986 , \22917 );
nor \U$37417 ( \37761 , \37759 , \37760 );
xnor \U$37418 ( \37762 , \37761 , \22767 );
and \U$37419 ( \37763 , \37758 , \37762 );
and \U$37420 ( \37764 , \31792 , \22651 );
and \U$37421 ( \37765 , \31172 , \22649 );
nor \U$37422 ( \37766 , \37764 , \37765 );
xnor \U$37423 ( \37767 , \37766 , \22495 );
and \U$37424 ( \37768 , \37762 , \37767 );
and \U$37425 ( \37769 , \37758 , \37767 );
or \U$37426 ( \37770 , \37763 , \37768 , \37769 );
xor \U$37427 ( \37771 , \37543 , \37547 );
xor \U$37428 ( \37772 , \37771 , \37552 );
and \U$37429 ( \37773 , \37770 , \37772 );
xor \U$37430 ( \37774 , \37559 , \37561 );
and \U$37431 ( \37775 , \37772 , \37774 );
and \U$37432 ( \37776 , \37770 , \37774 );
or \U$37433 ( \37777 , \37773 , \37775 , \37776 );
and \U$37434 ( \37778 , \37753 , \37777 );
and \U$37435 ( \37779 , \37701 , \37777 );
or \U$37436 ( \37780 , \37754 , \37778 , \37779 );
xor \U$37437 ( \37781 , \37494 , \37498 );
xor \U$37438 ( \37782 , \37781 , \22266 );
xor \U$37439 ( \37783 , \37506 , \37510 );
xor \U$37440 ( \37784 , \37783 , \37515 );
and \U$37441 ( \37785 , \37782 , \37784 );
xor \U$37442 ( \37786 , \37523 , \37527 );
xor \U$37443 ( \37787 , \37786 , \37532 );
and \U$37444 ( \37788 , \37784 , \37787 );
and \U$37445 ( \37789 , \37782 , \37787 );
or \U$37446 ( \37790 , \37785 , \37788 , \37789 );
xor \U$37447 ( \37791 , \37442 , \37446 );
xor \U$37448 ( \37792 , \37791 , \37451 );
xor \U$37449 ( \37793 , \37458 , \37462 );
xor \U$37450 ( \37794 , \37793 , \37467 );
and \U$37451 ( \37795 , \37792 , \37794 );
xor \U$37452 ( \37796 , \37475 , \37479 );
xor \U$37453 ( \37797 , \37796 , \37484 );
and \U$37454 ( \37798 , \37794 , \37797 );
and \U$37455 ( \37799 , \37792 , \37797 );
or \U$37456 ( \37800 , \37795 , \37798 , \37799 );
and \U$37457 ( \37801 , \37790 , \37800 );
xor \U$37458 ( \37802 , \37211 , \37215 );
xor \U$37459 ( \37803 , \37802 , \37220 );
and \U$37460 ( \37804 , \37800 , \37803 );
and \U$37461 ( \37805 , \37790 , \37803 );
or \U$37462 ( \37806 , \37801 , \37804 , \37805 );
and \U$37463 ( \37807 , \37780 , \37806 );
xor \U$37464 ( \37808 , \37555 , \37562 );
xor \U$37465 ( \37809 , \37808 , \37567 );
xor \U$37466 ( \37810 , \37575 , \37577 );
xor \U$37467 ( \37811 , \37810 , \37580 );
and \U$37468 ( \37812 , \37809 , \37811 );
xor \U$37469 ( \37813 , \37585 , \37587 );
xor \U$37470 ( \37814 , \37813 , \37590 );
and \U$37471 ( \37815 , \37811 , \37814 );
and \U$37472 ( \37816 , \37809 , \37814 );
or \U$37473 ( \37817 , \37812 , \37815 , \37816 );
and \U$37474 ( \37818 , \37806 , \37817 );
and \U$37475 ( \37819 , \37780 , \37817 );
or \U$37476 ( \37820 , \37807 , \37818 , \37819 );
xor \U$37477 ( \37821 , \37223 , \37239 );
xor \U$37478 ( \37822 , \37821 , \37256 );
xor \U$37479 ( \37823 , \37583 , \37593 );
xor \U$37480 ( \37824 , \37823 , \37596 );
and \U$37481 ( \37825 , \37822 , \37824 );
xor \U$37482 ( \37826 , \37602 , \37604 );
xor \U$37483 ( \37827 , \37826 , \37607 );
and \U$37484 ( \37828 , \37824 , \37827 );
and \U$37485 ( \37829 , \37822 , \37827 );
or \U$37486 ( \37830 , \37825 , \37828 , \37829 );
and \U$37487 ( \37831 , \37820 , \37830 );
xor \U$37488 ( \37832 , \37259 , \37311 );
xor \U$37489 ( \37833 , \37832 , \37336 );
and \U$37490 ( \37834 , \37830 , \37833 );
and \U$37491 ( \37835 , \37820 , \37833 );
or \U$37492 ( \37836 , \37831 , \37834 , \37835 );
xor \U$37493 ( \37837 , \37573 , \37599 );
xor \U$37494 ( \37838 , \37837 , \37610 );
xor \U$37495 ( \37839 , \37615 , \37617 );
xor \U$37496 ( \37840 , \37839 , \37620 );
and \U$37497 ( \37841 , \37838 , \37840 );
and \U$37498 ( \37842 , \37836 , \37841 );
xor \U$37499 ( \37843 , \37389 , \37391 );
xor \U$37500 ( \37844 , \37843 , \37394 );
and \U$37501 ( \37845 , \37841 , \37844 );
and \U$37502 ( \37846 , \37836 , \37844 );
or \U$37503 ( \37847 , \37842 , \37845 , \37846 );
xor \U$37504 ( \37848 , \37339 , \37365 );
xor \U$37505 ( \37849 , \37848 , \37376 );
xor \U$37506 ( \37850 , \37613 , \37623 );
xor \U$37507 ( \37851 , \37850 , \37626 );
and \U$37508 ( \37852 , \37849 , \37851 );
and \U$37509 ( \37853 , \37847 , \37852 );
xor \U$37510 ( \37854 , \37629 , \37631 );
xor \U$37511 ( \37855 , \37854 , \37634 );
and \U$37512 ( \37856 , \37852 , \37855 );
and \U$37513 ( \37857 , \37847 , \37855 );
or \U$37514 ( \37858 , \37853 , \37856 , \37857 );
and \U$37515 ( \37859 , \37649 , \37858 );
xor \U$37516 ( \37860 , \37649 , \37858 );
xor \U$37517 ( \37861 , \37847 , \37852 );
xor \U$37518 ( \37862 , \37861 , \37855 );
and \U$37519 ( \37863 , \24506 , \28592 );
and \U$37520 ( \37864 , \24089 , \28590 );
nor \U$37521 ( \37865 , \37863 , \37864 );
xnor \U$37522 ( \37866 , \37865 , \28343 );
and \U$37523 ( \37867 , \24836 , \28063 );
and \U$37524 ( \37868 , \24714 , \28061 );
nor \U$37525 ( \37869 , \37867 , \37868 );
xnor \U$37526 ( \37870 , \37869 , \27803 );
and \U$37527 ( \37871 , \37866 , \37870 );
and \U$37528 ( \37872 , \25097 , \27569 );
and \U$37529 ( \37873 , \24841 , \27567 );
nor \U$37530 ( \37874 , \37872 , \37873 );
xnor \U$37531 ( \37875 , \37874 , \27254 );
and \U$37532 ( \37876 , \37870 , \37875 );
and \U$37533 ( \37877 , \37866 , \37875 );
or \U$37534 ( \37878 , \37871 , \37876 , \37877 );
and \U$37535 ( \37879 , \23466 , \30258 );
and \U$37536 ( \37880 , \23202 , \30256 );
nor \U$37537 ( \37881 , \37879 , \37880 );
xnor \U$37538 ( \37882 , \37881 , \29948 );
and \U$37539 ( \37883 , \23665 , \29721 );
and \U$37540 ( \37884 , \23491 , \29719 );
nor \U$37541 ( \37885 , \37883 , \37884 );
xnor \U$37542 ( \37886 , \37885 , \29350 );
and \U$37543 ( \37887 , \37882 , \37886 );
and \U$37544 ( \37888 , \23970 , \29159 );
and \U$37545 ( \37889 , \23832 , \29157 );
nor \U$37546 ( \37890 , \37888 , \37889 );
xnor \U$37547 ( \37891 , \37890 , \28841 );
and \U$37548 ( \37892 , \37886 , \37891 );
and \U$37549 ( \37893 , \37882 , \37891 );
or \U$37550 ( \37894 , \37887 , \37892 , \37893 );
and \U$37551 ( \37895 , \37878 , \37894 );
and \U$37552 ( \37896 , \22867 , \31639 );
and \U$37553 ( \37897 , \22624 , \31636 );
nor \U$37554 ( \37898 , \37896 , \37897 );
xnor \U$37555 ( \37899 , \37898 , \30584 );
and \U$37556 ( \37900 , \23058 , \30826 );
and \U$37557 ( \37901 , \22872 , \30824 );
nor \U$37558 ( \37902 , \37900 , \37901 );
xnor \U$37559 ( \37903 , \37902 , \30587 );
and \U$37560 ( \37904 , \37899 , \37903 );
and \U$37561 ( \37905 , \37903 , \22495 );
and \U$37562 ( \37906 , \37899 , \22495 );
or \U$37563 ( \37907 , \37904 , \37905 , \37906 );
and \U$37564 ( \37908 , \37894 , \37907 );
and \U$37565 ( \37909 , \37878 , \37907 );
or \U$37566 ( \37910 , \37895 , \37908 , \37909 );
and \U$37567 ( \37911 , \28528 , \24462 );
and \U$37568 ( \37912 , \28002 , \24460 );
nor \U$37569 ( \37913 , \37911 , \37912 );
xnor \U$37570 ( \37914 , \37913 , \24275 );
and \U$37571 ( \37915 , \29198 , \24149 );
and \U$37572 ( \37916 , \28952 , \24147 );
nor \U$37573 ( \37917 , \37915 , \37916 );
xnor \U$37574 ( \37918 , \37917 , \23944 );
and \U$37575 ( \37919 , \37914 , \37918 );
and \U$37576 ( \37920 , \29522 , \23743 );
and \U$37577 ( \37921 , \29203 , \23741 );
nor \U$37578 ( \37922 , \37920 , \37921 );
xnor \U$37579 ( \37923 , \37922 , \23594 );
and \U$37580 ( \37924 , \37918 , \37923 );
and \U$37581 ( \37925 , \37914 , \37923 );
or \U$37582 ( \37926 , \37919 , \37924 , \37925 );
and \U$37583 ( \37927 , \25596 , \27060 );
and \U$37584 ( \37928 , \25294 , \27058 );
nor \U$37585 ( \37929 , \37927 , \37928 );
xnor \U$37586 ( \37930 , \37929 , \26720 );
and \U$37587 ( \37931 , \26073 , \26471 );
and \U$37588 ( \37932 , \25604 , \26469 );
nor \U$37589 ( \37933 , \37931 , \37932 );
xnor \U$37590 ( \37934 , \37933 , \26230 );
and \U$37591 ( \37935 , \37930 , \37934 );
and \U$37592 ( \37936 , \26342 , \26005 );
and \U$37593 ( \37937 , \26078 , \26003 );
nor \U$37594 ( \37938 , \37936 , \37937 );
xnor \U$37595 ( \37939 , \37938 , \25817 );
and \U$37596 ( \37940 , \37934 , \37939 );
and \U$37597 ( \37941 , \37930 , \37939 );
or \U$37598 ( \37942 , \37935 , \37940 , \37941 );
and \U$37599 ( \37943 , \37926 , \37942 );
and \U$37600 ( \37944 , \26973 , \25631 );
and \U$37601 ( \37945 , \26601 , \25629 );
nor \U$37602 ( \37946 , \37944 , \37945 );
xnor \U$37603 ( \37947 , \37946 , \25399 );
and \U$37604 ( \37948 , \27325 , \25180 );
and \U$37605 ( \37949 , \26982 , \25178 );
nor \U$37606 ( \37950 , \37948 , \37949 );
xnor \U$37607 ( \37951 , \37950 , \25037 );
and \U$37608 ( \37952 , \37947 , \37951 );
and \U$37609 ( \37953 , \27830 , \24857 );
and \U$37610 ( \37954 , \27527 , \24855 );
nor \U$37611 ( \37955 , \37953 , \37954 );
xnor \U$37612 ( \37956 , \37955 , \24611 );
and \U$37613 ( \37957 , \37951 , \37956 );
and \U$37614 ( \37958 , \37947 , \37956 );
or \U$37615 ( \37959 , \37952 , \37957 , \37958 );
and \U$37616 ( \37960 , \37942 , \37959 );
and \U$37617 ( \37961 , \37926 , \37959 );
or \U$37618 ( \37962 , \37943 , \37960 , \37961 );
and \U$37619 ( \37963 , \37910 , \37962 );
and \U$37620 ( \37964 , \30375 , \23421 );
and \U$37621 ( \37965 , \29806 , \23419 );
nor \U$37622 ( \37966 , \37964 , \37965 );
xnor \U$37623 ( \37967 , \37966 , \23279 );
and \U$37624 ( \37968 , \30986 , \23125 );
and \U$37625 ( \37969 , \30383 , \23123 );
nor \U$37626 ( \37970 , \37968 , \37969 );
xnor \U$37627 ( \37971 , \37970 , \22988 );
and \U$37628 ( \37972 , \37967 , \37971 );
and \U$37629 ( \37973 , \31172 , \22919 );
and \U$37630 ( \37974 , \30991 , \22917 );
nor \U$37631 ( \37975 , \37973 , \37974 );
xnor \U$37632 ( \37976 , \37975 , \22767 );
and \U$37633 ( \37977 , \37971 , \37976 );
and \U$37634 ( \37978 , \37967 , \37976 );
or \U$37635 ( \37979 , \37972 , \37977 , \37978 );
xor \U$37636 ( \37980 , \37669 , \37673 );
xor \U$37637 ( \37981 , \37980 , \37678 );
and \U$37638 ( \37982 , \37979 , \37981 );
xor \U$37639 ( \37983 , \37758 , \37762 );
xor \U$37640 ( \37984 , \37983 , \37767 );
and \U$37641 ( \37985 , \37981 , \37984 );
and \U$37642 ( \37986 , \37979 , \37984 );
or \U$37643 ( \37987 , \37982 , \37985 , \37986 );
and \U$37644 ( \37988 , \37962 , \37987 );
and \U$37645 ( \37989 , \37910 , \37987 );
or \U$37646 ( \37990 , \37963 , \37988 , \37989 );
xor \U$37647 ( \37991 , \37653 , \37657 );
xor \U$37648 ( \37992 , \37991 , \37662 );
xor \U$37649 ( \37993 , \37705 , \37709 );
xor \U$37650 ( \37994 , \37993 , \37714 );
and \U$37651 ( \37995 , \37992 , \37994 );
xor \U$37652 ( \37996 , \37686 , \37690 );
xor \U$37653 ( \37997 , \37996 , \37695 );
and \U$37654 ( \37998 , \37994 , \37997 );
and \U$37655 ( \37999 , \37992 , \37997 );
or \U$37656 ( \38000 , \37995 , \37998 , \37999 );
xor \U$37657 ( \38001 , \37721 , \37725 );
xor \U$37658 ( \38002 , \38001 , \37730 );
xor \U$37659 ( \38003 , \37738 , \37742 );
xor \U$37660 ( \38004 , \38003 , \37747 );
and \U$37661 ( \38005 , \38002 , \38004 );
and \U$37662 ( \38006 , \38000 , \38005 );
xor \U$37663 ( \38007 , \37782 , \37784 );
xor \U$37664 ( \38008 , \38007 , \37787 );
and \U$37665 ( \38009 , \38005 , \38008 );
and \U$37666 ( \38010 , \38000 , \38008 );
or \U$37667 ( \38011 , \38006 , \38009 , \38010 );
and \U$37668 ( \38012 , \37990 , \38011 );
xor \U$37669 ( \38013 , \37665 , \37681 );
xor \U$37670 ( \38014 , \38013 , \37698 );
xor \U$37671 ( \38015 , \37792 , \37794 );
xor \U$37672 ( \38016 , \38015 , \37797 );
and \U$37673 ( \38017 , \38014 , \38016 );
xor \U$37674 ( \38018 , \37770 , \37772 );
xor \U$37675 ( \38019 , \38018 , \37774 );
and \U$37676 ( \38020 , \38016 , \38019 );
and \U$37677 ( \38021 , \38014 , \38019 );
or \U$37678 ( \38022 , \38017 , \38020 , \38021 );
and \U$37679 ( \38023 , \38011 , \38022 );
and \U$37680 ( \38024 , \37990 , \38022 );
or \U$37681 ( \38025 , \38012 , \38023 , \38024 );
xor \U$37682 ( \38026 , \37454 , \37470 );
xor \U$37683 ( \38027 , \38026 , \37487 );
xor \U$37684 ( \38028 , \37502 , \37518 );
xor \U$37685 ( \38029 , \38028 , \37535 );
and \U$37686 ( \38030 , \38027 , \38029 );
xor \U$37687 ( \38031 , \37809 , \37811 );
xor \U$37688 ( \38032 , \38031 , \37814 );
and \U$37689 ( \38033 , \38029 , \38032 );
and \U$37690 ( \38034 , \38027 , \38032 );
or \U$37691 ( \38035 , \38030 , \38033 , \38034 );
and \U$37692 ( \38036 , \38025 , \38035 );
xor \U$37693 ( \38037 , \37490 , \37538 );
xor \U$37694 ( \38038 , \38037 , \37570 );
and \U$37695 ( \38039 , \38035 , \38038 );
and \U$37696 ( \38040 , \38025 , \38038 );
or \U$37697 ( \38041 , \38036 , \38039 , \38040 );
xor \U$37698 ( \38042 , \37820 , \37830 );
xor \U$37699 ( \38043 , \38042 , \37833 );
and \U$37700 ( \38044 , \38041 , \38043 );
xor \U$37701 ( \38045 , \37838 , \37840 );
and \U$37702 ( \38046 , \38043 , \38045 );
and \U$37703 ( \38047 , \38041 , \38045 );
or \U$37704 ( \38048 , \38044 , \38046 , \38047 );
xor \U$37705 ( \38049 , \37836 , \37841 );
xor \U$37706 ( \38050 , \38049 , \37844 );
and \U$37707 ( \38051 , \38048 , \38050 );
xor \U$37708 ( \38052 , \37849 , \37851 );
and \U$37709 ( \38053 , \38050 , \38052 );
and \U$37710 ( \38054 , \38048 , \38052 );
or \U$37711 ( \38055 , \38051 , \38053 , \38054 );
and \U$37712 ( \38056 , \37862 , \38055 );
xor \U$37713 ( \38057 , \37862 , \38055 );
xor \U$37714 ( \38058 , \38048 , \38050 );
xor \U$37715 ( \38059 , \38058 , \38052 );
and \U$37716 ( \38060 , \22872 , \31639 );
and \U$37717 ( \38061 , \22867 , \31636 );
nor \U$37718 ( \38062 , \38060 , \38061 );
xnor \U$37719 ( \38063 , \38062 , \30584 );
and \U$37720 ( \38064 , \23202 , \30826 );
and \U$37721 ( \38065 , \23058 , \30824 );
nor \U$37722 ( \38066 , \38064 , \38065 );
xnor \U$37723 ( \38067 , \38066 , \30587 );
and \U$37724 ( \38068 , \38063 , \38067 );
and \U$37725 ( \38069 , \23491 , \30258 );
and \U$37726 ( \38070 , \23466 , \30256 );
nor \U$37727 ( \38071 , \38069 , \38070 );
xnor \U$37728 ( \38072 , \38071 , \29948 );
and \U$37729 ( \38073 , \38067 , \38072 );
and \U$37730 ( \38074 , \38063 , \38072 );
or \U$37731 ( \38075 , \38068 , \38073 , \38074 );
and \U$37732 ( \38076 , \23832 , \29721 );
and \U$37733 ( \38077 , \23665 , \29719 );
nor \U$37734 ( \38078 , \38076 , \38077 );
xnor \U$37735 ( \38079 , \38078 , \29350 );
and \U$37736 ( \38080 , \24089 , \29159 );
and \U$37737 ( \38081 , \23970 , \29157 );
nor \U$37738 ( \38082 , \38080 , \38081 );
xnor \U$37739 ( \38083 , \38082 , \28841 );
and \U$37740 ( \38084 , \38079 , \38083 );
and \U$37741 ( \38085 , \24714 , \28592 );
and \U$37742 ( \38086 , \24506 , \28590 );
nor \U$37743 ( \38087 , \38085 , \38086 );
xnor \U$37744 ( \38088 , \38087 , \28343 );
and \U$37745 ( \38089 , \38083 , \38088 );
and \U$37746 ( \38090 , \38079 , \38088 );
or \U$37747 ( \38091 , \38084 , \38089 , \38090 );
and \U$37748 ( \38092 , \38075 , \38091 );
and \U$37749 ( \38093 , \24841 , \28063 );
and \U$37750 ( \38094 , \24836 , \28061 );
nor \U$37751 ( \38095 , \38093 , \38094 );
xnor \U$37752 ( \38096 , \38095 , \27803 );
and \U$37753 ( \38097 , \25294 , \27569 );
and \U$37754 ( \38098 , \25097 , \27567 );
nor \U$37755 ( \38099 , \38097 , \38098 );
xnor \U$37756 ( \38100 , \38099 , \27254 );
and \U$37757 ( \38101 , \38096 , \38100 );
and \U$37758 ( \38102 , \25604 , \27060 );
and \U$37759 ( \38103 , \25596 , \27058 );
nor \U$37760 ( \38104 , \38102 , \38103 );
xnor \U$37761 ( \38105 , \38104 , \26720 );
and \U$37762 ( \38106 , \38100 , \38105 );
and \U$37763 ( \38107 , \38096 , \38105 );
or \U$37764 ( \38108 , \38101 , \38106 , \38107 );
and \U$37765 ( \38109 , \38091 , \38108 );
and \U$37766 ( \38110 , \38075 , \38108 );
or \U$37767 ( \38111 , \38092 , \38109 , \38110 );
and \U$37768 ( \38112 , \27527 , \25180 );
and \U$37769 ( \38113 , \27325 , \25178 );
nor \U$37770 ( \38114 , \38112 , \38113 );
xnor \U$37771 ( \38115 , \38114 , \25037 );
and \U$37772 ( \38116 , \28002 , \24857 );
and \U$37773 ( \38117 , \27830 , \24855 );
nor \U$37774 ( \38118 , \38116 , \38117 );
xnor \U$37775 ( \38119 , \38118 , \24611 );
and \U$37776 ( \38120 , \38115 , \38119 );
and \U$37777 ( \38121 , \28952 , \24462 );
and \U$37778 ( \38122 , \28528 , \24460 );
nor \U$37779 ( \38123 , \38121 , \38122 );
xnor \U$37780 ( \38124 , \38123 , \24275 );
and \U$37781 ( \38125 , \38119 , \38124 );
and \U$37782 ( \38126 , \38115 , \38124 );
or \U$37783 ( \38127 , \38120 , \38125 , \38126 );
and \U$37784 ( \38128 , \26078 , \26471 );
and \U$37785 ( \38129 , \26073 , \26469 );
nor \U$37786 ( \38130 , \38128 , \38129 );
xnor \U$37787 ( \38131 , \38130 , \26230 );
and \U$37788 ( \38132 , \26601 , \26005 );
and \U$37789 ( \38133 , \26342 , \26003 );
nor \U$37790 ( \38134 , \38132 , \38133 );
xnor \U$37791 ( \38135 , \38134 , \25817 );
and \U$37792 ( \38136 , \38131 , \38135 );
and \U$37793 ( \38137 , \26982 , \25631 );
and \U$37794 ( \38138 , \26973 , \25629 );
nor \U$37795 ( \38139 , \38137 , \38138 );
xnor \U$37796 ( \38140 , \38139 , \25399 );
and \U$37797 ( \38141 , \38135 , \38140 );
and \U$37798 ( \38142 , \38131 , \38140 );
or \U$37799 ( \38143 , \38136 , \38141 , \38142 );
and \U$37800 ( \38144 , \38127 , \38143 );
and \U$37801 ( \38145 , \29203 , \24149 );
and \U$37802 ( \38146 , \29198 , \24147 );
nor \U$37803 ( \38147 , \38145 , \38146 );
xnor \U$37804 ( \38148 , \38147 , \23944 );
and \U$37805 ( \38149 , \29806 , \23743 );
and \U$37806 ( \38150 , \29522 , \23741 );
nor \U$37807 ( \38151 , \38149 , \38150 );
xnor \U$37808 ( \38152 , \38151 , \23594 );
and \U$37809 ( \38153 , \38148 , \38152 );
and \U$37810 ( \38154 , \30383 , \23421 );
and \U$37811 ( \38155 , \30375 , \23419 );
nor \U$37812 ( \38156 , \38154 , \38155 );
xnor \U$37813 ( \38157 , \38156 , \23279 );
and \U$37814 ( \38158 , \38152 , \38157 );
and \U$37815 ( \38159 , \38148 , \38157 );
or \U$37816 ( \38160 , \38153 , \38158 , \38159 );
and \U$37817 ( \38161 , \38143 , \38160 );
and \U$37818 ( \38162 , \38127 , \38160 );
or \U$37819 ( \38163 , \38144 , \38161 , \38162 );
and \U$37820 ( \38164 , \38111 , \38163 );
nand \U$37821 ( \38165 , \31792 , \22649 );
xnor \U$37822 ( \38166 , \38165 , \22495 );
xor \U$37823 ( \38167 , \37914 , \37918 );
xor \U$37824 ( \38168 , \38167 , \37923 );
and \U$37825 ( \38169 , \38166 , \38168 );
xor \U$37826 ( \38170 , \37967 , \37971 );
xor \U$37827 ( \38171 , \38170 , \37976 );
and \U$37828 ( \38172 , \38168 , \38171 );
and \U$37829 ( \38173 , \38166 , \38171 );
or \U$37830 ( \38174 , \38169 , \38172 , \38173 );
and \U$37831 ( \38175 , \38163 , \38174 );
and \U$37832 ( \38176 , \38111 , \38174 );
or \U$37833 ( \38177 , \38164 , \38175 , \38176 );
xor \U$37834 ( \38178 , \37878 , \37894 );
xor \U$37835 ( \38179 , \38178 , \37907 );
xor \U$37836 ( \38180 , \37926 , \37942 );
xor \U$37837 ( \38181 , \38180 , \37959 );
and \U$37838 ( \38182 , \38179 , \38181 );
xor \U$37839 ( \38183 , \37979 , \37981 );
xor \U$37840 ( \38184 , \38183 , \37984 );
and \U$37841 ( \38185 , \38181 , \38184 );
and \U$37842 ( \38186 , \38179 , \38184 );
or \U$37843 ( \38187 , \38182 , \38185 , \38186 );
and \U$37844 ( \38188 , \38177 , \38187 );
xor \U$37845 ( \38189 , \37866 , \37870 );
xor \U$37846 ( \38190 , \38189 , \37875 );
xor \U$37847 ( \38191 , \37930 , \37934 );
xor \U$37848 ( \38192 , \38191 , \37939 );
and \U$37849 ( \38193 , \38190 , \38192 );
xor \U$37850 ( \38194 , \37947 , \37951 );
xor \U$37851 ( \38195 , \38194 , \37956 );
and \U$37852 ( \38196 , \38192 , \38195 );
and \U$37853 ( \38197 , \38190 , \38195 );
or \U$37854 ( \38198 , \38193 , \38196 , \38197 );
xor \U$37855 ( \38199 , \37992 , \37994 );
xor \U$37856 ( \38200 , \38199 , \37997 );
and \U$37857 ( \38201 , \38198 , \38200 );
xor \U$37858 ( \38202 , \38002 , \38004 );
and \U$37859 ( \38203 , \38200 , \38202 );
and \U$37860 ( \38204 , \38198 , \38202 );
or \U$37861 ( \38205 , \38201 , \38203 , \38204 );
and \U$37862 ( \38206 , \38187 , \38205 );
and \U$37863 ( \38207 , \38177 , \38205 );
or \U$37864 ( \38208 , \38188 , \38206 , \38207 );
xor \U$37865 ( \38209 , \37717 , \37733 );
xor \U$37866 ( \38210 , \38209 , \37750 );
xor \U$37867 ( \38211 , \38000 , \38005 );
xor \U$37868 ( \38212 , \38211 , \38008 );
and \U$37869 ( \38213 , \38210 , \38212 );
xor \U$37870 ( \38214 , \38014 , \38016 );
xor \U$37871 ( \38215 , \38214 , \38019 );
and \U$37872 ( \38216 , \38212 , \38215 );
and \U$37873 ( \38217 , \38210 , \38215 );
or \U$37874 ( \38218 , \38213 , \38216 , \38217 );
and \U$37875 ( \38219 , \38208 , \38218 );
xor \U$37876 ( \38220 , \37790 , \37800 );
xor \U$37877 ( \38221 , \38220 , \37803 );
and \U$37878 ( \38222 , \38218 , \38221 );
and \U$37879 ( \38223 , \38208 , \38221 );
or \U$37880 ( \38224 , \38219 , \38222 , \38223 );
xor \U$37881 ( \38225 , \37701 , \37753 );
xor \U$37882 ( \38226 , \38225 , \37777 );
xor \U$37883 ( \38227 , \37990 , \38011 );
xor \U$37884 ( \38228 , \38227 , \38022 );
and \U$37885 ( \38229 , \38226 , \38228 );
xor \U$37886 ( \38230 , \38027 , \38029 );
xor \U$37887 ( \38231 , \38230 , \38032 );
and \U$37888 ( \38232 , \38228 , \38231 );
and \U$37889 ( \38233 , \38226 , \38231 );
or \U$37890 ( \38234 , \38229 , \38232 , \38233 );
and \U$37891 ( \38235 , \38224 , \38234 );
xor \U$37892 ( \38236 , \37822 , \37824 );
xor \U$37893 ( \38237 , \38236 , \37827 );
and \U$37894 ( \38238 , \38234 , \38237 );
and \U$37895 ( \38239 , \38224 , \38237 );
or \U$37896 ( \38240 , \38235 , \38238 , \38239 );
xor \U$37897 ( \38241 , \37780 , \37806 );
xor \U$37898 ( \38242 , \38241 , \37817 );
xor \U$37899 ( \38243 , \38025 , \38035 );
xor \U$37900 ( \38244 , \38243 , \38038 );
and \U$37901 ( \38245 , \38242 , \38244 );
and \U$37902 ( \38246 , \38240 , \38245 );
xor \U$37903 ( \38247 , \38041 , \38043 );
xor \U$37904 ( \38248 , \38247 , \38045 );
and \U$37905 ( \38249 , \38245 , \38248 );
and \U$37906 ( \38250 , \38240 , \38248 );
or \U$37907 ( \38251 , \38246 , \38249 , \38250 );
and \U$37908 ( \38252 , \38059 , \38251 );
xor \U$37909 ( \38253 , \38059 , \38251 );
xor \U$37910 ( \38254 , \38240 , \38245 );
xor \U$37911 ( \38255 , \38254 , \38248 );
and \U$37912 ( \38256 , \23058 , \31639 );
and \U$37913 ( \38257 , \22872 , \31636 );
nor \U$37914 ( \38258 , \38256 , \38257 );
xnor \U$37915 ( \38259 , \38258 , \30584 );
and \U$37916 ( \38260 , \23466 , \30826 );
and \U$37917 ( \38261 , \23202 , \30824 );
nor \U$37918 ( \38262 , \38260 , \38261 );
xnor \U$37919 ( \38263 , \38262 , \30587 );
and \U$37920 ( \38264 , \38259 , \38263 );
and \U$37921 ( \38265 , \38263 , \22767 );
and \U$37922 ( \38266 , \38259 , \22767 );
or \U$37923 ( \38267 , \38264 , \38265 , \38266 );
and \U$37924 ( \38268 , \24836 , \28592 );
and \U$37925 ( \38269 , \24714 , \28590 );
nor \U$37926 ( \38270 , \38268 , \38269 );
xnor \U$37927 ( \38271 , \38270 , \28343 );
and \U$37928 ( \38272 , \25097 , \28063 );
and \U$37929 ( \38273 , \24841 , \28061 );
nor \U$37930 ( \38274 , \38272 , \38273 );
xnor \U$37931 ( \38275 , \38274 , \27803 );
and \U$37932 ( \38276 , \38271 , \38275 );
and \U$37933 ( \38277 , \25596 , \27569 );
and \U$37934 ( \38278 , \25294 , \27567 );
nor \U$37935 ( \38279 , \38277 , \38278 );
xnor \U$37936 ( \38280 , \38279 , \27254 );
and \U$37937 ( \38281 , \38275 , \38280 );
and \U$37938 ( \38282 , \38271 , \38280 );
or \U$37939 ( \38283 , \38276 , \38281 , \38282 );
and \U$37940 ( \38284 , \38267 , \38283 );
and \U$37941 ( \38285 , \23665 , \30258 );
and \U$37942 ( \38286 , \23491 , \30256 );
nor \U$37943 ( \38287 , \38285 , \38286 );
xnor \U$37944 ( \38288 , \38287 , \29948 );
and \U$37945 ( \38289 , \23970 , \29721 );
and \U$37946 ( \38290 , \23832 , \29719 );
nor \U$37947 ( \38291 , \38289 , \38290 );
xnor \U$37948 ( \38292 , \38291 , \29350 );
and \U$37949 ( \38293 , \38288 , \38292 );
and \U$37950 ( \38294 , \24506 , \29159 );
and \U$37951 ( \38295 , \24089 , \29157 );
nor \U$37952 ( \38296 , \38294 , \38295 );
xnor \U$37953 ( \38297 , \38296 , \28841 );
and \U$37954 ( \38298 , \38292 , \38297 );
and \U$37955 ( \38299 , \38288 , \38297 );
or \U$37956 ( \38300 , \38293 , \38298 , \38299 );
and \U$37957 ( \38301 , \38283 , \38300 );
and \U$37958 ( \38302 , \38267 , \38300 );
or \U$37959 ( \38303 , \38284 , \38301 , \38302 );
and \U$37960 ( \38304 , \30986 , \23421 );
and \U$37961 ( \38305 , \30383 , \23419 );
nor \U$37962 ( \38306 , \38304 , \38305 );
xnor \U$37963 ( \38307 , \38306 , \23279 );
and \U$37964 ( \38308 , \31172 , \23125 );
and \U$37965 ( \38309 , \30991 , \23123 );
nor \U$37966 ( \38310 , \38308 , \38309 );
xnor \U$37967 ( \38311 , \38310 , \22988 );
and \U$37968 ( \38312 , \38307 , \38311 );
nand \U$37969 ( \38313 , \31792 , \22917 );
xnor \U$37970 ( \38314 , \38313 , \22767 );
and \U$37971 ( \38315 , \38311 , \38314 );
and \U$37972 ( \38316 , \38307 , \38314 );
or \U$37973 ( \38317 , \38312 , \38315 , \38316 );
and \U$37974 ( \38318 , \30991 , \23125 );
and \U$37975 ( \38319 , \30986 , \23123 );
nor \U$37976 ( \38320 , \38318 , \38319 );
xnor \U$37977 ( \38321 , \38320 , \22988 );
and \U$37978 ( \38322 , \38317 , \38321 );
and \U$37979 ( \38323 , \31792 , \22919 );
and \U$37980 ( \38324 , \31172 , \22917 );
nor \U$37981 ( \38325 , \38323 , \38324 );
xnor \U$37982 ( \38326 , \38325 , \22767 );
and \U$37983 ( \38327 , \38321 , \38326 );
and \U$37984 ( \38328 , \38317 , \38326 );
or \U$37985 ( \38329 , \38322 , \38327 , \38328 );
and \U$37986 ( \38330 , \38303 , \38329 );
and \U$37987 ( \38331 , \26073 , \27060 );
and \U$37988 ( \38332 , \25604 , \27058 );
nor \U$37989 ( \38333 , \38331 , \38332 );
xnor \U$37990 ( \38334 , \38333 , \26720 );
and \U$37991 ( \38335 , \26342 , \26471 );
and \U$37992 ( \38336 , \26078 , \26469 );
nor \U$37993 ( \38337 , \38335 , \38336 );
xnor \U$37994 ( \38338 , \38337 , \26230 );
and \U$37995 ( \38339 , \38334 , \38338 );
and \U$37996 ( \38340 , \26973 , \26005 );
and \U$37997 ( \38341 , \26601 , \26003 );
nor \U$37998 ( \38342 , \38340 , \38341 );
xnor \U$37999 ( \38343 , \38342 , \25817 );
and \U$38000 ( \38344 , \38338 , \38343 );
and \U$38001 ( \38345 , \38334 , \38343 );
or \U$38002 ( \38346 , \38339 , \38344 , \38345 );
and \U$38003 ( \38347 , \29198 , \24462 );
and \U$38004 ( \38348 , \28952 , \24460 );
nor \U$38005 ( \38349 , \38347 , \38348 );
xnor \U$38006 ( \38350 , \38349 , \24275 );
and \U$38007 ( \38351 , \29522 , \24149 );
and \U$38008 ( \38352 , \29203 , \24147 );
nor \U$38009 ( \38353 , \38351 , \38352 );
xnor \U$38010 ( \38354 , \38353 , \23944 );
and \U$38011 ( \38355 , \38350 , \38354 );
and \U$38012 ( \38356 , \30375 , \23743 );
and \U$38013 ( \38357 , \29806 , \23741 );
nor \U$38014 ( \38358 , \38356 , \38357 );
xnor \U$38015 ( \38359 , \38358 , \23594 );
and \U$38016 ( \38360 , \38354 , \38359 );
and \U$38017 ( \38361 , \38350 , \38359 );
or \U$38018 ( \38362 , \38355 , \38360 , \38361 );
and \U$38019 ( \38363 , \38346 , \38362 );
and \U$38020 ( \38364 , \27325 , \25631 );
and \U$38021 ( \38365 , \26982 , \25629 );
nor \U$38022 ( \38366 , \38364 , \38365 );
xnor \U$38023 ( \38367 , \38366 , \25399 );
and \U$38024 ( \38368 , \27830 , \25180 );
and \U$38025 ( \38369 , \27527 , \25178 );
nor \U$38026 ( \38370 , \38368 , \38369 );
xnor \U$38027 ( \38371 , \38370 , \25037 );
and \U$38028 ( \38372 , \38367 , \38371 );
and \U$38029 ( \38373 , \28528 , \24857 );
and \U$38030 ( \38374 , \28002 , \24855 );
nor \U$38031 ( \38375 , \38373 , \38374 );
xnor \U$38032 ( \38376 , \38375 , \24611 );
and \U$38033 ( \38377 , \38371 , \38376 );
and \U$38034 ( \38378 , \38367 , \38376 );
or \U$38035 ( \38379 , \38372 , \38377 , \38378 );
and \U$38036 ( \38380 , \38362 , \38379 );
and \U$38037 ( \38381 , \38346 , \38379 );
or \U$38038 ( \38382 , \38363 , \38380 , \38381 );
and \U$38039 ( \38383 , \38329 , \38382 );
and \U$38040 ( \38384 , \38303 , \38382 );
or \U$38041 ( \38385 , \38330 , \38383 , \38384 );
xor \U$38042 ( \38386 , \38063 , \38067 );
xor \U$38043 ( \38387 , \38386 , \38072 );
xor \U$38044 ( \38388 , \38079 , \38083 );
xor \U$38045 ( \38389 , \38388 , \38088 );
and \U$38046 ( \38390 , \38387 , \38389 );
xor \U$38047 ( \38391 , \38096 , \38100 );
xor \U$38048 ( \38392 , \38391 , \38105 );
and \U$38049 ( \38393 , \38389 , \38392 );
and \U$38050 ( \38394 , \38387 , \38392 );
or \U$38051 ( \38395 , \38390 , \38393 , \38394 );
xor \U$38052 ( \38396 , \38115 , \38119 );
xor \U$38053 ( \38397 , \38396 , \38124 );
xor \U$38054 ( \38398 , \38131 , \38135 );
xor \U$38055 ( \38399 , \38398 , \38140 );
and \U$38056 ( \38400 , \38397 , \38399 );
xor \U$38057 ( \38401 , \38148 , \38152 );
xor \U$38058 ( \38402 , \38401 , \38157 );
and \U$38059 ( \38403 , \38399 , \38402 );
and \U$38060 ( \38404 , \38397 , \38402 );
or \U$38061 ( \38405 , \38400 , \38403 , \38404 );
and \U$38062 ( \38406 , \38395 , \38405 );
xor \U$38063 ( \38407 , \37882 , \37886 );
xor \U$38064 ( \38408 , \38407 , \37891 );
and \U$38065 ( \38409 , \38405 , \38408 );
and \U$38066 ( \38410 , \38395 , \38408 );
or \U$38067 ( \38411 , \38406 , \38409 , \38410 );
and \U$38068 ( \38412 , \38385 , \38411 );
xor \U$38069 ( \38413 , \37899 , \37903 );
xor \U$38070 ( \38414 , \38413 , \22495 );
xor \U$38071 ( \38415 , \38190 , \38192 );
xor \U$38072 ( \38416 , \38415 , \38195 );
and \U$38073 ( \38417 , \38414 , \38416 );
xor \U$38074 ( \38418 , \38166 , \38168 );
xor \U$38075 ( \38419 , \38418 , \38171 );
and \U$38076 ( \38420 , \38416 , \38419 );
and \U$38077 ( \38421 , \38414 , \38419 );
or \U$38078 ( \38422 , \38417 , \38420 , \38421 );
and \U$38079 ( \38423 , \38411 , \38422 );
and \U$38080 ( \38424 , \38385 , \38422 );
or \U$38081 ( \38425 , \38412 , \38423 , \38424 );
xor \U$38082 ( \38426 , \38111 , \38163 );
xor \U$38083 ( \38427 , \38426 , \38174 );
xor \U$38084 ( \38428 , \38179 , \38181 );
xor \U$38085 ( \38429 , \38428 , \38184 );
and \U$38086 ( \38430 , \38427 , \38429 );
xor \U$38087 ( \38431 , \38198 , \38200 );
xor \U$38088 ( \38432 , \38431 , \38202 );
and \U$38089 ( \38433 , \38429 , \38432 );
and \U$38090 ( \38434 , \38427 , \38432 );
or \U$38091 ( \38435 , \38430 , \38433 , \38434 );
and \U$38092 ( \38436 , \38425 , \38435 );
xor \U$38093 ( \38437 , \37910 , \37962 );
xor \U$38094 ( \38438 , \38437 , \37987 );
and \U$38095 ( \38439 , \38435 , \38438 );
and \U$38096 ( \38440 , \38425 , \38438 );
or \U$38097 ( \38441 , \38436 , \38439 , \38440 );
xor \U$38098 ( \38442 , \38177 , \38187 );
xor \U$38099 ( \38443 , \38442 , \38205 );
xor \U$38100 ( \38444 , \38210 , \38212 );
xor \U$38101 ( \38445 , \38444 , \38215 );
and \U$38102 ( \38446 , \38443 , \38445 );
and \U$38103 ( \38447 , \38441 , \38446 );
xor \U$38104 ( \38448 , \38226 , \38228 );
xor \U$38105 ( \38449 , \38448 , \38231 );
and \U$38106 ( \38450 , \38446 , \38449 );
and \U$38107 ( \38451 , \38441 , \38449 );
or \U$38108 ( \38452 , \38447 , \38450 , \38451 );
xor \U$38109 ( \38453 , \38224 , \38234 );
xor \U$38110 ( \38454 , \38453 , \38237 );
and \U$38111 ( \38455 , \38452 , \38454 );
xor \U$38112 ( \38456 , \38242 , \38244 );
and \U$38113 ( \38457 , \38454 , \38456 );
and \U$38114 ( \38458 , \38452 , \38456 );
or \U$38115 ( \38459 , \38455 , \38457 , \38458 );
and \U$38116 ( \38460 , \38255 , \38459 );
xor \U$38117 ( \38461 , \38255 , \38459 );
xor \U$38118 ( \38462 , \38452 , \38454 );
xor \U$38119 ( \38463 , \38462 , \38456 );
and \U$38120 ( \38464 , \29806 , \24149 );
and \U$38121 ( \38465 , \29522 , \24147 );
nor \U$38122 ( \38466 , \38464 , \38465 );
xnor \U$38123 ( \38467 , \38466 , \23944 );
and \U$38124 ( \38468 , \30383 , \23743 );
and \U$38125 ( \38469 , \30375 , \23741 );
nor \U$38126 ( \38470 , \38468 , \38469 );
xnor \U$38127 ( \38471 , \38470 , \23594 );
and \U$38128 ( \38472 , \38467 , \38471 );
and \U$38129 ( \38473 , \30991 , \23421 );
and \U$38130 ( \38474 , \30986 , \23419 );
nor \U$38131 ( \38475 , \38473 , \38474 );
xnor \U$38132 ( \38476 , \38475 , \23279 );
and \U$38133 ( \38477 , \38471 , \38476 );
and \U$38134 ( \38478 , \38467 , \38476 );
or \U$38135 ( \38479 , \38472 , \38477 , \38478 );
and \U$38136 ( \38480 , \26601 , \26471 );
and \U$38137 ( \38481 , \26342 , \26469 );
nor \U$38138 ( \38482 , \38480 , \38481 );
xnor \U$38139 ( \38483 , \38482 , \26230 );
and \U$38140 ( \38484 , \26982 , \26005 );
and \U$38141 ( \38485 , \26973 , \26003 );
nor \U$38142 ( \38486 , \38484 , \38485 );
xnor \U$38143 ( \38487 , \38486 , \25817 );
and \U$38144 ( \38488 , \38483 , \38487 );
and \U$38145 ( \38489 , \27527 , \25631 );
and \U$38146 ( \38490 , \27325 , \25629 );
nor \U$38147 ( \38491 , \38489 , \38490 );
xnor \U$38148 ( \38492 , \38491 , \25399 );
and \U$38149 ( \38493 , \38487 , \38492 );
and \U$38150 ( \38494 , \38483 , \38492 );
or \U$38151 ( \38495 , \38488 , \38493 , \38494 );
and \U$38152 ( \38496 , \38479 , \38495 );
and \U$38153 ( \38497 , \28002 , \25180 );
and \U$38154 ( \38498 , \27830 , \25178 );
nor \U$38155 ( \38499 , \38497 , \38498 );
xnor \U$38156 ( \38500 , \38499 , \25037 );
and \U$38157 ( \38501 , \28952 , \24857 );
and \U$38158 ( \38502 , \28528 , \24855 );
nor \U$38159 ( \38503 , \38501 , \38502 );
xnor \U$38160 ( \38504 , \38503 , \24611 );
and \U$38161 ( \38505 , \38500 , \38504 );
and \U$38162 ( \38506 , \29203 , \24462 );
and \U$38163 ( \38507 , \29198 , \24460 );
nor \U$38164 ( \38508 , \38506 , \38507 );
xnor \U$38165 ( \38509 , \38508 , \24275 );
and \U$38166 ( \38510 , \38504 , \38509 );
and \U$38167 ( \38511 , \38500 , \38509 );
or \U$38168 ( \38512 , \38505 , \38510 , \38511 );
and \U$38169 ( \38513 , \38495 , \38512 );
and \U$38170 ( \38514 , \38479 , \38512 );
or \U$38171 ( \38515 , \38496 , \38513 , \38514 );
and \U$38172 ( \38516 , \25294 , \28063 );
and \U$38173 ( \38517 , \25097 , \28061 );
nor \U$38174 ( \38518 , \38516 , \38517 );
xnor \U$38175 ( \38519 , \38518 , \27803 );
and \U$38176 ( \38520 , \25604 , \27569 );
and \U$38177 ( \38521 , \25596 , \27567 );
nor \U$38178 ( \38522 , \38520 , \38521 );
xnor \U$38179 ( \38523 , \38522 , \27254 );
and \U$38180 ( \38524 , \38519 , \38523 );
and \U$38181 ( \38525 , \26078 , \27060 );
and \U$38182 ( \38526 , \26073 , \27058 );
nor \U$38183 ( \38527 , \38525 , \38526 );
xnor \U$38184 ( \38528 , \38527 , \26720 );
and \U$38185 ( \38529 , \38523 , \38528 );
and \U$38186 ( \38530 , \38519 , \38528 );
or \U$38187 ( \38531 , \38524 , \38529 , \38530 );
and \U$38188 ( \38532 , \24089 , \29721 );
and \U$38189 ( \38533 , \23970 , \29719 );
nor \U$38190 ( \38534 , \38532 , \38533 );
xnor \U$38191 ( \38535 , \38534 , \29350 );
and \U$38192 ( \38536 , \24714 , \29159 );
and \U$38193 ( \38537 , \24506 , \29157 );
nor \U$38194 ( \38538 , \38536 , \38537 );
xnor \U$38195 ( \38539 , \38538 , \28841 );
and \U$38196 ( \38540 , \38535 , \38539 );
and \U$38197 ( \38541 , \24841 , \28592 );
and \U$38198 ( \38542 , \24836 , \28590 );
nor \U$38199 ( \38543 , \38541 , \38542 );
xnor \U$38200 ( \38544 , \38543 , \28343 );
and \U$38201 ( \38545 , \38539 , \38544 );
and \U$38202 ( \38546 , \38535 , \38544 );
or \U$38203 ( \38547 , \38540 , \38545 , \38546 );
and \U$38204 ( \38548 , \38531 , \38547 );
and \U$38205 ( \38549 , \23202 , \31639 );
and \U$38206 ( \38550 , \23058 , \31636 );
nor \U$38207 ( \38551 , \38549 , \38550 );
xnor \U$38208 ( \38552 , \38551 , \30584 );
and \U$38209 ( \38553 , \23491 , \30826 );
and \U$38210 ( \38554 , \23466 , \30824 );
nor \U$38211 ( \38555 , \38553 , \38554 );
xnor \U$38212 ( \38556 , \38555 , \30587 );
and \U$38213 ( \38557 , \38552 , \38556 );
and \U$38214 ( \38558 , \23832 , \30258 );
and \U$38215 ( \38559 , \23665 , \30256 );
nor \U$38216 ( \38560 , \38558 , \38559 );
xnor \U$38217 ( \38561 , \38560 , \29948 );
and \U$38218 ( \38562 , \38556 , \38561 );
and \U$38219 ( \38563 , \38552 , \38561 );
or \U$38220 ( \38564 , \38557 , \38562 , \38563 );
and \U$38221 ( \38565 , \38547 , \38564 );
and \U$38222 ( \38566 , \38531 , \38564 );
or \U$38223 ( \38567 , \38548 , \38565 , \38566 );
and \U$38224 ( \38568 , \38515 , \38567 );
xor \U$38225 ( \38569 , \38307 , \38311 );
xor \U$38226 ( \38570 , \38569 , \38314 );
xor \U$38227 ( \38571 , \38350 , \38354 );
xor \U$38228 ( \38572 , \38571 , \38359 );
and \U$38229 ( \38573 , \38570 , \38572 );
xor \U$38230 ( \38574 , \38367 , \38371 );
xor \U$38231 ( \38575 , \38574 , \38376 );
and \U$38232 ( \38576 , \38572 , \38575 );
and \U$38233 ( \38577 , \38570 , \38575 );
or \U$38234 ( \38578 , \38573 , \38576 , \38577 );
and \U$38235 ( \38579 , \38567 , \38578 );
and \U$38236 ( \38580 , \38515 , \38578 );
or \U$38237 ( \38581 , \38568 , \38579 , \38580 );
xor \U$38238 ( \38582 , \38267 , \38283 );
xor \U$38239 ( \38583 , \38582 , \38300 );
xor \U$38240 ( \38584 , \38317 , \38321 );
xor \U$38241 ( \38585 , \38584 , \38326 );
and \U$38242 ( \38586 , \38583 , \38585 );
xor \U$38243 ( \38587 , \38346 , \38362 );
xor \U$38244 ( \38588 , \38587 , \38379 );
and \U$38245 ( \38589 , \38585 , \38588 );
and \U$38246 ( \38590 , \38583 , \38588 );
or \U$38247 ( \38591 , \38586 , \38589 , \38590 );
and \U$38248 ( \38592 , \38581 , \38591 );
xor \U$38249 ( \38593 , \38334 , \38338 );
xor \U$38250 ( \38594 , \38593 , \38343 );
xor \U$38251 ( \38595 , \38271 , \38275 );
xor \U$38252 ( \38596 , \38595 , \38280 );
and \U$38253 ( \38597 , \38594 , \38596 );
xor \U$38254 ( \38598 , \38288 , \38292 );
xor \U$38255 ( \38599 , \38598 , \38297 );
and \U$38256 ( \38600 , \38596 , \38599 );
and \U$38257 ( \38601 , \38594 , \38599 );
or \U$38258 ( \38602 , \38597 , \38600 , \38601 );
xor \U$38259 ( \38603 , \38387 , \38389 );
xor \U$38260 ( \38604 , \38603 , \38392 );
and \U$38261 ( \38605 , \38602 , \38604 );
xor \U$38262 ( \38606 , \38397 , \38399 );
xor \U$38263 ( \38607 , \38606 , \38402 );
and \U$38264 ( \38608 , \38604 , \38607 );
and \U$38265 ( \38609 , \38602 , \38607 );
or \U$38266 ( \38610 , \38605 , \38608 , \38609 );
and \U$38267 ( \38611 , \38591 , \38610 );
and \U$38268 ( \38612 , \38581 , \38610 );
or \U$38269 ( \38613 , \38592 , \38611 , \38612 );
xor \U$38270 ( \38614 , \38075 , \38091 );
xor \U$38271 ( \38615 , \38614 , \38108 );
xor \U$38272 ( \38616 , \38127 , \38143 );
xor \U$38273 ( \38617 , \38616 , \38160 );
and \U$38274 ( \38618 , \38615 , \38617 );
xor \U$38275 ( \38619 , \38414 , \38416 );
xor \U$38276 ( \38620 , \38619 , \38419 );
and \U$38277 ( \38621 , \38617 , \38620 );
and \U$38278 ( \38622 , \38615 , \38620 );
or \U$38279 ( \38623 , \38618 , \38621 , \38622 );
and \U$38280 ( \38624 , \38613 , \38623 );
xor \U$38281 ( \38625 , \38427 , \38429 );
xor \U$38282 ( \38626 , \38625 , \38432 );
and \U$38283 ( \38627 , \38623 , \38626 );
and \U$38284 ( \38628 , \38613 , \38626 );
or \U$38285 ( \38629 , \38624 , \38627 , \38628 );
xor \U$38286 ( \38630 , \38425 , \38435 );
xor \U$38287 ( \38631 , \38630 , \38438 );
and \U$38288 ( \38632 , \38629 , \38631 );
xor \U$38289 ( \38633 , \38443 , \38445 );
and \U$38290 ( \38634 , \38631 , \38633 );
and \U$38291 ( \38635 , \38629 , \38633 );
or \U$38292 ( \38636 , \38632 , \38634 , \38635 );
xor \U$38293 ( \38637 , \38208 , \38218 );
xor \U$38294 ( \38638 , \38637 , \38221 );
and \U$38295 ( \38639 , \38636 , \38638 );
xor \U$38296 ( \38640 , \38441 , \38446 );
xor \U$38297 ( \38641 , \38640 , \38449 );
and \U$38298 ( \38642 , \38638 , \38641 );
and \U$38299 ( \38643 , \38636 , \38641 );
or \U$38300 ( \38644 , \38639 , \38642 , \38643 );
and \U$38301 ( \38645 , \38463 , \38644 );
xor \U$38302 ( \38646 , \38463 , \38644 );
xor \U$38303 ( \38647 , \38636 , \38638 );
xor \U$38304 ( \38648 , \38647 , \38641 );
and \U$38305 ( \38649 , \25097 , \28592 );
and \U$38306 ( \38650 , \24841 , \28590 );
nor \U$38307 ( \38651 , \38649 , \38650 );
xnor \U$38308 ( \38652 , \38651 , \28343 );
and \U$38309 ( \38653 , \25596 , \28063 );
and \U$38310 ( \38654 , \25294 , \28061 );
nor \U$38311 ( \38655 , \38653 , \38654 );
xnor \U$38312 ( \38656 , \38655 , \27803 );
and \U$38313 ( \38657 , \38652 , \38656 );
and \U$38314 ( \38658 , \26073 , \27569 );
and \U$38315 ( \38659 , \25604 , \27567 );
nor \U$38316 ( \38660 , \38658 , \38659 );
xnor \U$38317 ( \38661 , \38660 , \27254 );
and \U$38318 ( \38662 , \38656 , \38661 );
and \U$38319 ( \38663 , \38652 , \38661 );
or \U$38320 ( \38664 , \38657 , \38662 , \38663 );
and \U$38321 ( \38665 , \23970 , \30258 );
and \U$38322 ( \38666 , \23832 , \30256 );
nor \U$38323 ( \38667 , \38665 , \38666 );
xnor \U$38324 ( \38668 , \38667 , \29948 );
and \U$38325 ( \38669 , \24506 , \29721 );
and \U$38326 ( \38670 , \24089 , \29719 );
nor \U$38327 ( \38671 , \38669 , \38670 );
xnor \U$38328 ( \38672 , \38671 , \29350 );
and \U$38329 ( \38673 , \38668 , \38672 );
and \U$38330 ( \38674 , \24836 , \29159 );
and \U$38331 ( \38675 , \24714 , \29157 );
nor \U$38332 ( \38676 , \38674 , \38675 );
xnor \U$38333 ( \38677 , \38676 , \28841 );
and \U$38334 ( \38678 , \38672 , \38677 );
and \U$38335 ( \38679 , \38668 , \38677 );
or \U$38336 ( \38680 , \38673 , \38678 , \38679 );
and \U$38337 ( \38681 , \38664 , \38680 );
and \U$38338 ( \38682 , \23466 , \31639 );
and \U$38339 ( \38683 , \23202 , \31636 );
nor \U$38340 ( \38684 , \38682 , \38683 );
xnor \U$38341 ( \38685 , \38684 , \30584 );
and \U$38342 ( \38686 , \23665 , \30826 );
and \U$38343 ( \38687 , \23491 , \30824 );
nor \U$38344 ( \38688 , \38686 , \38687 );
xnor \U$38345 ( \38689 , \38688 , \30587 );
and \U$38346 ( \38690 , \38685 , \38689 );
and \U$38347 ( \38691 , \38689 , \22988 );
and \U$38348 ( \38692 , \38685 , \22988 );
or \U$38349 ( \38693 , \38690 , \38691 , \38692 );
and \U$38350 ( \38694 , \38680 , \38693 );
and \U$38351 ( \38695 , \38664 , \38693 );
or \U$38352 ( \38696 , \38681 , \38694 , \38695 );
and \U$38353 ( \38697 , \29522 , \24462 );
and \U$38354 ( \38698 , \29203 , \24460 );
nor \U$38355 ( \38699 , \38697 , \38698 );
xnor \U$38356 ( \38700 , \38699 , \24275 );
and \U$38357 ( \38701 , \30375 , \24149 );
and \U$38358 ( \38702 , \29806 , \24147 );
nor \U$38359 ( \38703 , \38701 , \38702 );
xnor \U$38360 ( \38704 , \38703 , \23944 );
and \U$38361 ( \38705 , \38700 , \38704 );
and \U$38362 ( \38706 , \30986 , \23743 );
and \U$38363 ( \38707 , \30383 , \23741 );
nor \U$38364 ( \38708 , \38706 , \38707 );
xnor \U$38365 ( \38709 , \38708 , \23594 );
and \U$38366 ( \38710 , \38704 , \38709 );
and \U$38367 ( \38711 , \38700 , \38709 );
or \U$38368 ( \38712 , \38705 , \38710 , \38711 );
and \U$38369 ( \38713 , \26342 , \27060 );
and \U$38370 ( \38714 , \26078 , \27058 );
nor \U$38371 ( \38715 , \38713 , \38714 );
xnor \U$38372 ( \38716 , \38715 , \26720 );
and \U$38373 ( \38717 , \26973 , \26471 );
and \U$38374 ( \38718 , \26601 , \26469 );
nor \U$38375 ( \38719 , \38717 , \38718 );
xnor \U$38376 ( \38720 , \38719 , \26230 );
and \U$38377 ( \38721 , \38716 , \38720 );
and \U$38378 ( \38722 , \27325 , \26005 );
and \U$38379 ( \38723 , \26982 , \26003 );
nor \U$38380 ( \38724 , \38722 , \38723 );
xnor \U$38381 ( \38725 , \38724 , \25817 );
and \U$38382 ( \38726 , \38720 , \38725 );
and \U$38383 ( \38727 , \38716 , \38725 );
or \U$38384 ( \38728 , \38721 , \38726 , \38727 );
and \U$38385 ( \38729 , \38712 , \38728 );
and \U$38386 ( \38730 , \27830 , \25631 );
and \U$38387 ( \38731 , \27527 , \25629 );
nor \U$38388 ( \38732 , \38730 , \38731 );
xnor \U$38389 ( \38733 , \38732 , \25399 );
and \U$38390 ( \38734 , \28528 , \25180 );
and \U$38391 ( \38735 , \28002 , \25178 );
nor \U$38392 ( \38736 , \38734 , \38735 );
xnor \U$38393 ( \38737 , \38736 , \25037 );
and \U$38394 ( \38738 , \38733 , \38737 );
and \U$38395 ( \38739 , \29198 , \24857 );
and \U$38396 ( \38740 , \28952 , \24855 );
nor \U$38397 ( \38741 , \38739 , \38740 );
xnor \U$38398 ( \38742 , \38741 , \24611 );
and \U$38399 ( \38743 , \38737 , \38742 );
and \U$38400 ( \38744 , \38733 , \38742 );
or \U$38401 ( \38745 , \38738 , \38743 , \38744 );
and \U$38402 ( \38746 , \38728 , \38745 );
and \U$38403 ( \38747 , \38712 , \38745 );
or \U$38404 ( \38748 , \38729 , \38746 , \38747 );
and \U$38405 ( \38749 , \38696 , \38748 );
and \U$38406 ( \38750 , \31792 , \23125 );
and \U$38407 ( \38751 , \31172 , \23123 );
nor \U$38408 ( \38752 , \38750 , \38751 );
xnor \U$38409 ( \38753 , \38752 , \22988 );
xor \U$38410 ( \38754 , \38467 , \38471 );
xor \U$38411 ( \38755 , \38754 , \38476 );
and \U$38412 ( \38756 , \38753 , \38755 );
xor \U$38413 ( \38757 , \38500 , \38504 );
xor \U$38414 ( \38758 , \38757 , \38509 );
and \U$38415 ( \38759 , \38755 , \38758 );
and \U$38416 ( \38760 , \38753 , \38758 );
or \U$38417 ( \38761 , \38756 , \38759 , \38760 );
and \U$38418 ( \38762 , \38748 , \38761 );
and \U$38419 ( \38763 , \38696 , \38761 );
or \U$38420 ( \38764 , \38749 , \38762 , \38763 );
xor \U$38421 ( \38765 , \38519 , \38523 );
xor \U$38422 ( \38766 , \38765 , \38528 );
xor \U$38423 ( \38767 , \38483 , \38487 );
xor \U$38424 ( \38768 , \38767 , \38492 );
and \U$38425 ( \38769 , \38766 , \38768 );
xor \U$38426 ( \38770 , \38535 , \38539 );
xor \U$38427 ( \38771 , \38770 , \38544 );
and \U$38428 ( \38772 , \38768 , \38771 );
and \U$38429 ( \38773 , \38766 , \38771 );
or \U$38430 ( \38774 , \38769 , \38772 , \38773 );
xor \U$38431 ( \38775 , \38259 , \38263 );
xor \U$38432 ( \38776 , \38775 , \22767 );
and \U$38433 ( \38777 , \38774 , \38776 );
xor \U$38434 ( \38778 , \38594 , \38596 );
xor \U$38435 ( \38779 , \38778 , \38599 );
and \U$38436 ( \38780 , \38776 , \38779 );
and \U$38437 ( \38781 , \38774 , \38779 );
or \U$38438 ( \38782 , \38777 , \38780 , \38781 );
and \U$38439 ( \38783 , \38764 , \38782 );
xor \U$38440 ( \38784 , \38479 , \38495 );
xor \U$38441 ( \38785 , \38784 , \38512 );
xor \U$38442 ( \38786 , \38531 , \38547 );
xor \U$38443 ( \38787 , \38786 , \38564 );
and \U$38444 ( \38788 , \38785 , \38787 );
xor \U$38445 ( \38789 , \38570 , \38572 );
xor \U$38446 ( \38790 , \38789 , \38575 );
and \U$38447 ( \38791 , \38787 , \38790 );
and \U$38448 ( \38792 , \38785 , \38790 );
or \U$38449 ( \38793 , \38788 , \38791 , \38792 );
and \U$38450 ( \38794 , \38782 , \38793 );
and \U$38451 ( \38795 , \38764 , \38793 );
or \U$38452 ( \38796 , \38783 , \38794 , \38795 );
xor \U$38453 ( \38797 , \38515 , \38567 );
xor \U$38454 ( \38798 , \38797 , \38578 );
xor \U$38455 ( \38799 , \38583 , \38585 );
xor \U$38456 ( \38800 , \38799 , \38588 );
and \U$38457 ( \38801 , \38798 , \38800 );
xor \U$38458 ( \38802 , \38602 , \38604 );
xor \U$38459 ( \38803 , \38802 , \38607 );
and \U$38460 ( \38804 , \38800 , \38803 );
and \U$38461 ( \38805 , \38798 , \38803 );
or \U$38462 ( \38806 , \38801 , \38804 , \38805 );
and \U$38463 ( \38807 , \38796 , \38806 );
xor \U$38464 ( \38808 , \38395 , \38405 );
xor \U$38465 ( \38809 , \38808 , \38408 );
and \U$38466 ( \38810 , \38806 , \38809 );
and \U$38467 ( \38811 , \38796 , \38809 );
or \U$38468 ( \38812 , \38807 , \38810 , \38811 );
xor \U$38469 ( \38813 , \38303 , \38329 );
xor \U$38470 ( \38814 , \38813 , \38382 );
xor \U$38471 ( \38815 , \38581 , \38591 );
xor \U$38472 ( \38816 , \38815 , \38610 );
and \U$38473 ( \38817 , \38814 , \38816 );
xor \U$38474 ( \38818 , \38615 , \38617 );
xor \U$38475 ( \38819 , \38818 , \38620 );
and \U$38476 ( \38820 , \38816 , \38819 );
and \U$38477 ( \38821 , \38814 , \38819 );
or \U$38478 ( \38822 , \38817 , \38820 , \38821 );
and \U$38479 ( \38823 , \38812 , \38822 );
xor \U$38480 ( \38824 , \38385 , \38411 );
xor \U$38481 ( \38825 , \38824 , \38422 );
and \U$38482 ( \38826 , \38822 , \38825 );
and \U$38483 ( \38827 , \38812 , \38825 );
or \U$38484 ( \38828 , \38823 , \38826 , \38827 );
xor \U$38485 ( \38829 , \38629 , \38631 );
xor \U$38486 ( \38830 , \38829 , \38633 );
and \U$38487 ( \38831 , \38828 , \38830 );
and \U$38488 ( \38832 , \38648 , \38831 );
xor \U$38489 ( \38833 , \38648 , \38831 );
xor \U$38490 ( \38834 , \38828 , \38830 );
and \U$38491 ( \38835 , \23491 , \31639 );
and \U$38492 ( \38836 , \23466 , \31636 );
nor \U$38493 ( \38837 , \38835 , \38836 );
xnor \U$38494 ( \38838 , \38837 , \30584 );
and \U$38495 ( \38839 , \23832 , \30826 );
and \U$38496 ( \38840 , \23665 , \30824 );
nor \U$38497 ( \38841 , \38839 , \38840 );
xnor \U$38498 ( \38842 , \38841 , \30587 );
and \U$38499 ( \38843 , \38838 , \38842 );
and \U$38500 ( \38844 , \24089 , \30258 );
and \U$38501 ( \38845 , \23970 , \30256 );
nor \U$38502 ( \38846 , \38844 , \38845 );
xnor \U$38503 ( \38847 , \38846 , \29948 );
and \U$38504 ( \38848 , \38842 , \38847 );
and \U$38505 ( \38849 , \38838 , \38847 );
or \U$38506 ( \38850 , \38843 , \38848 , \38849 );
and \U$38507 ( \38851 , \24714 , \29721 );
and \U$38508 ( \38852 , \24506 , \29719 );
nor \U$38509 ( \38853 , \38851 , \38852 );
xnor \U$38510 ( \38854 , \38853 , \29350 );
and \U$38511 ( \38855 , \24841 , \29159 );
and \U$38512 ( \38856 , \24836 , \29157 );
nor \U$38513 ( \38857 , \38855 , \38856 );
xnor \U$38514 ( \38858 , \38857 , \28841 );
and \U$38515 ( \38859 , \38854 , \38858 );
and \U$38516 ( \38860 , \25294 , \28592 );
and \U$38517 ( \38861 , \25097 , \28590 );
nor \U$38518 ( \38862 , \38860 , \38861 );
xnor \U$38519 ( \38863 , \38862 , \28343 );
and \U$38520 ( \38864 , \38858 , \38863 );
and \U$38521 ( \38865 , \38854 , \38863 );
or \U$38522 ( \38866 , \38859 , \38864 , \38865 );
and \U$38523 ( \38867 , \38850 , \38866 );
and \U$38524 ( \38868 , \25604 , \28063 );
and \U$38525 ( \38869 , \25596 , \28061 );
nor \U$38526 ( \38870 , \38868 , \38869 );
xnor \U$38527 ( \38871 , \38870 , \27803 );
and \U$38528 ( \38872 , \26078 , \27569 );
and \U$38529 ( \38873 , \26073 , \27567 );
nor \U$38530 ( \38874 , \38872 , \38873 );
xnor \U$38531 ( \38875 , \38874 , \27254 );
and \U$38532 ( \38876 , \38871 , \38875 );
and \U$38533 ( \38877 , \26601 , \27060 );
and \U$38534 ( \38878 , \26342 , \27058 );
nor \U$38535 ( \38879 , \38877 , \38878 );
xnor \U$38536 ( \38880 , \38879 , \26720 );
and \U$38537 ( \38881 , \38875 , \38880 );
and \U$38538 ( \38882 , \38871 , \38880 );
or \U$38539 ( \38883 , \38876 , \38881 , \38882 );
and \U$38540 ( \38884 , \38866 , \38883 );
and \U$38541 ( \38885 , \38850 , \38883 );
or \U$38542 ( \38886 , \38867 , \38884 , \38885 );
and \U$38543 ( \38887 , \30383 , \24149 );
and \U$38544 ( \38888 , \30375 , \24147 );
nor \U$38545 ( \38889 , \38887 , \38888 );
xnor \U$38546 ( \38890 , \38889 , \23944 );
and \U$38547 ( \38891 , \30991 , \23743 );
and \U$38548 ( \38892 , \30986 , \23741 );
nor \U$38549 ( \38893 , \38891 , \38892 );
xnor \U$38550 ( \38894 , \38893 , \23594 );
and \U$38551 ( \38895 , \38890 , \38894 );
and \U$38552 ( \38896 , \31792 , \23421 );
and \U$38553 ( \38897 , \31172 , \23419 );
nor \U$38554 ( \38898 , \38896 , \38897 );
xnor \U$38555 ( \38899 , \38898 , \23279 );
and \U$38556 ( \38900 , \38894 , \38899 );
and \U$38557 ( \38901 , \38890 , \38899 );
or \U$38558 ( \38902 , \38895 , \38900 , \38901 );
and \U$38559 ( \38903 , \28952 , \25180 );
and \U$38560 ( \38904 , \28528 , \25178 );
nor \U$38561 ( \38905 , \38903 , \38904 );
xnor \U$38562 ( \38906 , \38905 , \25037 );
and \U$38563 ( \38907 , \29203 , \24857 );
and \U$38564 ( \38908 , \29198 , \24855 );
nor \U$38565 ( \38909 , \38907 , \38908 );
xnor \U$38566 ( \38910 , \38909 , \24611 );
and \U$38567 ( \38911 , \38906 , \38910 );
and \U$38568 ( \38912 , \29806 , \24462 );
and \U$38569 ( \38913 , \29522 , \24460 );
nor \U$38570 ( \38914 , \38912 , \38913 );
xnor \U$38571 ( \38915 , \38914 , \24275 );
and \U$38572 ( \38916 , \38910 , \38915 );
and \U$38573 ( \38917 , \38906 , \38915 );
or \U$38574 ( \38918 , \38911 , \38916 , \38917 );
and \U$38575 ( \38919 , \38902 , \38918 );
and \U$38576 ( \38920 , \26982 , \26471 );
and \U$38577 ( \38921 , \26973 , \26469 );
nor \U$38578 ( \38922 , \38920 , \38921 );
xnor \U$38579 ( \38923 , \38922 , \26230 );
and \U$38580 ( \38924 , \27527 , \26005 );
and \U$38581 ( \38925 , \27325 , \26003 );
nor \U$38582 ( \38926 , \38924 , \38925 );
xnor \U$38583 ( \38927 , \38926 , \25817 );
and \U$38584 ( \38928 , \38923 , \38927 );
and \U$38585 ( \38929 , \28002 , \25631 );
and \U$38586 ( \38930 , \27830 , \25629 );
nor \U$38587 ( \38931 , \38929 , \38930 );
xnor \U$38588 ( \38932 , \38931 , \25399 );
and \U$38589 ( \38933 , \38927 , \38932 );
and \U$38590 ( \38934 , \38923 , \38932 );
or \U$38591 ( \38935 , \38928 , \38933 , \38934 );
and \U$38592 ( \38936 , \38918 , \38935 );
and \U$38593 ( \38937 , \38902 , \38935 );
or \U$38594 ( \38938 , \38919 , \38936 , \38937 );
and \U$38595 ( \38939 , \38886 , \38938 );
and \U$38596 ( \38940 , \31172 , \23421 );
and \U$38597 ( \38941 , \30991 , \23419 );
nor \U$38598 ( \38942 , \38940 , \38941 );
xnor \U$38599 ( \38943 , \38942 , \23279 );
nand \U$38600 ( \38944 , \31792 , \23123 );
xnor \U$38601 ( \38945 , \38944 , \22988 );
and \U$38602 ( \38946 , \38943 , \38945 );
xor \U$38603 ( \38947 , \38700 , \38704 );
xor \U$38604 ( \38948 , \38947 , \38709 );
and \U$38605 ( \38949 , \38945 , \38948 );
and \U$38606 ( \38950 , \38943 , \38948 );
or \U$38607 ( \38951 , \38946 , \38949 , \38950 );
and \U$38608 ( \38952 , \38938 , \38951 );
and \U$38609 ( \38953 , \38886 , \38951 );
or \U$38610 ( \38954 , \38939 , \38952 , \38953 );
xor \U$38611 ( \38955 , \38652 , \38656 );
xor \U$38612 ( \38956 , \38955 , \38661 );
xor \U$38613 ( \38957 , \38716 , \38720 );
xor \U$38614 ( \38958 , \38957 , \38725 );
and \U$38615 ( \38959 , \38956 , \38958 );
xor \U$38616 ( \38960 , \38733 , \38737 );
xor \U$38617 ( \38961 , \38960 , \38742 );
and \U$38618 ( \38962 , \38958 , \38961 );
and \U$38619 ( \38963 , \38956 , \38961 );
or \U$38620 ( \38964 , \38959 , \38962 , \38963 );
xor \U$38621 ( \38965 , \38668 , \38672 );
xor \U$38622 ( \38966 , \38965 , \38677 );
xor \U$38623 ( \38967 , \38685 , \38689 );
xor \U$38624 ( \38968 , \38967 , \22988 );
and \U$38625 ( \38969 , \38966 , \38968 );
and \U$38626 ( \38970 , \38964 , \38969 );
xor \U$38627 ( \38971 , \38552 , \38556 );
xor \U$38628 ( \38972 , \38971 , \38561 );
and \U$38629 ( \38973 , \38969 , \38972 );
and \U$38630 ( \38974 , \38964 , \38972 );
or \U$38631 ( \38975 , \38970 , \38973 , \38974 );
and \U$38632 ( \38976 , \38954 , \38975 );
xor \U$38633 ( \38977 , \38712 , \38728 );
xor \U$38634 ( \38978 , \38977 , \38745 );
xor \U$38635 ( \38979 , \38766 , \38768 );
xor \U$38636 ( \38980 , \38979 , \38771 );
and \U$38637 ( \38981 , \38978 , \38980 );
xor \U$38638 ( \38982 , \38753 , \38755 );
xor \U$38639 ( \38983 , \38982 , \38758 );
and \U$38640 ( \38984 , \38980 , \38983 );
and \U$38641 ( \38985 , \38978 , \38983 );
or \U$38642 ( \38986 , \38981 , \38984 , \38985 );
and \U$38643 ( \38987 , \38975 , \38986 );
and \U$38644 ( \38988 , \38954 , \38986 );
or \U$38645 ( \38989 , \38976 , \38987 , \38988 );
xor \U$38646 ( \38990 , \38696 , \38748 );
xor \U$38647 ( \38991 , \38990 , \38761 );
xor \U$38648 ( \38992 , \38774 , \38776 );
xor \U$38649 ( \38993 , \38992 , \38779 );
and \U$38650 ( \38994 , \38991 , \38993 );
xor \U$38651 ( \38995 , \38785 , \38787 );
xor \U$38652 ( \38996 , \38995 , \38790 );
and \U$38653 ( \38997 , \38993 , \38996 );
and \U$38654 ( \38998 , \38991 , \38996 );
or \U$38655 ( \38999 , \38994 , \38997 , \38998 );
and \U$38656 ( \39000 , \38989 , \38999 );
xor \U$38657 ( \39001 , \38798 , \38800 );
xor \U$38658 ( \39002 , \39001 , \38803 );
and \U$38659 ( \39003 , \38999 , \39002 );
and \U$38660 ( \39004 , \38989 , \39002 );
or \U$38661 ( \39005 , \39000 , \39003 , \39004 );
xor \U$38662 ( \39006 , \38796 , \38806 );
xor \U$38663 ( \39007 , \39006 , \38809 );
and \U$38664 ( \39008 , \39005 , \39007 );
xor \U$38665 ( \39009 , \38814 , \38816 );
xor \U$38666 ( \39010 , \39009 , \38819 );
and \U$38667 ( \39011 , \39007 , \39010 );
and \U$38668 ( \39012 , \39005 , \39010 );
or \U$38669 ( \39013 , \39008 , \39011 , \39012 );
xor \U$38670 ( \39014 , \38812 , \38822 );
xor \U$38671 ( \39015 , \39014 , \38825 );
and \U$38672 ( \39016 , \39013 , \39015 );
xor \U$38673 ( \39017 , \38613 , \38623 );
xor \U$38674 ( \39018 , \39017 , \38626 );
and \U$38675 ( \39019 , \39015 , \39018 );
and \U$38676 ( \39020 , \39013 , \39018 );
or \U$38677 ( \39021 , \39016 , \39019 , \39020 );
and \U$38678 ( \39022 , \38834 , \39021 );
xor \U$38679 ( \39023 , \38834 , \39021 );
xor \U$38680 ( \39024 , \39013 , \39015 );
xor \U$38681 ( \39025 , \39024 , \39018 );
and \U$38682 ( \39026 , \23665 , \31639 );
and \U$38683 ( \39027 , \23491 , \31636 );
nor \U$38684 ( \39028 , \39026 , \39027 );
xnor \U$38685 ( \39029 , \39028 , \30584 );
and \U$38686 ( \39030 , \23970 , \30826 );
and \U$38687 ( \39031 , \23832 , \30824 );
nor \U$38688 ( \39032 , \39030 , \39031 );
xnor \U$38689 ( \39033 , \39032 , \30587 );
and \U$38690 ( \39034 , \39029 , \39033 );
and \U$38691 ( \39035 , \39033 , \23279 );
and \U$38692 ( \39036 , \39029 , \23279 );
or \U$38693 ( \39037 , \39034 , \39035 , \39036 );
and \U$38694 ( \39038 , \24506 , \30258 );
and \U$38695 ( \39039 , \24089 , \30256 );
nor \U$38696 ( \39040 , \39038 , \39039 );
xnor \U$38697 ( \39041 , \39040 , \29948 );
and \U$38698 ( \39042 , \24836 , \29721 );
and \U$38699 ( \39043 , \24714 , \29719 );
nor \U$38700 ( \39044 , \39042 , \39043 );
xnor \U$38701 ( \39045 , \39044 , \29350 );
and \U$38702 ( \39046 , \39041 , \39045 );
and \U$38703 ( \39047 , \25097 , \29159 );
and \U$38704 ( \39048 , \24841 , \29157 );
nor \U$38705 ( \39049 , \39047 , \39048 );
xnor \U$38706 ( \39050 , \39049 , \28841 );
and \U$38707 ( \39051 , \39045 , \39050 );
and \U$38708 ( \39052 , \39041 , \39050 );
or \U$38709 ( \39053 , \39046 , \39051 , \39052 );
and \U$38710 ( \39054 , \39037 , \39053 );
and \U$38711 ( \39055 , \25596 , \28592 );
and \U$38712 ( \39056 , \25294 , \28590 );
nor \U$38713 ( \39057 , \39055 , \39056 );
xnor \U$38714 ( \39058 , \39057 , \28343 );
and \U$38715 ( \39059 , \26073 , \28063 );
and \U$38716 ( \39060 , \25604 , \28061 );
nor \U$38717 ( \39061 , \39059 , \39060 );
xnor \U$38718 ( \39062 , \39061 , \27803 );
and \U$38719 ( \39063 , \39058 , \39062 );
and \U$38720 ( \39064 , \26342 , \27569 );
and \U$38721 ( \39065 , \26078 , \27567 );
nor \U$38722 ( \39066 , \39064 , \39065 );
xnor \U$38723 ( \39067 , \39066 , \27254 );
and \U$38724 ( \39068 , \39062 , \39067 );
and \U$38725 ( \39069 , \39058 , \39067 );
or \U$38726 ( \39070 , \39063 , \39068 , \39069 );
and \U$38727 ( \39071 , \39053 , \39070 );
and \U$38728 ( \39072 , \39037 , \39070 );
or \U$38729 ( \39073 , \39054 , \39071 , \39072 );
and \U$38730 ( \39074 , \26973 , \27060 );
and \U$38731 ( \39075 , \26601 , \27058 );
nor \U$38732 ( \39076 , \39074 , \39075 );
xnor \U$38733 ( \39077 , \39076 , \26720 );
and \U$38734 ( \39078 , \27325 , \26471 );
and \U$38735 ( \39079 , \26982 , \26469 );
nor \U$38736 ( \39080 , \39078 , \39079 );
xnor \U$38737 ( \39081 , \39080 , \26230 );
and \U$38738 ( \39082 , \39077 , \39081 );
and \U$38739 ( \39083 , \27830 , \26005 );
and \U$38740 ( \39084 , \27527 , \26003 );
nor \U$38741 ( \39085 , \39083 , \39084 );
xnor \U$38742 ( \39086 , \39085 , \25817 );
and \U$38743 ( \39087 , \39081 , \39086 );
and \U$38744 ( \39088 , \39077 , \39086 );
or \U$38745 ( \39089 , \39082 , \39087 , \39088 );
and \U$38746 ( \39090 , \28528 , \25631 );
and \U$38747 ( \39091 , \28002 , \25629 );
nor \U$38748 ( \39092 , \39090 , \39091 );
xnor \U$38749 ( \39093 , \39092 , \25399 );
and \U$38750 ( \39094 , \29198 , \25180 );
and \U$38751 ( \39095 , \28952 , \25178 );
nor \U$38752 ( \39096 , \39094 , \39095 );
xnor \U$38753 ( \39097 , \39096 , \25037 );
and \U$38754 ( \39098 , \39093 , \39097 );
and \U$38755 ( \39099 , \29522 , \24857 );
and \U$38756 ( \39100 , \29203 , \24855 );
nor \U$38757 ( \39101 , \39099 , \39100 );
xnor \U$38758 ( \39102 , \39101 , \24611 );
and \U$38759 ( \39103 , \39097 , \39102 );
and \U$38760 ( \39104 , \39093 , \39102 );
or \U$38761 ( \39105 , \39098 , \39103 , \39104 );
and \U$38762 ( \39106 , \39089 , \39105 );
and \U$38763 ( \39107 , \30375 , \24462 );
and \U$38764 ( \39108 , \29806 , \24460 );
nor \U$38765 ( \39109 , \39107 , \39108 );
xnor \U$38766 ( \39110 , \39109 , \24275 );
and \U$38767 ( \39111 , \30986 , \24149 );
and \U$38768 ( \39112 , \30383 , \24147 );
nor \U$38769 ( \39113 , \39111 , \39112 );
xnor \U$38770 ( \39114 , \39113 , \23944 );
and \U$38771 ( \39115 , \39110 , \39114 );
and \U$38772 ( \39116 , \31172 , \23743 );
and \U$38773 ( \39117 , \30991 , \23741 );
nor \U$38774 ( \39118 , \39116 , \39117 );
xnor \U$38775 ( \39119 , \39118 , \23594 );
and \U$38776 ( \39120 , \39114 , \39119 );
and \U$38777 ( \39121 , \39110 , \39119 );
or \U$38778 ( \39122 , \39115 , \39120 , \39121 );
and \U$38779 ( \39123 , \39105 , \39122 );
and \U$38780 ( \39124 , \39089 , \39122 );
or \U$38781 ( \39125 , \39106 , \39123 , \39124 );
and \U$38782 ( \39126 , \39073 , \39125 );
xor \U$38783 ( \39127 , \38890 , \38894 );
xor \U$38784 ( \39128 , \39127 , \38899 );
xor \U$38785 ( \39129 , \38906 , \38910 );
xor \U$38786 ( \39130 , \39129 , \38915 );
and \U$38787 ( \39131 , \39128 , \39130 );
xor \U$38788 ( \39132 , \38923 , \38927 );
xor \U$38789 ( \39133 , \39132 , \38932 );
and \U$38790 ( \39134 , \39130 , \39133 );
and \U$38791 ( \39135 , \39128 , \39133 );
or \U$38792 ( \39136 , \39131 , \39134 , \39135 );
and \U$38793 ( \39137 , \39125 , \39136 );
and \U$38794 ( \39138 , \39073 , \39136 );
or \U$38795 ( \39139 , \39126 , \39137 , \39138 );
xor \U$38796 ( \39140 , \38850 , \38866 );
xor \U$38797 ( \39141 , \39140 , \38883 );
xor \U$38798 ( \39142 , \38902 , \38918 );
xor \U$38799 ( \39143 , \39142 , \38935 );
and \U$38800 ( \39144 , \39141 , \39143 );
xor \U$38801 ( \39145 , \38943 , \38945 );
xor \U$38802 ( \39146 , \39145 , \38948 );
and \U$38803 ( \39147 , \39143 , \39146 );
and \U$38804 ( \39148 , \39141 , \39146 );
or \U$38805 ( \39149 , \39144 , \39147 , \39148 );
and \U$38806 ( \39150 , \39139 , \39149 );
xor \U$38807 ( \39151 , \38838 , \38842 );
xor \U$38808 ( \39152 , \39151 , \38847 );
xor \U$38809 ( \39153 , \38854 , \38858 );
xor \U$38810 ( \39154 , \39153 , \38863 );
and \U$38811 ( \39155 , \39152 , \39154 );
xor \U$38812 ( \39156 , \38871 , \38875 );
xor \U$38813 ( \39157 , \39156 , \38880 );
and \U$38814 ( \39158 , \39154 , \39157 );
and \U$38815 ( \39159 , \39152 , \39157 );
or \U$38816 ( \39160 , \39155 , \39158 , \39159 );
xor \U$38817 ( \39161 , \38956 , \38958 );
xor \U$38818 ( \39162 , \39161 , \38961 );
and \U$38819 ( \39163 , \39160 , \39162 );
xor \U$38820 ( \39164 , \38966 , \38968 );
and \U$38821 ( \39165 , \39162 , \39164 );
and \U$38822 ( \39166 , \39160 , \39164 );
or \U$38823 ( \39167 , \39163 , \39165 , \39166 );
and \U$38824 ( \39168 , \39149 , \39167 );
and \U$38825 ( \39169 , \39139 , \39167 );
or \U$38826 ( \39170 , \39150 , \39168 , \39169 );
xor \U$38827 ( \39171 , \38664 , \38680 );
xor \U$38828 ( \39172 , \39171 , \38693 );
xor \U$38829 ( \39173 , \38964 , \38969 );
xor \U$38830 ( \39174 , \39173 , \38972 );
and \U$38831 ( \39175 , \39172 , \39174 );
xor \U$38832 ( \39176 , \38978 , \38980 );
xor \U$38833 ( \39177 , \39176 , \38983 );
and \U$38834 ( \39178 , \39174 , \39177 );
and \U$38835 ( \39179 , \39172 , \39177 );
or \U$38836 ( \39180 , \39175 , \39178 , \39179 );
and \U$38837 ( \39181 , \39170 , \39180 );
xor \U$38838 ( \39182 , \38991 , \38993 );
xor \U$38839 ( \39183 , \39182 , \38996 );
and \U$38840 ( \39184 , \39180 , \39183 );
and \U$38841 ( \39185 , \39170 , \39183 );
or \U$38842 ( \39186 , \39181 , \39184 , \39185 );
xor \U$38843 ( \39187 , \38764 , \38782 );
xor \U$38844 ( \39188 , \39187 , \38793 );
and \U$38845 ( \39189 , \39186 , \39188 );
xor \U$38846 ( \39190 , \38989 , \38999 );
xor \U$38847 ( \39191 , \39190 , \39002 );
and \U$38848 ( \39192 , \39188 , \39191 );
and \U$38849 ( \39193 , \39186 , \39191 );
or \U$38850 ( \39194 , \39189 , \39192 , \39193 );
xor \U$38851 ( \39195 , \39005 , \39007 );
xor \U$38852 ( \39196 , \39195 , \39010 );
and \U$38853 ( \39197 , \39194 , \39196 );
and \U$38854 ( \39198 , \39025 , \39197 );
xor \U$38855 ( \39199 , \39025 , \39197 );
xor \U$38856 ( \39200 , \39194 , \39196 );
and \U$38857 ( \39201 , \26078 , \28063 );
and \U$38858 ( \39202 , \26073 , \28061 );
nor \U$38859 ( \39203 , \39201 , \39202 );
xnor \U$38860 ( \39204 , \39203 , \27803 );
and \U$38861 ( \39205 , \26601 , \27569 );
and \U$38862 ( \39206 , \26342 , \27567 );
nor \U$38863 ( \39207 , \39205 , \39206 );
xnor \U$38864 ( \39208 , \39207 , \27254 );
and \U$38865 ( \39209 , \39204 , \39208 );
and \U$38866 ( \39210 , \26982 , \27060 );
and \U$38867 ( \39211 , \26973 , \27058 );
nor \U$38868 ( \39212 , \39210 , \39211 );
xnor \U$38869 ( \39213 , \39212 , \26720 );
and \U$38870 ( \39214 , \39208 , \39213 );
and \U$38871 ( \39215 , \39204 , \39213 );
or \U$38872 ( \39216 , \39209 , \39214 , \39215 );
and \U$38873 ( \39217 , \23832 , \31639 );
and \U$38874 ( \39218 , \23665 , \31636 );
nor \U$38875 ( \39219 , \39217 , \39218 );
xnor \U$38876 ( \39220 , \39219 , \30584 );
and \U$38877 ( \39221 , \24089 , \30826 );
and \U$38878 ( \39222 , \23970 , \30824 );
nor \U$38879 ( \39223 , \39221 , \39222 );
xnor \U$38880 ( \39224 , \39223 , \30587 );
and \U$38881 ( \39225 , \39220 , \39224 );
and \U$38882 ( \39226 , \24714 , \30258 );
and \U$38883 ( \39227 , \24506 , \30256 );
nor \U$38884 ( \39228 , \39226 , \39227 );
xnor \U$38885 ( \39229 , \39228 , \29948 );
and \U$38886 ( \39230 , \39224 , \39229 );
and \U$38887 ( \39231 , \39220 , \39229 );
or \U$38888 ( \39232 , \39225 , \39230 , \39231 );
and \U$38889 ( \39233 , \39216 , \39232 );
and \U$38890 ( \39234 , \24841 , \29721 );
and \U$38891 ( \39235 , \24836 , \29719 );
nor \U$38892 ( \39236 , \39234 , \39235 );
xnor \U$38893 ( \39237 , \39236 , \29350 );
and \U$38894 ( \39238 , \25294 , \29159 );
and \U$38895 ( \39239 , \25097 , \29157 );
nor \U$38896 ( \39240 , \39238 , \39239 );
xnor \U$38897 ( \39241 , \39240 , \28841 );
and \U$38898 ( \39242 , \39237 , \39241 );
and \U$38899 ( \39243 , \25604 , \28592 );
and \U$38900 ( \39244 , \25596 , \28590 );
nor \U$38901 ( \39245 , \39243 , \39244 );
xnor \U$38902 ( \39246 , \39245 , \28343 );
and \U$38903 ( \39247 , \39241 , \39246 );
and \U$38904 ( \39248 , \39237 , \39246 );
or \U$38905 ( \39249 , \39242 , \39247 , \39248 );
and \U$38906 ( \39250 , \39232 , \39249 );
and \U$38907 ( \39251 , \39216 , \39249 );
or \U$38908 ( \39252 , \39233 , \39250 , \39251 );
and \U$38909 ( \39253 , \29203 , \25180 );
and \U$38910 ( \39254 , \29198 , \25178 );
nor \U$38911 ( \39255 , \39253 , \39254 );
xnor \U$38912 ( \39256 , \39255 , \25037 );
and \U$38913 ( \39257 , \29806 , \24857 );
and \U$38914 ( \39258 , \29522 , \24855 );
nor \U$38915 ( \39259 , \39257 , \39258 );
xnor \U$38916 ( \39260 , \39259 , \24611 );
and \U$38917 ( \39261 , \39256 , \39260 );
and \U$38918 ( \39262 , \30383 , \24462 );
and \U$38919 ( \39263 , \30375 , \24460 );
nor \U$38920 ( \39264 , \39262 , \39263 );
xnor \U$38921 ( \39265 , \39264 , \24275 );
and \U$38922 ( \39266 , \39260 , \39265 );
and \U$38923 ( \39267 , \39256 , \39265 );
or \U$38924 ( \39268 , \39261 , \39266 , \39267 );
and \U$38925 ( \39269 , \27527 , \26471 );
and \U$38926 ( \39270 , \27325 , \26469 );
nor \U$38927 ( \39271 , \39269 , \39270 );
xnor \U$38928 ( \39272 , \39271 , \26230 );
and \U$38929 ( \39273 , \28002 , \26005 );
and \U$38930 ( \39274 , \27830 , \26003 );
nor \U$38931 ( \39275 , \39273 , \39274 );
xnor \U$38932 ( \39276 , \39275 , \25817 );
and \U$38933 ( \39277 , \39272 , \39276 );
and \U$38934 ( \39278 , \28952 , \25631 );
and \U$38935 ( \39279 , \28528 , \25629 );
nor \U$38936 ( \39280 , \39278 , \39279 );
xnor \U$38937 ( \39281 , \39280 , \25399 );
and \U$38938 ( \39282 , \39276 , \39281 );
and \U$38939 ( \39283 , \39272 , \39281 );
or \U$38940 ( \39284 , \39277 , \39282 , \39283 );
and \U$38941 ( \39285 , \39268 , \39284 );
and \U$38942 ( \39286 , \30991 , \24149 );
and \U$38943 ( \39287 , \30986 , \24147 );
nor \U$38944 ( \39288 , \39286 , \39287 );
xnor \U$38945 ( \39289 , \39288 , \23944 );
and \U$38946 ( \39290 , \31792 , \23743 );
and \U$38947 ( \39291 , \31172 , \23741 );
nor \U$38948 ( \39292 , \39290 , \39291 );
xnor \U$38949 ( \39293 , \39292 , \23594 );
and \U$38950 ( \39294 , \39289 , \39293 );
and \U$38951 ( \39295 , \39284 , \39294 );
and \U$38952 ( \39296 , \39268 , \39294 );
or \U$38953 ( \39297 , \39285 , \39295 , \39296 );
and \U$38954 ( \39298 , \39252 , \39297 );
nand \U$38955 ( \39299 , \31792 , \23419 );
xnor \U$38956 ( \39300 , \39299 , \23279 );
xor \U$38957 ( \39301 , \39093 , \39097 );
xor \U$38958 ( \39302 , \39301 , \39102 );
and \U$38959 ( \39303 , \39300 , \39302 );
xor \U$38960 ( \39304 , \39110 , \39114 );
xor \U$38961 ( \39305 , \39304 , \39119 );
and \U$38962 ( \39306 , \39302 , \39305 );
and \U$38963 ( \39307 , \39300 , \39305 );
or \U$38964 ( \39308 , \39303 , \39306 , \39307 );
and \U$38965 ( \39309 , \39297 , \39308 );
and \U$38966 ( \39310 , \39252 , \39308 );
or \U$38967 ( \39311 , \39298 , \39309 , \39310 );
xor \U$38968 ( \39312 , \39041 , \39045 );
xor \U$38969 ( \39313 , \39312 , \39050 );
xor \U$38970 ( \39314 , \39077 , \39081 );
xor \U$38971 ( \39315 , \39314 , \39086 );
and \U$38972 ( \39316 , \39313 , \39315 );
xor \U$38973 ( \39317 , \39058 , \39062 );
xor \U$38974 ( \39318 , \39317 , \39067 );
and \U$38975 ( \39319 , \39315 , \39318 );
and \U$38976 ( \39320 , \39313 , \39318 );
or \U$38977 ( \39321 , \39316 , \39319 , \39320 );
xor \U$38978 ( \39322 , \39128 , \39130 );
xor \U$38979 ( \39323 , \39322 , \39133 );
and \U$38980 ( \39324 , \39321 , \39323 );
xor \U$38981 ( \39325 , \39152 , \39154 );
xor \U$38982 ( \39326 , \39325 , \39157 );
and \U$38983 ( \39327 , \39323 , \39326 );
and \U$38984 ( \39328 , \39321 , \39326 );
or \U$38985 ( \39329 , \39324 , \39327 , \39328 );
and \U$38986 ( \39330 , \39311 , \39329 );
xor \U$38987 ( \39331 , \39037 , \39053 );
xor \U$38988 ( \39332 , \39331 , \39070 );
xor \U$38989 ( \39333 , \39089 , \39105 );
xor \U$38990 ( \39334 , \39333 , \39122 );
and \U$38991 ( \39335 , \39332 , \39334 );
and \U$38992 ( \39336 , \39329 , \39335 );
and \U$38993 ( \39337 , \39311 , \39335 );
or \U$38994 ( \39338 , \39330 , \39336 , \39337 );
xor \U$38995 ( \39339 , \39073 , \39125 );
xor \U$38996 ( \39340 , \39339 , \39136 );
xor \U$38997 ( \39341 , \39141 , \39143 );
xor \U$38998 ( \39342 , \39341 , \39146 );
and \U$38999 ( \39343 , \39340 , \39342 );
xor \U$39000 ( \39344 , \39160 , \39162 );
xor \U$39001 ( \39345 , \39344 , \39164 );
and \U$39002 ( \39346 , \39342 , \39345 );
and \U$39003 ( \39347 , \39340 , \39345 );
or \U$39004 ( \39348 , \39343 , \39346 , \39347 );
and \U$39005 ( \39349 , \39338 , \39348 );
xor \U$39006 ( \39350 , \38886 , \38938 );
xor \U$39007 ( \39351 , \39350 , \38951 );
and \U$39008 ( \39352 , \39348 , \39351 );
and \U$39009 ( \39353 , \39338 , \39351 );
or \U$39010 ( \39354 , \39349 , \39352 , \39353 );
xor \U$39011 ( \39355 , \39139 , \39149 );
xor \U$39012 ( \39356 , \39355 , \39167 );
xor \U$39013 ( \39357 , \39172 , \39174 );
xor \U$39014 ( \39358 , \39357 , \39177 );
and \U$39015 ( \39359 , \39356 , \39358 );
and \U$39016 ( \39360 , \39354 , \39359 );
xor \U$39017 ( \39361 , \38954 , \38975 );
xor \U$39018 ( \39362 , \39361 , \38986 );
and \U$39019 ( \39363 , \39359 , \39362 );
and \U$39020 ( \39364 , \39354 , \39362 );
or \U$39021 ( \39365 , \39360 , \39363 , \39364 );
xor \U$39022 ( \39366 , \39186 , \39188 );
xor \U$39023 ( \39367 , \39366 , \39191 );
and \U$39024 ( \39368 , \39365 , \39367 );
and \U$39025 ( \39369 , \39200 , \39368 );
xor \U$39026 ( \39370 , \39200 , \39368 );
xor \U$39027 ( \39371 , \39365 , \39367 );
xor \U$39028 ( \39372 , \39354 , \39359 );
xor \U$39029 ( \39373 , \39372 , \39362 );
xor \U$39030 ( \39374 , \39170 , \39180 );
xor \U$39031 ( \39375 , \39374 , \39183 );
and \U$39032 ( \39376 , \39373 , \39375 );
and \U$39033 ( \39377 , \39371 , \39376 );
xor \U$39034 ( \39378 , \39371 , \39376 );
xor \U$39035 ( \39379 , \39373 , \39375 );
and \U$39036 ( \39380 , \29198 , \25631 );
and \U$39037 ( \39381 , \28952 , \25629 );
nor \U$39038 ( \39382 , \39380 , \39381 );
xnor \U$39039 ( \39383 , \39382 , \25399 );
and \U$39040 ( \39384 , \29522 , \25180 );
and \U$39041 ( \39385 , \29203 , \25178 );
nor \U$39042 ( \39386 , \39384 , \39385 );
xnor \U$39043 ( \39387 , \39386 , \25037 );
and \U$39044 ( \39388 , \39383 , \39387 );
and \U$39045 ( \39389 , \30375 , \24857 );
and \U$39046 ( \39390 , \29806 , \24855 );
nor \U$39047 ( \39391 , \39389 , \39390 );
xnor \U$39048 ( \39392 , \39391 , \24611 );
and \U$39049 ( \39393 , \39387 , \39392 );
and \U$39050 ( \39394 , \39383 , \39392 );
or \U$39051 ( \39395 , \39388 , \39393 , \39394 );
and \U$39052 ( \39396 , \30986 , \24462 );
and \U$39053 ( \39397 , \30383 , \24460 );
nor \U$39054 ( \39398 , \39396 , \39397 );
xnor \U$39055 ( \39399 , \39398 , \24275 );
and \U$39056 ( \39400 , \31172 , \24149 );
and \U$39057 ( \39401 , \30991 , \24147 );
nor \U$39058 ( \39402 , \39400 , \39401 );
xnor \U$39059 ( \39403 , \39402 , \23944 );
and \U$39060 ( \39404 , \39399 , \39403 );
nand \U$39061 ( \39405 , \31792 , \23741 );
xnor \U$39062 ( \39406 , \39405 , \23594 );
and \U$39063 ( \39407 , \39403 , \39406 );
and \U$39064 ( \39408 , \39399 , \39406 );
or \U$39065 ( \39409 , \39404 , \39407 , \39408 );
and \U$39066 ( \39410 , \39395 , \39409 );
and \U$39067 ( \39411 , \27325 , \27060 );
and \U$39068 ( \39412 , \26982 , \27058 );
nor \U$39069 ( \39413 , \39411 , \39412 );
xnor \U$39070 ( \39414 , \39413 , \26720 );
and \U$39071 ( \39415 , \27830 , \26471 );
and \U$39072 ( \39416 , \27527 , \26469 );
nor \U$39073 ( \39417 , \39415 , \39416 );
xnor \U$39074 ( \39418 , \39417 , \26230 );
and \U$39075 ( \39419 , \39414 , \39418 );
and \U$39076 ( \39420 , \28528 , \26005 );
and \U$39077 ( \39421 , \28002 , \26003 );
nor \U$39078 ( \39422 , \39420 , \39421 );
xnor \U$39079 ( \39423 , \39422 , \25817 );
and \U$39080 ( \39424 , \39418 , \39423 );
and \U$39081 ( \39425 , \39414 , \39423 );
or \U$39082 ( \39426 , \39419 , \39424 , \39425 );
and \U$39083 ( \39427 , \39409 , \39426 );
and \U$39084 ( \39428 , \39395 , \39426 );
or \U$39085 ( \39429 , \39410 , \39427 , \39428 );
and \U$39086 ( \39430 , \26073 , \28592 );
and \U$39087 ( \39431 , \25604 , \28590 );
nor \U$39088 ( \39432 , \39430 , \39431 );
xnor \U$39089 ( \39433 , \39432 , \28343 );
and \U$39090 ( \39434 , \26342 , \28063 );
and \U$39091 ( \39435 , \26078 , \28061 );
nor \U$39092 ( \39436 , \39434 , \39435 );
xnor \U$39093 ( \39437 , \39436 , \27803 );
and \U$39094 ( \39438 , \39433 , \39437 );
and \U$39095 ( \39439 , \26973 , \27569 );
and \U$39096 ( \39440 , \26601 , \27567 );
nor \U$39097 ( \39441 , \39439 , \39440 );
xnor \U$39098 ( \39442 , \39441 , \27254 );
and \U$39099 ( \39443 , \39437 , \39442 );
and \U$39100 ( \39444 , \39433 , \39442 );
or \U$39101 ( \39445 , \39438 , \39443 , \39444 );
and \U$39102 ( \39446 , \23970 , \31639 );
and \U$39103 ( \39447 , \23832 , \31636 );
nor \U$39104 ( \39448 , \39446 , \39447 );
xnor \U$39105 ( \39449 , \39448 , \30584 );
and \U$39106 ( \39450 , \24506 , \30826 );
and \U$39107 ( \39451 , \24089 , \30824 );
nor \U$39108 ( \39452 , \39450 , \39451 );
xnor \U$39109 ( \39453 , \39452 , \30587 );
and \U$39110 ( \39454 , \39449 , \39453 );
and \U$39111 ( \39455 , \39453 , \23594 );
and \U$39112 ( \39456 , \39449 , \23594 );
or \U$39113 ( \39457 , \39454 , \39455 , \39456 );
and \U$39114 ( \39458 , \39445 , \39457 );
and \U$39115 ( \39459 , \24836 , \30258 );
and \U$39116 ( \39460 , \24714 , \30256 );
nor \U$39117 ( \39461 , \39459 , \39460 );
xnor \U$39118 ( \39462 , \39461 , \29948 );
and \U$39119 ( \39463 , \25097 , \29721 );
and \U$39120 ( \39464 , \24841 , \29719 );
nor \U$39121 ( \39465 , \39463 , \39464 );
xnor \U$39122 ( \39466 , \39465 , \29350 );
and \U$39123 ( \39467 , \39462 , \39466 );
and \U$39124 ( \39468 , \25596 , \29159 );
and \U$39125 ( \39469 , \25294 , \29157 );
nor \U$39126 ( \39470 , \39468 , \39469 );
xnor \U$39127 ( \39471 , \39470 , \28841 );
and \U$39128 ( \39472 , \39466 , \39471 );
and \U$39129 ( \39473 , \39462 , \39471 );
or \U$39130 ( \39474 , \39467 , \39472 , \39473 );
and \U$39131 ( \39475 , \39457 , \39474 );
and \U$39132 ( \39476 , \39445 , \39474 );
or \U$39133 ( \39477 , \39458 , \39475 , \39476 );
and \U$39134 ( \39478 , \39429 , \39477 );
xor \U$39135 ( \39479 , \39256 , \39260 );
xor \U$39136 ( \39480 , \39479 , \39265 );
xor \U$39137 ( \39481 , \39272 , \39276 );
xor \U$39138 ( \39482 , \39481 , \39281 );
and \U$39139 ( \39483 , \39480 , \39482 );
xor \U$39140 ( \39484 , \39289 , \39293 );
and \U$39141 ( \39485 , \39482 , \39484 );
and \U$39142 ( \39486 , \39480 , \39484 );
or \U$39143 ( \39487 , \39483 , \39485 , \39486 );
and \U$39144 ( \39488 , \39477 , \39487 );
and \U$39145 ( \39489 , \39429 , \39487 );
or \U$39146 ( \39490 , \39478 , \39488 , \39489 );
xor \U$39147 ( \39491 , \39204 , \39208 );
xor \U$39148 ( \39492 , \39491 , \39213 );
xor \U$39149 ( \39493 , \39220 , \39224 );
xor \U$39150 ( \39494 , \39493 , \39229 );
and \U$39151 ( \39495 , \39492 , \39494 );
xor \U$39152 ( \39496 , \39237 , \39241 );
xor \U$39153 ( \39497 , \39496 , \39246 );
and \U$39154 ( \39498 , \39494 , \39497 );
and \U$39155 ( \39499 , \39492 , \39497 );
or \U$39156 ( \39500 , \39495 , \39498 , \39499 );
xor \U$39157 ( \39501 , \39029 , \39033 );
xor \U$39158 ( \39502 , \39501 , \23279 );
and \U$39159 ( \39503 , \39500 , \39502 );
xor \U$39160 ( \39504 , \39313 , \39315 );
xor \U$39161 ( \39505 , \39504 , \39318 );
and \U$39162 ( \39506 , \39502 , \39505 );
and \U$39163 ( \39507 , \39500 , \39505 );
or \U$39164 ( \39508 , \39503 , \39506 , \39507 );
and \U$39165 ( \39509 , \39490 , \39508 );
xor \U$39166 ( \39510 , \39216 , \39232 );
xor \U$39167 ( \39511 , \39510 , \39249 );
xor \U$39168 ( \39512 , \39268 , \39284 );
xor \U$39169 ( \39513 , \39512 , \39294 );
and \U$39170 ( \39514 , \39511 , \39513 );
xor \U$39171 ( \39515 , \39300 , \39302 );
xor \U$39172 ( \39516 , \39515 , \39305 );
and \U$39173 ( \39517 , \39513 , \39516 );
and \U$39174 ( \39518 , \39511 , \39516 );
or \U$39175 ( \39519 , \39514 , \39517 , \39518 );
and \U$39176 ( \39520 , \39508 , \39519 );
and \U$39177 ( \39521 , \39490 , \39519 );
or \U$39178 ( \39522 , \39509 , \39520 , \39521 );
xor \U$39179 ( \39523 , \39252 , \39297 );
xor \U$39180 ( \39524 , \39523 , \39308 );
xor \U$39181 ( \39525 , \39321 , \39323 );
xor \U$39182 ( \39526 , \39525 , \39326 );
and \U$39183 ( \39527 , \39524 , \39526 );
xor \U$39184 ( \39528 , \39332 , \39334 );
and \U$39185 ( \39529 , \39526 , \39528 );
and \U$39186 ( \39530 , \39524 , \39528 );
or \U$39187 ( \39531 , \39527 , \39529 , \39530 );
and \U$39188 ( \39532 , \39522 , \39531 );
xor \U$39189 ( \39533 , \39340 , \39342 );
xor \U$39190 ( \39534 , \39533 , \39345 );
and \U$39191 ( \39535 , \39531 , \39534 );
and \U$39192 ( \39536 , \39522 , \39534 );
or \U$39193 ( \39537 , \39532 , \39535 , \39536 );
xor \U$39194 ( \39538 , \39338 , \39348 );
xor \U$39195 ( \39539 , \39538 , \39351 );
and \U$39196 ( \39540 , \39537 , \39539 );
xor \U$39197 ( \39541 , \39356 , \39358 );
and \U$39198 ( \39542 , \39539 , \39541 );
and \U$39199 ( \39543 , \39537 , \39541 );
or \U$39200 ( \39544 , \39540 , \39542 , \39543 );
and \U$39201 ( \39545 , \39379 , \39544 );
xor \U$39202 ( \39546 , \39379 , \39544 );
xor \U$39203 ( \39547 , \39537 , \39539 );
xor \U$39204 ( \39548 , \39547 , \39541 );
and \U$39205 ( \39549 , \25294 , \29721 );
and \U$39206 ( \39550 , \25097 , \29719 );
nor \U$39207 ( \39551 , \39549 , \39550 );
xnor \U$39208 ( \39552 , \39551 , \29350 );
and \U$39209 ( \39553 , \25604 , \29159 );
and \U$39210 ( \39554 , \25596 , \29157 );
nor \U$39211 ( \39555 , \39553 , \39554 );
xnor \U$39212 ( \39556 , \39555 , \28841 );
and \U$39213 ( \39557 , \39552 , \39556 );
and \U$39214 ( \39558 , \26078 , \28592 );
and \U$39215 ( \39559 , \26073 , \28590 );
nor \U$39216 ( \39560 , \39558 , \39559 );
xnor \U$39217 ( \39561 , \39560 , \28343 );
and \U$39218 ( \39562 , \39556 , \39561 );
and \U$39219 ( \39563 , \39552 , \39561 );
or \U$39220 ( \39564 , \39557 , \39562 , \39563 );
and \U$39221 ( \39565 , \24089 , \31639 );
and \U$39222 ( \39566 , \23970 , \31636 );
nor \U$39223 ( \39567 , \39565 , \39566 );
xnor \U$39224 ( \39568 , \39567 , \30584 );
and \U$39225 ( \39569 , \24714 , \30826 );
and \U$39226 ( \39570 , \24506 , \30824 );
nor \U$39227 ( \39571 , \39569 , \39570 );
xnor \U$39228 ( \39572 , \39571 , \30587 );
and \U$39229 ( \39573 , \39568 , \39572 );
and \U$39230 ( \39574 , \24841 , \30258 );
and \U$39231 ( \39575 , \24836 , \30256 );
nor \U$39232 ( \39576 , \39574 , \39575 );
xnor \U$39233 ( \39577 , \39576 , \29948 );
and \U$39234 ( \39578 , \39572 , \39577 );
and \U$39235 ( \39579 , \39568 , \39577 );
or \U$39236 ( \39580 , \39573 , \39578 , \39579 );
and \U$39237 ( \39581 , \39564 , \39580 );
and \U$39238 ( \39582 , \26601 , \28063 );
and \U$39239 ( \39583 , \26342 , \28061 );
nor \U$39240 ( \39584 , \39582 , \39583 );
xnor \U$39241 ( \39585 , \39584 , \27803 );
and \U$39242 ( \39586 , \26982 , \27569 );
and \U$39243 ( \39587 , \26973 , \27567 );
nor \U$39244 ( \39588 , \39586 , \39587 );
xnor \U$39245 ( \39589 , \39588 , \27254 );
and \U$39246 ( \39590 , \39585 , \39589 );
and \U$39247 ( \39591 , \27527 , \27060 );
and \U$39248 ( \39592 , \27325 , \27058 );
nor \U$39249 ( \39593 , \39591 , \39592 );
xnor \U$39250 ( \39594 , \39593 , \26720 );
and \U$39251 ( \39595 , \39589 , \39594 );
and \U$39252 ( \39596 , \39585 , \39594 );
or \U$39253 ( \39597 , \39590 , \39595 , \39596 );
and \U$39254 ( \39598 , \39580 , \39597 );
and \U$39255 ( \39599 , \39564 , \39597 );
or \U$39256 ( \39600 , \39581 , \39598 , \39599 );
xor \U$39257 ( \39601 , \39383 , \39387 );
xor \U$39258 ( \39602 , \39601 , \39392 );
xor \U$39259 ( \39603 , \39433 , \39437 );
xor \U$39260 ( \39604 , \39603 , \39442 );
and \U$39261 ( \39605 , \39602 , \39604 );
xor \U$39262 ( \39606 , \39414 , \39418 );
xor \U$39263 ( \39607 , \39606 , \39423 );
and \U$39264 ( \39608 , \39604 , \39607 );
and \U$39265 ( \39609 , \39602 , \39607 );
or \U$39266 ( \39610 , \39605 , \39608 , \39609 );
and \U$39267 ( \39611 , \39600 , \39610 );
and \U$39268 ( \39612 , \28002 , \26471 );
and \U$39269 ( \39613 , \27830 , \26469 );
nor \U$39270 ( \39614 , \39612 , \39613 );
xnor \U$39271 ( \39615 , \39614 , \26230 );
and \U$39272 ( \39616 , \28952 , \26005 );
and \U$39273 ( \39617 , \28528 , \26003 );
nor \U$39274 ( \39618 , \39616 , \39617 );
xnor \U$39275 ( \39619 , \39618 , \25817 );
and \U$39276 ( \39620 , \39615 , \39619 );
and \U$39277 ( \39621 , \29203 , \25631 );
and \U$39278 ( \39622 , \29198 , \25629 );
nor \U$39279 ( \39623 , \39621 , \39622 );
xnor \U$39280 ( \39624 , \39623 , \25399 );
and \U$39281 ( \39625 , \39619 , \39624 );
and \U$39282 ( \39626 , \39615 , \39624 );
or \U$39283 ( \39627 , \39620 , \39625 , \39626 );
and \U$39284 ( \39628 , \29806 , \25180 );
and \U$39285 ( \39629 , \29522 , \25178 );
nor \U$39286 ( \39630 , \39628 , \39629 );
xnor \U$39287 ( \39631 , \39630 , \25037 );
and \U$39288 ( \39632 , \30383 , \24857 );
and \U$39289 ( \39633 , \30375 , \24855 );
nor \U$39290 ( \39634 , \39632 , \39633 );
xnor \U$39291 ( \39635 , \39634 , \24611 );
and \U$39292 ( \39636 , \39631 , \39635 );
and \U$39293 ( \39637 , \30991 , \24462 );
and \U$39294 ( \39638 , \30986 , \24460 );
nor \U$39295 ( \39639 , \39637 , \39638 );
xnor \U$39296 ( \39640 , \39639 , \24275 );
and \U$39297 ( \39641 , \39635 , \39640 );
and \U$39298 ( \39642 , \39631 , \39640 );
or \U$39299 ( \39643 , \39636 , \39641 , \39642 );
and \U$39300 ( \39644 , \39627 , \39643 );
xor \U$39301 ( \39645 , \39399 , \39403 );
xor \U$39302 ( \39646 , \39645 , \39406 );
and \U$39303 ( \39647 , \39643 , \39646 );
and \U$39304 ( \39648 , \39627 , \39646 );
or \U$39305 ( \39649 , \39644 , \39647 , \39648 );
and \U$39306 ( \39650 , \39610 , \39649 );
and \U$39307 ( \39651 , \39600 , \39649 );
or \U$39308 ( \39652 , \39611 , \39650 , \39651 );
xor \U$39309 ( \39653 , \39395 , \39409 );
xor \U$39310 ( \39654 , \39653 , \39426 );
xor \U$39311 ( \39655 , \39492 , \39494 );
xor \U$39312 ( \39656 , \39655 , \39497 );
and \U$39313 ( \39657 , \39654 , \39656 );
xor \U$39314 ( \39658 , \39480 , \39482 );
xor \U$39315 ( \39659 , \39658 , \39484 );
and \U$39316 ( \39660 , \39656 , \39659 );
and \U$39317 ( \39661 , \39654 , \39659 );
or \U$39318 ( \39662 , \39657 , \39660 , \39661 );
and \U$39319 ( \39663 , \39652 , \39662 );
xor \U$39320 ( \39664 , \39511 , \39513 );
xor \U$39321 ( \39665 , \39664 , \39516 );
and \U$39322 ( \39666 , \39662 , \39665 );
and \U$39323 ( \39667 , \39652 , \39665 );
or \U$39324 ( \39668 , \39663 , \39666 , \39667 );
xor \U$39325 ( \39669 , \39490 , \39508 );
xor \U$39326 ( \39670 , \39669 , \39519 );
and \U$39327 ( \39671 , \39668 , \39670 );
xor \U$39328 ( \39672 , \39524 , \39526 );
xor \U$39329 ( \39673 , \39672 , \39528 );
and \U$39330 ( \39674 , \39670 , \39673 );
and \U$39331 ( \39675 , \39668 , \39673 );
or \U$39332 ( \39676 , \39671 , \39674 , \39675 );
xor \U$39333 ( \39677 , \39311 , \39329 );
xor \U$39334 ( \39678 , \39677 , \39335 );
and \U$39335 ( \39679 , \39676 , \39678 );
xor \U$39336 ( \39680 , \39522 , \39531 );
xor \U$39337 ( \39681 , \39680 , \39534 );
and \U$39338 ( \39682 , \39678 , \39681 );
and \U$39339 ( \39683 , \39676 , \39681 );
or \U$39340 ( \39684 , \39679 , \39682 , \39683 );
and \U$39341 ( \39685 , \39548 , \39684 );
xor \U$39342 ( \39686 , \39548 , \39684 );
xor \U$39343 ( \39687 , \39676 , \39678 );
xor \U$39344 ( \39688 , \39687 , \39681 );
and \U$39345 ( \39689 , \25097 , \30258 );
and \U$39346 ( \39690 , \24841 , \30256 );
nor \U$39347 ( \39691 , \39689 , \39690 );
xnor \U$39348 ( \39692 , \39691 , \29948 );
and \U$39349 ( \39693 , \25596 , \29721 );
and \U$39350 ( \39694 , \25294 , \29719 );
nor \U$39351 ( \39695 , \39693 , \39694 );
xnor \U$39352 ( \39696 , \39695 , \29350 );
and \U$39353 ( \39697 , \39692 , \39696 );
and \U$39354 ( \39698 , \26073 , \29159 );
and \U$39355 ( \39699 , \25604 , \29157 );
nor \U$39356 ( \39700 , \39698 , \39699 );
xnor \U$39357 ( \39701 , \39700 , \28841 );
and \U$39358 ( \39702 , \39696 , \39701 );
and \U$39359 ( \39703 , \39692 , \39701 );
or \U$39360 ( \39704 , \39697 , \39702 , \39703 );
and \U$39361 ( \39705 , \26342 , \28592 );
and \U$39362 ( \39706 , \26078 , \28590 );
nor \U$39363 ( \39707 , \39705 , \39706 );
xnor \U$39364 ( \39708 , \39707 , \28343 );
and \U$39365 ( \39709 , \26973 , \28063 );
and \U$39366 ( \39710 , \26601 , \28061 );
nor \U$39367 ( \39711 , \39709 , \39710 );
xnor \U$39368 ( \39712 , \39711 , \27803 );
and \U$39369 ( \39713 , \39708 , \39712 );
and \U$39370 ( \39714 , \27325 , \27569 );
and \U$39371 ( \39715 , \26982 , \27567 );
nor \U$39372 ( \39716 , \39714 , \39715 );
xnor \U$39373 ( \39717 , \39716 , \27254 );
and \U$39374 ( \39718 , \39712 , \39717 );
and \U$39375 ( \39719 , \39708 , \39717 );
or \U$39376 ( \39720 , \39713 , \39718 , \39719 );
and \U$39377 ( \39721 , \39704 , \39720 );
and \U$39378 ( \39722 , \24506 , \31639 );
and \U$39379 ( \39723 , \24089 , \31636 );
nor \U$39380 ( \39724 , \39722 , \39723 );
xnor \U$39381 ( \39725 , \39724 , \30584 );
and \U$39382 ( \39726 , \24836 , \30826 );
and \U$39383 ( \39727 , \24714 , \30824 );
nor \U$39384 ( \39728 , \39726 , \39727 );
xnor \U$39385 ( \39729 , \39728 , \30587 );
and \U$39386 ( \39730 , \39725 , \39729 );
and \U$39387 ( \39731 , \39729 , \23944 );
and \U$39388 ( \39732 , \39725 , \23944 );
or \U$39389 ( \39733 , \39730 , \39731 , \39732 );
and \U$39390 ( \39734 , \39720 , \39733 );
and \U$39391 ( \39735 , \39704 , \39733 );
or \U$39392 ( \39736 , \39721 , \39734 , \39735 );
and \U$39393 ( \39737 , \29522 , \25631 );
and \U$39394 ( \39738 , \29203 , \25629 );
nor \U$39395 ( \39739 , \39737 , \39738 );
xnor \U$39396 ( \39740 , \39739 , \25399 );
and \U$39397 ( \39741 , \30375 , \25180 );
and \U$39398 ( \39742 , \29806 , \25178 );
nor \U$39399 ( \39743 , \39741 , \39742 );
xnor \U$39400 ( \39744 , \39743 , \25037 );
and \U$39401 ( \39745 , \39740 , \39744 );
and \U$39402 ( \39746 , \30986 , \24857 );
and \U$39403 ( \39747 , \30383 , \24855 );
nor \U$39404 ( \39748 , \39746 , \39747 );
xnor \U$39405 ( \39749 , \39748 , \24611 );
and \U$39406 ( \39750 , \39744 , \39749 );
and \U$39407 ( \39751 , \39740 , \39749 );
or \U$39408 ( \39752 , \39745 , \39750 , \39751 );
and \U$39409 ( \39753 , \27830 , \27060 );
and \U$39410 ( \39754 , \27527 , \27058 );
nor \U$39411 ( \39755 , \39753 , \39754 );
xnor \U$39412 ( \39756 , \39755 , \26720 );
and \U$39413 ( \39757 , \28528 , \26471 );
and \U$39414 ( \39758 , \28002 , \26469 );
nor \U$39415 ( \39759 , \39757 , \39758 );
xnor \U$39416 ( \39760 , \39759 , \26230 );
and \U$39417 ( \39761 , \39756 , \39760 );
and \U$39418 ( \39762 , \29198 , \26005 );
and \U$39419 ( \39763 , \28952 , \26003 );
nor \U$39420 ( \39764 , \39762 , \39763 );
xnor \U$39421 ( \39765 , \39764 , \25817 );
and \U$39422 ( \39766 , \39760 , \39765 );
and \U$39423 ( \39767 , \39756 , \39765 );
or \U$39424 ( \39768 , \39761 , \39766 , \39767 );
and \U$39425 ( \39769 , \39752 , \39768 );
and \U$39426 ( \39770 , \31792 , \24149 );
and \U$39427 ( \39771 , \31172 , \24147 );
nor \U$39428 ( \39772 , \39770 , \39771 );
xnor \U$39429 ( \39773 , \39772 , \23944 );
and \U$39430 ( \39774 , \39768 , \39773 );
and \U$39431 ( \39775 , \39752 , \39773 );
or \U$39432 ( \39776 , \39769 , \39774 , \39775 );
and \U$39433 ( \39777 , \39736 , \39776 );
xor \U$39434 ( \39778 , \39615 , \39619 );
xor \U$39435 ( \39779 , \39778 , \39624 );
xor \U$39436 ( \39780 , \39631 , \39635 );
xor \U$39437 ( \39781 , \39780 , \39640 );
and \U$39438 ( \39782 , \39779 , \39781 );
xor \U$39439 ( \39783 , \39585 , \39589 );
xor \U$39440 ( \39784 , \39783 , \39594 );
and \U$39441 ( \39785 , \39781 , \39784 );
and \U$39442 ( \39786 , \39779 , \39784 );
or \U$39443 ( \39787 , \39782 , \39785 , \39786 );
and \U$39444 ( \39788 , \39776 , \39787 );
and \U$39445 ( \39789 , \39736 , \39787 );
or \U$39446 ( \39790 , \39777 , \39788 , \39789 );
xor \U$39447 ( \39791 , \39449 , \39453 );
xor \U$39448 ( \39792 , \39791 , \23594 );
xor \U$39449 ( \39793 , \39462 , \39466 );
xor \U$39450 ( \39794 , \39793 , \39471 );
and \U$39451 ( \39795 , \39792 , \39794 );
xor \U$39452 ( \39796 , \39602 , \39604 );
xor \U$39453 ( \39797 , \39796 , \39607 );
and \U$39454 ( \39798 , \39794 , \39797 );
and \U$39455 ( \39799 , \39792 , \39797 );
or \U$39456 ( \39800 , \39795 , \39798 , \39799 );
and \U$39457 ( \39801 , \39790 , \39800 );
xor \U$39458 ( \39802 , \39564 , \39580 );
xor \U$39459 ( \39803 , \39802 , \39597 );
xor \U$39460 ( \39804 , \39627 , \39643 );
xor \U$39461 ( \39805 , \39804 , \39646 );
and \U$39462 ( \39806 , \39803 , \39805 );
and \U$39463 ( \39807 , \39800 , \39806 );
and \U$39464 ( \39808 , \39790 , \39806 );
or \U$39465 ( \39809 , \39801 , \39807 , \39808 );
xor \U$39466 ( \39810 , \39445 , \39457 );
xor \U$39467 ( \39811 , \39810 , \39474 );
xor \U$39468 ( \39812 , \39600 , \39610 );
xor \U$39469 ( \39813 , \39812 , \39649 );
and \U$39470 ( \39814 , \39811 , \39813 );
xor \U$39471 ( \39815 , \39654 , \39656 );
xor \U$39472 ( \39816 , \39815 , \39659 );
and \U$39473 ( \39817 , \39813 , \39816 );
and \U$39474 ( \39818 , \39811 , \39816 );
or \U$39475 ( \39819 , \39814 , \39817 , \39818 );
and \U$39476 ( \39820 , \39809 , \39819 );
xor \U$39477 ( \39821 , \39500 , \39502 );
xor \U$39478 ( \39822 , \39821 , \39505 );
and \U$39479 ( \39823 , \39819 , \39822 );
and \U$39480 ( \39824 , \39809 , \39822 );
or \U$39481 ( \39825 , \39820 , \39823 , \39824 );
xor \U$39482 ( \39826 , \39429 , \39477 );
xor \U$39483 ( \39827 , \39826 , \39487 );
xor \U$39484 ( \39828 , \39652 , \39662 );
xor \U$39485 ( \39829 , \39828 , \39665 );
and \U$39486 ( \39830 , \39827 , \39829 );
and \U$39487 ( \39831 , \39825 , \39830 );
xor \U$39488 ( \39832 , \39668 , \39670 );
xor \U$39489 ( \39833 , \39832 , \39673 );
and \U$39490 ( \39834 , \39830 , \39833 );
and \U$39491 ( \39835 , \39825 , \39833 );
or \U$39492 ( \39836 , \39831 , \39834 , \39835 );
and \U$39493 ( \39837 , \39688 , \39836 );
xor \U$39494 ( \39838 , \39688 , \39836 );
xor \U$39495 ( \39839 , \39825 , \39830 );
xor \U$39496 ( \39840 , \39839 , \39833 );
and \U$39497 ( \39841 , \26982 , \28063 );
and \U$39498 ( \39842 , \26973 , \28061 );
nor \U$39499 ( \39843 , \39841 , \39842 );
xnor \U$39500 ( \39844 , \39843 , \27803 );
and \U$39501 ( \39845 , \27527 , \27569 );
and \U$39502 ( \39846 , \27325 , \27567 );
nor \U$39503 ( \39847 , \39845 , \39846 );
xnor \U$39504 ( \39848 , \39847 , \27254 );
and \U$39505 ( \39849 , \39844 , \39848 );
and \U$39506 ( \39850 , \28002 , \27060 );
and \U$39507 ( \39851 , \27830 , \27058 );
nor \U$39508 ( \39852 , \39850 , \39851 );
xnor \U$39509 ( \39853 , \39852 , \26720 );
and \U$39510 ( \39854 , \39848 , \39853 );
and \U$39511 ( \39855 , \39844 , \39853 );
or \U$39512 ( \39856 , \39849 , \39854 , \39855 );
and \U$39513 ( \39857 , \25604 , \29721 );
and \U$39514 ( \39858 , \25596 , \29719 );
nor \U$39515 ( \39859 , \39857 , \39858 );
xnor \U$39516 ( \39860 , \39859 , \29350 );
and \U$39517 ( \39861 , \26078 , \29159 );
and \U$39518 ( \39862 , \26073 , \29157 );
nor \U$39519 ( \39863 , \39861 , \39862 );
xnor \U$39520 ( \39864 , \39863 , \28841 );
and \U$39521 ( \39865 , \39860 , \39864 );
and \U$39522 ( \39866 , \26601 , \28592 );
and \U$39523 ( \39867 , \26342 , \28590 );
nor \U$39524 ( \39868 , \39866 , \39867 );
xnor \U$39525 ( \39869 , \39868 , \28343 );
and \U$39526 ( \39870 , \39864 , \39869 );
and \U$39527 ( \39871 , \39860 , \39869 );
or \U$39528 ( \39872 , \39865 , \39870 , \39871 );
and \U$39529 ( \39873 , \39856 , \39872 );
and \U$39530 ( \39874 , \24714 , \31639 );
and \U$39531 ( \39875 , \24506 , \31636 );
nor \U$39532 ( \39876 , \39874 , \39875 );
xnor \U$39533 ( \39877 , \39876 , \30584 );
and \U$39534 ( \39878 , \24841 , \30826 );
and \U$39535 ( \39879 , \24836 , \30824 );
nor \U$39536 ( \39880 , \39878 , \39879 );
xnor \U$39537 ( \39881 , \39880 , \30587 );
and \U$39538 ( \39882 , \39877 , \39881 );
and \U$39539 ( \39883 , \25294 , \30258 );
and \U$39540 ( \39884 , \25097 , \30256 );
nor \U$39541 ( \39885 , \39883 , \39884 );
xnor \U$39542 ( \39886 , \39885 , \29948 );
and \U$39543 ( \39887 , \39881 , \39886 );
and \U$39544 ( \39888 , \39877 , \39886 );
or \U$39545 ( \39889 , \39882 , \39887 , \39888 );
and \U$39546 ( \39890 , \39872 , \39889 );
and \U$39547 ( \39891 , \39856 , \39889 );
or \U$39548 ( \39892 , \39873 , \39890 , \39891 );
and \U$39549 ( \39893 , \30383 , \25180 );
and \U$39550 ( \39894 , \30375 , \25178 );
nor \U$39551 ( \39895 , \39893 , \39894 );
xnor \U$39552 ( \39896 , \39895 , \25037 );
and \U$39553 ( \39897 , \30991 , \24857 );
and \U$39554 ( \39898 , \30986 , \24855 );
nor \U$39555 ( \39899 , \39897 , \39898 );
xnor \U$39556 ( \39900 , \39899 , \24611 );
and \U$39557 ( \39901 , \39896 , \39900 );
and \U$39558 ( \39902 , \31792 , \24462 );
and \U$39559 ( \39903 , \31172 , \24460 );
nor \U$39560 ( \39904 , \39902 , \39903 );
xnor \U$39561 ( \39905 , \39904 , \24275 );
and \U$39562 ( \39906 , \39900 , \39905 );
and \U$39563 ( \39907 , \39896 , \39905 );
or \U$39564 ( \39908 , \39901 , \39906 , \39907 );
and \U$39565 ( \39909 , \28952 , \26471 );
and \U$39566 ( \39910 , \28528 , \26469 );
nor \U$39567 ( \39911 , \39909 , \39910 );
xnor \U$39568 ( \39912 , \39911 , \26230 );
and \U$39569 ( \39913 , \29203 , \26005 );
and \U$39570 ( \39914 , \29198 , \26003 );
nor \U$39571 ( \39915 , \39913 , \39914 );
xnor \U$39572 ( \39916 , \39915 , \25817 );
and \U$39573 ( \39917 , \39912 , \39916 );
and \U$39574 ( \39918 , \29806 , \25631 );
and \U$39575 ( \39919 , \29522 , \25629 );
nor \U$39576 ( \39920 , \39918 , \39919 );
xnor \U$39577 ( \39921 , \39920 , \25399 );
and \U$39578 ( \39922 , \39916 , \39921 );
and \U$39579 ( \39923 , \39912 , \39921 );
or \U$39580 ( \39924 , \39917 , \39922 , \39923 );
and \U$39581 ( \39925 , \39908 , \39924 );
and \U$39582 ( \39926 , \31172 , \24462 );
and \U$39583 ( \39927 , \30991 , \24460 );
nor \U$39584 ( \39928 , \39926 , \39927 );
xnor \U$39585 ( \39929 , \39928 , \24275 );
and \U$39586 ( \39930 , \39924 , \39929 );
and \U$39587 ( \39931 , \39908 , \39929 );
or \U$39588 ( \39932 , \39925 , \39930 , \39931 );
and \U$39589 ( \39933 , \39892 , \39932 );
nand \U$39590 ( \39934 , \31792 , \24147 );
xnor \U$39591 ( \39935 , \39934 , \23944 );
xor \U$39592 ( \39936 , \39740 , \39744 );
xor \U$39593 ( \39937 , \39936 , \39749 );
and \U$39594 ( \39938 , \39935 , \39937 );
xor \U$39595 ( \39939 , \39756 , \39760 );
xor \U$39596 ( \39940 , \39939 , \39765 );
and \U$39597 ( \39941 , \39937 , \39940 );
and \U$39598 ( \39942 , \39935 , \39940 );
or \U$39599 ( \39943 , \39938 , \39941 , \39942 );
and \U$39600 ( \39944 , \39932 , \39943 );
and \U$39601 ( \39945 , \39892 , \39943 );
or \U$39602 ( \39946 , \39933 , \39944 , \39945 );
xor \U$39603 ( \39947 , \39692 , \39696 );
xor \U$39604 ( \39948 , \39947 , \39701 );
xor \U$39605 ( \39949 , \39708 , \39712 );
xor \U$39606 ( \39950 , \39949 , \39717 );
and \U$39607 ( \39951 , \39948 , \39950 );
xor \U$39608 ( \39952 , \39725 , \39729 );
xor \U$39609 ( \39953 , \39952 , \23944 );
and \U$39610 ( \39954 , \39950 , \39953 );
and \U$39611 ( \39955 , \39948 , \39953 );
or \U$39612 ( \39956 , \39951 , \39954 , \39955 );
xor \U$39613 ( \39957 , \39552 , \39556 );
xor \U$39614 ( \39958 , \39957 , \39561 );
and \U$39615 ( \39959 , \39956 , \39958 );
xor \U$39616 ( \39960 , \39568 , \39572 );
xor \U$39617 ( \39961 , \39960 , \39577 );
and \U$39618 ( \39962 , \39958 , \39961 );
and \U$39619 ( \39963 , \39956 , \39961 );
or \U$39620 ( \39964 , \39959 , \39962 , \39963 );
and \U$39621 ( \39965 , \39946 , \39964 );
xor \U$39622 ( \39966 , \39704 , \39720 );
xor \U$39623 ( \39967 , \39966 , \39733 );
xor \U$39624 ( \39968 , \39752 , \39768 );
xor \U$39625 ( \39969 , \39968 , \39773 );
and \U$39626 ( \39970 , \39967 , \39969 );
xor \U$39627 ( \39971 , \39779 , \39781 );
xor \U$39628 ( \39972 , \39971 , \39784 );
and \U$39629 ( \39973 , \39969 , \39972 );
and \U$39630 ( \39974 , \39967 , \39972 );
or \U$39631 ( \39975 , \39970 , \39973 , \39974 );
and \U$39632 ( \39976 , \39964 , \39975 );
and \U$39633 ( \39977 , \39946 , \39975 );
or \U$39634 ( \39978 , \39965 , \39976 , \39977 );
xor \U$39635 ( \39979 , \39736 , \39776 );
xor \U$39636 ( \39980 , \39979 , \39787 );
xor \U$39637 ( \39981 , \39792 , \39794 );
xor \U$39638 ( \39982 , \39981 , \39797 );
and \U$39639 ( \39983 , \39980 , \39982 );
xor \U$39640 ( \39984 , \39803 , \39805 );
and \U$39641 ( \39985 , \39982 , \39984 );
and \U$39642 ( \39986 , \39980 , \39984 );
or \U$39643 ( \39987 , \39983 , \39985 , \39986 );
and \U$39644 ( \39988 , \39978 , \39987 );
xor \U$39645 ( \39989 , \39811 , \39813 );
xor \U$39646 ( \39990 , \39989 , \39816 );
and \U$39647 ( \39991 , \39987 , \39990 );
and \U$39648 ( \39992 , \39978 , \39990 );
or \U$39649 ( \39993 , \39988 , \39991 , \39992 );
xor \U$39650 ( \39994 , \39809 , \39819 );
xor \U$39651 ( \39995 , \39994 , \39822 );
and \U$39652 ( \39996 , \39993 , \39995 );
xor \U$39653 ( \39997 , \39827 , \39829 );
and \U$39654 ( \39998 , \39995 , \39997 );
and \U$39655 ( \39999 , \39993 , \39997 );
or \U$39656 ( \40000 , \39996 , \39998 , \39999 );
and \U$39657 ( \40001 , \39840 , \40000 );
xor \U$39658 ( \40002 , \39840 , \40000 );
xor \U$39659 ( \40003 , \39993 , \39995 );
xor \U$39660 ( \40004 , \40003 , \39997 );
and \U$39661 ( \40005 , \26973 , \28592 );
and \U$39662 ( \40006 , \26601 , \28590 );
nor \U$39663 ( \40007 , \40005 , \40006 );
xnor \U$39664 ( \40008 , \40007 , \28343 );
and \U$39665 ( \40009 , \27325 , \28063 );
and \U$39666 ( \40010 , \26982 , \28061 );
nor \U$39667 ( \40011 , \40009 , \40010 );
xnor \U$39668 ( \40012 , \40011 , \27803 );
and \U$39669 ( \40013 , \40008 , \40012 );
and \U$39670 ( \40014 , \27830 , \27569 );
and \U$39671 ( \40015 , \27527 , \27567 );
nor \U$39672 ( \40016 , \40014 , \40015 );
xnor \U$39673 ( \40017 , \40016 , \27254 );
and \U$39674 ( \40018 , \40012 , \40017 );
and \U$39675 ( \40019 , \40008 , \40017 );
or \U$39676 ( \40020 , \40013 , \40018 , \40019 );
and \U$39677 ( \40021 , \25596 , \30258 );
and \U$39678 ( \40022 , \25294 , \30256 );
nor \U$39679 ( \40023 , \40021 , \40022 );
xnor \U$39680 ( \40024 , \40023 , \29948 );
and \U$39681 ( \40025 , \26073 , \29721 );
and \U$39682 ( \40026 , \25604 , \29719 );
nor \U$39683 ( \40027 , \40025 , \40026 );
xnor \U$39684 ( \40028 , \40027 , \29350 );
and \U$39685 ( \40029 , \40024 , \40028 );
and \U$39686 ( \40030 , \26342 , \29159 );
and \U$39687 ( \40031 , \26078 , \29157 );
nor \U$39688 ( \40032 , \40030 , \40031 );
xnor \U$39689 ( \40033 , \40032 , \28841 );
and \U$39690 ( \40034 , \40028 , \40033 );
and \U$39691 ( \40035 , \40024 , \40033 );
or \U$39692 ( \40036 , \40029 , \40034 , \40035 );
and \U$39693 ( \40037 , \40020 , \40036 );
and \U$39694 ( \40038 , \24836 , \31639 );
and \U$39695 ( \40039 , \24714 , \31636 );
nor \U$39696 ( \40040 , \40038 , \40039 );
xnor \U$39697 ( \40041 , \40040 , \30584 );
and \U$39698 ( \40042 , \25097 , \30826 );
and \U$39699 ( \40043 , \24841 , \30824 );
nor \U$39700 ( \40044 , \40042 , \40043 );
xnor \U$39701 ( \40045 , \40044 , \30587 );
and \U$39702 ( \40046 , \40041 , \40045 );
and \U$39703 ( \40047 , \40045 , \24275 );
and \U$39704 ( \40048 , \40041 , \24275 );
or \U$39705 ( \40049 , \40046 , \40047 , \40048 );
and \U$39706 ( \40050 , \40036 , \40049 );
and \U$39707 ( \40051 , \40020 , \40049 );
or \U$39708 ( \40052 , \40037 , \40050 , \40051 );
and \U$39709 ( \40053 , \28528 , \27060 );
and \U$39710 ( \40054 , \28002 , \27058 );
nor \U$39711 ( \40055 , \40053 , \40054 );
xnor \U$39712 ( \40056 , \40055 , \26720 );
and \U$39713 ( \40057 , \29198 , \26471 );
and \U$39714 ( \40058 , \28952 , \26469 );
nor \U$39715 ( \40059 , \40057 , \40058 );
xnor \U$39716 ( \40060 , \40059 , \26230 );
and \U$39717 ( \40061 , \40056 , \40060 );
and \U$39718 ( \40062 , \29522 , \26005 );
and \U$39719 ( \40063 , \29203 , \26003 );
nor \U$39720 ( \40064 , \40062 , \40063 );
xnor \U$39721 ( \40065 , \40064 , \25817 );
and \U$39722 ( \40066 , \40060 , \40065 );
and \U$39723 ( \40067 , \40056 , \40065 );
or \U$39724 ( \40068 , \40061 , \40066 , \40067 );
and \U$39725 ( \40069 , \30375 , \25631 );
and \U$39726 ( \40070 , \29806 , \25629 );
nor \U$39727 ( \40071 , \40069 , \40070 );
xnor \U$39728 ( \40072 , \40071 , \25399 );
and \U$39729 ( \40073 , \30986 , \25180 );
and \U$39730 ( \40074 , \30383 , \25178 );
nor \U$39731 ( \40075 , \40073 , \40074 );
xnor \U$39732 ( \40076 , \40075 , \25037 );
and \U$39733 ( \40077 , \40072 , \40076 );
and \U$39734 ( \40078 , \31172 , \24857 );
and \U$39735 ( \40079 , \30991 , \24855 );
nor \U$39736 ( \40080 , \40078 , \40079 );
xnor \U$39737 ( \40081 , \40080 , \24611 );
and \U$39738 ( \40082 , \40076 , \40081 );
and \U$39739 ( \40083 , \40072 , \40081 );
or \U$39740 ( \40084 , \40077 , \40082 , \40083 );
and \U$39741 ( \40085 , \40068 , \40084 );
xor \U$39742 ( \40086 , \39896 , \39900 );
xor \U$39743 ( \40087 , \40086 , \39905 );
and \U$39744 ( \40088 , \40084 , \40087 );
and \U$39745 ( \40089 , \40068 , \40087 );
or \U$39746 ( \40090 , \40085 , \40088 , \40089 );
and \U$39747 ( \40091 , \40052 , \40090 );
xor \U$39748 ( \40092 , \39844 , \39848 );
xor \U$39749 ( \40093 , \40092 , \39853 );
xor \U$39750 ( \40094 , \39860 , \39864 );
xor \U$39751 ( \40095 , \40094 , \39869 );
and \U$39752 ( \40096 , \40093 , \40095 );
xor \U$39753 ( \40097 , \39912 , \39916 );
xor \U$39754 ( \40098 , \40097 , \39921 );
and \U$39755 ( \40099 , \40095 , \40098 );
and \U$39756 ( \40100 , \40093 , \40098 );
or \U$39757 ( \40101 , \40096 , \40099 , \40100 );
and \U$39758 ( \40102 , \40090 , \40101 );
and \U$39759 ( \40103 , \40052 , \40101 );
or \U$39760 ( \40104 , \40091 , \40102 , \40103 );
xor \U$39761 ( \40105 , \39908 , \39924 );
xor \U$39762 ( \40106 , \40105 , \39929 );
xor \U$39763 ( \40107 , \39948 , \39950 );
xor \U$39764 ( \40108 , \40107 , \39953 );
and \U$39765 ( \40109 , \40106 , \40108 );
xor \U$39766 ( \40110 , \39935 , \39937 );
xor \U$39767 ( \40111 , \40110 , \39940 );
and \U$39768 ( \40112 , \40108 , \40111 );
and \U$39769 ( \40113 , \40106 , \40111 );
or \U$39770 ( \40114 , \40109 , \40112 , \40113 );
and \U$39771 ( \40115 , \40104 , \40114 );
xor \U$39772 ( \40116 , \39967 , \39969 );
xor \U$39773 ( \40117 , \40116 , \39972 );
and \U$39774 ( \40118 , \40114 , \40117 );
and \U$39775 ( \40119 , \40104 , \40117 );
or \U$39776 ( \40120 , \40115 , \40118 , \40119 );
xor \U$39777 ( \40121 , \39892 , \39932 );
xor \U$39778 ( \40122 , \40121 , \39943 );
xor \U$39779 ( \40123 , \39956 , \39958 );
xor \U$39780 ( \40124 , \40123 , \39961 );
and \U$39781 ( \40125 , \40122 , \40124 );
and \U$39782 ( \40126 , \40120 , \40125 );
xor \U$39783 ( \40127 , \39980 , \39982 );
xor \U$39784 ( \40128 , \40127 , \39984 );
and \U$39785 ( \40129 , \40125 , \40128 );
and \U$39786 ( \40130 , \40120 , \40128 );
or \U$39787 ( \40131 , \40126 , \40129 , \40130 );
xor \U$39788 ( \40132 , \39790 , \39800 );
xor \U$39789 ( \40133 , \40132 , \39806 );
and \U$39790 ( \40134 , \40131 , \40133 );
xor \U$39791 ( \40135 , \39978 , \39987 );
xor \U$39792 ( \40136 , \40135 , \39990 );
and \U$39793 ( \40137 , \40133 , \40136 );
and \U$39794 ( \40138 , \40131 , \40136 );
or \U$39795 ( \40139 , \40134 , \40137 , \40138 );
and \U$39796 ( \40140 , \40004 , \40139 );
xor \U$39797 ( \40141 , \40004 , \40139 );
xor \U$39798 ( \40142 , \40131 , \40133 );
xor \U$39799 ( \40143 , \40142 , \40136 );
and \U$39800 ( \40144 , \24841 , \31639 );
and \U$39801 ( \40145 , \24836 , \31636 );
nor \U$39802 ( \40146 , \40144 , \40145 );
xnor \U$39803 ( \40147 , \40146 , \30584 );
and \U$39804 ( \40148 , \25294 , \30826 );
and \U$39805 ( \40149 , \25097 , \30824 );
nor \U$39806 ( \40150 , \40148 , \40149 );
xnor \U$39807 ( \40151 , \40150 , \30587 );
and \U$39808 ( \40152 , \40147 , \40151 );
and \U$39809 ( \40153 , \25604 , \30258 );
and \U$39810 ( \40154 , \25596 , \30256 );
nor \U$39811 ( \40155 , \40153 , \40154 );
xnor \U$39812 ( \40156 , \40155 , \29948 );
and \U$39813 ( \40157 , \40151 , \40156 );
and \U$39814 ( \40158 , \40147 , \40156 );
or \U$39815 ( \40159 , \40152 , \40157 , \40158 );
and \U$39816 ( \40160 , \27527 , \28063 );
and \U$39817 ( \40161 , \27325 , \28061 );
nor \U$39818 ( \40162 , \40160 , \40161 );
xnor \U$39819 ( \40163 , \40162 , \27803 );
and \U$39820 ( \40164 , \28002 , \27569 );
and \U$39821 ( \40165 , \27830 , \27567 );
nor \U$39822 ( \40166 , \40164 , \40165 );
xnor \U$39823 ( \40167 , \40166 , \27254 );
and \U$39824 ( \40168 , \40163 , \40167 );
and \U$39825 ( \40169 , \28952 , \27060 );
and \U$39826 ( \40170 , \28528 , \27058 );
nor \U$39827 ( \40171 , \40169 , \40170 );
xnor \U$39828 ( \40172 , \40171 , \26720 );
and \U$39829 ( \40173 , \40167 , \40172 );
and \U$39830 ( \40174 , \40163 , \40172 );
or \U$39831 ( \40175 , \40168 , \40173 , \40174 );
and \U$39832 ( \40176 , \40159 , \40175 );
and \U$39833 ( \40177 , \26078 , \29721 );
and \U$39834 ( \40178 , \26073 , \29719 );
nor \U$39835 ( \40179 , \40177 , \40178 );
xnor \U$39836 ( \40180 , \40179 , \29350 );
and \U$39837 ( \40181 , \26601 , \29159 );
and \U$39838 ( \40182 , \26342 , \29157 );
nor \U$39839 ( \40183 , \40181 , \40182 );
xnor \U$39840 ( \40184 , \40183 , \28841 );
and \U$39841 ( \40185 , \40180 , \40184 );
and \U$39842 ( \40186 , \26982 , \28592 );
and \U$39843 ( \40187 , \26973 , \28590 );
nor \U$39844 ( \40188 , \40186 , \40187 );
xnor \U$39845 ( \40189 , \40188 , \28343 );
and \U$39846 ( \40190 , \40184 , \40189 );
and \U$39847 ( \40191 , \40180 , \40189 );
or \U$39848 ( \40192 , \40185 , \40190 , \40191 );
and \U$39849 ( \40193 , \40175 , \40192 );
and \U$39850 ( \40194 , \40159 , \40192 );
or \U$39851 ( \40195 , \40176 , \40193 , \40194 );
xor \U$39852 ( \40196 , \40008 , \40012 );
xor \U$39853 ( \40197 , \40196 , \40017 );
xor \U$39854 ( \40198 , \40024 , \40028 );
xor \U$39855 ( \40199 , \40198 , \40033 );
and \U$39856 ( \40200 , \40197 , \40199 );
xor \U$39857 ( \40201 , \40056 , \40060 );
xor \U$39858 ( \40202 , \40201 , \40065 );
and \U$39859 ( \40203 , \40199 , \40202 );
and \U$39860 ( \40204 , \40197 , \40202 );
or \U$39861 ( \40205 , \40200 , \40203 , \40204 );
and \U$39862 ( \40206 , \40195 , \40205 );
and \U$39863 ( \40207 , \29203 , \26471 );
and \U$39864 ( \40208 , \29198 , \26469 );
nor \U$39865 ( \40209 , \40207 , \40208 );
xnor \U$39866 ( \40210 , \40209 , \26230 );
and \U$39867 ( \40211 , \29806 , \26005 );
and \U$39868 ( \40212 , \29522 , \26003 );
nor \U$39869 ( \40213 , \40211 , \40212 );
xnor \U$39870 ( \40214 , \40213 , \25817 );
and \U$39871 ( \40215 , \40210 , \40214 );
and \U$39872 ( \40216 , \30383 , \25631 );
and \U$39873 ( \40217 , \30375 , \25629 );
nor \U$39874 ( \40218 , \40216 , \40217 );
xnor \U$39875 ( \40219 , \40218 , \25399 );
and \U$39876 ( \40220 , \40214 , \40219 );
and \U$39877 ( \40221 , \40210 , \40219 );
or \U$39878 ( \40222 , \40215 , \40220 , \40221 );
nand \U$39879 ( \40223 , \31792 , \24460 );
xnor \U$39880 ( \40224 , \40223 , \24275 );
and \U$39881 ( \40225 , \40222 , \40224 );
xor \U$39882 ( \40226 , \40072 , \40076 );
xor \U$39883 ( \40227 , \40226 , \40081 );
and \U$39884 ( \40228 , \40224 , \40227 );
and \U$39885 ( \40229 , \40222 , \40227 );
or \U$39886 ( \40230 , \40225 , \40228 , \40229 );
and \U$39887 ( \40231 , \40205 , \40230 );
and \U$39888 ( \40232 , \40195 , \40230 );
or \U$39889 ( \40233 , \40206 , \40231 , \40232 );
xor \U$39890 ( \40234 , \39877 , \39881 );
xor \U$39891 ( \40235 , \40234 , \39886 );
xor \U$39892 ( \40236 , \40068 , \40084 );
xor \U$39893 ( \40237 , \40236 , \40087 );
and \U$39894 ( \40238 , \40235 , \40237 );
xor \U$39895 ( \40239 , \40093 , \40095 );
xor \U$39896 ( \40240 , \40239 , \40098 );
and \U$39897 ( \40241 , \40237 , \40240 );
and \U$39898 ( \40242 , \40235 , \40240 );
or \U$39899 ( \40243 , \40238 , \40241 , \40242 );
and \U$39900 ( \40244 , \40233 , \40243 );
xor \U$39901 ( \40245 , \39856 , \39872 );
xor \U$39902 ( \40246 , \40245 , \39889 );
and \U$39903 ( \40247 , \40243 , \40246 );
and \U$39904 ( \40248 , \40233 , \40246 );
or \U$39905 ( \40249 , \40244 , \40247 , \40248 );
xor \U$39906 ( \40250 , \40104 , \40114 );
xor \U$39907 ( \40251 , \40250 , \40117 );
and \U$39908 ( \40252 , \40249 , \40251 );
xor \U$39909 ( \40253 , \40122 , \40124 );
and \U$39910 ( \40254 , \40251 , \40253 );
and \U$39911 ( \40255 , \40249 , \40253 );
or \U$39912 ( \40256 , \40252 , \40254 , \40255 );
xor \U$39913 ( \40257 , \39946 , \39964 );
xor \U$39914 ( \40258 , \40257 , \39975 );
and \U$39915 ( \40259 , \40256 , \40258 );
xor \U$39916 ( \40260 , \40120 , \40125 );
xor \U$39917 ( \40261 , \40260 , \40128 );
and \U$39918 ( \40262 , \40258 , \40261 );
and \U$39919 ( \40263 , \40256 , \40261 );
or \U$39920 ( \40264 , \40259 , \40262 , \40263 );
and \U$39921 ( \40265 , \40143 , \40264 );
xor \U$39922 ( \40266 , \40143 , \40264 );
xor \U$39923 ( \40267 , \40256 , \40258 );
xor \U$39924 ( \40268 , \40267 , \40261 );
and \U$39925 ( \40269 , \29198 , \27060 );
and \U$39926 ( \40270 , \28952 , \27058 );
nor \U$39927 ( \40271 , \40269 , \40270 );
xnor \U$39928 ( \40272 , \40271 , \26720 );
and \U$39929 ( \40273 , \29522 , \26471 );
and \U$39930 ( \40274 , \29203 , \26469 );
nor \U$39931 ( \40275 , \40273 , \40274 );
xnor \U$39932 ( \40276 , \40275 , \26230 );
and \U$39933 ( \40277 , \40272 , \40276 );
and \U$39934 ( \40278 , \30375 , \26005 );
and \U$39935 ( \40279 , \29806 , \26003 );
nor \U$39936 ( \40280 , \40278 , \40279 );
xnor \U$39937 ( \40281 , \40280 , \25817 );
and \U$39938 ( \40282 , \40276 , \40281 );
and \U$39939 ( \40283 , \40272 , \40281 );
or \U$39940 ( \40284 , \40277 , \40282 , \40283 );
and \U$39941 ( \40285 , \30986 , \25631 );
and \U$39942 ( \40286 , \30383 , \25629 );
nor \U$39943 ( \40287 , \40285 , \40286 );
xnor \U$39944 ( \40288 , \40287 , \25399 );
and \U$39945 ( \40289 , \31172 , \25180 );
and \U$39946 ( \40290 , \30991 , \25178 );
nor \U$39947 ( \40291 , \40289 , \40290 );
xnor \U$39948 ( \40292 , \40291 , \25037 );
and \U$39949 ( \40293 , \40288 , \40292 );
nand \U$39950 ( \40294 , \31792 , \24855 );
xnor \U$39951 ( \40295 , \40294 , \24611 );
and \U$39952 ( \40296 , \40292 , \40295 );
and \U$39953 ( \40297 , \40288 , \40295 );
or \U$39954 ( \40298 , \40293 , \40296 , \40297 );
and \U$39955 ( \40299 , \40284 , \40298 );
and \U$39956 ( \40300 , \30991 , \25180 );
and \U$39957 ( \40301 , \30986 , \25178 );
nor \U$39958 ( \40302 , \40300 , \40301 );
xnor \U$39959 ( \40303 , \40302 , \25037 );
and \U$39960 ( \40304 , \40298 , \40303 );
and \U$39961 ( \40305 , \40284 , \40303 );
or \U$39962 ( \40306 , \40299 , \40304 , \40305 );
and \U$39963 ( \40307 , \27325 , \28592 );
and \U$39964 ( \40308 , \26982 , \28590 );
nor \U$39965 ( \40309 , \40307 , \40308 );
xnor \U$39966 ( \40310 , \40309 , \28343 );
and \U$39967 ( \40311 , \27830 , \28063 );
and \U$39968 ( \40312 , \27527 , \28061 );
nor \U$39969 ( \40313 , \40311 , \40312 );
xnor \U$39970 ( \40314 , \40313 , \27803 );
and \U$39971 ( \40315 , \40310 , \40314 );
and \U$39972 ( \40316 , \28528 , \27569 );
and \U$39973 ( \40317 , \28002 , \27567 );
nor \U$39974 ( \40318 , \40316 , \40317 );
xnor \U$39975 ( \40319 , \40318 , \27254 );
and \U$39976 ( \40320 , \40314 , \40319 );
and \U$39977 ( \40321 , \40310 , \40319 );
or \U$39978 ( \40322 , \40315 , \40320 , \40321 );
and \U$39979 ( \40323 , \25097 , \31639 );
and \U$39980 ( \40324 , \24841 , \31636 );
nor \U$39981 ( \40325 , \40323 , \40324 );
xnor \U$39982 ( \40326 , \40325 , \30584 );
and \U$39983 ( \40327 , \25596 , \30826 );
and \U$39984 ( \40328 , \25294 , \30824 );
nor \U$39985 ( \40329 , \40327 , \40328 );
xnor \U$39986 ( \40330 , \40329 , \30587 );
and \U$39987 ( \40331 , \40326 , \40330 );
and \U$39988 ( \40332 , \40330 , \24611 );
and \U$39989 ( \40333 , \40326 , \24611 );
or \U$39990 ( \40334 , \40331 , \40332 , \40333 );
and \U$39991 ( \40335 , \40322 , \40334 );
and \U$39992 ( \40336 , \26073 , \30258 );
and \U$39993 ( \40337 , \25604 , \30256 );
nor \U$39994 ( \40338 , \40336 , \40337 );
xnor \U$39995 ( \40339 , \40338 , \29948 );
and \U$39996 ( \40340 , \26342 , \29721 );
and \U$39997 ( \40341 , \26078 , \29719 );
nor \U$39998 ( \40342 , \40340 , \40341 );
xnor \U$39999 ( \40343 , \40342 , \29350 );
and \U$40000 ( \40344 , \40339 , \40343 );
and \U$40001 ( \40345 , \26973 , \29159 );
and \U$40002 ( \40346 , \26601 , \29157 );
nor \U$40003 ( \40347 , \40345 , \40346 );
xnor \U$40004 ( \40348 , \40347 , \28841 );
and \U$40005 ( \40349 , \40343 , \40348 );
and \U$40006 ( \40350 , \40339 , \40348 );
or \U$40007 ( \40351 , \40344 , \40349 , \40350 );
and \U$40008 ( \40352 , \40334 , \40351 );
and \U$40009 ( \40353 , \40322 , \40351 );
or \U$40010 ( \40354 , \40335 , \40352 , \40353 );
and \U$40011 ( \40355 , \40306 , \40354 );
and \U$40012 ( \40356 , \31792 , \24857 );
and \U$40013 ( \40357 , \31172 , \24855 );
nor \U$40014 ( \40358 , \40356 , \40357 );
xnor \U$40015 ( \40359 , \40358 , \24611 );
xor \U$40016 ( \40360 , \40210 , \40214 );
xor \U$40017 ( \40361 , \40360 , \40219 );
and \U$40018 ( \40362 , \40359 , \40361 );
xor \U$40019 ( \40363 , \40163 , \40167 );
xor \U$40020 ( \40364 , \40363 , \40172 );
and \U$40021 ( \40365 , \40361 , \40364 );
and \U$40022 ( \40366 , \40359 , \40364 );
or \U$40023 ( \40367 , \40362 , \40365 , \40366 );
and \U$40024 ( \40368 , \40354 , \40367 );
and \U$40025 ( \40369 , \40306 , \40367 );
or \U$40026 ( \40370 , \40355 , \40368 , \40369 );
xor \U$40027 ( \40371 , \40041 , \40045 );
xor \U$40028 ( \40372 , \40371 , \24275 );
xor \U$40029 ( \40373 , \40197 , \40199 );
xor \U$40030 ( \40374 , \40373 , \40202 );
and \U$40031 ( \40375 , \40372 , \40374 );
xor \U$40032 ( \40376 , \40222 , \40224 );
xor \U$40033 ( \40377 , \40376 , \40227 );
and \U$40034 ( \40378 , \40374 , \40377 );
and \U$40035 ( \40379 , \40372 , \40377 );
or \U$40036 ( \40380 , \40375 , \40378 , \40379 );
and \U$40037 ( \40381 , \40370 , \40380 );
xor \U$40038 ( \40382 , \40020 , \40036 );
xor \U$40039 ( \40383 , \40382 , \40049 );
and \U$40040 ( \40384 , \40380 , \40383 );
and \U$40041 ( \40385 , \40370 , \40383 );
or \U$40042 ( \40386 , \40381 , \40384 , \40385 );
xor \U$40043 ( \40387 , \40195 , \40205 );
xor \U$40044 ( \40388 , \40387 , \40230 );
xor \U$40045 ( \40389 , \40235 , \40237 );
xor \U$40046 ( \40390 , \40389 , \40240 );
and \U$40047 ( \40391 , \40388 , \40390 );
and \U$40048 ( \40392 , \40386 , \40391 );
xor \U$40049 ( \40393 , \40106 , \40108 );
xor \U$40050 ( \40394 , \40393 , \40111 );
and \U$40051 ( \40395 , \40391 , \40394 );
and \U$40052 ( \40396 , \40386 , \40394 );
or \U$40053 ( \40397 , \40392 , \40395 , \40396 );
xor \U$40054 ( \40398 , \40052 , \40090 );
xor \U$40055 ( \40399 , \40398 , \40101 );
xor \U$40056 ( \40400 , \40233 , \40243 );
xor \U$40057 ( \40401 , \40400 , \40246 );
and \U$40058 ( \40402 , \40399 , \40401 );
and \U$40059 ( \40403 , \40397 , \40402 );
xor \U$40060 ( \40404 , \40249 , \40251 );
xor \U$40061 ( \40405 , \40404 , \40253 );
and \U$40062 ( \40406 , \40402 , \40405 );
and \U$40063 ( \40407 , \40397 , \40405 );
or \U$40064 ( \40408 , \40403 , \40406 , \40407 );
and \U$40065 ( \40409 , \40268 , \40408 );
xor \U$40066 ( \40410 , \40268 , \40408 );
xor \U$40067 ( \40411 , \40397 , \40402 );
xor \U$40068 ( \40412 , \40411 , \40405 );
and \U$40069 ( \40413 , \26601 , \29721 );
and \U$40070 ( \40414 , \26342 , \29719 );
nor \U$40071 ( \40415 , \40413 , \40414 );
xnor \U$40072 ( \40416 , \40415 , \29350 );
and \U$40073 ( \40417 , \26982 , \29159 );
and \U$40074 ( \40418 , \26973 , \29157 );
nor \U$40075 ( \40419 , \40417 , \40418 );
xnor \U$40076 ( \40420 , \40419 , \28841 );
and \U$40077 ( \40421 , \40416 , \40420 );
and \U$40078 ( \40422 , \27527 , \28592 );
and \U$40079 ( \40423 , \27325 , \28590 );
nor \U$40080 ( \40424 , \40422 , \40423 );
xnor \U$40081 ( \40425 , \40424 , \28343 );
and \U$40082 ( \40426 , \40420 , \40425 );
and \U$40083 ( \40427 , \40416 , \40425 );
or \U$40084 ( \40428 , \40421 , \40426 , \40427 );
and \U$40085 ( \40429 , \25294 , \31639 );
and \U$40086 ( \40430 , \25097 , \31636 );
nor \U$40087 ( \40431 , \40429 , \40430 );
xnor \U$40088 ( \40432 , \40431 , \30584 );
and \U$40089 ( \40433 , \25604 , \30826 );
and \U$40090 ( \40434 , \25596 , \30824 );
nor \U$40091 ( \40435 , \40433 , \40434 );
xnor \U$40092 ( \40436 , \40435 , \30587 );
and \U$40093 ( \40437 , \40432 , \40436 );
and \U$40094 ( \40438 , \26078 , \30258 );
and \U$40095 ( \40439 , \26073 , \30256 );
nor \U$40096 ( \40440 , \40438 , \40439 );
xnor \U$40097 ( \40441 , \40440 , \29948 );
and \U$40098 ( \40442 , \40436 , \40441 );
and \U$40099 ( \40443 , \40432 , \40441 );
or \U$40100 ( \40444 , \40437 , \40442 , \40443 );
and \U$40101 ( \40445 , \40428 , \40444 );
and \U$40102 ( \40446 , \28002 , \28063 );
and \U$40103 ( \40447 , \27830 , \28061 );
nor \U$40104 ( \40448 , \40446 , \40447 );
xnor \U$40105 ( \40449 , \40448 , \27803 );
and \U$40106 ( \40450 , \28952 , \27569 );
and \U$40107 ( \40451 , \28528 , \27567 );
nor \U$40108 ( \40452 , \40450 , \40451 );
xnor \U$40109 ( \40453 , \40452 , \27254 );
and \U$40110 ( \40454 , \40449 , \40453 );
and \U$40111 ( \40455 , \29203 , \27060 );
and \U$40112 ( \40456 , \29198 , \27058 );
nor \U$40113 ( \40457 , \40455 , \40456 );
xnor \U$40114 ( \40458 , \40457 , \26720 );
and \U$40115 ( \40459 , \40453 , \40458 );
and \U$40116 ( \40460 , \40449 , \40458 );
or \U$40117 ( \40461 , \40454 , \40459 , \40460 );
and \U$40118 ( \40462 , \40444 , \40461 );
and \U$40119 ( \40463 , \40428 , \40461 );
or \U$40120 ( \40464 , \40445 , \40462 , \40463 );
xor \U$40121 ( \40465 , \40310 , \40314 );
xor \U$40122 ( \40466 , \40465 , \40319 );
xor \U$40123 ( \40467 , \40326 , \40330 );
xor \U$40124 ( \40468 , \40467 , \24611 );
and \U$40125 ( \40469 , \40466 , \40468 );
xor \U$40126 ( \40470 , \40339 , \40343 );
xor \U$40127 ( \40471 , \40470 , \40348 );
and \U$40128 ( \40472 , \40468 , \40471 );
and \U$40129 ( \40473 , \40466 , \40471 );
or \U$40130 ( \40474 , \40469 , \40472 , \40473 );
and \U$40131 ( \40475 , \40464 , \40474 );
and \U$40132 ( \40476 , \29806 , \26471 );
and \U$40133 ( \40477 , \29522 , \26469 );
nor \U$40134 ( \40478 , \40476 , \40477 );
xnor \U$40135 ( \40479 , \40478 , \26230 );
and \U$40136 ( \40480 , \30383 , \26005 );
and \U$40137 ( \40481 , \30375 , \26003 );
nor \U$40138 ( \40482 , \40480 , \40481 );
xnor \U$40139 ( \40483 , \40482 , \25817 );
and \U$40140 ( \40484 , \40479 , \40483 );
and \U$40141 ( \40485 , \30991 , \25631 );
and \U$40142 ( \40486 , \30986 , \25629 );
nor \U$40143 ( \40487 , \40485 , \40486 );
xnor \U$40144 ( \40488 , \40487 , \25399 );
and \U$40145 ( \40489 , \40483 , \40488 );
and \U$40146 ( \40490 , \40479 , \40488 );
or \U$40147 ( \40491 , \40484 , \40489 , \40490 );
xor \U$40148 ( \40492 , \40272 , \40276 );
xor \U$40149 ( \40493 , \40492 , \40281 );
and \U$40150 ( \40494 , \40491 , \40493 );
xor \U$40151 ( \40495 , \40288 , \40292 );
xor \U$40152 ( \40496 , \40495 , \40295 );
and \U$40153 ( \40497 , \40493 , \40496 );
and \U$40154 ( \40498 , \40491 , \40496 );
or \U$40155 ( \40499 , \40494 , \40497 , \40498 );
and \U$40156 ( \40500 , \40474 , \40499 );
and \U$40157 ( \40501 , \40464 , \40499 );
or \U$40158 ( \40502 , \40475 , \40500 , \40501 );
xor \U$40159 ( \40503 , \40147 , \40151 );
xor \U$40160 ( \40504 , \40503 , \40156 );
xor \U$40161 ( \40505 , \40180 , \40184 );
xor \U$40162 ( \40506 , \40505 , \40189 );
and \U$40163 ( \40507 , \40504 , \40506 );
xor \U$40164 ( \40508 , \40359 , \40361 );
xor \U$40165 ( \40509 , \40508 , \40364 );
and \U$40166 ( \40510 , \40506 , \40509 );
and \U$40167 ( \40511 , \40504 , \40509 );
or \U$40168 ( \40512 , \40507 , \40510 , \40511 );
and \U$40169 ( \40513 , \40502 , \40512 );
xor \U$40170 ( \40514 , \40159 , \40175 );
xor \U$40171 ( \40515 , \40514 , \40192 );
and \U$40172 ( \40516 , \40512 , \40515 );
and \U$40173 ( \40517 , \40502 , \40515 );
or \U$40174 ( \40518 , \40513 , \40516 , \40517 );
xor \U$40175 ( \40519 , \40370 , \40380 );
xor \U$40176 ( \40520 , \40519 , \40383 );
and \U$40177 ( \40521 , \40518 , \40520 );
xor \U$40178 ( \40522 , \40388 , \40390 );
and \U$40179 ( \40523 , \40520 , \40522 );
and \U$40180 ( \40524 , \40518 , \40522 );
or \U$40181 ( \40525 , \40521 , \40523 , \40524 );
xor \U$40182 ( \40526 , \40386 , \40391 );
xor \U$40183 ( \40527 , \40526 , \40394 );
and \U$40184 ( \40528 , \40525 , \40527 );
xor \U$40185 ( \40529 , \40399 , \40401 );
and \U$40186 ( \40530 , \40527 , \40529 );
and \U$40187 ( \40531 , \40525 , \40529 );
or \U$40188 ( \40532 , \40528 , \40530 , \40531 );
and \U$40189 ( \40533 , \40412 , \40532 );
xor \U$40190 ( \40534 , \40412 , \40532 );
xor \U$40191 ( \40535 , \40525 , \40527 );
xor \U$40192 ( \40536 , \40535 , \40529 );
and \U$40193 ( \40537 , \26342 , \30258 );
and \U$40194 ( \40538 , \26078 , \30256 );
nor \U$40195 ( \40539 , \40537 , \40538 );
xnor \U$40196 ( \40540 , \40539 , \29948 );
and \U$40197 ( \40541 , \26973 , \29721 );
and \U$40198 ( \40542 , \26601 , \29719 );
nor \U$40199 ( \40543 , \40541 , \40542 );
xnor \U$40200 ( \40544 , \40543 , \29350 );
and \U$40201 ( \40545 , \40540 , \40544 );
and \U$40202 ( \40546 , \27325 , \29159 );
and \U$40203 ( \40547 , \26982 , \29157 );
nor \U$40204 ( \40548 , \40546 , \40547 );
xnor \U$40205 ( \40549 , \40548 , \28841 );
and \U$40206 ( \40550 , \40544 , \40549 );
and \U$40207 ( \40551 , \40540 , \40549 );
or \U$40208 ( \40552 , \40545 , \40550 , \40551 );
and \U$40209 ( \40553 , \25596 , \31639 );
and \U$40210 ( \40554 , \25294 , \31636 );
nor \U$40211 ( \40555 , \40553 , \40554 );
xnor \U$40212 ( \40556 , \40555 , \30584 );
and \U$40213 ( \40557 , \26073 , \30826 );
and \U$40214 ( \40558 , \25604 , \30824 );
nor \U$40215 ( \40559 , \40557 , \40558 );
xnor \U$40216 ( \40560 , \40559 , \30587 );
and \U$40217 ( \40561 , \40556 , \40560 );
and \U$40218 ( \40562 , \40560 , \25037 );
and \U$40219 ( \40563 , \40556 , \25037 );
or \U$40220 ( \40564 , \40561 , \40562 , \40563 );
and \U$40221 ( \40565 , \40552 , \40564 );
and \U$40222 ( \40566 , \27830 , \28592 );
and \U$40223 ( \40567 , \27527 , \28590 );
nor \U$40224 ( \40568 , \40566 , \40567 );
xnor \U$40225 ( \40569 , \40568 , \28343 );
and \U$40226 ( \40570 , \28528 , \28063 );
and \U$40227 ( \40571 , \28002 , \28061 );
nor \U$40228 ( \40572 , \40570 , \40571 );
xnor \U$40229 ( \40573 , \40572 , \27803 );
and \U$40230 ( \40574 , \40569 , \40573 );
and \U$40231 ( \40575 , \29198 , \27569 );
and \U$40232 ( \40576 , \28952 , \27567 );
nor \U$40233 ( \40577 , \40575 , \40576 );
xnor \U$40234 ( \40578 , \40577 , \27254 );
and \U$40235 ( \40579 , \40573 , \40578 );
and \U$40236 ( \40580 , \40569 , \40578 );
or \U$40237 ( \40581 , \40574 , \40579 , \40580 );
and \U$40238 ( \40582 , \40564 , \40581 );
and \U$40239 ( \40583 , \40552 , \40581 );
or \U$40240 ( \40584 , \40565 , \40582 , \40583 );
and \U$40241 ( \40585 , \29522 , \27060 );
and \U$40242 ( \40586 , \29203 , \27058 );
nor \U$40243 ( \40587 , \40585 , \40586 );
xnor \U$40244 ( \40588 , \40587 , \26720 );
and \U$40245 ( \40589 , \30375 , \26471 );
and \U$40246 ( \40590 , \29806 , \26469 );
nor \U$40247 ( \40591 , \40589 , \40590 );
xnor \U$40248 ( \40592 , \40591 , \26230 );
and \U$40249 ( \40593 , \40588 , \40592 );
and \U$40250 ( \40594 , \30986 , \26005 );
and \U$40251 ( \40595 , \30383 , \26003 );
nor \U$40252 ( \40596 , \40594 , \40595 );
xnor \U$40253 ( \40597 , \40596 , \25817 );
and \U$40254 ( \40598 , \40592 , \40597 );
and \U$40255 ( \40599 , \40588 , \40597 );
or \U$40256 ( \40600 , \40593 , \40598 , \40599 );
and \U$40257 ( \40601 , \31172 , \25631 );
and \U$40258 ( \40602 , \30991 , \25629 );
nor \U$40259 ( \40603 , \40601 , \40602 );
xnor \U$40260 ( \40604 , \40603 , \25399 );
nand \U$40261 ( \40605 , \31792 , \25178 );
xnor \U$40262 ( \40606 , \40605 , \25037 );
and \U$40263 ( \40607 , \40604 , \40606 );
and \U$40264 ( \40608 , \40600 , \40607 );
and \U$40265 ( \40609 , \31792 , \25180 );
and \U$40266 ( \40610 , \31172 , \25178 );
nor \U$40267 ( \40611 , \40609 , \40610 );
xnor \U$40268 ( \40612 , \40611 , \25037 );
and \U$40269 ( \40613 , \40607 , \40612 );
and \U$40270 ( \40614 , \40600 , \40612 );
or \U$40271 ( \40615 , \40608 , \40613 , \40614 );
and \U$40272 ( \40616 , \40584 , \40615 );
xor \U$40273 ( \40617 , \40416 , \40420 );
xor \U$40274 ( \40618 , \40617 , \40425 );
xor \U$40275 ( \40619 , \40479 , \40483 );
xor \U$40276 ( \40620 , \40619 , \40488 );
and \U$40277 ( \40621 , \40618 , \40620 );
xor \U$40278 ( \40622 , \40449 , \40453 );
xor \U$40279 ( \40623 , \40622 , \40458 );
and \U$40280 ( \40624 , \40620 , \40623 );
and \U$40281 ( \40625 , \40618 , \40623 );
or \U$40282 ( \40626 , \40621 , \40624 , \40625 );
and \U$40283 ( \40627 , \40615 , \40626 );
and \U$40284 ( \40628 , \40584 , \40626 );
or \U$40285 ( \40629 , \40616 , \40627 , \40628 );
xor \U$40286 ( \40630 , \40428 , \40444 );
xor \U$40287 ( \40631 , \40630 , \40461 );
xor \U$40288 ( \40632 , \40466 , \40468 );
xor \U$40289 ( \40633 , \40632 , \40471 );
and \U$40290 ( \40634 , \40631 , \40633 );
xor \U$40291 ( \40635 , \40491 , \40493 );
xor \U$40292 ( \40636 , \40635 , \40496 );
and \U$40293 ( \40637 , \40633 , \40636 );
and \U$40294 ( \40638 , \40631 , \40636 );
or \U$40295 ( \40639 , \40634 , \40637 , \40638 );
and \U$40296 ( \40640 , \40629 , \40639 );
xor \U$40297 ( \40641 , \40284 , \40298 );
xor \U$40298 ( \40642 , \40641 , \40303 );
and \U$40299 ( \40643 , \40639 , \40642 );
and \U$40300 ( \40644 , \40629 , \40642 );
or \U$40301 ( \40645 , \40640 , \40643 , \40644 );
xor \U$40302 ( \40646 , \40322 , \40334 );
xor \U$40303 ( \40647 , \40646 , \40351 );
xor \U$40304 ( \40648 , \40464 , \40474 );
xor \U$40305 ( \40649 , \40648 , \40499 );
and \U$40306 ( \40650 , \40647 , \40649 );
xor \U$40307 ( \40651 , \40504 , \40506 );
xor \U$40308 ( \40652 , \40651 , \40509 );
and \U$40309 ( \40653 , \40649 , \40652 );
and \U$40310 ( \40654 , \40647 , \40652 );
or \U$40311 ( \40655 , \40650 , \40653 , \40654 );
and \U$40312 ( \40656 , \40645 , \40655 );
xor \U$40313 ( \40657 , \40372 , \40374 );
xor \U$40314 ( \40658 , \40657 , \40377 );
and \U$40315 ( \40659 , \40655 , \40658 );
and \U$40316 ( \40660 , \40645 , \40658 );
or \U$40317 ( \40661 , \40656 , \40659 , \40660 );
xor \U$40318 ( \40662 , \40306 , \40354 );
xor \U$40319 ( \40663 , \40662 , \40367 );
xor \U$40320 ( \40664 , \40502 , \40512 );
xor \U$40321 ( \40665 , \40664 , \40515 );
and \U$40322 ( \40666 , \40663 , \40665 );
and \U$40323 ( \40667 , \40661 , \40666 );
xor \U$40324 ( \40668 , \40518 , \40520 );
xor \U$40325 ( \40669 , \40668 , \40522 );
and \U$40326 ( \40670 , \40666 , \40669 );
and \U$40327 ( \40671 , \40661 , \40669 );
or \U$40328 ( \40672 , \40667 , \40670 , \40671 );
and \U$40329 ( \40673 , \40536 , \40672 );
xor \U$40330 ( \40674 , \40536 , \40672 );
xor \U$40331 ( \40675 , \40661 , \40666 );
xor \U$40332 ( \40676 , \40675 , \40669 );
and \U$40333 ( \40677 , \26982 , \29721 );
and \U$40334 ( \40678 , \26973 , \29719 );
nor \U$40335 ( \40679 , \40677 , \40678 );
xnor \U$40336 ( \40680 , \40679 , \29350 );
and \U$40337 ( \40681 , \27527 , \29159 );
and \U$40338 ( \40682 , \27325 , \29157 );
nor \U$40339 ( \40683 , \40681 , \40682 );
xnor \U$40340 ( \40684 , \40683 , \28841 );
and \U$40341 ( \40685 , \40680 , \40684 );
and \U$40342 ( \40686 , \28002 , \28592 );
and \U$40343 ( \40687 , \27830 , \28590 );
nor \U$40344 ( \40688 , \40686 , \40687 );
xnor \U$40345 ( \40689 , \40688 , \28343 );
and \U$40346 ( \40690 , \40684 , \40689 );
and \U$40347 ( \40691 , \40680 , \40689 );
or \U$40348 ( \40692 , \40685 , \40690 , \40691 );
and \U$40349 ( \40693 , \28952 , \28063 );
and \U$40350 ( \40694 , \28528 , \28061 );
nor \U$40351 ( \40695 , \40693 , \40694 );
xnor \U$40352 ( \40696 , \40695 , \27803 );
and \U$40353 ( \40697 , \29203 , \27569 );
and \U$40354 ( \40698 , \29198 , \27567 );
nor \U$40355 ( \40699 , \40697 , \40698 );
xnor \U$40356 ( \40700 , \40699 , \27254 );
and \U$40357 ( \40701 , \40696 , \40700 );
and \U$40358 ( \40702 , \29806 , \27060 );
and \U$40359 ( \40703 , \29522 , \27058 );
nor \U$40360 ( \40704 , \40702 , \40703 );
xnor \U$40361 ( \40705 , \40704 , \26720 );
and \U$40362 ( \40706 , \40700 , \40705 );
and \U$40363 ( \40707 , \40696 , \40705 );
or \U$40364 ( \40708 , \40701 , \40706 , \40707 );
and \U$40365 ( \40709 , \40692 , \40708 );
and \U$40366 ( \40710 , \25604 , \31639 );
and \U$40367 ( \40711 , \25596 , \31636 );
nor \U$40368 ( \40712 , \40710 , \40711 );
xnor \U$40369 ( \40713 , \40712 , \30584 );
and \U$40370 ( \40714 , \26078 , \30826 );
and \U$40371 ( \40715 , \26073 , \30824 );
nor \U$40372 ( \40716 , \40714 , \40715 );
xnor \U$40373 ( \40717 , \40716 , \30587 );
and \U$40374 ( \40718 , \40713 , \40717 );
and \U$40375 ( \40719 , \26601 , \30258 );
and \U$40376 ( \40720 , \26342 , \30256 );
nor \U$40377 ( \40721 , \40719 , \40720 );
xnor \U$40378 ( \40722 , \40721 , \29948 );
and \U$40379 ( \40723 , \40717 , \40722 );
and \U$40380 ( \40724 , \40713 , \40722 );
or \U$40381 ( \40725 , \40718 , \40723 , \40724 );
and \U$40382 ( \40726 , \40708 , \40725 );
and \U$40383 ( \40727 , \40692 , \40725 );
or \U$40384 ( \40728 , \40709 , \40726 , \40727 );
xor \U$40385 ( \40729 , \40540 , \40544 );
xor \U$40386 ( \40730 , \40729 , \40549 );
xor \U$40387 ( \40731 , \40556 , \40560 );
xor \U$40388 ( \40732 , \40731 , \25037 );
and \U$40389 ( \40733 , \40730 , \40732 );
xor \U$40390 ( \40734 , \40569 , \40573 );
xor \U$40391 ( \40735 , \40734 , \40578 );
and \U$40392 ( \40736 , \40732 , \40735 );
and \U$40393 ( \40737 , \40730 , \40735 );
or \U$40394 ( \40738 , \40733 , \40736 , \40737 );
and \U$40395 ( \40739 , \40728 , \40738 );
and \U$40396 ( \40740 , \30383 , \26471 );
and \U$40397 ( \40741 , \30375 , \26469 );
nor \U$40398 ( \40742 , \40740 , \40741 );
xnor \U$40399 ( \40743 , \40742 , \26230 );
and \U$40400 ( \40744 , \30991 , \26005 );
and \U$40401 ( \40745 , \30986 , \26003 );
nor \U$40402 ( \40746 , \40744 , \40745 );
xnor \U$40403 ( \40747 , \40746 , \25817 );
and \U$40404 ( \40748 , \40743 , \40747 );
and \U$40405 ( \40749 , \31792 , \25631 );
and \U$40406 ( \40750 , \31172 , \25629 );
nor \U$40407 ( \40751 , \40749 , \40750 );
xnor \U$40408 ( \40752 , \40751 , \25399 );
and \U$40409 ( \40753 , \40747 , \40752 );
and \U$40410 ( \40754 , \40743 , \40752 );
or \U$40411 ( \40755 , \40748 , \40753 , \40754 );
xor \U$40412 ( \40756 , \40588 , \40592 );
xor \U$40413 ( \40757 , \40756 , \40597 );
and \U$40414 ( \40758 , \40755 , \40757 );
xor \U$40415 ( \40759 , \40604 , \40606 );
and \U$40416 ( \40760 , \40757 , \40759 );
and \U$40417 ( \40761 , \40755 , \40759 );
or \U$40418 ( \40762 , \40758 , \40760 , \40761 );
and \U$40419 ( \40763 , \40738 , \40762 );
and \U$40420 ( \40764 , \40728 , \40762 );
or \U$40421 ( \40765 , \40739 , \40763 , \40764 );
xor \U$40422 ( \40766 , \40432 , \40436 );
xor \U$40423 ( \40767 , \40766 , \40441 );
xor \U$40424 ( \40768 , \40600 , \40607 );
xor \U$40425 ( \40769 , \40768 , \40612 );
and \U$40426 ( \40770 , \40767 , \40769 );
xor \U$40427 ( \40771 , \40618 , \40620 );
xor \U$40428 ( \40772 , \40771 , \40623 );
and \U$40429 ( \40773 , \40769 , \40772 );
and \U$40430 ( \40774 , \40767 , \40772 );
or \U$40431 ( \40775 , \40770 , \40773 , \40774 );
and \U$40432 ( \40776 , \40765 , \40775 );
xor \U$40433 ( \40777 , \40631 , \40633 );
xor \U$40434 ( \40778 , \40777 , \40636 );
and \U$40435 ( \40779 , \40775 , \40778 );
and \U$40436 ( \40780 , \40765 , \40778 );
or \U$40437 ( \40781 , \40776 , \40779 , \40780 );
xor \U$40438 ( \40782 , \40629 , \40639 );
xor \U$40439 ( \40783 , \40782 , \40642 );
and \U$40440 ( \40784 , \40781 , \40783 );
xor \U$40441 ( \40785 , \40647 , \40649 );
xor \U$40442 ( \40786 , \40785 , \40652 );
and \U$40443 ( \40787 , \40783 , \40786 );
and \U$40444 ( \40788 , \40781 , \40786 );
or \U$40445 ( \40789 , \40784 , \40787 , \40788 );
xor \U$40446 ( \40790 , \40645 , \40655 );
xor \U$40447 ( \40791 , \40790 , \40658 );
and \U$40448 ( \40792 , \40789 , \40791 );
xor \U$40449 ( \40793 , \40663 , \40665 );
and \U$40450 ( \40794 , \40791 , \40793 );
and \U$40451 ( \40795 , \40789 , \40793 );
or \U$40452 ( \40796 , \40792 , \40794 , \40795 );
and \U$40453 ( \40797 , \40676 , \40796 );
xor \U$40454 ( \40798 , \40676 , \40796 );
xor \U$40455 ( \40799 , \40789 , \40791 );
xor \U$40456 ( \40800 , \40799 , \40793 );
and \U$40457 ( \40801 , \26973 , \30258 );
and \U$40458 ( \40802 , \26601 , \30256 );
nor \U$40459 ( \40803 , \40801 , \40802 );
xnor \U$40460 ( \40804 , \40803 , \29948 );
and \U$40461 ( \40805 , \27325 , \29721 );
and \U$40462 ( \40806 , \26982 , \29719 );
nor \U$40463 ( \40807 , \40805 , \40806 );
xnor \U$40464 ( \40808 , \40807 , \29350 );
and \U$40465 ( \40809 , \40804 , \40808 );
and \U$40466 ( \40810 , \27830 , \29159 );
and \U$40467 ( \40811 , \27527 , \29157 );
nor \U$40468 ( \40812 , \40810 , \40811 );
xnor \U$40469 ( \40813 , \40812 , \28841 );
and \U$40470 ( \40814 , \40808 , \40813 );
and \U$40471 ( \40815 , \40804 , \40813 );
or \U$40472 ( \40816 , \40809 , \40814 , \40815 );
and \U$40473 ( \40817 , \28528 , \28592 );
and \U$40474 ( \40818 , \28002 , \28590 );
nor \U$40475 ( \40819 , \40817 , \40818 );
xnor \U$40476 ( \40820 , \40819 , \28343 );
and \U$40477 ( \40821 , \29198 , \28063 );
and \U$40478 ( \40822 , \28952 , \28061 );
nor \U$40479 ( \40823 , \40821 , \40822 );
xnor \U$40480 ( \40824 , \40823 , \27803 );
and \U$40481 ( \40825 , \40820 , \40824 );
and \U$40482 ( \40826 , \29522 , \27569 );
and \U$40483 ( \40827 , \29203 , \27567 );
nor \U$40484 ( \40828 , \40826 , \40827 );
xnor \U$40485 ( \40829 , \40828 , \27254 );
and \U$40486 ( \40830 , \40824 , \40829 );
and \U$40487 ( \40831 , \40820 , \40829 );
or \U$40488 ( \40832 , \40825 , \40830 , \40831 );
and \U$40489 ( \40833 , \40816 , \40832 );
and \U$40490 ( \40834 , \26073 , \31639 );
and \U$40491 ( \40835 , \25604 , \31636 );
nor \U$40492 ( \40836 , \40834 , \40835 );
xnor \U$40493 ( \40837 , \40836 , \30584 );
and \U$40494 ( \40838 , \26342 , \30826 );
and \U$40495 ( \40839 , \26078 , \30824 );
nor \U$40496 ( \40840 , \40838 , \40839 );
xnor \U$40497 ( \40841 , \40840 , \30587 );
and \U$40498 ( \40842 , \40837 , \40841 );
and \U$40499 ( \40843 , \40841 , \25399 );
and \U$40500 ( \40844 , \40837 , \25399 );
or \U$40501 ( \40845 , \40842 , \40843 , \40844 );
and \U$40502 ( \40846 , \40832 , \40845 );
and \U$40503 ( \40847 , \40816 , \40845 );
or \U$40504 ( \40848 , \40833 , \40846 , \40847 );
and \U$40505 ( \40849 , \30375 , \27060 );
and \U$40506 ( \40850 , \29806 , \27058 );
nor \U$40507 ( \40851 , \40849 , \40850 );
xnor \U$40508 ( \40852 , \40851 , \26720 );
and \U$40509 ( \40853 , \30986 , \26471 );
and \U$40510 ( \40854 , \30383 , \26469 );
nor \U$40511 ( \40855 , \40853 , \40854 );
xnor \U$40512 ( \40856 , \40855 , \26230 );
and \U$40513 ( \40857 , \40852 , \40856 );
and \U$40514 ( \40858 , \31172 , \26005 );
and \U$40515 ( \40859 , \30991 , \26003 );
nor \U$40516 ( \40860 , \40858 , \40859 );
xnor \U$40517 ( \40861 , \40860 , \25817 );
and \U$40518 ( \40862 , \40856 , \40861 );
and \U$40519 ( \40863 , \40852 , \40861 );
or \U$40520 ( \40864 , \40857 , \40862 , \40863 );
xor \U$40521 ( \40865 , \40696 , \40700 );
xor \U$40522 ( \40866 , \40865 , \40705 );
and \U$40523 ( \40867 , \40864 , \40866 );
xor \U$40524 ( \40868 , \40743 , \40747 );
xor \U$40525 ( \40869 , \40868 , \40752 );
and \U$40526 ( \40870 , \40866 , \40869 );
and \U$40527 ( \40871 , \40864 , \40869 );
or \U$40528 ( \40872 , \40867 , \40870 , \40871 );
and \U$40529 ( \40873 , \40848 , \40872 );
xor \U$40530 ( \40874 , \40680 , \40684 );
xor \U$40531 ( \40875 , \40874 , \40689 );
xor \U$40532 ( \40876 , \40713 , \40717 );
xor \U$40533 ( \40877 , \40876 , \40722 );
and \U$40534 ( \40878 , \40875 , \40877 );
and \U$40535 ( \40879 , \40872 , \40878 );
and \U$40536 ( \40880 , \40848 , \40878 );
or \U$40537 ( \40881 , \40873 , \40879 , \40880 );
xor \U$40538 ( \40882 , \40692 , \40708 );
xor \U$40539 ( \40883 , \40882 , \40725 );
xor \U$40540 ( \40884 , \40730 , \40732 );
xor \U$40541 ( \40885 , \40884 , \40735 );
and \U$40542 ( \40886 , \40883 , \40885 );
xor \U$40543 ( \40887 , \40755 , \40757 );
xor \U$40544 ( \40888 , \40887 , \40759 );
and \U$40545 ( \40889 , \40885 , \40888 );
and \U$40546 ( \40890 , \40883 , \40888 );
or \U$40547 ( \40891 , \40886 , \40889 , \40890 );
and \U$40548 ( \40892 , \40881 , \40891 );
xor \U$40549 ( \40893 , \40552 , \40564 );
xor \U$40550 ( \40894 , \40893 , \40581 );
and \U$40551 ( \40895 , \40891 , \40894 );
and \U$40552 ( \40896 , \40881 , \40894 );
or \U$40553 ( \40897 , \40892 , \40895 , \40896 );
xor \U$40554 ( \40898 , \40728 , \40738 );
xor \U$40555 ( \40899 , \40898 , \40762 );
xor \U$40556 ( \40900 , \40767 , \40769 );
xor \U$40557 ( \40901 , \40900 , \40772 );
and \U$40558 ( \40902 , \40899 , \40901 );
and \U$40559 ( \40903 , \40897 , \40902 );
xor \U$40560 ( \40904 , \40584 , \40615 );
xor \U$40561 ( \40905 , \40904 , \40626 );
and \U$40562 ( \40906 , \40902 , \40905 );
and \U$40563 ( \40907 , \40897 , \40905 );
or \U$40564 ( \40908 , \40903 , \40906 , \40907 );
xor \U$40565 ( \40909 , \40781 , \40783 );
xor \U$40566 ( \40910 , \40909 , \40786 );
and \U$40567 ( \40911 , \40908 , \40910 );
and \U$40568 ( \40912 , \40800 , \40911 );
xor \U$40569 ( \40913 , \40800 , \40911 );
xor \U$40570 ( \40914 , \40908 , \40910 );
xor \U$40571 ( \40915 , \40897 , \40902 );
xor \U$40572 ( \40916 , \40915 , \40905 );
xor \U$40573 ( \40917 , \40765 , \40775 );
xor \U$40574 ( \40918 , \40917 , \40778 );
and \U$40575 ( \40919 , \40916 , \40918 );
and \U$40576 ( \40920 , \40914 , \40919 );
xor \U$40577 ( \40921 , \40914 , \40919 );
xor \U$40578 ( \40922 , \40916 , \40918 );
and \U$40579 ( \40923 , \26078 , \31639 );
and \U$40580 ( \40924 , \26073 , \31636 );
nor \U$40581 ( \40925 , \40923 , \40924 );
xnor \U$40582 ( \40926 , \40925 , \30584 );
and \U$40583 ( \40927 , \26601 , \30826 );
and \U$40584 ( \40928 , \26342 , \30824 );
nor \U$40585 ( \40929 , \40927 , \40928 );
xnor \U$40586 ( \40930 , \40929 , \30587 );
and \U$40587 ( \40931 , \40926 , \40930 );
and \U$40588 ( \40932 , \26982 , \30258 );
and \U$40589 ( \40933 , \26973 , \30256 );
nor \U$40590 ( \40934 , \40932 , \40933 );
xnor \U$40591 ( \40935 , \40934 , \29948 );
and \U$40592 ( \40936 , \40930 , \40935 );
and \U$40593 ( \40937 , \40926 , \40935 );
or \U$40594 ( \40938 , \40931 , \40936 , \40937 );
and \U$40595 ( \40939 , \29203 , \28063 );
and \U$40596 ( \40940 , \29198 , \28061 );
nor \U$40597 ( \40941 , \40939 , \40940 );
xnor \U$40598 ( \40942 , \40941 , \27803 );
and \U$40599 ( \40943 , \29806 , \27569 );
and \U$40600 ( \40944 , \29522 , \27567 );
nor \U$40601 ( \40945 , \40943 , \40944 );
xnor \U$40602 ( \40946 , \40945 , \27254 );
and \U$40603 ( \40947 , \40942 , \40946 );
and \U$40604 ( \40948 , \30383 , \27060 );
and \U$40605 ( \40949 , \30375 , \27058 );
nor \U$40606 ( \40950 , \40948 , \40949 );
xnor \U$40607 ( \40951 , \40950 , \26720 );
and \U$40608 ( \40952 , \40946 , \40951 );
and \U$40609 ( \40953 , \40942 , \40951 );
or \U$40610 ( \40954 , \40947 , \40952 , \40953 );
and \U$40611 ( \40955 , \40938 , \40954 );
and \U$40612 ( \40956 , \27527 , \29721 );
and \U$40613 ( \40957 , \27325 , \29719 );
nor \U$40614 ( \40958 , \40956 , \40957 );
xnor \U$40615 ( \40959 , \40958 , \29350 );
and \U$40616 ( \40960 , \28002 , \29159 );
and \U$40617 ( \40961 , \27830 , \29157 );
nor \U$40618 ( \40962 , \40960 , \40961 );
xnor \U$40619 ( \40963 , \40962 , \28841 );
and \U$40620 ( \40964 , \40959 , \40963 );
and \U$40621 ( \40965 , \28952 , \28592 );
and \U$40622 ( \40966 , \28528 , \28590 );
nor \U$40623 ( \40967 , \40965 , \40966 );
xnor \U$40624 ( \40968 , \40967 , \28343 );
and \U$40625 ( \40969 , \40963 , \40968 );
and \U$40626 ( \40970 , \40959 , \40968 );
or \U$40627 ( \40971 , \40964 , \40969 , \40970 );
and \U$40628 ( \40972 , \40954 , \40971 );
and \U$40629 ( \40973 , \40938 , \40971 );
or \U$40630 ( \40974 , \40955 , \40972 , \40973 );
nand \U$40631 ( \40975 , \31792 , \25629 );
xnor \U$40632 ( \40976 , \40975 , \25399 );
xor \U$40633 ( \40977 , \40820 , \40824 );
xor \U$40634 ( \40978 , \40977 , \40829 );
and \U$40635 ( \40979 , \40976 , \40978 );
xor \U$40636 ( \40980 , \40852 , \40856 );
xor \U$40637 ( \40981 , \40980 , \40861 );
and \U$40638 ( \40982 , \40978 , \40981 );
and \U$40639 ( \40983 , \40976 , \40981 );
or \U$40640 ( \40984 , \40979 , \40982 , \40983 );
and \U$40641 ( \40985 , \40974 , \40984 );
xor \U$40642 ( \40986 , \40804 , \40808 );
xor \U$40643 ( \40987 , \40986 , \40813 );
xor \U$40644 ( \40988 , \40837 , \40841 );
xor \U$40645 ( \40989 , \40988 , \25399 );
and \U$40646 ( \40990 , \40987 , \40989 );
and \U$40647 ( \40991 , \40984 , \40990 );
and \U$40648 ( \40992 , \40974 , \40990 );
or \U$40649 ( \40993 , \40985 , \40991 , \40992 );
xor \U$40650 ( \40994 , \40816 , \40832 );
xor \U$40651 ( \40995 , \40994 , \40845 );
xor \U$40652 ( \40996 , \40864 , \40866 );
xor \U$40653 ( \40997 , \40996 , \40869 );
and \U$40654 ( \40998 , \40995 , \40997 );
xor \U$40655 ( \40999 , \40875 , \40877 );
and \U$40656 ( \41000 , \40997 , \40999 );
and \U$40657 ( \41001 , \40995 , \40999 );
or \U$40658 ( \41002 , \40998 , \41000 , \41001 );
and \U$40659 ( \41003 , \40993 , \41002 );
xor \U$40660 ( \41004 , \40883 , \40885 );
xor \U$40661 ( \41005 , \41004 , \40888 );
and \U$40662 ( \41006 , \41002 , \41005 );
and \U$40663 ( \41007 , \40993 , \41005 );
or \U$40664 ( \41008 , \41003 , \41006 , \41007 );
xor \U$40665 ( \41009 , \40881 , \40891 );
xor \U$40666 ( \41010 , \41009 , \40894 );
and \U$40667 ( \41011 , \41008 , \41010 );
xor \U$40668 ( \41012 , \40899 , \40901 );
and \U$40669 ( \41013 , \41010 , \41012 );
and \U$40670 ( \41014 , \41008 , \41012 );
or \U$40671 ( \41015 , \41011 , \41013 , \41014 );
and \U$40672 ( \41016 , \40922 , \41015 );
xor \U$40673 ( \41017 , \40922 , \41015 );
xor \U$40674 ( \41018 , \41008 , \41010 );
xor \U$40675 ( \41019 , \41018 , \41012 );
and \U$40676 ( \41020 , \30986 , \27060 );
and \U$40677 ( \41021 , \30383 , \27058 );
nor \U$40678 ( \41022 , \41020 , \41021 );
xnor \U$40679 ( \41023 , \41022 , \26720 );
and \U$40680 ( \41024 , \31172 , \26471 );
and \U$40681 ( \41025 , \30991 , \26469 );
nor \U$40682 ( \41026 , \41024 , \41025 );
xnor \U$40683 ( \41027 , \41026 , \26230 );
and \U$40684 ( \41028 , \41023 , \41027 );
nand \U$40685 ( \41029 , \31792 , \26003 );
xnor \U$40686 ( \41030 , \41029 , \25817 );
and \U$40687 ( \41031 , \41027 , \41030 );
and \U$40688 ( \41032 , \41023 , \41030 );
or \U$40689 ( \41033 , \41028 , \41031 , \41032 );
and \U$40690 ( \41034 , \30991 , \26471 );
and \U$40691 ( \41035 , \30986 , \26469 );
nor \U$40692 ( \41036 , \41034 , \41035 );
xnor \U$40693 ( \41037 , \41036 , \26230 );
and \U$40694 ( \41038 , \41033 , \41037 );
and \U$40695 ( \41039 , \31792 , \26005 );
and \U$40696 ( \41040 , \31172 , \26003 );
nor \U$40697 ( \41041 , \41039 , \41040 );
xnor \U$40698 ( \41042 , \41041 , \25817 );
and \U$40699 ( \41043 , \41037 , \41042 );
and \U$40700 ( \41044 , \41033 , \41042 );
or \U$40701 ( \41045 , \41038 , \41043 , \41044 );
and \U$40702 ( \41046 , \26342 , \31639 );
and \U$40703 ( \41047 , \26078 , \31636 );
nor \U$40704 ( \41048 , \41046 , \41047 );
xnor \U$40705 ( \41049 , \41048 , \30584 );
and \U$40706 ( \41050 , \26973 , \30826 );
and \U$40707 ( \41051 , \26601 , \30824 );
nor \U$40708 ( \41052 , \41050 , \41051 );
xnor \U$40709 ( \41053 , \41052 , \30587 );
and \U$40710 ( \41054 , \41049 , \41053 );
and \U$40711 ( \41055 , \41053 , \25817 );
and \U$40712 ( \41056 , \41049 , \25817 );
or \U$40713 ( \41057 , \41054 , \41055 , \41056 );
and \U$40714 ( \41058 , \27325 , \30258 );
and \U$40715 ( \41059 , \26982 , \30256 );
nor \U$40716 ( \41060 , \41058 , \41059 );
xnor \U$40717 ( \41061 , \41060 , \29948 );
and \U$40718 ( \41062 , \27830 , \29721 );
and \U$40719 ( \41063 , \27527 , \29719 );
nor \U$40720 ( \41064 , \41062 , \41063 );
xnor \U$40721 ( \41065 , \41064 , \29350 );
and \U$40722 ( \41066 , \41061 , \41065 );
and \U$40723 ( \41067 , \28528 , \29159 );
and \U$40724 ( \41068 , \28002 , \29157 );
nor \U$40725 ( \41069 , \41067 , \41068 );
xnor \U$40726 ( \41070 , \41069 , \28841 );
and \U$40727 ( \41071 , \41065 , \41070 );
and \U$40728 ( \41072 , \41061 , \41070 );
or \U$40729 ( \41073 , \41066 , \41071 , \41072 );
and \U$40730 ( \41074 , \41057 , \41073 );
and \U$40731 ( \41075 , \29198 , \28592 );
and \U$40732 ( \41076 , \28952 , \28590 );
nor \U$40733 ( \41077 , \41075 , \41076 );
xnor \U$40734 ( \41078 , \41077 , \28343 );
and \U$40735 ( \41079 , \29522 , \28063 );
and \U$40736 ( \41080 , \29203 , \28061 );
nor \U$40737 ( \41081 , \41079 , \41080 );
xnor \U$40738 ( \41082 , \41081 , \27803 );
and \U$40739 ( \41083 , \41078 , \41082 );
and \U$40740 ( \41084 , \30375 , \27569 );
and \U$40741 ( \41085 , \29806 , \27567 );
nor \U$40742 ( \41086 , \41084 , \41085 );
xnor \U$40743 ( \41087 , \41086 , \27254 );
and \U$40744 ( \41088 , \41082 , \41087 );
and \U$40745 ( \41089 , \41078 , \41087 );
or \U$40746 ( \41090 , \41083 , \41088 , \41089 );
and \U$40747 ( \41091 , \41073 , \41090 );
and \U$40748 ( \41092 , \41057 , \41090 );
or \U$40749 ( \41093 , \41074 , \41091 , \41092 );
and \U$40750 ( \41094 , \41045 , \41093 );
xor \U$40751 ( \41095 , \40926 , \40930 );
xor \U$40752 ( \41096 , \41095 , \40935 );
xor \U$40753 ( \41097 , \40942 , \40946 );
xor \U$40754 ( \41098 , \41097 , \40951 );
and \U$40755 ( \41099 , \41096 , \41098 );
xor \U$40756 ( \41100 , \40959 , \40963 );
xor \U$40757 ( \41101 , \41100 , \40968 );
and \U$40758 ( \41102 , \41098 , \41101 );
and \U$40759 ( \41103 , \41096 , \41101 );
or \U$40760 ( \41104 , \41099 , \41102 , \41103 );
and \U$40761 ( \41105 , \41093 , \41104 );
and \U$40762 ( \41106 , \41045 , \41104 );
or \U$40763 ( \41107 , \41094 , \41105 , \41106 );
xor \U$40764 ( \41108 , \40938 , \40954 );
xor \U$40765 ( \41109 , \41108 , \40971 );
xor \U$40766 ( \41110 , \40976 , \40978 );
xor \U$40767 ( \41111 , \41110 , \40981 );
and \U$40768 ( \41112 , \41109 , \41111 );
xor \U$40769 ( \41113 , \40987 , \40989 );
and \U$40770 ( \41114 , \41111 , \41113 );
and \U$40771 ( \41115 , \41109 , \41113 );
or \U$40772 ( \41116 , \41112 , \41114 , \41115 );
and \U$40773 ( \41117 , \41107 , \41116 );
xor \U$40774 ( \41118 , \40995 , \40997 );
xor \U$40775 ( \41119 , \41118 , \40999 );
and \U$40776 ( \41120 , \41116 , \41119 );
and \U$40777 ( \41121 , \41107 , \41119 );
or \U$40778 ( \41122 , \41117 , \41120 , \41121 );
xor \U$40779 ( \41123 , \40848 , \40872 );
xor \U$40780 ( \41124 , \41123 , \40878 );
and \U$40781 ( \41125 , \41122 , \41124 );
xor \U$40782 ( \41126 , \40993 , \41002 );
xor \U$40783 ( \41127 , \41126 , \41005 );
and \U$40784 ( \41128 , \41124 , \41127 );
and \U$40785 ( \41129 , \41122 , \41127 );
or \U$40786 ( \41130 , \41125 , \41128 , \41129 );
and \U$40787 ( \41131 , \41019 , \41130 );
xor \U$40788 ( \41132 , \41019 , \41130 );
xor \U$40789 ( \41133 , \41122 , \41124 );
xor \U$40790 ( \41134 , \41133 , \41127 );
and \U$40791 ( \41135 , \29806 , \28063 );
and \U$40792 ( \41136 , \29522 , \28061 );
nor \U$40793 ( \41137 , \41135 , \41136 );
xnor \U$40794 ( \41138 , \41137 , \27803 );
and \U$40795 ( \41139 , \30383 , \27569 );
and \U$40796 ( \41140 , \30375 , \27567 );
nor \U$40797 ( \41141 , \41139 , \41140 );
xnor \U$40798 ( \41142 , \41141 , \27254 );
and \U$40799 ( \41143 , \41138 , \41142 );
and \U$40800 ( \41144 , \30991 , \27060 );
and \U$40801 ( \41145 , \30986 , \27058 );
nor \U$40802 ( \41146 , \41144 , \41145 );
xnor \U$40803 ( \41147 , \41146 , \26720 );
and \U$40804 ( \41148 , \41142 , \41147 );
and \U$40805 ( \41149 , \41138 , \41147 );
or \U$40806 ( \41150 , \41143 , \41148 , \41149 );
and \U$40807 ( \41151 , \26601 , \31639 );
and \U$40808 ( \41152 , \26342 , \31636 );
nor \U$40809 ( \41153 , \41151 , \41152 );
xnor \U$40810 ( \41154 , \41153 , \30584 );
and \U$40811 ( \41155 , \26982 , \30826 );
and \U$40812 ( \41156 , \26973 , \30824 );
nor \U$40813 ( \41157 , \41155 , \41156 );
xnor \U$40814 ( \41158 , \41157 , \30587 );
and \U$40815 ( \41159 , \41154 , \41158 );
and \U$40816 ( \41160 , \27527 , \30258 );
and \U$40817 ( \41161 , \27325 , \30256 );
nor \U$40818 ( \41162 , \41160 , \41161 );
xnor \U$40819 ( \41163 , \41162 , \29948 );
and \U$40820 ( \41164 , \41158 , \41163 );
and \U$40821 ( \41165 , \41154 , \41163 );
or \U$40822 ( \41166 , \41159 , \41164 , \41165 );
and \U$40823 ( \41167 , \41150 , \41166 );
and \U$40824 ( \41168 , \28002 , \29721 );
and \U$40825 ( \41169 , \27830 , \29719 );
nor \U$40826 ( \41170 , \41168 , \41169 );
xnor \U$40827 ( \41171 , \41170 , \29350 );
and \U$40828 ( \41172 , \28952 , \29159 );
and \U$40829 ( \41173 , \28528 , \29157 );
nor \U$40830 ( \41174 , \41172 , \41173 );
xnor \U$40831 ( \41175 , \41174 , \28841 );
and \U$40832 ( \41176 , \41171 , \41175 );
and \U$40833 ( \41177 , \29203 , \28592 );
and \U$40834 ( \41178 , \29198 , \28590 );
nor \U$40835 ( \41179 , \41177 , \41178 );
xnor \U$40836 ( \41180 , \41179 , \28343 );
and \U$40837 ( \41181 , \41175 , \41180 );
and \U$40838 ( \41182 , \41171 , \41180 );
or \U$40839 ( \41183 , \41176 , \41181 , \41182 );
and \U$40840 ( \41184 , \41166 , \41183 );
and \U$40841 ( \41185 , \41150 , \41183 );
or \U$40842 ( \41186 , \41167 , \41184 , \41185 );
xor \U$40843 ( \41187 , \41061 , \41065 );
xor \U$40844 ( \41188 , \41187 , \41070 );
xor \U$40845 ( \41189 , \41023 , \41027 );
xor \U$40846 ( \41190 , \41189 , \41030 );
and \U$40847 ( \41191 , \41188 , \41190 );
xor \U$40848 ( \41192 , \41078 , \41082 );
xor \U$40849 ( \41193 , \41192 , \41087 );
and \U$40850 ( \41194 , \41190 , \41193 );
and \U$40851 ( \41195 , \41188 , \41193 );
or \U$40852 ( \41196 , \41191 , \41194 , \41195 );
and \U$40853 ( \41197 , \41186 , \41196 );
xor \U$40854 ( \41198 , \41096 , \41098 );
xor \U$40855 ( \41199 , \41198 , \41101 );
and \U$40856 ( \41200 , \41196 , \41199 );
and \U$40857 ( \41201 , \41186 , \41199 );
or \U$40858 ( \41202 , \41197 , \41200 , \41201 );
xor \U$40859 ( \41203 , \41045 , \41093 );
xor \U$40860 ( \41204 , \41203 , \41104 );
and \U$40861 ( \41205 , \41202 , \41204 );
xor \U$40862 ( \41206 , \41109 , \41111 );
xor \U$40863 ( \41207 , \41206 , \41113 );
and \U$40864 ( \41208 , \41204 , \41207 );
and \U$40865 ( \41209 , \41202 , \41207 );
or \U$40866 ( \41210 , \41205 , \41208 , \41209 );
xor \U$40867 ( \41211 , \40974 , \40984 );
xor \U$40868 ( \41212 , \41211 , \40990 );
and \U$40869 ( \41213 , \41210 , \41212 );
xor \U$40870 ( \41214 , \41107 , \41116 );
xor \U$40871 ( \41215 , \41214 , \41119 );
and \U$40872 ( \41216 , \41212 , \41215 );
and \U$40873 ( \41217 , \41210 , \41215 );
or \U$40874 ( \41218 , \41213 , \41216 , \41217 );
and \U$40875 ( \41219 , \41134 , \41218 );
xor \U$40876 ( \41220 , \41134 , \41218 );
xor \U$40877 ( \41221 , \41210 , \41212 );
xor \U$40878 ( \41222 , \41221 , \41215 );
and \U$40879 ( \41223 , \26973 , \31639 );
and \U$40880 ( \41224 , \26601 , \31636 );
nor \U$40881 ( \41225 , \41223 , \41224 );
xnor \U$40882 ( \41226 , \41225 , \30584 );
and \U$40883 ( \41227 , \27325 , \30826 );
and \U$40884 ( \41228 , \26982 , \30824 );
nor \U$40885 ( \41229 , \41227 , \41228 );
xnor \U$40886 ( \41230 , \41229 , \30587 );
and \U$40887 ( \41231 , \41226 , \41230 );
and \U$40888 ( \41232 , \41230 , \26230 );
and \U$40889 ( \41233 , \41226 , \26230 );
or \U$40890 ( \41234 , \41231 , \41232 , \41233 );
and \U$40891 ( \41235 , \29522 , \28592 );
and \U$40892 ( \41236 , \29203 , \28590 );
nor \U$40893 ( \41237 , \41235 , \41236 );
xnor \U$40894 ( \41238 , \41237 , \28343 );
and \U$40895 ( \41239 , \30375 , \28063 );
and \U$40896 ( \41240 , \29806 , \28061 );
nor \U$40897 ( \41241 , \41239 , \41240 );
xnor \U$40898 ( \41242 , \41241 , \27803 );
and \U$40899 ( \41243 , \41238 , \41242 );
and \U$40900 ( \41244 , \30986 , \27569 );
and \U$40901 ( \41245 , \30383 , \27567 );
nor \U$40902 ( \41246 , \41244 , \41245 );
xnor \U$40903 ( \41247 , \41246 , \27254 );
and \U$40904 ( \41248 , \41242 , \41247 );
and \U$40905 ( \41249 , \41238 , \41247 );
or \U$40906 ( \41250 , \41243 , \41248 , \41249 );
and \U$40907 ( \41251 , \41234 , \41250 );
and \U$40908 ( \41252 , \27830 , \30258 );
and \U$40909 ( \41253 , \27527 , \30256 );
nor \U$40910 ( \41254 , \41252 , \41253 );
xnor \U$40911 ( \41255 , \41254 , \29948 );
and \U$40912 ( \41256 , \28528 , \29721 );
and \U$40913 ( \41257 , \28002 , \29719 );
nor \U$40914 ( \41258 , \41256 , \41257 );
xnor \U$40915 ( \41259 , \41258 , \29350 );
and \U$40916 ( \41260 , \41255 , \41259 );
and \U$40917 ( \41261 , \29198 , \29159 );
and \U$40918 ( \41262 , \28952 , \29157 );
nor \U$40919 ( \41263 , \41261 , \41262 );
xnor \U$40920 ( \41264 , \41263 , \28841 );
and \U$40921 ( \41265 , \41259 , \41264 );
and \U$40922 ( \41266 , \41255 , \41264 );
or \U$40923 ( \41267 , \41260 , \41265 , \41266 );
and \U$40924 ( \41268 , \41250 , \41267 );
and \U$40925 ( \41269 , \41234 , \41267 );
or \U$40926 ( \41270 , \41251 , \41268 , \41269 );
and \U$40927 ( \41271 , \31792 , \26471 );
and \U$40928 ( \41272 , \31172 , \26469 );
nor \U$40929 ( \41273 , \41271 , \41272 );
xnor \U$40930 ( \41274 , \41273 , \26230 );
xor \U$40931 ( \41275 , \41138 , \41142 );
xor \U$40932 ( \41276 , \41275 , \41147 );
and \U$40933 ( \41277 , \41274 , \41276 );
xor \U$40934 ( \41278 , \41171 , \41175 );
xor \U$40935 ( \41279 , \41278 , \41180 );
and \U$40936 ( \41280 , \41276 , \41279 );
and \U$40937 ( \41281 , \41274 , \41279 );
or \U$40938 ( \41282 , \41277 , \41280 , \41281 );
and \U$40939 ( \41283 , \41270 , \41282 );
xor \U$40940 ( \41284 , \41049 , \41053 );
xor \U$40941 ( \41285 , \41284 , \25817 );
and \U$40942 ( \41286 , \41282 , \41285 );
and \U$40943 ( \41287 , \41270 , \41285 );
or \U$40944 ( \41288 , \41283 , \41286 , \41287 );
xor \U$40945 ( \41289 , \41150 , \41166 );
xor \U$40946 ( \41290 , \41289 , \41183 );
xor \U$40947 ( \41291 , \41188 , \41190 );
xor \U$40948 ( \41292 , \41291 , \41193 );
and \U$40949 ( \41293 , \41290 , \41292 );
and \U$40950 ( \41294 , \41288 , \41293 );
xor \U$40951 ( \41295 , \41033 , \41037 );
xor \U$40952 ( \41296 , \41295 , \41042 );
and \U$40953 ( \41297 , \41293 , \41296 );
and \U$40954 ( \41298 , \41288 , \41296 );
or \U$40955 ( \41299 , \41294 , \41297 , \41298 );
xor \U$40956 ( \41300 , \41057 , \41073 );
xor \U$40957 ( \41301 , \41300 , \41090 );
xor \U$40958 ( \41302 , \41186 , \41196 );
xor \U$40959 ( \41303 , \41302 , \41199 );
and \U$40960 ( \41304 , \41301 , \41303 );
and \U$40961 ( \41305 , \41299 , \41304 );
xor \U$40962 ( \41306 , \41202 , \41204 );
xor \U$40963 ( \41307 , \41306 , \41207 );
and \U$40964 ( \41308 , \41304 , \41307 );
and \U$40965 ( \41309 , \41299 , \41307 );
or \U$40966 ( \41310 , \41305 , \41308 , \41309 );
and \U$40967 ( \41311 , \41222 , \41310 );
xor \U$40968 ( \41312 , \41222 , \41310 );
xor \U$40969 ( \41313 , \41299 , \41304 );
xor \U$40970 ( \41314 , \41313 , \41307 );
and \U$40971 ( \41315 , \28952 , \29721 );
and \U$40972 ( \41316 , \28528 , \29719 );
nor \U$40973 ( \41317 , \41315 , \41316 );
xnor \U$40974 ( \41318 , \41317 , \29350 );
and \U$40975 ( \41319 , \29203 , \29159 );
and \U$40976 ( \41320 , \29198 , \29157 );
nor \U$40977 ( \41321 , \41319 , \41320 );
xnor \U$40978 ( \41322 , \41321 , \28841 );
and \U$40979 ( \41323 , \41318 , \41322 );
and \U$40980 ( \41324 , \29806 , \28592 );
and \U$40981 ( \41325 , \29522 , \28590 );
nor \U$40982 ( \41326 , \41324 , \41325 );
xnor \U$40983 ( \41327 , \41326 , \28343 );
and \U$40984 ( \41328 , \41322 , \41327 );
and \U$40985 ( \41329 , \41318 , \41327 );
or \U$40986 ( \41330 , \41323 , \41328 , \41329 );
and \U$40987 ( \41331 , \26982 , \31639 );
and \U$40988 ( \41332 , \26973 , \31636 );
nor \U$40989 ( \41333 , \41331 , \41332 );
xnor \U$40990 ( \41334 , \41333 , \30584 );
and \U$40991 ( \41335 , \27527 , \30826 );
and \U$40992 ( \41336 , \27325 , \30824 );
nor \U$40993 ( \41337 , \41335 , \41336 );
xnor \U$40994 ( \41338 , \41337 , \30587 );
and \U$40995 ( \41339 , \41334 , \41338 );
and \U$40996 ( \41340 , \28002 , \30258 );
and \U$40997 ( \41341 , \27830 , \30256 );
nor \U$40998 ( \41342 , \41340 , \41341 );
xnor \U$40999 ( \41343 , \41342 , \29948 );
and \U$41000 ( \41344 , \41338 , \41343 );
and \U$41001 ( \41345 , \41334 , \41343 );
or \U$41002 ( \41346 , \41339 , \41344 , \41345 );
and \U$41003 ( \41347 , \41330 , \41346 );
and \U$41004 ( \41348 , \30383 , \28063 );
and \U$41005 ( \41349 , \30375 , \28061 );
nor \U$41006 ( \41350 , \41348 , \41349 );
xnor \U$41007 ( \41351 , \41350 , \27803 );
and \U$41008 ( \41352 , \30991 , \27569 );
and \U$41009 ( \41353 , \30986 , \27567 );
nor \U$41010 ( \41354 , \41352 , \41353 );
xnor \U$41011 ( \41355 , \41354 , \27254 );
and \U$41012 ( \41356 , \41351 , \41355 );
and \U$41013 ( \41357 , \31792 , \27060 );
and \U$41014 ( \41358 , \31172 , \27058 );
nor \U$41015 ( \41359 , \41357 , \41358 );
xnor \U$41016 ( \41360 , \41359 , \26720 );
and \U$41017 ( \41361 , \41355 , \41360 );
and \U$41018 ( \41362 , \41351 , \41360 );
or \U$41019 ( \41363 , \41356 , \41361 , \41362 );
and \U$41020 ( \41364 , \41346 , \41363 );
and \U$41021 ( \41365 , \41330 , \41363 );
or \U$41022 ( \41366 , \41347 , \41364 , \41365 );
and \U$41023 ( \41367 , \31172 , \27060 );
and \U$41024 ( \41368 , \30991 , \27058 );
nor \U$41025 ( \41369 , \41367 , \41368 );
xnor \U$41026 ( \41370 , \41369 , \26720 );
nand \U$41027 ( \41371 , \31792 , \26469 );
xnor \U$41028 ( \41372 , \41371 , \26230 );
and \U$41029 ( \41373 , \41370 , \41372 );
xor \U$41030 ( \41374 , \41238 , \41242 );
xor \U$41031 ( \41375 , \41374 , \41247 );
and \U$41032 ( \41376 , \41372 , \41375 );
and \U$41033 ( \41377 , \41370 , \41375 );
or \U$41034 ( \41378 , \41373 , \41376 , \41377 );
and \U$41035 ( \41379 , \41366 , \41378 );
xor \U$41036 ( \41380 , \41154 , \41158 );
xor \U$41037 ( \41381 , \41380 , \41163 );
and \U$41038 ( \41382 , \41378 , \41381 );
and \U$41039 ( \41383 , \41366 , \41381 );
or \U$41040 ( \41384 , \41379 , \41382 , \41383 );
xor \U$41041 ( \41385 , \41270 , \41282 );
xor \U$41042 ( \41386 , \41385 , \41285 );
and \U$41043 ( \41387 , \41384 , \41386 );
xor \U$41044 ( \41388 , \41290 , \41292 );
and \U$41045 ( \41389 , \41386 , \41388 );
and \U$41046 ( \41390 , \41384 , \41388 );
or \U$41047 ( \41391 , \41387 , \41389 , \41390 );
xor \U$41048 ( \41392 , \41288 , \41293 );
xor \U$41049 ( \41393 , \41392 , \41296 );
and \U$41050 ( \41394 , \41391 , \41393 );
xor \U$41051 ( \41395 , \41301 , \41303 );
and \U$41052 ( \41396 , \41393 , \41395 );
and \U$41053 ( \41397 , \41391 , \41395 );
or \U$41054 ( \41398 , \41394 , \41396 , \41397 );
and \U$41055 ( \41399 , \41314 , \41398 );
xor \U$41056 ( \41400 , \41314 , \41398 );
xor \U$41057 ( \41401 , \41391 , \41393 );
xor \U$41058 ( \41402 , \41401 , \41395 );
and \U$41059 ( \41403 , \28528 , \30258 );
and \U$41060 ( \41404 , \28002 , \30256 );
nor \U$41061 ( \41405 , \41403 , \41404 );
xnor \U$41062 ( \41406 , \41405 , \29948 );
and \U$41063 ( \41407 , \29198 , \29721 );
and \U$41064 ( \41408 , \28952 , \29719 );
nor \U$41065 ( \41409 , \41407 , \41408 );
xnor \U$41066 ( \41410 , \41409 , \29350 );
and \U$41067 ( \41411 , \41406 , \41410 );
and \U$41068 ( \41412 , \29522 , \29159 );
and \U$41069 ( \41413 , \29203 , \29157 );
nor \U$41070 ( \41414 , \41412 , \41413 );
xnor \U$41071 ( \41415 , \41414 , \28841 );
and \U$41072 ( \41416 , \41410 , \41415 );
and \U$41073 ( \41417 , \41406 , \41415 );
or \U$41074 ( \41418 , \41411 , \41416 , \41417 );
and \U$41075 ( \41419 , \27325 , \31639 );
and \U$41076 ( \41420 , \26982 , \31636 );
nor \U$41077 ( \41421 , \41419 , \41420 );
xnor \U$41078 ( \41422 , \41421 , \30584 );
and \U$41079 ( \41423 , \27830 , \30826 );
and \U$41080 ( \41424 , \27527 , \30824 );
nor \U$41081 ( \41425 , \41423 , \41424 );
xnor \U$41082 ( \41426 , \41425 , \30587 );
and \U$41083 ( \41427 , \41422 , \41426 );
and \U$41084 ( \41428 , \41426 , \26720 );
and \U$41085 ( \41429 , \41422 , \26720 );
or \U$41086 ( \41430 , \41427 , \41428 , \41429 );
and \U$41087 ( \41431 , \41418 , \41430 );
and \U$41088 ( \41432 , \30375 , \28592 );
and \U$41089 ( \41433 , \29806 , \28590 );
nor \U$41090 ( \41434 , \41432 , \41433 );
xnor \U$41091 ( \41435 , \41434 , \28343 );
and \U$41092 ( \41436 , \30986 , \28063 );
and \U$41093 ( \41437 , \30383 , \28061 );
nor \U$41094 ( \41438 , \41436 , \41437 );
xnor \U$41095 ( \41439 , \41438 , \27803 );
and \U$41096 ( \41440 , \41435 , \41439 );
and \U$41097 ( \41441 , \31172 , \27569 );
and \U$41098 ( \41442 , \30991 , \27567 );
nor \U$41099 ( \41443 , \41441 , \41442 );
xnor \U$41100 ( \41444 , \41443 , \27254 );
and \U$41101 ( \41445 , \41439 , \41444 );
and \U$41102 ( \41446 , \41435 , \41444 );
or \U$41103 ( \41447 , \41440 , \41445 , \41446 );
and \U$41104 ( \41448 , \41430 , \41447 );
and \U$41105 ( \41449 , \41418 , \41447 );
or \U$41106 ( \41450 , \41431 , \41448 , \41449 );
xor \U$41107 ( \41451 , \41318 , \41322 );
xor \U$41108 ( \41452 , \41451 , \41327 );
xor \U$41109 ( \41453 , \41334 , \41338 );
xor \U$41110 ( \41454 , \41453 , \41343 );
and \U$41111 ( \41455 , \41452 , \41454 );
xor \U$41112 ( \41456 , \41351 , \41355 );
xor \U$41113 ( \41457 , \41456 , \41360 );
and \U$41114 ( \41458 , \41454 , \41457 );
and \U$41115 ( \41459 , \41452 , \41457 );
or \U$41116 ( \41460 , \41455 , \41458 , \41459 );
and \U$41117 ( \41461 , \41450 , \41460 );
xor \U$41118 ( \41462 , \41255 , \41259 );
xor \U$41119 ( \41463 , \41462 , \41264 );
and \U$41120 ( \41464 , \41460 , \41463 );
and \U$41121 ( \41465 , \41450 , \41463 );
or \U$41122 ( \41466 , \41461 , \41464 , \41465 );
xor \U$41123 ( \41467 , \41226 , \41230 );
xor \U$41124 ( \41468 , \41467 , \26230 );
xor \U$41125 ( \41469 , \41330 , \41346 );
xor \U$41126 ( \41470 , \41469 , \41363 );
and \U$41127 ( \41471 , \41468 , \41470 );
xor \U$41128 ( \41472 , \41370 , \41372 );
xor \U$41129 ( \41473 , \41472 , \41375 );
and \U$41130 ( \41474 , \41470 , \41473 );
and \U$41131 ( \41475 , \41468 , \41473 );
or \U$41132 ( \41476 , \41471 , \41474 , \41475 );
and \U$41133 ( \41477 , \41466 , \41476 );
xor \U$41134 ( \41478 , \41274 , \41276 );
xor \U$41135 ( \41479 , \41478 , \41279 );
and \U$41136 ( \41480 , \41476 , \41479 );
and \U$41137 ( \41481 , \41466 , \41479 );
or \U$41138 ( \41482 , \41477 , \41480 , \41481 );
xor \U$41139 ( \41483 , \41234 , \41250 );
xor \U$41140 ( \41484 , \41483 , \41267 );
xor \U$41141 ( \41485 , \41366 , \41378 );
xor \U$41142 ( \41486 , \41485 , \41381 );
and \U$41143 ( \41487 , \41484 , \41486 );
and \U$41144 ( \41488 , \41482 , \41487 );
xor \U$41145 ( \41489 , \41384 , \41386 );
xor \U$41146 ( \41490 , \41489 , \41388 );
and \U$41147 ( \41491 , \41487 , \41490 );
and \U$41148 ( \41492 , \41482 , \41490 );
or \U$41149 ( \41493 , \41488 , \41491 , \41492 );
and \U$41150 ( \41494 , \41402 , \41493 );
xor \U$41151 ( \41495 , \41402 , \41493 );
xor \U$41152 ( \41496 , \41482 , \41487 );
xor \U$41153 ( \41497 , \41496 , \41490 );
and \U$41154 ( \41498 , \27527 , \31639 );
and \U$41155 ( \41499 , \27325 , \31636 );
nor \U$41156 ( \41500 , \41498 , \41499 );
xnor \U$41157 ( \41501 , \41500 , \30584 );
and \U$41158 ( \41502 , \28002 , \30826 );
and \U$41159 ( \41503 , \27830 , \30824 );
nor \U$41160 ( \41504 , \41502 , \41503 );
xnor \U$41161 ( \41505 , \41504 , \30587 );
and \U$41162 ( \41506 , \41501 , \41505 );
and \U$41163 ( \41507 , \28952 , \30258 );
and \U$41164 ( \41508 , \28528 , \30256 );
nor \U$41165 ( \41509 , \41507 , \41508 );
xnor \U$41166 ( \41510 , \41509 , \29948 );
and \U$41167 ( \41511 , \41505 , \41510 );
and \U$41168 ( \41512 , \41501 , \41510 );
or \U$41169 ( \41513 , \41506 , \41511 , \41512 );
and \U$41170 ( \41514 , \29203 , \29721 );
and \U$41171 ( \41515 , \29198 , \29719 );
nor \U$41172 ( \41516 , \41514 , \41515 );
xnor \U$41173 ( \41517 , \41516 , \29350 );
and \U$41174 ( \41518 , \29806 , \29159 );
and \U$41175 ( \41519 , \29522 , \29157 );
nor \U$41176 ( \41520 , \41518 , \41519 );
xnor \U$41177 ( \41521 , \41520 , \28841 );
and \U$41178 ( \41522 , \41517 , \41521 );
and \U$41179 ( \41523 , \30383 , \28592 );
and \U$41180 ( \41524 , \30375 , \28590 );
nor \U$41181 ( \41525 , \41523 , \41524 );
xnor \U$41182 ( \41526 , \41525 , \28343 );
and \U$41183 ( \41527 , \41521 , \41526 );
and \U$41184 ( \41528 , \41517 , \41526 );
or \U$41185 ( \41529 , \41522 , \41527 , \41528 );
and \U$41186 ( \41530 , \41513 , \41529 );
and \U$41187 ( \41531 , \30991 , \28063 );
and \U$41188 ( \41532 , \30986 , \28061 );
nor \U$41189 ( \41533 , \41531 , \41532 );
xnor \U$41190 ( \41534 , \41533 , \27803 );
and \U$41191 ( \41535 , \31792 , \27569 );
and \U$41192 ( \41536 , \31172 , \27567 );
nor \U$41193 ( \41537 , \41535 , \41536 );
xnor \U$41194 ( \41538 , \41537 , \27254 );
and \U$41195 ( \41539 , \41534 , \41538 );
and \U$41196 ( \41540 , \41529 , \41539 );
and \U$41197 ( \41541 , \41513 , \41539 );
or \U$41198 ( \41542 , \41530 , \41540 , \41541 );
nand \U$41199 ( \41543 , \31792 , \27058 );
xnor \U$41200 ( \41544 , \41543 , \26720 );
xor \U$41201 ( \41545 , \41406 , \41410 );
xor \U$41202 ( \41546 , \41545 , \41415 );
and \U$41203 ( \41547 , \41544 , \41546 );
xor \U$41204 ( \41548 , \41435 , \41439 );
xor \U$41205 ( \41549 , \41548 , \41444 );
and \U$41206 ( \41550 , \41546 , \41549 );
and \U$41207 ( \41551 , \41544 , \41549 );
or \U$41208 ( \41552 , \41547 , \41550 , \41551 );
and \U$41209 ( \41553 , \41542 , \41552 );
xor \U$41210 ( \41554 , \41452 , \41454 );
xor \U$41211 ( \41555 , \41554 , \41457 );
and \U$41212 ( \41556 , \41552 , \41555 );
and \U$41213 ( \41557 , \41542 , \41555 );
or \U$41214 ( \41558 , \41553 , \41556 , \41557 );
xor \U$41215 ( \41559 , \41450 , \41460 );
xor \U$41216 ( \41560 , \41559 , \41463 );
and \U$41217 ( \41561 , \41558 , \41560 );
xor \U$41218 ( \41562 , \41468 , \41470 );
xor \U$41219 ( \41563 , \41562 , \41473 );
and \U$41220 ( \41564 , \41560 , \41563 );
and \U$41221 ( \41565 , \41558 , \41563 );
or \U$41222 ( \41566 , \41561 , \41564 , \41565 );
xor \U$41223 ( \41567 , \41466 , \41476 );
xor \U$41224 ( \41568 , \41567 , \41479 );
and \U$41225 ( \41569 , \41566 , \41568 );
xor \U$41226 ( \41570 , \41484 , \41486 );
and \U$41227 ( \41571 , \41568 , \41570 );
and \U$41228 ( \41572 , \41566 , \41570 );
or \U$41229 ( \41573 , \41569 , \41571 , \41572 );
and \U$41230 ( \41574 , \41497 , \41573 );
xor \U$41231 ( \41575 , \41497 , \41573 );
xor \U$41232 ( \41576 , \41566 , \41568 );
xor \U$41233 ( \41577 , \41576 , \41570 );
and \U$41234 ( \41578 , \30986 , \28592 );
and \U$41235 ( \41579 , \30383 , \28590 );
nor \U$41236 ( \41580 , \41578 , \41579 );
xnor \U$41237 ( \41581 , \41580 , \28343 );
and \U$41238 ( \41582 , \31172 , \28063 );
and \U$41239 ( \41583 , \30991 , \28061 );
nor \U$41240 ( \41584 , \41582 , \41583 );
xnor \U$41241 ( \41585 , \41584 , \27803 );
and \U$41242 ( \41586 , \41581 , \41585 );
nand \U$41243 ( \41587 , \31792 , \27567 );
xnor \U$41244 ( \41588 , \41587 , \27254 );
and \U$41245 ( \41589 , \41585 , \41588 );
and \U$41246 ( \41590 , \41581 , \41588 );
or \U$41247 ( \41591 , \41586 , \41589 , \41590 );
and \U$41248 ( \41592 , \27830 , \31639 );
and \U$41249 ( \41593 , \27527 , \31636 );
nor \U$41250 ( \41594 , \41592 , \41593 );
xnor \U$41251 ( \41595 , \41594 , \30584 );
and \U$41252 ( \41596 , \28528 , \30826 );
and \U$41253 ( \41597 , \28002 , \30824 );
nor \U$41254 ( \41598 , \41596 , \41597 );
xnor \U$41255 ( \41599 , \41598 , \30587 );
and \U$41256 ( \41600 , \41595 , \41599 );
and \U$41257 ( \41601 , \41599 , \27254 );
and \U$41258 ( \41602 , \41595 , \27254 );
or \U$41259 ( \41603 , \41600 , \41601 , \41602 );
and \U$41260 ( \41604 , \41591 , \41603 );
and \U$41261 ( \41605 , \29198 , \30258 );
and \U$41262 ( \41606 , \28952 , \30256 );
nor \U$41263 ( \41607 , \41605 , \41606 );
xnor \U$41264 ( \41608 , \41607 , \29948 );
and \U$41265 ( \41609 , \29522 , \29721 );
and \U$41266 ( \41610 , \29203 , \29719 );
nor \U$41267 ( \41611 , \41609 , \41610 );
xnor \U$41268 ( \41612 , \41611 , \29350 );
and \U$41269 ( \41613 , \41608 , \41612 );
and \U$41270 ( \41614 , \30375 , \29159 );
and \U$41271 ( \41615 , \29806 , \29157 );
nor \U$41272 ( \41616 , \41614 , \41615 );
xnor \U$41273 ( \41617 , \41616 , \28841 );
and \U$41274 ( \41618 , \41612 , \41617 );
and \U$41275 ( \41619 , \41608 , \41617 );
or \U$41276 ( \41620 , \41613 , \41618 , \41619 );
and \U$41277 ( \41621 , \41603 , \41620 );
and \U$41278 ( \41622 , \41591 , \41620 );
or \U$41279 ( \41623 , \41604 , \41621 , \41622 );
xor \U$41280 ( \41624 , \41501 , \41505 );
xor \U$41281 ( \41625 , \41624 , \41510 );
xor \U$41282 ( \41626 , \41517 , \41521 );
xor \U$41283 ( \41627 , \41626 , \41526 );
and \U$41284 ( \41628 , \41625 , \41627 );
xor \U$41285 ( \41629 , \41534 , \41538 );
and \U$41286 ( \41630 , \41627 , \41629 );
and \U$41287 ( \41631 , \41625 , \41629 );
or \U$41288 ( \41632 , \41628 , \41630 , \41631 );
and \U$41289 ( \41633 , \41623 , \41632 );
xor \U$41290 ( \41634 , \41422 , \41426 );
xor \U$41291 ( \41635 , \41634 , \26720 );
and \U$41292 ( \41636 , \41632 , \41635 );
and \U$41293 ( \41637 , \41623 , \41635 );
or \U$41294 ( \41638 , \41633 , \41636 , \41637 );
xor \U$41295 ( \41639 , \41513 , \41529 );
xor \U$41296 ( \41640 , \41639 , \41539 );
xor \U$41297 ( \41641 , \41544 , \41546 );
xor \U$41298 ( \41642 , \41641 , \41549 );
and \U$41299 ( \41643 , \41640 , \41642 );
and \U$41300 ( \41644 , \41638 , \41643 );
xor \U$41301 ( \41645 , \41418 , \41430 );
xor \U$41302 ( \41646 , \41645 , \41447 );
and \U$41303 ( \41647 , \41643 , \41646 );
and \U$41304 ( \41648 , \41638 , \41646 );
or \U$41305 ( \41649 , \41644 , \41647 , \41648 );
xor \U$41306 ( \41650 , \41558 , \41560 );
xor \U$41307 ( \41651 , \41650 , \41563 );
and \U$41308 ( \41652 , \41649 , \41651 );
and \U$41309 ( \41653 , \41577 , \41652 );
xor \U$41310 ( \41654 , \41577 , \41652 );
xor \U$41311 ( \41655 , \41649 , \41651 );
xor \U$41312 ( \41656 , \41638 , \41643 );
xor \U$41313 ( \41657 , \41656 , \41646 );
xor \U$41314 ( \41658 , \41542 , \41552 );
xor \U$41315 ( \41659 , \41658 , \41555 );
and \U$41316 ( \41660 , \41657 , \41659 );
and \U$41317 ( \41661 , \41655 , \41660 );
xor \U$41318 ( \41662 , \41655 , \41660 );
xor \U$41319 ( \41663 , \41657 , \41659 );
and \U$41320 ( \41664 , \28002 , \31639 );
and \U$41321 ( \41665 , \27830 , \31636 );
nor \U$41322 ( \41666 , \41664 , \41665 );
xnor \U$41323 ( \41667 , \41666 , \30584 );
and \U$41324 ( \41668 , \28952 , \30826 );
and \U$41325 ( \41669 , \28528 , \30824 );
nor \U$41326 ( \41670 , \41668 , \41669 );
xnor \U$41327 ( \41671 , \41670 , \30587 );
and \U$41328 ( \41672 , \41667 , \41671 );
and \U$41329 ( \41673 , \29203 , \30258 );
and \U$41330 ( \41674 , \29198 , \30256 );
nor \U$41331 ( \41675 , \41673 , \41674 );
xnor \U$41332 ( \41676 , \41675 , \29948 );
and \U$41333 ( \41677 , \41671 , \41676 );
and \U$41334 ( \41678 , \41667 , \41676 );
or \U$41335 ( \41679 , \41672 , \41677 , \41678 );
and \U$41336 ( \41680 , \29806 , \29721 );
and \U$41337 ( \41681 , \29522 , \29719 );
nor \U$41338 ( \41682 , \41680 , \41681 );
xnor \U$41339 ( \41683 , \41682 , \29350 );
and \U$41340 ( \41684 , \30383 , \29159 );
and \U$41341 ( \41685 , \30375 , \29157 );
nor \U$41342 ( \41686 , \41684 , \41685 );
xnor \U$41343 ( \41687 , \41686 , \28841 );
and \U$41344 ( \41688 , \41683 , \41687 );
and \U$41345 ( \41689 , \30991 , \28592 );
and \U$41346 ( \41690 , \30986 , \28590 );
nor \U$41347 ( \41691 , \41689 , \41690 );
xnor \U$41348 ( \41692 , \41691 , \28343 );
and \U$41349 ( \41693 , \41687 , \41692 );
and \U$41350 ( \41694 , \41683 , \41692 );
or \U$41351 ( \41695 , \41688 , \41693 , \41694 );
and \U$41352 ( \41696 , \41679 , \41695 );
xor \U$41353 ( \41697 , \41581 , \41585 );
xor \U$41354 ( \41698 , \41697 , \41588 );
and \U$41355 ( \41699 , \41695 , \41698 );
and \U$41356 ( \41700 , \41679 , \41698 );
or \U$41357 ( \41701 , \41696 , \41699 , \41700 );
xor \U$41358 ( \41702 , \41595 , \41599 );
xor \U$41359 ( \41703 , \41702 , \27254 );
xor \U$41360 ( \41704 , \41608 , \41612 );
xor \U$41361 ( \41705 , \41704 , \41617 );
and \U$41362 ( \41706 , \41703 , \41705 );
and \U$41363 ( \41707 , \41701 , \41706 );
xor \U$41364 ( \41708 , \41625 , \41627 );
xor \U$41365 ( \41709 , \41708 , \41629 );
and \U$41366 ( \41710 , \41706 , \41709 );
and \U$41367 ( \41711 , \41701 , \41709 );
or \U$41368 ( \41712 , \41707 , \41710 , \41711 );
xor \U$41369 ( \41713 , \41623 , \41632 );
xor \U$41370 ( \41714 , \41713 , \41635 );
and \U$41371 ( \41715 , \41712 , \41714 );
xor \U$41372 ( \41716 , \41640 , \41642 );
and \U$41373 ( \41717 , \41714 , \41716 );
and \U$41374 ( \41718 , \41712 , \41716 );
or \U$41375 ( \41719 , \41715 , \41717 , \41718 );
and \U$41376 ( \41720 , \41663 , \41719 );
xor \U$41377 ( \41721 , \41663 , \41719 );
xor \U$41378 ( \41722 , \41712 , \41714 );
xor \U$41379 ( \41723 , \41722 , \41716 );
and \U$41380 ( \41724 , \28528 , \31639 );
and \U$41381 ( \41725 , \28002 , \31636 );
nor \U$41382 ( \41726 , \41724 , \41725 );
xnor \U$41383 ( \41727 , \41726 , \30584 );
and \U$41384 ( \41728 , \29198 , \30826 );
and \U$41385 ( \41729 , \28952 , \30824 );
nor \U$41386 ( \41730 , \41728 , \41729 );
xnor \U$41387 ( \41731 , \41730 , \30587 );
and \U$41388 ( \41732 , \41727 , \41731 );
and \U$41389 ( \41733 , \41731 , \27803 );
and \U$41390 ( \41734 , \41727 , \27803 );
or \U$41391 ( \41735 , \41732 , \41733 , \41734 );
and \U$41392 ( \41736 , \29522 , \30258 );
and \U$41393 ( \41737 , \29203 , \30256 );
nor \U$41394 ( \41738 , \41736 , \41737 );
xnor \U$41395 ( \41739 , \41738 , \29948 );
and \U$41396 ( \41740 , \30375 , \29721 );
and \U$41397 ( \41741 , \29806 , \29719 );
nor \U$41398 ( \41742 , \41740 , \41741 );
xnor \U$41399 ( \41743 , \41742 , \29350 );
and \U$41400 ( \41744 , \41739 , \41743 );
and \U$41401 ( \41745 , \30986 , \29159 );
and \U$41402 ( \41746 , \30383 , \29157 );
nor \U$41403 ( \41747 , \41745 , \41746 );
xnor \U$41404 ( \41748 , \41747 , \28841 );
and \U$41405 ( \41749 , \41743 , \41748 );
and \U$41406 ( \41750 , \41739 , \41748 );
or \U$41407 ( \41751 , \41744 , \41749 , \41750 );
and \U$41408 ( \41752 , \41735 , \41751 );
and \U$41409 ( \41753 , \31792 , \28063 );
and \U$41410 ( \41754 , \31172 , \28061 );
nor \U$41411 ( \41755 , \41753 , \41754 );
xnor \U$41412 ( \41756 , \41755 , \27803 );
and \U$41413 ( \41757 , \41751 , \41756 );
and \U$41414 ( \41758 , \41735 , \41756 );
or \U$41415 ( \41759 , \41752 , \41757 , \41758 );
xor \U$41416 ( \41760 , \41679 , \41695 );
xor \U$41417 ( \41761 , \41760 , \41698 );
and \U$41418 ( \41762 , \41759 , \41761 );
xor \U$41419 ( \41763 , \41703 , \41705 );
and \U$41420 ( \41764 , \41761 , \41763 );
and \U$41421 ( \41765 , \41759 , \41763 );
or \U$41422 ( \41766 , \41762 , \41764 , \41765 );
xor \U$41423 ( \41767 , \41591 , \41603 );
xor \U$41424 ( \41768 , \41767 , \41620 );
and \U$41425 ( \41769 , \41766 , \41768 );
xor \U$41426 ( \41770 , \41701 , \41706 );
xor \U$41427 ( \41771 , \41770 , \41709 );
and \U$41428 ( \41772 , \41768 , \41771 );
and \U$41429 ( \41773 , \41766 , \41771 );
or \U$41430 ( \41774 , \41769 , \41772 , \41773 );
and \U$41431 ( \41775 , \41723 , \41774 );
xor \U$41432 ( \41776 , \41723 , \41774 );
xor \U$41433 ( \41777 , \41766 , \41768 );
xor \U$41434 ( \41778 , \41777 , \41771 );
and \U$41435 ( \41779 , \30383 , \29721 );
and \U$41436 ( \41780 , \30375 , \29719 );
nor \U$41437 ( \41781 , \41779 , \41780 );
xnor \U$41438 ( \41782 , \41781 , \29350 );
and \U$41439 ( \41783 , \30991 , \29159 );
and \U$41440 ( \41784 , \30986 , \29157 );
nor \U$41441 ( \41785 , \41783 , \41784 );
xnor \U$41442 ( \41786 , \41785 , \28841 );
and \U$41443 ( \41787 , \41782 , \41786 );
and \U$41444 ( \41788 , \31792 , \28592 );
and \U$41445 ( \41789 , \31172 , \28590 );
nor \U$41446 ( \41790 , \41788 , \41789 );
xnor \U$41447 ( \41791 , \41790 , \28343 );
and \U$41448 ( \41792 , \41786 , \41791 );
and \U$41449 ( \41793 , \41782 , \41791 );
or \U$41450 ( \41794 , \41787 , \41792 , \41793 );
and \U$41451 ( \41795 , \28952 , \31639 );
and \U$41452 ( \41796 , \28528 , \31636 );
nor \U$41453 ( \41797 , \41795 , \41796 );
xnor \U$41454 ( \41798 , \41797 , \30584 );
and \U$41455 ( \41799 , \29203 , \30826 );
and \U$41456 ( \41800 , \29198 , \30824 );
nor \U$41457 ( \41801 , \41799 , \41800 );
xnor \U$41458 ( \41802 , \41801 , \30587 );
and \U$41459 ( \41803 , \41798 , \41802 );
and \U$41460 ( \41804 , \29806 , \30258 );
and \U$41461 ( \41805 , \29522 , \30256 );
nor \U$41462 ( \41806 , \41804 , \41805 );
xnor \U$41463 ( \41807 , \41806 , \29948 );
and \U$41464 ( \41808 , \41802 , \41807 );
and \U$41465 ( \41809 , \41798 , \41807 );
or \U$41466 ( \41810 , \41803 , \41808 , \41809 );
and \U$41467 ( \41811 , \41794 , \41810 );
and \U$41468 ( \41812 , \31172 , \28592 );
and \U$41469 ( \41813 , \30991 , \28590 );
nor \U$41470 ( \41814 , \41812 , \41813 );
xnor \U$41471 ( \41815 , \41814 , \28343 );
and \U$41472 ( \41816 , \41810 , \41815 );
and \U$41473 ( \41817 , \41794 , \41815 );
or \U$41474 ( \41818 , \41811 , \41816 , \41817 );
nand \U$41475 ( \41819 , \31792 , \28061 );
xnor \U$41476 ( \41820 , \41819 , \27803 );
xor \U$41477 ( \41821 , \41727 , \41731 );
xor \U$41478 ( \41822 , \41821 , \27803 );
and \U$41479 ( \41823 , \41820 , \41822 );
xor \U$41480 ( \41824 , \41739 , \41743 );
xor \U$41481 ( \41825 , \41824 , \41748 );
and \U$41482 ( \41826 , \41822 , \41825 );
and \U$41483 ( \41827 , \41820 , \41825 );
or \U$41484 ( \41828 , \41823 , \41826 , \41827 );
and \U$41485 ( \41829 , \41818 , \41828 );
xor \U$41486 ( \41830 , \41683 , \41687 );
xor \U$41487 ( \41831 , \41830 , \41692 );
and \U$41488 ( \41832 , \41828 , \41831 );
and \U$41489 ( \41833 , \41818 , \41831 );
or \U$41490 ( \41834 , \41829 , \41832 , \41833 );
xor \U$41491 ( \41835 , \41667 , \41671 );
xor \U$41492 ( \41836 , \41835 , \41676 );
xor \U$41493 ( \41837 , \41735 , \41751 );
xor \U$41494 ( \41838 , \41837 , \41756 );
and \U$41495 ( \41839 , \41836 , \41838 );
and \U$41496 ( \41840 , \41834 , \41839 );
xor \U$41497 ( \41841 , \41759 , \41761 );
xor \U$41498 ( \41842 , \41841 , \41763 );
and \U$41499 ( \41843 , \41839 , \41842 );
and \U$41500 ( \41844 , \41834 , \41842 );
or \U$41501 ( \41845 , \41840 , \41843 , \41844 );
and \U$41502 ( \41846 , \41778 , \41845 );
xor \U$41503 ( \41847 , \41778 , \41845 );
xor \U$41504 ( \41848 , \41834 , \41839 );
xor \U$41505 ( \41849 , \41848 , \41842 );
and \U$41506 ( \41850 , \30375 , \30258 );
and \U$41507 ( \41851 , \29806 , \30256 );
nor \U$41508 ( \41852 , \41850 , \41851 );
xnor \U$41509 ( \41853 , \41852 , \29948 );
and \U$41510 ( \41854 , \30986 , \29721 );
and \U$41511 ( \41855 , \30383 , \29719 );
nor \U$41512 ( \41856 , \41854 , \41855 );
xnor \U$41513 ( \41857 , \41856 , \29350 );
and \U$41514 ( \41858 , \41853 , \41857 );
and \U$41515 ( \41859 , \31172 , \29159 );
and \U$41516 ( \41860 , \30991 , \29157 );
nor \U$41517 ( \41861 , \41859 , \41860 );
xnor \U$41518 ( \41862 , \41861 , \28841 );
and \U$41519 ( \41863 , \41857 , \41862 );
and \U$41520 ( \41864 , \41853 , \41862 );
or \U$41521 ( \41865 , \41858 , \41863 , \41864 );
and \U$41522 ( \41866 , \29198 , \31639 );
and \U$41523 ( \41867 , \28952 , \31636 );
nor \U$41524 ( \41868 , \41866 , \41867 );
xnor \U$41525 ( \41869 , \41868 , \30584 );
and \U$41526 ( \41870 , \29522 , \30826 );
and \U$41527 ( \41871 , \29203 , \30824 );
nor \U$41528 ( \41872 , \41870 , \41871 );
xnor \U$41529 ( \41873 , \41872 , \30587 );
and \U$41530 ( \41874 , \41869 , \41873 );
and \U$41531 ( \41875 , \41873 , \28343 );
and \U$41532 ( \41876 , \41869 , \28343 );
or \U$41533 ( \41877 , \41874 , \41875 , \41876 );
and \U$41534 ( \41878 , \41865 , \41877 );
xor \U$41535 ( \41879 , \41782 , \41786 );
xor \U$41536 ( \41880 , \41879 , \41791 );
and \U$41537 ( \41881 , \41877 , \41880 );
and \U$41538 ( \41882 , \41865 , \41880 );
or \U$41539 ( \41883 , \41878 , \41881 , \41882 );
xor \U$41540 ( \41884 , \41794 , \41810 );
xor \U$41541 ( \41885 , \41884 , \41815 );
and \U$41542 ( \41886 , \41883 , \41885 );
xor \U$41543 ( \41887 , \41820 , \41822 );
xor \U$41544 ( \41888 , \41887 , \41825 );
and \U$41545 ( \41889 , \41885 , \41888 );
and \U$41546 ( \41890 , \41883 , \41888 );
or \U$41547 ( \41891 , \41886 , \41889 , \41890 );
xor \U$41548 ( \41892 , \41818 , \41828 );
xor \U$41549 ( \41893 , \41892 , \41831 );
and \U$41550 ( \41894 , \41891 , \41893 );
xor \U$41551 ( \41895 , \41836 , \41838 );
and \U$41552 ( \41896 , \41893 , \41895 );
and \U$41553 ( \41897 , \41891 , \41895 );
or \U$41554 ( \41898 , \41894 , \41896 , \41897 );
and \U$41555 ( \41899 , \41849 , \41898 );
xor \U$41556 ( \41900 , \41849 , \41898 );
xor \U$41557 ( \41901 , \41891 , \41893 );
xor \U$41558 ( \41902 , \41901 , \41895 );
and \U$41559 ( \41903 , \29203 , \31639 );
and \U$41560 ( \41904 , \29198 , \31636 );
nor \U$41561 ( \41905 , \41903 , \41904 );
xnor \U$41562 ( \41906 , \41905 , \30584 );
and \U$41563 ( \41907 , \29806 , \30826 );
and \U$41564 ( \41908 , \29522 , \30824 );
nor \U$41565 ( \41909 , \41907 , \41908 );
xnor \U$41566 ( \41910 , \41909 , \30587 );
and \U$41567 ( \41911 , \41906 , \41910 );
and \U$41568 ( \41912 , \30383 , \30258 );
and \U$41569 ( \41913 , \30375 , \30256 );
nor \U$41570 ( \41914 , \41912 , \41913 );
xnor \U$41571 ( \41915 , \41914 , \29948 );
and \U$41572 ( \41916 , \41910 , \41915 );
and \U$41573 ( \41917 , \41906 , \41915 );
or \U$41574 ( \41918 , \41911 , \41916 , \41917 );
nand \U$41575 ( \41919 , \31792 , \28590 );
xnor \U$41576 ( \41920 , \41919 , \28343 );
and \U$41577 ( \41921 , \41918 , \41920 );
xor \U$41578 ( \41922 , \41853 , \41857 );
xor \U$41579 ( \41923 , \41922 , \41862 );
and \U$41580 ( \41924 , \41920 , \41923 );
and \U$41581 ( \41925 , \41918 , \41923 );
or \U$41582 ( \41926 , \41921 , \41924 , \41925 );
xor \U$41583 ( \41927 , \41798 , \41802 );
xor \U$41584 ( \41928 , \41927 , \41807 );
and \U$41585 ( \41929 , \41926 , \41928 );
xor \U$41586 ( \41930 , \41865 , \41877 );
xor \U$41587 ( \41931 , \41930 , \41880 );
and \U$41588 ( \41932 , \41928 , \41931 );
and \U$41589 ( \41933 , \41926 , \41931 );
or \U$41590 ( \41934 , \41929 , \41932 , \41933 );
xor \U$41591 ( \41935 , \41883 , \41885 );
xor \U$41592 ( \41936 , \41935 , \41888 );
and \U$41593 ( \41937 , \41934 , \41936 );
and \U$41594 ( \41938 , \41902 , \41937 );
xor \U$41595 ( \41939 , \41902 , \41937 );
xor \U$41596 ( \41940 , \41934 , \41936 );
and \U$41597 ( \41941 , \30986 , \30258 );
and \U$41598 ( \41942 , \30383 , \30256 );
nor \U$41599 ( \41943 , \41941 , \41942 );
xnor \U$41600 ( \41944 , \41943 , \29948 );
and \U$41601 ( \41945 , \31172 , \29721 );
and \U$41602 ( \41946 , \30991 , \29719 );
nor \U$41603 ( \41947 , \41945 , \41946 );
xnor \U$41604 ( \41948 , \41947 , \29350 );
and \U$41605 ( \41949 , \41944 , \41948 );
nand \U$41606 ( \41950 , \31792 , \29157 );
xnor \U$41607 ( \41951 , \41950 , \28841 );
and \U$41608 ( \41952 , \41948 , \41951 );
and \U$41609 ( \41953 , \41944 , \41951 );
or \U$41610 ( \41954 , \41949 , \41952 , \41953 );
and \U$41611 ( \41955 , \29522 , \31639 );
and \U$41612 ( \41956 , \29203 , \31636 );
nor \U$41613 ( \41957 , \41955 , \41956 );
xnor \U$41614 ( \41958 , \41957 , \30584 );
and \U$41615 ( \41959 , \30375 , \30826 );
and \U$41616 ( \41960 , \29806 , \30824 );
nor \U$41617 ( \41961 , \41959 , \41960 );
xnor \U$41618 ( \41962 , \41961 , \30587 );
and \U$41619 ( \41963 , \41958 , \41962 );
and \U$41620 ( \41964 , \41962 , \28841 );
and \U$41621 ( \41965 , \41958 , \28841 );
or \U$41622 ( \41966 , \41963 , \41964 , \41965 );
and \U$41623 ( \41967 , \41954 , \41966 );
and \U$41624 ( \41968 , \30991 , \29721 );
and \U$41625 ( \41969 , \30986 , \29719 );
nor \U$41626 ( \41970 , \41968 , \41969 );
xnor \U$41627 ( \41971 , \41970 , \29350 );
and \U$41628 ( \41972 , \41966 , \41971 );
and \U$41629 ( \41973 , \41954 , \41971 );
or \U$41630 ( \41974 , \41967 , \41972 , \41973 );
and \U$41631 ( \41975 , \31792 , \29159 );
and \U$41632 ( \41976 , \31172 , \29157 );
nor \U$41633 ( \41977 , \41975 , \41976 );
xnor \U$41634 ( \41978 , \41977 , \28841 );
xor \U$41635 ( \41979 , \41906 , \41910 );
xor \U$41636 ( \41980 , \41979 , \41915 );
and \U$41637 ( \41981 , \41978 , \41980 );
and \U$41638 ( \41982 , \41974 , \41981 );
xor \U$41639 ( \41983 , \41869 , \41873 );
xor \U$41640 ( \41984 , \41983 , \28343 );
and \U$41641 ( \41985 , \41981 , \41984 );
and \U$41642 ( \41986 , \41974 , \41984 );
or \U$41643 ( \41987 , \41982 , \41985 , \41986 );
xor \U$41644 ( \41988 , \41926 , \41928 );
xor \U$41645 ( \41989 , \41988 , \41931 );
and \U$41646 ( \41990 , \41987 , \41989 );
and \U$41647 ( \41991 , \41940 , \41990 );
xor \U$41648 ( \41992 , \41940 , \41990 );
xor \U$41649 ( \41993 , \41987 , \41989 );
xor \U$41650 ( \41994 , \41918 , \41920 );
xor \U$41651 ( \41995 , \41994 , \41923 );
xor \U$41652 ( \41996 , \41974 , \41981 );
xor \U$41653 ( \41997 , \41996 , \41984 );
and \U$41654 ( \41998 , \41995 , \41997 );
and \U$41655 ( \41999 , \41993 , \41998 );
xor \U$41656 ( \42000 , \41993 , \41998 );
xor \U$41657 ( \42001 , \41995 , \41997 );
and \U$41658 ( \42002 , \29806 , \31639 );
and \U$41659 ( \42003 , \29522 , \31636 );
nor \U$41660 ( \42004 , \42002 , \42003 );
xnor \U$41661 ( \42005 , \42004 , \30584 );
and \U$41662 ( \42006 , \30383 , \30826 );
and \U$41663 ( \42007 , \30375 , \30824 );
nor \U$41664 ( \42008 , \42006 , \42007 );
xnor \U$41665 ( \42009 , \42008 , \30587 );
and \U$41666 ( \42010 , \42005 , \42009 );
and \U$41667 ( \42011 , \30991 , \30258 );
and \U$41668 ( \42012 , \30986 , \30256 );
nor \U$41669 ( \42013 , \42011 , \42012 );
xnor \U$41670 ( \42014 , \42013 , \29948 );
and \U$41671 ( \42015 , \42009 , \42014 );
and \U$41672 ( \42016 , \42005 , \42014 );
or \U$41673 ( \42017 , \42010 , \42015 , \42016 );
xor \U$41674 ( \42018 , \41944 , \41948 );
xor \U$41675 ( \42019 , \42018 , \41951 );
and \U$41676 ( \42020 , \42017 , \42019 );
xor \U$41677 ( \42021 , \41958 , \41962 );
xor \U$41678 ( \42022 , \42021 , \28841 );
and \U$41679 ( \42023 , \42019 , \42022 );
and \U$41680 ( \42024 , \42017 , \42022 );
or \U$41681 ( \42025 , \42020 , \42023 , \42024 );
xor \U$41682 ( \42026 , \41954 , \41966 );
xor \U$41683 ( \42027 , \42026 , \41971 );
and \U$41684 ( \42028 , \42025 , \42027 );
xor \U$41685 ( \42029 , \41978 , \41980 );
and \U$41686 ( \42030 , \42027 , \42029 );
and \U$41687 ( \42031 , \42025 , \42029 );
or \U$41688 ( \42032 , \42028 , \42030 , \42031 );
and \U$41689 ( \42033 , \42001 , \42032 );
xor \U$41690 ( \42034 , \42001 , \42032 );
xor \U$41691 ( \42035 , \42025 , \42027 );
xor \U$41692 ( \42036 , \42035 , \42029 );
and \U$41693 ( \42037 , \30375 , \31639 );
and \U$41694 ( \42038 , \29806 , \31636 );
nor \U$41695 ( \42039 , \42037 , \42038 );
xnor \U$41696 ( \42040 , \42039 , \30584 );
and \U$41697 ( \42041 , \30986 , \30826 );
and \U$41698 ( \42042 , \30383 , \30824 );
nor \U$41699 ( \42043 , \42041 , \42042 );
xnor \U$41700 ( \42044 , \42043 , \30587 );
and \U$41701 ( \42045 , \42040 , \42044 );
and \U$41702 ( \42046 , \42044 , \29350 );
and \U$41703 ( \42047 , \42040 , \29350 );
or \U$41704 ( \42048 , \42045 , \42046 , \42047 );
and \U$41705 ( \42049 , \31172 , \30258 );
and \U$41706 ( \42050 , \30991 , \30256 );
nor \U$41707 ( \42051 , \42049 , \42050 );
xnor \U$41708 ( \42052 , \42051 , \29948 );
nand \U$41709 ( \42053 , \31792 , \29719 );
xnor \U$41710 ( \42054 , \42053 , \29350 );
and \U$41711 ( \42055 , \42052 , \42054 );
and \U$41712 ( \42056 , \42048 , \42055 );
and \U$41713 ( \42057 , \31792 , \29721 );
and \U$41714 ( \42058 , \31172 , \29719 );
nor \U$41715 ( \42059 , \42057 , \42058 );
xnor \U$41716 ( \42060 , \42059 , \29350 );
and \U$41717 ( \42061 , \42055 , \42060 );
and \U$41718 ( \42062 , \42048 , \42060 );
or \U$41719 ( \42063 , \42056 , \42061 , \42062 );
xor \U$41720 ( \42064 , \42017 , \42019 );
xor \U$41721 ( \42065 , \42064 , \42022 );
and \U$41722 ( \42066 , \42063 , \42065 );
and \U$41723 ( \42067 , \42036 , \42066 );
xor \U$41724 ( \42068 , \42036 , \42066 );
xor \U$41725 ( \42069 , \42063 , \42065 );
xor \U$41726 ( \42070 , \42005 , \42009 );
xor \U$41727 ( \42071 , \42070 , \42014 );
xor \U$41728 ( \42072 , \42048 , \42055 );
xor \U$41729 ( \42073 , \42072 , \42060 );
and \U$41730 ( \42074 , \42071 , \42073 );
and \U$41731 ( \42075 , \42069 , \42074 );
xor \U$41732 ( \42076 , \42069 , \42074 );
xor \U$41733 ( \42077 , \42071 , \42073 );
and \U$41734 ( \42078 , \30383 , \31639 );
and \U$41735 ( \42079 , \30375 , \31636 );
nor \U$41736 ( \42080 , \42078 , \42079 );
xnor \U$41737 ( \42081 , \42080 , \30584 );
and \U$41738 ( \42082 , \30991 , \30826 );
and \U$41739 ( \42083 , \30986 , \30824 );
nor \U$41740 ( \42084 , \42082 , \42083 );
xnor \U$41741 ( \42085 , \42084 , \30587 );
and \U$41742 ( \42086 , \42081 , \42085 );
and \U$41743 ( \42087 , \31792 , \30258 );
and \U$41744 ( \42088 , \31172 , \30256 );
nor \U$41745 ( \42089 , \42087 , \42088 );
xnor \U$41746 ( \42090 , \42089 , \29948 );
and \U$41747 ( \42091 , \42085 , \42090 );
and \U$41748 ( \42092 , \42081 , \42090 );
or \U$41749 ( \42093 , \42086 , \42091 , \42092 );
xor \U$41750 ( \42094 , \42040 , \42044 );
xor \U$41751 ( \42095 , \42094 , \29350 );
and \U$41752 ( \42096 , \42093 , \42095 );
xor \U$41753 ( \42097 , \42052 , \42054 );
and \U$41754 ( \42098 , \42095 , \42097 );
and \U$41755 ( \42099 , \42093 , \42097 );
or \U$41756 ( \42100 , \42096 , \42098 , \42099 );
and \U$41757 ( \42101 , \42077 , \42100 );
xor \U$41758 ( \42102 , \42077 , \42100 );
xor \U$41759 ( \42103 , \42093 , \42095 );
xor \U$41760 ( \42104 , \42103 , \42097 );
and \U$41761 ( \42105 , \30986 , \31639 );
and \U$41762 ( \42106 , \30383 , \31636 );
nor \U$41763 ( \42107 , \42105 , \42106 );
xnor \U$41764 ( \42108 , \42107 , \30584 );
and \U$41765 ( \42109 , \31172 , \30826 );
and \U$41766 ( \42110 , \30991 , \30824 );
nor \U$41767 ( \42111 , \42109 , \42110 );
xnor \U$41768 ( \42112 , \42111 , \30587 );
and \U$41769 ( \42113 , \42108 , \42112 );
and \U$41770 ( \42114 , \42112 , \29948 );
and \U$41771 ( \42115 , \42108 , \29948 );
or \U$41772 ( \42116 , \42113 , \42114 , \42115 );
xor \U$41773 ( \42117 , \42081 , \42085 );
xor \U$41774 ( \42118 , \42117 , \42090 );
and \U$41775 ( \42119 , \42116 , \42118 );
and \U$41776 ( \42120 , \42104 , \42119 );
xor \U$41777 ( \42121 , \42104 , \42119 );
xor \U$41778 ( \42122 , \42116 , \42118 );
nand \U$41779 ( \42123 , \31792 , \30256 );
xnor \U$41780 ( \42124 , \42123 , \29948 );
xor \U$41781 ( \42125 , \42108 , \42112 );
xor \U$41782 ( \42126 , \42125 , \29948 );
and \U$41783 ( \42127 , \42124 , \42126 );
and \U$41784 ( \42128 , \42122 , \42127 );
xor \U$41785 ( \42129 , \42122 , \42127 );
xor \U$41786 ( \42130 , \42124 , \42126 );
and \U$41787 ( \42131 , \30991 , \31639 );
and \U$41788 ( \42132 , \30986 , \31636 );
nor \U$41789 ( \42133 , \42131 , \42132 );
xnor \U$41790 ( \42134 , \42133 , \30584 );
and \U$41791 ( \42135 , \31792 , \30826 );
and \U$41792 ( \42136 , \31172 , \30824 );
nor \U$41793 ( \42137 , \42135 , \42136 );
xnor \U$41794 ( \42138 , \42137 , \30587 );
and \U$41795 ( \42139 , \42134 , \42138 );
and \U$41796 ( \42140 , \42130 , \42139 );
xor \U$41797 ( \42141 , \42130 , \42139 );
xor \U$41798 ( \42142 , \42134 , \42138 );
and \U$41799 ( \42143 , \31172 , \31639 );
and \U$41800 ( \42144 , \30991 , \31636 );
nor \U$41801 ( \42145 , \42143 , \42144 );
xnor \U$41802 ( \42146 , \42145 , \30584 );
and \U$41803 ( \42147 , \42146 , \30587 );
and \U$41804 ( \42148 , \42142 , \42147 );
xor \U$41805 ( \42149 , \42142 , \42147 );
nand \U$41806 ( \42150 , \31792 , \30824 );
xnor \U$41807 ( \42151 , \42150 , \30587 );
xor \U$41808 ( \42152 , \42146 , \30587 );
and \U$41809 ( \42153 , \42151 , \42152 );
xor \U$41810 ( \42154 , \42151 , \42152 );
and \U$41811 ( \42155 , \31792 , \31639 );
and \U$41812 ( \42156 , \31172 , \31636 );
nor \U$41813 ( \42157 , \42155 , \42156 );
xnor \U$41814 ( \42158 , \42157 , \30584 );
nand \U$41815 ( \42159 , \31792 , \31636 );
xnor \U$41816 ( \42160 , \42159 , \30584 );
and \U$41817 ( \42161 , \42160 , \30584 );
and \U$41818 ( \42162 , \42158 , \42161 );
and \U$41819 ( \42163 , \42154 , \42162 );
or \U$41820 ( \42164 , \42153 , \42163 );
and \U$41821 ( \42165 , \42149 , \42164 );
or \U$41822 ( \42166 , \42148 , \42165 );
and \U$41823 ( \42167 , \42141 , \42166 );
or \U$41824 ( \42168 , \42140 , \42167 );
and \U$41825 ( \42169 , \42129 , \42168 );
or \U$41826 ( \42170 , \42128 , \42169 );
and \U$41827 ( \42171 , \42121 , \42170 );
or \U$41828 ( \42172 , \42120 , \42171 );
and \U$41829 ( \42173 , \42102 , \42172 );
or \U$41830 ( \42174 , \42101 , \42173 );
and \U$41831 ( \42175 , \42076 , \42174 );
or \U$41832 ( \42176 , \42075 , \42175 );
and \U$41833 ( \42177 , \42068 , \42176 );
or \U$41834 ( \42178 , \42067 , \42177 );
and \U$41835 ( \42179 , \42034 , \42178 );
or \U$41836 ( \42180 , \42033 , \42179 );
and \U$41837 ( \42181 , \42000 , \42180 );
or \U$41838 ( \42182 , \41999 , \42181 );
and \U$41839 ( \42183 , \41992 , \42182 );
or \U$41840 ( \42184 , \41991 , \42183 );
and \U$41841 ( \42185 , \41939 , \42184 );
or \U$41842 ( \42186 , \41938 , \42185 );
and \U$41843 ( \42187 , \41900 , \42186 );
or \U$41844 ( \42188 , \41899 , \42187 );
and \U$41845 ( \42189 , \41847 , \42188 );
or \U$41846 ( \42190 , \41846 , \42189 );
and \U$41847 ( \42191 , \41776 , \42190 );
or \U$41848 ( \42192 , \41775 , \42191 );
and \U$41849 ( \42193 , \41721 , \42192 );
or \U$41850 ( \42194 , \41720 , \42193 );
and \U$41851 ( \42195 , \41662 , \42194 );
or \U$41852 ( \42196 , \41661 , \42195 );
and \U$41853 ( \42197 , \41654 , \42196 );
or \U$41854 ( \42198 , \41653 , \42197 );
and \U$41855 ( \42199 , \41575 , \42198 );
or \U$41856 ( \42200 , \41574 , \42199 );
and \U$41857 ( \42201 , \41495 , \42200 );
or \U$41858 ( \42202 , \41494 , \42201 );
and \U$41859 ( \42203 , \41400 , \42202 );
or \U$41860 ( \42204 , \41399 , \42203 );
and \U$41861 ( \42205 , \41312 , \42204 );
or \U$41862 ( \42206 , \41311 , \42205 );
and \U$41863 ( \42207 , \41220 , \42206 );
or \U$41864 ( \42208 , \41219 , \42207 );
and \U$41865 ( \42209 , \41132 , \42208 );
or \U$41866 ( \42210 , \41131 , \42209 );
and \U$41867 ( \42211 , \41017 , \42210 );
or \U$41868 ( \42212 , \41016 , \42211 );
and \U$41869 ( \42213 , \40921 , \42212 );
or \U$41870 ( \42214 , \40920 , \42213 );
and \U$41871 ( \42215 , \40913 , \42214 );
or \U$41872 ( \42216 , \40912 , \42215 );
and \U$41873 ( \42217 , \40798 , \42216 );
or \U$41874 ( \42218 , \40797 , \42217 );
and \U$41875 ( \42219 , \40674 , \42218 );
or \U$41876 ( \42220 , \40673 , \42219 );
and \U$41877 ( \42221 , \40534 , \42220 );
or \U$41878 ( \42222 , \40533 , \42221 );
and \U$41879 ( \42223 , \40410 , \42222 );
or \U$41880 ( \42224 , \40409 , \42223 );
and \U$41881 ( \42225 , \40266 , \42224 );
or \U$41882 ( \42226 , \40265 , \42225 );
and \U$41883 ( \42227 , \40141 , \42226 );
or \U$41884 ( \42228 , \40140 , \42227 );
and \U$41885 ( \42229 , \40002 , \42228 );
or \U$41886 ( \42230 , \40001 , \42229 );
and \U$41887 ( \42231 , \39838 , \42230 );
or \U$41888 ( \42232 , \39837 , \42231 );
and \U$41889 ( \42233 , \39686 , \42232 );
or \U$41890 ( \42234 , \39685 , \42233 );
and \U$41891 ( \42235 , \39546 , \42234 );
or \U$41892 ( \42236 , \39545 , \42235 );
and \U$41893 ( \42237 , \39378 , \42236 );
or \U$41894 ( \42238 , \39377 , \42237 );
and \U$41895 ( \42239 , \39370 , \42238 );
or \U$41896 ( \42240 , \39369 , \42239 );
and \U$41897 ( \42241 , \39199 , \42240 );
or \U$41898 ( \42242 , \39198 , \42241 );
and \U$41899 ( \42243 , \39023 , \42242 );
or \U$41900 ( \42244 , \39022 , \42243 );
and \U$41901 ( \42245 , \38833 , \42244 );
or \U$41902 ( \42246 , \38832 , \42245 );
and \U$41903 ( \42247 , \38646 , \42246 );
or \U$41904 ( \42248 , \38645 , \42247 );
and \U$41905 ( \42249 , \38461 , \42248 );
or \U$41906 ( \42250 , \38460 , \42249 );
and \U$41907 ( \42251 , \38253 , \42250 );
or \U$41908 ( \42252 , \38252 , \42251 );
and \U$41909 ( \42253 , \38057 , \42252 );
or \U$41910 ( \42254 , \38056 , \42253 );
and \U$41911 ( \42255 , \37860 , \42254 );
or \U$41912 ( \42256 , \37859 , \42255 );
and \U$41913 ( \42257 , \37647 , \42256 );
or \U$41914 ( \42258 , \37646 , \42257 );
and \U$41915 ( \42259 , \37436 , \42258 );
or \U$41916 ( \42260 , \37435 , \42259 );
and \U$41917 ( \42261 , \37205 , \42260 );
or \U$41918 ( \42262 , \37204 , \42261 );
and \U$41919 ( \42263 , \36975 , \42262 );
or \U$41920 ( \42264 , \36974 , \42263 );
and \U$41921 ( \42265 , \36756 , \42264 );
or \U$41922 ( \42266 , \36755 , \42265 );
and \U$41923 ( \42267 , \36531 , \42266 );
or \U$41924 ( \42268 , \36530 , \42267 );
and \U$41925 ( \42269 , \36281 , \42268 );
or \U$41926 ( \42270 , \36280 , \42269 );
and \U$41927 ( \42271 , \36051 , \42270 );
or \U$41928 ( \42272 , \36050 , \42271 );
and \U$41929 ( \42273 , \35805 , \42272 );
or \U$41930 ( \42274 , \35804 , \42273 );
and \U$41931 ( \42275 , \35797 , \42274 );
or \U$41932 ( \42276 , \35796 , \42275 );
and \U$41933 ( \42277 , \35536 , \42276 );
or \U$41934 ( \42278 , \35535 , \42277 );
and \U$41935 ( \42279 , \35274 , \42278 );
or \U$41936 ( \42280 , \35273 , \42279 );
and \U$41937 ( \42281 , \35004 , \42280 );
or \U$41938 ( \42282 , \35003 , \42281 );
and \U$41939 ( \42283 , \34727 , \42282 );
or \U$41940 ( \42284 , \34726 , \42283 );
and \U$41941 ( \42285 , \34451 , \42284 );
or \U$41942 ( \42286 , \34450 , \42285 );
and \U$41943 ( \42287 , \34180 , \42286 );
or \U$41944 ( \42288 , \34179 , \42287 );
and \U$41945 ( \42289 , \33877 , \42288 );
or \U$41946 ( \42290 , \33876 , \42289 );
and \U$41947 ( \42291 , \33598 , \42290 );
or \U$41948 ( \42292 , \33597 , \42291 );
and \U$41949 ( \42293 , \33313 , \42292 );
or \U$41950 ( \42294 , \33312 , \42293 );
and \U$41951 ( \42295 , \32997 , \42294 );
or \U$41952 ( \42296 , \32996 , \42295 );
and \U$41953 ( \42297 , \32697 , \42296 );
or \U$41954 ( \42298 , \32696 , \42297 );
and \U$41955 ( \42299 , \32381 , \42298 );
or \U$41956 ( \42300 , \32380 , \42299 );
and \U$41957 ( \42301 , \32063 , \42300 );
or \U$41958 ( \42302 , \32062 , \42301 );
and \U$41959 ( \42303 , \31752 , \42302 );
or \U$41960 ( \42304 , \31751 , \42303 );
and \U$41961 ( \42305 , \31439 , \42304 );
or \U$41962 ( \42306 , \31438 , \42305 );
and \U$41963 ( \42307 , \31123 , \42306 );
or \U$41964 ( \42308 , \31122 , \42307 );
and \U$41965 ( \42309 , \30805 , \42308 );
or \U$41966 ( \42310 , \30804 , \42309 );
and \U$41967 ( \42311 , \30496 , \42310 );
or \U$41968 ( \42312 , \30495 , \42311 );
and \U$41969 ( \42313 , \30200 , \42312 );
or \U$41970 ( \42314 , \30199 , \42313 );
and \U$41971 ( \42315 , \29899 , \42314 );
or \U$41972 ( \42316 , \29898 , \42315 );
and \U$41973 ( \42317 , \29611 , \42316 );
or \U$41974 ( \42318 , \29610 , \42317 );
and \U$41975 ( \42319 , \29328 , \42318 );
or \U$41976 ( \42320 , \29327 , \42319 );
and \U$41977 ( \42321 , \29033 , \42320 );
or \U$41978 ( \42322 , \29032 , \42321 );
and \U$41979 ( \42323 , \28767 , \42322 );
or \U$41980 ( \42324 , \28766 , \42323 );
and \U$41981 ( \42325 , \28501 , \42324 );
or \U$41982 ( \42326 , \28500 , \42325 );
and \U$41983 ( \42327 , \28240 , \42326 );
or \U$41984 ( \42328 , \28239 , \42327 );
and \U$41985 ( \42329 , \27975 , \42328 );
or \U$41986 ( \42330 , \27974 , \42329 );
and \U$41987 ( \42331 , \27712 , \42330 );
or \U$41988 ( \42332 , \27711 , \42331 );
and \U$41989 ( \42333 , \27455 , \42332 );
or \U$41990 ( \42334 , \27454 , \42333 );
and \U$41991 ( \42335 , \27199 , \42334 );
or \U$41992 ( \42336 , \27198 , \42335 );
and \U$41993 ( \42337 , \26946 , \42336 );
or \U$41994 ( \42338 , \26945 , \42337 );
and \U$41995 ( \42339 , \26698 , \42338 );
or \U$41996 ( \42340 , \26697 , \42339 );
and \U$41997 ( \42341 , \26466 , \42340 );
or \U$41998 ( \42342 , \26465 , \42341 );
and \U$41999 ( \42343 , \26223 , \42342 );
or \U$42000 ( \42344 , \26222 , \42343 );
and \U$42001 ( \42345 , \25794 , \42344 );
or \U$42002 ( \42346 , \25793 , \42345 );
and \U$42003 ( \42347 , \25584 , \42346 );
or \U$42004 ( \42348 , \25583 , \42347 );
and \U$42005 ( \42349 , \25377 , \42348 );
or \U$42006 ( \42350 , \25376 , \42349 );
and \U$42007 ( \42351 , \25175 , \42350 );
or \U$42008 ( \42352 , \25174 , \42351 );
and \U$42009 ( \42353 , \24979 , \42352 );
or \U$42010 ( \42354 , \24978 , \42353 );
and \U$42011 ( \42355 , \24782 , \42354 );
or \U$42012 ( \42356 , \24781 , \42355 );
and \U$42013 ( \42357 , \24605 , \42356 );
or \U$42014 ( \42358 , \24604 , \42357 );
and \U$42015 ( \42359 , \24424 , \42358 );
or \U$42016 ( \42360 , \24423 , \42359 );
and \U$42017 ( \42361 , \24253 , \42360 );
or \U$42018 ( \42362 , \24252 , \42361 );
and \U$42019 ( \42363 , \24078 , \42362 );
or \U$42020 ( \42364 , \24077 , \42363 );
and \U$42021 ( \42365 , \23905 , \42364 );
or \U$42022 ( \42366 , \23904 , \42365 );
and \U$42023 ( \42367 , \23738 , \42366 );
or \U$42024 ( \42368 , \23737 , \42367 );
and \U$42025 ( \42369 , \23572 , \42368 );
or \U$42026 ( \42370 , \23571 , \42369 );
and \U$42027 ( \42371 , \23399 , \42370 );
or \U$42028 ( \42372 , \23398 , \42371 );
and \U$42029 ( \42373 , \23119 , \42372 );
or \U$42030 ( \42374 , \23118 , \42373 );
and \U$42031 ( \42375 , \22982 , \42374 );
or \U$42032 ( \42376 , \22981 , \42375 );
and \U$42033 ( \42377 , \22849 , \42376 );
or \U$42034 ( \42378 , \22848 , \42377 );
and \U$42035 ( \42379 , \22728 , \42378 );
or \U$42036 ( \42380 , \22727 , \42379 );
and \U$42037 ( \42381 , \22605 , \42380 );
or \U$42038 ( \42382 , \22604 , \42381 );
and \U$42039 ( \42383 , \22489 , \42382 );
or \U$42040 ( \42384 , \22488 , \42383 );
and \U$42041 ( \42385 , \22374 , \42384 );
or \U$42042 ( \42386 , \22373 , \42385 );
and \U$42043 ( \42387 , \22260 , \42386 );
or \U$42044 ( \42388 , \22259 , \42387 );
and \U$42045 ( \42389 , \22146 , \42388 );
or \U$42046 ( \42390 , \22145 , \42389 );
and \U$42047 ( \42391 , \21964 , \42390 );
or \U$42048 ( \42392 , \21963 , \42391 );
and \U$42049 ( \42393 , \21885 , \42392 );
or \U$42050 ( \42394 , \21884 , \42393 );
and \U$42051 ( \42395 , \21802 , \42394 );
or \U$42052 ( \42396 , \21801 , \42395 );
xor \U$42053 ( \42397 , \21721 , \42396 );
buf gac83_GF_PartitionCandidate( \42398_nGac83 , \42397 );
buf \U$42054 ( \42399 , \42398_nGac83 );
xor \U$42055 ( \42400 , \21371 , \42399 );
xor \U$42056 ( \42401 , \774 , \21366 );
buf gabce_GF_PartitionCandidate( \42402_nGabce , \42401 );
buf \U$42057 ( \42403 , \42402_nGabce );
xor \U$42058 ( \42404 , \21802 , \42394 );
buf gac0d_GF_PartitionCandidate( \42405_nGac0d , \42404 );
buf \U$42059 ( \42406 , \42405_nGac0d );
and \U$42060 ( \42407 , \42403 , \42406 );
xor \U$42061 ( \42408 , \857 , \21364 );
buf gab43_GF_PartitionCandidate( \42409_nGab43 , \42408 );
buf \U$42062 ( \42410 , \42409_nGab43 );
xor \U$42063 ( \42411 , \21885 , \42392 );
buf gab87_GF_PartitionCandidate( \42412_nGab87 , \42411 );
buf \U$42064 ( \42413 , \42412_nGab87 );
and \U$42065 ( \42414 , \42410 , \42413 );
xor \U$42066 ( \42415 , \936 , \21362 );
buf gaab0_GF_PartitionCandidate( \42416_nGaab0 , \42415 );
buf \U$42067 ( \42417 , \42416_nGaab0 );
xor \U$42068 ( \42418 , \21964 , \42390 );
buf gaaf7_GF_PartitionCandidate( \42419_nGaaf7 , \42418 );
buf \U$42069 ( \42420 , \42419_nGaaf7 );
and \U$42070 ( \42421 , \42417 , \42420 );
xor \U$42071 ( \42422 , \1118 , \21360 );
buf gaa15_GF_PartitionCandidate( \42423_nGaa15 , \42422 );
buf \U$42072 ( \42424 , \42423_nGaa15 );
xor \U$42073 ( \42425 , \22146 , \42388 );
buf gaa61_GF_PartitionCandidate( \42426_nGaa61 , \42425 );
buf \U$42074 ( \42427 , \42426_nGaa61 );
and \U$42075 ( \42428 , \42424 , \42427 );
xor \U$42076 ( \42429 , \1232 , \21358 );
buf ga96e_GF_PartitionCandidate( \42430_nGa96e , \42429 );
buf \U$42077 ( \42431 , \42430_nGa96e );
xor \U$42078 ( \42432 , \22260 , \42386 );
buf ga9c1_GF_PartitionCandidate( \42433_nGa9c1 , \42432 );
buf \U$42079 ( \42434 , \42433_nGa9c1 );
and \U$42080 ( \42435 , \42431 , \42434 );
xor \U$42081 ( \42436 , \1346 , \21356 );
buf ga8be_GF_PartitionCandidate( \42437_nGa8be , \42436 );
buf \U$42082 ( \42438 , \42437_nGa8be );
xor \U$42083 ( \42439 , \22374 , \42384 );
buf ga913_GF_PartitionCandidate( \42440_nGa913 , \42439 );
buf \U$42084 ( \42441 , \42440_nGa913 );
and \U$42085 ( \42442 , \42438 , \42441 );
xor \U$42086 ( \42443 , \1461 , \21354 );
buf ga804_GF_PartitionCandidate( \42444_nGa804 , \42443 );
buf \U$42087 ( \42445 , \42444_nGa804 );
xor \U$42088 ( \42446 , \22489 , \42382 );
buf ga861_GF_PartitionCandidate( \42447_nGa861 , \42446 );
buf \U$42089 ( \42448 , \42447_nGa861 );
and \U$42090 ( \42449 , \42445 , \42448 );
xor \U$42091 ( \42450 , \1577 , \21352 );
buf ga740_GF_PartitionCandidate( \42451_nGa740 , \42450 );
buf \U$42092 ( \42452 , \42451_nGa740 );
xor \U$42093 ( \42453 , \22605 , \42380 );
buf ga79f_GF_PartitionCandidate( \42454_nGa79f , \42453 );
buf \U$42094 ( \42455 , \42454_nGa79f );
and \U$42095 ( \42456 , \42452 , \42455 );
xor \U$42096 ( \42457 , \1700 , \21350 );
buf ga672_GF_PartitionCandidate( \42458_nGa672 , \42457 );
buf \U$42097 ( \42459 , \42458_nGa672 );
xor \U$42098 ( \42460 , \22728 , \42378 );
buf ga6d9_GF_PartitionCandidate( \42461_nGa6d9 , \42460 );
buf \U$42099 ( \42462 , \42461_nGa6d9 );
and \U$42100 ( \42463 , \42459 , \42462 );
xor \U$42101 ( \42464 , \1821 , \21348 );
buf ga59a_GF_PartitionCandidate( \42465_nGa59a , \42464 );
buf \U$42102 ( \42466 , \42465_nGa59a );
xor \U$42103 ( \42467 , \22849 , \42376 );
buf ga603_GF_PartitionCandidate( \42468_nGa603 , \42467 );
buf \U$42104 ( \42469 , \42468_nGa603 );
and \U$42105 ( \42470 , \42466 , \42469 );
xor \U$42106 ( \42471 , \1954 , \21346 );
buf ga4bb_GF_PartitionCandidate( \42472_nGa4bb , \42471 );
buf \U$42107 ( \42473 , \42472_nGa4bb );
xor \U$42108 ( \42474 , \22982 , \42374 );
buf ga529_GF_PartitionCandidate( \42475_nGa529 , \42474 );
buf \U$42109 ( \42476 , \42475_nGa529 );
and \U$42110 ( \42477 , \42473 , \42476 );
xor \U$42111 ( \42478 , \2091 , \21344 );
buf ga3d1_GF_PartitionCandidate( \42479_nGa3d1 , \42478 );
buf \U$42112 ( \42480 , \42479_nGa3d1 );
xor \U$42113 ( \42481 , \23119 , \42372 );
buf ga445_GF_PartitionCandidate( \42482_nGa445 , \42481 );
buf \U$42114 ( \42483 , \42482_nGa445 );
and \U$42115 ( \42484 , \42480 , \42483 );
xor \U$42116 ( \42485 , \2371 , \21342 );
buf ga2da_GF_PartitionCandidate( \42486_nGa2da , \42485 );
buf \U$42117 ( \42487 , \42486_nGa2da );
xor \U$42118 ( \42488 , \23399 , \42370 );
buf ga355_GF_PartitionCandidate( \42489_nGa355 , \42488 );
buf \U$42119 ( \42490 , \42489_nGa355 );
and \U$42120 ( \42491 , \42487 , \42490 );
xor \U$42121 ( \42492 , \2544 , \21340 );
buf ga1d7_GF_PartitionCandidate( \42493_nGa1d7 , \42492 );
buf \U$42122 ( \42494 , \42493_nGa1d7 );
xor \U$42123 ( \42495 , \23572 , \42368 );
buf ga257_GF_PartitionCandidate( \42496_nGa257 , \42495 );
buf \U$42124 ( \42497 , \42496_nGa257 );
and \U$42125 ( \42498 , \42494 , \42497 );
xor \U$42126 ( \42499 , \2710 , \21338 );
buf ga0c9_GF_PartitionCandidate( \42500_nGa0c9 , \42499 );
buf \U$42127 ( \42501 , \42500_nGa0c9 );
xor \U$42128 ( \42502 , \23738 , \42366 );
buf ga14f_GF_PartitionCandidate( \42503_nGa14f , \42502 );
buf \U$42129 ( \42504 , \42503_nGa14f );
and \U$42130 ( \42505 , \42501 , \42504 );
xor \U$42131 ( \42506 , \2877 , \21336 );
buf g9fb4_GF_PartitionCandidate( \42507_nG9fb4 , \42506 );
buf \U$42132 ( \42508 , \42507_nG9fb4 );
xor \U$42133 ( \42509 , \23905 , \42364 );
buf ga03b_GF_PartitionCandidate( \42510_nGa03b , \42509 );
buf \U$42134 ( \42511 , \42510_nGa03b );
and \U$42135 ( \42512 , \42508 , \42511 );
xor \U$42136 ( \42513 , \3050 , \21334 );
buf g9e96_GF_PartitionCandidate( \42514_nG9e96 , \42513 );
buf \U$42137 ( \42515 , \42514_nG9e96 );
xor \U$42138 ( \42516 , \24078 , \42362 );
buf g9f25_GF_PartitionCandidate( \42517_nG9f25 , \42516 );
buf \U$42139 ( \42518 , \42517_nG9f25 );
and \U$42140 ( \42519 , \42515 , \42518 );
xor \U$42141 ( \42520 , \3225 , \21332 );
buf g9d6b_GF_PartitionCandidate( \42521_nG9d6b , \42520 );
buf \U$42142 ( \42522 , \42521_nG9d6b );
xor \U$42143 ( \42523 , \24253 , \42360 );
buf g9dff_GF_PartitionCandidate( \42524_nG9dff , \42523 );
buf \U$42144 ( \42525 , \42524_nG9dff );
and \U$42145 ( \42526 , \42522 , \42525 );
xor \U$42146 ( \42527 , \3396 , \21330 );
buf g9c34_GF_PartitionCandidate( \42528_nG9c34 , \42527 );
buf \U$42147 ( \42529 , \42528_nG9c34 );
xor \U$42148 ( \42530 , \24424 , \42358 );
buf g9ccf_GF_PartitionCandidate( \42531_nG9ccf , \42530 );
buf \U$42149 ( \42532 , \42531_nG9ccf );
and \U$42150 ( \42533 , \42529 , \42532 );
xor \U$42151 ( \42534 , \3577 , \21328 );
buf g9af1_GF_PartitionCandidate( \42535_nG9af1 , \42534 );
buf \U$42152 ( \42536 , \42535_nG9af1 );
xor \U$42153 ( \42537 , \24605 , \42356 );
buf g9b91_GF_PartitionCandidate( \42538_nG9b91 , \42537 );
buf \U$42154 ( \42539 , \42538_nG9b91 );
and \U$42155 ( \42540 , \42536 , \42539 );
xor \U$42156 ( \42541 , \3754 , \21326 );
buf g99a6_GF_PartitionCandidate( \42542_nG99a6 , \42541 );
buf \U$42157 ( \42543 , \42542_nG99a6 );
xor \U$42158 ( \42544 , \24782 , \42354 );
buf g9a49_GF_PartitionCandidate( \42545_nG9a49 , \42544 );
buf \U$42159 ( \42546 , \42545_nG9a49 );
and \U$42160 ( \42547 , \42543 , \42546 );
xor \U$42161 ( \42548 , \3951 , \21324 );
buf g9856_GF_PartitionCandidate( \42549_nG9856 , \42548 );
buf \U$42162 ( \42550 , \42549_nG9856 );
xor \U$42163 ( \42551 , \24979 , \42352 );
buf g98fb_GF_PartitionCandidate( \42552_nG98fb , \42551 );
buf \U$42164 ( \42553 , \42552_nG98fb );
and \U$42165 ( \42554 , \42550 , \42553 );
xor \U$42166 ( \42555 , \4147 , \21322 );
buf g96ff_GF_PartitionCandidate( \42556_nG96ff , \42555 );
buf \U$42167 ( \42557 , \42556_nG96ff );
xor \U$42168 ( \42558 , \25175 , \42350 );
buf g97a9_GF_PartitionCandidate( \42559_nG97a9 , \42558 );
buf \U$42169 ( \42560 , \42559_nG97a9 );
and \U$42170 ( \42561 , \42557 , \42560 );
xor \U$42171 ( \42562 , \4349 , \21320 );
buf g95a0_GF_PartitionCandidate( \42563_nG95a0 , \42562 );
buf \U$42172 ( \42564 , \42563_nG95a0 );
xor \U$42173 ( \42565 , \25377 , \42348 );
buf g964d_GF_PartitionCandidate( \42566_nG964d , \42565 );
buf \U$42174 ( \42567 , \42566_nG964d );
and \U$42175 ( \42568 , \42564 , \42567 );
xor \U$42176 ( \42569 , \4556 , \21318 );
buf g9436_GF_PartitionCandidate( \42570_nG9436 , \42569 );
buf \U$42177 ( \42571 , \42570_nG9436 );
xor \U$42178 ( \42572 , \25584 , \42346 );
buf g94eb_GF_PartitionCandidate( \42573_nG94eb , \42572 );
buf \U$42179 ( \42574 , \42573_nG94eb );
and \U$42180 ( \42575 , \42571 , \42574 );
xor \U$42181 ( \42576 , \4766 , \21316 );
buf g92bf_GF_PartitionCandidate( \42577_nG92bf , \42576 );
buf \U$42182 ( \42578 , \42577_nG92bf );
xor \U$42183 ( \42579 , \25794 , \42344 );
buf g9379_GF_PartitionCandidate( \42580_nG9379 , \42579 );
buf \U$42184 ( \42581 , \42580_nG9379 );
and \U$42185 ( \42582 , \42578 , \42581 );
xor \U$42186 ( \42583 , \5195 , \21314 );
buf g913c_GF_PartitionCandidate( \42584_nG913c , \42583 );
buf \U$42187 ( \42585 , \42584_nG913c );
xor \U$42188 ( \42586 , \26223 , \42342 );
buf g91fd_GF_PartitionCandidate( \42587_nG91fd , \42586 );
buf \U$42189 ( \42588 , \42587_nG91fd );
and \U$42190 ( \42589 , \42585 , \42588 );
xor \U$42191 ( \42590 , \5438 , \21312 );
buf g8fb0_GF_PartitionCandidate( \42591_nG8fb0 , \42590 );
buf \U$42192 ( \42592 , \42591_nG8fb0 );
xor \U$42193 ( \42593 , \26466 , \42340 );
buf g9073_GF_PartitionCandidate( \42594_nG9073 , \42593 );
buf \U$42194 ( \42595 , \42594_nG9073 );
and \U$42195 ( \42596 , \42592 , \42595 );
xor \U$42196 ( \42597 , \5670 , \21310 );
buf g8e1a_GF_PartitionCandidate( \42598_nG8e1a , \42597 );
buf \U$42197 ( \42599 , \42598_nG8e1a );
xor \U$42198 ( \42600 , \26698 , \42338 );
buf g8ee5_GF_PartitionCandidate( \42601_nG8ee5 , \42600 );
buf \U$42199 ( \42602 , \42601_nG8ee5 );
and \U$42200 ( \42603 , \42599 , \42602 );
xor \U$42201 ( \42604 , \5918 , \21308 );
buf g8c7a_GF_PartitionCandidate( \42605_nG8c7a , \42604 );
buf \U$42202 ( \42606 , \42605_nG8c7a );
xor \U$42203 ( \42607 , \26946 , \42336 );
buf g8d47_GF_PartitionCandidate( \42608_nG8d47 , \42607 );
buf \U$42204 ( \42609 , \42608_nG8d47 );
and \U$42205 ( \42610 , \42606 , \42609 );
xor \U$42206 ( \42611 , \6171 , \21306 );
buf g8ad0_GF_PartitionCandidate( \42612_nG8ad0 , \42611 );
buf \U$42207 ( \42613 , \42612_nG8ad0 );
xor \U$42208 ( \42614 , \27199 , \42334 );
buf g8ba5_GF_PartitionCandidate( \42615_nG8ba5 , \42614 );
buf \U$42209 ( \42616 , \42615_nG8ba5 );
and \U$42210 ( \42617 , \42613 , \42616 );
xor \U$42211 ( \42618 , \6427 , \21304 );
buf g8919_GF_PartitionCandidate( \42619_nG8919 , \42618 );
buf \U$42212 ( \42620 , \42619_nG8919 );
xor \U$42213 ( \42621 , \27455 , \42332 );
buf g89f3_GF_PartitionCandidate( \42622_nG89f3 , \42621 );
buf \U$42214 ( \42623 , \42622_nG89f3 );
and \U$42215 ( \42624 , \42620 , \42623 );
xor \U$42216 ( \42625 , \6684 , \21302 );
buf g8757_GF_PartitionCandidate( \42626_nG8757 , \42625 );
buf \U$42217 ( \42627 , \42626_nG8757 );
xor \U$42218 ( \42628 , \27712 , \42330 );
buf g8837_GF_PartitionCandidate( \42629_nG8837 , \42628 );
buf \U$42219 ( \42630 , \42629_nG8837 );
and \U$42220 ( \42631 , \42627 , \42630 );
xor \U$42221 ( \42632 , \6947 , \21300 );
buf g858b_GF_PartitionCandidate( \42633_nG858b , \42632 );
buf \U$42222 ( \42634 , \42633_nG858b );
xor \U$42223 ( \42635 , \27975 , \42328 );
buf g866f_GF_PartitionCandidate( \42636_nG866f , \42635 );
buf \U$42224 ( \42637 , \42636_nG866f );
and \U$42225 ( \42638 , \42634 , \42637 );
xor \U$42226 ( \42639 , \7212 , \21298 );
buf g83b4_GF_PartitionCandidate( \42640_nG83b4 , \42639 );
buf \U$42227 ( \42641 , \42640_nG83b4 );
xor \U$42228 ( \42642 , \28240 , \42326 );
buf g849f_GF_PartitionCandidate( \42643_nG849f , \42642 );
buf \U$42229 ( \42644 , \42643_nG849f );
and \U$42230 ( \42645 , \42641 , \42644 );
xor \U$42231 ( \42646 , \7473 , \21296 );
buf g81d4_GF_PartitionCandidate( \42647_nG81d4 , \42646 );
buf \U$42232 ( \42648 , \42647_nG81d4 );
xor \U$42233 ( \42649 , \28501 , \42324 );
buf g82c1_GF_PartitionCandidate( \42650_nG82c1 , \42649 );
buf \U$42234 ( \42651 , \42650_nG82c1 );
and \U$42235 ( \42652 , \42648 , \42651 );
xor \U$42236 ( \42653 , \7739 , \21294 );
buf g7fea_GF_PartitionCandidate( \42654_nG7fea , \42653 );
buf \U$42237 ( \42655 , \42654_nG7fea );
xor \U$42238 ( \42656 , \28767 , \42322 );
buf g80df_GF_PartitionCandidate( \42657_nG80df , \42656 );
buf \U$42239 ( \42658 , \42657_nG80df );
and \U$42240 ( \42659 , \42655 , \42658 );
xor \U$42241 ( \42660 , \8005 , \21292 );
buf g7df3_GF_PartitionCandidate( \42661_nG7df3 , \42660 );
buf \U$42242 ( \42662 , \42661_nG7df3 );
xor \U$42243 ( \42663 , \29033 , \42320 );
buf g7eed_GF_PartitionCandidate( \42664_nG7eed , \42663 );
buf \U$42244 ( \42665 , \42664_nG7eed );
and \U$42245 ( \42666 , \42662 , \42665 );
xor \U$42246 ( \42667 , \8300 , \21290 );
buf g7bf4_GF_PartitionCandidate( \42668_nG7bf4 , \42667 );
buf \U$42247 ( \42669 , \42668_nG7bf4 );
xor \U$42248 ( \42670 , \29328 , \42318 );
buf g7cf1_GF_PartitionCandidate( \42671_nG7cf1 , \42670 );
buf \U$42249 ( \42672 , \42671_nG7cf1 );
and \U$42250 ( \42673 , \42669 , \42672 );
xor \U$42251 ( \42674 , \8583 , \21288 );
buf g79f0_GF_PartitionCandidate( \42675_nG79f0 , \42674 );
buf \U$42252 ( \42676 , \42675_nG79f0 );
xor \U$42253 ( \42677 , \29611 , \42316 );
buf g7aef_GF_PartitionCandidate( \42678_nG7aef , \42677 );
buf \U$42254 ( \42679 , \42678_nG7aef );
and \U$42255 ( \42680 , \42676 , \42679 );
xor \U$42256 ( \42681 , \8871 , \21286 );
buf g77e5_GF_PartitionCandidate( \42682_nG77e5 , \42681 );
buf \U$42257 ( \42683 , \42682_nG77e5 );
xor \U$42258 ( \42684 , \29899 , \42314 );
buf g78e9_GF_PartitionCandidate( \42685_nG78e9 , \42684 );
buf \U$42259 ( \42686 , \42685_nG78e9 );
and \U$42260 ( \42687 , \42683 , \42686 );
xor \U$42261 ( \42688 , \9172 , \21284 );
buf g75cf_GF_PartitionCandidate( \42689_nG75cf , \42688 );
buf \U$42262 ( \42690 , \42689_nG75cf );
xor \U$42263 ( \42691 , \30200 , \42312 );
buf g76d9_GF_PartitionCandidate( \42692_nG76d9 , \42691 );
buf \U$42264 ( \42693 , \42692_nG76d9 );
and \U$42265 ( \42694 , \42690 , \42693 );
xor \U$42266 ( \42695 , \9468 , \21282 );
buf g73af_GF_PartitionCandidate( \42696_nG73af , \42695 );
buf \U$42267 ( \42697 , \42696_nG73af );
xor \U$42268 ( \42698 , \30496 , \42310 );
buf g74bd_GF_PartitionCandidate( \42699_nG74bd , \42698 );
buf \U$42269 ( \42700 , \42699_nG74bd );
and \U$42270 ( \42701 , \42697 , \42700 );
xor \U$42271 ( \42702 , \9777 , \21280 );
buf g7188_GF_PartitionCandidate( \42703_nG7188 , \42702 );
buf \U$42272 ( \42704 , \42703_nG7188 );
xor \U$42273 ( \42705 , \30805 , \42308 );
buf g7299_GF_PartitionCandidate( \42706_nG7299 , \42705 );
buf \U$42274 ( \42707 , \42706_nG7299 );
and \U$42275 ( \42708 , \42704 , \42707 );
xor \U$42276 ( \42709 , \10095 , \21278 );
buf g6f56_GF_PartitionCandidate( \42710_nG6f56 , \42709 );
buf \U$42277 ( \42711 , \42710_nG6f56 );
xor \U$42278 ( \42712 , \31123 , \42306 );
buf g706f_GF_PartitionCandidate( \42713_nG706f , \42712 );
buf \U$42279 ( \42714 , \42713_nG706f );
and \U$42280 ( \42715 , \42711 , \42714 );
xor \U$42281 ( \42716 , \10411 , \21276 );
buf g6d1a_GF_PartitionCandidate( \42717_nG6d1a , \42716 );
buf \U$42282 ( \42718 , \42717_nG6d1a );
xor \U$42283 ( \42719 , \31439 , \42304 );
buf g6e35_GF_PartitionCandidate( \42720_nG6e35 , \42719 );
buf \U$42284 ( \42721 , \42720_nG6e35 );
and \U$42285 ( \42722 , \42718 , \42721 );
xor \U$42286 ( \42723 , \10724 , \21274 );
buf g6ad4_GF_PartitionCandidate( \42724_nG6ad4 , \42723 );
buf \U$42287 ( \42725 , \42724_nG6ad4 );
xor \U$42288 ( \42726 , \31752 , \42302 );
buf g6bf7_GF_PartitionCandidate( \42727_nG6bf7 , \42726 );
buf \U$42289 ( \42728 , \42727_nG6bf7 );
and \U$42290 ( \42729 , \42725 , \42728 );
xor \U$42291 ( \42730 , \11035 , \21272 );
buf g6881_GF_PartitionCandidate( \42731_nG6881 , \42730 );
buf \U$42292 ( \42732 , \42731_nG6881 );
xor \U$42293 ( \42733 , \32063 , \42300 );
buf g69a9_GF_PartitionCandidate( \42734_nG69a9 , \42733 );
buf \U$42294 ( \42735 , \42734_nG69a9 );
and \U$42295 ( \42736 , \42732 , \42735 );
xor \U$42296 ( \42737 , \11353 , \21270 );
buf g6622_GF_PartitionCandidate( \42738_nG6622 , \42737 );
buf \U$42297 ( \42739 , \42738_nG6622 );
xor \U$42298 ( \42740 , \32381 , \42298 );
buf g6751_GF_PartitionCandidate( \42741_nG6751 , \42740 );
buf \U$42299 ( \42742 , \42741_nG6751 );
and \U$42300 ( \42743 , \42739 , \42742 );
xor \U$42301 ( \42744 , \11669 , \21268 );
buf g63b7_GF_PartitionCandidate( \42745_nG63b7 , \42744 );
buf \U$42302 ( \42746 , \42745_nG63b7 );
xor \U$42303 ( \42747 , \32697 , \42296 );
buf g64eb_GF_PartitionCandidate( \42748_nG64eb , \42747 );
buf \U$42304 ( \42749 , \42748_nG64eb );
and \U$42305 ( \42750 , \42746 , \42749 );
xor \U$42306 ( \42751 , \11969 , \21266 );
buf g6144_GF_PartitionCandidate( \42752_nG6144 , \42751 );
buf \U$42307 ( \42753 , \42752_nG6144 );
xor \U$42308 ( \42754 , \32997 , \42294 );
buf g627b_GF_PartitionCandidate( \42755_nG627b , \42754 );
buf \U$42309 ( \42756 , \42755_nG627b );
and \U$42310 ( \42757 , \42753 , \42756 );
xor \U$42311 ( \42758 , \12285 , \21264 );
buf g5ec9_GF_PartitionCandidate( \42759_nG5ec9 , \42758 );
buf \U$42312 ( \42760 , \42759_nG5ec9 );
xor \U$42313 ( \42761 , \33313 , \42292 );
buf g6005_GF_PartitionCandidate( \42762_nG6005 , \42761 );
buf \U$42314 ( \42763 , \42762_nG6005 );
and \U$42315 ( \42764 , \42760 , \42763 );
xor \U$42316 ( \42765 , \12570 , \21262 );
buf g5c48_GF_PartitionCandidate( \42766_nG5c48 , \42765 );
buf \U$42317 ( \42767 , \42766_nG5c48 );
xor \U$42318 ( \42768 , \33598 , \42290 );
buf g5d85_GF_PartitionCandidate( \42769_nG5d85 , \42768 );
buf \U$42319 ( \42770 , \42769_nG5d85 );
and \U$42320 ( \42771 , \42767 , \42770 );
xor \U$42321 ( \42772 , \12849 , \21260 );
buf g59c5_GF_PartitionCandidate( \42773_nG59c5 , \42772 );
buf \U$42322 ( \42774 , \42773_nG59c5 );
xor \U$42323 ( \42775 , \33877 , \42288 );
buf g5b03_GF_PartitionCandidate( \42776_nG5b03 , \42775 );
buf \U$42324 ( \42777 , \42776_nG5b03 );
and \U$42325 ( \42778 , \42774 , \42777 );
xor \U$42326 ( \42779 , \13152 , \21258 );
buf g5740_GF_PartitionCandidate( \42780_nG5740 , \42779 );
buf \U$42327 ( \42781 , \42780_nG5740 );
xor \U$42328 ( \42782 , \34180 , \42286 );
buf g587f_GF_PartitionCandidate( \42783_nG587f , \42782 );
buf \U$42329 ( \42784 , \42783_nG587f );
and \U$42330 ( \42785 , \42781 , \42784 );
xor \U$42331 ( \42786 , \13423 , \21256 );
buf g54b8_GF_PartitionCandidate( \42787_nG54b8 , \42786 );
buf \U$42332 ( \42788 , \42787_nG54b8 );
xor \U$42333 ( \42789 , \34451 , \42284 );
buf g55f9_GF_PartitionCandidate( \42790_nG55f9 , \42789 );
buf \U$42334 ( \42791 , \42790_nG55f9 );
and \U$42335 ( \42792 , \42788 , \42791 );
xor \U$42336 ( \42793 , \13699 , \21254 );
buf g5231_GF_PartitionCandidate( \42794_nG5231 , \42793 );
buf \U$42337 ( \42795 , \42794_nG5231 );
xor \U$42338 ( \42796 , \34727 , \42282 );
buf g536f_GF_PartitionCandidate( \42797_nG536f , \42796 );
buf \U$42339 ( \42798 , \42797_nG536f );
and \U$42340 ( \42799 , \42795 , \42798 );
xor \U$42341 ( \42800 , \13976 , \21252 );
buf g4fb4_GF_PartitionCandidate( \42801_nG4fb4 , \42800 );
buf \U$42342 ( \42802 , \42801_nG4fb4 );
xor \U$42343 ( \42803 , \35004 , \42280 );
buf g50eb_GF_PartitionCandidate( \42804_nG50eb , \42803 );
buf \U$42344 ( \42805 , \42804_nG50eb );
and \U$42345 ( \42806 , \42802 , \42805 );
xor \U$42346 ( \42807 , \14246 , \21250 );
buf g4d41_GF_PartitionCandidate( \42808_nG4d41 , \42807 );
buf \U$42347 ( \42809 , \42808_nG4d41 );
xor \U$42348 ( \42810 , \35274 , \42278 );
buf g4e75_GF_PartitionCandidate( \42811_nG4e75 , \42810 );
buf \U$42349 ( \42812 , \42811_nG4e75 );
and \U$42350 ( \42813 , \42809 , \42812 );
xor \U$42351 ( \42814 , \14508 , \21248 );
buf g4ad8_GF_PartitionCandidate( \42815_nG4ad8 , \42814 );
buf \U$42352 ( \42816 , \42815_nG4ad8 );
xor \U$42353 ( \42817 , \35536 , \42276 );
buf g4c05_GF_PartitionCandidate( \42818_nG4c05 , \42817 );
buf \U$42354 ( \42819 , \42818_nG4c05 );
and \U$42355 ( \42820 , \42816 , \42819 );
xor \U$42356 ( \42821 , \14769 , \21246 );
buf g4879_GF_PartitionCandidate( \42822_nG4879 , \42821 );
buf \U$42357 ( \42823 , \42822_nG4879 );
xor \U$42358 ( \42824 , \35797 , \42274 );
buf g49a3_GF_PartitionCandidate( \42825_nG49a3 , \42824 );
buf \U$42359 ( \42826 , \42825_nG49a3 );
and \U$42360 ( \42827 , \42823 , \42826 );
xor \U$42361 ( \42828 , \14777 , \21244 );
buf g4624_GF_PartitionCandidate( \42829_nG4624 , \42828 );
buf \U$42362 ( \42830 , \42829_nG4624 );
xor \U$42363 ( \42831 , \35805 , \42272 );
buf g4747_GF_PartitionCandidate( \42832_nG4747 , \42831 );
buf \U$42364 ( \42833 , \42832_nG4747 );
and \U$42365 ( \42834 , \42830 , \42833 );
xor \U$42366 ( \42835 , \15023 , \21242 );
buf g43d9_GF_PartitionCandidate( \42836_nG43d9 , \42835 );
buf \U$42367 ( \42837 , \42836_nG43d9 );
xor \U$42368 ( \42838 , \36051 , \42270 );
buf g44f9_GF_PartitionCandidate( \42839_nG44f9 , \42838 );
buf \U$42369 ( \42840 , \42839_nG44f9 );
and \U$42370 ( \42841 , \42837 , \42840 );
xor \U$42371 ( \42842 , \15253 , \21240 );
buf g4198_GF_PartitionCandidate( \42843_nG4198 , \42842 );
buf \U$42372 ( \42844 , \42843_nG4198 );
xor \U$42373 ( \42845 , \36281 , \42268 );
buf g42b1_GF_PartitionCandidate( \42846_nG42b1 , \42845 );
buf \U$42374 ( \42847 , \42846_nG42b1 );
and \U$42375 ( \42848 , \42844 , \42847 );
xor \U$42376 ( \42849 , \15503 , \21238 );
buf g3f61_GF_PartitionCandidate( \42850_nG3f61 , \42849 );
buf \U$42377 ( \42851 , \42850_nG3f61 );
xor \U$42378 ( \42852 , \36531 , \42266 );
buf g4077_GF_PartitionCandidate( \42853_nG4077 , \42852 );
buf \U$42379 ( \42854 , \42853_nG4077 );
and \U$42380 ( \42855 , \42851 , \42854 );
xor \U$42381 ( \42856 , \15728 , \21236 );
buf g3d34_GF_PartitionCandidate( \42857_nG3d34 , \42856 );
buf \U$42382 ( \42858 , \42857_nG3d34 );
xor \U$42383 ( \42859 , \36756 , \42264 );
buf g3e43_GF_PartitionCandidate( \42860_nG3e43 , \42859 );
buf \U$42384 ( \42861 , \42860_nG3e43 );
and \U$42385 ( \42862 , \42858 , \42861 );
xor \U$42386 ( \42863 , \15947 , \21234 );
buf g3b11_GF_PartitionCandidate( \42864_nG3b11 , \42863 );
buf \U$42387 ( \42865 , \42864_nG3b11 );
xor \U$42388 ( \42866 , \36975 , \42262 );
buf g3c1d_GF_PartitionCandidate( \42867_nG3c1d , \42866 );
buf \U$42389 ( \42868 , \42867_nG3c1d );
and \U$42390 ( \42869 , \42865 , \42868 );
xor \U$42391 ( \42870 , \16177 , \21232 );
buf g38f8_GF_PartitionCandidate( \42871_nG38f8 , \42870 );
buf \U$42392 ( \42872 , \42871_nG38f8 );
xor \U$42393 ( \42873 , \37205 , \42260 );
buf g39fd_GF_PartitionCandidate( \42874_nG39fd , \42873 );
buf \U$42394 ( \42875 , \42874_nG39fd );
and \U$42395 ( \42876 , \42872 , \42875 );
xor \U$42396 ( \42877 , \16408 , \21230 );
buf g36e9_GF_PartitionCandidate( \42878_nG36e9 , \42877 );
buf \U$42397 ( \42879 , \42878_nG36e9 );
xor \U$42398 ( \42880 , \37436 , \42258 );
buf g37eb_GF_PartitionCandidate( \42881_nG37eb , \42880 );
buf \U$42399 ( \42882 , \42881_nG37eb );
and \U$42400 ( \42883 , \42879 , \42882 );
xor \U$42401 ( \42884 , \16619 , \21228 );
buf g34e4_GF_PartitionCandidate( \42885_nG34e4 , \42884 );
buf \U$42402 ( \42886 , \42885_nG34e4 );
xor \U$42403 ( \42887 , \37647 , \42256 );
buf g35df_GF_PartitionCandidate( \42888_nG35df , \42887 );
buf \U$42404 ( \42889 , \42888_nG35df );
and \U$42405 ( \42890 , \42886 , \42889 );
xor \U$42406 ( \42891 , \16832 , \21226 );
buf g32e9_GF_PartitionCandidate( \42892_nG32e9 , \42891 );
buf \U$42407 ( \42893 , \42892_nG32e9 );
xor \U$42408 ( \42894 , \37860 , \42254 );
buf g33e1_GF_PartitionCandidate( \42895_nG33e1 , \42894 );
buf \U$42409 ( \42896 , \42895_nG33e1 );
and \U$42410 ( \42897 , \42893 , \42896 );
xor \U$42411 ( \42898 , \17029 , \21224 );
buf g30f8_GF_PartitionCandidate( \42899_nG30f8 , \42898 );
buf \U$42412 ( \42900 , \42899_nG30f8 );
xor \U$42413 ( \42901 , \38057 , \42252 );
buf g31e9_GF_PartitionCandidate( \42902_nG31e9 , \42901 );
buf \U$42414 ( \42903 , \42902_nG31e9 );
and \U$42415 ( \42904 , \42900 , \42903 );
xor \U$42416 ( \42905 , \17225 , \21222 );
buf g2f11_GF_PartitionCandidate( \42906_nG2f11 , \42905 );
buf \U$42417 ( \42907 , \42906_nG2f11 );
xor \U$42418 ( \42908 , \38253 , \42250 );
buf g2fff_GF_PartitionCandidate( \42909_nG2fff , \42908 );
buf \U$42419 ( \42910 , \42909_nG2fff );
and \U$42420 ( \42911 , \42907 , \42910 );
xor \U$42421 ( \42912 , \17433 , \21220 );
buf g2d34_GF_PartitionCandidate( \42913_nG2d34 , \42912 );
buf \U$42422 ( \42914 , \42913_nG2d34 );
xor \U$42423 ( \42915 , \38461 , \42248 );
buf g2e1b_GF_PartitionCandidate( \42916_nG2e1b , \42915 );
buf \U$42424 ( \42917 , \42916_nG2e1b );
and \U$42425 ( \42918 , \42914 , \42917 );
xor \U$42426 ( \42919 , \17618 , \21218 );
buf g2b5e_GF_PartitionCandidate( \42920_nG2b5e , \42919 );
buf \U$42427 ( \42921 , \42920_nG2b5e );
xor \U$42428 ( \42922 , \38646 , \42246 );
buf g2c45_GF_PartitionCandidate( \42923_nG2c45 , \42922 );
buf \U$42429 ( \42924 , \42923_nG2c45 );
and \U$42430 ( \42925 , \42921 , \42924 );
xor \U$42431 ( \42926 , \17805 , \21216 );
buf g2993_GF_PartitionCandidate( \42927_nG2993 , \42926 );
buf \U$42432 ( \42928 , \42927_nG2993 );
xor \U$42433 ( \42929 , \38833 , \42244 );
buf g2a6f_GF_PartitionCandidate( \42930_nG2a6f , \42929 );
buf \U$42434 ( \42931 , \42930_nG2a6f );
and \U$42435 ( \42932 , \42928 , \42931 );
xor \U$42436 ( \42933 , \17995 , \21214 );
buf g27d5_GF_PartitionCandidate( \42934_nG27d5 , \42933 );
buf \U$42437 ( \42935 , \42934_nG27d5 );
xor \U$42438 ( \42936 , \39023 , \42242 );
buf g28af_GF_PartitionCandidate( \42937_nG28af , \42936 );
buf \U$42439 ( \42938 , \42937_nG28af );
and \U$42440 ( \42939 , \42935 , \42938 );
xor \U$42441 ( \42940 , \18171 , \21212 );
buf g2620_GF_PartitionCandidate( \42941_nG2620 , \42940 );
buf \U$42442 ( \42942 , \42941_nG2620 );
xor \U$42443 ( \42943 , \39199 , \42240 );
buf g26f3_GF_PartitionCandidate( \42944_nG26f3 , \42943 );
buf \U$42444 ( \42945 , \42944_nG26f3 );
and \U$42445 ( \42946 , \42942 , \42945 );
xor \U$42446 ( \42947 , \18342 , \21210 );
buf g2475_GF_PartitionCandidate( \42948_nG2475 , \42947 );
buf \U$42447 ( \42949 , \42948_nG2475 );
xor \U$42448 ( \42950 , \39370 , \42238 );
buf g2545_GF_PartitionCandidate( \42951_nG2545 , \42950 );
buf \U$42449 ( \42952 , \42951_nG2545 );
and \U$42450 ( \42953 , \42949 , \42952 );
xor \U$42451 ( \42954 , \18350 , \21208 );
buf g22d4_GF_PartitionCandidate( \42955_nG22d4 , \42954 );
buf \U$42452 ( \42956 , \42955_nG22d4 );
xor \U$42453 ( \42957 , \39378 , \42236 );
buf g239d_GF_PartitionCandidate( \42958_nG239d , \42957 );
buf \U$42454 ( \42959 , \42958_nG239d );
and \U$42455 ( \42960 , \42956 , \42959 );
xor \U$42456 ( \42961 , \18518 , \21206 );
buf g213d_GF_PartitionCandidate( \42962_nG213d , \42961 );
buf \U$42457 ( \42963 , \42962_nG213d );
xor \U$42458 ( \42964 , \39546 , \42234 );
buf g2203_GF_PartitionCandidate( \42965_nG2203 , \42964 );
buf \U$42459 ( \42966 , \42965_nG2203 );
and \U$42460 ( \42967 , \42963 , \42966 );
xor \U$42461 ( \42968 , \18658 , \21204 );
buf g1fb0_GF_PartitionCandidate( \42969_nG1fb0 , \42968 );
buf \U$42462 ( \42970 , \42969_nG1fb0 );
xor \U$42463 ( \42971 , \39686 , \42232 );
buf g206f_GF_PartitionCandidate( \42972_nG206f , \42971 );
buf \U$42464 ( \42973 , \42972_nG206f );
and \U$42465 ( \42974 , \42970 , \42973 );
xor \U$42466 ( \42975 , \18810 , \21202 );
buf g1e2d_GF_PartitionCandidate( \42976_nG1e2d , \42975 );
buf \U$42467 ( \42977 , \42976_nG1e2d );
xor \U$42468 ( \42978 , \39838 , \42230 );
buf g1ee9_GF_PartitionCandidate( \42979_nG1ee9 , \42978 );
buf \U$42469 ( \42980 , \42979_nG1ee9 );
and \U$42470 ( \42981 , \42977 , \42980 );
xor \U$42471 ( \42982 , \18974 , \21200 );
buf g1cb4_GF_PartitionCandidate( \42983_nG1cb4 , \42982 );
buf \U$42472 ( \42984 , \42983_nG1cb4 );
xor \U$42473 ( \42985 , \40002 , \42228 );
buf g1d69_GF_PartitionCandidate( \42986_nG1d69 , \42985 );
buf \U$42474 ( \42987 , \42986_nG1d69 );
and \U$42475 ( \42988 , \42984 , \42987 );
xor \U$42476 ( \42989 , \19113 , \21198 );
buf g1b45_GF_PartitionCandidate( \42990_nG1b45 , \42989 );
buf \U$42477 ( \42991 , \42990_nG1b45 );
xor \U$42478 ( \42992 , \40141 , \42226 );
buf g1bf7_GF_PartitionCandidate( \42993_nG1bf7 , \42992 );
buf \U$42479 ( \42994 , \42993_nG1bf7 );
and \U$42480 ( \42995 , \42991 , \42994 );
xor \U$42481 ( \42996 , \19238 , \21196 );
buf g19e0_GF_PartitionCandidate( \42997_nG19e0 , \42996 );
buf \U$42482 ( \42998 , \42997_nG19e0 );
xor \U$42483 ( \42999 , \40266 , \42224 );
buf g1a8b_GF_PartitionCandidate( \43000_nG1a8b , \42999 );
buf \U$42484 ( \43001 , \43000_nG1a8b );
and \U$42485 ( \43002 , \42998 , \43001 );
xor \U$42486 ( \43003 , \19382 , \21194 );
buf g1885_GF_PartitionCandidate( \43004_nG1885 , \43003 );
buf \U$42487 ( \43005 , \43004_nG1885 );
xor \U$42488 ( \43006 , \40410 , \42222 );
buf g192d_GF_PartitionCandidate( \43007_nG192d , \43006 );
buf \U$42489 ( \43008 , \43007_nG192d );
and \U$42490 ( \43009 , \43005 , \43008 );
xor \U$42491 ( \43010 , \19506 , \21192 );
buf g1734_GF_PartitionCandidate( \43011_nG1734 , \43010 );
buf \U$42492 ( \43012 , \43011_nG1734 );
xor \U$42493 ( \43013 , \40534 , \42220 );
buf g17d5_GF_PartitionCandidate( \43014_nG17d5 , \43013 );
buf \U$42494 ( \43015 , \43014_nG17d5 );
and \U$42495 ( \43016 , \43012 , \43015 );
xor \U$42496 ( \43017 , \19646 , \21190 );
buf g15ed_GF_PartitionCandidate( \43018_nG15ed , \43017 );
buf \U$42497 ( \43019 , \43018_nG15ed );
xor \U$42498 ( \43020 , \40674 , \42218 );
buf g168b_GF_PartitionCandidate( \43021_nG168b , \43020 );
buf \U$42499 ( \43022 , \43021_nG168b );
and \U$42500 ( \43023 , \43019 , \43022 );
xor \U$42501 ( \43024 , \19770 , \21188 );
buf g14b0_GF_PartitionCandidate( \43025_nG14b0 , \43024 );
buf \U$42502 ( \43026 , \43025_nG14b0 );
xor \U$42503 ( \43027 , \40798 , \42216 );
buf g1547_GF_PartitionCandidate( \43028_nG1547 , \43027 );
buf \U$42504 ( \43029 , \43028_nG1547 );
and \U$42505 ( \43030 , \43026 , \43029 );
xor \U$42506 ( \43031 , \19885 , \21186 );
buf g137d_GF_PartitionCandidate( \43032_nG137d , \43031 );
buf \U$42507 ( \43033 , \43032_nG137d );
xor \U$42508 ( \43034 , \40913 , \42214 );
buf g1411_GF_PartitionCandidate( \43035_nG1411 , \43034 );
buf \U$42509 ( \43036 , \43035_nG1411 );
and \U$42510 ( \43037 , \43033 , \43036 );
xor \U$42511 ( \43038 , \19893 , \21184 );
buf g1254_GF_PartitionCandidate( \43039_nG1254 , \43038 );
buf \U$42512 ( \43040 , \43039_nG1254 );
xor \U$42513 ( \43041 , \40921 , \42212 );
buf g12e1_GF_PartitionCandidate( \43042_nG12e1 , \43041 );
buf \U$42514 ( \43043 , \43042_nG12e1 );
and \U$42515 ( \43044 , \43040 , \43043 );
xor \U$42516 ( \43045 , \19989 , \21182 );
buf g1135_GF_PartitionCandidate( \43046_nG1135 , \43045 );
buf \U$42517 ( \43047 , \43046_nG1135 );
xor \U$42518 ( \43048 , \41017 , \42210 );
buf g11bf_GF_PartitionCandidate( \43049_nG11bf , \43048 );
buf \U$42519 ( \43050 , \43049_nG11bf );
and \U$42520 ( \43051 , \43047 , \43050 );
xor \U$42521 ( \43052 , \20104 , \21180 );
buf g1020_GF_PartitionCandidate( \43053_nG1020 , \43052 );
buf \U$42522 ( \43054 , \43053_nG1020 );
xor \U$42523 ( \43055 , \41132 , \42208 );
buf g10a3_GF_PartitionCandidate( \43056_nG10a3 , \43055 );
buf \U$42524 ( \43057 , \43056_nG10a3 );
and \U$42525 ( \43058 , \43054 , \43057 );
xor \U$42526 ( \43059 , \20192 , \21178 );
buf gf15_GF_PartitionCandidate( \43060_nGf15 , \43059 );
buf \U$42527 ( \43061 , \43060_nGf15 );
xor \U$42528 ( \43062 , \41220 , \42206 );
buf gf95_GF_PartitionCandidate( \43063_nGf95 , \43062 );
buf \U$42529 ( \43064 , \43063_nGf95 );
and \U$42530 ( \43065 , \43061 , \43064 );
xor \U$42531 ( \43066 , \20284 , \21176 );
buf ge14_GF_PartitionCandidate( \43067_nGe14 , \43066 );
buf \U$42532 ( \43068 , \43067_nGe14 );
xor \U$42533 ( \43069 , \41312 , \42204 );
buf ge8d_GF_PartitionCandidate( \43070_nGe8d , \43069 );
buf \U$42534 ( \43071 , \43070_nGe8d );
and \U$42535 ( \43072 , \43068 , \43071 );
xor \U$42536 ( \43073 , \20372 , \21174 );
buf gd1d_GF_PartitionCandidate( \43074_nGd1d , \43073 );
buf \U$42537 ( \43075 , \43074_nGd1d );
xor \U$42538 ( \43076 , \41400 , \42202 );
buf gd93_GF_PartitionCandidate( \43077_nGd93 , \43076 );
buf \U$42539 ( \43078 , \43077_nGd93 );
and \U$42540 ( \43079 , \43075 , \43078 );
xor \U$42541 ( \43080 , \20467 , \21172 );
buf gc30_GF_PartitionCandidate( \43081_nGc30 , \43080 );
buf \U$42542 ( \43082 , \43081_nGc30 );
xor \U$42543 ( \43083 , \41495 , \42200 );
buf gc9f_GF_PartitionCandidate( \43084_nGc9f , \43083 );
buf \U$42544 ( \43085 , \43084_nGc9f );
and \U$42545 ( \43086 , \43082 , \43085 );
xor \U$42546 ( \43087 , \20547 , \21170 );
buf gb4d_GF_PartitionCandidate( \43088_nGb4d , \43087 );
buf \U$42547 ( \43089 , \43088_nGb4d );
xor \U$42548 ( \43090 , \41575 , \42198 );
buf gbb9_GF_PartitionCandidate( \43091_nGbb9 , \43090 );
buf \U$42549 ( \43092 , \43091_nGbb9 );
and \U$42550 ( \43093 , \43089 , \43092 );
xor \U$42551 ( \43094 , \20626 , \21168 );
buf ga74_GF_PartitionCandidate( \43095_nGa74 , \43094 );
buf \U$42552 ( \43096 , \43095_nGa74 );
xor \U$42553 ( \43097 , \41654 , \42196 );
buf gad9_GF_PartitionCandidate( \43098_nGad9 , \43097 );
buf \U$42554 ( \43099 , \43098_nGad9 );
and \U$42555 ( \43100 , \43096 , \43099 );
xor \U$42556 ( \43101 , \20634 , \21166 );
buf g9a5_GF_PartitionCandidate( \43102_nG9a5 , \43101 );
buf \U$42557 ( \43103 , \43102_nG9a5 );
xor \U$42558 ( \43104 , \41662 , \42194 );
buf ga07_GF_PartitionCandidate( \43105_nGa07 , \43104 );
buf \U$42559 ( \43106 , \43105_nGa07 );
and \U$42560 ( \43107 , \43103 , \43106 );
xor \U$42561 ( \43108 , \20693 , \21164 );
buf g8e0_GF_PartitionCandidate( \43109_nG8e0 , \43108 );
buf \U$42562 ( \43110 , \43109_nG8e0 );
xor \U$42563 ( \43111 , \41721 , \42192 );
buf g93b_GF_PartitionCandidate( \43112_nG93b , \43111 );
buf \U$42564 ( \43113 , \43112_nG93b );
and \U$42565 ( \43114 , \43110 , \43113 );
xor \U$42566 ( \43115 , \20748 , \21162 );
buf g825_GF_PartitionCandidate( \43116_nG825 , \43115 );
buf \U$42567 ( \43117 , \43116_nG825 );
xor \U$42568 ( \43118 , \41776 , \42190 );
buf g87d_GF_PartitionCandidate( \43119_nG87d , \43118 );
buf \U$42569 ( \43120 , \43119_nG87d );
and \U$42570 ( \43121 , \43117 , \43120 );
xor \U$42571 ( \43122 , \20819 , \21160 );
buf g774_GF_PartitionCandidate( \43123_nG774 , \43122 );
buf \U$42572 ( \43124 , \43123_nG774 );
xor \U$42573 ( \43125 , \41847 , \42188 );
buf g7c5_GF_PartitionCandidate( \43126_nG7c5 , \43125 );
buf \U$42574 ( \43127 , \43126_nG7c5 );
and \U$42575 ( \43128 , \43124 , \43127 );
xor \U$42576 ( \43129 , \20872 , \21158 );
buf g6cd_GF_PartitionCandidate( \43130_nG6cd , \43129 );
buf \U$42577 ( \43131 , \43130_nG6cd );
xor \U$42578 ( \43132 , \41900 , \42186 );
buf g71b_GF_PartitionCandidate( \43133_nG71b , \43132 );
buf \U$42579 ( \43134 , \43133_nG71b );
and \U$42580 ( \43135 , \43131 , \43134 );
xor \U$42581 ( \43136 , \20911 , \21156 );
buf g630_GF_PartitionCandidate( \43137_nG630 , \43136 );
buf \U$42582 ( \43138 , \43137_nG630 );
xor \U$42583 ( \43139 , \41939 , \42184 );
buf g677_GF_PartitionCandidate( \43140_nG677 , \43139 );
buf \U$42584 ( \43141 , \43140_nG677 );
and \U$42585 ( \43142 , \43138 , \43141 );
xor \U$42586 ( \43143 , \20964 , \21154 );
buf g59d_GF_PartitionCandidate( \43144_nG59d , \43143 );
buf \U$42587 ( \43145 , \43144_nG59d );
xor \U$42588 ( \43146 , \41992 , \42182 );
buf g5e1_GF_PartitionCandidate( \43147_nG5e1 , \43146 );
buf \U$42589 ( \43148 , \43147_nG5e1 );
and \U$42590 ( \43149 , \43145 , \43148 );
xor \U$42591 ( \43150 , \20972 , \21152 );
buf g514_GF_PartitionCandidate( \43151_nG514 , \43150 );
buf \U$42592 ( \43152 , \43151_nG514 );
xor \U$42593 ( \43153 , \42000 , \42180 );
buf g551_GF_PartitionCandidate( \43154_nG551 , \43153 );
buf \U$42594 ( \43155 , \43154_nG551 );
and \U$42595 ( \43156 , \43152 , \43155 );
xor \U$42596 ( \43157 , \21006 , \21150 );
buf g495_GF_PartitionCandidate( \43158_nG495 , \43157 );
buf \U$42597 ( \43159 , \43158_nG495 );
xor \U$42598 ( \43160 , \42034 , \42178 );
buf g4cf_GF_PartitionCandidate( \43161_nG4cf , \43160 );
buf \U$42599 ( \43162 , \43161_nG4cf );
and \U$42600 ( \43163 , \43159 , \43162 );
xor \U$42601 ( \43164 , \21040 , \21148 );
buf g420_GF_PartitionCandidate( \43165_nG420 , \43164 );
buf \U$42602 ( \43166 , \43165_nG420 );
xor \U$42603 ( \43167 , \42068 , \42176 );
buf g453_GF_PartitionCandidate( \43168_nG453 , \43167 );
buf \U$42604 ( \43169 , \43168_nG453 );
and \U$42605 ( \43170 , \43166 , \43169 );
xor \U$42606 ( \43171 , \21048 , \21146 );
buf g3b5_GF_PartitionCandidate( \43172_nG3b5 , \43171 );
buf \U$42607 ( \43173 , \43172_nG3b5 );
xor \U$42608 ( \43174 , \42076 , \42174 );
buf g3e5_GF_PartitionCandidate( \43175_nG3e5 , \43174 );
buf \U$42609 ( \43176 , \43175_nG3e5 );
and \U$42610 ( \43177 , \43173 , \43176 );
xor \U$42611 ( \43178 , \21074 , \21144 );
buf g354_GF_PartitionCandidate( \43179_nG354 , \43178 );
buf \U$42612 ( \43180 , \43179_nG354 );
xor \U$42613 ( \43181 , \42102 , \42172 );
buf g37d_GF_PartitionCandidate( \43182_nG37d , \43181 );
buf \U$42614 ( \43183 , \43182_nG37d );
and \U$42615 ( \43184 , \43180 , \43183 );
xor \U$42616 ( \43185 , \21093 , \21142 );
buf g2fd_GF_PartitionCandidate( \43186_nG2fd , \43185 );
buf \U$42617 ( \43187 , \43186_nG2fd );
xor \U$42618 ( \43188 , \42121 , \42170 );
buf g323_GF_PartitionCandidate( \43189_nG323 , \43188 );
buf \U$42619 ( \43190 , \43189_nG323 );
and \U$42620 ( \43191 , \43187 , \43190 );
xor \U$42621 ( \43192 , \21101 , \21140 );
buf g2b0_GF_PartitionCandidate( \43193_nG2b0 , \43192 );
buf \U$42622 ( \43194 , \43193_nG2b0 );
xor \U$42623 ( \43195 , \42129 , \42168 );
buf g2cf_GF_PartitionCandidate( \43196_nG2cf , \43195 );
buf \U$42624 ( \43197 , \43196_nG2cf );
and \U$42625 ( \43198 , \43194 , \43197 );
xor \U$42626 ( \43199 , \21113 , \21138 );
buf g26d_GF_PartitionCandidate( \43200_nG26d , \43199 );
buf \U$42627 ( \43201 , \43200_nG26d );
xor \U$42628 ( \43202 , \42141 , \42166 );
buf g289_GF_PartitionCandidate( \43203_nG289 , \43202 );
buf \U$42629 ( \43204 , \43203_nG289 );
and \U$42630 ( \43205 , \43201 , \43204 );
xor \U$42631 ( \43206 , \21121 , \21136 );
buf g234_GF_PartitionCandidate( \43207_nG234 , \43206 );
buf \U$42632 ( \43208 , \43207_nG234 );
xor \U$42633 ( \43209 , \42149 , \42164 );
buf g249_GF_PartitionCandidate( \43210_nG249 , \43209 );
buf \U$42634 ( \43211 , \43210_nG249 );
and \U$42635 ( \43212 , \43208 , \43211 );
xor \U$42636 ( \43213 , \21126 , \21134 );
buf g204_GF_PartitionCandidate( \43214_nG204 , \43213 );
buf \U$42637 ( \43215 , \43214_nG204 );
xor \U$42638 ( \43216 , \42154 , \42162 );
buf g217_GF_PartitionCandidate( \43217_nG217 , \43216 );
buf \U$42639 ( \43218 , \43217_nG217 );
and \U$42640 ( \43219 , \43215 , \43218 );
xor \U$42641 ( \43220 , \21130 , \21133 );
buf g1e0_GF_PartitionCandidate( \43221_nG1e0 , \43220 );
buf \U$42642 ( \43222 , \43221_nG1e0 );
xor \U$42643 ( \43223 , \42158 , \42161 );
buf g1ec_GF_PartitionCandidate( \43224_nG1ec , \43223 );
buf \U$42644 ( \43225 , \43224_nG1ec );
and \U$42645 ( \43226 , \43222 , \43225 );
xor \U$42646 ( \43227 , \21132 , \9556 );
buf g189_GF_PartitionCandidate( \43228_nG189 , \43227 );
buf \U$42647 ( \43229 , \43228_nG189 );
xor \U$42648 ( \43230 , \42160 , \30584 );
buf g191_GF_PartitionCandidate( \43231_nG191 , \43230 );
buf \U$42649 ( \43232 , \43231_nG191 );
and \U$42650 ( \43233 , \43229 , \43232 );
and \U$42651 ( \43234 , \43225 , \43233 );
and \U$42652 ( \43235 , \43222 , \43233 );
or \U$42653 ( \43236 , \43226 , \43234 , \43235 );
and \U$42654 ( \43237 , \43218 , \43236 );
and \U$42655 ( \43238 , \43215 , \43236 );
or \U$42656 ( \43239 , \43219 , \43237 , \43238 );
and \U$42657 ( \43240 , \43211 , \43239 );
and \U$42658 ( \43241 , \43208 , \43239 );
or \U$42659 ( \43242 , \43212 , \43240 , \43241 );
and \U$42660 ( \43243 , \43204 , \43242 );
and \U$42661 ( \43244 , \43201 , \43242 );
or \U$42662 ( \43245 , \43205 , \43243 , \43244 );
and \U$42663 ( \43246 , \43197 , \43245 );
and \U$42664 ( \43247 , \43194 , \43245 );
or \U$42665 ( \43248 , \43198 , \43246 , \43247 );
and \U$42666 ( \43249 , \43190 , \43248 );
and \U$42667 ( \43250 , \43187 , \43248 );
or \U$42668 ( \43251 , \43191 , \43249 , \43250 );
and \U$42669 ( \43252 , \43183 , \43251 );
and \U$42670 ( \43253 , \43180 , \43251 );
or \U$42671 ( \43254 , \43184 , \43252 , \43253 );
and \U$42672 ( \43255 , \43176 , \43254 );
and \U$42673 ( \43256 , \43173 , \43254 );
or \U$42674 ( \43257 , \43177 , \43255 , \43256 );
and \U$42675 ( \43258 , \43169 , \43257 );
and \U$42676 ( \43259 , \43166 , \43257 );
or \U$42677 ( \43260 , \43170 , \43258 , \43259 );
and \U$42678 ( \43261 , \43162 , \43260 );
and \U$42679 ( \43262 , \43159 , \43260 );
or \U$42680 ( \43263 , \43163 , \43261 , \43262 );
and \U$42681 ( \43264 , \43155 , \43263 );
and \U$42682 ( \43265 , \43152 , \43263 );
or \U$42683 ( \43266 , \43156 , \43264 , \43265 );
and \U$42684 ( \43267 , \43148 , \43266 );
and \U$42685 ( \43268 , \43145 , \43266 );
or \U$42686 ( \43269 , \43149 , \43267 , \43268 );
and \U$42687 ( \43270 , \43141 , \43269 );
and \U$42688 ( \43271 , \43138 , \43269 );
or \U$42689 ( \43272 , \43142 , \43270 , \43271 );
and \U$42690 ( \43273 , \43134 , \43272 );
and \U$42691 ( \43274 , \43131 , \43272 );
or \U$42692 ( \43275 , \43135 , \43273 , \43274 );
and \U$42693 ( \43276 , \43127 , \43275 );
and \U$42694 ( \43277 , \43124 , \43275 );
or \U$42695 ( \43278 , \43128 , \43276 , \43277 );
and \U$42696 ( \43279 , \43120 , \43278 );
and \U$42697 ( \43280 , \43117 , \43278 );
or \U$42698 ( \43281 , \43121 , \43279 , \43280 );
and \U$42699 ( \43282 , \43113 , \43281 );
and \U$42700 ( \43283 , \43110 , \43281 );
or \U$42701 ( \43284 , \43114 , \43282 , \43283 );
and \U$42702 ( \43285 , \43106 , \43284 );
and \U$42703 ( \43286 , \43103 , \43284 );
or \U$42704 ( \43287 , \43107 , \43285 , \43286 );
and \U$42705 ( \43288 , \43099 , \43287 );
and \U$42706 ( \43289 , \43096 , \43287 );
or \U$42707 ( \43290 , \43100 , \43288 , \43289 );
and \U$42708 ( \43291 , \43092 , \43290 );
and \U$42709 ( \43292 , \43089 , \43290 );
or \U$42710 ( \43293 , \43093 , \43291 , \43292 );
and \U$42711 ( \43294 , \43085 , \43293 );
and \U$42712 ( \43295 , \43082 , \43293 );
or \U$42713 ( \43296 , \43086 , \43294 , \43295 );
and \U$42714 ( \43297 , \43078 , \43296 );
and \U$42715 ( \43298 , \43075 , \43296 );
or \U$42716 ( \43299 , \43079 , \43297 , \43298 );
and \U$42717 ( \43300 , \43071 , \43299 );
and \U$42718 ( \43301 , \43068 , \43299 );
or \U$42719 ( \43302 , \43072 , \43300 , \43301 );
and \U$42720 ( \43303 , \43064 , \43302 );
and \U$42721 ( \43304 , \43061 , \43302 );
or \U$42722 ( \43305 , \43065 , \43303 , \43304 );
and \U$42723 ( \43306 , \43057 , \43305 );
and \U$42724 ( \43307 , \43054 , \43305 );
or \U$42725 ( \43308 , \43058 , \43306 , \43307 );
and \U$42726 ( \43309 , \43050 , \43308 );
and \U$42727 ( \43310 , \43047 , \43308 );
or \U$42728 ( \43311 , \43051 , \43309 , \43310 );
and \U$42729 ( \43312 , \43043 , \43311 );
and \U$42730 ( \43313 , \43040 , \43311 );
or \U$42731 ( \43314 , \43044 , \43312 , \43313 );
and \U$42732 ( \43315 , \43036 , \43314 );
and \U$42733 ( \43316 , \43033 , \43314 );
or \U$42734 ( \43317 , \43037 , \43315 , \43316 );
and \U$42735 ( \43318 , \43029 , \43317 );
and \U$42736 ( \43319 , \43026 , \43317 );
or \U$42737 ( \43320 , \43030 , \43318 , \43319 );
and \U$42738 ( \43321 , \43022 , \43320 );
and \U$42739 ( \43322 , \43019 , \43320 );
or \U$42740 ( \43323 , \43023 , \43321 , \43322 );
and \U$42741 ( \43324 , \43015 , \43323 );
and \U$42742 ( \43325 , \43012 , \43323 );
or \U$42743 ( \43326 , \43016 , \43324 , \43325 );
and \U$42744 ( \43327 , \43008 , \43326 );
and \U$42745 ( \43328 , \43005 , \43326 );
or \U$42746 ( \43329 , \43009 , \43327 , \43328 );
and \U$42747 ( \43330 , \43001 , \43329 );
and \U$42748 ( \43331 , \42998 , \43329 );
or \U$42749 ( \43332 , \43002 , \43330 , \43331 );
and \U$42750 ( \43333 , \42994 , \43332 );
and \U$42751 ( \43334 , \42991 , \43332 );
or \U$42752 ( \43335 , \42995 , \43333 , \43334 );
and \U$42753 ( \43336 , \42987 , \43335 );
and \U$42754 ( \43337 , \42984 , \43335 );
or \U$42755 ( \43338 , \42988 , \43336 , \43337 );
and \U$42756 ( \43339 , \42980 , \43338 );
and \U$42757 ( \43340 , \42977 , \43338 );
or \U$42758 ( \43341 , \42981 , \43339 , \43340 );
and \U$42759 ( \43342 , \42973 , \43341 );
and \U$42760 ( \43343 , \42970 , \43341 );
or \U$42761 ( \43344 , \42974 , \43342 , \43343 );
and \U$42762 ( \43345 , \42966 , \43344 );
and \U$42763 ( \43346 , \42963 , \43344 );
or \U$42764 ( \43347 , \42967 , \43345 , \43346 );
and \U$42765 ( \43348 , \42959 , \43347 );
and \U$42766 ( \43349 , \42956 , \43347 );
or \U$42767 ( \43350 , \42960 , \43348 , \43349 );
and \U$42768 ( \43351 , \42952 , \43350 );
and \U$42769 ( \43352 , \42949 , \43350 );
or \U$42770 ( \43353 , \42953 , \43351 , \43352 );
and \U$42771 ( \43354 , \42945 , \43353 );
and \U$42772 ( \43355 , \42942 , \43353 );
or \U$42773 ( \43356 , \42946 , \43354 , \43355 );
and \U$42774 ( \43357 , \42938 , \43356 );
and \U$42775 ( \43358 , \42935 , \43356 );
or \U$42776 ( \43359 , \42939 , \43357 , \43358 );
and \U$42777 ( \43360 , \42931 , \43359 );
and \U$42778 ( \43361 , \42928 , \43359 );
or \U$42779 ( \43362 , \42932 , \43360 , \43361 );
and \U$42780 ( \43363 , \42924 , \43362 );
and \U$42781 ( \43364 , \42921 , \43362 );
or \U$42782 ( \43365 , \42925 , \43363 , \43364 );
and \U$42783 ( \43366 , \42917 , \43365 );
and \U$42784 ( \43367 , \42914 , \43365 );
or \U$42785 ( \43368 , \42918 , \43366 , \43367 );
and \U$42786 ( \43369 , \42910 , \43368 );
and \U$42787 ( \43370 , \42907 , \43368 );
or \U$42788 ( \43371 , \42911 , \43369 , \43370 );
and \U$42789 ( \43372 , \42903 , \43371 );
and \U$42790 ( \43373 , \42900 , \43371 );
or \U$42791 ( \43374 , \42904 , \43372 , \43373 );
and \U$42792 ( \43375 , \42896 , \43374 );
and \U$42793 ( \43376 , \42893 , \43374 );
or \U$42794 ( \43377 , \42897 , \43375 , \43376 );
and \U$42795 ( \43378 , \42889 , \43377 );
and \U$42796 ( \43379 , \42886 , \43377 );
or \U$42797 ( \43380 , \42890 , \43378 , \43379 );
and \U$42798 ( \43381 , \42882 , \43380 );
and \U$42799 ( \43382 , \42879 , \43380 );
or \U$42800 ( \43383 , \42883 , \43381 , \43382 );
and \U$42801 ( \43384 , \42875 , \43383 );
and \U$42802 ( \43385 , \42872 , \43383 );
or \U$42803 ( \43386 , \42876 , \43384 , \43385 );
and \U$42804 ( \43387 , \42868 , \43386 );
and \U$42805 ( \43388 , \42865 , \43386 );
or \U$42806 ( \43389 , \42869 , \43387 , \43388 );
and \U$42807 ( \43390 , \42861 , \43389 );
and \U$42808 ( \43391 , \42858 , \43389 );
or \U$42809 ( \43392 , \42862 , \43390 , \43391 );
and \U$42810 ( \43393 , \42854 , \43392 );
and \U$42811 ( \43394 , \42851 , \43392 );
or \U$42812 ( \43395 , \42855 , \43393 , \43394 );
and \U$42813 ( \43396 , \42847 , \43395 );
and \U$42814 ( \43397 , \42844 , \43395 );
or \U$42815 ( \43398 , \42848 , \43396 , \43397 );
and \U$42816 ( \43399 , \42840 , \43398 );
and \U$42817 ( \43400 , \42837 , \43398 );
or \U$42818 ( \43401 , \42841 , \43399 , \43400 );
and \U$42819 ( \43402 , \42833 , \43401 );
and \U$42820 ( \43403 , \42830 , \43401 );
or \U$42821 ( \43404 , \42834 , \43402 , \43403 );
and \U$42822 ( \43405 , \42826 , \43404 );
and \U$42823 ( \43406 , \42823 , \43404 );
or \U$42824 ( \43407 , \42827 , \43405 , \43406 );
and \U$42825 ( \43408 , \42819 , \43407 );
and \U$42826 ( \43409 , \42816 , \43407 );
or \U$42827 ( \43410 , \42820 , \43408 , \43409 );
and \U$42828 ( \43411 , \42812 , \43410 );
and \U$42829 ( \43412 , \42809 , \43410 );
or \U$42830 ( \43413 , \42813 , \43411 , \43412 );
and \U$42831 ( \43414 , \42805 , \43413 );
and \U$42832 ( \43415 , \42802 , \43413 );
or \U$42833 ( \43416 , \42806 , \43414 , \43415 );
and \U$42834 ( \43417 , \42798 , \43416 );
and \U$42835 ( \43418 , \42795 , \43416 );
or \U$42836 ( \43419 , \42799 , \43417 , \43418 );
and \U$42837 ( \43420 , \42791 , \43419 );
and \U$42838 ( \43421 , \42788 , \43419 );
or \U$42839 ( \43422 , \42792 , \43420 , \43421 );
and \U$42840 ( \43423 , \42784 , \43422 );
and \U$42841 ( \43424 , \42781 , \43422 );
or \U$42842 ( \43425 , \42785 , \43423 , \43424 );
and \U$42843 ( \43426 , \42777 , \43425 );
and \U$42844 ( \43427 , \42774 , \43425 );
or \U$42845 ( \43428 , \42778 , \43426 , \43427 );
and \U$42846 ( \43429 , \42770 , \43428 );
and \U$42847 ( \43430 , \42767 , \43428 );
or \U$42848 ( \43431 , \42771 , \43429 , \43430 );
and \U$42849 ( \43432 , \42763 , \43431 );
and \U$42850 ( \43433 , \42760 , \43431 );
or \U$42851 ( \43434 , \42764 , \43432 , \43433 );
and \U$42852 ( \43435 , \42756 , \43434 );
and \U$42853 ( \43436 , \42753 , \43434 );
or \U$42854 ( \43437 , \42757 , \43435 , \43436 );
and \U$42855 ( \43438 , \42749 , \43437 );
and \U$42856 ( \43439 , \42746 , \43437 );
or \U$42857 ( \43440 , \42750 , \43438 , \43439 );
and \U$42858 ( \43441 , \42742 , \43440 );
and \U$42859 ( \43442 , \42739 , \43440 );
or \U$42860 ( \43443 , \42743 , \43441 , \43442 );
and \U$42861 ( \43444 , \42735 , \43443 );
and \U$42862 ( \43445 , \42732 , \43443 );
or \U$42863 ( \43446 , \42736 , \43444 , \43445 );
and \U$42864 ( \43447 , \42728 , \43446 );
and \U$42865 ( \43448 , \42725 , \43446 );
or \U$42866 ( \43449 , \42729 , \43447 , \43448 );
and \U$42867 ( \43450 , \42721 , \43449 );
and \U$42868 ( \43451 , \42718 , \43449 );
or \U$42869 ( \43452 , \42722 , \43450 , \43451 );
and \U$42870 ( \43453 , \42714 , \43452 );
and \U$42871 ( \43454 , \42711 , \43452 );
or \U$42872 ( \43455 , \42715 , \43453 , \43454 );
and \U$42873 ( \43456 , \42707 , \43455 );
and \U$42874 ( \43457 , \42704 , \43455 );
or \U$42875 ( \43458 , \42708 , \43456 , \43457 );
and \U$42876 ( \43459 , \42700 , \43458 );
and \U$42877 ( \43460 , \42697 , \43458 );
or \U$42878 ( \43461 , \42701 , \43459 , \43460 );
and \U$42879 ( \43462 , \42693 , \43461 );
and \U$42880 ( \43463 , \42690 , \43461 );
or \U$42881 ( \43464 , \42694 , \43462 , \43463 );
and \U$42882 ( \43465 , \42686 , \43464 );
and \U$42883 ( \43466 , \42683 , \43464 );
or \U$42884 ( \43467 , \42687 , \43465 , \43466 );
and \U$42885 ( \43468 , \42679 , \43467 );
and \U$42886 ( \43469 , \42676 , \43467 );
or \U$42887 ( \43470 , \42680 , \43468 , \43469 );
and \U$42888 ( \43471 , \42672 , \43470 );
and \U$42889 ( \43472 , \42669 , \43470 );
or \U$42890 ( \43473 , \42673 , \43471 , \43472 );
and \U$42891 ( \43474 , \42665 , \43473 );
and \U$42892 ( \43475 , \42662 , \43473 );
or \U$42893 ( \43476 , \42666 , \43474 , \43475 );
and \U$42894 ( \43477 , \42658 , \43476 );
and \U$42895 ( \43478 , \42655 , \43476 );
or \U$42896 ( \43479 , \42659 , \43477 , \43478 );
and \U$42897 ( \43480 , \42651 , \43479 );
and \U$42898 ( \43481 , \42648 , \43479 );
or \U$42899 ( \43482 , \42652 , \43480 , \43481 );
and \U$42900 ( \43483 , \42644 , \43482 );
and \U$42901 ( \43484 , \42641 , \43482 );
or \U$42902 ( \43485 , \42645 , \43483 , \43484 );
and \U$42903 ( \43486 , \42637 , \43485 );
and \U$42904 ( \43487 , \42634 , \43485 );
or \U$42905 ( \43488 , \42638 , \43486 , \43487 );
and \U$42906 ( \43489 , \42630 , \43488 );
and \U$42907 ( \43490 , \42627 , \43488 );
or \U$42908 ( \43491 , \42631 , \43489 , \43490 );
and \U$42909 ( \43492 , \42623 , \43491 );
and \U$42910 ( \43493 , \42620 , \43491 );
or \U$42911 ( \43494 , \42624 , \43492 , \43493 );
and \U$42912 ( \43495 , \42616 , \43494 );
and \U$42913 ( \43496 , \42613 , \43494 );
or \U$42914 ( \43497 , \42617 , \43495 , \43496 );
and \U$42915 ( \43498 , \42609 , \43497 );
and \U$42916 ( \43499 , \42606 , \43497 );
or \U$42917 ( \43500 , \42610 , \43498 , \43499 );
and \U$42918 ( \43501 , \42602 , \43500 );
and \U$42919 ( \43502 , \42599 , \43500 );
or \U$42920 ( \43503 , \42603 , \43501 , \43502 );
and \U$42921 ( \43504 , \42595 , \43503 );
and \U$42922 ( \43505 , \42592 , \43503 );
or \U$42923 ( \43506 , \42596 , \43504 , \43505 );
and \U$42924 ( \43507 , \42588 , \43506 );
and \U$42925 ( \43508 , \42585 , \43506 );
or \U$42926 ( \43509 , \42589 , \43507 , \43508 );
and \U$42927 ( \43510 , \42581 , \43509 );
and \U$42928 ( \43511 , \42578 , \43509 );
or \U$42929 ( \43512 , \42582 , \43510 , \43511 );
and \U$42930 ( \43513 , \42574 , \43512 );
and \U$42931 ( \43514 , \42571 , \43512 );
or \U$42932 ( \43515 , \42575 , \43513 , \43514 );
and \U$42933 ( \43516 , \42567 , \43515 );
and \U$42934 ( \43517 , \42564 , \43515 );
or \U$42935 ( \43518 , \42568 , \43516 , \43517 );
and \U$42936 ( \43519 , \42560 , \43518 );
and \U$42937 ( \43520 , \42557 , \43518 );
or \U$42938 ( \43521 , \42561 , \43519 , \43520 );
and \U$42939 ( \43522 , \42553 , \43521 );
and \U$42940 ( \43523 , \42550 , \43521 );
or \U$42941 ( \43524 , \42554 , \43522 , \43523 );
and \U$42942 ( \43525 , \42546 , \43524 );
and \U$42943 ( \43526 , \42543 , \43524 );
or \U$42944 ( \43527 , \42547 , \43525 , \43526 );
and \U$42945 ( \43528 , \42539 , \43527 );
and \U$42946 ( \43529 , \42536 , \43527 );
or \U$42947 ( \43530 , \42540 , \43528 , \43529 );
and \U$42948 ( \43531 , \42532 , \43530 );
and \U$42949 ( \43532 , \42529 , \43530 );
or \U$42950 ( \43533 , \42533 , \43531 , \43532 );
and \U$42951 ( \43534 , \42525 , \43533 );
and \U$42952 ( \43535 , \42522 , \43533 );
or \U$42953 ( \43536 , \42526 , \43534 , \43535 );
and \U$42954 ( \43537 , \42518 , \43536 );
and \U$42955 ( \43538 , \42515 , \43536 );
or \U$42956 ( \43539 , \42519 , \43537 , \43538 );
and \U$42957 ( \43540 , \42511 , \43539 );
and \U$42958 ( \43541 , \42508 , \43539 );
or \U$42959 ( \43542 , \42512 , \43540 , \43541 );
and \U$42960 ( \43543 , \42504 , \43542 );
and \U$42961 ( \43544 , \42501 , \43542 );
or \U$42962 ( \43545 , \42505 , \43543 , \43544 );
and \U$42963 ( \43546 , \42497 , \43545 );
and \U$42964 ( \43547 , \42494 , \43545 );
or \U$42965 ( \43548 , \42498 , \43546 , \43547 );
and \U$42966 ( \43549 , \42490 , \43548 );
and \U$42967 ( \43550 , \42487 , \43548 );
or \U$42968 ( \43551 , \42491 , \43549 , \43550 );
and \U$42969 ( \43552 , \42483 , \43551 );
and \U$42970 ( \43553 , \42480 , \43551 );
or \U$42971 ( \43554 , \42484 , \43552 , \43553 );
and \U$42972 ( \43555 , \42476 , \43554 );
and \U$42973 ( \43556 , \42473 , \43554 );
or \U$42974 ( \43557 , \42477 , \43555 , \43556 );
and \U$42975 ( \43558 , \42469 , \43557 );
and \U$42976 ( \43559 , \42466 , \43557 );
or \U$42977 ( \43560 , \42470 , \43558 , \43559 );
and \U$42978 ( \43561 , \42462 , \43560 );
and \U$42979 ( \43562 , \42459 , \43560 );
or \U$42980 ( \43563 , \42463 , \43561 , \43562 );
and \U$42981 ( \43564 , \42455 , \43563 );
and \U$42982 ( \43565 , \42452 , \43563 );
or \U$42983 ( \43566 , \42456 , \43564 , \43565 );
and \U$42984 ( \43567 , \42448 , \43566 );
and \U$42985 ( \43568 , \42445 , \43566 );
or \U$42986 ( \43569 , \42449 , \43567 , \43568 );
and \U$42987 ( \43570 , \42441 , \43569 );
and \U$42988 ( \43571 , \42438 , \43569 );
or \U$42989 ( \43572 , \42442 , \43570 , \43571 );
and \U$42990 ( \43573 , \42434 , \43572 );
and \U$42991 ( \43574 , \42431 , \43572 );
or \U$42992 ( \43575 , \42435 , \43573 , \43574 );
and \U$42993 ( \43576 , \42427 , \43575 );
and \U$42994 ( \43577 , \42424 , \43575 );
or \U$42995 ( \43578 , \42428 , \43576 , \43577 );
and \U$42996 ( \43579 , \42420 , \43578 );
and \U$42997 ( \43580 , \42417 , \43578 );
or \U$42998 ( \43581 , \42421 , \43579 , \43580 );
and \U$42999 ( \43582 , \42413 , \43581 );
and \U$43000 ( \43583 , \42410 , \43581 );
or \U$43001 ( \43584 , \42414 , \43582 , \43583 );
and \U$43002 ( \43585 , \42406 , \43584 );
and \U$43003 ( \43586 , \42403 , \43584 );
or \U$43004 ( \43587 , \42407 , \43585 , \43586 );
xor \U$43005 ( \43588 , \42400 , \43587 );
buf gac8b_GF_PartitionCandidate( \43589_nGac8b , \43588 );
xor \U$43006 ( \43590 , RIbb333f0_193, RIbb33468_194);
xor \U$43007 ( \43591 , RIbb334e0_195, RIbb33558_196);
xor \U$43008 ( \43592 , \43590 , \43591 );
xor \U$43009 ( \43593 , RIbb335d0_197, RIbb33648_198);
xor \U$43010 ( \43594 , RIbb336c0_199, RIbb33738_200);
xor \U$43011 ( \43595 , \43593 , \43594 );
xor \U$43012 ( \43596 , \43592 , \43595 );
xor \U$43013 ( \43597 , RIbb337b0_201, RIbb33828_202);
xor \U$43014 ( \43598 , RIbb338a0_203, RIbb33918_204);
xor \U$43015 ( \43599 , \43597 , \43598 );
xor \U$43016 ( \43600 , RIbb33990_205, RIbb33a08_206);
xor \U$43017 ( \43601 , RIbb33a80_207, RIbb33af8_208);
xor \U$43018 ( \43602 , \43600 , \43601 );
xor \U$43019 ( \43603 , \43599 , \43602 );
xor \U$43020 ( \43604 , \43596 , \43603 );
xor \U$43021 ( \43605 , RIbb33b70_209, RIbb33be8_210);
xor \U$43022 ( \43606 , RIbb33c60_211, RIbb33cd8_212);
xor \U$43023 ( \43607 , \43605 , \43606 );
xor \U$43024 ( \43608 , RIbb33d50_213, RIbb33dc8_214);
xor \U$43025 ( \43609 , RIbb33e40_215, RIbb33eb8_216);
xor \U$43026 ( \43610 , \43608 , \43609 );
xor \U$43027 ( \43611 , \43607 , \43610 );
xor \U$43028 ( \43612 , RIbb33f30_217, RIbb33fa8_218);
xor \U$43029 ( \43613 , RIbb34020_219, RIbb34098_220);
xor \U$43030 ( \43614 , \43612 , \43613 );
xor \U$43031 ( \43615 , RIbb34110_221, RIbb34188_222);
xor \U$43032 ( \43616 , RIbb34200_223, RIbb34278_224);
xor \U$43033 ( \43617 , \43615 , \43616 );
xor \U$43034 ( \43618 , \43614 , \43617 );
xor \U$43035 ( \43619 , \43611 , \43618 );
xor \U$43036 ( \43620 , \43604 , \43619 );
xor \U$43037 ( \43621 , RIbb342f0_225, RIbb34368_226);
xor \U$43038 ( \43622 , RIbb343e0_227, RIbb34458_228);
xor \U$43039 ( \43623 , \43621 , \43622 );
xor \U$43040 ( \43624 , RIbb344d0_229, RIbb34548_230);
xor \U$43041 ( \43625 , RIbb345c0_231, RIbb34638_232);
xor \U$43042 ( \43626 , \43624 , \43625 );
xor \U$43043 ( \43627 , \43623 , \43626 );
xor \U$43044 ( \43628 , RIbb346b0_233, RIbb34728_234);
xor \U$43045 ( \43629 , RIbb347a0_235, RIbb34818_236);
xor \U$43046 ( \43630 , \43628 , \43629 );
xor \U$43047 ( \43631 , RIbb34890_237, RIbb34908_238);
xor \U$43048 ( \43632 , RIbb34980_239, RIbb349f8_240);
xor \U$43049 ( \43633 , \43631 , \43632 );
xor \U$43050 ( \43634 , \43630 , \43633 );
xor \U$43051 ( \43635 , \43627 , \43634 );
xor \U$43052 ( \43636 , RIbb34a70_241, RIbb34ae8_242);
xor \U$43053 ( \43637 , RIbb34b60_243, RIbb34bd8_244);
xor \U$43054 ( \43638 , \43636 , \43637 );
xor \U$43055 ( \43639 , RIbb34c50_245, RIbb34cc8_246);
xor \U$43056 ( \43640 , RIbb34d40_247, RIbb34db8_248);
xor \U$43057 ( \43641 , \43639 , \43640 );
xor \U$43058 ( \43642 , \43638 , \43641 );
xor \U$43059 ( \43643 , RIbb34e30_249, RIbb34ea8_250);
xor \U$43060 ( \43644 , RIbb34f20_251, RIbb34f98_252);
xor \U$43061 ( \43645 , \43643 , \43644 );
xor \U$43062 ( \43646 , RIbb35010_253, RIbb35088_254);
xor \U$43063 ( \43647 , RIbb35100_255, RIbb35178_256);
xor \U$43064 ( \43648 , \43646 , \43647 );
xor \U$43065 ( \43649 , \43645 , \43648 );
xor \U$43066 ( \43650 , \43642 , \43649 );
xor \U$43067 ( \43651 , \43635 , \43650 );
xor \U$43068 ( \43652 , \43620 , \43651 );
not \U$43069 ( \43653 , \43652 );
_DC gac8c ( \43654_nGac8c , \43589_nGac8b , \43653 );
buf \U$43070 ( \43655 , \43654_nGac8c );
xor \U$43071 ( \43656 , \42403 , \42406 );
xor \U$43072 ( \43657 , \43656 , \43584 );
buf gac15_GF_PartitionCandidate( \43658_nGac15 , \43657 );
_DC gac16 ( \43659_nGac16 , \43658_nGac15 , \43653 );
buf \U$43073 ( \43660 , \43659_nGac16 );
xor \U$43074 ( \43661 , \42417 , \42420 );
xor \U$43075 ( \43662 , \43661 , \43578 );
buf gaaff_GF_PartitionCandidate( \43663_nGaaff , \43662 );
_DC gab00 ( \43664_nGab00 , \43663_nGaaff , \43653 );
buf \U$43076 ( \43665 , \43664_nGab00 );
xor \U$43077 ( \43666 , \42438 , \42441 );
xor \U$43078 ( \43667 , \43666 , \43569 );
buf ga91b_GF_PartitionCandidate( \43668_nGa91b , \43667 );
_DC ga91c ( \43669_nGa91c , \43668_nGa91b , \43653 );
buf \U$43079 ( \43670 , \43669_nGa91c );
xor \U$43080 ( \43671 , \42452 , \42455 );
xor \U$43081 ( \43672 , \43671 , \43563 );
buf ga7a7_GF_PartitionCandidate( \43673_nGa7a7 , \43672 );
_DC ga7a8 ( \43674_nGa7a8 , \43673_nGa7a7 , \43653 );
buf \U$43082 ( \43675 , \43674_nGa7a8 );
xor \U$43083 ( \43676 , \42508 , \42511 );
xor \U$43084 ( \43677 , \43676 , \43539 );
buf ga043_GF_PartitionCandidate( \43678_nGa043 , \43677 );
_DC ga044 ( \43679_nGa044 , \43678_nGa043 , \43653 );
buf \U$43085 ( \43680 , \43679_nGa044 );
xor \U$43086 ( \43681 , \42529 , \42532 );
xor \U$43087 ( \43682 , \43681 , \43530 );
buf g9cd7_GF_PartitionCandidate( \43683_nG9cd7 , \43682 );
_DC g9cd8 ( \43684_nG9cd8 , \43683_nG9cd7 , \43653 );
buf \U$43088 ( \43685 , \43684_nG9cd8 );
xor \U$43089 ( \43686 , \42536 , \42539 );
xor \U$43090 ( \43687 , \43686 , \43527 );
buf g9b99_GF_PartitionCandidate( \43688_nG9b99 , \43687 );
_DC g9b9a ( \43689_nG9b9a , \43688_nG9b99 , \43653 );
buf \U$43091 ( \43690 , \43689_nG9b9a );
xor \U$43092 ( \43691 , \42550 , \42553 );
xor \U$43093 ( \43692 , \43691 , \43521 );
buf g9903_GF_PartitionCandidate( \43693_nG9903 , \43692 );
_DC g9904 ( \43694_nG9904 , \43693_nG9903 , \43653 );
buf \U$43094 ( \43695 , \43694_nG9904 );
xor \U$43095 ( \43696 , \42571 , \42574 );
xor \U$43096 ( \43697 , \43696 , \43512 );
buf g94f3_GF_PartitionCandidate( \43698_nG94f3 , \43697 );
_DC g94f4 ( \43699_nG94f4 , \43698_nG94f3 , \43653 );
buf \U$43097 ( \43700 , \43699_nG94f4 );
xor \U$43098 ( \43701 , \42578 , \42581 );
xor \U$43099 ( \43702 , \43701 , \43509 );
buf g9381_GF_PartitionCandidate( \43703_nG9381 , \43702 );
_DC g9382 ( \43704_nG9382 , \43703_nG9381 , \43653 );
buf \U$43100 ( \43705 , \43704_nG9382 );
xor \U$43101 ( \43706 , \42585 , \42588 );
xor \U$43102 ( \43707 , \43706 , \43506 );
buf g9205_GF_PartitionCandidate( \43708_nG9205 , \43707 );
_DC g9206 ( \43709_nG9206 , \43708_nG9205 , \43653 );
buf \U$43103 ( \43710 , \43709_nG9206 );
xor \U$43104 ( \43711 , \42592 , \42595 );
xor \U$43105 ( \43712 , \43711 , \43503 );
buf g907b_GF_PartitionCandidate( \43713_nG907b , \43712 );
_DC g907c ( \43714_nG907c , \43713_nG907b , \43653 );
buf \U$43106 ( \43715 , \43714_nG907c );
xor \U$43107 ( \43716 , \42606 , \42609 );
xor \U$43108 ( \43717 , \43716 , \43497 );
buf g8d4f_GF_PartitionCandidate( \43718_nG8d4f , \43717 );
_DC g8d50 ( \43719_nG8d50 , \43718_nG8d4f , \43653 );
buf \U$43109 ( \43720 , \43719_nG8d50 );
xor \U$43110 ( \43721 , \42613 , \42616 );
xor \U$43111 ( \43722 , \43721 , \43494 );
buf g8bad_GF_PartitionCandidate( \43723_nG8bad , \43722 );
_DC g8bae ( \43724_nG8bae , \43723_nG8bad , \43653 );
buf \U$43112 ( \43725 , \43724_nG8bae );
xor \U$43113 ( \43726 , \42620 , \42623 );
xor \U$43114 ( \43727 , \43726 , \43491 );
buf g89fb_GF_PartitionCandidate( \43728_nG89fb , \43727 );
_DC g89fc ( \43729_nG89fc , \43728_nG89fb , \43653 );
buf \U$43115 ( \43730 , \43729_nG89fc );
xor \U$43116 ( \43731 , \42634 , \42637 );
xor \U$43117 ( \43732 , \43731 , \43485 );
buf g8677_GF_PartitionCandidate( \43733_nG8677 , \43732 );
_DC g8678 ( \43734_nG8678 , \43733_nG8677 , \43653 );
buf \U$43118 ( \43735 , \43734_nG8678 );
xor \U$43119 ( \43736 , \42641 , \42644 );
xor \U$43120 ( \43737 , \43736 , \43482 );
buf g84a7_GF_PartitionCandidate( \43738_nG84a7 , \43737 );
_DC g84a8 ( \43739_nG84a8 , \43738_nG84a7 , \43653 );
buf \U$43121 ( \43740 , \43739_nG84a8 );
xor \U$43122 ( \43741 , \42655 , \42658 );
xor \U$43123 ( \43742 , \43741 , \43476 );
buf g80e7_GF_PartitionCandidate( \43743_nG80e7 , \43742 );
_DC g80e8 ( \43744_nG80e8 , \43743_nG80e7 , \43653 );
buf \U$43124 ( \43745 , \43744_nG80e8 );
xor \U$43125 ( \43746 , \42662 , \42665 );
xor \U$43126 ( \43747 , \43746 , \43473 );
buf g7ef5_GF_PartitionCandidate( \43748_nG7ef5 , \43747 );
_DC g7ef6 ( \43749_nG7ef6 , \43748_nG7ef5 , \43653 );
buf \U$43127 ( \43750 , \43749_nG7ef6 );
xor \U$43128 ( \43751 , \42669 , \42672 );
xor \U$43129 ( \43752 , \43751 , \43470 );
buf g7cf9_GF_PartitionCandidate( \43753_nG7cf9 , \43752 );
_DC g7cfa ( \43754_nG7cfa , \43753_nG7cf9 , \43653 );
buf \U$43130 ( \43755 , \43754_nG7cfa );
xor \U$43131 ( \43756 , \42676 , \42679 );
xor \U$43132 ( \43757 , \43756 , \43467 );
buf g7af7_GF_PartitionCandidate( \43758_nG7af7 , \43757 );
_DC g7af8 ( \43759_nG7af8 , \43758_nG7af7 , \43653 );
buf \U$43133 ( \43760 , \43759_nG7af8 );
xor \U$43134 ( \43761 , \42704 , \42707 );
xor \U$43135 ( \43762 , \43761 , \43455 );
buf g72a1_GF_PartitionCandidate( \43763_nG72a1 , \43762 );
_DC g72a2 ( \43764_nG72a2 , \43763_nG72a1 , \43653 );
buf \U$43136 ( \43765 , \43764_nG72a2 );
xor \U$43137 ( \43766 , \42711 , \42714 );
xor \U$43138 ( \43767 , \43766 , \43452 );
buf g7077_GF_PartitionCandidate( \43768_nG7077 , \43767 );
_DC g7078 ( \43769_nG7078 , \43768_nG7077 , \43653 );
buf \U$43139 ( \43770 , \43769_nG7078 );
xor \U$43140 ( \43771 , \42718 , \42721 );
xor \U$43141 ( \43772 , \43771 , \43449 );
buf g6e3d_GF_PartitionCandidate( \43773_nG6e3d , \43772 );
_DC g6e3e ( \43774_nG6e3e , \43773_nG6e3d , \43653 );
buf \U$43142 ( \43775 , \43774_nG6e3e );
xor \U$43143 ( \43776 , \42725 , \42728 );
xor \U$43144 ( \43777 , \43776 , \43446 );
buf g6bff_GF_PartitionCandidate( \43778_nG6bff , \43777 );
_DC g6c00 ( \43779_nG6c00 , \43778_nG6bff , \43653 );
buf \U$43145 ( \43780 , \43779_nG6c00 );
xor \U$43146 ( \43781 , \42732 , \42735 );
xor \U$43147 ( \43782 , \43781 , \43443 );
buf g69b1_GF_PartitionCandidate( \43783_nG69b1 , \43782 );
_DC g69b2 ( \43784_nG69b2 , \43783_nG69b1 , \43653 );
buf \U$43148 ( \43785 , \43784_nG69b2 );
xor \U$43149 ( \43786 , \42746 , \42749 );
xor \U$43150 ( \43787 , \43786 , \43437 );
buf g64f3_GF_PartitionCandidate( \43788_nG64f3 , \43787 );
_DC g64f4 ( \43789_nG64f4 , \43788_nG64f3 , \43653 );
buf \U$43151 ( \43790 , \43789_nG64f4 );
xor \U$43152 ( \43791 , \42760 , \42763 );
xor \U$43153 ( \43792 , \43791 , \43431 );
buf g600d_GF_PartitionCandidate( \43793_nG600d , \43792 );
_DC g600e ( \43794_nG600e , \43793_nG600d , \43653 );
buf \U$43154 ( \43795 , \43794_nG600e );
xor \U$43155 ( \43796 , \42767 , \42770 );
xor \U$43156 ( \43797 , \43796 , \43428 );
buf g5d8d_GF_PartitionCandidate( \43798_nG5d8d , \43797 );
_DC g5d8e ( \43799_nG5d8e , \43798_nG5d8d , \43653 );
buf \U$43157 ( \43800 , \43799_nG5d8e );
xor \U$43158 ( \43801 , \42774 , \42777 );
xor \U$43159 ( \43802 , \43801 , \43425 );
buf g5b0b_GF_PartitionCandidate( \43803_nG5b0b , \43802 );
_DC g5b0c ( \43804_nG5b0c , \43803_nG5b0b , \43653 );
buf \U$43160 ( \43805 , \43804_nG5b0c );
xor \U$43161 ( \43806 , \42781 , \42784 );
xor \U$43162 ( \43807 , \43806 , \43422 );
buf g5887_GF_PartitionCandidate( \43808_nG5887 , \43807 );
_DC g5888 ( \43809_nG5888 , \43808_nG5887 , \43653 );
buf \U$43163 ( \43810 , \43809_nG5888 );
xor \U$43164 ( \43811 , \42788 , \42791 );
xor \U$43165 ( \43812 , \43811 , \43419 );
buf g5601_GF_PartitionCandidate( \43813_nG5601 , \43812 );
_DC g5602 ( \43814_nG5602 , \43813_nG5601 , \43653 );
buf \U$43166 ( \43815 , \43814_nG5602 );
xor \U$43167 ( \43816 , \42802 , \42805 );
xor \U$43168 ( \43817 , \43816 , \43413 );
buf g50f3_GF_PartitionCandidate( \43818_nG50f3 , \43817 );
_DC g50f4 ( \43819_nG50f4 , \43818_nG50f3 , \43653 );
buf \U$43169 ( \43820 , \43819_nG50f4 );
xor \U$43170 ( \43821 , \42809 , \42812 );
xor \U$43171 ( \43822 , \43821 , \43410 );
buf g4e7d_GF_PartitionCandidate( \43823_nG4e7d , \43822 );
_DC g4e7e ( \43824_nG4e7e , \43823_nG4e7d , \43653 );
buf \U$43172 ( \43825 , \43824_nG4e7e );
xor \U$43173 ( \43826 , \42816 , \42819 );
xor \U$43174 ( \43827 , \43826 , \43407 );
buf g4c0d_GF_PartitionCandidate( \43828_nG4c0d , \43827 );
_DC g4c0e ( \43829_nG4c0e , \43828_nG4c0d , \43653 );
buf \U$43175 ( \43830 , \43829_nG4c0e );
xor \U$43176 ( \43831 , \42823 , \42826 );
xor \U$43177 ( \43832 , \43831 , \43404 );
buf g49ab_GF_PartitionCandidate( \43833_nG49ab , \43832 );
_DC g49ac ( \43834_nG49ac , \43833_nG49ab , \43653 );
buf \U$43178 ( \43835 , \43834_nG49ac );
xor \U$43179 ( \43836 , \42830 , \42833 );
xor \U$43180 ( \43837 , \43836 , \43401 );
buf g474f_GF_PartitionCandidate( \43838_nG474f , \43837 );
_DC g4750 ( \43839_nG4750 , \43838_nG474f , \43653 );
buf \U$43181 ( \43840 , \43839_nG4750 );
xor \U$43182 ( \43841 , \42837 , \42840 );
xor \U$43183 ( \43842 , \43841 , \43398 );
buf g4501_GF_PartitionCandidate( \43843_nG4501 , \43842 );
_DC g4502 ( \43844_nG4502 , \43843_nG4501 , \43653 );
buf \U$43184 ( \43845 , \43844_nG4502 );
xor \U$43185 ( \43846 , \42844 , \42847 );
xor \U$43186 ( \43847 , \43846 , \43395 );
buf g42b9_GF_PartitionCandidate( \43848_nG42b9 , \43847 );
_DC g42ba ( \43849_nG42ba , \43848_nG42b9 , \43653 );
buf \U$43187 ( \43850 , \43849_nG42ba );
xor \U$43188 ( \43851 , \42851 , \42854 );
xor \U$43189 ( \43852 , \43851 , \43392 );
buf g407f_GF_PartitionCandidate( \43853_nG407f , \43852 );
_DC g4080 ( \43854_nG4080 , \43853_nG407f , \43653 );
buf \U$43190 ( \43855 , \43854_nG4080 );
xor \U$43191 ( \43856 , \42858 , \42861 );
xor \U$43192 ( \43857 , \43856 , \43389 );
buf g3e4b_GF_PartitionCandidate( \43858_nG3e4b , \43857 );
_DC g3e4c ( \43859_nG3e4c , \43858_nG3e4b , \43653 );
buf \U$43193 ( \43860 , \43859_nG3e4c );
xor \U$43194 ( \43861 , \42865 , \42868 );
xor \U$43195 ( \43862 , \43861 , \43386 );
buf g3c25_GF_PartitionCandidate( \43863_nG3c25 , \43862 );
_DC g3c26 ( \43864_nG3c26 , \43863_nG3c25 , \43653 );
buf \U$43196 ( \43865 , \43864_nG3c26 );
xor \U$43197 ( \43866 , \42872 , \42875 );
xor \U$43198 ( \43867 , \43866 , \43383 );
buf g3a05_GF_PartitionCandidate( \43868_nG3a05 , \43867 );
_DC g3a06 ( \43869_nG3a06 , \43868_nG3a05 , \43653 );
buf \U$43199 ( \43870 , \43869_nG3a06 );
xor \U$43200 ( \43871 , \42879 , \42882 );
xor \U$43201 ( \43872 , \43871 , \43380 );
buf g37f3_GF_PartitionCandidate( \43873_nG37f3 , \43872 );
_DC g37f4 ( \43874_nG37f4 , \43873_nG37f3 , \43653 );
buf \U$43202 ( \43875 , \43874_nG37f4 );
xor \U$43203 ( \43876 , \42886 , \42889 );
xor \U$43204 ( \43877 , \43876 , \43377 );
buf g35e7_GF_PartitionCandidate( \43878_nG35e7 , \43877 );
_DC g35e8 ( \43879_nG35e8 , \43878_nG35e7 , \43653 );
buf \U$43205 ( \43880 , \43879_nG35e8 );
xor \U$43206 ( \43881 , \42893 , \42896 );
xor \U$43207 ( \43882 , \43881 , \43374 );
buf g33e9_GF_PartitionCandidate( \43883_nG33e9 , \43882 );
_DC g33ea ( \43884_nG33ea , \43883_nG33e9 , \43653 );
buf \U$43208 ( \43885 , \43884_nG33ea );
xor \U$43209 ( \43886 , \42900 , \42903 );
xor \U$43210 ( \43887 , \43886 , \43371 );
buf g31f1_GF_PartitionCandidate( \43888_nG31f1 , \43887 );
_DC g31f2 ( \43889_nG31f2 , \43888_nG31f1 , \43653 );
buf \U$43211 ( \43890 , \43889_nG31f2 );
xor \U$43212 ( \43891 , \42907 , \42910 );
xor \U$43213 ( \43892 , \43891 , \43368 );
buf g3007_GF_PartitionCandidate( \43893_nG3007 , \43892 );
_DC g3008 ( \43894_nG3008 , \43893_nG3007 , \43653 );
buf \U$43214 ( \43895 , \43894_nG3008 );
xor \U$43215 ( \43896 , \42914 , \42917 );
xor \U$43216 ( \43897 , \43896 , \43365 );
buf g2e23_GF_PartitionCandidate( \43898_nG2e23 , \43897 );
_DC g2e24 ( \43899_nG2e24 , \43898_nG2e23 , \43653 );
buf \U$43217 ( \43900 , \43899_nG2e24 );
xor \U$43218 ( \43901 , \42921 , \42924 );
xor \U$43219 ( \43902 , \43901 , \43362 );
buf g2c4d_GF_PartitionCandidate( \43903_nG2c4d , \43902 );
_DC g2c4e ( \43904_nG2c4e , \43903_nG2c4d , \43653 );
buf \U$43220 ( \43905 , \43904_nG2c4e );
xor \U$43221 ( \43906 , \42928 , \42931 );
xor \U$43222 ( \43907 , \43906 , \43359 );
buf g2a77_GF_PartitionCandidate( \43908_nG2a77 , \43907 );
_DC g2a78 ( \43909_nG2a78 , \43908_nG2a77 , \43653 );
buf \U$43223 ( \43910 , \43909_nG2a78 );
xor \U$43224 ( \43911 , \42935 , \42938 );
xor \U$43225 ( \43912 , \43911 , \43356 );
buf g28b7_GF_PartitionCandidate( \43913_nG28b7 , \43912 );
_DC g28b8 ( \43914_nG28b8 , \43913_nG28b7 , \43653 );
buf \U$43226 ( \43915 , \43914_nG28b8 );
xor \U$43227 ( \43916 , \42942 , \42945 );
xor \U$43228 ( \43917 , \43916 , \43353 );
buf g26fb_GF_PartitionCandidate( \43918_nG26fb , \43917 );
_DC g26fc ( \43919_nG26fc , \43918_nG26fb , \43653 );
buf \U$43229 ( \43920 , \43919_nG26fc );
xor \U$43230 ( \43921 , \42949 , \42952 );
xor \U$43231 ( \43922 , \43921 , \43350 );
buf g254d_GF_PartitionCandidate( \43923_nG254d , \43922 );
_DC g254e ( \43924_nG254e , \43923_nG254d , \43653 );
buf \U$43232 ( \43925 , \43924_nG254e );
xor \U$43233 ( \43926 , \42956 , \42959 );
xor \U$43234 ( \43927 , \43926 , \43347 );
buf g23a5_GF_PartitionCandidate( \43928_nG23a5 , \43927 );
_DC g23a6 ( \43929_nG23a6 , \43928_nG23a5 , \43653 );
buf \U$43235 ( \43930 , \43929_nG23a6 );
xor \U$43236 ( \43931 , \42963 , \42966 );
xor \U$43237 ( \43932 , \43931 , \43344 );
buf g220b_GF_PartitionCandidate( \43933_nG220b , \43932 );
_DC g220c ( \43934_nG220c , \43933_nG220b , \43653 );
buf \U$43238 ( \43935 , \43934_nG220c );
xor \U$43239 ( \43936 , \42970 , \42973 );
xor \U$43240 ( \43937 , \43936 , \43341 );
buf g2077_GF_PartitionCandidate( \43938_nG2077 , \43937 );
_DC g2078 ( \43939_nG2078 , \43938_nG2077 , \43653 );
buf \U$43241 ( \43940 , \43939_nG2078 );
xor \U$43242 ( \43941 , \42977 , \42980 );
xor \U$43243 ( \43942 , \43941 , \43338 );
buf g1ef1_GF_PartitionCandidate( \43943_nG1ef1 , \43942 );
_DC g1ef2 ( \43944_nG1ef2 , \43943_nG1ef1 , \43653 );
buf \U$43244 ( \43945 , \43944_nG1ef2 );
xor \U$43245 ( \43946 , \42984 , \42987 );
xor \U$43246 ( \43947 , \43946 , \43335 );
buf g1d71_GF_PartitionCandidate( \43948_nG1d71 , \43947 );
_DC g1d72 ( \43949_nG1d72 , \43948_nG1d71 , \43653 );
buf \U$43247 ( \43950 , \43949_nG1d72 );
xor \U$43248 ( \43951 , \42991 , \42994 );
xor \U$43249 ( \43952 , \43951 , \43332 );
buf g1bff_GF_PartitionCandidate( \43953_nG1bff , \43952 );
_DC g1c00 ( \43954_nG1c00 , \43953_nG1bff , \43653 );
buf \U$43250 ( \43955 , \43954_nG1c00 );
xor \U$43251 ( \43956 , \42998 , \43001 );
xor \U$43252 ( \43957 , \43956 , \43329 );
buf g1a93_GF_PartitionCandidate( \43958_nG1a93 , \43957 );
_DC g1a94 ( \43959_nG1a94 , \43958_nG1a93 , \43653 );
buf \U$43253 ( \43960 , \43959_nG1a94 );
xor \U$43254 ( \43961 , \43005 , \43008 );
xor \U$43255 ( \43962 , \43961 , \43326 );
buf g1935_GF_PartitionCandidate( \43963_nG1935 , \43962 );
_DC g1936 ( \43964_nG1936 , \43963_nG1935 , \43653 );
buf \U$43256 ( \43965 , \43964_nG1936 );
xor \U$43257 ( \43966 , \43012 , \43015 );
xor \U$43258 ( \43967 , \43966 , \43323 );
buf g17dd_GF_PartitionCandidate( \43968_nG17dd , \43967 );
_DC g17de ( \43969_nG17de , \43968_nG17dd , \43653 );
buf \U$43259 ( \43970 , \43969_nG17de );
xor \U$43260 ( \43971 , \43019 , \43022 );
xor \U$43261 ( \43972 , \43971 , \43320 );
buf g1693_GF_PartitionCandidate( \43973_nG1693 , \43972 );
_DC g1694 ( \43974_nG1694 , \43973_nG1693 , \43653 );
buf \U$43262 ( \43975 , \43974_nG1694 );
xor \U$43263 ( \43976 , \43026 , \43029 );
xor \U$43264 ( \43977 , \43976 , \43317 );
buf g154f_GF_PartitionCandidate( \43978_nG154f , \43977 );
_DC g1550 ( \43979_nG1550 , \43978_nG154f , \43653 );
buf \U$43265 ( \43980 , \43979_nG1550 );
xor \U$43266 ( \43981 , \43033 , \43036 );
xor \U$43267 ( \43982 , \43981 , \43314 );
buf g1419_GF_PartitionCandidate( \43983_nG1419 , \43982 );
_DC g141a ( \43984_nG141a , \43983_nG1419 , \43653 );
buf \U$43268 ( \43985 , \43984_nG141a );
xor \U$43269 ( \43986 , \43040 , \43043 );
xor \U$43270 ( \43987 , \43986 , \43311 );
buf g12e9_GF_PartitionCandidate( \43988_nG12e9 , \43987 );
_DC g12ea ( \43989_nG12ea , \43988_nG12e9 , \43653 );
buf \U$43271 ( \43990 , \43989_nG12ea );
xor \U$43272 ( \43991 , \43047 , \43050 );
xor \U$43273 ( \43992 , \43991 , \43308 );
buf g11c7_GF_PartitionCandidate( \43993_nG11c7 , \43992 );
_DC g11c8 ( \43994_nG11c8 , \43993_nG11c7 , \43653 );
buf \U$43274 ( \43995 , \43994_nG11c8 );
xor \U$43275 ( \43996 , \43054 , \43057 );
xor \U$43276 ( \43997 , \43996 , \43305 );
buf g10ab_GF_PartitionCandidate( \43998_nG10ab , \43997 );
_DC g10ac ( \43999_nG10ac , \43998_nG10ab , \43653 );
buf \U$43277 ( \44000 , \43999_nG10ac );
xor \U$43278 ( \44001 , \43061 , \43064 );
xor \U$43279 ( \44002 , \44001 , \43302 );
buf gf9d_GF_PartitionCandidate( \44003_nGf9d , \44002 );
_DC gf9e ( \44004_nGf9e , \44003_nGf9d , \43653 );
buf \U$43280 ( \44005 , \44004_nGf9e );
xor \U$43281 ( \44006 , \43068 , \43071 );
xor \U$43282 ( \44007 , \44006 , \43299 );
buf ge95_GF_PartitionCandidate( \44008_nGe95 , \44007 );
_DC ge96 ( \44009_nGe96 , \44008_nGe95 , \43653 );
buf \U$43283 ( \44010 , \44009_nGe96 );
xor \U$43284 ( \44011 , \43075 , \43078 );
xor \U$43285 ( \44012 , \44011 , \43296 );
buf gd9b_GF_PartitionCandidate( \44013_nGd9b , \44012 );
_DC gd9c ( \44014_nGd9c , \44013_nGd9b , \43653 );
buf \U$43286 ( \44015 , \44014_nGd9c );
xor \U$43287 ( \44016 , \43082 , \43085 );
xor \U$43288 ( \44017 , \44016 , \43293 );
buf gca7_GF_PartitionCandidate( \44018_nGca7 , \44017 );
_DC gca8 ( \44019_nGca8 , \44018_nGca7 , \43653 );
buf \U$43289 ( \44020 , \44019_nGca8 );
xor \U$43290 ( \44021 , \43089 , \43092 );
xor \U$43291 ( \44022 , \44021 , \43290 );
buf gbc1_GF_PartitionCandidate( \44023_nGbc1 , \44022 );
_DC gbc2 ( \44024_nGbc2 , \44023_nGbc1 , \43653 );
buf \U$43292 ( \44025 , \44024_nGbc2 );
xor \U$43293 ( \44026 , \43096 , \43099 );
xor \U$43294 ( \44027 , \44026 , \43287 );
buf gae1_GF_PartitionCandidate( \44028_nGae1 , \44027 );
_DC gae2 ( \44029_nGae2 , \44028_nGae1 , \43653 );
buf \U$43295 ( \44030 , \44029_nGae2 );
xor \U$43296 ( \44031 , \43103 , \43106 );
xor \U$43297 ( \44032 , \44031 , \43284 );
buf ga0f_GF_PartitionCandidate( \44033_nGa0f , \44032 );
_DC ga10 ( \44034_nGa10 , \44033_nGa0f , \43653 );
buf \U$43298 ( \44035 , \44034_nGa10 );
xor \U$43299 ( \44036 , \43110 , \43113 );
xor \U$43300 ( \44037 , \44036 , \43281 );
buf g943_GF_PartitionCandidate( \44038_nG943 , \44037 );
_DC g944 ( \44039_nG944 , \44038_nG943 , \43653 );
buf \U$43301 ( \44040 , \44039_nG944 );
xor \U$43302 ( \44041 , \43117 , \43120 );
xor \U$43303 ( \44042 , \44041 , \43278 );
buf g885_GF_PartitionCandidate( \44043_nG885 , \44042 );
_DC g886 ( \44044_nG886 , \44043_nG885 , \43653 );
buf \U$43304 ( \44045 , \44044_nG886 );
xor \U$43305 ( \44046 , \43124 , \43127 );
xor \U$43306 ( \44047 , \44046 , \43275 );
buf g7cd_GF_PartitionCandidate( \44048_nG7cd , \44047 );
_DC g7ce ( \44049_nG7ce , \44048_nG7cd , \43653 );
buf \U$43307 ( \44050 , \44049_nG7ce );
xor \U$43308 ( \44051 , \43131 , \43134 );
xor \U$43309 ( \44052 , \44051 , \43272 );
buf g723_GF_PartitionCandidate( \44053_nG723 , \44052 );
_DC g724 ( \44054_nG724 , \44053_nG723 , \43653 );
buf \U$43310 ( \44055 , \44054_nG724 );
xor \U$43311 ( \44056 , \43138 , \43141 );
xor \U$43312 ( \44057 , \44056 , \43269 );
buf g67f_GF_PartitionCandidate( \44058_nG67f , \44057 );
_DC g680 ( \44059_nG680 , \44058_nG67f , \43653 );
buf \U$43313 ( \44060 , \44059_nG680 );
xor \U$43314 ( \44061 , \43145 , \43148 );
xor \U$43315 ( \44062 , \44061 , \43266 );
buf g5e9_GF_PartitionCandidate( \44063_nG5e9 , \44062 );
_DC g5ea ( \44064_nG5ea , \44063_nG5e9 , \43653 );
buf \U$43316 ( \44065 , \44064_nG5ea );
xor \U$43317 ( \44066 , \43152 , \43155 );
xor \U$43318 ( \44067 , \44066 , \43263 );
buf g559_GF_PartitionCandidate( \44068_nG559 , \44067 );
_DC g55a ( \44069_nG55a , \44068_nG559 , \43653 );
buf \U$43319 ( \44070 , \44069_nG55a );
xor \U$43320 ( \44071 , \43159 , \43162 );
xor \U$43321 ( \44072 , \44071 , \43260 );
buf g4d7_GF_PartitionCandidate( \44073_nG4d7 , \44072 );
_DC g4d8 ( \44074_nG4d8 , \44073_nG4d7 , \43653 );
buf \U$43322 ( \44075 , \44074_nG4d8 );
endmodule

