//
// Conformal-LEC Version 20.10-d130 (26-Jun-2020)
//
module top(RIb559478_125,RIb55f760_53,RIb55f6e8_54,RIb55f670_55,RIb5594f0_124,RIb559388_127,RIb55f850_51,RIb55f7d8_52,RIb559400_126,
        RIb559310_128,RIb55f8c8_50,RIb55f940_49,RIb55da50_115,RIb55f2b0_63,RIb55f238_64,RIb55dac8_114,RIb55d960_117,RIb55f3a0_61,RIb55f328_62,
        RIb55d9d8_116,RIb55d870_119,RIb55f490_59,RIb55f418_60,RIb55d8e8_118,RIb55d780_121,RIb55f580_57,RIb55f508_58,RIb55d7f8_120,RIb55d690_123,
        RIb55f5f8_56,RIb55d708_122,RIb55db40_113,RIb55dbb8_112,RIb55fa30_47,RIb55f9b8_48,RIb55dc30_111,RIb55dca8_110,RIb55fb20_45,RIb55faa8_46,
        RIb55dd20_109,RIb55dd98_108,RIb55fc10_43,RIb55fb98_44,RIb55de10_107,RIb55fc88_42,RIb55fd00_41,RIb55de88_106,RIb55df00_105,RIb55df78_104,
        RIb55fdf0_39,RIb55fd78_40,RIb55dff0_103,RIb55e068_102,RIb55fee0_37,RIb55fe68_38,RIb55e0e0_101,RIb55e158_100,RIb55ffd0_35,RIb55ff58_36,
        RIb55e1d0_99,RIb55e248_98,RIb5600c0_33,RIb560048_34,RIb55e2c0_97,RIb55e338_96,RIb5601b0_31,RIb560138_32,RIb55e3b0_95,RIb55e428_94,
        RIb5602a0_29,RIb560228_30,RIb55e4a0_93,RIb560318_28,RIb560390_27,RIb55e518_92,RIb55e590_91,RIb55e608_90,RIb560480_25,RIb560408_26,
        RIb55e680_89,RIb55e6f8_88,RIb560570_23,RIb5604f8_24,RIb55e770_87,RIb55e7e8_86,RIb560660_21,RIb5605e8_22,RIb55e860_85,RIb55e8d8_84,
        RIb560750_19,RIb5606d8_20,RIb55e950_83,RIb55e9c8_82,RIb560840_17,RIb5607c8_18,RIb55ea40_81,RIb5608b8_16,RIb560930_15,RIb55eab8_80,
        RIb55eb30_79,RIb5609a8_14,RIb560a20_13,RIb55eba8_78,RIb55ec20_77,RIb560a98_12,RIb560b10_11,RIb55ec98_76,RIb55ed10_75,RIb55ed88_74,
        RIb560c00_9,RIb560b88_10,RIb55ee00_73,RIb560c78_8,RIb560cf0_7,RIb55ee78_72,RIb55eef0_71,RIb55ef68_70,RIb560de0_5,RIb560d68_6,
        RIb55efe0_69,RIb55f058_68,RIb560ed0_3,RIb560e58_4,RIb55f0d0_67,RIb560f48_2,RIb560fc0_1,RIb55f148_66,RIb55f1c0_65,R_81_7e072f0);
input RIb559478_125,RIb55f760_53,RIb55f6e8_54,RIb55f670_55,RIb5594f0_124,RIb559388_127,RIb55f850_51,RIb55f7d8_52,RIb559400_126,
        RIb559310_128,RIb55f8c8_50,RIb55f940_49,RIb55da50_115,RIb55f2b0_63,RIb55f238_64,RIb55dac8_114,RIb55d960_117,RIb55f3a0_61,RIb55f328_62,
        RIb55d9d8_116,RIb55d870_119,RIb55f490_59,RIb55f418_60,RIb55d8e8_118,RIb55d780_121,RIb55f580_57,RIb55f508_58,RIb55d7f8_120,RIb55d690_123,
        RIb55f5f8_56,RIb55d708_122,RIb55db40_113,RIb55dbb8_112,RIb55fa30_47,RIb55f9b8_48,RIb55dc30_111,RIb55dca8_110,RIb55fb20_45,RIb55faa8_46,
        RIb55dd20_109,RIb55dd98_108,RIb55fc10_43,RIb55fb98_44,RIb55de10_107,RIb55fc88_42,RIb55fd00_41,RIb55de88_106,RIb55df00_105,RIb55df78_104,
        RIb55fdf0_39,RIb55fd78_40,RIb55dff0_103,RIb55e068_102,RIb55fee0_37,RIb55fe68_38,RIb55e0e0_101,RIb55e158_100,RIb55ffd0_35,RIb55ff58_36,
        RIb55e1d0_99,RIb55e248_98,RIb5600c0_33,RIb560048_34,RIb55e2c0_97,RIb55e338_96,RIb5601b0_31,RIb560138_32,RIb55e3b0_95,RIb55e428_94,
        RIb5602a0_29,RIb560228_30,RIb55e4a0_93,RIb560318_28,RIb560390_27,RIb55e518_92,RIb55e590_91,RIb55e608_90,RIb560480_25,RIb560408_26,
        RIb55e680_89,RIb55e6f8_88,RIb560570_23,RIb5604f8_24,RIb55e770_87,RIb55e7e8_86,RIb560660_21,RIb5605e8_22,RIb55e860_85,RIb55e8d8_84,
        RIb560750_19,RIb5606d8_20,RIb55e950_83,RIb55e9c8_82,RIb560840_17,RIb5607c8_18,RIb55ea40_81,RIb5608b8_16,RIb560930_15,RIb55eab8_80,
        RIb55eb30_79,RIb5609a8_14,RIb560a20_13,RIb55eba8_78,RIb55ec20_77,RIb560a98_12,RIb560b10_11,RIb55ec98_76,RIb55ed10_75,RIb55ed88_74,
        RIb560c00_9,RIb560b88_10,RIb55ee00_73,RIb560c78_8,RIb560cf0_7,RIb55ee78_72,RIb55eef0_71,RIb55ef68_70,RIb560de0_5,RIb560d68_6,
        RIb55efe0_69,RIb55f058_68,RIb560ed0_3,RIb560e58_4,RIb55f0d0_67,RIb560f48_2,RIb560fc0_1,RIb55f148_66,RIb55f1c0_65;
output R_81_7e072f0;

wire \130 , \131_N$1 , \132_ZERO , \133_ONE , \134 , \135 , \136 , \137 , \138 ,
         \139 , \140 , \141 , \142 , \143 , \144 , \145 , \146 , \147 , \148 ,
         \149 , \150 , \151 , \152 , \153 , \154 , \155 , \156 , \157 , \158 ,
         \159 , \160 , \161 , \162 , \163 , \164 , \165 , \166 , \167 , \168 ,
         \169 , \170 , \171 , \172 , \173 , \174 , \175 , \176 , \177 , \178 ,
         \179 , \180 , \181 , \182 , \183 , \184 , \185 , \186 , \187 , \188 ,
         \189 , \190 , \191 , \192 , \193 , \194 , \195 , \196 , \197 , \198 ,
         \199 , \200 , \201 , \202 , \203 , \204 , \205 , \206 , \207 , \208 ,
         \209 , \210 , \211 , \212 , \213 , \214 , \215 , \216 , \217 , \218 ,
         \219 , \220 , \221 , \222 , \223 , \224 , \225 , \226 , \227 , \228 ,
         \229 , \230 , \231 , \232 , \233 , \234 , \235 , \236 , \237 , \238 ,
         \239 , \240 , \241 , \242 , \243 , \244 , \245 , \246 , \247 , \248 ,
         \249 , \250 , \251 , \252 , \253 , \254 , \255 , \256 , \257 , \258 ,
         \259 , \260 , \261 , \262 , \263 , \264 , \265 , \266 , \267 , \268 ,
         \269 , \270 , \271 , \272 , \273 , \274 , \275 , \276 , \277 , \278 ,
         \279 , \280 , \281 , \282 , \283 , \284 , \285 , \286 , \287 , \288 ,
         \289 , \290 , \291 , \292 , \293 , \294 , \295 , \296 , \297 , \298 ,
         \299 , \300 , \301 , \302 , \303 , \304 , \305 , \306 , \307 , \308 ,
         \309 , \310 , \311 , \312 , \313 , \314 , \315 , \316 , \317 , \318 ,
         \319 , \320 , \321 , \322 , \323 , \324 , \325 , \326 , \327 , \328 ,
         \329 , \330 , \331 , \332 , \333 , \334 , \335 , \336 , \337 , \338 ,
         \339 , \340 , \341 , \342 , \343 , \344 , \345 , \346 , \347 , \348 ,
         \349 , \350 , \351 , \352 , \353 , \354 , \355 , \356 , \357 , \358 ,
         \359 , \360 , \361 , \362 , \363 , \364 , \365 , \366 , \367 , \368 ,
         \369 , \370 , \371 , \372 , \373 , \374 , \375 , \376 , \377 , \378 ,
         \379 , \380 , \381 , \382 , \383 , \384 , \385 , \386 , \387 , \388 ,
         \389 , \390 , \391 , \392 , \393 , \394 , \395 , \396 , \397 , \398 ,
         \399 , \400 , \401 , \402 , \403 , \404 , \405 , \406 , \407 , \408 ,
         \409 , \410 , \411 , \412 , \413 , \414 , \415 , \416 , \417 , \418 ,
         \419 , \420 , \421 , \422 , \423 , \424 , \425 , \426 , \427 , \428 ,
         \429 , \430 , \431 , \432 , \433 , \434 , \435 , \436 , \437 , \438 ,
         \439 , \440 , \441 , \442 , \443 , \444 , \445 , \446 , \447 , \448 ,
         \449 , \450 , \451 , \452 , \453 , \454 , \455 , \456 , \457 , \458 ,
         \459 , \460 , \461 , \462 , \463 , \464 , \465 , \466 , \467 , \468 ,
         \469 , \470 , \471 , \472 , \473 , \474 , \475 , \476 , \477 , \478 ,
         \479 , \480 , \481 , \482 , \483 , \484 , \485 , \486 , \487 , \488 ,
         \489 , \490 , \491 , \492 , \493 , \494 , \495 , \496 , \497 , \498 ,
         \499 , \500 , \501 , \502 , \503 , \504 , \505 , \506 , \507 , \508 ,
         \509 , \510 , \511 , \512 , \513 , \514 , \515 , \516 , \517 , \518 ,
         \519 , \520 , \521 , \522 , \523 , \524 , \525 , \526 , \527 , \528 ,
         \529 , \530 , \531 , \532 , \533 , \534 , \535 , \536 , \537 , \538 ,
         \539 , \540 , \541 , \542 , \543 , \544 , \545 , \546 , \547 , \548 ,
         \549 , \550 , \551 , \552 , \553 , \554 , \555 , \556 , \557 , \558 ,
         \559 , \560 , \561 , \562 , \563 , \564 , \565 , \566 , \567 , \568 ,
         \569 , \570 , \571 , \572 , \573 , \574 , \575 , \576 , \577 , \578 ,
         \579 , \580 , \581 , \582 , \583 , \584 , \585 , \586 , \587 , \588 ,
         \589 , \590 , \591 , \592 , \593 , \594 , \595 , \596 , \597 , \598 ,
         \599 , \600 , \601 , \602 , \603 , \604 , \605 , \606 , \607 , \608 ,
         \609 , \610 , \611 , \612 , \613 , \614 , \615 , \616 , \617 , \618 ,
         \619 , \620 , \621 , \622 , \623 , \624 , \625 , \626 , \627 , \628 ,
         \629 , \630 , \631 , \632 , \633 , \634 , \635 , \636 , \637 , \638 ,
         \639 , \640 , \641 , \642 , \643 , \644 , \645 , \646 , \647 , \648 ,
         \649 , \650 , \651 , \652 , \653 , \654 , \655 , \656 , \657 , \658 ,
         \659 , \660 , \661 , \662 , \663 , \664 , \665 , \666 , \667 , \668 ,
         \669 , \670 , \671 , \672 , \673 , \674 , \675 , \676 , \677 , \678 ,
         \679 , \680 , \681 , \682 , \683 , \684 , \685 , \686 , \687 , \688 ,
         \689 , \690 , \691 , \692 , \693 , \694 , \695 , \696 , \697 , \698 ,
         \699 , \700 , \701 , \702 , \703 , \704 , \705 , \706 , \707 , \708 ,
         \709 , \710 , \711 , \712 , \713 , \714 , \715 , \716 , \717 , \718 ,
         \719 , \720 , \721 , \722 , \723 , \724 , \725 , \726 , \727 , \728 ,
         \729 , \730 , \731 , \732 , \733 , \734 , \735 , \736 , \737 , \738 ,
         \739 , \740 , \741 , \742 , \743 , \744 , \745 , \746 , \747 , \748 ,
         \749 , \750 , \751 , \752 , \753 , \754 , \755 , \756 , \757 , \758 ,
         \759 , \760 , \761 , \762 , \763 , \764 , \765 , \766 , \767 , \768 ,
         \769 , \770 , \771 , \772 , \773 , \774 , \775 , \776 , \777 , \778 ,
         \779 , \780 , \781 , \782 , \783 , \784 , \785 , \786 , \787 , \788 ,
         \789 , \790 , \791 , \792 , \793 , \794 , \795 , \796 , \797 , \798 ,
         \799 , \800 , \801 , \802 , \803 , \804 , \805 , \806 , \807 , \808 ,
         \809 , \810 , \811 , \812 , \813 , \814 , \815 , \816 , \817 , \818 ,
         \819 , \820 , \821 , \822 , \823 , \824 , \825 , \826 , \827 , \828 ,
         \829 , \830 , \831 , \832 , \833 , \834 , \835 , \836 , \837 , \838 ,
         \839 , \840 , \841 , \842 , \843 , \844 , \845 , \846 , \847 , \848 ,
         \849 , \850 , \851 , \852 , \853 , \854 , \855 , \856 , \857 , \858 ,
         \859 , \860 , \861 , \862 , \863 , \864 , \865 , \866 , \867 , \868 ,
         \869 , \870 , \871 , \872 , \873 , \874 , \875 , \876 , \877 , \878 ,
         \879 , \880 , \881 , \882 , \883 , \884 , \885 , \886 , \887 , \888 ,
         \889 , \890 , \891 , \892 , \893 , \894 , \895 , \896 , \897 , \898 ,
         \899 , \900 , \901 , \902 , \903 , \904 , \905 , \906 , \907 , \908 ,
         \909 , \910 , \911 , \912 , \913 , \914 , \915 , \916 , \917 , \918 ,
         \919 , \920 , \921 , \922 , \923 , \924 , \925 , \926 , \927 , \928 ,
         \929 , \930 , \931 , \932 , \933 , \934 , \935 , \936 , \937 , \938 ,
         \939 , \940 , \941 , \942 , \943 , \944 , \945 , \946 , \947 , \948 ,
         \949 , \950 , \951 , \952 , \953 , \954 , \955 , \956 , \957 , \958 ,
         \959 , \960 , \961 , \962 , \963 , \964 , \965 , \966 , \967 , \968 ,
         \969 , \970 , \971 , \972 , \973 , \974 , \975 , \976 , \977 , \978 ,
         \979 , \980 , \981 , \982 , \983 , \984 , \985 , \986 , \987 , \988 ,
         \989 , \990 , \991 , \992 , \993 , \994 , \995 , \996 , \997 , \998 ,
         \999 , \1000 , \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 , \1008 ,
         \1009 , \1010 , \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 , \1018 ,
         \1019 , \1020 , \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 , \1028 ,
         \1029 , \1030 , \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 , \1038 ,
         \1039 , \1040 , \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 , \1048 ,
         \1049 , \1050 , \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 , \1058 ,
         \1059 , \1060 , \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 , \1068 ,
         \1069_nG5577 , \1070 , \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 , \1078 ,
         \1079 , \1080 , \1081 , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 , \1088 ,
         \1089 , \1090 , \1091 , \1092 , \1093 , \1094 , \1095 , \1096 , \1097 , \1098 ,
         \1099 , \1100 , \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 , \1108 ,
         \1109 , \1110 , \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117 , \1118 ,
         \1119 , \1120 , \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 , \1128 ,
         \1129 , \1130 , \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 , \1138 ,
         \1139 , \1140 , \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 , \1148 ,
         \1149 , \1150 , \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 , \1158 ,
         \1159 , \1160 , \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 , \1168 ,
         \1169 , \1170_nG5575 , \1171 , \1172 , \1173 , \1174 , \1175 , \1176 , \1177 , \1178 ,
         \1179 , \1180 , \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 , \1188 ,
         \1189 , \1190 , \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 , \1198 ,
         \1199 , \1200 , \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 , \1208 ,
         \1209 , \1210 , \1211 , \1212 , \1213 , \1214 , \1215 , \1216 , \1217 , \1218 ,
         \1219 , \1220 , \1221 , \1222 , \1223 , \1224 , \1225 , \1226 , \1227 , \1228 ,
         \1229 , \1230 , \1231 , \1232 , \1233 , \1234 , \1235 , \1236 , \1237 , \1238 ,
         \1239 , \1240 , \1241 , \1242 , \1243 , \1244 , \1245 , \1246 , \1247 , \1248 ,
         \1249 , \1250 , \1251 , \1252 , \1253 , \1254 , \1255 , \1256 , \1257 , \1258 ,
         \1259 , \1260 , \1261 , \1262 , \1263 , \1264 , \1265 , \1266 , \1267 , \1268 ,
         \1269 , \1270 , \1271 , \1272 , \1273 , \1274 , \1275 , \1276 , \1277 , \1278_nG5573 ,
         \1279 , \1280 , \1281 , \1282 , \1283 , \1284 , \1285 , \1286 , \1287 , \1288 ,
         \1289 , \1290 , \1291 , \1292 , \1293 , \1294 , \1295 , \1296 , \1297 , \1298 ,
         \1299 , \1300 , \1301 , \1302 , \1303 , \1304 , \1305 , \1306 , \1307 , \1308 ,
         \1309 , \1310 , \1311 , \1312 , \1313 , \1314 , \1315 , \1316 , \1317 , \1318 ,
         \1319 , \1320 , \1321 , \1322 , \1323 , \1324 , \1325 , \1326 , \1327 , \1328 ,
         \1329 , \1330 , \1331 , \1332 , \1333 , \1334 , \1335 , \1336 , \1337 , \1338 ,
         \1339 , \1340 , \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 ,
         \1349 , \1350 , \1351 , \1352 , \1353 , \1354 , \1355 , \1356 , \1357 , \1358 ,
         \1359 , \1360 , \1361 , \1362 , \1363 , \1364 , \1365 , \1366 , \1367 , \1368 ,
         \1369 , \1370 , \1371 , \1372 , \1373 , \1374 , \1375 , \1376 , \1377 , \1378 ,
         \1379 , \1380 , \1381 , \1382 , \1383 , \1384 , \1385 , \1386 , \1387 , \1388 ,
         \1389_nG5571 , \1390 , \1391 , \1392 , \1393 , \1394 , \1395 , \1396 , \1397 , \1398 ,
         \1399 , \1400 , \1401 , \1402 , \1403 , \1404 , \1405 , \1406 , \1407 , \1408 ,
         \1409 , \1410 , \1411 , \1412 , \1413 , \1414 , \1415 , \1416 , \1417 , \1418 ,
         \1419 , \1420 , \1421 , \1422 , \1423 , \1424 , \1425 , \1426 , \1427 , \1428 ,
         \1429 , \1430 , \1431 , \1432 , \1433 , \1434 , \1435 , \1436 , \1437 , \1438 ,
         \1439 , \1440 , \1441 , \1442 , \1443 , \1444 , \1445 , \1446 , \1447 , \1448 ,
         \1449 , \1450 , \1451 , \1452 , \1453 , \1454 , \1455 , \1456 , \1457 , \1458 ,
         \1459 , \1460 , \1461 , \1462 , \1463 , \1464 , \1465 , \1466 , \1467 , \1468 ,
         \1469 , \1470 , \1471 , \1472 , \1473 , \1474 , \1475 , \1476 , \1477 , \1478 ,
         \1479 , \1480 , \1481 , \1482 , \1483 , \1484 , \1485 , \1486 , \1487 , \1488 ,
         \1489 , \1490 , \1491 , \1492 , \1493 , \1494 , \1495 , \1496 , \1497 , \1498 ,
         \1499 , \1500 , \1501 , \1502 , \1503 , \1504 , \1505 , \1506 , \1507_nG556f , \1508 ,
         \1509 , \1510 , \1511 , \1512 , \1513 , \1514 , \1515 , \1516 , \1517 , \1518 ,
         \1519 , \1520 , \1521 , \1522 , \1523 , \1524 , \1525 , \1526 , \1527 , \1528 ,
         \1529 , \1530 , \1531 , \1532 , \1533 , \1534 , \1535 , \1536 , \1537 , \1538 ,
         \1539 , \1540 , \1541 , \1542 , \1543 , \1544 , \1545 , \1546 , \1547 , \1548 ,
         \1549 , \1550 , \1551 , \1552 , \1553 , \1554 , \1555 , \1556 , \1557 , \1558 ,
         \1559 , \1560 , \1561 , \1562 , \1563 , \1564 , \1565 , \1566 , \1567 , \1568 ,
         \1569 , \1570 , \1571 , \1572 , \1573 , \1574 , \1575 , \1576 , \1577 , \1578 ,
         \1579 , \1580 , \1581 , \1582 , \1583 , \1584 , \1585 , \1586 , \1587 , \1588 ,
         \1589 , \1590 , \1591 , \1592 , \1593 , \1594 , \1595 , \1596 , \1597 , \1598 ,
         \1599 , \1600 , \1601 , \1602 , \1603 , \1604 , \1605 , \1606 , \1607 , \1608 ,
         \1609 , \1610 , \1611 , \1612 , \1613 , \1614 , \1615 , \1616 , \1617 , \1618 ,
         \1619 , \1620 , \1621 , \1622 , \1623 , \1624 , \1625 , \1626 , \1627 , \1628_nG556d ,
         \1629 , \1630 , \1631 , \1632 , \1633 , \1634 , \1635 , \1636 , \1637 , \1638 ,
         \1639 , \1640 , \1641 , \1642 , \1643 , \1644 , \1645 , \1646 , \1647 , \1648 ,
         \1649 , \1650 , \1651 , \1652 , \1653 , \1654 , \1655 , \1656 , \1657 , \1658 ,
         \1659 , \1660 , \1661 , \1662 , \1663 , \1664 , \1665 , \1666 , \1667 , \1668 ,
         \1669 , \1670 , \1671 , \1672 , \1673 , \1674 , \1675 , \1676 , \1677 , \1678 ,
         \1679 , \1680 , \1681 , \1682 , \1683 , \1684 , \1685 , \1686 , \1687 , \1688 ,
         \1689 , \1690 , \1691 , \1692 , \1693 , \1694 , \1695 , \1696 , \1697 , \1698 ,
         \1699 , \1700 , \1701 , \1702 , \1703 , \1704 , \1705 , \1706 , \1707 , \1708 ,
         \1709 , \1710 , \1711 , \1712 , \1713 , \1714 , \1715 , \1716 , \1717 , \1718 ,
         \1719 , \1720 , \1721 , \1722 , \1723 , \1724 , \1725 , \1726 , \1727 , \1728 ,
         \1729 , \1730 , \1731 , \1732 , \1733 , \1734 , \1735 , \1736 , \1737 , \1738 ,
         \1739 , \1740 , \1741 , \1742 , \1743 , \1744 , \1745 , \1746 , \1747 , \1748 ,
         \1749 , \1750 , \1751 , \1752 , \1753 , \1754 , \1755 , \1756_nG556b , \1757 , \1758 ,
         \1759 , \1760 , \1761 , \1762 , \1763 , \1764 , \1765 , \1766 , \1767 , \1768 ,
         \1769 , \1770 , \1771 , \1772 , \1773 , \1774 , \1775 , \1776 , \1777 , \1778 ,
         \1779 , \1780 , \1781 , \1782 , \1783 , \1784 , \1785 , \1786 , \1787 , \1788 ,
         \1789 , \1790 , \1791 , \1792 , \1793 , \1794 , \1795 , \1796 , \1797 , \1798 ,
         \1799 , \1800 , \1801 , \1802 , \1803 , \1804 , \1805 , \1806 , \1807 , \1808 ,
         \1809 , \1810 , \1811 , \1812 , \1813 , \1814 , \1815 , \1816 , \1817 , \1818 ,
         \1819 , \1820 , \1821 , \1822 , \1823 , \1824 , \1825 , \1826 , \1827 , \1828 ,
         \1829 , \1830 , \1831 , \1832 , \1833 , \1834 , \1835 , \1836 , \1837 , \1838 ,
         \1839 , \1840 , \1841 , \1842 , \1843 , \1844 , \1845 , \1846 , \1847 , \1848 ,
         \1849 , \1850 , \1851 , \1852 , \1853 , \1854 , \1855 , \1856 , \1857 , \1858 ,
         \1859 , \1860 , \1861 , \1862 , \1863 , \1864 , \1865 , \1866 , \1867 , \1868 ,
         \1869 , \1870 , \1871 , \1872 , \1873 , \1874 , \1875 , \1876 , \1877 , \1878 ,
         \1879 , \1880 , \1881 , \1882 , \1883 , \1884 , \1885 , \1886 , \1887_nG5569 , \1888 ,
         \1889 , \1890 , \1891 , \1892 , \1893 , \1894 , \1895 , \1896 , \1897 , \1898 ,
         \1899 , \1900 , \1901 , \1902 , \1903 , \1904 , \1905 , \1906 , \1907 , \1908 ,
         \1909 , \1910 , \1911 , \1912 , \1913 , \1914 , \1915 , \1916 , \1917 , \1918 ,
         \1919 , \1920 , \1921 , \1922 , \1923 , \1924 , \1925 , \1926 , \1927 , \1928 ,
         \1929 , \1930 , \1931 , \1932 , \1933 , \1934 , \1935 , \1936 , \1937 , \1938 ,
         \1939 , \1940 , \1941 , \1942 , \1943 , \1944 , \1945 , \1946 , \1947 , \1948 ,
         \1949 , \1950 , \1951 , \1952 , \1953 , \1954 , \1955 , \1956 , \1957 , \1958 ,
         \1959 , \1960 , \1961 , \1962 , \1963 , \1964 , \1965 , \1966 , \1967 , \1968 ,
         \1969 , \1970 , \1971 , \1972 , \1973 , \1974 , \1975 , \1976 , \1977 , \1978 ,
         \1979 , \1980 , \1981 , \1982 , \1983 , \1984 , \1985 , \1986 , \1987 , \1988 ,
         \1989 , \1990 , \1991 , \1992 , \1993 , \1994 , \1995 , \1996 , \1997 , \1998 ,
         \1999 , \2000 , \2001 , \2002 , \2003 , \2004 , \2005 , \2006 , \2007 , \2008 ,
         \2009 , \2010 , \2011 , \2012 , \2013 , \2014 , \2015 , \2016 , \2017 , \2018 ,
         \2019 , \2020 , \2021 , \2022 , \2023 , \2024 , \2025_nG5567 , \2026 , \2027 , \2028 ,
         \2029 , \2030 , \2031 , \2032 , \2033 , \2034 , \2035 , \2036 , \2037 , \2038 ,
         \2039 , \2040 , \2041 , \2042 , \2043 , \2044 , \2045 , \2046 , \2047 , \2048 ,
         \2049 , \2050 , \2051 , \2052 , \2053 , \2054 , \2055 , \2056 , \2057 , \2058 ,
         \2059 , \2060 , \2061 , \2062 , \2063 , \2064 , \2065 , \2066 , \2067 , \2068 ,
         \2069 , \2070 , \2071 , \2072 , \2073 , \2074 , \2075 , \2076 , \2077 , \2078 ,
         \2079 , \2080 , \2081 , \2082 , \2083 , \2084 , \2085 , \2086 , \2087 , \2088 ,
         \2089 , \2090 , \2091 , \2092 , \2093 , \2094 , \2095 , \2096 , \2097 , \2098 ,
         \2099 , \2100 , \2101 , \2102 , \2103 , \2104 , \2105 , \2106 , \2107 , \2108 ,
         \2109 , \2110 , \2111 , \2112 , \2113 , \2114 , \2115 , \2116 , \2117 , \2118 ,
         \2119 , \2120 , \2121 , \2122 , \2123 , \2124 , \2125 , \2126 , \2127 , \2128 ,
         \2129 , \2130 , \2131 , \2132 , \2133 , \2134 , \2135 , \2136 , \2137 , \2138 ,
         \2139 , \2140 , \2141 , \2142 , \2143 , \2144 , \2145 , \2146 , \2147 , \2148 ,
         \2149 , \2150 , \2151 , \2152 , \2153 , \2154 , \2155 , \2156 , \2157 , \2158 ,
         \2159 , \2160 , \2161 , \2162 , \2163 , \2164 , \2165 , \2166_nG5565 , \2167 , \2168 ,
         \2169 , \2170 , \2171 , \2172 , \2173 , \2174 , \2175 , \2176 , \2177 , \2178 ,
         \2179 , \2180 , \2181 , \2182 , \2183 , \2184 , \2185 , \2186 , \2187 , \2188 ,
         \2189 , \2190 , \2191 , \2192 , \2193 , \2194 , \2195 , \2196 , \2197 , \2198 ,
         \2199 , \2200 , \2201 , \2202 , \2203 , \2204 , \2205 , \2206 , \2207 , \2208 ,
         \2209 , \2210 , \2211 , \2212 , \2213 , \2214 , \2215 , \2216 , \2217 , \2218 ,
         \2219 , \2220 , \2221 , \2222 , \2223 , \2224 , \2225 , \2226 , \2227 , \2228 ,
         \2229 , \2230 , \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 , \2238 ,
         \2239 , \2240 , \2241 , \2242 , \2243 , \2244 , \2245 , \2246 , \2247 , \2248 ,
         \2249 , \2250 , \2251 , \2252 , \2253 , \2254 , \2255 , \2256 , \2257 , \2258 ,
         \2259 , \2260 , \2261 , \2262 , \2263 , \2264 , \2265 , \2266 , \2267 , \2268 ,
         \2269 , \2270 , \2271 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 , \2278 ,
         \2279 , \2280 , \2281 , \2282 , \2283 , \2284 , \2285 , \2286 , \2287 , \2288 ,
         \2289 , \2290 , \2291 , \2292 , \2293 , \2294 , \2295 , \2296 , \2297 , \2298 ,
         \2299 , \2300 , \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 , \2308 ,
         \2309 , \2310 , \2311 , \2312 , \2313 , \2314_nG5563 , \2315 , \2316 , \2317 , \2318 ,
         \2319 , \2320 , \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 , \2328 ,
         \2329 , \2330 , \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 , \2338 ,
         \2339 , \2340 , \2341 , \2342 , \2343 , \2344 , \2345 , \2346 , \2347 , \2348 ,
         \2349 , \2350 , \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 , \2358 ,
         \2359 , \2360 , \2361 , \2362 , \2363 , \2364 , \2365 , \2366 , \2367 , \2368 ,
         \2369 , \2370 , \2371 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 , \2378 ,
         \2379 , \2380 , \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 , \2388 ,
         \2389 , \2390 , \2391 , \2392 , \2393 , \2394 , \2395 , \2396 , \2397 , \2398 ,
         \2399 , \2400 , \2401 , \2402 , \2403 , \2404 , \2405 , \2406 , \2407 , \2408 ,
         \2409 , \2410 , \2411 , \2412 , \2413 , \2414 , \2415 , \2416 , \2417 , \2418 ,
         \2419 , \2420 , \2421 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 , \2428 ,
         \2429 , \2430 , \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 , \2438 ,
         \2439 , \2440 , \2441 , \2442 , \2443 , \2444 , \2445 , \2446 , \2447 , \2448 ,
         \2449 , \2450 , \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 , \2458 ,
         \2459 , \2460 , \2461 , \2462 , \2463 , \2464 , \2465_nG5561 , \2466 , \2467 , \2468 ,
         \2469 , \2470 , \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 , \2478 ,
         \2479 , \2480 , \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 , \2488 ,
         \2489 , \2490 , \2491 , \2492 , \2493 , \2494 , \2495 , \2496 , \2497 , \2498 ,
         \2499 , \2500 , \2501 , \2502 , \2503 , \2504 , \2505 , \2506 , \2507 , \2508 ,
         \2509 , \2510 , \2511 , \2512 , \2513 , \2514 , \2515 , \2516 , \2517 , \2518 ,
         \2519 , \2520 , \2521 , \2522 , \2523 , \2524 , \2525 , \2526 , \2527 , \2528 ,
         \2529 , \2530 , \2531 , \2532 , \2533 , \2534 , \2535 , \2536 , \2537 , \2538 ,
         \2539 , \2540 , \2541 , \2542 , \2543 , \2544 , \2545 , \2546 , \2547 , \2548 ,
         \2549 , \2550 , \2551 , \2552 , \2553 , \2554 , \2555 , \2556 , \2557 , \2558 ,
         \2559 , \2560 , \2561 , \2562 , \2563 , \2564 , \2565 , \2566 , \2567 , \2568 ,
         \2569 , \2570 , \2571 , \2572 , \2573 , \2574 , \2575 , \2576 , \2577 , \2578 ,
         \2579 , \2580 , \2581 , \2582 , \2583 , \2584 , \2585 , \2586 , \2587 , \2588 ,
         \2589 , \2590 , \2591 , \2592 , \2593 , \2594 , \2595 , \2596 , \2597 , \2598 ,
         \2599 , \2600 , \2601 , \2602 , \2603 , \2604 , \2605 , \2606 , \2607 , \2608 ,
         \2609 , \2610 , \2611 , \2612 , \2613 , \2614 , \2615 , \2616 , \2617 , \2618 ,
         \2619 , \2620 , \2621 , \2622 , \2623_nG555f , \2624 , \2625 , \2626 , \2627 , \2628 ,
         \2629 , \2630 , \2631 , \2632 , \2633 , \2634 , \2635 , \2636 , \2637 , \2638 ,
         \2639 , \2640 , \2641 , \2642 , \2643 , \2644 , \2645 , \2646 , \2647 , \2648 ,
         \2649 , \2650 , \2651 , \2652 , \2653 , \2654 , \2655 , \2656 , \2657 , \2658 ,
         \2659 , \2660 , \2661 , \2662 , \2663 , \2664 , \2665 , \2666 , \2667 , \2668 ,
         \2669 , \2670 , \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 , \2678 ,
         \2679 , \2680 , \2681 , \2682 , \2683 , \2684 , \2685 , \2686 , \2687 , \2688 ,
         \2689 , \2690 , \2691 , \2692 , \2693 , \2694 , \2695 , \2696 , \2697 , \2698 ,
         \2699 , \2700 , \2701 , \2702 , \2703 , \2704 , \2705 , \2706 , \2707 , \2708 ,
         \2709 , \2710 , \2711 , \2712 , \2713 , \2714 , \2715 , \2716 , \2717 , \2718 ,
         \2719 , \2720 , \2721 , \2722 , \2723 , \2724 , \2725 , \2726 , \2727 , \2728 ,
         \2729 , \2730 , \2731 , \2732 , \2733 , \2734 , \2735 , \2736 , \2737 , \2738 ,
         \2739 , \2740 , \2741 , \2742 , \2743 , \2744 , \2745 , \2746 , \2747 , \2748 ,
         \2749 , \2750 , \2751 , \2752 , \2753 , \2754 , \2755 , \2756 , \2757 , \2758 ,
         \2759 , \2760 , \2761 , \2762 , \2763 , \2764 , \2765 , \2766 , \2767 , \2768 ,
         \2769 , \2770 , \2771 , \2772 , \2773 , \2774 , \2775 , \2776 , \2777 , \2778 ,
         \2779 , \2780 , \2781 , \2782 , \2783 , \2784_nG555d , \2785 , \2786 , \2787 , \2788 ,
         \2789 , \2790 , \2791 , \2792 , \2793 , \2794 , \2795 , \2796 , \2797 , \2798 ,
         \2799 , \2800 , \2801 , \2802 , \2803 , \2804 , \2805 , \2806 , \2807 , \2808 ,
         \2809 , \2810 , \2811 , \2812 , \2813 , \2814 , \2815 , \2816 , \2817 , \2818 ,
         \2819 , \2820 , \2821 , \2822 , \2823 , \2824 , \2825 , \2826 , \2827 , \2828 ,
         \2829 , \2830 , \2831 , \2832 , \2833 , \2834 , \2835 , \2836 , \2837 , \2838 ,
         \2839 , \2840 , \2841 , \2842 , \2843 , \2844 , \2845 , \2846 , \2847 , \2848 ,
         \2849 , \2850 , \2851 , \2852 , \2853 , \2854 , \2855 , \2856 , \2857 , \2858 ,
         \2859 , \2860 , \2861 , \2862 , \2863 , \2864 , \2865 , \2866 , \2867 , \2868 ,
         \2869 , \2870 , \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 , \2878 ,
         \2879 , \2880 , \2881 , \2882 , \2883 , \2884 , \2885 , \2886 , \2887 , \2888 ,
         \2889 , \2890 , \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 , \2898 ,
         \2899 , \2900 , \2901 , \2902 , \2903 , \2904 , \2905 , \2906 , \2907 , \2908 ,
         \2909 , \2910 , \2911 , \2912 , \2913 , \2914 , \2915 , \2916 , \2917 , \2918 ,
         \2919 , \2920 , \2921 , \2922 , \2923 , \2924 , \2925 , \2926 , \2927 , \2928 ,
         \2929 , \2930 , \2931 , \2932 , \2933 , \2934 , \2935 , \2936 , \2937 , \2938 ,
         \2939 , \2940 , \2941 , \2942 , \2943 , \2944 , \2945 , \2946 , \2947 , \2948 ,
         \2949 , \2950 , \2951 , \2952_nG555b , \2953 , \2954 , \2955 , \2956 , \2957 , \2958 ,
         \2959 , \2960 , \2961 , \2962 , \2963 , \2964 , \2965 , \2966 , \2967 , \2968 ,
         \2969 , \2970 , \2971 , \2972 , \2973 , \2974 , \2975 , \2976 , \2977 , \2978 ,
         \2979 , \2980 , \2981 , \2982 , \2983 , \2984 , \2985 , \2986 , \2987 , \2988 ,
         \2989 , \2990 , \2991 , \2992 , \2993 , \2994 , \2995 , \2996 , \2997 , \2998 ,
         \2999 , \3000 , \3001 , \3002 , \3003 , \3004 , \3005 , \3006 , \3007 , \3008 ,
         \3009 , \3010 , \3011 , \3012 , \3013 , \3014 , \3015 , \3016 , \3017 , \3018 ,
         \3019 , \3020 , \3021 , \3022 , \3023 , \3024 , \3025 , \3026 , \3027 , \3028 ,
         \3029 , \3030 , \3031 , \3032 , \3033 , \3034 , \3035 , \3036 , \3037 , \3038 ,
         \3039 , \3040 , \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 , \3048 ,
         \3049 , \3050 , \3051 , \3052 , \3053 , \3054 , \3055 , \3056 , \3057 , \3058 ,
         \3059 , \3060 , \3061 , \3062 , \3063 , \3064 , \3065 , \3066 , \3067 , \3068 ,
         \3069 , \3070 , \3071 , \3072 , \3073 , \3074 , \3075 , \3076 , \3077 , \3078 ,
         \3079 , \3080 , \3081 , \3082 , \3083 , \3084 , \3085 , \3086 , \3087 , \3088 ,
         \3089 , \3090 , \3091 , \3092 , \3093 , \3094 , \3095 , \3096 , \3097 , \3098 ,
         \3099 , \3100 , \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 , \3108 ,
         \3109 , \3110 , \3111 , \3112 , \3113 , \3114 , \3115 , \3116 , \3117 , \3118 ,
         \3119 , \3120 , \3121 , \3122 , \3123_nG5559 , \3124 , \3125 , \3126 , \3127 , \3128 ,
         \3129 , \3130 , \3131 , \3132 , \3133 , \3134 , \3135 , \3136 , \3137 , \3138 ,
         \3139 , \3140 , \3141 , \3142 , \3143 , \3144 , \3145 , \3146 , \3147 , \3148 ,
         \3149 , \3150 , \3151 , \3152 , \3153 , \3154 , \3155 , \3156 , \3157 , \3158 ,
         \3159 , \3160 , \3161 , \3162 , \3163 , \3164 , \3165 , \3166 , \3167 , \3168 ,
         \3169 , \3170 , \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 , \3178 ,
         \3179 , \3180 , \3181 , \3182 , \3183 , \3184 , \3185 , \3186 , \3187 , \3188 ,
         \3189 , \3190 , \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 , \3198 ,
         \3199 , \3200 , \3201 , \3202 , \3203 , \3204 , \3205 , \3206 , \3207 , \3208 ,
         \3209 , \3210 , \3211 , \3212 , \3213 , \3214 , \3215 , \3216 , \3217 , \3218 ,
         \3219 , \3220 , \3221 , \3222 , \3223 , \3224 , \3225 , \3226 , \3227 , \3228 ,
         \3229 , \3230 , \3231 , \3232 , \3233 , \3234 , \3235 , \3236 , \3237 , \3238 ,
         \3239 , \3240 , \3241 , \3242 , \3243 , \3244 , \3245 , \3246 , \3247 , \3248 ,
         \3249 , \3250 , \3251 , \3252 , \3253 , \3254 , \3255 , \3256 , \3257 , \3258 ,
         \3259 , \3260 , \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 , \3268 ,
         \3269 , \3270 , \3271 , \3272 , \3273 , \3274 , \3275 , \3276 , \3277 , \3278 ,
         \3279 , \3280 , \3281 , \3282 , \3283 , \3284 , \3285 , \3286 , \3287 , \3288 ,
         \3289 , \3290 , \3291 , \3292 , \3293 , \3294 , \3295 , \3296 , \3297 , \3298 ,
         \3299 , \3300 , \3301_nG5557 , \3302 , \3303 , \3304 , \3305 , \3306 , \3307 , \3308 ,
         \3309 , \3310 , \3311 , \3312 , \3313 , \3314 , \3315 , \3316 , \3317 , \3318 ,
         \3319 , \3320 , \3321 , \3322 , \3323 , \3324 , \3325 , \3326 , \3327 , \3328 ,
         \3329 , \3330 , \3331 , \3332 , \3333 , \3334 , \3335 , \3336 , \3337 , \3338 ,
         \3339 , \3340 , \3341 , \3342 , \3343 , \3344 , \3345 , \3346 , \3347 , \3348 ,
         \3349 , \3350 , \3351 , \3352 , \3353 , \3354 , \3355 , \3356 , \3357 , \3358 ,
         \3359 , \3360 , \3361 , \3362 , \3363 , \3364 , \3365 , \3366 , \3367 , \3368 ,
         \3369 , \3370 , \3371 , \3372 , \3373 , \3374 , \3375 , \3376 , \3377 , \3378 ,
         \3379 , \3380 , \3381 , \3382 , \3383 , \3384 , \3385 , \3386 , \3387 , \3388 ,
         \3389 , \3390 , \3391 , \3392 , \3393 , \3394 , \3395 , \3396 , \3397 , \3398 ,
         \3399 , \3400 , \3401 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 , \3408 ,
         \3409 , \3410 , \3411 , \3412 , \3413 , \3414 , \3415 , \3416 , \3417 , \3418 ,
         \3419 , \3420 , \3421 , \3422 , \3423 , \3424 , \3425 , \3426 , \3427 , \3428 ,
         \3429 , \3430 , \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 , \3438 ,
         \3439 , \3440 , \3441 , \3442 , \3443 , \3444 , \3445 , \3446 , \3447 , \3448 ,
         \3449 , \3450 , \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 , \3458 ,
         \3459 , \3460 , \3461 , \3462 , \3463 , \3464 , \3465 , \3466 , \3467 , \3468 ,
         \3469 , \3470 , \3471 , \3472 , \3473 , \3474 , \3475 , \3476 , \3477 , \3478 ,
         \3479 , \3480 , \3481 , \3482_nG5555 , \3483 , \3484 , \3485 , \3486 , \3487 , \3488 ,
         \3489 , \3490 , \3491 , \3492 , \3493 , \3494 , \3495 , \3496 , \3497 , \3498 ,
         \3499 , \3500 , \3501 , \3502 , \3503 , \3504 , \3505 , \3506 , \3507 , \3508 ,
         \3509 , \3510 , \3511 , \3512 , \3513 , \3514 , \3515 , \3516 , \3517 , \3518 ,
         \3519 , \3520 , \3521 , \3522 , \3523 , \3524 , \3525 , \3526 , \3527 , \3528 ,
         \3529 , \3530 , \3531 , \3532 , \3533 , \3534 , \3535 , \3536 , \3537 , \3538 ,
         \3539 , \3540 , \3541 , \3542 , \3543 , \3544 , \3545 , \3546 , \3547 , \3548 ,
         \3549 , \3550 , \3551 , \3552 , \3553 , \3554 , \3555 , \3556 , \3557 , \3558 ,
         \3559 , \3560 , \3561 , \3562 , \3563 , \3564 , \3565 , \3566 , \3567 , \3568 ,
         \3569 , \3570 , \3571 , \3572 , \3573 , \3574 , \3575 , \3576 , \3577 , \3578 ,
         \3579 , \3580 , \3581 , \3582 , \3583 , \3584 , \3585 , \3586 , \3587 , \3588 ,
         \3589 , \3590 , \3591 , \3592 , \3593 , \3594 , \3595 , \3596 , \3597 , \3598 ,
         \3599 , \3600 , \3601 , \3602 , \3603 , \3604 , \3605 , \3606 , \3607 , \3608 ,
         \3609 , \3610 , \3611 , \3612 , \3613 , \3614 , \3615 , \3616 , \3617 , \3618 ,
         \3619 , \3620 , \3621 , \3622 , \3623 , \3624 , \3625 , \3626 , \3627 , \3628 ,
         \3629 , \3630 , \3631 , \3632 , \3633 , \3634 , \3635 , \3636 , \3637 , \3638 ,
         \3639 , \3640 , \3641 , \3642 , \3643 , \3644 , \3645 , \3646 , \3647 , \3648 ,
         \3649 , \3650 , \3651 , \3652 , \3653 , \3654 , \3655 , \3656 , \3657 , \3658 ,
         \3659 , \3660 , \3661 , \3662 , \3663 , \3664 , \3665 , \3666 , \3667 , \3668 ,
         \3669 , \3670_nG5553 , \3671 , \3672 , \3673 , \3674 , \3675 , \3676 , \3677 , \3678 ,
         \3679 , \3680 , \3681 , \3682 , \3683 , \3684 , \3685 , \3686 , \3687 , \3688 ,
         \3689 , \3690 , \3691 , \3692 , \3693 , \3694 , \3695 , \3696 , \3697 , \3698 ,
         \3699 , \3700 , \3701 , \3702 , \3703 , \3704 , \3705 , \3706 , \3707 , \3708 ,
         \3709 , \3710 , \3711 , \3712 , \3713 , \3714 , \3715 , \3716 , \3717 , \3718 ,
         \3719 , \3720 , \3721 , \3722 , \3723 , \3724 , \3725 , \3726 , \3727 , \3728 ,
         \3729 , \3730 , \3731 , \3732 , \3733 , \3734 , \3735 , \3736 , \3737 , \3738 ,
         \3739 , \3740 , \3741 , \3742 , \3743 , \3744 , \3745 , \3746 , \3747 , \3748 ,
         \3749 , \3750 , \3751 , \3752 , \3753 , \3754 , \3755 , \3756 , \3757 , \3758 ,
         \3759 , \3760 , \3761 , \3762 , \3763 , \3764 , \3765 , \3766 , \3767 , \3768 ,
         \3769 , \3770 , \3771 , \3772 , \3773 , \3774 , \3775 , \3776 , \3777 , \3778 ,
         \3779 , \3780 , \3781 , \3782 , \3783 , \3784 , \3785 , \3786 , \3787 , \3788 ,
         \3789 , \3790 , \3791 , \3792 , \3793 , \3794 , \3795 , \3796 , \3797 , \3798 ,
         \3799 , \3800 , \3801 , \3802 , \3803 , \3804 , \3805 , \3806 , \3807 , \3808 ,
         \3809 , \3810 , \3811 , \3812 , \3813 , \3814 , \3815 , \3816 , \3817 , \3818 ,
         \3819 , \3820 , \3821 , \3822 , \3823 , \3824 , \3825 , \3826 , \3827 , \3828 ,
         \3829 , \3830 , \3831 , \3832 , \3833 , \3834 , \3835 , \3836 , \3837 , \3838 ,
         \3839 , \3840 , \3841 , \3842 , \3843 , \3844 , \3845 , \3846 , \3847 , \3848 ,
         \3849 , \3850 , \3851 , \3852 , \3853 , \3854 , \3855 , \3856 , \3857 , \3858 ,
         \3859 , \3860 , \3861_nG5551 , \3862 , \3863 , \3864 , \3865 , \3866 , \3867 , \3868 ,
         \3869 , \3870 , \3871 , \3872 , \3873 , \3874 , \3875 , \3876 , \3877 , \3878 ,
         \3879 , \3880 , \3881 , \3882 , \3883 , \3884 , \3885 , \3886 , \3887 , \3888 ,
         \3889 , \3890 , \3891 , \3892 , \3893 , \3894 , \3895 , \3896 , \3897 , \3898 ,
         \3899 , \3900 , \3901 , \3902 , \3903 , \3904 , \3905 , \3906 , \3907 , \3908 ,
         \3909 , \3910 , \3911 , \3912 , \3913 , \3914 , \3915 , \3916 , \3917 , \3918 ,
         \3919 , \3920 , \3921 , \3922 , \3923 , \3924 , \3925 , \3926 , \3927 , \3928 ,
         \3929 , \3930 , \3931 , \3932 , \3933 , \3934 , \3935 , \3936 , \3937 , \3938 ,
         \3939 , \3940 , \3941 , \3942 , \3943 , \3944 , \3945 , \3946 , \3947 , \3948 ,
         \3949 , \3950 , \3951 , \3952 , \3953 , \3954 , \3955 , \3956 , \3957 , \3958 ,
         \3959 , \3960 , \3961 , \3962 , \3963 , \3964 , \3965 , \3966 , \3967 , \3968 ,
         \3969 , \3970 , \3971 , \3972 , \3973 , \3974 , \3975 , \3976 , \3977 , \3978 ,
         \3979 , \3980 , \3981 , \3982 , \3983 , \3984 , \3985 , \3986 , \3987 , \3988 ,
         \3989 , \3990 , \3991 , \3992 , \3993 , \3994 , \3995 , \3996 , \3997 , \3998 ,
         \3999 , \4000 , \4001 , \4002 , \4003 , \4004 , \4005 , \4006 , \4007 , \4008 ,
         \4009 , \4010 , \4011 , \4012 , \4013 , \4014 , \4015 , \4016 , \4017 , \4018 ,
         \4019 , \4020 , \4021 , \4022 , \4023 , \4024 , \4025 , \4026 , \4027 , \4028 ,
         \4029 , \4030 , \4031 , \4032 , \4033 , \4034 , \4035 , \4036 , \4037 , \4038 ,
         \4039 , \4040 , \4041 , \4042 , \4043 , \4044 , \4045 , \4046 , \4047 , \4048 ,
         \4049 , \4050 , \4051 , \4052 , \4053 , \4054 , \4055 , \4056 , \4057 , \4058 ,
         \4059_nG554f , \4060 , \4061 , \4062 , \4063 , \4064 , \4065 , \4066 , \4067 , \4068 ,
         \4069 , \4070 , \4071 , \4072 , \4073 , \4074 , \4075 , \4076 , \4077 , \4078 ,
         \4079 , \4080 , \4081 , \4082 , \4083 , \4084 , \4085 , \4086 , \4087 , \4088 ,
         \4089 , \4090 , \4091 , \4092 , \4093 , \4094 , \4095 , \4096 , \4097 , \4098 ,
         \4099 , \4100 , \4101 , \4102 , \4103 , \4104 , \4105 , \4106 , \4107 , \4108 ,
         \4109 , \4110 , \4111 , \4112 , \4113 , \4114 , \4115 , \4116 , \4117 , \4118 ,
         \4119 , \4120 , \4121 , \4122 , \4123 , \4124 , \4125 , \4126 , \4127 , \4128 ,
         \4129 , \4130 , \4131 , \4132 , \4133 , \4134 , \4135 , \4136 , \4137 , \4138 ,
         \4139 , \4140 , \4141 , \4142 , \4143 , \4144 , \4145 , \4146 , \4147 , \4148 ,
         \4149 , \4150 , \4151 , \4152 , \4153 , \4154 , \4155 , \4156 , \4157 , \4158 ,
         \4159 , \4160 , \4161 , \4162 , \4163 , \4164 , \4165 , \4166 , \4167 , \4168 ,
         \4169 , \4170 , \4171 , \4172 , \4173 , \4174 , \4175 , \4176 , \4177 , \4178 ,
         \4179 , \4180 , \4181 , \4182 , \4183 , \4184 , \4185 , \4186 , \4187 , \4188 ,
         \4189 , \4190 , \4191 , \4192 , \4193 , \4194 , \4195 , \4196 , \4197 , \4198 ,
         \4199 , \4200 , \4201 , \4202 , \4203 , \4204 , \4205 , \4206 , \4207 , \4208 ,
         \4209 , \4210 , \4211 , \4212 , \4213 , \4214 , \4215 , \4216 , \4217 , \4218 ,
         \4219 , \4220 , \4221 , \4222 , \4223 , \4224 , \4225 , \4226 , \4227 , \4228 ,
         \4229 , \4230 , \4231 , \4232 , \4233 , \4234 , \4235 , \4236 , \4237 , \4238 ,
         \4239 , \4240 , \4241 , \4242 , \4243 , \4244 , \4245 , \4246 , \4247 , \4248 ,
         \4249 , \4250 , \4251 , \4252 , \4253 , \4254 , \4255 , \4256 , \4257 , \4258 ,
         \4259 , \4260_nG554d , \4261 , \4262 , \4263 , \4264 , \4265 , \4266 , \4267 , \4268 ,
         \4269 , \4270 , \4271 , \4272 , \4273 , \4274 , \4275 , \4276 , \4277 , \4278 ,
         \4279 , \4280 , \4281 , \4282 , \4283 , \4284 , \4285 , \4286 , \4287 , \4288 ,
         \4289 , \4290 , \4291 , \4292 , \4293 , \4294 , \4295 , \4296 , \4297 , \4298 ,
         \4299 , \4300 , \4301 , \4302 , \4303 , \4304 , \4305 , \4306 , \4307 , \4308 ,
         \4309 , \4310 , \4311 , \4312 , \4313 , \4314 , \4315 , \4316 , \4317 , \4318 ,
         \4319 , \4320 , \4321 , \4322 , \4323 , \4324 , \4325 , \4326 , \4327 , \4328 ,
         \4329 , \4330 , \4331 , \4332 , \4333 , \4334 , \4335 , \4336 , \4337 , \4338 ,
         \4339 , \4340 , \4341 , \4342 , \4343 , \4344 , \4345 , \4346 , \4347 , \4348 ,
         \4349 , \4350 , \4351 , \4352 , \4353 , \4354 , \4355 , \4356 , \4357 , \4358 ,
         \4359 , \4360 , \4361 , \4362 , \4363 , \4364 , \4365 , \4366 , \4367 , \4368 ,
         \4369 , \4370 , \4371 , \4372 , \4373 , \4374 , \4375 , \4376 , \4377 , \4378 ,
         \4379 , \4380 , \4381 , \4382 , \4383 , \4384 , \4385 , \4386 , \4387 , \4388 ,
         \4389 , \4390 , \4391 , \4392 , \4393 , \4394 , \4395 , \4396 , \4397 , \4398 ,
         \4399 , \4400 , \4401 , \4402 , \4403 , \4404 , \4405 , \4406 , \4407 , \4408 ,
         \4409 , \4410 , \4411 , \4412 , \4413 , \4414 , \4415 , \4416 , \4417 , \4418 ,
         \4419 , \4420 , \4421 , \4422 , \4423 , \4424 , \4425 , \4426 , \4427 , \4428 ,
         \4429 , \4430 , \4431 , \4432 , \4433 , \4434 , \4435 , \4436 , \4437 , \4438 ,
         \4439 , \4440 , \4441 , \4442 , \4443 , \4444 , \4445 , \4446 , \4447 , \4448 ,
         \4449 , \4450 , \4451 , \4452 , \4453 , \4454 , \4455 , \4456 , \4457 , \4458 ,
         \4459 , \4460 , \4461 , \4462 , \4463 , \4464 , \4465 , \4466 , \4467 , \4468_nG554b ,
         \4469 , \4470 , \4471 , \4472 , \4473 , \4474 , \4475 , \4476 , \4477 , \4478 ,
         \4479 , \4480 , \4481 , \4482 , \4483 , \4484 , \4485 , \4486 , \4487 , \4488 ,
         \4489 , \4490 , \4491 , \4492 , \4493 , \4494 , \4495 , \4496 , \4497 , \4498 ,
         \4499 , \4500 , \4501 , \4502 , \4503 , \4504 , \4505 , \4506 , \4507 , \4508 ,
         \4509 , \4510 , \4511 , \4512 , \4513 , \4514 , \4515 , \4516 , \4517 , \4518 ,
         \4519 , \4520 , \4521 , \4522 , \4523 , \4524 , \4525 , \4526 , \4527 , \4528 ,
         \4529 , \4530 , \4531 , \4532 , \4533 , \4534 , \4535 , \4536 , \4537 , \4538 ,
         \4539 , \4540 , \4541 , \4542 , \4543 , \4544 , \4545 , \4546 , \4547 , \4548 ,
         \4549 , \4550 , \4551 , \4552 , \4553 , \4554 , \4555 , \4556 , \4557 , \4558 ,
         \4559 , \4560 , \4561 , \4562 , \4563 , \4564 , \4565 , \4566 , \4567 , \4568 ,
         \4569 , \4570 , \4571 , \4572 , \4573 , \4574 , \4575 , \4576 , \4577 , \4578 ,
         \4579 , \4580 , \4581 , \4582 , \4583 , \4584 , \4585 , \4586 , \4587 , \4588 ,
         \4589 , \4590 , \4591 , \4592 , \4593 , \4594 , \4595 , \4596 , \4597 , \4598 ,
         \4599 , \4600 , \4601 , \4602 , \4603 , \4604 , \4605 , \4606 , \4607 , \4608 ,
         \4609 , \4610 , \4611 , \4612 , \4613 , \4614 , \4615 , \4616 , \4617 , \4618 ,
         \4619 , \4620 , \4621 , \4622 , \4623 , \4624 , \4625 , \4626 , \4627 , \4628 ,
         \4629 , \4630 , \4631 , \4632 , \4633 , \4634 , \4635 , \4636 , \4637 , \4638 ,
         \4639 , \4640 , \4641 , \4642 , \4643 , \4644 , \4645 , \4646 , \4647 , \4648 ,
         \4649 , \4650 , \4651 , \4652 , \4653 , \4654 , \4655 , \4656 , \4657 , \4658 ,
         \4659 , \4660 , \4661 , \4662 , \4663 , \4664 , \4665 , \4666 , \4667 , \4668 ,
         \4669 , \4670 , \4671 , \4672 , \4673 , \4674 , \4675 , \4676 , \4677 , \4678 ,
         \4679_nG5549 , \4680 , \4681 , \4682 , \4683 , \4684 , \4685 , \4686 , \4687 , \4688 ,
         \4689 , \4690 , \4691 , \4692 , \4693 , \4694 , \4695 , \4696 , \4697 , \4698 ,
         \4699 , \4700 , \4701 , \4702 , \4703 , \4704 , \4705 , \4706 , \4707 , \4708 ,
         \4709 , \4710 , \4711 , \4712 , \4713 , \4714 , \4715 , \4716 , \4717 , \4718 ,
         \4719 , \4720 , \4721 , \4722 , \4723 , \4724 , \4725 , \4726 , \4727 , \4728 ,
         \4729 , \4730 , \4731 , \4732 , \4733 , \4734 , \4735 , \4736 , \4737 , \4738 ,
         \4739 , \4740 , \4741 , \4742 , \4743 , \4744 , \4745 , \4746 , \4747 , \4748 ,
         \4749 , \4750 , \4751 , \4752 , \4753 , \4754 , \4755 , \4756 , \4757 , \4758 ,
         \4759 , \4760 , \4761 , \4762 , \4763 , \4764 , \4765 , \4766 , \4767 , \4768 ,
         \4769 , \4770 , \4771 , \4772 , \4773 , \4774 , \4775 , \4776 , \4777 , \4778 ,
         \4779 , \4780 , \4781 , \4782 , \4783 , \4784 , \4785 , \4786 , \4787 , \4788 ,
         \4789 , \4790 , \4791 , \4792 , \4793 , \4794 , \4795 , \4796 , \4797 , \4798 ,
         \4799 , \4800 , \4801 , \4802 , \4803 , \4804 , \4805 , \4806 , \4807 , \4808 ,
         \4809 , \4810 , \4811 , \4812 , \4813 , \4814 , \4815 , \4816 , \4817 , \4818 ,
         \4819 , \4820 , \4821 , \4822 , \4823 , \4824 , \4825 , \4826 , \4827 , \4828 ,
         \4829 , \4830 , \4831 , \4832 , \4833 , \4834 , \4835 , \4836 , \4837 , \4838 ,
         \4839 , \4840 , \4841 , \4842 , \4843 , \4844 , \4845 , \4846 , \4847 , \4848 ,
         \4849 , \4850 , \4851 , \4852 , \4853 , \4854 , \4855 , \4856 , \4857 , \4858 ,
         \4859 , \4860 , \4861 , \4862 , \4863 , \4864 , \4865 , \4866 , \4867 , \4868 ,
         \4869 , \4870 , \4871 , \4872 , \4873 , \4874 , \4875 , \4876 , \4877 , \4878 ,
         \4879 , \4880 , \4881 , \4882 , \4883 , \4884 , \4885 , \4886 , \4887 , \4888 ,
         \4889 , \4890 , \4891 , \4892 , \4893 , \4894 , \4895 , \4896 , \4897_nG5547 , \4898 ,
         \4899 , \4900 , \4901 , \4902 , \4903 , \4904 , \4905 , \4906 , \4907 , \4908 ,
         \4909 , \4910 , \4911 , \4912 , \4913 , \4914 , \4915 , \4916 , \4917 , \4918 ,
         \4919 , \4920 , \4921 , \4922 , \4923 , \4924 , \4925 , \4926 , \4927 , \4928 ,
         \4929 , \4930 , \4931 , \4932 , \4933 , \4934 , \4935 , \4936 , \4937 , \4938 ,
         \4939 , \4940 , \4941 , \4942 , \4943 , \4944 , \4945 , \4946 , \4947 , \4948 ,
         \4949 , \4950 , \4951 , \4952 , \4953 , \4954 , \4955 , \4956 , \4957 , \4958 ,
         \4959 , \4960 , \4961 , \4962 , \4963 , \4964 , \4965 , \4966 , \4967 , \4968 ,
         \4969 , \4970 , \4971 , \4972 , \4973 , \4974 , \4975 , \4976 , \4977 , \4978 ,
         \4979 , \4980 , \4981 , \4982 , \4983 , \4984 , \4985 , \4986 , \4987 , \4988 ,
         \4989 , \4990 , \4991 , \4992 , \4993 , \4994 , \4995 , \4996 , \4997 , \4998 ,
         \4999 , \5000 , \5001 , \5002 , \5003 , \5004 , \5005 , \5006 , \5007 , \5008 ,
         \5009 , \5010 , \5011 , \5012 , \5013 , \5014 , \5015 , \5016 , \5017 , \5018 ,
         \5019 , \5020 , \5021 , \5022 , \5023 , \5024 , \5025 , \5026 , \5027 , \5028 ,
         \5029 , \5030 , \5031 , \5032 , \5033 , \5034 , \5035 , \5036 , \5037 , \5038 ,
         \5039 , \5040 , \5041 , \5042 , \5043 , \5044 , \5045 , \5046 , \5047 , \5048 ,
         \5049 , \5050 , \5051 , \5052 , \5053 , \5054 , \5055 , \5056 , \5057 , \5058 ,
         \5059 , \5060 , \5061 , \5062 , \5063 , \5064 , \5065 , \5066 , \5067 , \5068 ,
         \5069 , \5070 , \5071 , \5072 , \5073 , \5074 , \5075 , \5076 , \5077 , \5078 ,
         \5079 , \5080 , \5081 , \5082 , \5083 , \5084 , \5085 , \5086 , \5087 , \5088 ,
         \5089 , \5090 , \5091 , \5092 , \5093 , \5094 , \5095 , \5096 , \5097 , \5098 ,
         \5099 , \5100 , \5101 , \5102 , \5103 , \5104 , \5105 , \5106 , \5107 , \5108 ,
         \5109 , \5110 , \5111 , \5112 , \5113 , \5114 , \5115 , \5116 , \5117_nG5545 , \5118 ,
         \5119 , \5120 , \5121 , \5122 , \5123 , \5124 , \5125 , \5126 , \5127 , \5128 ,
         \5129 , \5130 , \5131 , \5132 , \5133 , \5134 , \5135 , \5136 , \5137 , \5138 ,
         \5139 , \5140 , \5141 , \5142 , \5143 , \5144 , \5145 , \5146 , \5147 , \5148 ,
         \5149 , \5150 , \5151 , \5152 , \5153 , \5154 , \5155 , \5156 , \5157 , \5158 ,
         \5159 , \5160 , \5161 , \5162 , \5163 , \5164 , \5165 , \5166 , \5167 , \5168 ,
         \5169 , \5170 , \5171 , \5172 , \5173 , \5174 , \5175 , \5176 , \5177 , \5178 ,
         \5179 , \5180 , \5181 , \5182 , \5183 , \5184 , \5185 , \5186 , \5187 , \5188 ,
         \5189 , \5190 , \5191 , \5192 , \5193 , \5194 , \5195 , \5196 , \5197 , \5198 ,
         \5199 , \5200 , \5201 , \5202 , \5203 , \5204 , \5205 , \5206 , \5207 , \5208 ,
         \5209 , \5210 , \5211 , \5212 , \5213 , \5214 , \5215 , \5216 , \5217 , \5218 ,
         \5219 , \5220 , \5221 , \5222 , \5223 , \5224 , \5225 , \5226 , \5227 , \5228 ,
         \5229 , \5230 , \5231 , \5232 , \5233 , \5234 , \5235 , \5236 , \5237 , \5238 ,
         \5239 , \5240 , \5241 , \5242 , \5243 , \5244 , \5245 , \5246 , \5247 , \5248 ,
         \5249 , \5250 , \5251 , \5252 , \5253 , \5254 , \5255 , \5256 , \5257 , \5258 ,
         \5259 , \5260 , \5261 , \5262 , \5263 , \5264 , \5265 , \5266 , \5267 , \5268 ,
         \5269 , \5270 , \5271 , \5272 , \5273 , \5274 , \5275 , \5276 , \5277 , \5278 ,
         \5279 , \5280 , \5281 , \5282 , \5283 , \5284 , \5285 , \5286 , \5287 , \5288 ,
         \5289 , \5290 , \5291 , \5292 , \5293 , \5294 , \5295 , \5296 , \5297 , \5298 ,
         \5299 , \5300 , \5301 , \5302 , \5303 , \5304 , \5305 , \5306 , \5307 , \5308 ,
         \5309 , \5310 , \5311 , \5312 , \5313 , \5314 , \5315 , \5316 , \5317 , \5318 ,
         \5319 , \5320 , \5321 , \5322 , \5323 , \5324 , \5325 , \5326 , \5327 , \5328 ,
         \5329 , \5330 , \5331 , \5332 , \5333 , \5334 , \5335 , \5336 , \5337 , \5338 ,
         \5339 , \5340 , \5341 , \5342 , \5343 , \5344 , \5345 , \5346 , \5347 , \5348_nG5543 ,
         \5349 , \5350 , \5351 , \5352 , \5353 , \5354 , \5355 , \5356 , \5357 , \5358 ,
         \5359 , \5360 , \5361 , \5362 , \5363 , \5364 , \5365 , \5366 , \5367 , \5368 ,
         \5369 , \5370 , \5371 , \5372 , \5373 , \5374 , \5375 , \5376 , \5377 , \5378 ,
         \5379 , \5380 , \5381 , \5382 , \5383 , \5384 , \5385 , \5386 , \5387 , \5388 ,
         \5389 , \5390 , \5391 , \5392 , \5393 , \5394 , \5395 , \5396 , \5397 , \5398 ,
         \5399 , \5400 , \5401 , \5402 , \5403 , \5404 , \5405 , \5406 , \5407 , \5408 ,
         \5409 , \5410 , \5411 , \5412 , \5413 , \5414 , \5415 , \5416 , \5417 , \5418 ,
         \5419 , \5420 , \5421 , \5422 , \5423 , \5424 , \5425 , \5426 , \5427 , \5428 ,
         \5429 , \5430 , \5431 , \5432 , \5433 , \5434 , \5435 , \5436 , \5437 , \5438 ,
         \5439 , \5440 , \5441 , \5442 , \5443 , \5444 , \5445 , \5446 , \5447 , \5448 ,
         \5449 , \5450 , \5451 , \5452 , \5453 , \5454 , \5455 , \5456 , \5457 , \5458 ,
         \5459 , \5460 , \5461 , \5462 , \5463 , \5464 , \5465 , \5466 , \5467 , \5468 ,
         \5469 , \5470 , \5471 , \5472 , \5473 , \5474 , \5475 , \5476 , \5477 , \5478 ,
         \5479 , \5480 , \5481 , \5482 , \5483 , \5484 , \5485 , \5486 , \5487 , \5488 ,
         \5489 , \5490 , \5491 , \5492 , \5493 , \5494 , \5495 , \5496 , \5497 , \5498 ,
         \5499 , \5500 , \5501 , \5502 , \5503 , \5504 , \5505 , \5506 , \5507 , \5508 ,
         \5509 , \5510 , \5511 , \5512 , \5513 , \5514 , \5515 , \5516 , \5517 , \5518 ,
         \5519 , \5520 , \5521 , \5522 , \5523 , \5524 , \5525 , \5526 , \5527 , \5528 ,
         \5529 , \5530 , \5531 , \5532 , \5533 , \5534 , \5535 , \5536 , \5537 , \5538 ,
         \5539 , \5540 , \5541 , \5542 , \5543 , \5544 , \5545 , \5546 , \5547 , \5548 ,
         \5549 , \5550 , \5551 , \5552 , \5553 , \5554 , \5555 , \5556 , \5557 , \5558 ,
         \5559 , \5560 , \5561 , \5562 , \5563 , \5564 , \5565 , \5566 , \5567 , \5568 ,
         \5569 , \5570 , \5571 , \5572 , \5573 , \5574 , \5575 , \5576 , \5577 , \5578 ,
         \5579_nG5541 , \5580 , \5581 , \5582 , \5583 , \5584 , \5585 , \5586 , \5587 , \5588 ,
         \5589 , \5590 , \5591 , \5592 , \5593 , \5594 , \5595 , \5596 , \5597 , \5598 ,
         \5599 , \5600 , \5601 , \5602 , \5603 , \5604 , \5605 , \5606 , \5607 , \5608 ,
         \5609 , \5610 , \5611 , \5612 , \5613 , \5614 , \5615 , \5616 , \5617 , \5618 ,
         \5619 , \5620 , \5621 , \5622 , \5623 , \5624 , \5625 , \5626 , \5627 , \5628 ,
         \5629 , \5630 , \5631 , \5632 , \5633 , \5634 , \5635 , \5636 , \5637 , \5638 ,
         \5639 , \5640 , \5641 , \5642 , \5643 , \5644 , \5645 , \5646 , \5647 , \5648 ,
         \5649 , \5650 , \5651 , \5652 , \5653 , \5654 , \5655 , \5656 , \5657 , \5658 ,
         \5659 , \5660 , \5661 , \5662 , \5663 , \5664 , \5665 , \5666 , \5667 , \5668 ,
         \5669 , \5670 , \5671 , \5672 , \5673 , \5674 , \5675 , \5676 , \5677 , \5678 ,
         \5679 , \5680 , \5681 , \5682 , \5683 , \5684 , \5685 , \5686 , \5687 , \5688 ,
         \5689 , \5690 , \5691 , \5692 , \5693 , \5694 , \5695 , \5696 , \5697 , \5698 ,
         \5699 , \5700 , \5701 , \5702 , \5703 , \5704 , \5705 , \5706 , \5707 , \5708 ,
         \5709 , \5710 , \5711 , \5712 , \5713 , \5714 , \5715 , \5716 , \5717 , \5718 ,
         \5719 , \5720 , \5721 , \5722 , \5723 , \5724 , \5725 , \5726 , \5727 , \5728 ,
         \5729 , \5730 , \5731 , \5732 , \5733 , \5734 , \5735 , \5736 , \5737 , \5738 ,
         \5739 , \5740 , \5741 , \5742 , \5743 , \5744 , \5745 , \5746 , \5747 , \5748 ,
         \5749 , \5750 , \5751 , \5752 , \5753 , \5754 , \5755 , \5756 , \5757 , \5758 ,
         \5759 , \5760 , \5761 , \5762 , \5763 , \5764 , \5765 , \5766 , \5767 , \5768 ,
         \5769 , \5770 , \5771 , \5772 , \5773 , \5774 , \5775 , \5776 , \5777 , \5778 ,
         \5779 , \5780 , \5781 , \5782 , \5783 , \5784 , \5785 , \5786 , \5787 , \5788 ,
         \5789 , \5790 , \5791 , \5792 , \5793 , \5794 , \5795 , \5796 , \5797 , \5798 ,
         \5799 , \5800 , \5801 , \5802 , \5803 , \5804 , \5805 , \5806 , \5807 , \5808 ,
         \5809 , \5810 , \5811 , \5812 , \5813 , \5814 , \5815 , \5816 , \5817_nG553f , \5818 ,
         \5819 , \5820 , \5821 , \5822 , \5823 , \5824 , \5825 , \5826 , \5827 , \5828 ,
         \5829 , \5830 , \5831 , \5832 , \5833 , \5834 , \5835 , \5836 , \5837 , \5838 ,
         \5839 , \5840 , \5841 , \5842 , \5843 , \5844 , \5845 , \5846 , \5847 , \5848 ,
         \5849 , \5850 , \5851 , \5852 , \5853 , \5854 , \5855 , \5856 , \5857 , \5858 ,
         \5859 , \5860 , \5861 , \5862 , \5863 , \5864 , \5865 , \5866 , \5867 , \5868 ,
         \5869 , \5870 , \5871 , \5872 , \5873 , \5874 , \5875 , \5876 , \5877 , \5878 ,
         \5879 , \5880 , \5881 , \5882 , \5883 , \5884 , \5885 , \5886 , \5887 , \5888 ,
         \5889 , \5890 , \5891 , \5892 , \5893 , \5894 , \5895 , \5896 , \5897 , \5898 ,
         \5899 , \5900 , \5901 , \5902 , \5903 , \5904 , \5905 , \5906 , \5907 , \5908 ,
         \5909 , \5910 , \5911 , \5912 , \5913 , \5914 , \5915 , \5916 , \5917 , \5918 ,
         \5919 , \5920 , \5921 , \5922 , \5923 , \5924 , \5925 , \5926 , \5927 , \5928 ,
         \5929 , \5930 , \5931 , \5932 , \5933 , \5934 , \5935 , \5936 , \5937 , \5938 ,
         \5939 , \5940 , \5941 , \5942 , \5943 , \5944 , \5945 , \5946 , \5947 , \5948 ,
         \5949 , \5950 , \5951 , \5952 , \5953 , \5954 , \5955 , \5956 , \5957 , \5958 ,
         \5959 , \5960 , \5961 , \5962 , \5963 , \5964 , \5965 , \5966 , \5967 , \5968 ,
         \5969 , \5970 , \5971 , \5972 , \5973 , \5974 , \5975 , \5976 , \5977 , \5978 ,
         \5979 , \5980 , \5981 , \5982 , \5983 , \5984 , \5985 , \5986 , \5987 , \5988 ,
         \5989 , \5990 , \5991 , \5992 , \5993 , \5994 , \5995 , \5996 , \5997 , \5998 ,
         \5999 , \6000 , \6001 , \6002 , \6003 , \6004 , \6005 , \6006 , \6007 , \6008 ,
         \6009 , \6010 , \6011 , \6012 , \6013 , \6014 , \6015 , \6016 , \6017 , \6018 ,
         \6019 , \6020 , \6021 , \6022 , \6023 , \6024 , \6025 , \6026 , \6027 , \6028 ,
         \6029 , \6030 , \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 , \6038 ,
         \6039 , \6040 , \6041 , \6042 , \6043 , \6044 , \6045 , \6046 , \6047 , \6048 ,
         \6049 , \6050 , \6051 , \6052 , \6053 , \6054 , \6055 , \6056 , \6057 , \6058_nG553d ,
         \6059 , \6060 , \6061 , \6062 , \6063 , \6064 , \6065 , \6066 , \6067 , \6068 ,
         \6069 , \6070 , \6071 , \6072 , \6073 , \6074 , \6075 , \6076 , \6077 , \6078 ,
         \6079 , \6080 , \6081 , \6082 , \6083 , \6084 , \6085 , \6086 , \6087 , \6088 ,
         \6089 , \6090 , \6091 , \6092 , \6093 , \6094 , \6095 , \6096 , \6097 , \6098 ,
         \6099 , \6100 , \6101 , \6102 , \6103 , \6104 , \6105 , \6106 , \6107 , \6108 ,
         \6109 , \6110 , \6111 , \6112 , \6113 , \6114 , \6115 , \6116 , \6117 , \6118 ,
         \6119 , \6120 , \6121 , \6122 , \6123 , \6124 , \6125 , \6126 , \6127 , \6128 ,
         \6129 , \6130 , \6131 , \6132 , \6133 , \6134 , \6135 , \6136 , \6137 , \6138 ,
         \6139 , \6140 , \6141 , \6142 , \6143 , \6144 , \6145 , \6146 , \6147 , \6148 ,
         \6149 , \6150 , \6151 , \6152 , \6153 , \6154 , \6155 , \6156 , \6157 , \6158 ,
         \6159 , \6160 , \6161 , \6162 , \6163 , \6164 , \6165 , \6166 , \6167 , \6168 ,
         \6169 , \6170 , \6171 , \6172 , \6173 , \6174 , \6175 , \6176 , \6177 , \6178 ,
         \6179 , \6180 , \6181 , \6182 , \6183 , \6184 , \6185 , \6186 , \6187 , \6188 ,
         \6189 , \6190 , \6191 , \6192 , \6193 , \6194 , \6195 , \6196 , \6197 , \6198 ,
         \6199 , \6200 , \6201 , \6202 , \6203 , \6204 , \6205 , \6206 , \6207 , \6208 ,
         \6209 , \6210 , \6211 , \6212 , \6213 , \6214 , \6215 , \6216 , \6217 , \6218 ,
         \6219 , \6220 , \6221 , \6222 , \6223 , \6224 , \6225 , \6226 , \6227 , \6228 ,
         \6229 , \6230 , \6231 , \6232 , \6233 , \6234 , \6235 , \6236 , \6237 , \6238 ,
         \6239 , \6240 , \6241 , \6242 , \6243 , \6244 , \6245 , \6246 , \6247 , \6248 ,
         \6249 , \6250 , \6251 , \6252 , \6253 , \6254 , \6255 , \6256 , \6257 , \6258 ,
         \6259 , \6260 , \6261 , \6262 , \6263 , \6264 , \6265 , \6266 , \6267 , \6268 ,
         \6269 , \6270 , \6271 , \6272 , \6273 , \6274 , \6275 , \6276 , \6277 , \6278 ,
         \6279 , \6280 , \6281 , \6282 , \6283 , \6284 , \6285 , \6286 , \6287 , \6288 ,
         \6289 , \6290 , \6291 , \6292 , \6293 , \6294 , \6295 , \6296 , \6297 , \6298 ,
         \6299 , \6300 , \6301 , \6302 , \6303 , \6304 , \6305 , \6306_nG553b , \6307 , \6308 ,
         \6309 , \6310 , \6311 , \6312 , \6313 , \6314 , \6315 , \6316 , \6317 , \6318 ,
         \6319 , \6320 , \6321 , \6322 , \6323 , \6324 , \6325 , \6326 , \6327 , \6328 ,
         \6329 , \6330 , \6331 , \6332 , \6333 , \6334 , \6335 , \6336 , \6337 , \6338 ,
         \6339 , \6340 , \6341 , \6342 , \6343 , \6344 , \6345 , \6346 , \6347 , \6348 ,
         \6349 , \6350 , \6351 , \6352 , \6353 , \6354 , \6355 , \6356 , \6357 , \6358 ,
         \6359 , \6360 , \6361 , \6362 , \6363 , \6364 , \6365 , \6366 , \6367 , \6368 ,
         \6369 , \6370 , \6371 , \6372 , \6373 , \6374 , \6375 , \6376 , \6377 , \6378 ,
         \6379 , \6380 , \6381 , \6382 , \6383 , \6384 , \6385 , \6386 , \6387 , \6388 ,
         \6389 , \6390 , \6391 , \6392 , \6393 , \6394 , \6395 , \6396 , \6397 , \6398 ,
         \6399 , \6400 , \6401 , \6402 , \6403 , \6404 , \6405 , \6406 , \6407 , \6408 ,
         \6409 , \6410 , \6411 , \6412 , \6413 , \6414 , \6415 , \6416 , \6417 , \6418 ,
         \6419 , \6420 , \6421 , \6422 , \6423 , \6424 , \6425 , \6426 , \6427 , \6428 ,
         \6429 , \6430 , \6431 , \6432 , \6433 , \6434 , \6435 , \6436 , \6437 , \6438 ,
         \6439 , \6440 , \6441 , \6442 , \6443 , \6444 , \6445 , \6446 , \6447 , \6448 ,
         \6449 , \6450 , \6451 , \6452 , \6453 , \6454 , \6455 , \6456 , \6457 , \6458 ,
         \6459 , \6460 , \6461 , \6462 , \6463 , \6464 , \6465 , \6466 , \6467 , \6468 ,
         \6469 , \6470 , \6471 , \6472 , \6473 , \6474 , \6475 , \6476 , \6477 , \6478 ,
         \6479 , \6480 , \6481 , \6482 , \6483 , \6484 , \6485 , \6486 , \6487 , \6488 ,
         \6489 , \6490 , \6491 , \6492 , \6493 , \6494 , \6495 , \6496 , \6497 , \6498 ,
         \6499 , \6500 , \6501 , \6502 , \6503 , \6504 , \6505 , \6506 , \6507 , \6508 ,
         \6509 , \6510 , \6511 , \6512 , \6513 , \6514 , \6515 , \6516 , \6517 , \6518 ,
         \6519 , \6520 , \6521 , \6522 , \6523 , \6524 , \6525 , \6526 , \6527 , \6528 ,
         \6529 , \6530 , \6531 , \6532 , \6533 , \6534 , \6535 , \6536 , \6537 , \6538 ,
         \6539 , \6540 , \6541 , \6542 , \6543 , \6544 , \6545 , \6546 , \6547 , \6548 ,
         \6549 , \6550 , \6551 , \6552 , \6553 , \6554 , \6555 , \6556 , \6557_nG5539 , \6558 ,
         \6559 , \6560 , \6561 , \6562 , \6563 , \6564 , \6565 , \6566 , \6567 , \6568 ,
         \6569 , \6570 , \6571 , \6572 , \6573 , \6574 , \6575 , \6576 , \6577 , \6578 ,
         \6579 , \6580 , \6581 , \6582 , \6583 , \6584 , \6585 , \6586 , \6587 , \6588 ,
         \6589 , \6590 , \6591 , \6592 , \6593 , \6594 , \6595 , \6596 , \6597 , \6598 ,
         \6599 , \6600 , \6601 , \6602 , \6603 , \6604 , \6605 , \6606 , \6607 , \6608 ,
         \6609 , \6610 , \6611 , \6612 , \6613 , \6614 , \6615 , \6616 , \6617 , \6618 ,
         \6619 , \6620 , \6621 , \6622 , \6623 , \6624 , \6625 , \6626 , \6627 , \6628 ,
         \6629 , \6630 , \6631 , \6632 , \6633 , \6634 , \6635 , \6636 , \6637 , \6638 ,
         \6639 , \6640 , \6641 , \6642 , \6643 , \6644 , \6645 , \6646 , \6647 , \6648 ,
         \6649 , \6650 , \6651 , \6652 , \6653 , \6654 , \6655 , \6656 , \6657 , \6658 ,
         \6659 , \6660 , \6661 , \6662 , \6663 , \6664 , \6665 , \6666 , \6667 , \6668 ,
         \6669 , \6670 , \6671 , \6672 , \6673 , \6674 , \6675 , \6676 , \6677 , \6678 ,
         \6679 , \6680 , \6681 , \6682 , \6683 , \6684 , \6685 , \6686 , \6687 , \6688 ,
         \6689 , \6690 , \6691 , \6692 , \6693 , \6694 , \6695 , \6696 , \6697 , \6698 ,
         \6699 , \6700 , \6701 , \6702 , \6703 , \6704 , \6705 , \6706 , \6707 , \6708 ,
         \6709 , \6710 , \6711 , \6712 , \6713 , \6714 , \6715 , \6716 , \6717 , \6718 ,
         \6719 , \6720 , \6721 , \6722 , \6723 , \6724 , \6725 , \6726 , \6727 , \6728 ,
         \6729 , \6730 , \6731 , \6732 , \6733 , \6734 , \6735 , \6736 , \6737 , \6738 ,
         \6739 , \6740 , \6741 , \6742 , \6743 , \6744 , \6745 , \6746 , \6747 , \6748 ,
         \6749 , \6750 , \6751 , \6752 , \6753 , \6754 , \6755 , \6756 , \6757 , \6758 ,
         \6759 , \6760 , \6761 , \6762 , \6763 , \6764 , \6765 , \6766 , \6767 , \6768 ,
         \6769 , \6770 , \6771 , \6772 , \6773 , \6774 , \6775 , \6776 , \6777 , \6778 ,
         \6779 , \6780 , \6781 , \6782 , \6783 , \6784 , \6785 , \6786 , \6787 , \6788 ,
         \6789 , \6790 , \6791 , \6792 , \6793 , \6794 , \6795 , \6796 , \6797 , \6798 ,
         \6799 , \6800 , \6801 , \6802 , \6803 , \6804 , \6805 , \6806 , \6807 , \6808 ,
         \6809 , \6810 , \6811 , \6812 , \6813 , \6814 , \6815_nG5537 , \6816 , \6817 , \6818 ,
         \6819 , \6820 , \6821 , \6822 , \6823 , \6824 , \6825 , \6826 , \6827 , \6828 ,
         \6829 , \6830 , \6831 , \6832 , \6833 , \6834 , \6835 , \6836 , \6837 , \6838 ,
         \6839 , \6840 , \6841 , \6842 , \6843 , \6844 , \6845 , \6846 , \6847 , \6848 ,
         \6849 , \6850 , \6851 , \6852 , \6853 , \6854 , \6855 , \6856 , \6857 , \6858 ,
         \6859 , \6860 , \6861 , \6862 , \6863 , \6864 , \6865 , \6866 , \6867 , \6868 ,
         \6869 , \6870 , \6871 , \6872 , \6873 , \6874 , \6875 , \6876 , \6877 , \6878 ,
         \6879 , \6880 , \6881 , \6882 , \6883 , \6884 , \6885 , \6886 , \6887 , \6888 ,
         \6889 , \6890 , \6891 , \6892 , \6893 , \6894 , \6895 , \6896 , \6897 , \6898 ,
         \6899 , \6900 , \6901 , \6902 , \6903 , \6904 , \6905 , \6906 , \6907 , \6908 ,
         \6909 , \6910 , \6911 , \6912 , \6913 , \6914 , \6915 , \6916 , \6917 , \6918 ,
         \6919 , \6920 , \6921 , \6922 , \6923 , \6924 , \6925 , \6926 , \6927 , \6928 ,
         \6929 , \6930 , \6931 , \6932 , \6933 , \6934 , \6935 , \6936 , \6937 , \6938 ,
         \6939 , \6940 , \6941 , \6942 , \6943 , \6944 , \6945 , \6946 , \6947 , \6948 ,
         \6949 , \6950 , \6951 , \6952 , \6953 , \6954 , \6955 , \6956 , \6957 , \6958 ,
         \6959 , \6960 , \6961 , \6962 , \6963 , \6964 , \6965 , \6966 , \6967 , \6968 ,
         \6969 , \6970 , \6971 , \6972 , \6973 , \6974 , \6975 , \6976 , \6977 , \6978 ,
         \6979 , \6980 , \6981 , \6982 , \6983 , \6984 , \6985 , \6986 , \6987 , \6988 ,
         \6989 , \6990 , \6991 , \6992 , \6993 , \6994 , \6995 , \6996 , \6997 , \6998 ,
         \6999 , \7000 , \7001 , \7002 , \7003 , \7004 , \7005 , \7006 , \7007 , \7008 ,
         \7009 , \7010 , \7011 , \7012 , \7013 , \7014 , \7015 , \7016 , \7017 , \7018 ,
         \7019 , \7020 , \7021 , \7022 , \7023 , \7024 , \7025 , \7026 , \7027 , \7028 ,
         \7029 , \7030 , \7031 , \7032 , \7033 , \7034 , \7035 , \7036 , \7037 , \7038 ,
         \7039 , \7040 , \7041 , \7042 , \7043 , \7044 , \7045 , \7046 , \7047 , \7048 ,
         \7049 , \7050 , \7051 , \7052 , \7053 , \7054 , \7055 , \7056 , \7057 , \7058 ,
         \7059 , \7060 , \7061 , \7062 , \7063 , \7064 , \7065 , \7066 , \7067 , \7068 ,
         \7069 , \7070 , \7071 , \7072 , \7073 , \7074 , \7075 , \7076_nG5535 , \7077 , \7078 ,
         \7079 , \7080 , \7081 , \7082 , \7083 , \7084 , \7085 , \7086 , \7087 , \7088 ,
         \7089 , \7090 , \7091 , \7092 , \7093 , \7094 , \7095 , \7096 , \7097 , \7098 ,
         \7099 , \7100 , \7101 , \7102 , \7103 , \7104 , \7105 , \7106 , \7107 , \7108 ,
         \7109 , \7110 , \7111 , \7112 , \7113 , \7114 , \7115 , \7116 , \7117 , \7118 ,
         \7119 , \7120 , \7121 , \7122 , \7123 , \7124 , \7125 , \7126 , \7127 , \7128 ,
         \7129 , \7130 , \7131 , \7132 , \7133 , \7134 , \7135 , \7136 , \7137 , \7138 ,
         \7139 , \7140 , \7141 , \7142 , \7143 , \7144 , \7145 , \7146 , \7147 , \7148 ,
         \7149 , \7150 , \7151 , \7152 , \7153 , \7154 , \7155 , \7156 , \7157 , \7158 ,
         \7159 , \7160 , \7161 , \7162 , \7163 , \7164 , \7165 , \7166 , \7167 , \7168 ,
         \7169 , \7170 , \7171 , \7172 , \7173 , \7174 , \7175 , \7176 , \7177 , \7178 ,
         \7179 , \7180 , \7181 , \7182 , \7183 , \7184 , \7185 , \7186 , \7187 , \7188 ,
         \7189 , \7190 , \7191 , \7192 , \7193 , \7194 , \7195 , \7196 , \7197 , \7198 ,
         \7199 , \7200 , \7201 , \7202 , \7203 , \7204 , \7205 , \7206 , \7207 , \7208 ,
         \7209 , \7210 , \7211 , \7212 , \7213 , \7214 , \7215 , \7216 , \7217 , \7218 ,
         \7219 , \7220 , \7221 , \7222 , \7223 , \7224 , \7225 , \7226 , \7227 , \7228 ,
         \7229 , \7230 , \7231 , \7232 , \7233 , \7234 , \7235 , \7236 , \7237 , \7238 ,
         \7239 , \7240 , \7241 , \7242 , \7243 , \7244 , \7245 , \7246 , \7247 , \7248 ,
         \7249 , \7250 , \7251 , \7252 , \7253 , \7254 , \7255 , \7256 , \7257 , \7258 ,
         \7259 , \7260 , \7261 , \7262 , \7263 , \7264 , \7265 , \7266 , \7267 , \7268 ,
         \7269 , \7270 , \7271 , \7272 , \7273 , \7274 , \7275 , \7276 , \7277 , \7278 ,
         \7279 , \7280 , \7281 , \7282 , \7283 , \7284 , \7285 , \7286 , \7287 , \7288 ,
         \7289 , \7290 , \7291 , \7292 , \7293 , \7294 , \7295 , \7296 , \7297 , \7298 ,
         \7299 , \7300 , \7301 , \7302 , \7303 , \7304 , \7305 , \7306 , \7307 , \7308 ,
         \7309 , \7310 , \7311 , \7312 , \7313 , \7314 , \7315 , \7316 , \7317 , \7318 ,
         \7319 , \7320 , \7321 , \7322 , \7323 , \7324 , \7325 , \7326 , \7327 , \7328 ,
         \7329 , \7330 , \7331 , \7332 , \7333 , \7334 , \7335 , \7336 , \7337 , \7338 ,
         \7339 , \7340 , \7341 , \7342 , \7343 , \7344_nG5533 , \7345 , \7346 , \7347 , \7348 ,
         \7349 , \7350 , \7351 , \7352 , \7353 , \7354 , \7355 , \7356 , \7357 , \7358 ,
         \7359 , \7360 , \7361 , \7362 , \7363 , \7364 , \7365 , \7366 , \7367 , \7368 ,
         \7369 , \7370 , \7371 , \7372 , \7373 , \7374 , \7375 , \7376 , \7377 , \7378 ,
         \7379 , \7380 , \7381 , \7382 , \7383 , \7384 , \7385 , \7386 , \7387 , \7388 ,
         \7389 , \7390 , \7391 , \7392 , \7393 , \7394 , \7395 , \7396 , \7397 , \7398 ,
         \7399 , \7400 , \7401 , \7402 , \7403 , \7404 , \7405 , \7406 , \7407 , \7408 ,
         \7409 , \7410 , \7411 , \7412 , \7413 , \7414 , \7415 , \7416 , \7417 , \7418 ,
         \7419 , \7420 , \7421 , \7422 , \7423 , \7424 , \7425 , \7426 , \7427 , \7428 ,
         \7429 , \7430 , \7431 , \7432 , \7433 , \7434 , \7435 , \7436 , \7437 , \7438 ,
         \7439 , \7440 , \7441 , \7442 , \7443 , \7444 , \7445 , \7446 , \7447 , \7448 ,
         \7449 , \7450 , \7451 , \7452 , \7453 , \7454 , \7455 , \7456 , \7457 , \7458 ,
         \7459 , \7460 , \7461 , \7462 , \7463 , \7464 , \7465 , \7466 , \7467 , \7468 ,
         \7469 , \7470 , \7471 , \7472 , \7473 , \7474 , \7475 , \7476 , \7477 , \7478 ,
         \7479 , \7480 , \7481 , \7482 , \7483 , \7484 , \7485 , \7486 , \7487 , \7488 ,
         \7489 , \7490 , \7491 , \7492 , \7493 , \7494 , \7495 , \7496 , \7497 , \7498 ,
         \7499 , \7500 , \7501 , \7502 , \7503 , \7504 , \7505 , \7506 , \7507 , \7508 ,
         \7509 , \7510 , \7511 , \7512 , \7513 , \7514 , \7515 , \7516 , \7517 , \7518 ,
         \7519 , \7520 , \7521 , \7522 , \7523 , \7524 , \7525 , \7526 , \7527 , \7528 ,
         \7529 , \7530 , \7531 , \7532 , \7533 , \7534 , \7535 , \7536 , \7537 , \7538 ,
         \7539 , \7540 , \7541 , \7542 , \7543 , \7544 , \7545 , \7546 , \7547 , \7548 ,
         \7549 , \7550 , \7551 , \7552 , \7553 , \7554 , \7555 , \7556 , \7557 , \7558 ,
         \7559 , \7560 , \7561 , \7562 , \7563 , \7564 , \7565 , \7566 , \7567 , \7568 ,
         \7569 , \7570 , \7571 , \7572 , \7573 , \7574 , \7575 , \7576 , \7577 , \7578 ,
         \7579 , \7580 , \7581 , \7582 , \7583 , \7584 , \7585 , \7586 , \7587 , \7588 ,
         \7589 , \7590 , \7591 , \7592 , \7593 , \7594 , \7595 , \7596 , \7597 , \7598 ,
         \7599 , \7600 , \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 , \7608 ,
         \7609 , \7610 , \7611 , \7612 , \7613 , \7614 , \7615_nG5531 , \7616 , \7617 , \7618 ,
         \7619 , \7620 , \7621 , \7622 , \7623 , \7624 , \7625 , \7626 , \7627 , \7628 ,
         \7629 , \7630 , \7631 , \7632 , \7633 , \7634 , \7635 , \7636 , \7637 , \7638 ,
         \7639 , \7640 , \7641 , \7642 , \7643 , \7644 , \7645 , \7646 , \7647 , \7648 ,
         \7649 , \7650 , \7651 , \7652 , \7653 , \7654 , \7655 , \7656 , \7657 , \7658 ,
         \7659 , \7660 , \7661 , \7662 , \7663 , \7664 , \7665 , \7666 , \7667 , \7668 ,
         \7669 , \7670 , \7671 , \7672 , \7673 , \7674 , \7675 , \7676 , \7677 , \7678 ,
         \7679 , \7680 , \7681 , \7682 , \7683 , \7684 , \7685 , \7686 , \7687 , \7688 ,
         \7689 , \7690 , \7691 , \7692 , \7693 , \7694 , \7695 , \7696 , \7697 , \7698 ,
         \7699 , \7700 , \7701 , \7702 , \7703 , \7704 , \7705 , \7706 , \7707 , \7708 ,
         \7709 , \7710 , \7711 , \7712 , \7713 , \7714 , \7715 , \7716 , \7717 , \7718 ,
         \7719 , \7720 , \7721 , \7722 , \7723 , \7724 , \7725 , \7726 , \7727 , \7728 ,
         \7729 , \7730 , \7731 , \7732 , \7733 , \7734 , \7735 , \7736 , \7737 , \7738 ,
         \7739 , \7740 , \7741 , \7742 , \7743 , \7744 , \7745 , \7746 , \7747 , \7748 ,
         \7749 , \7750 , \7751 , \7752 , \7753 , \7754 , \7755 , \7756 , \7757 , \7758 ,
         \7759 , \7760 , \7761 , \7762 , \7763 , \7764 , \7765 , \7766 , \7767 , \7768 ,
         \7769 , \7770 , \7771 , \7772 , \7773 , \7774 , \7775 , \7776 , \7777 , \7778 ,
         \7779 , \7780 , \7781 , \7782 , \7783 , \7784 , \7785 , \7786 , \7787 , \7788 ,
         \7789 , \7790 , \7791 , \7792 , \7793 , \7794 , \7795 , \7796 , \7797 , \7798 ,
         \7799 , \7800 , \7801 , \7802 , \7803 , \7804 , \7805 , \7806 , \7807 , \7808 ,
         \7809 , \7810 , \7811 , \7812 , \7813 , \7814 , \7815 , \7816 , \7817 , \7818 ,
         \7819 , \7820 , \7821 , \7822 , \7823 , \7824 , \7825 , \7826 , \7827 , \7828 ,
         \7829 , \7830 , \7831 , \7832 , \7833 , \7834 , \7835 , \7836 , \7837 , \7838 ,
         \7839 , \7840 , \7841 , \7842 , \7843 , \7844 , \7845 , \7846 , \7847 , \7848 ,
         \7849 , \7850 , \7851 , \7852 , \7853 , \7854 , \7855 , \7856 , \7857 , \7858 ,
         \7859 , \7860 , \7861 , \7862 , \7863 , \7864 , \7865 , \7866 , \7867 , \7868 ,
         \7869 , \7870 , \7871 , \7872 , \7873 , \7874 , \7875 , \7876 , \7877 , \7878 ,
         \7879 , \7880 , \7881 , \7882 , \7883 , \7884 , \7885 , \7886 , \7887 , \7888 ,
         \7889 , \7890 , \7891 , \7892 , \7893_nG552f , \7894 , \7895 , \7896 , \7897 , \7898 ,
         \7899 , \7900 , \7901 , \7902 , \7903 , \7904 , \7905 , \7906 , \7907 , \7908 ,
         \7909 , \7910 , \7911 , \7912 , \7913 , \7914 , \7915 , \7916 , \7917 , \7918 ,
         \7919 , \7920 , \7921 , \7922 , \7923 , \7924 , \7925 , \7926 , \7927 , \7928 ,
         \7929 , \7930 , \7931 , \7932 , \7933 , \7934 , \7935 , \7936 , \7937 , \7938 ,
         \7939 , \7940 , \7941 , \7942 , \7943 , \7944 , \7945 , \7946 , \7947 , \7948 ,
         \7949 , \7950 , \7951 , \7952 , \7953 , \7954 , \7955 , \7956 , \7957 , \7958 ,
         \7959 , \7960 , \7961 , \7962 , \7963 , \7964 , \7965 , \7966 , \7967 , \7968 ,
         \7969 , \7970 , \7971 , \7972 , \7973 , \7974 , \7975 , \7976 , \7977 , \7978 ,
         \7979 , \7980 , \7981 , \7982 , \7983 , \7984 , \7985 , \7986 , \7987 , \7988 ,
         \7989 , \7990 , \7991 , \7992 , \7993 , \7994 , \7995 , \7996 , \7997 , \7998 ,
         \7999 , \8000 , \8001 , \8002 , \8003 , \8004 , \8005 , \8006 , \8007 , \8008 ,
         \8009 , \8010 , \8011 , \8012 , \8013 , \8014 , \8015 , \8016 , \8017 , \8018 ,
         \8019 , \8020 , \8021 , \8022 , \8023 , \8024 , \8025 , \8026 , \8027 , \8028 ,
         \8029 , \8030 , \8031 , \8032 , \8033 , \8034 , \8035 , \8036 , \8037 , \8038 ,
         \8039 , \8040 , \8041 , \8042 , \8043 , \8044 , \8045 , \8046 , \8047 , \8048 ,
         \8049 , \8050 , \8051 , \8052 , \8053 , \8054 , \8055 , \8056 , \8057 , \8058 ,
         \8059 , \8060 , \8061 , \8062 , \8063 , \8064 , \8065 , \8066 , \8067 , \8068 ,
         \8069 , \8070 , \8071 , \8072 , \8073 , \8074 , \8075 , \8076 , \8077 , \8078 ,
         \8079 , \8080 , \8081 , \8082 , \8083 , \8084 , \8085 , \8086 , \8087 , \8088 ,
         \8089 , \8090 , \8091 , \8092 , \8093 , \8094 , \8095 , \8096 , \8097 , \8098 ,
         \8099 , \8100 , \8101 , \8102 , \8103 , \8104 , \8105 , \8106 , \8107 , \8108 ,
         \8109 , \8110 , \8111 , \8112 , \8113 , \8114 , \8115 , \8116 , \8117 , \8118 ,
         \8119 , \8120 , \8121 , \8122 , \8123 , \8124 , \8125 , \8126 , \8127 , \8128 ,
         \8129 , \8130 , \8131 , \8132 , \8133 , \8134 , \8135 , \8136 , \8137 , \8138 ,
         \8139 , \8140 , \8141 , \8142 , \8143 , \8144 , \8145 , \8146 , \8147 , \8148 ,
         \8149 , \8150 , \8151 , \8152 , \8153 , \8154 , \8155 , \8156 , \8157 , \8158 ,
         \8159 , \8160 , \8161 , \8162 , \8163 , \8164 , \8165 , \8166 , \8167 , \8168 ,
         \8169 , \8170 , \8171 , \8172 , \8173 , \8174_nG552d , \8175 , \8176 , \8177 , \8178 ,
         \8179 , \8180 , \8181 , \8182 , \8183 , \8184 , \8185 , \8186 , \8187 , \8188 ,
         \8189 , \8190 , \8191 , \8192 , \8193 , \8194 , \8195 , \8196 , \8197 , \8198 ,
         \8199 , \8200 , \8201 , \8202 , \8203 , \8204 , \8205 , \8206 , \8207 , \8208 ,
         \8209 , \8210 , \8211 , \8212 , \8213 , \8214 , \8215 , \8216 , \8217 , \8218 ,
         \8219 , \8220 , \8221 , \8222 , \8223 , \8224 , \8225 , \8226 , \8227 , \8228 ,
         \8229 , \8230 , \8231 , \8232 , \8233 , \8234 , \8235 , \8236 , \8237 , \8238 ,
         \8239 , \8240 , \8241 , \8242 , \8243 , \8244 , \8245 , \8246 , \8247 , \8248 ,
         \8249 , \8250 , \8251 , \8252 , \8253 , \8254 , \8255 , \8256 , \8257 , \8258 ,
         \8259 , \8260 , \8261 , \8262 , \8263 , \8264 , \8265 , \8266 , \8267 , \8268 ,
         \8269 , \8270 , \8271 , \8272 , \8273 , \8274 , \8275 , \8276 , \8277 , \8278 ,
         \8279 , \8280 , \8281 , \8282 , \8283 , \8284 , \8285 , \8286 , \8287 , \8288 ,
         \8289 , \8290 , \8291 , \8292 , \8293 , \8294 , \8295 , \8296 , \8297 , \8298 ,
         \8299 , \8300 , \8301 , \8302 , \8303 , \8304 , \8305 , \8306 , \8307 , \8308 ,
         \8309 , \8310 , \8311 , \8312 , \8313 , \8314 , \8315 , \8316 , \8317 , \8318 ,
         \8319 , \8320 , \8321 , \8322 , \8323 , \8324 , \8325 , \8326 , \8327 , \8328 ,
         \8329 , \8330 , \8331 , \8332 , \8333 , \8334 , \8335 , \8336 , \8337 , \8338 ,
         \8339 , \8340 , \8341 , \8342 , \8343 , \8344 , \8345 , \8346 , \8347 , \8348 ,
         \8349 , \8350 , \8351 , \8352 , \8353 , \8354 , \8355 , \8356 , \8357 , \8358 ,
         \8359 , \8360 , \8361 , \8362 , \8363 , \8364 , \8365 , \8366 , \8367 , \8368 ,
         \8369 , \8370 , \8371 , \8372 , \8373 , \8374 , \8375 , \8376 , \8377 , \8378 ,
         \8379 , \8380 , \8381 , \8382 , \8383 , \8384 , \8385 , \8386 , \8387 , \8388 ,
         \8389 , \8390 , \8391 , \8392 , \8393 , \8394 , \8395 , \8396 , \8397 , \8398 ,
         \8399 , \8400 , \8401 , \8402 , \8403 , \8404 , \8405 , \8406 , \8407 , \8408 ,
         \8409 , \8410 , \8411 , \8412 , \8413 , \8414 , \8415 , \8416 , \8417 , \8418 ,
         \8419 , \8420 , \8421 , \8422 , \8423 , \8424 , \8425 , \8426 , \8427 , \8428 ,
         \8429 , \8430 , \8431 , \8432 , \8433 , \8434 , \8435 , \8436 , \8437 , \8438 ,
         \8439 , \8440 , \8441 , \8442 , \8443 , \8444 , \8445 , \8446 , \8447 , \8448 ,
         \8449 , \8450 , \8451 , \8452 , \8453 , \8454 , \8455 , \8456 , \8457 , \8458 ,
         \8459 , \8460 , \8461 , \8462_nG552b , \8463 , \8464 , \8465 , \8466 , \8467 , \8468 ,
         \8469 , \8470 , \8471 , \8472 , \8473 , \8474 , \8475 , \8476 , \8477 , \8478 ,
         \8479 , \8480 , \8481 , \8482 , \8483 , \8484 , \8485 , \8486 , \8487 , \8488 ,
         \8489 , \8490 , \8491 , \8492 , \8493 , \8494 , \8495 , \8496 , \8497 , \8498 ,
         \8499 , \8500 , \8501 , \8502 , \8503 , \8504 , \8505 , \8506 , \8507 , \8508 ,
         \8509 , \8510 , \8511 , \8512 , \8513 , \8514 , \8515 , \8516 , \8517 , \8518 ,
         \8519 , \8520 , \8521 , \8522 , \8523 , \8524 , \8525 , \8526 , \8527 , \8528 ,
         \8529 , \8530 , \8531 , \8532 , \8533 , \8534 , \8535 , \8536 , \8537 , \8538 ,
         \8539 , \8540 , \8541 , \8542 , \8543 , \8544 , \8545 , \8546 , \8547 , \8548 ,
         \8549 , \8550 , \8551 , \8552 , \8553 , \8554 , \8555 , \8556 , \8557 , \8558 ,
         \8559 , \8560 , \8561 , \8562 , \8563 , \8564 , \8565 , \8566 , \8567 , \8568 ,
         \8569 , \8570 , \8571 , \8572 , \8573 , \8574 , \8575 , \8576 , \8577 , \8578 ,
         \8579 , \8580 , \8581 , \8582 , \8583 , \8584 , \8585 , \8586 , \8587 , \8588 ,
         \8589 , \8590 , \8591 , \8592 , \8593 , \8594 , \8595 , \8596 , \8597 , \8598 ,
         \8599 , \8600 , \8601 , \8602 , \8603 , \8604 , \8605 , \8606 , \8607 , \8608 ,
         \8609 , \8610 , \8611 , \8612 , \8613 , \8614 , \8615 , \8616 , \8617 , \8618 ,
         \8619 , \8620 , \8621 , \8622 , \8623 , \8624 , \8625 , \8626 , \8627 , \8628 ,
         \8629 , \8630 , \8631 , \8632 , \8633 , \8634 , \8635 , \8636 , \8637 , \8638 ,
         \8639 , \8640 , \8641 , \8642 , \8643 , \8644 , \8645 , \8646 , \8647 , \8648 ,
         \8649 , \8650 , \8651 , \8652 , \8653 , \8654 , \8655 , \8656 , \8657 , \8658 ,
         \8659 , \8660 , \8661 , \8662 , \8663 , \8664 , \8665 , \8666 , \8667 , \8668 ,
         \8669 , \8670 , \8671 , \8672 , \8673 , \8674 , \8675 , \8676 , \8677 , \8678 ,
         \8679 , \8680 , \8681 , \8682 , \8683 , \8684 , \8685 , \8686 , \8687 , \8688 ,
         \8689 , \8690 , \8691 , \8692 , \8693 , \8694 , \8695 , \8696 , \8697 , \8698 ,
         \8699 , \8700 , \8701 , \8702 , \8703 , \8704 , \8705 , \8706 , \8707 , \8708 ,
         \8709 , \8710 , \8711 , \8712 , \8713 , \8714 , \8715 , \8716 , \8717 , \8718 ,
         \8719 , \8720 , \8721 , \8722 , \8723 , \8724 , \8725 , \8726 , \8727 , \8728 ,
         \8729 , \8730 , \8731 , \8732 , \8733 , \8734 , \8735 , \8736 , \8737 , \8738 ,
         \8739 , \8740 , \8741 , \8742 , \8743 , \8744 , \8745 , \8746 , \8747 , \8748 ,
         \8749 , \8750 , \8751 , \8752 , \8753_nG5529 , \8754 , \8755 , \8756 , \8757 , \8758 ,
         \8759 , \8760 , \8761 , \8762 , \8763 , \8764 , \8765 , \8766 , \8767 , \8768 ,
         \8769 , \8770 , \8771 , \8772 , \8773 , \8774 , \8775 , \8776 , \8777 , \8778 ,
         \8779 , \8780 , \8781 , \8782 , \8783 , \8784 , \8785 , \8786 , \8787 , \8788 ,
         \8789 , \8790 , \8791 , \8792 , \8793 , \8794 , \8795 , \8796 , \8797 , \8798 ,
         \8799 , \8800 , \8801 , \8802 , \8803 , \8804 , \8805 , \8806 , \8807 , \8808 ,
         \8809 , \8810 , \8811 , \8812 , \8813 , \8814 , \8815 , \8816 , \8817 , \8818 ,
         \8819 , \8820 , \8821 , \8822 , \8823 , \8824 , \8825 , \8826 , \8827 , \8828 ,
         \8829 , \8830 , \8831 , \8832 , \8833 , \8834 , \8835 , \8836 , \8837 , \8838 ,
         \8839 , \8840 , \8841 , \8842 , \8843 , \8844 , \8845 , \8846 , \8847 , \8848 ,
         \8849 , \8850 , \8851 , \8852 , \8853 , \8854 , \8855 , \8856 , \8857 , \8858 ,
         \8859 , \8860 , \8861 , \8862 , \8863 , \8864 , \8865 , \8866 , \8867 , \8868 ,
         \8869 , \8870 , \8871 , \8872 , \8873 , \8874 , \8875 , \8876 , \8877 , \8878 ,
         \8879 , \8880 , \8881 , \8882 , \8883 , \8884 , \8885 , \8886 , \8887 , \8888 ,
         \8889 , \8890 , \8891 , \8892 , \8893 , \8894 , \8895 , \8896 , \8897 , \8898 ,
         \8899 , \8900 , \8901 , \8902 , \8903 , \8904 , \8905 , \8906 , \8907 , \8908 ,
         \8909 , \8910 , \8911 , \8912 , \8913 , \8914 , \8915 , \8916 , \8917 , \8918 ,
         \8919 , \8920 , \8921 , \8922 , \8923 , \8924 , \8925 , \8926 , \8927 , \8928 ,
         \8929 , \8930 , \8931 , \8932 , \8933 , \8934 , \8935 , \8936 , \8937 , \8938 ,
         \8939 , \8940 , \8941 , \8942 , \8943 , \8944 , \8945 , \8946 , \8947 , \8948 ,
         \8949 , \8950 , \8951 , \8952 , \8953 , \8954 , \8955 , \8956 , \8957 , \8958 ,
         \8959 , \8960 , \8961 , \8962 , \8963 , \8964 , \8965 , \8966 , \8967 , \8968 ,
         \8969 , \8970 , \8971 , \8972 , \8973 , \8974 , \8975 , \8976 , \8977 , \8978 ,
         \8979 , \8980 , \8981 , \8982 , \8983 , \8984 , \8985 , \8986 , \8987 , \8988 ,
         \8989 , \8990 , \8991 , \8992 , \8993 , \8994 , \8995 , \8996 , \8997 , \8998 ,
         \8999 , \9000 , \9001 , \9002 , \9003 , \9004 , \9005 , \9006 , \9007 , \9008 ,
         \9009 , \9010 , \9011 , \9012 , \9013 , \9014 , \9015 , \9016 , \9017 , \9018 ,
         \9019 , \9020 , \9021 , \9022 , \9023 , \9024 , \9025 , \9026 , \9027 , \9028 ,
         \9029 , \9030 , \9031 , \9032 , \9033 , \9034 , \9035 , \9036 , \9037 , \9038 ,
         \9039 , \9040 , \9041 , \9042 , \9043 , \9044 , \9045 , \9046 , \9047 , \9048 ,
         \9049 , \9050 , \9051_nG5527 , \9052 , \9053 , \9054 , \9055 , \9056 , \9057 , \9058 ,
         \9059 , \9060 , \9061 , \9062 , \9063 , \9064 , \9065 , \9066 , \9067 , \9068 ,
         \9069 , \9070 , \9071 , \9072 , \9073 , \9074 , \9075 , \9076 , \9077 , \9078 ,
         \9079 , \9080 , \9081 , \9082 , \9083 , \9084 , \9085 , \9086 , \9087 , \9088 ,
         \9089 , \9090 , \9091 , \9092 , \9093 , \9094 , \9095 , \9096 , \9097 , \9098 ,
         \9099 , \9100 , \9101 , \9102 , \9103 , \9104 , \9105 , \9106 , \9107 , \9108 ,
         \9109 , \9110 , \9111 , \9112 , \9113 , \9114 , \9115 , \9116 , \9117 , \9118 ,
         \9119 , \9120 , \9121 , \9122 , \9123 , \9124 , \9125 , \9126 , \9127 , \9128 ,
         \9129 , \9130 , \9131 , \9132 , \9133 , \9134 , \9135 , \9136 , \9137 , \9138 ,
         \9139 , \9140 , \9141 , \9142 , \9143 , \9144 , \9145 , \9146 , \9147 , \9148 ,
         \9149 , \9150 , \9151 , \9152 , \9153 , \9154 , \9155 , \9156 , \9157 , \9158 ,
         \9159 , \9160 , \9161 , \9162 , \9163 , \9164 , \9165 , \9166 , \9167 , \9168 ,
         \9169 , \9170 , \9171 , \9172 , \9173 , \9174 , \9175 , \9176 , \9177 , \9178 ,
         \9179 , \9180 , \9181 , \9182 , \9183 , \9184 , \9185 , \9186 , \9187 , \9188 ,
         \9189 , \9190 , \9191 , \9192 , \9193 , \9194 , \9195 , \9196 , \9197 , \9198 ,
         \9199 , \9200 , \9201 , \9202 , \9203 , \9204 , \9205 , \9206 , \9207 , \9208 ,
         \9209 , \9210 , \9211 , \9212 , \9213 , \9214 , \9215 , \9216 , \9217 , \9218 ,
         \9219 , \9220 , \9221 , \9222 , \9223 , \9224 , \9225 , \9226 , \9227 , \9228 ,
         \9229 , \9230 , \9231 , \9232 , \9233 , \9234 , \9235 , \9236 , \9237 , \9238 ,
         \9239 , \9240 , \9241 , \9242 , \9243 , \9244 , \9245 , \9246 , \9247 , \9248 ,
         \9249 , \9250 , \9251 , \9252 , \9253 , \9254 , \9255 , \9256 , \9257 , \9258 ,
         \9259 , \9260 , \9261 , \9262 , \9263 , \9264 , \9265 , \9266 , \9267 , \9268 ,
         \9269 , \9270 , \9271 , \9272 , \9273 , \9274 , \9275 , \9276 , \9277 , \9278 ,
         \9279 , \9280 , \9281 , \9282 , \9283 , \9284 , \9285 , \9286 , \9287 , \9288 ,
         \9289 , \9290 , \9291 , \9292 , \9293 , \9294 , \9295 , \9296 , \9297 , \9298 ,
         \9299 , \9300 , \9301 , \9302 , \9303 , \9304 , \9305 , \9306 , \9307 , \9308 ,
         \9309 , \9310 , \9311 , \9312 , \9313 , \9314 , \9315 , \9316 , \9317 , \9318 ,
         \9319 , \9320 , \9321 , \9322 , \9323 , \9324 , \9325 , \9326 , \9327 , \9328 ,
         \9329 , \9330 , \9331 , \9332 , \9333 , \9334 , \9335 , \9336 , \9337 , \9338 ,
         \9339 , \9340 , \9341 , \9342 , \9343 , \9344 , \9345 , \9346 , \9347 , \9348 ,
         \9349 , \9350 , \9351 , \9352_nG5525 , \9353 , \9354 , \9355 , \9356 , \9357 , \9358 ,
         \9359 , \9360 , \9361 , \9362 , \9363 , \9364 , \9365 , \9366 , \9367 , \9368 ,
         \9369 , \9370 , \9371 , \9372 , \9373 , \9374 , \9375 , \9376 , \9377 , \9378 ,
         \9379 , \9380 , \9381 , \9382 , \9383 , \9384 , \9385 , \9386 , \9387 , \9388 ,
         \9389 , \9390 , \9391 , \9392 , \9393 , \9394 , \9395 , \9396 , \9397 , \9398 ,
         \9399 , \9400 , \9401 , \9402 , \9403 , \9404 , \9405 , \9406 , \9407 , \9408 ,
         \9409 , \9410 , \9411 , \9412 , \9413 , \9414 , \9415 , \9416 , \9417 , \9418 ,
         \9419 , \9420 , \9421 , \9422 , \9423 , \9424 , \9425 , \9426 , \9427 , \9428 ,
         \9429 , \9430 , \9431 , \9432 , \9433 , \9434 , \9435 , \9436 , \9437 , \9438 ,
         \9439 , \9440 , \9441 , \9442 , \9443 , \9444 , \9445 , \9446 , \9447 , \9448 ,
         \9449 , \9450 , \9451 , \9452 , \9453 , \9454 , \9455 , \9456 , \9457 , \9458 ,
         \9459 , \9460 , \9461 , \9462 , \9463 , \9464 , \9465 , \9466 , \9467 , \9468 ,
         \9469 , \9470 , \9471 , \9472 , \9473 , \9474 , \9475 , \9476 , \9477 , \9478 ,
         \9479 , \9480 , \9481 , \9482 , \9483 , \9484 , \9485 , \9486 , \9487 , \9488 ,
         \9489 , \9490 , \9491 , \9492 , \9493 , \9494 , \9495 , \9496 , \9497 , \9498 ,
         \9499 , \9500 , \9501 , \9502 , \9503 , \9504 , \9505 , \9506 , \9507 , \9508 ,
         \9509 , \9510 , \9511 , \9512 , \9513 , \9514 , \9515 , \9516 , \9517 , \9518 ,
         \9519 , \9520 , \9521 , \9522 , \9523 , \9524 , \9525 , \9526 , \9527 , \9528 ,
         \9529 , \9530 , \9531 , \9532 , \9533 , \9534 , \9535 , \9536 , \9537 , \9538 ,
         \9539 , \9540 , \9541 , \9542 , \9543 , \9544 , \9545 , \9546 , \9547 , \9548 ,
         \9549 , \9550 , \9551 , \9552 , \9553 , \9554 , \9555 , \9556 , \9557 , \9558 ,
         \9559 , \9560 , \9561 , \9562 , \9563 , \9564 , \9565 , \9566 , \9567 , \9568 ,
         \9569 , \9570 , \9571 , \9572 , \9573 , \9574 , \9575 , \9576 , \9577 , \9578 ,
         \9579 , \9580 , \9581 , \9582 , \9583 , \9584 , \9585 , \9586 , \9587 , \9588 ,
         \9589 , \9590 , \9591 , \9592 , \9593 , \9594 , \9595 , \9596 , \9597 , \9598 ,
         \9599 , \9600 , \9601 , \9602 , \9603 , \9604 , \9605 , \9606 , \9607 , \9608 ,
         \9609 , \9610 , \9611 , \9612 , \9613 , \9614 , \9615 , \9616 , \9617 , \9618 ,
         \9619 , \9620 , \9621 , \9622 , \9623 , \9624 , \9625 , \9626 , \9627 , \9628 ,
         \9629 , \9630 , \9631 , \9632 , \9633 , \9634 , \9635 , \9636 , \9637 , \9638 ,
         \9639 , \9640 , \9641 , \9642 , \9643 , \9644 , \9645 , \9646 , \9647 , \9648 ,
         \9649 , \9650 , \9651 , \9652 , \9653 , \9654 , \9655 , \9656 , \9657 , \9658 ,
         \9659 , \9660_nG5523 , \9661 , \9662 , \9663 , \9664 , \9665 , \9666 , \9667 , \9668 ,
         \9669 , \9670 , \9671 , \9672 , \9673 , \9674 , \9675 , \9676 , \9677 , \9678 ,
         \9679 , \9680 , \9681 , \9682 , \9683 , \9684 , \9685 , \9686 , \9687 , \9688 ,
         \9689 , \9690 , \9691 , \9692 , \9693 , \9694 , \9695 , \9696 , \9697 , \9698 ,
         \9699 , \9700 , \9701 , \9702 , \9703 , \9704 , \9705 , \9706 , \9707 , \9708 ,
         \9709 , \9710 , \9711 , \9712 , \9713 , \9714 , \9715 , \9716 , \9717 , \9718 ,
         \9719 , \9720 , \9721 , \9722 , \9723 , \9724 , \9725 , \9726 , \9727 , \9728 ,
         \9729 , \9730 , \9731 , \9732 , \9733 , \9734 , \9735 , \9736 , \9737 , \9738 ,
         \9739 , \9740 , \9741 , \9742 , \9743 , \9744 , \9745 , \9746 , \9747 , \9748 ,
         \9749 , \9750 , \9751 , \9752 , \9753 , \9754 , \9755 , \9756 , \9757 , \9758 ,
         \9759 , \9760 , \9761 , \9762 , \9763 , \9764 , \9765 , \9766 , \9767 , \9768 ,
         \9769 , \9770 , \9771 , \9772 , \9773 , \9774 , \9775 , \9776 , \9777 , \9778 ,
         \9779 , \9780 , \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 , \9788 ,
         \9789 , \9790 , \9791 , \9792 , \9793 , \9794 , \9795 , \9796 , \9797 , \9798 ,
         \9799 , \9800 , \9801 , \9802 , \9803 , \9804 , \9805 , \9806 , \9807 , \9808 ,
         \9809 , \9810 , \9811 , \9812 , \9813 , \9814 , \9815 , \9816 , \9817 , \9818 ,
         \9819 , \9820 , \9821 , \9822 , \9823 , \9824 , \9825 , \9826 , \9827 , \9828 ,
         \9829 , \9830 , \9831 , \9832 , \9833 , \9834 , \9835 , \9836 , \9837 , \9838 ,
         \9839 , \9840 , \9841 , \9842 , \9843 , \9844 , \9845 , \9846 , \9847 , \9848 ,
         \9849 , \9850 , \9851 , \9852 , \9853 , \9854 , \9855 , \9856 , \9857 , \9858 ,
         \9859 , \9860 , \9861 , \9862 , \9863 , \9864 , \9865 , \9866 , \9867 , \9868 ,
         \9869 , \9870 , \9871 , \9872 , \9873 , \9874 , \9875 , \9876 , \9877 , \9878 ,
         \9879 , \9880 , \9881 , \9882 , \9883 , \9884 , \9885 , \9886 , \9887 , \9888 ,
         \9889 , \9890 , \9891 , \9892 , \9893 , \9894 , \9895 , \9896 , \9897 , \9898 ,
         \9899 , \9900 , \9901 , \9902 , \9903 , \9904 , \9905 , \9906 , \9907 , \9908 ,
         \9909 , \9910 , \9911 , \9912 , \9913 , \9914 , \9915 , \9916 , \9917 , \9918 ,
         \9919 , \9920 , \9921 , \9922 , \9923 , \9924 , \9925 , \9926 , \9927 , \9928 ,
         \9929 , \9930 , \9931 , \9932 , \9933 , \9934 , \9935 , \9936 , \9937 , \9938 ,
         \9939 , \9940 , \9941 , \9942 , \9943 , \9944 , \9945 , \9946 , \9947 , \9948 ,
         \9949 , \9950 , \9951 , \9952 , \9953 , \9954 , \9955 , \9956 , \9957 , \9958 ,
         \9959 , \9960 , \9961 , \9962 , \9963 , \9964 , \9965 , \9966 , \9967 , \9968 ,
         \9969 , \9970 , \9971_nG5521 , \9972 , \9973 , \9974 , \9975 , \9976 , \9977 , \9978 ,
         \9979 , \9980 , \9981 , \9982 , \9983 , \9984 , \9985 , \9986 , \9987 , \9988 ,
         \9989 , \9990 , \9991 , \9992 , \9993 , \9994 , \9995 , \9996 , \9997 , \9998 ,
         \9999 , \10000 , \10001 , \10002 , \10003 , \10004 , \10005 , \10006 , \10007 , \10008 ,
         \10009 , \10010 , \10011 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 , \10018 ,
         \10019 , \10020 , \10021 , \10022 , \10023 , \10024 , \10025 , \10026 , \10027 , \10028 ,
         \10029 , \10030 , \10031 , \10032 , \10033 , \10034 , \10035 , \10036 , \10037 , \10038 ,
         \10039 , \10040 , \10041 , \10042 , \10043 , \10044 , \10045 , \10046 , \10047 , \10048 ,
         \10049 , \10050 , \10051 , \10052 , \10053 , \10054 , \10055 , \10056 , \10057 , \10058 ,
         \10059 , \10060 , \10061 , \10062 , \10063 , \10064 , \10065 , \10066 , \10067 , \10068 ,
         \10069 , \10070 , \10071 , \10072 , \10073 , \10074 , \10075 , \10076 , \10077 , \10078 ,
         \10079 , \10080 , \10081 , \10082 , \10083 , \10084 , \10085 , \10086 , \10087 , \10088 ,
         \10089 , \10090 , \10091 , \10092 , \10093 , \10094 , \10095 , \10096 , \10097 , \10098 ,
         \10099 , \10100 , \10101 , \10102 , \10103 , \10104 , \10105 , \10106 , \10107 , \10108 ,
         \10109 , \10110 , \10111 , \10112 , \10113 , \10114 , \10115 , \10116 , \10117 , \10118 ,
         \10119 , \10120 , \10121 , \10122 , \10123 , \10124 , \10125 , \10126 , \10127 , \10128 ,
         \10129 , \10130 , \10131 , \10132 , \10133 , \10134 , \10135 , \10136 , \10137 , \10138 ,
         \10139 , \10140 , \10141 , \10142 , \10143 , \10144 , \10145 , \10146 , \10147 , \10148 ,
         \10149 , \10150 , \10151 , \10152 , \10153 , \10154 , \10155 , \10156 , \10157 , \10158 ,
         \10159 , \10160 , \10161 , \10162 , \10163 , \10164 , \10165 , \10166 , \10167 , \10168 ,
         \10169 , \10170 , \10171 , \10172 , \10173 , \10174 , \10175 , \10176 , \10177 , \10178 ,
         \10179 , \10180 , \10181 , \10182 , \10183 , \10184 , \10185 , \10186 , \10187 , \10188 ,
         \10189 , \10190 , \10191 , \10192 , \10193 , \10194 , \10195 , \10196 , \10197 , \10198 ,
         \10199 , \10200 , \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10207 , \10208 ,
         \10209 , \10210 , \10211 , \10212 , \10213 , \10214 , \10215 , \10216 , \10217 , \10218 ,
         \10219 , \10220 , \10221 , \10222 , \10223 , \10224 , \10225 , \10226 , \10227 , \10228 ,
         \10229 , \10230 , \10231 , \10232 , \10233 , \10234 , \10235 , \10236 , \10237 , \10238 ,
         \10239 , \10240 , \10241 , \10242 , \10243 , \10244 , \10245 , \10246 , \10247 , \10248 ,
         \10249 , \10250 , \10251 , \10252 , \10253 , \10254 , \10255 , \10256 , \10257 , \10258 ,
         \10259 , \10260 , \10261 , \10262 , \10263 , \10264 , \10265 , \10266 , \10267 , \10268 ,
         \10269 , \10270 , \10271 , \10272 , \10273 , \10274 , \10275 , \10276 , \10277 , \10278 ,
         \10279 , \10280 , \10281 , \10282 , \10283 , \10284 , \10285 , \10286 , \10287 , \10288 ,
         \10289_nG551f , \10290 , \10291 , \10292 , \10293 , \10294 , \10295 , \10296 , \10297 , \10298 ,
         \10299 , \10300 , \10301 , \10302 , \10303 , \10304 , \10305 , \10306 , \10307 , \10308 ,
         \10309 , \10310 , \10311 , \10312 , \10313 , \10314 , \10315 , \10316 , \10317 , \10318 ,
         \10319 , \10320 , \10321 , \10322 , \10323 , \10324 , \10325 , \10326 , \10327 , \10328 ,
         \10329 , \10330 , \10331 , \10332 , \10333 , \10334 , \10335 , \10336 , \10337 , \10338 ,
         \10339 , \10340 , \10341 , \10342 , \10343 , \10344 , \10345 , \10346 , \10347 , \10348 ,
         \10349 , \10350 , \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 , \10358 ,
         \10359 , \10360 , \10361 , \10362 , \10363 , \10364 , \10365 , \10366 , \10367 , \10368 ,
         \10369 , \10370 , \10371 , \10372 , \10373 , \10374 , \10375 , \10376 , \10377 , \10378 ,
         \10379 , \10380 , \10381 , \10382 , \10383 , \10384 , \10385 , \10386 , \10387 , \10388 ,
         \10389 , \10390 , \10391 , \10392 , \10393 , \10394 , \10395 , \10396 , \10397 , \10398 ,
         \10399 , \10400 , \10401 , \10402 , \10403 , \10404 , \10405 , \10406 , \10407 , \10408 ,
         \10409 , \10410 , \10411 , \10412 , \10413 , \10414 , \10415 , \10416 , \10417 , \10418 ,
         \10419 , \10420 , \10421 , \10422 , \10423 , \10424 , \10425 , \10426 , \10427 , \10428 ,
         \10429 , \10430 , \10431 , \10432 , \10433 , \10434 , \10435 , \10436 , \10437 , \10438 ,
         \10439 , \10440 , \10441 , \10442 , \10443 , \10444 , \10445 , \10446 , \10447 , \10448 ,
         \10449 , \10450 , \10451 , \10452 , \10453 , \10454 , \10455 , \10456 , \10457 , \10458 ,
         \10459 , \10460 , \10461 , \10462 , \10463 , \10464 , \10465 , \10466 , \10467 , \10468 ,
         \10469 , \10470 , \10471 , \10472 , \10473 , \10474 , \10475 , \10476 , \10477 , \10478 ,
         \10479 , \10480 , \10481 , \10482 , \10483 , \10484 , \10485 , \10486 , \10487 , \10488 ,
         \10489 , \10490 , \10491 , \10492 , \10493 , \10494 , \10495 , \10496 , \10497 , \10498 ,
         \10499 , \10500 , \10501 , \10502 , \10503 , \10504 , \10505 , \10506 , \10507 , \10508 ,
         \10509 , \10510 , \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 , \10518 ,
         \10519 , \10520 , \10521 , \10522 , \10523 , \10524 , \10525 , \10526 , \10527 , \10528 ,
         \10529 , \10530 , \10531 , \10532 , \10533 , \10534 , \10535 , \10536 , \10537 , \10538 ,
         \10539 , \10540 , \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 , \10548 ,
         \10549 , \10550 , \10551 , \10552 , \10553 , \10554 , \10555 , \10556 , \10557 , \10558 ,
         \10559 , \10560 , \10561 , \10562 , \10563 , \10564 , \10565 , \10566 , \10567 , \10568 ,
         \10569 , \10570 , \10571 , \10572 , \10573 , \10574 , \10575 , \10576 , \10577 , \10578 ,
         \10579 , \10580 , \10581 , \10582 , \10583 , \10584 , \10585 , \10586 , \10587 , \10588 ,
         \10589 , \10590 , \10591 , \10592 , \10593 , \10594 , \10595 , \10596 , \10597 , \10598 ,
         \10599 , \10600 , \10601 , \10602 , \10603 , \10604 , \10605 , \10606 , \10607 , \10608 ,
         \10609 , \10610_nG551d , \10611 , \10612 , \10613 , \10614 , \10615 , \10616 , \10617 , \10618 ,
         \10619 , \10620 , \10621 , \10622 , \10623 , \10624 , \10625 , \10626 , \10627 , \10628 ,
         \10629 , \10630 , \10631 , \10632 , \10633 , \10634 , \10635 , \10636 , \10637 , \10638 ,
         \10639 , \10640 , \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 , \10648 ,
         \10649 , \10650 , \10651 , \10652 , \10653 , \10654 , \10655 , \10656 , \10657 , \10658 ,
         \10659 , \10660 , \10661 , \10662 , \10663 , \10664 , \10665 , \10666 , \10667 , \10668 ,
         \10669 , \10670 , \10671 , \10672 , \10673 , \10674 , \10675 , \10676 , \10677 , \10678 ,
         \10679 , \10680 , \10681 , \10682 , \10683 , \10684 , \10685 , \10686 , \10687 , \10688 ,
         \10689 , \10690 , \10691 , \10692 , \10693 , \10694 , \10695 , \10696 , \10697 , \10698 ,
         \10699 , \10700 , \10701 , \10702 , \10703 , \10704 , \10705 , \10706 , \10707 , \10708 ,
         \10709 , \10710 , \10711 , \10712 , \10713 , \10714 , \10715 , \10716 , \10717 , \10718 ,
         \10719 , \10720 , \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 , \10728 ,
         \10729 , \10730 , \10731 , \10732 , \10733 , \10734 , \10735 , \10736 , \10737 , \10738 ,
         \10739 , \10740 , \10741 , \10742 , \10743 , \10744 , \10745 , \10746 , \10747 , \10748 ,
         \10749 , \10750 , \10751 , \10752 , \10753 , \10754 , \10755 , \10756 , \10757 , \10758 ,
         \10759 , \10760 , \10761 , \10762 , \10763 , \10764 , \10765 , \10766 , \10767 , \10768 ,
         \10769 , \10770 , \10771 , \10772 , \10773 , \10774 , \10775 , \10776 , \10777 , \10778 ,
         \10779 , \10780 , \10781 , \10782 , \10783 , \10784 , \10785 , \10786 , \10787 , \10788 ,
         \10789 , \10790 , \10791 , \10792 , \10793 , \10794 , \10795 , \10796 , \10797 , \10798 ,
         \10799 , \10800 , \10801 , \10802 , \10803 , \10804 , \10805 , \10806 , \10807 , \10808 ,
         \10809 , \10810 , \10811 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 , \10818 ,
         \10819 , \10820 , \10821 , \10822 , \10823 , \10824 , \10825 , \10826 , \10827 , \10828 ,
         \10829 , \10830 , \10831 , \10832 , \10833 , \10834 , \10835 , \10836 , \10837 , \10838 ,
         \10839 , \10840 , \10841 , \10842 , \10843 , \10844 , \10845 , \10846 , \10847 , \10848 ,
         \10849 , \10850 , \10851 , \10852 , \10853 , \10854 , \10855 , \10856 , \10857 , \10858 ,
         \10859 , \10860 , \10861 , \10862 , \10863 , \10864 , \10865 , \10866 , \10867 , \10868 ,
         \10869 , \10870 , \10871 , \10872 , \10873 , \10874 , \10875 , \10876 , \10877 , \10878 ,
         \10879 , \10880 , \10881 , \10882 , \10883 , \10884 , \10885 , \10886 , \10887 , \10888 ,
         \10889 , \10890 , \10891 , \10892 , \10893 , \10894 , \10895 , \10896 , \10897 , \10898 ,
         \10899 , \10900 , \10901 , \10902 , \10903 , \10904 , \10905 , \10906 , \10907 , \10908 ,
         \10909 , \10910 , \10911 , \10912 , \10913 , \10914 , \10915 , \10916 , \10917 , \10918 ,
         \10919 , \10920 , \10921 , \10922 , \10923 , \10924 , \10925 , \10926 , \10927 , \10928 ,
         \10929_nG551b , \10930 , \10931 , \10932 , \10933 , \10934 , \10935 , \10936 , \10937 , \10938 ,
         \10939 , \10940 , \10941 , \10942 , \10943 , \10944 , \10945 , \10946 , \10947 , \10948 ,
         \10949 , \10950 , \10951 , \10952 , \10953 , \10954 , \10955 , \10956 , \10957 , \10958 ,
         \10959 , \10960 , \10961 , \10962 , \10963 , \10964 , \10965 , \10966 , \10967 , \10968 ,
         \10969 , \10970 , \10971 , \10972 , \10973 , \10974 , \10975 , \10976 , \10977 , \10978 ,
         \10979 , \10980 , \10981 , \10982 , \10983 , \10984 , \10985 , \10986 , \10987 , \10988 ,
         \10989 , \10990 , \10991 , \10992 , \10993 , \10994 , \10995 , \10996 , \10997 , \10998 ,
         \10999 , \11000 , \11001 , \11002 , \11003 , \11004 , \11005 , \11006 , \11007 , \11008 ,
         \11009 , \11010 , \11011 , \11012 , \11013 , \11014 , \11015 , \11016 , \11017 , \11018 ,
         \11019 , \11020 , \11021 , \11022 , \11023 , \11024 , \11025 , \11026 , \11027 , \11028 ,
         \11029 , \11030 , \11031 , \11032 , \11033 , \11034 , \11035 , \11036 , \11037 , \11038 ,
         \11039 , \11040 , \11041 , \11042 , \11043 , \11044 , \11045 , \11046 , \11047 , \11048 ,
         \11049 , \11050 , \11051 , \11052 , \11053 , \11054 , \11055 , \11056 , \11057 , \11058 ,
         \11059 , \11060 , \11061 , \11062 , \11063 , \11064 , \11065 , \11066 , \11067 , \11068 ,
         \11069 , \11070 , \11071 , \11072 , \11073 , \11074 , \11075 , \11076 , \11077 , \11078 ,
         \11079 , \11080 , \11081 , \11082 , \11083 , \11084 , \11085 , \11086 , \11087 , \11088 ,
         \11089 , \11090 , \11091 , \11092 , \11093 , \11094 , \11095 , \11096 , \11097 , \11098 ,
         \11099 , \11100 , \11101 , \11102 , \11103 , \11104 , \11105 , \11106 , \11107 , \11108 ,
         \11109 , \11110 , \11111 , \11112 , \11113 , \11114 , \11115 , \11116 , \11117 , \11118 ,
         \11119 , \11120 , \11121 , \11122 , \11123 , \11124 , \11125 , \11126 , \11127 , \11128 ,
         \11129 , \11130 , \11131 , \11132 , \11133 , \11134 , \11135 , \11136 , \11137 , \11138 ,
         \11139 , \11140 , \11141 , \11142 , \11143 , \11144 , \11145 , \11146 , \11147 , \11148 ,
         \11149 , \11150 , \11151 , \11152 , \11153 , \11154 , \11155 , \11156 , \11157 , \11158 ,
         \11159 , \11160 , \11161 , \11162 , \11163 , \11164 , \11165 , \11166 , \11167 , \11168 ,
         \11169 , \11170 , \11171 , \11172 , \11173 , \11174 , \11175 , \11176 , \11177 , \11178 ,
         \11179 , \11180 , \11181 , \11182 , \11183 , \11184 , \11185 , \11186 , \11187 , \11188 ,
         \11189 , \11190 , \11191 , \11192 , \11193 , \11194 , \11195 , \11196 , \11197 , \11198 ,
         \11199 , \11200 , \11201 , \11202 , \11203 , \11204 , \11205 , \11206 , \11207 , \11208 ,
         \11209 , \11210 , \11211 , \11212 , \11213 , \11214 , \11215 , \11216 , \11217 , \11218 ,
         \11219 , \11220 , \11221 , \11222 , \11223 , \11224 , \11225 , \11226 , \11227 , \11228 ,
         \11229 , \11230 , \11231 , \11232 , \11233 , \11234 , \11235 , \11236 , \11237 , \11238 ,
         \11239 , \11240 , \11241 , \11242 , \11243 , \11244 , \11245 , \11246 , \11247_nG5519 , \11248 ,
         \11249 , \11250 , \11251 , \11252 , \11253 , \11254 , \11255 , \11256 , \11257 , \11258 ,
         \11259 , \11260 , \11261 , \11262 , \11263 , \11264 , \11265 , \11266 , \11267 , \11268 ,
         \11269 , \11270 , \11271 , \11272 , \11273 , \11274 , \11275 , \11276 , \11277 , \11278 ,
         \11279 , \11280 , \11281 , \11282 , \11283 , \11284 , \11285 , \11286 , \11287 , \11288 ,
         \11289 , \11290 , \11291 , \11292 , \11293 , \11294 , \11295 , \11296 , \11297 , \11298 ,
         \11299 , \11300 , \11301 , \11302 , \11303 , \11304 , \11305 , \11306 , \11307 , \11308 ,
         \11309 , \11310 , \11311 , \11312 , \11313 , \11314 , \11315 , \11316 , \11317 , \11318 ,
         \11319 , \11320 , \11321 , \11322 , \11323 , \11324 , \11325 , \11326 , \11327 , \11328 ,
         \11329 , \11330 , \11331 , \11332 , \11333 , \11334 , \11335 , \11336 , \11337 , \11338 ,
         \11339 , \11340 , \11341 , \11342 , \11343 , \11344 , \11345 , \11346 , \11347 , \11348 ,
         \11349 , \11350 , \11351 , \11352 , \11353 , \11354 , \11355 , \11356 , \11357 , \11358 ,
         \11359 , \11360 , \11361 , \11362 , \11363 , \11364 , \11365 , \11366 , \11367 , \11368 ,
         \11369 , \11370 , \11371 , \11372 , \11373 , \11374 , \11375 , \11376 , \11377 , \11378 ,
         \11379 , \11380 , \11381 , \11382 , \11383 , \11384 , \11385 , \11386 , \11387 , \11388 ,
         \11389 , \11390 , \11391 , \11392 , \11393 , \11394 , \11395 , \11396 , \11397 , \11398 ,
         \11399 , \11400 , \11401 , \11402 , \11403 , \11404 , \11405 , \11406 , \11407 , \11408 ,
         \11409 , \11410 , \11411 , \11412 , \11413 , \11414 , \11415 , \11416 , \11417 , \11418 ,
         \11419 , \11420 , \11421 , \11422 , \11423 , \11424 , \11425 , \11426 , \11427 , \11428 ,
         \11429 , \11430 , \11431 , \11432 , \11433 , \11434 , \11435 , \11436 , \11437 , \11438 ,
         \11439 , \11440 , \11441 , \11442 , \11443 , \11444 , \11445 , \11446 , \11447 , \11448 ,
         \11449 , \11450 , \11451 , \11452 , \11453 , \11454 , \11455 , \11456 , \11457 , \11458 ,
         \11459 , \11460 , \11461 , \11462 , \11463 , \11464 , \11465 , \11466 , \11467 , \11468 ,
         \11469 , \11470 , \11471 , \11472 , \11473 , \11474 , \11475 , \11476 , \11477 , \11478 ,
         \11479 , \11480 , \11481 , \11482 , \11483 , \11484 , \11485 , \11486 , \11487 , \11488 ,
         \11489 , \11490 , \11491 , \11492 , \11493 , \11494 , \11495 , \11496 , \11497 , \11498 ,
         \11499 , \11500 , \11501 , \11502 , \11503 , \11504 , \11505 , \11506 , \11507 , \11508 ,
         \11509 , \11510 , \11511 , \11512 , \11513 , \11514 , \11515 , \11516 , \11517 , \11518 ,
         \11519 , \11520 , \11521 , \11522 , \11523 , \11524 , \11525 , \11526 , \11527 , \11528 ,
         \11529 , \11530 , \11531 , \11532 , \11533 , \11534 , \11535 , \11536 , \11537 , \11538 ,
         \11539 , \11540 , \11541 , \11542 , \11543 , \11544 , \11545 , \11546 , \11547 , \11548 ,
         \11549 , \11550 , \11551 , \11552 , \11553 , \11554 , \11555 , \11556 , \11557 , \11558 ,
         \11559 , \11560 , \11561 , \11562 , \11563 , \11564_nG5517 , \11565 , \11566 , \11567 , \11568 ,
         \11569 , \11570 , \11571 , \11572 , \11573 , \11574 , \11575 , \11576 , \11577 , \11578 ,
         \11579 , \11580 , \11581 , \11582 , \11583 , \11584 , \11585 , \11586 , \11587 , \11588 ,
         \11589 , \11590 , \11591 , \11592 , \11593 , \11594 , \11595 , \11596 , \11597 , \11598 ,
         \11599 , \11600 , \11601 , \11602 , \11603 , \11604 , \11605 , \11606 , \11607 , \11608 ,
         \11609 , \11610 , \11611 , \11612 , \11613 , \11614 , \11615 , \11616 , \11617 , \11618 ,
         \11619 , \11620 , \11621 , \11622 , \11623 , \11624 , \11625 , \11626 , \11627 , \11628 ,
         \11629 , \11630 , \11631 , \11632 , \11633 , \11634 , \11635 , \11636 , \11637 , \11638 ,
         \11639 , \11640 , \11641 , \11642 , \11643 , \11644 , \11645 , \11646 , \11647 , \11648 ,
         \11649 , \11650 , \11651 , \11652 , \11653 , \11654 , \11655 , \11656 , \11657 , \11658 ,
         \11659 , \11660 , \11661 , \11662 , \11663 , \11664 , \11665 , \11666 , \11667 , \11668 ,
         \11669 , \11670 , \11671 , \11672 , \11673 , \11674 , \11675 , \11676 , \11677 , \11678 ,
         \11679 , \11680 , \11681 , \11682 , \11683 , \11684 , \11685 , \11686 , \11687 , \11688 ,
         \11689 , \11690 , \11691 , \11692 , \11693 , \11694 , \11695 , \11696 , \11697 , \11698 ,
         \11699 , \11700 , \11701 , \11702 , \11703 , \11704 , \11705 , \11706 , \11707 , \11708 ,
         \11709 , \11710 , \11711 , \11712 , \11713 , \11714 , \11715 , \11716 , \11717 , \11718 ,
         \11719 , \11720 , \11721 , \11722 , \11723 , \11724 , \11725 , \11726 , \11727 , \11728 ,
         \11729 , \11730 , \11731 , \11732 , \11733 , \11734 , \11735 , \11736 , \11737 , \11738 ,
         \11739 , \11740 , \11741 , \11742 , \11743 , \11744 , \11745 , \11746 , \11747 , \11748 ,
         \11749 , \11750 , \11751 , \11752 , \11753 , \11754 , \11755 , \11756 , \11757 , \11758 ,
         \11759 , \11760 , \11761 , \11762 , \11763 , \11764 , \11765 , \11766 , \11767 , \11768 ,
         \11769 , \11770 , \11771 , \11772 , \11773 , \11774 , \11775 , \11776 , \11777 , \11778 ,
         \11779 , \11780 , \11781 , \11782 , \11783 , \11784 , \11785 , \11786 , \11787 , \11788 ,
         \11789 , \11790 , \11791 , \11792 , \11793 , \11794 , \11795 , \11796 , \11797 , \11798 ,
         \11799 , \11800 , \11801 , \11802 , \11803 , \11804 , \11805 , \11806 , \11807 , \11808 ,
         \11809 , \11810 , \11811 , \11812 , \11813 , \11814 , \11815 , \11816 , \11817 , \11818 ,
         \11819 , \11820 , \11821 , \11822 , \11823 , \11824 , \11825 , \11826 , \11827 , \11828 ,
         \11829 , \11830 , \11831 , \11832 , \11833 , \11834 , \11835 , \11836 , \11837 , \11838 ,
         \11839 , \11840 , \11841 , \11842 , \11843 , \11844 , \11845 , \11846 , \11847 , \11848 ,
         \11849 , \11850 , \11851 , \11852 , \11853 , \11854 , \11855 , \11856 , \11857 , \11858 ,
         \11859 , \11860 , \11861 , \11862 , \11863 , \11864 , \11865 , \11866 , \11867 , \11868 ,
         \11869 , \11870 , \11871 , \11872 , \11873 , \11874 , \11875 , \11876 , \11877 , \11878 ,
         \11879 , \11880_nG5515 , \11881 , \11882 , \11883 , \11884 , \11885 , \11886 , \11887 , \11888 ,
         \11889 , \11890 , \11891 , \11892 , \11893 , \11894 , \11895 , \11896 , \11897 , \11898 ,
         \11899 , \11900 , \11901 , \11902 , \11903 , \11904 , \11905 , \11906 , \11907 , \11908 ,
         \11909 , \11910 , \11911 , \11912 , \11913 , \11914 , \11915 , \11916 , \11917 , \11918 ,
         \11919 , \11920 , \11921 , \11922 , \11923 , \11924 , \11925 , \11926 , \11927 , \11928 ,
         \11929 , \11930 , \11931 , \11932 , \11933 , \11934 , \11935 , \11936 , \11937 , \11938 ,
         \11939 , \11940 , \11941 , \11942 , \11943 , \11944 , \11945 , \11946 , \11947 , \11948 ,
         \11949 , \11950 , \11951 , \11952 , \11953 , \11954 , \11955 , \11956 , \11957 , \11958 ,
         \11959 , \11960 , \11961 , \11962 , \11963 , \11964 , \11965 , \11966 , \11967 , \11968 ,
         \11969 , \11970 , \11971 , \11972 , \11973 , \11974 , \11975 , \11976 , \11977 , \11978 ,
         \11979 , \11980 , \11981 , \11982 , \11983 , \11984 , \11985 , \11986 , \11987 , \11988 ,
         \11989 , \11990 , \11991 , \11992 , \11993 , \11994 , \11995 , \11996 , \11997 , \11998 ,
         \11999 , \12000 , \12001 , \12002 , \12003 , \12004 , \12005 , \12006 , \12007 , \12008 ,
         \12009 , \12010 , \12011 , \12012 , \12013 , \12014 , \12015 , \12016 , \12017 , \12018 ,
         \12019 , \12020 , \12021 , \12022 , \12023 , \12024 , \12025 , \12026 , \12027 , \12028 ,
         \12029 , \12030 , \12031 , \12032 , \12033 , \12034 , \12035 , \12036 , \12037 , \12038 ,
         \12039 , \12040 , \12041 , \12042 , \12043 , \12044 , \12045 , \12046 , \12047 , \12048 ,
         \12049 , \12050 , \12051 , \12052 , \12053 , \12054 , \12055 , \12056 , \12057 , \12058 ,
         \12059 , \12060 , \12061 , \12062 , \12063 , \12064 , \12065 , \12066 , \12067 , \12068 ,
         \12069 , \12070 , \12071 , \12072 , \12073 , \12074 , \12075 , \12076 , \12077 , \12078 ,
         \12079 , \12080 , \12081 , \12082 , \12083 , \12084 , \12085 , \12086 , \12087 , \12088 ,
         \12089 , \12090 , \12091 , \12092 , \12093 , \12094 , \12095 , \12096 , \12097 , \12098 ,
         \12099 , \12100 , \12101 , \12102 , \12103 , \12104 , \12105 , \12106 , \12107 , \12108 ,
         \12109 , \12110 , \12111 , \12112 , \12113 , \12114 , \12115 , \12116 , \12117 , \12118 ,
         \12119 , \12120 , \12121 , \12122 , \12123 , \12124 , \12125 , \12126 , \12127 , \12128 ,
         \12129 , \12130 , \12131 , \12132 , \12133 , \12134 , \12135 , \12136 , \12137 , \12138 ,
         \12139 , \12140 , \12141 , \12142 , \12143 , \12144 , \12145 , \12146 , \12147 , \12148 ,
         \12149 , \12150 , \12151 , \12152 , \12153 , \12154 , \12155 , \12156 , \12157 , \12158 ,
         \12159 , \12160 , \12161 , \12162 , \12163 , \12164 , \12165 , \12166 , \12167 , \12168 ,
         \12169 , \12170 , \12171 , \12172 , \12173 , \12174 , \12175 , \12176 , \12177 , \12178 ,
         \12179 , \12180 , \12181 , \12182 , \12183 , \12184 , \12185 , \12186 , \12187 , \12188 ,
         \12189 , \12190 , \12191_nG5513 , \12192 , \12193 , \12194 , \12195 , \12196 , \12197 , \12198 ,
         \12199 , \12200 , \12201 , \12202 , \12203 , \12204 , \12205 , \12206 , \12207 , \12208 ,
         \12209 , \12210 , \12211 , \12212 , \12213 , \12214 , \12215 , \12216 , \12217 , \12218 ,
         \12219 , \12220 , \12221 , \12222 , \12223 , \12224 , \12225 , \12226 , \12227 , \12228 ,
         \12229 , \12230 , \12231 , \12232 , \12233 , \12234 , \12235 , \12236 , \12237 , \12238 ,
         \12239 , \12240 , \12241 , \12242 , \12243 , \12244 , \12245 , \12246 , \12247 , \12248 ,
         \12249 , \12250 , \12251 , \12252 , \12253 , \12254 , \12255 , \12256 , \12257 , \12258 ,
         \12259 , \12260 , \12261 , \12262 , \12263 , \12264 , \12265 , \12266 , \12267 , \12268 ,
         \12269 , \12270 , \12271 , \12272 , \12273 , \12274 , \12275 , \12276 , \12277 , \12278 ,
         \12279 , \12280 , \12281 , \12282 , \12283 , \12284 , \12285 , \12286 , \12287 , \12288 ,
         \12289 , \12290 , \12291 , \12292 , \12293 , \12294 , \12295 , \12296 , \12297 , \12298 ,
         \12299 , \12300 , \12301 , \12302 , \12303 , \12304 , \12305 , \12306 , \12307 , \12308 ,
         \12309 , \12310 , \12311 , \12312 , \12313 , \12314 , \12315 , \12316 , \12317 , \12318 ,
         \12319 , \12320 , \12321 , \12322 , \12323 , \12324 , \12325 , \12326 , \12327 , \12328 ,
         \12329 , \12330 , \12331 , \12332 , \12333 , \12334 , \12335 , \12336 , \12337 , \12338 ,
         \12339 , \12340 , \12341 , \12342 , \12343 , \12344 , \12345 , \12346 , \12347 , \12348 ,
         \12349 , \12350 , \12351 , \12352 , \12353 , \12354 , \12355 , \12356 , \12357 , \12358 ,
         \12359 , \12360 , \12361 , \12362 , \12363 , \12364 , \12365 , \12366 , \12367 , \12368 ,
         \12369 , \12370 , \12371 , \12372 , \12373 , \12374 , \12375 , \12376 , \12377 , \12378 ,
         \12379 , \12380 , \12381 , \12382 , \12383 , \12384 , \12385 , \12386 , \12387 , \12388 ,
         \12389 , \12390 , \12391 , \12392 , \12393 , \12394 , \12395 , \12396 , \12397 , \12398 ,
         \12399 , \12400 , \12401 , \12402 , \12403 , \12404 , \12405 , \12406 , \12407 , \12408 ,
         \12409 , \12410 , \12411 , \12412 , \12413 , \12414 , \12415 , \12416 , \12417 , \12418 ,
         \12419 , \12420 , \12421 , \12422 , \12423 , \12424 , \12425 , \12426 , \12427 , \12428 ,
         \12429 , \12430 , \12431 , \12432 , \12433 , \12434 , \12435 , \12436 , \12437 , \12438 ,
         \12439 , \12440 , \12441 , \12442 , \12443 , \12444 , \12445 , \12446 , \12447 , \12448 ,
         \12449 , \12450 , \12451 , \12452 , \12453 , \12454 , \12455 , \12456 , \12457 , \12458 ,
         \12459 , \12460 , \12461 , \12462 , \12463 , \12464 , \12465 , \12466 , \12467 , \12468 ,
         \12469 , \12470 , \12471 , \12472 , \12473 , \12474 , \12475 , \12476 , \12477 , \12478 ,
         \12479 , \12480 , \12481 , \12482 , \12483 , \12484 , \12485 , \12486 , \12487 , \12488 ,
         \12489 , \12490 , \12491 , \12492 , \12493 , \12494 , \12495 , \12496 , \12497 , \12498 ,
         \12499_nG5511 , \12500 , \12501 , \12502 , \12503 , \12504 , \12505 , \12506 , \12507 , \12508 ,
         \12509 , \12510 , \12511 , \12512 , \12513 , \12514 , \12515 , \12516 , \12517 , \12518 ,
         \12519 , \12520 , \12521 , \12522 , \12523 , \12524 , \12525 , \12526 , \12527 , \12528 ,
         \12529 , \12530 , \12531 , \12532 , \12533 , \12534 , \12535 , \12536 , \12537 , \12538 ,
         \12539 , \12540 , \12541 , \12542 , \12543 , \12544 , \12545 , \12546 , \12547 , \12548 ,
         \12549 , \12550 , \12551 , \12552 , \12553 , \12554 , \12555 , \12556 , \12557 , \12558 ,
         \12559 , \12560 , \12561 , \12562 , \12563 , \12564 , \12565 , \12566 , \12567 , \12568 ,
         \12569 , \12570 , \12571 , \12572 , \12573 , \12574 , \12575 , \12576 , \12577 , \12578 ,
         \12579 , \12580 , \12581 , \12582 , \12583 , \12584 , \12585 , \12586 , \12587 , \12588 ,
         \12589 , \12590 , \12591 , \12592 , \12593 , \12594 , \12595 , \12596 , \12597 , \12598 ,
         \12599 , \12600 , \12601 , \12602 , \12603 , \12604 , \12605 , \12606 , \12607 , \12608 ,
         \12609 , \12610 , \12611 , \12612 , \12613 , \12614 , \12615 , \12616 , \12617 , \12618 ,
         \12619 , \12620 , \12621 , \12622 , \12623 , \12624 , \12625 , \12626 , \12627 , \12628 ,
         \12629 , \12630 , \12631 , \12632 , \12633 , \12634 , \12635 , \12636 , \12637 , \12638 ,
         \12639 , \12640 , \12641 , \12642 , \12643 , \12644 , \12645 , \12646 , \12647 , \12648 ,
         \12649 , \12650 , \12651 , \12652 , \12653 , \12654 , \12655 , \12656 , \12657 , \12658 ,
         \12659 , \12660 , \12661 , \12662 , \12663 , \12664 , \12665 , \12666 , \12667 , \12668 ,
         \12669 , \12670 , \12671 , \12672 , \12673 , \12674 , \12675 , \12676 , \12677 , \12678 ,
         \12679 , \12680 , \12681 , \12682 , \12683 , \12684 , \12685 , \12686 , \12687 , \12688 ,
         \12689 , \12690 , \12691 , \12692 , \12693 , \12694 , \12695 , \12696 , \12697 , \12698 ,
         \12699 , \12700 , \12701 , \12702 , \12703 , \12704 , \12705 , \12706 , \12707 , \12708 ,
         \12709 , \12710 , \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 , \12718 ,
         \12719 , \12720 , \12721 , \12722 , \12723 , \12724 , \12725 , \12726 , \12727 , \12728 ,
         \12729 , \12730 , \12731 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 , \12738 ,
         \12739 , \12740 , \12741 , \12742 , \12743 , \12744 , \12745 , \12746 , \12747 , \12748 ,
         \12749 , \12750 , \12751 , \12752 , \12753 , \12754 , \12755 , \12756 , \12757 , \12758 ,
         \12759 , \12760 , \12761 , \12762 , \12763 , \12764 , \12765 , \12766 , \12767 , \12768 ,
         \12769 , \12770 , \12771 , \12772 , \12773 , \12774 , \12775 , \12776 , \12777 , \12778 ,
         \12779 , \12780 , \12781 , \12782 , \12783 , \12784 , \12785 , \12786 , \12787 , \12788 ,
         \12789 , \12790 , \12791 , \12792 , \12793 , \12794 , \12795 , \12796 , \12797 , \12798 ,
         \12799 , \12800 , \12801 , \12802_nG550f , \12803 , \12804 , \12805 , \12806 , \12807 , \12808 ,
         \12809 , \12810 , \12811 , \12812 , \12813 , \12814 , \12815 , \12816 , \12817 , \12818 ,
         \12819 , \12820 , \12821 , \12822 , \12823 , \12824 , \12825 , \12826 , \12827 , \12828 ,
         \12829 , \12830 , \12831 , \12832 , \12833 , \12834 , \12835 , \12836 , \12837 , \12838 ,
         \12839 , \12840 , \12841 , \12842 , \12843 , \12844 , \12845 , \12846 , \12847 , \12848 ,
         \12849 , \12850 , \12851 , \12852 , \12853 , \12854 , \12855 , \12856 , \12857 , \12858 ,
         \12859 , \12860 , \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 , \12868 ,
         \12869 , \12870 , \12871 , \12872 , \12873 , \12874 , \12875 , \12876 , \12877 , \12878 ,
         \12879 , \12880 , \12881 , \12882 , \12883 , \12884 , \12885 , \12886 , \12887 , \12888 ,
         \12889 , \12890 , \12891 , \12892 , \12893 , \12894 , \12895 , \12896 , \12897 , \12898 ,
         \12899 , \12900 , \12901 , \12902 , \12903 , \12904 , \12905 , \12906 , \12907 , \12908 ,
         \12909 , \12910 , \12911 , \12912 , \12913 , \12914 , \12915 , \12916 , \12917 , \12918 ,
         \12919 , \12920 , \12921 , \12922 , \12923 , \12924 , \12925 , \12926 , \12927 , \12928 ,
         \12929 , \12930 , \12931 , \12932 , \12933 , \12934 , \12935 , \12936 , \12937 , \12938 ,
         \12939 , \12940 , \12941 , \12942 , \12943 , \12944 , \12945 , \12946 , \12947 , \12948 ,
         \12949 , \12950 , \12951 , \12952 , \12953 , \12954 , \12955 , \12956 , \12957 , \12958 ,
         \12959 , \12960 , \12961 , \12962 , \12963 , \12964 , \12965 , \12966 , \12967 , \12968 ,
         \12969 , \12970 , \12971 , \12972 , \12973 , \12974 , \12975 , \12976 , \12977 , \12978 ,
         \12979 , \12980 , \12981 , \12982 , \12983 , \12984 , \12985 , \12986 , \12987 , \12988 ,
         \12989 , \12990 , \12991 , \12992 , \12993 , \12994 , \12995 , \12996 , \12997 , \12998 ,
         \12999 , \13000 , \13001 , \13002 , \13003 , \13004 , \13005 , \13006 , \13007 , \13008 ,
         \13009 , \13010 , \13011 , \13012 , \13013 , \13014 , \13015 , \13016 , \13017 , \13018 ,
         \13019 , \13020 , \13021 , \13022 , \13023 , \13024 , \13025 , \13026 , \13027 , \13028 ,
         \13029 , \13030 , \13031 , \13032 , \13033 , \13034 , \13035 , \13036 , \13037 , \13038 ,
         \13039 , \13040 , \13041 , \13042 , \13043 , \13044 , \13045 , \13046 , \13047 , \13048 ,
         \13049 , \13050 , \13051 , \13052 , \13053 , \13054 , \13055 , \13056 , \13057 , \13058 ,
         \13059 , \13060 , \13061 , \13062 , \13063 , \13064 , \13065 , \13066 , \13067 , \13068 ,
         \13069 , \13070 , \13071 , \13072 , \13073 , \13074 , \13075 , \13076 , \13077 , \13078 ,
         \13079 , \13080 , \13081 , \13082 , \13083 , \13084 , \13085 , \13086 , \13087 , \13088 ,
         \13089 , \13090 , \13091 , \13092 , \13093 , \13094 , \13095 , \13096 , \13097 , \13098_nG550d ,
         \13099 , \13100 , \13101 , \13102 , \13103 , \13104 , \13105 , \13106 , \13107 , \13108 ,
         \13109 , \13110 , \13111 , \13112 , \13113 , \13114 , \13115 , \13116 , \13117 , \13118 ,
         \13119 , \13120 , \13121 , \13122 , \13123 , \13124 , \13125 , \13126 , \13127 , \13128 ,
         \13129 , \13130 , \13131 , \13132 , \13133 , \13134 , \13135 , \13136 , \13137 , \13138 ,
         \13139 , \13140 , \13141 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 , \13148 ,
         \13149 , \13150 , \13151 , \13152 , \13153 , \13154 , \13155 , \13156 , \13157 , \13158 ,
         \13159 , \13160 , \13161 , \13162 , \13163 , \13164 , \13165 , \13166 , \13167 , \13168 ,
         \13169 , \13170 , \13171 , \13172 , \13173 , \13174 , \13175 , \13176 , \13177 , \13178 ,
         \13179 , \13180 , \13181 , \13182 , \13183 , \13184 , \13185 , \13186 , \13187 , \13188 ,
         \13189 , \13190 , \13191 , \13192 , \13193 , \13194 , \13195 , \13196 , \13197 , \13198 ,
         \13199 , \13200 , \13201 , \13202 , \13203 , \13204 , \13205 , \13206 , \13207 , \13208 ,
         \13209 , \13210 , \13211 , \13212 , \13213 , \13214 , \13215 , \13216 , \13217 , \13218 ,
         \13219 , \13220 , \13221 , \13222 , \13223 , \13224 , \13225 , \13226 , \13227 , \13228 ,
         \13229 , \13230 , \13231 , \13232 , \13233 , \13234 , \13235 , \13236 , \13237 , \13238 ,
         \13239 , \13240 , \13241 , \13242 , \13243 , \13244 , \13245 , \13246 , \13247 , \13248 ,
         \13249 , \13250 , \13251 , \13252 , \13253 , \13254 , \13255 , \13256 , \13257 , \13258 ,
         \13259 , \13260 , \13261 , \13262 , \13263 , \13264 , \13265 , \13266 , \13267 , \13268 ,
         \13269 , \13270 , \13271 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 , \13278 ,
         \13279 , \13280 , \13281 , \13282 , \13283 , \13284 , \13285 , \13286 , \13287 , \13288 ,
         \13289 , \13290 , \13291 , \13292 , \13293 , \13294 , \13295 , \13296 , \13297 , \13298 ,
         \13299 , \13300 , \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 , \13308 ,
         \13309 , \13310 , \13311 , \13312 , \13313 , \13314 , \13315 , \13316 , \13317 , \13318 ,
         \13319 , \13320 , \13321 , \13322 , \13323 , \13324 , \13325 , \13326 , \13327 , \13328 ,
         \13329 , \13330 , \13331 , \13332 , \13333 , \13334 , \13335 , \13336 , \13337 , \13338 ,
         \13339 , \13340 , \13341 , \13342 , \13343 , \13344 , \13345 , \13346 , \13347 , \13348 ,
         \13349 , \13350 , \13351 , \13352 , \13353 , \13354 , \13355 , \13356 , \13357 , \13358 ,
         \13359 , \13360 , \13361 , \13362 , \13363 , \13364 , \13365 , \13366 , \13367 , \13368 ,
         \13369 , \13370 , \13371 , \13372 , \13373 , \13374 , \13375 , \13376 , \13377 , \13378 ,
         \13379 , \13380 , \13381 , \13382 , \13383 , \13384 , \13385 , \13386 , \13387 , \13388 ,
         \13389_nG550b , \13390 , \13391 , \13392 , \13393 , \13394 , \13395 , \13396 , \13397 , \13398 ,
         \13399 , \13400 , \13401 , \13402 , \13403 , \13404 , \13405 , \13406 , \13407 , \13408 ,
         \13409 , \13410 , \13411 , \13412 , \13413 , \13414 , \13415 , \13416 , \13417 , \13418 ,
         \13419 , \13420 , \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 , \13428 ,
         \13429 , \13430 , \13431 , \13432 , \13433 , \13434 , \13435 , \13436 , \13437 , \13438 ,
         \13439 , \13440 , \13441 , \13442 , \13443 , \13444 , \13445 , \13446 , \13447 , \13448 ,
         \13449 , \13450 , \13451 , \13452 , \13453 , \13454 , \13455 , \13456 , \13457 , \13458 ,
         \13459 , \13460 , \13461 , \13462 , \13463 , \13464 , \13465 , \13466 , \13467 , \13468 ,
         \13469 , \13470 , \13471 , \13472 , \13473 , \13474 , \13475 , \13476 , \13477 , \13478 ,
         \13479 , \13480 , \13481 , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 , \13488 ,
         \13489 , \13490 , \13491 , \13492 , \13493 , \13494 , \13495 , \13496 , \13497 , \13498 ,
         \13499 , \13500 , \13501 , \13502 , \13503 , \13504 , \13505 , \13506 , \13507 , \13508 ,
         \13509 , \13510 , \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 , \13518 ,
         \13519 , \13520 , \13521 , \13522 , \13523 , \13524 , \13525 , \13526 , \13527 , \13528 ,
         \13529 , \13530 , \13531 , \13532 , \13533 , \13534 , \13535 , \13536 , \13537 , \13538 ,
         \13539 , \13540 , \13541 , \13542 , \13543 , \13544 , \13545 , \13546 , \13547 , \13548 ,
         \13549 , \13550 , \13551 , \13552 , \13553 , \13554 , \13555 , \13556 , \13557 , \13558 ,
         \13559 , \13560 , \13561 , \13562 , \13563 , \13564 , \13565 , \13566 , \13567 , \13568 ,
         \13569 , \13570 , \13571 , \13572 , \13573 , \13574 , \13575 , \13576 , \13577 , \13578 ,
         \13579 , \13580 , \13581 , \13582 , \13583 , \13584 , \13585 , \13586 , \13587 , \13588 ,
         \13589 , \13590 , \13591 , \13592 , \13593 , \13594 , \13595 , \13596 , \13597 , \13598 ,
         \13599 , \13600 , \13601 , \13602 , \13603 , \13604 , \13605 , \13606 , \13607 , \13608 ,
         \13609 , \13610 , \13611 , \13612 , \13613 , \13614 , \13615 , \13616 , \13617 , \13618 ,
         \13619 , \13620 , \13621 , \13622 , \13623 , \13624 , \13625 , \13626 , \13627 , \13628 ,
         \13629 , \13630 , \13631 , \13632 , \13633 , \13634 , \13635 , \13636 , \13637 , \13638 ,
         \13639 , \13640 , \13641 , \13642 , \13643 , \13644 , \13645 , \13646 , \13647 , \13648 ,
         \13649 , \13650 , \13651 , \13652 , \13653 , \13654 , \13655 , \13656 , \13657 , \13658 ,
         \13659 , \13660 , \13661 , \13662 , \13663 , \13664 , \13665 , \13666 , \13667 , \13668 ,
         \13669 , \13670 , \13671 , \13672_nG5509 , \13673 , \13674 , \13675 , \13676 , \13677 , \13678 ,
         \13679 , \13680 , \13681 , \13682 , \13683 , \13684 , \13685 , \13686 , \13687 , \13688 ,
         \13689 , \13690 , \13691 , \13692 , \13693 , \13694 , \13695 , \13696 , \13697 , \13698 ,
         \13699 , \13700 , \13701 , \13702 , \13703 , \13704 , \13705 , \13706 , \13707 , \13708 ,
         \13709 , \13710 , \13711 , \13712 , \13713 , \13714 , \13715 , \13716 , \13717 , \13718 ,
         \13719 , \13720 , \13721 , \13722 , \13723 , \13724 , \13725 , \13726 , \13727 , \13728 ,
         \13729 , \13730 , \13731 , \13732 , \13733 , \13734 , \13735 , \13736 , \13737 , \13738 ,
         \13739 , \13740 , \13741 , \13742 , \13743 , \13744 , \13745 , \13746 , \13747 , \13748 ,
         \13749 , \13750 , \13751 , \13752 , \13753 , \13754 , \13755 , \13756 , \13757 , \13758 ,
         \13759 , \13760 , \13761 , \13762 , \13763 , \13764 , \13765 , \13766 , \13767 , \13768 ,
         \13769 , \13770 , \13771 , \13772 , \13773 , \13774 , \13775 , \13776 , \13777 , \13778 ,
         \13779 , \13780 , \13781 , \13782 , \13783 , \13784 , \13785 , \13786 , \13787 , \13788 ,
         \13789 , \13790 , \13791 , \13792 , \13793 , \13794 , \13795 , \13796 , \13797 , \13798 ,
         \13799 , \13800 , \13801 , \13802 , \13803 , \13804 , \13805 , \13806 , \13807 , \13808 ,
         \13809 , \13810 , \13811 , \13812 , \13813 , \13814 , \13815 , \13816 , \13817 , \13818 ,
         \13819 , \13820 , \13821 , \13822 , \13823 , \13824 , \13825 , \13826 , \13827 , \13828 ,
         \13829 , \13830 , \13831 , \13832 , \13833 , \13834 , \13835 , \13836 , \13837 , \13838 ,
         \13839 , \13840 , \13841 , \13842 , \13843 , \13844 , \13845 , \13846 , \13847 , \13848 ,
         \13849 , \13850 , \13851 , \13852 , \13853 , \13854 , \13855 , \13856 , \13857 , \13858 ,
         \13859 , \13860 , \13861 , \13862 , \13863 , \13864 , \13865 , \13866 , \13867 , \13868 ,
         \13869 , \13870 , \13871 , \13872 , \13873 , \13874 , \13875 , \13876 , \13877 , \13878 ,
         \13879 , \13880 , \13881 , \13882 , \13883 , \13884 , \13885 , \13886 , \13887 , \13888 ,
         \13889 , \13890 , \13891 , \13892 , \13893 , \13894 , \13895 , \13896 , \13897 , \13898 ,
         \13899 , \13900 , \13901 , \13902 , \13903 , \13904 , \13905 , \13906 , \13907 , \13908 ,
         \13909 , \13910 , \13911 , \13912 , \13913 , \13914 , \13915 , \13916 , \13917 , \13918 ,
         \13919 , \13920 , \13921 , \13922 , \13923 , \13924 , \13925 , \13926 , \13927 , \13928 ,
         \13929 , \13930 , \13931 , \13932 , \13933 , \13934 , \13935 , \13936 , \13937 , \13938 ,
         \13939 , \13940 , \13941 , \13942 , \13943 , \13944 , \13945 , \13946 , \13947 , \13948 ,
         \13949 , \13950 , \13951 , \13952 , \13953_nG5507 , \13954 , \13955 , \13956 , \13957 , \13958 ,
         \13959 , \13960 , \13961 , \13962 , \13963 , \13964 , \13965 , \13966 , \13967 , \13968 ,
         \13969 , \13970 , \13971 , \13972 , \13973 , \13974 , \13975 , \13976 , \13977 , \13978 ,
         \13979 , \13980 , \13981 , \13982 , \13983 , \13984 , \13985 , \13986 , \13987 , \13988 ,
         \13989 , \13990 , \13991 , \13992 , \13993 , \13994 , \13995 , \13996 , \13997 , \13998 ,
         \13999 , \14000 , \14001 , \14002 , \14003 , \14004 , \14005 , \14006 , \14007 , \14008 ,
         \14009 , \14010 , \14011 , \14012 , \14013 , \14014 , \14015 , \14016 , \14017 , \14018 ,
         \14019 , \14020 , \14021 , \14022 , \14023 , \14024 , \14025 , \14026 , \14027 , \14028 ,
         \14029 , \14030 , \14031 , \14032 , \14033 , \14034 , \14035 , \14036 , \14037 , \14038 ,
         \14039 , \14040 , \14041 , \14042 , \14043 , \14044 , \14045 , \14046 , \14047 , \14048 ,
         \14049 , \14050 , \14051 , \14052 , \14053 , \14054 , \14055 , \14056 , \14057 , \14058 ,
         \14059 , \14060 , \14061 , \14062 , \14063 , \14064 , \14065 , \14066 , \14067 , \14068 ,
         \14069 , \14070 , \14071 , \14072 , \14073 , \14074 , \14075 , \14076 , \14077 , \14078 ,
         \14079 , \14080 , \14081 , \14082 , \14083 , \14084 , \14085 , \14086 , \14087 , \14088 ,
         \14089 , \14090 , \14091 , \14092 , \14093 , \14094 , \14095 , \14096 , \14097 , \14098 ,
         \14099 , \14100 , \14101 , \14102 , \14103 , \14104 , \14105 , \14106 , \14107 , \14108 ,
         \14109 , \14110 , \14111 , \14112 , \14113 , \14114 , \14115 , \14116 , \14117 , \14118 ,
         \14119 , \14120 , \14121 , \14122 , \14123 , \14124 , \14125 , \14126 , \14127 , \14128 ,
         \14129 , \14130 , \14131 , \14132 , \14133 , \14134 , \14135 , \14136 , \14137 , \14138 ,
         \14139 , \14140 , \14141 , \14142 , \14143 , \14144 , \14145 , \14146 , \14147 , \14148 ,
         \14149 , \14150 , \14151 , \14152 , \14153 , \14154 , \14155 , \14156 , \14157 , \14158 ,
         \14159 , \14160 , \14161 , \14162 , \14163 , \14164 , \14165 , \14166 , \14167 , \14168 ,
         \14169 , \14170 , \14171 , \14172 , \14173 , \14174 , \14175 , \14176 , \14177 , \14178 ,
         \14179 , \14180 , \14181 , \14182 , \14183 , \14184 , \14185 , \14186 , \14187 , \14188 ,
         \14189 , \14190 , \14191 , \14192 , \14193 , \14194 , \14195 , \14196 , \14197 , \14198 ,
         \14199 , \14200 , \14201 , \14202 , \14203 , \14204 , \14205 , \14206 , \14207 , \14208 ,
         \14209 , \14210 , \14211 , \14212 , \14213 , \14214 , \14215 , \14216 , \14217 , \14218 ,
         \14219 , \14220 , \14221 , \14222 , \14223 , \14224 , \14225 , \14226_nG5505 , \14227 , \14228 ,
         \14229 , \14230 , \14231 , \14232 , \14233 , \14234 , \14235 , \14236 , \14237 , \14238 ,
         \14239 , \14240 , \14241 , \14242 , \14243 , \14244 , \14245 , \14246 , \14247 , \14248 ,
         \14249 , \14250 , \14251 , \14252 , \14253 , \14254 , \14255 , \14256 , \14257 , \14258 ,
         \14259 , \14260 , \14261 , \14262 , \14263 , \14264 , \14265 , \14266 , \14267 , \14268 ,
         \14269 , \14270 , \14271 , \14272 , \14273 , \14274 , \14275 , \14276 , \14277 , \14278 ,
         \14279 , \14280 , \14281 , \14282 , \14283 , \14284 , \14285 , \14286 , \14287 , \14288 ,
         \14289 , \14290 , \14291 , \14292 , \14293 , \14294 , \14295 , \14296 , \14297 , \14298 ,
         \14299 , \14300 , \14301 , \14302 , \14303 , \14304 , \14305 , \14306 , \14307 , \14308 ,
         \14309 , \14310 , \14311 , \14312 , \14313 , \14314 , \14315 , \14316 , \14317 , \14318 ,
         \14319 , \14320 , \14321 , \14322 , \14323 , \14324 , \14325 , \14326 , \14327 , \14328 ,
         \14329 , \14330 , \14331 , \14332 , \14333 , \14334 , \14335 , \14336 , \14337 , \14338 ,
         \14339 , \14340 , \14341 , \14342 , \14343 , \14344 , \14345 , \14346 , \14347 , \14348 ,
         \14349 , \14350 , \14351 , \14352 , \14353 , \14354 , \14355 , \14356 , \14357 , \14358 ,
         \14359 , \14360 , \14361 , \14362 , \14363 , \14364 , \14365 , \14366 , \14367 , \14368 ,
         \14369 , \14370 , \14371 , \14372 , \14373 , \14374 , \14375 , \14376 , \14377 , \14378 ,
         \14379 , \14380 , \14381 , \14382 , \14383 , \14384 , \14385 , \14386 , \14387 , \14388 ,
         \14389 , \14390 , \14391 , \14392 , \14393 , \14394 , \14395 , \14396 , \14397 , \14398 ,
         \14399 , \14400 , \14401 , \14402 , \14403 , \14404 , \14405 , \14406 , \14407 , \14408 ,
         \14409 , \14410 , \14411 , \14412 , \14413 , \14414 , \14415 , \14416 , \14417 , \14418 ,
         \14419 , \14420 , \14421 , \14422 , \14423 , \14424 , \14425 , \14426 , \14427 , \14428 ,
         \14429 , \14430 , \14431 , \14432 , \14433 , \14434 , \14435 , \14436 , \14437 , \14438 ,
         \14439 , \14440 , \14441 , \14442 , \14443 , \14444 , \14445 , \14446 , \14447 , \14448 ,
         \14449 , \14450 , \14451 , \14452 , \14453 , \14454 , \14455 , \14456 , \14457 , \14458 ,
         \14459 , \14460 , \14461 , \14462 , \14463 , \14464 , \14465 , \14466 , \14467 , \14468 ,
         \14469 , \14470 , \14471 , \14472 , \14473 , \14474 , \14475 , \14476 , \14477 , \14478 ,
         \14479 , \14480 , \14481 , \14482 , \14483 , \14484 , \14485 , \14486 , \14487 , \14488 ,
         \14489 , \14490 , \14491 , \14492 , \14493 , \14494 , \14495 , \14496_nG5503 , \14497 , \14498 ,
         \14499 , \14500 , \14501 , \14502 , \14503 , \14504 , \14505 , \14506 , \14507 , \14508 ,
         \14509 , \14510 , \14511 , \14512 , \14513 , \14514 , \14515 , \14516 , \14517 , \14518 ,
         \14519 , \14520 , \14521 , \14522 , \14523 , \14524 , \14525 , \14526 , \14527 , \14528 ,
         \14529 , \14530 , \14531 , \14532 , \14533 , \14534 , \14535 , \14536 , \14537 , \14538 ,
         \14539 , \14540 , \14541 , \14542 , \14543 , \14544 , \14545 , \14546 , \14547 , \14548 ,
         \14549 , \14550 , \14551 , \14552 , \14553 , \14554 , \14555 , \14556 , \14557 , \14558 ,
         \14559 , \14560 , \14561 , \14562 , \14563 , \14564 , \14565 , \14566 , \14567 , \14568 ,
         \14569 , \14570 , \14571 , \14572 , \14573 , \14574 , \14575 , \14576 , \14577 , \14578 ,
         \14579 , \14580 , \14581 , \14582 , \14583 , \14584 , \14585 , \14586 , \14587 , \14588 ,
         \14589 , \14590 , \14591 , \14592 , \14593 , \14594 , \14595 , \14596 , \14597 , \14598 ,
         \14599 , \14600 , \14601 , \14602 , \14603 , \14604 , \14605 , \14606 , \14607 , \14608 ,
         \14609 , \14610 , \14611 , \14612 , \14613 , \14614 , \14615 , \14616 , \14617 , \14618 ,
         \14619 , \14620 , \14621 , \14622 , \14623 , \14624 , \14625 , \14626 , \14627 , \14628 ,
         \14629 , \14630 , \14631 , \14632 , \14633 , \14634 , \14635 , \14636 , \14637 , \14638 ,
         \14639 , \14640 , \14641 , \14642 , \14643 , \14644 , \14645 , \14646 , \14647 , \14648 ,
         \14649 , \14650 , \14651 , \14652 , \14653 , \14654 , \14655 , \14656 , \14657 , \14658 ,
         \14659 , \14660 , \14661 , \14662 , \14663 , \14664 , \14665 , \14666 , \14667 , \14668 ,
         \14669 , \14670 , \14671 , \14672 , \14673 , \14674 , \14675 , \14676 , \14677 , \14678 ,
         \14679 , \14680 , \14681 , \14682 , \14683 , \14684 , \14685 , \14686 , \14687 , \14688 ,
         \14689 , \14690 , \14691 , \14692 , \14693 , \14694 , \14695 , \14696 , \14697 , \14698 ,
         \14699 , \14700 , \14701 , \14702 , \14703 , \14704 , \14705 , \14706 , \14707 , \14708 ,
         \14709 , \14710 , \14711 , \14712 , \14713 , \14714 , \14715 , \14716 , \14717 , \14718 ,
         \14719 , \14720 , \14721 , \14722 , \14723 , \14724 , \14725 , \14726 , \14727 , \14728 ,
         \14729 , \14730 , \14731 , \14732 , \14733 , \14734 , \14735 , \14736 , \14737 , \14738 ,
         \14739 , \14740 , \14741 , \14742 , \14743 , \14744 , \14745 , \14746 , \14747 , \14748 ,
         \14749 , \14750 , \14751 , \14752 , \14753 , \14754 , \14755 , \14756 , \14757 , \14758 ,
         \14759 , \14760 , \14761 , \14762_nG5501 , \14763 , \14764 , \14765 , \14766 , \14767 , \14768 ,
         \14769 , \14770 , \14771 , \14772 , \14773 , \14774 , \14775 , \14776 , \14777 , \14778 ,
         \14779 , \14780 , \14781 , \14782 , \14783 , \14784 , \14785 , \14786 , \14787 , \14788 ,
         \14789 , \14790 , \14791 , \14792 , \14793 , \14794 , \14795 , \14796 , \14797 , \14798 ,
         \14799 , \14800 , \14801 , \14802 , \14803 , \14804 , \14805 , \14806 , \14807 , \14808 ,
         \14809 , \14810 , \14811 , \14812 , \14813 , \14814 , \14815 , \14816 , \14817 , \14818 ,
         \14819 , \14820 , \14821 , \14822 , \14823 , \14824 , \14825 , \14826 , \14827 , \14828 ,
         \14829 , \14830 , \14831 , \14832 , \14833 , \14834 , \14835 , \14836 , \14837 , \14838 ,
         \14839 , \14840 , \14841 , \14842 , \14843 , \14844 , \14845 , \14846 , \14847 , \14848 ,
         \14849 , \14850 , \14851 , \14852 , \14853 , \14854 , \14855 , \14856 , \14857 , \14858 ,
         \14859 , \14860 , \14861 , \14862 , \14863 , \14864 , \14865 , \14866 , \14867 , \14868 ,
         \14869 , \14870 , \14871 , \14872 , \14873 , \14874 , \14875 , \14876 , \14877 , \14878 ,
         \14879 , \14880 , \14881 , \14882 , \14883 , \14884 , \14885 , \14886 , \14887 , \14888 ,
         \14889 , \14890 , \14891 , \14892 , \14893 , \14894 , \14895 , \14896 , \14897 , \14898 ,
         \14899 , \14900 , \14901 , \14902 , \14903 , \14904 , \14905 , \14906 , \14907 , \14908 ,
         \14909 , \14910 , \14911 , \14912 , \14913 , \14914 , \14915 , \14916 , \14917 , \14918 ,
         \14919 , \14920 , \14921 , \14922 , \14923 , \14924 , \14925 , \14926 , \14927 , \14928 ,
         \14929 , \14930 , \14931 , \14932 , \14933 , \14934 , \14935 , \14936 , \14937 , \14938 ,
         \14939 , \14940 , \14941 , \14942 , \14943 , \14944 , \14945 , \14946 , \14947 , \14948 ,
         \14949 , \14950 , \14951 , \14952 , \14953 , \14954 , \14955 , \14956 , \14957 , \14958 ,
         \14959 , \14960 , \14961 , \14962 , \14963 , \14964 , \14965 , \14966 , \14967 , \14968 ,
         \14969 , \14970 , \14971 , \14972 , \14973 , \14974 , \14975 , \14976 , \14977 , \14978 ,
         \14979 , \14980 , \14981 , \14982 , \14983 , \14984 , \14985 , \14986 , \14987 , \14988 ,
         \14989 , \14990 , \14991 , \14992 , \14993 , \14994 , \14995 , \14996 , \14997 , \14998 ,
         \14999 , \15000 , \15001 , \15002 , \15003 , \15004 , \15005 , \15006 , \15007 , \15008 ,
         \15009 , \15010 , \15011 , \15012 , \15013 , \15014 , \15015 , \15016 , \15017 , \15018 ,
         \15019 , \15020 , \15021 , \15022_nG54ff , \15023 , \15024 , \15025 , \15026 , \15027 , \15028 ,
         \15029 , \15030 , \15031 , \15032 , \15033 , \15034 , \15035 , \15036 , \15037 , \15038 ,
         \15039 , \15040 , \15041 , \15042 , \15043 , \15044 , \15045 , \15046 , \15047 , \15048 ,
         \15049 , \15050 , \15051 , \15052 , \15053 , \15054 , \15055 , \15056 , \15057 , \15058 ,
         \15059 , \15060 , \15061 , \15062 , \15063 , \15064 , \15065 , \15066 , \15067 , \15068 ,
         \15069 , \15070 , \15071 , \15072 , \15073 , \15074 , \15075 , \15076 , \15077 , \15078 ,
         \15079 , \15080 , \15081 , \15082 , \15083 , \15084 , \15085 , \15086 , \15087 , \15088 ,
         \15089 , \15090 , \15091 , \15092 , \15093 , \15094 , \15095 , \15096 , \15097 , \15098 ,
         \15099 , \15100 , \15101 , \15102 , \15103 , \15104 , \15105 , \15106 , \15107 , \15108 ,
         \15109 , \15110 , \15111 , \15112 , \15113 , \15114 , \15115 , \15116 , \15117 , \15118 ,
         \15119 , \15120 , \15121 , \15122 , \15123 , \15124 , \15125 , \15126 , \15127 , \15128 ,
         \15129 , \15130 , \15131 , \15132 , \15133 , \15134 , \15135 , \15136 , \15137 , \15138 ,
         \15139 , \15140 , \15141 , \15142 , \15143 , \15144 , \15145 , \15146 , \15147 , \15148 ,
         \15149 , \15150 , \15151 , \15152 , \15153 , \15154 , \15155 , \15156 , \15157 , \15158 ,
         \15159 , \15160 , \15161 , \15162 , \15163 , \15164 , \15165 , \15166 , \15167 , \15168 ,
         \15169 , \15170 , \15171 , \15172 , \15173 , \15174 , \15175 , \15176 , \15177 , \15178 ,
         \15179 , \15180 , \15181 , \15182 , \15183 , \15184 , \15185 , \15186 , \15187 , \15188 ,
         \15189 , \15190 , \15191 , \15192 , \15193 , \15194 , \15195 , \15196 , \15197 , \15198 ,
         \15199 , \15200 , \15201 , \15202 , \15203 , \15204 , \15205 , \15206 , \15207 , \15208 ,
         \15209 , \15210 , \15211 , \15212 , \15213 , \15214 , \15215 , \15216 , \15217 , \15218 ,
         \15219 , \15220 , \15221 , \15222 , \15223 , \15224 , \15225 , \15226 , \15227 , \15228 ,
         \15229 , \15230 , \15231 , \15232 , \15233 , \15234 , \15235 , \15236 , \15237 , \15238 ,
         \15239 , \15240 , \15241 , \15242 , \15243 , \15244 , \15245 , \15246 , \15247 , \15248 ,
         \15249 , \15250 , \15251 , \15252 , \15253 , \15254 , \15255 , \15256 , \15257 , \15258 ,
         \15259 , \15260 , \15261 , \15262 , \15263 , \15264 , \15265 , \15266 , \15267 , \15268 ,
         \15269 , \15270 , \15271 , \15272 , \15273 , \15274 , \15275 , \15276 , \15277_nG54fd , \15278 ,
         \15279 , \15280 , \15281 , \15282 , \15283 , \15284 , \15285 , \15286 , \15287 , \15288 ,
         \15289 , \15290 , \15291 , \15292 , \15293 , \15294 , \15295 , \15296 , \15297 , \15298 ,
         \15299 , \15300 , \15301 , \15302 , \15303 , \15304 , \15305 , \15306 , \15307 , \15308 ,
         \15309 , \15310 , \15311 , \15312 , \15313 , \15314 , \15315 , \15316 , \15317 , \15318 ,
         \15319 , \15320 , \15321 , \15322 , \15323 , \15324 , \15325 , \15326 , \15327 , \15328 ,
         \15329 , \15330 , \15331 , \15332 , \15333 , \15334 , \15335 , \15336 , \15337 , \15338 ,
         \15339 , \15340 , \15341 , \15342 , \15343 , \15344 , \15345 , \15346 , \15347 , \15348 ,
         \15349 , \15350 , \15351 , \15352 , \15353 , \15354 , \15355 , \15356 , \15357 , \15358 ,
         \15359 , \15360 , \15361 , \15362 , \15363 , \15364 , \15365 , \15366 , \15367 , \15368 ,
         \15369 , \15370 , \15371 , \15372 , \15373 , \15374 , \15375 , \15376 , \15377 , \15378 ,
         \15379 , \15380 , \15381 , \15382 , \15383 , \15384 , \15385 , \15386 , \15387 , \15388 ,
         \15389 , \15390 , \15391 , \15392 , \15393 , \15394 , \15395 , \15396 , \15397 , \15398 ,
         \15399 , \15400 , \15401 , \15402 , \15403 , \15404 , \15405 , \15406 , \15407 , \15408 ,
         \15409 , \15410 , \15411 , \15412 , \15413 , \15414 , \15415 , \15416 , \15417 , \15418 ,
         \15419 , \15420 , \15421 , \15422 , \15423 , \15424 , \15425 , \15426 , \15427 , \15428 ,
         \15429 , \15430 , \15431 , \15432 , \15433 , \15434 , \15435 , \15436 , \15437 , \15438 ,
         \15439 , \15440 , \15441 , \15442 , \15443 , \15444 , \15445 , \15446 , \15447 , \15448 ,
         \15449 , \15450 , \15451 , \15452 , \15453 , \15454 , \15455 , \15456 , \15457 , \15458 ,
         \15459 , \15460 , \15461 , \15462 , \15463 , \15464 , \15465 , \15466 , \15467 , \15468 ,
         \15469 , \15470 , \15471 , \15472 , \15473 , \15474 , \15475 , \15476 , \15477 , \15478 ,
         \15479 , \15480 , \15481 , \15482 , \15483 , \15484 , \15485 , \15486 , \15487 , \15488 ,
         \15489 , \15490 , \15491 , \15492 , \15493 , \15494 , \15495 , \15496 , \15497 , \15498 ,
         \15499 , \15500 , \15501 , \15502 , \15503 , \15504 , \15505 , \15506 , \15507 , \15508 ,
         \15509 , \15510 , \15511 , \15512 , \15513 , \15514 , \15515 , \15516 , \15517 , \15518 ,
         \15519 , \15520 , \15521 , \15522 , \15523 , \15524 , \15525 , \15526 , \15527 , \15528 ,
         \15529 , \15530_nG54fb , \15531 , \15532 , \15533 , \15534 , \15535 , \15536 , \15537 , \15538 ,
         \15539 , \15540 , \15541 , \15542 , \15543 , \15544 , \15545 , \15546 , \15547 , \15548 ,
         \15549 , \15550 , \15551 , \15552 , \15553 , \15554 , \15555 , \15556 , \15557 , \15558 ,
         \15559 , \15560 , \15561 , \15562 , \15563 , \15564 , \15565 , \15566 , \15567 , \15568 ,
         \15569 , \15570 , \15571 , \15572 , \15573 , \15574 , \15575 , \15576 , \15577 , \15578 ,
         \15579 , \15580 , \15581 , \15582 , \15583 , \15584 , \15585 , \15586 , \15587 , \15588 ,
         \15589 , \15590 , \15591 , \15592 , \15593 , \15594 , \15595 , \15596 , \15597 , \15598 ,
         \15599 , \15600 , \15601 , \15602 , \15603 , \15604 , \15605 , \15606 , \15607 , \15608 ,
         \15609 , \15610 , \15611 , \15612 , \15613 , \15614 , \15615 , \15616 , \15617 , \15618 ,
         \15619 , \15620 , \15621 , \15622 , \15623 , \15624 , \15625 , \15626 , \15627 , \15628 ,
         \15629 , \15630 , \15631 , \15632 , \15633 , \15634 , \15635 , \15636 , \15637 , \15638 ,
         \15639 , \15640 , \15641 , \15642 , \15643 , \15644 , \15645 , \15646 , \15647 , \15648 ,
         \15649 , \15650 , \15651 , \15652 , \15653 , \15654 , \15655 , \15656 , \15657 , \15658 ,
         \15659 , \15660 , \15661 , \15662 , \15663 , \15664 , \15665 , \15666 , \15667 , \15668 ,
         \15669 , \15670 , \15671 , \15672 , \15673 , \15674 , \15675 , \15676 , \15677 , \15678 ,
         \15679 , \15680 , \15681 , \15682 , \15683 , \15684 , \15685 , \15686 , \15687 , \15688 ,
         \15689 , \15690 , \15691 , \15692 , \15693 , \15694 , \15695 , \15696 , \15697 , \15698 ,
         \15699 , \15700 , \15701 , \15702 , \15703 , \15704 , \15705 , \15706 , \15707 , \15708 ,
         \15709 , \15710 , \15711 , \15712 , \15713 , \15714 , \15715 , \15716 , \15717 , \15718 ,
         \15719 , \15720 , \15721 , \15722 , \15723 , \15724 , \15725 , \15726 , \15727 , \15728 ,
         \15729 , \15730 , \15731 , \15732 , \15733 , \15734 , \15735 , \15736 , \15737 , \15738 ,
         \15739 , \15740 , \15741 , \15742 , \15743 , \15744 , \15745 , \15746 , \15747 , \15748 ,
         \15749 , \15750 , \15751 , \15752 , \15753 , \15754 , \15755 , \15756 , \15757 , \15758 ,
         \15759 , \15760 , \15761 , \15762 , \15763 , \15764 , \15765 , \15766 , \15767 , \15768 ,
         \15769 , \15770 , \15771 , \15772 , \15773 , \15774 , \15775 , \15776 , \15777 , \15778 ,
         \15779 , \15780_nG54f9 , \15781 , \15782 , \15783 , \15784 , \15785 , \15786 , \15787 , \15788 ,
         \15789 , \15790 , \15791 , \15792 , \15793 , \15794 , \15795 , \15796 , \15797 , \15798 ,
         \15799 , \15800 , \15801 , \15802 , \15803 , \15804 , \15805 , \15806 , \15807 , \15808 ,
         \15809 , \15810 , \15811 , \15812 , \15813 , \15814 , \15815 , \15816 , \15817 , \15818 ,
         \15819 , \15820 , \15821 , \15822 , \15823 , \15824 , \15825 , \15826 , \15827 , \15828 ,
         \15829 , \15830 , \15831 , \15832 , \15833 , \15834 , \15835 , \15836 , \15837 , \15838 ,
         \15839 , \15840 , \15841 , \15842 , \15843 , \15844 , \15845 , \15846 , \15847 , \15848 ,
         \15849 , \15850 , \15851 , \15852 , \15853 , \15854 , \15855 , \15856 , \15857 , \15858 ,
         \15859 , \15860 , \15861 , \15862 , \15863 , \15864 , \15865 , \15866 , \15867 , \15868 ,
         \15869 , \15870 , \15871 , \15872 , \15873 , \15874 , \15875 , \15876 , \15877 , \15878 ,
         \15879 , \15880 , \15881 , \15882 , \15883 , \15884 , \15885 , \15886 , \15887 , \15888 ,
         \15889 , \15890 , \15891 , \15892 , \15893 , \15894 , \15895 , \15896 , \15897 , \15898 ,
         \15899 , \15900 , \15901 , \15902 , \15903 , \15904 , \15905 , \15906 , \15907 , \15908 ,
         \15909 , \15910 , \15911 , \15912 , \15913 , \15914 , \15915 , \15916 , \15917 , \15918 ,
         \15919 , \15920 , \15921 , \15922 , \15923 , \15924 , \15925 , \15926 , \15927 , \15928 ,
         \15929 , \15930 , \15931 , \15932 , \15933 , \15934 , \15935 , \15936 , \15937 , \15938 ,
         \15939 , \15940 , \15941 , \15942 , \15943 , \15944 , \15945 , \15946 , \15947 , \15948 ,
         \15949 , \15950 , \15951 , \15952 , \15953 , \15954 , \15955 , \15956 , \15957 , \15958 ,
         \15959 , \15960 , \15961 , \15962 , \15963 , \15964 , \15965 , \15966 , \15967 , \15968 ,
         \15969 , \15970 , \15971 , \15972 , \15973 , \15974 , \15975 , \15976 , \15977 , \15978 ,
         \15979 , \15980 , \15981 , \15982 , \15983 , \15984 , \15985 , \15986 , \15987 , \15988 ,
         \15989 , \15990 , \15991 , \15992 , \15993 , \15994 , \15995 , \15996 , \15997 , \15998 ,
         \15999 , \16000 , \16001 , \16002 , \16003 , \16004 , \16005 , \16006 , \16007 , \16008 ,
         \16009 , \16010 , \16011 , \16012 , \16013 , \16014 , \16015 , \16016 , \16017 , \16018 ,
         \16019 , \16020 , \16021 , \16022 , \16023 , \16024 , \16025 , \16026_nG54f7 , \16027 , \16028 ,
         \16029 , \16030 , \16031 , \16032 , \16033 , \16034 , \16035 , \16036 , \16037 , \16038 ,
         \16039 , \16040 , \16041 , \16042 , \16043 , \16044 , \16045 , \16046 , \16047 , \16048 ,
         \16049 , \16050 , \16051 , \16052 , \16053 , \16054 , \16055 , \16056 , \16057 , \16058 ,
         \16059 , \16060 , \16061 , \16062 , \16063 , \16064 , \16065 , \16066 , \16067 , \16068 ,
         \16069 , \16070 , \16071 , \16072 , \16073 , \16074 , \16075 , \16076 , \16077 , \16078 ,
         \16079 , \16080 , \16081 , \16082 , \16083 , \16084 , \16085 , \16086 , \16087 , \16088 ,
         \16089 , \16090 , \16091 , \16092 , \16093 , \16094 , \16095 , \16096 , \16097 , \16098 ,
         \16099 , \16100 , \16101 , \16102 , \16103 , \16104 , \16105 , \16106 , \16107 , \16108 ,
         \16109 , \16110 , \16111 , \16112 , \16113 , \16114 , \16115 , \16116 , \16117 , \16118 ,
         \16119 , \16120 , \16121 , \16122 , \16123 , \16124 , \16125 , \16126 , \16127 , \16128 ,
         \16129 , \16130 , \16131 , \16132 , \16133 , \16134 , \16135 , \16136 , \16137 , \16138 ,
         \16139 , \16140 , \16141 , \16142 , \16143 , \16144 , \16145 , \16146 , \16147 , \16148 ,
         \16149 , \16150 , \16151 , \16152 , \16153 , \16154 , \16155 , \16156 , \16157 , \16158 ,
         \16159 , \16160 , \16161 , \16162 , \16163 , \16164 , \16165 , \16166 , \16167 , \16168 ,
         \16169 , \16170 , \16171 , \16172 , \16173 , \16174 , \16175 , \16176 , \16177 , \16178 ,
         \16179 , \16180 , \16181 , \16182 , \16183 , \16184 , \16185 , \16186 , \16187 , \16188 ,
         \16189 , \16190 , \16191 , \16192 , \16193 , \16194 , \16195 , \16196 , \16197 , \16198 ,
         \16199 , \16200 , \16201 , \16202 , \16203 , \16204 , \16205 , \16206 , \16207 , \16208 ,
         \16209 , \16210 , \16211 , \16212 , \16213 , \16214 , \16215 , \16216 , \16217 , \16218 ,
         \16219 , \16220 , \16221 , \16222 , \16223 , \16224 , \16225 , \16226 , \16227 , \16228 ,
         \16229 , \16230 , \16231 , \16232 , \16233 , \16234 , \16235 , \16236 , \16237 , \16238 ,
         \16239 , \16240 , \16241 , \16242 , \16243 , \16244 , \16245 , \16246 , \16247 , \16248 ,
         \16249 , \16250 , \16251 , \16252 , \16253 , \16254 , \16255 , \16256 , \16257 , \16258 ,
         \16259 , \16260 , \16261 , \16262 , \16263_nG54f5 , \16264 , \16265 , \16266 , \16267 , \16268 ,
         \16269 , \16270 , \16271 , \16272 , \16273 , \16274 , \16275 , \16276 , \16277 , \16278 ,
         \16279 , \16280 , \16281 , \16282 , \16283 , \16284 , \16285 , \16286 , \16287 , \16288 ,
         \16289 , \16290 , \16291 , \16292 , \16293 , \16294 , \16295 , \16296 , \16297 , \16298 ,
         \16299 , \16300 , \16301 , \16302 , \16303 , \16304 , \16305 , \16306 , \16307 , \16308 ,
         \16309 , \16310 , \16311 , \16312 , \16313 , \16314 , \16315 , \16316 , \16317 , \16318 ,
         \16319 , \16320 , \16321 , \16322 , \16323 , \16324 , \16325 , \16326 , \16327 , \16328 ,
         \16329 , \16330 , \16331 , \16332 , \16333 , \16334 , \16335 , \16336 , \16337 , \16338 ,
         \16339 , \16340 , \16341 , \16342 , \16343 , \16344 , \16345 , \16346 , \16347 , \16348 ,
         \16349 , \16350 , \16351 , \16352 , \16353 , \16354 , \16355 , \16356 , \16357 , \16358 ,
         \16359 , \16360 , \16361 , \16362 , \16363 , \16364 , \16365 , \16366 , \16367 , \16368 ,
         \16369 , \16370 , \16371 , \16372 , \16373 , \16374 , \16375 , \16376 , \16377 , \16378 ,
         \16379 , \16380 , \16381 , \16382 , \16383 , \16384 , \16385 , \16386 , \16387 , \16388 ,
         \16389 , \16390 , \16391 , \16392 , \16393 , \16394 , \16395 , \16396 , \16397 , \16398 ,
         \16399 , \16400 , \16401 , \16402 , \16403 , \16404 , \16405 , \16406 , \16407 , \16408 ,
         \16409 , \16410 , \16411 , \16412 , \16413 , \16414 , \16415 , \16416 , \16417 , \16418 ,
         \16419 , \16420 , \16421 , \16422 , \16423 , \16424 , \16425 , \16426 , \16427 , \16428 ,
         \16429 , \16430 , \16431 , \16432 , \16433 , \16434 , \16435 , \16436 , \16437 , \16438 ,
         \16439 , \16440 , \16441 , \16442 , \16443 , \16444 , \16445 , \16446 , \16447 , \16448 ,
         \16449 , \16450 , \16451 , \16452 , \16453 , \16454 , \16455 , \16456 , \16457 , \16458 ,
         \16459 , \16460 , \16461 , \16462 , \16463 , \16464 , \16465 , \16466 , \16467 , \16468 ,
         \16469 , \16470 , \16471 , \16472 , \16473 , \16474 , \16475 , \16476 , \16477 , \16478 ,
         \16479 , \16480 , \16481 , \16482 , \16483 , \16484 , \16485 , \16486 , \16487 , \16488 ,
         \16489 , \16490 , \16491 , \16492 , \16493 , \16494 , \16495 , \16496 , \16497 , \16498_nG54f3 ,
         \16499 , \16500 , \16501 , \16502 , \16503 , \16504 , \16505 , \16506 , \16507 , \16508 ,
         \16509 , \16510 , \16511 , \16512 , \16513 , \16514 , \16515 , \16516 , \16517 , \16518 ,
         \16519 , \16520 , \16521 , \16522 , \16523 , \16524 , \16525 , \16526 , \16527 , \16528 ,
         \16529 , \16530 , \16531 , \16532 , \16533 , \16534 , \16535 , \16536 , \16537 , \16538 ,
         \16539 , \16540 , \16541 , \16542 , \16543 , \16544 , \16545 , \16546 , \16547 , \16548 ,
         \16549 , \16550 , \16551 , \16552 , \16553 , \16554 , \16555 , \16556 , \16557 , \16558 ,
         \16559 , \16560 , \16561 , \16562 , \16563 , \16564 , \16565 , \16566 , \16567 , \16568 ,
         \16569 , \16570 , \16571 , \16572 , \16573 , \16574 , \16575 , \16576 , \16577 , \16578 ,
         \16579 , \16580 , \16581 , \16582 , \16583 , \16584 , \16585 , \16586 , \16587 , \16588 ,
         \16589 , \16590 , \16591 , \16592 , \16593 , \16594 , \16595 , \16596 , \16597 , \16598 ,
         \16599 , \16600 , \16601 , \16602 , \16603 , \16604 , \16605 , \16606 , \16607 , \16608 ,
         \16609 , \16610 , \16611 , \16612 , \16613 , \16614 , \16615 , \16616 , \16617 , \16618 ,
         \16619 , \16620 , \16621 , \16622 , \16623 , \16624 , \16625 , \16626 , \16627 , \16628 ,
         \16629 , \16630 , \16631 , \16632 , \16633 , \16634 , \16635 , \16636 , \16637 , \16638 ,
         \16639 , \16640 , \16641 , \16642 , \16643 , \16644 , \16645 , \16646 , \16647 , \16648 ,
         \16649 , \16650 , \16651 , \16652 , \16653 , \16654 , \16655 , \16656 , \16657 , \16658 ,
         \16659 , \16660 , \16661 , \16662 , \16663 , \16664 , \16665 , \16666 , \16667 , \16668 ,
         \16669 , \16670 , \16671 , \16672 , \16673 , \16674 , \16675 , \16676 , \16677 , \16678 ,
         \16679 , \16680 , \16681 , \16682 , \16683 , \16684 , \16685 , \16686 , \16687 , \16688 ,
         \16689 , \16690 , \16691 , \16692 , \16693 , \16694 , \16695 , \16696 , \16697 , \16698 ,
         \16699 , \16700 , \16701 , \16702 , \16703 , \16704 , \16705 , \16706 , \16707 , \16708 ,
         \16709 , \16710 , \16711 , \16712 , \16713 , \16714 , \16715 , \16716 , \16717 , \16718 ,
         \16719 , \16720 , \16721 , \16722 , \16723 , \16724 , \16725 , \16726_nG54f1 , \16727 , \16728 ,
         \16729 , \16730 , \16731 , \16732 , \16733 , \16734 , \16735 , \16736 , \16737 , \16738 ,
         \16739 , \16740 , \16741 , \16742 , \16743 , \16744 , \16745 , \16746 , \16747 , \16748 ,
         \16749 , \16750 , \16751 , \16752 , \16753 , \16754 , \16755 , \16756 , \16757 , \16758 ,
         \16759 , \16760 , \16761 , \16762 , \16763 , \16764 , \16765 , \16766 , \16767 , \16768 ,
         \16769 , \16770 , \16771 , \16772 , \16773 , \16774 , \16775 , \16776 , \16777 , \16778 ,
         \16779 , \16780 , \16781 , \16782 , \16783 , \16784 , \16785 , \16786 , \16787 , \16788 ,
         \16789 , \16790 , \16791 , \16792 , \16793 , \16794 , \16795 , \16796 , \16797 , \16798 ,
         \16799 , \16800 , \16801 , \16802 , \16803 , \16804 , \16805 , \16806 , \16807 , \16808 ,
         \16809 , \16810 , \16811 , \16812 , \16813 , \16814 , \16815 , \16816 , \16817 , \16818 ,
         \16819 , \16820 , \16821 , \16822 , \16823 , \16824 , \16825 , \16826 , \16827 , \16828 ,
         \16829 , \16830 , \16831 , \16832 , \16833 , \16834 , \16835 , \16836 , \16837 , \16838 ,
         \16839 , \16840 , \16841 , \16842 , \16843 , \16844 , \16845 , \16846 , \16847 , \16848 ,
         \16849 , \16850 , \16851 , \16852 , \16853 , \16854 , \16855 , \16856 , \16857 , \16858 ,
         \16859 , \16860 , \16861 , \16862 , \16863 , \16864 , \16865 , \16866 , \16867 , \16868 ,
         \16869 , \16870 , \16871 , \16872 , \16873 , \16874 , \16875 , \16876 , \16877 , \16878 ,
         \16879 , \16880 , \16881 , \16882 , \16883 , \16884 , \16885 , \16886 , \16887 , \16888 ,
         \16889 , \16890 , \16891 , \16892 , \16893 , \16894 , \16895 , \16896 , \16897 , \16898 ,
         \16899 , \16900 , \16901 , \16902 , \16903 , \16904 , \16905 , \16906 , \16907 , \16908 ,
         \16909 , \16910 , \16911 , \16912 , \16913 , \16914 , \16915 , \16916 , \16917 , \16918 ,
         \16919 , \16920 , \16921 , \16922 , \16923 , \16924 , \16925 , \16926 , \16927 , \16928 ,
         \16929 , \16930 , \16931 , \16932 , \16933 , \16934 , \16935 , \16936 , \16937 , \16938 ,
         \16939 , \16940 , \16941 , \16942 , \16943 , \16944 , \16945 , \16946 , \16947 , \16948 ,
         \16949 , \16950_nG54ef , \16951 , \16952 , \16953 , \16954 , \16955 , \16956 , \16957 , \16958 ,
         \16959 , \16960 , \16961 , \16962 , \16963 , \16964 , \16965 , \16966 , \16967 , \16968 ,
         \16969 , \16970 , \16971 , \16972 , \16973 , \16974 , \16975 , \16976 , \16977 , \16978 ,
         \16979 , \16980 , \16981 , \16982 , \16983 , \16984 , \16985 , \16986 , \16987 , \16988 ,
         \16989 , \16990 , \16991 , \16992 , \16993 , \16994 , \16995 , \16996 , \16997 , \16998 ,
         \16999 , \17000 , \17001 , \17002 , \17003 , \17004 , \17005 , \17006 , \17007 , \17008 ,
         \17009 , \17010 , \17011 , \17012 , \17013 , \17014 , \17015 , \17016 , \17017 , \17018 ,
         \17019 , \17020 , \17021 , \17022 , \17023 , \17024 , \17025 , \17026 , \17027 , \17028 ,
         \17029 , \17030 , \17031 , \17032 , \17033 , \17034 , \17035 , \17036 , \17037 , \17038 ,
         \17039 , \17040 , \17041 , \17042 , \17043 , \17044 , \17045 , \17046 , \17047 , \17048 ,
         \17049 , \17050 , \17051 , \17052 , \17053 , \17054 , \17055 , \17056 , \17057 , \17058 ,
         \17059 , \17060 , \17061 , \17062 , \17063 , \17064 , \17065 , \17066 , \17067 , \17068 ,
         \17069 , \17070 , \17071 , \17072 , \17073 , \17074 , \17075 , \17076 , \17077 , \17078 ,
         \17079 , \17080 , \17081 , \17082 , \17083 , \17084 , \17085 , \17086 , \17087 , \17088 ,
         \17089 , \17090 , \17091 , \17092 , \17093 , \17094 , \17095 , \17096 , \17097 , \17098 ,
         \17099 , \17100 , \17101 , \17102 , \17103 , \17104 , \17105 , \17106 , \17107 , \17108 ,
         \17109 , \17110 , \17111 , \17112 , \17113 , \17114 , \17115 , \17116 , \17117 , \17118 ,
         \17119 , \17120 , \17121 , \17122 , \17123 , \17124 , \17125 , \17126 , \17127 , \17128 ,
         \17129 , \17130 , \17131 , \17132 , \17133 , \17134 , \17135 , \17136 , \17137 , \17138 ,
         \17139 , \17140 , \17141 , \17142 , \17143 , \17144 , \17145 , \17146 , \17147 , \17148 ,
         \17149 , \17150 , \17151 , \17152 , \17153 , \17154 , \17155 , \17156 , \17157 , \17158 ,
         \17159 , \17160 , \17161 , \17162 , \17163 , \17164 , \17165 , \17166 , \17167 , \17168_nG54ed ,
         \17169 , \17170 , \17171 , \17172 , \17173 , \17174 , \17175 , \17176 , \17177 , \17178 ,
         \17179 , \17180 , \17181 , \17182 , \17183 , \17184 , \17185 , \17186 , \17187 , \17188 ,
         \17189 , \17190 , \17191 , \17192 , \17193 , \17194 , \17195 , \17196 , \17197 , \17198 ,
         \17199 , \17200 , \17201 , \17202 , \17203 , \17204 , \17205 , \17206 , \17207 , \17208 ,
         \17209 , \17210 , \17211 , \17212 , \17213 , \17214 , \17215 , \17216 , \17217 , \17218 ,
         \17219 , \17220 , \17221 , \17222 , \17223 , \17224 , \17225 , \17226 , \17227 , \17228 ,
         \17229 , \17230 , \17231 , \17232 , \17233 , \17234 , \17235 , \17236 , \17237 , \17238 ,
         \17239 , \17240 , \17241 , \17242 , \17243 , \17244 , \17245 , \17246 , \17247 , \17248 ,
         \17249 , \17250 , \17251 , \17252 , \17253 , \17254 , \17255 , \17256 , \17257 , \17258 ,
         \17259 , \17260 , \17261 , \17262 , \17263 , \17264 , \17265 , \17266 , \17267 , \17268 ,
         \17269 , \17270 , \17271 , \17272 , \17273 , \17274 , \17275 , \17276 , \17277 , \17278 ,
         \17279 , \17280 , \17281 , \17282 , \17283 , \17284 , \17285 , \17286 , \17287 , \17288 ,
         \17289 , \17290 , \17291 , \17292 , \17293 , \17294 , \17295 , \17296 , \17297 , \17298 ,
         \17299 , \17300 , \17301 , \17302 , \17303 , \17304 , \17305 , \17306 , \17307 , \17308 ,
         \17309 , \17310 , \17311 , \17312 , \17313 , \17314 , \17315 , \17316 , \17317 , \17318 ,
         \17319 , \17320 , \17321 , \17322 , \17323 , \17324 , \17325 , \17326 , \17327 , \17328 ,
         \17329 , \17330 , \17331 , \17332 , \17333 , \17334 , \17335 , \17336 , \17337 , \17338 ,
         \17339 , \17340 , \17341 , \17342 , \17343 , \17344 , \17345 , \17346 , \17347 , \17348 ,
         \17349 , \17350 , \17351 , \17352 , \17353 , \17354 , \17355 , \17356 , \17357 , \17358 ,
         \17359 , \17360 , \17361 , \17362 , \17363 , \17364 , \17365 , \17366 , \17367 , \17368 ,
         \17369 , \17370 , \17371 , \17372 , \17373 , \17374 , \17375 , \17376 , \17377 , \17378 ,
         \17379 , \17380 , \17381_nG54eb , \17382 , \17383 , \17384 , \17385 , \17386 , \17387 , \17388 ,
         \17389 , \17390 , \17391 , \17392 , \17393 , \17394 , \17395 , \17396 , \17397 , \17398 ,
         \17399 , \17400 , \17401 , \17402 , \17403 , \17404 , \17405 , \17406 , \17407 , \17408 ,
         \17409 , \17410 , \17411 , \17412 , \17413 , \17414 , \17415 , \17416 , \17417 , \17418 ,
         \17419 , \17420 , \17421 , \17422 , \17423 , \17424 , \17425 , \17426 , \17427 , \17428 ,
         \17429 , \17430 , \17431 , \17432 , \17433 , \17434 , \17435 , \17436 , \17437 , \17438 ,
         \17439 , \17440 , \17441 , \17442 , \17443 , \17444 , \17445 , \17446 , \17447 , \17448 ,
         \17449 , \17450 , \17451 , \17452 , \17453 , \17454 , \17455 , \17456 , \17457 , \17458 ,
         \17459 , \17460 , \17461 , \17462 , \17463 , \17464 , \17465 , \17466 , \17467 , \17468 ,
         \17469 , \17470 , \17471 , \17472 , \17473 , \17474 , \17475 , \17476 , \17477 , \17478 ,
         \17479 , \17480 , \17481 , \17482 , \17483 , \17484 , \17485 , \17486 , \17487 , \17488 ,
         \17489 , \17490 , \17491 , \17492 , \17493 , \17494 , \17495 , \17496 , \17497 , \17498 ,
         \17499 , \17500 , \17501 , \17502 , \17503 , \17504 , \17505 , \17506 , \17507 , \17508 ,
         \17509 , \17510 , \17511 , \17512 , \17513 , \17514 , \17515 , \17516 , \17517 , \17518 ,
         \17519 , \17520 , \17521 , \17522 , \17523 , \17524 , \17525 , \17526 , \17527 , \17528 ,
         \17529 , \17530 , \17531 , \17532 , \17533 , \17534 , \17535 , \17536 , \17537 , \17538 ,
         \17539 , \17540 , \17541 , \17542 , \17543 , \17544 , \17545 , \17546 , \17547 , \17548 ,
         \17549 , \17550 , \17551 , \17552 , \17553 , \17554 , \17555 , \17556 , \17557 , \17558 ,
         \17559 , \17560 , \17561 , \17562 , \17563 , \17564 , \17565 , \17566 , \17567 , \17568 ,
         \17569 , \17570 , \17571 , \17572 , \17573 , \17574 , \17575 , \17576 , \17577 , \17578 ,
         \17579 , \17580 , \17581 , \17582 , \17583 , \17584 , \17585 , \17586_nG54e9 , \17587 , \17588 ,
         \17589 , \17590 , \17591 , \17592 , \17593 , \17594 , \17595 , \17596 , \17597 , \17598 ,
         \17599 , \17600 , \17601 , \17602 , \17603 , \17604 , \17605 , \17606 , \17607 , \17608 ,
         \17609 , \17610 , \17611 , \17612 , \17613 , \17614 , \17615 , \17616 , \17617 , \17618 ,
         \17619 , \17620 , \17621 , \17622 , \17623 , \17624 , \17625 , \17626 , \17627 , \17628 ,
         \17629 , \17630 , \17631 , \17632 , \17633 , \17634 , \17635 , \17636 , \17637 , \17638 ,
         \17639 , \17640 , \17641 , \17642 , \17643 , \17644 , \17645 , \17646 , \17647 , \17648 ,
         \17649 , \17650 , \17651 , \17652 , \17653 , \17654 , \17655 , \17656 , \17657 , \17658 ,
         \17659 , \17660 , \17661 , \17662 , \17663 , \17664 , \17665 , \17666 , \17667 , \17668 ,
         \17669 , \17670 , \17671 , \17672 , \17673 , \17674 , \17675 , \17676 , \17677 , \17678 ,
         \17679 , \17680 , \17681 , \17682 , \17683 , \17684 , \17685 , \17686 , \17687 , \17688 ,
         \17689 , \17690 , \17691 , \17692 , \17693 , \17694 , \17695 , \17696 , \17697 , \17698 ,
         \17699 , \17700 , \17701 , \17702 , \17703 , \17704 , \17705 , \17706 , \17707 , \17708 ,
         \17709 , \17710 , \17711 , \17712 , \17713 , \17714 , \17715 , \17716 , \17717 , \17718 ,
         \17719 , \17720 , \17721 , \17722 , \17723 , \17724 , \17725 , \17726 , \17727 , \17728 ,
         \17729 , \17730 , \17731 , \17732 , \17733 , \17734 , \17735 , \17736 , \17737 , \17738 ,
         \17739 , \17740 , \17741 , \17742 , \17743 , \17744 , \17745 , \17746 , \17747 , \17748 ,
         \17749 , \17750 , \17751 , \17752 , \17753 , \17754 , \17755 , \17756 , \17757 , \17758 ,
         \17759 , \17760 , \17761 , \17762 , \17763 , \17764 , \17765 , \17766 , \17767 , \17768 ,
         \17769 , \17770 , \17771 , \17772 , \17773 , \17774 , \17775 , \17776 , \17777 , \17778 ,
         \17779 , \17780 , \17781 , \17782 , \17783 , \17784 , \17785 , \17786 , \17787 , \17788 ,
         \17789_nG54e7 , \17790 , \17791 , \17792 , \17793 , \17794 , \17795 , \17796 , \17797 , \17798 ,
         \17799 , \17800 , \17801 , \17802 , \17803 , \17804 , \17805 , \17806 , \17807 , \17808 ,
         \17809 , \17810 , \17811 , \17812 , \17813 , \17814 , \17815 , \17816 , \17817 , \17818 ,
         \17819 , \17820 , \17821 , \17822 , \17823 , \17824 , \17825 , \17826 , \17827 , \17828 ,
         \17829 , \17830 , \17831 , \17832 , \17833 , \17834 , \17835 , \17836 , \17837 , \17838 ,
         \17839 , \17840 , \17841 , \17842 , \17843 , \17844 , \17845 , \17846 , \17847 , \17848 ,
         \17849 , \17850 , \17851 , \17852 , \17853 , \17854 , \17855 , \17856 , \17857 , \17858 ,
         \17859 , \17860 , \17861 , \17862 , \17863 , \17864 , \17865 , \17866 , \17867 , \17868 ,
         \17869 , \17870 , \17871 , \17872 , \17873 , \17874 , \17875 , \17876 , \17877 , \17878 ,
         \17879 , \17880 , \17881 , \17882 , \17883 , \17884 , \17885 , \17886 , \17887 , \17888 ,
         \17889 , \17890 , \17891 , \17892 , \17893 , \17894 , \17895 , \17896 , \17897 , \17898 ,
         \17899 , \17900 , \17901 , \17902 , \17903 , \17904 , \17905 , \17906 , \17907 , \17908 ,
         \17909 , \17910 , \17911 , \17912 , \17913 , \17914 , \17915 , \17916 , \17917 , \17918 ,
         \17919 , \17920 , \17921 , \17922 , \17923 , \17924 , \17925 , \17926 , \17927 , \17928 ,
         \17929 , \17930 , \17931 , \17932 , \17933 , \17934 , \17935 , \17936 , \17937 , \17938 ,
         \17939 , \17940 , \17941 , \17942 , \17943 , \17944 , \17945 , \17946 , \17947 , \17948 ,
         \17949 , \17950 , \17951 , \17952 , \17953 , \17954 , \17955 , \17956 , \17957 , \17958 ,
         \17959 , \17960 , \17961 , \17962 , \17963 , \17964 , \17965 , \17966 , \17967 , \17968 ,
         \17969 , \17970 , \17971 , \17972 , \17973 , \17974 , \17975 , \17976 , \17977 , \17978 ,
         \17979 , \17980 , \17981 , \17982 , \17983 , \17984_nG54e5 , \17985 , \17986 , \17987 , \17988 ,
         \17989 , \17990 , \17991 , \17992 , \17993 , \17994 , \17995 , \17996 , \17997 , \17998 ,
         \17999 , \18000 , \18001 , \18002 , \18003 , \18004 , \18005 , \18006 , \18007 , \18008 ,
         \18009 , \18010 , \18011 , \18012 , \18013 , \18014 , \18015 , \18016 , \18017 , \18018 ,
         \18019 , \18020 , \18021 , \18022 , \18023 , \18024 , \18025 , \18026 , \18027 , \18028 ,
         \18029 , \18030 , \18031 , \18032 , \18033 , \18034 , \18035 , \18036 , \18037 , \18038 ,
         \18039 , \18040 , \18041 , \18042 , \18043 , \18044 , \18045 , \18046 , \18047 , \18048 ,
         \18049 , \18050 , \18051 , \18052 , \18053 , \18054 , \18055 , \18056 , \18057 , \18058 ,
         \18059 , \18060 , \18061 , \18062 , \18063 , \18064 , \18065 , \18066 , \18067 , \18068 ,
         \18069 , \18070 , \18071 , \18072 , \18073 , \18074 , \18075 , \18076 , \18077 , \18078 ,
         \18079 , \18080 , \18081 , \18082 , \18083 , \18084 , \18085 , \18086 , \18087 , \18088 ,
         \18089 , \18090 , \18091 , \18092 , \18093 , \18094 , \18095 , \18096 , \18097 , \18098 ,
         \18099 , \18100 , \18101 , \18102 , \18103 , \18104 , \18105 , \18106 , \18107 , \18108 ,
         \18109 , \18110 , \18111 , \18112 , \18113 , \18114 , \18115 , \18116 , \18117 , \18118 ,
         \18119 , \18120 , \18121 , \18122 , \18123 , \18124 , \18125 , \18126 , \18127 , \18128 ,
         \18129 , \18130 , \18131 , \18132 , \18133 , \18134 , \18135 , \18136 , \18137 , \18138 ,
         \18139 , \18140 , \18141 , \18142 , \18143 , \18144 , \18145 , \18146 , \18147 , \18148 ,
         \18149 , \18150 , \18151 , \18152 , \18153 , \18154 , \18155 , \18156 , \18157 , \18158 ,
         \18159 , \18160 , \18161 , \18162 , \18163 , \18164 , \18165 , \18166 , \18167 , \18168 ,
         \18169 , \18170 , \18171 , \18172 , \18173 , \18174 , \18175 , \18176 , \18177_nG54e3 , \18178 ,
         \18179 , \18180 , \18181 , \18182 , \18183 , \18184 , \18185 , \18186 , \18187 , \18188 ,
         \18189 , \18190 , \18191 , \18192 , \18193 , \18194 , \18195 , \18196 , \18197 , \18198 ,
         \18199 , \18200 , \18201 , \18202 , \18203 , \18204 , \18205 , \18206 , \18207 , \18208 ,
         \18209 , \18210 , \18211 , \18212 , \18213 , \18214 , \18215 , \18216 , \18217 , \18218 ,
         \18219 , \18220 , \18221 , \18222 , \18223 , \18224 , \18225 , \18226 , \18227 , \18228 ,
         \18229 , \18230 , \18231 , \18232 , \18233 , \18234 , \18235 , \18236 , \18237 , \18238 ,
         \18239 , \18240 , \18241 , \18242 , \18243 , \18244 , \18245 , \18246 , \18247 , \18248 ,
         \18249 , \18250 , \18251 , \18252 , \18253 , \18254 , \18255 , \18256 , \18257 , \18258 ,
         \18259 , \18260 , \18261 , \18262 , \18263 , \18264 , \18265 , \18266 , \18267 , \18268 ,
         \18269 , \18270 , \18271 , \18272 , \18273 , \18274 , \18275 , \18276 , \18277 , \18278 ,
         \18279 , \18280 , \18281 , \18282 , \18283 , \18284 , \18285 , \18286 , \18287 , \18288 ,
         \18289 , \18290 , \18291 , \18292 , \18293 , \18294 , \18295 , \18296 , \18297 , \18298 ,
         \18299 , \18300 , \18301 , \18302 , \18303 , \18304 , \18305 , \18306 , \18307 , \18308 ,
         \18309 , \18310 , \18311 , \18312 , \18313 , \18314 , \18315 , \18316 , \18317 , \18318 ,
         \18319 , \18320 , \18321 , \18322 , \18323 , \18324 , \18325 , \18326 , \18327 , \18328 ,
         \18329 , \18330 , \18331 , \18332 , \18333 , \18334 , \18335 , \18336 , \18337 , \18338 ,
         \18339 , \18340 , \18341 , \18342 , \18343 , \18344 , \18345 , \18346 , \18347 , \18348 ,
         \18349 , \18350 , \18351 , \18352 , \18353 , \18354 , \18355 , \18356 , \18357 , \18358 ,
         \18359 , \18360 , \18361 , \18362 , \18363_nG54e1 , \18364 , \18365 , \18366 , \18367 , \18368 ,
         \18369 , \18370 , \18371 , \18372 , \18373 , \18374 , \18375 , \18376 , \18377 , \18378 ,
         \18379 , \18380 , \18381 , \18382 , \18383 , \18384 , \18385 , \18386 , \18387 , \18388 ,
         \18389 , \18390 , \18391 , \18392 , \18393 , \18394 , \18395 , \18396 , \18397 , \18398 ,
         \18399 , \18400 , \18401 , \18402 , \18403 , \18404 , \18405 , \18406 , \18407 , \18408 ,
         \18409 , \18410 , \18411 , \18412 , \18413 , \18414 , \18415 , \18416 , \18417 , \18418 ,
         \18419 , \18420 , \18421 , \18422 , \18423 , \18424 , \18425 , \18426 , \18427 , \18428 ,
         \18429 , \18430 , \18431 , \18432 , \18433 , \18434 , \18435 , \18436 , \18437 , \18438 ,
         \18439 , \18440 , \18441 , \18442 , \18443 , \18444 , \18445 , \18446 , \18447 , \18448 ,
         \18449 , \18450 , \18451 , \18452 , \18453 , \18454 , \18455 , \18456 , \18457 , \18458 ,
         \18459 , \18460 , \18461 , \18462 , \18463 , \18464 , \18465 , \18466 , \18467 , \18468 ,
         \18469 , \18470 , \18471 , \18472 , \18473 , \18474 , \18475 , \18476 , \18477 , \18478 ,
         \18479 , \18480 , \18481 , \18482 , \18483 , \18484 , \18485 , \18486 , \18487 , \18488 ,
         \18489 , \18490 , \18491 , \18492 , \18493 , \18494 , \18495 , \18496 , \18497 , \18498 ,
         \18499 , \18500 , \18501 , \18502 , \18503 , \18504 , \18505 , \18506 , \18507 , \18508 ,
         \18509 , \18510 , \18511 , \18512 , \18513 , \18514 , \18515 , \18516 , \18517 , \18518 ,
         \18519 , \18520 , \18521 , \18522 , \18523 , \18524 , \18525 , \18526 , \18527 , \18528 ,
         \18529 , \18530 , \18531 , \18532 , \18533 , \18534 , \18535 , \18536 , \18537 , \18538 ,
         \18539 , \18540 , \18541 , \18542 , \18543 , \18544_nG54df , \18545 , \18546 , \18547 , \18548 ,
         \18549 , \18550 , \18551 , \18552 , \18553 , \18554 , \18555 , \18556 , \18557 , \18558 ,
         \18559 , \18560 , \18561 , \18562 , \18563 , \18564 , \18565 , \18566 , \18567 , \18568 ,
         \18569 , \18570 , \18571 , \18572 , \18573 , \18574 , \18575 , \18576 , \18577 , \18578 ,
         \18579 , \18580 , \18581 , \18582 , \18583 , \18584 , \18585 , \18586 , \18587 , \18588 ,
         \18589 , \18590 , \18591 , \18592 , \18593 , \18594 , \18595 , \18596 , \18597 , \18598 ,
         \18599 , \18600 , \18601 , \18602 , \18603 , \18604 , \18605 , \18606 , \18607 , \18608 ,
         \18609 , \18610 , \18611 , \18612 , \18613 , \18614 , \18615 , \18616 , \18617 , \18618 ,
         \18619 , \18620 , \18621 , \18622 , \18623 , \18624 , \18625 , \18626 , \18627 , \18628 ,
         \18629 , \18630 , \18631 , \18632 , \18633 , \18634 , \18635 , \18636 , \18637 , \18638 ,
         \18639 , \18640 , \18641 , \18642 , \18643 , \18644 , \18645 , \18646 , \18647 , \18648 ,
         \18649 , \18650 , \18651 , \18652 , \18653 , \18654 , \18655 , \18656 , \18657 , \18658 ,
         \18659 , \18660 , \18661 , \18662 , \18663 , \18664 , \18665 , \18666 , \18667 , \18668 ,
         \18669 , \18670 , \18671 , \18672 , \18673 , \18674 , \18675 , \18676 , \18677 , \18678 ,
         \18679 , \18680 , \18681 , \18682 , \18683 , \18684 , \18685 , \18686 , \18687 , \18688 ,
         \18689 , \18690 , \18691 , \18692 , \18693 , \18694 , \18695 , \18696 , \18697 , \18698 ,
         \18699 , \18700 , \18701 , \18702 , \18703 , \18704 , \18705 , \18706 , \18707 , \18708 ,
         \18709 , \18710 , \18711 , \18712 , \18713 , \18714 , \18715 , \18716 , \18717_nG54dd , \18718 ,
         \18719 , \18720 , \18721 , \18722 , \18723 , \18724 , \18725 , \18726 , \18727 , \18728 ,
         \18729 , \18730 , \18731 , \18732 , \18733 , \18734 , \18735 , \18736 , \18737 , \18738 ,
         \18739 , \18740 , \18741 , \18742 , \18743 , \18744 , \18745 , \18746 , \18747 , \18748 ,
         \18749 , \18750 , \18751 , \18752 , \18753 , \18754 , \18755 , \18756 , \18757 , \18758 ,
         \18759 , \18760 , \18761 , \18762 , \18763 , \18764 , \18765 , \18766 , \18767 , \18768 ,
         \18769 , \18770 , \18771 , \18772 , \18773 , \18774 , \18775 , \18776 , \18777 , \18778 ,
         \18779 , \18780 , \18781 , \18782 , \18783 , \18784 , \18785 , \18786 , \18787 , \18788 ,
         \18789 , \18790 , \18791 , \18792 , \18793 , \18794 , \18795 , \18796 , \18797 , \18798 ,
         \18799 , \18800 , \18801 , \18802 , \18803 , \18804 , \18805 , \18806 , \18807 , \18808 ,
         \18809 , \18810 , \18811 , \18812 , \18813 , \18814 , \18815 , \18816 , \18817 , \18818 ,
         \18819 , \18820 , \18821 , \18822 , \18823 , \18824 , \18825 , \18826 , \18827 , \18828 ,
         \18829 , \18830 , \18831 , \18832 , \18833 , \18834 , \18835 , \18836 , \18837 , \18838 ,
         \18839 , \18840 , \18841 , \18842 , \18843 , \18844 , \18845 , \18846 , \18847 , \18848 ,
         \18849 , \18850 , \18851 , \18852 , \18853 , \18854 , \18855 , \18856 , \18857 , \18858 ,
         \18859 , \18860 , \18861 , \18862 , \18863 , \18864 , \18865 , \18866 , \18867 , \18868 ,
         \18869 , \18870 , \18871 , \18872 , \18873 , \18874 , \18875 , \18876 , \18877 , \18878 ,
         \18879 , \18880 , \18881 , \18882 , \18883 , \18884 , \18885 , \18886 , \18887_nG54db , \18888 ,
         \18889 , \18890 , \18891 , \18892 , \18893 , \18894 , \18895 , \18896 , \18897 , \18898 ,
         \18899 , \18900 , \18901 , \18902 , \18903 , \18904 , \18905 , \18906 , \18907 , \18908 ,
         \18909 , \18910 , \18911 , \18912 , \18913 , \18914 , \18915 , \18916 , \18917 , \18918 ,
         \18919 , \18920 , \18921 , \18922 , \18923 , \18924 , \18925 , \18926 , \18927 , \18928 ,
         \18929 , \18930 , \18931 , \18932 , \18933 , \18934 , \18935 , \18936 , \18937 , \18938 ,
         \18939 , \18940 , \18941 , \18942 , \18943 , \18944 , \18945 , \18946 , \18947 , \18948 ,
         \18949 , \18950 , \18951 , \18952 , \18953 , \18954 , \18955 , \18956 , \18957 , \18958 ,
         \18959 , \18960 , \18961 , \18962 , \18963 , \18964 , \18965 , \18966 , \18967 , \18968 ,
         \18969 , \18970 , \18971 , \18972 , \18973 , \18974 , \18975 , \18976 , \18977 , \18978 ,
         \18979 , \18980 , \18981 , \18982 , \18983 , \18984 , \18985 , \18986 , \18987 , \18988 ,
         \18989 , \18990 , \18991 , \18992 , \18993 , \18994 , \18995 , \18996 , \18997 , \18998 ,
         \18999 , \19000 , \19001 , \19002 , \19003 , \19004 , \19005 , \19006 , \19007 , \19008 ,
         \19009 , \19010 , \19011 , \19012 , \19013 , \19014 , \19015 , \19016 , \19017 , \19018 ,
         \19019 , \19020 , \19021 , \19022 , \19023 , \19024 , \19025 , \19026 , \19027 , \19028 ,
         \19029 , \19030 , \19031 , \19032 , \19033 , \19034 , \19035 , \19036 , \19037 , \19038 ,
         \19039 , \19040 , \19041 , \19042 , \19043 , \19044 , \19045 , \19046 , \19047 , \19048 ,
         \19049 , \19050 , \19051 , \19052_nG54d9 , \19053 , \19054 , \19055 , \19056 , \19057 , \19058 ,
         \19059 , \19060 , \19061 , \19062 , \19063 , \19064 , \19065 , \19066 , \19067 , \19068 ,
         \19069 , \19070 , \19071 , \19072 , \19073 , \19074 , \19075 , \19076 , \19077 , \19078 ,
         \19079 , \19080 , \19081 , \19082 , \19083 , \19084 , \19085 , \19086 , \19087 , \19088 ,
         \19089 , \19090 , \19091 , \19092 , \19093 , \19094 , \19095 , \19096 , \19097 , \19098 ,
         \19099 , \19100 , \19101 , \19102 , \19103 , \19104 , \19105 , \19106 , \19107 , \19108 ,
         \19109 , \19110 , \19111 , \19112 , \19113 , \19114 , \19115 , \19116 , \19117 , \19118 ,
         \19119 , \19120 , \19121 , \19122 , \19123 , \19124 , \19125 , \19126 , \19127 , \19128 ,
         \19129 , \19130 , \19131 , \19132 , \19133 , \19134 , \19135 , \19136 , \19137 , \19138 ,
         \19139 , \19140 , \19141 , \19142 , \19143 , \19144 , \19145 , \19146 , \19147 , \19148 ,
         \19149 , \19150 , \19151 , \19152 , \19153 , \19154 , \19155 , \19156 , \19157 , \19158 ,
         \19159 , \19160 , \19161 , \19162 , \19163 , \19164 , \19165 , \19166 , \19167 , \19168 ,
         \19169 , \19170 , \19171 , \19172 , \19173 , \19174 , \19175 , \19176 , \19177 , \19178 ,
         \19179 , \19180 , \19181 , \19182 , \19183 , \19184 , \19185 , \19186 , \19187 , \19188 ,
         \19189 , \19190 , \19191 , \19192 , \19193 , \19194 , \19195 , \19196 , \19197 , \19198 ,
         \19199 , \19200 , \19201 , \19202 , \19203 , \19204 , \19205 , \19206 , \19207 , \19208 ,
         \19209 , \19210 , \19211 , \19212 , \19213 , \19214 , \19215_nG54d7 , \19216 , \19217 , \19218 ,
         \19219 , \19220 , \19221 , \19222 , \19223 , \19224 , \19225 , \19226 , \19227 , \19228 ,
         \19229 , \19230 , \19231 , \19232 , \19233 , \19234 , \19235 , \19236 , \19237 , \19238 ,
         \19239 , \19240 , \19241 , \19242 , \19243 , \19244 , \19245 , \19246 , \19247 , \19248 ,
         \19249 , \19250 , \19251 , \19252 , \19253 , \19254 , \19255 , \19256 , \19257 , \19258 ,
         \19259 , \19260 , \19261 , \19262 , \19263 , \19264 , \19265 , \19266 , \19267 , \19268 ,
         \19269 , \19270 , \19271 , \19272 , \19273 , \19274 , \19275 , \19276 , \19277 , \19278 ,
         \19279 , \19280 , \19281 , \19282 , \19283 , \19284 , \19285 , \19286 , \19287 , \19288 ,
         \19289 , \19290 , \19291 , \19292 , \19293 , \19294 , \19295 , \19296 , \19297 , \19298 ,
         \19299 , \19300 , \19301 , \19302 , \19303 , \19304 , \19305 , \19306 , \19307 , \19308 ,
         \19309 , \19310 , \19311 , \19312 , \19313 , \19314 , \19315 , \19316 , \19317 , \19318 ,
         \19319 , \19320 , \19321 , \19322 , \19323 , \19324 , \19325 , \19326 , \19327 , \19328 ,
         \19329 , \19330 , \19331 , \19332 , \19333 , \19334 , \19335 , \19336 , \19337 , \19338 ,
         \19339 , \19340 , \19341 , \19342 , \19343 , \19344 , \19345 , \19346 , \19347 , \19348 ,
         \19349 , \19350 , \19351 , \19352 , \19353 , \19354 , \19355 , \19356 , \19357 , \19358 ,
         \19359 , \19360 , \19361 , \19362 , \19363 , \19364 , \19365 , \19366 , \19367 , \19368 ,
         \19369 , \19370 , \19371 , \19372 , \19373 , \19374 , \19375_nG54d5 , \19376 , \19377 , \19378 ,
         \19379 , \19380 , \19381 , \19382 , \19383 , \19384 , \19385 , \19386 , \19387 , \19388 ,
         \19389 , \19390 , \19391 , \19392 , \19393 , \19394 , \19395 , \19396 , \19397 , \19398 ,
         \19399 , \19400 , \19401 , \19402 , \19403 , \19404 , \19405 , \19406 , \19407 , \19408 ,
         \19409 , \19410 , \19411 , \19412 , \19413 , \19414 , \19415 , \19416 , \19417 , \19418 ,
         \19419 , \19420 , \19421 , \19422 , \19423 , \19424 , \19425 , \19426 , \19427 , \19428 ,
         \19429 , \19430 , \19431 , \19432 , \19433 , \19434 , \19435 , \19436 , \19437 , \19438 ,
         \19439 , \19440 , \19441 , \19442 , \19443 , \19444 , \19445 , \19446 , \19447 , \19448 ,
         \19449 , \19450 , \19451 , \19452 , \19453 , \19454 , \19455 , \19456 , \19457 , \19458 ,
         \19459 , \19460 , \19461 , \19462 , \19463 , \19464 , \19465 , \19466 , \19467 , \19468 ,
         \19469 , \19470 , \19471 , \19472 , \19473 , \19474 , \19475 , \19476 , \19477 , \19478 ,
         \19479 , \19480 , \19481 , \19482 , \19483 , \19484 , \19485 , \19486 , \19487 , \19488 ,
         \19489 , \19490 , \19491 , \19492 , \19493 , \19494 , \19495 , \19496 , \19497 , \19498 ,
         \19499 , \19500 , \19501 , \19502 , \19503 , \19504 , \19505 , \19506 , \19507 , \19508 ,
         \19509 , \19510 , \19511 , \19512 , \19513 , \19514 , \19515 , \19516 , \19517 , \19518 ,
         \19519 , \19520 , \19521 , \19522 , \19523 , \19524 , \19525 , \19526 , \19527 , \19528 ,
         \19529 , \19530_nG54d3 , \19531 , \19532 , \19533 , \19534 , \19535 , \19536 , \19537 , \19538 ,
         \19539 , \19540 , \19541 , \19542 , \19543 , \19544 , \19545 , \19546 , \19547 , \19548 ,
         \19549 , \19550 , \19551 , \19552 , \19553 , \19554 , \19555 , \19556 , \19557 , \19558 ,
         \19559 , \19560 , \19561 , \19562 , \19563 , \19564 , \19565 , \19566 , \19567 , \19568 ,
         \19569 , \19570 , \19571 , \19572 , \19573 , \19574 , \19575 , \19576 , \19577 , \19578 ,
         \19579 , \19580 , \19581 , \19582 , \19583 , \19584 , \19585 , \19586 , \19587 , \19588 ,
         \19589 , \19590 , \19591 , \19592 , \19593 , \19594 , \19595 , \19596 , \19597 , \19598 ,
         \19599 , \19600 , \19601 , \19602 , \19603 , \19604 , \19605 , \19606 , \19607 , \19608 ,
         \19609 , \19610 , \19611 , \19612 , \19613 , \19614 , \19615 , \19616 , \19617 , \19618 ,
         \19619 , \19620 , \19621 , \19622 , \19623 , \19624 , \19625 , \19626 , \19627 , \19628 ,
         \19629 , \19630 , \19631 , \19632 , \19633 , \19634 , \19635 , \19636 , \19637 , \19638 ,
         \19639 , \19640 , \19641 , \19642 , \19643 , \19644 , \19645 , \19646 , \19647 , \19648 ,
         \19649 , \19650 , \19651 , \19652 , \19653 , \19654 , \19655 , \19656 , \19657 , \19658 ,
         \19659 , \19660 , \19661 , \19662 , \19663 , \19664 , \19665 , \19666 , \19667 , \19668 ,
         \19669 , \19670 , \19671 , \19672 , \19673 , \19674 , \19675 , \19676 , \19677 , \19678_nG54d1 ,
         \19679 , \19680 , \19681 , \19682 , \19683 , \19684 , \19685 , \19686 , \19687 , \19688 ,
         \19689 , \19690 , \19691 , \19692 , \19693 , \19694 , \19695 , \19696 , \19697 , \19698 ,
         \19699 , \19700 , \19701 , \19702 , \19703 , \19704 , \19705 , \19706 , \19707 , \19708 ,
         \19709 , \19710 , \19711 , \19712 , \19713 , \19714 , \19715 , \19716 , \19717 , \19718 ,
         \19719 , \19720 , \19721 , \19722 , \19723 , \19724 , \19725 , \19726 , \19727 , \19728 ,
         \19729 , \19730 , \19731 , \19732 , \19733 , \19734 , \19735 , \19736 , \19737 , \19738 ,
         \19739 , \19740 , \19741 , \19742 , \19743 , \19744 , \19745 , \19746 , \19747 , \19748 ,
         \19749 , \19750 , \19751 , \19752 , \19753 , \19754 , \19755 , \19756 , \19757 , \19758 ,
         \19759 , \19760 , \19761 , \19762 , \19763 , \19764 , \19765 , \19766 , \19767 , \19768 ,
         \19769 , \19770 , \19771 , \19772 , \19773 , \19774 , \19775 , \19776 , \19777 , \19778 ,
         \19779 , \19780 , \19781 , \19782 , \19783 , \19784 , \19785 , \19786 , \19787 , \19788 ,
         \19789 , \19790 , \19791 , \19792 , \19793 , \19794 , \19795 , \19796 , \19797 , \19798 ,
         \19799 , \19800 , \19801 , \19802 , \19803 , \19804 , \19805 , \19806 , \19807 , \19808 ,
         \19809 , \19810 , \19811 , \19812 , \19813 , \19814 , \19815 , \19816 , \19817 , \19818 ,
         \19819 , \19820 , \19821_nG54cf , \19822 , \19823 , \19824 , \19825 , \19826 , \19827 , \19828 ,
         \19829 , \19830 , \19831 , \19832 , \19833 , \19834 , \19835 , \19836 , \19837 , \19838 ,
         \19839 , \19840 , \19841 , \19842 , \19843 , \19844 , \19845 , \19846 , \19847 , \19848 ,
         \19849 , \19850 , \19851 , \19852 , \19853 , \19854 , \19855 , \19856 , \19857 , \19858 ,
         \19859 , \19860 , \19861 , \19862 , \19863 , \19864 , \19865 , \19866 , \19867 , \19868 ,
         \19869 , \19870 , \19871 , \19872 , \19873 , \19874 , \19875 , \19876 , \19877 , \19878 ,
         \19879 , \19880 , \19881 , \19882 , \19883 , \19884 , \19885 , \19886 , \19887 , \19888 ,
         \19889 , \19890 , \19891 , \19892 , \19893 , \19894 , \19895 , \19896 , \19897 , \19898 ,
         \19899 , \19900 , \19901 , \19902 , \19903 , \19904 , \19905 , \19906 , \19907 , \19908 ,
         \19909 , \19910 , \19911 , \19912 , \19913 , \19914 , \19915 , \19916 , \19917 , \19918 ,
         \19919 , \19920 , \19921 , \19922 , \19923 , \19924 , \19925 , \19926 , \19927 , \19928 ,
         \19929 , \19930 , \19931 , \19932 , \19933 , \19934 , \19935 , \19936 , \19937 , \19938 ,
         \19939 , \19940 , \19941 , \19942 , \19943 , \19944 , \19945 , \19946 , \19947 , \19948 ,
         \19949 , \19950 , \19951 , \19952 , \19953 , \19954 , \19955 , \19956_nG54cd , \19957 , \19958 ,
         \19959 , \19960 , \19961 , \19962 , \19963 , \19964 , \19965 , \19966 , \19967 , \19968 ,
         \19969 , \19970 , \19971 , \19972 , \19973 , \19974 , \19975 , \19976 , \19977 , \19978 ,
         \19979 , \19980 , \19981 , \19982 , \19983 , \19984 , \19985 , \19986 , \19987 , \19988 ,
         \19989 , \19990 , \19991 , \19992 , \19993 , \19994 , \19995 , \19996 , \19997 , \19998 ,
         \19999 , \20000 , \20001 , \20002 , \20003 , \20004 , \20005 , \20006 , \20007 , \20008 ,
         \20009 , \20010 , \20011 , \20012 , \20013 , \20014 , \20015 , \20016 , \20017 , \20018 ,
         \20019 , \20020 , \20021 , \20022 , \20023 , \20024 , \20025 , \20026 , \20027 , \20028 ,
         \20029 , \20030 , \20031 , \20032 , \20033 , \20034 , \20035 , \20036 , \20037 , \20038 ,
         \20039 , \20040 , \20041 , \20042 , \20043 , \20044 , \20045 , \20046 , \20047 , \20048 ,
         \20049 , \20050 , \20051 , \20052 , \20053 , \20054 , \20055 , \20056 , \20057 , \20058 ,
         \20059 , \20060 , \20061 , \20062 , \20063 , \20064 , \20065 , \20066 , \20067 , \20068 ,
         \20069 , \20070 , \20071 , \20072 , \20073 , \20074 , \20075 , \20076 , \20077 , \20078 ,
         \20079 , \20080 , \20081 , \20082 , \20083 , \20084 , \20085 , \20086 , \20087 , \20088 ,
         \20089 , \20090_nG54cb , \20091 , \20092 , \20093 , \20094 , \20095 , \20096 , \20097 , \20098 ,
         \20099 , \20100 , \20101 , \20102 , \20103 , \20104 , \20105 , \20106 , \20107 , \20108 ,
         \20109 , \20110 , \20111 , \20112 , \20113 , \20114 , \20115 , \20116 , \20117 , \20118 ,
         \20119 , \20120 , \20121 , \20122 , \20123 , \20124 , \20125 , \20126 , \20127 , \20128 ,
         \20129 , \20130 , \20131 , \20132 , \20133 , \20134 , \20135 , \20136 , \20137 , \20138 ,
         \20139 , \20140 , \20141 , \20142 , \20143 , \20144 , \20145 , \20146 , \20147 , \20148 ,
         \20149 , \20150 , \20151 , \20152 , \20153 , \20154 , \20155 , \20156 , \20157 , \20158 ,
         \20159 , \20160 , \20161 , \20162 , \20163 , \20164 , \20165 , \20166 , \20167 , \20168 ,
         \20169 , \20170 , \20171 , \20172 , \20173 , \20174 , \20175 , \20176 , \20177 , \20178 ,
         \20179 , \20180 , \20181 , \20182 , \20183 , \20184 , \20185 , \20186 , \20187 , \20188 ,
         \20189 , \20190 , \20191 , \20192 , \20193 , \20194 , \20195 , \20196 , \20197 , \20198 ,
         \20199 , \20200 , \20201 , \20202 , \20203 , \20204 , \20205 , \20206 , \20207 , \20208 ,
         \20209 , \20210 , \20211 , \20212 , \20213 , \20214 , \20215 , \20216 , \20217 , \20218_nG54c9 ,
         \20219 , \20220 , \20221 , \20222 , \20223 , \20224 , \20225 , \20226 , \20227 , \20228 ,
         \20229 , \20230 , \20231 , \20232 , \20233 , \20234 , \20235 , \20236 , \20237 , \20238 ,
         \20239 , \20240 , \20241 , \20242 , \20243 , \20244 , \20245 , \20246 , \20247 , \20248 ,
         \20249 , \20250 , \20251 , \20252 , \20253 , \20254 , \20255 , \20256 , \20257 , \20258 ,
         \20259 , \20260 , \20261 , \20262 , \20263 , \20264 , \20265 , \20266 , \20267 , \20268 ,
         \20269 , \20270 , \20271 , \20272 , \20273 , \20274 , \20275 , \20276 , \20277 , \20278 ,
         \20279 , \20280 , \20281 , \20282 , \20283 , \20284 , \20285 , \20286 , \20287 , \20288 ,
         \20289 , \20290 , \20291 , \20292 , \20293 , \20294 , \20295 , \20296 , \20297 , \20298 ,
         \20299 , \20300 , \20301 , \20302 , \20303 , \20304 , \20305 , \20306 , \20307 , \20308 ,
         \20309 , \20310 , \20311 , \20312 , \20313 , \20314 , \20315 , \20316 , \20317 , \20318 ,
         \20319 , \20320 , \20321 , \20322 , \20323 , \20324 , \20325 , \20326 , \20327 , \20328 ,
         \20329 , \20330 , \20331 , \20332 , \20333 , \20334 , \20335 , \20336 , \20337 , \20338 ,
         \20339 , \20340 , \20341_nG54c7 , \20342 , \20343 , \20344 , \20345 , \20346 , \20347 , \20348 ,
         \20349 , \20350 , \20351 , \20352 , \20353 , \20354 , \20355 , \20356 , \20357 , \20358 ,
         \20359 , \20360 , \20361 , \20362 , \20363 , \20364 , \20365 , \20366 , \20367 , \20368 ,
         \20369 , \20370 , \20371 , \20372 , \20373 , \20374 , \20375 , \20376 , \20377 , \20378 ,
         \20379 , \20380 , \20381 , \20382 , \20383 , \20384 , \20385 , \20386 , \20387 , \20388 ,
         \20389 , \20390 , \20391 , \20392 , \20393 , \20394 , \20395 , \20396 , \20397 , \20398 ,
         \20399 , \20400 , \20401 , \20402 , \20403 , \20404 , \20405 , \20406 , \20407 , \20408 ,
         \20409 , \20410 , \20411 , \20412 , \20413 , \20414 , \20415 , \20416 , \20417 , \20418 ,
         \20419 , \20420 , \20421 , \20422 , \20423 , \20424 , \20425 , \20426 , \20427 , \20428 ,
         \20429 , \20430 , \20431 , \20432 , \20433 , \20434 , \20435 , \20436 , \20437 , \20438 ,
         \20439 , \20440 , \20441 , \20442 , \20443 , \20444 , \20445 , \20446 , \20447 , \20448 ,
         \20449 , \20450 , \20451 , \20452 , \20453 , \20454 , \20455 , \20456 , \20457_nG54c5 , \20458 ,
         \20459 , \20460 , \20461 , \20462 , \20463 , \20464 , \20465 , \20466 , \20467 , \20468 ,
         \20469 , \20470 , \20471 , \20472 , \20473 , \20474 , \20475 , \20476 , \20477 , \20478 ,
         \20479 , \20480 , \20481 , \20482 , \20483 , \20484 , \20485 , \20486 , \20487 , \20488 ,
         \20489 , \20490 , \20491 , \20492 , \20493 , \20494 , \20495 , \20496 , \20497 , \20498 ,
         \20499 , \20500 , \20501 , \20502 , \20503 , \20504 , \20505 , \20506 , \20507 , \20508 ,
         \20509 , \20510 , \20511 , \20512 , \20513 , \20514 , \20515 , \20516 , \20517 , \20518 ,
         \20519 , \20520 , \20521 , \20522 , \20523 , \20524 , \20525 , \20526 , \20527 , \20528 ,
         \20529 , \20530 , \20531 , \20532 , \20533 , \20534 , \20535 , \20536 , \20537 , \20538 ,
         \20539 , \20540 , \20541 , \20542 , \20543 , \20544 , \20545 , \20546 , \20547 , \20548 ,
         \20549 , \20550 , \20551 , \20552 , \20553 , \20554 , \20555 , \20556 , \20557 , \20558 ,
         \20559 , \20560 , \20561 , \20562 , \20563 , \20564 , \20565 , \20566 , \20567_nG54c3 , \20568 ,
         \20569 , \20570 , \20571 , \20572 , \20573 , \20574 , \20575 , \20576 , \20577 , \20578 ,
         \20579 , \20580 , \20581 , \20582 , \20583 , \20584 , \20585 , \20586 , \20587 , \20588 ,
         \20589 , \20590 , \20591 , \20592 , \20593 , \20594 , \20595 , \20596 , \20597 , \20598 ,
         \20599 , \20600 , \20601 , \20602 , \20603 , \20604 , \20605 , \20606 , \20607 , \20608 ,
         \20609 , \20610 , \20611 , \20612 , \20613 , \20614 , \20615 , \20616 , \20617 , \20618 ,
         \20619 , \20620 , \20621 , \20622 , \20623 , \20624 , \20625 , \20626 , \20627 , \20628 ,
         \20629 , \20630 , \20631 , \20632 , \20633 , \20634 , \20635 , \20636 , \20637 , \20638 ,
         \20639 , \20640 , \20641 , \20642 , \20643 , \20644 , \20645 , \20646 , \20647 , \20648 ,
         \20649 , \20650 , \20651 , \20652 , \20653 , \20654 , \20655 , \20656 , \20657 , \20658 ,
         \20659 , \20660 , \20661 , \20662 , \20663 , \20664 , \20665 , \20666 , \20667 , \20668 ,
         \20669 , \20670 , \20671 , \20672_nG54c1 , \20673 , \20674 , \20675 , \20676 , \20677 , \20678 ,
         \20679 , \20680 , \20681 , \20682 , \20683 , \20684 , \20685 , \20686 , \20687 , \20688 ,
         \20689 , \20690 , \20691 , \20692 , \20693 , \20694 , \20695 , \20696 , \20697 , \20698 ,
         \20699 , \20700 , \20701 , \20702 , \20703 , \20704 , \20705 , \20706 , \20707 , \20708 ,
         \20709 , \20710 , \20711 , \20712 , \20713 , \20714 , \20715 , \20716 , \20717 , \20718 ,
         \20719 , \20720 , \20721 , \20722 , \20723 , \20724 , \20725 , \20726 , \20727 , \20728 ,
         \20729 , \20730 , \20731 , \20732 , \20733 , \20734 , \20735 , \20736 , \20737 , \20738 ,
         \20739 , \20740 , \20741 , \20742 , \20743 , \20744 , \20745 , \20746 , \20747 , \20748 ,
         \20749 , \20750 , \20751 , \20752 , \20753 , \20754 , \20755 , \20756 , \20757 , \20758 ,
         \20759 , \20760 , \20761 , \20762 , \20763 , \20764 , \20765 , \20766 , \20767 , \20768 ,
         \20769 , \20770 , \20771 , \20772 , \20773 , \20774 , \20775_nG54bf , \20776 , \20777 , \20778 ,
         \20779 , \20780 , \20781 , \20782 , \20783 , \20784 , \20785 , \20786 , \20787 , \20788 ,
         \20789 , \20790 , \20791 , \20792 , \20793 , \20794 , \20795 , \20796 , \20797 , \20798 ,
         \20799 , \20800 , \20801 , \20802 , \20803 , \20804 , \20805 , \20806 , \20807 , \20808 ,
         \20809 , \20810 , \20811 , \20812 , \20813 , \20814 , \20815 , \20816 , \20817 , \20818 ,
         \20819 , \20820 , \20821 , \20822 , \20823 , \20824 , \20825 , \20826 , \20827 , \20828 ,
         \20829 , \20830 , \20831 , \20832 , \20833 , \20834 , \20835 , \20836 , \20837 , \20838 ,
         \20839 , \20840 , \20841 , \20842 , \20843 , \20844 , \20845 , \20846 , \20847 , \20848 ,
         \20849 , \20850 , \20851 , \20852 , \20853 , \20854 , \20855 , \20856 , \20857 , \20858 ,
         \20859 , \20860 , \20861 , \20862 , \20863 , \20864 , \20865 , \20866 , \20867 , \20868 ,
         \20869 , \20870_nG54bd , \20871 , \20872 , \20873 , \20874 , \20875 , \20876 , \20877 , \20878 ,
         \20879 , \20880 , \20881 , \20882 , \20883 , \20884 , \20885 , \20886 , \20887 , \20888 ,
         \20889 , \20890 , \20891 , \20892 , \20893 , \20894 , \20895 , \20896 , \20897 , \20898 ,
         \20899 , \20900 , \20901 , \20902 , \20903 , \20904 , \20905 , \20906 , \20907 , \20908 ,
         \20909 , \20910 , \20911 , \20912 , \20913 , \20914 , \20915 , \20916 , \20917 , \20918 ,
         \20919 , \20920 , \20921 , \20922 , \20923 , \20924 , \20925 , \20926 , \20927 , \20928 ,
         \20929 , \20930 , \20931 , \20932 , \20933 , \20934 , \20935 , \20936 , \20937 , \20938 ,
         \20939 , \20940 , \20941 , \20942 , \20943 , \20944 , \20945 , \20946 , \20947 , \20948 ,
         \20949 , \20950 , \20951 , \20952 , \20953 , \20954 , \20955 , \20956 , \20957 , \20958 ,
         \20959 , \20960 , \20961 , \20962 , \20963_nG54bb , \20964 , \20965 , \20966 , \20967 , \20968 ,
         \20969 , \20970 , \20971 , \20972 , \20973 , \20974 , \20975 , \20976 , \20977 , \20978 ,
         \20979 , \20980 , \20981 , \20982 , \20983 , \20984 , \20985 , \20986 , \20987 , \20988 ,
         \20989 , \20990 , \20991 , \20992 , \20993 , \20994 , \20995 , \20996 , \20997 , \20998 ,
         \20999 , \21000 , \21001 , \21002 , \21003 , \21004 , \21005 , \21006 , \21007 , \21008 ,
         \21009 , \21010 , \21011 , \21012 , \21013 , \21014 , \21015 , \21016 , \21017 , \21018 ,
         \21019 , \21020 , \21021 , \21022 , \21023 , \21024 , \21025 , \21026 , \21027 , \21028 ,
         \21029 , \21030 , \21031 , \21032 , \21033 , \21034 , \21035 , \21036 , \21037 , \21038 ,
         \21039 , \21040 , \21041 , \21042 , \21043 , \21044 , \21045 , \21046 , \21047 , \21048_nG54b9 ,
         \21049 , \21050 , \21051 , \21052 , \21053 , \21054 , \21055 , \21056 , \21057 , \21058 ,
         \21059 , \21060 , \21061 , \21062 , \21063 , \21064 , \21065 , \21066 , \21067 , \21068 ,
         \21069 , \21070 , \21071 , \21072 , \21073 , \21074 , \21075 , \21076 , \21077 , \21078 ,
         \21079 , \21080 , \21081 , \21082 , \21083 , \21084 , \21085 , \21086 , \21087 , \21088 ,
         \21089 , \21090 , \21091 , \21092 , \21093 , \21094 , \21095 , \21096 , \21097 , \21098 ,
         \21099 , \21100 , \21101 , \21102 , \21103 , \21104 , \21105 , \21106 , \21107 , \21108 ,
         \21109 , \21110 , \21111 , \21112 , \21113 , \21114 , \21115 , \21116 , \21117 , \21118 ,
         \21119 , \21120 , \21121 , \21122 , \21123 , \21124 , \21125 , \21126 , \21127 , \21128 ,
         \21129 , \21130 , \21131_nG54b7 , \21132 , \21133 , \21134 , \21135 , \21136 , \21137 , \21138 ,
         \21139 , \21140 , \21141 , \21142 , \21143 , \21144 , \21145 , \21146 , \21147 , \21148 ,
         \21149 , \21150 , \21151 , \21152 , \21153 , \21154 , \21155 , \21156 , \21157 , \21158 ,
         \21159 , \21160 , \21161 , \21162 , \21163 , \21164 , \21165 , \21166 , \21167 , \21168 ,
         \21169 , \21170 , \21171 , \21172 , \21173 , \21174 , \21175 , \21176 , \21177 , \21178 ,
         \21179 , \21180 , \21181 , \21182 , \21183 , \21184 , \21185 , \21186 , \21187 , \21188 ,
         \21189 , \21190 , \21191 , \21192 , \21193 , \21194 , \21195 , \21196 , \21197 , \21198 ,
         \21199 , \21200 , \21201 , \21202 , \21203 , \21204 , \21205 , \21206 , \21207_nG54b5 , \21208 ,
         \21209 , \21210 , \21211 , \21212 , \21213 , \21214 , \21215 , \21216 , \21217 , \21218 ,
         \21219 , \21220 , \21221 , \21222 , \21223 , \21224 , \21225 , \21226 , \21227 , \21228 ,
         \21229 , \21230 , \21231 , \21232 , \21233 , \21234 , \21235 , \21236 , \21237 , \21238 ,
         \21239 , \21240 , \21241 , \21242 , \21243 , \21244 , \21245 , \21246 , \21247 , \21248 ,
         \21249 , \21250 , \21251 , \21252 , \21253 , \21254 , \21255 , \21256 , \21257 , \21258 ,
         \21259 , \21260 , \21261 , \21262 , \21263 , \21264 , \21265 , \21266 , \21267 , \21268 ,
         \21269 , \21270 , \21271 , \21272 , \21273 , \21274 , \21275 , \21276 , \21277 , \21278_nG54b3 ,
         \21279 , \21280 , \21281 , \21282 , \21283 , \21284 , \21285 , \21286 , \21287 , \21288 ,
         \21289 , \21290 , \21291 , \21292 , \21293 , \21294 , \21295 , \21296 , \21297 , \21298 ,
         \21299 , \21300 , \21301 , \21302 , \21303 , \21304 , \21305 , \21306 , \21307 , \21308 ,
         \21309 , \21310 , \21311 , \21312 , \21313 , \21314 , \21315 , \21316 , \21317 , \21318 ,
         \21319 , \21320 , \21321 , \21322 , \21323 , \21324 , \21325 , \21326 , \21327 , \21328 ,
         \21329 , \21330 , \21331 , \21332 , \21333 , \21334 , \21335 , \21336 , \21337 , \21338 ,
         \21339 , \21340 , \21341 , \21342 , \21343 , \21344 , \21345 , \21346_nG54b1 , \21347 , \21348 ,
         \21349 , \21350 , \21351 , \21352 , \21353 , \21354 , \21355 , \21356 , \21357 , \21358 ,
         \21359 , \21360 , \21361 , \21362 , \21363 , \21364 , \21365 , \21366 , \21367 , \21368 ,
         \21369 , \21370 , \21371 , \21372 , \21373 , \21374 , \21375 , \21376 , \21377 , \21378 ,
         \21379 , \21380 , \21381 , \21382 , \21383 , \21384 , \21385 , \21386 , \21387 , \21388 ,
         \21389 , \21390 , \21391 , \21392 , \21393 , \21394 , \21395 , \21396 , \21397 , \21398 ,
         \21399 , \21400 , \21401 , \21402 , \21403 , \21404 , \21405 , \21406 , \21407 , \21408 ,
         \21409_nG54af , \21410 , \21411 , \21412 , \21413 , \21414 , \21415 , \21416 , \21417 , \21418 ,
         \21419 , \21420 , \21421 , \21422 , \21423 , \21424 , \21425 , \21426 , \21427 , \21428 ,
         \21429 , \21430 , \21431 , \21432 , \21433 , \21434 , \21435 , \21436 , \21437 , \21438 ,
         \21439 , \21440 , \21441 , \21442 , \21443 , \21444 , \21445 , \21446 , \21447 , \21448 ,
         \21449 , \21450 , \21451 , \21452 , \21453 , \21454 , \21455 , \21456 , \21457 , \21458 ,
         \21459 , \21460 , \21461 , \21462 , \21463 , \21464_nG54ad , \21465 , \21466 , \21467 , \21468 ,
         \21469 , \21470 , \21471 , \21472 , \21473 , \21474 , \21475 , \21476 , \21477 , \21478 ,
         \21479 , \21480 , \21481 , \21482 , \21483 , \21484 , \21485 , \21486 , \21487 , \21488 ,
         \21489 , \21490 , \21491 , \21492 , \21493 , \21494 , \21495 , \21496 , \21497 , \21498 ,
         \21499 , \21500 , \21501 , \21502 , \21503 , \21504 , \21505 , \21506 , \21507 , \21508 ,
         \21509 , \21510 , \21511 , \21512 , \21513 , \21514 , \21515 , \21516 , \21517_nG54ab , \21518 ,
         \21519 , \21520 , \21521 , \21522 , \21523 , \21524 , \21525 , \21526 , \21527 , \21528 ,
         \21529 , \21530 , \21531 , \21532 , \21533 , \21534 , \21535 , \21536 , \21537 , \21538 ,
         \21539 , \21540 , \21541 , \21542 , \21543 , \21544 , \21545 , \21546 , \21547 , \21548 ,
         \21549 , \21550 , \21551 , \21552 , \21553 , \21554 , \21555 , \21556 , \21557 , \21558 ,
         \21559 , \21560 , \21561 , \21562 , \21563_nG54a9 , \21564 , \21565 , \21566 , \21567 , \21568 ,
         \21569 , \21570 , \21571 , \21572 , \21573 , \21574 , \21575 , \21576 , \21577 , \21578 ,
         \21579 , \21580 , \21581 , \21582 , \21583 , \21584 , \21585 , \21586 , \21587 , \21588 ,
         \21589 , \21590 , \21591 , \21592 , \21593 , \21594 , \21595 , \21596 , \21597 , \21598 ,
         \21599 , \21600 , \21601 , \21602 , \21603 , \21604_nG54a7 , \21605 , \21606 , \21607 , \21608 ,
         \21609 , \21610 , \21611 , \21612 , \21613 , \21614 , \21615 , \21616 , \21617 , \21618 ,
         \21619 , \21620 , \21621 , \21622 , \21623 , \21624 , \21625 , \21626 , \21627 , \21628 ,
         \21629 , \21630 , \21631 , \21632 , \21633 , \21634 , \21635 , \21636 , \21637 , \21638 ,
         \21639 , \21640 , \21641 , \21642_nG54a5 , \21643 , \21644 , \21645 , \21646 , \21647 , \21648 ,
         \21649 , \21650 , \21651 , \21652 , \21653 , \21654 , \21655 , \21656 , \21657 , \21658 ,
         \21659 , \21660 , \21661 , \21662 , \21663 , \21664 , \21665 , \21666 , \21667 , \21668 ,
         \21669 , \21670 , \21671 , \21672 , \21673 , \21674 , \21675_nG54a3 , \21676 , \21677 , \21678 ,
         \21679 , \21680 , \21681 , \21682 , \21683 , \21684 , \21685 , \21686 , \21687 , \21688 ,
         \21689 , \21690 , \21691 , \21692 , \21693 , \21694 , \21695 , \21696 , \21697 , \21698 ,
         \21699 , \21700 , \21701_nG54a1 , \21702 , \21703 , \21704 , \21705 , \21706 , \21707 , \21708 ,
         \21709 , \21710 , \21711 , \21712 , \21713 , \21714 , \21715 , \21716 , \21717 , \21718 ,
         \21719 , \21720 , \21721 , \21722_nG549f , \21723 , \21724 , \21725 , \21726 , \21727 , \21728 ,
         \21729 , \21730 , \21731 , \21732 , \21733 , \21734 , \21735_nG549d , \21736 , \21737 , \21738_nG557b ,
         \21739 , \21740 , \21741_nG5579 , \21742 , \21743 , \21744_nG5583 , \21745 , \21746 , \21747_nG5581 , \21748 ,
         \21749 , \21750_nG557f , \21751 , \21752 , \21753_nG557d , \21754 , \21755 , \21756_nG5587 , \21757 , \21758 ,
         \21759_nG5585 , \21760 , \21761 , \21762_nG5589 , \21763 , \21764 , \21765_nG558b , \21766 , \21767 , \21768_nG558f ,
         \21769 , \21770 , \21771_nG558d , \21772 , \21773 , \21774_nG5599 , \21775 , \21776 , \21777_nG5597 , \21778 ,
         \21779 , \21780_nG5595 , \21781 , \21782 , \21783_nG5593 , \21784 , \21785 , \21786_nG5591 , \21787 , \21788 ,
         \21789_nG559b , \21790 , \21791 , \21792 , \21793 , \21794 , \21795 , \21796 , \21797 , \21798 ,
         \21799 , \21800 , \21801 , \21802 , \21803 , \21804 , \21805 , \21806 , \21807 , \21808 ,
         \21809 , \21810 , \21811 , \21812 , \21813 , \21814 , \21815 , \21816 , \21817 , \21818 ,
         \21819 , \21820 , \21821 , \21822 , \21823 , \21824 , \21825 , \21826 , \21827 , \21828 ,
         \21829 , \21830 , \21831 , \21832 , \21833 , \21834 , \21835 , \21836 , \21837 , \21838 ,
         \21839 , \21840 , \21841 , \21842 , \21843 , \21844 , \21845 , \21846 , \21847 , \21848 ,
         \21849 , \21850 , \21851 , \21852 , \21853 , \21854 , \21855 , \21856 , \21857 , \21858 ,
         \21859 , \21860 , \21861 , \21862 , \21863 , \21864 , \21865 , \21866 , \21867 , \21868 ,
         \21869 , \21870 , \21871 , \21872 , \21873 , \21874 , \21875 , \21876 , \21877 , \21878 ,
         \21879 , \21880 , \21881 , \21882 , \21883 , \21884 , \21885 , \21886 , \21887 , \21888 ,
         \21889 , \21890 , \21891 , \21892 , \21893 , \21894 , \21895 , \21896 , \21897 , \21898 ,
         \21899 , \21900 , \21901 , \21902 , \21903 , \21904 , \21905 , \21906 , \21907 , \21908 ,
         \21909 , \21910 , \21911 , \21912 , \21913 , \21914 , \21915 , \21916 , \21917 , \21918 ,
         \21919 , \21920 , \21921 , \21922 , \21923 , \21924 , \21925 , \21926 , \21927 , \21928 ,
         \21929 , \21930 , \21931 , \21932 , \21933 , \21934 , \21935 , \21936 , \21937 , \21938 ,
         \21939 , \21940 , \21941 , \21942 , \21943 , \21944_nG56b6 , \21945 ;
buf \U$labaj2214 ( R_81_7e072f0, \21945 );
buf \U$2 ( \134 , RIb559478_125);
buf \U$3 ( \135 , RIb55f760_53);
buf \U$4 ( \136 , RIb55f6e8_54);
xor \U$5 ( \137 , \135 , \136 );
buf \U$6 ( \138 , RIb55f670_55);
xor \U$7 ( \139 , \136 , \138 );
not \U$8 ( \140 , \139 );
and \U$9 ( \141 , \137 , \140 );
and \U$10 ( \142 , \134 , \141 );
buf \U$11 ( \143 , RIb5594f0_124);
and \U$12 ( \144 , \143 , \139 );
nor \U$13 ( \145 , \142 , \144 );
and \U$14 ( \146 , \136 , \138 );
not \U$15 ( \147 , \146 );
and \U$16 ( \148 , \135 , \147 );
xnor \U$17 ( \149 , \145 , \148 );
buf \U$18 ( \150 , RIb559388_127);
buf \U$19 ( \151 , RIb55f850_51);
buf \U$20 ( \152 , RIb55f7d8_52);
xor \U$21 ( \153 , \151 , \152 );
xor \U$22 ( \154 , \152 , \135 );
not \U$23 ( \155 , \154 );
and \U$24 ( \156 , \153 , \155 );
and \U$25 ( \157 , \150 , \156 );
buf \U$26 ( \158 , RIb559400_126);
and \U$27 ( \159 , \158 , \154 );
nor \U$28 ( \160 , \157 , \159 );
and \U$29 ( \161 , \152 , \135 );
not \U$30 ( \162 , \161 );
and \U$31 ( \163 , \151 , \162 );
xnor \U$32 ( \164 , \160 , \163 );
and \U$33 ( \165 , \149 , \164 );
buf \U$34 ( \166 , RIb559310_128);
buf \U$35 ( \167 , RIb55f8c8_50);
xor \U$36 ( \168 , \167 , \151 );
nand \U$37 ( \169 , \166 , \168 );
buf \U$38 ( \170 , RIb55f940_49);
and \U$39 ( \171 , \167 , \151 );
not \U$40 ( \172 , \171 );
and \U$41 ( \173 , \170 , \172 );
xnor \U$42 ( \174 , \169 , \173 );
and \U$43 ( \175 , \164 , \174 );
and \U$44 ( \176 , \149 , \174 );
or \U$45 ( \177 , \165 , \175 , \176 );
buf \U$46 ( \178 , RIb55da50_115);
buf \U$47 ( \179 , RIb55f2b0_63);
buf \U$48 ( \180 , RIb55f238_64);
xor \U$49 ( \181 , \179 , \180 );
not \U$50 ( \182 , \180 );
and \U$51 ( \183 , \181 , \182 );
and \U$52 ( \184 , \178 , \183 );
buf \U$53 ( \185 , RIb55dac8_114);
and \U$54 ( \186 , \185 , \180 );
nor \U$55 ( \187 , \184 , \186 );
xnor \U$56 ( \188 , \187 , \179 );
buf \U$57 ( \189 , RIb55d960_117);
buf \U$58 ( \190 , RIb55f3a0_61);
buf \U$59 ( \191 , RIb55f328_62);
xor \U$60 ( \192 , \190 , \191 );
xor \U$61 ( \193 , \191 , \179 );
not \U$62 ( \194 , \193 );
and \U$63 ( \195 , \192 , \194 );
and \U$64 ( \196 , \189 , \195 );
buf \U$65 ( \197 , RIb55d9d8_116);
and \U$66 ( \198 , \197 , \193 );
nor \U$67 ( \199 , \196 , \198 );
and \U$68 ( \200 , \191 , \179 );
not \U$69 ( \201 , \200 );
and \U$70 ( \202 , \190 , \201 );
xnor \U$71 ( \203 , \199 , \202 );
and \U$72 ( \204 , \188 , \203 );
and \U$73 ( \205 , \203 , \173 );
and \U$74 ( \206 , \188 , \173 );
or \U$75 ( \207 , \204 , \205 , \206 );
and \U$76 ( \208 , \177 , \207 );
buf \U$77 ( \209 , RIb55d870_119);
buf \U$78 ( \210 , RIb55f490_59);
buf \U$79 ( \211 , RIb55f418_60);
xor \U$80 ( \212 , \210 , \211 );
xor \U$81 ( \213 , \211 , \190 );
not \U$82 ( \214 , \213 );
and \U$83 ( \215 , \212 , \214 );
and \U$84 ( \216 , \209 , \215 );
buf \U$85 ( \217 , RIb55d8e8_118);
and \U$86 ( \218 , \217 , \213 );
nor \U$87 ( \219 , \216 , \218 );
and \U$88 ( \220 , \211 , \190 );
not \U$89 ( \221 , \220 );
and \U$90 ( \222 , \210 , \221 );
xnor \U$91 ( \223 , \219 , \222 );
buf \U$92 ( \224 , RIb55d780_121);
buf \U$93 ( \225 , RIb55f580_57);
buf \U$94 ( \226 , RIb55f508_58);
xor \U$95 ( \227 , \225 , \226 );
xor \U$96 ( \228 , \226 , \210 );
not \U$97 ( \229 , \228 );
and \U$98 ( \230 , \227 , \229 );
and \U$99 ( \231 , \224 , \230 );
buf \U$100 ( \232 , RIb55d7f8_120);
and \U$101 ( \233 , \232 , \228 );
nor \U$102 ( \234 , \231 , \233 );
and \U$103 ( \235 , \226 , \210 );
not \U$104 ( \236 , \235 );
and \U$105 ( \237 , \225 , \236 );
xnor \U$106 ( \238 , \234 , \237 );
and \U$107 ( \239 , \223 , \238 );
buf \U$108 ( \240 , RIb55d690_123);
buf \U$109 ( \241 , RIb55f5f8_56);
xor \U$110 ( \242 , \138 , \241 );
xor \U$111 ( \243 , \241 , \225 );
not \U$112 ( \244 , \243 );
and \U$113 ( \245 , \242 , \244 );
and \U$114 ( \246 , \240 , \245 );
buf \U$115 ( \247 , RIb55d708_122);
and \U$116 ( \248 , \247 , \243 );
nor \U$117 ( \249 , \246 , \248 );
and \U$118 ( \250 , \241 , \225 );
not \U$119 ( \251 , \250 );
and \U$120 ( \252 , \138 , \251 );
xnor \U$121 ( \253 , \249 , \252 );
and \U$122 ( \254 , \238 , \253 );
and \U$123 ( \255 , \223 , \253 );
or \U$124 ( \256 , \239 , \254 , \255 );
and \U$125 ( \257 , \207 , \256 );
and \U$126 ( \258 , \177 , \256 );
or \U$127 ( \259 , \208 , \257 , \258 );
and \U$128 ( \260 , \185 , \183 );
buf \U$129 ( \261 , RIb55db40_113);
and \U$130 ( \262 , \261 , \180 );
nor \U$131 ( \263 , \260 , \262 );
xnor \U$132 ( \264 , \263 , \179 );
and \U$133 ( \265 , \197 , \195 );
and \U$134 ( \266 , \178 , \193 );
nor \U$135 ( \267 , \265 , \266 );
xnor \U$136 ( \268 , \267 , \202 );
xor \U$137 ( \269 , \264 , \268 );
and \U$138 ( \270 , \217 , \215 );
and \U$139 ( \271 , \189 , \213 );
nor \U$140 ( \272 , \270 , \271 );
xnor \U$141 ( \273 , \272 , \222 );
xor \U$142 ( \274 , \269 , \273 );
and \U$143 ( \275 , \232 , \230 );
and \U$144 ( \276 , \209 , \228 );
nor \U$145 ( \277 , \275 , \276 );
xnor \U$146 ( \278 , \277 , \237 );
and \U$147 ( \279 , \247 , \245 );
and \U$148 ( \280 , \224 , \243 );
nor \U$149 ( \281 , \279 , \280 );
xnor \U$150 ( \282 , \281 , \252 );
xor \U$151 ( \283 , \278 , \282 );
and \U$152 ( \284 , \143 , \141 );
and \U$153 ( \285 , \240 , \139 );
nor \U$154 ( \286 , \284 , \285 );
xnor \U$155 ( \287 , \286 , \148 );
xor \U$156 ( \288 , \283 , \287 );
and \U$157 ( \289 , \274 , \288 );
and \U$158 ( \290 , \158 , \156 );
and \U$159 ( \291 , \134 , \154 );
nor \U$160 ( \292 , \290 , \291 );
xnor \U$161 ( \293 , \292 , \163 );
xor \U$162 ( \294 , \170 , \167 );
not \U$163 ( \295 , \168 );
and \U$164 ( \296 , \294 , \295 );
and \U$165 ( \297 , \166 , \296 );
and \U$166 ( \298 , \150 , \168 );
nor \U$167 ( \299 , \297 , \298 );
xnor \U$168 ( \300 , \299 , \173 );
xor \U$169 ( \301 , \293 , \300 );
and \U$170 ( \302 , \288 , \301 );
and \U$171 ( \303 , \274 , \301 );
or \U$172 ( \304 , \289 , \302 , \303 );
and \U$173 ( \305 , \259 , \304 );
and \U$174 ( \306 , \261 , \183 );
buf \U$175 ( \307 , RIb55dbb8_112);
and \U$176 ( \308 , \307 , \180 );
nor \U$177 ( \309 , \306 , \308 );
xnor \U$178 ( \310 , \309 , \179 );
and \U$179 ( \311 , \178 , \195 );
and \U$180 ( \312 , \185 , \193 );
nor \U$181 ( \313 , \311 , \312 );
xnor \U$182 ( \314 , \313 , \202 );
xor \U$183 ( \315 , \310 , \314 );
buf \U$184 ( \316 , RIb55fa30_47);
buf \U$185 ( \317 , RIb55f9b8_48);
and \U$186 ( \318 , \317 , \170 );
not \U$187 ( \319 , \318 );
and \U$188 ( \320 , \316 , \319 );
xor \U$189 ( \321 , \315 , \320 );
and \U$190 ( \322 , \304 , \321 );
and \U$191 ( \323 , \259 , \321 );
or \U$192 ( \324 , \305 , \322 , \323 );
and \U$193 ( \325 , \264 , \268 );
and \U$194 ( \326 , \268 , \273 );
and \U$195 ( \327 , \264 , \273 );
or \U$196 ( \328 , \325 , \326 , \327 );
and \U$197 ( \329 , \278 , \282 );
and \U$198 ( \330 , \282 , \287 );
and \U$199 ( \331 , \278 , \287 );
or \U$200 ( \332 , \329 , \330 , \331 );
xor \U$201 ( \333 , \328 , \332 );
and \U$202 ( \334 , \293 , \300 );
xor \U$203 ( \335 , \333 , \334 );
xor \U$204 ( \336 , \317 , \170 );
nand \U$205 ( \337 , \166 , \336 );
xnor \U$206 ( \338 , \337 , \320 );
and \U$207 ( \339 , \189 , \215 );
and \U$208 ( \340 , \197 , \213 );
nor \U$209 ( \341 , \339 , \340 );
xnor \U$210 ( \342 , \341 , \222 );
and \U$211 ( \343 , \209 , \230 );
and \U$212 ( \344 , \217 , \228 );
nor \U$213 ( \345 , \343 , \344 );
xnor \U$214 ( \346 , \345 , \237 );
xor \U$215 ( \347 , \342 , \346 );
and \U$216 ( \348 , \224 , \245 );
and \U$217 ( \349 , \232 , \243 );
nor \U$218 ( \350 , \348 , \349 );
xnor \U$219 ( \351 , \350 , \252 );
xor \U$220 ( \352 , \347 , \351 );
xor \U$221 ( \353 , \338 , \352 );
and \U$222 ( \354 , \240 , \141 );
and \U$223 ( \355 , \247 , \139 );
nor \U$224 ( \356 , \354 , \355 );
xnor \U$225 ( \357 , \356 , \148 );
and \U$226 ( \358 , \134 , \156 );
and \U$227 ( \359 , \143 , \154 );
nor \U$228 ( \360 , \358 , \359 );
xnor \U$229 ( \361 , \360 , \163 );
xor \U$230 ( \362 , \357 , \361 );
and \U$231 ( \363 , \150 , \296 );
and \U$232 ( \364 , \158 , \168 );
nor \U$233 ( \365 , \363 , \364 );
xnor \U$234 ( \366 , \365 , \173 );
xor \U$235 ( \367 , \362 , \366 );
xor \U$236 ( \368 , \353 , \367 );
and \U$237 ( \369 , \335 , \368 );
and \U$238 ( \370 , \324 , \369 );
and \U$239 ( \371 , \342 , \346 );
and \U$240 ( \372 , \346 , \351 );
and \U$241 ( \373 , \342 , \351 );
or \U$242 ( \374 , \371 , \372 , \373 );
and \U$243 ( \375 , \310 , \314 );
and \U$244 ( \376 , \314 , \320 );
and \U$245 ( \377 , \310 , \320 );
or \U$246 ( \378 , \375 , \376 , \377 );
xor \U$247 ( \379 , \374 , \378 );
and \U$248 ( \380 , \357 , \361 );
and \U$249 ( \381 , \361 , \366 );
and \U$250 ( \382 , \357 , \366 );
or \U$251 ( \383 , \380 , \381 , \382 );
xor \U$252 ( \384 , \379 , \383 );
and \U$253 ( \385 , \369 , \384 );
and \U$254 ( \386 , \324 , \384 );
or \U$255 ( \387 , \370 , \385 , \386 );
and \U$256 ( \388 , \328 , \332 );
and \U$257 ( \389 , \332 , \334 );
and \U$258 ( \390 , \328 , \334 );
or \U$259 ( \391 , \388 , \389 , \390 );
and \U$260 ( \392 , \338 , \352 );
and \U$261 ( \393 , \352 , \367 );
and \U$262 ( \394 , \338 , \367 );
or \U$263 ( \395 , \392 , \393 , \394 );
and \U$264 ( \396 , \391 , \395 );
and \U$265 ( \397 , \217 , \230 );
and \U$266 ( \398 , \189 , \228 );
nor \U$267 ( \399 , \397 , \398 );
xnor \U$268 ( \400 , \399 , \237 );
and \U$269 ( \401 , \232 , \245 );
and \U$270 ( \402 , \209 , \243 );
nor \U$271 ( \403 , \401 , \402 );
xnor \U$272 ( \404 , \403 , \252 );
xor \U$273 ( \405 , \400 , \404 );
and \U$274 ( \406 , \247 , \141 );
and \U$275 ( \407 , \224 , \139 );
nor \U$276 ( \408 , \406 , \407 );
xnor \U$277 ( \409 , \408 , \148 );
xor \U$278 ( \410 , \405 , \409 );
and \U$279 ( \411 , \307 , \183 );
buf \U$280 ( \412 , RIb55dc30_111);
and \U$281 ( \413 , \412 , \180 );
nor \U$282 ( \414 , \411 , \413 );
xnor \U$283 ( \415 , \414 , \179 );
and \U$284 ( \416 , \185 , \195 );
and \U$285 ( \417 , \261 , \193 );
nor \U$286 ( \418 , \416 , \417 );
xnor \U$287 ( \419 , \418 , \202 );
xor \U$288 ( \420 , \415 , \419 );
and \U$289 ( \421 , \197 , \215 );
and \U$290 ( \422 , \178 , \213 );
nor \U$291 ( \423 , \421 , \422 );
xnor \U$292 ( \424 , \423 , \222 );
xor \U$293 ( \425 , \420 , \424 );
xor \U$294 ( \426 , \410 , \425 );
and \U$295 ( \427 , \143 , \156 );
and \U$296 ( \428 , \240 , \154 );
nor \U$297 ( \429 , \427 , \428 );
xnor \U$298 ( \430 , \429 , \163 );
and \U$299 ( \431 , \158 , \296 );
and \U$300 ( \432 , \134 , \168 );
nor \U$301 ( \433 , \431 , \432 );
xnor \U$302 ( \434 , \433 , \173 );
xor \U$303 ( \435 , \430 , \434 );
xor \U$304 ( \436 , \316 , \317 );
not \U$305 ( \437 , \336 );
and \U$306 ( \438 , \436 , \437 );
and \U$307 ( \439 , \166 , \438 );
and \U$308 ( \440 , \150 , \336 );
nor \U$309 ( \441 , \439 , \440 );
xnor \U$310 ( \442 , \441 , \320 );
xor \U$311 ( \443 , \435 , \442 );
xor \U$312 ( \444 , \426 , \443 );
and \U$313 ( \445 , \395 , \444 );
and \U$314 ( \446 , \391 , \444 );
or \U$315 ( \447 , \396 , \445 , \446 );
and \U$316 ( \448 , \374 , \378 );
and \U$317 ( \449 , \378 , \383 );
and \U$318 ( \450 , \374 , \383 );
or \U$319 ( \451 , \448 , \449 , \450 );
and \U$320 ( \452 , \410 , \425 );
and \U$321 ( \453 , \425 , \443 );
and \U$322 ( \454 , \410 , \443 );
or \U$323 ( \455 , \452 , \453 , \454 );
xor \U$324 ( \456 , \451 , \455 );
and \U$325 ( \457 , \178 , \215 );
and \U$326 ( \458 , \185 , \213 );
nor \U$327 ( \459 , \457 , \458 );
xnor \U$328 ( \460 , \459 , \222 );
and \U$329 ( \461 , \189 , \230 );
and \U$330 ( \462 , \197 , \228 );
nor \U$331 ( \463 , \461 , \462 );
xnor \U$332 ( \464 , \463 , \237 );
xor \U$333 ( \465 , \460 , \464 );
and \U$334 ( \466 , \209 , \245 );
and \U$335 ( \467 , \217 , \243 );
nor \U$336 ( \468 , \466 , \467 );
xnor \U$337 ( \469 , \468 , \252 );
xor \U$338 ( \470 , \465 , \469 );
xor \U$339 ( \471 , \456 , \470 );
xor \U$340 ( \472 , \447 , \471 );
and \U$341 ( \473 , \412 , \183 );
buf \U$342 ( \474 , RIb55dca8_110);
and \U$343 ( \475 , \474 , \180 );
nor \U$344 ( \476 , \473 , \475 );
xnor \U$345 ( \477 , \476 , \179 );
and \U$346 ( \478 , \261 , \195 );
and \U$347 ( \479 , \307 , \193 );
nor \U$348 ( \480 , \478 , \479 );
xnor \U$349 ( \481 , \480 , \202 );
xor \U$350 ( \482 , \477 , \481 );
buf \U$351 ( \483 , RIb55fb20_45);
buf \U$352 ( \484 , RIb55faa8_46);
and \U$353 ( \485 , \484 , \316 );
not \U$354 ( \486 , \485 );
and \U$355 ( \487 , \483 , \486 );
xor \U$356 ( \488 , \482 , \487 );
and \U$357 ( \489 , \400 , \404 );
and \U$358 ( \490 , \404 , \409 );
and \U$359 ( \491 , \400 , \409 );
or \U$360 ( \492 , \489 , \490 , \491 );
and \U$361 ( \493 , \415 , \419 );
and \U$362 ( \494 , \419 , \424 );
and \U$363 ( \495 , \415 , \424 );
or \U$364 ( \496 , \493 , \494 , \495 );
xor \U$365 ( \497 , \492 , \496 );
and \U$366 ( \498 , \430 , \434 );
and \U$367 ( \499 , \434 , \442 );
and \U$368 ( \500 , \430 , \442 );
or \U$369 ( \501 , \498 , \499 , \500 );
xor \U$370 ( \502 , \497 , \501 );
xor \U$371 ( \503 , \488 , \502 );
and \U$372 ( \504 , \150 , \438 );
and \U$373 ( \505 , \158 , \336 );
nor \U$374 ( \506 , \504 , \505 );
xnor \U$375 ( \507 , \506 , \320 );
xor \U$376 ( \508 , \484 , \316 );
nand \U$377 ( \509 , \166 , \508 );
xnor \U$378 ( \510 , \509 , \487 );
xor \U$379 ( \511 , \507 , \510 );
and \U$380 ( \512 , \224 , \141 );
and \U$381 ( \513 , \232 , \139 );
nor \U$382 ( \514 , \512 , \513 );
xnor \U$383 ( \515 , \514 , \148 );
and \U$384 ( \516 , \240 , \156 );
and \U$385 ( \517 , \247 , \154 );
nor \U$386 ( \518 , \516 , \517 );
xnor \U$387 ( \519 , \518 , \163 );
xor \U$388 ( \520 , \515 , \519 );
and \U$389 ( \521 , \134 , \296 );
and \U$390 ( \522 , \143 , \168 );
nor \U$391 ( \523 , \521 , \522 );
xnor \U$392 ( \524 , \523 , \173 );
xor \U$393 ( \525 , \520 , \524 );
xor \U$394 ( \526 , \511 , \525 );
xor \U$395 ( \527 , \503 , \526 );
xor \U$396 ( \528 , \472 , \527 );
xor \U$397 ( \529 , \387 , \528 );
xor \U$398 ( \530 , \324 , \369 );
xor \U$399 ( \531 , \530 , \384 );
xor \U$400 ( \532 , \391 , \395 );
xor \U$401 ( \533 , \532 , \444 );
and \U$402 ( \534 , \531 , \533 );
xor \U$403 ( \535 , \529 , \534 );
xor \U$404 ( \536 , \531 , \533 );
and \U$405 ( \537 , \197 , \183 );
and \U$406 ( \538 , \178 , \180 );
nor \U$407 ( \539 , \537 , \538 );
xnor \U$408 ( \540 , \539 , \179 );
and \U$409 ( \541 , \217 , \195 );
and \U$410 ( \542 , \189 , \193 );
nor \U$411 ( \543 , \541 , \542 );
xnor \U$412 ( \544 , \543 , \202 );
and \U$413 ( \545 , \540 , \544 );
and \U$414 ( \546 , \232 , \215 );
and \U$415 ( \547 , \209 , \213 );
nor \U$416 ( \548 , \546 , \547 );
xnor \U$417 ( \549 , \548 , \222 );
and \U$418 ( \550 , \544 , \549 );
and \U$419 ( \551 , \540 , \549 );
or \U$420 ( \552 , \545 , \550 , \551 );
and \U$421 ( \553 , \247 , \230 );
and \U$422 ( \554 , \224 , \228 );
nor \U$423 ( \555 , \553 , \554 );
xnor \U$424 ( \556 , \555 , \237 );
and \U$425 ( \557 , \143 , \245 );
and \U$426 ( \558 , \240 , \243 );
nor \U$427 ( \559 , \557 , \558 );
xnor \U$428 ( \560 , \559 , \252 );
and \U$429 ( \561 , \556 , \560 );
and \U$430 ( \562 , \158 , \141 );
and \U$431 ( \563 , \134 , \139 );
nor \U$432 ( \564 , \562 , \563 );
xnor \U$433 ( \565 , \564 , \148 );
and \U$434 ( \566 , \560 , \565 );
and \U$435 ( \567 , \556 , \565 );
or \U$436 ( \568 , \561 , \566 , \567 );
and \U$437 ( \569 , \552 , \568 );
xor \U$438 ( \570 , \149 , \164 );
xor \U$439 ( \571 , \570 , \174 );
and \U$440 ( \572 , \568 , \571 );
and \U$441 ( \573 , \552 , \571 );
or \U$442 ( \574 , \569 , \572 , \573 );
xor \U$443 ( \575 , \188 , \203 );
xor \U$444 ( \576 , \575 , \173 );
xor \U$445 ( \577 , \223 , \238 );
xor \U$446 ( \578 , \577 , \253 );
and \U$447 ( \579 , \576 , \578 );
and \U$448 ( \580 , \574 , \579 );
xor \U$449 ( \581 , \274 , \288 );
xor \U$450 ( \582 , \581 , \301 );
and \U$451 ( \583 , \579 , \582 );
and \U$452 ( \584 , \574 , \582 );
or \U$453 ( \585 , \580 , \583 , \584 );
xor \U$454 ( \586 , \259 , \304 );
xor \U$455 ( \587 , \586 , \321 );
and \U$456 ( \588 , \585 , \587 );
xor \U$457 ( \589 , \335 , \368 );
and \U$458 ( \590 , \587 , \589 );
and \U$459 ( \591 , \585 , \589 );
or \U$460 ( \592 , \588 , \590 , \591 );
and \U$461 ( \593 , \536 , \592 );
xor \U$462 ( \594 , \536 , \592 );
xor \U$463 ( \595 , \585 , \587 );
xor \U$464 ( \596 , \595 , \589 );
and \U$465 ( \597 , \189 , \183 );
and \U$466 ( \598 , \197 , \180 );
nor \U$467 ( \599 , \597 , \598 );
xnor \U$468 ( \600 , \599 , \179 );
and \U$469 ( \601 , \209 , \195 );
and \U$470 ( \602 , \217 , \193 );
nor \U$471 ( \603 , \601 , \602 );
xnor \U$472 ( \604 , \603 , \202 );
and \U$473 ( \605 , \600 , \604 );
and \U$474 ( \606 , \604 , \163 );
and \U$475 ( \607 , \600 , \163 );
or \U$476 ( \608 , \605 , \606 , \607 );
and \U$477 ( \609 , \224 , \215 );
and \U$478 ( \610 , \232 , \213 );
nor \U$479 ( \611 , \609 , \610 );
xnor \U$480 ( \612 , \611 , \222 );
and \U$481 ( \613 , \240 , \230 );
and \U$482 ( \614 , \247 , \228 );
nor \U$483 ( \615 , \613 , \614 );
xnor \U$484 ( \616 , \615 , \237 );
and \U$485 ( \617 , \612 , \616 );
and \U$486 ( \618 , \134 , \245 );
and \U$487 ( \619 , \143 , \243 );
nor \U$488 ( \620 , \618 , \619 );
xnor \U$489 ( \621 , \620 , \252 );
and \U$490 ( \622 , \616 , \621 );
and \U$491 ( \623 , \612 , \621 );
or \U$492 ( \624 , \617 , \622 , \623 );
and \U$493 ( \625 , \608 , \624 );
and \U$494 ( \626 , \166 , \156 );
and \U$495 ( \627 , \150 , \154 );
nor \U$496 ( \628 , \626 , \627 );
xnor \U$497 ( \629 , \628 , \163 );
and \U$498 ( \630 , \624 , \629 );
and \U$499 ( \631 , \608 , \629 );
or \U$500 ( \632 , \625 , \630 , \631 );
xor \U$501 ( \633 , \552 , \568 );
xor \U$502 ( \634 , \633 , \571 );
and \U$503 ( \635 , \632 , \634 );
xor \U$504 ( \636 , \576 , \578 );
and \U$505 ( \637 , \634 , \636 );
and \U$506 ( \638 , \632 , \636 );
or \U$507 ( \639 , \635 , \637 , \638 );
xor \U$508 ( \640 , \177 , \207 );
xor \U$509 ( \641 , \640 , \256 );
and \U$510 ( \642 , \639 , \641 );
xor \U$511 ( \643 , \574 , \579 );
xor \U$512 ( \644 , \643 , \582 );
and \U$513 ( \645 , \641 , \644 );
and \U$514 ( \646 , \639 , \644 );
or \U$515 ( \647 , \642 , \645 , \646 );
and \U$516 ( \648 , \596 , \647 );
xor \U$517 ( \649 , \596 , \647 );
xor \U$518 ( \650 , \639 , \641 );
xor \U$519 ( \651 , \650 , \644 );
and \U$520 ( \652 , \143 , \230 );
and \U$521 ( \653 , \240 , \228 );
nor \U$522 ( \654 , \652 , \653 );
xnor \U$523 ( \655 , \654 , \237 );
and \U$524 ( \656 , \158 , \245 );
and \U$525 ( \657 , \134 , \243 );
nor \U$526 ( \658 , \656 , \657 );
xnor \U$527 ( \659 , \658 , \252 );
and \U$528 ( \660 , \655 , \659 );
and \U$529 ( \661 , \166 , \141 );
and \U$530 ( \662 , \150 , \139 );
nor \U$531 ( \663 , \661 , \662 );
xnor \U$532 ( \664 , \663 , \148 );
and \U$533 ( \665 , \659 , \664 );
and \U$534 ( \666 , \655 , \664 );
or \U$535 ( \667 , \660 , \665 , \666 );
and \U$536 ( \668 , \217 , \183 );
and \U$537 ( \669 , \189 , \180 );
nor \U$538 ( \670 , \668 , \669 );
xnor \U$539 ( \671 , \670 , \179 );
and \U$540 ( \672 , \232 , \195 );
and \U$541 ( \673 , \209 , \193 );
nor \U$542 ( \674 , \672 , \673 );
xnor \U$543 ( \675 , \674 , \202 );
and \U$544 ( \676 , \671 , \675 );
and \U$545 ( \677 , \247 , \215 );
and \U$546 ( \678 , \224 , \213 );
nor \U$547 ( \679 , \677 , \678 );
xnor \U$548 ( \680 , \679 , \222 );
and \U$549 ( \681 , \675 , \680 );
and \U$550 ( \682 , \671 , \680 );
or \U$551 ( \683 , \676 , \681 , \682 );
and \U$552 ( \684 , \667 , \683 );
and \U$553 ( \685 , \150 , \141 );
and \U$554 ( \686 , \158 , \139 );
nor \U$555 ( \687 , \685 , \686 );
xnor \U$556 ( \688 , \687 , \148 );
and \U$557 ( \689 , \683 , \688 );
and \U$558 ( \690 , \667 , \688 );
or \U$559 ( \691 , \684 , \689 , \690 );
nand \U$560 ( \692 , \166 , \154 );
xnor \U$561 ( \693 , \692 , \163 );
xor \U$562 ( \694 , \600 , \604 );
xor \U$563 ( \695 , \694 , \163 );
and \U$564 ( \696 , \693 , \695 );
xor \U$565 ( \697 , \612 , \616 );
xor \U$566 ( \698 , \697 , \621 );
and \U$567 ( \699 , \695 , \698 );
and \U$568 ( \700 , \693 , \698 );
or \U$569 ( \701 , \696 , \699 , \700 );
and \U$570 ( \702 , \691 , \701 );
xor \U$571 ( \703 , \556 , \560 );
xor \U$572 ( \704 , \703 , \565 );
and \U$573 ( \705 , \701 , \704 );
and \U$574 ( \706 , \691 , \704 );
or \U$575 ( \707 , \702 , \705 , \706 );
xor \U$576 ( \708 , \540 , \544 );
xor \U$577 ( \709 , \708 , \549 );
xor \U$578 ( \710 , \608 , \624 );
xor \U$579 ( \711 , \710 , \629 );
and \U$580 ( \712 , \709 , \711 );
and \U$581 ( \713 , \707 , \712 );
xor \U$582 ( \714 , \632 , \634 );
xor \U$583 ( \715 , \714 , \636 );
and \U$584 ( \716 , \712 , \715 );
and \U$585 ( \717 , \707 , \715 );
or \U$586 ( \718 , \713 , \716 , \717 );
and \U$587 ( \719 , \651 , \718 );
xor \U$588 ( \720 , \651 , \718 );
xor \U$589 ( \721 , \707 , \712 );
xor \U$590 ( \722 , \721 , \715 );
and \U$591 ( \723 , \240 , \215 );
and \U$592 ( \724 , \247 , \213 );
nor \U$593 ( \725 , \723 , \724 );
xnor \U$594 ( \726 , \725 , \222 );
and \U$595 ( \727 , \134 , \230 );
and \U$596 ( \728 , \143 , \228 );
nor \U$597 ( \729 , \727 , \728 );
xnor \U$598 ( \730 , \729 , \237 );
and \U$599 ( \731 , \726 , \730 );
and \U$600 ( \732 , \150 , \245 );
and \U$601 ( \733 , \158 , \243 );
nor \U$602 ( \734 , \732 , \733 );
xnor \U$603 ( \735 , \734 , \252 );
and \U$604 ( \736 , \730 , \735 );
and \U$605 ( \737 , \726 , \735 );
or \U$606 ( \738 , \731 , \736 , \737 );
and \U$607 ( \739 , \209 , \183 );
and \U$608 ( \740 , \217 , \180 );
nor \U$609 ( \741 , \739 , \740 );
xnor \U$610 ( \742 , \741 , \179 );
and \U$611 ( \743 , \224 , \195 );
and \U$612 ( \744 , \232 , \193 );
nor \U$613 ( \745 , \743 , \744 );
xnor \U$614 ( \746 , \745 , \202 );
and \U$615 ( \747 , \742 , \746 );
and \U$616 ( \748 , \746 , \148 );
and \U$617 ( \749 , \742 , \148 );
or \U$618 ( \750 , \747 , \748 , \749 );
and \U$619 ( \751 , \738 , \750 );
xor \U$620 ( \752 , \655 , \659 );
xor \U$621 ( \753 , \752 , \664 );
and \U$622 ( \754 , \750 , \753 );
and \U$623 ( \755 , \738 , \753 );
or \U$624 ( \756 , \751 , \754 , \755 );
xor \U$625 ( \757 , \667 , \683 );
xor \U$626 ( \758 , \757 , \688 );
and \U$627 ( \759 , \756 , \758 );
xor \U$628 ( \760 , \693 , \695 );
xor \U$629 ( \761 , \760 , \698 );
and \U$630 ( \762 , \758 , \761 );
and \U$631 ( \763 , \756 , \761 );
or \U$632 ( \764 , \759 , \762 , \763 );
xor \U$633 ( \765 , \691 , \701 );
xor \U$634 ( \766 , \765 , \704 );
and \U$635 ( \767 , \764 , \766 );
xor \U$636 ( \768 , \709 , \711 );
and \U$637 ( \769 , \766 , \768 );
and \U$638 ( \770 , \764 , \768 );
or \U$639 ( \771 , \767 , \769 , \770 );
and \U$640 ( \772 , \722 , \771 );
xor \U$641 ( \773 , \722 , \771 );
xor \U$642 ( \774 , \764 , \766 );
xor \U$643 ( \775 , \774 , \768 );
and \U$644 ( \776 , \232 , \183 );
and \U$645 ( \777 , \209 , \180 );
nor \U$646 ( \778 , \776 , \777 );
xnor \U$647 ( \779 , \778 , \179 );
and \U$648 ( \780 , \247 , \195 );
and \U$649 ( \781 , \224 , \193 );
nor \U$650 ( \782 , \780 , \781 );
xnor \U$651 ( \783 , \782 , \202 );
and \U$652 ( \784 , \779 , \783 );
and \U$653 ( \785 , \143 , \215 );
and \U$654 ( \786 , \240 , \213 );
nor \U$655 ( \787 , \785 , \786 );
xnor \U$656 ( \788 , \787 , \222 );
and \U$657 ( \789 , \783 , \788 );
and \U$658 ( \790 , \779 , \788 );
or \U$659 ( \791 , \784 , \789 , \790 );
nand \U$660 ( \792 , \166 , \139 );
xnor \U$661 ( \793 , \792 , \148 );
and \U$662 ( \794 , \791 , \793 );
xor \U$663 ( \795 , \726 , \730 );
xor \U$664 ( \796 , \795 , \735 );
and \U$665 ( \797 , \793 , \796 );
and \U$666 ( \798 , \791 , \796 );
or \U$667 ( \799 , \794 , \797 , \798 );
xor \U$668 ( \800 , \671 , \675 );
xor \U$669 ( \801 , \800 , \680 );
and \U$670 ( \802 , \799 , \801 );
xor \U$671 ( \803 , \738 , \750 );
xor \U$672 ( \804 , \803 , \753 );
and \U$673 ( \805 , \801 , \804 );
and \U$674 ( \806 , \799 , \804 );
or \U$675 ( \807 , \802 , \805 , \806 );
xor \U$676 ( \808 , \756 , \758 );
xor \U$677 ( \809 , \808 , \761 );
and \U$678 ( \810 , \807 , \809 );
and \U$679 ( \811 , \775 , \810 );
xor \U$680 ( \812 , \775 , \810 );
xor \U$681 ( \813 , \807 , \809 );
and \U$682 ( \814 , \134 , \215 );
and \U$683 ( \815 , \143 , \213 );
nor \U$684 ( \816 , \814 , \815 );
xnor \U$685 ( \817 , \816 , \222 );
and \U$686 ( \818 , \150 , \230 );
and \U$687 ( \819 , \158 , \228 );
nor \U$688 ( \820 , \818 , \819 );
xnor \U$689 ( \821 , \820 , \237 );
and \U$690 ( \822 , \817 , \821 );
nand \U$691 ( \823 , \166 , \243 );
xnor \U$692 ( \824 , \823 , \252 );
and \U$693 ( \825 , \821 , \824 );
and \U$694 ( \826 , \817 , \824 );
or \U$695 ( \827 , \822 , \825 , \826 );
and \U$696 ( \828 , \224 , \183 );
and \U$697 ( \829 , \232 , \180 );
nor \U$698 ( \830 , \828 , \829 );
xnor \U$699 ( \831 , \830 , \179 );
and \U$700 ( \832 , \240 , \195 );
and \U$701 ( \833 , \247 , \193 );
nor \U$702 ( \834 , \832 , \833 );
xnor \U$703 ( \835 , \834 , \202 );
and \U$704 ( \836 , \831 , \835 );
and \U$705 ( \837 , \835 , \252 );
and \U$706 ( \838 , \831 , \252 );
or \U$707 ( \839 , \836 , \837 , \838 );
and \U$708 ( \840 , \827 , \839 );
and \U$709 ( \841 , \158 , \230 );
and \U$710 ( \842 , \134 , \228 );
nor \U$711 ( \843 , \841 , \842 );
xnor \U$712 ( \844 , \843 , \237 );
and \U$713 ( \845 , \839 , \844 );
and \U$714 ( \846 , \827 , \844 );
or \U$715 ( \847 , \840 , \845 , \846 );
and \U$716 ( \848 , \166 , \245 );
and \U$717 ( \849 , \150 , \243 );
nor \U$718 ( \850 , \848 , \849 );
xnor \U$719 ( \851 , \850 , \252 );
xor \U$720 ( \852 , \779 , \783 );
xor \U$721 ( \853 , \852 , \788 );
and \U$722 ( \854 , \851 , \853 );
and \U$723 ( \855 , \847 , \854 );
xor \U$724 ( \856 , \742 , \746 );
xor \U$725 ( \857 , \856 , \148 );
and \U$726 ( \858 , \854 , \857 );
and \U$727 ( \859 , \847 , \857 );
or \U$728 ( \860 , \855 , \858 , \859 );
xor \U$729 ( \861 , \799 , \801 );
xor \U$730 ( \862 , \861 , \804 );
and \U$731 ( \863 , \860 , \862 );
and \U$732 ( \864 , \813 , \863 );
xor \U$733 ( \865 , \813 , \863 );
xor \U$734 ( \866 , \860 , \862 );
xor \U$735 ( \867 , \791 , \793 );
xor \U$736 ( \868 , \867 , \796 );
xor \U$737 ( \869 , \847 , \854 );
xor \U$738 ( \870 , \869 , \857 );
and \U$739 ( \871 , \868 , \870 );
and \U$740 ( \872 , \866 , \871 );
xor \U$741 ( \873 , \866 , \871 );
xor \U$742 ( \874 , \868 , \870 );
and \U$743 ( \875 , \247 , \183 );
and \U$744 ( \876 , \224 , \180 );
nor \U$745 ( \877 , \875 , \876 );
xnor \U$746 ( \878 , \877 , \179 );
and \U$747 ( \879 , \143 , \195 );
and \U$748 ( \880 , \240 , \193 );
nor \U$749 ( \881 , \879 , \880 );
xnor \U$750 ( \882 , \881 , \202 );
and \U$751 ( \883 , \878 , \882 );
and \U$752 ( \884 , \158 , \215 );
and \U$753 ( \885 , \134 , \213 );
nor \U$754 ( \886 , \884 , \885 );
xnor \U$755 ( \887 , \886 , \222 );
and \U$756 ( \888 , \882 , \887 );
and \U$757 ( \889 , \878 , \887 );
or \U$758 ( \890 , \883 , \888 , \889 );
xor \U$759 ( \891 , \817 , \821 );
xor \U$760 ( \892 , \891 , \824 );
and \U$761 ( \893 , \890 , \892 );
xor \U$762 ( \894 , \831 , \835 );
xor \U$763 ( \895 , \894 , \252 );
and \U$764 ( \896 , \892 , \895 );
and \U$765 ( \897 , \890 , \895 );
or \U$766 ( \898 , \893 , \896 , \897 );
xor \U$767 ( \899 , \827 , \839 );
xor \U$768 ( \900 , \899 , \844 );
and \U$769 ( \901 , \898 , \900 );
xor \U$770 ( \902 , \851 , \853 );
and \U$771 ( \903 , \900 , \902 );
and \U$772 ( \904 , \898 , \902 );
or \U$773 ( \905 , \901 , \903 , \904 );
and \U$774 ( \906 , \874 , \905 );
xor \U$775 ( \907 , \874 , \905 );
xor \U$776 ( \908 , \898 , \900 );
xor \U$777 ( \909 , \908 , \902 );
and \U$778 ( \910 , \240 , \183 );
and \U$779 ( \911 , \247 , \180 );
nor \U$780 ( \912 , \910 , \911 );
xnor \U$781 ( \913 , \912 , \179 );
and \U$782 ( \914 , \134 , \195 );
and \U$783 ( \915 , \143 , \193 );
nor \U$784 ( \916 , \914 , \915 );
xnor \U$785 ( \917 , \916 , \202 );
and \U$786 ( \918 , \913 , \917 );
and \U$787 ( \919 , \917 , \237 );
and \U$788 ( \920 , \913 , \237 );
or \U$789 ( \921 , \918 , \919 , \920 );
and \U$790 ( \922 , \150 , \215 );
and \U$791 ( \923 , \158 , \213 );
nor \U$792 ( \924 , \922 , \923 );
xnor \U$793 ( \925 , \924 , \222 );
nand \U$794 ( \926 , \166 , \228 );
xnor \U$795 ( \927 , \926 , \237 );
and \U$796 ( \928 , \925 , \927 );
and \U$797 ( \929 , \921 , \928 );
and \U$798 ( \930 , \166 , \230 );
and \U$799 ( \931 , \150 , \228 );
nor \U$800 ( \932 , \930 , \931 );
xnor \U$801 ( \933 , \932 , \237 );
and \U$802 ( \934 , \928 , \933 );
and \U$803 ( \935 , \921 , \933 );
or \U$804 ( \936 , \929 , \934 , \935 );
xor \U$805 ( \937 , \890 , \892 );
xor \U$806 ( \938 , \937 , \895 );
and \U$807 ( \939 , \936 , \938 );
and \U$808 ( \940 , \909 , \939 );
xor \U$809 ( \941 , \909 , \939 );
xor \U$810 ( \942 , \936 , \938 );
xor \U$811 ( \943 , \878 , \882 );
xor \U$812 ( \944 , \943 , \887 );
xor \U$813 ( \945 , \921 , \928 );
xor \U$814 ( \946 , \945 , \933 );
and \U$815 ( \947 , \944 , \946 );
and \U$816 ( \948 , \942 , \947 );
xor \U$817 ( \949 , \942 , \947 );
xor \U$818 ( \950 , \944 , \946 );
and \U$819 ( \951 , \143 , \183 );
and \U$820 ( \952 , \240 , \180 );
nor \U$821 ( \953 , \951 , \952 );
xnor \U$822 ( \954 , \953 , \179 );
and \U$823 ( \955 , \158 , \195 );
and \U$824 ( \956 , \134 , \193 );
nor \U$825 ( \957 , \955 , \956 );
xnor \U$826 ( \958 , \957 , \202 );
and \U$827 ( \959 , \954 , \958 );
and \U$828 ( \960 , \166 , \215 );
and \U$829 ( \961 , \150 , \213 );
nor \U$830 ( \962 , \960 , \961 );
xnor \U$831 ( \963 , \962 , \222 );
and \U$832 ( \964 , \958 , \963 );
and \U$833 ( \965 , \954 , \963 );
or \U$834 ( \966 , \959 , \964 , \965 );
xor \U$835 ( \967 , \913 , \917 );
xor \U$836 ( \968 , \967 , \237 );
and \U$837 ( \969 , \966 , \968 );
xor \U$838 ( \970 , \925 , \927 );
and \U$839 ( \971 , \968 , \970 );
and \U$840 ( \972 , \966 , \970 );
or \U$841 ( \973 , \969 , \971 , \972 );
and \U$842 ( \974 , \950 , \973 );
xor \U$843 ( \975 , \950 , \973 );
xor \U$844 ( \976 , \966 , \968 );
xor \U$845 ( \977 , \976 , \970 );
and \U$846 ( \978 , \134 , \183 );
and \U$847 ( \979 , \143 , \180 );
nor \U$848 ( \980 , \978 , \979 );
xnor \U$849 ( \981 , \980 , \179 );
and \U$850 ( \982 , \150 , \195 );
and \U$851 ( \983 , \158 , \193 );
nor \U$852 ( \984 , \982 , \983 );
xnor \U$853 ( \985 , \984 , \202 );
and \U$854 ( \986 , \981 , \985 );
and \U$855 ( \987 , \985 , \222 );
and \U$856 ( \988 , \981 , \222 );
or \U$857 ( \989 , \986 , \987 , \988 );
xor \U$858 ( \990 , \954 , \958 );
xor \U$859 ( \991 , \990 , \963 );
and \U$860 ( \992 , \989 , \991 );
and \U$861 ( \993 , \977 , \992 );
xor \U$862 ( \994 , \977 , \992 );
xor \U$863 ( \995 , \989 , \991 );
nand \U$864 ( \996 , \166 , \213 );
xnor \U$865 ( \997 , \996 , \222 );
xor \U$866 ( \998 , \981 , \985 );
xor \U$867 ( \999 , \998 , \222 );
and \U$868 ( \1000 , \997 , \999 );
and \U$869 ( \1001 , \995 , \1000 );
xor \U$870 ( \1002 , \995 , \1000 );
xor \U$871 ( \1003 , \997 , \999 );
and \U$872 ( \1004 , \158 , \183 );
and \U$873 ( \1005 , \134 , \180 );
nor \U$874 ( \1006 , \1004 , \1005 );
xnor \U$875 ( \1007 , \1006 , \179 );
and \U$876 ( \1008 , \166 , \195 );
and \U$877 ( \1009 , \150 , \193 );
nor \U$878 ( \1010 , \1008 , \1009 );
xnor \U$879 ( \1011 , \1010 , \202 );
and \U$880 ( \1012 , \1007 , \1011 );
and \U$881 ( \1013 , \1003 , \1012 );
xor \U$882 ( \1014 , \1003 , \1012 );
xor \U$883 ( \1015 , \1007 , \1011 );
and \U$884 ( \1016 , \150 , \183 );
and \U$885 ( \1017 , \158 , \180 );
nor \U$886 ( \1018 , \1016 , \1017 );
xnor \U$887 ( \1019 , \1018 , \179 );
and \U$888 ( \1020 , \1019 , \202 );
and \U$889 ( \1021 , \1015 , \1020 );
xor \U$890 ( \1022 , \1015 , \1020 );
nand \U$891 ( \1023 , \166 , \193 );
xnor \U$892 ( \1024 , \1023 , \202 );
xor \U$893 ( \1025 , \1019 , \202 );
and \U$894 ( \1026 , \1024 , \1025 );
xor \U$895 ( \1027 , \1024 , \1025 );
and \U$896 ( \1028 , \166 , \183 );
and \U$897 ( \1029 , \150 , \180 );
nor \U$898 ( \1030 , \1028 , \1029 );
xnor \U$899 ( \1031 , \1030 , \179 );
nand \U$900 ( \1032 , \166 , \180 );
xnor \U$901 ( \1033 , \1032 , \179 );
and \U$902 ( \1034 , \1033 , \179 );
and \U$903 ( \1035 , \1031 , \1034 );
and \U$904 ( \1036 , \1027 , \1035 );
or \U$905 ( \1037 , \1026 , \1036 );
and \U$906 ( \1038 , \1022 , \1037 );
or \U$907 ( \1039 , \1021 , \1038 );
and \U$908 ( \1040 , \1014 , \1039 );
or \U$909 ( \1041 , \1013 , \1040 );
and \U$910 ( \1042 , \1002 , \1041 );
or \U$911 ( \1043 , \1001 , \1042 );
and \U$912 ( \1044 , \994 , \1043 );
or \U$913 ( \1045 , \993 , \1044 );
and \U$914 ( \1046 , \975 , \1045 );
or \U$915 ( \1047 , \974 , \1046 );
and \U$916 ( \1048 , \949 , \1047 );
or \U$917 ( \1049 , \948 , \1048 );
and \U$918 ( \1050 , \941 , \1049 );
or \U$919 ( \1051 , \940 , \1050 );
and \U$920 ( \1052 , \907 , \1051 );
or \U$921 ( \1053 , \906 , \1052 );
and \U$922 ( \1054 , \873 , \1053 );
or \U$923 ( \1055 , \872 , \1054 );
and \U$924 ( \1056 , \865 , \1055 );
or \U$925 ( \1057 , \864 , \1056 );
and \U$926 ( \1058 , \812 , \1057 );
or \U$927 ( \1059 , \811 , \1058 );
and \U$928 ( \1060 , \773 , \1059 );
or \U$929 ( \1061 , \772 , \1060 );
and \U$930 ( \1062 , \720 , \1061 );
or \U$931 ( \1063 , \719 , \1062 );
and \U$932 ( \1064 , \649 , \1063 );
or \U$933 ( \1065 , \648 , \1064 );
and \U$934 ( \1066 , \594 , \1065 );
or \U$935 ( \1067 , \593 , \1066 );
xor \U$936 ( \1068 , \535 , \1067 );
buf g5577_GF_PartitionCandidate( \1069_nG5577 , \1068 );
buf \U$937 ( \1070 , \1069_nG5577 );
and \U$938 ( \1071 , \447 , \471 );
and \U$939 ( \1072 , \471 , \527 );
and \U$940 ( \1073 , \447 , \527 );
or \U$941 ( \1074 , \1071 , \1072 , \1073 );
and \U$942 ( \1075 , \451 , \455 );
and \U$943 ( \1076 , \455 , \470 );
and \U$944 ( \1077 , \451 , \470 );
or \U$945 ( \1078 , \1075 , \1076 , \1077 );
and \U$946 ( \1079 , \488 , \502 );
and \U$947 ( \1080 , \502 , \526 );
and \U$948 ( \1081 , \488 , \526 );
or \U$949 ( \1082 , \1079 , \1080 , \1081 );
xor \U$950 ( \1083 , \1078 , \1082 );
xor \U$951 ( \1084 , \483 , \484 );
not \U$952 ( \1085 , \508 );
and \U$953 ( \1086 , \1084 , \1085 );
and \U$954 ( \1087 , \166 , \1086 );
and \U$955 ( \1088 , \150 , \508 );
nor \U$956 ( \1089 , \1087 , \1088 );
xnor \U$957 ( \1090 , \1089 , \487 );
and \U$958 ( \1091 , \247 , \156 );
and \U$959 ( \1092 , \224 , \154 );
nor \U$960 ( \1093 , \1091 , \1092 );
xnor \U$961 ( \1094 , \1093 , \163 );
and \U$962 ( \1095 , \143 , \296 );
and \U$963 ( \1096 , \240 , \168 );
nor \U$964 ( \1097 , \1095 , \1096 );
xnor \U$965 ( \1098 , \1097 , \173 );
xor \U$966 ( \1099 , \1094 , \1098 );
and \U$967 ( \1100 , \158 , \438 );
and \U$968 ( \1101 , \134 , \336 );
nor \U$969 ( \1102 , \1100 , \1101 );
xnor \U$970 ( \1103 , \1102 , \320 );
xor \U$971 ( \1104 , \1099 , \1103 );
xor \U$972 ( \1105 , \1090 , \1104 );
and \U$973 ( \1106 , \197 , \230 );
and \U$974 ( \1107 , \178 , \228 );
nor \U$975 ( \1108 , \1106 , \1107 );
xnor \U$976 ( \1109 , \1108 , \237 );
and \U$977 ( \1110 , \217 , \245 );
and \U$978 ( \1111 , \189 , \243 );
nor \U$979 ( \1112 , \1110 , \1111 );
xnor \U$980 ( \1113 , \1112 , \252 );
xor \U$981 ( \1114 , \1109 , \1113 );
and \U$982 ( \1115 , \232 , \141 );
and \U$983 ( \1116 , \209 , \139 );
nor \U$984 ( \1117 , \1115 , \1116 );
xnor \U$985 ( \1118 , \1117 , \148 );
xor \U$986 ( \1119 , \1114 , \1118 );
xor \U$987 ( \1120 , \1105 , \1119 );
xor \U$988 ( \1121 , \1083 , \1120 );
xor \U$989 ( \1122 , \1074 , \1121 );
and \U$990 ( \1123 , \477 , \481 );
and \U$991 ( \1124 , \481 , \487 );
and \U$992 ( \1125 , \477 , \487 );
or \U$993 ( \1126 , \1123 , \1124 , \1125 );
and \U$994 ( \1127 , \515 , \519 );
and \U$995 ( \1128 , \519 , \524 );
and \U$996 ( \1129 , \515 , \524 );
or \U$997 ( \1130 , \1127 , \1128 , \1129 );
xor \U$998 ( \1131 , \1126 , \1130 );
and \U$999 ( \1132 , \460 , \464 );
and \U$1000 ( \1133 , \464 , \469 );
and \U$1001 ( \1134 , \460 , \469 );
or \U$1002 ( \1135 , \1132 , \1133 , \1134 );
xor \U$1003 ( \1136 , \1131 , \1135 );
and \U$1004 ( \1137 , \492 , \496 );
and \U$1005 ( \1138 , \496 , \501 );
and \U$1006 ( \1139 , \492 , \501 );
or \U$1007 ( \1140 , \1137 , \1138 , \1139 );
and \U$1008 ( \1141 , \507 , \510 );
and \U$1009 ( \1142 , \510 , \525 );
and \U$1010 ( \1143 , \507 , \525 );
or \U$1011 ( \1144 , \1141 , \1142 , \1143 );
xor \U$1012 ( \1145 , \1140 , \1144 );
and \U$1013 ( \1146 , \474 , \183 );
buf \U$1014 ( \1147 , RIb55dd20_109);
and \U$1015 ( \1148 , \1147 , \180 );
nor \U$1016 ( \1149 , \1146 , \1148 );
xnor \U$1017 ( \1150 , \1149 , \179 );
and \U$1018 ( \1151 , \307 , \195 );
and \U$1019 ( \1152 , \412 , \193 );
nor \U$1020 ( \1153 , \1151 , \1152 );
xnor \U$1021 ( \1154 , \1153 , \202 );
xor \U$1022 ( \1155 , \1150 , \1154 );
and \U$1023 ( \1156 , \185 , \215 );
and \U$1024 ( \1157 , \261 , \213 );
nor \U$1025 ( \1158 , \1156 , \1157 );
xnor \U$1026 ( \1159 , \1158 , \222 );
xor \U$1027 ( \1160 , \1155 , \1159 );
xor \U$1028 ( \1161 , \1145 , \1160 );
xor \U$1029 ( \1162 , \1136 , \1161 );
xor \U$1030 ( \1163 , \1122 , \1162 );
and \U$1031 ( \1164 , \387 , \528 );
xor \U$1032 ( \1165 , \1163 , \1164 );
and \U$1033 ( \1166 , \529 , \534 );
and \U$1034 ( \1167 , \535 , \1067 );
or \U$1035 ( \1168 , \1166 , \1167 );
xor \U$1036 ( \1169 , \1165 , \1168 );
buf g5575_GF_PartitionCandidate( \1170_nG5575 , \1169 );
buf \U$1037 ( \1171 , \1170_nG5575 );
and \U$1038 ( \1172 , \1078 , \1082 );
and \U$1039 ( \1173 , \1082 , \1120 );
and \U$1040 ( \1174 , \1078 , \1120 );
or \U$1041 ( \1175 , \1172 , \1173 , \1174 );
and \U$1042 ( \1176 , \1136 , \1161 );
xor \U$1043 ( \1177 , \1175 , \1176 );
and \U$1044 ( \1178 , \1140 , \1144 );
and \U$1045 ( \1179 , \1144 , \1160 );
and \U$1046 ( \1180 , \1140 , \1160 );
or \U$1047 ( \1181 , \1178 , \1179 , \1180 );
and \U$1048 ( \1182 , \1126 , \1130 );
and \U$1049 ( \1183 , \1130 , \1135 );
and \U$1050 ( \1184 , \1126 , \1135 );
or \U$1051 ( \1185 , \1182 , \1183 , \1184 );
and \U$1052 ( \1186 , \1090 , \1104 );
and \U$1053 ( \1187 , \1104 , \1119 );
and \U$1054 ( \1188 , \1090 , \1119 );
or \U$1055 ( \1189 , \1186 , \1187 , \1188 );
xor \U$1056 ( \1190 , \1185 , \1189 );
and \U$1057 ( \1191 , \1147 , \183 );
buf \U$1058 ( \1192 , RIb55dd98_108);
and \U$1059 ( \1193 , \1192 , \180 );
nor \U$1060 ( \1194 , \1191 , \1193 );
xnor \U$1061 ( \1195 , \1194 , \179 );
and \U$1062 ( \1196 , \412 , \195 );
and \U$1063 ( \1197 , \474 , \193 );
nor \U$1064 ( \1198 , \1196 , \1197 );
xnor \U$1065 ( \1199 , \1198 , \202 );
xor \U$1066 ( \1200 , \1195 , \1199 );
buf \U$1067 ( \1201 , RIb55fc10_43);
buf \U$1068 ( \1202 , RIb55fb98_44);
and \U$1069 ( \1203 , \1202 , \483 );
not \U$1070 ( \1204 , \1203 );
and \U$1071 ( \1205 , \1201 , \1204 );
xor \U$1072 ( \1206 , \1200 , \1205 );
xor \U$1073 ( \1207 , \1190 , \1206 );
xor \U$1074 ( \1208 , \1181 , \1207 );
and \U$1075 ( \1209 , \1094 , \1098 );
and \U$1076 ( \1210 , \1098 , \1103 );
and \U$1077 ( \1211 , \1094 , \1103 );
or \U$1078 ( \1212 , \1209 , \1210 , \1211 );
and \U$1079 ( \1213 , \1150 , \1154 );
and \U$1080 ( \1214 , \1154 , \1159 );
and \U$1081 ( \1215 , \1150 , \1159 );
or \U$1082 ( \1216 , \1213 , \1214 , \1215 );
xor \U$1083 ( \1217 , \1212 , \1216 );
and \U$1084 ( \1218 , \1109 , \1113 );
and \U$1085 ( \1219 , \1113 , \1118 );
and \U$1086 ( \1220 , \1109 , \1118 );
or \U$1087 ( \1221 , \1218 , \1219 , \1220 );
xor \U$1088 ( \1222 , \1217 , \1221 );
and \U$1089 ( \1223 , \261 , \215 );
and \U$1090 ( \1224 , \307 , \213 );
nor \U$1091 ( \1225 , \1223 , \1224 );
xnor \U$1092 ( \1226 , \1225 , \222 );
and \U$1093 ( \1227 , \178 , \230 );
and \U$1094 ( \1228 , \185 , \228 );
nor \U$1095 ( \1229 , \1227 , \1228 );
xnor \U$1096 ( \1230 , \1229 , \237 );
xor \U$1097 ( \1231 , \1226 , \1230 );
and \U$1098 ( \1232 , \189 , \245 );
and \U$1099 ( \1233 , \197 , \243 );
nor \U$1100 ( \1234 , \1232 , \1233 );
xnor \U$1101 ( \1235 , \1234 , \252 );
xor \U$1102 ( \1236 , \1231 , \1235 );
and \U$1103 ( \1237 , \134 , \438 );
and \U$1104 ( \1238 , \143 , \336 );
nor \U$1105 ( \1239 , \1237 , \1238 );
xnor \U$1106 ( \1240 , \1239 , \320 );
and \U$1107 ( \1241 , \150 , \1086 );
and \U$1108 ( \1242 , \158 , \508 );
nor \U$1109 ( \1243 , \1241 , \1242 );
xnor \U$1110 ( \1244 , \1243 , \487 );
xor \U$1111 ( \1245 , \1240 , \1244 );
xor \U$1112 ( \1246 , \1202 , \483 );
nand \U$1113 ( \1247 , \166 , \1246 );
xnor \U$1114 ( \1248 , \1247 , \1205 );
xor \U$1115 ( \1249 , \1245 , \1248 );
xor \U$1116 ( \1250 , \1236 , \1249 );
and \U$1117 ( \1251 , \209 , \141 );
and \U$1118 ( \1252 , \217 , \139 );
nor \U$1119 ( \1253 , \1251 , \1252 );
xnor \U$1120 ( \1254 , \1253 , \148 );
and \U$1121 ( \1255 , \224 , \156 );
and \U$1122 ( \1256 , \232 , \154 );
nor \U$1123 ( \1257 , \1255 , \1256 );
xnor \U$1124 ( \1258 , \1257 , \163 );
xor \U$1125 ( \1259 , \1254 , \1258 );
and \U$1126 ( \1260 , \240 , \296 );
and \U$1127 ( \1261 , \247 , \168 );
nor \U$1128 ( \1262 , \1260 , \1261 );
xnor \U$1129 ( \1263 , \1262 , \173 );
xor \U$1130 ( \1264 , \1259 , \1263 );
xor \U$1131 ( \1265 , \1250 , \1264 );
xor \U$1132 ( \1266 , \1222 , \1265 );
xor \U$1133 ( \1267 , \1208 , \1266 );
xor \U$1134 ( \1268 , \1177 , \1267 );
and \U$1135 ( \1269 , \1074 , \1121 );
and \U$1136 ( \1270 , \1121 , \1162 );
and \U$1137 ( \1271 , \1074 , \1162 );
or \U$1138 ( \1272 , \1269 , \1270 , \1271 );
xor \U$1139 ( \1273 , \1268 , \1272 );
and \U$1140 ( \1274 , \1163 , \1164 );
and \U$1141 ( \1275 , \1165 , \1168 );
or \U$1142 ( \1276 , \1274 , \1275 );
xor \U$1143 ( \1277 , \1273 , \1276 );
buf g5573_GF_PartitionCandidate( \1278_nG5573 , \1277 );
buf \U$1144 ( \1279 , \1278_nG5573 );
and \U$1145 ( \1280 , \1181 , \1207 );
and \U$1146 ( \1281 , \1207 , \1266 );
and \U$1147 ( \1282 , \1181 , \1266 );
or \U$1148 ( \1283 , \1280 , \1281 , \1282 );
and \U$1149 ( \1284 , \1185 , \1189 );
and \U$1150 ( \1285 , \1189 , \1206 );
and \U$1151 ( \1286 , \1185 , \1206 );
or \U$1152 ( \1287 , \1284 , \1285 , \1286 );
and \U$1153 ( \1288 , \1222 , \1265 );
xor \U$1154 ( \1289 , \1287 , \1288 );
and \U$1155 ( \1290 , \1240 , \1244 );
and \U$1156 ( \1291 , \1244 , \1248 );
and \U$1157 ( \1292 , \1240 , \1248 );
or \U$1158 ( \1293 , \1290 , \1291 , \1292 );
and \U$1159 ( \1294 , \158 , \1086 );
and \U$1160 ( \1295 , \134 , \508 );
nor \U$1161 ( \1296 , \1294 , \1295 );
xnor \U$1162 ( \1297 , \1296 , \487 );
xor \U$1163 ( \1298 , \1293 , \1297 );
xor \U$1164 ( \1299 , \1201 , \1202 );
not \U$1165 ( \1300 , \1246 );
and \U$1166 ( \1301 , \1299 , \1300 );
and \U$1167 ( \1302 , \166 , \1301 );
and \U$1168 ( \1303 , \150 , \1246 );
nor \U$1169 ( \1304 , \1302 , \1303 );
xnor \U$1170 ( \1305 , \1304 , \1205 );
xor \U$1171 ( \1306 , \1298 , \1305 );
xor \U$1172 ( \1307 , \1289 , \1306 );
xor \U$1173 ( \1308 , \1283 , \1307 );
and \U$1174 ( \1309 , \1195 , \1199 );
and \U$1175 ( \1310 , \1199 , \1205 );
and \U$1176 ( \1311 , \1195 , \1205 );
or \U$1177 ( \1312 , \1309 , \1310 , \1311 );
and \U$1178 ( \1313 , \1226 , \1230 );
and \U$1179 ( \1314 , \1230 , \1235 );
and \U$1180 ( \1315 , \1226 , \1235 );
or \U$1181 ( \1316 , \1313 , \1314 , \1315 );
xor \U$1182 ( \1317 , \1312 , \1316 );
and \U$1183 ( \1318 , \1254 , \1258 );
and \U$1184 ( \1319 , \1258 , \1263 );
and \U$1185 ( \1320 , \1254 , \1263 );
or \U$1186 ( \1321 , \1318 , \1319 , \1320 );
xor \U$1187 ( \1322 , \1317 , \1321 );
and \U$1188 ( \1323 , \1212 , \1216 );
and \U$1189 ( \1324 , \1216 , \1221 );
and \U$1190 ( \1325 , \1212 , \1221 );
or \U$1191 ( \1326 , \1323 , \1324 , \1325 );
and \U$1192 ( \1327 , \1236 , \1249 );
and \U$1193 ( \1328 , \1249 , \1264 );
and \U$1194 ( \1329 , \1236 , \1264 );
or \U$1195 ( \1330 , \1327 , \1328 , \1329 );
xor \U$1196 ( \1331 , \1326 , \1330 );
and \U$1197 ( \1332 , \1192 , \183 );
buf \U$1198 ( \1333 , RIb55de10_107);
and \U$1199 ( \1334 , \1333 , \180 );
nor \U$1200 ( \1335 , \1332 , \1334 );
xnor \U$1201 ( \1336 , \1335 , \179 );
and \U$1202 ( \1337 , \474 , \195 );
and \U$1203 ( \1338 , \1147 , \193 );
nor \U$1204 ( \1339 , \1337 , \1338 );
xnor \U$1205 ( \1340 , \1339 , \202 );
xor \U$1206 ( \1341 , \1336 , \1340 );
and \U$1207 ( \1342 , \307 , \215 );
and \U$1208 ( \1343 , \412 , \213 );
nor \U$1209 ( \1344 , \1342 , \1343 );
xnor \U$1210 ( \1345 , \1344 , \222 );
xor \U$1211 ( \1346 , \1341 , \1345 );
and \U$1212 ( \1347 , \232 , \156 );
and \U$1213 ( \1348 , \209 , \154 );
nor \U$1214 ( \1349 , \1347 , \1348 );
xnor \U$1215 ( \1350 , \1349 , \163 );
and \U$1216 ( \1351 , \247 , \296 );
and \U$1217 ( \1352 , \224 , \168 );
nor \U$1218 ( \1353 , \1351 , \1352 );
xnor \U$1219 ( \1354 , \1353 , \173 );
xor \U$1220 ( \1355 , \1350 , \1354 );
and \U$1221 ( \1356 , \143 , \438 );
and \U$1222 ( \1357 , \240 , \336 );
nor \U$1223 ( \1358 , \1356 , \1357 );
xnor \U$1224 ( \1359 , \1358 , \320 );
xor \U$1225 ( \1360 , \1355 , \1359 );
xor \U$1226 ( \1361 , \1346 , \1360 );
and \U$1227 ( \1362 , \185 , \230 );
and \U$1228 ( \1363 , \261 , \228 );
nor \U$1229 ( \1364 , \1362 , \1363 );
xnor \U$1230 ( \1365 , \1364 , \237 );
and \U$1231 ( \1366 , \197 , \245 );
and \U$1232 ( \1367 , \178 , \243 );
nor \U$1233 ( \1368 , \1366 , \1367 );
xnor \U$1234 ( \1369 , \1368 , \252 );
xor \U$1235 ( \1370 , \1365 , \1369 );
and \U$1236 ( \1371 , \217 , \141 );
and \U$1237 ( \1372 , \189 , \139 );
nor \U$1238 ( \1373 , \1371 , \1372 );
xnor \U$1239 ( \1374 , \1373 , \148 );
xor \U$1240 ( \1375 , \1370 , \1374 );
xor \U$1241 ( \1376 , \1361 , \1375 );
xor \U$1242 ( \1377 , \1331 , \1376 );
xor \U$1243 ( \1378 , \1322 , \1377 );
xor \U$1244 ( \1379 , \1308 , \1378 );
and \U$1245 ( \1380 , \1175 , \1176 );
and \U$1246 ( \1381 , \1176 , \1267 );
and \U$1247 ( \1382 , \1175 , \1267 );
or \U$1248 ( \1383 , \1380 , \1381 , \1382 );
xor \U$1249 ( \1384 , \1379 , \1383 );
and \U$1250 ( \1385 , \1268 , \1272 );
and \U$1251 ( \1386 , \1273 , \1276 );
or \U$1252 ( \1387 , \1385 , \1386 );
xor \U$1253 ( \1388 , \1384 , \1387 );
buf g5571_GF_PartitionCandidate( \1389_nG5571 , \1388 );
buf \U$1254 ( \1390 , \1389_nG5571 );
and \U$1255 ( \1391 , \1287 , \1288 );
and \U$1256 ( \1392 , \1288 , \1306 );
and \U$1257 ( \1393 , \1287 , \1306 );
or \U$1258 ( \1394 , \1391 , \1392 , \1393 );
and \U$1259 ( \1395 , \1322 , \1377 );
xor \U$1260 ( \1396 , \1394 , \1395 );
and \U$1261 ( \1397 , \1326 , \1330 );
and \U$1262 ( \1398 , \1330 , \1376 );
and \U$1263 ( \1399 , \1326 , \1376 );
or \U$1264 ( \1400 , \1397 , \1398 , \1399 );
and \U$1265 ( \1401 , \1293 , \1297 );
and \U$1266 ( \1402 , \1297 , \1305 );
and \U$1267 ( \1403 , \1293 , \1305 );
or \U$1268 ( \1404 , \1401 , \1402 , \1403 );
and \U$1269 ( \1405 , \1312 , \1316 );
and \U$1270 ( \1406 , \1316 , \1321 );
and \U$1271 ( \1407 , \1312 , \1321 );
or \U$1272 ( \1408 , \1405 , \1406 , \1407 );
xor \U$1273 ( \1409 , \1404 , \1408 );
and \U$1274 ( \1410 , \1346 , \1360 );
and \U$1275 ( \1411 , \1360 , \1375 );
and \U$1276 ( \1412 , \1346 , \1375 );
or \U$1277 ( \1413 , \1410 , \1411 , \1412 );
xor \U$1278 ( \1414 , \1409 , \1413 );
xor \U$1279 ( \1415 , \1400 , \1414 );
and \U$1280 ( \1416 , \1336 , \1340 );
and \U$1281 ( \1417 , \1340 , \1345 );
and \U$1282 ( \1418 , \1336 , \1345 );
or \U$1283 ( \1419 , \1416 , \1417 , \1418 );
and \U$1284 ( \1420 , \1350 , \1354 );
and \U$1285 ( \1421 , \1354 , \1359 );
and \U$1286 ( \1422 , \1350 , \1359 );
or \U$1287 ( \1423 , \1420 , \1421 , \1422 );
xor \U$1288 ( \1424 , \1419 , \1423 );
and \U$1289 ( \1425 , \1365 , \1369 );
and \U$1290 ( \1426 , \1369 , \1374 );
and \U$1291 ( \1427 , \1365 , \1374 );
or \U$1292 ( \1428 , \1425 , \1426 , \1427 );
xor \U$1293 ( \1429 , \1424 , \1428 );
buf \U$1294 ( \1430 , RIb55fc88_42);
xor \U$1295 ( \1431 , \1430 , \1201 );
nand \U$1296 ( \1432 , \166 , \1431 );
buf \U$1297 ( \1433 , RIb55fd00_41);
and \U$1298 ( \1434 , \1430 , \1201 );
not \U$1299 ( \1435 , \1434 );
and \U$1300 ( \1436 , \1433 , \1435 );
xnor \U$1301 ( \1437 , \1432 , \1436 );
and \U$1302 ( \1438 , \189 , \141 );
and \U$1303 ( \1439 , \197 , \139 );
nor \U$1304 ( \1440 , \1438 , \1439 );
xnor \U$1305 ( \1441 , \1440 , \148 );
and \U$1306 ( \1442 , \209 , \156 );
and \U$1307 ( \1443 , \217 , \154 );
nor \U$1308 ( \1444 , \1442 , \1443 );
xnor \U$1309 ( \1445 , \1444 , \163 );
xor \U$1310 ( \1446 , \1441 , \1445 );
and \U$1311 ( \1447 , \224 , \296 );
and \U$1312 ( \1448 , \232 , \168 );
nor \U$1313 ( \1449 , \1447 , \1448 );
xnor \U$1314 ( \1450 , \1449 , \173 );
xor \U$1315 ( \1451 , \1446 , \1450 );
xor \U$1316 ( \1452 , \1437 , \1451 );
and \U$1317 ( \1453 , \240 , \438 );
and \U$1318 ( \1454 , \247 , \336 );
nor \U$1319 ( \1455 , \1453 , \1454 );
xnor \U$1320 ( \1456 , \1455 , \320 );
and \U$1321 ( \1457 , \134 , \1086 );
and \U$1322 ( \1458 , \143 , \508 );
nor \U$1323 ( \1459 , \1457 , \1458 );
xnor \U$1324 ( \1460 , \1459 , \487 );
xor \U$1325 ( \1461 , \1456 , \1460 );
and \U$1326 ( \1462 , \150 , \1301 );
and \U$1327 ( \1463 , \158 , \1246 );
nor \U$1328 ( \1464 , \1462 , \1463 );
xnor \U$1329 ( \1465 , \1464 , \1205 );
xor \U$1330 ( \1466 , \1461 , \1465 );
xor \U$1331 ( \1467 , \1452 , \1466 );
xor \U$1332 ( \1468 , \1429 , \1467 );
and \U$1333 ( \1469 , \412 , \215 );
and \U$1334 ( \1470 , \474 , \213 );
nor \U$1335 ( \1471 , \1469 , \1470 );
xnor \U$1336 ( \1472 , \1471 , \222 );
and \U$1337 ( \1473 , \261 , \230 );
and \U$1338 ( \1474 , \307 , \228 );
nor \U$1339 ( \1475 , \1473 , \1474 );
xnor \U$1340 ( \1476 , \1475 , \237 );
xor \U$1341 ( \1477 , \1472 , \1476 );
and \U$1342 ( \1478 , \178 , \245 );
and \U$1343 ( \1479 , \185 , \243 );
nor \U$1344 ( \1480 , \1478 , \1479 );
xnor \U$1345 ( \1481 , \1480 , \252 );
xor \U$1346 ( \1482 , \1477 , \1481 );
and \U$1347 ( \1483 , \1333 , \183 );
buf \U$1348 ( \1484 , RIb55de88_106);
and \U$1349 ( \1485 , \1484 , \180 );
nor \U$1350 ( \1486 , \1483 , \1485 );
xnor \U$1351 ( \1487 , \1486 , \179 );
and \U$1352 ( \1488 , \1147 , \195 );
and \U$1353 ( \1489 , \1192 , \193 );
nor \U$1354 ( \1490 , \1488 , \1489 );
xnor \U$1355 ( \1491 , \1490 , \202 );
xor \U$1356 ( \1492 , \1487 , \1491 );
xor \U$1357 ( \1493 , \1492 , \1436 );
xor \U$1358 ( \1494 , \1482 , \1493 );
xor \U$1359 ( \1495 , \1468 , \1494 );
xor \U$1360 ( \1496 , \1415 , \1495 );
xor \U$1361 ( \1497 , \1396 , \1496 );
and \U$1362 ( \1498 , \1283 , \1307 );
and \U$1363 ( \1499 , \1307 , \1378 );
and \U$1364 ( \1500 , \1283 , \1378 );
or \U$1365 ( \1501 , \1498 , \1499 , \1500 );
xor \U$1366 ( \1502 , \1497 , \1501 );
and \U$1367 ( \1503 , \1379 , \1383 );
and \U$1368 ( \1504 , \1384 , \1387 );
or \U$1369 ( \1505 , \1503 , \1504 );
xor \U$1370 ( \1506 , \1502 , \1505 );
buf g556f_GF_PartitionCandidate( \1507_nG556f , \1506 );
buf \U$1371 ( \1508 , \1507_nG556f );
and \U$1372 ( \1509 , \1400 , \1414 );
and \U$1373 ( \1510 , \1414 , \1495 );
and \U$1374 ( \1511 , \1400 , \1495 );
or \U$1375 ( \1512 , \1509 , \1510 , \1511 );
and \U$1376 ( \1513 , \1419 , \1423 );
and \U$1377 ( \1514 , \1423 , \1428 );
and \U$1378 ( \1515 , \1419 , \1428 );
or \U$1379 ( \1516 , \1513 , \1514 , \1515 );
and \U$1380 ( \1517 , \1437 , \1451 );
and \U$1381 ( \1518 , \1451 , \1466 );
and \U$1382 ( \1519 , \1437 , \1466 );
or \U$1383 ( \1520 , \1517 , \1518 , \1519 );
xor \U$1384 ( \1521 , \1516 , \1520 );
and \U$1385 ( \1522 , \1482 , \1493 );
xor \U$1386 ( \1523 , \1521 , \1522 );
xor \U$1387 ( \1524 , \1512 , \1523 );
and \U$1388 ( \1525 , \1404 , \1408 );
and \U$1389 ( \1526 , \1408 , \1413 );
and \U$1390 ( \1527 , \1404 , \1413 );
or \U$1391 ( \1528 , \1525 , \1526 , \1527 );
and \U$1392 ( \1529 , \1429 , \1467 );
and \U$1393 ( \1530 , \1467 , \1494 );
and \U$1394 ( \1531 , \1429 , \1494 );
or \U$1395 ( \1532 , \1529 , \1530 , \1531 );
xor \U$1396 ( \1533 , \1528 , \1532 );
and \U$1397 ( \1534 , \1472 , \1476 );
and \U$1398 ( \1535 , \1476 , \1481 );
and \U$1399 ( \1536 , \1472 , \1481 );
or \U$1400 ( \1537 , \1534 , \1535 , \1536 );
and \U$1401 ( \1538 , \1441 , \1445 );
and \U$1402 ( \1539 , \1445 , \1450 );
and \U$1403 ( \1540 , \1441 , \1450 );
or \U$1404 ( \1541 , \1538 , \1539 , \1540 );
xor \U$1405 ( \1542 , \1537 , \1541 );
and \U$1406 ( \1543 , \1487 , \1491 );
and \U$1407 ( \1544 , \1491 , \1436 );
and \U$1408 ( \1545 , \1487 , \1436 );
or \U$1409 ( \1546 , \1543 , \1544 , \1545 );
xor \U$1410 ( \1547 , \1542 , \1546 );
and \U$1411 ( \1548 , \1456 , \1460 );
and \U$1412 ( \1549 , \1460 , \1465 );
and \U$1413 ( \1550 , \1456 , \1465 );
or \U$1414 ( \1551 , \1548 , \1549 , \1550 );
and \U$1415 ( \1552 , \217 , \156 );
and \U$1416 ( \1553 , \189 , \154 );
nor \U$1417 ( \1554 , \1552 , \1553 );
xnor \U$1418 ( \1555 , \1554 , \163 );
and \U$1419 ( \1556 , \232 , \296 );
and \U$1420 ( \1557 , \209 , \168 );
nor \U$1421 ( \1558 , \1556 , \1557 );
xnor \U$1422 ( \1559 , \1558 , \173 );
xor \U$1423 ( \1560 , \1555 , \1559 );
and \U$1424 ( \1561 , \247 , \438 );
and \U$1425 ( \1562 , \224 , \336 );
nor \U$1426 ( \1563 , \1561 , \1562 );
xnor \U$1427 ( \1564 , \1563 , \320 );
xor \U$1428 ( \1565 , \1560 , \1564 );
xor \U$1429 ( \1566 , \1551 , \1565 );
and \U$1430 ( \1567 , \143 , \1086 );
and \U$1431 ( \1568 , \240 , \508 );
nor \U$1432 ( \1569 , \1567 , \1568 );
xnor \U$1433 ( \1570 , \1569 , \487 );
and \U$1434 ( \1571 , \158 , \1301 );
and \U$1435 ( \1572 , \134 , \1246 );
nor \U$1436 ( \1573 , \1571 , \1572 );
xnor \U$1437 ( \1574 , \1573 , \1205 );
xor \U$1438 ( \1575 , \1570 , \1574 );
xor \U$1439 ( \1576 , \1433 , \1430 );
not \U$1440 ( \1577 , \1431 );
and \U$1441 ( \1578 , \1576 , \1577 );
and \U$1442 ( \1579 , \166 , \1578 );
and \U$1443 ( \1580 , \150 , \1431 );
nor \U$1444 ( \1581 , \1579 , \1580 );
xnor \U$1445 ( \1582 , \1581 , \1436 );
xor \U$1446 ( \1583 , \1575 , \1582 );
xor \U$1447 ( \1584 , \1566 , \1583 );
xor \U$1448 ( \1585 , \1547 , \1584 );
and \U$1449 ( \1586 , \307 , \230 );
and \U$1450 ( \1587 , \412 , \228 );
nor \U$1451 ( \1588 , \1586 , \1587 );
xnor \U$1452 ( \1589 , \1588 , \237 );
and \U$1453 ( \1590 , \185 , \245 );
and \U$1454 ( \1591 , \261 , \243 );
nor \U$1455 ( \1592 , \1590 , \1591 );
xnor \U$1456 ( \1593 , \1592 , \252 );
xor \U$1457 ( \1594 , \1589 , \1593 );
and \U$1458 ( \1595 , \197 , \141 );
and \U$1459 ( \1596 , \178 , \139 );
nor \U$1460 ( \1597 , \1595 , \1596 );
xnor \U$1461 ( \1598 , \1597 , \148 );
xor \U$1462 ( \1599 , \1594 , \1598 );
and \U$1463 ( \1600 , \1484 , \183 );
buf \U$1464 ( \1601 , RIb55df00_105);
and \U$1465 ( \1602 , \1601 , \180 );
nor \U$1466 ( \1603 , \1600 , \1602 );
xnor \U$1467 ( \1604 , \1603 , \179 );
and \U$1468 ( \1605 , \1192 , \195 );
and \U$1469 ( \1606 , \1333 , \193 );
nor \U$1470 ( \1607 , \1605 , \1606 );
xnor \U$1471 ( \1608 , \1607 , \202 );
xor \U$1472 ( \1609 , \1604 , \1608 );
and \U$1473 ( \1610 , \474 , \215 );
and \U$1474 ( \1611 , \1147 , \213 );
nor \U$1475 ( \1612 , \1610 , \1611 );
xnor \U$1476 ( \1613 , \1612 , \222 );
xor \U$1477 ( \1614 , \1609 , \1613 );
xor \U$1478 ( \1615 , \1599 , \1614 );
xor \U$1479 ( \1616 , \1585 , \1615 );
xor \U$1480 ( \1617 , \1533 , \1616 );
xor \U$1481 ( \1618 , \1524 , \1617 );
and \U$1482 ( \1619 , \1394 , \1395 );
and \U$1483 ( \1620 , \1395 , \1496 );
and \U$1484 ( \1621 , \1394 , \1496 );
or \U$1485 ( \1622 , \1619 , \1620 , \1621 );
xor \U$1486 ( \1623 , \1618 , \1622 );
and \U$1487 ( \1624 , \1497 , \1501 );
and \U$1488 ( \1625 , \1502 , \1505 );
or \U$1489 ( \1626 , \1624 , \1625 );
xor \U$1490 ( \1627 , \1623 , \1626 );
buf g556d_GF_PartitionCandidate( \1628_nG556d , \1627 );
buf \U$1491 ( \1629 , \1628_nG556d );
and \U$1492 ( \1630 , \1528 , \1532 );
and \U$1493 ( \1631 , \1532 , \1616 );
and \U$1494 ( \1632 , \1528 , \1616 );
or \U$1495 ( \1633 , \1630 , \1631 , \1632 );
and \U$1496 ( \1634 , \1537 , \1541 );
and \U$1497 ( \1635 , \1541 , \1546 );
and \U$1498 ( \1636 , \1537 , \1546 );
or \U$1499 ( \1637 , \1634 , \1635 , \1636 );
and \U$1500 ( \1638 , \1551 , \1565 );
and \U$1501 ( \1639 , \1565 , \1583 );
and \U$1502 ( \1640 , \1551 , \1583 );
or \U$1503 ( \1641 , \1638 , \1639 , \1640 );
xor \U$1504 ( \1642 , \1637 , \1641 );
and \U$1505 ( \1643 , \1599 , \1614 );
xor \U$1506 ( \1644 , \1642 , \1643 );
xor \U$1507 ( \1645 , \1633 , \1644 );
and \U$1508 ( \1646 , \1516 , \1520 );
and \U$1509 ( \1647 , \1520 , \1522 );
and \U$1510 ( \1648 , \1516 , \1522 );
or \U$1511 ( \1649 , \1646 , \1647 , \1648 );
and \U$1512 ( \1650 , \1547 , \1584 );
and \U$1513 ( \1651 , \1584 , \1615 );
and \U$1514 ( \1652 , \1547 , \1615 );
or \U$1515 ( \1653 , \1650 , \1651 , \1652 );
xor \U$1516 ( \1654 , \1649 , \1653 );
and \U$1517 ( \1655 , \1589 , \1593 );
and \U$1518 ( \1656 , \1593 , \1598 );
and \U$1519 ( \1657 , \1589 , \1598 );
or \U$1520 ( \1658 , \1655 , \1656 , \1657 );
and \U$1521 ( \1659 , \1555 , \1559 );
and \U$1522 ( \1660 , \1559 , \1564 );
and \U$1523 ( \1661 , \1555 , \1564 );
or \U$1524 ( \1662 , \1659 , \1660 , \1661 );
xor \U$1525 ( \1663 , \1658 , \1662 );
and \U$1526 ( \1664 , \1604 , \1608 );
and \U$1527 ( \1665 , \1608 , \1613 );
and \U$1528 ( \1666 , \1604 , \1613 );
or \U$1529 ( \1667 , \1664 , \1665 , \1666 );
xor \U$1530 ( \1668 , \1663 , \1667 );
and \U$1531 ( \1669 , \1147 , \215 );
and \U$1532 ( \1670 , \1192 , \213 );
nor \U$1533 ( \1671 , \1669 , \1670 );
xnor \U$1534 ( \1672 , \1671 , \222 );
and \U$1535 ( \1673 , \412 , \230 );
and \U$1536 ( \1674 , \474 , \228 );
nor \U$1537 ( \1675 , \1673 , \1674 );
xnor \U$1538 ( \1676 , \1675 , \237 );
xor \U$1539 ( \1677 , \1672 , \1676 );
and \U$1540 ( \1678 , \261 , \245 );
and \U$1541 ( \1679 , \307 , \243 );
nor \U$1542 ( \1680 , \1678 , \1679 );
xnor \U$1543 ( \1681 , \1680 , \252 );
xor \U$1544 ( \1682 , \1677 , \1681 );
and \U$1545 ( \1683 , \1601 , \183 );
buf \U$1546 ( \1684 , RIb55df78_104);
and \U$1547 ( \1685 , \1684 , \180 );
nor \U$1548 ( \1686 , \1683 , \1685 );
xnor \U$1549 ( \1687 , \1686 , \179 );
and \U$1550 ( \1688 , \1333 , \195 );
and \U$1551 ( \1689 , \1484 , \193 );
nor \U$1552 ( \1690 , \1688 , \1689 );
xnor \U$1553 ( \1691 , \1690 , \202 );
xor \U$1554 ( \1692 , \1687 , \1691 );
buf \U$1555 ( \1693 , RIb55fdf0_39);
buf \U$1556 ( \1694 , RIb55fd78_40);
and \U$1557 ( \1695 , \1694 , \1433 );
not \U$1558 ( \1696 , \1695 );
and \U$1559 ( \1697 , \1693 , \1696 );
xor \U$1560 ( \1698 , \1692 , \1697 );
xor \U$1561 ( \1699 , \1682 , \1698 );
and \U$1562 ( \1700 , \178 , \141 );
and \U$1563 ( \1701 , \185 , \139 );
nor \U$1564 ( \1702 , \1700 , \1701 );
xnor \U$1565 ( \1703 , \1702 , \148 );
and \U$1566 ( \1704 , \189 , \156 );
and \U$1567 ( \1705 , \197 , \154 );
nor \U$1568 ( \1706 , \1704 , \1705 );
xnor \U$1569 ( \1707 , \1706 , \163 );
xor \U$1570 ( \1708 , \1703 , \1707 );
and \U$1571 ( \1709 , \209 , \296 );
and \U$1572 ( \1710 , \217 , \168 );
nor \U$1573 ( \1711 , \1709 , \1710 );
xnor \U$1574 ( \1712 , \1711 , \173 );
xor \U$1575 ( \1713 , \1708 , \1712 );
xor \U$1576 ( \1714 , \1699 , \1713 );
xor \U$1577 ( \1715 , \1668 , \1714 );
and \U$1578 ( \1716 , \1570 , \1574 );
and \U$1579 ( \1717 , \1574 , \1582 );
and \U$1580 ( \1718 , \1570 , \1582 );
or \U$1581 ( \1719 , \1716 , \1717 , \1718 );
and \U$1582 ( \1720 , \224 , \438 );
and \U$1583 ( \1721 , \232 , \336 );
nor \U$1584 ( \1722 , \1720 , \1721 );
xnor \U$1585 ( \1723 , \1722 , \320 );
and \U$1586 ( \1724 , \240 , \1086 );
and \U$1587 ( \1725 , \247 , \508 );
nor \U$1588 ( \1726 , \1724 , \1725 );
xnor \U$1589 ( \1727 , \1726 , \487 );
xor \U$1590 ( \1728 , \1723 , \1727 );
and \U$1591 ( \1729 , \134 , \1301 );
and \U$1592 ( \1730 , \143 , \1246 );
nor \U$1593 ( \1731 , \1729 , \1730 );
xnor \U$1594 ( \1732 , \1731 , \1205 );
xor \U$1595 ( \1733 , \1728 , \1732 );
xor \U$1596 ( \1734 , \1719 , \1733 );
and \U$1597 ( \1735 , \150 , \1578 );
and \U$1598 ( \1736 , \158 , \1431 );
nor \U$1599 ( \1737 , \1735 , \1736 );
xnor \U$1600 ( \1738 , \1737 , \1436 );
xor \U$1601 ( \1739 , \1694 , \1433 );
nand \U$1602 ( \1740 , \166 , \1739 );
xnor \U$1603 ( \1741 , \1740 , \1697 );
xor \U$1604 ( \1742 , \1738 , \1741 );
xor \U$1605 ( \1743 , \1734 , \1742 );
xor \U$1606 ( \1744 , \1715 , \1743 );
xor \U$1607 ( \1745 , \1654 , \1744 );
xor \U$1608 ( \1746 , \1645 , \1745 );
and \U$1609 ( \1747 , \1512 , \1523 );
and \U$1610 ( \1748 , \1523 , \1617 );
and \U$1611 ( \1749 , \1512 , \1617 );
or \U$1612 ( \1750 , \1747 , \1748 , \1749 );
xor \U$1613 ( \1751 , \1746 , \1750 );
and \U$1614 ( \1752 , \1618 , \1622 );
and \U$1615 ( \1753 , \1623 , \1626 );
or \U$1616 ( \1754 , \1752 , \1753 );
xor \U$1617 ( \1755 , \1751 , \1754 );
buf g556b_GF_PartitionCandidate( \1756_nG556b , \1755 );
buf \U$1618 ( \1757 , \1756_nG556b );
and \U$1619 ( \1758 , \1649 , \1653 );
and \U$1620 ( \1759 , \1653 , \1744 );
and \U$1621 ( \1760 , \1649 , \1744 );
or \U$1622 ( \1761 , \1758 , \1759 , \1760 );
and \U$1623 ( \1762 , \1637 , \1641 );
and \U$1624 ( \1763 , \1641 , \1643 );
and \U$1625 ( \1764 , \1637 , \1643 );
or \U$1626 ( \1765 , \1762 , \1763 , \1764 );
and \U$1627 ( \1766 , \1668 , \1714 );
and \U$1628 ( \1767 , \1714 , \1743 );
and \U$1629 ( \1768 , \1668 , \1743 );
or \U$1630 ( \1769 , \1766 , \1767 , \1768 );
xor \U$1631 ( \1770 , \1765 , \1769 );
and \U$1632 ( \1771 , \1672 , \1676 );
and \U$1633 ( \1772 , \1676 , \1681 );
and \U$1634 ( \1773 , \1672 , \1681 );
or \U$1635 ( \1774 , \1771 , \1772 , \1773 );
and \U$1636 ( \1775 , \1687 , \1691 );
and \U$1637 ( \1776 , \1691 , \1697 );
and \U$1638 ( \1777 , \1687 , \1697 );
or \U$1639 ( \1778 , \1775 , \1776 , \1777 );
xor \U$1640 ( \1779 , \1774 , \1778 );
and \U$1641 ( \1780 , \1703 , \1707 );
and \U$1642 ( \1781 , \1707 , \1712 );
and \U$1643 ( \1782 , \1703 , \1712 );
or \U$1644 ( \1783 , \1780 , \1781 , \1782 );
xor \U$1645 ( \1784 , \1779 , \1783 );
xor \U$1646 ( \1785 , \1770 , \1784 );
xor \U$1647 ( \1786 , \1761 , \1785 );
and \U$1648 ( \1787 , \1658 , \1662 );
and \U$1649 ( \1788 , \1662 , \1667 );
and \U$1650 ( \1789 , \1658 , \1667 );
or \U$1651 ( \1790 , \1787 , \1788 , \1789 );
and \U$1652 ( \1791 , \1682 , \1698 );
and \U$1653 ( \1792 , \1698 , \1713 );
and \U$1654 ( \1793 , \1682 , \1713 );
or \U$1655 ( \1794 , \1791 , \1792 , \1793 );
xor \U$1656 ( \1795 , \1790 , \1794 );
and \U$1657 ( \1796 , \1719 , \1733 );
and \U$1658 ( \1797 , \1733 , \1742 );
and \U$1659 ( \1798 , \1719 , \1742 );
or \U$1660 ( \1799 , \1796 , \1797 , \1798 );
xor \U$1661 ( \1800 , \1795 , \1799 );
and \U$1662 ( \1801 , \1684 , \183 );
buf \U$1663 ( \1802 , RIb55dff0_103);
and \U$1664 ( \1803 , \1802 , \180 );
nor \U$1665 ( \1804 , \1801 , \1803 );
xnor \U$1666 ( \1805 , \1804 , \179 );
and \U$1667 ( \1806 , \1484 , \195 );
and \U$1668 ( \1807 , \1601 , \193 );
nor \U$1669 ( \1808 , \1806 , \1807 );
xnor \U$1670 ( \1809 , \1808 , \202 );
xor \U$1671 ( \1810 , \1805 , \1809 );
and \U$1672 ( \1811 , \1192 , \215 );
and \U$1673 ( \1812 , \1333 , \213 );
nor \U$1674 ( \1813 , \1811 , \1812 );
xnor \U$1675 ( \1814 , \1813 , \222 );
xor \U$1676 ( \1815 , \1810 , \1814 );
and \U$1677 ( \1816 , \1723 , \1727 );
and \U$1678 ( \1817 , \1727 , \1732 );
and \U$1679 ( \1818 , \1723 , \1732 );
or \U$1680 ( \1819 , \1816 , \1817 , \1818 );
and \U$1681 ( \1820 , \1738 , \1741 );
xor \U$1682 ( \1821 , \1819 , \1820 );
xor \U$1683 ( \1822 , \1693 , \1694 );
not \U$1684 ( \1823 , \1739 );
and \U$1685 ( \1824 , \1822 , \1823 );
and \U$1686 ( \1825 , \166 , \1824 );
and \U$1687 ( \1826 , \150 , \1739 );
nor \U$1688 ( \1827 , \1825 , \1826 );
xnor \U$1689 ( \1828 , \1827 , \1697 );
xor \U$1690 ( \1829 , \1821 , \1828 );
xor \U$1691 ( \1830 , \1815 , \1829 );
and \U$1692 ( \1831 , \474 , \230 );
and \U$1693 ( \1832 , \1147 , \228 );
nor \U$1694 ( \1833 , \1831 , \1832 );
xnor \U$1695 ( \1834 , \1833 , \237 );
and \U$1696 ( \1835 , \307 , \245 );
and \U$1697 ( \1836 , \412 , \243 );
nor \U$1698 ( \1837 , \1835 , \1836 );
xnor \U$1699 ( \1838 , \1837 , \252 );
xor \U$1700 ( \1839 , \1834 , \1838 );
and \U$1701 ( \1840 , \185 , \141 );
and \U$1702 ( \1841 , \261 , \139 );
nor \U$1703 ( \1842 , \1840 , \1841 );
xnor \U$1704 ( \1843 , \1842 , \148 );
xor \U$1705 ( \1844 , \1839 , \1843 );
and \U$1706 ( \1845 , \247 , \1086 );
and \U$1707 ( \1846 , \224 , \508 );
nor \U$1708 ( \1847 , \1845 , \1846 );
xnor \U$1709 ( \1848 , \1847 , \487 );
and \U$1710 ( \1849 , \143 , \1301 );
and \U$1711 ( \1850 , \240 , \1246 );
nor \U$1712 ( \1851 , \1849 , \1850 );
xnor \U$1713 ( \1852 , \1851 , \1205 );
xor \U$1714 ( \1853 , \1848 , \1852 );
and \U$1715 ( \1854 , \158 , \1578 );
and \U$1716 ( \1855 , \134 , \1431 );
nor \U$1717 ( \1856 , \1854 , \1855 );
xnor \U$1718 ( \1857 , \1856 , \1436 );
xor \U$1719 ( \1858 , \1853 , \1857 );
xor \U$1720 ( \1859 , \1844 , \1858 );
and \U$1721 ( \1860 , \197 , \156 );
and \U$1722 ( \1861 , \178 , \154 );
nor \U$1723 ( \1862 , \1860 , \1861 );
xnor \U$1724 ( \1863 , \1862 , \163 );
and \U$1725 ( \1864 , \217 , \296 );
and \U$1726 ( \1865 , \189 , \168 );
nor \U$1727 ( \1866 , \1864 , \1865 );
xnor \U$1728 ( \1867 , \1866 , \173 );
xor \U$1729 ( \1868 , \1863 , \1867 );
and \U$1730 ( \1869 , \232 , \438 );
and \U$1731 ( \1870 , \209 , \336 );
nor \U$1732 ( \1871 , \1869 , \1870 );
xnor \U$1733 ( \1872 , \1871 , \320 );
xor \U$1734 ( \1873 , \1868 , \1872 );
xor \U$1735 ( \1874 , \1859 , \1873 );
xor \U$1736 ( \1875 , \1830 , \1874 );
xor \U$1737 ( \1876 , \1800 , \1875 );
xor \U$1738 ( \1877 , \1786 , \1876 );
and \U$1739 ( \1878 , \1633 , \1644 );
and \U$1740 ( \1879 , \1644 , \1745 );
and \U$1741 ( \1880 , \1633 , \1745 );
or \U$1742 ( \1881 , \1878 , \1879 , \1880 );
xor \U$1743 ( \1882 , \1877 , \1881 );
and \U$1744 ( \1883 , \1746 , \1750 );
and \U$1745 ( \1884 , \1751 , \1754 );
or \U$1746 ( \1885 , \1883 , \1884 );
xor \U$1747 ( \1886 , \1882 , \1885 );
buf g5569_GF_PartitionCandidate( \1887_nG5569 , \1886 );
buf \U$1748 ( \1888 , \1887_nG5569 );
and \U$1749 ( \1889 , \1765 , \1769 );
and \U$1750 ( \1890 , \1769 , \1784 );
and \U$1751 ( \1891 , \1765 , \1784 );
or \U$1752 ( \1892 , \1889 , \1890 , \1891 );
and \U$1753 ( \1893 , \1800 , \1875 );
xor \U$1754 ( \1894 , \1892 , \1893 );
and \U$1755 ( \1895 , \1774 , \1778 );
and \U$1756 ( \1896 , \1778 , \1783 );
and \U$1757 ( \1897 , \1774 , \1783 );
or \U$1758 ( \1898 , \1895 , \1896 , \1897 );
and \U$1759 ( \1899 , \1819 , \1820 );
and \U$1760 ( \1900 , \1820 , \1828 );
and \U$1761 ( \1901 , \1819 , \1828 );
or \U$1762 ( \1902 , \1899 , \1900 , \1901 );
xor \U$1763 ( \1903 , \1898 , \1902 );
and \U$1764 ( \1904 , \1844 , \1858 );
and \U$1765 ( \1905 , \1858 , \1873 );
and \U$1766 ( \1906 , \1844 , \1873 );
or \U$1767 ( \1907 , \1904 , \1905 , \1906 );
xor \U$1768 ( \1908 , \1903 , \1907 );
xor \U$1769 ( \1909 , \1894 , \1908 );
and \U$1770 ( \1910 , \1790 , \1794 );
and \U$1771 ( \1911 , \1794 , \1799 );
and \U$1772 ( \1912 , \1790 , \1799 );
or \U$1773 ( \1913 , \1910 , \1911 , \1912 );
and \U$1774 ( \1914 , \1815 , \1829 );
and \U$1775 ( \1915 , \1829 , \1874 );
and \U$1776 ( \1916 , \1815 , \1874 );
or \U$1777 ( \1917 , \1914 , \1915 , \1916 );
xor \U$1778 ( \1918 , \1913 , \1917 );
and \U$1779 ( \1919 , \1834 , \1838 );
and \U$1780 ( \1920 , \1838 , \1843 );
and \U$1781 ( \1921 , \1834 , \1843 );
or \U$1782 ( \1922 , \1919 , \1920 , \1921 );
and \U$1783 ( \1923 , \1805 , \1809 );
and \U$1784 ( \1924 , \1809 , \1814 );
and \U$1785 ( \1925 , \1805 , \1814 );
or \U$1786 ( \1926 , \1923 , \1924 , \1925 );
xor \U$1787 ( \1927 , \1922 , \1926 );
and \U$1788 ( \1928 , \1863 , \1867 );
and \U$1789 ( \1929 , \1867 , \1872 );
and \U$1790 ( \1930 , \1863 , \1872 );
or \U$1791 ( \1931 , \1928 , \1929 , \1930 );
xor \U$1792 ( \1932 , \1927 , \1931 );
and \U$1793 ( \1933 , \261 , \141 );
and \U$1794 ( \1934 , \307 , \139 );
nor \U$1795 ( \1935 , \1933 , \1934 );
xnor \U$1796 ( \1936 , \1935 , \148 );
and \U$1797 ( \1937 , \178 , \156 );
and \U$1798 ( \1938 , \185 , \154 );
nor \U$1799 ( \1939 , \1937 , \1938 );
xnor \U$1800 ( \1940 , \1939 , \163 );
xor \U$1801 ( \1941 , \1936 , \1940 );
and \U$1802 ( \1942 , \189 , \296 );
and \U$1803 ( \1943 , \197 , \168 );
nor \U$1804 ( \1944 , \1942 , \1943 );
xnor \U$1805 ( \1945 , \1944 , \173 );
xor \U$1806 ( \1946 , \1941 , \1945 );
and \U$1807 ( \1947 , \1802 , \183 );
buf \U$1808 ( \1948 , RIb55e068_102);
and \U$1809 ( \1949 , \1948 , \180 );
nor \U$1810 ( \1950 , \1947 , \1949 );
xnor \U$1811 ( \1951 , \1950 , \179 );
and \U$1812 ( \1952 , \1601 , \195 );
and \U$1813 ( \1953 , \1684 , \193 );
nor \U$1814 ( \1954 , \1952 , \1953 );
xnor \U$1815 ( \1955 , \1954 , \202 );
xor \U$1816 ( \1956 , \1951 , \1955 );
buf \U$1817 ( \1957 , RIb55fee0_37);
buf \U$1818 ( \1958 , RIb55fe68_38);
and \U$1819 ( \1959 , \1958 , \1693 );
not \U$1820 ( \1960 , \1959 );
and \U$1821 ( \1961 , \1957 , \1960 );
xor \U$1822 ( \1962 , \1956 , \1961 );
xor \U$1823 ( \1963 , \1946 , \1962 );
and \U$1824 ( \1964 , \1333 , \215 );
and \U$1825 ( \1965 , \1484 , \213 );
nor \U$1826 ( \1966 , \1964 , \1965 );
xnor \U$1827 ( \1967 , \1966 , \222 );
and \U$1828 ( \1968 , \1147 , \230 );
and \U$1829 ( \1969 , \1192 , \228 );
nor \U$1830 ( \1970 , \1968 , \1969 );
xnor \U$1831 ( \1971 , \1970 , \237 );
xor \U$1832 ( \1972 , \1967 , \1971 );
and \U$1833 ( \1973 , \412 , \245 );
and \U$1834 ( \1974 , \474 , \243 );
nor \U$1835 ( \1975 , \1973 , \1974 );
xnor \U$1836 ( \1976 , \1975 , \252 );
xor \U$1837 ( \1977 , \1972 , \1976 );
xor \U$1838 ( \1978 , \1963 , \1977 );
xor \U$1839 ( \1979 , \1932 , \1978 );
and \U$1840 ( \1980 , \1848 , \1852 );
and \U$1841 ( \1981 , \1852 , \1857 );
and \U$1842 ( \1982 , \1848 , \1857 );
or \U$1843 ( \1983 , \1980 , \1981 , \1982 );
and \U$1844 ( \1984 , \209 , \438 );
and \U$1845 ( \1985 , \217 , \336 );
nor \U$1846 ( \1986 , \1984 , \1985 );
xnor \U$1847 ( \1987 , \1986 , \320 );
and \U$1848 ( \1988 , \224 , \1086 );
and \U$1849 ( \1989 , \232 , \508 );
nor \U$1850 ( \1990 , \1988 , \1989 );
xnor \U$1851 ( \1991 , \1990 , \487 );
xor \U$1852 ( \1992 , \1987 , \1991 );
and \U$1853 ( \1993 , \240 , \1301 );
and \U$1854 ( \1994 , \247 , \1246 );
nor \U$1855 ( \1995 , \1993 , \1994 );
xnor \U$1856 ( \1996 , \1995 , \1205 );
xor \U$1857 ( \1997 , \1992 , \1996 );
xor \U$1858 ( \1998 , \1983 , \1997 );
and \U$1859 ( \1999 , \134 , \1578 );
and \U$1860 ( \2000 , \143 , \1431 );
nor \U$1861 ( \2001 , \1999 , \2000 );
xnor \U$1862 ( \2002 , \2001 , \1436 );
and \U$1863 ( \2003 , \150 , \1824 );
and \U$1864 ( \2004 , \158 , \1739 );
nor \U$1865 ( \2005 , \2003 , \2004 );
xnor \U$1866 ( \2006 , \2005 , \1697 );
xor \U$1867 ( \2007 , \2002 , \2006 );
xor \U$1868 ( \2008 , \1958 , \1693 );
nand \U$1869 ( \2009 , \166 , \2008 );
xnor \U$1870 ( \2010 , \2009 , \1961 );
xor \U$1871 ( \2011 , \2007 , \2010 );
xor \U$1872 ( \2012 , \1998 , \2011 );
xor \U$1873 ( \2013 , \1979 , \2012 );
xor \U$1874 ( \2014 , \1918 , \2013 );
xor \U$1875 ( \2015 , \1909 , \2014 );
and \U$1876 ( \2016 , \1761 , \1785 );
and \U$1877 ( \2017 , \1785 , \1876 );
and \U$1878 ( \2018 , \1761 , \1876 );
or \U$1879 ( \2019 , \2016 , \2017 , \2018 );
xor \U$1880 ( \2020 , \2015 , \2019 );
and \U$1881 ( \2021 , \1877 , \1881 );
and \U$1882 ( \2022 , \1882 , \1885 );
or \U$1883 ( \2023 , \2021 , \2022 );
xor \U$1884 ( \2024 , \2020 , \2023 );
buf g5567_GF_PartitionCandidate( \2025_nG5567 , \2024 );
buf \U$1885 ( \2026 , \2025_nG5567 );
and \U$1886 ( \2027 , \1892 , \1893 );
and \U$1887 ( \2028 , \1893 , \1908 );
and \U$1888 ( \2029 , \1892 , \1908 );
or \U$1889 ( \2030 , \2027 , \2028 , \2029 );
and \U$1890 ( \2031 , \1913 , \1917 );
and \U$1891 ( \2032 , \1917 , \2013 );
and \U$1892 ( \2033 , \1913 , \2013 );
or \U$1893 ( \2034 , \2031 , \2032 , \2033 );
and \U$1894 ( \2035 , \1898 , \1902 );
and \U$1895 ( \2036 , \1902 , \1907 );
and \U$1896 ( \2037 , \1898 , \1907 );
or \U$1897 ( \2038 , \2035 , \2036 , \2037 );
and \U$1898 ( \2039 , \1932 , \1978 );
and \U$1899 ( \2040 , \1978 , \2012 );
and \U$1900 ( \2041 , \1932 , \2012 );
or \U$1901 ( \2042 , \2039 , \2040 , \2041 );
xor \U$1902 ( \2043 , \2038 , \2042 );
and \U$1903 ( \2044 , \1987 , \1991 );
and \U$1904 ( \2045 , \1991 , \1996 );
and \U$1905 ( \2046 , \1987 , \1996 );
or \U$1906 ( \2047 , \2044 , \2045 , \2046 );
and \U$1907 ( \2048 , \2002 , \2006 );
and \U$1908 ( \2049 , \2006 , \2010 );
and \U$1909 ( \2050 , \2002 , \2010 );
or \U$1910 ( \2051 , \2048 , \2049 , \2050 );
xor \U$1911 ( \2052 , \2047 , \2051 );
and \U$1912 ( \2053 , \158 , \1824 );
and \U$1913 ( \2054 , \134 , \1739 );
nor \U$1914 ( \2055 , \2053 , \2054 );
xnor \U$1915 ( \2056 , \2055 , \1697 );
xor \U$1916 ( \2057 , \2052 , \2056 );
xor \U$1917 ( \2058 , \2043 , \2057 );
xor \U$1918 ( \2059 , \2034 , \2058 );
and \U$1919 ( \2060 , \1936 , \1940 );
and \U$1920 ( \2061 , \1940 , \1945 );
and \U$1921 ( \2062 , \1936 , \1945 );
or \U$1922 ( \2063 , \2060 , \2061 , \2062 );
and \U$1923 ( \2064 , \1951 , \1955 );
and \U$1924 ( \2065 , \1955 , \1961 );
and \U$1925 ( \2066 , \1951 , \1961 );
or \U$1926 ( \2067 , \2064 , \2065 , \2066 );
xor \U$1927 ( \2068 , \2063 , \2067 );
and \U$1928 ( \2069 , \1967 , \1971 );
and \U$1929 ( \2070 , \1971 , \1976 );
and \U$1930 ( \2071 , \1967 , \1976 );
or \U$1931 ( \2072 , \2069 , \2070 , \2071 );
xor \U$1932 ( \2073 , \2068 , \2072 );
and \U$1933 ( \2074 , \1922 , \1926 );
and \U$1934 ( \2075 , \1926 , \1931 );
and \U$1935 ( \2076 , \1922 , \1931 );
or \U$1936 ( \2077 , \2074 , \2075 , \2076 );
and \U$1937 ( \2078 , \1946 , \1962 );
and \U$1938 ( \2079 , \1962 , \1977 );
and \U$1939 ( \2080 , \1946 , \1977 );
or \U$1940 ( \2081 , \2078 , \2079 , \2080 );
xor \U$1941 ( \2082 , \2077 , \2081 );
and \U$1942 ( \2083 , \1983 , \1997 );
and \U$1943 ( \2084 , \1997 , \2011 );
and \U$1944 ( \2085 , \1983 , \2011 );
or \U$1945 ( \2086 , \2083 , \2084 , \2085 );
xor \U$1946 ( \2087 , \2082 , \2086 );
xor \U$1947 ( \2088 , \2073 , \2087 );
and \U$1948 ( \2089 , \1948 , \183 );
buf \U$1949 ( \2090 , RIb55e0e0_101);
and \U$1950 ( \2091 , \2090 , \180 );
nor \U$1951 ( \2092 , \2089 , \2091 );
xnor \U$1952 ( \2093 , \2092 , \179 );
and \U$1953 ( \2094 , \1684 , \195 );
and \U$1954 ( \2095 , \1802 , \193 );
nor \U$1955 ( \2096 , \2094 , \2095 );
xnor \U$1956 ( \2097 , \2096 , \202 );
xor \U$1957 ( \2098 , \2093 , \2097 );
and \U$1958 ( \2099 , \1484 , \215 );
and \U$1959 ( \2100 , \1601 , \213 );
nor \U$1960 ( \2101 , \2099 , \2100 );
xnor \U$1961 ( \2102 , \2101 , \222 );
xor \U$1962 ( \2103 , \2098 , \2102 );
and \U$1963 ( \2104 , \1192 , \230 );
and \U$1964 ( \2105 , \1333 , \228 );
nor \U$1965 ( \2106 , \2104 , \2105 );
xnor \U$1966 ( \2107 , \2106 , \237 );
and \U$1967 ( \2108 , \474 , \245 );
and \U$1968 ( \2109 , \1147 , \243 );
nor \U$1969 ( \2110 , \2108 , \2109 );
xnor \U$1970 ( \2111 , \2110 , \252 );
xor \U$1971 ( \2112 , \2107 , \2111 );
and \U$1972 ( \2113 , \307 , \141 );
and \U$1973 ( \2114 , \412 , \139 );
nor \U$1974 ( \2115 , \2113 , \2114 );
xnor \U$1975 ( \2116 , \2115 , \148 );
xor \U$1976 ( \2117 , \2112 , \2116 );
xor \U$1977 ( \2118 , \2103 , \2117 );
xor \U$1978 ( \2119 , \1957 , \1958 );
not \U$1979 ( \2120 , \2008 );
and \U$1980 ( \2121 , \2119 , \2120 );
and \U$1981 ( \2122 , \166 , \2121 );
and \U$1982 ( \2123 , \150 , \2008 );
nor \U$1983 ( \2124 , \2122 , \2123 );
xnor \U$1984 ( \2125 , \2124 , \1961 );
and \U$1985 ( \2126 , \232 , \1086 );
and \U$1986 ( \2127 , \209 , \508 );
nor \U$1987 ( \2128 , \2126 , \2127 );
xnor \U$1988 ( \2129 , \2128 , \487 );
and \U$1989 ( \2130 , \247 , \1301 );
and \U$1990 ( \2131 , \224 , \1246 );
nor \U$1991 ( \2132 , \2130 , \2131 );
xnor \U$1992 ( \2133 , \2132 , \1205 );
xor \U$1993 ( \2134 , \2129 , \2133 );
and \U$1994 ( \2135 , \143 , \1578 );
and \U$1995 ( \2136 , \240 , \1431 );
nor \U$1996 ( \2137 , \2135 , \2136 );
xnor \U$1997 ( \2138 , \2137 , \1436 );
xor \U$1998 ( \2139 , \2134 , \2138 );
xor \U$1999 ( \2140 , \2125 , \2139 );
and \U$2000 ( \2141 , \185 , \156 );
and \U$2001 ( \2142 , \261 , \154 );
nor \U$2002 ( \2143 , \2141 , \2142 );
xnor \U$2003 ( \2144 , \2143 , \163 );
and \U$2004 ( \2145 , \197 , \296 );
and \U$2005 ( \2146 , \178 , \168 );
nor \U$2006 ( \2147 , \2145 , \2146 );
xnor \U$2007 ( \2148 , \2147 , \173 );
xor \U$2008 ( \2149 , \2144 , \2148 );
and \U$2009 ( \2150 , \217 , \438 );
and \U$2010 ( \2151 , \189 , \336 );
nor \U$2011 ( \2152 , \2150 , \2151 );
xnor \U$2012 ( \2153 , \2152 , \320 );
xor \U$2013 ( \2154 , \2149 , \2153 );
xor \U$2014 ( \2155 , \2140 , \2154 );
xor \U$2015 ( \2156 , \2118 , \2155 );
xor \U$2016 ( \2157 , \2088 , \2156 );
xor \U$2017 ( \2158 , \2059 , \2157 );
xor \U$2018 ( \2159 , \2030 , \2158 );
and \U$2019 ( \2160 , \1909 , \2014 );
xor \U$2020 ( \2161 , \2159 , \2160 );
and \U$2021 ( \2162 , \2015 , \2019 );
and \U$2022 ( \2163 , \2020 , \2023 );
or \U$2023 ( \2164 , \2162 , \2163 );
xor \U$2024 ( \2165 , \2161 , \2164 );
buf g5565_GF_PartitionCandidate( \2166_nG5565 , \2165 );
buf \U$2025 ( \2167 , \2166_nG5565 );
and \U$2026 ( \2168 , \2034 , \2058 );
and \U$2027 ( \2169 , \2058 , \2157 );
and \U$2028 ( \2170 , \2034 , \2157 );
or \U$2029 ( \2171 , \2168 , \2169 , \2170 );
and \U$2030 ( \2172 , \2038 , \2042 );
and \U$2031 ( \2173 , \2042 , \2057 );
and \U$2032 ( \2174 , \2038 , \2057 );
or \U$2033 ( \2175 , \2172 , \2173 , \2174 );
and \U$2034 ( \2176 , \2073 , \2087 );
and \U$2035 ( \2177 , \2087 , \2156 );
and \U$2036 ( \2178 , \2073 , \2156 );
or \U$2037 ( \2179 , \2176 , \2177 , \2178 );
xor \U$2038 ( \2180 , \2175 , \2179 );
and \U$2039 ( \2181 , \2090 , \183 );
buf \U$2040 ( \2182 , RIb55e158_100);
and \U$2041 ( \2183 , \2182 , \180 );
nor \U$2042 ( \2184 , \2181 , \2183 );
xnor \U$2043 ( \2185 , \2184 , \179 );
and \U$2044 ( \2186 , \1802 , \195 );
and \U$2045 ( \2187 , \1948 , \193 );
nor \U$2046 ( \2188 , \2186 , \2187 );
xnor \U$2047 ( \2189 , \2188 , \202 );
xor \U$2048 ( \2190 , \2185 , \2189 );
buf \U$2049 ( \2191 , RIb55ffd0_35);
buf \U$2050 ( \2192 , RIb55ff58_36);
and \U$2051 ( \2193 , \2192 , \1957 );
not \U$2052 ( \2194 , \2193 );
and \U$2053 ( \2195 , \2191 , \2194 );
xor \U$2054 ( \2196 , \2190 , \2195 );
and \U$2055 ( \2197 , \412 , \141 );
and \U$2056 ( \2198 , \474 , \139 );
nor \U$2057 ( \2199 , \2197 , \2198 );
xnor \U$2058 ( \2200 , \2199 , \148 );
and \U$2059 ( \2201 , \261 , \156 );
and \U$2060 ( \2202 , \307 , \154 );
nor \U$2061 ( \2203 , \2201 , \2202 );
xnor \U$2062 ( \2204 , \2203 , \163 );
xor \U$2063 ( \2205 , \2200 , \2204 );
and \U$2064 ( \2206 , \178 , \296 );
and \U$2065 ( \2207 , \185 , \168 );
nor \U$2066 ( \2208 , \2206 , \2207 );
xnor \U$2067 ( \2209 , \2208 , \173 );
xor \U$2068 ( \2210 , \2205 , \2209 );
and \U$2069 ( \2211 , \1601 , \215 );
and \U$2070 ( \2212 , \1684 , \213 );
nor \U$2071 ( \2213 , \2211 , \2212 );
xnor \U$2072 ( \2214 , \2213 , \222 );
and \U$2073 ( \2215 , \1333 , \230 );
and \U$2074 ( \2216 , \1484 , \228 );
nor \U$2075 ( \2217 , \2215 , \2216 );
xnor \U$2076 ( \2218 , \2217 , \237 );
xor \U$2077 ( \2219 , \2214 , \2218 );
and \U$2078 ( \2220 , \1147 , \245 );
and \U$2079 ( \2221 , \1192 , \243 );
nor \U$2080 ( \2222 , \2220 , \2221 );
xnor \U$2081 ( \2223 , \2222 , \252 );
xor \U$2082 ( \2224 , \2219 , \2223 );
xor \U$2083 ( \2225 , \2210 , \2224 );
and \U$2084 ( \2226 , \189 , \438 );
and \U$2085 ( \2227 , \197 , \336 );
nor \U$2086 ( \2228 , \2226 , \2227 );
xnor \U$2087 ( \2229 , \2228 , \320 );
and \U$2088 ( \2230 , \209 , \1086 );
and \U$2089 ( \2231 , \217 , \508 );
nor \U$2090 ( \2232 , \2230 , \2231 );
xnor \U$2091 ( \2233 , \2232 , \487 );
xor \U$2092 ( \2234 , \2229 , \2233 );
and \U$2093 ( \2235 , \224 , \1301 );
and \U$2094 ( \2236 , \232 , \1246 );
nor \U$2095 ( \2237 , \2235 , \2236 );
xnor \U$2096 ( \2238 , \2237 , \1205 );
xor \U$2097 ( \2239 , \2234 , \2238 );
xor \U$2098 ( \2240 , \2225 , \2239 );
xor \U$2099 ( \2241 , \2196 , \2240 );
and \U$2100 ( \2242 , \2129 , \2133 );
and \U$2101 ( \2243 , \2133 , \2138 );
and \U$2102 ( \2244 , \2129 , \2138 );
or \U$2103 ( \2245 , \2242 , \2243 , \2244 );
xor \U$2104 ( \2246 , \2192 , \1957 );
nand \U$2105 ( \2247 , \166 , \2246 );
xnor \U$2106 ( \2248 , \2247 , \2195 );
xor \U$2107 ( \2249 , \2245 , \2248 );
and \U$2108 ( \2250 , \240 , \1578 );
and \U$2109 ( \2251 , \247 , \1431 );
nor \U$2110 ( \2252 , \2250 , \2251 );
xnor \U$2111 ( \2253 , \2252 , \1436 );
and \U$2112 ( \2254 , \134 , \1824 );
and \U$2113 ( \2255 , \143 , \1739 );
nor \U$2114 ( \2256 , \2254 , \2255 );
xnor \U$2115 ( \2257 , \2256 , \1697 );
xor \U$2116 ( \2258 , \2253 , \2257 );
and \U$2117 ( \2259 , \150 , \2121 );
and \U$2118 ( \2260 , \158 , \2008 );
nor \U$2119 ( \2261 , \2259 , \2260 );
xnor \U$2120 ( \2262 , \2261 , \1961 );
xor \U$2121 ( \2263 , \2258 , \2262 );
xor \U$2122 ( \2264 , \2249 , \2263 );
xor \U$2123 ( \2265 , \2241 , \2264 );
xor \U$2124 ( \2266 , \2180 , \2265 );
xor \U$2125 ( \2267 , \2171 , \2266 );
and \U$2126 ( \2268 , \2047 , \2051 );
and \U$2127 ( \2269 , \2051 , \2056 );
and \U$2128 ( \2270 , \2047 , \2056 );
or \U$2129 ( \2271 , \2268 , \2269 , \2270 );
and \U$2130 ( \2272 , \2063 , \2067 );
and \U$2131 ( \2273 , \2067 , \2072 );
and \U$2132 ( \2274 , \2063 , \2072 );
or \U$2133 ( \2275 , \2272 , \2273 , \2274 );
xor \U$2134 ( \2276 , \2271 , \2275 );
and \U$2135 ( \2277 , \2125 , \2139 );
and \U$2136 ( \2278 , \2139 , \2154 );
and \U$2137 ( \2279 , \2125 , \2154 );
or \U$2138 ( \2280 , \2277 , \2278 , \2279 );
xor \U$2139 ( \2281 , \2276 , \2280 );
and \U$2140 ( \2282 , \2077 , \2081 );
and \U$2141 ( \2283 , \2081 , \2086 );
and \U$2142 ( \2284 , \2077 , \2086 );
or \U$2143 ( \2285 , \2282 , \2283 , \2284 );
and \U$2144 ( \2286 , \2103 , \2117 );
and \U$2145 ( \2287 , \2117 , \2155 );
and \U$2146 ( \2288 , \2103 , \2155 );
or \U$2147 ( \2289 , \2286 , \2287 , \2288 );
xor \U$2148 ( \2290 , \2285 , \2289 );
and \U$2149 ( \2291 , \2093 , \2097 );
and \U$2150 ( \2292 , \2097 , \2102 );
and \U$2151 ( \2293 , \2093 , \2102 );
or \U$2152 ( \2294 , \2291 , \2292 , \2293 );
and \U$2153 ( \2295 , \2144 , \2148 );
and \U$2154 ( \2296 , \2148 , \2153 );
and \U$2155 ( \2297 , \2144 , \2153 );
or \U$2156 ( \2298 , \2295 , \2296 , \2297 );
xor \U$2157 ( \2299 , \2294 , \2298 );
and \U$2158 ( \2300 , \2107 , \2111 );
and \U$2159 ( \2301 , \2111 , \2116 );
and \U$2160 ( \2302 , \2107 , \2116 );
or \U$2161 ( \2303 , \2300 , \2301 , \2302 );
xor \U$2162 ( \2304 , \2299 , \2303 );
xor \U$2163 ( \2305 , \2290 , \2304 );
xor \U$2164 ( \2306 , \2281 , \2305 );
xor \U$2165 ( \2307 , \2267 , \2306 );
and \U$2166 ( \2308 , \2030 , \2158 );
xor \U$2167 ( \2309 , \2307 , \2308 );
and \U$2168 ( \2310 , \2159 , \2160 );
and \U$2169 ( \2311 , \2161 , \2164 );
or \U$2170 ( \2312 , \2310 , \2311 );
xor \U$2171 ( \2313 , \2309 , \2312 );
buf g5563_GF_PartitionCandidate( \2314_nG5563 , \2313 );
buf \U$2172 ( \2315 , \2314_nG5563 );
and \U$2173 ( \2316 , \2175 , \2179 );
and \U$2174 ( \2317 , \2179 , \2265 );
and \U$2175 ( \2318 , \2175 , \2265 );
or \U$2176 ( \2319 , \2316 , \2317 , \2318 );
and \U$2177 ( \2320 , \2281 , \2305 );
xor \U$2178 ( \2321 , \2319 , \2320 );
and \U$2179 ( \2322 , \2285 , \2289 );
and \U$2180 ( \2323 , \2289 , \2304 );
and \U$2181 ( \2324 , \2285 , \2304 );
or \U$2182 ( \2325 , \2322 , \2323 , \2324 );
and \U$2183 ( \2326 , \2271 , \2275 );
and \U$2184 ( \2327 , \2275 , \2280 );
and \U$2185 ( \2328 , \2271 , \2280 );
or \U$2186 ( \2329 , \2326 , \2327 , \2328 );
and \U$2187 ( \2330 , \2196 , \2240 );
and \U$2188 ( \2331 , \2240 , \2264 );
and \U$2189 ( \2332 , \2196 , \2264 );
or \U$2190 ( \2333 , \2330 , \2331 , \2332 );
xor \U$2191 ( \2334 , \2329 , \2333 );
and \U$2192 ( \2335 , \2200 , \2204 );
and \U$2193 ( \2336 , \2204 , \2209 );
and \U$2194 ( \2337 , \2200 , \2209 );
or \U$2195 ( \2338 , \2335 , \2336 , \2337 );
and \U$2196 ( \2339 , \2214 , \2218 );
and \U$2197 ( \2340 , \2218 , \2223 );
and \U$2198 ( \2341 , \2214 , \2223 );
or \U$2199 ( \2342 , \2339 , \2340 , \2341 );
xor \U$2200 ( \2343 , \2338 , \2342 );
and \U$2201 ( \2344 , \2185 , \2189 );
and \U$2202 ( \2345 , \2189 , \2195 );
and \U$2203 ( \2346 , \2185 , \2195 );
or \U$2204 ( \2347 , \2344 , \2345 , \2346 );
xor \U$2205 ( \2348 , \2343 , \2347 );
xor \U$2206 ( \2349 , \2334 , \2348 );
xor \U$2207 ( \2350 , \2325 , \2349 );
and \U$2208 ( \2351 , \2294 , \2298 );
and \U$2209 ( \2352 , \2298 , \2303 );
and \U$2210 ( \2353 , \2294 , \2303 );
or \U$2211 ( \2354 , \2351 , \2352 , \2353 );
and \U$2212 ( \2355 , \2210 , \2224 );
and \U$2213 ( \2356 , \2224 , \2239 );
and \U$2214 ( \2357 , \2210 , \2239 );
or \U$2215 ( \2358 , \2355 , \2356 , \2357 );
xor \U$2216 ( \2359 , \2354 , \2358 );
and \U$2217 ( \2360 , \2245 , \2248 );
and \U$2218 ( \2361 , \2248 , \2263 );
and \U$2219 ( \2362 , \2245 , \2263 );
or \U$2220 ( \2363 , \2360 , \2361 , \2362 );
xor \U$2221 ( \2364 , \2359 , \2363 );
and \U$2222 ( \2365 , \2182 , \183 );
buf \U$2223 ( \2366 , RIb55e1d0_99);
and \U$2224 ( \2367 , \2366 , \180 );
nor \U$2225 ( \2368 , \2365 , \2367 );
xnor \U$2226 ( \2369 , \2368 , \179 );
and \U$2227 ( \2370 , \1948 , \195 );
and \U$2228 ( \2371 , \2090 , \193 );
nor \U$2229 ( \2372 , \2370 , \2371 );
xnor \U$2230 ( \2373 , \2372 , \202 );
xor \U$2231 ( \2374 , \2369 , \2373 );
and \U$2232 ( \2375 , \1684 , \215 );
and \U$2233 ( \2376 , \1802 , \213 );
nor \U$2234 ( \2377 , \2375 , \2376 );
xnor \U$2235 ( \2378 , \2377 , \222 );
xor \U$2236 ( \2379 , \2374 , \2378 );
and \U$2237 ( \2380 , \2229 , \2233 );
and \U$2238 ( \2381 , \2233 , \2238 );
and \U$2239 ( \2382 , \2229 , \2238 );
or \U$2240 ( \2383 , \2380 , \2381 , \2382 );
and \U$2241 ( \2384 , \2253 , \2257 );
and \U$2242 ( \2385 , \2257 , \2262 );
and \U$2243 ( \2386 , \2253 , \2262 );
or \U$2244 ( \2387 , \2384 , \2385 , \2386 );
xor \U$2245 ( \2388 , \2383 , \2387 );
and \U$2246 ( \2389 , \143 , \1824 );
and \U$2247 ( \2390 , \240 , \1739 );
nor \U$2248 ( \2391 , \2389 , \2390 );
xnor \U$2249 ( \2392 , \2391 , \1697 );
and \U$2250 ( \2393 , \158 , \2121 );
and \U$2251 ( \2394 , \134 , \2008 );
nor \U$2252 ( \2395 , \2393 , \2394 );
xnor \U$2253 ( \2396 , \2395 , \1961 );
xor \U$2254 ( \2397 , \2392 , \2396 );
xor \U$2255 ( \2398 , \2191 , \2192 );
not \U$2256 ( \2399 , \2246 );
and \U$2257 ( \2400 , \2398 , \2399 );
and \U$2258 ( \2401 , \166 , \2400 );
and \U$2259 ( \2402 , \150 , \2246 );
nor \U$2260 ( \2403 , \2401 , \2402 );
xnor \U$2261 ( \2404 , \2403 , \2195 );
xor \U$2262 ( \2405 , \2397 , \2404 );
xor \U$2263 ( \2406 , \2388 , \2405 );
xor \U$2264 ( \2407 , \2379 , \2406 );
and \U$2265 ( \2408 , \307 , \156 );
and \U$2266 ( \2409 , \412 , \154 );
nor \U$2267 ( \2410 , \2408 , \2409 );
xnor \U$2268 ( \2411 , \2410 , \163 );
and \U$2269 ( \2412 , \185 , \296 );
and \U$2270 ( \2413 , \261 , \168 );
nor \U$2271 ( \2414 , \2412 , \2413 );
xnor \U$2272 ( \2415 , \2414 , \173 );
xor \U$2273 ( \2416 , \2411 , \2415 );
and \U$2274 ( \2417 , \197 , \438 );
and \U$2275 ( \2418 , \178 , \336 );
nor \U$2276 ( \2419 , \2417 , \2418 );
xnor \U$2277 ( \2420 , \2419 , \320 );
xor \U$2278 ( \2421 , \2416 , \2420 );
and \U$2279 ( \2422 , \1484 , \230 );
and \U$2280 ( \2423 , \1601 , \228 );
nor \U$2281 ( \2424 , \2422 , \2423 );
xnor \U$2282 ( \2425 , \2424 , \237 );
and \U$2283 ( \2426 , \1192 , \245 );
and \U$2284 ( \2427 , \1333 , \243 );
nor \U$2285 ( \2428 , \2426 , \2427 );
xnor \U$2286 ( \2429 , \2428 , \252 );
xor \U$2287 ( \2430 , \2425 , \2429 );
and \U$2288 ( \2431 , \474 , \141 );
and \U$2289 ( \2432 , \1147 , \139 );
nor \U$2290 ( \2433 , \2431 , \2432 );
xnor \U$2291 ( \2434 , \2433 , \148 );
xor \U$2292 ( \2435 , \2430 , \2434 );
xor \U$2293 ( \2436 , \2421 , \2435 );
and \U$2294 ( \2437 , \217 , \1086 );
and \U$2295 ( \2438 , \189 , \508 );
nor \U$2296 ( \2439 , \2437 , \2438 );
xnor \U$2297 ( \2440 , \2439 , \487 );
and \U$2298 ( \2441 , \232 , \1301 );
and \U$2299 ( \2442 , \209 , \1246 );
nor \U$2300 ( \2443 , \2441 , \2442 );
xnor \U$2301 ( \2444 , \2443 , \1205 );
xor \U$2302 ( \2445 , \2440 , \2444 );
and \U$2303 ( \2446 , \247 , \1578 );
and \U$2304 ( \2447 , \224 , \1431 );
nor \U$2305 ( \2448 , \2446 , \2447 );
xnor \U$2306 ( \2449 , \2448 , \1436 );
xor \U$2307 ( \2450 , \2445 , \2449 );
xor \U$2308 ( \2451 , \2436 , \2450 );
xor \U$2309 ( \2452 , \2407 , \2451 );
xor \U$2310 ( \2453 , \2364 , \2452 );
xor \U$2311 ( \2454 , \2350 , \2453 );
xor \U$2312 ( \2455 , \2321 , \2454 );
and \U$2313 ( \2456 , \2171 , \2266 );
and \U$2314 ( \2457 , \2266 , \2306 );
and \U$2315 ( \2458 , \2171 , \2306 );
or \U$2316 ( \2459 , \2456 , \2457 , \2458 );
xor \U$2317 ( \2460 , \2455 , \2459 );
and \U$2318 ( \2461 , \2307 , \2308 );
and \U$2319 ( \2462 , \2309 , \2312 );
or \U$2320 ( \2463 , \2461 , \2462 );
xor \U$2321 ( \2464 , \2460 , \2463 );
buf g5561_GF_PartitionCandidate( \2465_nG5561 , \2464 );
buf \U$2322 ( \2466 , \2465_nG5561 );
and \U$2323 ( \2467 , \2325 , \2349 );
and \U$2324 ( \2468 , \2349 , \2453 );
and \U$2325 ( \2469 , \2325 , \2453 );
or \U$2326 ( \2470 , \2467 , \2468 , \2469 );
and \U$2327 ( \2471 , \2329 , \2333 );
and \U$2328 ( \2472 , \2333 , \2348 );
and \U$2329 ( \2473 , \2329 , \2348 );
or \U$2330 ( \2474 , \2471 , \2472 , \2473 );
and \U$2331 ( \2475 , \2364 , \2452 );
xor \U$2332 ( \2476 , \2474 , \2475 );
and \U$2333 ( \2477 , \2392 , \2396 );
and \U$2334 ( \2478 , \2396 , \2404 );
and \U$2335 ( \2479 , \2392 , \2404 );
or \U$2336 ( \2480 , \2477 , \2478 , \2479 );
and \U$2337 ( \2481 , \2440 , \2444 );
and \U$2338 ( \2482 , \2444 , \2449 );
and \U$2339 ( \2483 , \2440 , \2449 );
or \U$2340 ( \2484 , \2481 , \2482 , \2483 );
xor \U$2341 ( \2485 , \2480 , \2484 );
and \U$2342 ( \2486 , \150 , \2400 );
and \U$2343 ( \2487 , \158 , \2246 );
nor \U$2344 ( \2488 , \2486 , \2487 );
xnor \U$2345 ( \2489 , \2488 , \2195 );
xor \U$2346 ( \2490 , \2485 , \2489 );
and \U$2347 ( \2491 , \1802 , \215 );
and \U$2348 ( \2492 , \1948 , \213 );
nor \U$2349 ( \2493 , \2491 , \2492 );
xnor \U$2350 ( \2494 , \2493 , \222 );
and \U$2351 ( \2495 , \1601 , \230 );
and \U$2352 ( \2496 , \1684 , \228 );
nor \U$2353 ( \2497 , \2495 , \2496 );
xnor \U$2354 ( \2498 , \2497 , \237 );
xor \U$2355 ( \2499 , \2494 , \2498 );
and \U$2356 ( \2500 , \1333 , \245 );
and \U$2357 ( \2501 , \1484 , \243 );
nor \U$2358 ( \2502 , \2500 , \2501 );
xnor \U$2359 ( \2503 , \2502 , \252 );
xor \U$2360 ( \2504 , \2499 , \2503 );
and \U$2361 ( \2505 , \1147 , \141 );
and \U$2362 ( \2506 , \1192 , \139 );
nor \U$2363 ( \2507 , \2505 , \2506 );
xnor \U$2364 ( \2508 , \2507 , \148 );
and \U$2365 ( \2509 , \412 , \156 );
and \U$2366 ( \2510 , \474 , \154 );
nor \U$2367 ( \2511 , \2509 , \2510 );
xnor \U$2368 ( \2512 , \2511 , \163 );
xor \U$2369 ( \2513 , \2508 , \2512 );
and \U$2370 ( \2514 , \261 , \296 );
and \U$2371 ( \2515 , \307 , \168 );
nor \U$2372 ( \2516 , \2514 , \2515 );
xnor \U$2373 ( \2517 , \2516 , \173 );
xor \U$2374 ( \2518 , \2513 , \2517 );
xor \U$2375 ( \2519 , \2504 , \2518 );
and \U$2376 ( \2520 , \2366 , \183 );
buf \U$2377 ( \2521 , RIb55e248_98);
and \U$2378 ( \2522 , \2521 , \180 );
nor \U$2379 ( \2523 , \2520 , \2522 );
xnor \U$2380 ( \2524 , \2523 , \179 );
and \U$2381 ( \2525 , \2090 , \195 );
and \U$2382 ( \2526 , \2182 , \193 );
nor \U$2383 ( \2527 , \2525 , \2526 );
xnor \U$2384 ( \2528 , \2527 , \202 );
xor \U$2385 ( \2529 , \2524 , \2528 );
buf \U$2386 ( \2530 , RIb5600c0_33);
buf \U$2387 ( \2531 , RIb560048_34);
and \U$2388 ( \2532 , \2531 , \2191 );
not \U$2389 ( \2533 , \2532 );
and \U$2390 ( \2534 , \2530 , \2533 );
xor \U$2391 ( \2535 , \2529 , \2534 );
xor \U$2392 ( \2536 , \2519 , \2535 );
xor \U$2393 ( \2537 , \2490 , \2536 );
xor \U$2394 ( \2538 , \2531 , \2191 );
nand \U$2395 ( \2539 , \166 , \2538 );
xnor \U$2396 ( \2540 , \2539 , \2534 );
and \U$2397 ( \2541 , \224 , \1578 );
and \U$2398 ( \2542 , \232 , \1431 );
nor \U$2399 ( \2543 , \2541 , \2542 );
xnor \U$2400 ( \2544 , \2543 , \1436 );
and \U$2401 ( \2545 , \240 , \1824 );
and \U$2402 ( \2546 , \247 , \1739 );
nor \U$2403 ( \2547 , \2545 , \2546 );
xnor \U$2404 ( \2548 , \2547 , \1697 );
xor \U$2405 ( \2549 , \2544 , \2548 );
and \U$2406 ( \2550 , \134 , \2121 );
and \U$2407 ( \2551 , \143 , \2008 );
nor \U$2408 ( \2552 , \2550 , \2551 );
xnor \U$2409 ( \2553 , \2552 , \1961 );
xor \U$2410 ( \2554 , \2549 , \2553 );
xor \U$2411 ( \2555 , \2540 , \2554 );
and \U$2412 ( \2556 , \178 , \438 );
and \U$2413 ( \2557 , \185 , \336 );
nor \U$2414 ( \2558 , \2556 , \2557 );
xnor \U$2415 ( \2559 , \2558 , \320 );
and \U$2416 ( \2560 , \189 , \1086 );
and \U$2417 ( \2561 , \197 , \508 );
nor \U$2418 ( \2562 , \2560 , \2561 );
xnor \U$2419 ( \2563 , \2562 , \487 );
xor \U$2420 ( \2564 , \2559 , \2563 );
and \U$2421 ( \2565 , \209 , \1301 );
and \U$2422 ( \2566 , \217 , \1246 );
nor \U$2423 ( \2567 , \2565 , \2566 );
xnor \U$2424 ( \2568 , \2567 , \1205 );
xor \U$2425 ( \2569 , \2564 , \2568 );
xor \U$2426 ( \2570 , \2555 , \2569 );
xor \U$2427 ( \2571 , \2537 , \2570 );
xor \U$2428 ( \2572 , \2476 , \2571 );
xor \U$2429 ( \2573 , \2470 , \2572 );
and \U$2430 ( \2574 , \2338 , \2342 );
and \U$2431 ( \2575 , \2342 , \2347 );
and \U$2432 ( \2576 , \2338 , \2347 );
or \U$2433 ( \2577 , \2574 , \2575 , \2576 );
and \U$2434 ( \2578 , \2383 , \2387 );
and \U$2435 ( \2579 , \2387 , \2405 );
and \U$2436 ( \2580 , \2383 , \2405 );
or \U$2437 ( \2581 , \2578 , \2579 , \2580 );
xor \U$2438 ( \2582 , \2577 , \2581 );
and \U$2439 ( \2583 , \2421 , \2435 );
and \U$2440 ( \2584 , \2435 , \2450 );
and \U$2441 ( \2585 , \2421 , \2450 );
or \U$2442 ( \2586 , \2583 , \2584 , \2585 );
xor \U$2443 ( \2587 , \2582 , \2586 );
and \U$2444 ( \2588 , \2354 , \2358 );
and \U$2445 ( \2589 , \2358 , \2363 );
and \U$2446 ( \2590 , \2354 , \2363 );
or \U$2447 ( \2591 , \2588 , \2589 , \2590 );
and \U$2448 ( \2592 , \2379 , \2406 );
and \U$2449 ( \2593 , \2406 , \2451 );
and \U$2450 ( \2594 , \2379 , \2451 );
or \U$2451 ( \2595 , \2592 , \2593 , \2594 );
xor \U$2452 ( \2596 , \2591 , \2595 );
and \U$2453 ( \2597 , \2411 , \2415 );
and \U$2454 ( \2598 , \2415 , \2420 );
and \U$2455 ( \2599 , \2411 , \2420 );
or \U$2456 ( \2600 , \2597 , \2598 , \2599 );
and \U$2457 ( \2601 , \2425 , \2429 );
and \U$2458 ( \2602 , \2429 , \2434 );
and \U$2459 ( \2603 , \2425 , \2434 );
or \U$2460 ( \2604 , \2601 , \2602 , \2603 );
xor \U$2461 ( \2605 , \2600 , \2604 );
and \U$2462 ( \2606 , \2369 , \2373 );
and \U$2463 ( \2607 , \2373 , \2378 );
and \U$2464 ( \2608 , \2369 , \2378 );
or \U$2465 ( \2609 , \2606 , \2607 , \2608 );
xor \U$2466 ( \2610 , \2605 , \2609 );
xor \U$2467 ( \2611 , \2596 , \2610 );
xor \U$2468 ( \2612 , \2587 , \2611 );
xor \U$2469 ( \2613 , \2573 , \2612 );
and \U$2470 ( \2614 , \2319 , \2320 );
and \U$2471 ( \2615 , \2320 , \2454 );
and \U$2472 ( \2616 , \2319 , \2454 );
or \U$2473 ( \2617 , \2614 , \2615 , \2616 );
xor \U$2474 ( \2618 , \2613 , \2617 );
and \U$2475 ( \2619 , \2455 , \2459 );
and \U$2476 ( \2620 , \2460 , \2463 );
or \U$2477 ( \2621 , \2619 , \2620 );
xor \U$2478 ( \2622 , \2618 , \2621 );
buf g555f_GF_PartitionCandidate( \2623_nG555f , \2622 );
buf \U$2479 ( \2624 , \2623_nG555f );
and \U$2480 ( \2625 , \2474 , \2475 );
and \U$2481 ( \2626 , \2475 , \2571 );
and \U$2482 ( \2627 , \2474 , \2571 );
or \U$2483 ( \2628 , \2625 , \2626 , \2627 );
and \U$2484 ( \2629 , \2587 , \2611 );
xor \U$2485 ( \2630 , \2628 , \2629 );
and \U$2486 ( \2631 , \2591 , \2595 );
and \U$2487 ( \2632 , \2595 , \2610 );
and \U$2488 ( \2633 , \2591 , \2610 );
or \U$2489 ( \2634 , \2631 , \2632 , \2633 );
and \U$2490 ( \2635 , \2577 , \2581 );
and \U$2491 ( \2636 , \2581 , \2586 );
and \U$2492 ( \2637 , \2577 , \2586 );
or \U$2493 ( \2638 , \2635 , \2636 , \2637 );
and \U$2494 ( \2639 , \2490 , \2536 );
and \U$2495 ( \2640 , \2536 , \2570 );
and \U$2496 ( \2641 , \2490 , \2570 );
or \U$2497 ( \2642 , \2639 , \2640 , \2641 );
xor \U$2498 ( \2643 , \2638 , \2642 );
and \U$2499 ( \2644 , \2494 , \2498 );
and \U$2500 ( \2645 , \2498 , \2503 );
and \U$2501 ( \2646 , \2494 , \2503 );
or \U$2502 ( \2647 , \2644 , \2645 , \2646 );
and \U$2503 ( \2648 , \2508 , \2512 );
and \U$2504 ( \2649 , \2512 , \2517 );
and \U$2505 ( \2650 , \2508 , \2517 );
or \U$2506 ( \2651 , \2648 , \2649 , \2650 );
xor \U$2507 ( \2652 , \2647 , \2651 );
and \U$2508 ( \2653 , \2524 , \2528 );
and \U$2509 ( \2654 , \2528 , \2534 );
and \U$2510 ( \2655 , \2524 , \2534 );
or \U$2511 ( \2656 , \2653 , \2654 , \2655 );
xor \U$2512 ( \2657 , \2652 , \2656 );
and \U$2513 ( \2658 , \2544 , \2548 );
and \U$2514 ( \2659 , \2548 , \2553 );
and \U$2515 ( \2660 , \2544 , \2553 );
or \U$2516 ( \2661 , \2658 , \2659 , \2660 );
and \U$2517 ( \2662 , \2559 , \2563 );
and \U$2518 ( \2663 , \2563 , \2568 );
and \U$2519 ( \2664 , \2559 , \2568 );
or \U$2520 ( \2665 , \2662 , \2663 , \2664 );
xor \U$2521 ( \2666 , \2661 , \2665 );
xor \U$2522 ( \2667 , \2530 , \2531 );
not \U$2523 ( \2668 , \2538 );
and \U$2524 ( \2669 , \2667 , \2668 );
and \U$2525 ( \2670 , \166 , \2669 );
and \U$2526 ( \2671 , \150 , \2538 );
nor \U$2527 ( \2672 , \2670 , \2671 );
xnor \U$2528 ( \2673 , \2672 , \2534 );
xor \U$2529 ( \2674 , \2666 , \2673 );
xor \U$2530 ( \2675 , \2657 , \2674 );
and \U$2531 ( \2676 , \197 , \1086 );
and \U$2532 ( \2677 , \178 , \508 );
nor \U$2533 ( \2678 , \2676 , \2677 );
xnor \U$2534 ( \2679 , \2678 , \487 );
and \U$2535 ( \2680 , \217 , \1301 );
and \U$2536 ( \2681 , \189 , \1246 );
nor \U$2537 ( \2682 , \2680 , \2681 );
xnor \U$2538 ( \2683 , \2682 , \1205 );
xor \U$2539 ( \2684 , \2679 , \2683 );
and \U$2540 ( \2685 , \232 , \1578 );
and \U$2541 ( \2686 , \209 , \1431 );
nor \U$2542 ( \2687 , \2685 , \2686 );
xnor \U$2543 ( \2688 , \2687 , \1436 );
xor \U$2544 ( \2689 , \2684 , \2688 );
and \U$2545 ( \2690 , \247 , \1824 );
and \U$2546 ( \2691 , \224 , \1739 );
nor \U$2547 ( \2692 , \2690 , \2691 );
xnor \U$2548 ( \2693 , \2692 , \1697 );
and \U$2549 ( \2694 , \143 , \2121 );
and \U$2550 ( \2695 , \240 , \2008 );
nor \U$2551 ( \2696 , \2694 , \2695 );
xnor \U$2552 ( \2697 , \2696 , \1961 );
xor \U$2553 ( \2698 , \2693 , \2697 );
and \U$2554 ( \2699 , \158 , \2400 );
and \U$2555 ( \2700 , \134 , \2246 );
nor \U$2556 ( \2701 , \2699 , \2700 );
xnor \U$2557 ( \2702 , \2701 , \2195 );
xor \U$2558 ( \2703 , \2698 , \2702 );
xor \U$2559 ( \2704 , \2689 , \2703 );
and \U$2560 ( \2705 , \474 , \156 );
and \U$2561 ( \2706 , \1147 , \154 );
nor \U$2562 ( \2707 , \2705 , \2706 );
xnor \U$2563 ( \2708 , \2707 , \163 );
and \U$2564 ( \2709 , \307 , \296 );
and \U$2565 ( \2710 , \412 , \168 );
nor \U$2566 ( \2711 , \2709 , \2710 );
xnor \U$2567 ( \2712 , \2711 , \173 );
xor \U$2568 ( \2713 , \2708 , \2712 );
and \U$2569 ( \2714 , \185 , \438 );
and \U$2570 ( \2715 , \261 , \336 );
nor \U$2571 ( \2716 , \2714 , \2715 );
xnor \U$2572 ( \2717 , \2716 , \320 );
xor \U$2573 ( \2718 , \2713 , \2717 );
xor \U$2574 ( \2719 , \2704 , \2718 );
xor \U$2575 ( \2720 , \2675 , \2719 );
xor \U$2576 ( \2721 , \2643 , \2720 );
xor \U$2577 ( \2722 , \2634 , \2721 );
and \U$2578 ( \2723 , \2600 , \2604 );
and \U$2579 ( \2724 , \2604 , \2609 );
and \U$2580 ( \2725 , \2600 , \2609 );
or \U$2581 ( \2726 , \2723 , \2724 , \2725 );
and \U$2582 ( \2727 , \2480 , \2484 );
and \U$2583 ( \2728 , \2484 , \2489 );
and \U$2584 ( \2729 , \2480 , \2489 );
or \U$2585 ( \2730 , \2727 , \2728 , \2729 );
xor \U$2586 ( \2731 , \2726 , \2730 );
and \U$2587 ( \2732 , \2540 , \2554 );
and \U$2588 ( \2733 , \2554 , \2569 );
and \U$2589 ( \2734 , \2540 , \2569 );
or \U$2590 ( \2735 , \2732 , \2733 , \2734 );
xor \U$2591 ( \2736 , \2731 , \2735 );
and \U$2592 ( \2737 , \2504 , \2518 );
and \U$2593 ( \2738 , \2518 , \2535 );
and \U$2594 ( \2739 , \2504 , \2535 );
or \U$2595 ( \2740 , \2737 , \2738 , \2739 );
and \U$2596 ( \2741 , \1684 , \230 );
and \U$2597 ( \2742 , \1802 , \228 );
nor \U$2598 ( \2743 , \2741 , \2742 );
xnor \U$2599 ( \2744 , \2743 , \237 );
and \U$2600 ( \2745 , \1484 , \245 );
and \U$2601 ( \2746 , \1601 , \243 );
nor \U$2602 ( \2747 , \2745 , \2746 );
xnor \U$2603 ( \2748 , \2747 , \252 );
xor \U$2604 ( \2749 , \2744 , \2748 );
and \U$2605 ( \2750 , \1192 , \141 );
and \U$2606 ( \2751 , \1333 , \139 );
nor \U$2607 ( \2752 , \2750 , \2751 );
xnor \U$2608 ( \2753 , \2752 , \148 );
xor \U$2609 ( \2754 , \2749 , \2753 );
xor \U$2610 ( \2755 , \2740 , \2754 );
and \U$2611 ( \2756 , \2521 , \183 );
buf \U$2612 ( \2757 , RIb55e2c0_97);
and \U$2613 ( \2758 , \2757 , \180 );
nor \U$2614 ( \2759 , \2756 , \2758 );
xnor \U$2615 ( \2760 , \2759 , \179 );
and \U$2616 ( \2761 , \2182 , \195 );
and \U$2617 ( \2762 , \2366 , \193 );
nor \U$2618 ( \2763 , \2761 , \2762 );
xnor \U$2619 ( \2764 , \2763 , \202 );
xor \U$2620 ( \2765 , \2760 , \2764 );
and \U$2621 ( \2766 , \1948 , \215 );
and \U$2622 ( \2767 , \2090 , \213 );
nor \U$2623 ( \2768 , \2766 , \2767 );
xnor \U$2624 ( \2769 , \2768 , \222 );
xor \U$2625 ( \2770 , \2765 , \2769 );
xor \U$2626 ( \2771 , \2755 , \2770 );
xor \U$2627 ( \2772 , \2736 , \2771 );
xor \U$2628 ( \2773 , \2722 , \2772 );
xor \U$2629 ( \2774 , \2630 , \2773 );
and \U$2630 ( \2775 , \2470 , \2572 );
and \U$2631 ( \2776 , \2572 , \2612 );
and \U$2632 ( \2777 , \2470 , \2612 );
or \U$2633 ( \2778 , \2775 , \2776 , \2777 );
xor \U$2634 ( \2779 , \2774 , \2778 );
and \U$2635 ( \2780 , \2613 , \2617 );
and \U$2636 ( \2781 , \2618 , \2621 );
or \U$2637 ( \2782 , \2780 , \2781 );
xor \U$2638 ( \2783 , \2779 , \2782 );
buf g555d_GF_PartitionCandidate( \2784_nG555d , \2783 );
buf \U$2639 ( \2785 , \2784_nG555d );
and \U$2640 ( \2786 , \2634 , \2721 );
and \U$2641 ( \2787 , \2721 , \2772 );
and \U$2642 ( \2788 , \2634 , \2772 );
or \U$2643 ( \2789 , \2786 , \2787 , \2788 );
and \U$2644 ( \2790 , \2726 , \2730 );
and \U$2645 ( \2791 , \2730 , \2735 );
and \U$2646 ( \2792 , \2726 , \2735 );
or \U$2647 ( \2793 , \2790 , \2791 , \2792 );
and \U$2648 ( \2794 , \2740 , \2754 );
and \U$2649 ( \2795 , \2754 , \2770 );
and \U$2650 ( \2796 , \2740 , \2770 );
or \U$2651 ( \2797 , \2794 , \2795 , \2796 );
xor \U$2652 ( \2798 , \2793 , \2797 );
and \U$2653 ( \2799 , \2657 , \2674 );
and \U$2654 ( \2800 , \2674 , \2719 );
and \U$2655 ( \2801 , \2657 , \2719 );
or \U$2656 ( \2802 , \2799 , \2800 , \2801 );
xor \U$2657 ( \2803 , \2798 , \2802 );
xor \U$2658 ( \2804 , \2789 , \2803 );
and \U$2659 ( \2805 , \2638 , \2642 );
and \U$2660 ( \2806 , \2642 , \2720 );
and \U$2661 ( \2807 , \2638 , \2720 );
or \U$2662 ( \2808 , \2805 , \2806 , \2807 );
and \U$2663 ( \2809 , \2736 , \2771 );
xor \U$2664 ( \2810 , \2808 , \2809 );
and \U$2665 ( \2811 , \2647 , \2651 );
and \U$2666 ( \2812 , \2651 , \2656 );
and \U$2667 ( \2813 , \2647 , \2656 );
or \U$2668 ( \2814 , \2811 , \2812 , \2813 );
and \U$2669 ( \2815 , \2661 , \2665 );
and \U$2670 ( \2816 , \2665 , \2673 );
and \U$2671 ( \2817 , \2661 , \2673 );
or \U$2672 ( \2818 , \2815 , \2816 , \2817 );
xor \U$2673 ( \2819 , \2814 , \2818 );
and \U$2674 ( \2820 , \2689 , \2703 );
and \U$2675 ( \2821 , \2703 , \2718 );
and \U$2676 ( \2822 , \2689 , \2718 );
or \U$2677 ( \2823 , \2820 , \2821 , \2822 );
xor \U$2678 ( \2824 , \2819 , \2823 );
and \U$2679 ( \2825 , \2757 , \183 );
buf \U$2680 ( \2826 , RIb55e338_96);
and \U$2681 ( \2827 , \2826 , \180 );
nor \U$2682 ( \2828 , \2825 , \2827 );
xnor \U$2683 ( \2829 , \2828 , \179 );
and \U$2684 ( \2830 , \2366 , \195 );
and \U$2685 ( \2831 , \2521 , \193 );
nor \U$2686 ( \2832 , \2830 , \2831 );
xnor \U$2687 ( \2833 , \2832 , \202 );
xor \U$2688 ( \2834 , \2829 , \2833 );
buf \U$2689 ( \2835 , RIb5601b0_31);
buf \U$2690 ( \2836 , RIb560138_32);
and \U$2691 ( \2837 , \2836 , \2530 );
not \U$2692 ( \2838 , \2837 );
and \U$2693 ( \2839 , \2835 , \2838 );
xor \U$2694 ( \2840 , \2834 , \2839 );
and \U$2695 ( \2841 , \2090 , \215 );
and \U$2696 ( \2842 , \2182 , \213 );
nor \U$2697 ( \2843 , \2841 , \2842 );
xnor \U$2698 ( \2844 , \2843 , \222 );
and \U$2699 ( \2845 , \1802 , \230 );
and \U$2700 ( \2846 , \1948 , \228 );
nor \U$2701 ( \2847 , \2845 , \2846 );
xnor \U$2702 ( \2848 , \2847 , \237 );
xor \U$2703 ( \2849 , \2844 , \2848 );
and \U$2704 ( \2850 , \1601 , \245 );
and \U$2705 ( \2851 , \1684 , \243 );
nor \U$2706 ( \2852 , \2850 , \2851 );
xnor \U$2707 ( \2853 , \2852 , \252 );
xor \U$2708 ( \2854 , \2849 , \2853 );
xor \U$2709 ( \2855 , \2840 , \2854 );
and \U$2710 ( \2856 , \209 , \1578 );
and \U$2711 ( \2857 , \217 , \1431 );
nor \U$2712 ( \2858 , \2856 , \2857 );
xnor \U$2713 ( \2859 , \2858 , \1436 );
and \U$2714 ( \2860 , \224 , \1824 );
and \U$2715 ( \2861 , \232 , \1739 );
nor \U$2716 ( \2862 , \2860 , \2861 );
xnor \U$2717 ( \2863 , \2862 , \1697 );
xor \U$2718 ( \2864 , \2859 , \2863 );
and \U$2719 ( \2865 , \240 , \2121 );
and \U$2720 ( \2866 , \247 , \2008 );
nor \U$2721 ( \2867 , \2865 , \2866 );
xnor \U$2722 ( \2868 , \2867 , \1961 );
xor \U$2723 ( \2869 , \2864 , \2868 );
and \U$2724 ( \2870 , \1333 , \141 );
and \U$2725 ( \2871 , \1484 , \139 );
nor \U$2726 ( \2872 , \2870 , \2871 );
xnor \U$2727 ( \2873 , \2872 , \148 );
and \U$2728 ( \2874 , \1147 , \156 );
and \U$2729 ( \2875 , \1192 , \154 );
nor \U$2730 ( \2876 , \2874 , \2875 );
xnor \U$2731 ( \2877 , \2876 , \163 );
xor \U$2732 ( \2878 , \2873 , \2877 );
and \U$2733 ( \2879 , \412 , \296 );
and \U$2734 ( \2880 , \474 , \168 );
nor \U$2735 ( \2881 , \2879 , \2880 );
xnor \U$2736 ( \2882 , \2881 , \173 );
xor \U$2737 ( \2883 , \2878 , \2882 );
xor \U$2738 ( \2884 , \2869 , \2883 );
and \U$2739 ( \2885 , \261 , \438 );
and \U$2740 ( \2886 , \307 , \336 );
nor \U$2741 ( \2887 , \2885 , \2886 );
xnor \U$2742 ( \2888 , \2887 , \320 );
and \U$2743 ( \2889 , \178 , \1086 );
and \U$2744 ( \2890 , \185 , \508 );
nor \U$2745 ( \2891 , \2889 , \2890 );
xnor \U$2746 ( \2892 , \2891 , \487 );
xor \U$2747 ( \2893 , \2888 , \2892 );
and \U$2748 ( \2894 , \189 , \1301 );
and \U$2749 ( \2895 , \197 , \1246 );
nor \U$2750 ( \2896 , \2894 , \2895 );
xnor \U$2751 ( \2897 , \2896 , \1205 );
xor \U$2752 ( \2898 , \2893 , \2897 );
xor \U$2753 ( \2899 , \2884 , \2898 );
xor \U$2754 ( \2900 , \2855 , \2899 );
xor \U$2755 ( \2901 , \2824 , \2900 );
and \U$2756 ( \2902 , \2744 , \2748 );
and \U$2757 ( \2903 , \2748 , \2753 );
and \U$2758 ( \2904 , \2744 , \2753 );
or \U$2759 ( \2905 , \2902 , \2903 , \2904 );
and \U$2760 ( \2906 , \2760 , \2764 );
and \U$2761 ( \2907 , \2764 , \2769 );
and \U$2762 ( \2908 , \2760 , \2769 );
or \U$2763 ( \2909 , \2906 , \2907 , \2908 );
xor \U$2764 ( \2910 , \2905 , \2909 );
and \U$2765 ( \2911 , \2708 , \2712 );
and \U$2766 ( \2912 , \2712 , \2717 );
and \U$2767 ( \2913 , \2708 , \2717 );
or \U$2768 ( \2914 , \2911 , \2912 , \2913 );
xor \U$2769 ( \2915 , \2910 , \2914 );
and \U$2770 ( \2916 , \2679 , \2683 );
and \U$2771 ( \2917 , \2683 , \2688 );
and \U$2772 ( \2918 , \2679 , \2688 );
or \U$2773 ( \2919 , \2916 , \2917 , \2918 );
and \U$2774 ( \2920 , \2693 , \2697 );
and \U$2775 ( \2921 , \2697 , \2702 );
and \U$2776 ( \2922 , \2693 , \2702 );
or \U$2777 ( \2923 , \2920 , \2921 , \2922 );
xor \U$2778 ( \2924 , \2919 , \2923 );
and \U$2779 ( \2925 , \134 , \2400 );
and \U$2780 ( \2926 , \143 , \2246 );
nor \U$2781 ( \2927 , \2925 , \2926 );
xnor \U$2782 ( \2928 , \2927 , \2195 );
and \U$2783 ( \2929 , \150 , \2669 );
and \U$2784 ( \2930 , \158 , \2538 );
nor \U$2785 ( \2931 , \2929 , \2930 );
xnor \U$2786 ( \2932 , \2931 , \2534 );
xor \U$2787 ( \2933 , \2928 , \2932 );
xor \U$2788 ( \2934 , \2836 , \2530 );
nand \U$2789 ( \2935 , \166 , \2934 );
xnor \U$2790 ( \2936 , \2935 , \2839 );
xor \U$2791 ( \2937 , \2933 , \2936 );
xor \U$2792 ( \2938 , \2924 , \2937 );
xor \U$2793 ( \2939 , \2915 , \2938 );
xor \U$2794 ( \2940 , \2901 , \2939 );
xor \U$2795 ( \2941 , \2810 , \2940 );
xor \U$2796 ( \2942 , \2804 , \2941 );
and \U$2797 ( \2943 , \2628 , \2629 );
and \U$2798 ( \2944 , \2629 , \2773 );
and \U$2799 ( \2945 , \2628 , \2773 );
or \U$2800 ( \2946 , \2943 , \2944 , \2945 );
xor \U$2801 ( \2947 , \2942 , \2946 );
and \U$2802 ( \2948 , \2774 , \2778 );
and \U$2803 ( \2949 , \2779 , \2782 );
or \U$2804 ( \2950 , \2948 , \2949 );
xor \U$2805 ( \2951 , \2947 , \2950 );
buf g555b_GF_PartitionCandidate( \2952_nG555b , \2951 );
buf \U$2806 ( \2953 , \2952_nG555b );
and \U$2807 ( \2954 , \2808 , \2809 );
and \U$2808 ( \2955 , \2809 , \2940 );
and \U$2809 ( \2956 , \2808 , \2940 );
or \U$2810 ( \2957 , \2954 , \2955 , \2956 );
and \U$2811 ( \2958 , \2814 , \2818 );
and \U$2812 ( \2959 , \2818 , \2823 );
and \U$2813 ( \2960 , \2814 , \2823 );
or \U$2814 ( \2961 , \2958 , \2959 , \2960 );
and \U$2815 ( \2962 , \2840 , \2854 );
and \U$2816 ( \2963 , \2854 , \2899 );
and \U$2817 ( \2964 , \2840 , \2899 );
or \U$2818 ( \2965 , \2962 , \2963 , \2964 );
xor \U$2819 ( \2966 , \2961 , \2965 );
and \U$2820 ( \2967 , \2915 , \2938 );
xor \U$2821 ( \2968 , \2966 , \2967 );
xor \U$2822 ( \2969 , \2957 , \2968 );
and \U$2823 ( \2970 , \2793 , \2797 );
and \U$2824 ( \2971 , \2797 , \2802 );
and \U$2825 ( \2972 , \2793 , \2802 );
or \U$2826 ( \2973 , \2970 , \2971 , \2972 );
and \U$2827 ( \2974 , \2824 , \2900 );
and \U$2828 ( \2975 , \2900 , \2939 );
and \U$2829 ( \2976 , \2824 , \2939 );
or \U$2830 ( \2977 , \2974 , \2975 , \2976 );
xor \U$2831 ( \2978 , \2973 , \2977 );
and \U$2832 ( \2979 , \2873 , \2877 );
and \U$2833 ( \2980 , \2877 , \2882 );
and \U$2834 ( \2981 , \2873 , \2882 );
or \U$2835 ( \2982 , \2979 , \2980 , \2981 );
and \U$2836 ( \2983 , \2829 , \2833 );
and \U$2837 ( \2984 , \2833 , \2839 );
and \U$2838 ( \2985 , \2829 , \2839 );
or \U$2839 ( \2986 , \2983 , \2984 , \2985 );
xor \U$2840 ( \2987 , \2982 , \2986 );
and \U$2841 ( \2988 , \2844 , \2848 );
and \U$2842 ( \2989 , \2848 , \2853 );
and \U$2843 ( \2990 , \2844 , \2853 );
or \U$2844 ( \2991 , \2988 , \2989 , \2990 );
xor \U$2845 ( \2992 , \2987 , \2991 );
and \U$2846 ( \2993 , \2905 , \2909 );
and \U$2847 ( \2994 , \2909 , \2914 );
and \U$2848 ( \2995 , \2905 , \2914 );
or \U$2849 ( \2996 , \2993 , \2994 , \2995 );
and \U$2850 ( \2997 , \2869 , \2883 );
and \U$2851 ( \2998 , \2883 , \2898 );
and \U$2852 ( \2999 , \2869 , \2898 );
or \U$2853 ( \3000 , \2997 , \2998 , \2999 );
xor \U$2854 ( \3001 , \2996 , \3000 );
and \U$2855 ( \3002 , \2919 , \2923 );
and \U$2856 ( \3003 , \2923 , \2937 );
and \U$2857 ( \3004 , \2919 , \2937 );
or \U$2858 ( \3005 , \3002 , \3003 , \3004 );
xor \U$2859 ( \3006 , \3001 , \3005 );
xor \U$2860 ( \3007 , \2992 , \3006 );
and \U$2861 ( \3008 , \2859 , \2863 );
and \U$2862 ( \3009 , \2863 , \2868 );
and \U$2863 ( \3010 , \2859 , \2868 );
or \U$2864 ( \3011 , \3008 , \3009 , \3010 );
and \U$2865 ( \3012 , \2928 , \2932 );
and \U$2866 ( \3013 , \2932 , \2936 );
and \U$2867 ( \3014 , \2928 , \2936 );
or \U$2868 ( \3015 , \3012 , \3013 , \3014 );
xor \U$2869 ( \3016 , \3011 , \3015 );
and \U$2870 ( \3017 , \2888 , \2892 );
and \U$2871 ( \3018 , \2892 , \2897 );
and \U$2872 ( \3019 , \2888 , \2897 );
or \U$2873 ( \3020 , \3017 , \3018 , \3019 );
xor \U$2874 ( \3021 , \3016 , \3020 );
and \U$2875 ( \3022 , \1192 , \156 );
and \U$2876 ( \3023 , \1333 , \154 );
nor \U$2877 ( \3024 , \3022 , \3023 );
xnor \U$2878 ( \3025 , \3024 , \163 );
and \U$2879 ( \3026 , \474 , \296 );
and \U$2880 ( \3027 , \1147 , \168 );
nor \U$2881 ( \3028 , \3026 , \3027 );
xnor \U$2882 ( \3029 , \3028 , \173 );
xor \U$2883 ( \3030 , \3025 , \3029 );
and \U$2884 ( \3031 , \307 , \438 );
and \U$2885 ( \3032 , \412 , \336 );
nor \U$2886 ( \3033 , \3031 , \3032 );
xnor \U$2887 ( \3034 , \3033 , \320 );
xor \U$2888 ( \3035 , \3030 , \3034 );
and \U$2889 ( \3036 , \2826 , \183 );
buf \U$2890 ( \3037 , RIb55e3b0_95);
and \U$2891 ( \3038 , \3037 , \180 );
nor \U$2892 ( \3039 , \3036 , \3038 );
xnor \U$2893 ( \3040 , \3039 , \179 );
and \U$2894 ( \3041 , \2521 , \195 );
and \U$2895 ( \3042 , \2757 , \193 );
nor \U$2896 ( \3043 , \3041 , \3042 );
xnor \U$2897 ( \3044 , \3043 , \202 );
xor \U$2898 ( \3045 , \3040 , \3044 );
and \U$2899 ( \3046 , \2182 , \215 );
and \U$2900 ( \3047 , \2366 , \213 );
nor \U$2901 ( \3048 , \3046 , \3047 );
xnor \U$2902 ( \3049 , \3048 , \222 );
xor \U$2903 ( \3050 , \3045 , \3049 );
xor \U$2904 ( \3051 , \3035 , \3050 );
and \U$2905 ( \3052 , \1948 , \230 );
and \U$2906 ( \3053 , \2090 , \228 );
nor \U$2907 ( \3054 , \3052 , \3053 );
xnor \U$2908 ( \3055 , \3054 , \237 );
and \U$2909 ( \3056 , \1684 , \245 );
and \U$2910 ( \3057 , \1802 , \243 );
nor \U$2911 ( \3058 , \3056 , \3057 );
xnor \U$2912 ( \3059 , \3058 , \252 );
xor \U$2913 ( \3060 , \3055 , \3059 );
and \U$2914 ( \3061 , \1484 , \141 );
and \U$2915 ( \3062 , \1601 , \139 );
nor \U$2916 ( \3063 , \3061 , \3062 );
xnor \U$2917 ( \3064 , \3063 , \148 );
xor \U$2918 ( \3065 , \3060 , \3064 );
xor \U$2919 ( \3066 , \3051 , \3065 );
xor \U$2920 ( \3067 , \3021 , \3066 );
and \U$2921 ( \3068 , \232 , \1824 );
and \U$2922 ( \3069 , \209 , \1739 );
nor \U$2923 ( \3070 , \3068 , \3069 );
xnor \U$2924 ( \3071 , \3070 , \1697 );
and \U$2925 ( \3072 , \247 , \2121 );
and \U$2926 ( \3073 , \224 , \2008 );
nor \U$2927 ( \3074 , \3072 , \3073 );
xnor \U$2928 ( \3075 , \3074 , \1961 );
xor \U$2929 ( \3076 , \3071 , \3075 );
and \U$2930 ( \3077 , \143 , \2400 );
and \U$2931 ( \3078 , \240 , \2246 );
nor \U$2932 ( \3079 , \3077 , \3078 );
xnor \U$2933 ( \3080 , \3079 , \2195 );
xor \U$2934 ( \3081 , \3076 , \3080 );
and \U$2935 ( \3082 , \185 , \1086 );
and \U$2936 ( \3083 , \261 , \508 );
nor \U$2937 ( \3084 , \3082 , \3083 );
xnor \U$2938 ( \3085 , \3084 , \487 );
and \U$2939 ( \3086 , \197 , \1301 );
and \U$2940 ( \3087 , \178 , \1246 );
nor \U$2941 ( \3088 , \3086 , \3087 );
xnor \U$2942 ( \3089 , \3088 , \1205 );
xor \U$2943 ( \3090 , \3085 , \3089 );
and \U$2944 ( \3091 , \217 , \1578 );
and \U$2945 ( \3092 , \189 , \1431 );
nor \U$2946 ( \3093 , \3091 , \3092 );
xnor \U$2947 ( \3094 , \3093 , \1436 );
xor \U$2948 ( \3095 , \3090 , \3094 );
xor \U$2949 ( \3096 , \3081 , \3095 );
and \U$2950 ( \3097 , \158 , \2669 );
and \U$2951 ( \3098 , \134 , \2538 );
nor \U$2952 ( \3099 , \3097 , \3098 );
xnor \U$2953 ( \3100 , \3099 , \2534 );
xor \U$2954 ( \3101 , \2835 , \2836 );
not \U$2955 ( \3102 , \2934 );
and \U$2956 ( \3103 , \3101 , \3102 );
and \U$2957 ( \3104 , \166 , \3103 );
and \U$2958 ( \3105 , \150 , \2934 );
nor \U$2959 ( \3106 , \3104 , \3105 );
xnor \U$2960 ( \3107 , \3106 , \2839 );
xor \U$2961 ( \3108 , \3100 , \3107 );
xor \U$2962 ( \3109 , \3096 , \3108 );
xor \U$2963 ( \3110 , \3067 , \3109 );
xor \U$2964 ( \3111 , \3007 , \3110 );
xor \U$2965 ( \3112 , \2978 , \3111 );
xor \U$2966 ( \3113 , \2969 , \3112 );
and \U$2967 ( \3114 , \2789 , \2803 );
and \U$2968 ( \3115 , \2803 , \2941 );
and \U$2969 ( \3116 , \2789 , \2941 );
or \U$2970 ( \3117 , \3114 , \3115 , \3116 );
xor \U$2971 ( \3118 , \3113 , \3117 );
and \U$2972 ( \3119 , \2942 , \2946 );
and \U$2973 ( \3120 , \2947 , \2950 );
or \U$2974 ( \3121 , \3119 , \3120 );
xor \U$2975 ( \3122 , \3118 , \3121 );
buf g5559_GF_PartitionCandidate( \3123_nG5559 , \3122 );
buf \U$2976 ( \3124 , \3123_nG5559 );
and \U$2977 ( \3125 , \2973 , \2977 );
and \U$2978 ( \3126 , \2977 , \3111 );
and \U$2979 ( \3127 , \2973 , \3111 );
or \U$2980 ( \3128 , \3125 , \3126 , \3127 );
and \U$2981 ( \3129 , \2961 , \2965 );
and \U$2982 ( \3130 , \2965 , \2967 );
and \U$2983 ( \3131 , \2961 , \2967 );
or \U$2984 ( \3132 , \3129 , \3130 , \3131 );
and \U$2985 ( \3133 , \2992 , \3006 );
and \U$2986 ( \3134 , \3006 , \3110 );
and \U$2987 ( \3135 , \2992 , \3110 );
or \U$2988 ( \3136 , \3133 , \3134 , \3135 );
xor \U$2989 ( \3137 , \3132 , \3136 );
and \U$2990 ( \3138 , \3035 , \3050 );
and \U$2991 ( \3139 , \3050 , \3065 );
and \U$2992 ( \3140 , \3035 , \3065 );
or \U$2993 ( \3141 , \3138 , \3139 , \3140 );
and \U$2994 ( \3142 , \3037 , \183 );
buf \U$2995 ( \3143 , RIb55e428_94);
and \U$2996 ( \3144 , \3143 , \180 );
nor \U$2997 ( \3145 , \3142 , \3144 );
xnor \U$2998 ( \3146 , \3145 , \179 );
and \U$2999 ( \3147 , \2757 , \195 );
and \U$3000 ( \3148 , \2826 , \193 );
nor \U$3001 ( \3149 , \3147 , \3148 );
xnor \U$3002 ( \3150 , \3149 , \202 );
xor \U$3003 ( \3151 , \3146 , \3150 );
buf \U$3004 ( \3152 , RIb5602a0_29);
buf \U$3005 ( \3153 , RIb560228_30);
and \U$3006 ( \3154 , \3153 , \2835 );
not \U$3007 ( \3155 , \3154 );
and \U$3008 ( \3156 , \3152 , \3155 );
xor \U$3009 ( \3157 , \3151 , \3156 );
xor \U$3010 ( \3158 , \3141 , \3157 );
and \U$3011 ( \3159 , \2366 , \215 );
and \U$3012 ( \3160 , \2521 , \213 );
nor \U$3013 ( \3161 , \3159 , \3160 );
xnor \U$3014 ( \3162 , \3161 , \222 );
and \U$3015 ( \3163 , \2090 , \230 );
and \U$3016 ( \3164 , \2182 , \228 );
nor \U$3017 ( \3165 , \3163 , \3164 );
xnor \U$3018 ( \3166 , \3165 , \237 );
xor \U$3019 ( \3167 , \3162 , \3166 );
and \U$3020 ( \3168 , \1802 , \245 );
and \U$3021 ( \3169 , \1948 , \243 );
nor \U$3022 ( \3170 , \3168 , \3169 );
xnor \U$3023 ( \3171 , \3170 , \252 );
xor \U$3024 ( \3172 , \3167 , \3171 );
and \U$3025 ( \3173 , \412 , \438 );
and \U$3026 ( \3174 , \474 , \336 );
nor \U$3027 ( \3175 , \3173 , \3174 );
xnor \U$3028 ( \3176 , \3175 , \320 );
and \U$3029 ( \3177 , \261 , \1086 );
and \U$3030 ( \3178 , \307 , \508 );
nor \U$3031 ( \3179 , \3177 , \3178 );
xnor \U$3032 ( \3180 , \3179 , \487 );
xor \U$3033 ( \3181 , \3176 , \3180 );
and \U$3034 ( \3182 , \178 , \1301 );
and \U$3035 ( \3183 , \185 , \1246 );
nor \U$3036 ( \3184 , \3182 , \3183 );
xnor \U$3037 ( \3185 , \3184 , \1205 );
xor \U$3038 ( \3186 , \3181 , \3185 );
xor \U$3039 ( \3187 , \3172 , \3186 );
and \U$3040 ( \3188 , \1601 , \141 );
and \U$3041 ( \3189 , \1684 , \139 );
nor \U$3042 ( \3190 , \3188 , \3189 );
xnor \U$3043 ( \3191 , \3190 , \148 );
and \U$3044 ( \3192 , \1333 , \156 );
and \U$3045 ( \3193 , \1484 , \154 );
nor \U$3046 ( \3194 , \3192 , \3193 );
xnor \U$3047 ( \3195 , \3194 , \163 );
xor \U$3048 ( \3196 , \3191 , \3195 );
and \U$3049 ( \3197 , \1147 , \296 );
and \U$3050 ( \3198 , \1192 , \168 );
nor \U$3051 ( \3199 , \3197 , \3198 );
xnor \U$3052 ( \3200 , \3199 , \173 );
xor \U$3053 ( \3201 , \3196 , \3200 );
xor \U$3054 ( \3202 , \3187 , \3201 );
xor \U$3055 ( \3203 , \3158 , \3202 );
xor \U$3056 ( \3204 , \3137 , \3203 );
xor \U$3057 ( \3205 , \3128 , \3204 );
and \U$3058 ( \3206 , \3011 , \3015 );
and \U$3059 ( \3207 , \3015 , \3020 );
and \U$3060 ( \3208 , \3011 , \3020 );
or \U$3061 ( \3209 , \3206 , \3207 , \3208 );
and \U$3062 ( \3210 , \2982 , \2986 );
and \U$3063 ( \3211 , \2986 , \2991 );
and \U$3064 ( \3212 , \2982 , \2991 );
or \U$3065 ( \3213 , \3210 , \3211 , \3212 );
xor \U$3066 ( \3214 , \3209 , \3213 );
and \U$3067 ( \3215 , \3081 , \3095 );
and \U$3068 ( \3216 , \3095 , \3108 );
and \U$3069 ( \3217 , \3081 , \3108 );
or \U$3070 ( \3218 , \3215 , \3216 , \3217 );
xor \U$3071 ( \3219 , \3214 , \3218 );
and \U$3072 ( \3220 , \2996 , \3000 );
and \U$3073 ( \3221 , \3000 , \3005 );
and \U$3074 ( \3222 , \2996 , \3005 );
or \U$3075 ( \3223 , \3220 , \3221 , \3222 );
and \U$3076 ( \3224 , \3021 , \3066 );
and \U$3077 ( \3225 , \3066 , \3109 );
and \U$3078 ( \3226 , \3021 , \3109 );
or \U$3079 ( \3227 , \3224 , \3225 , \3226 );
xor \U$3080 ( \3228 , \3223 , \3227 );
and \U$3081 ( \3229 , \3025 , \3029 );
and \U$3082 ( \3230 , \3029 , \3034 );
and \U$3083 ( \3231 , \3025 , \3034 );
or \U$3084 ( \3232 , \3229 , \3230 , \3231 );
and \U$3085 ( \3233 , \3040 , \3044 );
and \U$3086 ( \3234 , \3044 , \3049 );
and \U$3087 ( \3235 , \3040 , \3049 );
or \U$3088 ( \3236 , \3233 , \3234 , \3235 );
xor \U$3089 ( \3237 , \3232 , \3236 );
and \U$3090 ( \3238 , \3055 , \3059 );
and \U$3091 ( \3239 , \3059 , \3064 );
and \U$3092 ( \3240 , \3055 , \3064 );
or \U$3093 ( \3241 , \3238 , \3239 , \3240 );
xor \U$3094 ( \3242 , \3237 , \3241 );
and \U$3095 ( \3243 , \3071 , \3075 );
and \U$3096 ( \3244 , \3075 , \3080 );
and \U$3097 ( \3245 , \3071 , \3080 );
or \U$3098 ( \3246 , \3243 , \3244 , \3245 );
and \U$3099 ( \3247 , \3085 , \3089 );
and \U$3100 ( \3248 , \3089 , \3094 );
and \U$3101 ( \3249 , \3085 , \3094 );
or \U$3102 ( \3250 , \3247 , \3248 , \3249 );
xor \U$3103 ( \3251 , \3246 , \3250 );
and \U$3104 ( \3252 , \3100 , \3107 );
xor \U$3105 ( \3253 , \3251 , \3252 );
xor \U$3106 ( \3254 , \3242 , \3253 );
xor \U$3107 ( \3255 , \3153 , \2835 );
nand \U$3108 ( \3256 , \166 , \3255 );
xnor \U$3109 ( \3257 , \3256 , \3156 );
and \U$3110 ( \3258 , \189 , \1578 );
and \U$3111 ( \3259 , \197 , \1431 );
nor \U$3112 ( \3260 , \3258 , \3259 );
xnor \U$3113 ( \3261 , \3260 , \1436 );
and \U$3114 ( \3262 , \209 , \1824 );
and \U$3115 ( \3263 , \217 , \1739 );
nor \U$3116 ( \3264 , \3262 , \3263 );
xnor \U$3117 ( \3265 , \3264 , \1697 );
xor \U$3118 ( \3266 , \3261 , \3265 );
and \U$3119 ( \3267 , \224 , \2121 );
and \U$3120 ( \3268 , \232 , \2008 );
nor \U$3121 ( \3269 , \3267 , \3268 );
xnor \U$3122 ( \3270 , \3269 , \1961 );
xor \U$3123 ( \3271 , \3266 , \3270 );
xor \U$3124 ( \3272 , \3257 , \3271 );
and \U$3125 ( \3273 , \240 , \2400 );
and \U$3126 ( \3274 , \247 , \2246 );
nor \U$3127 ( \3275 , \3273 , \3274 );
xnor \U$3128 ( \3276 , \3275 , \2195 );
and \U$3129 ( \3277 , \134 , \2669 );
and \U$3130 ( \3278 , \143 , \2538 );
nor \U$3131 ( \3279 , \3277 , \3278 );
xnor \U$3132 ( \3280 , \3279 , \2534 );
xor \U$3133 ( \3281 , \3276 , \3280 );
and \U$3134 ( \3282 , \150 , \3103 );
and \U$3135 ( \3283 , \158 , \2934 );
nor \U$3136 ( \3284 , \3282 , \3283 );
xnor \U$3137 ( \3285 , \3284 , \2839 );
xor \U$3138 ( \3286 , \3281 , \3285 );
xor \U$3139 ( \3287 , \3272 , \3286 );
xor \U$3140 ( \3288 , \3254 , \3287 );
xor \U$3141 ( \3289 , \3228 , \3288 );
xor \U$3142 ( \3290 , \3219 , \3289 );
xor \U$3143 ( \3291 , \3205 , \3290 );
and \U$3144 ( \3292 , \2957 , \2968 );
and \U$3145 ( \3293 , \2968 , \3112 );
and \U$3146 ( \3294 , \2957 , \3112 );
or \U$3147 ( \3295 , \3292 , \3293 , \3294 );
xor \U$3148 ( \3296 , \3291 , \3295 );
and \U$3149 ( \3297 , \3113 , \3117 );
and \U$3150 ( \3298 , \3118 , \3121 );
or \U$3151 ( \3299 , \3297 , \3298 );
xor \U$3152 ( \3300 , \3296 , \3299 );
buf g5557_GF_PartitionCandidate( \3301_nG5557 , \3300 );
buf \U$3153 ( \3302 , \3301_nG5557 );
and \U$3154 ( \3303 , \3132 , \3136 );
and \U$3155 ( \3304 , \3136 , \3203 );
and \U$3156 ( \3305 , \3132 , \3203 );
or \U$3157 ( \3306 , \3303 , \3304 , \3305 );
and \U$3158 ( \3307 , \3219 , \3289 );
xor \U$3159 ( \3308 , \3306 , \3307 );
and \U$3160 ( \3309 , \3223 , \3227 );
and \U$3161 ( \3310 , \3227 , \3288 );
and \U$3162 ( \3311 , \3223 , \3288 );
or \U$3163 ( \3312 , \3309 , \3310 , \3311 );
and \U$3164 ( \3313 , \3209 , \3213 );
and \U$3165 ( \3314 , \3213 , \3218 );
and \U$3166 ( \3315 , \3209 , \3218 );
or \U$3167 ( \3316 , \3313 , \3314 , \3315 );
and \U$3168 ( \3317 , \3141 , \3157 );
and \U$3169 ( \3318 , \3157 , \3202 );
and \U$3170 ( \3319 , \3141 , \3202 );
or \U$3171 ( \3320 , \3317 , \3318 , \3319 );
xor \U$3172 ( \3321 , \3316 , \3320 );
and \U$3173 ( \3322 , \3242 , \3253 );
and \U$3174 ( \3323 , \3253 , \3287 );
and \U$3175 ( \3324 , \3242 , \3287 );
or \U$3176 ( \3325 , \3322 , \3323 , \3324 );
xor \U$3177 ( \3326 , \3321 , \3325 );
xor \U$3178 ( \3327 , \3312 , \3326 );
and \U$3179 ( \3328 , \3232 , \3236 );
and \U$3180 ( \3329 , \3236 , \3241 );
and \U$3181 ( \3330 , \3232 , \3241 );
or \U$3182 ( \3331 , \3328 , \3329 , \3330 );
and \U$3183 ( \3332 , \3246 , \3250 );
and \U$3184 ( \3333 , \3250 , \3252 );
and \U$3185 ( \3334 , \3246 , \3252 );
or \U$3186 ( \3335 , \3332 , \3333 , \3334 );
xor \U$3187 ( \3336 , \3331 , \3335 );
and \U$3188 ( \3337 , \3257 , \3271 );
and \U$3189 ( \3338 , \3271 , \3286 );
and \U$3190 ( \3339 , \3257 , \3286 );
or \U$3191 ( \3340 , \3337 , \3338 , \3339 );
xor \U$3192 ( \3341 , \3336 , \3340 );
and \U$3193 ( \3342 , \3172 , \3186 );
and \U$3194 ( \3343 , \3186 , \3201 );
and \U$3195 ( \3344 , \3172 , \3201 );
or \U$3196 ( \3345 , \3342 , \3343 , \3344 );
and \U$3197 ( \3346 , \143 , \2669 );
and \U$3198 ( \3347 , \240 , \2538 );
nor \U$3199 ( \3348 , \3346 , \3347 );
xnor \U$3200 ( \3349 , \3348 , \2534 );
and \U$3201 ( \3350 , \158 , \3103 );
and \U$3202 ( \3351 , \134 , \2934 );
nor \U$3203 ( \3352 , \3350 , \3351 );
xnor \U$3204 ( \3353 , \3352 , \2839 );
xor \U$3205 ( \3354 , \3349 , \3353 );
xor \U$3206 ( \3355 , \3152 , \3153 );
not \U$3207 ( \3356 , \3255 );
and \U$3208 ( \3357 , \3355 , \3356 );
and \U$3209 ( \3358 , \166 , \3357 );
and \U$3210 ( \3359 , \150 , \3255 );
nor \U$3211 ( \3360 , \3358 , \3359 );
xnor \U$3212 ( \3361 , \3360 , \3156 );
xor \U$3213 ( \3362 , \3354 , \3361 );
and \U$3214 ( \3363 , \217 , \1824 );
and \U$3215 ( \3364 , \189 , \1739 );
nor \U$3216 ( \3365 , \3363 , \3364 );
xnor \U$3217 ( \3366 , \3365 , \1697 );
and \U$3218 ( \3367 , \232 , \2121 );
and \U$3219 ( \3368 , \209 , \2008 );
nor \U$3220 ( \3369 , \3367 , \3368 );
xnor \U$3221 ( \3370 , \3369 , \1961 );
xor \U$3222 ( \3371 , \3366 , \3370 );
and \U$3223 ( \3372 , \247 , \2400 );
and \U$3224 ( \3373 , \224 , \2246 );
nor \U$3225 ( \3374 , \3372 , \3373 );
xnor \U$3226 ( \3375 , \3374 , \2195 );
xor \U$3227 ( \3376 , \3371 , \3375 );
xor \U$3228 ( \3377 , \3362 , \3376 );
and \U$3229 ( \3378 , \307 , \1086 );
and \U$3230 ( \3379 , \412 , \508 );
nor \U$3231 ( \3380 , \3378 , \3379 );
xnor \U$3232 ( \3381 , \3380 , \487 );
and \U$3233 ( \3382 , \185 , \1301 );
and \U$3234 ( \3383 , \261 , \1246 );
nor \U$3235 ( \3384 , \3382 , \3383 );
xnor \U$3236 ( \3385 , \3384 , \1205 );
xor \U$3237 ( \3386 , \3381 , \3385 );
and \U$3238 ( \3387 , \197 , \1578 );
and \U$3239 ( \3388 , \178 , \1431 );
nor \U$3240 ( \3389 , \3387 , \3388 );
xnor \U$3241 ( \3390 , \3389 , \1436 );
xor \U$3242 ( \3391 , \3386 , \3390 );
xor \U$3243 ( \3392 , \3377 , \3391 );
xor \U$3244 ( \3393 , \3345 , \3392 );
and \U$3245 ( \3394 , \3143 , \183 );
buf \U$3246 ( \3395 , RIb55e4a0_93);
and \U$3247 ( \3396 , \3395 , \180 );
nor \U$3248 ( \3397 , \3394 , \3396 );
xnor \U$3249 ( \3398 , \3397 , \179 );
and \U$3250 ( \3399 , \2826 , \195 );
and \U$3251 ( \3400 , \3037 , \193 );
nor \U$3252 ( \3401 , \3399 , \3400 );
xnor \U$3253 ( \3402 , \3401 , \202 );
xor \U$3254 ( \3403 , \3398 , \3402 );
and \U$3255 ( \3404 , \2521 , \215 );
and \U$3256 ( \3405 , \2757 , \213 );
nor \U$3257 ( \3406 , \3404 , \3405 );
xnor \U$3258 ( \3407 , \3406 , \222 );
xor \U$3259 ( \3408 , \3403 , \3407 );
and \U$3260 ( \3409 , \2182 , \230 );
and \U$3261 ( \3410 , \2366 , \228 );
nor \U$3262 ( \3411 , \3409 , \3410 );
xnor \U$3263 ( \3412 , \3411 , \237 );
and \U$3264 ( \3413 , \1948 , \245 );
and \U$3265 ( \3414 , \2090 , \243 );
nor \U$3266 ( \3415 , \3413 , \3414 );
xnor \U$3267 ( \3416 , \3415 , \252 );
xor \U$3268 ( \3417 , \3412 , \3416 );
and \U$3269 ( \3418 , \1684 , \141 );
and \U$3270 ( \3419 , \1802 , \139 );
nor \U$3271 ( \3420 , \3418 , \3419 );
xnor \U$3272 ( \3421 , \3420 , \148 );
xor \U$3273 ( \3422 , \3417 , \3421 );
xor \U$3274 ( \3423 , \3408 , \3422 );
and \U$3275 ( \3424 , \1484 , \156 );
and \U$3276 ( \3425 , \1601 , \154 );
nor \U$3277 ( \3426 , \3424 , \3425 );
xnor \U$3278 ( \3427 , \3426 , \163 );
and \U$3279 ( \3428 , \1192 , \296 );
and \U$3280 ( \3429 , \1333 , \168 );
nor \U$3281 ( \3430 , \3428 , \3429 );
xnor \U$3282 ( \3431 , \3430 , \173 );
xor \U$3283 ( \3432 , \3427 , \3431 );
and \U$3284 ( \3433 , \474 , \438 );
and \U$3285 ( \3434 , \1147 , \336 );
nor \U$3286 ( \3435 , \3433 , \3434 );
xnor \U$3287 ( \3436 , \3435 , \320 );
xor \U$3288 ( \3437 , \3432 , \3436 );
xor \U$3289 ( \3438 , \3423 , \3437 );
xor \U$3290 ( \3439 , \3393 , \3438 );
xor \U$3291 ( \3440 , \3341 , \3439 );
and \U$3292 ( \3441 , \3146 , \3150 );
and \U$3293 ( \3442 , \3150 , \3156 );
and \U$3294 ( \3443 , \3146 , \3156 );
or \U$3295 ( \3444 , \3441 , \3442 , \3443 );
and \U$3296 ( \3445 , \3162 , \3166 );
and \U$3297 ( \3446 , \3166 , \3171 );
and \U$3298 ( \3447 , \3162 , \3171 );
or \U$3299 ( \3448 , \3445 , \3446 , \3447 );
xor \U$3300 ( \3449 , \3444 , \3448 );
and \U$3301 ( \3450 , \3191 , \3195 );
and \U$3302 ( \3451 , \3195 , \3200 );
and \U$3303 ( \3452 , \3191 , \3200 );
or \U$3304 ( \3453 , \3450 , \3451 , \3452 );
xor \U$3305 ( \3454 , \3449 , \3453 );
and \U$3306 ( \3455 , \3176 , \3180 );
and \U$3307 ( \3456 , \3180 , \3185 );
and \U$3308 ( \3457 , \3176 , \3185 );
or \U$3309 ( \3458 , \3455 , \3456 , \3457 );
and \U$3310 ( \3459 , \3261 , \3265 );
and \U$3311 ( \3460 , \3265 , \3270 );
and \U$3312 ( \3461 , \3261 , \3270 );
or \U$3313 ( \3462 , \3459 , \3460 , \3461 );
xor \U$3314 ( \3463 , \3458 , \3462 );
and \U$3315 ( \3464 , \3276 , \3280 );
and \U$3316 ( \3465 , \3280 , \3285 );
and \U$3317 ( \3466 , \3276 , \3285 );
or \U$3318 ( \3467 , \3464 , \3465 , \3466 );
xor \U$3319 ( \3468 , \3463 , \3467 );
xor \U$3320 ( \3469 , \3454 , \3468 );
xor \U$3321 ( \3470 , \3440 , \3469 );
xor \U$3322 ( \3471 , \3327 , \3470 );
xor \U$3323 ( \3472 , \3308 , \3471 );
and \U$3324 ( \3473 , \3128 , \3204 );
and \U$3325 ( \3474 , \3204 , \3290 );
and \U$3326 ( \3475 , \3128 , \3290 );
or \U$3327 ( \3476 , \3473 , \3474 , \3475 );
xor \U$3328 ( \3477 , \3472 , \3476 );
and \U$3329 ( \3478 , \3291 , \3295 );
and \U$3330 ( \3479 , \3296 , \3299 );
or \U$3331 ( \3480 , \3478 , \3479 );
xor \U$3332 ( \3481 , \3477 , \3480 );
buf g5555_GF_PartitionCandidate( \3482_nG5555 , \3481 );
buf \U$3333 ( \3483 , \3482_nG5555 );
and \U$3334 ( \3484 , \3312 , \3326 );
and \U$3335 ( \3485 , \3326 , \3470 );
and \U$3336 ( \3486 , \3312 , \3470 );
or \U$3337 ( \3487 , \3484 , \3485 , \3486 );
and \U$3338 ( \3488 , \3331 , \3335 );
and \U$3339 ( \3489 , \3335 , \3340 );
and \U$3340 ( \3490 , \3331 , \3340 );
or \U$3341 ( \3491 , \3488 , \3489 , \3490 );
and \U$3342 ( \3492 , \3345 , \3392 );
and \U$3343 ( \3493 , \3392 , \3438 );
and \U$3344 ( \3494 , \3345 , \3438 );
or \U$3345 ( \3495 , \3492 , \3493 , \3494 );
xor \U$3346 ( \3496 , \3491 , \3495 );
and \U$3347 ( \3497 , \3454 , \3468 );
xor \U$3348 ( \3498 , \3496 , \3497 );
xor \U$3349 ( \3499 , \3487 , \3498 );
and \U$3350 ( \3500 , \3316 , \3320 );
and \U$3351 ( \3501 , \3320 , \3325 );
and \U$3352 ( \3502 , \3316 , \3325 );
or \U$3353 ( \3503 , \3500 , \3501 , \3502 );
and \U$3354 ( \3504 , \3341 , \3439 );
and \U$3355 ( \3505 , \3439 , \3469 );
and \U$3356 ( \3506 , \3341 , \3469 );
or \U$3357 ( \3507 , \3504 , \3505 , \3506 );
xor \U$3358 ( \3508 , \3503 , \3507 );
and \U$3359 ( \3509 , \3444 , \3448 );
and \U$3360 ( \3510 , \3448 , \3453 );
and \U$3361 ( \3511 , \3444 , \3453 );
or \U$3362 ( \3512 , \3509 , \3510 , \3511 );
and \U$3363 ( \3513 , \3458 , \3462 );
and \U$3364 ( \3514 , \3462 , \3467 );
and \U$3365 ( \3515 , \3458 , \3467 );
or \U$3366 ( \3516 , \3513 , \3514 , \3515 );
xor \U$3367 ( \3517 , \3512 , \3516 );
and \U$3368 ( \3518 , \3362 , \3376 );
and \U$3369 ( \3519 , \3376 , \3391 );
and \U$3370 ( \3520 , \3362 , \3391 );
or \U$3371 ( \3521 , \3518 , \3519 , \3520 );
xor \U$3372 ( \3522 , \3517 , \3521 );
and \U$3373 ( \3523 , \3398 , \3402 );
and \U$3374 ( \3524 , \3402 , \3407 );
and \U$3375 ( \3525 , \3398 , \3407 );
or \U$3376 ( \3526 , \3523 , \3524 , \3525 );
and \U$3377 ( \3527 , \3412 , \3416 );
and \U$3378 ( \3528 , \3416 , \3421 );
and \U$3379 ( \3529 , \3412 , \3421 );
or \U$3380 ( \3530 , \3527 , \3528 , \3529 );
xor \U$3381 ( \3531 , \3526 , \3530 );
and \U$3382 ( \3532 , \3427 , \3431 );
and \U$3383 ( \3533 , \3431 , \3436 );
and \U$3384 ( \3534 , \3427 , \3436 );
or \U$3385 ( \3535 , \3532 , \3533 , \3534 );
xor \U$3386 ( \3536 , \3531 , \3535 );
and \U$3387 ( \3537 , \3349 , \3353 );
and \U$3388 ( \3538 , \3353 , \3361 );
and \U$3389 ( \3539 , \3349 , \3361 );
or \U$3390 ( \3540 , \3537 , \3538 , \3539 );
and \U$3391 ( \3541 , \3366 , \3370 );
and \U$3392 ( \3542 , \3370 , \3375 );
and \U$3393 ( \3543 , \3366 , \3375 );
or \U$3394 ( \3544 , \3541 , \3542 , \3543 );
xor \U$3395 ( \3545 , \3540 , \3544 );
and \U$3396 ( \3546 , \3381 , \3385 );
and \U$3397 ( \3547 , \3385 , \3390 );
and \U$3398 ( \3548 , \3381 , \3390 );
or \U$3399 ( \3549 , \3546 , \3547 , \3548 );
xor \U$3400 ( \3550 , \3545 , \3549 );
xor \U$3401 ( \3551 , \3536 , \3550 );
and \U$3402 ( \3552 , \150 , \3357 );
and \U$3403 ( \3553 , \158 , \3255 );
nor \U$3404 ( \3554 , \3552 , \3553 );
xnor \U$3405 ( \3555 , \3554 , \3156 );
buf \U$3406 ( \3556 , RIb560318_28);
xor \U$3407 ( \3557 , \3556 , \3152 );
nand \U$3408 ( \3558 , \166 , \3557 );
buf \U$3409 ( \3559 , RIb560390_27);
and \U$3410 ( \3560 , \3556 , \3152 );
not \U$3411 ( \3561 , \3560 );
and \U$3412 ( \3562 , \3559 , \3561 );
xnor \U$3413 ( \3563 , \3558 , \3562 );
xor \U$3414 ( \3564 , \3555 , \3563 );
and \U$3415 ( \3565 , \224 , \2400 );
and \U$3416 ( \3566 , \232 , \2246 );
nor \U$3417 ( \3567 , \3565 , \3566 );
xnor \U$3418 ( \3568 , \3567 , \2195 );
and \U$3419 ( \3569 , \240 , \2669 );
and \U$3420 ( \3570 , \247 , \2538 );
nor \U$3421 ( \3571 , \3569 , \3570 );
xnor \U$3422 ( \3572 , \3571 , \2534 );
xor \U$3423 ( \3573 , \3568 , \3572 );
and \U$3424 ( \3574 , \134 , \3103 );
and \U$3425 ( \3575 , \143 , \2934 );
nor \U$3426 ( \3576 , \3574 , \3575 );
xnor \U$3427 ( \3577 , \3576 , \2839 );
xor \U$3428 ( \3578 , \3573 , \3577 );
xor \U$3429 ( \3579 , \3564 , \3578 );
xor \U$3430 ( \3580 , \3551 , \3579 );
xor \U$3431 ( \3581 , \3522 , \3580 );
and \U$3432 ( \3582 , \3408 , \3422 );
and \U$3433 ( \3583 , \3422 , \3437 );
and \U$3434 ( \3584 , \3408 , \3437 );
or \U$3435 ( \3585 , \3582 , \3583 , \3584 );
and \U$3436 ( \3586 , \1802 , \141 );
and \U$3437 ( \3587 , \1948 , \139 );
nor \U$3438 ( \3588 , \3586 , \3587 );
xnor \U$3439 ( \3589 , \3588 , \148 );
and \U$3440 ( \3590 , \1601 , \156 );
and \U$3441 ( \3591 , \1684 , \154 );
nor \U$3442 ( \3592 , \3590 , \3591 );
xnor \U$3443 ( \3593 , \3592 , \163 );
xor \U$3444 ( \3594 , \3589 , \3593 );
and \U$3445 ( \3595 , \1333 , \296 );
and \U$3446 ( \3596 , \1484 , \168 );
nor \U$3447 ( \3597 , \3595 , \3596 );
xnor \U$3448 ( \3598 , \3597 , \173 );
xor \U$3449 ( \3599 , \3594 , \3598 );
and \U$3450 ( \3600 , \1147 , \438 );
and \U$3451 ( \3601 , \1192 , \336 );
nor \U$3452 ( \3602 , \3600 , \3601 );
xnor \U$3453 ( \3603 , \3602 , \320 );
and \U$3454 ( \3604 , \412 , \1086 );
and \U$3455 ( \3605 , \474 , \508 );
nor \U$3456 ( \3606 , \3604 , \3605 );
xnor \U$3457 ( \3607 , \3606 , \487 );
xor \U$3458 ( \3608 , \3603 , \3607 );
and \U$3459 ( \3609 , \261 , \1301 );
and \U$3460 ( \3610 , \307 , \1246 );
nor \U$3461 ( \3611 , \3609 , \3610 );
xnor \U$3462 ( \3612 , \3611 , \1205 );
xor \U$3463 ( \3613 , \3608 , \3612 );
xor \U$3464 ( \3614 , \3599 , \3613 );
and \U$3465 ( \3615 , \178 , \1578 );
and \U$3466 ( \3616 , \185 , \1431 );
nor \U$3467 ( \3617 , \3615 , \3616 );
xnor \U$3468 ( \3618 , \3617 , \1436 );
and \U$3469 ( \3619 , \189 , \1824 );
and \U$3470 ( \3620 , \197 , \1739 );
nor \U$3471 ( \3621 , \3619 , \3620 );
xnor \U$3472 ( \3622 , \3621 , \1697 );
xor \U$3473 ( \3623 , \3618 , \3622 );
and \U$3474 ( \3624 , \209 , \2121 );
and \U$3475 ( \3625 , \217 , \2008 );
nor \U$3476 ( \3626 , \3624 , \3625 );
xnor \U$3477 ( \3627 , \3626 , \1961 );
xor \U$3478 ( \3628 , \3623 , \3627 );
xor \U$3479 ( \3629 , \3614 , \3628 );
xor \U$3480 ( \3630 , \3585 , \3629 );
and \U$3481 ( \3631 , \2757 , \215 );
and \U$3482 ( \3632 , \2826 , \213 );
nor \U$3483 ( \3633 , \3631 , \3632 );
xnor \U$3484 ( \3634 , \3633 , \222 );
and \U$3485 ( \3635 , \2366 , \230 );
and \U$3486 ( \3636 , \2521 , \228 );
nor \U$3487 ( \3637 , \3635 , \3636 );
xnor \U$3488 ( \3638 , \3637 , \237 );
xor \U$3489 ( \3639 , \3634 , \3638 );
and \U$3490 ( \3640 , \2090 , \245 );
and \U$3491 ( \3641 , \2182 , \243 );
nor \U$3492 ( \3642 , \3640 , \3641 );
xnor \U$3493 ( \3643 , \3642 , \252 );
xor \U$3494 ( \3644 , \3639 , \3643 );
and \U$3495 ( \3645 , \3395 , \183 );
buf \U$3496 ( \3646 , RIb55e518_92);
and \U$3497 ( \3647 , \3646 , \180 );
nor \U$3498 ( \3648 , \3645 , \3647 );
xnor \U$3499 ( \3649 , \3648 , \179 );
and \U$3500 ( \3650 , \3037 , \195 );
and \U$3501 ( \3651 , \3143 , \193 );
nor \U$3502 ( \3652 , \3650 , \3651 );
xnor \U$3503 ( \3653 , \3652 , \202 );
xor \U$3504 ( \3654 , \3649 , \3653 );
xor \U$3505 ( \3655 , \3654 , \3562 );
xor \U$3506 ( \3656 , \3644 , \3655 );
xor \U$3507 ( \3657 , \3630 , \3656 );
xor \U$3508 ( \3658 , \3581 , \3657 );
xor \U$3509 ( \3659 , \3508 , \3658 );
xor \U$3510 ( \3660 , \3499 , \3659 );
and \U$3511 ( \3661 , \3306 , \3307 );
and \U$3512 ( \3662 , \3307 , \3471 );
and \U$3513 ( \3663 , \3306 , \3471 );
or \U$3514 ( \3664 , \3661 , \3662 , \3663 );
xor \U$3515 ( \3665 , \3660 , \3664 );
and \U$3516 ( \3666 , \3472 , \3476 );
and \U$3517 ( \3667 , \3477 , \3480 );
or \U$3518 ( \3668 , \3666 , \3667 );
xor \U$3519 ( \3669 , \3665 , \3668 );
buf g5553_GF_PartitionCandidate( \3670_nG5553 , \3669 );
buf \U$3520 ( \3671 , \3670_nG5553 );
and \U$3521 ( \3672 , \3503 , \3507 );
and \U$3522 ( \3673 , \3507 , \3658 );
and \U$3523 ( \3674 , \3503 , \3658 );
or \U$3524 ( \3675 , \3672 , \3673 , \3674 );
and \U$3525 ( \3676 , \3491 , \3495 );
and \U$3526 ( \3677 , \3495 , \3497 );
and \U$3527 ( \3678 , \3491 , \3497 );
or \U$3528 ( \3679 , \3676 , \3677 , \3678 );
and \U$3529 ( \3680 , \3522 , \3580 );
and \U$3530 ( \3681 , \3580 , \3657 );
and \U$3531 ( \3682 , \3522 , \3657 );
or \U$3532 ( \3683 , \3680 , \3681 , \3682 );
xor \U$3533 ( \3684 , \3679 , \3683 );
and \U$3534 ( \3685 , \3526 , \3530 );
and \U$3535 ( \3686 , \3530 , \3535 );
and \U$3536 ( \3687 , \3526 , \3535 );
or \U$3537 ( \3688 , \3685 , \3686 , \3687 );
and \U$3538 ( \3689 , \3540 , \3544 );
and \U$3539 ( \3690 , \3544 , \3549 );
and \U$3540 ( \3691 , \3540 , \3549 );
or \U$3541 ( \3692 , \3689 , \3690 , \3691 );
xor \U$3542 ( \3693 , \3688 , \3692 );
and \U$3543 ( \3694 , \3555 , \3563 );
and \U$3544 ( \3695 , \3563 , \3578 );
and \U$3545 ( \3696 , \3555 , \3578 );
or \U$3546 ( \3697 , \3694 , \3695 , \3696 );
xor \U$3547 ( \3698 , \3693 , \3697 );
xor \U$3548 ( \3699 , \3684 , \3698 );
xor \U$3549 ( \3700 , \3675 , \3699 );
and \U$3550 ( \3701 , \3512 , \3516 );
and \U$3551 ( \3702 , \3516 , \3521 );
and \U$3552 ( \3703 , \3512 , \3521 );
or \U$3553 ( \3704 , \3701 , \3702 , \3703 );
and \U$3554 ( \3705 , \3536 , \3550 );
and \U$3555 ( \3706 , \3550 , \3579 );
and \U$3556 ( \3707 , \3536 , \3579 );
or \U$3557 ( \3708 , \3705 , \3706 , \3707 );
xor \U$3558 ( \3709 , \3704 , \3708 );
and \U$3559 ( \3710 , \3585 , \3629 );
and \U$3560 ( \3711 , \3629 , \3656 );
and \U$3561 ( \3712 , \3585 , \3656 );
or \U$3562 ( \3713 , \3710 , \3711 , \3712 );
xor \U$3563 ( \3714 , \3709 , \3713 );
and \U$3564 ( \3715 , \3589 , \3593 );
and \U$3565 ( \3716 , \3593 , \3598 );
and \U$3566 ( \3717 , \3589 , \3598 );
or \U$3567 ( \3718 , \3715 , \3716 , \3717 );
and \U$3568 ( \3719 , \3634 , \3638 );
and \U$3569 ( \3720 , \3638 , \3643 );
and \U$3570 ( \3721 , \3634 , \3643 );
or \U$3571 ( \3722 , \3719 , \3720 , \3721 );
xor \U$3572 ( \3723 , \3718 , \3722 );
and \U$3573 ( \3724 , \3649 , \3653 );
and \U$3574 ( \3725 , \3653 , \3562 );
and \U$3575 ( \3726 , \3649 , \3562 );
or \U$3576 ( \3727 , \3724 , \3725 , \3726 );
xor \U$3577 ( \3728 , \3723 , \3727 );
and \U$3578 ( \3729 , \3599 , \3613 );
and \U$3579 ( \3730 , \3613 , \3628 );
and \U$3580 ( \3731 , \3599 , \3628 );
or \U$3581 ( \3732 , \3729 , \3730 , \3731 );
and \U$3582 ( \3733 , \3644 , \3655 );
xor \U$3583 ( \3734 , \3732 , \3733 );
and \U$3584 ( \3735 , \3646 , \183 );
buf \U$3585 ( \3736 , RIb55e590_91);
and \U$3586 ( \3737 , \3736 , \180 );
nor \U$3587 ( \3738 , \3735 , \3737 );
xnor \U$3588 ( \3739 , \3738 , \179 );
and \U$3589 ( \3740 , \3143 , \195 );
and \U$3590 ( \3741 , \3395 , \193 );
nor \U$3591 ( \3742 , \3740 , \3741 );
xnor \U$3592 ( \3743 , \3742 , \202 );
xor \U$3593 ( \3744 , \3739 , \3743 );
and \U$3594 ( \3745 , \2826 , \215 );
and \U$3595 ( \3746 , \3037 , \213 );
nor \U$3596 ( \3747 , \3745 , \3746 );
xnor \U$3597 ( \3748 , \3747 , \222 );
xor \U$3598 ( \3749 , \3744 , \3748 );
xor \U$3599 ( \3750 , \3734 , \3749 );
xor \U$3600 ( \3751 , \3728 , \3750 );
and \U$3601 ( \3752 , \3568 , \3572 );
and \U$3602 ( \3753 , \3572 , \3577 );
and \U$3603 ( \3754 , \3568 , \3577 );
or \U$3604 ( \3755 , \3752 , \3753 , \3754 );
and \U$3605 ( \3756 , \3603 , \3607 );
and \U$3606 ( \3757 , \3607 , \3612 );
and \U$3607 ( \3758 , \3603 , \3612 );
or \U$3608 ( \3759 , \3756 , \3757 , \3758 );
xor \U$3609 ( \3760 , \3755 , \3759 );
and \U$3610 ( \3761 , \3618 , \3622 );
and \U$3611 ( \3762 , \3622 , \3627 );
and \U$3612 ( \3763 , \3618 , \3627 );
or \U$3613 ( \3764 , \3761 , \3762 , \3763 );
xor \U$3614 ( \3765 , \3760 , \3764 );
and \U$3615 ( \3766 , \1684 , \156 );
and \U$3616 ( \3767 , \1802 , \154 );
nor \U$3617 ( \3768 , \3766 , \3767 );
xnor \U$3618 ( \3769 , \3768 , \163 );
and \U$3619 ( \3770 , \1484 , \296 );
and \U$3620 ( \3771 , \1601 , \168 );
nor \U$3621 ( \3772 , \3770 , \3771 );
xnor \U$3622 ( \3773 , \3772 , \173 );
xor \U$3623 ( \3774 , \3769 , \3773 );
and \U$3624 ( \3775 , \1192 , \438 );
and \U$3625 ( \3776 , \1333 , \336 );
nor \U$3626 ( \3777 , \3775 , \3776 );
xnor \U$3627 ( \3778 , \3777 , \320 );
xor \U$3628 ( \3779 , \3774 , \3778 );
and \U$3629 ( \3780 , \474 , \1086 );
and \U$3630 ( \3781 , \1147 , \508 );
nor \U$3631 ( \3782 , \3780 , \3781 );
xnor \U$3632 ( \3783 , \3782 , \487 );
and \U$3633 ( \3784 , \307 , \1301 );
and \U$3634 ( \3785 , \412 , \1246 );
nor \U$3635 ( \3786 , \3784 , \3785 );
xnor \U$3636 ( \3787 , \3786 , \1205 );
xor \U$3637 ( \3788 , \3783 , \3787 );
and \U$3638 ( \3789 , \185 , \1578 );
and \U$3639 ( \3790 , \261 , \1431 );
nor \U$3640 ( \3791 , \3789 , \3790 );
xnor \U$3641 ( \3792 , \3791 , \1436 );
xor \U$3642 ( \3793 , \3788 , \3792 );
xor \U$3643 ( \3794 , \3779 , \3793 );
and \U$3644 ( \3795 , \2521 , \230 );
and \U$3645 ( \3796 , \2757 , \228 );
nor \U$3646 ( \3797 , \3795 , \3796 );
xnor \U$3647 ( \3798 , \3797 , \237 );
and \U$3648 ( \3799 , \2182 , \245 );
and \U$3649 ( \3800 , \2366 , \243 );
nor \U$3650 ( \3801 , \3799 , \3800 );
xnor \U$3651 ( \3802 , \3801 , \252 );
xor \U$3652 ( \3803 , \3798 , \3802 );
and \U$3653 ( \3804 , \1948 , \141 );
and \U$3654 ( \3805 , \2090 , \139 );
nor \U$3655 ( \3806 , \3804 , \3805 );
xnor \U$3656 ( \3807 , \3806 , \148 );
xor \U$3657 ( \3808 , \3803 , \3807 );
xor \U$3658 ( \3809 , \3794 , \3808 );
xor \U$3659 ( \3810 , \3765 , \3809 );
xor \U$3660 ( \3811 , \3559 , \3556 );
not \U$3661 ( \3812 , \3557 );
and \U$3662 ( \3813 , \3811 , \3812 );
and \U$3663 ( \3814 , \166 , \3813 );
and \U$3664 ( \3815 , \150 , \3557 );
nor \U$3665 ( \3816 , \3814 , \3815 );
xnor \U$3666 ( \3817 , \3816 , \3562 );
and \U$3667 ( \3818 , \247 , \2669 );
and \U$3668 ( \3819 , \224 , \2538 );
nor \U$3669 ( \3820 , \3818 , \3819 );
xnor \U$3670 ( \3821 , \3820 , \2534 );
and \U$3671 ( \3822 , \143 , \3103 );
and \U$3672 ( \3823 , \240 , \2934 );
nor \U$3673 ( \3824 , \3822 , \3823 );
xnor \U$3674 ( \3825 , \3824 , \2839 );
xor \U$3675 ( \3826 , \3821 , \3825 );
and \U$3676 ( \3827 , \158 , \3357 );
and \U$3677 ( \3828 , \134 , \3255 );
nor \U$3678 ( \3829 , \3827 , \3828 );
xnor \U$3679 ( \3830 , \3829 , \3156 );
xor \U$3680 ( \3831 , \3826 , \3830 );
xor \U$3681 ( \3832 , \3817 , \3831 );
and \U$3682 ( \3833 , \197 , \1824 );
and \U$3683 ( \3834 , \178 , \1739 );
nor \U$3684 ( \3835 , \3833 , \3834 );
xnor \U$3685 ( \3836 , \3835 , \1697 );
and \U$3686 ( \3837 , \217 , \2121 );
and \U$3687 ( \3838 , \189 , \2008 );
nor \U$3688 ( \3839 , \3837 , \3838 );
xnor \U$3689 ( \3840 , \3839 , \1961 );
xor \U$3690 ( \3841 , \3836 , \3840 );
and \U$3691 ( \3842 , \232 , \2400 );
and \U$3692 ( \3843 , \209 , \2246 );
nor \U$3693 ( \3844 , \3842 , \3843 );
xnor \U$3694 ( \3845 , \3844 , \2195 );
xor \U$3695 ( \3846 , \3841 , \3845 );
xor \U$3696 ( \3847 , \3832 , \3846 );
xor \U$3697 ( \3848 , \3810 , \3847 );
xor \U$3698 ( \3849 , \3751 , \3848 );
xor \U$3699 ( \3850 , \3714 , \3849 );
xor \U$3700 ( \3851 , \3700 , \3850 );
and \U$3701 ( \3852 , \3487 , \3498 );
and \U$3702 ( \3853 , \3498 , \3659 );
and \U$3703 ( \3854 , \3487 , \3659 );
or \U$3704 ( \3855 , \3852 , \3853 , \3854 );
xor \U$3705 ( \3856 , \3851 , \3855 );
and \U$3706 ( \3857 , \3660 , \3664 );
and \U$3707 ( \3858 , \3665 , \3668 );
or \U$3708 ( \3859 , \3857 , \3858 );
xor \U$3709 ( \3860 , \3856 , \3859 );
buf g5551_GF_PartitionCandidate( \3861_nG5551 , \3860 );
buf \U$3710 ( \3862 , \3861_nG5551 );
and \U$3711 ( \3863 , \3679 , \3683 );
and \U$3712 ( \3864 , \3683 , \3698 );
and \U$3713 ( \3865 , \3679 , \3698 );
or \U$3714 ( \3866 , \3863 , \3864 , \3865 );
and \U$3715 ( \3867 , \3714 , \3849 );
xor \U$3716 ( \3868 , \3866 , \3867 );
and \U$3717 ( \3869 , \3688 , \3692 );
and \U$3718 ( \3870 , \3692 , \3697 );
and \U$3719 ( \3871 , \3688 , \3697 );
or \U$3720 ( \3872 , \3869 , \3870 , \3871 );
and \U$3721 ( \3873 , \3732 , \3733 );
and \U$3722 ( \3874 , \3733 , \3749 );
and \U$3723 ( \3875 , \3732 , \3749 );
or \U$3724 ( \3876 , \3873 , \3874 , \3875 );
xor \U$3725 ( \3877 , \3872 , \3876 );
and \U$3726 ( \3878 , \3765 , \3809 );
and \U$3727 ( \3879 , \3809 , \3847 );
and \U$3728 ( \3880 , \3765 , \3847 );
or \U$3729 ( \3881 , \3878 , \3879 , \3880 );
xor \U$3730 ( \3882 , \3877 , \3881 );
xor \U$3731 ( \3883 , \3868 , \3882 );
and \U$3732 ( \3884 , \3704 , \3708 );
and \U$3733 ( \3885 , \3708 , \3713 );
and \U$3734 ( \3886 , \3704 , \3713 );
or \U$3735 ( \3887 , \3884 , \3885 , \3886 );
and \U$3736 ( \3888 , \3728 , \3750 );
and \U$3737 ( \3889 , \3750 , \3848 );
and \U$3738 ( \3890 , \3728 , \3848 );
or \U$3739 ( \3891 , \3888 , \3889 , \3890 );
xor \U$3740 ( \3892 , \3887 , \3891 );
and \U$3741 ( \3893 , \3718 , \3722 );
and \U$3742 ( \3894 , \3722 , \3727 );
and \U$3743 ( \3895 , \3718 , \3727 );
or \U$3744 ( \3896 , \3893 , \3894 , \3895 );
and \U$3745 ( \3897 , \3755 , \3759 );
and \U$3746 ( \3898 , \3759 , \3764 );
and \U$3747 ( \3899 , \3755 , \3764 );
or \U$3748 ( \3900 , \3897 , \3898 , \3899 );
xor \U$3749 ( \3901 , \3896 , \3900 );
and \U$3750 ( \3902 , \3817 , \3831 );
and \U$3751 ( \3903 , \3831 , \3846 );
and \U$3752 ( \3904 , \3817 , \3846 );
or \U$3753 ( \3905 , \3902 , \3903 , \3904 );
xor \U$3754 ( \3906 , \3901 , \3905 );
and \U$3755 ( \3907 , \3779 , \3793 );
and \U$3756 ( \3908 , \3793 , \3808 );
and \U$3757 ( \3909 , \3779 , \3808 );
or \U$3758 ( \3910 , \3907 , \3908 , \3909 );
and \U$3759 ( \3911 , \3736 , \183 );
buf \U$3760 ( \3912 , RIb55e608_90);
and \U$3761 ( \3913 , \3912 , \180 );
nor \U$3762 ( \3914 , \3911 , \3913 );
xnor \U$3763 ( \3915 , \3914 , \179 );
and \U$3764 ( \3916 , \3395 , \195 );
and \U$3765 ( \3917 , \3646 , \193 );
nor \U$3766 ( \3918 , \3916 , \3917 );
xnor \U$3767 ( \3919 , \3918 , \202 );
xor \U$3768 ( \3920 , \3915 , \3919 );
buf \U$3769 ( \3921 , RIb560480_25);
buf \U$3770 ( \3922 , RIb560408_26);
and \U$3771 ( \3923 , \3922 , \3559 );
not \U$3772 ( \3924 , \3923 );
and \U$3773 ( \3925 , \3921 , \3924 );
xor \U$3774 ( \3926 , \3920 , \3925 );
xor \U$3775 ( \3927 , \3910 , \3926 );
and \U$3776 ( \3928 , \1333 , \438 );
and \U$3777 ( \3929 , \1484 , \336 );
nor \U$3778 ( \3930 , \3928 , \3929 );
xnor \U$3779 ( \3931 , \3930 , \320 );
and \U$3780 ( \3932 , \1147 , \1086 );
and \U$3781 ( \3933 , \1192 , \508 );
nor \U$3782 ( \3934 , \3932 , \3933 );
xnor \U$3783 ( \3935 , \3934 , \487 );
xor \U$3784 ( \3936 , \3931 , \3935 );
and \U$3785 ( \3937 , \412 , \1301 );
and \U$3786 ( \3938 , \474 , \1246 );
nor \U$3787 ( \3939 , \3937 , \3938 );
xnor \U$3788 ( \3940 , \3939 , \1205 );
xor \U$3789 ( \3941 , \3936 , \3940 );
and \U$3790 ( \3942 , \2090 , \141 );
and \U$3791 ( \3943 , \2182 , \139 );
nor \U$3792 ( \3944 , \3942 , \3943 );
xnor \U$3793 ( \3945 , \3944 , \148 );
and \U$3794 ( \3946 , \1802 , \156 );
and \U$3795 ( \3947 , \1948 , \154 );
nor \U$3796 ( \3948 , \3946 , \3947 );
xnor \U$3797 ( \3949 , \3948 , \163 );
xor \U$3798 ( \3950 , \3945 , \3949 );
and \U$3799 ( \3951 , \1601 , \296 );
and \U$3800 ( \3952 , \1684 , \168 );
nor \U$3801 ( \3953 , \3951 , \3952 );
xnor \U$3802 ( \3954 , \3953 , \173 );
xor \U$3803 ( \3955 , \3950 , \3954 );
xor \U$3804 ( \3956 , \3941 , \3955 );
and \U$3805 ( \3957 , \3037 , \215 );
and \U$3806 ( \3958 , \3143 , \213 );
nor \U$3807 ( \3959 , \3957 , \3958 );
xnor \U$3808 ( \3960 , \3959 , \222 );
and \U$3809 ( \3961 , \2757 , \230 );
and \U$3810 ( \3962 , \2826 , \228 );
nor \U$3811 ( \3963 , \3961 , \3962 );
xnor \U$3812 ( \3964 , \3963 , \237 );
xor \U$3813 ( \3965 , \3960 , \3964 );
and \U$3814 ( \3966 , \2366 , \245 );
and \U$3815 ( \3967 , \2521 , \243 );
nor \U$3816 ( \3968 , \3966 , \3967 );
xnor \U$3817 ( \3969 , \3968 , \252 );
xor \U$3818 ( \3970 , \3965 , \3969 );
xor \U$3819 ( \3971 , \3956 , \3970 );
xor \U$3820 ( \3972 , \3927 , \3971 );
xor \U$3821 ( \3973 , \3906 , \3972 );
and \U$3822 ( \3974 , \3821 , \3825 );
and \U$3823 ( \3975 , \3825 , \3830 );
and \U$3824 ( \3976 , \3821 , \3830 );
or \U$3825 ( \3977 , \3974 , \3975 , \3976 );
and \U$3826 ( \3978 , \3783 , \3787 );
and \U$3827 ( \3979 , \3787 , \3792 );
and \U$3828 ( \3980 , \3783 , \3792 );
or \U$3829 ( \3981 , \3978 , \3979 , \3980 );
xor \U$3830 ( \3982 , \3977 , \3981 );
and \U$3831 ( \3983 , \3836 , \3840 );
and \U$3832 ( \3984 , \3840 , \3845 );
and \U$3833 ( \3985 , \3836 , \3845 );
or \U$3834 ( \3986 , \3983 , \3984 , \3985 );
xor \U$3835 ( \3987 , \3982 , \3986 );
and \U$3836 ( \3988 , \3769 , \3773 );
and \U$3837 ( \3989 , \3773 , \3778 );
and \U$3838 ( \3990 , \3769 , \3778 );
or \U$3839 ( \3991 , \3988 , \3989 , \3990 );
and \U$3840 ( \3992 , \3798 , \3802 );
and \U$3841 ( \3993 , \3802 , \3807 );
and \U$3842 ( \3994 , \3798 , \3807 );
or \U$3843 ( \3995 , \3992 , \3993 , \3994 );
xor \U$3844 ( \3996 , \3991 , \3995 );
and \U$3845 ( \3997 , \3739 , \3743 );
and \U$3846 ( \3998 , \3743 , \3748 );
and \U$3847 ( \3999 , \3739 , \3748 );
or \U$3848 ( \4000 , \3997 , \3998 , \3999 );
xor \U$3849 ( \4001 , \3996 , \4000 );
xor \U$3850 ( \4002 , \3987 , \4001 );
and \U$3851 ( \4003 , \134 , \3357 );
and \U$3852 ( \4004 , \143 , \3255 );
nor \U$3853 ( \4005 , \4003 , \4004 );
xnor \U$3854 ( \4006 , \4005 , \3156 );
and \U$3855 ( \4007 , \150 , \3813 );
and \U$3856 ( \4008 , \158 , \3557 );
nor \U$3857 ( \4009 , \4007 , \4008 );
xnor \U$3858 ( \4010 , \4009 , \3562 );
xor \U$3859 ( \4011 , \4006 , \4010 );
xor \U$3860 ( \4012 , \3922 , \3559 );
nand \U$3861 ( \4013 , \166 , \4012 );
xnor \U$3862 ( \4014 , \4013 , \3925 );
xor \U$3863 ( \4015 , \4011 , \4014 );
and \U$3864 ( \4016 , \209 , \2400 );
and \U$3865 ( \4017 , \217 , \2246 );
nor \U$3866 ( \4018 , \4016 , \4017 );
xnor \U$3867 ( \4019 , \4018 , \2195 );
and \U$3868 ( \4020 , \224 , \2669 );
and \U$3869 ( \4021 , \232 , \2538 );
nor \U$3870 ( \4022 , \4020 , \4021 );
xnor \U$3871 ( \4023 , \4022 , \2534 );
xor \U$3872 ( \4024 , \4019 , \4023 );
and \U$3873 ( \4025 , \240 , \3103 );
and \U$3874 ( \4026 , \247 , \2934 );
nor \U$3875 ( \4027 , \4025 , \4026 );
xnor \U$3876 ( \4028 , \4027 , \2839 );
xor \U$3877 ( \4029 , \4024 , \4028 );
xor \U$3878 ( \4030 , \4015 , \4029 );
and \U$3879 ( \4031 , \261 , \1578 );
and \U$3880 ( \4032 , \307 , \1431 );
nor \U$3881 ( \4033 , \4031 , \4032 );
xnor \U$3882 ( \4034 , \4033 , \1436 );
and \U$3883 ( \4035 , \178 , \1824 );
and \U$3884 ( \4036 , \185 , \1739 );
nor \U$3885 ( \4037 , \4035 , \4036 );
xnor \U$3886 ( \4038 , \4037 , \1697 );
xor \U$3887 ( \4039 , \4034 , \4038 );
and \U$3888 ( \4040 , \189 , \2121 );
and \U$3889 ( \4041 , \197 , \2008 );
nor \U$3890 ( \4042 , \4040 , \4041 );
xnor \U$3891 ( \4043 , \4042 , \1961 );
xor \U$3892 ( \4044 , \4039 , \4043 );
xor \U$3893 ( \4045 , \4030 , \4044 );
xor \U$3894 ( \4046 , \4002 , \4045 );
xor \U$3895 ( \4047 , \3973 , \4046 );
xor \U$3896 ( \4048 , \3892 , \4047 );
xor \U$3897 ( \4049 , \3883 , \4048 );
and \U$3898 ( \4050 , \3675 , \3699 );
and \U$3899 ( \4051 , \3699 , \3850 );
and \U$3900 ( \4052 , \3675 , \3850 );
or \U$3901 ( \4053 , \4050 , \4051 , \4052 );
xor \U$3902 ( \4054 , \4049 , \4053 );
and \U$3903 ( \4055 , \3851 , \3855 );
and \U$3904 ( \4056 , \3856 , \3859 );
or \U$3905 ( \4057 , \4055 , \4056 );
xor \U$3906 ( \4058 , \4054 , \4057 );
buf g554f_GF_PartitionCandidate( \4059_nG554f , \4058 );
buf \U$3907 ( \4060 , \4059_nG554f );
and \U$3908 ( \4061 , \3866 , \3867 );
and \U$3909 ( \4062 , \3867 , \3882 );
and \U$3910 ( \4063 , \3866 , \3882 );
or \U$3911 ( \4064 , \4061 , \4062 , \4063 );
and \U$3912 ( \4065 , \3887 , \3891 );
and \U$3913 ( \4066 , \3891 , \4047 );
and \U$3914 ( \4067 , \3887 , \4047 );
or \U$3915 ( \4068 , \4065 , \4066 , \4067 );
and \U$3916 ( \4069 , \3896 , \3900 );
and \U$3917 ( \4070 , \3900 , \3905 );
and \U$3918 ( \4071 , \3896 , \3905 );
or \U$3919 ( \4072 , \4069 , \4070 , \4071 );
and \U$3920 ( \4073 , \3910 , \3926 );
and \U$3921 ( \4074 , \3926 , \3971 );
and \U$3922 ( \4075 , \3910 , \3971 );
or \U$3923 ( \4076 , \4073 , \4074 , \4075 );
xor \U$3924 ( \4077 , \4072 , \4076 );
and \U$3925 ( \4078 , \3987 , \4001 );
and \U$3926 ( \4079 , \4001 , \4045 );
and \U$3927 ( \4080 , \3987 , \4045 );
or \U$3928 ( \4081 , \4078 , \4079 , \4080 );
xor \U$3929 ( \4082 , \4077 , \4081 );
xor \U$3930 ( \4083 , \4068 , \4082 );
and \U$3931 ( \4084 , \3872 , \3876 );
and \U$3932 ( \4085 , \3876 , \3881 );
and \U$3933 ( \4086 , \3872 , \3881 );
or \U$3934 ( \4087 , \4084 , \4085 , \4086 );
and \U$3935 ( \4088 , \3906 , \3972 );
and \U$3936 ( \4089 , \3972 , \4046 );
and \U$3937 ( \4090 , \3906 , \4046 );
or \U$3938 ( \4091 , \4088 , \4089 , \4090 );
xor \U$3939 ( \4092 , \4087 , \4091 );
and \U$3940 ( \4093 , \3977 , \3981 );
and \U$3941 ( \4094 , \3981 , \3986 );
and \U$3942 ( \4095 , \3977 , \3986 );
or \U$3943 ( \4096 , \4093 , \4094 , \4095 );
and \U$3944 ( \4097 , \3991 , \3995 );
and \U$3945 ( \4098 , \3995 , \4000 );
and \U$3946 ( \4099 , \3991 , \4000 );
or \U$3947 ( \4100 , \4097 , \4098 , \4099 );
xor \U$3948 ( \4101 , \4096 , \4100 );
and \U$3949 ( \4102 , \4015 , \4029 );
and \U$3950 ( \4103 , \4029 , \4044 );
and \U$3951 ( \4104 , \4015 , \4044 );
or \U$3952 ( \4105 , \4102 , \4103 , \4104 );
xor \U$3953 ( \4106 , \4101 , \4105 );
and \U$3954 ( \4107 , \3915 , \3919 );
and \U$3955 ( \4108 , \3919 , \3925 );
and \U$3956 ( \4109 , \3915 , \3925 );
or \U$3957 ( \4110 , \4107 , \4108 , \4109 );
and \U$3958 ( \4111 , \3945 , \3949 );
and \U$3959 ( \4112 , \3949 , \3954 );
and \U$3960 ( \4113 , \3945 , \3954 );
or \U$3961 ( \4114 , \4111 , \4112 , \4113 );
xor \U$3962 ( \4115 , \4110 , \4114 );
and \U$3963 ( \4116 , \3960 , \3964 );
and \U$3964 ( \4117 , \3964 , \3969 );
and \U$3965 ( \4118 , \3960 , \3969 );
or \U$3966 ( \4119 , \4116 , \4117 , \4118 );
xor \U$3967 ( \4120 , \4115 , \4119 );
and \U$3968 ( \4121 , \4006 , \4010 );
and \U$3969 ( \4122 , \4010 , \4014 );
and \U$3970 ( \4123 , \4006 , \4014 );
or \U$3971 ( \4124 , \4121 , \4122 , \4123 );
and \U$3972 ( \4125 , \158 , \3813 );
and \U$3973 ( \4126 , \134 , \3557 );
nor \U$3974 ( \4127 , \4125 , \4126 );
xnor \U$3975 ( \4128 , \4127 , \3562 );
xor \U$3976 ( \4129 , \4124 , \4128 );
xor \U$3977 ( \4130 , \3921 , \3922 );
not \U$3978 ( \4131 , \4012 );
and \U$3979 ( \4132 , \4130 , \4131 );
and \U$3980 ( \4133 , \166 , \4132 );
and \U$3981 ( \4134 , \150 , \4012 );
nor \U$3982 ( \4135 , \4133 , \4134 );
xnor \U$3983 ( \4136 , \4135 , \3925 );
xor \U$3984 ( \4137 , \4129 , \4136 );
xor \U$3985 ( \4138 , \4120 , \4137 );
and \U$3986 ( \4139 , \3931 , \3935 );
and \U$3987 ( \4140 , \3935 , \3940 );
and \U$3988 ( \4141 , \3931 , \3940 );
or \U$3989 ( \4142 , \4139 , \4140 , \4141 );
and \U$3990 ( \4143 , \4019 , \4023 );
and \U$3991 ( \4144 , \4023 , \4028 );
and \U$3992 ( \4145 , \4019 , \4028 );
or \U$3993 ( \4146 , \4143 , \4144 , \4145 );
xor \U$3994 ( \4147 , \4142 , \4146 );
and \U$3995 ( \4148 , \4034 , \4038 );
and \U$3996 ( \4149 , \4038 , \4043 );
and \U$3997 ( \4150 , \4034 , \4043 );
or \U$3998 ( \4151 , \4148 , \4149 , \4150 );
xor \U$3999 ( \4152 , \4147 , \4151 );
xor \U$4000 ( \4153 , \4138 , \4152 );
xor \U$4001 ( \4154 , \4106 , \4153 );
and \U$4002 ( \4155 , \3941 , \3955 );
and \U$4003 ( \4156 , \3955 , \3970 );
and \U$4004 ( \4157 , \3941 , \3970 );
or \U$4005 ( \4158 , \4155 , \4156 , \4157 );
and \U$4006 ( \4159 , \3912 , \183 );
buf \U$4007 ( \4160 , RIb55e680_89);
and \U$4008 ( \4161 , \4160 , \180 );
nor \U$4009 ( \4162 , \4159 , \4161 );
xnor \U$4010 ( \4163 , \4162 , \179 );
and \U$4011 ( \4164 , \3646 , \195 );
and \U$4012 ( \4165 , \3736 , \193 );
nor \U$4013 ( \4166 , \4164 , \4165 );
xnor \U$4014 ( \4167 , \4166 , \202 );
xor \U$4015 ( \4168 , \4163 , \4167 );
and \U$4016 ( \4169 , \3143 , \215 );
and \U$4017 ( \4170 , \3395 , \213 );
nor \U$4018 ( \4171 , \4169 , \4170 );
xnor \U$4019 ( \4172 , \4171 , \222 );
xor \U$4020 ( \4173 , \4168 , \4172 );
and \U$4021 ( \4174 , \2826 , \230 );
and \U$4022 ( \4175 , \3037 , \228 );
nor \U$4023 ( \4176 , \4174 , \4175 );
xnor \U$4024 ( \4177 , \4176 , \237 );
and \U$4025 ( \4178 , \2521 , \245 );
and \U$4026 ( \4179 , \2757 , \243 );
nor \U$4027 ( \4180 , \4178 , \4179 );
xnor \U$4028 ( \4181 , \4180 , \252 );
xor \U$4029 ( \4182 , \4177 , \4181 );
and \U$4030 ( \4183 , \2182 , \141 );
and \U$4031 ( \4184 , \2366 , \139 );
nor \U$4032 ( \4185 , \4183 , \4184 );
xnor \U$4033 ( \4186 , \4185 , \148 );
xor \U$4034 ( \4187 , \4182 , \4186 );
xor \U$4035 ( \4188 , \4173 , \4187 );
and \U$4036 ( \4189 , \1948 , \156 );
and \U$4037 ( \4190 , \2090 , \154 );
nor \U$4038 ( \4191 , \4189 , \4190 );
xnor \U$4039 ( \4192 , \4191 , \163 );
and \U$4040 ( \4193 , \1684 , \296 );
and \U$4041 ( \4194 , \1802 , \168 );
nor \U$4042 ( \4195 , \4193 , \4194 );
xnor \U$4043 ( \4196 , \4195 , \173 );
xor \U$4044 ( \4197 , \4192 , \4196 );
and \U$4045 ( \4198 , \1484 , \438 );
and \U$4046 ( \4199 , \1601 , \336 );
nor \U$4047 ( \4200 , \4198 , \4199 );
xnor \U$4048 ( \4201 , \4200 , \320 );
xor \U$4049 ( \4202 , \4197 , \4201 );
xor \U$4050 ( \4203 , \4188 , \4202 );
xor \U$4051 ( \4204 , \4158 , \4203 );
and \U$4052 ( \4205 , \185 , \1824 );
and \U$4053 ( \4206 , \261 , \1739 );
nor \U$4054 ( \4207 , \4205 , \4206 );
xnor \U$4055 ( \4208 , \4207 , \1697 );
and \U$4056 ( \4209 , \197 , \2121 );
and \U$4057 ( \4210 , \178 , \2008 );
nor \U$4058 ( \4211 , \4209 , \4210 );
xnor \U$4059 ( \4212 , \4211 , \1961 );
xor \U$4060 ( \4213 , \4208 , \4212 );
and \U$4061 ( \4214 , \217 , \2400 );
and \U$4062 ( \4215 , \189 , \2246 );
nor \U$4063 ( \4216 , \4214 , \4215 );
xnor \U$4064 ( \4217 , \4216 , \2195 );
xor \U$4065 ( \4218 , \4213 , \4217 );
and \U$4066 ( \4219 , \1192 , \1086 );
and \U$4067 ( \4220 , \1333 , \508 );
nor \U$4068 ( \4221 , \4219 , \4220 );
xnor \U$4069 ( \4222 , \4221 , \487 );
and \U$4070 ( \4223 , \474 , \1301 );
and \U$4071 ( \4224 , \1147 , \1246 );
nor \U$4072 ( \4225 , \4223 , \4224 );
xnor \U$4073 ( \4226 , \4225 , \1205 );
xor \U$4074 ( \4227 , \4222 , \4226 );
and \U$4075 ( \4228 , \307 , \1578 );
and \U$4076 ( \4229 , \412 , \1431 );
nor \U$4077 ( \4230 , \4228 , \4229 );
xnor \U$4078 ( \4231 , \4230 , \1436 );
xor \U$4079 ( \4232 , \4227 , \4231 );
xor \U$4080 ( \4233 , \4218 , \4232 );
and \U$4081 ( \4234 , \232 , \2669 );
and \U$4082 ( \4235 , \209 , \2538 );
nor \U$4083 ( \4236 , \4234 , \4235 );
xnor \U$4084 ( \4237 , \4236 , \2534 );
and \U$4085 ( \4238 , \247 , \3103 );
and \U$4086 ( \4239 , \224 , \2934 );
nor \U$4087 ( \4240 , \4238 , \4239 );
xnor \U$4088 ( \4241 , \4240 , \2839 );
xor \U$4089 ( \4242 , \4237 , \4241 );
and \U$4090 ( \4243 , \143 , \3357 );
and \U$4091 ( \4244 , \240 , \3255 );
nor \U$4092 ( \4245 , \4243 , \4244 );
xnor \U$4093 ( \4246 , \4245 , \3156 );
xor \U$4094 ( \4247 , \4242 , \4246 );
xor \U$4095 ( \4248 , \4233 , \4247 );
xor \U$4096 ( \4249 , \4204 , \4248 );
xor \U$4097 ( \4250 , \4154 , \4249 );
xor \U$4098 ( \4251 , \4092 , \4250 );
xor \U$4099 ( \4252 , \4083 , \4251 );
xor \U$4100 ( \4253 , \4064 , \4252 );
and \U$4101 ( \4254 , \3883 , \4048 );
xor \U$4102 ( \4255 , \4253 , \4254 );
and \U$4103 ( \4256 , \4049 , \4053 );
and \U$4104 ( \4257 , \4054 , \4057 );
or \U$4105 ( \4258 , \4256 , \4257 );
xor \U$4106 ( \4259 , \4255 , \4258 );
buf g554d_GF_PartitionCandidate( \4260_nG554d , \4259 );
buf \U$4107 ( \4261 , \4260_nG554d );
and \U$4108 ( \4262 , \4068 , \4082 );
and \U$4109 ( \4263 , \4082 , \4251 );
and \U$4110 ( \4264 , \4068 , \4251 );
or \U$4111 ( \4265 , \4262 , \4263 , \4264 );
and \U$4112 ( \4266 , \4087 , \4091 );
and \U$4113 ( \4267 , \4091 , \4250 );
and \U$4114 ( \4268 , \4087 , \4250 );
or \U$4115 ( \4269 , \4266 , \4267 , \4268 );
and \U$4116 ( \4270 , \4072 , \4076 );
and \U$4117 ( \4271 , \4076 , \4081 );
and \U$4118 ( \4272 , \4072 , \4081 );
or \U$4119 ( \4273 , \4270 , \4271 , \4272 );
and \U$4120 ( \4274 , \4106 , \4153 );
and \U$4121 ( \4275 , \4153 , \4249 );
and \U$4122 ( \4276 , \4106 , \4249 );
or \U$4123 ( \4277 , \4274 , \4275 , \4276 );
xor \U$4124 ( \4278 , \4273 , \4277 );
and \U$4125 ( \4279 , \4173 , \4187 );
and \U$4126 ( \4280 , \4187 , \4202 );
and \U$4127 ( \4281 , \4173 , \4202 );
or \U$4128 ( \4282 , \4279 , \4280 , \4281 );
and \U$4129 ( \4283 , \4218 , \4232 );
and \U$4130 ( \4284 , \4232 , \4247 );
and \U$4131 ( \4285 , \4218 , \4247 );
or \U$4132 ( \4286 , \4283 , \4284 , \4285 );
xor \U$4133 ( \4287 , \4282 , \4286 );
and \U$4134 ( \4288 , \3395 , \215 );
and \U$4135 ( \4289 , \3646 , \213 );
nor \U$4136 ( \4290 , \4288 , \4289 );
xnor \U$4137 ( \4291 , \4290 , \222 );
and \U$4138 ( \4292 , \3037 , \230 );
and \U$4139 ( \4293 , \3143 , \228 );
nor \U$4140 ( \4294 , \4292 , \4293 );
xnor \U$4141 ( \4295 , \4294 , \237 );
xor \U$4142 ( \4296 , \4291 , \4295 );
and \U$4143 ( \4297 , \2757 , \245 );
and \U$4144 ( \4298 , \2826 , \243 );
nor \U$4145 ( \4299 , \4297 , \4298 );
xnor \U$4146 ( \4300 , \4299 , \252 );
xor \U$4147 ( \4301 , \4296 , \4300 );
xor \U$4148 ( \4302 , \4287 , \4301 );
xor \U$4149 ( \4303 , \4278 , \4302 );
xor \U$4150 ( \4304 , \4269 , \4303 );
and \U$4151 ( \4305 , \4110 , \4114 );
and \U$4152 ( \4306 , \4114 , \4119 );
and \U$4153 ( \4307 , \4110 , \4119 );
or \U$4154 ( \4308 , \4305 , \4306 , \4307 );
and \U$4155 ( \4309 , \4124 , \4128 );
and \U$4156 ( \4310 , \4128 , \4136 );
and \U$4157 ( \4311 , \4124 , \4136 );
or \U$4158 ( \4312 , \4309 , \4310 , \4311 );
xor \U$4159 ( \4313 , \4308 , \4312 );
and \U$4160 ( \4314 , \4142 , \4146 );
and \U$4161 ( \4315 , \4146 , \4151 );
and \U$4162 ( \4316 , \4142 , \4151 );
or \U$4163 ( \4317 , \4314 , \4315 , \4316 );
xor \U$4164 ( \4318 , \4313 , \4317 );
and \U$4165 ( \4319 , \4096 , \4100 );
and \U$4166 ( \4320 , \4100 , \4105 );
and \U$4167 ( \4321 , \4096 , \4105 );
or \U$4168 ( \4322 , \4319 , \4320 , \4321 );
and \U$4169 ( \4323 , \4120 , \4137 );
and \U$4170 ( \4324 , \4137 , \4152 );
and \U$4171 ( \4325 , \4120 , \4152 );
or \U$4172 ( \4326 , \4323 , \4324 , \4325 );
xor \U$4173 ( \4327 , \4322 , \4326 );
and \U$4174 ( \4328 , \4158 , \4203 );
and \U$4175 ( \4329 , \4203 , \4248 );
and \U$4176 ( \4330 , \4158 , \4248 );
or \U$4177 ( \4331 , \4328 , \4329 , \4330 );
xor \U$4178 ( \4332 , \4327 , \4331 );
xor \U$4179 ( \4333 , \4318 , \4332 );
and \U$4180 ( \4334 , \4163 , \4167 );
and \U$4181 ( \4335 , \4167 , \4172 );
and \U$4182 ( \4336 , \4163 , \4172 );
or \U$4183 ( \4337 , \4334 , \4335 , \4336 );
and \U$4184 ( \4338 , \4177 , \4181 );
and \U$4185 ( \4339 , \4181 , \4186 );
and \U$4186 ( \4340 , \4177 , \4186 );
or \U$4187 ( \4341 , \4338 , \4339 , \4340 );
xor \U$4188 ( \4342 , \4337 , \4341 );
and \U$4189 ( \4343 , \4192 , \4196 );
and \U$4190 ( \4344 , \4196 , \4201 );
and \U$4191 ( \4345 , \4192 , \4201 );
or \U$4192 ( \4346 , \4343 , \4344 , \4345 );
xor \U$4193 ( \4347 , \4342 , \4346 );
and \U$4194 ( \4348 , \4208 , \4212 );
and \U$4195 ( \4349 , \4212 , \4217 );
and \U$4196 ( \4350 , \4208 , \4217 );
or \U$4197 ( \4351 , \4348 , \4349 , \4350 );
and \U$4198 ( \4352 , \4222 , \4226 );
and \U$4199 ( \4353 , \4226 , \4231 );
and \U$4200 ( \4354 , \4222 , \4231 );
or \U$4201 ( \4355 , \4352 , \4353 , \4354 );
xor \U$4202 ( \4356 , \4351 , \4355 );
and \U$4203 ( \4357 , \4237 , \4241 );
and \U$4204 ( \4358 , \4241 , \4246 );
and \U$4205 ( \4359 , \4237 , \4246 );
or \U$4206 ( \4360 , \4357 , \4358 , \4359 );
xor \U$4207 ( \4361 , \4356 , \4360 );
xor \U$4208 ( \4362 , \4347 , \4361 );
and \U$4209 ( \4363 , \4160 , \183 );
buf \U$4210 ( \4364 , RIb55e6f8_88);
and \U$4211 ( \4365 , \4364 , \180 );
nor \U$4212 ( \4366 , \4363 , \4365 );
xnor \U$4213 ( \4367 , \4366 , \179 );
and \U$4214 ( \4368 , \3736 , \195 );
and \U$4215 ( \4369 , \3912 , \193 );
nor \U$4216 ( \4370 , \4368 , \4369 );
xnor \U$4217 ( \4371 , \4370 , \202 );
xor \U$4218 ( \4372 , \4367 , \4371 );
buf \U$4219 ( \4373 , RIb560570_23);
buf \U$4220 ( \4374 , RIb5604f8_24);
and \U$4221 ( \4375 , \4374 , \3921 );
not \U$4222 ( \4376 , \4375 );
and \U$4223 ( \4377 , \4373 , \4376 );
xor \U$4224 ( \4378 , \4372 , \4377 );
and \U$4225 ( \4379 , \2366 , \141 );
and \U$4226 ( \4380 , \2521 , \139 );
nor \U$4227 ( \4381 , \4379 , \4380 );
xnor \U$4228 ( \4382 , \4381 , \148 );
and \U$4229 ( \4383 , \2090 , \156 );
and \U$4230 ( \4384 , \2182 , \154 );
nor \U$4231 ( \4385 , \4383 , \4384 );
xnor \U$4232 ( \4386 , \4385 , \163 );
xor \U$4233 ( \4387 , \4382 , \4386 );
and \U$4234 ( \4388 , \1802 , \296 );
and \U$4235 ( \4389 , \1948 , \168 );
nor \U$4236 ( \4390 , \4388 , \4389 );
xnor \U$4237 ( \4391 , \4390 , \173 );
xor \U$4238 ( \4392 , \4387 , \4391 );
and \U$4239 ( \4393 , \1601 , \438 );
and \U$4240 ( \4394 , \1684 , \336 );
nor \U$4241 ( \4395 , \4393 , \4394 );
xnor \U$4242 ( \4396 , \4395 , \320 );
and \U$4243 ( \4397 , \1333 , \1086 );
and \U$4244 ( \4398 , \1484 , \508 );
nor \U$4245 ( \4399 , \4397 , \4398 );
xnor \U$4246 ( \4400 , \4399 , \487 );
xor \U$4247 ( \4401 , \4396 , \4400 );
and \U$4248 ( \4402 , \1147 , \1301 );
and \U$4249 ( \4403 , \1192 , \1246 );
nor \U$4250 ( \4404 , \4402 , \4403 );
xnor \U$4251 ( \4405 , \4404 , \1205 );
xor \U$4252 ( \4406 , \4401 , \4405 );
xor \U$4253 ( \4407 , \4392 , \4406 );
and \U$4254 ( \4408 , \412 , \1578 );
and \U$4255 ( \4409 , \474 , \1431 );
nor \U$4256 ( \4410 , \4408 , \4409 );
xnor \U$4257 ( \4411 , \4410 , \1436 );
and \U$4258 ( \4412 , \261 , \1824 );
and \U$4259 ( \4413 , \307 , \1739 );
nor \U$4260 ( \4414 , \4412 , \4413 );
xnor \U$4261 ( \4415 , \4414 , \1697 );
xor \U$4262 ( \4416 , \4411 , \4415 );
and \U$4263 ( \4417 , \178 , \2121 );
and \U$4264 ( \4418 , \185 , \2008 );
nor \U$4265 ( \4419 , \4417 , \4418 );
xnor \U$4266 ( \4420 , \4419 , \1961 );
xor \U$4267 ( \4421 , \4416 , \4420 );
xor \U$4268 ( \4422 , \4407 , \4421 );
xor \U$4269 ( \4423 , \4378 , \4422 );
xor \U$4270 ( \4424 , \4374 , \3921 );
nand \U$4271 ( \4425 , \166 , \4424 );
xnor \U$4272 ( \4426 , \4425 , \4377 );
and \U$4273 ( \4427 , \189 , \2400 );
and \U$4274 ( \4428 , \197 , \2246 );
nor \U$4275 ( \4429 , \4427 , \4428 );
xnor \U$4276 ( \4430 , \4429 , \2195 );
and \U$4277 ( \4431 , \209 , \2669 );
and \U$4278 ( \4432 , \217 , \2538 );
nor \U$4279 ( \4433 , \4431 , \4432 );
xnor \U$4280 ( \4434 , \4433 , \2534 );
xor \U$4281 ( \4435 , \4430 , \4434 );
and \U$4282 ( \4436 , \224 , \3103 );
and \U$4283 ( \4437 , \232 , \2934 );
nor \U$4284 ( \4438 , \4436 , \4437 );
xnor \U$4285 ( \4439 , \4438 , \2839 );
xor \U$4286 ( \4440 , \4435 , \4439 );
xor \U$4287 ( \4441 , \4426 , \4440 );
and \U$4288 ( \4442 , \240 , \3357 );
and \U$4289 ( \4443 , \247 , \3255 );
nor \U$4290 ( \4444 , \4442 , \4443 );
xnor \U$4291 ( \4445 , \4444 , \3156 );
and \U$4292 ( \4446 , \134 , \3813 );
and \U$4293 ( \4447 , \143 , \3557 );
nor \U$4294 ( \4448 , \4446 , \4447 );
xnor \U$4295 ( \4449 , \4448 , \3562 );
xor \U$4296 ( \4450 , \4445 , \4449 );
and \U$4297 ( \4451 , \150 , \4132 );
and \U$4298 ( \4452 , \158 , \4012 );
nor \U$4299 ( \4453 , \4451 , \4452 );
xnor \U$4300 ( \4454 , \4453 , \3925 );
xor \U$4301 ( \4455 , \4450 , \4454 );
xor \U$4302 ( \4456 , \4441 , \4455 );
xor \U$4303 ( \4457 , \4423 , \4456 );
xor \U$4304 ( \4458 , \4362 , \4457 );
xor \U$4305 ( \4459 , \4333 , \4458 );
xor \U$4306 ( \4460 , \4304 , \4459 );
xor \U$4307 ( \4461 , \4265 , \4460 );
and \U$4308 ( \4462 , \4064 , \4252 );
xor \U$4309 ( \4463 , \4461 , \4462 );
and \U$4310 ( \4464 , \4253 , \4254 );
and \U$4311 ( \4465 , \4255 , \4258 );
or \U$4312 ( \4466 , \4464 , \4465 );
xor \U$4313 ( \4467 , \4463 , \4466 );
buf g554b_GF_PartitionCandidate( \4468_nG554b , \4467 );
buf \U$4314 ( \4469 , \4468_nG554b );
and \U$4315 ( \4470 , \4269 , \4303 );
and \U$4316 ( \4471 , \4303 , \4459 );
and \U$4317 ( \4472 , \4269 , \4459 );
or \U$4318 ( \4473 , \4470 , \4471 , \4472 );
and \U$4319 ( \4474 , \4273 , \4277 );
and \U$4320 ( \4475 , \4277 , \4302 );
and \U$4321 ( \4476 , \4273 , \4302 );
or \U$4322 ( \4477 , \4474 , \4475 , \4476 );
and \U$4323 ( \4478 , \4318 , \4332 );
and \U$4324 ( \4479 , \4332 , \4458 );
and \U$4325 ( \4480 , \4318 , \4458 );
or \U$4326 ( \4481 , \4478 , \4479 , \4480 );
xor \U$4327 ( \4482 , \4477 , \4481 );
and \U$4328 ( \4483 , \4308 , \4312 );
and \U$4329 ( \4484 , \4312 , \4317 );
and \U$4330 ( \4485 , \4308 , \4317 );
or \U$4331 ( \4486 , \4483 , \4484 , \4485 );
and \U$4332 ( \4487 , \4282 , \4286 );
and \U$4333 ( \4488 , \4286 , \4301 );
and \U$4334 ( \4489 , \4282 , \4301 );
or \U$4335 ( \4490 , \4487 , \4488 , \4489 );
xor \U$4336 ( \4491 , \4486 , \4490 );
and \U$4337 ( \4492 , \4378 , \4422 );
and \U$4338 ( \4493 , \4422 , \4456 );
and \U$4339 ( \4494 , \4378 , \4456 );
or \U$4340 ( \4495 , \4492 , \4493 , \4494 );
xor \U$4341 ( \4496 , \4491 , \4495 );
xor \U$4342 ( \4497 , \4482 , \4496 );
xor \U$4343 ( \4498 , \4473 , \4497 );
and \U$4344 ( \4499 , \4322 , \4326 );
and \U$4345 ( \4500 , \4326 , \4331 );
and \U$4346 ( \4501 , \4322 , \4331 );
or \U$4347 ( \4502 , \4499 , \4500 , \4501 );
and \U$4348 ( \4503 , \4347 , \4361 );
and \U$4349 ( \4504 , \4361 , \4457 );
and \U$4350 ( \4505 , \4347 , \4457 );
or \U$4351 ( \4506 , \4503 , \4504 , \4505 );
xor \U$4352 ( \4507 , \4502 , \4506 );
and \U$4353 ( \4508 , \4337 , \4341 );
and \U$4354 ( \4509 , \4341 , \4346 );
and \U$4355 ( \4510 , \4337 , \4346 );
or \U$4356 ( \4511 , \4508 , \4509 , \4510 );
and \U$4357 ( \4512 , \4351 , \4355 );
and \U$4358 ( \4513 , \4355 , \4360 );
and \U$4359 ( \4514 , \4351 , \4360 );
or \U$4360 ( \4515 , \4512 , \4513 , \4514 );
xor \U$4361 ( \4516 , \4511 , \4515 );
and \U$4362 ( \4517 , \4426 , \4440 );
and \U$4363 ( \4518 , \4440 , \4455 );
and \U$4364 ( \4519 , \4426 , \4455 );
or \U$4365 ( \4520 , \4517 , \4518 , \4519 );
xor \U$4366 ( \4521 , \4516 , \4520 );
and \U$4367 ( \4522 , \4382 , \4386 );
and \U$4368 ( \4523 , \4386 , \4391 );
and \U$4369 ( \4524 , \4382 , \4391 );
or \U$4370 ( \4525 , \4522 , \4523 , \4524 );
and \U$4371 ( \4526 , \4291 , \4295 );
and \U$4372 ( \4527 , \4295 , \4300 );
and \U$4373 ( \4528 , \4291 , \4300 );
or \U$4374 ( \4529 , \4526 , \4527 , \4528 );
xor \U$4375 ( \4530 , \4525 , \4529 );
and \U$4376 ( \4531 , \4367 , \4371 );
and \U$4377 ( \4532 , \4371 , \4377 );
and \U$4378 ( \4533 , \4367 , \4377 );
or \U$4379 ( \4534 , \4531 , \4532 , \4533 );
xor \U$4380 ( \4535 , \4530 , \4534 );
and \U$4381 ( \4536 , \4430 , \4434 );
and \U$4382 ( \4537 , \4434 , \4439 );
and \U$4383 ( \4538 , \4430 , \4439 );
or \U$4384 ( \4539 , \4536 , \4537 , \4538 );
and \U$4385 ( \4540 , \4396 , \4400 );
and \U$4386 ( \4541 , \4400 , \4405 );
and \U$4387 ( \4542 , \4396 , \4405 );
or \U$4388 ( \4543 , \4540 , \4541 , \4542 );
xor \U$4389 ( \4544 , \4539 , \4543 );
and \U$4390 ( \4545 , \4411 , \4415 );
and \U$4391 ( \4546 , \4415 , \4420 );
and \U$4392 ( \4547 , \4411 , \4420 );
or \U$4393 ( \4548 , \4545 , \4546 , \4547 );
xor \U$4394 ( \4549 , \4544 , \4548 );
xor \U$4395 ( \4550 , \4535 , \4549 );
and \U$4396 ( \4551 , \4445 , \4449 );
and \U$4397 ( \4552 , \4449 , \4454 );
and \U$4398 ( \4553 , \4445 , \4454 );
or \U$4399 ( \4554 , \4551 , \4552 , \4553 );
and \U$4400 ( \4555 , \217 , \2669 );
and \U$4401 ( \4556 , \189 , \2538 );
nor \U$4402 ( \4557 , \4555 , \4556 );
xnor \U$4403 ( \4558 , \4557 , \2534 );
and \U$4404 ( \4559 , \232 , \3103 );
and \U$4405 ( \4560 , \209 , \2934 );
nor \U$4406 ( \4561 , \4559 , \4560 );
xnor \U$4407 ( \4562 , \4561 , \2839 );
xor \U$4408 ( \4563 , \4558 , \4562 );
and \U$4409 ( \4564 , \247 , \3357 );
and \U$4410 ( \4565 , \224 , \3255 );
nor \U$4411 ( \4566 , \4564 , \4565 );
xnor \U$4412 ( \4567 , \4566 , \3156 );
xor \U$4413 ( \4568 , \4563 , \4567 );
xor \U$4414 ( \4569 , \4554 , \4568 );
and \U$4415 ( \4570 , \143 , \3813 );
and \U$4416 ( \4571 , \240 , \3557 );
nor \U$4417 ( \4572 , \4570 , \4571 );
xnor \U$4418 ( \4573 , \4572 , \3562 );
and \U$4419 ( \4574 , \158 , \4132 );
and \U$4420 ( \4575 , \134 , \4012 );
nor \U$4421 ( \4576 , \4574 , \4575 );
xnor \U$4422 ( \4577 , \4576 , \3925 );
xor \U$4423 ( \4578 , \4573 , \4577 );
xor \U$4424 ( \4579 , \4373 , \4374 );
not \U$4425 ( \4580 , \4424 );
and \U$4426 ( \4581 , \4579 , \4580 );
and \U$4427 ( \4582 , \166 , \4581 );
and \U$4428 ( \4583 , \150 , \4424 );
nor \U$4429 ( \4584 , \4582 , \4583 );
xnor \U$4430 ( \4585 , \4584 , \4377 );
xor \U$4431 ( \4586 , \4578 , \4585 );
xor \U$4432 ( \4587 , \4569 , \4586 );
xor \U$4433 ( \4588 , \4550 , \4587 );
xor \U$4434 ( \4589 , \4521 , \4588 );
and \U$4435 ( \4590 , \4392 , \4406 );
and \U$4436 ( \4591 , \4406 , \4421 );
and \U$4437 ( \4592 , \4392 , \4421 );
or \U$4438 ( \4593 , \4590 , \4591 , \4592 );
and \U$4439 ( \4594 , \307 , \1824 );
and \U$4440 ( \4595 , \412 , \1739 );
nor \U$4441 ( \4596 , \4594 , \4595 );
xnor \U$4442 ( \4597 , \4596 , \1697 );
and \U$4443 ( \4598 , \185 , \2121 );
and \U$4444 ( \4599 , \261 , \2008 );
nor \U$4445 ( \4600 , \4598 , \4599 );
xnor \U$4446 ( \4601 , \4600 , \1961 );
xor \U$4447 ( \4602 , \4597 , \4601 );
and \U$4448 ( \4603 , \197 , \2400 );
and \U$4449 ( \4604 , \178 , \2246 );
nor \U$4450 ( \4605 , \4603 , \4604 );
xnor \U$4451 ( \4606 , \4605 , \2195 );
xor \U$4452 ( \4607 , \4602 , \4606 );
and \U$4453 ( \4608 , \2182 , \156 );
and \U$4454 ( \4609 , \2366 , \154 );
nor \U$4455 ( \4610 , \4608 , \4609 );
xnor \U$4456 ( \4611 , \4610 , \163 );
and \U$4457 ( \4612 , \1948 , \296 );
and \U$4458 ( \4613 , \2090 , \168 );
nor \U$4459 ( \4614 , \4612 , \4613 );
xnor \U$4460 ( \4615 , \4614 , \173 );
xor \U$4461 ( \4616 , \4611 , \4615 );
and \U$4462 ( \4617 , \1684 , \438 );
and \U$4463 ( \4618 , \1802 , \336 );
nor \U$4464 ( \4619 , \4617 , \4618 );
xnor \U$4465 ( \4620 , \4619 , \320 );
xor \U$4466 ( \4621 , \4616 , \4620 );
xor \U$4467 ( \4622 , \4607 , \4621 );
and \U$4468 ( \4623 , \1484 , \1086 );
and \U$4469 ( \4624 , \1601 , \508 );
nor \U$4470 ( \4625 , \4623 , \4624 );
xnor \U$4471 ( \4626 , \4625 , \487 );
and \U$4472 ( \4627 , \1192 , \1301 );
and \U$4473 ( \4628 , \1333 , \1246 );
nor \U$4474 ( \4629 , \4627 , \4628 );
xnor \U$4475 ( \4630 , \4629 , \1205 );
xor \U$4476 ( \4631 , \4626 , \4630 );
and \U$4477 ( \4632 , \474 , \1578 );
and \U$4478 ( \4633 , \1147 , \1431 );
nor \U$4479 ( \4634 , \4632 , \4633 );
xnor \U$4480 ( \4635 , \4634 , \1436 );
xor \U$4481 ( \4636 , \4631 , \4635 );
xor \U$4482 ( \4637 , \4622 , \4636 );
xor \U$4483 ( \4638 , \4593 , \4637 );
and \U$4484 ( \4639 , \3143 , \230 );
and \U$4485 ( \4640 , \3395 , \228 );
nor \U$4486 ( \4641 , \4639 , \4640 );
xnor \U$4487 ( \4642 , \4641 , \237 );
and \U$4488 ( \4643 , \2826 , \245 );
and \U$4489 ( \4644 , \3037 , \243 );
nor \U$4490 ( \4645 , \4643 , \4644 );
xnor \U$4491 ( \4646 , \4645 , \252 );
xor \U$4492 ( \4647 , \4642 , \4646 );
and \U$4493 ( \4648 , \2521 , \141 );
and \U$4494 ( \4649 , \2757 , \139 );
nor \U$4495 ( \4650 , \4648 , \4649 );
xnor \U$4496 ( \4651 , \4650 , \148 );
xor \U$4497 ( \4652 , \4647 , \4651 );
and \U$4498 ( \4653 , \4364 , \183 );
buf \U$4499 ( \4654 , RIb55e770_87);
and \U$4500 ( \4655 , \4654 , \180 );
nor \U$4501 ( \4656 , \4653 , \4655 );
xnor \U$4502 ( \4657 , \4656 , \179 );
and \U$4503 ( \4658 , \3912 , \195 );
and \U$4504 ( \4659 , \4160 , \193 );
nor \U$4505 ( \4660 , \4658 , \4659 );
xnor \U$4506 ( \4661 , \4660 , \202 );
xor \U$4507 ( \4662 , \4657 , \4661 );
and \U$4508 ( \4663 , \3646 , \215 );
and \U$4509 ( \4664 , \3736 , \213 );
nor \U$4510 ( \4665 , \4663 , \4664 );
xnor \U$4511 ( \4666 , \4665 , \222 );
xor \U$4512 ( \4667 , \4662 , \4666 );
xor \U$4513 ( \4668 , \4652 , \4667 );
xor \U$4514 ( \4669 , \4638 , \4668 );
xor \U$4515 ( \4670 , \4589 , \4669 );
xor \U$4516 ( \4671 , \4507 , \4670 );
xor \U$4517 ( \4672 , \4498 , \4671 );
and \U$4518 ( \4673 , \4265 , \4460 );
xor \U$4519 ( \4674 , \4672 , \4673 );
and \U$4520 ( \4675 , \4461 , \4462 );
and \U$4521 ( \4676 , \4463 , \4466 );
or \U$4522 ( \4677 , \4675 , \4676 );
xor \U$4523 ( \4678 , \4674 , \4677 );
buf g5549_GF_PartitionCandidate( \4679_nG5549 , \4678 );
buf \U$4524 ( \4680 , \4679_nG5549 );
and \U$4525 ( \4681 , \4477 , \4481 );
and \U$4526 ( \4682 , \4481 , \4496 );
and \U$4527 ( \4683 , \4477 , \4496 );
or \U$4528 ( \4684 , \4681 , \4682 , \4683 );
and \U$4529 ( \4685 , \4502 , \4506 );
and \U$4530 ( \4686 , \4506 , \4670 );
and \U$4531 ( \4687 , \4502 , \4670 );
or \U$4532 ( \4688 , \4685 , \4686 , \4687 );
and \U$4533 ( \4689 , \4486 , \4490 );
and \U$4534 ( \4690 , \4490 , \4495 );
and \U$4535 ( \4691 , \4486 , \4495 );
or \U$4536 ( \4692 , \4689 , \4690 , \4691 );
and \U$4537 ( \4693 , \4521 , \4588 );
and \U$4538 ( \4694 , \4588 , \4669 );
and \U$4539 ( \4695 , \4521 , \4669 );
or \U$4540 ( \4696 , \4693 , \4694 , \4695 );
xor \U$4541 ( \4697 , \4692 , \4696 );
and \U$4542 ( \4698 , \4525 , \4529 );
and \U$4543 ( \4699 , \4529 , \4534 );
and \U$4544 ( \4700 , \4525 , \4534 );
or \U$4545 ( \4701 , \4698 , \4699 , \4700 );
and \U$4546 ( \4702 , \4539 , \4543 );
and \U$4547 ( \4703 , \4543 , \4548 );
and \U$4548 ( \4704 , \4539 , \4548 );
or \U$4549 ( \4705 , \4702 , \4703 , \4704 );
xor \U$4550 ( \4706 , \4701 , \4705 );
and \U$4551 ( \4707 , \4554 , \4568 );
and \U$4552 ( \4708 , \4568 , \4586 );
and \U$4553 ( \4709 , \4554 , \4586 );
or \U$4554 ( \4710 , \4707 , \4708 , \4709 );
xor \U$4555 ( \4711 , \4706 , \4710 );
xor \U$4556 ( \4712 , \4697 , \4711 );
xor \U$4557 ( \4713 , \4688 , \4712 );
and \U$4558 ( \4714 , \4511 , \4515 );
and \U$4559 ( \4715 , \4515 , \4520 );
and \U$4560 ( \4716 , \4511 , \4520 );
or \U$4561 ( \4717 , \4714 , \4715 , \4716 );
and \U$4562 ( \4718 , \4535 , \4549 );
and \U$4563 ( \4719 , \4549 , \4587 );
and \U$4564 ( \4720 , \4535 , \4587 );
or \U$4565 ( \4721 , \4718 , \4719 , \4720 );
xor \U$4566 ( \4722 , \4717 , \4721 );
and \U$4567 ( \4723 , \4593 , \4637 );
and \U$4568 ( \4724 , \4637 , \4668 );
and \U$4569 ( \4725 , \4593 , \4668 );
or \U$4570 ( \4726 , \4723 , \4724 , \4725 );
xor \U$4571 ( \4727 , \4722 , \4726 );
and \U$4572 ( \4728 , \4611 , \4615 );
and \U$4573 ( \4729 , \4615 , \4620 );
and \U$4574 ( \4730 , \4611 , \4620 );
or \U$4575 ( \4731 , \4728 , \4729 , \4730 );
and \U$4576 ( \4732 , \4642 , \4646 );
and \U$4577 ( \4733 , \4646 , \4651 );
and \U$4578 ( \4734 , \4642 , \4651 );
or \U$4579 ( \4735 , \4732 , \4733 , \4734 );
xor \U$4580 ( \4736 , \4731 , \4735 );
and \U$4581 ( \4737 , \4657 , \4661 );
and \U$4582 ( \4738 , \4661 , \4666 );
and \U$4583 ( \4739 , \4657 , \4666 );
or \U$4584 ( \4740 , \4737 , \4738 , \4739 );
xor \U$4585 ( \4741 , \4736 , \4740 );
and \U$4586 ( \4742 , \4607 , \4621 );
and \U$4587 ( \4743 , \4621 , \4636 );
and \U$4588 ( \4744 , \4607 , \4636 );
or \U$4589 ( \4745 , \4742 , \4743 , \4744 );
and \U$4590 ( \4746 , \4652 , \4667 );
xor \U$4591 ( \4747 , \4745 , \4746 );
and \U$4592 ( \4748 , \4654 , \183 );
buf \U$4593 ( \4749 , RIb55e7e8_86);
and \U$4594 ( \4750 , \4749 , \180 );
nor \U$4595 ( \4751 , \4748 , \4750 );
xnor \U$4596 ( \4752 , \4751 , \179 );
and \U$4597 ( \4753 , \4160 , \195 );
and \U$4598 ( \4754 , \4364 , \193 );
nor \U$4599 ( \4755 , \4753 , \4754 );
xnor \U$4600 ( \4756 , \4755 , \202 );
xor \U$4601 ( \4757 , \4752 , \4756 );
buf \U$4602 ( \4758 , RIb560660_21);
buf \U$4603 ( \4759 , RIb5605e8_22);
and \U$4604 ( \4760 , \4759 , \4373 );
not \U$4605 ( \4761 , \4760 );
and \U$4606 ( \4762 , \4758 , \4761 );
xor \U$4607 ( \4763 , \4757 , \4762 );
and \U$4608 ( \4764 , \2757 , \141 );
and \U$4609 ( \4765 , \2826 , \139 );
nor \U$4610 ( \4766 , \4764 , \4765 );
xnor \U$4611 ( \4767 , \4766 , \148 );
and \U$4612 ( \4768 , \2366 , \156 );
and \U$4613 ( \4769 , \2521 , \154 );
nor \U$4614 ( \4770 , \4768 , \4769 );
xnor \U$4615 ( \4771 , \4770 , \163 );
xor \U$4616 ( \4772 , \4767 , \4771 );
and \U$4617 ( \4773 , \2090 , \296 );
and \U$4618 ( \4774 , \2182 , \168 );
nor \U$4619 ( \4775 , \4773 , \4774 );
xnor \U$4620 ( \4776 , \4775 , \173 );
xor \U$4621 ( \4777 , \4772 , \4776 );
xor \U$4622 ( \4778 , \4763 , \4777 );
and \U$4623 ( \4779 , \3736 , \215 );
and \U$4624 ( \4780 , \3912 , \213 );
nor \U$4625 ( \4781 , \4779 , \4780 );
xnor \U$4626 ( \4782 , \4781 , \222 );
and \U$4627 ( \4783 , \3395 , \230 );
and \U$4628 ( \4784 , \3646 , \228 );
nor \U$4629 ( \4785 , \4783 , \4784 );
xnor \U$4630 ( \4786 , \4785 , \237 );
xor \U$4631 ( \4787 , \4782 , \4786 );
and \U$4632 ( \4788 , \3037 , \245 );
and \U$4633 ( \4789 , \3143 , \243 );
nor \U$4634 ( \4790 , \4788 , \4789 );
xnor \U$4635 ( \4791 , \4790 , \252 );
xor \U$4636 ( \4792 , \4787 , \4791 );
xor \U$4637 ( \4793 , \4778 , \4792 );
xor \U$4638 ( \4794 , \4747 , \4793 );
xor \U$4639 ( \4795 , \4741 , \4794 );
and \U$4640 ( \4796 , \4597 , \4601 );
and \U$4641 ( \4797 , \4601 , \4606 );
and \U$4642 ( \4798 , \4597 , \4606 );
or \U$4643 ( \4799 , \4796 , \4797 , \4798 );
and \U$4644 ( \4800 , \4558 , \4562 );
and \U$4645 ( \4801 , \4562 , \4567 );
and \U$4646 ( \4802 , \4558 , \4567 );
or \U$4647 ( \4803 , \4800 , \4801 , \4802 );
xor \U$4648 ( \4804 , \4799 , \4803 );
and \U$4649 ( \4805 , \4626 , \4630 );
and \U$4650 ( \4806 , \4630 , \4635 );
and \U$4651 ( \4807 , \4626 , \4635 );
or \U$4652 ( \4808 , \4805 , \4806 , \4807 );
xor \U$4653 ( \4809 , \4804 , \4808 );
and \U$4654 ( \4810 , \178 , \2400 );
and \U$4655 ( \4811 , \185 , \2246 );
nor \U$4656 ( \4812 , \4810 , \4811 );
xnor \U$4657 ( \4813 , \4812 , \2195 );
and \U$4658 ( \4814 , \189 , \2669 );
and \U$4659 ( \4815 , \197 , \2538 );
nor \U$4660 ( \4816 , \4814 , \4815 );
xnor \U$4661 ( \4817 , \4816 , \2534 );
xor \U$4662 ( \4818 , \4813 , \4817 );
and \U$4663 ( \4819 , \209 , \3103 );
and \U$4664 ( \4820 , \217 , \2934 );
nor \U$4665 ( \4821 , \4819 , \4820 );
xnor \U$4666 ( \4822 , \4821 , \2839 );
xor \U$4667 ( \4823 , \4818 , \4822 );
and \U$4668 ( \4824 , \1802 , \438 );
and \U$4669 ( \4825 , \1948 , \336 );
nor \U$4670 ( \4826 , \4824 , \4825 );
xnor \U$4671 ( \4827 , \4826 , \320 );
and \U$4672 ( \4828 , \1601 , \1086 );
and \U$4673 ( \4829 , \1684 , \508 );
nor \U$4674 ( \4830 , \4828 , \4829 );
xnor \U$4675 ( \4831 , \4830 , \487 );
xor \U$4676 ( \4832 , \4827 , \4831 );
and \U$4677 ( \4833 , \1333 , \1301 );
and \U$4678 ( \4834 , \1484 , \1246 );
nor \U$4679 ( \4835 , \4833 , \4834 );
xnor \U$4680 ( \4836 , \4835 , \1205 );
xor \U$4681 ( \4837 , \4832 , \4836 );
xor \U$4682 ( \4838 , \4823 , \4837 );
and \U$4683 ( \4839 , \1147 , \1578 );
and \U$4684 ( \4840 , \1192 , \1431 );
nor \U$4685 ( \4841 , \4839 , \4840 );
xnor \U$4686 ( \4842 , \4841 , \1436 );
and \U$4687 ( \4843 , \412 , \1824 );
and \U$4688 ( \4844 , \474 , \1739 );
nor \U$4689 ( \4845 , \4843 , \4844 );
xnor \U$4690 ( \4846 , \4845 , \1697 );
xor \U$4691 ( \4847 , \4842 , \4846 );
and \U$4692 ( \4848 , \261 , \2121 );
and \U$4693 ( \4849 , \307 , \2008 );
nor \U$4694 ( \4850 , \4848 , \4849 );
xnor \U$4695 ( \4851 , \4850 , \1961 );
xor \U$4696 ( \4852 , \4847 , \4851 );
xor \U$4697 ( \4853 , \4838 , \4852 );
xor \U$4698 ( \4854 , \4809 , \4853 );
and \U$4699 ( \4855 , \4573 , \4577 );
and \U$4700 ( \4856 , \4577 , \4585 );
and \U$4701 ( \4857 , \4573 , \4585 );
or \U$4702 ( \4858 , \4855 , \4856 , \4857 );
and \U$4703 ( \4859 , \224 , \3357 );
and \U$4704 ( \4860 , \232 , \3255 );
nor \U$4705 ( \4861 , \4859 , \4860 );
xnor \U$4706 ( \4862 , \4861 , \3156 );
and \U$4707 ( \4863 , \240 , \3813 );
and \U$4708 ( \4864 , \247 , \3557 );
nor \U$4709 ( \4865 , \4863 , \4864 );
xnor \U$4710 ( \4866 , \4865 , \3562 );
xor \U$4711 ( \4867 , \4862 , \4866 );
and \U$4712 ( \4868 , \134 , \4132 );
and \U$4713 ( \4869 , \143 , \4012 );
nor \U$4714 ( \4870 , \4868 , \4869 );
xnor \U$4715 ( \4871 , \4870 , \3925 );
xor \U$4716 ( \4872 , \4867 , \4871 );
xor \U$4717 ( \4873 , \4858 , \4872 );
and \U$4718 ( \4874 , \150 , \4581 );
and \U$4719 ( \4875 , \158 , \4424 );
nor \U$4720 ( \4876 , \4874 , \4875 );
xnor \U$4721 ( \4877 , \4876 , \4377 );
xor \U$4722 ( \4878 , \4759 , \4373 );
nand \U$4723 ( \4879 , \166 , \4878 );
xnor \U$4724 ( \4880 , \4879 , \4762 );
xor \U$4725 ( \4881 , \4877 , \4880 );
xor \U$4726 ( \4882 , \4873 , \4881 );
xor \U$4727 ( \4883 , \4854 , \4882 );
xor \U$4728 ( \4884 , \4795 , \4883 );
xor \U$4729 ( \4885 , \4727 , \4884 );
xor \U$4730 ( \4886 , \4713 , \4885 );
xor \U$4731 ( \4887 , \4684 , \4886 );
and \U$4732 ( \4888 , \4473 , \4497 );
and \U$4733 ( \4889 , \4497 , \4671 );
and \U$4734 ( \4890 , \4473 , \4671 );
or \U$4735 ( \4891 , \4888 , \4889 , \4890 );
xor \U$4736 ( \4892 , \4887 , \4891 );
and \U$4737 ( \4893 , \4672 , \4673 );
and \U$4738 ( \4894 , \4674 , \4677 );
or \U$4739 ( \4895 , \4893 , \4894 );
xor \U$4740 ( \4896 , \4892 , \4895 );
buf g5547_GF_PartitionCandidate( \4897_nG5547 , \4896 );
buf \U$4741 ( \4898 , \4897_nG5547 );
and \U$4742 ( \4899 , \4688 , \4712 );
and \U$4743 ( \4900 , \4712 , \4885 );
and \U$4744 ( \4901 , \4688 , \4885 );
or \U$4745 ( \4902 , \4899 , \4900 , \4901 );
and \U$4746 ( \4903 , \4717 , \4721 );
and \U$4747 ( \4904 , \4721 , \4726 );
and \U$4748 ( \4905 , \4717 , \4726 );
or \U$4749 ( \4906 , \4903 , \4904 , \4905 );
and \U$4750 ( \4907 , \4741 , \4794 );
and \U$4751 ( \4908 , \4794 , \4883 );
and \U$4752 ( \4909 , \4741 , \4883 );
or \U$4753 ( \4910 , \4907 , \4908 , \4909 );
xor \U$4754 ( \4911 , \4906 , \4910 );
and \U$4755 ( \4912 , \4763 , \4777 );
and \U$4756 ( \4913 , \4777 , \4792 );
and \U$4757 ( \4914 , \4763 , \4792 );
or \U$4758 ( \4915 , \4912 , \4913 , \4914 );
and \U$4759 ( \4916 , \4823 , \4837 );
and \U$4760 ( \4917 , \4837 , \4852 );
and \U$4761 ( \4918 , \4823 , \4852 );
or \U$4762 ( \4919 , \4916 , \4917 , \4918 );
xor \U$4763 ( \4920 , \4915 , \4919 );
and \U$4764 ( \4921 , \4749 , \183 );
buf \U$4765 ( \4922 , RIb55e860_85);
and \U$4766 ( \4923 , \4922 , \180 );
nor \U$4767 ( \4924 , \4921 , \4923 );
xnor \U$4768 ( \4925 , \4924 , \179 );
and \U$4769 ( \4926 , \4364 , \195 );
and \U$4770 ( \4927 , \4654 , \193 );
nor \U$4771 ( \4928 , \4926 , \4927 );
xnor \U$4772 ( \4929 , \4928 , \202 );
xor \U$4773 ( \4930 , \4925 , \4929 );
and \U$4774 ( \4931 , \3912 , \215 );
and \U$4775 ( \4932 , \4160 , \213 );
nor \U$4776 ( \4933 , \4931 , \4932 );
xnor \U$4777 ( \4934 , \4933 , \222 );
xor \U$4778 ( \4935 , \4930 , \4934 );
xor \U$4779 ( \4936 , \4920 , \4935 );
xor \U$4780 ( \4937 , \4911 , \4936 );
xor \U$4781 ( \4938 , \4902 , \4937 );
and \U$4782 ( \4939 , \4692 , \4696 );
and \U$4783 ( \4940 , \4696 , \4711 );
and \U$4784 ( \4941 , \4692 , \4711 );
or \U$4785 ( \4942 , \4939 , \4940 , \4941 );
and \U$4786 ( \4943 , \4727 , \4884 );
xor \U$4787 ( \4944 , \4942 , \4943 );
and \U$4788 ( \4945 , \4799 , \4803 );
and \U$4789 ( \4946 , \4803 , \4808 );
and \U$4790 ( \4947 , \4799 , \4808 );
or \U$4791 ( \4948 , \4945 , \4946 , \4947 );
and \U$4792 ( \4949 , \4731 , \4735 );
and \U$4793 ( \4950 , \4735 , \4740 );
and \U$4794 ( \4951 , \4731 , \4740 );
or \U$4795 ( \4952 , \4949 , \4950 , \4951 );
xor \U$4796 ( \4953 , \4948 , \4952 );
and \U$4797 ( \4954 , \4858 , \4872 );
and \U$4798 ( \4955 , \4872 , \4881 );
and \U$4799 ( \4956 , \4858 , \4881 );
or \U$4800 ( \4957 , \4954 , \4955 , \4956 );
xor \U$4801 ( \4958 , \4953 , \4957 );
and \U$4802 ( \4959 , \4701 , \4705 );
and \U$4803 ( \4960 , \4705 , \4710 );
and \U$4804 ( \4961 , \4701 , \4710 );
or \U$4805 ( \4962 , \4959 , \4960 , \4961 );
and \U$4806 ( \4963 , \4745 , \4746 );
and \U$4807 ( \4964 , \4746 , \4793 );
and \U$4808 ( \4965 , \4745 , \4793 );
or \U$4809 ( \4966 , \4963 , \4964 , \4965 );
xor \U$4810 ( \4967 , \4962 , \4966 );
and \U$4811 ( \4968 , \4809 , \4853 );
and \U$4812 ( \4969 , \4853 , \4882 );
and \U$4813 ( \4970 , \4809 , \4882 );
or \U$4814 ( \4971 , \4968 , \4969 , \4970 );
xor \U$4815 ( \4972 , \4967 , \4971 );
xor \U$4816 ( \4973 , \4958 , \4972 );
and \U$4817 ( \4974 , \4813 , \4817 );
and \U$4818 ( \4975 , \4817 , \4822 );
and \U$4819 ( \4976 , \4813 , \4822 );
or \U$4820 ( \4977 , \4974 , \4975 , \4976 );
and \U$4821 ( \4978 , \4827 , \4831 );
and \U$4822 ( \4979 , \4831 , \4836 );
and \U$4823 ( \4980 , \4827 , \4836 );
or \U$4824 ( \4981 , \4978 , \4979 , \4980 );
xor \U$4825 ( \4982 , \4977 , \4981 );
and \U$4826 ( \4983 , \4842 , \4846 );
and \U$4827 ( \4984 , \4846 , \4851 );
and \U$4828 ( \4985 , \4842 , \4851 );
or \U$4829 ( \4986 , \4983 , \4984 , \4985 );
xor \U$4830 ( \4987 , \4982 , \4986 );
and \U$4831 ( \4988 , \4752 , \4756 );
and \U$4832 ( \4989 , \4756 , \4762 );
and \U$4833 ( \4990 , \4752 , \4762 );
or \U$4834 ( \4991 , \4988 , \4989 , \4990 );
and \U$4835 ( \4992 , \4767 , \4771 );
and \U$4836 ( \4993 , \4771 , \4776 );
and \U$4837 ( \4994 , \4767 , \4776 );
or \U$4838 ( \4995 , \4992 , \4993 , \4994 );
xor \U$4839 ( \4996 , \4991 , \4995 );
and \U$4840 ( \4997 , \4782 , \4786 );
and \U$4841 ( \4998 , \4786 , \4791 );
and \U$4842 ( \4999 , \4782 , \4791 );
or \U$4843 ( \5000 , \4997 , \4998 , \4999 );
xor \U$4844 ( \5001 , \4996 , \5000 );
xor \U$4845 ( \5002 , \4987 , \5001 );
and \U$4846 ( \5003 , \4862 , \4866 );
and \U$4847 ( \5004 , \4866 , \4871 );
and \U$4848 ( \5005 , \4862 , \4871 );
or \U$4849 ( \5006 , \5003 , \5004 , \5005 );
and \U$4850 ( \5007 , \4877 , \4880 );
xor \U$4851 ( \5008 , \5006 , \5007 );
xor \U$4852 ( \5009 , \4758 , \4759 );
not \U$4853 ( \5010 , \4878 );
and \U$4854 ( \5011 , \5009 , \5010 );
and \U$4855 ( \5012 , \166 , \5011 );
and \U$4856 ( \5013 , \150 , \4878 );
nor \U$4857 ( \5014 , \5012 , \5013 );
xnor \U$4858 ( \5015 , \5014 , \4762 );
xor \U$4859 ( \5016 , \5008 , \5015 );
and \U$4860 ( \5017 , \3646 , \230 );
and \U$4861 ( \5018 , \3736 , \228 );
nor \U$4862 ( \5019 , \5017 , \5018 );
xnor \U$4863 ( \5020 , \5019 , \237 );
and \U$4864 ( \5021 , \3143 , \245 );
and \U$4865 ( \5022 , \3395 , \243 );
nor \U$4866 ( \5023 , \5021 , \5022 );
xnor \U$4867 ( \5024 , \5023 , \252 );
xor \U$4868 ( \5025 , \5020 , \5024 );
and \U$4869 ( \5026 , \2826 , \141 );
and \U$4870 ( \5027 , \3037 , \139 );
nor \U$4871 ( \5028 , \5026 , \5027 );
xnor \U$4872 ( \5029 , \5028 , \148 );
xor \U$4873 ( \5030 , \5025 , \5029 );
and \U$4874 ( \5031 , \1684 , \1086 );
and \U$4875 ( \5032 , \1802 , \508 );
nor \U$4876 ( \5033 , \5031 , \5032 );
xnor \U$4877 ( \5034 , \5033 , \487 );
and \U$4878 ( \5035 , \1484 , \1301 );
and \U$4879 ( \5036 , \1601 , \1246 );
nor \U$4880 ( \5037 , \5035 , \5036 );
xnor \U$4881 ( \5038 , \5037 , \1205 );
xor \U$4882 ( \5039 , \5034 , \5038 );
and \U$4883 ( \5040 , \1192 , \1578 );
and \U$4884 ( \5041 , \1333 , \1431 );
nor \U$4885 ( \5042 , \5040 , \5041 );
xnor \U$4886 ( \5043 , \5042 , \1436 );
xor \U$4887 ( \5044 , \5039 , \5043 );
xor \U$4888 ( \5045 , \5030 , \5044 );
and \U$4889 ( \5046 , \2521 , \156 );
and \U$4890 ( \5047 , \2757 , \154 );
nor \U$4891 ( \5048 , \5046 , \5047 );
xnor \U$4892 ( \5049 , \5048 , \163 );
and \U$4893 ( \5050 , \2182 , \296 );
and \U$4894 ( \5051 , \2366 , \168 );
nor \U$4895 ( \5052 , \5050 , \5051 );
xnor \U$4896 ( \5053 , \5052 , \173 );
xor \U$4897 ( \5054 , \5049 , \5053 );
and \U$4898 ( \5055 , \1948 , \438 );
and \U$4899 ( \5056 , \2090 , \336 );
nor \U$4900 ( \5057 , \5055 , \5056 );
xnor \U$4901 ( \5058 , \5057 , \320 );
xor \U$4902 ( \5059 , \5054 , \5058 );
xor \U$4903 ( \5060 , \5045 , \5059 );
xor \U$4904 ( \5061 , \5016 , \5060 );
and \U$4905 ( \5062 , \474 , \1824 );
and \U$4906 ( \5063 , \1147 , \1739 );
nor \U$4907 ( \5064 , \5062 , \5063 );
xnor \U$4908 ( \5065 , \5064 , \1697 );
and \U$4909 ( \5066 , \307 , \2121 );
and \U$4910 ( \5067 , \412 , \2008 );
nor \U$4911 ( \5068 , \5066 , \5067 );
xnor \U$4912 ( \5069 , \5068 , \1961 );
xor \U$4913 ( \5070 , \5065 , \5069 );
and \U$4914 ( \5071 , \185 , \2400 );
and \U$4915 ( \5072 , \261 , \2246 );
nor \U$4916 ( \5073 , \5071 , \5072 );
xnor \U$4917 ( \5074 , \5073 , \2195 );
xor \U$4918 ( \5075 , \5070 , \5074 );
and \U$4919 ( \5076 , \247 , \3813 );
and \U$4920 ( \5077 , \224 , \3557 );
nor \U$4921 ( \5078 , \5076 , \5077 );
xnor \U$4922 ( \5079 , \5078 , \3562 );
and \U$4923 ( \5080 , \143 , \4132 );
and \U$4924 ( \5081 , \240 , \4012 );
nor \U$4925 ( \5082 , \5080 , \5081 );
xnor \U$4926 ( \5083 , \5082 , \3925 );
xor \U$4927 ( \5084 , \5079 , \5083 );
and \U$4928 ( \5085 , \158 , \4581 );
and \U$4929 ( \5086 , \134 , \4424 );
nor \U$4930 ( \5087 , \5085 , \5086 );
xnor \U$4931 ( \5088 , \5087 , \4377 );
xor \U$4932 ( \5089 , \5084 , \5088 );
xor \U$4933 ( \5090 , \5075 , \5089 );
and \U$4934 ( \5091 , \197 , \2669 );
and \U$4935 ( \5092 , \178 , \2538 );
nor \U$4936 ( \5093 , \5091 , \5092 );
xnor \U$4937 ( \5094 , \5093 , \2534 );
and \U$4938 ( \5095 , \217 , \3103 );
and \U$4939 ( \5096 , \189 , \2934 );
nor \U$4940 ( \5097 , \5095 , \5096 );
xnor \U$4941 ( \5098 , \5097 , \2839 );
xor \U$4942 ( \5099 , \5094 , \5098 );
and \U$4943 ( \5100 , \232 , \3357 );
and \U$4944 ( \5101 , \209 , \3255 );
nor \U$4945 ( \5102 , \5100 , \5101 );
xnor \U$4946 ( \5103 , \5102 , \3156 );
xor \U$4947 ( \5104 , \5099 , \5103 );
xor \U$4948 ( \5105 , \5090 , \5104 );
xor \U$4949 ( \5106 , \5061 , \5105 );
xor \U$4950 ( \5107 , \5002 , \5106 );
xor \U$4951 ( \5108 , \4973 , \5107 );
xor \U$4952 ( \5109 , \4944 , \5108 );
xor \U$4953 ( \5110 , \4938 , \5109 );
and \U$4954 ( \5111 , \4684 , \4886 );
xor \U$4955 ( \5112 , \5110 , \5111 );
and \U$4956 ( \5113 , \4887 , \4891 );
and \U$4957 ( \5114 , \4892 , \4895 );
or \U$4958 ( \5115 , \5113 , \5114 );
xor \U$4959 ( \5116 , \5112 , \5115 );
buf g5545_GF_PartitionCandidate( \5117_nG5545 , \5116 );
buf \U$4960 ( \5118 , \5117_nG5545 );
and \U$4961 ( \5119 , \4942 , \4943 );
and \U$4962 ( \5120 , \4943 , \5108 );
and \U$4963 ( \5121 , \4942 , \5108 );
or \U$4964 ( \5122 , \5119 , \5120 , \5121 );
and \U$4965 ( \5123 , \4906 , \4910 );
and \U$4966 ( \5124 , \4910 , \4936 );
and \U$4967 ( \5125 , \4906 , \4936 );
or \U$4968 ( \5126 , \5123 , \5124 , \5125 );
and \U$4969 ( \5127 , \4958 , \4972 );
and \U$4970 ( \5128 , \4972 , \5107 );
and \U$4971 ( \5129 , \4958 , \5107 );
or \U$4972 ( \5130 , \5127 , \5128 , \5129 );
xor \U$4973 ( \5131 , \5126 , \5130 );
and \U$4974 ( \5132 , \4925 , \4929 );
and \U$4975 ( \5133 , \4929 , \4934 );
and \U$4976 ( \5134 , \4925 , \4934 );
or \U$4977 ( \5135 , \5132 , \5133 , \5134 );
and \U$4978 ( \5136 , \5020 , \5024 );
and \U$4979 ( \5137 , \5024 , \5029 );
and \U$4980 ( \5138 , \5020 , \5029 );
or \U$4981 ( \5139 , \5136 , \5137 , \5138 );
xor \U$4982 ( \5140 , \5135 , \5139 );
and \U$4983 ( \5141 , \5049 , \5053 );
and \U$4984 ( \5142 , \5053 , \5058 );
and \U$4985 ( \5143 , \5049 , \5058 );
or \U$4986 ( \5144 , \5141 , \5142 , \5143 );
xor \U$4987 ( \5145 , \5140 , \5144 );
and \U$4988 ( \5146 , \5030 , \5044 );
and \U$4989 ( \5147 , \5044 , \5059 );
and \U$4990 ( \5148 , \5030 , \5059 );
or \U$4991 ( \5149 , \5146 , \5147 , \5148 );
and \U$4992 ( \5150 , \5075 , \5089 );
and \U$4993 ( \5151 , \5089 , \5104 );
and \U$4994 ( \5152 , \5075 , \5104 );
or \U$4995 ( \5153 , \5150 , \5151 , \5152 );
xor \U$4996 ( \5154 , \5149 , \5153 );
and \U$4997 ( \5155 , \4922 , \183 );
buf \U$4998 ( \5156 , RIb55e8d8_84);
and \U$4999 ( \5157 , \5156 , \180 );
nor \U$5000 ( \5158 , \5155 , \5157 );
xnor \U$5001 ( \5159 , \5158 , \179 );
and \U$5002 ( \5160 , \4654 , \195 );
and \U$5003 ( \5161 , \4749 , \193 );
nor \U$5004 ( \5162 , \5160 , \5161 );
xnor \U$5005 ( \5163 , \5162 , \202 );
xor \U$5006 ( \5164 , \5159 , \5163 );
buf \U$5007 ( \5165 , RIb560750_19);
buf \U$5008 ( \5166 , RIb5606d8_20);
and \U$5009 ( \5167 , \5166 , \4758 );
not \U$5010 ( \5168 , \5167 );
and \U$5011 ( \5169 , \5165 , \5168 );
xor \U$5012 ( \5170 , \5164 , \5169 );
and \U$5013 ( \5171 , \3037 , \141 );
and \U$5014 ( \5172 , \3143 , \139 );
nor \U$5015 ( \5173 , \5171 , \5172 );
xnor \U$5016 ( \5174 , \5173 , \148 );
and \U$5017 ( \5175 , \2757 , \156 );
and \U$5018 ( \5176 , \2826 , \154 );
nor \U$5019 ( \5177 , \5175 , \5176 );
xnor \U$5020 ( \5178 , \5177 , \163 );
xor \U$5021 ( \5179 , \5174 , \5178 );
and \U$5022 ( \5180 , \2366 , \296 );
and \U$5023 ( \5181 , \2521 , \168 );
nor \U$5024 ( \5182 , \5180 , \5181 );
xnor \U$5025 ( \5183 , \5182 , \173 );
xor \U$5026 ( \5184 , \5179 , \5183 );
xor \U$5027 ( \5185 , \5170 , \5184 );
and \U$5028 ( \5186 , \4160 , \215 );
and \U$5029 ( \5187 , \4364 , \213 );
nor \U$5030 ( \5188 , \5186 , \5187 );
xnor \U$5031 ( \5189 , \5188 , \222 );
and \U$5032 ( \5190 , \3736 , \230 );
and \U$5033 ( \5191 , \3912 , \228 );
nor \U$5034 ( \5192 , \5190 , \5191 );
xnor \U$5035 ( \5193 , \5192 , \237 );
xor \U$5036 ( \5194 , \5189 , \5193 );
and \U$5037 ( \5195 , \3395 , \245 );
and \U$5038 ( \5196 , \3646 , \243 );
nor \U$5039 ( \5197 , \5195 , \5196 );
xnor \U$5040 ( \5198 , \5197 , \252 );
xor \U$5041 ( \5199 , \5194 , \5198 );
xor \U$5042 ( \5200 , \5185 , \5199 );
xor \U$5043 ( \5201 , \5154 , \5200 );
xor \U$5044 ( \5202 , \5145 , \5201 );
and \U$5045 ( \5203 , \5065 , \5069 );
and \U$5046 ( \5204 , \5069 , \5074 );
and \U$5047 ( \5205 , \5065 , \5074 );
or \U$5048 ( \5206 , \5203 , \5204 , \5205 );
and \U$5049 ( \5207 , \5094 , \5098 );
and \U$5050 ( \5208 , \5098 , \5103 );
and \U$5051 ( \5209 , \5094 , \5103 );
or \U$5052 ( \5210 , \5207 , \5208 , \5209 );
xor \U$5053 ( \5211 , \5206 , \5210 );
and \U$5054 ( \5212 , \5034 , \5038 );
and \U$5055 ( \5213 , \5038 , \5043 );
and \U$5056 ( \5214 , \5034 , \5043 );
or \U$5057 ( \5215 , \5212 , \5213 , \5214 );
xor \U$5058 ( \5216 , \5211 , \5215 );
and \U$5059 ( \5217 , \2090 , \438 );
and \U$5060 ( \5218 , \2182 , \336 );
nor \U$5061 ( \5219 , \5217 , \5218 );
xnor \U$5062 ( \5220 , \5219 , \320 );
and \U$5063 ( \5221 , \1802 , \1086 );
and \U$5064 ( \5222 , \1948 , \508 );
nor \U$5065 ( \5223 , \5221 , \5222 );
xnor \U$5066 ( \5224 , \5223 , \487 );
xor \U$5067 ( \5225 , \5220 , \5224 );
and \U$5068 ( \5226 , \1601 , \1301 );
and \U$5069 ( \5227 , \1684 , \1246 );
nor \U$5070 ( \5228 , \5226 , \5227 );
xnor \U$5071 ( \5229 , \5228 , \1205 );
xor \U$5072 ( \5230 , \5225 , \5229 );
and \U$5073 ( \5231 , \1333 , \1578 );
and \U$5074 ( \5232 , \1484 , \1431 );
nor \U$5075 ( \5233 , \5231 , \5232 );
xnor \U$5076 ( \5234 , \5233 , \1436 );
and \U$5077 ( \5235 , \1147 , \1824 );
and \U$5078 ( \5236 , \1192 , \1739 );
nor \U$5079 ( \5237 , \5235 , \5236 );
xnor \U$5080 ( \5238 , \5237 , \1697 );
xor \U$5081 ( \5239 , \5234 , \5238 );
and \U$5082 ( \5240 , \412 , \2121 );
and \U$5083 ( \5241 , \474 , \2008 );
nor \U$5084 ( \5242 , \5240 , \5241 );
xnor \U$5085 ( \5243 , \5242 , \1961 );
xor \U$5086 ( \5244 , \5239 , \5243 );
xor \U$5087 ( \5245 , \5230 , \5244 );
and \U$5088 ( \5246 , \261 , \2400 );
and \U$5089 ( \5247 , \307 , \2246 );
nor \U$5090 ( \5248 , \5246 , \5247 );
xnor \U$5091 ( \5249 , \5248 , \2195 );
and \U$5092 ( \5250 , \178 , \2669 );
and \U$5093 ( \5251 , \185 , \2538 );
nor \U$5094 ( \5252 , \5250 , \5251 );
xnor \U$5095 ( \5253 , \5252 , \2534 );
xor \U$5096 ( \5254 , \5249 , \5253 );
and \U$5097 ( \5255 , \189 , \3103 );
and \U$5098 ( \5256 , \197 , \2934 );
nor \U$5099 ( \5257 , \5255 , \5256 );
xnor \U$5100 ( \5258 , \5257 , \2839 );
xor \U$5101 ( \5259 , \5254 , \5258 );
xor \U$5102 ( \5260 , \5245 , \5259 );
xor \U$5103 ( \5261 , \5216 , \5260 );
and \U$5104 ( \5262 , \5079 , \5083 );
and \U$5105 ( \5263 , \5083 , \5088 );
and \U$5106 ( \5264 , \5079 , \5088 );
or \U$5107 ( \5265 , \5262 , \5263 , \5264 );
and \U$5108 ( \5266 , \134 , \4581 );
and \U$5109 ( \5267 , \143 , \4424 );
nor \U$5110 ( \5268 , \5266 , \5267 );
xnor \U$5111 ( \5269 , \5268 , \4377 );
and \U$5112 ( \5270 , \150 , \5011 );
and \U$5113 ( \5271 , \158 , \4878 );
nor \U$5114 ( \5272 , \5270 , \5271 );
xnor \U$5115 ( \5273 , \5272 , \4762 );
xor \U$5116 ( \5274 , \5269 , \5273 );
xor \U$5117 ( \5275 , \5166 , \4758 );
nand \U$5118 ( \5276 , \166 , \5275 );
xnor \U$5119 ( \5277 , \5276 , \5169 );
xor \U$5120 ( \5278 , \5274 , \5277 );
xor \U$5121 ( \5279 , \5265 , \5278 );
and \U$5122 ( \5280 , \209 , \3357 );
and \U$5123 ( \5281 , \217 , \3255 );
nor \U$5124 ( \5282 , \5280 , \5281 );
xnor \U$5125 ( \5283 , \5282 , \3156 );
and \U$5126 ( \5284 , \224 , \3813 );
and \U$5127 ( \5285 , \232 , \3557 );
nor \U$5128 ( \5286 , \5284 , \5285 );
xnor \U$5129 ( \5287 , \5286 , \3562 );
xor \U$5130 ( \5288 , \5283 , \5287 );
and \U$5131 ( \5289 , \240 , \4132 );
and \U$5132 ( \5290 , \247 , \4012 );
nor \U$5133 ( \5291 , \5289 , \5290 );
xnor \U$5134 ( \5292 , \5291 , \3925 );
xor \U$5135 ( \5293 , \5288 , \5292 );
xor \U$5136 ( \5294 , \5279 , \5293 );
xor \U$5137 ( \5295 , \5261 , \5294 );
xor \U$5138 ( \5296 , \5202 , \5295 );
xor \U$5139 ( \5297 , \5131 , \5296 );
xor \U$5140 ( \5298 , \5122 , \5297 );
and \U$5141 ( \5299 , \4948 , \4952 );
and \U$5142 ( \5300 , \4952 , \4957 );
and \U$5143 ( \5301 , \4948 , \4957 );
or \U$5144 ( \5302 , \5299 , \5300 , \5301 );
and \U$5145 ( \5303 , \4915 , \4919 );
and \U$5146 ( \5304 , \4919 , \4935 );
and \U$5147 ( \5305 , \4915 , \4935 );
or \U$5148 ( \5306 , \5303 , \5304 , \5305 );
xor \U$5149 ( \5307 , \5302 , \5306 );
and \U$5150 ( \5308 , \5016 , \5060 );
and \U$5151 ( \5309 , \5060 , \5105 );
and \U$5152 ( \5310 , \5016 , \5105 );
or \U$5153 ( \5311 , \5308 , \5309 , \5310 );
xor \U$5154 ( \5312 , \5307 , \5311 );
and \U$5155 ( \5313 , \4962 , \4966 );
and \U$5156 ( \5314 , \4966 , \4971 );
and \U$5157 ( \5315 , \4962 , \4971 );
or \U$5158 ( \5316 , \5313 , \5314 , \5315 );
and \U$5159 ( \5317 , \4987 , \5001 );
and \U$5160 ( \5318 , \5001 , \5106 );
and \U$5161 ( \5319 , \4987 , \5106 );
or \U$5162 ( \5320 , \5317 , \5318 , \5319 );
xor \U$5163 ( \5321 , \5316 , \5320 );
and \U$5164 ( \5322 , \4977 , \4981 );
and \U$5165 ( \5323 , \4981 , \4986 );
and \U$5166 ( \5324 , \4977 , \4986 );
or \U$5167 ( \5325 , \5322 , \5323 , \5324 );
and \U$5168 ( \5326 , \4991 , \4995 );
and \U$5169 ( \5327 , \4995 , \5000 );
and \U$5170 ( \5328 , \4991 , \5000 );
or \U$5171 ( \5329 , \5326 , \5327 , \5328 );
xor \U$5172 ( \5330 , \5325 , \5329 );
and \U$5173 ( \5331 , \5006 , \5007 );
and \U$5174 ( \5332 , \5007 , \5015 );
and \U$5175 ( \5333 , \5006 , \5015 );
or \U$5176 ( \5334 , \5331 , \5332 , \5333 );
xor \U$5177 ( \5335 , \5330 , \5334 );
xor \U$5178 ( \5336 , \5321 , \5335 );
xor \U$5179 ( \5337 , \5312 , \5336 );
xor \U$5180 ( \5338 , \5298 , \5337 );
and \U$5181 ( \5339 , \4902 , \4937 );
and \U$5182 ( \5340 , \4937 , \5109 );
and \U$5183 ( \5341 , \4902 , \5109 );
or \U$5184 ( \5342 , \5339 , \5340 , \5341 );
xor \U$5185 ( \5343 , \5338 , \5342 );
and \U$5186 ( \5344 , \5110 , \5111 );
and \U$5187 ( \5345 , \5112 , \5115 );
or \U$5188 ( \5346 , \5344 , \5345 );
xor \U$5189 ( \5347 , \5343 , \5346 );
buf g5543_GF_PartitionCandidate( \5348_nG5543 , \5347 );
buf \U$5190 ( \5349 , \5348_nG5543 );
and \U$5191 ( \5350 , \5126 , \5130 );
and \U$5192 ( \5351 , \5130 , \5296 );
and \U$5193 ( \5352 , \5126 , \5296 );
or \U$5194 ( \5353 , \5350 , \5351 , \5352 );
and \U$5195 ( \5354 , \5312 , \5336 );
xor \U$5196 ( \5355 , \5353 , \5354 );
and \U$5197 ( \5356 , \5316 , \5320 );
and \U$5198 ( \5357 , \5320 , \5335 );
and \U$5199 ( \5358 , \5316 , \5335 );
or \U$5200 ( \5359 , \5356 , \5357 , \5358 );
and \U$5201 ( \5360 , \5302 , \5306 );
and \U$5202 ( \5361 , \5306 , \5311 );
and \U$5203 ( \5362 , \5302 , \5311 );
or \U$5204 ( \5363 , \5360 , \5361 , \5362 );
and \U$5205 ( \5364 , \5145 , \5201 );
and \U$5206 ( \5365 , \5201 , \5295 );
and \U$5207 ( \5366 , \5145 , \5295 );
or \U$5208 ( \5367 , \5364 , \5365 , \5366 );
xor \U$5209 ( \5368 , \5363 , \5367 );
and \U$5210 ( \5369 , \5135 , \5139 );
and \U$5211 ( \5370 , \5139 , \5144 );
and \U$5212 ( \5371 , \5135 , \5144 );
or \U$5213 ( \5372 , \5369 , \5370 , \5371 );
and \U$5214 ( \5373 , \5206 , \5210 );
and \U$5215 ( \5374 , \5210 , \5215 );
and \U$5216 ( \5375 , \5206 , \5215 );
or \U$5217 ( \5376 , \5373 , \5374 , \5375 );
xor \U$5218 ( \5377 , \5372 , \5376 );
and \U$5219 ( \5378 , \5265 , \5278 );
and \U$5220 ( \5379 , \5278 , \5293 );
and \U$5221 ( \5380 , \5265 , \5293 );
or \U$5222 ( \5381 , \5378 , \5379 , \5380 );
xor \U$5223 ( \5382 , \5377 , \5381 );
xor \U$5224 ( \5383 , \5368 , \5382 );
xor \U$5225 ( \5384 , \5359 , \5383 );
and \U$5226 ( \5385 , \5325 , \5329 );
and \U$5227 ( \5386 , \5329 , \5334 );
and \U$5228 ( \5387 , \5325 , \5334 );
or \U$5229 ( \5388 , \5385 , \5386 , \5387 );
and \U$5230 ( \5389 , \5149 , \5153 );
and \U$5231 ( \5390 , \5153 , \5200 );
and \U$5232 ( \5391 , \5149 , \5200 );
or \U$5233 ( \5392 , \5389 , \5390 , \5391 );
xor \U$5234 ( \5393 , \5388 , \5392 );
and \U$5235 ( \5394 , \5216 , \5260 );
and \U$5236 ( \5395 , \5260 , \5294 );
and \U$5237 ( \5396 , \5216 , \5294 );
or \U$5238 ( \5397 , \5394 , \5395 , \5396 );
xor \U$5239 ( \5398 , \5393 , \5397 );
and \U$5240 ( \5399 , \5159 , \5163 );
and \U$5241 ( \5400 , \5163 , \5169 );
and \U$5242 ( \5401 , \5159 , \5169 );
or \U$5243 ( \5402 , \5399 , \5400 , \5401 );
and \U$5244 ( \5403 , \5174 , \5178 );
and \U$5245 ( \5404 , \5178 , \5183 );
and \U$5246 ( \5405 , \5174 , \5183 );
or \U$5247 ( \5406 , \5403 , \5404 , \5405 );
xor \U$5248 ( \5407 , \5402 , \5406 );
and \U$5249 ( \5408 , \5189 , \5193 );
and \U$5250 ( \5409 , \5193 , \5198 );
and \U$5251 ( \5410 , \5189 , \5198 );
or \U$5252 ( \5411 , \5408 , \5409 , \5410 );
xor \U$5253 ( \5412 , \5407 , \5411 );
and \U$5254 ( \5413 , \5220 , \5224 );
and \U$5255 ( \5414 , \5224 , \5229 );
and \U$5256 ( \5415 , \5220 , \5229 );
or \U$5257 ( \5416 , \5413 , \5414 , \5415 );
and \U$5258 ( \5417 , \5234 , \5238 );
and \U$5259 ( \5418 , \5238 , \5243 );
and \U$5260 ( \5419 , \5234 , \5243 );
or \U$5261 ( \5420 , \5417 , \5418 , \5419 );
xor \U$5262 ( \5421 , \5416 , \5420 );
and \U$5263 ( \5422 , \5249 , \5253 );
and \U$5264 ( \5423 , \5253 , \5258 );
and \U$5265 ( \5424 , \5249 , \5258 );
or \U$5266 ( \5425 , \5422 , \5423 , \5424 );
xor \U$5267 ( \5426 , \5421 , \5425 );
xor \U$5268 ( \5427 , \5412 , \5426 );
and \U$5269 ( \5428 , \5269 , \5273 );
and \U$5270 ( \5429 , \5273 , \5277 );
and \U$5271 ( \5430 , \5269 , \5277 );
or \U$5272 ( \5431 , \5428 , \5429 , \5430 );
and \U$5273 ( \5432 , \5283 , \5287 );
and \U$5274 ( \5433 , \5287 , \5292 );
and \U$5275 ( \5434 , \5283 , \5292 );
or \U$5276 ( \5435 , \5432 , \5433 , \5434 );
xor \U$5277 ( \5436 , \5431 , \5435 );
and \U$5278 ( \5437 , \158 , \5011 );
and \U$5279 ( \5438 , \134 , \4878 );
nor \U$5280 ( \5439 , \5437 , \5438 );
xnor \U$5281 ( \5440 , \5439 , \4762 );
xor \U$5282 ( \5441 , \5436 , \5440 );
xor \U$5283 ( \5442 , \5427 , \5441 );
and \U$5284 ( \5443 , \5230 , \5244 );
and \U$5285 ( \5444 , \5244 , \5259 );
and \U$5286 ( \5445 , \5230 , \5259 );
or \U$5287 ( \5446 , \5443 , \5444 , \5445 );
and \U$5288 ( \5447 , \5170 , \5184 );
and \U$5289 ( \5448 , \5184 , \5199 );
and \U$5290 ( \5449 , \5170 , \5199 );
or \U$5291 ( \5450 , \5447 , \5448 , \5449 );
xor \U$5292 ( \5451 , \5446 , \5450 );
and \U$5293 ( \5452 , \3912 , \230 );
and \U$5294 ( \5453 , \4160 , \228 );
nor \U$5295 ( \5454 , \5452 , \5453 );
xnor \U$5296 ( \5455 , \5454 , \237 );
and \U$5297 ( \5456 , \3646 , \245 );
and \U$5298 ( \5457 , \3736 , \243 );
nor \U$5299 ( \5458 , \5456 , \5457 );
xnor \U$5300 ( \5459 , \5458 , \252 );
xor \U$5301 ( \5460 , \5455 , \5459 );
and \U$5302 ( \5461 , \3143 , \141 );
and \U$5303 ( \5462 , \3395 , \139 );
nor \U$5304 ( \5463 , \5461 , \5462 );
xnor \U$5305 ( \5464 , \5463 , \148 );
xor \U$5306 ( \5465 , \5460 , \5464 );
xor \U$5307 ( \5466 , \5451 , \5465 );
xor \U$5308 ( \5467 , \5442 , \5466 );
and \U$5309 ( \5468 , \5156 , \183 );
buf \U$5310 ( \5469 , RIb55e950_83);
and \U$5311 ( \5470 , \5469 , \180 );
nor \U$5312 ( \5471 , \5468 , \5470 );
xnor \U$5313 ( \5472 , \5471 , \179 );
and \U$5314 ( \5473 , \4749 , \195 );
and \U$5315 ( \5474 , \4922 , \193 );
nor \U$5316 ( \5475 , \5473 , \5474 );
xnor \U$5317 ( \5476 , \5475 , \202 );
xor \U$5318 ( \5477 , \5472 , \5476 );
and \U$5319 ( \5478 , \4364 , \215 );
and \U$5320 ( \5479 , \4654 , \213 );
nor \U$5321 ( \5480 , \5478 , \5479 );
xnor \U$5322 ( \5481 , \5480 , \222 );
xor \U$5323 ( \5482 , \5477 , \5481 );
xor \U$5324 ( \5483 , \5165 , \5166 );
not \U$5325 ( \5484 , \5275 );
and \U$5326 ( \5485 , \5483 , \5484 );
and \U$5327 ( \5486 , \166 , \5485 );
and \U$5328 ( \5487 , \150 , \5275 );
nor \U$5329 ( \5488 , \5486 , \5487 );
xnor \U$5330 ( \5489 , \5488 , \5169 );
and \U$5331 ( \5490 , \185 , \2669 );
and \U$5332 ( \5491 , \261 , \2538 );
nor \U$5333 ( \5492 , \5490 , \5491 );
xnor \U$5334 ( \5493 , \5492 , \2534 );
and \U$5335 ( \5494 , \197 , \3103 );
and \U$5336 ( \5495 , \178 , \2934 );
nor \U$5337 ( \5496 , \5494 , \5495 );
xnor \U$5338 ( \5497 , \5496 , \2839 );
xor \U$5339 ( \5498 , \5493 , \5497 );
and \U$5340 ( \5499 , \217 , \3357 );
and \U$5341 ( \5500 , \189 , \3255 );
nor \U$5342 ( \5501 , \5499 , \5500 );
xnor \U$5343 ( \5502 , \5501 , \3156 );
xor \U$5344 ( \5503 , \5498 , \5502 );
xor \U$5345 ( \5504 , \5489 , \5503 );
and \U$5346 ( \5505 , \232 , \3813 );
and \U$5347 ( \5506 , \209 , \3557 );
nor \U$5348 ( \5507 , \5505 , \5506 );
xnor \U$5349 ( \5508 , \5507 , \3562 );
and \U$5350 ( \5509 , \247 , \4132 );
and \U$5351 ( \5510 , \224 , \4012 );
nor \U$5352 ( \5511 , \5509 , \5510 );
xnor \U$5353 ( \5512 , \5511 , \3925 );
xor \U$5354 ( \5513 , \5508 , \5512 );
and \U$5355 ( \5514 , \143 , \4581 );
and \U$5356 ( \5515 , \240 , \4424 );
nor \U$5357 ( \5516 , \5514 , \5515 );
xnor \U$5358 ( \5517 , \5516 , \4377 );
xor \U$5359 ( \5518 , \5513 , \5517 );
xor \U$5360 ( \5519 , \5504 , \5518 );
xor \U$5361 ( \5520 , \5482 , \5519 );
and \U$5362 ( \5521 , \1948 , \1086 );
and \U$5363 ( \5522 , \2090 , \508 );
nor \U$5364 ( \5523 , \5521 , \5522 );
xnor \U$5365 ( \5524 , \5523 , \487 );
and \U$5366 ( \5525 , \1684 , \1301 );
and \U$5367 ( \5526 , \1802 , \1246 );
nor \U$5368 ( \5527 , \5525 , \5526 );
xnor \U$5369 ( \5528 , \5527 , \1205 );
xor \U$5370 ( \5529 , \5524 , \5528 );
and \U$5371 ( \5530 , \1484 , \1578 );
and \U$5372 ( \5531 , \1601 , \1431 );
nor \U$5373 ( \5532 , \5530 , \5531 );
xnor \U$5374 ( \5533 , \5532 , \1436 );
xor \U$5375 ( \5534 , \5529 , \5533 );
and \U$5376 ( \5535 , \1192 , \1824 );
and \U$5377 ( \5536 , \1333 , \1739 );
nor \U$5378 ( \5537 , \5535 , \5536 );
xnor \U$5379 ( \5538 , \5537 , \1697 );
and \U$5380 ( \5539 , \474 , \2121 );
and \U$5381 ( \5540 , \1147 , \2008 );
nor \U$5382 ( \5541 , \5539 , \5540 );
xnor \U$5383 ( \5542 , \5541 , \1961 );
xor \U$5384 ( \5543 , \5538 , \5542 );
and \U$5385 ( \5544 , \307 , \2400 );
and \U$5386 ( \5545 , \412 , \2246 );
nor \U$5387 ( \5546 , \5544 , \5545 );
xnor \U$5388 ( \5547 , \5546 , \2195 );
xor \U$5389 ( \5548 , \5543 , \5547 );
xor \U$5390 ( \5549 , \5534 , \5548 );
and \U$5391 ( \5550 , \2826 , \156 );
and \U$5392 ( \5551 , \3037 , \154 );
nor \U$5393 ( \5552 , \5550 , \5551 );
xnor \U$5394 ( \5553 , \5552 , \163 );
and \U$5395 ( \5554 , \2521 , \296 );
and \U$5396 ( \5555 , \2757 , \168 );
nor \U$5397 ( \5556 , \5554 , \5555 );
xnor \U$5398 ( \5557 , \5556 , \173 );
xor \U$5399 ( \5558 , \5553 , \5557 );
and \U$5400 ( \5559 , \2182 , \438 );
and \U$5401 ( \5560 , \2366 , \336 );
nor \U$5402 ( \5561 , \5559 , \5560 );
xnor \U$5403 ( \5562 , \5561 , \320 );
xor \U$5404 ( \5563 , \5558 , \5562 );
xor \U$5405 ( \5564 , \5549 , \5563 );
xor \U$5406 ( \5565 , \5520 , \5564 );
xor \U$5407 ( \5566 , \5467 , \5565 );
xor \U$5408 ( \5567 , \5398 , \5566 );
xor \U$5409 ( \5568 , \5384 , \5567 );
xor \U$5410 ( \5569 , \5355 , \5568 );
and \U$5411 ( \5570 , \5122 , \5297 );
and \U$5412 ( \5571 , \5297 , \5337 );
and \U$5413 ( \5572 , \5122 , \5337 );
or \U$5414 ( \5573 , \5570 , \5571 , \5572 );
xor \U$5415 ( \5574 , \5569 , \5573 );
and \U$5416 ( \5575 , \5338 , \5342 );
and \U$5417 ( \5576 , \5343 , \5346 );
or \U$5418 ( \5577 , \5575 , \5576 );
xor \U$5419 ( \5578 , \5574 , \5577 );
buf g5541_GF_PartitionCandidate( \5579_nG5541 , \5578 );
buf \U$5420 ( \5580 , \5579_nG5541 );
and \U$5421 ( \5581 , \5359 , \5383 );
and \U$5422 ( \5582 , \5383 , \5567 );
and \U$5423 ( \5583 , \5359 , \5567 );
or \U$5424 ( \5584 , \5581 , \5582 , \5583 );
and \U$5425 ( \5585 , \5363 , \5367 );
and \U$5426 ( \5586 , \5367 , \5382 );
and \U$5427 ( \5587 , \5363 , \5382 );
or \U$5428 ( \5588 , \5585 , \5586 , \5587 );
and \U$5429 ( \5589 , \5398 , \5566 );
xor \U$5430 ( \5590 , \5588 , \5589 );
and \U$5431 ( \5591 , \5412 , \5426 );
and \U$5432 ( \5592 , \5426 , \5441 );
and \U$5433 ( \5593 , \5412 , \5441 );
or \U$5434 ( \5594 , \5591 , \5592 , \5593 );
and \U$5435 ( \5595 , \5524 , \5528 );
and \U$5436 ( \5596 , \5528 , \5533 );
and \U$5437 ( \5597 , \5524 , \5533 );
or \U$5438 ( \5598 , \5595 , \5596 , \5597 );
and \U$5439 ( \5599 , \5538 , \5542 );
and \U$5440 ( \5600 , \5542 , \5547 );
and \U$5441 ( \5601 , \5538 , \5547 );
or \U$5442 ( \5602 , \5599 , \5600 , \5601 );
xor \U$5443 ( \5603 , \5598 , \5602 );
and \U$5444 ( \5604 , \5493 , \5497 );
and \U$5445 ( \5605 , \5497 , \5502 );
and \U$5446 ( \5606 , \5493 , \5502 );
or \U$5447 ( \5607 , \5604 , \5605 , \5606 );
xor \U$5448 ( \5608 , \5603 , \5607 );
xor \U$5449 ( \5609 , \5594 , \5608 );
and \U$5450 ( \5610 , \5455 , \5459 );
and \U$5451 ( \5611 , \5459 , \5464 );
and \U$5452 ( \5612 , \5455 , \5464 );
or \U$5453 ( \5613 , \5610 , \5611 , \5612 );
and \U$5454 ( \5614 , \5553 , \5557 );
and \U$5455 ( \5615 , \5557 , \5562 );
and \U$5456 ( \5616 , \5553 , \5562 );
or \U$5457 ( \5617 , \5614 , \5615 , \5616 );
xor \U$5458 ( \5618 , \5613 , \5617 );
and \U$5459 ( \5619 , \5472 , \5476 );
and \U$5460 ( \5620 , \5476 , \5481 );
and \U$5461 ( \5621 , \5472 , \5481 );
or \U$5462 ( \5622 , \5619 , \5620 , \5621 );
xor \U$5463 ( \5623 , \5618 , \5622 );
xor \U$5464 ( \5624 , \5609 , \5623 );
xor \U$5465 ( \5625 , \5590 , \5624 );
xor \U$5466 ( \5626 , \5584 , \5625 );
and \U$5467 ( \5627 , \5372 , \5376 );
and \U$5468 ( \5628 , \5376 , \5381 );
and \U$5469 ( \5629 , \5372 , \5381 );
or \U$5470 ( \5630 , \5627 , \5628 , \5629 );
and \U$5471 ( \5631 , \5446 , \5450 );
and \U$5472 ( \5632 , \5450 , \5465 );
and \U$5473 ( \5633 , \5446 , \5465 );
or \U$5474 ( \5634 , \5631 , \5632 , \5633 );
xor \U$5475 ( \5635 , \5630 , \5634 );
and \U$5476 ( \5636 , \5482 , \5519 );
and \U$5477 ( \5637 , \5519 , \5564 );
and \U$5478 ( \5638 , \5482 , \5564 );
or \U$5479 ( \5639 , \5636 , \5637 , \5638 );
xor \U$5480 ( \5640 , \5635 , \5639 );
and \U$5481 ( \5641 , \5388 , \5392 );
and \U$5482 ( \5642 , \5392 , \5397 );
and \U$5483 ( \5643 , \5388 , \5397 );
or \U$5484 ( \5644 , \5641 , \5642 , \5643 );
and \U$5485 ( \5645 , \5442 , \5466 );
and \U$5486 ( \5646 , \5466 , \5565 );
and \U$5487 ( \5647 , \5442 , \5565 );
or \U$5488 ( \5648 , \5645 , \5646 , \5647 );
xor \U$5489 ( \5649 , \5644 , \5648 );
and \U$5490 ( \5650 , \5402 , \5406 );
and \U$5491 ( \5651 , \5406 , \5411 );
and \U$5492 ( \5652 , \5402 , \5411 );
or \U$5493 ( \5653 , \5650 , \5651 , \5652 );
and \U$5494 ( \5654 , \5416 , \5420 );
and \U$5495 ( \5655 , \5420 , \5425 );
and \U$5496 ( \5656 , \5416 , \5425 );
or \U$5497 ( \5657 , \5654 , \5655 , \5656 );
xor \U$5498 ( \5658 , \5653 , \5657 );
and \U$5499 ( \5659 , \5431 , \5435 );
and \U$5500 ( \5660 , \5435 , \5440 );
and \U$5501 ( \5661 , \5431 , \5440 );
or \U$5502 ( \5662 , \5659 , \5660 , \5661 );
xor \U$5503 ( \5663 , \5658 , \5662 );
and \U$5504 ( \5664 , \5489 , \5503 );
and \U$5505 ( \5665 , \5503 , \5518 );
and \U$5506 ( \5666 , \5489 , \5518 );
or \U$5507 ( \5667 , \5664 , \5665 , \5666 );
and \U$5508 ( \5668 , \5534 , \5548 );
and \U$5509 ( \5669 , \5548 , \5563 );
and \U$5510 ( \5670 , \5534 , \5563 );
or \U$5511 ( \5671 , \5668 , \5669 , \5670 );
xor \U$5512 ( \5672 , \5667 , \5671 );
and \U$5513 ( \5673 , \5469 , \183 );
buf \U$5514 ( \5674 , RIb55e9c8_82);
and \U$5515 ( \5675 , \5674 , \180 );
nor \U$5516 ( \5676 , \5673 , \5675 );
xnor \U$5517 ( \5677 , \5676 , \179 );
and \U$5518 ( \5678 , \4922 , \195 );
and \U$5519 ( \5679 , \5156 , \193 );
nor \U$5520 ( \5680 , \5678 , \5679 );
xnor \U$5521 ( \5681 , \5680 , \202 );
xor \U$5522 ( \5682 , \5677 , \5681 );
buf \U$5523 ( \5683 , RIb560840_17);
buf \U$5524 ( \5684 , RIb5607c8_18);
and \U$5525 ( \5685 , \5684 , \5165 );
not \U$5526 ( \5686 , \5685 );
and \U$5527 ( \5687 , \5683 , \5686 );
xor \U$5528 ( \5688 , \5682 , \5687 );
xor \U$5529 ( \5689 , \5672 , \5688 );
xor \U$5530 ( \5690 , \5663 , \5689 );
and \U$5531 ( \5691 , \5508 , \5512 );
and \U$5532 ( \5692 , \5512 , \5517 );
and \U$5533 ( \5693 , \5508 , \5517 );
or \U$5534 ( \5694 , \5691 , \5692 , \5693 );
xor \U$5535 ( \5695 , \5684 , \5165 );
nand \U$5536 ( \5696 , \166 , \5695 );
xnor \U$5537 ( \5697 , \5696 , \5687 );
xor \U$5538 ( \5698 , \5694 , \5697 );
and \U$5539 ( \5699 , \240 , \4581 );
and \U$5540 ( \5700 , \247 , \4424 );
nor \U$5541 ( \5701 , \5699 , \5700 );
xnor \U$5542 ( \5702 , \5701 , \4377 );
and \U$5543 ( \5703 , \134 , \5011 );
and \U$5544 ( \5704 , \143 , \4878 );
nor \U$5545 ( \5705 , \5703 , \5704 );
xnor \U$5546 ( \5706 , \5705 , \4762 );
xor \U$5547 ( \5707 , \5702 , \5706 );
and \U$5548 ( \5708 , \150 , \5485 );
and \U$5549 ( \5709 , \158 , \5275 );
nor \U$5550 ( \5710 , \5708 , \5709 );
xnor \U$5551 ( \5711 , \5710 , \5169 );
xor \U$5552 ( \5712 , \5707 , \5711 );
xor \U$5553 ( \5713 , \5698 , \5712 );
and \U$5554 ( \5714 , \412 , \2400 );
and \U$5555 ( \5715 , \474 , \2246 );
nor \U$5556 ( \5716 , \5714 , \5715 );
xnor \U$5557 ( \5717 , \5716 , \2195 );
and \U$5558 ( \5718 , \261 , \2669 );
and \U$5559 ( \5719 , \307 , \2538 );
nor \U$5560 ( \5720 , \5718 , \5719 );
xnor \U$5561 ( \5721 , \5720 , \2534 );
xor \U$5562 ( \5722 , \5717 , \5721 );
and \U$5563 ( \5723 , \178 , \3103 );
and \U$5564 ( \5724 , \185 , \2934 );
nor \U$5565 ( \5725 , \5723 , \5724 );
xnor \U$5566 ( \5726 , \5725 , \2839 );
xor \U$5567 ( \5727 , \5722 , \5726 );
and \U$5568 ( \5728 , \189 , \3357 );
and \U$5569 ( \5729 , \197 , \3255 );
nor \U$5570 ( \5730 , \5728 , \5729 );
xnor \U$5571 ( \5731 , \5730 , \3156 );
and \U$5572 ( \5732 , \209 , \3813 );
and \U$5573 ( \5733 , \217 , \3557 );
nor \U$5574 ( \5734 , \5732 , \5733 );
xnor \U$5575 ( \5735 , \5734 , \3562 );
xor \U$5576 ( \5736 , \5731 , \5735 );
and \U$5577 ( \5737 , \224 , \4132 );
and \U$5578 ( \5738 , \232 , \4012 );
nor \U$5579 ( \5739 , \5737 , \5738 );
xnor \U$5580 ( \5740 , \5739 , \3925 );
xor \U$5581 ( \5741 , \5736 , \5740 );
xor \U$5582 ( \5742 , \5727 , \5741 );
and \U$5583 ( \5743 , \1601 , \1578 );
and \U$5584 ( \5744 , \1684 , \1431 );
nor \U$5585 ( \5745 , \5743 , \5744 );
xnor \U$5586 ( \5746 , \5745 , \1436 );
and \U$5587 ( \5747 , \1333 , \1824 );
and \U$5588 ( \5748 , \1484 , \1739 );
nor \U$5589 ( \5749 , \5747 , \5748 );
xnor \U$5590 ( \5750 , \5749 , \1697 );
xor \U$5591 ( \5751 , \5746 , \5750 );
and \U$5592 ( \5752 , \1147 , \2121 );
and \U$5593 ( \5753 , \1192 , \2008 );
nor \U$5594 ( \5754 , \5752 , \5753 );
xnor \U$5595 ( \5755 , \5754 , \1961 );
xor \U$5596 ( \5756 , \5751 , \5755 );
xor \U$5597 ( \5757 , \5742 , \5756 );
xor \U$5598 ( \5758 , \5713 , \5757 );
and \U$5599 ( \5759 , \4654 , \215 );
and \U$5600 ( \5760 , \4749 , \213 );
nor \U$5601 ( \5761 , \5759 , \5760 );
xnor \U$5602 ( \5762 , \5761 , \222 );
and \U$5603 ( \5763 , \4160 , \230 );
and \U$5604 ( \5764 , \4364 , \228 );
nor \U$5605 ( \5765 , \5763 , \5764 );
xnor \U$5606 ( \5766 , \5765 , \237 );
xor \U$5607 ( \5767 , \5762 , \5766 );
and \U$5608 ( \5768 , \3736 , \245 );
and \U$5609 ( \5769 , \3912 , \243 );
nor \U$5610 ( \5770 , \5768 , \5769 );
xnor \U$5611 ( \5771 , \5770 , \252 );
xor \U$5612 ( \5772 , \5767 , \5771 );
and \U$5613 ( \5773 , \2366 , \438 );
and \U$5614 ( \5774 , \2521 , \336 );
nor \U$5615 ( \5775 , \5773 , \5774 );
xnor \U$5616 ( \5776 , \5775 , \320 );
and \U$5617 ( \5777 , \2090 , \1086 );
and \U$5618 ( \5778 , \2182 , \508 );
nor \U$5619 ( \5779 , \5777 , \5778 );
xnor \U$5620 ( \5780 , \5779 , \487 );
xor \U$5621 ( \5781 , \5776 , \5780 );
and \U$5622 ( \5782 , \1802 , \1301 );
and \U$5623 ( \5783 , \1948 , \1246 );
nor \U$5624 ( \5784 , \5782 , \5783 );
xnor \U$5625 ( \5785 , \5784 , \1205 );
xor \U$5626 ( \5786 , \5781 , \5785 );
xor \U$5627 ( \5787 , \5772 , \5786 );
and \U$5628 ( \5788 , \3395 , \141 );
and \U$5629 ( \5789 , \3646 , \139 );
nor \U$5630 ( \5790 , \5788 , \5789 );
xnor \U$5631 ( \5791 , \5790 , \148 );
and \U$5632 ( \5792 , \3037 , \156 );
and \U$5633 ( \5793 , \3143 , \154 );
nor \U$5634 ( \5794 , \5792 , \5793 );
xnor \U$5635 ( \5795 , \5794 , \163 );
xor \U$5636 ( \5796 , \5791 , \5795 );
and \U$5637 ( \5797 , \2757 , \296 );
and \U$5638 ( \5798 , \2826 , \168 );
nor \U$5639 ( \5799 , \5797 , \5798 );
xnor \U$5640 ( \5800 , \5799 , \173 );
xor \U$5641 ( \5801 , \5796 , \5800 );
xor \U$5642 ( \5802 , \5787 , \5801 );
xor \U$5643 ( \5803 , \5758 , \5802 );
xor \U$5644 ( \5804 , \5690 , \5803 );
xor \U$5645 ( \5805 , \5649 , \5804 );
xor \U$5646 ( \5806 , \5640 , \5805 );
xor \U$5647 ( \5807 , \5626 , \5806 );
and \U$5648 ( \5808 , \5353 , \5354 );
and \U$5649 ( \5809 , \5354 , \5568 );
and \U$5650 ( \5810 , \5353 , \5568 );
or \U$5651 ( \5811 , \5808 , \5809 , \5810 );
xor \U$5652 ( \5812 , \5807 , \5811 );
and \U$5653 ( \5813 , \5569 , \5573 );
and \U$5654 ( \5814 , \5574 , \5577 );
or \U$5655 ( \5815 , \5813 , \5814 );
xor \U$5656 ( \5816 , \5812 , \5815 );
buf g553f_GF_PartitionCandidate( \5817_nG553f , \5816 );
buf \U$5657 ( \5818 , \5817_nG553f );
and \U$5658 ( \5819 , \5588 , \5589 );
and \U$5659 ( \5820 , \5589 , \5624 );
and \U$5660 ( \5821 , \5588 , \5624 );
or \U$5661 ( \5822 , \5819 , \5820 , \5821 );
and \U$5662 ( \5823 , \5640 , \5805 );
xor \U$5663 ( \5824 , \5822 , \5823 );
and \U$5664 ( \5825 , \5644 , \5648 );
and \U$5665 ( \5826 , \5648 , \5804 );
and \U$5666 ( \5827 , \5644 , \5804 );
or \U$5667 ( \5828 , \5825 , \5826 , \5827 );
and \U$5668 ( \5829 , \5630 , \5634 );
and \U$5669 ( \5830 , \5634 , \5639 );
and \U$5670 ( \5831 , \5630 , \5639 );
or \U$5671 ( \5832 , \5829 , \5830 , \5831 );
and \U$5672 ( \5833 , \5594 , \5608 );
and \U$5673 ( \5834 , \5608 , \5623 );
and \U$5674 ( \5835 , \5594 , \5623 );
or \U$5675 ( \5836 , \5833 , \5834 , \5835 );
xor \U$5676 ( \5837 , \5832 , \5836 );
and \U$5677 ( \5838 , \5663 , \5689 );
and \U$5678 ( \5839 , \5689 , \5803 );
and \U$5679 ( \5840 , \5663 , \5803 );
or \U$5680 ( \5841 , \5838 , \5839 , \5840 );
xor \U$5681 ( \5842 , \5837 , \5841 );
xor \U$5682 ( \5843 , \5828 , \5842 );
and \U$5683 ( \5844 , \5653 , \5657 );
and \U$5684 ( \5845 , \5657 , \5662 );
and \U$5685 ( \5846 , \5653 , \5662 );
or \U$5686 ( \5847 , \5844 , \5845 , \5846 );
and \U$5687 ( \5848 , \5667 , \5671 );
and \U$5688 ( \5849 , \5671 , \5688 );
and \U$5689 ( \5850 , \5667 , \5688 );
or \U$5690 ( \5851 , \5848 , \5849 , \5850 );
xor \U$5691 ( \5852 , \5847 , \5851 );
and \U$5692 ( \5853 , \5713 , \5757 );
and \U$5693 ( \5854 , \5757 , \5802 );
and \U$5694 ( \5855 , \5713 , \5802 );
or \U$5695 ( \5856 , \5853 , \5854 , \5855 );
xor \U$5696 ( \5857 , \5852 , \5856 );
and \U$5697 ( \5858 , \5717 , \5721 );
and \U$5698 ( \5859 , \5721 , \5726 );
and \U$5699 ( \5860 , \5717 , \5726 );
or \U$5700 ( \5861 , \5858 , \5859 , \5860 );
and \U$5701 ( \5862 , \5746 , \5750 );
and \U$5702 ( \5863 , \5750 , \5755 );
and \U$5703 ( \5864 , \5746 , \5755 );
or \U$5704 ( \5865 , \5862 , \5863 , \5864 );
xor \U$5705 ( \5866 , \5861 , \5865 );
and \U$5706 ( \5867 , \5776 , \5780 );
and \U$5707 ( \5868 , \5780 , \5785 );
and \U$5708 ( \5869 , \5776 , \5785 );
or \U$5709 ( \5870 , \5867 , \5868 , \5869 );
xor \U$5710 ( \5871 , \5866 , \5870 );
and \U$5711 ( \5872 , \5762 , \5766 );
and \U$5712 ( \5873 , \5766 , \5771 );
and \U$5713 ( \5874 , \5762 , \5771 );
or \U$5714 ( \5875 , \5872 , \5873 , \5874 );
and \U$5715 ( \5876 , \5677 , \5681 );
and \U$5716 ( \5877 , \5681 , \5687 );
and \U$5717 ( \5878 , \5677 , \5687 );
or \U$5718 ( \5879 , \5876 , \5877 , \5878 );
xor \U$5719 ( \5880 , \5875 , \5879 );
and \U$5720 ( \5881 , \5791 , \5795 );
and \U$5721 ( \5882 , \5795 , \5800 );
and \U$5722 ( \5883 , \5791 , \5800 );
or \U$5723 ( \5884 , \5881 , \5882 , \5883 );
xor \U$5724 ( \5885 , \5880 , \5884 );
xor \U$5725 ( \5886 , \5871 , \5885 );
and \U$5726 ( \5887 , \217 , \3813 );
and \U$5727 ( \5888 , \189 , \3557 );
nor \U$5728 ( \5889 , \5887 , \5888 );
xnor \U$5729 ( \5890 , \5889 , \3562 );
and \U$5730 ( \5891 , \232 , \4132 );
and \U$5731 ( \5892 , \209 , \4012 );
nor \U$5732 ( \5893 , \5891 , \5892 );
xnor \U$5733 ( \5894 , \5893 , \3925 );
xor \U$5734 ( \5895 , \5890 , \5894 );
and \U$5735 ( \5896 , \247 , \4581 );
and \U$5736 ( \5897 , \224 , \4424 );
nor \U$5737 ( \5898 , \5896 , \5897 );
xnor \U$5738 ( \5899 , \5898 , \4377 );
xor \U$5739 ( \5900 , \5895 , \5899 );
and \U$5740 ( \5901 , \1484 , \1824 );
and \U$5741 ( \5902 , \1601 , \1739 );
nor \U$5742 ( \5903 , \5901 , \5902 );
xnor \U$5743 ( \5904 , \5903 , \1697 );
and \U$5744 ( \5905 , \1192 , \2121 );
and \U$5745 ( \5906 , \1333 , \2008 );
nor \U$5746 ( \5907 , \5905 , \5906 );
xnor \U$5747 ( \5908 , \5907 , \1961 );
xor \U$5748 ( \5909 , \5904 , \5908 );
and \U$5749 ( \5910 , \474 , \2400 );
and \U$5750 ( \5911 , \1147 , \2246 );
nor \U$5751 ( \5912 , \5910 , \5911 );
xnor \U$5752 ( \5913 , \5912 , \2195 );
xor \U$5753 ( \5914 , \5909 , \5913 );
xor \U$5754 ( \5915 , \5900 , \5914 );
and \U$5755 ( \5916 , \307 , \2669 );
and \U$5756 ( \5917 , \412 , \2538 );
nor \U$5757 ( \5918 , \5916 , \5917 );
xnor \U$5758 ( \5919 , \5918 , \2534 );
and \U$5759 ( \5920 , \185 , \3103 );
and \U$5760 ( \5921 , \261 , \2934 );
nor \U$5761 ( \5922 , \5920 , \5921 );
xnor \U$5762 ( \5923 , \5922 , \2839 );
xor \U$5763 ( \5924 , \5919 , \5923 );
and \U$5764 ( \5925 , \197 , \3357 );
and \U$5765 ( \5926 , \178 , \3255 );
nor \U$5766 ( \5927 , \5925 , \5926 );
xnor \U$5767 ( \5928 , \5927 , \3156 );
xor \U$5768 ( \5929 , \5924 , \5928 );
xor \U$5769 ( \5930 , \5915 , \5929 );
and \U$5770 ( \5931 , \4364 , \230 );
and \U$5771 ( \5932 , \4654 , \228 );
nor \U$5772 ( \5933 , \5931 , \5932 );
xnor \U$5773 ( \5934 , \5933 , \237 );
and \U$5774 ( \5935 , \3912 , \245 );
and \U$5775 ( \5936 , \4160 , \243 );
nor \U$5776 ( \5937 , \5935 , \5936 );
xnor \U$5777 ( \5938 , \5937 , \252 );
xor \U$5778 ( \5939 , \5934 , \5938 );
and \U$5779 ( \5940 , \3646 , \141 );
and \U$5780 ( \5941 , \3736 , \139 );
nor \U$5781 ( \5942 , \5940 , \5941 );
xnor \U$5782 ( \5943 , \5942 , \148 );
xor \U$5783 ( \5944 , \5939 , \5943 );
and \U$5784 ( \5945 , \2182 , \1086 );
and \U$5785 ( \5946 , \2366 , \508 );
nor \U$5786 ( \5947 , \5945 , \5946 );
xnor \U$5787 ( \5948 , \5947 , \487 );
and \U$5788 ( \5949 , \1948 , \1301 );
and \U$5789 ( \5950 , \2090 , \1246 );
nor \U$5790 ( \5951 , \5949 , \5950 );
xnor \U$5791 ( \5952 , \5951 , \1205 );
xor \U$5792 ( \5953 , \5948 , \5952 );
and \U$5793 ( \5954 , \1684 , \1578 );
and \U$5794 ( \5955 , \1802 , \1431 );
nor \U$5795 ( \5956 , \5954 , \5955 );
xnor \U$5796 ( \5957 , \5956 , \1436 );
xor \U$5797 ( \5958 , \5953 , \5957 );
xor \U$5798 ( \5959 , \5944 , \5958 );
and \U$5799 ( \5960 , \3143 , \156 );
and \U$5800 ( \5961 , \3395 , \154 );
nor \U$5801 ( \5962 , \5960 , \5961 );
xnor \U$5802 ( \5963 , \5962 , \163 );
and \U$5803 ( \5964 , \2826 , \296 );
and \U$5804 ( \5965 , \3037 , \168 );
nor \U$5805 ( \5966 , \5964 , \5965 );
xnor \U$5806 ( \5967 , \5966 , \173 );
xor \U$5807 ( \5968 , \5963 , \5967 );
and \U$5808 ( \5969 , \2521 , \438 );
and \U$5809 ( \5970 , \2757 , \336 );
nor \U$5810 ( \5971 , \5969 , \5970 );
xnor \U$5811 ( \5972 , \5971 , \320 );
xor \U$5812 ( \5973 , \5968 , \5972 );
xor \U$5813 ( \5974 , \5959 , \5973 );
xor \U$5814 ( \5975 , \5930 , \5974 );
and \U$5815 ( \5976 , \5731 , \5735 );
and \U$5816 ( \5977 , \5735 , \5740 );
and \U$5817 ( \5978 , \5731 , \5740 );
or \U$5818 ( \5979 , \5976 , \5977 , \5978 );
and \U$5819 ( \5980 , \5702 , \5706 );
and \U$5820 ( \5981 , \5706 , \5711 );
and \U$5821 ( \5982 , \5702 , \5711 );
or \U$5822 ( \5983 , \5980 , \5981 , \5982 );
xor \U$5823 ( \5984 , \5979 , \5983 );
and \U$5824 ( \5985 , \143 , \5011 );
and \U$5825 ( \5986 , \240 , \4878 );
nor \U$5826 ( \5987 , \5985 , \5986 );
xnor \U$5827 ( \5988 , \5987 , \4762 );
and \U$5828 ( \5989 , \158 , \5485 );
and \U$5829 ( \5990 , \134 , \5275 );
nor \U$5830 ( \5991 , \5989 , \5990 );
xnor \U$5831 ( \5992 , \5991 , \5169 );
xor \U$5832 ( \5993 , \5988 , \5992 );
xor \U$5833 ( \5994 , \5683 , \5684 );
not \U$5834 ( \5995 , \5695 );
and \U$5835 ( \5996 , \5994 , \5995 );
and \U$5836 ( \5997 , \166 , \5996 );
and \U$5837 ( \5998 , \150 , \5695 );
nor \U$5838 ( \5999 , \5997 , \5998 );
xnor \U$5839 ( \6000 , \5999 , \5687 );
xor \U$5840 ( \6001 , \5993 , \6000 );
xor \U$5841 ( \6002 , \5984 , \6001 );
xor \U$5842 ( \6003 , \5975 , \6002 );
xor \U$5843 ( \6004 , \5886 , \6003 );
xor \U$5844 ( \6005 , \5857 , \6004 );
and \U$5845 ( \6006 , \5598 , \5602 );
and \U$5846 ( \6007 , \5602 , \5607 );
and \U$5847 ( \6008 , \5598 , \5607 );
or \U$5848 ( \6009 , \6006 , \6007 , \6008 );
and \U$5849 ( \6010 , \5613 , \5617 );
and \U$5850 ( \6011 , \5617 , \5622 );
and \U$5851 ( \6012 , \5613 , \5622 );
or \U$5852 ( \6013 , \6010 , \6011 , \6012 );
xor \U$5853 ( \6014 , \6009 , \6013 );
and \U$5854 ( \6015 , \5694 , \5697 );
and \U$5855 ( \6016 , \5697 , \5712 );
and \U$5856 ( \6017 , \5694 , \5712 );
or \U$5857 ( \6018 , \6015 , \6016 , \6017 );
xor \U$5858 ( \6019 , \6014 , \6018 );
and \U$5859 ( \6020 , \5727 , \5741 );
and \U$5860 ( \6021 , \5741 , \5756 );
and \U$5861 ( \6022 , \5727 , \5756 );
or \U$5862 ( \6023 , \6020 , \6021 , \6022 );
and \U$5863 ( \6024 , \5772 , \5786 );
and \U$5864 ( \6025 , \5786 , \5801 );
and \U$5865 ( \6026 , \5772 , \5801 );
or \U$5866 ( \6027 , \6024 , \6025 , \6026 );
xor \U$5867 ( \6028 , \6023 , \6027 );
and \U$5868 ( \6029 , \5674 , \183 );
buf \U$5869 ( \6030 , RIb55ea40_81);
and \U$5870 ( \6031 , \6030 , \180 );
nor \U$5871 ( \6032 , \6029 , \6031 );
xnor \U$5872 ( \6033 , \6032 , \179 );
and \U$5873 ( \6034 , \5156 , \195 );
and \U$5874 ( \6035 , \5469 , \193 );
nor \U$5875 ( \6036 , \6034 , \6035 );
xnor \U$5876 ( \6037 , \6036 , \202 );
xor \U$5877 ( \6038 , \6033 , \6037 );
and \U$5878 ( \6039 , \4749 , \215 );
and \U$5879 ( \6040 , \4922 , \213 );
nor \U$5880 ( \6041 , \6039 , \6040 );
xnor \U$5881 ( \6042 , \6041 , \222 );
xor \U$5882 ( \6043 , \6038 , \6042 );
xor \U$5883 ( \6044 , \6028 , \6043 );
xor \U$5884 ( \6045 , \6019 , \6044 );
xor \U$5885 ( \6046 , \6005 , \6045 );
xor \U$5886 ( \6047 , \5843 , \6046 );
xor \U$5887 ( \6048 , \5824 , \6047 );
and \U$5888 ( \6049 , \5584 , \5625 );
and \U$5889 ( \6050 , \5625 , \5806 );
and \U$5890 ( \6051 , \5584 , \5806 );
or \U$5891 ( \6052 , \6049 , \6050 , \6051 );
xor \U$5892 ( \6053 , \6048 , \6052 );
and \U$5893 ( \6054 , \5807 , \5811 );
and \U$5894 ( \6055 , \5812 , \5815 );
or \U$5895 ( \6056 , \6054 , \6055 );
xor \U$5896 ( \6057 , \6053 , \6056 );
buf g553d_GF_PartitionCandidate( \6058_nG553d , \6057 );
buf \U$5897 ( \6059 , \6058_nG553d );
and \U$5898 ( \6060 , \5828 , \5842 );
and \U$5899 ( \6061 , \5842 , \6046 );
and \U$5900 ( \6062 , \5828 , \6046 );
or \U$5901 ( \6063 , \6060 , \6061 , \6062 );
and \U$5902 ( \6064 , \5847 , \5851 );
and \U$5903 ( \6065 , \5851 , \5856 );
and \U$5904 ( \6066 , \5847 , \5856 );
or \U$5905 ( \6067 , \6064 , \6065 , \6066 );
and \U$5906 ( \6068 , \5871 , \5885 );
and \U$5907 ( \6069 , \5885 , \6003 );
and \U$5908 ( \6070 , \5871 , \6003 );
or \U$5909 ( \6071 , \6068 , \6069 , \6070 );
xor \U$5910 ( \6072 , \6067 , \6071 );
and \U$5911 ( \6073 , \6019 , \6044 );
xor \U$5912 ( \6074 , \6072 , \6073 );
xor \U$5913 ( \6075 , \6063 , \6074 );
and \U$5914 ( \6076 , \5832 , \5836 );
and \U$5915 ( \6077 , \5836 , \5841 );
and \U$5916 ( \6078 , \5832 , \5841 );
or \U$5917 ( \6079 , \6076 , \6077 , \6078 );
and \U$5918 ( \6080 , \5857 , \6004 );
and \U$5919 ( \6081 , \6004 , \6045 );
and \U$5920 ( \6082 , \5857 , \6045 );
or \U$5921 ( \6083 , \6080 , \6081 , \6082 );
xor \U$5922 ( \6084 , \6079 , \6083 );
and \U$5923 ( \6085 , \6009 , \6013 );
and \U$5924 ( \6086 , \6013 , \6018 );
and \U$5925 ( \6087 , \6009 , \6018 );
or \U$5926 ( \6088 , \6085 , \6086 , \6087 );
and \U$5927 ( \6089 , \6023 , \6027 );
and \U$5928 ( \6090 , \6027 , \6043 );
and \U$5929 ( \6091 , \6023 , \6043 );
or \U$5930 ( \6092 , \6089 , \6090 , \6091 );
xor \U$5931 ( \6093 , \6088 , \6092 );
and \U$5932 ( \6094 , \5930 , \5974 );
and \U$5933 ( \6095 , \5974 , \6002 );
and \U$5934 ( \6096 , \5930 , \6002 );
or \U$5935 ( \6097 , \6094 , \6095 , \6096 );
xor \U$5936 ( \6098 , \6093 , \6097 );
and \U$5937 ( \6099 , \6033 , \6037 );
and \U$5938 ( \6100 , \6037 , \6042 );
and \U$5939 ( \6101 , \6033 , \6042 );
or \U$5940 ( \6102 , \6099 , \6100 , \6101 );
and \U$5941 ( \6103 , \5934 , \5938 );
and \U$5942 ( \6104 , \5938 , \5943 );
and \U$5943 ( \6105 , \5934 , \5943 );
or \U$5944 ( \6106 , \6103 , \6104 , \6105 );
xor \U$5945 ( \6107 , \6102 , \6106 );
and \U$5946 ( \6108 , \5963 , \5967 );
and \U$5947 ( \6109 , \5967 , \5972 );
and \U$5948 ( \6110 , \5963 , \5972 );
or \U$5949 ( \6111 , \6108 , \6109 , \6110 );
xor \U$5950 ( \6112 , \6107 , \6111 );
and \U$5951 ( \6113 , \5904 , \5908 );
and \U$5952 ( \6114 , \5908 , \5913 );
and \U$5953 ( \6115 , \5904 , \5913 );
or \U$5954 ( \6116 , \6113 , \6114 , \6115 );
and \U$5955 ( \6117 , \5919 , \5923 );
and \U$5956 ( \6118 , \5923 , \5928 );
and \U$5957 ( \6119 , \5919 , \5928 );
or \U$5958 ( \6120 , \6117 , \6118 , \6119 );
xor \U$5959 ( \6121 , \6116 , \6120 );
and \U$5960 ( \6122 , \5948 , \5952 );
and \U$5961 ( \6123 , \5952 , \5957 );
and \U$5962 ( \6124 , \5948 , \5957 );
or \U$5963 ( \6125 , \6122 , \6123 , \6124 );
xor \U$5964 ( \6126 , \6121 , \6125 );
xor \U$5965 ( \6127 , \6112 , \6126 );
and \U$5966 ( \6128 , \5890 , \5894 );
and \U$5967 ( \6129 , \5894 , \5899 );
and \U$5968 ( \6130 , \5890 , \5899 );
or \U$5969 ( \6131 , \6128 , \6129 , \6130 );
and \U$5970 ( \6132 , \5988 , \5992 );
and \U$5971 ( \6133 , \5992 , \6000 );
and \U$5972 ( \6134 , \5988 , \6000 );
or \U$5973 ( \6135 , \6132 , \6133 , \6134 );
xor \U$5974 ( \6136 , \6131 , \6135 );
and \U$5975 ( \6137 , \150 , \5996 );
and \U$5976 ( \6138 , \158 , \5695 );
nor \U$5977 ( \6139 , \6137 , \6138 );
xnor \U$5978 ( \6140 , \6139 , \5687 );
xor \U$5979 ( \6141 , \6136 , \6140 );
buf \U$5980 ( \6142 , RIb5608b8_16);
xor \U$5981 ( \6143 , \6142 , \5683 );
nand \U$5982 ( \6144 , \166 , \6143 );
buf \U$5983 ( \6145 , RIb560930_15);
and \U$5984 ( \6146 , \6142 , \5683 );
not \U$5985 ( \6147 , \6146 );
and \U$5986 ( \6148 , \6145 , \6147 );
xnor \U$5987 ( \6149 , \6144 , \6148 );
and \U$5988 ( \6150 , \178 , \3357 );
and \U$5989 ( \6151 , \185 , \3255 );
nor \U$5990 ( \6152 , \6150 , \6151 );
xnor \U$5991 ( \6153 , \6152 , \3156 );
and \U$5992 ( \6154 , \189 , \3813 );
and \U$5993 ( \6155 , \197 , \3557 );
nor \U$5994 ( \6156 , \6154 , \6155 );
xnor \U$5995 ( \6157 , \6156 , \3562 );
xor \U$5996 ( \6158 , \6153 , \6157 );
and \U$5997 ( \6159 , \209 , \4132 );
and \U$5998 ( \6160 , \217 , \4012 );
nor \U$5999 ( \6161 , \6159 , \6160 );
xnor \U$6000 ( \6162 , \6161 , \3925 );
xor \U$6001 ( \6163 , \6158 , \6162 );
xor \U$6002 ( \6164 , \6149 , \6163 );
and \U$6003 ( \6165 , \224 , \4581 );
and \U$6004 ( \6166 , \232 , \4424 );
nor \U$6005 ( \6167 , \6165 , \6166 );
xnor \U$6006 ( \6168 , \6167 , \4377 );
and \U$6007 ( \6169 , \240 , \5011 );
and \U$6008 ( \6170 , \247 , \4878 );
nor \U$6009 ( \6171 , \6169 , \6170 );
xnor \U$6010 ( \6172 , \6171 , \4762 );
xor \U$6011 ( \6173 , \6168 , \6172 );
and \U$6012 ( \6174 , \134 , \5485 );
and \U$6013 ( \6175 , \143 , \5275 );
nor \U$6014 ( \6176 , \6174 , \6175 );
xnor \U$6015 ( \6177 , \6176 , \5169 );
xor \U$6016 ( \6178 , \6173 , \6177 );
xor \U$6017 ( \6179 , \6164 , \6178 );
xor \U$6018 ( \6180 , \6141 , \6179 );
and \U$6019 ( \6181 , \1802 , \1578 );
and \U$6020 ( \6182 , \1948 , \1431 );
nor \U$6021 ( \6183 , \6181 , \6182 );
xnor \U$6022 ( \6184 , \6183 , \1436 );
and \U$6023 ( \6185 , \1601 , \1824 );
and \U$6024 ( \6186 , \1684 , \1739 );
nor \U$6025 ( \6187 , \6185 , \6186 );
xnor \U$6026 ( \6188 , \6187 , \1697 );
xor \U$6027 ( \6189 , \6184 , \6188 );
and \U$6028 ( \6190 , \1333 , \2121 );
and \U$6029 ( \6191 , \1484 , \2008 );
nor \U$6030 ( \6192 , \6190 , \6191 );
xnor \U$6031 ( \6193 , \6192 , \1961 );
xor \U$6032 ( \6194 , \6189 , \6193 );
and \U$6033 ( \6195 , \2757 , \438 );
and \U$6034 ( \6196 , \2826 , \336 );
nor \U$6035 ( \6197 , \6195 , \6196 );
xnor \U$6036 ( \6198 , \6197 , \320 );
and \U$6037 ( \6199 , \2366 , \1086 );
and \U$6038 ( \6200 , \2521 , \508 );
nor \U$6039 ( \6201 , \6199 , \6200 );
xnor \U$6040 ( \6202 , \6201 , \487 );
xor \U$6041 ( \6203 , \6198 , \6202 );
and \U$6042 ( \6204 , \2090 , \1301 );
and \U$6043 ( \6205 , \2182 , \1246 );
nor \U$6044 ( \6206 , \6204 , \6205 );
xnor \U$6045 ( \6207 , \6206 , \1205 );
xor \U$6046 ( \6208 , \6203 , \6207 );
xor \U$6047 ( \6209 , \6194 , \6208 );
and \U$6048 ( \6210 , \1147 , \2400 );
and \U$6049 ( \6211 , \1192 , \2246 );
nor \U$6050 ( \6212 , \6210 , \6211 );
xnor \U$6051 ( \6213 , \6212 , \2195 );
and \U$6052 ( \6214 , \412 , \2669 );
and \U$6053 ( \6215 , \474 , \2538 );
nor \U$6054 ( \6216 , \6214 , \6215 );
xnor \U$6055 ( \6217 , \6216 , \2534 );
xor \U$6056 ( \6218 , \6213 , \6217 );
and \U$6057 ( \6219 , \261 , \3103 );
and \U$6058 ( \6220 , \307 , \2934 );
nor \U$6059 ( \6221 , \6219 , \6220 );
xnor \U$6060 ( \6222 , \6221 , \2839 );
xor \U$6061 ( \6223 , \6218 , \6222 );
xor \U$6062 ( \6224 , \6209 , \6223 );
xor \U$6063 ( \6225 , \6180 , \6224 );
xor \U$6064 ( \6226 , \6127 , \6225 );
xor \U$6065 ( \6227 , \6098 , \6226 );
and \U$6066 ( \6228 , \5861 , \5865 );
and \U$6067 ( \6229 , \5865 , \5870 );
and \U$6068 ( \6230 , \5861 , \5870 );
or \U$6069 ( \6231 , \6228 , \6229 , \6230 );
and \U$6070 ( \6232 , \5875 , \5879 );
and \U$6071 ( \6233 , \5879 , \5884 );
and \U$6072 ( \6234 , \5875 , \5884 );
or \U$6073 ( \6235 , \6232 , \6233 , \6234 );
xor \U$6074 ( \6236 , \6231 , \6235 );
and \U$6075 ( \6237 , \5979 , \5983 );
and \U$6076 ( \6238 , \5983 , \6001 );
and \U$6077 ( \6239 , \5979 , \6001 );
or \U$6078 ( \6240 , \6237 , \6238 , \6239 );
xor \U$6079 ( \6241 , \6236 , \6240 );
and \U$6080 ( \6242 , \5900 , \5914 );
and \U$6081 ( \6243 , \5914 , \5929 );
and \U$6082 ( \6244 , \5900 , \5929 );
or \U$6083 ( \6245 , \6242 , \6243 , \6244 );
and \U$6084 ( \6246 , \5944 , \5958 );
and \U$6085 ( \6247 , \5958 , \5973 );
and \U$6086 ( \6248 , \5944 , \5973 );
or \U$6087 ( \6249 , \6246 , \6247 , \6248 );
xor \U$6088 ( \6250 , \6245 , \6249 );
and \U$6089 ( \6251 , \3736 , \141 );
and \U$6090 ( \6252 , \3912 , \139 );
nor \U$6091 ( \6253 , \6251 , \6252 );
xnor \U$6092 ( \6254 , \6253 , \148 );
and \U$6093 ( \6255 , \3395 , \156 );
and \U$6094 ( \6256 , \3646 , \154 );
nor \U$6095 ( \6257 , \6255 , \6256 );
xnor \U$6096 ( \6258 , \6257 , \163 );
xor \U$6097 ( \6259 , \6254 , \6258 );
and \U$6098 ( \6260 , \3037 , \296 );
and \U$6099 ( \6261 , \3143 , \168 );
nor \U$6100 ( \6262 , \6260 , \6261 );
xnor \U$6101 ( \6263 , \6262 , \173 );
xor \U$6102 ( \6264 , \6259 , \6263 );
and \U$6103 ( \6265 , \4922 , \215 );
and \U$6104 ( \6266 , \5156 , \213 );
nor \U$6105 ( \6267 , \6265 , \6266 );
xnor \U$6106 ( \6268 , \6267 , \222 );
and \U$6107 ( \6269 , \4654 , \230 );
and \U$6108 ( \6270 , \4749 , \228 );
nor \U$6109 ( \6271 , \6269 , \6270 );
xnor \U$6110 ( \6272 , \6271 , \237 );
xor \U$6111 ( \6273 , \6268 , \6272 );
and \U$6112 ( \6274 , \4160 , \245 );
and \U$6113 ( \6275 , \4364 , \243 );
nor \U$6114 ( \6276 , \6274 , \6275 );
xnor \U$6115 ( \6277 , \6276 , \252 );
xor \U$6116 ( \6278 , \6273 , \6277 );
xor \U$6117 ( \6279 , \6264 , \6278 );
and \U$6118 ( \6280 , \6030 , \183 );
buf \U$6119 ( \6281 , RIb55eab8_80);
and \U$6120 ( \6282 , \6281 , \180 );
nor \U$6121 ( \6283 , \6280 , \6282 );
xnor \U$6122 ( \6284 , \6283 , \179 );
and \U$6123 ( \6285 , \5469 , \195 );
and \U$6124 ( \6286 , \5674 , \193 );
nor \U$6125 ( \6287 , \6285 , \6286 );
xnor \U$6126 ( \6288 , \6287 , \202 );
xor \U$6127 ( \6289 , \6284 , \6288 );
xor \U$6128 ( \6290 , \6289 , \6148 );
xor \U$6129 ( \6291 , \6279 , \6290 );
xor \U$6130 ( \6292 , \6250 , \6291 );
xor \U$6131 ( \6293 , \6241 , \6292 );
xor \U$6132 ( \6294 , \6227 , \6293 );
xor \U$6133 ( \6295 , \6084 , \6294 );
xor \U$6134 ( \6296 , \6075 , \6295 );
and \U$6135 ( \6297 , \5822 , \5823 );
and \U$6136 ( \6298 , \5823 , \6047 );
and \U$6137 ( \6299 , \5822 , \6047 );
or \U$6138 ( \6300 , \6297 , \6298 , \6299 );
xor \U$6139 ( \6301 , \6296 , \6300 );
and \U$6140 ( \6302 , \6048 , \6052 );
and \U$6141 ( \6303 , \6053 , \6056 );
or \U$6142 ( \6304 , \6302 , \6303 );
xor \U$6143 ( \6305 , \6301 , \6304 );
buf g553b_GF_PartitionCandidate( \6306_nG553b , \6305 );
buf \U$6144 ( \6307 , \6306_nG553b );
and \U$6145 ( \6308 , \6079 , \6083 );
and \U$6146 ( \6309 , \6083 , \6294 );
and \U$6147 ( \6310 , \6079 , \6294 );
or \U$6148 ( \6311 , \6308 , \6309 , \6310 );
and \U$6149 ( \6312 , \6088 , \6092 );
and \U$6150 ( \6313 , \6092 , \6097 );
and \U$6151 ( \6314 , \6088 , \6097 );
or \U$6152 ( \6315 , \6312 , \6313 , \6314 );
and \U$6153 ( \6316 , \6112 , \6126 );
and \U$6154 ( \6317 , \6126 , \6225 );
and \U$6155 ( \6318 , \6112 , \6225 );
or \U$6156 ( \6319 , \6316 , \6317 , \6318 );
xor \U$6157 ( \6320 , \6315 , \6319 );
and \U$6158 ( \6321 , \6241 , \6292 );
xor \U$6159 ( \6322 , \6320 , \6321 );
xor \U$6160 ( \6323 , \6311 , \6322 );
and \U$6161 ( \6324 , \6067 , \6071 );
and \U$6162 ( \6325 , \6071 , \6073 );
and \U$6163 ( \6326 , \6067 , \6073 );
or \U$6164 ( \6327 , \6324 , \6325 , \6326 );
and \U$6165 ( \6328 , \6098 , \6226 );
and \U$6166 ( \6329 , \6226 , \6293 );
and \U$6167 ( \6330 , \6098 , \6293 );
or \U$6168 ( \6331 , \6328 , \6329 , \6330 );
xor \U$6169 ( \6332 , \6327 , \6331 );
and \U$6170 ( \6333 , \6131 , \6135 );
and \U$6171 ( \6334 , \6135 , \6140 );
and \U$6172 ( \6335 , \6131 , \6140 );
or \U$6173 ( \6336 , \6333 , \6334 , \6335 );
and \U$6174 ( \6337 , \6102 , \6106 );
and \U$6175 ( \6338 , \6106 , \6111 );
and \U$6176 ( \6339 , \6102 , \6111 );
or \U$6177 ( \6340 , \6337 , \6338 , \6339 );
xor \U$6178 ( \6341 , \6336 , \6340 );
and \U$6179 ( \6342 , \6116 , \6120 );
and \U$6180 ( \6343 , \6120 , \6125 );
and \U$6181 ( \6344 , \6116 , \6125 );
or \U$6182 ( \6345 , \6342 , \6343 , \6344 );
xor \U$6183 ( \6346 , \6341 , \6345 );
and \U$6184 ( \6347 , \6231 , \6235 );
and \U$6185 ( \6348 , \6235 , \6240 );
and \U$6186 ( \6349 , \6231 , \6240 );
or \U$6187 ( \6350 , \6347 , \6348 , \6349 );
and \U$6188 ( \6351 , \6245 , \6249 );
and \U$6189 ( \6352 , \6249 , \6291 );
and \U$6190 ( \6353 , \6245 , \6291 );
or \U$6191 ( \6354 , \6351 , \6352 , \6353 );
xor \U$6192 ( \6355 , \6350 , \6354 );
and \U$6193 ( \6356 , \6141 , \6179 );
and \U$6194 ( \6357 , \6179 , \6224 );
and \U$6195 ( \6358 , \6141 , \6224 );
or \U$6196 ( \6359 , \6356 , \6357 , \6358 );
xor \U$6197 ( \6360 , \6355 , \6359 );
xor \U$6198 ( \6361 , \6346 , \6360 );
and \U$6199 ( \6362 , \6264 , \6278 );
and \U$6200 ( \6363 , \6278 , \6290 );
and \U$6201 ( \6364 , \6264 , \6290 );
or \U$6202 ( \6365 , \6362 , \6363 , \6364 );
and \U$6203 ( \6366 , \6149 , \6163 );
and \U$6204 ( \6367 , \6163 , \6178 );
and \U$6205 ( \6368 , \6149 , \6178 );
or \U$6206 ( \6369 , \6366 , \6367 , \6368 );
xor \U$6207 ( \6370 , \6365 , \6369 );
and \U$6208 ( \6371 , \6194 , \6208 );
and \U$6209 ( \6372 , \6208 , \6223 );
and \U$6210 ( \6373 , \6194 , \6223 );
or \U$6211 ( \6374 , \6371 , \6372 , \6373 );
xor \U$6212 ( \6375 , \6370 , \6374 );
and \U$6213 ( \6376 , \6254 , \6258 );
and \U$6214 ( \6377 , \6258 , \6263 );
and \U$6215 ( \6378 , \6254 , \6263 );
or \U$6216 ( \6379 , \6376 , \6377 , \6378 );
and \U$6217 ( \6380 , \6268 , \6272 );
and \U$6218 ( \6381 , \6272 , \6277 );
and \U$6219 ( \6382 , \6268 , \6277 );
or \U$6220 ( \6383 , \6380 , \6381 , \6382 );
xor \U$6221 ( \6384 , \6379 , \6383 );
and \U$6222 ( \6385 , \6284 , \6288 );
and \U$6223 ( \6386 , \6288 , \6148 );
and \U$6224 ( \6387 , \6284 , \6148 );
or \U$6225 ( \6388 , \6385 , \6386 , \6387 );
xor \U$6226 ( \6389 , \6384 , \6388 );
and \U$6227 ( \6390 , \6153 , \6157 );
and \U$6228 ( \6391 , \6157 , \6162 );
and \U$6229 ( \6392 , \6153 , \6162 );
or \U$6230 ( \6393 , \6390 , \6391 , \6392 );
and \U$6231 ( \6394 , \6168 , \6172 );
and \U$6232 ( \6395 , \6172 , \6177 );
and \U$6233 ( \6396 , \6168 , \6177 );
or \U$6234 ( \6397 , \6394 , \6395 , \6396 );
xor \U$6235 ( \6398 , \6393 , \6397 );
xor \U$6236 ( \6399 , \6145 , \6142 );
not \U$6237 ( \6400 , \6143 );
and \U$6238 ( \6401 , \6399 , \6400 );
and \U$6239 ( \6402 , \166 , \6401 );
and \U$6240 ( \6403 , \150 , \6143 );
nor \U$6241 ( \6404 , \6402 , \6403 );
xnor \U$6242 ( \6405 , \6404 , \6148 );
xor \U$6243 ( \6406 , \6398 , \6405 );
xor \U$6244 ( \6407 , \6389 , \6406 );
and \U$6245 ( \6408 , \6184 , \6188 );
and \U$6246 ( \6409 , \6188 , \6193 );
and \U$6247 ( \6410 , \6184 , \6193 );
or \U$6248 ( \6411 , \6408 , \6409 , \6410 );
and \U$6249 ( \6412 , \6198 , \6202 );
and \U$6250 ( \6413 , \6202 , \6207 );
and \U$6251 ( \6414 , \6198 , \6207 );
or \U$6252 ( \6415 , \6412 , \6413 , \6414 );
xor \U$6253 ( \6416 , \6411 , \6415 );
and \U$6254 ( \6417 , \6213 , \6217 );
and \U$6255 ( \6418 , \6217 , \6222 );
and \U$6256 ( \6419 , \6213 , \6222 );
or \U$6257 ( \6420 , \6417 , \6418 , \6419 );
xor \U$6258 ( \6421 , \6416 , \6420 );
xor \U$6259 ( \6422 , \6407 , \6421 );
xor \U$6260 ( \6423 , \6375 , \6422 );
and \U$6261 ( \6424 , \247 , \5011 );
and \U$6262 ( \6425 , \224 , \4878 );
nor \U$6263 ( \6426 , \6424 , \6425 );
xnor \U$6264 ( \6427 , \6426 , \4762 );
and \U$6265 ( \6428 , \143 , \5485 );
and \U$6266 ( \6429 , \240 , \5275 );
nor \U$6267 ( \6430 , \6428 , \6429 );
xnor \U$6268 ( \6431 , \6430 , \5169 );
xor \U$6269 ( \6432 , \6427 , \6431 );
and \U$6270 ( \6433 , \158 , \5996 );
and \U$6271 ( \6434 , \134 , \5695 );
nor \U$6272 ( \6435 , \6433 , \6434 );
xnor \U$6273 ( \6436 , \6435 , \5687 );
xor \U$6274 ( \6437 , \6432 , \6436 );
and \U$6275 ( \6438 , \474 , \2669 );
and \U$6276 ( \6439 , \1147 , \2538 );
nor \U$6277 ( \6440 , \6438 , \6439 );
xnor \U$6278 ( \6441 , \6440 , \2534 );
and \U$6279 ( \6442 , \307 , \3103 );
and \U$6280 ( \6443 , \412 , \2934 );
nor \U$6281 ( \6444 , \6442 , \6443 );
xnor \U$6282 ( \6445 , \6444 , \2839 );
xor \U$6283 ( \6446 , \6441 , \6445 );
and \U$6284 ( \6447 , \185 , \3357 );
and \U$6285 ( \6448 , \261 , \3255 );
nor \U$6286 ( \6449 , \6447 , \6448 );
xnor \U$6287 ( \6450 , \6449 , \3156 );
xor \U$6288 ( \6451 , \6446 , \6450 );
xor \U$6289 ( \6452 , \6437 , \6451 );
and \U$6290 ( \6453 , \197 , \3813 );
and \U$6291 ( \6454 , \178 , \3557 );
nor \U$6292 ( \6455 , \6453 , \6454 );
xnor \U$6293 ( \6456 , \6455 , \3562 );
and \U$6294 ( \6457 , \217 , \4132 );
and \U$6295 ( \6458 , \189 , \4012 );
nor \U$6296 ( \6459 , \6457 , \6458 );
xnor \U$6297 ( \6460 , \6459 , \3925 );
xor \U$6298 ( \6461 , \6456 , \6460 );
and \U$6299 ( \6462 , \232 , \4581 );
and \U$6300 ( \6463 , \209 , \4424 );
nor \U$6301 ( \6464 , \6462 , \6463 );
xnor \U$6302 ( \6465 , \6464 , \4377 );
xor \U$6303 ( \6466 , \6461 , \6465 );
xor \U$6304 ( \6467 , \6452 , \6466 );
and \U$6305 ( \6468 , \1684 , \1824 );
and \U$6306 ( \6469 , \1802 , \1739 );
nor \U$6307 ( \6470 , \6468 , \6469 );
xnor \U$6308 ( \6471 , \6470 , \1697 );
and \U$6309 ( \6472 , \1484 , \2121 );
and \U$6310 ( \6473 , \1601 , \2008 );
nor \U$6311 ( \6474 , \6472 , \6473 );
xnor \U$6312 ( \6475 , \6474 , \1961 );
xor \U$6313 ( \6476 , \6471 , \6475 );
and \U$6314 ( \6477 , \1192 , \2400 );
and \U$6315 ( \6478 , \1333 , \2246 );
nor \U$6316 ( \6479 , \6477 , \6478 );
xnor \U$6317 ( \6480 , \6479 , \2195 );
xor \U$6318 ( \6481 , \6476 , \6480 );
and \U$6319 ( \6482 , \2521 , \1086 );
and \U$6320 ( \6483 , \2757 , \508 );
nor \U$6321 ( \6484 , \6482 , \6483 );
xnor \U$6322 ( \6485 , \6484 , \487 );
and \U$6323 ( \6486 , \2182 , \1301 );
and \U$6324 ( \6487 , \2366 , \1246 );
nor \U$6325 ( \6488 , \6486 , \6487 );
xnor \U$6326 ( \6489 , \6488 , \1205 );
xor \U$6327 ( \6490 , \6485 , \6489 );
and \U$6328 ( \6491 , \1948 , \1578 );
and \U$6329 ( \6492 , \2090 , \1431 );
nor \U$6330 ( \6493 , \6491 , \6492 );
xnor \U$6331 ( \6494 , \6493 , \1436 );
xor \U$6332 ( \6495 , \6490 , \6494 );
xor \U$6333 ( \6496 , \6481 , \6495 );
and \U$6334 ( \6497 , \3646 , \156 );
and \U$6335 ( \6498 , \3736 , \154 );
nor \U$6336 ( \6499 , \6497 , \6498 );
xnor \U$6337 ( \6500 , \6499 , \163 );
and \U$6338 ( \6501 , \3143 , \296 );
and \U$6339 ( \6502 , \3395 , \168 );
nor \U$6340 ( \6503 , \6501 , \6502 );
xnor \U$6341 ( \6504 , \6503 , \173 );
xor \U$6342 ( \6505 , \6500 , \6504 );
and \U$6343 ( \6506 , \2826 , \438 );
and \U$6344 ( \6507 , \3037 , \336 );
nor \U$6345 ( \6508 , \6506 , \6507 );
xnor \U$6346 ( \6509 , \6508 , \320 );
xor \U$6347 ( \6510 , \6505 , \6509 );
xor \U$6348 ( \6511 , \6496 , \6510 );
xor \U$6349 ( \6512 , \6467 , \6511 );
and \U$6350 ( \6513 , \6281 , \183 );
buf \U$6351 ( \6514 , RIb55eb30_79);
and \U$6352 ( \6515 , \6514 , \180 );
nor \U$6353 ( \6516 , \6513 , \6515 );
xnor \U$6354 ( \6517 , \6516 , \179 );
and \U$6355 ( \6518 , \5674 , \195 );
and \U$6356 ( \6519 , \6030 , \193 );
nor \U$6357 ( \6520 , \6518 , \6519 );
xnor \U$6358 ( \6521 , \6520 , \202 );
xor \U$6359 ( \6522 , \6517 , \6521 );
and \U$6360 ( \6523 , \5156 , \215 );
and \U$6361 ( \6524 , \5469 , \213 );
nor \U$6362 ( \6525 , \6523 , \6524 );
xnor \U$6363 ( \6526 , \6525 , \222 );
xor \U$6364 ( \6527 , \6522 , \6526 );
and \U$6365 ( \6528 , \4749 , \230 );
and \U$6366 ( \6529 , \4922 , \228 );
nor \U$6367 ( \6530 , \6528 , \6529 );
xnor \U$6368 ( \6531 , \6530 , \237 );
and \U$6369 ( \6532 , \4364 , \245 );
and \U$6370 ( \6533 , \4654 , \243 );
nor \U$6371 ( \6534 , \6532 , \6533 );
xnor \U$6372 ( \6535 , \6534 , \252 );
xor \U$6373 ( \6536 , \6531 , \6535 );
and \U$6374 ( \6537 , \3912 , \141 );
and \U$6375 ( \6538 , \4160 , \139 );
nor \U$6376 ( \6539 , \6537 , \6538 );
xnor \U$6377 ( \6540 , \6539 , \148 );
xor \U$6378 ( \6541 , \6536 , \6540 );
xor \U$6379 ( \6542 , \6527 , \6541 );
xor \U$6380 ( \6543 , \6512 , \6542 );
xor \U$6381 ( \6544 , \6423 , \6543 );
xor \U$6382 ( \6545 , \6361 , \6544 );
xor \U$6383 ( \6546 , \6332 , \6545 );
xor \U$6384 ( \6547 , \6323 , \6546 );
and \U$6385 ( \6548 , \6063 , \6074 );
and \U$6386 ( \6549 , \6074 , \6295 );
and \U$6387 ( \6550 , \6063 , \6295 );
or \U$6388 ( \6551 , \6548 , \6549 , \6550 );
xor \U$6389 ( \6552 , \6547 , \6551 );
and \U$6390 ( \6553 , \6296 , \6300 );
and \U$6391 ( \6554 , \6301 , \6304 );
or \U$6392 ( \6555 , \6553 , \6554 );
xor \U$6393 ( \6556 , \6552 , \6555 );
buf g5539_GF_PartitionCandidate( \6557_nG5539 , \6556 );
buf \U$6394 ( \6558 , \6557_nG5539 );
and \U$6395 ( \6559 , \6327 , \6331 );
and \U$6396 ( \6560 , \6331 , \6545 );
and \U$6397 ( \6561 , \6327 , \6545 );
or \U$6398 ( \6562 , \6559 , \6560 , \6561 );
and \U$6399 ( \6563 , \6350 , \6354 );
and \U$6400 ( \6564 , \6354 , \6359 );
and \U$6401 ( \6565 , \6350 , \6359 );
or \U$6402 ( \6566 , \6563 , \6564 , \6565 );
and \U$6403 ( \6567 , \6375 , \6422 );
and \U$6404 ( \6568 , \6422 , \6543 );
and \U$6405 ( \6569 , \6375 , \6543 );
or \U$6406 ( \6570 , \6567 , \6568 , \6569 );
xor \U$6407 ( \6571 , \6566 , \6570 );
and \U$6408 ( \6572 , \6437 , \6451 );
and \U$6409 ( \6573 , \6451 , \6466 );
and \U$6410 ( \6574 , \6437 , \6466 );
or \U$6411 ( \6575 , \6572 , \6573 , \6574 );
and \U$6412 ( \6576 , \6481 , \6495 );
and \U$6413 ( \6577 , \6495 , \6510 );
and \U$6414 ( \6578 , \6481 , \6510 );
or \U$6415 ( \6579 , \6576 , \6577 , \6578 );
xor \U$6416 ( \6580 , \6575 , \6579 );
and \U$6417 ( \6581 , \6527 , \6541 );
xor \U$6418 ( \6582 , \6580 , \6581 );
xor \U$6419 ( \6583 , \6571 , \6582 );
xor \U$6420 ( \6584 , \6562 , \6583 );
and \U$6421 ( \6585 , \6315 , \6319 );
and \U$6422 ( \6586 , \6319 , \6321 );
and \U$6423 ( \6587 , \6315 , \6321 );
or \U$6424 ( \6588 , \6585 , \6586 , \6587 );
and \U$6425 ( \6589 , \6346 , \6360 );
and \U$6426 ( \6590 , \6360 , \6544 );
and \U$6427 ( \6591 , \6346 , \6544 );
or \U$6428 ( \6592 , \6589 , \6590 , \6591 );
xor \U$6429 ( \6593 , \6588 , \6592 );
and \U$6430 ( \6594 , \6379 , \6383 );
and \U$6431 ( \6595 , \6383 , \6388 );
and \U$6432 ( \6596 , \6379 , \6388 );
or \U$6433 ( \6597 , \6594 , \6595 , \6596 );
and \U$6434 ( \6598 , \6393 , \6397 );
and \U$6435 ( \6599 , \6397 , \6405 );
and \U$6436 ( \6600 , \6393 , \6405 );
or \U$6437 ( \6601 , \6598 , \6599 , \6600 );
xor \U$6438 ( \6602 , \6597 , \6601 );
and \U$6439 ( \6603 , \6411 , \6415 );
and \U$6440 ( \6604 , \6415 , \6420 );
and \U$6441 ( \6605 , \6411 , \6420 );
or \U$6442 ( \6606 , \6603 , \6604 , \6605 );
xor \U$6443 ( \6607 , \6602 , \6606 );
and \U$6444 ( \6608 , \6365 , \6369 );
and \U$6445 ( \6609 , \6369 , \6374 );
and \U$6446 ( \6610 , \6365 , \6374 );
or \U$6447 ( \6611 , \6608 , \6609 , \6610 );
and \U$6448 ( \6612 , \6336 , \6340 );
and \U$6449 ( \6613 , \6340 , \6345 );
and \U$6450 ( \6614 , \6336 , \6345 );
or \U$6451 ( \6615 , \6612 , \6613 , \6614 );
xor \U$6452 ( \6616 , \6611 , \6615 );
and \U$6453 ( \6617 , \6467 , \6511 );
and \U$6454 ( \6618 , \6511 , \6542 );
and \U$6455 ( \6619 , \6467 , \6542 );
or \U$6456 ( \6620 , \6617 , \6618 , \6619 );
xor \U$6457 ( \6621 , \6616 , \6620 );
xor \U$6458 ( \6622 , \6607 , \6621 );
and \U$6459 ( \6623 , \6389 , \6406 );
and \U$6460 ( \6624 , \6406 , \6421 );
and \U$6461 ( \6625 , \6389 , \6421 );
or \U$6462 ( \6626 , \6623 , \6624 , \6625 );
and \U$6463 ( \6627 , \6500 , \6504 );
and \U$6464 ( \6628 , \6504 , \6509 );
and \U$6465 ( \6629 , \6500 , \6509 );
or \U$6466 ( \6630 , \6627 , \6628 , \6629 );
and \U$6467 ( \6631 , \6517 , \6521 );
and \U$6468 ( \6632 , \6521 , \6526 );
and \U$6469 ( \6633 , \6517 , \6526 );
or \U$6470 ( \6634 , \6631 , \6632 , \6633 );
xor \U$6471 ( \6635 , \6630 , \6634 );
and \U$6472 ( \6636 , \6531 , \6535 );
and \U$6473 ( \6637 , \6535 , \6540 );
and \U$6474 ( \6638 , \6531 , \6540 );
or \U$6475 ( \6639 , \6636 , \6637 , \6638 );
xor \U$6476 ( \6640 , \6635 , \6639 );
and \U$6477 ( \6641 , \6471 , \6475 );
and \U$6478 ( \6642 , \6475 , \6480 );
and \U$6479 ( \6643 , \6471 , \6480 );
or \U$6480 ( \6644 , \6641 , \6642 , \6643 );
and \U$6481 ( \6645 , \6485 , \6489 );
and \U$6482 ( \6646 , \6489 , \6494 );
and \U$6483 ( \6647 , \6485 , \6494 );
or \U$6484 ( \6648 , \6645 , \6646 , \6647 );
xor \U$6485 ( \6649 , \6644 , \6648 );
and \U$6486 ( \6650 , \6441 , \6445 );
and \U$6487 ( \6651 , \6445 , \6450 );
and \U$6488 ( \6652 , \6441 , \6450 );
or \U$6489 ( \6653 , \6650 , \6651 , \6652 );
xor \U$6490 ( \6654 , \6649 , \6653 );
xor \U$6491 ( \6655 , \6640 , \6654 );
and \U$6492 ( \6656 , \6427 , \6431 );
and \U$6493 ( \6657 , \6431 , \6436 );
and \U$6494 ( \6658 , \6427 , \6436 );
or \U$6495 ( \6659 , \6656 , \6657 , \6658 );
and \U$6496 ( \6660 , \6456 , \6460 );
and \U$6497 ( \6661 , \6460 , \6465 );
and \U$6498 ( \6662 , \6456 , \6465 );
or \U$6499 ( \6663 , \6660 , \6661 , \6662 );
xor \U$6500 ( \6664 , \6659 , \6663 );
and \U$6501 ( \6665 , \134 , \5996 );
and \U$6502 ( \6666 , \143 , \5695 );
nor \U$6503 ( \6667 , \6665 , \6666 );
xnor \U$6504 ( \6668 , \6667 , \5687 );
and \U$6505 ( \6669 , \150 , \6401 );
and \U$6506 ( \6670 , \158 , \6143 );
nor \U$6507 ( \6671 , \6669 , \6670 );
xnor \U$6508 ( \6672 , \6671 , \6148 );
xor \U$6509 ( \6673 , \6668 , \6672 );
buf \U$6510 ( \6674 , RIb5609a8_14);
xor \U$6511 ( \6675 , \6674 , \6145 );
nand \U$6512 ( \6676 , \166 , \6675 );
buf \U$6513 ( \6677 , RIb560a20_13);
and \U$6514 ( \6678 , \6674 , \6145 );
not \U$6515 ( \6679 , \6678 );
and \U$6516 ( \6680 , \6677 , \6679 );
xnor \U$6517 ( \6681 , \6676 , \6680 );
xor \U$6518 ( \6682 , \6673 , \6681 );
xor \U$6519 ( \6683 , \6664 , \6682 );
xor \U$6520 ( \6684 , \6655 , \6683 );
xor \U$6521 ( \6685 , \6626 , \6684 );
and \U$6522 ( \6686 , \261 , \3357 );
and \U$6523 ( \6687 , \307 , \3255 );
nor \U$6524 ( \6688 , \6686 , \6687 );
xnor \U$6525 ( \6689 , \6688 , \3156 );
and \U$6526 ( \6690 , \178 , \3813 );
and \U$6527 ( \6691 , \185 , \3557 );
nor \U$6528 ( \6692 , \6690 , \6691 );
xnor \U$6529 ( \6693 , \6692 , \3562 );
xor \U$6530 ( \6694 , \6689 , \6693 );
and \U$6531 ( \6695 , \189 , \4132 );
and \U$6532 ( \6696 , \197 , \4012 );
nor \U$6533 ( \6697 , \6695 , \6696 );
xnor \U$6534 ( \6698 , \6697 , \3925 );
xor \U$6535 ( \6699 , \6694 , \6698 );
and \U$6536 ( \6700 , \1333 , \2400 );
and \U$6537 ( \6701 , \1484 , \2246 );
nor \U$6538 ( \6702 , \6700 , \6701 );
xnor \U$6539 ( \6703 , \6702 , \2195 );
and \U$6540 ( \6704 , \1147 , \2669 );
and \U$6541 ( \6705 , \1192 , \2538 );
nor \U$6542 ( \6706 , \6704 , \6705 );
xnor \U$6543 ( \6707 , \6706 , \2534 );
xor \U$6544 ( \6708 , \6703 , \6707 );
and \U$6545 ( \6709 , \412 , \3103 );
and \U$6546 ( \6710 , \474 , \2934 );
nor \U$6547 ( \6711 , \6709 , \6710 );
xnor \U$6548 ( \6712 , \6711 , \2839 );
xor \U$6549 ( \6713 , \6708 , \6712 );
xor \U$6550 ( \6714 , \6699 , \6713 );
and \U$6551 ( \6715 , \209 , \4581 );
and \U$6552 ( \6716 , \217 , \4424 );
nor \U$6553 ( \6717 , \6715 , \6716 );
xnor \U$6554 ( \6718 , \6717 , \4377 );
and \U$6555 ( \6719 , \224 , \5011 );
and \U$6556 ( \6720 , \232 , \4878 );
nor \U$6557 ( \6721 , \6719 , \6720 );
xnor \U$6558 ( \6722 , \6721 , \4762 );
xor \U$6559 ( \6723 , \6718 , \6722 );
and \U$6560 ( \6724 , \240 , \5485 );
and \U$6561 ( \6725 , \247 , \5275 );
nor \U$6562 ( \6726 , \6724 , \6725 );
xnor \U$6563 ( \6727 , \6726 , \5169 );
xor \U$6564 ( \6728 , \6723 , \6727 );
xor \U$6565 ( \6729 , \6714 , \6728 );
and \U$6566 ( \6730 , \2090 , \1578 );
and \U$6567 ( \6731 , \2182 , \1431 );
nor \U$6568 ( \6732 , \6730 , \6731 );
xnor \U$6569 ( \6733 , \6732 , \1436 );
and \U$6570 ( \6734 , \1802 , \1824 );
and \U$6571 ( \6735 , \1948 , \1739 );
nor \U$6572 ( \6736 , \6734 , \6735 );
xnor \U$6573 ( \6737 , \6736 , \1697 );
xor \U$6574 ( \6738 , \6733 , \6737 );
and \U$6575 ( \6739 , \1601 , \2121 );
and \U$6576 ( \6740 , \1684 , \2008 );
nor \U$6577 ( \6741 , \6739 , \6740 );
xnor \U$6578 ( \6742 , \6741 , \1961 );
xor \U$6579 ( \6743 , \6738 , \6742 );
and \U$6580 ( \6744 , \3037 , \438 );
and \U$6581 ( \6745 , \3143 , \336 );
nor \U$6582 ( \6746 , \6744 , \6745 );
xnor \U$6583 ( \6747 , \6746 , \320 );
and \U$6584 ( \6748 , \2757 , \1086 );
and \U$6585 ( \6749 , \2826 , \508 );
nor \U$6586 ( \6750 , \6748 , \6749 );
xnor \U$6587 ( \6751 , \6750 , \487 );
xor \U$6588 ( \6752 , \6747 , \6751 );
and \U$6589 ( \6753 , \2366 , \1301 );
and \U$6590 ( \6754 , \2521 , \1246 );
nor \U$6591 ( \6755 , \6753 , \6754 );
xnor \U$6592 ( \6756 , \6755 , \1205 );
xor \U$6593 ( \6757 , \6752 , \6756 );
xor \U$6594 ( \6758 , \6743 , \6757 );
and \U$6595 ( \6759 , \4160 , \141 );
and \U$6596 ( \6760 , \4364 , \139 );
nor \U$6597 ( \6761 , \6759 , \6760 );
xnor \U$6598 ( \6762 , \6761 , \148 );
and \U$6599 ( \6763 , \3736 , \156 );
and \U$6600 ( \6764 , \3912 , \154 );
nor \U$6601 ( \6765 , \6763 , \6764 );
xnor \U$6602 ( \6766 , \6765 , \163 );
xor \U$6603 ( \6767 , \6762 , \6766 );
and \U$6604 ( \6768 , \3395 , \296 );
and \U$6605 ( \6769 , \3646 , \168 );
nor \U$6606 ( \6770 , \6768 , \6769 );
xnor \U$6607 ( \6771 , \6770 , \173 );
xor \U$6608 ( \6772 , \6767 , \6771 );
xor \U$6609 ( \6773 , \6758 , \6772 );
xor \U$6610 ( \6774 , \6729 , \6773 );
and \U$6611 ( \6775 , \5469 , \215 );
and \U$6612 ( \6776 , \5674 , \213 );
nor \U$6613 ( \6777 , \6775 , \6776 );
xnor \U$6614 ( \6778 , \6777 , \222 );
and \U$6615 ( \6779 , \4922 , \230 );
and \U$6616 ( \6780 , \5156 , \228 );
nor \U$6617 ( \6781 , \6779 , \6780 );
xnor \U$6618 ( \6782 , \6781 , \237 );
xor \U$6619 ( \6783 , \6778 , \6782 );
and \U$6620 ( \6784 , \4654 , \245 );
and \U$6621 ( \6785 , \4749 , \243 );
nor \U$6622 ( \6786 , \6784 , \6785 );
xnor \U$6623 ( \6787 , \6786 , \252 );
xor \U$6624 ( \6788 , \6783 , \6787 );
and \U$6625 ( \6789 , \6514 , \183 );
buf \U$6626 ( \6790 , RIb55eba8_78);
and \U$6627 ( \6791 , \6790 , \180 );
nor \U$6628 ( \6792 , \6789 , \6791 );
xnor \U$6629 ( \6793 , \6792 , \179 );
and \U$6630 ( \6794 , \6030 , \195 );
and \U$6631 ( \6795 , \6281 , \193 );
nor \U$6632 ( \6796 , \6794 , \6795 );
xnor \U$6633 ( \6797 , \6796 , \202 );
xor \U$6634 ( \6798 , \6793 , \6797 );
xor \U$6635 ( \6799 , \6798 , \6680 );
xor \U$6636 ( \6800 , \6788 , \6799 );
xor \U$6637 ( \6801 , \6774 , \6800 );
xor \U$6638 ( \6802 , \6685 , \6801 );
xor \U$6639 ( \6803 , \6622 , \6802 );
xor \U$6640 ( \6804 , \6593 , \6803 );
xor \U$6641 ( \6805 , \6584 , \6804 );
and \U$6642 ( \6806 , \6311 , \6322 );
and \U$6643 ( \6807 , \6322 , \6546 );
and \U$6644 ( \6808 , \6311 , \6546 );
or \U$6645 ( \6809 , \6806 , \6807 , \6808 );
xor \U$6646 ( \6810 , \6805 , \6809 );
and \U$6647 ( \6811 , \6547 , \6551 );
and \U$6648 ( \6812 , \6552 , \6555 );
or \U$6649 ( \6813 , \6811 , \6812 );
xor \U$6650 ( \6814 , \6810 , \6813 );
buf g5537_GF_PartitionCandidate( \6815_nG5537 , \6814 );
buf \U$6651 ( \6816 , \6815_nG5537 );
and \U$6652 ( \6817 , \6588 , \6592 );
and \U$6653 ( \6818 , \6592 , \6803 );
and \U$6654 ( \6819 , \6588 , \6803 );
or \U$6655 ( \6820 , \6817 , \6818 , \6819 );
and \U$6656 ( \6821 , \6611 , \6615 );
and \U$6657 ( \6822 , \6615 , \6620 );
and \U$6658 ( \6823 , \6611 , \6620 );
or \U$6659 ( \6824 , \6821 , \6822 , \6823 );
and \U$6660 ( \6825 , \6626 , \6684 );
and \U$6661 ( \6826 , \6684 , \6801 );
and \U$6662 ( \6827 , \6626 , \6801 );
or \U$6663 ( \6828 , \6825 , \6826 , \6827 );
xor \U$6664 ( \6829 , \6824 , \6828 );
and \U$6665 ( \6830 , \6699 , \6713 );
and \U$6666 ( \6831 , \6713 , \6728 );
and \U$6667 ( \6832 , \6699 , \6728 );
or \U$6668 ( \6833 , \6830 , \6831 , \6832 );
and \U$6669 ( \6834 , \6743 , \6757 );
and \U$6670 ( \6835 , \6757 , \6772 );
and \U$6671 ( \6836 , \6743 , \6772 );
or \U$6672 ( \6837 , \6834 , \6835 , \6836 );
xor \U$6673 ( \6838 , \6833 , \6837 );
and \U$6674 ( \6839 , \6788 , \6799 );
xor \U$6675 ( \6840 , \6838 , \6839 );
xor \U$6676 ( \6841 , \6829 , \6840 );
xor \U$6677 ( \6842 , \6820 , \6841 );
and \U$6678 ( \6843 , \6566 , \6570 );
and \U$6679 ( \6844 , \6570 , \6582 );
and \U$6680 ( \6845 , \6566 , \6582 );
or \U$6681 ( \6846 , \6843 , \6844 , \6845 );
and \U$6682 ( \6847 , \6607 , \6621 );
and \U$6683 ( \6848 , \6621 , \6802 );
and \U$6684 ( \6849 , \6607 , \6802 );
or \U$6685 ( \6850 , \6847 , \6848 , \6849 );
xor \U$6686 ( \6851 , \6846 , \6850 );
and \U$6687 ( \6852 , \6630 , \6634 );
and \U$6688 ( \6853 , \6634 , \6639 );
and \U$6689 ( \6854 , \6630 , \6639 );
or \U$6690 ( \6855 , \6852 , \6853 , \6854 );
and \U$6691 ( \6856 , \6644 , \6648 );
and \U$6692 ( \6857 , \6648 , \6653 );
and \U$6693 ( \6858 , \6644 , \6653 );
or \U$6694 ( \6859 , \6856 , \6857 , \6858 );
xor \U$6695 ( \6860 , \6855 , \6859 );
and \U$6696 ( \6861 , \6659 , \6663 );
and \U$6697 ( \6862 , \6663 , \6682 );
and \U$6698 ( \6863 , \6659 , \6682 );
or \U$6699 ( \6864 , \6861 , \6862 , \6863 );
xor \U$6700 ( \6865 , \6860 , \6864 );
and \U$6701 ( \6866 , \6597 , \6601 );
and \U$6702 ( \6867 , \6601 , \6606 );
and \U$6703 ( \6868 , \6597 , \6606 );
or \U$6704 ( \6869 , \6866 , \6867 , \6868 );
and \U$6705 ( \6870 , \6575 , \6579 );
and \U$6706 ( \6871 , \6579 , \6581 );
and \U$6707 ( \6872 , \6575 , \6581 );
or \U$6708 ( \6873 , \6870 , \6871 , \6872 );
xor \U$6709 ( \6874 , \6869 , \6873 );
and \U$6710 ( \6875 , \6729 , \6773 );
and \U$6711 ( \6876 , \6773 , \6800 );
and \U$6712 ( \6877 , \6729 , \6800 );
or \U$6713 ( \6878 , \6875 , \6876 , \6877 );
xor \U$6714 ( \6879 , \6874 , \6878 );
xor \U$6715 ( \6880 , \6865 , \6879 );
and \U$6716 ( \6881 , \6640 , \6654 );
and \U$6717 ( \6882 , \6654 , \6683 );
and \U$6718 ( \6883 , \6640 , \6683 );
or \U$6719 ( \6884 , \6881 , \6882 , \6883 );
and \U$6720 ( \6885 , \6733 , \6737 );
and \U$6721 ( \6886 , \6737 , \6742 );
and \U$6722 ( \6887 , \6733 , \6742 );
or \U$6723 ( \6888 , \6885 , \6886 , \6887 );
and \U$6724 ( \6889 , \6747 , \6751 );
and \U$6725 ( \6890 , \6751 , \6756 );
and \U$6726 ( \6891 , \6747 , \6756 );
or \U$6727 ( \6892 , \6889 , \6890 , \6891 );
xor \U$6728 ( \6893 , \6888 , \6892 );
and \U$6729 ( \6894 , \6703 , \6707 );
and \U$6730 ( \6895 , \6707 , \6712 );
and \U$6731 ( \6896 , \6703 , \6712 );
or \U$6732 ( \6897 , \6894 , \6895 , \6896 );
xor \U$6733 ( \6898 , \6893 , \6897 );
and \U$6734 ( \6899 , \6762 , \6766 );
and \U$6735 ( \6900 , \6766 , \6771 );
and \U$6736 ( \6901 , \6762 , \6771 );
or \U$6737 ( \6902 , \6899 , \6900 , \6901 );
and \U$6738 ( \6903 , \6778 , \6782 );
and \U$6739 ( \6904 , \6782 , \6787 );
and \U$6740 ( \6905 , \6778 , \6787 );
or \U$6741 ( \6906 , \6903 , \6904 , \6905 );
xor \U$6742 ( \6907 , \6902 , \6906 );
and \U$6743 ( \6908 , \6793 , \6797 );
and \U$6744 ( \6909 , \6797 , \6680 );
and \U$6745 ( \6910 , \6793 , \6680 );
or \U$6746 ( \6911 , \6908 , \6909 , \6910 );
xor \U$6747 ( \6912 , \6907 , \6911 );
xor \U$6748 ( \6913 , \6898 , \6912 );
and \U$6749 ( \6914 , \6689 , \6693 );
and \U$6750 ( \6915 , \6693 , \6698 );
and \U$6751 ( \6916 , \6689 , \6698 );
or \U$6752 ( \6917 , \6914 , \6915 , \6916 );
and \U$6753 ( \6918 , \6668 , \6672 );
and \U$6754 ( \6919 , \6672 , \6681 );
and \U$6755 ( \6920 , \6668 , \6681 );
or \U$6756 ( \6921 , \6918 , \6919 , \6920 );
xor \U$6757 ( \6922 , \6917 , \6921 );
and \U$6758 ( \6923 , \6718 , \6722 );
and \U$6759 ( \6924 , \6722 , \6727 );
and \U$6760 ( \6925 , \6718 , \6727 );
or \U$6761 ( \6926 , \6923 , \6924 , \6925 );
xor \U$6762 ( \6927 , \6922 , \6926 );
xor \U$6763 ( \6928 , \6913 , \6927 );
xor \U$6764 ( \6929 , \6884 , \6928 );
and \U$6765 ( \6930 , \3912 , \156 );
and \U$6766 ( \6931 , \4160 , \154 );
nor \U$6767 ( \6932 , \6930 , \6931 );
xnor \U$6768 ( \6933 , \6932 , \163 );
and \U$6769 ( \6934 , \3646 , \296 );
and \U$6770 ( \6935 , \3736 , \168 );
nor \U$6771 ( \6936 , \6934 , \6935 );
xnor \U$6772 ( \6937 , \6936 , \173 );
xor \U$6773 ( \6938 , \6933 , \6937 );
and \U$6774 ( \6939 , \3143 , \438 );
and \U$6775 ( \6940 , \3395 , \336 );
nor \U$6776 ( \6941 , \6939 , \6940 );
xnor \U$6777 ( \6942 , \6941 , \320 );
xor \U$6778 ( \6943 , \6938 , \6942 );
and \U$6779 ( \6944 , \6790 , \183 );
buf \U$6780 ( \6945 , RIb55ec20_77);
and \U$6781 ( \6946 , \6945 , \180 );
nor \U$6782 ( \6947 , \6944 , \6946 );
xnor \U$6783 ( \6948 , \6947 , \179 );
and \U$6784 ( \6949 , \6281 , \195 );
and \U$6785 ( \6950 , \6514 , \193 );
nor \U$6786 ( \6951 , \6949 , \6950 );
xnor \U$6787 ( \6952 , \6951 , \202 );
xor \U$6788 ( \6953 , \6948 , \6952 );
and \U$6789 ( \6954 , \5674 , \215 );
and \U$6790 ( \6955 , \6030 , \213 );
nor \U$6791 ( \6956 , \6954 , \6955 );
xnor \U$6792 ( \6957 , \6956 , \222 );
xor \U$6793 ( \6958 , \6953 , \6957 );
xor \U$6794 ( \6959 , \6943 , \6958 );
and \U$6795 ( \6960 , \5156 , \230 );
and \U$6796 ( \6961 , \5469 , \228 );
nor \U$6797 ( \6962 , \6960 , \6961 );
xnor \U$6798 ( \6963 , \6962 , \237 );
and \U$6799 ( \6964 , \4749 , \245 );
and \U$6800 ( \6965 , \4922 , \243 );
nor \U$6801 ( \6966 , \6964 , \6965 );
xnor \U$6802 ( \6967 , \6966 , \252 );
xor \U$6803 ( \6968 , \6963 , \6967 );
and \U$6804 ( \6969 , \4364 , \141 );
and \U$6805 ( \6970 , \4654 , \139 );
nor \U$6806 ( \6971 , \6969 , \6970 );
xnor \U$6807 ( \6972 , \6971 , \148 );
xor \U$6808 ( \6973 , \6968 , \6972 );
xor \U$6809 ( \6974 , \6959 , \6973 );
and \U$6810 ( \6975 , \1948 , \1824 );
and \U$6811 ( \6976 , \2090 , \1739 );
nor \U$6812 ( \6977 , \6975 , \6976 );
xnor \U$6813 ( \6978 , \6977 , \1697 );
and \U$6814 ( \6979 , \1684 , \2121 );
and \U$6815 ( \6980 , \1802 , \2008 );
nor \U$6816 ( \6981 , \6979 , \6980 );
xnor \U$6817 ( \6982 , \6981 , \1961 );
xor \U$6818 ( \6983 , \6978 , \6982 );
and \U$6819 ( \6984 , \1484 , \2400 );
and \U$6820 ( \6985 , \1601 , \2246 );
nor \U$6821 ( \6986 , \6984 , \6985 );
xnor \U$6822 ( \6987 , \6986 , \2195 );
xor \U$6823 ( \6988 , \6983 , \6987 );
and \U$6824 ( \6989 , \2826 , \1086 );
and \U$6825 ( \6990 , \3037 , \508 );
nor \U$6826 ( \6991 , \6989 , \6990 );
xnor \U$6827 ( \6992 , \6991 , \487 );
and \U$6828 ( \6993 , \2521 , \1301 );
and \U$6829 ( \6994 , \2757 , \1246 );
nor \U$6830 ( \6995 , \6993 , \6994 );
xnor \U$6831 ( \6996 , \6995 , \1205 );
xor \U$6832 ( \6997 , \6992 , \6996 );
and \U$6833 ( \6998 , \2182 , \1578 );
and \U$6834 ( \6999 , \2366 , \1431 );
nor \U$6835 ( \7000 , \6998 , \6999 );
xnor \U$6836 ( \7001 , \7000 , \1436 );
xor \U$6837 ( \7002 , \6997 , \7001 );
xor \U$6838 ( \7003 , \6988 , \7002 );
and \U$6839 ( \7004 , \1192 , \2669 );
and \U$6840 ( \7005 , \1333 , \2538 );
nor \U$6841 ( \7006 , \7004 , \7005 );
xnor \U$6842 ( \7007 , \7006 , \2534 );
and \U$6843 ( \7008 , \474 , \3103 );
and \U$6844 ( \7009 , \1147 , \2934 );
nor \U$6845 ( \7010 , \7008 , \7009 );
xnor \U$6846 ( \7011 , \7010 , \2839 );
xor \U$6847 ( \7012 , \7007 , \7011 );
and \U$6848 ( \7013 , \307 , \3357 );
and \U$6849 ( \7014 , \412 , \3255 );
nor \U$6850 ( \7015 , \7013 , \7014 );
xnor \U$6851 ( \7016 , \7015 , \3156 );
xor \U$6852 ( \7017 , \7012 , \7016 );
xor \U$6853 ( \7018 , \7003 , \7017 );
xor \U$6854 ( \7019 , \6974 , \7018 );
and \U$6855 ( \7020 , \232 , \5011 );
and \U$6856 ( \7021 , \209 , \4878 );
nor \U$6857 ( \7022 , \7020 , \7021 );
xnor \U$6858 ( \7023 , \7022 , \4762 );
and \U$6859 ( \7024 , \247 , \5485 );
and \U$6860 ( \7025 , \224 , \5275 );
nor \U$6861 ( \7026 , \7024 , \7025 );
xnor \U$6862 ( \7027 , \7026 , \5169 );
xor \U$6863 ( \7028 , \7023 , \7027 );
and \U$6864 ( \7029 , \143 , \5996 );
and \U$6865 ( \7030 , \240 , \5695 );
nor \U$6866 ( \7031 , \7029 , \7030 );
xnor \U$6867 ( \7032 , \7031 , \5687 );
xor \U$6868 ( \7033 , \7028 , \7032 );
and \U$6869 ( \7034 , \185 , \3813 );
and \U$6870 ( \7035 , \261 , \3557 );
nor \U$6871 ( \7036 , \7034 , \7035 );
xnor \U$6872 ( \7037 , \7036 , \3562 );
and \U$6873 ( \7038 , \197 , \4132 );
and \U$6874 ( \7039 , \178 , \4012 );
nor \U$6875 ( \7040 , \7038 , \7039 );
xnor \U$6876 ( \7041 , \7040 , \3925 );
xor \U$6877 ( \7042 , \7037 , \7041 );
and \U$6878 ( \7043 , \217 , \4581 );
and \U$6879 ( \7044 , \189 , \4424 );
nor \U$6880 ( \7045 , \7043 , \7044 );
xnor \U$6881 ( \7046 , \7045 , \4377 );
xor \U$6882 ( \7047 , \7042 , \7046 );
xor \U$6883 ( \7048 , \7033 , \7047 );
and \U$6884 ( \7049 , \158 , \6401 );
and \U$6885 ( \7050 , \134 , \6143 );
nor \U$6886 ( \7051 , \7049 , \7050 );
xnor \U$6887 ( \7052 , \7051 , \6148 );
xor \U$6888 ( \7053 , \6677 , \6674 );
not \U$6889 ( \7054 , \6675 );
and \U$6890 ( \7055 , \7053 , \7054 );
and \U$6891 ( \7056 , \166 , \7055 );
and \U$6892 ( \7057 , \150 , \6675 );
nor \U$6893 ( \7058 , \7056 , \7057 );
xnor \U$6894 ( \7059 , \7058 , \6680 );
xor \U$6895 ( \7060 , \7052 , \7059 );
xor \U$6896 ( \7061 , \7048 , \7060 );
xor \U$6897 ( \7062 , \7019 , \7061 );
xor \U$6898 ( \7063 , \6929 , \7062 );
xor \U$6899 ( \7064 , \6880 , \7063 );
xor \U$6900 ( \7065 , \6851 , \7064 );
xor \U$6901 ( \7066 , \6842 , \7065 );
and \U$6902 ( \7067 , \6562 , \6583 );
and \U$6903 ( \7068 , \6583 , \6804 );
and \U$6904 ( \7069 , \6562 , \6804 );
or \U$6905 ( \7070 , \7067 , \7068 , \7069 );
xor \U$6906 ( \7071 , \7066 , \7070 );
and \U$6907 ( \7072 , \6805 , \6809 );
and \U$6908 ( \7073 , \6810 , \6813 );
or \U$6909 ( \7074 , \7072 , \7073 );
xor \U$6910 ( \7075 , \7071 , \7074 );
buf g5535_GF_PartitionCandidate( \7076_nG5535 , \7075 );
buf \U$6911 ( \7077 , \7076_nG5535 );
and \U$6912 ( \7078 , \6846 , \6850 );
and \U$6913 ( \7079 , \6850 , \7064 );
and \U$6914 ( \7080 , \6846 , \7064 );
or \U$6915 ( \7081 , \7078 , \7079 , \7080 );
and \U$6916 ( \7082 , \6824 , \6828 );
and \U$6917 ( \7083 , \6828 , \6840 );
and \U$6918 ( \7084 , \6824 , \6840 );
or \U$6919 ( \7085 , \7082 , \7083 , \7084 );
and \U$6920 ( \7086 , \6865 , \6879 );
and \U$6921 ( \7087 , \6879 , \7063 );
and \U$6922 ( \7088 , \6865 , \7063 );
or \U$6923 ( \7089 , \7086 , \7087 , \7088 );
xor \U$6924 ( \7090 , \7085 , \7089 );
and \U$6925 ( \7091 , \6898 , \6912 );
and \U$6926 ( \7092 , \6912 , \6927 );
and \U$6927 ( \7093 , \6898 , \6927 );
or \U$6928 ( \7094 , \7091 , \7092 , \7093 );
and \U$6929 ( \7095 , \6933 , \6937 );
and \U$6930 ( \7096 , \6937 , \6942 );
and \U$6931 ( \7097 , \6933 , \6942 );
or \U$6932 ( \7098 , \7095 , \7096 , \7097 );
and \U$6933 ( \7099 , \6948 , \6952 );
and \U$6934 ( \7100 , \6952 , \6957 );
and \U$6935 ( \7101 , \6948 , \6957 );
or \U$6936 ( \7102 , \7099 , \7100 , \7101 );
xor \U$6937 ( \7103 , \7098 , \7102 );
and \U$6938 ( \7104 , \6963 , \6967 );
and \U$6939 ( \7105 , \6967 , \6972 );
and \U$6940 ( \7106 , \6963 , \6972 );
or \U$6941 ( \7107 , \7104 , \7105 , \7106 );
xor \U$6942 ( \7108 , \7103 , \7107 );
xor \U$6943 ( \7109 , \7094 , \7108 );
and \U$6944 ( \7110 , \6978 , \6982 );
and \U$6945 ( \7111 , \6982 , \6987 );
and \U$6946 ( \7112 , \6978 , \6987 );
or \U$6947 ( \7113 , \7110 , \7111 , \7112 );
and \U$6948 ( \7114 , \6992 , \6996 );
and \U$6949 ( \7115 , \6996 , \7001 );
and \U$6950 ( \7116 , \6992 , \7001 );
or \U$6951 ( \7117 , \7114 , \7115 , \7116 );
xor \U$6952 ( \7118 , \7113 , \7117 );
and \U$6953 ( \7119 , \7007 , \7011 );
and \U$6954 ( \7120 , \7011 , \7016 );
and \U$6955 ( \7121 , \7007 , \7016 );
or \U$6956 ( \7122 , \7119 , \7120 , \7121 );
xor \U$6957 ( \7123 , \7118 , \7122 );
and \U$6958 ( \7124 , \7023 , \7027 );
and \U$6959 ( \7125 , \7027 , \7032 );
and \U$6960 ( \7126 , \7023 , \7032 );
or \U$6961 ( \7127 , \7124 , \7125 , \7126 );
and \U$6962 ( \7128 , \7037 , \7041 );
and \U$6963 ( \7129 , \7041 , \7046 );
and \U$6964 ( \7130 , \7037 , \7046 );
or \U$6965 ( \7131 , \7128 , \7129 , \7130 );
xor \U$6966 ( \7132 , \7127 , \7131 );
and \U$6967 ( \7133 , \7052 , \7059 );
xor \U$6968 ( \7134 , \7132 , \7133 );
xor \U$6969 ( \7135 , \7123 , \7134 );
buf \U$6970 ( \7136 , RIb560a98_12);
xor \U$6971 ( \7137 , \7136 , \6677 );
nand \U$6972 ( \7138 , \166 , \7137 );
buf \U$6973 ( \7139 , RIb560b10_11);
and \U$6974 ( \7140 , \7136 , \6677 );
not \U$6975 ( \7141 , \7140 );
and \U$6976 ( \7142 , \7139 , \7141 );
xnor \U$6977 ( \7143 , \7138 , \7142 );
and \U$6978 ( \7144 , \240 , \5996 );
and \U$6979 ( \7145 , \247 , \5695 );
nor \U$6980 ( \7146 , \7144 , \7145 );
xnor \U$6981 ( \7147 , \7146 , \5687 );
and \U$6982 ( \7148 , \134 , \6401 );
and \U$6983 ( \7149 , \143 , \6143 );
nor \U$6984 ( \7150 , \7148 , \7149 );
xnor \U$6985 ( \7151 , \7150 , \6148 );
xor \U$6986 ( \7152 , \7147 , \7151 );
and \U$6987 ( \7153 , \150 , \7055 );
and \U$6988 ( \7154 , \158 , \6675 );
nor \U$6989 ( \7155 , \7153 , \7154 );
xnor \U$6990 ( \7156 , \7155 , \6680 );
xor \U$6991 ( \7157 , \7152 , \7156 );
xor \U$6992 ( \7158 , \7143 , \7157 );
and \U$6993 ( \7159 , \189 , \4581 );
and \U$6994 ( \7160 , \197 , \4424 );
nor \U$6995 ( \7161 , \7159 , \7160 );
xnor \U$6996 ( \7162 , \7161 , \4377 );
and \U$6997 ( \7163 , \209 , \5011 );
and \U$6998 ( \7164 , \217 , \4878 );
nor \U$6999 ( \7165 , \7163 , \7164 );
xnor \U$7000 ( \7166 , \7165 , \4762 );
xor \U$7001 ( \7167 , \7162 , \7166 );
and \U$7002 ( \7168 , \224 , \5485 );
and \U$7003 ( \7169 , \232 , \5275 );
nor \U$7004 ( \7170 , \7168 , \7169 );
xnor \U$7005 ( \7171 , \7170 , \5169 );
xor \U$7006 ( \7172 , \7167 , \7171 );
xor \U$7007 ( \7173 , \7158 , \7172 );
xor \U$7008 ( \7174 , \7135 , \7173 );
xor \U$7009 ( \7175 , \7109 , \7174 );
xor \U$7010 ( \7176 , \7090 , \7175 );
xor \U$7011 ( \7177 , \7081 , \7176 );
and \U$7012 ( \7178 , \6855 , \6859 );
and \U$7013 ( \7179 , \6859 , \6864 );
and \U$7014 ( \7180 , \6855 , \6864 );
or \U$7015 ( \7181 , \7178 , \7179 , \7180 );
and \U$7016 ( \7182 , \6833 , \6837 );
and \U$7017 ( \7183 , \6837 , \6839 );
and \U$7018 ( \7184 , \6833 , \6839 );
or \U$7019 ( \7185 , \7182 , \7183 , \7184 );
xor \U$7020 ( \7186 , \7181 , \7185 );
and \U$7021 ( \7187 , \6974 , \7018 );
and \U$7022 ( \7188 , \7018 , \7061 );
and \U$7023 ( \7189 , \6974 , \7061 );
or \U$7024 ( \7190 , \7187 , \7188 , \7189 );
xor \U$7025 ( \7191 , \7186 , \7190 );
and \U$7026 ( \7192 , \6869 , \6873 );
and \U$7027 ( \7193 , \6873 , \6878 );
and \U$7028 ( \7194 , \6869 , \6878 );
or \U$7029 ( \7195 , \7192 , \7193 , \7194 );
and \U$7030 ( \7196 , \6884 , \6928 );
and \U$7031 ( \7197 , \6928 , \7062 );
and \U$7032 ( \7198 , \6884 , \7062 );
or \U$7033 ( \7199 , \7196 , \7197 , \7198 );
xor \U$7034 ( \7200 , \7195 , \7199 );
and \U$7035 ( \7201 , \6888 , \6892 );
and \U$7036 ( \7202 , \6892 , \6897 );
and \U$7037 ( \7203 , \6888 , \6897 );
or \U$7038 ( \7204 , \7201 , \7202 , \7203 );
and \U$7039 ( \7205 , \6902 , \6906 );
and \U$7040 ( \7206 , \6906 , \6911 );
and \U$7041 ( \7207 , \6902 , \6911 );
or \U$7042 ( \7208 , \7205 , \7206 , \7207 );
xor \U$7043 ( \7209 , \7204 , \7208 );
and \U$7044 ( \7210 , \6917 , \6921 );
and \U$7045 ( \7211 , \6921 , \6926 );
and \U$7046 ( \7212 , \6917 , \6926 );
or \U$7047 ( \7213 , \7210 , \7211 , \7212 );
xor \U$7048 ( \7214 , \7209 , \7213 );
and \U$7049 ( \7215 , \6943 , \6958 );
and \U$7050 ( \7216 , \6958 , \6973 );
and \U$7051 ( \7217 , \6943 , \6973 );
or \U$7052 ( \7218 , \7215 , \7216 , \7217 );
and \U$7053 ( \7219 , \6988 , \7002 );
and \U$7054 ( \7220 , \7002 , \7017 );
and \U$7055 ( \7221 , \6988 , \7017 );
or \U$7056 ( \7222 , \7219 , \7220 , \7221 );
xor \U$7057 ( \7223 , \7218 , \7222 );
and \U$7058 ( \7224 , \7033 , \7047 );
and \U$7059 ( \7225 , \7047 , \7060 );
and \U$7060 ( \7226 , \7033 , \7060 );
or \U$7061 ( \7227 , \7224 , \7225 , \7226 );
xor \U$7062 ( \7228 , \7223 , \7227 );
xor \U$7063 ( \7229 , \7214 , \7228 );
and \U$7064 ( \7230 , \6945 , \183 );
buf \U$7065 ( \7231 , RIb55ec98_76);
and \U$7066 ( \7232 , \7231 , \180 );
nor \U$7067 ( \7233 , \7230 , \7232 );
xnor \U$7068 ( \7234 , \7233 , \179 );
and \U$7069 ( \7235 , \6514 , \195 );
and \U$7070 ( \7236 , \6790 , \193 );
nor \U$7071 ( \7237 , \7235 , \7236 );
xnor \U$7072 ( \7238 , \7237 , \202 );
xor \U$7073 ( \7239 , \7234 , \7238 );
xor \U$7074 ( \7240 , \7239 , \7142 );
and \U$7075 ( \7241 , \6030 , \215 );
and \U$7076 ( \7242 , \6281 , \213 );
nor \U$7077 ( \7243 , \7241 , \7242 );
xnor \U$7078 ( \7244 , \7243 , \222 );
and \U$7079 ( \7245 , \5469 , \230 );
and \U$7080 ( \7246 , \5674 , \228 );
nor \U$7081 ( \7247 , \7245 , \7246 );
xnor \U$7082 ( \7248 , \7247 , \237 );
xor \U$7083 ( \7249 , \7244 , \7248 );
and \U$7084 ( \7250 , \4922 , \245 );
and \U$7085 ( \7251 , \5156 , \243 );
nor \U$7086 ( \7252 , \7250 , \7251 );
xnor \U$7087 ( \7253 , \7252 , \252 );
xor \U$7088 ( \7254 , \7249 , \7253 );
and \U$7089 ( \7255 , \4654 , \141 );
and \U$7090 ( \7256 , \4749 , \139 );
nor \U$7091 ( \7257 , \7255 , \7256 );
xnor \U$7092 ( \7258 , \7257 , \148 );
and \U$7093 ( \7259 , \4160 , \156 );
and \U$7094 ( \7260 , \4364 , \154 );
nor \U$7095 ( \7261 , \7259 , \7260 );
xnor \U$7096 ( \7262 , \7261 , \163 );
xor \U$7097 ( \7263 , \7258 , \7262 );
and \U$7098 ( \7264 , \3736 , \296 );
and \U$7099 ( \7265 , \3912 , \168 );
nor \U$7100 ( \7266 , \7264 , \7265 );
xnor \U$7101 ( \7267 , \7266 , \173 );
xor \U$7102 ( \7268 , \7263 , \7267 );
xor \U$7103 ( \7269 , \7254 , \7268 );
and \U$7104 ( \7270 , \3395 , \438 );
and \U$7105 ( \7271 , \3646 , \336 );
nor \U$7106 ( \7272 , \7270 , \7271 );
xnor \U$7107 ( \7273 , \7272 , \320 );
and \U$7108 ( \7274 , \3037 , \1086 );
and \U$7109 ( \7275 , \3143 , \508 );
nor \U$7110 ( \7276 , \7274 , \7275 );
xnor \U$7111 ( \7277 , \7276 , \487 );
xor \U$7112 ( \7278 , \7273 , \7277 );
and \U$7113 ( \7279 , \2757 , \1301 );
and \U$7114 ( \7280 , \2826 , \1246 );
nor \U$7115 ( \7281 , \7279 , \7280 );
xnor \U$7116 ( \7282 , \7281 , \1205 );
xor \U$7117 ( \7283 , \7278 , \7282 );
xor \U$7118 ( \7284 , \7269 , \7283 );
xor \U$7119 ( \7285 , \7240 , \7284 );
and \U$7120 ( \7286 , \412 , \3357 );
and \U$7121 ( \7287 , \474 , \3255 );
nor \U$7122 ( \7288 , \7286 , \7287 );
xnor \U$7123 ( \7289 , \7288 , \3156 );
and \U$7124 ( \7290 , \261 , \3813 );
and \U$7125 ( \7291 , \307 , \3557 );
nor \U$7126 ( \7292 , \7290 , \7291 );
xnor \U$7127 ( \7293 , \7292 , \3562 );
xor \U$7128 ( \7294 , \7289 , \7293 );
and \U$7129 ( \7295 , \178 , \4132 );
and \U$7130 ( \7296 , \185 , \4012 );
nor \U$7131 ( \7297 , \7295 , \7296 );
xnor \U$7132 ( \7298 , \7297 , \3925 );
xor \U$7133 ( \7299 , \7294 , \7298 );
and \U$7134 ( \7300 , \1601 , \2400 );
and \U$7135 ( \7301 , \1684 , \2246 );
nor \U$7136 ( \7302 , \7300 , \7301 );
xnor \U$7137 ( \7303 , \7302 , \2195 );
and \U$7138 ( \7304 , \1333 , \2669 );
and \U$7139 ( \7305 , \1484 , \2538 );
nor \U$7140 ( \7306 , \7304 , \7305 );
xnor \U$7141 ( \7307 , \7306 , \2534 );
xor \U$7142 ( \7308 , \7303 , \7307 );
and \U$7143 ( \7309 , \1147 , \3103 );
and \U$7144 ( \7310 , \1192 , \2934 );
nor \U$7145 ( \7311 , \7309 , \7310 );
xnor \U$7146 ( \7312 , \7311 , \2839 );
xor \U$7147 ( \7313 , \7308 , \7312 );
xor \U$7148 ( \7314 , \7299 , \7313 );
and \U$7149 ( \7315 , \2366 , \1578 );
and \U$7150 ( \7316 , \2521 , \1431 );
nor \U$7151 ( \7317 , \7315 , \7316 );
xnor \U$7152 ( \7318 , \7317 , \1436 );
and \U$7153 ( \7319 , \2090 , \1824 );
and \U$7154 ( \7320 , \2182 , \1739 );
nor \U$7155 ( \7321 , \7319 , \7320 );
xnor \U$7156 ( \7322 , \7321 , \1697 );
xor \U$7157 ( \7323 , \7318 , \7322 );
and \U$7158 ( \7324 , \1802 , \2121 );
and \U$7159 ( \7325 , \1948 , \2008 );
nor \U$7160 ( \7326 , \7324 , \7325 );
xnor \U$7161 ( \7327 , \7326 , \1961 );
xor \U$7162 ( \7328 , \7323 , \7327 );
xor \U$7163 ( \7329 , \7314 , \7328 );
xor \U$7164 ( \7330 , \7285 , \7329 );
xor \U$7165 ( \7331 , \7229 , \7330 );
xor \U$7166 ( \7332 , \7200 , \7331 );
xor \U$7167 ( \7333 , \7191 , \7332 );
xor \U$7168 ( \7334 , \7177 , \7333 );
and \U$7169 ( \7335 , \6820 , \6841 );
and \U$7170 ( \7336 , \6841 , \7065 );
and \U$7171 ( \7337 , \6820 , \7065 );
or \U$7172 ( \7338 , \7335 , \7336 , \7337 );
xor \U$7173 ( \7339 , \7334 , \7338 );
and \U$7174 ( \7340 , \7066 , \7070 );
and \U$7175 ( \7341 , \7071 , \7074 );
or \U$7176 ( \7342 , \7340 , \7341 );
xor \U$7177 ( \7343 , \7339 , \7342 );
buf g5533_GF_PartitionCandidate( \7344_nG5533 , \7343 );
buf \U$7178 ( \7345 , \7344_nG5533 );
and \U$7179 ( \7346 , \7085 , \7089 );
and \U$7180 ( \7347 , \7089 , \7175 );
and \U$7181 ( \7348 , \7085 , \7175 );
or \U$7182 ( \7349 , \7346 , \7347 , \7348 );
and \U$7183 ( \7350 , \7191 , \7332 );
xor \U$7184 ( \7351 , \7349 , \7350 );
and \U$7185 ( \7352 , \7195 , \7199 );
and \U$7186 ( \7353 , \7199 , \7331 );
and \U$7187 ( \7354 , \7195 , \7331 );
or \U$7188 ( \7355 , \7352 , \7353 , \7354 );
and \U$7189 ( \7356 , \7181 , \7185 );
and \U$7190 ( \7357 , \7185 , \7190 );
and \U$7191 ( \7358 , \7181 , \7190 );
or \U$7192 ( \7359 , \7356 , \7357 , \7358 );
and \U$7193 ( \7360 , \7094 , \7108 );
and \U$7194 ( \7361 , \7108 , \7174 );
and \U$7195 ( \7362 , \7094 , \7174 );
or \U$7196 ( \7363 , \7360 , \7361 , \7362 );
xor \U$7197 ( \7364 , \7359 , \7363 );
and \U$7198 ( \7365 , \7214 , \7228 );
and \U$7199 ( \7366 , \7228 , \7330 );
and \U$7200 ( \7367 , \7214 , \7330 );
or \U$7201 ( \7368 , \7365 , \7366 , \7367 );
xor \U$7202 ( \7369 , \7364 , \7368 );
xor \U$7203 ( \7370 , \7355 , \7369 );
and \U$7204 ( \7371 , \7204 , \7208 );
and \U$7205 ( \7372 , \7208 , \7213 );
and \U$7206 ( \7373 , \7204 , \7213 );
or \U$7207 ( \7374 , \7371 , \7372 , \7373 );
and \U$7208 ( \7375 , \7218 , \7222 );
and \U$7209 ( \7376 , \7222 , \7227 );
and \U$7210 ( \7377 , \7218 , \7227 );
or \U$7211 ( \7378 , \7375 , \7376 , \7377 );
xor \U$7212 ( \7379 , \7374 , \7378 );
and \U$7213 ( \7380 , \7240 , \7284 );
and \U$7214 ( \7381 , \7284 , \7329 );
and \U$7215 ( \7382 , \7240 , \7329 );
or \U$7216 ( \7383 , \7380 , \7381 , \7382 );
xor \U$7217 ( \7384 , \7379 , \7383 );
and \U$7218 ( \7385 , \7123 , \7134 );
and \U$7219 ( \7386 , \7134 , \7173 );
and \U$7220 ( \7387 , \7123 , \7173 );
or \U$7221 ( \7388 , \7385 , \7386 , \7387 );
and \U$7222 ( \7389 , \7303 , \7307 );
and \U$7223 ( \7390 , \7307 , \7312 );
and \U$7224 ( \7391 , \7303 , \7312 );
or \U$7225 ( \7392 , \7389 , \7390 , \7391 );
and \U$7226 ( \7393 , \7273 , \7277 );
and \U$7227 ( \7394 , \7277 , \7282 );
and \U$7228 ( \7395 , \7273 , \7282 );
or \U$7229 ( \7396 , \7393 , \7394 , \7395 );
xor \U$7230 ( \7397 , \7392 , \7396 );
and \U$7231 ( \7398 , \7318 , \7322 );
and \U$7232 ( \7399 , \7322 , \7327 );
and \U$7233 ( \7400 , \7318 , \7327 );
or \U$7234 ( \7401 , \7398 , \7399 , \7400 );
xor \U$7235 ( \7402 , \7397 , \7401 );
and \U$7236 ( \7403 , \7244 , \7248 );
and \U$7237 ( \7404 , \7248 , \7253 );
and \U$7238 ( \7405 , \7244 , \7253 );
or \U$7239 ( \7406 , \7403 , \7404 , \7405 );
and \U$7240 ( \7407 , \7234 , \7238 );
and \U$7241 ( \7408 , \7238 , \7142 );
and \U$7242 ( \7409 , \7234 , \7142 );
or \U$7243 ( \7410 , \7407 , \7408 , \7409 );
xor \U$7244 ( \7411 , \7406 , \7410 );
and \U$7245 ( \7412 , \7258 , \7262 );
and \U$7246 ( \7413 , \7262 , \7267 );
and \U$7247 ( \7414 , \7258 , \7267 );
or \U$7248 ( \7415 , \7412 , \7413 , \7414 );
xor \U$7249 ( \7416 , \7411 , \7415 );
xor \U$7250 ( \7417 , \7402 , \7416 );
and \U$7251 ( \7418 , \7147 , \7151 );
and \U$7252 ( \7419 , \7151 , \7156 );
and \U$7253 ( \7420 , \7147 , \7156 );
or \U$7254 ( \7421 , \7418 , \7419 , \7420 );
and \U$7255 ( \7422 , \7289 , \7293 );
and \U$7256 ( \7423 , \7293 , \7298 );
and \U$7257 ( \7424 , \7289 , \7298 );
or \U$7258 ( \7425 , \7422 , \7423 , \7424 );
xor \U$7259 ( \7426 , \7421 , \7425 );
and \U$7260 ( \7427 , \7162 , \7166 );
and \U$7261 ( \7428 , \7166 , \7171 );
and \U$7262 ( \7429 , \7162 , \7171 );
or \U$7263 ( \7430 , \7427 , \7428 , \7429 );
xor \U$7264 ( \7431 , \7426 , \7430 );
xor \U$7265 ( \7432 , \7417 , \7431 );
xor \U$7266 ( \7433 , \7388 , \7432 );
and \U$7267 ( \7434 , \1484 , \2669 );
and \U$7268 ( \7435 , \1601 , \2538 );
nor \U$7269 ( \7436 , \7434 , \7435 );
xnor \U$7270 ( \7437 , \7436 , \2534 );
and \U$7271 ( \7438 , \1192 , \3103 );
and \U$7272 ( \7439 , \1333 , \2934 );
nor \U$7273 ( \7440 , \7438 , \7439 );
xnor \U$7274 ( \7441 , \7440 , \2839 );
xor \U$7275 ( \7442 , \7437 , \7441 );
and \U$7276 ( \7443 , \474 , \3357 );
and \U$7277 ( \7444 , \1147 , \3255 );
nor \U$7278 ( \7445 , \7443 , \7444 );
xnor \U$7279 ( \7446 , \7445 , \3156 );
xor \U$7280 ( \7447 , \7442 , \7446 );
and \U$7281 ( \7448 , \2182 , \1824 );
and \U$7282 ( \7449 , \2366 , \1739 );
nor \U$7283 ( \7450 , \7448 , \7449 );
xnor \U$7284 ( \7451 , \7450 , \1697 );
and \U$7285 ( \7452 , \1948 , \2121 );
and \U$7286 ( \7453 , \2090 , \2008 );
nor \U$7287 ( \7454 , \7452 , \7453 );
xnor \U$7288 ( \7455 , \7454 , \1961 );
xor \U$7289 ( \7456 , \7451 , \7455 );
and \U$7290 ( \7457 , \1684 , \2400 );
and \U$7291 ( \7458 , \1802 , \2246 );
nor \U$7292 ( \7459 , \7457 , \7458 );
xnor \U$7293 ( \7460 , \7459 , \2195 );
xor \U$7294 ( \7461 , \7456 , \7460 );
xor \U$7295 ( \7462 , \7447 , \7461 );
and \U$7296 ( \7463 , \3143 , \1086 );
and \U$7297 ( \7464 , \3395 , \508 );
nor \U$7298 ( \7465 , \7463 , \7464 );
xnor \U$7299 ( \7466 , \7465 , \487 );
and \U$7300 ( \7467 , \2826 , \1301 );
and \U$7301 ( \7468 , \3037 , \1246 );
nor \U$7302 ( \7469 , \7467 , \7468 );
xnor \U$7303 ( \7470 , \7469 , \1205 );
xor \U$7304 ( \7471 , \7466 , \7470 );
and \U$7305 ( \7472 , \2521 , \1578 );
and \U$7306 ( \7473 , \2757 , \1431 );
nor \U$7307 ( \7474 , \7472 , \7473 );
xnor \U$7308 ( \7475 , \7474 , \1436 );
xor \U$7309 ( \7476 , \7471 , \7475 );
xor \U$7310 ( \7477 , \7462 , \7476 );
and \U$7311 ( \7478 , \143 , \6401 );
and \U$7312 ( \7479 , \240 , \6143 );
nor \U$7313 ( \7480 , \7478 , \7479 );
xnor \U$7314 ( \7481 , \7480 , \6148 );
and \U$7315 ( \7482 , \158 , \7055 );
and \U$7316 ( \7483 , \134 , \6675 );
nor \U$7317 ( \7484 , \7482 , \7483 );
xnor \U$7318 ( \7485 , \7484 , \6680 );
xor \U$7319 ( \7486 , \7481 , \7485 );
xor \U$7320 ( \7487 , \7139 , \7136 );
not \U$7321 ( \7488 , \7137 );
and \U$7322 ( \7489 , \7487 , \7488 );
and \U$7323 ( \7490 , \166 , \7489 );
and \U$7324 ( \7491 , \150 , \7137 );
nor \U$7325 ( \7492 , \7490 , \7491 );
xnor \U$7326 ( \7493 , \7492 , \7142 );
xor \U$7327 ( \7494 , \7486 , \7493 );
and \U$7328 ( \7495 , \307 , \3813 );
and \U$7329 ( \7496 , \412 , \3557 );
nor \U$7330 ( \7497 , \7495 , \7496 );
xnor \U$7331 ( \7498 , \7497 , \3562 );
and \U$7332 ( \7499 , \185 , \4132 );
and \U$7333 ( \7500 , \261 , \4012 );
nor \U$7334 ( \7501 , \7499 , \7500 );
xnor \U$7335 ( \7502 , \7501 , \3925 );
xor \U$7336 ( \7503 , \7498 , \7502 );
and \U$7337 ( \7504 , \197 , \4581 );
and \U$7338 ( \7505 , \178 , \4424 );
nor \U$7339 ( \7506 , \7504 , \7505 );
xnor \U$7340 ( \7507 , \7506 , \4377 );
xor \U$7341 ( \7508 , \7503 , \7507 );
xor \U$7342 ( \7509 , \7494 , \7508 );
and \U$7343 ( \7510 , \217 , \5011 );
and \U$7344 ( \7511 , \189 , \4878 );
nor \U$7345 ( \7512 , \7510 , \7511 );
xnor \U$7346 ( \7513 , \7512 , \4762 );
and \U$7347 ( \7514 , \232 , \5485 );
and \U$7348 ( \7515 , \209 , \5275 );
nor \U$7349 ( \7516 , \7514 , \7515 );
xnor \U$7350 ( \7517 , \7516 , \5169 );
xor \U$7351 ( \7518 , \7513 , \7517 );
and \U$7352 ( \7519 , \247 , \5996 );
and \U$7353 ( \7520 , \224 , \5695 );
nor \U$7354 ( \7521 , \7519 , \7520 );
xnor \U$7355 ( \7522 , \7521 , \5687 );
xor \U$7356 ( \7523 , \7518 , \7522 );
xor \U$7357 ( \7524 , \7509 , \7523 );
xor \U$7358 ( \7525 , \7477 , \7524 );
and \U$7359 ( \7526 , \5674 , \230 );
and \U$7360 ( \7527 , \6030 , \228 );
nor \U$7361 ( \7528 , \7526 , \7527 );
xnor \U$7362 ( \7529 , \7528 , \237 );
and \U$7363 ( \7530 , \5156 , \245 );
and \U$7364 ( \7531 , \5469 , \243 );
nor \U$7365 ( \7532 , \7530 , \7531 );
xnor \U$7366 ( \7533 , \7532 , \252 );
xor \U$7367 ( \7534 , \7529 , \7533 );
and \U$7368 ( \7535 , \4749 , \141 );
and \U$7369 ( \7536 , \4922 , \139 );
nor \U$7370 ( \7537 , \7535 , \7536 );
xnor \U$7371 ( \7538 , \7537 , \148 );
xor \U$7372 ( \7539 , \7534 , \7538 );
and \U$7373 ( \7540 , \4364 , \156 );
and \U$7374 ( \7541 , \4654 , \154 );
nor \U$7375 ( \7542 , \7540 , \7541 );
xnor \U$7376 ( \7543 , \7542 , \163 );
and \U$7377 ( \7544 , \3912 , \296 );
and \U$7378 ( \7545 , \4160 , \168 );
nor \U$7379 ( \7546 , \7544 , \7545 );
xnor \U$7380 ( \7547 , \7546 , \173 );
xor \U$7381 ( \7548 , \7543 , \7547 );
and \U$7382 ( \7549 , \3646 , \438 );
and \U$7383 ( \7550 , \3736 , \336 );
nor \U$7384 ( \7551 , \7549 , \7550 );
xnor \U$7385 ( \7552 , \7551 , \320 );
xor \U$7386 ( \7553 , \7548 , \7552 );
xor \U$7387 ( \7554 , \7539 , \7553 );
and \U$7388 ( \7555 , \7231 , \183 );
buf \U$7389 ( \7556 , RIb55ed10_75);
and \U$7390 ( \7557 , \7556 , \180 );
nor \U$7391 ( \7558 , \7555 , \7557 );
xnor \U$7392 ( \7559 , \7558 , \179 );
and \U$7393 ( \7560 , \6790 , \195 );
and \U$7394 ( \7561 , \6945 , \193 );
nor \U$7395 ( \7562 , \7560 , \7561 );
xnor \U$7396 ( \7563 , \7562 , \202 );
xor \U$7397 ( \7564 , \7559 , \7563 );
and \U$7398 ( \7565 , \6281 , \215 );
and \U$7399 ( \7566 , \6514 , \213 );
nor \U$7400 ( \7567 , \7565 , \7566 );
xnor \U$7401 ( \7568 , \7567 , \222 );
xor \U$7402 ( \7569 , \7564 , \7568 );
xor \U$7403 ( \7570 , \7554 , \7569 );
xor \U$7404 ( \7571 , \7525 , \7570 );
xor \U$7405 ( \7572 , \7433 , \7571 );
xor \U$7406 ( \7573 , \7384 , \7572 );
and \U$7407 ( \7574 , \7113 , \7117 );
and \U$7408 ( \7575 , \7117 , \7122 );
and \U$7409 ( \7576 , \7113 , \7122 );
or \U$7410 ( \7577 , \7574 , \7575 , \7576 );
and \U$7411 ( \7578 , \7127 , \7131 );
and \U$7412 ( \7579 , \7131 , \7133 );
and \U$7413 ( \7580 , \7127 , \7133 );
or \U$7414 ( \7581 , \7578 , \7579 , \7580 );
xor \U$7415 ( \7582 , \7577 , \7581 );
and \U$7416 ( \7583 , \7098 , \7102 );
and \U$7417 ( \7584 , \7102 , \7107 );
and \U$7418 ( \7585 , \7098 , \7107 );
or \U$7419 ( \7586 , \7583 , \7584 , \7585 );
xor \U$7420 ( \7587 , \7582 , \7586 );
and \U$7421 ( \7588 , \7254 , \7268 );
and \U$7422 ( \7589 , \7268 , \7283 );
and \U$7423 ( \7590 , \7254 , \7283 );
or \U$7424 ( \7591 , \7588 , \7589 , \7590 );
and \U$7425 ( \7592 , \7143 , \7157 );
and \U$7426 ( \7593 , \7157 , \7172 );
and \U$7427 ( \7594 , \7143 , \7172 );
or \U$7428 ( \7595 , \7592 , \7593 , \7594 );
xor \U$7429 ( \7596 , \7591 , \7595 );
and \U$7430 ( \7597 , \7299 , \7313 );
and \U$7431 ( \7598 , \7313 , \7328 );
and \U$7432 ( \7599 , \7299 , \7328 );
or \U$7433 ( \7600 , \7597 , \7598 , \7599 );
xor \U$7434 ( \7601 , \7596 , \7600 );
xor \U$7435 ( \7602 , \7587 , \7601 );
xor \U$7436 ( \7603 , \7573 , \7602 );
xor \U$7437 ( \7604 , \7370 , \7603 );
xor \U$7438 ( \7605 , \7351 , \7604 );
and \U$7439 ( \7606 , \7081 , \7176 );
and \U$7440 ( \7607 , \7176 , \7333 );
and \U$7441 ( \7608 , \7081 , \7333 );
or \U$7442 ( \7609 , \7606 , \7607 , \7608 );
xor \U$7443 ( \7610 , \7605 , \7609 );
and \U$7444 ( \7611 , \7334 , \7338 );
and \U$7445 ( \7612 , \7339 , \7342 );
or \U$7446 ( \7613 , \7611 , \7612 );
xor \U$7447 ( \7614 , \7610 , \7613 );
buf g5531_GF_PartitionCandidate( \7615_nG5531 , \7614 );
buf \U$7448 ( \7616 , \7615_nG5531 );
and \U$7449 ( \7617 , \7355 , \7369 );
and \U$7450 ( \7618 , \7369 , \7603 );
and \U$7451 ( \7619 , \7355 , \7603 );
or \U$7452 ( \7620 , \7617 , \7618 , \7619 );
and \U$7453 ( \7621 , \7374 , \7378 );
and \U$7454 ( \7622 , \7378 , \7383 );
and \U$7455 ( \7623 , \7374 , \7383 );
or \U$7456 ( \7624 , \7621 , \7622 , \7623 );
and \U$7457 ( \7625 , \7388 , \7432 );
and \U$7458 ( \7626 , \7432 , \7571 );
and \U$7459 ( \7627 , \7388 , \7571 );
or \U$7460 ( \7628 , \7625 , \7626 , \7627 );
xor \U$7461 ( \7629 , \7624 , \7628 );
and \U$7462 ( \7630 , \7587 , \7601 );
xor \U$7463 ( \7631 , \7629 , \7630 );
xor \U$7464 ( \7632 , \7620 , \7631 );
and \U$7465 ( \7633 , \7359 , \7363 );
and \U$7466 ( \7634 , \7363 , \7368 );
and \U$7467 ( \7635 , \7359 , \7368 );
or \U$7468 ( \7636 , \7633 , \7634 , \7635 );
and \U$7469 ( \7637 , \7384 , \7572 );
and \U$7470 ( \7638 , \7572 , \7602 );
and \U$7471 ( \7639 , \7384 , \7602 );
or \U$7472 ( \7640 , \7637 , \7638 , \7639 );
xor \U$7473 ( \7641 , \7636 , \7640 );
and \U$7474 ( \7642 , \7577 , \7581 );
and \U$7475 ( \7643 , \7581 , \7586 );
and \U$7476 ( \7644 , \7577 , \7586 );
or \U$7477 ( \7645 , \7642 , \7643 , \7644 );
and \U$7478 ( \7646 , \7591 , \7595 );
and \U$7479 ( \7647 , \7595 , \7600 );
and \U$7480 ( \7648 , \7591 , \7600 );
or \U$7481 ( \7649 , \7646 , \7647 , \7648 );
xor \U$7482 ( \7650 , \7645 , \7649 );
and \U$7483 ( \7651 , \7477 , \7524 );
and \U$7484 ( \7652 , \7524 , \7570 );
and \U$7485 ( \7653 , \7477 , \7570 );
or \U$7486 ( \7654 , \7651 , \7652 , \7653 );
xor \U$7487 ( \7655 , \7650 , \7654 );
and \U$7488 ( \7656 , \7447 , \7461 );
and \U$7489 ( \7657 , \7461 , \7476 );
and \U$7490 ( \7658 , \7447 , \7476 );
or \U$7491 ( \7659 , \7656 , \7657 , \7658 );
and \U$7492 ( \7660 , \7494 , \7508 );
and \U$7493 ( \7661 , \7508 , \7523 );
and \U$7494 ( \7662 , \7494 , \7523 );
or \U$7495 ( \7663 , \7660 , \7661 , \7662 );
xor \U$7496 ( \7664 , \7659 , \7663 );
and \U$7497 ( \7665 , \7539 , \7553 );
and \U$7498 ( \7666 , \7553 , \7569 );
and \U$7499 ( \7667 , \7539 , \7569 );
or \U$7500 ( \7668 , \7665 , \7666 , \7667 );
xor \U$7501 ( \7669 , \7664 , \7668 );
and \U$7502 ( \7670 , \7392 , \7396 );
and \U$7503 ( \7671 , \7396 , \7401 );
and \U$7504 ( \7672 , \7392 , \7401 );
or \U$7505 ( \7673 , \7670 , \7671 , \7672 );
and \U$7506 ( \7674 , \7406 , \7410 );
and \U$7507 ( \7675 , \7410 , \7415 );
and \U$7508 ( \7676 , \7406 , \7415 );
or \U$7509 ( \7677 , \7674 , \7675 , \7676 );
xor \U$7510 ( \7678 , \7673 , \7677 );
and \U$7511 ( \7679 , \7421 , \7425 );
and \U$7512 ( \7680 , \7425 , \7430 );
and \U$7513 ( \7681 , \7421 , \7430 );
or \U$7514 ( \7682 , \7679 , \7680 , \7681 );
xor \U$7515 ( \7683 , \7678 , \7682 );
xor \U$7516 ( \7684 , \7669 , \7683 );
and \U$7517 ( \7685 , \6514 , \215 );
and \U$7518 ( \7686 , \6790 , \213 );
nor \U$7519 ( \7687 , \7685 , \7686 );
xnor \U$7520 ( \7688 , \7687 , \222 );
and \U$7521 ( \7689 , \6030 , \230 );
and \U$7522 ( \7690 , \6281 , \228 );
nor \U$7523 ( \7691 , \7689 , \7690 );
xnor \U$7524 ( \7692 , \7691 , \237 );
xor \U$7525 ( \7693 , \7688 , \7692 );
and \U$7526 ( \7694 , \5469 , \245 );
and \U$7527 ( \7695 , \5674 , \243 );
nor \U$7528 ( \7696 , \7694 , \7695 );
xnor \U$7529 ( \7697 , \7696 , \252 );
xor \U$7530 ( \7698 , \7693 , \7697 );
and \U$7531 ( \7699 , \7556 , \183 );
buf \U$7532 ( \7700 , RIb55ed88_74);
and \U$7533 ( \7701 , \7700 , \180 );
nor \U$7534 ( \7702 , \7699 , \7701 );
xnor \U$7535 ( \7703 , \7702 , \179 );
and \U$7536 ( \7704 , \6945 , \195 );
and \U$7537 ( \7705 , \7231 , \193 );
nor \U$7538 ( \7706 , \7704 , \7705 );
xnor \U$7539 ( \7707 , \7706 , \202 );
xor \U$7540 ( \7708 , \7703 , \7707 );
buf \U$7541 ( \7709 , RIb560c00_9);
buf \U$7542 ( \7710 , RIb560b88_10);
and \U$7543 ( \7711 , \7710 , \7139 );
not \U$7544 ( \7712 , \7711 );
and \U$7545 ( \7713 , \7709 , \7712 );
xor \U$7546 ( \7714 , \7708 , \7713 );
xor \U$7547 ( \7715 , \7698 , \7714 );
and \U$7548 ( \7716 , \4922 , \141 );
and \U$7549 ( \7717 , \5156 , \139 );
nor \U$7550 ( \7718 , \7716 , \7717 );
xnor \U$7551 ( \7719 , \7718 , \148 );
and \U$7552 ( \7720 , \4654 , \156 );
and \U$7553 ( \7721 , \4749 , \154 );
nor \U$7554 ( \7722 , \7720 , \7721 );
xnor \U$7555 ( \7723 , \7722 , \163 );
xor \U$7556 ( \7724 , \7719 , \7723 );
and \U$7557 ( \7725 , \4160 , \296 );
and \U$7558 ( \7726 , \4364 , \168 );
nor \U$7559 ( \7727 , \7725 , \7726 );
xnor \U$7560 ( \7728 , \7727 , \173 );
xor \U$7561 ( \7729 , \7724 , \7728 );
and \U$7562 ( \7730 , \2757 , \1578 );
and \U$7563 ( \7731 , \2826 , \1431 );
nor \U$7564 ( \7732 , \7730 , \7731 );
xnor \U$7565 ( \7733 , \7732 , \1436 );
and \U$7566 ( \7734 , \2366 , \1824 );
and \U$7567 ( \7735 , \2521 , \1739 );
nor \U$7568 ( \7736 , \7734 , \7735 );
xnor \U$7569 ( \7737 , \7736 , \1697 );
xor \U$7570 ( \7738 , \7733 , \7737 );
and \U$7571 ( \7739 , \2090 , \2121 );
and \U$7572 ( \7740 , \2182 , \2008 );
nor \U$7573 ( \7741 , \7739 , \7740 );
xnor \U$7574 ( \7742 , \7741 , \1961 );
xor \U$7575 ( \7743 , \7738 , \7742 );
xor \U$7576 ( \7744 , \7729 , \7743 );
and \U$7577 ( \7745 , \3736 , \438 );
and \U$7578 ( \7746 , \3912 , \336 );
nor \U$7579 ( \7747 , \7745 , \7746 );
xnor \U$7580 ( \7748 , \7747 , \320 );
and \U$7581 ( \7749 , \3395 , \1086 );
and \U$7582 ( \7750 , \3646 , \508 );
nor \U$7583 ( \7751 , \7749 , \7750 );
xnor \U$7584 ( \7752 , \7751 , \487 );
xor \U$7585 ( \7753 , \7748 , \7752 );
and \U$7586 ( \7754 , \3037 , \1301 );
and \U$7587 ( \7755 , \3143 , \1246 );
nor \U$7588 ( \7756 , \7754 , \7755 );
xnor \U$7589 ( \7757 , \7756 , \1205 );
xor \U$7590 ( \7758 , \7753 , \7757 );
xor \U$7591 ( \7759 , \7744 , \7758 );
xor \U$7592 ( \7760 , \7715 , \7759 );
xor \U$7593 ( \7761 , \7684 , \7760 );
xor \U$7594 ( \7762 , \7655 , \7761 );
and \U$7595 ( \7763 , \7402 , \7416 );
and \U$7596 ( \7764 , \7416 , \7431 );
and \U$7597 ( \7765 , \7402 , \7431 );
or \U$7598 ( \7766 , \7763 , \7764 , \7765 );
and \U$7599 ( \7767 , \7481 , \7485 );
and \U$7600 ( \7768 , \7485 , \7493 );
and \U$7601 ( \7769 , \7481 , \7493 );
or \U$7602 ( \7770 , \7767 , \7768 , \7769 );
and \U$7603 ( \7771 , \7498 , \7502 );
and \U$7604 ( \7772 , \7502 , \7507 );
and \U$7605 ( \7773 , \7498 , \7507 );
or \U$7606 ( \7774 , \7771 , \7772 , \7773 );
xor \U$7607 ( \7775 , \7770 , \7774 );
and \U$7608 ( \7776 , \7513 , \7517 );
and \U$7609 ( \7777 , \7517 , \7522 );
and \U$7610 ( \7778 , \7513 , \7522 );
or \U$7611 ( \7779 , \7776 , \7777 , \7778 );
xor \U$7612 ( \7780 , \7775 , \7779 );
and \U$7613 ( \7781 , \1802 , \2400 );
and \U$7614 ( \7782 , \1948 , \2246 );
nor \U$7615 ( \7783 , \7781 , \7782 );
xnor \U$7616 ( \7784 , \7783 , \2195 );
and \U$7617 ( \7785 , \1601 , \2669 );
and \U$7618 ( \7786 , \1684 , \2538 );
nor \U$7619 ( \7787 , \7785 , \7786 );
xnor \U$7620 ( \7788 , \7787 , \2534 );
xor \U$7621 ( \7789 , \7784 , \7788 );
and \U$7622 ( \7790 , \1333 , \3103 );
and \U$7623 ( \7791 , \1484 , \2934 );
nor \U$7624 ( \7792 , \7790 , \7791 );
xnor \U$7625 ( \7793 , \7792 , \2839 );
xor \U$7626 ( \7794 , \7789 , \7793 );
and \U$7627 ( \7795 , \1147 , \3357 );
and \U$7628 ( \7796 , \1192 , \3255 );
nor \U$7629 ( \7797 , \7795 , \7796 );
xnor \U$7630 ( \7798 , \7797 , \3156 );
and \U$7631 ( \7799 , \412 , \3813 );
and \U$7632 ( \7800 , \474 , \3557 );
nor \U$7633 ( \7801 , \7799 , \7800 );
xnor \U$7634 ( \7802 , \7801 , \3562 );
xor \U$7635 ( \7803 , \7798 , \7802 );
and \U$7636 ( \7804 , \261 , \4132 );
and \U$7637 ( \7805 , \307 , \4012 );
nor \U$7638 ( \7806 , \7804 , \7805 );
xnor \U$7639 ( \7807 , \7806 , \3925 );
xor \U$7640 ( \7808 , \7803 , \7807 );
xor \U$7641 ( \7809 , \7794 , \7808 );
and \U$7642 ( \7810 , \178 , \4581 );
and \U$7643 ( \7811 , \185 , \4424 );
nor \U$7644 ( \7812 , \7810 , \7811 );
xnor \U$7645 ( \7813 , \7812 , \4377 );
and \U$7646 ( \7814 , \189 , \5011 );
and \U$7647 ( \7815 , \197 , \4878 );
nor \U$7648 ( \7816 , \7814 , \7815 );
xnor \U$7649 ( \7817 , \7816 , \4762 );
xor \U$7650 ( \7818 , \7813 , \7817 );
and \U$7651 ( \7819 , \209 , \5485 );
and \U$7652 ( \7820 , \217 , \5275 );
nor \U$7653 ( \7821 , \7819 , \7820 );
xnor \U$7654 ( \7822 , \7821 , \5169 );
xor \U$7655 ( \7823 , \7818 , \7822 );
xor \U$7656 ( \7824 , \7809 , \7823 );
xor \U$7657 ( \7825 , \7780 , \7824 );
and \U$7658 ( \7826 , \150 , \7489 );
and \U$7659 ( \7827 , \158 , \7137 );
nor \U$7660 ( \7828 , \7826 , \7827 );
xnor \U$7661 ( \7829 , \7828 , \7142 );
xor \U$7662 ( \7830 , \7710 , \7139 );
nand \U$7663 ( \7831 , \166 , \7830 );
xnor \U$7664 ( \7832 , \7831 , \7713 );
xor \U$7665 ( \7833 , \7829 , \7832 );
and \U$7666 ( \7834 , \224 , \5996 );
and \U$7667 ( \7835 , \232 , \5695 );
nor \U$7668 ( \7836 , \7834 , \7835 );
xnor \U$7669 ( \7837 , \7836 , \5687 );
and \U$7670 ( \7838 , \240 , \6401 );
and \U$7671 ( \7839 , \247 , \6143 );
nor \U$7672 ( \7840 , \7838 , \7839 );
xnor \U$7673 ( \7841 , \7840 , \6148 );
xor \U$7674 ( \7842 , \7837 , \7841 );
and \U$7675 ( \7843 , \134 , \7055 );
and \U$7676 ( \7844 , \143 , \6675 );
nor \U$7677 ( \7845 , \7843 , \7844 );
xnor \U$7678 ( \7846 , \7845 , \6680 );
xor \U$7679 ( \7847 , \7842 , \7846 );
xor \U$7680 ( \7848 , \7833 , \7847 );
xor \U$7681 ( \7849 , \7825 , \7848 );
xor \U$7682 ( \7850 , \7766 , \7849 );
and \U$7683 ( \7851 , \7529 , \7533 );
and \U$7684 ( \7852 , \7533 , \7538 );
and \U$7685 ( \7853 , \7529 , \7538 );
or \U$7686 ( \7854 , \7851 , \7852 , \7853 );
and \U$7687 ( \7855 , \7543 , \7547 );
and \U$7688 ( \7856 , \7547 , \7552 );
and \U$7689 ( \7857 , \7543 , \7552 );
or \U$7690 ( \7858 , \7855 , \7856 , \7857 );
xor \U$7691 ( \7859 , \7854 , \7858 );
and \U$7692 ( \7860 , \7559 , \7563 );
and \U$7693 ( \7861 , \7563 , \7568 );
and \U$7694 ( \7862 , \7559 , \7568 );
or \U$7695 ( \7863 , \7860 , \7861 , \7862 );
xor \U$7696 ( \7864 , \7859 , \7863 );
and \U$7697 ( \7865 , \7437 , \7441 );
and \U$7698 ( \7866 , \7441 , \7446 );
and \U$7699 ( \7867 , \7437 , \7446 );
or \U$7700 ( \7868 , \7865 , \7866 , \7867 );
and \U$7701 ( \7869 , \7451 , \7455 );
and \U$7702 ( \7870 , \7455 , \7460 );
and \U$7703 ( \7871 , \7451 , \7460 );
or \U$7704 ( \7872 , \7869 , \7870 , \7871 );
xor \U$7705 ( \7873 , \7868 , \7872 );
and \U$7706 ( \7874 , \7466 , \7470 );
and \U$7707 ( \7875 , \7470 , \7475 );
and \U$7708 ( \7876 , \7466 , \7475 );
or \U$7709 ( \7877 , \7874 , \7875 , \7876 );
xor \U$7710 ( \7878 , \7873 , \7877 );
xor \U$7711 ( \7879 , \7864 , \7878 );
xor \U$7712 ( \7880 , \7850 , \7879 );
xor \U$7713 ( \7881 , \7762 , \7880 );
xor \U$7714 ( \7882 , \7641 , \7881 );
xor \U$7715 ( \7883 , \7632 , \7882 );
and \U$7716 ( \7884 , \7349 , \7350 );
and \U$7717 ( \7885 , \7350 , \7604 );
and \U$7718 ( \7886 , \7349 , \7604 );
or \U$7719 ( \7887 , \7884 , \7885 , \7886 );
xor \U$7720 ( \7888 , \7883 , \7887 );
and \U$7721 ( \7889 , \7605 , \7609 );
and \U$7722 ( \7890 , \7610 , \7613 );
or \U$7723 ( \7891 , \7889 , \7890 );
xor \U$7724 ( \7892 , \7888 , \7891 );
buf g552f_GF_PartitionCandidate( \7893_nG552f , \7892 );
buf \U$7725 ( \7894 , \7893_nG552f );
and \U$7726 ( \7895 , \7636 , \7640 );
and \U$7727 ( \7896 , \7640 , \7881 );
and \U$7728 ( \7897 , \7636 , \7881 );
or \U$7729 ( \7898 , \7895 , \7896 , \7897 );
and \U$7730 ( \7899 , \7624 , \7628 );
and \U$7731 ( \7900 , \7628 , \7630 );
and \U$7732 ( \7901 , \7624 , \7630 );
or \U$7733 ( \7902 , \7899 , \7900 , \7901 );
and \U$7734 ( \7903 , \7655 , \7761 );
and \U$7735 ( \7904 , \7761 , \7880 );
and \U$7736 ( \7905 , \7655 , \7880 );
or \U$7737 ( \7906 , \7903 , \7904 , \7905 );
xor \U$7738 ( \7907 , \7902 , \7906 );
and \U$7739 ( \7908 , \7659 , \7663 );
and \U$7740 ( \7909 , \7663 , \7668 );
and \U$7741 ( \7910 , \7659 , \7668 );
or \U$7742 ( \7911 , \7908 , \7909 , \7910 );
and \U$7743 ( \7912 , \7673 , \7677 );
and \U$7744 ( \7913 , \7677 , \7682 );
and \U$7745 ( \7914 , \7673 , \7682 );
or \U$7746 ( \7915 , \7912 , \7913 , \7914 );
xor \U$7747 ( \7916 , \7911 , \7915 );
and \U$7748 ( \7917 , \7698 , \7714 );
and \U$7749 ( \7918 , \7714 , \7759 );
and \U$7750 ( \7919 , \7698 , \7759 );
or \U$7751 ( \7920 , \7917 , \7918 , \7919 );
xor \U$7752 ( \7921 , \7916 , \7920 );
xor \U$7753 ( \7922 , \7907 , \7921 );
xor \U$7754 ( \7923 , \7898 , \7922 );
and \U$7755 ( \7924 , \7645 , \7649 );
and \U$7756 ( \7925 , \7649 , \7654 );
and \U$7757 ( \7926 , \7645 , \7654 );
or \U$7758 ( \7927 , \7924 , \7925 , \7926 );
and \U$7759 ( \7928 , \7669 , \7683 );
and \U$7760 ( \7929 , \7683 , \7760 );
and \U$7761 ( \7930 , \7669 , \7760 );
or \U$7762 ( \7931 , \7928 , \7929 , \7930 );
xor \U$7763 ( \7932 , \7927 , \7931 );
and \U$7764 ( \7933 , \7766 , \7849 );
and \U$7765 ( \7934 , \7849 , \7879 );
and \U$7766 ( \7935 , \7766 , \7879 );
or \U$7767 ( \7936 , \7933 , \7934 , \7935 );
xor \U$7768 ( \7937 , \7932 , \7936 );
and \U$7769 ( \7938 , \7770 , \7774 );
and \U$7770 ( \7939 , \7774 , \7779 );
and \U$7771 ( \7940 , \7770 , \7779 );
or \U$7772 ( \7941 , \7938 , \7939 , \7940 );
and \U$7773 ( \7942 , \7854 , \7858 );
and \U$7774 ( \7943 , \7858 , \7863 );
and \U$7775 ( \7944 , \7854 , \7863 );
or \U$7776 ( \7945 , \7942 , \7943 , \7944 );
xor \U$7777 ( \7946 , \7941 , \7945 );
and \U$7778 ( \7947 , \7868 , \7872 );
and \U$7779 ( \7948 , \7872 , \7877 );
and \U$7780 ( \7949 , \7868 , \7877 );
or \U$7781 ( \7950 , \7947 , \7948 , \7949 );
xor \U$7782 ( \7951 , \7946 , \7950 );
and \U$7783 ( \7952 , \7780 , \7824 );
and \U$7784 ( \7953 , \7824 , \7848 );
and \U$7785 ( \7954 , \7780 , \7848 );
or \U$7786 ( \7955 , \7952 , \7953 , \7954 );
and \U$7787 ( \7956 , \7864 , \7878 );
xor \U$7788 ( \7957 , \7955 , \7956 );
and \U$7789 ( \7958 , \7719 , \7723 );
and \U$7790 ( \7959 , \7723 , \7728 );
and \U$7791 ( \7960 , \7719 , \7728 );
or \U$7792 ( \7961 , \7958 , \7959 , \7960 );
and \U$7793 ( \7962 , \7688 , \7692 );
and \U$7794 ( \7963 , \7692 , \7697 );
and \U$7795 ( \7964 , \7688 , \7697 );
or \U$7796 ( \7965 , \7962 , \7963 , \7964 );
xor \U$7797 ( \7966 , \7961 , \7965 );
and \U$7798 ( \7967 , \7703 , \7707 );
and \U$7799 ( \7968 , \7707 , \7713 );
and \U$7800 ( \7969 , \7703 , \7713 );
or \U$7801 ( \7970 , \7967 , \7968 , \7969 );
xor \U$7802 ( \7971 , \7966 , \7970 );
xor \U$7803 ( \7972 , \7957 , \7971 );
xor \U$7804 ( \7973 , \7951 , \7972 );
and \U$7805 ( \7974 , \7794 , \7808 );
and \U$7806 ( \7975 , \7808 , \7823 );
and \U$7807 ( \7976 , \7794 , \7823 );
or \U$7808 ( \7977 , \7974 , \7975 , \7976 );
and \U$7809 ( \7978 , \7829 , \7832 );
and \U$7810 ( \7979 , \7832 , \7847 );
and \U$7811 ( \7980 , \7829 , \7847 );
or \U$7812 ( \7981 , \7978 , \7979 , \7980 );
xor \U$7813 ( \7982 , \7977 , \7981 );
and \U$7814 ( \7983 , \7729 , \7743 );
and \U$7815 ( \7984 , \7743 , \7758 );
and \U$7816 ( \7985 , \7729 , \7758 );
or \U$7817 ( \7986 , \7983 , \7984 , \7985 );
xor \U$7818 ( \7987 , \7982 , \7986 );
and \U$7819 ( \7988 , \7837 , \7841 );
and \U$7820 ( \7989 , \7841 , \7846 );
and \U$7821 ( \7990 , \7837 , \7846 );
or \U$7822 ( \7991 , \7988 , \7989 , \7990 );
and \U$7823 ( \7992 , \7798 , \7802 );
and \U$7824 ( \7993 , \7802 , \7807 );
and \U$7825 ( \7994 , \7798 , \7807 );
or \U$7826 ( \7995 , \7992 , \7993 , \7994 );
xor \U$7827 ( \7996 , \7991 , \7995 );
and \U$7828 ( \7997 , \7813 , \7817 );
and \U$7829 ( \7998 , \7817 , \7822 );
and \U$7830 ( \7999 , \7813 , \7822 );
or \U$7831 ( \8000 , \7997 , \7998 , \7999 );
xor \U$7832 ( \8001 , \7996 , \8000 );
and \U$7833 ( \8002 , \7784 , \7788 );
and \U$7834 ( \8003 , \7788 , \7793 );
and \U$7835 ( \8004 , \7784 , \7793 );
or \U$7836 ( \8005 , \8002 , \8003 , \8004 );
and \U$7837 ( \8006 , \7733 , \7737 );
and \U$7838 ( \8007 , \7737 , \7742 );
and \U$7839 ( \8008 , \7733 , \7742 );
or \U$7840 ( \8009 , \8006 , \8007 , \8008 );
xor \U$7841 ( \8010 , \8005 , \8009 );
and \U$7842 ( \8011 , \7748 , \7752 );
and \U$7843 ( \8012 , \7752 , \7757 );
and \U$7844 ( \8013 , \7748 , \7757 );
or \U$7845 ( \8014 , \8011 , \8012 , \8013 );
xor \U$7846 ( \8015 , \8010 , \8014 );
xor \U$7847 ( \8016 , \8001 , \8015 );
xor \U$7848 ( \8017 , \7709 , \7710 );
not \U$7849 ( \8018 , \7830 );
and \U$7850 ( \8019 , \8017 , \8018 );
and \U$7851 ( \8020 , \166 , \8019 );
and \U$7852 ( \8021 , \150 , \7830 );
nor \U$7853 ( \8022 , \8020 , \8021 );
xnor \U$7854 ( \8023 , \8022 , \7713 );
and \U$7855 ( \8024 , \247 , \6401 );
and \U$7856 ( \8025 , \224 , \6143 );
nor \U$7857 ( \8026 , \8024 , \8025 );
xnor \U$7858 ( \8027 , \8026 , \6148 );
and \U$7859 ( \8028 , \143 , \7055 );
and \U$7860 ( \8029 , \240 , \6675 );
nor \U$7861 ( \8030 , \8028 , \8029 );
xnor \U$7862 ( \8031 , \8030 , \6680 );
xor \U$7863 ( \8032 , \8027 , \8031 );
and \U$7864 ( \8033 , \158 , \7489 );
and \U$7865 ( \8034 , \134 , \7137 );
nor \U$7866 ( \8035 , \8033 , \8034 );
xnor \U$7867 ( \8036 , \8035 , \7142 );
xor \U$7868 ( \8037 , \8032 , \8036 );
xor \U$7869 ( \8038 , \8023 , \8037 );
and \U$7870 ( \8039 , \197 , \5011 );
and \U$7871 ( \8040 , \178 , \4878 );
nor \U$7872 ( \8041 , \8039 , \8040 );
xnor \U$7873 ( \8042 , \8041 , \4762 );
and \U$7874 ( \8043 , \217 , \5485 );
and \U$7875 ( \8044 , \189 , \5275 );
nor \U$7876 ( \8045 , \8043 , \8044 );
xnor \U$7877 ( \8046 , \8045 , \5169 );
xor \U$7878 ( \8047 , \8042 , \8046 );
and \U$7879 ( \8048 , \232 , \5996 );
and \U$7880 ( \8049 , \209 , \5695 );
nor \U$7881 ( \8050 , \8048 , \8049 );
xnor \U$7882 ( \8051 , \8050 , \5687 );
xor \U$7883 ( \8052 , \8047 , \8051 );
xor \U$7884 ( \8053 , \8038 , \8052 );
xor \U$7885 ( \8054 , \8016 , \8053 );
xor \U$7886 ( \8055 , \7987 , \8054 );
and \U$7887 ( \8056 , \7700 , \183 );
buf \U$7888 ( \8057 , RIb55ee00_73);
and \U$7889 ( \8058 , \8057 , \180 );
nor \U$7890 ( \8059 , \8056 , \8058 );
xnor \U$7891 ( \8060 , \8059 , \179 );
and \U$7892 ( \8061 , \7231 , \195 );
and \U$7893 ( \8062 , \7556 , \193 );
nor \U$7894 ( \8063 , \8061 , \8062 );
xnor \U$7895 ( \8064 , \8063 , \202 );
xor \U$7896 ( \8065 , \8060 , \8064 );
and \U$7897 ( \8066 , \6790 , \215 );
and \U$7898 ( \8067 , \6945 , \213 );
nor \U$7899 ( \8068 , \8066 , \8067 );
xnor \U$7900 ( \8069 , \8068 , \222 );
xor \U$7901 ( \8070 , \8065 , \8069 );
and \U$7902 ( \8071 , \1684 , \2669 );
and \U$7903 ( \8072 , \1802 , \2538 );
nor \U$7904 ( \8073 , \8071 , \8072 );
xnor \U$7905 ( \8074 , \8073 , \2534 );
and \U$7906 ( \8075 , \1484 , \3103 );
and \U$7907 ( \8076 , \1601 , \2934 );
nor \U$7908 ( \8077 , \8075 , \8076 );
xnor \U$7909 ( \8078 , \8077 , \2839 );
xor \U$7910 ( \8079 , \8074 , \8078 );
and \U$7911 ( \8080 , \1192 , \3357 );
and \U$7912 ( \8081 , \1333 , \3255 );
nor \U$7913 ( \8082 , \8080 , \8081 );
xnor \U$7914 ( \8083 , \8082 , \3156 );
xor \U$7915 ( \8084 , \8079 , \8083 );
and \U$7916 ( \8085 , \2521 , \1824 );
and \U$7917 ( \8086 , \2757 , \1739 );
nor \U$7918 ( \8087 , \8085 , \8086 );
xnor \U$7919 ( \8088 , \8087 , \1697 );
and \U$7920 ( \8089 , \2182 , \2121 );
and \U$7921 ( \8090 , \2366 , \2008 );
nor \U$7922 ( \8091 , \8089 , \8090 );
xnor \U$7923 ( \8092 , \8091 , \1961 );
xor \U$7924 ( \8093 , \8088 , \8092 );
and \U$7925 ( \8094 , \1948 , \2400 );
and \U$7926 ( \8095 , \2090 , \2246 );
nor \U$7927 ( \8096 , \8094 , \8095 );
xnor \U$7928 ( \8097 , \8096 , \2195 );
xor \U$7929 ( \8098 , \8093 , \8097 );
xor \U$7930 ( \8099 , \8084 , \8098 );
and \U$7931 ( \8100 , \474 , \3813 );
and \U$7932 ( \8101 , \1147 , \3557 );
nor \U$7933 ( \8102 , \8100 , \8101 );
xnor \U$7934 ( \8103 , \8102 , \3562 );
and \U$7935 ( \8104 , \307 , \4132 );
and \U$7936 ( \8105 , \412 , \4012 );
nor \U$7937 ( \8106 , \8104 , \8105 );
xnor \U$7938 ( \8107 , \8106 , \3925 );
xor \U$7939 ( \8108 , \8103 , \8107 );
and \U$7940 ( \8109 , \185 , \4581 );
and \U$7941 ( \8110 , \261 , \4424 );
nor \U$7942 ( \8111 , \8109 , \8110 );
xnor \U$7943 ( \8112 , \8111 , \4377 );
xor \U$7944 ( \8113 , \8108 , \8112 );
xor \U$7945 ( \8114 , \8099 , \8113 );
xor \U$7946 ( \8115 , \8070 , \8114 );
and \U$7947 ( \8116 , \3646 , \1086 );
and \U$7948 ( \8117 , \3736 , \508 );
nor \U$7949 ( \8118 , \8116 , \8117 );
xnor \U$7950 ( \8119 , \8118 , \487 );
and \U$7951 ( \8120 , \3143 , \1301 );
and \U$7952 ( \8121 , \3395 , \1246 );
nor \U$7953 ( \8122 , \8120 , \8121 );
xnor \U$7954 ( \8123 , \8122 , \1205 );
xor \U$7955 ( \8124 , \8119 , \8123 );
and \U$7956 ( \8125 , \2826 , \1578 );
and \U$7957 ( \8126 , \3037 , \1431 );
nor \U$7958 ( \8127 , \8125 , \8126 );
xnor \U$7959 ( \8128 , \8127 , \1436 );
xor \U$7960 ( \8129 , \8124 , \8128 );
and \U$7961 ( \8130 , \4749 , \156 );
and \U$7962 ( \8131 , \4922 , \154 );
nor \U$7963 ( \8132 , \8130 , \8131 );
xnor \U$7964 ( \8133 , \8132 , \163 );
and \U$7965 ( \8134 , \4364 , \296 );
and \U$7966 ( \8135 , \4654 , \168 );
nor \U$7967 ( \8136 , \8134 , \8135 );
xnor \U$7968 ( \8137 , \8136 , \173 );
xor \U$7969 ( \8138 , \8133 , \8137 );
and \U$7970 ( \8139 , \3912 , \438 );
and \U$7971 ( \8140 , \4160 , \336 );
nor \U$7972 ( \8141 , \8139 , \8140 );
xnor \U$7973 ( \8142 , \8141 , \320 );
xor \U$7974 ( \8143 , \8138 , \8142 );
xor \U$7975 ( \8144 , \8129 , \8143 );
and \U$7976 ( \8145 , \6281 , \230 );
and \U$7977 ( \8146 , \6514 , \228 );
nor \U$7978 ( \8147 , \8145 , \8146 );
xnor \U$7979 ( \8148 , \8147 , \237 );
and \U$7980 ( \8149 , \5674 , \245 );
and \U$7981 ( \8150 , \6030 , \243 );
nor \U$7982 ( \8151 , \8149 , \8150 );
xnor \U$7983 ( \8152 , \8151 , \252 );
xor \U$7984 ( \8153 , \8148 , \8152 );
and \U$7985 ( \8154 , \5156 , \141 );
and \U$7986 ( \8155 , \5469 , \139 );
nor \U$7987 ( \8156 , \8154 , \8155 );
xnor \U$7988 ( \8157 , \8156 , \148 );
xor \U$7989 ( \8158 , \8153 , \8157 );
xor \U$7990 ( \8159 , \8144 , \8158 );
xor \U$7991 ( \8160 , \8115 , \8159 );
xor \U$7992 ( \8161 , \8055 , \8160 );
xor \U$7993 ( \8162 , \7973 , \8161 );
xor \U$7994 ( \8163 , \7937 , \8162 );
xor \U$7995 ( \8164 , \7923 , \8163 );
and \U$7996 ( \8165 , \7620 , \7631 );
and \U$7997 ( \8166 , \7631 , \7882 );
and \U$7998 ( \8167 , \7620 , \7882 );
or \U$7999 ( \8168 , \8165 , \8166 , \8167 );
xor \U$8000 ( \8169 , \8164 , \8168 );
and \U$8001 ( \8170 , \7883 , \7887 );
and \U$8002 ( \8171 , \7888 , \7891 );
or \U$8003 ( \8172 , \8170 , \8171 );
xor \U$8004 ( \8173 , \8169 , \8172 );
buf g552d_GF_PartitionCandidate( \8174_nG552d , \8173 );
buf \U$8005 ( \8175 , \8174_nG552d );
and \U$8006 ( \8176 , \7902 , \7906 );
and \U$8007 ( \8177 , \7906 , \7921 );
and \U$8008 ( \8178 , \7902 , \7921 );
or \U$8009 ( \8179 , \8176 , \8177 , \8178 );
and \U$8010 ( \8180 , \7937 , \8162 );
xor \U$8011 ( \8181 , \8179 , \8180 );
and \U$8012 ( \8182 , \7911 , \7915 );
and \U$8013 ( \8183 , \7915 , \7920 );
and \U$8014 ( \8184 , \7911 , \7920 );
or \U$8015 ( \8185 , \8182 , \8183 , \8184 );
and \U$8016 ( \8186 , \7955 , \7956 );
and \U$8017 ( \8187 , \7956 , \7971 );
and \U$8018 ( \8188 , \7955 , \7971 );
or \U$8019 ( \8189 , \8186 , \8187 , \8188 );
xor \U$8020 ( \8190 , \8185 , \8189 );
and \U$8021 ( \8191 , \7987 , \8054 );
and \U$8022 ( \8192 , \8054 , \8160 );
and \U$8023 ( \8193 , \7987 , \8160 );
or \U$8024 ( \8194 , \8191 , \8192 , \8193 );
xor \U$8025 ( \8195 , \8190 , \8194 );
xor \U$8026 ( \8196 , \8181 , \8195 );
and \U$8027 ( \8197 , \7927 , \7931 );
and \U$8028 ( \8198 , \7931 , \7936 );
and \U$8029 ( \8199 , \7927 , \7936 );
or \U$8030 ( \8200 , \8197 , \8198 , \8199 );
and \U$8031 ( \8201 , \7951 , \7972 );
and \U$8032 ( \8202 , \7972 , \8161 );
and \U$8033 ( \8203 , \7951 , \8161 );
or \U$8034 ( \8204 , \8201 , \8202 , \8203 );
xor \U$8035 ( \8205 , \8200 , \8204 );
and \U$8036 ( \8206 , \7977 , \7981 );
and \U$8037 ( \8207 , \7981 , \7986 );
and \U$8038 ( \8208 , \7977 , \7986 );
or \U$8039 ( \8209 , \8206 , \8207 , \8208 );
and \U$8040 ( \8210 , \7941 , \7945 );
and \U$8041 ( \8211 , \7945 , \7950 );
and \U$8042 ( \8212 , \7941 , \7950 );
or \U$8043 ( \8213 , \8210 , \8211 , \8212 );
xor \U$8044 ( \8214 , \8209 , \8213 );
and \U$8045 ( \8215 , \8070 , \8114 );
and \U$8046 ( \8216 , \8114 , \8159 );
and \U$8047 ( \8217 , \8070 , \8159 );
or \U$8048 ( \8218 , \8215 , \8216 , \8217 );
xor \U$8049 ( \8219 , \8214 , \8218 );
and \U$8050 ( \8220 , \8001 , \8015 );
and \U$8051 ( \8221 , \8015 , \8053 );
and \U$8052 ( \8222 , \8001 , \8053 );
or \U$8053 ( \8223 , \8220 , \8221 , \8222 );
and \U$8054 ( \8224 , \8133 , \8137 );
and \U$8055 ( \8225 , \8137 , \8142 );
and \U$8056 ( \8226 , \8133 , \8142 );
or \U$8057 ( \8227 , \8224 , \8225 , \8226 );
and \U$8058 ( \8228 , \8060 , \8064 );
and \U$8059 ( \8229 , \8064 , \8069 );
and \U$8060 ( \8230 , \8060 , \8069 );
or \U$8061 ( \8231 , \8228 , \8229 , \8230 );
xor \U$8062 ( \8232 , \8227 , \8231 );
and \U$8063 ( \8233 , \8148 , \8152 );
and \U$8064 ( \8234 , \8152 , \8157 );
and \U$8065 ( \8235 , \8148 , \8157 );
or \U$8066 ( \8236 , \8233 , \8234 , \8235 );
xor \U$8067 ( \8237 , \8232 , \8236 );
xor \U$8068 ( \8238 , \8223 , \8237 );
and \U$8069 ( \8239 , \8119 , \8123 );
and \U$8070 ( \8240 , \8123 , \8128 );
and \U$8071 ( \8241 , \8119 , \8128 );
or \U$8072 ( \8242 , \8239 , \8240 , \8241 );
and \U$8073 ( \8243 , \8074 , \8078 );
and \U$8074 ( \8244 , \8078 , \8083 );
and \U$8075 ( \8245 , \8074 , \8083 );
or \U$8076 ( \8246 , \8243 , \8244 , \8245 );
xor \U$8077 ( \8247 , \8242 , \8246 );
and \U$8078 ( \8248 , \8088 , \8092 );
and \U$8079 ( \8249 , \8092 , \8097 );
and \U$8080 ( \8250 , \8088 , \8097 );
or \U$8081 ( \8251 , \8248 , \8249 , \8250 );
xor \U$8082 ( \8252 , \8247 , \8251 );
and \U$8083 ( \8253 , \8027 , \8031 );
and \U$8084 ( \8254 , \8031 , \8036 );
and \U$8085 ( \8255 , \8027 , \8036 );
or \U$8086 ( \8256 , \8253 , \8254 , \8255 );
and \U$8087 ( \8257 , \8042 , \8046 );
and \U$8088 ( \8258 , \8046 , \8051 );
and \U$8089 ( \8259 , \8042 , \8051 );
or \U$8090 ( \8260 , \8257 , \8258 , \8259 );
xor \U$8091 ( \8261 , \8256 , \8260 );
and \U$8092 ( \8262 , \8103 , \8107 );
and \U$8093 ( \8263 , \8107 , \8112 );
and \U$8094 ( \8264 , \8103 , \8112 );
or \U$8095 ( \8265 , \8262 , \8263 , \8264 );
xor \U$8096 ( \8266 , \8261 , \8265 );
xor \U$8097 ( \8267 , \8252 , \8266 );
and \U$8098 ( \8268 , \261 , \4581 );
and \U$8099 ( \8269 , \307 , \4424 );
nor \U$8100 ( \8270 , \8268 , \8269 );
xnor \U$8101 ( \8271 , \8270 , \4377 );
and \U$8102 ( \8272 , \178 , \5011 );
and \U$8103 ( \8273 , \185 , \4878 );
nor \U$8104 ( \8274 , \8272 , \8273 );
xnor \U$8105 ( \8275 , \8274 , \4762 );
xor \U$8106 ( \8276 , \8271 , \8275 );
and \U$8107 ( \8277 , \189 , \5485 );
and \U$8108 ( \8278 , \197 , \5275 );
nor \U$8109 ( \8279 , \8277 , \8278 );
xnor \U$8110 ( \8280 , \8279 , \5169 );
xor \U$8111 ( \8281 , \8276 , \8280 );
and \U$8112 ( \8282 , \134 , \7489 );
and \U$8113 ( \8283 , \143 , \7137 );
nor \U$8114 ( \8284 , \8282 , \8283 );
xnor \U$8115 ( \8285 , \8284 , \7142 );
and \U$8116 ( \8286 , \150 , \8019 );
and \U$8117 ( \8287 , \158 , \7830 );
nor \U$8118 ( \8288 , \8286 , \8287 );
xnor \U$8119 ( \8289 , \8288 , \7713 );
xor \U$8120 ( \8290 , \8285 , \8289 );
buf \U$8121 ( \8291 , RIb560c78_8);
xor \U$8122 ( \8292 , \8291 , \7709 );
nand \U$8123 ( \8293 , \166 , \8292 );
buf \U$8124 ( \8294 , RIb560cf0_7);
and \U$8125 ( \8295 , \8291 , \7709 );
not \U$8126 ( \8296 , \8295 );
and \U$8127 ( \8297 , \8294 , \8296 );
xnor \U$8128 ( \8298 , \8293 , \8297 );
xor \U$8129 ( \8299 , \8290 , \8298 );
xor \U$8130 ( \8300 , \8281 , \8299 );
and \U$8131 ( \8301 , \209 , \5996 );
and \U$8132 ( \8302 , \217 , \5695 );
nor \U$8133 ( \8303 , \8301 , \8302 );
xnor \U$8134 ( \8304 , \8303 , \5687 );
and \U$8135 ( \8305 , \224 , \6401 );
and \U$8136 ( \8306 , \232 , \6143 );
nor \U$8137 ( \8307 , \8305 , \8306 );
xnor \U$8138 ( \8308 , \8307 , \6148 );
xor \U$8139 ( \8309 , \8304 , \8308 );
and \U$8140 ( \8310 , \240 , \7055 );
and \U$8141 ( \8311 , \247 , \6675 );
nor \U$8142 ( \8312 , \8310 , \8311 );
xnor \U$8143 ( \8313 , \8312 , \6680 );
xor \U$8144 ( \8314 , \8309 , \8313 );
xor \U$8145 ( \8315 , \8300 , \8314 );
xor \U$8146 ( \8316 , \8267 , \8315 );
xor \U$8147 ( \8317 , \8238 , \8316 );
xor \U$8148 ( \8318 , \8219 , \8317 );
and \U$8149 ( \8319 , \8084 , \8098 );
and \U$8150 ( \8320 , \8098 , \8113 );
and \U$8151 ( \8321 , \8084 , \8113 );
or \U$8152 ( \8322 , \8319 , \8320 , \8321 );
and \U$8153 ( \8323 , \8129 , \8143 );
and \U$8154 ( \8324 , \8143 , \8158 );
and \U$8155 ( \8325 , \8129 , \8158 );
or \U$8156 ( \8326 , \8323 , \8324 , \8325 );
xor \U$8157 ( \8327 , \8322 , \8326 );
and \U$8158 ( \8328 , \8023 , \8037 );
and \U$8159 ( \8329 , \8037 , \8052 );
and \U$8160 ( \8330 , \8023 , \8052 );
or \U$8161 ( \8331 , \8328 , \8329 , \8330 );
xor \U$8162 ( \8332 , \8327 , \8331 );
and \U$8163 ( \8333 , \7961 , \7965 );
and \U$8164 ( \8334 , \7965 , \7970 );
and \U$8165 ( \8335 , \7961 , \7970 );
or \U$8166 ( \8336 , \8333 , \8334 , \8335 );
and \U$8167 ( \8337 , \7991 , \7995 );
and \U$8168 ( \8338 , \7995 , \8000 );
and \U$8169 ( \8339 , \7991 , \8000 );
or \U$8170 ( \8340 , \8337 , \8338 , \8339 );
xor \U$8171 ( \8341 , \8336 , \8340 );
and \U$8172 ( \8342 , \8005 , \8009 );
and \U$8173 ( \8343 , \8009 , \8014 );
and \U$8174 ( \8344 , \8005 , \8014 );
or \U$8175 ( \8345 , \8342 , \8343 , \8344 );
xor \U$8176 ( \8346 , \8341 , \8345 );
xor \U$8177 ( \8347 , \8332 , \8346 );
and \U$8178 ( \8348 , \8057 , \183 );
buf \U$8179 ( \8349 , RIb55ee78_72);
and \U$8180 ( \8350 , \8349 , \180 );
nor \U$8181 ( \8351 , \8348 , \8350 );
xnor \U$8182 ( \8352 , \8351 , \179 );
and \U$8183 ( \8353 , \7556 , \195 );
and \U$8184 ( \8354 , \7700 , \193 );
nor \U$8185 ( \8355 , \8353 , \8354 );
xnor \U$8186 ( \8356 , \8355 , \202 );
xor \U$8187 ( \8357 , \8352 , \8356 );
xor \U$8188 ( \8358 , \8357 , \8297 );
and \U$8189 ( \8359 , \6945 , \215 );
and \U$8190 ( \8360 , \7231 , \213 );
nor \U$8191 ( \8361 , \8359 , \8360 );
xnor \U$8192 ( \8362 , \8361 , \222 );
and \U$8193 ( \8363 , \6514 , \230 );
and \U$8194 ( \8364 , \6790 , \228 );
nor \U$8195 ( \8365 , \8363 , \8364 );
xnor \U$8196 ( \8366 , \8365 , \237 );
xor \U$8197 ( \8367 , \8362 , \8366 );
and \U$8198 ( \8368 , \6030 , \245 );
and \U$8199 ( \8369 , \6281 , \243 );
nor \U$8200 ( \8370 , \8368 , \8369 );
xnor \U$8201 ( \8371 , \8370 , \252 );
xor \U$8202 ( \8372 , \8367 , \8371 );
and \U$8203 ( \8373 , \5469 , \141 );
and \U$8204 ( \8374 , \5674 , \139 );
nor \U$8205 ( \8375 , \8373 , \8374 );
xnor \U$8206 ( \8376 , \8375 , \148 );
and \U$8207 ( \8377 , \4922 , \156 );
and \U$8208 ( \8378 , \5156 , \154 );
nor \U$8209 ( \8379 , \8377 , \8378 );
xnor \U$8210 ( \8380 , \8379 , \163 );
xor \U$8211 ( \8381 , \8376 , \8380 );
and \U$8212 ( \8382 , \4654 , \296 );
and \U$8213 ( \8383 , \4749 , \168 );
nor \U$8214 ( \8384 , \8382 , \8383 );
xnor \U$8215 ( \8385 , \8384 , \173 );
xor \U$8216 ( \8386 , \8381 , \8385 );
xor \U$8217 ( \8387 , \8372 , \8386 );
and \U$8218 ( \8388 , \4160 , \438 );
and \U$8219 ( \8389 , \4364 , \336 );
nor \U$8220 ( \8390 , \8388 , \8389 );
xnor \U$8221 ( \8391 , \8390 , \320 );
and \U$8222 ( \8392 , \3736 , \1086 );
and \U$8223 ( \8393 , \3912 , \508 );
nor \U$8224 ( \8394 , \8392 , \8393 );
xnor \U$8225 ( \8395 , \8394 , \487 );
xor \U$8226 ( \8396 , \8391 , \8395 );
and \U$8227 ( \8397 , \3395 , \1301 );
and \U$8228 ( \8398 , \3646 , \1246 );
nor \U$8229 ( \8399 , \8397 , \8398 );
xnor \U$8230 ( \8400 , \8399 , \1205 );
xor \U$8231 ( \8401 , \8396 , \8400 );
xor \U$8232 ( \8402 , \8387 , \8401 );
xor \U$8233 ( \8403 , \8358 , \8402 );
and \U$8234 ( \8404 , \2090 , \2400 );
and \U$8235 ( \8405 , \2182 , \2246 );
nor \U$8236 ( \8406 , \8404 , \8405 );
xnor \U$8237 ( \8407 , \8406 , \2195 );
and \U$8238 ( \8408 , \1802 , \2669 );
and \U$8239 ( \8409 , \1948 , \2538 );
nor \U$8240 ( \8410 , \8408 , \8409 );
xnor \U$8241 ( \8411 , \8410 , \2534 );
xor \U$8242 ( \8412 , \8407 , \8411 );
and \U$8243 ( \8413 , \1601 , \3103 );
and \U$8244 ( \8414 , \1684 , \2934 );
nor \U$8245 ( \8415 , \8413 , \8414 );
xnor \U$8246 ( \8416 , \8415 , \2839 );
xor \U$8247 ( \8417 , \8412 , \8416 );
and \U$8248 ( \8418 , \3037 , \1578 );
and \U$8249 ( \8419 , \3143 , \1431 );
nor \U$8250 ( \8420 , \8418 , \8419 );
xnor \U$8251 ( \8421 , \8420 , \1436 );
and \U$8252 ( \8422 , \2757 , \1824 );
and \U$8253 ( \8423 , \2826 , \1739 );
nor \U$8254 ( \8424 , \8422 , \8423 );
xnor \U$8255 ( \8425 , \8424 , \1697 );
xor \U$8256 ( \8426 , \8421 , \8425 );
and \U$8257 ( \8427 , \2366 , \2121 );
and \U$8258 ( \8428 , \2521 , \2008 );
nor \U$8259 ( \8429 , \8427 , \8428 );
xnor \U$8260 ( \8430 , \8429 , \1961 );
xor \U$8261 ( \8431 , \8426 , \8430 );
xor \U$8262 ( \8432 , \8417 , \8431 );
and \U$8263 ( \8433 , \1333 , \3357 );
and \U$8264 ( \8434 , \1484 , \3255 );
nor \U$8265 ( \8435 , \8433 , \8434 );
xnor \U$8266 ( \8436 , \8435 , \3156 );
and \U$8267 ( \8437 , \1147 , \3813 );
and \U$8268 ( \8438 , \1192 , \3557 );
nor \U$8269 ( \8439 , \8437 , \8438 );
xnor \U$8270 ( \8440 , \8439 , \3562 );
xor \U$8271 ( \8441 , \8436 , \8440 );
and \U$8272 ( \8442 , \412 , \4132 );
and \U$8273 ( \8443 , \474 , \4012 );
nor \U$8274 ( \8444 , \8442 , \8443 );
xnor \U$8275 ( \8445 , \8444 , \3925 );
xor \U$8276 ( \8446 , \8441 , \8445 );
xor \U$8277 ( \8447 , \8432 , \8446 );
xor \U$8278 ( \8448 , \8403 , \8447 );
xor \U$8279 ( \8449 , \8347 , \8448 );
xor \U$8280 ( \8450 , \8318 , \8449 );
xor \U$8281 ( \8451 , \8205 , \8450 );
xor \U$8282 ( \8452 , \8196 , \8451 );
and \U$8283 ( \8453 , \7898 , \7922 );
and \U$8284 ( \8454 , \7922 , \8163 );
and \U$8285 ( \8455 , \7898 , \8163 );
or \U$8286 ( \8456 , \8453 , \8454 , \8455 );
xor \U$8287 ( \8457 , \8452 , \8456 );
and \U$8288 ( \8458 , \8164 , \8168 );
and \U$8289 ( \8459 , \8169 , \8172 );
or \U$8290 ( \8460 , \8458 , \8459 );
xor \U$8291 ( \8461 , \8457 , \8460 );
buf g552b_GF_PartitionCandidate( \8462_nG552b , \8461 );
buf \U$8292 ( \8463 , \8462_nG552b );
and \U$8293 ( \8464 , \8179 , \8180 );
and \U$8294 ( \8465 , \8180 , \8195 );
and \U$8295 ( \8466 , \8179 , \8195 );
or \U$8296 ( \8467 , \8464 , \8465 , \8466 );
and \U$8297 ( \8468 , \8200 , \8204 );
and \U$8298 ( \8469 , \8204 , \8450 );
and \U$8299 ( \8470 , \8200 , \8450 );
or \U$8300 ( \8471 , \8468 , \8469 , \8470 );
and \U$8301 ( \8472 , \8209 , \8213 );
and \U$8302 ( \8473 , \8213 , \8218 );
and \U$8303 ( \8474 , \8209 , \8218 );
or \U$8304 ( \8475 , \8472 , \8473 , \8474 );
and \U$8305 ( \8476 , \8223 , \8237 );
and \U$8306 ( \8477 , \8237 , \8316 );
and \U$8307 ( \8478 , \8223 , \8316 );
or \U$8308 ( \8479 , \8476 , \8477 , \8478 );
xor \U$8309 ( \8480 , \8475 , \8479 );
and \U$8310 ( \8481 , \8332 , \8346 );
and \U$8311 ( \8482 , \8346 , \8448 );
and \U$8312 ( \8483 , \8332 , \8448 );
or \U$8313 ( \8484 , \8481 , \8482 , \8483 );
xor \U$8314 ( \8485 , \8480 , \8484 );
xor \U$8315 ( \8486 , \8471 , \8485 );
and \U$8316 ( \8487 , \8185 , \8189 );
and \U$8317 ( \8488 , \8189 , \8194 );
and \U$8318 ( \8489 , \8185 , \8194 );
or \U$8319 ( \8490 , \8487 , \8488 , \8489 );
and \U$8320 ( \8491 , \8219 , \8317 );
and \U$8321 ( \8492 , \8317 , \8449 );
and \U$8322 ( \8493 , \8219 , \8449 );
or \U$8323 ( \8494 , \8491 , \8492 , \8493 );
xor \U$8324 ( \8495 , \8490 , \8494 );
and \U$8325 ( \8496 , \8322 , \8326 );
and \U$8326 ( \8497 , \8326 , \8331 );
and \U$8327 ( \8498 , \8322 , \8331 );
or \U$8328 ( \8499 , \8496 , \8497 , \8498 );
and \U$8329 ( \8500 , \8336 , \8340 );
and \U$8330 ( \8501 , \8340 , \8345 );
and \U$8331 ( \8502 , \8336 , \8345 );
or \U$8332 ( \8503 , \8500 , \8501 , \8502 );
xor \U$8333 ( \8504 , \8499 , \8503 );
and \U$8334 ( \8505 , \8358 , \8402 );
and \U$8335 ( \8506 , \8402 , \8447 );
and \U$8336 ( \8507 , \8358 , \8447 );
or \U$8337 ( \8508 , \8505 , \8506 , \8507 );
xor \U$8338 ( \8509 , \8504 , \8508 );
and \U$8339 ( \8510 , \8252 , \8266 );
and \U$8340 ( \8511 , \8266 , \8315 );
and \U$8341 ( \8512 , \8252 , \8315 );
or \U$8342 ( \8513 , \8510 , \8511 , \8512 );
and \U$8343 ( \8514 , \8362 , \8366 );
and \U$8344 ( \8515 , \8366 , \8371 );
and \U$8345 ( \8516 , \8362 , \8371 );
or \U$8346 ( \8517 , \8514 , \8515 , \8516 );
and \U$8347 ( \8518 , \8376 , \8380 );
and \U$8348 ( \8519 , \8380 , \8385 );
and \U$8349 ( \8520 , \8376 , \8385 );
or \U$8350 ( \8521 , \8518 , \8519 , \8520 );
xor \U$8351 ( \8522 , \8517 , \8521 );
and \U$8352 ( \8523 , \8352 , \8356 );
and \U$8353 ( \8524 , \8356 , \8297 );
and \U$8354 ( \8525 , \8352 , \8297 );
or \U$8355 ( \8526 , \8523 , \8524 , \8525 );
xor \U$8356 ( \8527 , \8522 , \8526 );
xor \U$8357 ( \8528 , \8513 , \8527 );
and \U$8358 ( \8529 , \8285 , \8289 );
and \U$8359 ( \8530 , \8289 , \8298 );
and \U$8360 ( \8531 , \8285 , \8298 );
or \U$8361 ( \8532 , \8529 , \8530 , \8531 );
and \U$8362 ( \8533 , \158 , \8019 );
and \U$8363 ( \8534 , \134 , \7830 );
nor \U$8364 ( \8535 , \8533 , \8534 );
xnor \U$8365 ( \8536 , \8535 , \7713 );
xor \U$8366 ( \8537 , \8532 , \8536 );
xor \U$8367 ( \8538 , \8294 , \8291 );
not \U$8368 ( \8539 , \8292 );
and \U$8369 ( \8540 , \8538 , \8539 );
and \U$8370 ( \8541 , \166 , \8540 );
and \U$8371 ( \8542 , \150 , \8292 );
nor \U$8372 ( \8543 , \8541 , \8542 );
xnor \U$8373 ( \8544 , \8543 , \8297 );
xor \U$8374 ( \8545 , \8537 , \8544 );
and \U$8375 ( \8546 , \8407 , \8411 );
and \U$8376 ( \8547 , \8411 , \8416 );
and \U$8377 ( \8548 , \8407 , \8416 );
or \U$8378 ( \8549 , \8546 , \8547 , \8548 );
and \U$8379 ( \8550 , \8391 , \8395 );
and \U$8380 ( \8551 , \8395 , \8400 );
and \U$8381 ( \8552 , \8391 , \8400 );
or \U$8382 ( \8553 , \8550 , \8551 , \8552 );
xor \U$8383 ( \8554 , \8549 , \8553 );
and \U$8384 ( \8555 , \8421 , \8425 );
and \U$8385 ( \8556 , \8425 , \8430 );
and \U$8386 ( \8557 , \8421 , \8430 );
or \U$8387 ( \8558 , \8555 , \8556 , \8557 );
xor \U$8388 ( \8559 , \8554 , \8558 );
xor \U$8389 ( \8560 , \8545 , \8559 );
and \U$8390 ( \8561 , \8271 , \8275 );
and \U$8391 ( \8562 , \8275 , \8280 );
and \U$8392 ( \8563 , \8271 , \8280 );
or \U$8393 ( \8564 , \8561 , \8562 , \8563 );
and \U$8394 ( \8565 , \8304 , \8308 );
and \U$8395 ( \8566 , \8308 , \8313 );
and \U$8396 ( \8567 , \8304 , \8313 );
or \U$8397 ( \8568 , \8565 , \8566 , \8567 );
xor \U$8398 ( \8569 , \8564 , \8568 );
and \U$8399 ( \8570 , \8436 , \8440 );
and \U$8400 ( \8571 , \8440 , \8445 );
and \U$8401 ( \8572 , \8436 , \8445 );
or \U$8402 ( \8573 , \8570 , \8571 , \8572 );
xor \U$8403 ( \8574 , \8569 , \8573 );
xor \U$8404 ( \8575 , \8560 , \8574 );
xor \U$8405 ( \8576 , \8528 , \8575 );
xor \U$8406 ( \8577 , \8509 , \8576 );
and \U$8407 ( \8578 , \8372 , \8386 );
and \U$8408 ( \8579 , \8386 , \8401 );
and \U$8409 ( \8580 , \8372 , \8401 );
or \U$8410 ( \8581 , \8578 , \8579 , \8580 );
and \U$8411 ( \8582 , \8417 , \8431 );
and \U$8412 ( \8583 , \8431 , \8446 );
and \U$8413 ( \8584 , \8417 , \8446 );
or \U$8414 ( \8585 , \8582 , \8583 , \8584 );
xor \U$8415 ( \8586 , \8581 , \8585 );
and \U$8416 ( \8587 , \8281 , \8299 );
and \U$8417 ( \8588 , \8299 , \8314 );
and \U$8418 ( \8589 , \8281 , \8314 );
or \U$8419 ( \8590 , \8587 , \8588 , \8589 );
xor \U$8420 ( \8591 , \8586 , \8590 );
and \U$8421 ( \8592 , \8242 , \8246 );
and \U$8422 ( \8593 , \8246 , \8251 );
and \U$8423 ( \8594 , \8242 , \8251 );
or \U$8424 ( \8595 , \8592 , \8593 , \8594 );
and \U$8425 ( \8596 , \8256 , \8260 );
and \U$8426 ( \8597 , \8260 , \8265 );
and \U$8427 ( \8598 , \8256 , \8265 );
or \U$8428 ( \8599 , \8596 , \8597 , \8598 );
xor \U$8429 ( \8600 , \8595 , \8599 );
and \U$8430 ( \8601 , \8227 , \8231 );
and \U$8431 ( \8602 , \8231 , \8236 );
and \U$8432 ( \8603 , \8227 , \8236 );
or \U$8433 ( \8604 , \8601 , \8602 , \8603 );
xor \U$8434 ( \8605 , \8600 , \8604 );
xor \U$8435 ( \8606 , \8591 , \8605 );
and \U$8436 ( \8607 , \185 , \5011 );
and \U$8437 ( \8608 , \261 , \4878 );
nor \U$8438 ( \8609 , \8607 , \8608 );
xnor \U$8439 ( \8610 , \8609 , \4762 );
and \U$8440 ( \8611 , \197 , \5485 );
and \U$8441 ( \8612 , \178 , \5275 );
nor \U$8442 ( \8613 , \8611 , \8612 );
xnor \U$8443 ( \8614 , \8613 , \5169 );
xor \U$8444 ( \8615 , \8610 , \8614 );
and \U$8445 ( \8616 , \217 , \5996 );
and \U$8446 ( \8617 , \189 , \5695 );
nor \U$8447 ( \8618 , \8616 , \8617 );
xnor \U$8448 ( \8619 , \8618 , \5687 );
xor \U$8449 ( \8620 , \8615 , \8619 );
and \U$8450 ( \8621 , \232 , \6401 );
and \U$8451 ( \8622 , \209 , \6143 );
nor \U$8452 ( \8623 , \8621 , \8622 );
xnor \U$8453 ( \8624 , \8623 , \6148 );
and \U$8454 ( \8625 , \247 , \7055 );
and \U$8455 ( \8626 , \224 , \6675 );
nor \U$8456 ( \8627 , \8625 , \8626 );
xnor \U$8457 ( \8628 , \8627 , \6680 );
xor \U$8458 ( \8629 , \8624 , \8628 );
and \U$8459 ( \8630 , \143 , \7489 );
and \U$8460 ( \8631 , \240 , \7137 );
nor \U$8461 ( \8632 , \8630 , \8631 );
xnor \U$8462 ( \8633 , \8632 , \7142 );
xor \U$8463 ( \8634 , \8629 , \8633 );
xor \U$8464 ( \8635 , \8620 , \8634 );
and \U$8465 ( \8636 , \1192 , \3813 );
and \U$8466 ( \8637 , \1333 , \3557 );
nor \U$8467 ( \8638 , \8636 , \8637 );
xnor \U$8468 ( \8639 , \8638 , \3562 );
and \U$8469 ( \8640 , \474 , \4132 );
and \U$8470 ( \8641 , \1147 , \4012 );
nor \U$8471 ( \8642 , \8640 , \8641 );
xnor \U$8472 ( \8643 , \8642 , \3925 );
xor \U$8473 ( \8644 , \8639 , \8643 );
and \U$8474 ( \8645 , \307 , \4581 );
and \U$8475 ( \8646 , \412 , \4424 );
nor \U$8476 ( \8647 , \8645 , \8646 );
xnor \U$8477 ( \8648 , \8647 , \4377 );
xor \U$8478 ( \8649 , \8644 , \8648 );
xor \U$8479 ( \8650 , \8635 , \8649 );
and \U$8480 ( \8651 , \8349 , \183 );
buf \U$8481 ( \8652 , RIb55eef0_71);
and \U$8482 ( \8653 , \8652 , \180 );
nor \U$8483 ( \8654 , \8651 , \8653 );
xnor \U$8484 ( \8655 , \8654 , \179 );
and \U$8485 ( \8656 , \7700 , \195 );
and \U$8486 ( \8657 , \8057 , \193 );
nor \U$8487 ( \8658 , \8656 , \8657 );
xnor \U$8488 ( \8659 , \8658 , \202 );
xor \U$8489 ( \8660 , \8655 , \8659 );
and \U$8490 ( \8661 , \7231 , \215 );
and \U$8491 ( \8662 , \7556 , \213 );
nor \U$8492 ( \8663 , \8661 , \8662 );
xnor \U$8493 ( \8664 , \8663 , \222 );
xor \U$8494 ( \8665 , \8660 , \8664 );
and \U$8495 ( \8666 , \6790 , \230 );
and \U$8496 ( \8667 , \6945 , \228 );
nor \U$8497 ( \8668 , \8666 , \8667 );
xnor \U$8498 ( \8669 , \8668 , \237 );
and \U$8499 ( \8670 , \6281 , \245 );
and \U$8500 ( \8671 , \6514 , \243 );
nor \U$8501 ( \8672 , \8670 , \8671 );
xnor \U$8502 ( \8673 , \8672 , \252 );
xor \U$8503 ( \8674 , \8669 , \8673 );
and \U$8504 ( \8675 , \5674 , \141 );
and \U$8505 ( \8676 , \6030 , \139 );
nor \U$8506 ( \8677 , \8675 , \8676 );
xnor \U$8507 ( \8678 , \8677 , \148 );
xor \U$8508 ( \8679 , \8674 , \8678 );
xor \U$8509 ( \8680 , \8665 , \8679 );
and \U$8510 ( \8681 , \5156 , \156 );
and \U$8511 ( \8682 , \5469 , \154 );
nor \U$8512 ( \8683 , \8681 , \8682 );
xnor \U$8513 ( \8684 , \8683 , \163 );
and \U$8514 ( \8685 , \4749 , \296 );
and \U$8515 ( \8686 , \4922 , \168 );
nor \U$8516 ( \8687 , \8685 , \8686 );
xnor \U$8517 ( \8688 , \8687 , \173 );
xor \U$8518 ( \8689 , \8684 , \8688 );
and \U$8519 ( \8690 , \4364 , \438 );
and \U$8520 ( \8691 , \4654 , \336 );
nor \U$8521 ( \8692 , \8690 , \8691 );
xnor \U$8522 ( \8693 , \8692 , \320 );
xor \U$8523 ( \8694 , \8689 , \8693 );
xor \U$8524 ( \8695 , \8680 , \8694 );
xor \U$8525 ( \8696 , \8650 , \8695 );
and \U$8526 ( \8697 , \2826 , \1824 );
and \U$8527 ( \8698 , \3037 , \1739 );
nor \U$8528 ( \8699 , \8697 , \8698 );
xnor \U$8529 ( \8700 , \8699 , \1697 );
and \U$8530 ( \8701 , \2521 , \2121 );
and \U$8531 ( \8702 , \2757 , \2008 );
nor \U$8532 ( \8703 , \8701 , \8702 );
xnor \U$8533 ( \8704 , \8703 , \1961 );
xor \U$8534 ( \8705 , \8700 , \8704 );
and \U$8535 ( \8706 , \2182 , \2400 );
and \U$8536 ( \8707 , \2366 , \2246 );
nor \U$8537 ( \8708 , \8706 , \8707 );
xnor \U$8538 ( \8709 , \8708 , \2195 );
xor \U$8539 ( \8710 , \8705 , \8709 );
and \U$8540 ( \8711 , \1948 , \2669 );
and \U$8541 ( \8712 , \2090 , \2538 );
nor \U$8542 ( \8713 , \8711 , \8712 );
xnor \U$8543 ( \8714 , \8713 , \2534 );
and \U$8544 ( \8715 , \1684 , \3103 );
and \U$8545 ( \8716 , \1802 , \2934 );
nor \U$8546 ( \8717 , \8715 , \8716 );
xnor \U$8547 ( \8718 , \8717 , \2839 );
xor \U$8548 ( \8719 , \8714 , \8718 );
and \U$8549 ( \8720 , \1484 , \3357 );
and \U$8550 ( \8721 , \1601 , \3255 );
nor \U$8551 ( \8722 , \8720 , \8721 );
xnor \U$8552 ( \8723 , \8722 , \3156 );
xor \U$8553 ( \8724 , \8719 , \8723 );
xor \U$8554 ( \8725 , \8710 , \8724 );
and \U$8555 ( \8726 , \3912 , \1086 );
and \U$8556 ( \8727 , \4160 , \508 );
nor \U$8557 ( \8728 , \8726 , \8727 );
xnor \U$8558 ( \8729 , \8728 , \487 );
and \U$8559 ( \8730 , \3646 , \1301 );
and \U$8560 ( \8731 , \3736 , \1246 );
nor \U$8561 ( \8732 , \8730 , \8731 );
xnor \U$8562 ( \8733 , \8732 , \1205 );
xor \U$8563 ( \8734 , \8729 , \8733 );
and \U$8564 ( \8735 , \3143 , \1578 );
and \U$8565 ( \8736 , \3395 , \1431 );
nor \U$8566 ( \8737 , \8735 , \8736 );
xnor \U$8567 ( \8738 , \8737 , \1436 );
xor \U$8568 ( \8739 , \8734 , \8738 );
xor \U$8569 ( \8740 , \8725 , \8739 );
xor \U$8570 ( \8741 , \8696 , \8740 );
xor \U$8571 ( \8742 , \8606 , \8741 );
xor \U$8572 ( \8743 , \8577 , \8742 );
xor \U$8573 ( \8744 , \8495 , \8743 );
xor \U$8574 ( \8745 , \8486 , \8744 );
xor \U$8575 ( \8746 , \8467 , \8745 );
and \U$8576 ( \8747 , \8196 , \8451 );
xor \U$8577 ( \8748 , \8746 , \8747 );
and \U$8578 ( \8749 , \8452 , \8456 );
and \U$8579 ( \8750 , \8457 , \8460 );
or \U$8580 ( \8751 , \8749 , \8750 );
xor \U$8581 ( \8752 , \8748 , \8751 );
buf g5529_GF_PartitionCandidate( \8753_nG5529 , \8752 );
buf \U$8582 ( \8754 , \8753_nG5529 );
and \U$8583 ( \8755 , \8471 , \8485 );
and \U$8584 ( \8756 , \8485 , \8744 );
and \U$8585 ( \8757 , \8471 , \8744 );
or \U$8586 ( \8758 , \8755 , \8756 , \8757 );
and \U$8587 ( \8759 , \8490 , \8494 );
and \U$8588 ( \8760 , \8494 , \8743 );
and \U$8589 ( \8761 , \8490 , \8743 );
or \U$8590 ( \8762 , \8759 , \8760 , \8761 );
and \U$8591 ( \8763 , \8499 , \8503 );
and \U$8592 ( \8764 , \8503 , \8508 );
and \U$8593 ( \8765 , \8499 , \8508 );
or \U$8594 ( \8766 , \8763 , \8764 , \8765 );
and \U$8595 ( \8767 , \8513 , \8527 );
and \U$8596 ( \8768 , \8527 , \8575 );
and \U$8597 ( \8769 , \8513 , \8575 );
or \U$8598 ( \8770 , \8767 , \8768 , \8769 );
xor \U$8599 ( \8771 , \8766 , \8770 );
and \U$8600 ( \8772 , \8591 , \8605 );
and \U$8601 ( \8773 , \8605 , \8741 );
and \U$8602 ( \8774 , \8591 , \8741 );
or \U$8603 ( \8775 , \8772 , \8773 , \8774 );
xor \U$8604 ( \8776 , \8771 , \8775 );
xor \U$8605 ( \8777 , \8762 , \8776 );
and \U$8606 ( \8778 , \8475 , \8479 );
and \U$8607 ( \8779 , \8479 , \8484 );
and \U$8608 ( \8780 , \8475 , \8484 );
or \U$8609 ( \8781 , \8778 , \8779 , \8780 );
and \U$8610 ( \8782 , \8509 , \8576 );
and \U$8611 ( \8783 , \8576 , \8742 );
and \U$8612 ( \8784 , \8509 , \8742 );
or \U$8613 ( \8785 , \8782 , \8783 , \8784 );
xor \U$8614 ( \8786 , \8781 , \8785 );
and \U$8615 ( \8787 , \8581 , \8585 );
and \U$8616 ( \8788 , \8585 , \8590 );
and \U$8617 ( \8789 , \8581 , \8590 );
or \U$8618 ( \8790 , \8787 , \8788 , \8789 );
and \U$8619 ( \8791 , \8595 , \8599 );
and \U$8620 ( \8792 , \8599 , \8604 );
and \U$8621 ( \8793 , \8595 , \8604 );
or \U$8622 ( \8794 , \8791 , \8792 , \8793 );
xor \U$8623 ( \8795 , \8790 , \8794 );
and \U$8624 ( \8796 , \8650 , \8695 );
and \U$8625 ( \8797 , \8695 , \8740 );
and \U$8626 ( \8798 , \8650 , \8740 );
or \U$8627 ( \8799 , \8796 , \8797 , \8798 );
xor \U$8628 ( \8800 , \8795 , \8799 );
and \U$8629 ( \8801 , \8532 , \8536 );
and \U$8630 ( \8802 , \8536 , \8544 );
and \U$8631 ( \8803 , \8532 , \8544 );
or \U$8632 ( \8804 , \8801 , \8802 , \8803 );
and \U$8633 ( \8805 , \8620 , \8634 );
and \U$8634 ( \8806 , \8634 , \8649 );
and \U$8635 ( \8807 , \8620 , \8649 );
or \U$8636 ( \8808 , \8805 , \8806 , \8807 );
xor \U$8637 ( \8809 , \8804 , \8808 );
and \U$8638 ( \8810 , \8710 , \8724 );
and \U$8639 ( \8811 , \8724 , \8739 );
and \U$8640 ( \8812 , \8710 , \8739 );
or \U$8641 ( \8813 , \8810 , \8811 , \8812 );
xor \U$8642 ( \8814 , \8809 , \8813 );
and \U$8643 ( \8815 , \8517 , \8521 );
and \U$8644 ( \8816 , \8521 , \8526 );
and \U$8645 ( \8817 , \8517 , \8526 );
or \U$8646 ( \8818 , \8815 , \8816 , \8817 );
and \U$8647 ( \8819 , \8549 , \8553 );
and \U$8648 ( \8820 , \8553 , \8558 );
and \U$8649 ( \8821 , \8549 , \8558 );
or \U$8650 ( \8822 , \8819 , \8820 , \8821 );
xor \U$8651 ( \8823 , \8818 , \8822 );
and \U$8652 ( \8824 , \8564 , \8568 );
and \U$8653 ( \8825 , \8568 , \8573 );
and \U$8654 ( \8826 , \8564 , \8573 );
or \U$8655 ( \8827 , \8824 , \8825 , \8826 );
xor \U$8656 ( \8828 , \8823 , \8827 );
xor \U$8657 ( \8829 , \8814 , \8828 );
and \U$8658 ( \8830 , \8665 , \8679 );
and \U$8659 ( \8831 , \8679 , \8694 );
and \U$8660 ( \8832 , \8665 , \8694 );
or \U$8661 ( \8833 , \8830 , \8831 , \8832 );
and \U$8662 ( \8834 , \8652 , \183 );
buf \U$8663 ( \8835 , RIb55ef68_70);
and \U$8664 ( \8836 , \8835 , \180 );
nor \U$8665 ( \8837 , \8834 , \8836 );
xnor \U$8666 ( \8838 , \8837 , \179 );
and \U$8667 ( \8839 , \8057 , \195 );
and \U$8668 ( \8840 , \8349 , \193 );
nor \U$8669 ( \8841 , \8839 , \8840 );
xnor \U$8670 ( \8842 , \8841 , \202 );
xor \U$8671 ( \8843 , \8838 , \8842 );
buf \U$8672 ( \8844 , RIb560de0_5);
buf \U$8673 ( \8845 , RIb560d68_6);
and \U$8674 ( \8846 , \8845 , \8294 );
not \U$8675 ( \8847 , \8846 );
and \U$8676 ( \8848 , \8844 , \8847 );
xor \U$8677 ( \8849 , \8843 , \8848 );
xor \U$8678 ( \8850 , \8833 , \8849 );
and \U$8679 ( \8851 , \7556 , \215 );
and \U$8680 ( \8852 , \7700 , \213 );
nor \U$8681 ( \8853 , \8851 , \8852 );
xnor \U$8682 ( \8854 , \8853 , \222 );
and \U$8683 ( \8855 , \6945 , \230 );
and \U$8684 ( \8856 , \7231 , \228 );
nor \U$8685 ( \8857 , \8855 , \8856 );
xnor \U$8686 ( \8858 , \8857 , \237 );
xor \U$8687 ( \8859 , \8854 , \8858 );
and \U$8688 ( \8860 , \6514 , \245 );
and \U$8689 ( \8861 , \6790 , \243 );
nor \U$8690 ( \8862 , \8860 , \8861 );
xnor \U$8691 ( \8863 , \8862 , \252 );
xor \U$8692 ( \8864 , \8859 , \8863 );
xor \U$8693 ( \8865 , \8850 , \8864 );
xor \U$8694 ( \8866 , \8829 , \8865 );
xor \U$8695 ( \8867 , \8800 , \8866 );
and \U$8696 ( \8868 , \8545 , \8559 );
and \U$8697 ( \8869 , \8559 , \8574 );
and \U$8698 ( \8870 , \8545 , \8574 );
or \U$8699 ( \8871 , \8868 , \8869 , \8870 );
and \U$8700 ( \8872 , \8700 , \8704 );
and \U$8701 ( \8873 , \8704 , \8709 );
and \U$8702 ( \8874 , \8700 , \8709 );
or \U$8703 ( \8875 , \8872 , \8873 , \8874 );
and \U$8704 ( \8876 , \8714 , \8718 );
and \U$8705 ( \8877 , \8718 , \8723 );
and \U$8706 ( \8878 , \8714 , \8723 );
or \U$8707 ( \8879 , \8876 , \8877 , \8878 );
xor \U$8708 ( \8880 , \8875 , \8879 );
and \U$8709 ( \8881 , \8729 , \8733 );
and \U$8710 ( \8882 , \8733 , \8738 );
and \U$8711 ( \8883 , \8729 , \8738 );
or \U$8712 ( \8884 , \8881 , \8882 , \8883 );
xor \U$8713 ( \8885 , \8880 , \8884 );
and \U$8714 ( \8886 , \8610 , \8614 );
and \U$8715 ( \8887 , \8614 , \8619 );
and \U$8716 ( \8888 , \8610 , \8619 );
or \U$8717 ( \8889 , \8886 , \8887 , \8888 );
and \U$8718 ( \8890 , \8624 , \8628 );
and \U$8719 ( \8891 , \8628 , \8633 );
and \U$8720 ( \8892 , \8624 , \8633 );
or \U$8721 ( \8893 , \8890 , \8891 , \8892 );
xor \U$8722 ( \8894 , \8889 , \8893 );
and \U$8723 ( \8895 , \8639 , \8643 );
and \U$8724 ( \8896 , \8643 , \8648 );
and \U$8725 ( \8897 , \8639 , \8648 );
or \U$8726 ( \8898 , \8895 , \8896 , \8897 );
xor \U$8727 ( \8899 , \8894 , \8898 );
xor \U$8728 ( \8900 , \8885 , \8899 );
and \U$8729 ( \8901 , \8655 , \8659 );
and \U$8730 ( \8902 , \8659 , \8664 );
and \U$8731 ( \8903 , \8655 , \8664 );
or \U$8732 ( \8904 , \8901 , \8902 , \8903 );
and \U$8733 ( \8905 , \8669 , \8673 );
and \U$8734 ( \8906 , \8673 , \8678 );
and \U$8735 ( \8907 , \8669 , \8678 );
or \U$8736 ( \8908 , \8905 , \8906 , \8907 );
xor \U$8737 ( \8909 , \8904 , \8908 );
and \U$8738 ( \8910 , \8684 , \8688 );
and \U$8739 ( \8911 , \8688 , \8693 );
and \U$8740 ( \8912 , \8684 , \8693 );
or \U$8741 ( \8913 , \8910 , \8911 , \8912 );
xor \U$8742 ( \8914 , \8909 , \8913 );
xor \U$8743 ( \8915 , \8900 , \8914 );
xor \U$8744 ( \8916 , \8871 , \8915 );
and \U$8745 ( \8917 , \6030 , \141 );
and \U$8746 ( \8918 , \6281 , \139 );
nor \U$8747 ( \8919 , \8917 , \8918 );
xnor \U$8748 ( \8920 , \8919 , \148 );
and \U$8749 ( \8921 , \5469 , \156 );
and \U$8750 ( \8922 , \5674 , \154 );
nor \U$8751 ( \8923 , \8921 , \8922 );
xnor \U$8752 ( \8924 , \8923 , \163 );
xor \U$8753 ( \8925 , \8920 , \8924 );
and \U$8754 ( \8926 , \4922 , \296 );
and \U$8755 ( \8927 , \5156 , \168 );
nor \U$8756 ( \8928 , \8926 , \8927 );
xnor \U$8757 ( \8929 , \8928 , \173 );
xor \U$8758 ( \8930 , \8925 , \8929 );
and \U$8759 ( \8931 , \3395 , \1578 );
and \U$8760 ( \8932 , \3646 , \1431 );
nor \U$8761 ( \8933 , \8931 , \8932 );
xnor \U$8762 ( \8934 , \8933 , \1436 );
and \U$8763 ( \8935 , \3037 , \1824 );
and \U$8764 ( \8936 , \3143 , \1739 );
nor \U$8765 ( \8937 , \8935 , \8936 );
xnor \U$8766 ( \8938 , \8937 , \1697 );
xor \U$8767 ( \8939 , \8934 , \8938 );
and \U$8768 ( \8940 , \2757 , \2121 );
and \U$8769 ( \8941 , \2826 , \2008 );
nor \U$8770 ( \8942 , \8940 , \8941 );
xnor \U$8771 ( \8943 , \8942 , \1961 );
xor \U$8772 ( \8944 , \8939 , \8943 );
xor \U$8773 ( \8945 , \8930 , \8944 );
and \U$8774 ( \8946 , \4654 , \438 );
and \U$8775 ( \8947 , \4749 , \336 );
nor \U$8776 ( \8948 , \8946 , \8947 );
xnor \U$8777 ( \8949 , \8948 , \320 );
and \U$8778 ( \8950 , \4160 , \1086 );
and \U$8779 ( \8951 , \4364 , \508 );
nor \U$8780 ( \8952 , \8950 , \8951 );
xnor \U$8781 ( \8953 , \8952 , \487 );
xor \U$8782 ( \8954 , \8949 , \8953 );
and \U$8783 ( \8955 , \3736 , \1301 );
and \U$8784 ( \8956 , \3912 , \1246 );
nor \U$8785 ( \8957 , \8955 , \8956 );
xnor \U$8786 ( \8958 , \8957 , \1205 );
xor \U$8787 ( \8959 , \8954 , \8958 );
xor \U$8788 ( \8960 , \8945 , \8959 );
and \U$8789 ( \8961 , \2366 , \2400 );
and \U$8790 ( \8962 , \2521 , \2246 );
nor \U$8791 ( \8963 , \8961 , \8962 );
xnor \U$8792 ( \8964 , \8963 , \2195 );
and \U$8793 ( \8965 , \2090 , \2669 );
and \U$8794 ( \8966 , \2182 , \2538 );
nor \U$8795 ( \8967 , \8965 , \8966 );
xnor \U$8796 ( \8968 , \8967 , \2534 );
xor \U$8797 ( \8969 , \8964 , \8968 );
and \U$8798 ( \8970 , \1802 , \3103 );
and \U$8799 ( \8971 , \1948 , \2934 );
nor \U$8800 ( \8972 , \8970 , \8971 );
xnor \U$8801 ( \8973 , \8972 , \2839 );
xor \U$8802 ( \8974 , \8969 , \8973 );
and \U$8803 ( \8975 , \1601 , \3357 );
and \U$8804 ( \8976 , \1684 , \3255 );
nor \U$8805 ( \8977 , \8975 , \8976 );
xnor \U$8806 ( \8978 , \8977 , \3156 );
and \U$8807 ( \8979 , \1333 , \3813 );
and \U$8808 ( \8980 , \1484 , \3557 );
nor \U$8809 ( \8981 , \8979 , \8980 );
xnor \U$8810 ( \8982 , \8981 , \3562 );
xor \U$8811 ( \8983 , \8978 , \8982 );
and \U$8812 ( \8984 , \1147 , \4132 );
and \U$8813 ( \8985 , \1192 , \4012 );
nor \U$8814 ( \8986 , \8984 , \8985 );
xnor \U$8815 ( \8987 , \8986 , \3925 );
xor \U$8816 ( \8988 , \8983 , \8987 );
xor \U$8817 ( \8989 , \8974 , \8988 );
and \U$8818 ( \8990 , \412 , \4581 );
and \U$8819 ( \8991 , \474 , \4424 );
nor \U$8820 ( \8992 , \8990 , \8991 );
xnor \U$8821 ( \8993 , \8992 , \4377 );
and \U$8822 ( \8994 , \261 , \5011 );
and \U$8823 ( \8995 , \307 , \4878 );
nor \U$8824 ( \8996 , \8994 , \8995 );
xnor \U$8825 ( \8997 , \8996 , \4762 );
xor \U$8826 ( \8998 , \8993 , \8997 );
and \U$8827 ( \8999 , \178 , \5485 );
and \U$8828 ( \9000 , \185 , \5275 );
nor \U$8829 ( \9001 , \8999 , \9000 );
xnor \U$8830 ( \9002 , \9001 , \5169 );
xor \U$8831 ( \9003 , \8998 , \9002 );
xor \U$8832 ( \9004 , \8989 , \9003 );
xor \U$8833 ( \9005 , \8960 , \9004 );
xor \U$8834 ( \9006 , \8845 , \8294 );
nand \U$8835 ( \9007 , \166 , \9006 );
xnor \U$8836 ( \9008 , \9007 , \8848 );
and \U$8837 ( \9009 , \189 , \5996 );
and \U$8838 ( \9010 , \197 , \5695 );
nor \U$8839 ( \9011 , \9009 , \9010 );
xnor \U$8840 ( \9012 , \9011 , \5687 );
and \U$8841 ( \9013 , \209 , \6401 );
and \U$8842 ( \9014 , \217 , \6143 );
nor \U$8843 ( \9015 , \9013 , \9014 );
xnor \U$8844 ( \9016 , \9015 , \6148 );
xor \U$8845 ( \9017 , \9012 , \9016 );
and \U$8846 ( \9018 , \224 , \7055 );
and \U$8847 ( \9019 , \232 , \6675 );
nor \U$8848 ( \9020 , \9018 , \9019 );
xnor \U$8849 ( \9021 , \9020 , \6680 );
xor \U$8850 ( \9022 , \9017 , \9021 );
xor \U$8851 ( \9023 , \9008 , \9022 );
and \U$8852 ( \9024 , \240 , \7489 );
and \U$8853 ( \9025 , \247 , \7137 );
nor \U$8854 ( \9026 , \9024 , \9025 );
xnor \U$8855 ( \9027 , \9026 , \7142 );
and \U$8856 ( \9028 , \134 , \8019 );
and \U$8857 ( \9029 , \143 , \7830 );
nor \U$8858 ( \9030 , \9028 , \9029 );
xnor \U$8859 ( \9031 , \9030 , \7713 );
xor \U$8860 ( \9032 , \9027 , \9031 );
and \U$8861 ( \9033 , \150 , \8540 );
and \U$8862 ( \9034 , \158 , \8292 );
nor \U$8863 ( \9035 , \9033 , \9034 );
xnor \U$8864 ( \9036 , \9035 , \8297 );
xor \U$8865 ( \9037 , \9032 , \9036 );
xor \U$8866 ( \9038 , \9023 , \9037 );
xor \U$8867 ( \9039 , \9005 , \9038 );
xor \U$8868 ( \9040 , \8916 , \9039 );
xor \U$8869 ( \9041 , \8867 , \9040 );
xor \U$8870 ( \9042 , \8786 , \9041 );
xor \U$8871 ( \9043 , \8777 , \9042 );
xor \U$8872 ( \9044 , \8758 , \9043 );
and \U$8873 ( \9045 , \8467 , \8745 );
xor \U$8874 ( \9046 , \9044 , \9045 );
and \U$8875 ( \9047 , \8746 , \8747 );
and \U$8876 ( \9048 , \8748 , \8751 );
or \U$8877 ( \9049 , \9047 , \9048 );
xor \U$8878 ( \9050 , \9046 , \9049 );
buf g5527_GF_PartitionCandidate( \9051_nG5527 , \9050 );
buf \U$8879 ( \9052 , \9051_nG5527 );
and \U$8880 ( \9053 , \8762 , \8776 );
and \U$8881 ( \9054 , \8776 , \9042 );
and \U$8882 ( \9055 , \8762 , \9042 );
or \U$8883 ( \9056 , \9053 , \9054 , \9055 );
and \U$8884 ( \9057 , \8781 , \8785 );
and \U$8885 ( \9058 , \8785 , \9041 );
and \U$8886 ( \9059 , \8781 , \9041 );
or \U$8887 ( \9060 , \9057 , \9058 , \9059 );
and \U$8888 ( \9061 , \8766 , \8770 );
and \U$8889 ( \9062 , \8770 , \8775 );
and \U$8890 ( \9063 , \8766 , \8775 );
or \U$8891 ( \9064 , \9061 , \9062 , \9063 );
and \U$8892 ( \9065 , \8800 , \8866 );
and \U$8893 ( \9066 , \8866 , \9040 );
and \U$8894 ( \9067 , \8800 , \9040 );
or \U$8895 ( \9068 , \9065 , \9066 , \9067 );
xor \U$8896 ( \9069 , \9064 , \9068 );
and \U$8897 ( \9070 , \8885 , \8899 );
and \U$8898 ( \9071 , \8899 , \8914 );
and \U$8899 ( \9072 , \8885 , \8914 );
or \U$8900 ( \9073 , \9070 , \9071 , \9072 );
and \U$8901 ( \9074 , \8960 , \9004 );
and \U$8902 ( \9075 , \9004 , \9038 );
and \U$8903 ( \9076 , \8960 , \9038 );
or \U$8904 ( \9077 , \9074 , \9075 , \9076 );
xor \U$8905 ( \9078 , \9073 , \9077 );
and \U$8906 ( \9079 , \8964 , \8968 );
and \U$8907 ( \9080 , \8968 , \8973 );
and \U$8908 ( \9081 , \8964 , \8973 );
or \U$8909 ( \9082 , \9079 , \9080 , \9081 );
and \U$8910 ( \9083 , \8934 , \8938 );
and \U$8911 ( \9084 , \8938 , \8943 );
and \U$8912 ( \9085 , \8934 , \8943 );
or \U$8913 ( \9086 , \9083 , \9084 , \9085 );
xor \U$8914 ( \9087 , \9082 , \9086 );
and \U$8915 ( \9088 , \8949 , \8953 );
and \U$8916 ( \9089 , \8953 , \8958 );
and \U$8917 ( \9090 , \8949 , \8958 );
or \U$8918 ( \9091 , \9088 , \9089 , \9090 );
xor \U$8919 ( \9092 , \9087 , \9091 );
xor \U$8920 ( \9093 , \9078 , \9092 );
xor \U$8921 ( \9094 , \9069 , \9093 );
xor \U$8922 ( \9095 , \9060 , \9094 );
and \U$8923 ( \9096 , \8804 , \8808 );
and \U$8924 ( \9097 , \8808 , \8813 );
and \U$8925 ( \9098 , \8804 , \8813 );
or \U$8926 ( \9099 , \9096 , \9097 , \9098 );
and \U$8927 ( \9100 , \8818 , \8822 );
and \U$8928 ( \9101 , \8822 , \8827 );
and \U$8929 ( \9102 , \8818 , \8827 );
or \U$8930 ( \9103 , \9100 , \9101 , \9102 );
xor \U$8931 ( \9104 , \9099 , \9103 );
and \U$8932 ( \9105 , \8833 , \8849 );
and \U$8933 ( \9106 , \8849 , \8864 );
and \U$8934 ( \9107 , \8833 , \8864 );
or \U$8935 ( \9108 , \9105 , \9106 , \9107 );
xor \U$8936 ( \9109 , \9104 , \9108 );
and \U$8937 ( \9110 , \8790 , \8794 );
and \U$8938 ( \9111 , \8794 , \8799 );
and \U$8939 ( \9112 , \8790 , \8799 );
or \U$8940 ( \9113 , \9110 , \9111 , \9112 );
and \U$8941 ( \9114 , \8814 , \8828 );
and \U$8942 ( \9115 , \8828 , \8865 );
and \U$8943 ( \9116 , \8814 , \8865 );
or \U$8944 ( \9117 , \9114 , \9115 , \9116 );
xor \U$8945 ( \9118 , \9113 , \9117 );
and \U$8946 ( \9119 , \8871 , \8915 );
and \U$8947 ( \9120 , \8915 , \9039 );
and \U$8948 ( \9121 , \8871 , \9039 );
or \U$8949 ( \9122 , \9119 , \9120 , \9121 );
xor \U$8950 ( \9123 , \9118 , \9122 );
xor \U$8951 ( \9124 , \9109 , \9123 );
and \U$8952 ( \9125 , \8875 , \8879 );
and \U$8953 ( \9126 , \8879 , \8884 );
and \U$8954 ( \9127 , \8875 , \8884 );
or \U$8955 ( \9128 , \9125 , \9126 , \9127 );
and \U$8956 ( \9129 , \8889 , \8893 );
and \U$8957 ( \9130 , \8893 , \8898 );
and \U$8958 ( \9131 , \8889 , \8898 );
or \U$8959 ( \9132 , \9129 , \9130 , \9131 );
xor \U$8960 ( \9133 , \9128 , \9132 );
and \U$8961 ( \9134 , \8904 , \8908 );
and \U$8962 ( \9135 , \8908 , \8913 );
and \U$8963 ( \9136 , \8904 , \8913 );
or \U$8964 ( \9137 , \9134 , \9135 , \9136 );
xor \U$8965 ( \9138 , \9133 , \9137 );
and \U$8966 ( \9139 , \8930 , \8944 );
and \U$8967 ( \9140 , \8944 , \8959 );
and \U$8968 ( \9141 , \8930 , \8959 );
or \U$8969 ( \9142 , \9139 , \9140 , \9141 );
and \U$8970 ( \9143 , \8974 , \8988 );
and \U$8971 ( \9144 , \8988 , \9003 );
and \U$8972 ( \9145 , \8974 , \9003 );
or \U$8973 ( \9146 , \9143 , \9144 , \9145 );
xor \U$8974 ( \9147 , \9142 , \9146 );
and \U$8975 ( \9148 , \9008 , \9022 );
and \U$8976 ( \9149 , \9022 , \9037 );
and \U$8977 ( \9150 , \9008 , \9037 );
or \U$8978 ( \9151 , \9148 , \9149 , \9150 );
xor \U$8979 ( \9152 , \9147 , \9151 );
xor \U$8980 ( \9153 , \9138 , \9152 );
and \U$8981 ( \9154 , \8920 , \8924 );
and \U$8982 ( \9155 , \8924 , \8929 );
and \U$8983 ( \9156 , \8920 , \8929 );
or \U$8984 ( \9157 , \9154 , \9155 , \9156 );
and \U$8985 ( \9158 , \8838 , \8842 );
and \U$8986 ( \9159 , \8842 , \8848 );
and \U$8987 ( \9160 , \8838 , \8848 );
or \U$8988 ( \9161 , \9158 , \9159 , \9160 );
xor \U$8989 ( \9162 , \9157 , \9161 );
and \U$8990 ( \9163 , \8854 , \8858 );
and \U$8991 ( \9164 , \8858 , \8863 );
and \U$8992 ( \9165 , \8854 , \8863 );
or \U$8993 ( \9166 , \9163 , \9164 , \9165 );
xor \U$8994 ( \9167 , \9162 , \9166 );
and \U$8995 ( \9168 , \8835 , \183 );
buf \U$8996 ( \9169 , RIb55efe0_69);
and \U$8997 ( \9170 , \9169 , \180 );
nor \U$8998 ( \9171 , \9168 , \9170 );
xnor \U$8999 ( \9172 , \9171 , \179 );
and \U$9000 ( \9173 , \8349 , \195 );
and \U$9001 ( \9174 , \8652 , \193 );
nor \U$9002 ( \9175 , \9173 , \9174 );
xnor \U$9003 ( \9176 , \9175 , \202 );
xor \U$9004 ( \9177 , \9172 , \9176 );
and \U$9005 ( \9178 , \7700 , \215 );
and \U$9006 ( \9179 , \8057 , \213 );
nor \U$9007 ( \9180 , \9178 , \9179 );
xnor \U$9008 ( \9181 , \9180 , \222 );
xor \U$9009 ( \9182 , \9177 , \9181 );
and \U$9010 ( \9183 , \7231 , \230 );
and \U$9011 ( \9184 , \7556 , \228 );
nor \U$9012 ( \9185 , \9183 , \9184 );
xnor \U$9013 ( \9186 , \9185 , \237 );
and \U$9014 ( \9187 , \6790 , \245 );
and \U$9015 ( \9188 , \6945 , \243 );
nor \U$9016 ( \9189 , \9187 , \9188 );
xnor \U$9017 ( \9190 , \9189 , \252 );
xor \U$9018 ( \9191 , \9186 , \9190 );
and \U$9019 ( \9192 , \6281 , \141 );
and \U$9020 ( \9193 , \6514 , \139 );
nor \U$9021 ( \9194 , \9192 , \9193 );
xnor \U$9022 ( \9195 , \9194 , \148 );
xor \U$9023 ( \9196 , \9191 , \9195 );
xor \U$9024 ( \9197 , \9182 , \9196 );
and \U$9025 ( \9198 , \5674 , \156 );
and \U$9026 ( \9199 , \6030 , \154 );
nor \U$9027 ( \9200 , \9198 , \9199 );
xnor \U$9028 ( \9201 , \9200 , \163 );
and \U$9029 ( \9202 , \5156 , \296 );
and \U$9030 ( \9203 , \5469 , \168 );
nor \U$9031 ( \9204 , \9202 , \9203 );
xnor \U$9032 ( \9205 , \9204 , \173 );
xor \U$9033 ( \9206 , \9201 , \9205 );
and \U$9034 ( \9207 , \4749 , \438 );
and \U$9035 ( \9208 , \4922 , \336 );
nor \U$9036 ( \9209 , \9207 , \9208 );
xnor \U$9037 ( \9210 , \9209 , \320 );
xor \U$9038 ( \9211 , \9206 , \9210 );
and \U$9039 ( \9212 , \4364 , \1086 );
and \U$9040 ( \9213 , \4654 , \508 );
nor \U$9041 ( \9214 , \9212 , \9213 );
xnor \U$9042 ( \9215 , \9214 , \487 );
and \U$9043 ( \9216 , \3912 , \1301 );
and \U$9044 ( \9217 , \4160 , \1246 );
nor \U$9045 ( \9218 , \9216 , \9217 );
xnor \U$9046 ( \9219 , \9218 , \1205 );
xor \U$9047 ( \9220 , \9215 , \9219 );
and \U$9048 ( \9221 , \3646 , \1578 );
and \U$9049 ( \9222 , \3736 , \1431 );
nor \U$9050 ( \9223 , \9221 , \9222 );
xnor \U$9051 ( \9224 , \9223 , \1436 );
xor \U$9052 ( \9225 , \9220 , \9224 );
xor \U$9053 ( \9226 , \9211 , \9225 );
and \U$9054 ( \9227 , \3143 , \1824 );
and \U$9055 ( \9228 , \3395 , \1739 );
nor \U$9056 ( \9229 , \9227 , \9228 );
xnor \U$9057 ( \9230 , \9229 , \1697 );
and \U$9058 ( \9231 , \2826 , \2121 );
and \U$9059 ( \9232 , \3037 , \2008 );
nor \U$9060 ( \9233 , \9231 , \9232 );
xnor \U$9061 ( \9234 , \9233 , \1961 );
xor \U$9062 ( \9235 , \9230 , \9234 );
and \U$9063 ( \9236 , \2521 , \2400 );
and \U$9064 ( \9237 , \2757 , \2246 );
nor \U$9065 ( \9238 , \9236 , \9237 );
xnor \U$9066 ( \9239 , \9238 , \2195 );
xor \U$9067 ( \9240 , \9235 , \9239 );
xor \U$9068 ( \9241 , \9226 , \9240 );
xor \U$9069 ( \9242 , \9197 , \9241 );
xor \U$9070 ( \9243 , \9167 , \9242 );
and \U$9071 ( \9244 , \8978 , \8982 );
and \U$9072 ( \9245 , \8982 , \8987 );
and \U$9073 ( \9246 , \8978 , \8987 );
or \U$9074 ( \9247 , \9244 , \9245 , \9246 );
and \U$9075 ( \9248 , \8993 , \8997 );
and \U$9076 ( \9249 , \8997 , \9002 );
and \U$9077 ( \9250 , \8993 , \9002 );
or \U$9078 ( \9251 , \9248 , \9249 , \9250 );
xor \U$9079 ( \9252 , \9247 , \9251 );
and \U$9080 ( \9253 , \9012 , \9016 );
and \U$9081 ( \9254 , \9016 , \9021 );
and \U$9082 ( \9255 , \9012 , \9021 );
or \U$9083 ( \9256 , \9253 , \9254 , \9255 );
xor \U$9084 ( \9257 , \9252 , \9256 );
and \U$9085 ( \9258 , \2182 , \2669 );
and \U$9086 ( \9259 , \2366 , \2538 );
nor \U$9087 ( \9260 , \9258 , \9259 );
xnor \U$9088 ( \9261 , \9260 , \2534 );
and \U$9089 ( \9262 , \1948 , \3103 );
and \U$9090 ( \9263 , \2090 , \2934 );
nor \U$9091 ( \9264 , \9262 , \9263 );
xnor \U$9092 ( \9265 , \9264 , \2839 );
xor \U$9093 ( \9266 , \9261 , \9265 );
and \U$9094 ( \9267 , \1684 , \3357 );
and \U$9095 ( \9268 , \1802 , \3255 );
nor \U$9096 ( \9269 , \9267 , \9268 );
xnor \U$9097 ( \9270 , \9269 , \3156 );
xor \U$9098 ( \9271 , \9266 , \9270 );
and \U$9099 ( \9272 , \1484 , \3813 );
and \U$9100 ( \9273 , \1601 , \3557 );
nor \U$9101 ( \9274 , \9272 , \9273 );
xnor \U$9102 ( \9275 , \9274 , \3562 );
and \U$9103 ( \9276 , \1192 , \4132 );
and \U$9104 ( \9277 , \1333 , \4012 );
nor \U$9105 ( \9278 , \9276 , \9277 );
xnor \U$9106 ( \9279 , \9278 , \3925 );
xor \U$9107 ( \9280 , \9275 , \9279 );
and \U$9108 ( \9281 , \474 , \4581 );
and \U$9109 ( \9282 , \1147 , \4424 );
nor \U$9110 ( \9283 , \9281 , \9282 );
xnor \U$9111 ( \9284 , \9283 , \4377 );
xor \U$9112 ( \9285 , \9280 , \9284 );
xor \U$9113 ( \9286 , \9271 , \9285 );
and \U$9114 ( \9287 , \307 , \5011 );
and \U$9115 ( \9288 , \412 , \4878 );
nor \U$9116 ( \9289 , \9287 , \9288 );
xnor \U$9117 ( \9290 , \9289 , \4762 );
and \U$9118 ( \9291 , \185 , \5485 );
and \U$9119 ( \9292 , \261 , \5275 );
nor \U$9120 ( \9293 , \9291 , \9292 );
xnor \U$9121 ( \9294 , \9293 , \5169 );
xor \U$9122 ( \9295 , \9290 , \9294 );
and \U$9123 ( \9296 , \197 , \5996 );
and \U$9124 ( \9297 , \178 , \5695 );
nor \U$9125 ( \9298 , \9296 , \9297 );
xnor \U$9126 ( \9299 , \9298 , \5687 );
xor \U$9127 ( \9300 , \9295 , \9299 );
xor \U$9128 ( \9301 , \9286 , \9300 );
xor \U$9129 ( \9302 , \9257 , \9301 );
and \U$9130 ( \9303 , \9027 , \9031 );
and \U$9131 ( \9304 , \9031 , \9036 );
and \U$9132 ( \9305 , \9027 , \9036 );
or \U$9133 ( \9306 , \9303 , \9304 , \9305 );
and \U$9134 ( \9307 , \217 , \6401 );
and \U$9135 ( \9308 , \189 , \6143 );
nor \U$9136 ( \9309 , \9307 , \9308 );
xnor \U$9137 ( \9310 , \9309 , \6148 );
and \U$9138 ( \9311 , \232 , \7055 );
and \U$9139 ( \9312 , \209 , \6675 );
nor \U$9140 ( \9313 , \9311 , \9312 );
xnor \U$9141 ( \9314 , \9313 , \6680 );
xor \U$9142 ( \9315 , \9310 , \9314 );
and \U$9143 ( \9316 , \247 , \7489 );
and \U$9144 ( \9317 , \224 , \7137 );
nor \U$9145 ( \9318 , \9316 , \9317 );
xnor \U$9146 ( \9319 , \9318 , \7142 );
xor \U$9147 ( \9320 , \9315 , \9319 );
xor \U$9148 ( \9321 , \9306 , \9320 );
and \U$9149 ( \9322 , \143 , \8019 );
and \U$9150 ( \9323 , \240 , \7830 );
nor \U$9151 ( \9324 , \9322 , \9323 );
xnor \U$9152 ( \9325 , \9324 , \7713 );
and \U$9153 ( \9326 , \158 , \8540 );
and \U$9154 ( \9327 , \134 , \8292 );
nor \U$9155 ( \9328 , \9326 , \9327 );
xnor \U$9156 ( \9329 , \9328 , \8297 );
xor \U$9157 ( \9330 , \9325 , \9329 );
xor \U$9158 ( \9331 , \8844 , \8845 );
not \U$9159 ( \9332 , \9006 );
and \U$9160 ( \9333 , \9331 , \9332 );
and \U$9161 ( \9334 , \166 , \9333 );
and \U$9162 ( \9335 , \150 , \9006 );
nor \U$9163 ( \9336 , \9334 , \9335 );
xnor \U$9164 ( \9337 , \9336 , \8848 );
xor \U$9165 ( \9338 , \9330 , \9337 );
xor \U$9166 ( \9339 , \9321 , \9338 );
xor \U$9167 ( \9340 , \9302 , \9339 );
xor \U$9168 ( \9341 , \9243 , \9340 );
xor \U$9169 ( \9342 , \9153 , \9341 );
xor \U$9170 ( \9343 , \9124 , \9342 );
xor \U$9171 ( \9344 , \9095 , \9343 );
xor \U$9172 ( \9345 , \9056 , \9344 );
and \U$9173 ( \9346 , \8758 , \9043 );
xor \U$9174 ( \9347 , \9345 , \9346 );
and \U$9175 ( \9348 , \9044 , \9045 );
and \U$9176 ( \9349 , \9046 , \9049 );
or \U$9177 ( \9350 , \9348 , \9349 );
xor \U$9178 ( \9351 , \9347 , \9350 );
buf g5525_GF_PartitionCandidate( \9352_nG5525 , \9351 );
buf \U$9179 ( \9353 , \9352_nG5525 );
and \U$9180 ( \9354 , \9060 , \9094 );
and \U$9181 ( \9355 , \9094 , \9343 );
and \U$9182 ( \9356 , \9060 , \9343 );
or \U$9183 ( \9357 , \9354 , \9355 , \9356 );
and \U$9184 ( \9358 , \9064 , \9068 );
and \U$9185 ( \9359 , \9068 , \9093 );
and \U$9186 ( \9360 , \9064 , \9093 );
or \U$9187 ( \9361 , \9358 , \9359 , \9360 );
and \U$9188 ( \9362 , \9109 , \9123 );
and \U$9189 ( \9363 , \9123 , \9342 );
and \U$9190 ( \9364 , \9109 , \9342 );
or \U$9191 ( \9365 , \9362 , \9363 , \9364 );
xor \U$9192 ( \9366 , \9361 , \9365 );
and \U$9193 ( \9367 , \9099 , \9103 );
and \U$9194 ( \9368 , \9103 , \9108 );
and \U$9195 ( \9369 , \9099 , \9108 );
or \U$9196 ( \9370 , \9367 , \9368 , \9369 );
and \U$9197 ( \9371 , \9073 , \9077 );
and \U$9198 ( \9372 , \9077 , \9092 );
and \U$9199 ( \9373 , \9073 , \9092 );
or \U$9200 ( \9374 , \9371 , \9372 , \9373 );
xor \U$9201 ( \9375 , \9370 , \9374 );
and \U$9202 ( \9376 , \9167 , \9242 );
and \U$9203 ( \9377 , \9242 , \9340 );
and \U$9204 ( \9378 , \9167 , \9340 );
or \U$9205 ( \9379 , \9376 , \9377 , \9378 );
xor \U$9206 ( \9380 , \9375 , \9379 );
xor \U$9207 ( \9381 , \9366 , \9380 );
xor \U$9208 ( \9382 , \9357 , \9381 );
and \U$9209 ( \9383 , \9113 , \9117 );
and \U$9210 ( \9384 , \9117 , \9122 );
and \U$9211 ( \9385 , \9113 , \9122 );
or \U$9212 ( \9386 , \9383 , \9384 , \9385 );
and \U$9213 ( \9387 , \9138 , \9152 );
and \U$9214 ( \9388 , \9152 , \9341 );
and \U$9215 ( \9389 , \9138 , \9341 );
or \U$9216 ( \9390 , \9387 , \9388 , \9389 );
xor \U$9217 ( \9391 , \9386 , \9390 );
and \U$9218 ( \9392 , \9128 , \9132 );
and \U$9219 ( \9393 , \9132 , \9137 );
and \U$9220 ( \9394 , \9128 , \9137 );
or \U$9221 ( \9395 , \9392 , \9393 , \9394 );
and \U$9222 ( \9396 , \9142 , \9146 );
and \U$9223 ( \9397 , \9146 , \9151 );
and \U$9224 ( \9398 , \9142 , \9151 );
or \U$9225 ( \9399 , \9396 , \9397 , \9398 );
xor \U$9226 ( \9400 , \9395 , \9399 );
and \U$9227 ( \9401 , \9182 , \9196 );
and \U$9228 ( \9402 , \9196 , \9241 );
and \U$9229 ( \9403 , \9182 , \9241 );
or \U$9230 ( \9404 , \9401 , \9402 , \9403 );
xor \U$9231 ( \9405 , \9400 , \9404 );
and \U$9232 ( \9406 , \9271 , \9285 );
and \U$9233 ( \9407 , \9285 , \9300 );
and \U$9234 ( \9408 , \9271 , \9300 );
or \U$9235 ( \9409 , \9406 , \9407 , \9408 );
and \U$9236 ( \9410 , \9306 , \9320 );
and \U$9237 ( \9411 , \9320 , \9338 );
and \U$9238 ( \9412 , \9306 , \9338 );
or \U$9239 ( \9413 , \9410 , \9411 , \9412 );
xor \U$9240 ( \9414 , \9409 , \9413 );
and \U$9241 ( \9415 , \9211 , \9225 );
and \U$9242 ( \9416 , \9225 , \9240 );
and \U$9243 ( \9417 , \9211 , \9240 );
or \U$9244 ( \9418 , \9415 , \9416 , \9417 );
xor \U$9245 ( \9419 , \9414 , \9418 );
and \U$9246 ( \9420 , \9157 , \9161 );
and \U$9247 ( \9421 , \9161 , \9166 );
and \U$9248 ( \9422 , \9157 , \9166 );
or \U$9249 ( \9423 , \9420 , \9421 , \9422 );
and \U$9250 ( \9424 , \9082 , \9086 );
and \U$9251 ( \9425 , \9086 , \9091 );
and \U$9252 ( \9426 , \9082 , \9091 );
or \U$9253 ( \9427 , \9424 , \9425 , \9426 );
xor \U$9254 ( \9428 , \9423 , \9427 );
and \U$9255 ( \9429 , \9247 , \9251 );
and \U$9256 ( \9430 , \9251 , \9256 );
and \U$9257 ( \9431 , \9247 , \9256 );
or \U$9258 ( \9432 , \9429 , \9430 , \9431 );
xor \U$9259 ( \9433 , \9428 , \9432 );
xor \U$9260 ( \9434 , \9419 , \9433 );
and \U$9261 ( \9435 , \6514 , \141 );
and \U$9262 ( \9436 , \6790 , \139 );
nor \U$9263 ( \9437 , \9435 , \9436 );
xnor \U$9264 ( \9438 , \9437 , \148 );
and \U$9265 ( \9439 , \6030 , \156 );
and \U$9266 ( \9440 , \6281 , \154 );
nor \U$9267 ( \9441 , \9439 , \9440 );
xnor \U$9268 ( \9442 , \9441 , \163 );
xor \U$9269 ( \9443 , \9438 , \9442 );
and \U$9270 ( \9444 , \5469 , \296 );
and \U$9271 ( \9445 , \5674 , \168 );
nor \U$9272 ( \9446 , \9444 , \9445 );
xnor \U$9273 ( \9447 , \9446 , \173 );
xor \U$9274 ( \9448 , \9443 , \9447 );
and \U$9275 ( \9449 , \8057 , \215 );
and \U$9276 ( \9450 , \8349 , \213 );
nor \U$9277 ( \9451 , \9449 , \9450 );
xnor \U$9278 ( \9452 , \9451 , \222 );
and \U$9279 ( \9453 , \7556 , \230 );
and \U$9280 ( \9454 , \7700 , \228 );
nor \U$9281 ( \9455 , \9453 , \9454 );
xnor \U$9282 ( \9456 , \9455 , \237 );
xor \U$9283 ( \9457 , \9452 , \9456 );
and \U$9284 ( \9458 , \6945 , \245 );
and \U$9285 ( \9459 , \7231 , \243 );
nor \U$9286 ( \9460 , \9458 , \9459 );
xnor \U$9287 ( \9461 , \9460 , \252 );
xor \U$9288 ( \9462 , \9457 , \9461 );
xor \U$9289 ( \9463 , \9448 , \9462 );
and \U$9290 ( \9464 , \9169 , \183 );
buf \U$9291 ( \9465 , RIb55f058_68);
and \U$9292 ( \9466 , \9465 , \180 );
nor \U$9293 ( \9467 , \9464 , \9466 );
xnor \U$9294 ( \9468 , \9467 , \179 );
and \U$9295 ( \9469 , \8652 , \195 );
and \U$9296 ( \9470 , \8835 , \193 );
nor \U$9297 ( \9471 , \9469 , \9470 );
xnor \U$9298 ( \9472 , \9471 , \202 );
xor \U$9299 ( \9473 , \9468 , \9472 );
buf \U$9300 ( \9474 , RIb560ed0_3);
buf \U$9301 ( \9475 , RIb560e58_4);
and \U$9302 ( \9476 , \9475 , \8844 );
not \U$9303 ( \9477 , \9476 );
and \U$9304 ( \9478 , \9474 , \9477 );
xor \U$9305 ( \9479 , \9473 , \9478 );
xor \U$9306 ( \9480 , \9463 , \9479 );
and \U$9307 ( \9481 , \178 , \5996 );
and \U$9308 ( \9482 , \185 , \5695 );
nor \U$9309 ( \9483 , \9481 , \9482 );
xnor \U$9310 ( \9484 , \9483 , \5687 );
and \U$9311 ( \9485 , \189 , \6401 );
and \U$9312 ( \9486 , \197 , \6143 );
nor \U$9313 ( \9487 , \9485 , \9486 );
xnor \U$9314 ( \9488 , \9487 , \6148 );
xor \U$9315 ( \9489 , \9484 , \9488 );
and \U$9316 ( \9490 , \209 , \7055 );
and \U$9317 ( \9491 , \217 , \6675 );
nor \U$9318 ( \9492 , \9490 , \9491 );
xnor \U$9319 ( \9493 , \9492 , \6680 );
xor \U$9320 ( \9494 , \9489 , \9493 );
and \U$9321 ( \9495 , \1802 , \3357 );
and \U$9322 ( \9496 , \1948 , \3255 );
nor \U$9323 ( \9497 , \9495 , \9496 );
xnor \U$9324 ( \9498 , \9497 , \3156 );
and \U$9325 ( \9499 , \1601 , \3813 );
and \U$9326 ( \9500 , \1684 , \3557 );
nor \U$9327 ( \9501 , \9499 , \9500 );
xnor \U$9328 ( \9502 , \9501 , \3562 );
xor \U$9329 ( \9503 , \9498 , \9502 );
and \U$9330 ( \9504 , \1333 , \4132 );
and \U$9331 ( \9505 , \1484 , \4012 );
nor \U$9332 ( \9506 , \9504 , \9505 );
xnor \U$9333 ( \9507 , \9506 , \3925 );
xor \U$9334 ( \9508 , \9503 , \9507 );
xor \U$9335 ( \9509 , \9494 , \9508 );
and \U$9336 ( \9510 , \1147 , \4581 );
and \U$9337 ( \9511 , \1192 , \4424 );
nor \U$9338 ( \9512 , \9510 , \9511 );
xnor \U$9339 ( \9513 , \9512 , \4377 );
and \U$9340 ( \9514 , \412 , \5011 );
and \U$9341 ( \9515 , \474 , \4878 );
nor \U$9342 ( \9516 , \9514 , \9515 );
xnor \U$9343 ( \9517 , \9516 , \4762 );
xor \U$9344 ( \9518 , \9513 , \9517 );
and \U$9345 ( \9519 , \261 , \5485 );
and \U$9346 ( \9520 , \307 , \5275 );
nor \U$9347 ( \9521 , \9519 , \9520 );
xnor \U$9348 ( \9522 , \9521 , \5169 );
xor \U$9349 ( \9523 , \9518 , \9522 );
xor \U$9350 ( \9524 , \9509 , \9523 );
xor \U$9351 ( \9525 , \9480 , \9524 );
and \U$9352 ( \9526 , \4922 , \438 );
and \U$9353 ( \9527 , \5156 , \336 );
nor \U$9354 ( \9528 , \9526 , \9527 );
xnor \U$9355 ( \9529 , \9528 , \320 );
and \U$9356 ( \9530 , \4654 , \1086 );
and \U$9357 ( \9531 , \4749 , \508 );
nor \U$9358 ( \9532 , \9530 , \9531 );
xnor \U$9359 ( \9533 , \9532 , \487 );
xor \U$9360 ( \9534 , \9529 , \9533 );
and \U$9361 ( \9535 , \4160 , \1301 );
and \U$9362 ( \9536 , \4364 , \1246 );
nor \U$9363 ( \9537 , \9535 , \9536 );
xnor \U$9364 ( \9538 , \9537 , \1205 );
xor \U$9365 ( \9539 , \9534 , \9538 );
and \U$9366 ( \9540 , \3736 , \1578 );
and \U$9367 ( \9541 , \3912 , \1431 );
nor \U$9368 ( \9542 , \9540 , \9541 );
xnor \U$9369 ( \9543 , \9542 , \1436 );
and \U$9370 ( \9544 , \3395 , \1824 );
and \U$9371 ( \9545 , \3646 , \1739 );
nor \U$9372 ( \9546 , \9544 , \9545 );
xnor \U$9373 ( \9547 , \9546 , \1697 );
xor \U$9374 ( \9548 , \9543 , \9547 );
and \U$9375 ( \9549 , \3037 , \2121 );
and \U$9376 ( \9550 , \3143 , \2008 );
nor \U$9377 ( \9551 , \9549 , \9550 );
xnor \U$9378 ( \9552 , \9551 , \1961 );
xor \U$9379 ( \9553 , \9548 , \9552 );
xor \U$9380 ( \9554 , \9539 , \9553 );
and \U$9381 ( \9555 , \2757 , \2400 );
and \U$9382 ( \9556 , \2826 , \2246 );
nor \U$9383 ( \9557 , \9555 , \9556 );
xnor \U$9384 ( \9558 , \9557 , \2195 );
and \U$9385 ( \9559 , \2366 , \2669 );
and \U$9386 ( \9560 , \2521 , \2538 );
nor \U$9387 ( \9561 , \9559 , \9560 );
xnor \U$9388 ( \9562 , \9561 , \2534 );
xor \U$9389 ( \9563 , \9558 , \9562 );
and \U$9390 ( \9564 , \2090 , \3103 );
and \U$9391 ( \9565 , \2182 , \2934 );
nor \U$9392 ( \9566 , \9564 , \9565 );
xnor \U$9393 ( \9567 , \9566 , \2839 );
xor \U$9394 ( \9568 , \9563 , \9567 );
xor \U$9395 ( \9569 , \9554 , \9568 );
xor \U$9396 ( \9570 , \9525 , \9569 );
xor \U$9397 ( \9571 , \9434 , \9570 );
xor \U$9398 ( \9572 , \9405 , \9571 );
and \U$9399 ( \9573 , \9257 , \9301 );
and \U$9400 ( \9574 , \9301 , \9339 );
and \U$9401 ( \9575 , \9257 , \9339 );
or \U$9402 ( \9576 , \9573 , \9574 , \9575 );
and \U$9403 ( \9577 , \9201 , \9205 );
and \U$9404 ( \9578 , \9205 , \9210 );
and \U$9405 ( \9579 , \9201 , \9210 );
or \U$9406 ( \9580 , \9577 , \9578 , \9579 );
and \U$9407 ( \9581 , \9172 , \9176 );
and \U$9408 ( \9582 , \9176 , \9181 );
and \U$9409 ( \9583 , \9172 , \9181 );
or \U$9410 ( \9584 , \9581 , \9582 , \9583 );
xor \U$9411 ( \9585 , \9580 , \9584 );
and \U$9412 ( \9586 , \9186 , \9190 );
and \U$9413 ( \9587 , \9190 , \9195 );
and \U$9414 ( \9588 , \9186 , \9195 );
or \U$9415 ( \9589 , \9586 , \9587 , \9588 );
xor \U$9416 ( \9590 , \9585 , \9589 );
xor \U$9417 ( \9591 , \9576 , \9590 );
and \U$9418 ( \9592 , \9261 , \9265 );
and \U$9419 ( \9593 , \9265 , \9270 );
and \U$9420 ( \9594 , \9261 , \9270 );
or \U$9421 ( \9595 , \9592 , \9593 , \9594 );
and \U$9422 ( \9596 , \9215 , \9219 );
and \U$9423 ( \9597 , \9219 , \9224 );
and \U$9424 ( \9598 , \9215 , \9224 );
or \U$9425 ( \9599 , \9596 , \9597 , \9598 );
xor \U$9426 ( \9600 , \9595 , \9599 );
and \U$9427 ( \9601 , \9230 , \9234 );
and \U$9428 ( \9602 , \9234 , \9239 );
and \U$9429 ( \9603 , \9230 , \9239 );
or \U$9430 ( \9604 , \9601 , \9602 , \9603 );
xor \U$9431 ( \9605 , \9600 , \9604 );
and \U$9432 ( \9606 , \9275 , \9279 );
and \U$9433 ( \9607 , \9279 , \9284 );
and \U$9434 ( \9608 , \9275 , \9284 );
or \U$9435 ( \9609 , \9606 , \9607 , \9608 );
and \U$9436 ( \9610 , \9310 , \9314 );
and \U$9437 ( \9611 , \9314 , \9319 );
and \U$9438 ( \9612 , \9310 , \9319 );
or \U$9439 ( \9613 , \9610 , \9611 , \9612 );
xor \U$9440 ( \9614 , \9609 , \9613 );
and \U$9441 ( \9615 , \9290 , \9294 );
and \U$9442 ( \9616 , \9294 , \9299 );
and \U$9443 ( \9617 , \9290 , \9299 );
or \U$9444 ( \9618 , \9615 , \9616 , \9617 );
xor \U$9445 ( \9619 , \9614 , \9618 );
xor \U$9446 ( \9620 , \9605 , \9619 );
and \U$9447 ( \9621 , \9325 , \9329 );
and \U$9448 ( \9622 , \9329 , \9337 );
and \U$9449 ( \9623 , \9325 , \9337 );
or \U$9450 ( \9624 , \9621 , \9622 , \9623 );
and \U$9451 ( \9625 , \224 , \7489 );
and \U$9452 ( \9626 , \232 , \7137 );
nor \U$9453 ( \9627 , \9625 , \9626 );
xnor \U$9454 ( \9628 , \9627 , \7142 );
and \U$9455 ( \9629 , \240 , \8019 );
and \U$9456 ( \9630 , \247 , \7830 );
nor \U$9457 ( \9631 , \9629 , \9630 );
xnor \U$9458 ( \9632 , \9631 , \7713 );
xor \U$9459 ( \9633 , \9628 , \9632 );
and \U$9460 ( \9634 , \134 , \8540 );
and \U$9461 ( \9635 , \143 , \8292 );
nor \U$9462 ( \9636 , \9634 , \9635 );
xnor \U$9463 ( \9637 , \9636 , \8297 );
xor \U$9464 ( \9638 , \9633 , \9637 );
xor \U$9465 ( \9639 , \9624 , \9638 );
and \U$9466 ( \9640 , \150 , \9333 );
and \U$9467 ( \9641 , \158 , \9006 );
nor \U$9468 ( \9642 , \9640 , \9641 );
xnor \U$9469 ( \9643 , \9642 , \8848 );
xor \U$9470 ( \9644 , \9475 , \8844 );
nand \U$9471 ( \9645 , \166 , \9644 );
xnor \U$9472 ( \9646 , \9645 , \9478 );
xor \U$9473 ( \9647 , \9643 , \9646 );
xor \U$9474 ( \9648 , \9639 , \9647 );
xor \U$9475 ( \9649 , \9620 , \9648 );
xor \U$9476 ( \9650 , \9591 , \9649 );
xor \U$9477 ( \9651 , \9572 , \9650 );
xor \U$9478 ( \9652 , \9391 , \9651 );
xor \U$9479 ( \9653 , \9382 , \9652 );
and \U$9480 ( \9654 , \9056 , \9344 );
xor \U$9481 ( \9655 , \9653 , \9654 );
and \U$9482 ( \9656 , \9345 , \9346 );
and \U$9483 ( \9657 , \9347 , \9350 );
or \U$9484 ( \9658 , \9656 , \9657 );
xor \U$9485 ( \9659 , \9655 , \9658 );
buf g5523_GF_PartitionCandidate( \9660_nG5523 , \9659 );
buf \U$9486 ( \9661 , \9660_nG5523 );
and \U$9487 ( \9662 , \9361 , \9365 );
and \U$9488 ( \9663 , \9365 , \9380 );
and \U$9489 ( \9664 , \9361 , \9380 );
or \U$9490 ( \9665 , \9662 , \9663 , \9664 );
and \U$9491 ( \9666 , \9386 , \9390 );
and \U$9492 ( \9667 , \9390 , \9651 );
and \U$9493 ( \9668 , \9386 , \9651 );
or \U$9494 ( \9669 , \9666 , \9667 , \9668 );
and \U$9495 ( \9670 , \9395 , \9399 );
and \U$9496 ( \9671 , \9399 , \9404 );
and \U$9497 ( \9672 , \9395 , \9404 );
or \U$9498 ( \9673 , \9670 , \9671 , \9672 );
and \U$9499 ( \9674 , \9419 , \9433 );
and \U$9500 ( \9675 , \9433 , \9570 );
and \U$9501 ( \9676 , \9419 , \9570 );
or \U$9502 ( \9677 , \9674 , \9675 , \9676 );
xor \U$9503 ( \9678 , \9673 , \9677 );
and \U$9504 ( \9679 , \9576 , \9590 );
and \U$9505 ( \9680 , \9590 , \9649 );
and \U$9506 ( \9681 , \9576 , \9649 );
or \U$9507 ( \9682 , \9679 , \9680 , \9681 );
xor \U$9508 ( \9683 , \9678 , \9682 );
xor \U$9509 ( \9684 , \9669 , \9683 );
and \U$9510 ( \9685 , \9370 , \9374 );
and \U$9511 ( \9686 , \9374 , \9379 );
and \U$9512 ( \9687 , \9370 , \9379 );
or \U$9513 ( \9688 , \9685 , \9686 , \9687 );
and \U$9514 ( \9689 , \9405 , \9571 );
and \U$9515 ( \9690 , \9571 , \9650 );
and \U$9516 ( \9691 , \9405 , \9650 );
or \U$9517 ( \9692 , \9689 , \9690 , \9691 );
xor \U$9518 ( \9693 , \9688 , \9692 );
and \U$9519 ( \9694 , \9409 , \9413 );
and \U$9520 ( \9695 , \9413 , \9418 );
and \U$9521 ( \9696 , \9409 , \9418 );
or \U$9522 ( \9697 , \9694 , \9695 , \9696 );
and \U$9523 ( \9698 , \9423 , \9427 );
and \U$9524 ( \9699 , \9427 , \9432 );
and \U$9525 ( \9700 , \9423 , \9432 );
or \U$9526 ( \9701 , \9698 , \9699 , \9700 );
xor \U$9527 ( \9702 , \9697 , \9701 );
and \U$9528 ( \9703 , \9480 , \9524 );
and \U$9529 ( \9704 , \9524 , \9569 );
and \U$9530 ( \9705 , \9480 , \9569 );
or \U$9531 ( \9706 , \9703 , \9704 , \9705 );
xor \U$9532 ( \9707 , \9702 , \9706 );
and \U$9533 ( \9708 , \9605 , \9619 );
and \U$9534 ( \9709 , \9619 , \9648 );
and \U$9535 ( \9710 , \9605 , \9648 );
or \U$9536 ( \9711 , \9708 , \9709 , \9710 );
and \U$9537 ( \9712 , \9484 , \9488 );
and \U$9538 ( \9713 , \9488 , \9493 );
and \U$9539 ( \9714 , \9484 , \9493 );
or \U$9540 ( \9715 , \9712 , \9713 , \9714 );
and \U$9541 ( \9716 , \9498 , \9502 );
and \U$9542 ( \9717 , \9502 , \9507 );
and \U$9543 ( \9718 , \9498 , \9507 );
or \U$9544 ( \9719 , \9716 , \9717 , \9718 );
xor \U$9545 ( \9720 , \9715 , \9719 );
and \U$9546 ( \9721 , \9513 , \9517 );
and \U$9547 ( \9722 , \9517 , \9522 );
and \U$9548 ( \9723 , \9513 , \9522 );
or \U$9549 ( \9724 , \9721 , \9722 , \9723 );
xor \U$9550 ( \9725 , \9720 , \9724 );
and \U$9551 ( \9726 , \9438 , \9442 );
and \U$9552 ( \9727 , \9442 , \9447 );
and \U$9553 ( \9728 , \9438 , \9447 );
or \U$9554 ( \9729 , \9726 , \9727 , \9728 );
and \U$9555 ( \9730 , \9452 , \9456 );
and \U$9556 ( \9731 , \9456 , \9461 );
and \U$9557 ( \9732 , \9452 , \9461 );
or \U$9558 ( \9733 , \9730 , \9731 , \9732 );
xor \U$9559 ( \9734 , \9729 , \9733 );
and \U$9560 ( \9735 , \9468 , \9472 );
and \U$9561 ( \9736 , \9472 , \9478 );
and \U$9562 ( \9737 , \9468 , \9478 );
or \U$9563 ( \9738 , \9735 , \9736 , \9737 );
xor \U$9564 ( \9739 , \9734 , \9738 );
xor \U$9565 ( \9740 , \9725 , \9739 );
and \U$9566 ( \9741 , \9529 , \9533 );
and \U$9567 ( \9742 , \9533 , \9538 );
and \U$9568 ( \9743 , \9529 , \9538 );
or \U$9569 ( \9744 , \9741 , \9742 , \9743 );
and \U$9570 ( \9745 , \9543 , \9547 );
and \U$9571 ( \9746 , \9547 , \9552 );
and \U$9572 ( \9747 , \9543 , \9552 );
or \U$9573 ( \9748 , \9745 , \9746 , \9747 );
xor \U$9574 ( \9749 , \9744 , \9748 );
and \U$9575 ( \9750 , \9558 , \9562 );
and \U$9576 ( \9751 , \9562 , \9567 );
and \U$9577 ( \9752 , \9558 , \9567 );
or \U$9578 ( \9753 , \9750 , \9751 , \9752 );
xor \U$9579 ( \9754 , \9749 , \9753 );
xor \U$9580 ( \9755 , \9740 , \9754 );
xor \U$9581 ( \9756 , \9711 , \9755 );
and \U$9582 ( \9757 , \9628 , \9632 );
and \U$9583 ( \9758 , \9632 , \9637 );
and \U$9584 ( \9759 , \9628 , \9637 );
or \U$9585 ( \9760 , \9757 , \9758 , \9759 );
and \U$9586 ( \9761 , \9643 , \9646 );
xor \U$9587 ( \9762 , \9760 , \9761 );
xor \U$9588 ( \9763 , \9474 , \9475 );
not \U$9589 ( \9764 , \9644 );
and \U$9590 ( \9765 , \9763 , \9764 );
and \U$9591 ( \9766 , \166 , \9765 );
and \U$9592 ( \9767 , \150 , \9644 );
nor \U$9593 ( \9768 , \9766 , \9767 );
xnor \U$9594 ( \9769 , \9768 , \9478 );
xor \U$9595 ( \9770 , \9762 , \9769 );
and \U$9596 ( \9771 , \1684 , \3813 );
and \U$9597 ( \9772 , \1802 , \3557 );
nor \U$9598 ( \9773 , \9771 , \9772 );
xnor \U$9599 ( \9774 , \9773 , \3562 );
and \U$9600 ( \9775 , \1484 , \4132 );
and \U$9601 ( \9776 , \1601 , \4012 );
nor \U$9602 ( \9777 , \9775 , \9776 );
xnor \U$9603 ( \9778 , \9777 , \3925 );
xor \U$9604 ( \9779 , \9774 , \9778 );
and \U$9605 ( \9780 , \1192 , \4581 );
and \U$9606 ( \9781 , \1333 , \4424 );
nor \U$9607 ( \9782 , \9780 , \9781 );
xnor \U$9608 ( \9783 , \9782 , \4377 );
xor \U$9609 ( \9784 , \9779 , \9783 );
and \U$9610 ( \9785 , \2521 , \2669 );
and \U$9611 ( \9786 , \2757 , \2538 );
nor \U$9612 ( \9787 , \9785 , \9786 );
xnor \U$9613 ( \9788 , \9787 , \2534 );
and \U$9614 ( \9789 , \2182 , \3103 );
and \U$9615 ( \9790 , \2366 , \2934 );
nor \U$9616 ( \9791 , \9789 , \9790 );
xnor \U$9617 ( \9792 , \9791 , \2839 );
xor \U$9618 ( \9793 , \9788 , \9792 );
and \U$9619 ( \9794 , \1948 , \3357 );
and \U$9620 ( \9795 , \2090 , \3255 );
nor \U$9621 ( \9796 , \9794 , \9795 );
xnor \U$9622 ( \9797 , \9796 , \3156 );
xor \U$9623 ( \9798 , \9793 , \9797 );
xor \U$9624 ( \9799 , \9784 , \9798 );
and \U$9625 ( \9800 , \3646 , \1824 );
and \U$9626 ( \9801 , \3736 , \1739 );
nor \U$9627 ( \9802 , \9800 , \9801 );
xnor \U$9628 ( \9803 , \9802 , \1697 );
and \U$9629 ( \9804 , \3143 , \2121 );
and \U$9630 ( \9805 , \3395 , \2008 );
nor \U$9631 ( \9806 , \9804 , \9805 );
xnor \U$9632 ( \9807 , \9806 , \1961 );
xor \U$9633 ( \9808 , \9803 , \9807 );
and \U$9634 ( \9809 , \2826 , \2400 );
and \U$9635 ( \9810 , \3037 , \2246 );
nor \U$9636 ( \9811 , \9809 , \9810 );
xnor \U$9637 ( \9812 , \9811 , \2195 );
xor \U$9638 ( \9813 , \9808 , \9812 );
xor \U$9639 ( \9814 , \9799 , \9813 );
xor \U$9640 ( \9815 , \9770 , \9814 );
and \U$9641 ( \9816 , \474 , \5011 );
and \U$9642 ( \9817 , \1147 , \4878 );
nor \U$9643 ( \9818 , \9816 , \9817 );
xnor \U$9644 ( \9819 , \9818 , \4762 );
and \U$9645 ( \9820 , \307 , \5485 );
and \U$9646 ( \9821 , \412 , \5275 );
nor \U$9647 ( \9822 , \9820 , \9821 );
xnor \U$9648 ( \9823 , \9822 , \5169 );
xor \U$9649 ( \9824 , \9819 , \9823 );
and \U$9650 ( \9825 , \185 , \5996 );
and \U$9651 ( \9826 , \261 , \5695 );
nor \U$9652 ( \9827 , \9825 , \9826 );
xnor \U$9653 ( \9828 , \9827 , \5687 );
xor \U$9654 ( \9829 , \9824 , \9828 );
and \U$9655 ( \9830 , \197 , \6401 );
and \U$9656 ( \9831 , \178 , \6143 );
nor \U$9657 ( \9832 , \9830 , \9831 );
xnor \U$9658 ( \9833 , \9832 , \6148 );
and \U$9659 ( \9834 , \217 , \7055 );
and \U$9660 ( \9835 , \189 , \6675 );
nor \U$9661 ( \9836 , \9834 , \9835 );
xnor \U$9662 ( \9837 , \9836 , \6680 );
xor \U$9663 ( \9838 , \9833 , \9837 );
and \U$9664 ( \9839 , \232 , \7489 );
and \U$9665 ( \9840 , \209 , \7137 );
nor \U$9666 ( \9841 , \9839 , \9840 );
xnor \U$9667 ( \9842 , \9841 , \7142 );
xor \U$9668 ( \9843 , \9838 , \9842 );
xor \U$9669 ( \9844 , \9829 , \9843 );
and \U$9670 ( \9845 , \247 , \8019 );
and \U$9671 ( \9846 , \224 , \7830 );
nor \U$9672 ( \9847 , \9845 , \9846 );
xnor \U$9673 ( \9848 , \9847 , \7713 );
and \U$9674 ( \9849 , \143 , \8540 );
and \U$9675 ( \9850 , \240 , \8292 );
nor \U$9676 ( \9851 , \9849 , \9850 );
xnor \U$9677 ( \9852 , \9851 , \8297 );
xor \U$9678 ( \9853 , \9848 , \9852 );
and \U$9679 ( \9854 , \158 , \9333 );
and \U$9680 ( \9855 , \134 , \9006 );
nor \U$9681 ( \9856 , \9854 , \9855 );
xnor \U$9682 ( \9857 , \9856 , \8848 );
xor \U$9683 ( \9858 , \9853 , \9857 );
xor \U$9684 ( \9859 , \9844 , \9858 );
xor \U$9685 ( \9860 , \9815 , \9859 );
xor \U$9686 ( \9861 , \9756 , \9860 );
xor \U$9687 ( \9862 , \9707 , \9861 );
and \U$9688 ( \9863 , \9494 , \9508 );
and \U$9689 ( \9864 , \9508 , \9523 );
and \U$9690 ( \9865 , \9494 , \9523 );
or \U$9691 ( \9866 , \9863 , \9864 , \9865 );
and \U$9692 ( \9867 , \9539 , \9553 );
and \U$9693 ( \9868 , \9553 , \9568 );
and \U$9694 ( \9869 , \9539 , \9568 );
or \U$9695 ( \9870 , \9867 , \9868 , \9869 );
xor \U$9696 ( \9871 , \9866 , \9870 );
and \U$9697 ( \9872 , \9624 , \9638 );
and \U$9698 ( \9873 , \9638 , \9647 );
and \U$9699 ( \9874 , \9624 , \9647 );
or \U$9700 ( \9875 , \9872 , \9873 , \9874 );
xor \U$9701 ( \9876 , \9871 , \9875 );
and \U$9702 ( \9877 , \9595 , \9599 );
and \U$9703 ( \9878 , \9599 , \9604 );
and \U$9704 ( \9879 , \9595 , \9604 );
or \U$9705 ( \9880 , \9877 , \9878 , \9879 );
and \U$9706 ( \9881 , \9580 , \9584 );
and \U$9707 ( \9882 , \9584 , \9589 );
and \U$9708 ( \9883 , \9580 , \9589 );
or \U$9709 ( \9884 , \9881 , \9882 , \9883 );
xor \U$9710 ( \9885 , \9880 , \9884 );
and \U$9711 ( \9886 , \9609 , \9613 );
and \U$9712 ( \9887 , \9613 , \9618 );
and \U$9713 ( \9888 , \9609 , \9618 );
or \U$9714 ( \9889 , \9886 , \9887 , \9888 );
xor \U$9715 ( \9890 , \9885 , \9889 );
xor \U$9716 ( \9891 , \9876 , \9890 );
and \U$9717 ( \9892 , \9448 , \9462 );
and \U$9718 ( \9893 , \9462 , \9479 );
and \U$9719 ( \9894 , \9448 , \9479 );
or \U$9720 ( \9895 , \9892 , \9893 , \9894 );
and \U$9721 ( \9896 , \9465 , \183 );
buf \U$9722 ( \9897 , RIb55f0d0_67);
and \U$9723 ( \9898 , \9897 , \180 );
nor \U$9724 ( \9899 , \9896 , \9898 );
xnor \U$9725 ( \9900 , \9899 , \179 );
and \U$9726 ( \9901 , \8835 , \195 );
and \U$9727 ( \9902 , \9169 , \193 );
nor \U$9728 ( \9903 , \9901 , \9902 );
xnor \U$9729 ( \9904 , \9903 , \202 );
xor \U$9730 ( \9905 , \9900 , \9904 );
and \U$9731 ( \9906 , \8349 , \215 );
and \U$9732 ( \9907 , \8652 , \213 );
nor \U$9733 ( \9908 , \9906 , \9907 );
xnor \U$9734 ( \9909 , \9908 , \222 );
xor \U$9735 ( \9910 , \9905 , \9909 );
xor \U$9736 ( \9911 , \9895 , \9910 );
and \U$9737 ( \9912 , \7700 , \230 );
and \U$9738 ( \9913 , \8057 , \228 );
nor \U$9739 ( \9914 , \9912 , \9913 );
xnor \U$9740 ( \9915 , \9914 , \237 );
and \U$9741 ( \9916 , \7231 , \245 );
and \U$9742 ( \9917 , \7556 , \243 );
nor \U$9743 ( \9918 , \9916 , \9917 );
xnor \U$9744 ( \9919 , \9918 , \252 );
xor \U$9745 ( \9920 , \9915 , \9919 );
and \U$9746 ( \9921 , \6790 , \141 );
and \U$9747 ( \9922 , \6945 , \139 );
nor \U$9748 ( \9923 , \9921 , \9922 );
xnor \U$9749 ( \9924 , \9923 , \148 );
xor \U$9750 ( \9925 , \9920 , \9924 );
and \U$9751 ( \9926 , \4749 , \1086 );
and \U$9752 ( \9927 , \4922 , \508 );
nor \U$9753 ( \9928 , \9926 , \9927 );
xnor \U$9754 ( \9929 , \9928 , \487 );
and \U$9755 ( \9930 , \4364 , \1301 );
and \U$9756 ( \9931 , \4654 , \1246 );
nor \U$9757 ( \9932 , \9930 , \9931 );
xnor \U$9758 ( \9933 , \9932 , \1205 );
xor \U$9759 ( \9934 , \9929 , \9933 );
and \U$9760 ( \9935 , \3912 , \1578 );
and \U$9761 ( \9936 , \4160 , \1431 );
nor \U$9762 ( \9937 , \9935 , \9936 );
xnor \U$9763 ( \9938 , \9937 , \1436 );
xor \U$9764 ( \9939 , \9934 , \9938 );
xor \U$9765 ( \9940 , \9925 , \9939 );
and \U$9766 ( \9941 , \6281 , \156 );
and \U$9767 ( \9942 , \6514 , \154 );
nor \U$9768 ( \9943 , \9941 , \9942 );
xnor \U$9769 ( \9944 , \9943 , \163 );
and \U$9770 ( \9945 , \5674 , \296 );
and \U$9771 ( \9946 , \6030 , \168 );
nor \U$9772 ( \9947 , \9945 , \9946 );
xnor \U$9773 ( \9948 , \9947 , \173 );
xor \U$9774 ( \9949 , \9944 , \9948 );
and \U$9775 ( \9950 , \5156 , \438 );
and \U$9776 ( \9951 , \5469 , \336 );
nor \U$9777 ( \9952 , \9950 , \9951 );
xnor \U$9778 ( \9953 , \9952 , \320 );
xor \U$9779 ( \9954 , \9949 , \9953 );
xor \U$9780 ( \9955 , \9940 , \9954 );
xor \U$9781 ( \9956 , \9911 , \9955 );
xor \U$9782 ( \9957 , \9891 , \9956 );
xor \U$9783 ( \9958 , \9862 , \9957 );
xor \U$9784 ( \9959 , \9693 , \9958 );
xor \U$9785 ( \9960 , \9684 , \9959 );
xor \U$9786 ( \9961 , \9665 , \9960 );
and \U$9787 ( \9962 , \9357 , \9381 );
and \U$9788 ( \9963 , \9381 , \9652 );
and \U$9789 ( \9964 , \9357 , \9652 );
or \U$9790 ( \9965 , \9962 , \9963 , \9964 );
xor \U$9791 ( \9966 , \9961 , \9965 );
and \U$9792 ( \9967 , \9653 , \9654 );
and \U$9793 ( \9968 , \9655 , \9658 );
or \U$9794 ( \9969 , \9967 , \9968 );
xor \U$9795 ( \9970 , \9966 , \9969 );
buf g5521_GF_PartitionCandidate( \9971_nG5521 , \9970 );
buf \U$9796 ( \9972 , \9971_nG5521 );
and \U$9797 ( \9973 , \9669 , \9683 );
and \U$9798 ( \9974 , \9683 , \9959 );
and \U$9799 ( \9975 , \9669 , \9959 );
or \U$9800 ( \9976 , \9973 , \9974 , \9975 );
and \U$9801 ( \9977 , \9688 , \9692 );
and \U$9802 ( \9978 , \9692 , \9958 );
and \U$9803 ( \9979 , \9688 , \9958 );
or \U$9804 ( \9980 , \9977 , \9978 , \9979 );
and \U$9805 ( \9981 , \9673 , \9677 );
and \U$9806 ( \9982 , \9677 , \9682 );
and \U$9807 ( \9983 , \9673 , \9682 );
or \U$9808 ( \9984 , \9981 , \9982 , \9983 );
and \U$9809 ( \9985 , \9707 , \9861 );
and \U$9810 ( \9986 , \9861 , \9957 );
and \U$9811 ( \9987 , \9707 , \9957 );
or \U$9812 ( \9988 , \9985 , \9986 , \9987 );
xor \U$9813 ( \9989 , \9984 , \9988 );
and \U$9814 ( \9990 , \9725 , \9739 );
and \U$9815 ( \9991 , \9739 , \9754 );
and \U$9816 ( \9992 , \9725 , \9754 );
or \U$9817 ( \9993 , \9990 , \9991 , \9992 );
and \U$9818 ( \9994 , \9770 , \9814 );
and \U$9819 ( \9995 , \9814 , \9859 );
and \U$9820 ( \9996 , \9770 , \9859 );
or \U$9821 ( \9997 , \9994 , \9995 , \9996 );
xor \U$9822 ( \9998 , \9993 , \9997 );
and \U$9823 ( \9999 , \9929 , \9933 );
and \U$9824 ( \10000 , \9933 , \9938 );
and \U$9825 ( \10001 , \9929 , \9938 );
or \U$9826 ( \10002 , \9999 , \10000 , \10001 );
and \U$9827 ( \10003 , \9788 , \9792 );
and \U$9828 ( \10004 , \9792 , \9797 );
and \U$9829 ( \10005 , \9788 , \9797 );
or \U$9830 ( \10006 , \10003 , \10004 , \10005 );
xor \U$9831 ( \10007 , \10002 , \10006 );
and \U$9832 ( \10008 , \9803 , \9807 );
and \U$9833 ( \10009 , \9807 , \9812 );
and \U$9834 ( \10010 , \9803 , \9812 );
or \U$9835 ( \10011 , \10008 , \10009 , \10010 );
xor \U$9836 ( \10012 , \10007 , \10011 );
xor \U$9837 ( \10013 , \9998 , \10012 );
xor \U$9838 ( \10014 , \9989 , \10013 );
xor \U$9839 ( \10015 , \9980 , \10014 );
and \U$9840 ( \10016 , \9866 , \9870 );
and \U$9841 ( \10017 , \9870 , \9875 );
and \U$9842 ( \10018 , \9866 , \9875 );
or \U$9843 ( \10019 , \10016 , \10017 , \10018 );
and \U$9844 ( \10020 , \9880 , \9884 );
and \U$9845 ( \10021 , \9884 , \9889 );
and \U$9846 ( \10022 , \9880 , \9889 );
or \U$9847 ( \10023 , \10020 , \10021 , \10022 );
xor \U$9848 ( \10024 , \10019 , \10023 );
and \U$9849 ( \10025 , \9895 , \9910 );
and \U$9850 ( \10026 , \9910 , \9955 );
and \U$9851 ( \10027 , \9895 , \9955 );
or \U$9852 ( \10028 , \10025 , \10026 , \10027 );
xor \U$9853 ( \10029 , \10024 , \10028 );
and \U$9854 ( \10030 , \9697 , \9701 );
and \U$9855 ( \10031 , \9701 , \9706 );
and \U$9856 ( \10032 , \9697 , \9706 );
or \U$9857 ( \10033 , \10030 , \10031 , \10032 );
and \U$9858 ( \10034 , \9711 , \9755 );
and \U$9859 ( \10035 , \9755 , \9860 );
and \U$9860 ( \10036 , \9711 , \9860 );
or \U$9861 ( \10037 , \10034 , \10035 , \10036 );
xor \U$9862 ( \10038 , \10033 , \10037 );
and \U$9863 ( \10039 , \9876 , \9890 );
and \U$9864 ( \10040 , \9890 , \9956 );
and \U$9865 ( \10041 , \9876 , \9956 );
or \U$9866 ( \10042 , \10039 , \10040 , \10041 );
xor \U$9867 ( \10043 , \10038 , \10042 );
xor \U$9868 ( \10044 , \10029 , \10043 );
and \U$9869 ( \10045 , \9715 , \9719 );
and \U$9870 ( \10046 , \9719 , \9724 );
and \U$9871 ( \10047 , \9715 , \9724 );
or \U$9872 ( \10048 , \10045 , \10046 , \10047 );
and \U$9873 ( \10049 , \9729 , \9733 );
and \U$9874 ( \10050 , \9733 , \9738 );
and \U$9875 ( \10051 , \9729 , \9738 );
or \U$9876 ( \10052 , \10049 , \10050 , \10051 );
xor \U$9877 ( \10053 , \10048 , \10052 );
and \U$9878 ( \10054 , \9744 , \9748 );
and \U$9879 ( \10055 , \9748 , \9753 );
and \U$9880 ( \10056 , \9744 , \9753 );
or \U$9881 ( \10057 , \10054 , \10055 , \10056 );
xor \U$9882 ( \10058 , \10053 , \10057 );
and \U$9883 ( \10059 , \9760 , \9761 );
and \U$9884 ( \10060 , \9761 , \9769 );
and \U$9885 ( \10061 , \9760 , \9769 );
or \U$9886 ( \10062 , \10059 , \10060 , \10061 );
and \U$9887 ( \10063 , \9784 , \9798 );
and \U$9888 ( \10064 , \9798 , \9813 );
and \U$9889 ( \10065 , \9784 , \9813 );
or \U$9890 ( \10066 , \10063 , \10064 , \10065 );
xor \U$9891 ( \10067 , \10062 , \10066 );
and \U$9892 ( \10068 , \9829 , \9843 );
and \U$9893 ( \10069 , \9843 , \9858 );
and \U$9894 ( \10070 , \9829 , \9858 );
or \U$9895 ( \10071 , \10068 , \10069 , \10070 );
xor \U$9896 ( \10072 , \10067 , \10071 );
xor \U$9897 ( \10073 , \10058 , \10072 );
and \U$9898 ( \10074 , \9915 , \9919 );
and \U$9899 ( \10075 , \9919 , \9924 );
and \U$9900 ( \10076 , \9915 , \9924 );
or \U$9901 ( \10077 , \10074 , \10075 , \10076 );
and \U$9902 ( \10078 , \9900 , \9904 );
and \U$9903 ( \10079 , \9904 , \9909 );
and \U$9904 ( \10080 , \9900 , \9909 );
or \U$9905 ( \10081 , \10078 , \10079 , \10080 );
xor \U$9906 ( \10082 , \10077 , \10081 );
and \U$9907 ( \10083 , \9944 , \9948 );
and \U$9908 ( \10084 , \9948 , \9953 );
and \U$9909 ( \10085 , \9944 , \9953 );
or \U$9910 ( \10086 , \10083 , \10084 , \10085 );
xor \U$9911 ( \10087 , \10082 , \10086 );
and \U$9912 ( \10088 , \9819 , \9823 );
and \U$9913 ( \10089 , \9823 , \9828 );
and \U$9914 ( \10090 , \9819 , \9828 );
or \U$9915 ( \10091 , \10088 , \10089 , \10090 );
and \U$9916 ( \10092 , \9833 , \9837 );
and \U$9917 ( \10093 , \9837 , \9842 );
and \U$9918 ( \10094 , \9833 , \9842 );
or \U$9919 ( \10095 , \10092 , \10093 , \10094 );
xor \U$9920 ( \10096 , \10091 , \10095 );
and \U$9921 ( \10097 , \9774 , \9778 );
and \U$9922 ( \10098 , \9778 , \9783 );
and \U$9923 ( \10099 , \9774 , \9783 );
or \U$9924 ( \10100 , \10097 , \10098 , \10099 );
xor \U$9925 ( \10101 , \10096 , \10100 );
and \U$9926 ( \10102 , \9848 , \9852 );
and \U$9927 ( \10103 , \9852 , \9857 );
and \U$9928 ( \10104 , \9848 , \9857 );
or \U$9929 ( \10105 , \10102 , \10103 , \10104 );
and \U$9930 ( \10106 , \134 , \9333 );
and \U$9931 ( \10107 , \143 , \9006 );
nor \U$9932 ( \10108 , \10106 , \10107 );
xnor \U$9933 ( \10109 , \10108 , \8848 );
and \U$9934 ( \10110 , \150 , \9765 );
and \U$9935 ( \10111 , \158 , \9644 );
nor \U$9936 ( \10112 , \10110 , \10111 );
xnor \U$9937 ( \10113 , \10112 , \9478 );
xor \U$9938 ( \10114 , \10109 , \10113 );
buf \U$9939 ( \10115 , RIb560f48_2);
xor \U$9940 ( \10116 , \10115 , \9474 );
nand \U$9941 ( \10117 , \166 , \10116 );
buf \U$9942 ( \10118 , RIb560fc0_1);
and \U$9943 ( \10119 , \10115 , \9474 );
not \U$9944 ( \10120 , \10119 );
and \U$9945 ( \10121 , \10118 , \10120 );
xnor \U$9946 ( \10122 , \10117 , \10121 );
xor \U$9947 ( \10123 , \10114 , \10122 );
xor \U$9948 ( \10124 , \10105 , \10123 );
and \U$9949 ( \10125 , \209 , \7489 );
and \U$9950 ( \10126 , \217 , \7137 );
nor \U$9951 ( \10127 , \10125 , \10126 );
xnor \U$9952 ( \10128 , \10127 , \7142 );
and \U$9953 ( \10129 , \224 , \8019 );
and \U$9954 ( \10130 , \232 , \7830 );
nor \U$9955 ( \10131 , \10129 , \10130 );
xnor \U$9956 ( \10132 , \10131 , \7713 );
xor \U$9957 ( \10133 , \10128 , \10132 );
and \U$9958 ( \10134 , \240 , \8540 );
and \U$9959 ( \10135 , \247 , \8292 );
nor \U$9960 ( \10136 , \10134 , \10135 );
xnor \U$9961 ( \10137 , \10136 , \8297 );
xor \U$9962 ( \10138 , \10133 , \10137 );
xor \U$9963 ( \10139 , \10124 , \10138 );
xor \U$9964 ( \10140 , \10101 , \10139 );
and \U$9965 ( \10141 , \1333 , \4581 );
and \U$9966 ( \10142 , \1484 , \4424 );
nor \U$9967 ( \10143 , \10141 , \10142 );
xnor \U$9968 ( \10144 , \10143 , \4377 );
and \U$9969 ( \10145 , \1147 , \5011 );
and \U$9970 ( \10146 , \1192 , \4878 );
nor \U$9971 ( \10147 , \10145 , \10146 );
xnor \U$9972 ( \10148 , \10147 , \4762 );
xor \U$9973 ( \10149 , \10144 , \10148 );
and \U$9974 ( \10150 , \412 , \5485 );
and \U$9975 ( \10151 , \474 , \5275 );
nor \U$9976 ( \10152 , \10150 , \10151 );
xnor \U$9977 ( \10153 , \10152 , \5169 );
xor \U$9978 ( \10154 , \10149 , \10153 );
and \U$9979 ( \10155 , \2090 , \3357 );
and \U$9980 ( \10156 , \2182 , \3255 );
nor \U$9981 ( \10157 , \10155 , \10156 );
xnor \U$9982 ( \10158 , \10157 , \3156 );
and \U$9983 ( \10159 , \1802 , \3813 );
and \U$9984 ( \10160 , \1948 , \3557 );
nor \U$9985 ( \10161 , \10159 , \10160 );
xnor \U$9986 ( \10162 , \10161 , \3562 );
xor \U$9987 ( \10163 , \10158 , \10162 );
and \U$9988 ( \10164 , \1601 , \4132 );
and \U$9989 ( \10165 , \1684 , \4012 );
nor \U$9990 ( \10166 , \10164 , \10165 );
xnor \U$9991 ( \10167 , \10166 , \3925 );
xor \U$9992 ( \10168 , \10163 , \10167 );
xor \U$9993 ( \10169 , \10154 , \10168 );
and \U$9994 ( \10170 , \261 , \5996 );
and \U$9995 ( \10171 , \307 , \5695 );
nor \U$9996 ( \10172 , \10170 , \10171 );
xnor \U$9997 ( \10173 , \10172 , \5687 );
and \U$9998 ( \10174 , \178 , \6401 );
and \U$9999 ( \10175 , \185 , \6143 );
nor \U$10000 ( \10176 , \10174 , \10175 );
xnor \U$10001 ( \10177 , \10176 , \6148 );
xor \U$10002 ( \10178 , \10173 , \10177 );
and \U$10003 ( \10179 , \189 , \7055 );
and \U$10004 ( \10180 , \197 , \6675 );
nor \U$10005 ( \10181 , \10179 , \10180 );
xnor \U$10006 ( \10182 , \10181 , \6680 );
xor \U$10007 ( \10183 , \10178 , \10182 );
xor \U$10008 ( \10184 , \10169 , \10183 );
xor \U$10009 ( \10185 , \10140 , \10184 );
xor \U$10010 ( \10186 , \10087 , \10185 );
and \U$10011 ( \10187 , \9925 , \9939 );
and \U$10012 ( \10188 , \9939 , \9954 );
and \U$10013 ( \10189 , \9925 , \9954 );
or \U$10014 ( \10190 , \10187 , \10188 , \10189 );
and \U$10015 ( \10191 , \6945 , \141 );
and \U$10016 ( \10192 , \7231 , \139 );
nor \U$10017 ( \10193 , \10191 , \10192 );
xnor \U$10018 ( \10194 , \10193 , \148 );
and \U$10019 ( \10195 , \6514 , \156 );
and \U$10020 ( \10196 , \6790 , \154 );
nor \U$10021 ( \10197 , \10195 , \10196 );
xnor \U$10022 ( \10198 , \10197 , \163 );
xor \U$10023 ( \10199 , \10194 , \10198 );
and \U$10024 ( \10200 , \6030 , \296 );
and \U$10025 ( \10201 , \6281 , \168 );
nor \U$10026 ( \10202 , \10200 , \10201 );
xnor \U$10027 ( \10203 , \10202 , \173 );
xor \U$10028 ( \10204 , \10199 , \10203 );
and \U$10029 ( \10205 , \9897 , \183 );
buf \U$10030 ( \10206 , RIb55f148_66);
and \U$10031 ( \10207 , \10206 , \180 );
nor \U$10032 ( \10208 , \10205 , \10207 );
xnor \U$10033 ( \10209 , \10208 , \179 );
and \U$10034 ( \10210 , \9169 , \195 );
and \U$10035 ( \10211 , \9465 , \193 );
nor \U$10036 ( \10212 , \10210 , \10211 );
xnor \U$10037 ( \10213 , \10212 , \202 );
xor \U$10038 ( \10214 , \10209 , \10213 );
xor \U$10039 ( \10215 , \10214 , \10121 );
xor \U$10040 ( \10216 , \10204 , \10215 );
and \U$10041 ( \10217 , \8652 , \215 );
and \U$10042 ( \10218 , \8835 , \213 );
nor \U$10043 ( \10219 , \10217 , \10218 );
xnor \U$10044 ( \10220 , \10219 , \222 );
and \U$10045 ( \10221 , \8057 , \230 );
and \U$10046 ( \10222 , \8349 , \228 );
nor \U$10047 ( \10223 , \10221 , \10222 );
xnor \U$10048 ( \10224 , \10223 , \237 );
xor \U$10049 ( \10225 , \10220 , \10224 );
and \U$10050 ( \10226 , \7556 , \245 );
and \U$10051 ( \10227 , \7700 , \243 );
nor \U$10052 ( \10228 , \10226 , \10227 );
xnor \U$10053 ( \10229 , \10228 , \252 );
xor \U$10054 ( \10230 , \10225 , \10229 );
xor \U$10055 ( \10231 , \10216 , \10230 );
xor \U$10056 ( \10232 , \10190 , \10231 );
and \U$10057 ( \10233 , \4160 , \1578 );
and \U$10058 ( \10234 , \4364 , \1431 );
nor \U$10059 ( \10235 , \10233 , \10234 );
xnor \U$10060 ( \10236 , \10235 , \1436 );
and \U$10061 ( \10237 , \3736 , \1824 );
and \U$10062 ( \10238 , \3912 , \1739 );
nor \U$10063 ( \10239 , \10237 , \10238 );
xnor \U$10064 ( \10240 , \10239 , \1697 );
xor \U$10065 ( \10241 , \10236 , \10240 );
and \U$10066 ( \10242 , \3395 , \2121 );
and \U$10067 ( \10243 , \3646 , \2008 );
nor \U$10068 ( \10244 , \10242 , \10243 );
xnor \U$10069 ( \10245 , \10244 , \1961 );
xor \U$10070 ( \10246 , \10241 , \10245 );
and \U$10071 ( \10247 , \5469 , \438 );
and \U$10072 ( \10248 , \5674 , \336 );
nor \U$10073 ( \10249 , \10247 , \10248 );
xnor \U$10074 ( \10250 , \10249 , \320 );
and \U$10075 ( \10251 , \4922 , \1086 );
and \U$10076 ( \10252 , \5156 , \508 );
nor \U$10077 ( \10253 , \10251 , \10252 );
xnor \U$10078 ( \10254 , \10253 , \487 );
xor \U$10079 ( \10255 , \10250 , \10254 );
and \U$10080 ( \10256 , \4654 , \1301 );
and \U$10081 ( \10257 , \4749 , \1246 );
nor \U$10082 ( \10258 , \10256 , \10257 );
xnor \U$10083 ( \10259 , \10258 , \1205 );
xor \U$10084 ( \10260 , \10255 , \10259 );
xor \U$10085 ( \10261 , \10246 , \10260 );
and \U$10086 ( \10262 , \3037 , \2400 );
and \U$10087 ( \10263 , \3143 , \2246 );
nor \U$10088 ( \10264 , \10262 , \10263 );
xnor \U$10089 ( \10265 , \10264 , \2195 );
and \U$10090 ( \10266 , \2757 , \2669 );
and \U$10091 ( \10267 , \2826 , \2538 );
nor \U$10092 ( \10268 , \10266 , \10267 );
xnor \U$10093 ( \10269 , \10268 , \2534 );
xor \U$10094 ( \10270 , \10265 , \10269 );
and \U$10095 ( \10271 , \2366 , \3103 );
and \U$10096 ( \10272 , \2521 , \2934 );
nor \U$10097 ( \10273 , \10271 , \10272 );
xnor \U$10098 ( \10274 , \10273 , \2839 );
xor \U$10099 ( \10275 , \10270 , \10274 );
xor \U$10100 ( \10276 , \10261 , \10275 );
xor \U$10101 ( \10277 , \10232 , \10276 );
xor \U$10102 ( \10278 , \10186 , \10277 );
xor \U$10103 ( \10279 , \10073 , \10278 );
xor \U$10104 ( \10280 , \10044 , \10279 );
xor \U$10105 ( \10281 , \10015 , \10280 );
xor \U$10106 ( \10282 , \9976 , \10281 );
and \U$10107 ( \10283 , \9665 , \9960 );
xor \U$10108 ( \10284 , \10282 , \10283 );
and \U$10109 ( \10285 , \9961 , \9965 );
and \U$10110 ( \10286 , \9966 , \9969 );
or \U$10111 ( \10287 , \10285 , \10286 );
xor \U$10112 ( \10288 , \10284 , \10287 );
buf g551f_GF_PartitionCandidate( \10289_nG551f , \10288 );
buf \U$10113 ( \10290 , \10289_nG551f );
and \U$10114 ( \10291 , \9980 , \10014 );
and \U$10115 ( \10292 , \10014 , \10280 );
and \U$10116 ( \10293 , \9980 , \10280 );
or \U$10117 ( \10294 , \10291 , \10292 , \10293 );
and \U$10118 ( \10295 , \9984 , \9988 );
and \U$10119 ( \10296 , \9988 , \10013 );
and \U$10120 ( \10297 , \9984 , \10013 );
or \U$10121 ( \10298 , \10295 , \10296 , \10297 );
and \U$10122 ( \10299 , \10029 , \10043 );
and \U$10123 ( \10300 , \10043 , \10279 );
and \U$10124 ( \10301 , \10029 , \10279 );
or \U$10125 ( \10302 , \10299 , \10300 , \10301 );
xor \U$10126 ( \10303 , \10298 , \10302 );
and \U$10127 ( \10304 , \10019 , \10023 );
and \U$10128 ( \10305 , \10023 , \10028 );
and \U$10129 ( \10306 , \10019 , \10028 );
or \U$10130 ( \10307 , \10304 , \10305 , \10306 );
and \U$10131 ( \10308 , \9993 , \9997 );
and \U$10132 ( \10309 , \9997 , \10012 );
and \U$10133 ( \10310 , \9993 , \10012 );
or \U$10134 ( \10311 , \10308 , \10309 , \10310 );
xor \U$10135 ( \10312 , \10307 , \10311 );
and \U$10136 ( \10313 , \10087 , \10185 );
and \U$10137 ( \10314 , \10185 , \10277 );
and \U$10138 ( \10315 , \10087 , \10277 );
or \U$10139 ( \10316 , \10313 , \10314 , \10315 );
xor \U$10140 ( \10317 , \10312 , \10316 );
xor \U$10141 ( \10318 , \10303 , \10317 );
xor \U$10142 ( \10319 , \10294 , \10318 );
and \U$10143 ( \10320 , \10033 , \10037 );
and \U$10144 ( \10321 , \10037 , \10042 );
and \U$10145 ( \10322 , \10033 , \10042 );
or \U$10146 ( \10323 , \10320 , \10321 , \10322 );
and \U$10147 ( \10324 , \10058 , \10072 );
and \U$10148 ( \10325 , \10072 , \10278 );
and \U$10149 ( \10326 , \10058 , \10278 );
or \U$10150 ( \10327 , \10324 , \10325 , \10326 );
xor \U$10151 ( \10328 , \10323 , \10327 );
and \U$10152 ( \10329 , \10048 , \10052 );
and \U$10153 ( \10330 , \10052 , \10057 );
and \U$10154 ( \10331 , \10048 , \10057 );
or \U$10155 ( \10332 , \10329 , \10330 , \10331 );
and \U$10156 ( \10333 , \10062 , \10066 );
and \U$10157 ( \10334 , \10066 , \10071 );
and \U$10158 ( \10335 , \10062 , \10071 );
or \U$10159 ( \10336 , \10333 , \10334 , \10335 );
xor \U$10160 ( \10337 , \10332 , \10336 );
and \U$10161 ( \10338 , \10190 , \10231 );
and \U$10162 ( \10339 , \10231 , \10276 );
and \U$10163 ( \10340 , \10190 , \10276 );
or \U$10164 ( \10341 , \10338 , \10339 , \10340 );
xor \U$10165 ( \10342 , \10337 , \10341 );
and \U$10166 ( \10343 , \10101 , \10139 );
and \U$10167 ( \10344 , \10139 , \10184 );
and \U$10168 ( \10345 , \10101 , \10184 );
or \U$10169 ( \10346 , \10343 , \10344 , \10345 );
and \U$10170 ( \10347 , \10144 , \10148 );
and \U$10171 ( \10348 , \10148 , \10153 );
and \U$10172 ( \10349 , \10144 , \10153 );
or \U$10173 ( \10350 , \10347 , \10348 , \10349 );
and \U$10174 ( \10351 , \10158 , \10162 );
and \U$10175 ( \10352 , \10162 , \10167 );
and \U$10176 ( \10353 , \10158 , \10167 );
or \U$10177 ( \10354 , \10351 , \10352 , \10353 );
xor \U$10178 ( \10355 , \10350 , \10354 );
and \U$10179 ( \10356 , \10173 , \10177 );
and \U$10180 ( \10357 , \10177 , \10182 );
and \U$10181 ( \10358 , \10173 , \10182 );
or \U$10182 ( \10359 , \10356 , \10357 , \10358 );
xor \U$10183 ( \10360 , \10355 , \10359 );
and \U$10184 ( \10361 , \10194 , \10198 );
and \U$10185 ( \10362 , \10198 , \10203 );
and \U$10186 ( \10363 , \10194 , \10203 );
or \U$10187 ( \10364 , \10361 , \10362 , \10363 );
and \U$10188 ( \10365 , \10209 , \10213 );
and \U$10189 ( \10366 , \10213 , \10121 );
and \U$10190 ( \10367 , \10209 , \10121 );
or \U$10191 ( \10368 , \10365 , \10366 , \10367 );
xor \U$10192 ( \10369 , \10364 , \10368 );
and \U$10193 ( \10370 , \10220 , \10224 );
and \U$10194 ( \10371 , \10224 , \10229 );
and \U$10195 ( \10372 , \10220 , \10229 );
or \U$10196 ( \10373 , \10370 , \10371 , \10372 );
xor \U$10197 ( \10374 , \10369 , \10373 );
xor \U$10198 ( \10375 , \10360 , \10374 );
and \U$10199 ( \10376 , \10236 , \10240 );
and \U$10200 ( \10377 , \10240 , \10245 );
and \U$10201 ( \10378 , \10236 , \10245 );
or \U$10202 ( \10379 , \10376 , \10377 , \10378 );
and \U$10203 ( \10380 , \10250 , \10254 );
and \U$10204 ( \10381 , \10254 , \10259 );
and \U$10205 ( \10382 , \10250 , \10259 );
or \U$10206 ( \10383 , \10380 , \10381 , \10382 );
xor \U$10207 ( \10384 , \10379 , \10383 );
and \U$10208 ( \10385 , \10265 , \10269 );
and \U$10209 ( \10386 , \10269 , \10274 );
and \U$10210 ( \10387 , \10265 , \10274 );
or \U$10211 ( \10388 , \10385 , \10386 , \10387 );
xor \U$10212 ( \10389 , \10384 , \10388 );
xor \U$10213 ( \10390 , \10375 , \10389 );
xor \U$10214 ( \10391 , \10346 , \10390 );
and \U$10215 ( \10392 , \10109 , \10113 );
and \U$10216 ( \10393 , \10113 , \10122 );
and \U$10217 ( \10394 , \10109 , \10122 );
or \U$10218 ( \10395 , \10392 , \10393 , \10394 );
and \U$10219 ( \10396 , \10128 , \10132 );
and \U$10220 ( \10397 , \10132 , \10137 );
and \U$10221 ( \10398 , \10128 , \10137 );
or \U$10222 ( \10399 , \10396 , \10397 , \10398 );
xor \U$10223 ( \10400 , \10395 , \10399 );
and \U$10224 ( \10401 , \158 , \9765 );
and \U$10225 ( \10402 , \134 , \9644 );
nor \U$10226 ( \10403 , \10401 , \10402 );
xnor \U$10227 ( \10404 , \10403 , \9478 );
xor \U$10228 ( \10405 , \10400 , \10404 );
xor \U$10229 ( \10406 , \10118 , \10115 );
not \U$10230 ( \10407 , \10116 );
and \U$10231 ( \10408 , \10406 , \10407 );
and \U$10232 ( \10409 , \166 , \10408 );
and \U$10233 ( \10410 , \150 , \10116 );
nor \U$10234 ( \10411 , \10409 , \10410 );
xnor \U$10235 ( \10412 , \10411 , \10121 );
and \U$10236 ( \10413 , \185 , \6401 );
and \U$10237 ( \10414 , \261 , \6143 );
nor \U$10238 ( \10415 , \10413 , \10414 );
xnor \U$10239 ( \10416 , \10415 , \6148 );
and \U$10240 ( \10417 , \197 , \7055 );
and \U$10241 ( \10418 , \178 , \6675 );
nor \U$10242 ( \10419 , \10417 , \10418 );
xnor \U$10243 ( \10420 , \10419 , \6680 );
xor \U$10244 ( \10421 , \10416 , \10420 );
and \U$10245 ( \10422 , \217 , \7489 );
and \U$10246 ( \10423 , \189 , \7137 );
nor \U$10247 ( \10424 , \10422 , \10423 );
xnor \U$10248 ( \10425 , \10424 , \7142 );
xor \U$10249 ( \10426 , \10421 , \10425 );
xor \U$10250 ( \10427 , \10412 , \10426 );
and \U$10251 ( \10428 , \232 , \8019 );
and \U$10252 ( \10429 , \209 , \7830 );
nor \U$10253 ( \10430 , \10428 , \10429 );
xnor \U$10254 ( \10431 , \10430 , \7713 );
and \U$10255 ( \10432 , \247 , \8540 );
and \U$10256 ( \10433 , \224 , \8292 );
nor \U$10257 ( \10434 , \10432 , \10433 );
xnor \U$10258 ( \10435 , \10434 , \8297 );
xor \U$10259 ( \10436 , \10431 , \10435 );
and \U$10260 ( \10437 , \143 , \9333 );
and \U$10261 ( \10438 , \240 , \9006 );
nor \U$10262 ( \10439 , \10437 , \10438 );
xnor \U$10263 ( \10440 , \10439 , \8848 );
xor \U$10264 ( \10441 , \10436 , \10440 );
xor \U$10265 ( \10442 , \10427 , \10441 );
xor \U$10266 ( \10443 , \10405 , \10442 );
and \U$10267 ( \10444 , \1192 , \5011 );
and \U$10268 ( \10445 , \1333 , \4878 );
nor \U$10269 ( \10446 , \10444 , \10445 );
xnor \U$10270 ( \10447 , \10446 , \4762 );
and \U$10271 ( \10448 , \474 , \5485 );
and \U$10272 ( \10449 , \1147 , \5275 );
nor \U$10273 ( \10450 , \10448 , \10449 );
xnor \U$10274 ( \10451 , \10450 , \5169 );
xor \U$10275 ( \10452 , \10447 , \10451 );
and \U$10276 ( \10453 , \307 , \5996 );
and \U$10277 ( \10454 , \412 , \5695 );
nor \U$10278 ( \10455 , \10453 , \10454 );
xnor \U$10279 ( \10456 , \10455 , \5687 );
xor \U$10280 ( \10457 , \10452 , \10456 );
and \U$10281 ( \10458 , \1948 , \3813 );
and \U$10282 ( \10459 , \2090 , \3557 );
nor \U$10283 ( \10460 , \10458 , \10459 );
xnor \U$10284 ( \10461 , \10460 , \3562 );
and \U$10285 ( \10462 , \1684 , \4132 );
and \U$10286 ( \10463 , \1802 , \4012 );
nor \U$10287 ( \10464 , \10462 , \10463 );
xnor \U$10288 ( \10465 , \10464 , \3925 );
xor \U$10289 ( \10466 , \10461 , \10465 );
and \U$10290 ( \10467 , \1484 , \4581 );
and \U$10291 ( \10468 , \1601 , \4424 );
nor \U$10292 ( \10469 , \10467 , \10468 );
xnor \U$10293 ( \10470 , \10469 , \4377 );
xor \U$10294 ( \10471 , \10466 , \10470 );
xor \U$10295 ( \10472 , \10457 , \10471 );
and \U$10296 ( \10473 , \2826 , \2669 );
and \U$10297 ( \10474 , \3037 , \2538 );
nor \U$10298 ( \10475 , \10473 , \10474 );
xnor \U$10299 ( \10476 , \10475 , \2534 );
and \U$10300 ( \10477 , \2521 , \3103 );
and \U$10301 ( \10478 , \2757 , \2934 );
nor \U$10302 ( \10479 , \10477 , \10478 );
xnor \U$10303 ( \10480 , \10479 , \2839 );
xor \U$10304 ( \10481 , \10476 , \10480 );
and \U$10305 ( \10482 , \2182 , \3357 );
and \U$10306 ( \10483 , \2366 , \3255 );
nor \U$10307 ( \10484 , \10482 , \10483 );
xnor \U$10308 ( \10485 , \10484 , \3156 );
xor \U$10309 ( \10486 , \10481 , \10485 );
xor \U$10310 ( \10487 , \10472 , \10486 );
xor \U$10311 ( \10488 , \10443 , \10487 );
xor \U$10312 ( \10489 , \10391 , \10488 );
xor \U$10313 ( \10490 , \10342 , \10489 );
and \U$10314 ( \10491 , \10077 , \10081 );
and \U$10315 ( \10492 , \10081 , \10086 );
and \U$10316 ( \10493 , \10077 , \10086 );
or \U$10317 ( \10494 , \10491 , \10492 , \10493 );
and \U$10318 ( \10495 , \10091 , \10095 );
and \U$10319 ( \10496 , \10095 , \10100 );
and \U$10320 ( \10497 , \10091 , \10100 );
or \U$10321 ( \10498 , \10495 , \10496 , \10497 );
xor \U$10322 ( \10499 , \10494 , \10498 );
and \U$10323 ( \10500 , \10002 , \10006 );
and \U$10324 ( \10501 , \10006 , \10011 );
and \U$10325 ( \10502 , \10002 , \10011 );
or \U$10326 ( \10503 , \10500 , \10501 , \10502 );
xor \U$10327 ( \10504 , \10499 , \10503 );
and \U$10328 ( \10505 , \10246 , \10260 );
and \U$10329 ( \10506 , \10260 , \10275 );
and \U$10330 ( \10507 , \10246 , \10275 );
or \U$10331 ( \10508 , \10505 , \10506 , \10507 );
and \U$10332 ( \10509 , \10105 , \10123 );
and \U$10333 ( \10510 , \10123 , \10138 );
and \U$10334 ( \10511 , \10105 , \10138 );
or \U$10335 ( \10512 , \10509 , \10510 , \10511 );
xor \U$10336 ( \10513 , \10508 , \10512 );
and \U$10337 ( \10514 , \10154 , \10168 );
and \U$10338 ( \10515 , \10168 , \10183 );
and \U$10339 ( \10516 , \10154 , \10183 );
or \U$10340 ( \10517 , \10514 , \10515 , \10516 );
xor \U$10341 ( \10518 , \10513 , \10517 );
xor \U$10342 ( \10519 , \10504 , \10518 );
and \U$10343 ( \10520 , \10204 , \10215 );
and \U$10344 ( \10521 , \10215 , \10230 );
and \U$10345 ( \10522 , \10204 , \10230 );
or \U$10346 ( \10523 , \10520 , \10521 , \10522 );
and \U$10347 ( \10524 , \3912 , \1824 );
and \U$10348 ( \10525 , \4160 , \1739 );
nor \U$10349 ( \10526 , \10524 , \10525 );
xnor \U$10350 ( \10527 , \10526 , \1697 );
and \U$10351 ( \10528 , \3646 , \2121 );
and \U$10352 ( \10529 , \3736 , \2008 );
nor \U$10353 ( \10530 , \10528 , \10529 );
xnor \U$10354 ( \10531 , \10530 , \1961 );
xor \U$10355 ( \10532 , \10527 , \10531 );
and \U$10356 ( \10533 , \3143 , \2400 );
and \U$10357 ( \10534 , \3395 , \2246 );
nor \U$10358 ( \10535 , \10533 , \10534 );
xnor \U$10359 ( \10536 , \10535 , \2195 );
xor \U$10360 ( \10537 , \10532 , \10536 );
and \U$10361 ( \10538 , \5156 , \1086 );
and \U$10362 ( \10539 , \5469 , \508 );
nor \U$10363 ( \10540 , \10538 , \10539 );
xnor \U$10364 ( \10541 , \10540 , \487 );
and \U$10365 ( \10542 , \4749 , \1301 );
and \U$10366 ( \10543 , \4922 , \1246 );
nor \U$10367 ( \10544 , \10542 , \10543 );
xnor \U$10368 ( \10545 , \10544 , \1205 );
xor \U$10369 ( \10546 , \10541 , \10545 );
and \U$10370 ( \10547 , \4364 , \1578 );
and \U$10371 ( \10548 , \4654 , \1431 );
nor \U$10372 ( \10549 , \10547 , \10548 );
xnor \U$10373 ( \10550 , \10549 , \1436 );
xor \U$10374 ( \10551 , \10546 , \10550 );
xor \U$10375 ( \10552 , \10537 , \10551 );
and \U$10376 ( \10553 , \6790 , \156 );
and \U$10377 ( \10554 , \6945 , \154 );
nor \U$10378 ( \10555 , \10553 , \10554 );
xnor \U$10379 ( \10556 , \10555 , \163 );
and \U$10380 ( \10557 , \6281 , \296 );
and \U$10381 ( \10558 , \6514 , \168 );
nor \U$10382 ( \10559 , \10557 , \10558 );
xnor \U$10383 ( \10560 , \10559 , \173 );
xor \U$10384 ( \10561 , \10556 , \10560 );
and \U$10385 ( \10562 , \5674 , \438 );
and \U$10386 ( \10563 , \6030 , \336 );
nor \U$10387 ( \10564 , \10562 , \10563 );
xnor \U$10388 ( \10565 , \10564 , \320 );
xor \U$10389 ( \10566 , \10561 , \10565 );
xor \U$10390 ( \10567 , \10552 , \10566 );
xor \U$10391 ( \10568 , \10523 , \10567 );
and \U$10392 ( \10569 , \8349 , \230 );
and \U$10393 ( \10570 , \8652 , \228 );
nor \U$10394 ( \10571 , \10569 , \10570 );
xnor \U$10395 ( \10572 , \10571 , \237 );
and \U$10396 ( \10573 , \7700 , \245 );
and \U$10397 ( \10574 , \8057 , \243 );
nor \U$10398 ( \10575 , \10573 , \10574 );
xnor \U$10399 ( \10576 , \10575 , \252 );
xor \U$10400 ( \10577 , \10572 , \10576 );
and \U$10401 ( \10578 , \7231 , \141 );
and \U$10402 ( \10579 , \7556 , \139 );
nor \U$10403 ( \10580 , \10578 , \10579 );
xnor \U$10404 ( \10581 , \10580 , \148 );
xor \U$10405 ( \10582 , \10577 , \10581 );
and \U$10406 ( \10583 , \10206 , \183 );
buf \U$10407 ( \10584 , RIb55f1c0_65);
and \U$10408 ( \10585 , \10584 , \180 );
nor \U$10409 ( \10586 , \10583 , \10585 );
xnor \U$10410 ( \10587 , \10586 , \179 );
and \U$10411 ( \10588 , \9465 , \195 );
and \U$10412 ( \10589 , \9897 , \193 );
nor \U$10413 ( \10590 , \10588 , \10589 );
xnor \U$10414 ( \10591 , \10590 , \202 );
xor \U$10415 ( \10592 , \10587 , \10591 );
and \U$10416 ( \10593 , \8835 , \215 );
and \U$10417 ( \10594 , \9169 , \213 );
nor \U$10418 ( \10595 , \10593 , \10594 );
xnor \U$10419 ( \10596 , \10595 , \222 );
xor \U$10420 ( \10597 , \10592 , \10596 );
xor \U$10421 ( \10598 , \10582 , \10597 );
xor \U$10422 ( \10599 , \10568 , \10598 );
xor \U$10423 ( \10600 , \10519 , \10599 );
xor \U$10424 ( \10601 , \10490 , \10600 );
xor \U$10425 ( \10602 , \10328 , \10601 );
xor \U$10426 ( \10603 , \10319 , \10602 );
and \U$10427 ( \10604 , \9976 , \10281 );
xor \U$10428 ( \10605 , \10603 , \10604 );
and \U$10429 ( \10606 , \10282 , \10283 );
and \U$10430 ( \10607 , \10284 , \10287 );
or \U$10431 ( \10608 , \10606 , \10607 );
xor \U$10432 ( \10609 , \10605 , \10608 );
buf g551d_GF_PartitionCandidate( \10610_nG551d , \10609 );
buf \U$10433 ( \10611 , \10610_nG551d );
and \U$10434 ( \10612 , \10298 , \10302 );
and \U$10435 ( \10613 , \10302 , \10317 );
and \U$10436 ( \10614 , \10298 , \10317 );
or \U$10437 ( \10615 , \10612 , \10613 , \10614 );
and \U$10438 ( \10616 , \10323 , \10327 );
and \U$10439 ( \10617 , \10327 , \10601 );
and \U$10440 ( \10618 , \10323 , \10601 );
or \U$10441 ( \10619 , \10616 , \10617 , \10618 );
and \U$10442 ( \10620 , \10307 , \10311 );
and \U$10443 ( \10621 , \10311 , \10316 );
and \U$10444 ( \10622 , \10307 , \10316 );
or \U$10445 ( \10623 , \10620 , \10621 , \10622 );
and \U$10446 ( \10624 , \10342 , \10489 );
and \U$10447 ( \10625 , \10489 , \10600 );
and \U$10448 ( \10626 , \10342 , \10600 );
or \U$10449 ( \10627 , \10624 , \10625 , \10626 );
xor \U$10450 ( \10628 , \10623 , \10627 );
and \U$10451 ( \10629 , \10360 , \10374 );
and \U$10452 ( \10630 , \10374 , \10389 );
and \U$10453 ( \10631 , \10360 , \10389 );
or \U$10454 ( \10632 , \10629 , \10630 , \10631 );
and \U$10455 ( \10633 , \10405 , \10442 );
and \U$10456 ( \10634 , \10442 , \10487 );
and \U$10457 ( \10635 , \10405 , \10487 );
or \U$10458 ( \10636 , \10633 , \10634 , \10635 );
xor \U$10459 ( \10637 , \10632 , \10636 );
and \U$10460 ( \10638 , \10556 , \10560 );
and \U$10461 ( \10639 , \10560 , \10565 );
and \U$10462 ( \10640 , \10556 , \10565 );
or \U$10463 ( \10641 , \10638 , \10639 , \10640 );
and \U$10464 ( \10642 , \10572 , \10576 );
and \U$10465 ( \10643 , \10576 , \10581 );
and \U$10466 ( \10644 , \10572 , \10581 );
or \U$10467 ( \10645 , \10642 , \10643 , \10644 );
xor \U$10468 ( \10646 , \10641 , \10645 );
and \U$10469 ( \10647 , \10587 , \10591 );
and \U$10470 ( \10648 , \10591 , \10596 );
and \U$10471 ( \10649 , \10587 , \10596 );
or \U$10472 ( \10650 , \10647 , \10648 , \10649 );
xor \U$10473 ( \10651 , \10646 , \10650 );
xor \U$10474 ( \10652 , \10637 , \10651 );
xor \U$10475 ( \10653 , \10628 , \10652 );
xor \U$10476 ( \10654 , \10619 , \10653 );
and \U$10477 ( \10655 , \10494 , \10498 );
and \U$10478 ( \10656 , \10498 , \10503 );
and \U$10479 ( \10657 , \10494 , \10503 );
or \U$10480 ( \10658 , \10655 , \10656 , \10657 );
and \U$10481 ( \10659 , \10508 , \10512 );
and \U$10482 ( \10660 , \10512 , \10517 );
and \U$10483 ( \10661 , \10508 , \10517 );
or \U$10484 ( \10662 , \10659 , \10660 , \10661 );
xor \U$10485 ( \10663 , \10658 , \10662 );
and \U$10486 ( \10664 , \10523 , \10567 );
and \U$10487 ( \10665 , \10567 , \10598 );
and \U$10488 ( \10666 , \10523 , \10598 );
or \U$10489 ( \10667 , \10664 , \10665 , \10666 );
xor \U$10490 ( \10668 , \10663 , \10667 );
and \U$10491 ( \10669 , \10332 , \10336 );
and \U$10492 ( \10670 , \10336 , \10341 );
and \U$10493 ( \10671 , \10332 , \10341 );
or \U$10494 ( \10672 , \10669 , \10670 , \10671 );
and \U$10495 ( \10673 , \10346 , \10390 );
and \U$10496 ( \10674 , \10390 , \10488 );
and \U$10497 ( \10675 , \10346 , \10488 );
or \U$10498 ( \10676 , \10673 , \10674 , \10675 );
xor \U$10499 ( \10677 , \10672 , \10676 );
and \U$10500 ( \10678 , \10504 , \10518 );
and \U$10501 ( \10679 , \10518 , \10599 );
and \U$10502 ( \10680 , \10504 , \10599 );
or \U$10503 ( \10681 , \10678 , \10679 , \10680 );
xor \U$10504 ( \10682 , \10677 , \10681 );
xor \U$10505 ( \10683 , \10668 , \10682 );
and \U$10506 ( \10684 , \10395 , \10399 );
and \U$10507 ( \10685 , \10399 , \10404 );
and \U$10508 ( \10686 , \10395 , \10404 );
or \U$10509 ( \10687 , \10684 , \10685 , \10686 );
and \U$10510 ( \10688 , \10412 , \10426 );
and \U$10511 ( \10689 , \10426 , \10441 );
and \U$10512 ( \10690 , \10412 , \10441 );
or \U$10513 ( \10691 , \10688 , \10689 , \10690 );
xor \U$10514 ( \10692 , \10687 , \10691 );
and \U$10515 ( \10693 , \10457 , \10471 );
and \U$10516 ( \10694 , \10471 , \10486 );
and \U$10517 ( \10695 , \10457 , \10486 );
or \U$10518 ( \10696 , \10693 , \10694 , \10695 );
xor \U$10519 ( \10697 , \10692 , \10696 );
and \U$10520 ( \10698 , \10350 , \10354 );
and \U$10521 ( \10699 , \10354 , \10359 );
and \U$10522 ( \10700 , \10350 , \10359 );
or \U$10523 ( \10701 , \10698 , \10699 , \10700 );
and \U$10524 ( \10702 , \10364 , \10368 );
and \U$10525 ( \10703 , \10368 , \10373 );
and \U$10526 ( \10704 , \10364 , \10373 );
or \U$10527 ( \10705 , \10702 , \10703 , \10704 );
xor \U$10528 ( \10706 , \10701 , \10705 );
and \U$10529 ( \10707 , \10379 , \10383 );
and \U$10530 ( \10708 , \10383 , \10388 );
and \U$10531 ( \10709 , \10379 , \10388 );
or \U$10532 ( \10710 , \10707 , \10708 , \10709 );
xor \U$10533 ( \10711 , \10706 , \10710 );
xor \U$10534 ( \10712 , \10697 , \10711 );
and \U$10535 ( \10713 , \10527 , \10531 );
and \U$10536 ( \10714 , \10531 , \10536 );
and \U$10537 ( \10715 , \10527 , \10536 );
or \U$10538 ( \10716 , \10713 , \10714 , \10715 );
and \U$10539 ( \10717 , \10541 , \10545 );
and \U$10540 ( \10718 , \10545 , \10550 );
and \U$10541 ( \10719 , \10541 , \10550 );
or \U$10542 ( \10720 , \10717 , \10718 , \10719 );
xor \U$10543 ( \10721 , \10716 , \10720 );
and \U$10544 ( \10722 , \10476 , \10480 );
and \U$10545 ( \10723 , \10480 , \10485 );
and \U$10546 ( \10724 , \10476 , \10485 );
or \U$10547 ( \10725 , \10722 , \10723 , \10724 );
xor \U$10548 ( \10726 , \10721 , \10725 );
and \U$10549 ( \10727 , \10447 , \10451 );
and \U$10550 ( \10728 , \10451 , \10456 );
and \U$10551 ( \10729 , \10447 , \10456 );
or \U$10552 ( \10730 , \10727 , \10728 , \10729 );
and \U$10553 ( \10731 , \10461 , \10465 );
and \U$10554 ( \10732 , \10465 , \10470 );
and \U$10555 ( \10733 , \10461 , \10470 );
or \U$10556 ( \10734 , \10731 , \10732 , \10733 );
xor \U$10557 ( \10735 , \10730 , \10734 );
and \U$10558 ( \10736 , \10416 , \10420 );
and \U$10559 ( \10737 , \10420 , \10425 );
and \U$10560 ( \10738 , \10416 , \10425 );
or \U$10561 ( \10739 , \10736 , \10737 , \10738 );
xor \U$10562 ( \10740 , \10735 , \10739 );
xor \U$10563 ( \10741 , \10726 , \10740 );
and \U$10564 ( \10742 , \10431 , \10435 );
and \U$10565 ( \10743 , \10435 , \10440 );
and \U$10566 ( \10744 , \10431 , \10440 );
or \U$10567 ( \10745 , \10742 , \10743 , \10744 );
nand \U$10568 ( \10746 , \166 , \10118 );
not \U$10569 ( \10747 , \10746 );
xor \U$10570 ( \10748 , \10745 , \10747 );
and \U$10571 ( \10749 , \240 , \9333 );
and \U$10572 ( \10750 , \247 , \9006 );
nor \U$10573 ( \10751 , \10749 , \10750 );
xnor \U$10574 ( \10752 , \10751 , \8848 );
and \U$10575 ( \10753 , \134 , \9765 );
and \U$10576 ( \10754 , \143 , \9644 );
nor \U$10577 ( \10755 , \10753 , \10754 );
xnor \U$10578 ( \10756 , \10755 , \9478 );
xor \U$10579 ( \10757 , \10752 , \10756 );
and \U$10580 ( \10758 , \150 , \10408 );
and \U$10581 ( \10759 , \158 , \10116 );
nor \U$10582 ( \10760 , \10758 , \10759 );
xnor \U$10583 ( \10761 , \10760 , \10121 );
xor \U$10584 ( \10762 , \10757 , \10761 );
xor \U$10585 ( \10763 , \10748 , \10762 );
xor \U$10586 ( \10764 , \10741 , \10763 );
and \U$10587 ( \10765 , \9169 , \215 );
and \U$10588 ( \10766 , \9465 , \213 );
nor \U$10589 ( \10767 , \10765 , \10766 );
xnor \U$10590 ( \10768 , \10767 , \222 );
and \U$10591 ( \10769 , \8652 , \230 );
and \U$10592 ( \10770 , \8835 , \228 );
nor \U$10593 ( \10771 , \10769 , \10770 );
xnor \U$10594 ( \10772 , \10771 , \237 );
xor \U$10595 ( \10773 , \10768 , \10772 );
and \U$10596 ( \10774 , \8057 , \245 );
and \U$10597 ( \10775 , \8349 , \243 );
nor \U$10598 ( \10776 , \10774 , \10775 );
xnor \U$10599 ( \10777 , \10776 , \252 );
xor \U$10600 ( \10778 , \10773 , \10777 );
and \U$10601 ( \10779 , \7556 , \141 );
and \U$10602 ( \10780 , \7700 , \139 );
nor \U$10603 ( \10781 , \10779 , \10780 );
xnor \U$10604 ( \10782 , \10781 , \148 );
and \U$10605 ( \10783 , \6945 , \156 );
and \U$10606 ( \10784 , \7231 , \154 );
nor \U$10607 ( \10785 , \10783 , \10784 );
xnor \U$10608 ( \10786 , \10785 , \163 );
xor \U$10609 ( \10787 , \10782 , \10786 );
and \U$10610 ( \10788 , \6514 , \296 );
and \U$10611 ( \10789 , \6790 , \168 );
nor \U$10612 ( \10790 , \10788 , \10789 );
xnor \U$10613 ( \10791 , \10790 , \173 );
xor \U$10614 ( \10792 , \10787 , \10791 );
xor \U$10615 ( \10793 , \10778 , \10792 );
and \U$10616 ( \10794 , \6030 , \438 );
and \U$10617 ( \10795 , \6281 , \336 );
nor \U$10618 ( \10796 , \10794 , \10795 );
xnor \U$10619 ( \10797 , \10796 , \320 );
and \U$10620 ( \10798 , \5469 , \1086 );
and \U$10621 ( \10799 , \5674 , \508 );
nor \U$10622 ( \10800 , \10798 , \10799 );
xnor \U$10623 ( \10801 , \10800 , \487 );
xor \U$10624 ( \10802 , \10797 , \10801 );
and \U$10625 ( \10803 , \4922 , \1301 );
and \U$10626 ( \10804 , \5156 , \1246 );
nor \U$10627 ( \10805 , \10803 , \10804 );
xnor \U$10628 ( \10806 , \10805 , \1205 );
xor \U$10629 ( \10807 , \10802 , \10806 );
xor \U$10630 ( \10808 , \10793 , \10807 );
and \U$10631 ( \10809 , \1601 , \4581 );
and \U$10632 ( \10810 , \1684 , \4424 );
nor \U$10633 ( \10811 , \10809 , \10810 );
xnor \U$10634 ( \10812 , \10811 , \4377 );
and \U$10635 ( \10813 , \1333 , \5011 );
and \U$10636 ( \10814 , \1484 , \4878 );
nor \U$10637 ( \10815 , \10813 , \10814 );
xnor \U$10638 ( \10816 , \10815 , \4762 );
xor \U$10639 ( \10817 , \10812 , \10816 );
and \U$10640 ( \10818 , \1147 , \5485 );
and \U$10641 ( \10819 , \1192 , \5275 );
nor \U$10642 ( \10820 , \10818 , \10819 );
xnor \U$10643 ( \10821 , \10820 , \5169 );
xor \U$10644 ( \10822 , \10817 , \10821 );
and \U$10645 ( \10823 , \189 , \7489 );
and \U$10646 ( \10824 , \197 , \7137 );
nor \U$10647 ( \10825 , \10823 , \10824 );
xnor \U$10648 ( \10826 , \10825 , \7142 );
and \U$10649 ( \10827 , \209 , \8019 );
and \U$10650 ( \10828 , \217 , \7830 );
nor \U$10651 ( \10829 , \10827 , \10828 );
xnor \U$10652 ( \10830 , \10829 , \7713 );
xor \U$10653 ( \10831 , \10826 , \10830 );
and \U$10654 ( \10832 , \224 , \8540 );
and \U$10655 ( \10833 , \232 , \8292 );
nor \U$10656 ( \10834 , \10832 , \10833 );
xnor \U$10657 ( \10835 , \10834 , \8297 );
xor \U$10658 ( \10836 , \10831 , \10835 );
xor \U$10659 ( \10837 , \10822 , \10836 );
and \U$10660 ( \10838 , \412 , \5996 );
and \U$10661 ( \10839 , \474 , \5695 );
nor \U$10662 ( \10840 , \10838 , \10839 );
xnor \U$10663 ( \10841 , \10840 , \5687 );
and \U$10664 ( \10842 , \261 , \6401 );
and \U$10665 ( \10843 , \307 , \6143 );
nor \U$10666 ( \10844 , \10842 , \10843 );
xnor \U$10667 ( \10845 , \10844 , \6148 );
xor \U$10668 ( \10846 , \10841 , \10845 );
and \U$10669 ( \10847 , \178 , \7055 );
and \U$10670 ( \10848 , \185 , \6675 );
nor \U$10671 ( \10849 , \10847 , \10848 );
xnor \U$10672 ( \10850 , \10849 , \6680 );
xor \U$10673 ( \10851 , \10846 , \10850 );
xor \U$10674 ( \10852 , \10837 , \10851 );
xor \U$10675 ( \10853 , \10808 , \10852 );
and \U$10676 ( \10854 , \4654 , \1578 );
and \U$10677 ( \10855 , \4749 , \1431 );
nor \U$10678 ( \10856 , \10854 , \10855 );
xnor \U$10679 ( \10857 , \10856 , \1436 );
and \U$10680 ( \10858 , \4160 , \1824 );
and \U$10681 ( \10859 , \4364 , \1739 );
nor \U$10682 ( \10860 , \10858 , \10859 );
xnor \U$10683 ( \10861 , \10860 , \1697 );
xor \U$10684 ( \10862 , \10857 , \10861 );
and \U$10685 ( \10863 , \3736 , \2121 );
and \U$10686 ( \10864 , \3912 , \2008 );
nor \U$10687 ( \10865 , \10863 , \10864 );
xnor \U$10688 ( \10866 , \10865 , \1961 );
xor \U$10689 ( \10867 , \10862 , \10866 );
and \U$10690 ( \10868 , \3395 , \2400 );
and \U$10691 ( \10869 , \3646 , \2246 );
nor \U$10692 ( \10870 , \10868 , \10869 );
xnor \U$10693 ( \10871 , \10870 , \2195 );
and \U$10694 ( \10872 , \3037 , \2669 );
and \U$10695 ( \10873 , \3143 , \2538 );
nor \U$10696 ( \10874 , \10872 , \10873 );
xnor \U$10697 ( \10875 , \10874 , \2534 );
xor \U$10698 ( \10876 , \10871 , \10875 );
and \U$10699 ( \10877 , \2757 , \3103 );
and \U$10700 ( \10878 , \2826 , \2934 );
nor \U$10701 ( \10879 , \10877 , \10878 );
xnor \U$10702 ( \10880 , \10879 , \2839 );
xor \U$10703 ( \10881 , \10876 , \10880 );
xor \U$10704 ( \10882 , \10867 , \10881 );
and \U$10705 ( \10883 , \2366 , \3357 );
and \U$10706 ( \10884 , \2521 , \3255 );
nor \U$10707 ( \10885 , \10883 , \10884 );
xnor \U$10708 ( \10886 , \10885 , \3156 );
and \U$10709 ( \10887 , \2090 , \3813 );
and \U$10710 ( \10888 , \2182 , \3557 );
nor \U$10711 ( \10889 , \10887 , \10888 );
xnor \U$10712 ( \10890 , \10889 , \3562 );
xor \U$10713 ( \10891 , \10886 , \10890 );
and \U$10714 ( \10892 , \1802 , \4132 );
and \U$10715 ( \10893 , \1948 , \4012 );
nor \U$10716 ( \10894 , \10892 , \10893 );
xnor \U$10717 ( \10895 , \10894 , \3925 );
xor \U$10718 ( \10896 , \10891 , \10895 );
xor \U$10719 ( \10897 , \10882 , \10896 );
xor \U$10720 ( \10898 , \10853 , \10897 );
xor \U$10721 ( \10899 , \10764 , \10898 );
and \U$10722 ( \10900 , \10537 , \10551 );
and \U$10723 ( \10901 , \10551 , \10566 );
and \U$10724 ( \10902 , \10537 , \10566 );
or \U$10725 ( \10903 , \10900 , \10901 , \10902 );
and \U$10726 ( \10904 , \10582 , \10597 );
xor \U$10727 ( \10905 , \10903 , \10904 );
and \U$10728 ( \10906 , \10584 , \183 );
not \U$10729 ( \10907 , \10906 );
xnor \U$10730 ( \10908 , \10907 , \179 );
and \U$10731 ( \10909 , \9897 , \195 );
and \U$10732 ( \10910 , \10206 , \193 );
nor \U$10733 ( \10911 , \10909 , \10910 );
xnor \U$10734 ( \10912 , \10911 , \202 );
xor \U$10735 ( \10913 , \10908 , \10912 );
xor \U$10736 ( \10914 , \10905 , \10913 );
xor \U$10737 ( \10915 , \10899 , \10914 );
xor \U$10738 ( \10916 , \10712 , \10915 );
xor \U$10739 ( \10917 , \10683 , \10916 );
xor \U$10740 ( \10918 , \10654 , \10917 );
xor \U$10741 ( \10919 , \10615 , \10918 );
and \U$10742 ( \10920 , \10294 , \10318 );
and \U$10743 ( \10921 , \10318 , \10602 );
and \U$10744 ( \10922 , \10294 , \10602 );
or \U$10745 ( \10923 , \10920 , \10921 , \10922 );
xor \U$10746 ( \10924 , \10919 , \10923 );
and \U$10747 ( \10925 , \10603 , \10604 );
and \U$10748 ( \10926 , \10605 , \10608 );
or \U$10749 ( \10927 , \10925 , \10926 );
xor \U$10750 ( \10928 , \10924 , \10927 );
buf g551b_GF_PartitionCandidate( \10929_nG551b , \10928 );
buf \U$10751 ( \10930 , \10929_nG551b );
and \U$10752 ( \10931 , \10619 , \10653 );
and \U$10753 ( \10932 , \10653 , \10917 );
and \U$10754 ( \10933 , \10619 , \10917 );
or \U$10755 ( \10934 , \10931 , \10932 , \10933 );
and \U$10756 ( \10935 , \10623 , \10627 );
and \U$10757 ( \10936 , \10627 , \10652 );
and \U$10758 ( \10937 , \10623 , \10652 );
or \U$10759 ( \10938 , \10935 , \10936 , \10937 );
and \U$10760 ( \10939 , \10668 , \10682 );
and \U$10761 ( \10940 , \10682 , \10916 );
and \U$10762 ( \10941 , \10668 , \10916 );
or \U$10763 ( \10942 , \10939 , \10940 , \10941 );
xor \U$10764 ( \10943 , \10938 , \10942 );
and \U$10765 ( \10944 , \10716 , \10720 );
and \U$10766 ( \10945 , \10720 , \10725 );
and \U$10767 ( \10946 , \10716 , \10725 );
or \U$10768 ( \10947 , \10944 , \10945 , \10946 );
and \U$10769 ( \10948 , \10641 , \10645 );
and \U$10770 ( \10949 , \10645 , \10650 );
and \U$10771 ( \10950 , \10641 , \10650 );
or \U$10772 ( \10951 , \10948 , \10949 , \10950 );
xor \U$10773 ( \10952 , \10947 , \10951 );
and \U$10774 ( \10953 , \10730 , \10734 );
and \U$10775 ( \10954 , \10734 , \10739 );
and \U$10776 ( \10955 , \10730 , \10739 );
or \U$10777 ( \10956 , \10953 , \10954 , \10955 );
xor \U$10778 ( \10957 , \10952 , \10956 );
and \U$10779 ( \10958 , \10726 , \10740 );
and \U$10780 ( \10959 , \10740 , \10763 );
and \U$10781 ( \10960 , \10726 , \10763 );
or \U$10782 ( \10961 , \10958 , \10959 , \10960 );
and \U$10783 ( \10962 , \10808 , \10852 );
and \U$10784 ( \10963 , \10852 , \10897 );
and \U$10785 ( \10964 , \10808 , \10897 );
or \U$10786 ( \10965 , \10962 , \10963 , \10964 );
xor \U$10787 ( \10966 , \10961 , \10965 );
and \U$10788 ( \10967 , \10812 , \10816 );
and \U$10789 ( \10968 , \10816 , \10821 );
and \U$10790 ( \10969 , \10812 , \10821 );
or \U$10791 ( \10970 , \10967 , \10968 , \10969 );
and \U$10792 ( \10971 , \10841 , \10845 );
and \U$10793 ( \10972 , \10845 , \10850 );
and \U$10794 ( \10973 , \10841 , \10850 );
or \U$10795 ( \10974 , \10971 , \10972 , \10973 );
xor \U$10796 ( \10975 , \10970 , \10974 );
and \U$10797 ( \10976 , \10886 , \10890 );
and \U$10798 ( \10977 , \10890 , \10895 );
and \U$10799 ( \10978 , \10886 , \10895 );
or \U$10800 ( \10979 , \10976 , \10977 , \10978 );
xor \U$10801 ( \10980 , \10975 , \10979 );
and \U$10802 ( \10981 , \10857 , \10861 );
and \U$10803 ( \10982 , \10861 , \10866 );
and \U$10804 ( \10983 , \10857 , \10866 );
or \U$10805 ( \10984 , \10981 , \10982 , \10983 );
and \U$10806 ( \10985 , \10871 , \10875 );
and \U$10807 ( \10986 , \10875 , \10880 );
and \U$10808 ( \10987 , \10871 , \10880 );
or \U$10809 ( \10988 , \10985 , \10986 , \10987 );
xor \U$10810 ( \10989 , \10984 , \10988 );
and \U$10811 ( \10990 , \10797 , \10801 );
and \U$10812 ( \10991 , \10801 , \10806 );
and \U$10813 ( \10992 , \10797 , \10806 );
or \U$10814 ( \10993 , \10990 , \10991 , \10992 );
xor \U$10815 ( \10994 , \10989 , \10993 );
xor \U$10816 ( \10995 , \10980 , \10994 );
and \U$10817 ( \10996 , \10768 , \10772 );
and \U$10818 ( \10997 , \10772 , \10777 );
and \U$10819 ( \10998 , \10768 , \10777 );
or \U$10820 ( \10999 , \10996 , \10997 , \10998 );
and \U$10821 ( \11000 , \10782 , \10786 );
and \U$10822 ( \11001 , \10786 , \10791 );
and \U$10823 ( \11002 , \10782 , \10791 );
or \U$10824 ( \11003 , \11000 , \11001 , \11002 );
xor \U$10825 ( \11004 , \10999 , \11003 );
and \U$10826 ( \11005 , \10908 , \10912 );
xor \U$10827 ( \11006 , \11004 , \11005 );
xor \U$10828 ( \11007 , \10995 , \11006 );
xor \U$10829 ( \11008 , \10966 , \11007 );
xor \U$10830 ( \11009 , \10957 , \11008 );
and \U$10831 ( \11010 , \10822 , \10836 );
and \U$10832 ( \11011 , \10836 , \10851 );
and \U$10833 ( \11012 , \10822 , \10851 );
or \U$10834 ( \11013 , \11010 , \11011 , \11012 );
and \U$10835 ( \11014 , \10867 , \10881 );
and \U$10836 ( \11015 , \10881 , \10896 );
and \U$10837 ( \11016 , \10867 , \10896 );
or \U$10838 ( \11017 , \11014 , \11015 , \11016 );
xor \U$10839 ( \11018 , \11013 , \11017 );
and \U$10840 ( \11019 , \10745 , \10747 );
and \U$10841 ( \11020 , \10747 , \10762 );
and \U$10842 ( \11021 , \10745 , \10762 );
or \U$10843 ( \11022 , \11019 , \11020 , \11021 );
xor \U$10844 ( \11023 , \11018 , \11022 );
and \U$10845 ( \11024 , \1484 , \5011 );
and \U$10846 ( \11025 , \1601 , \4878 );
nor \U$10847 ( \11026 , \11024 , \11025 );
xnor \U$10848 ( \11027 , \11026 , \4762 );
and \U$10849 ( \11028 , \1192 , \5485 );
and \U$10850 ( \11029 , \1333 , \5275 );
nor \U$10851 ( \11030 , \11028 , \11029 );
xnor \U$10852 ( \11031 , \11030 , \5169 );
xor \U$10853 ( \11032 , \11027 , \11031 );
and \U$10854 ( \11033 , \474 , \5996 );
and \U$10855 ( \11034 , \1147 , \5695 );
nor \U$10856 ( \11035 , \11033 , \11034 );
xnor \U$10857 ( \11036 , \11035 , \5687 );
xor \U$10858 ( \11037 , \11032 , \11036 );
and \U$10859 ( \11038 , \2182 , \3813 );
and \U$10860 ( \11039 , \2366 , \3557 );
nor \U$10861 ( \11040 , \11038 , \11039 );
xnor \U$10862 ( \11041 , \11040 , \3562 );
and \U$10863 ( \11042 , \1948 , \4132 );
and \U$10864 ( \11043 , \2090 , \4012 );
nor \U$10865 ( \11044 , \11042 , \11043 );
xnor \U$10866 ( \11045 , \11044 , \3925 );
xor \U$10867 ( \11046 , \11041 , \11045 );
and \U$10868 ( \11047 , \1684 , \4581 );
and \U$10869 ( \11048 , \1802 , \4424 );
nor \U$10870 ( \11049 , \11047 , \11048 );
xnor \U$10871 ( \11050 , \11049 , \4377 );
xor \U$10872 ( \11051 , \11046 , \11050 );
xor \U$10873 ( \11052 , \11037 , \11051 );
and \U$10874 ( \11053 , \3143 , \2669 );
and \U$10875 ( \11054 , \3395 , \2538 );
nor \U$10876 ( \11055 , \11053 , \11054 );
xnor \U$10877 ( \11056 , \11055 , \2534 );
and \U$10878 ( \11057 , \2826 , \3103 );
and \U$10879 ( \11058 , \3037 , \2934 );
nor \U$10880 ( \11059 , \11057 , \11058 );
xnor \U$10881 ( \11060 , \11059 , \2839 );
xor \U$10882 ( \11061 , \11056 , \11060 );
and \U$10883 ( \11062 , \2521 , \3357 );
and \U$10884 ( \11063 , \2757 , \3255 );
nor \U$10885 ( \11064 , \11062 , \11063 );
xnor \U$10886 ( \11065 , \11064 , \3156 );
xor \U$10887 ( \11066 , \11061 , \11065 );
xor \U$10888 ( \11067 , \11052 , \11066 );
and \U$10889 ( \11068 , \217 , \8019 );
and \U$10890 ( \11069 , \189 , \7830 );
nor \U$10891 ( \11070 , \11068 , \11069 );
xnor \U$10892 ( \11071 , \11070 , \7713 );
and \U$10893 ( \11072 , \232 , \8540 );
and \U$10894 ( \11073 , \209 , \8292 );
nor \U$10895 ( \11074 , \11072 , \11073 );
xnor \U$10896 ( \11075 , \11074 , \8297 );
xor \U$10897 ( \11076 , \11071 , \11075 );
and \U$10898 ( \11077 , \247 , \9333 );
and \U$10899 ( \11078 , \224 , \9006 );
nor \U$10900 ( \11079 , \11077 , \11078 );
xnor \U$10901 ( \11080 , \11079 , \8848 );
xor \U$10902 ( \11081 , \11076 , \11080 );
and \U$10903 ( \11082 , \143 , \9765 );
and \U$10904 ( \11083 , \240 , \9644 );
nor \U$10905 ( \11084 , \11082 , \11083 );
xnor \U$10906 ( \11085 , \11084 , \9478 );
and \U$10907 ( \11086 , \158 , \10408 );
and \U$10908 ( \11087 , \134 , \10116 );
nor \U$10909 ( \11088 , \11086 , \11087 );
xnor \U$10910 ( \11089 , \11088 , \10121 );
xor \U$10911 ( \11090 , \11085 , \11089 );
and \U$10912 ( \11091 , \150 , \10118 );
xor \U$10913 ( \11092 , \11090 , \11091 );
xor \U$10914 ( \11093 , \11081 , \11092 );
and \U$10915 ( \11094 , \307 , \6401 );
and \U$10916 ( \11095 , \412 , \6143 );
nor \U$10917 ( \11096 , \11094 , \11095 );
xnor \U$10918 ( \11097 , \11096 , \6148 );
and \U$10919 ( \11098 , \185 , \7055 );
and \U$10920 ( \11099 , \261 , \6675 );
nor \U$10921 ( \11100 , \11098 , \11099 );
xnor \U$10922 ( \11101 , \11100 , \6680 );
xor \U$10923 ( \11102 , \11097 , \11101 );
and \U$10924 ( \11103 , \197 , \7489 );
and \U$10925 ( \11104 , \178 , \7137 );
nor \U$10926 ( \11105 , \11103 , \11104 );
xnor \U$10927 ( \11106 , \11105 , \7142 );
xor \U$10928 ( \11107 , \11102 , \11106 );
xor \U$10929 ( \11108 , \11093 , \11107 );
xor \U$10930 ( \11109 , \11067 , \11108 );
and \U$10931 ( \11110 , \10826 , \10830 );
and \U$10932 ( \11111 , \10830 , \10835 );
and \U$10933 ( \11112 , \10826 , \10835 );
or \U$10934 ( \11113 , \11110 , \11111 , \11112 );
and \U$10935 ( \11114 , \10752 , \10756 );
and \U$10936 ( \11115 , \10756 , \10761 );
and \U$10937 ( \11116 , \10752 , \10761 );
or \U$10938 ( \11117 , \11114 , \11115 , \11116 );
xnor \U$10939 ( \11118 , \11113 , \11117 );
xor \U$10940 ( \11119 , \11109 , \11118 );
xor \U$10941 ( \11120 , \11023 , \11119 );
and \U$10942 ( \11121 , \10778 , \10792 );
and \U$10943 ( \11122 , \10792 , \10807 );
and \U$10944 ( \11123 , \10778 , \10807 );
or \U$10945 ( \11124 , \11121 , \11122 , \11123 );
and \U$10946 ( \11125 , \4364 , \1824 );
and \U$10947 ( \11126 , \4654 , \1739 );
nor \U$10948 ( \11127 , \11125 , \11126 );
xnor \U$10949 ( \11128 , \11127 , \1697 );
and \U$10950 ( \11129 , \3912 , \2121 );
and \U$10951 ( \11130 , \4160 , \2008 );
nor \U$10952 ( \11131 , \11129 , \11130 );
xnor \U$10953 ( \11132 , \11131 , \1961 );
xor \U$10954 ( \11133 , \11128 , \11132 );
and \U$10955 ( \11134 , \3646 , \2400 );
and \U$10956 ( \11135 , \3736 , \2246 );
nor \U$10957 ( \11136 , \11134 , \11135 );
xnor \U$10958 ( \11137 , \11136 , \2195 );
xor \U$10959 ( \11138 , \11133 , \11137 );
and \U$10960 ( \11139 , \7231 , \156 );
and \U$10961 ( \11140 , \7556 , \154 );
nor \U$10962 ( \11141 , \11139 , \11140 );
xnor \U$10963 ( \11142 , \11141 , \163 );
and \U$10964 ( \11143 , \6790 , \296 );
and \U$10965 ( \11144 , \6945 , \168 );
nor \U$10966 ( \11145 , \11143 , \11144 );
xnor \U$10967 ( \11146 , \11145 , \173 );
xor \U$10968 ( \11147 , \11142 , \11146 );
and \U$10969 ( \11148 , \6281 , \438 );
and \U$10970 ( \11149 , \6514 , \336 );
nor \U$10971 ( \11150 , \11148 , \11149 );
xnor \U$10972 ( \11151 , \11150 , \320 );
xor \U$10973 ( \11152 , \11147 , \11151 );
xor \U$10974 ( \11153 , \11138 , \11152 );
and \U$10975 ( \11154 , \5674 , \1086 );
and \U$10976 ( \11155 , \6030 , \508 );
nor \U$10977 ( \11156 , \11154 , \11155 );
xnor \U$10978 ( \11157 , \11156 , \487 );
and \U$10979 ( \11158 , \5156 , \1301 );
and \U$10980 ( \11159 , \5469 , \1246 );
nor \U$10981 ( \11160 , \11158 , \11159 );
xnor \U$10982 ( \11161 , \11160 , \1205 );
xor \U$10983 ( \11162 , \11157 , \11161 );
and \U$10984 ( \11163 , \4749 , \1578 );
and \U$10985 ( \11164 , \4922 , \1431 );
nor \U$10986 ( \11165 , \11163 , \11164 );
xnor \U$10987 ( \11166 , \11165 , \1436 );
xor \U$10988 ( \11167 , \11162 , \11166 );
xor \U$10989 ( \11168 , \11153 , \11167 );
xor \U$10990 ( \11169 , \11124 , \11168 );
not \U$10991 ( \11170 , \179 );
and \U$10992 ( \11171 , \10206 , \195 );
and \U$10993 ( \11172 , \10584 , \193 );
nor \U$10994 ( \11173 , \11171 , \11172 );
xnor \U$10995 ( \11174 , \11173 , \202 );
xor \U$10996 ( \11175 , \11170 , \11174 );
and \U$10997 ( \11176 , \9465 , \215 );
and \U$10998 ( \11177 , \9897 , \213 );
nor \U$10999 ( \11178 , \11176 , \11177 );
xnor \U$11000 ( \11179 , \11178 , \222 );
xor \U$11001 ( \11180 , \11175 , \11179 );
and \U$11002 ( \11181 , \8835 , \230 );
and \U$11003 ( \11182 , \9169 , \228 );
nor \U$11004 ( \11183 , \11181 , \11182 );
xnor \U$11005 ( \11184 , \11183 , \237 );
and \U$11006 ( \11185 , \8349 , \245 );
and \U$11007 ( \11186 , \8652 , \243 );
nor \U$11008 ( \11187 , \11185 , \11186 );
xnor \U$11009 ( \11188 , \11187 , \252 );
xor \U$11010 ( \11189 , \11184 , \11188 );
and \U$11011 ( \11190 , \7700 , \141 );
and \U$11012 ( \11191 , \8057 , \139 );
nor \U$11013 ( \11192 , \11190 , \11191 );
xnor \U$11014 ( \11193 , \11192 , \148 );
xor \U$11015 ( \11194 , \11189 , \11193 );
xor \U$11016 ( \11195 , \11180 , \11194 );
xor \U$11017 ( \11196 , \11169 , \11195 );
xor \U$11018 ( \11197 , \11120 , \11196 );
xor \U$11019 ( \11198 , \11009 , \11197 );
xor \U$11020 ( \11199 , \10943 , \11198 );
xor \U$11021 ( \11200 , \10934 , \11199 );
and \U$11022 ( \11201 , \10658 , \10662 );
and \U$11023 ( \11202 , \10662 , \10667 );
and \U$11024 ( \11203 , \10658 , \10667 );
or \U$11025 ( \11204 , \11201 , \11202 , \11203 );
and \U$11026 ( \11205 , \10632 , \10636 );
and \U$11027 ( \11206 , \10636 , \10651 );
and \U$11028 ( \11207 , \10632 , \10651 );
or \U$11029 ( \11208 , \11205 , \11206 , \11207 );
xor \U$11030 ( \11209 , \11204 , \11208 );
and \U$11031 ( \11210 , \10764 , \10898 );
and \U$11032 ( \11211 , \10898 , \10914 );
and \U$11033 ( \11212 , \10764 , \10914 );
or \U$11034 ( \11213 , \11210 , \11211 , \11212 );
xor \U$11035 ( \11214 , \11209 , \11213 );
and \U$11036 ( \11215 , \10672 , \10676 );
and \U$11037 ( \11216 , \10676 , \10681 );
and \U$11038 ( \11217 , \10672 , \10681 );
or \U$11039 ( \11218 , \11215 , \11216 , \11217 );
and \U$11040 ( \11219 , \10697 , \10711 );
and \U$11041 ( \11220 , \10711 , \10915 );
and \U$11042 ( \11221 , \10697 , \10915 );
or \U$11043 ( \11222 , \11219 , \11220 , \11221 );
xor \U$11044 ( \11223 , \11218 , \11222 );
and \U$11045 ( \11224 , \10687 , \10691 );
and \U$11046 ( \11225 , \10691 , \10696 );
and \U$11047 ( \11226 , \10687 , \10696 );
or \U$11048 ( \11227 , \11224 , \11225 , \11226 );
and \U$11049 ( \11228 , \10701 , \10705 );
and \U$11050 ( \11229 , \10705 , \10710 );
and \U$11051 ( \11230 , \10701 , \10710 );
or \U$11052 ( \11231 , \11228 , \11229 , \11230 );
xor \U$11053 ( \11232 , \11227 , \11231 );
and \U$11054 ( \11233 , \10903 , \10904 );
and \U$11055 ( \11234 , \10904 , \10913 );
and \U$11056 ( \11235 , \10903 , \10913 );
or \U$11057 ( \11236 , \11233 , \11234 , \11235 );
xor \U$11058 ( \11237 , \11232 , \11236 );
xor \U$11059 ( \11238 , \11223 , \11237 );
xor \U$11060 ( \11239 , \11214 , \11238 );
xor \U$11061 ( \11240 , \11200 , \11239 );
and \U$11062 ( \11241 , \10615 , \10918 );
xor \U$11063 ( \11242 , \11240 , \11241 );
and \U$11064 ( \11243 , \10919 , \10923 );
and \U$11065 ( \11244 , \10924 , \10927 );
or \U$11066 ( \11245 , \11243 , \11244 );
xor \U$11067 ( \11246 , \11242 , \11245 );
buf g5519_GF_PartitionCandidate( \11247_nG5519 , \11246 );
buf \U$11068 ( \11248 , \11247_nG5519 );
and \U$11069 ( \11249 , \10938 , \10942 );
and \U$11070 ( \11250 , \10942 , \11198 );
and \U$11071 ( \11251 , \10938 , \11198 );
or \U$11072 ( \11252 , \11249 , \11250 , \11251 );
and \U$11073 ( \11253 , \11214 , \11238 );
xor \U$11074 ( \11254 , \11252 , \11253 );
and \U$11075 ( \11255 , \11218 , \11222 );
and \U$11076 ( \11256 , \11222 , \11237 );
and \U$11077 ( \11257 , \11218 , \11237 );
or \U$11078 ( \11258 , \11255 , \11256 , \11257 );
and \U$11079 ( \11259 , \11204 , \11208 );
and \U$11080 ( \11260 , \11208 , \11213 );
and \U$11081 ( \11261 , \11204 , \11213 );
or \U$11082 ( \11262 , \11259 , \11260 , \11261 );
and \U$11083 ( \11263 , \10957 , \11008 );
and \U$11084 ( \11264 , \11008 , \11197 );
and \U$11085 ( \11265 , \10957 , \11197 );
or \U$11086 ( \11266 , \11263 , \11264 , \11265 );
xor \U$11087 ( \11267 , \11262 , \11266 );
and \U$11088 ( \11268 , \10980 , \10994 );
and \U$11089 ( \11269 , \10994 , \11006 );
and \U$11090 ( \11270 , \10980 , \11006 );
or \U$11091 ( \11271 , \11268 , \11269 , \11270 );
and \U$11092 ( \11272 , \11067 , \11108 );
and \U$11093 ( \11273 , \11108 , \11118 );
and \U$11094 ( \11274 , \11067 , \11118 );
or \U$11095 ( \11275 , \11272 , \11273 , \11274 );
xor \U$11096 ( \11276 , \11271 , \11275 );
and \U$11097 ( \11277 , \11170 , \11174 );
and \U$11098 ( \11278 , \11174 , \11179 );
and \U$11099 ( \11279 , \11170 , \11179 );
or \U$11100 ( \11280 , \11277 , \11278 , \11279 );
and \U$11101 ( \11281 , \11184 , \11188 );
and \U$11102 ( \11282 , \11188 , \11193 );
and \U$11103 ( \11283 , \11184 , \11193 );
or \U$11104 ( \11284 , \11281 , \11282 , \11283 );
xor \U$11105 ( \11285 , \11280 , \11284 );
and \U$11106 ( \11286 , \11142 , \11146 );
and \U$11107 ( \11287 , \11146 , \11151 );
and \U$11108 ( \11288 , \11142 , \11151 );
or \U$11109 ( \11289 , \11286 , \11287 , \11288 );
xor \U$11110 ( \11290 , \11285 , \11289 );
xor \U$11111 ( \11291 , \11276 , \11290 );
xor \U$11112 ( \11292 , \11267 , \11291 );
xor \U$11113 ( \11293 , \11258 , \11292 );
and \U$11114 ( \11294 , \11013 , \11017 );
and \U$11115 ( \11295 , \11017 , \11022 );
and \U$11116 ( \11296 , \11013 , \11022 );
or \U$11117 ( \11297 , \11294 , \11295 , \11296 );
and \U$11118 ( \11298 , \10947 , \10951 );
and \U$11119 ( \11299 , \10951 , \10956 );
and \U$11120 ( \11300 , \10947 , \10956 );
or \U$11121 ( \11301 , \11298 , \11299 , \11300 );
xor \U$11122 ( \11302 , \11297 , \11301 );
and \U$11123 ( \11303 , \11124 , \11168 );
and \U$11124 ( \11304 , \11168 , \11195 );
and \U$11125 ( \11305 , \11124 , \11195 );
or \U$11126 ( \11306 , \11303 , \11304 , \11305 );
xor \U$11127 ( \11307 , \11302 , \11306 );
and \U$11128 ( \11308 , \11227 , \11231 );
and \U$11129 ( \11309 , \11231 , \11236 );
and \U$11130 ( \11310 , \11227 , \11236 );
or \U$11131 ( \11311 , \11308 , \11309 , \11310 );
and \U$11132 ( \11312 , \10961 , \10965 );
and \U$11133 ( \11313 , \10965 , \11007 );
and \U$11134 ( \11314 , \10961 , \11007 );
or \U$11135 ( \11315 , \11312 , \11313 , \11314 );
xor \U$11136 ( \11316 , \11311 , \11315 );
and \U$11137 ( \11317 , \11023 , \11119 );
and \U$11138 ( \11318 , \11119 , \11196 );
and \U$11139 ( \11319 , \11023 , \11196 );
or \U$11140 ( \11320 , \11317 , \11318 , \11319 );
xor \U$11141 ( \11321 , \11316 , \11320 );
xor \U$11142 ( \11322 , \11307 , \11321 );
and \U$11143 ( \11323 , \11037 , \11051 );
and \U$11144 ( \11324 , \11051 , \11066 );
and \U$11145 ( \11325 , \11037 , \11066 );
or \U$11146 ( \11326 , \11323 , \11324 , \11325 );
and \U$11147 ( \11327 , \11081 , \11092 );
and \U$11148 ( \11328 , \11092 , \11107 );
and \U$11149 ( \11329 , \11081 , \11107 );
or \U$11150 ( \11330 , \11327 , \11328 , \11329 );
xor \U$11151 ( \11331 , \11326 , \11330 );
or \U$11152 ( \11332 , \11113 , \11117 );
xor \U$11153 ( \11333 , \11331 , \11332 );
and \U$11154 ( \11334 , \10970 , \10974 );
and \U$11155 ( \11335 , \10974 , \10979 );
and \U$11156 ( \11336 , \10970 , \10979 );
or \U$11157 ( \11337 , \11334 , \11335 , \11336 );
and \U$11158 ( \11338 , \10984 , \10988 );
and \U$11159 ( \11339 , \10988 , \10993 );
and \U$11160 ( \11340 , \10984 , \10993 );
or \U$11161 ( \11341 , \11338 , \11339 , \11340 );
xor \U$11162 ( \11342 , \11337 , \11341 );
and \U$11163 ( \11343 , \10999 , \11003 );
and \U$11164 ( \11344 , \11003 , \11005 );
and \U$11165 ( \11345 , \10999 , \11005 );
or \U$11166 ( \11346 , \11343 , \11344 , \11345 );
xor \U$11167 ( \11347 , \11342 , \11346 );
xor \U$11168 ( \11348 , \11333 , \11347 );
and \U$11169 ( \11349 , \11138 , \11152 );
and \U$11170 ( \11350 , \11152 , \11167 );
and \U$11171 ( \11351 , \11138 , \11167 );
or \U$11172 ( \11352 , \11349 , \11350 , \11351 );
and \U$11173 ( \11353 , \11180 , \11194 );
xor \U$11174 ( \11354 , \11352 , \11353 );
and \U$11175 ( \11355 , \10584 , \195 );
not \U$11176 ( \11356 , \11355 );
xnor \U$11177 ( \11357 , \11356 , \202 );
and \U$11178 ( \11358 , \9897 , \215 );
and \U$11179 ( \11359 , \10206 , \213 );
nor \U$11180 ( \11360 , \11358 , \11359 );
xnor \U$11181 ( \11361 , \11360 , \222 );
xor \U$11182 ( \11362 , \11357 , \11361 );
and \U$11183 ( \11363 , \9169 , \230 );
and \U$11184 ( \11364 , \9465 , \228 );
nor \U$11185 ( \11365 , \11363 , \11364 );
xnor \U$11186 ( \11366 , \11365 , \237 );
xor \U$11187 ( \11367 , \11362 , \11366 );
xor \U$11188 ( \11368 , \11354 , \11367 );
and \U$11189 ( \11369 , \5469 , \1301 );
and \U$11190 ( \11370 , \5674 , \1246 );
nor \U$11191 ( \11371 , \11369 , \11370 );
xnor \U$11192 ( \11372 , \11371 , \1205 );
and \U$11193 ( \11373 , \4922 , \1578 );
and \U$11194 ( \11374 , \5156 , \1431 );
nor \U$11195 ( \11375 , \11373 , \11374 );
xnor \U$11196 ( \11376 , \11375 , \1436 );
xor \U$11197 ( \11377 , \11372 , \11376 );
and \U$11198 ( \11378 , \4654 , \1824 );
and \U$11199 ( \11379 , \4749 , \1739 );
nor \U$11200 ( \11380 , \11378 , \11379 );
xnor \U$11201 ( \11381 , \11380 , \1697 );
xor \U$11202 ( \11382 , \11377 , \11381 );
and \U$11203 ( \11383 , \6945 , \296 );
and \U$11204 ( \11384 , \7231 , \168 );
nor \U$11205 ( \11385 , \11383 , \11384 );
xnor \U$11206 ( \11386 , \11385 , \173 );
and \U$11207 ( \11387 , \6514 , \438 );
and \U$11208 ( \11388 , \6790 , \336 );
nor \U$11209 ( \11389 , \11387 , \11388 );
xnor \U$11210 ( \11390 , \11389 , \320 );
xor \U$11211 ( \11391 , \11386 , \11390 );
and \U$11212 ( \11392 , \6030 , \1086 );
and \U$11213 ( \11393 , \6281 , \508 );
nor \U$11214 ( \11394 , \11392 , \11393 );
xnor \U$11215 ( \11395 , \11394 , \487 );
xor \U$11216 ( \11396 , \11391 , \11395 );
xor \U$11217 ( \11397 , \11382 , \11396 );
and \U$11218 ( \11398 , \8652 , \245 );
and \U$11219 ( \11399 , \8835 , \243 );
nor \U$11220 ( \11400 , \11398 , \11399 );
xnor \U$11221 ( \11401 , \11400 , \252 );
and \U$11222 ( \11402 , \8057 , \141 );
and \U$11223 ( \11403 , \8349 , \139 );
nor \U$11224 ( \11404 , \11402 , \11403 );
xnor \U$11225 ( \11405 , \11404 , \148 );
xor \U$11226 ( \11406 , \11401 , \11405 );
and \U$11227 ( \11407 , \7556 , \156 );
and \U$11228 ( \11408 , \7700 , \154 );
nor \U$11229 ( \11409 , \11407 , \11408 );
xnor \U$11230 ( \11410 , \11409 , \163 );
xor \U$11231 ( \11411 , \11406 , \11410 );
xor \U$11232 ( \11412 , \11397 , \11411 );
and \U$11233 ( \11413 , \3037 , \3103 );
and \U$11234 ( \11414 , \3143 , \2934 );
nor \U$11235 ( \11415 , \11413 , \11414 );
xnor \U$11236 ( \11416 , \11415 , \2839 );
and \U$11237 ( \11417 , \2757 , \3357 );
and \U$11238 ( \11418 , \2826 , \3255 );
nor \U$11239 ( \11419 , \11417 , \11418 );
xnor \U$11240 ( \11420 , \11419 , \3156 );
xor \U$11241 ( \11421 , \11416 , \11420 );
and \U$11242 ( \11422 , \2366 , \3813 );
and \U$11243 ( \11423 , \2521 , \3557 );
nor \U$11244 ( \11424 , \11422 , \11423 );
xnor \U$11245 ( \11425 , \11424 , \3562 );
xor \U$11246 ( \11426 , \11421 , \11425 );
and \U$11247 ( \11427 , \4160 , \2121 );
and \U$11248 ( \11428 , \4364 , \2008 );
nor \U$11249 ( \11429 , \11427 , \11428 );
xnor \U$11250 ( \11430 , \11429 , \1961 );
and \U$11251 ( \11431 , \3736 , \2400 );
and \U$11252 ( \11432 , \3912 , \2246 );
nor \U$11253 ( \11433 , \11431 , \11432 );
xnor \U$11254 ( \11434 , \11433 , \2195 );
xor \U$11255 ( \11435 , \11430 , \11434 );
and \U$11256 ( \11436 , \3395 , \2669 );
and \U$11257 ( \11437 , \3646 , \2538 );
nor \U$11258 ( \11438 , \11436 , \11437 );
xnor \U$11259 ( \11439 , \11438 , \2534 );
xor \U$11260 ( \11440 , \11435 , \11439 );
xor \U$11261 ( \11441 , \11426 , \11440 );
and \U$11262 ( \11442 , \2090 , \4132 );
and \U$11263 ( \11443 , \2182 , \4012 );
nor \U$11264 ( \11444 , \11442 , \11443 );
xnor \U$11265 ( \11445 , \11444 , \3925 );
and \U$11266 ( \11446 , \1802 , \4581 );
and \U$11267 ( \11447 , \1948 , \4424 );
nor \U$11268 ( \11448 , \11446 , \11447 );
xnor \U$11269 ( \11449 , \11448 , \4377 );
xor \U$11270 ( \11450 , \11445 , \11449 );
and \U$11271 ( \11451 , \1601 , \5011 );
and \U$11272 ( \11452 , \1684 , \4878 );
nor \U$11273 ( \11453 , \11451 , \11452 );
xnor \U$11274 ( \11454 , \11453 , \4762 );
xor \U$11275 ( \11455 , \11450 , \11454 );
xor \U$11276 ( \11456 , \11441 , \11455 );
xor \U$11277 ( \11457 , \11412 , \11456 );
and \U$11278 ( \11458 , \261 , \7055 );
and \U$11279 ( \11459 , \307 , \6675 );
nor \U$11280 ( \11460 , \11458 , \11459 );
xnor \U$11281 ( \11461 , \11460 , \6680 );
and \U$11282 ( \11462 , \178 , \7489 );
and \U$11283 ( \11463 , \185 , \7137 );
nor \U$11284 ( \11464 , \11462 , \11463 );
xnor \U$11285 ( \11465 , \11464 , \7142 );
xor \U$11286 ( \11466 , \11461 , \11465 );
and \U$11287 ( \11467 , \189 , \8019 );
and \U$11288 ( \11468 , \197 , \7830 );
nor \U$11289 ( \11469 , \11467 , \11468 );
xnor \U$11290 ( \11470 , \11469 , \7713 );
xor \U$11291 ( \11471 , \11466 , \11470 );
and \U$11292 ( \11472 , \209 , \8540 );
and \U$11293 ( \11473 , \217 , \8292 );
nor \U$11294 ( \11474 , \11472 , \11473 );
xnor \U$11295 ( \11475 , \11474 , \8297 );
and \U$11296 ( \11476 , \224 , \9333 );
and \U$11297 ( \11477 , \232 , \9006 );
nor \U$11298 ( \11478 , \11476 , \11477 );
xnor \U$11299 ( \11479 , \11478 , \8848 );
xor \U$11300 ( \11480 , \11475 , \11479 );
and \U$11301 ( \11481 , \240 , \9765 );
and \U$11302 ( \11482 , \247 , \9644 );
nor \U$11303 ( \11483 , \11481 , \11482 );
xnor \U$11304 ( \11484 , \11483 , \9478 );
xor \U$11305 ( \11485 , \11480 , \11484 );
xor \U$11306 ( \11486 , \11471 , \11485 );
and \U$11307 ( \11487 , \1333 , \5485 );
and \U$11308 ( \11488 , \1484 , \5275 );
nor \U$11309 ( \11489 , \11487 , \11488 );
xnor \U$11310 ( \11490 , \11489 , \5169 );
and \U$11311 ( \11491 , \1147 , \5996 );
and \U$11312 ( \11492 , \1192 , \5695 );
nor \U$11313 ( \11493 , \11491 , \11492 );
xnor \U$11314 ( \11494 , \11493 , \5687 );
xor \U$11315 ( \11495 , \11490 , \11494 );
and \U$11316 ( \11496 , \412 , \6401 );
and \U$11317 ( \11497 , \474 , \6143 );
nor \U$11318 ( \11498 , \11496 , \11497 );
xnor \U$11319 ( \11499 , \11498 , \6148 );
xor \U$11320 ( \11500 , \11495 , \11499 );
xor \U$11321 ( \11501 , \11486 , \11500 );
xor \U$11322 ( \11502 , \11457 , \11501 );
xor \U$11323 ( \11503 , \11368 , \11502 );
and \U$11324 ( \11504 , \11027 , \11031 );
and \U$11325 ( \11505 , \11031 , \11036 );
and \U$11326 ( \11506 , \11027 , \11036 );
or \U$11327 ( \11507 , \11504 , \11505 , \11506 );
and \U$11328 ( \11508 , \11041 , \11045 );
and \U$11329 ( \11509 , \11045 , \11050 );
and \U$11330 ( \11510 , \11041 , \11050 );
or \U$11331 ( \11511 , \11508 , \11509 , \11510 );
xor \U$11332 ( \11512 , \11507 , \11511 );
and \U$11333 ( \11513 , \11097 , \11101 );
and \U$11334 ( \11514 , \11101 , \11106 );
and \U$11335 ( \11515 , \11097 , \11106 );
or \U$11336 ( \11516 , \11513 , \11514 , \11515 );
xor \U$11337 ( \11517 , \11512 , \11516 );
and \U$11338 ( \11518 , \11128 , \11132 );
and \U$11339 ( \11519 , \11132 , \11137 );
and \U$11340 ( \11520 , \11128 , \11137 );
or \U$11341 ( \11521 , \11518 , \11519 , \11520 );
and \U$11342 ( \11522 , \11056 , \11060 );
and \U$11343 ( \11523 , \11060 , \11065 );
and \U$11344 ( \11524 , \11056 , \11065 );
or \U$11345 ( \11525 , \11522 , \11523 , \11524 );
xor \U$11346 ( \11526 , \11521 , \11525 );
and \U$11347 ( \11527 , \11157 , \11161 );
and \U$11348 ( \11528 , \11161 , \11166 );
and \U$11349 ( \11529 , \11157 , \11166 );
or \U$11350 ( \11530 , \11527 , \11528 , \11529 );
xor \U$11351 ( \11531 , \11526 , \11530 );
xor \U$11352 ( \11532 , \11517 , \11531 );
and \U$11353 ( \11533 , \11071 , \11075 );
and \U$11354 ( \11534 , \11075 , \11080 );
and \U$11355 ( \11535 , \11071 , \11080 );
or \U$11356 ( \11536 , \11533 , \11534 , \11535 );
and \U$11357 ( \11537 , \11085 , \11089 );
and \U$11358 ( \11538 , \11089 , \11091 );
and \U$11359 ( \11539 , \11085 , \11091 );
or \U$11360 ( \11540 , \11537 , \11538 , \11539 );
xor \U$11361 ( \11541 , \11536 , \11540 );
and \U$11362 ( \11542 , \134 , \10408 );
and \U$11363 ( \11543 , \143 , \10116 );
nor \U$11364 ( \11544 , \11542 , \11543 );
xnor \U$11365 ( \11545 , \11544 , \10121 );
and \U$11366 ( \11546 , \158 , \10118 );
xnor \U$11367 ( \11547 , \11545 , \11546 );
xor \U$11368 ( \11548 , \11541 , \11547 );
xor \U$11369 ( \11549 , \11532 , \11548 );
xor \U$11370 ( \11550 , \11503 , \11549 );
xor \U$11371 ( \11551 , \11348 , \11550 );
xor \U$11372 ( \11552 , \11322 , \11551 );
xor \U$11373 ( \11553 , \11293 , \11552 );
xor \U$11374 ( \11554 , \11254 , \11553 );
and \U$11375 ( \11555 , \10934 , \11199 );
and \U$11376 ( \11556 , \11199 , \11239 );
and \U$11377 ( \11557 , \10934 , \11239 );
or \U$11378 ( \11558 , \11555 , \11556 , \11557 );
xor \U$11379 ( \11559 , \11554 , \11558 );
and \U$11380 ( \11560 , \11240 , \11241 );
and \U$11381 ( \11561 , \11242 , \11245 );
or \U$11382 ( \11562 , \11560 , \11561 );
xor \U$11383 ( \11563 , \11559 , \11562 );
buf g5517_GF_PartitionCandidate( \11564_nG5517 , \11563 );
buf \U$11384 ( \11565 , \11564_nG5517 );
and \U$11385 ( \11566 , \11258 , \11292 );
and \U$11386 ( \11567 , \11292 , \11552 );
and \U$11387 ( \11568 , \11258 , \11552 );
or \U$11388 ( \11569 , \11566 , \11567 , \11568 );
and \U$11389 ( \11570 , \11262 , \11266 );
and \U$11390 ( \11571 , \11266 , \11291 );
and \U$11391 ( \11572 , \11262 , \11291 );
or \U$11392 ( \11573 , \11570 , \11571 , \11572 );
and \U$11393 ( \11574 , \11307 , \11321 );
and \U$11394 ( \11575 , \11321 , \11551 );
and \U$11395 ( \11576 , \11307 , \11551 );
or \U$11396 ( \11577 , \11574 , \11575 , \11576 );
xor \U$11397 ( \11578 , \11573 , \11577 );
and \U$11398 ( \11579 , \11280 , \11284 );
and \U$11399 ( \11580 , \11284 , \11289 );
and \U$11400 ( \11581 , \11280 , \11289 );
or \U$11401 ( \11582 , \11579 , \11580 , \11581 );
and \U$11402 ( \11583 , \11507 , \11511 );
and \U$11403 ( \11584 , \11511 , \11516 );
and \U$11404 ( \11585 , \11507 , \11516 );
or \U$11405 ( \11586 , \11583 , \11584 , \11585 );
xor \U$11406 ( \11587 , \11582 , \11586 );
and \U$11407 ( \11588 , \11521 , \11525 );
and \U$11408 ( \11589 , \11525 , \11530 );
and \U$11409 ( \11590 , \11521 , \11530 );
or \U$11410 ( \11591 , \11588 , \11589 , \11590 );
xor \U$11411 ( \11592 , \11587 , \11591 );
and \U$11412 ( \11593 , \11412 , \11456 );
and \U$11413 ( \11594 , \11456 , \11501 );
and \U$11414 ( \11595 , \11412 , \11501 );
or \U$11415 ( \11596 , \11593 , \11594 , \11595 );
and \U$11416 ( \11597 , \11517 , \11531 );
and \U$11417 ( \11598 , \11531 , \11548 );
and \U$11418 ( \11599 , \11517 , \11548 );
or \U$11419 ( \11600 , \11597 , \11598 , \11599 );
xor \U$11420 ( \11601 , \11596 , \11600 );
and \U$11421 ( \11602 , \11386 , \11390 );
and \U$11422 ( \11603 , \11390 , \11395 );
and \U$11423 ( \11604 , \11386 , \11395 );
or \U$11424 ( \11605 , \11602 , \11603 , \11604 );
and \U$11425 ( \11606 , \11357 , \11361 );
and \U$11426 ( \11607 , \11361 , \11366 );
and \U$11427 ( \11608 , \11357 , \11366 );
or \U$11428 ( \11609 , \11606 , \11607 , \11608 );
xor \U$11429 ( \11610 , \11605 , \11609 );
and \U$11430 ( \11611 , \11401 , \11405 );
and \U$11431 ( \11612 , \11405 , \11410 );
and \U$11432 ( \11613 , \11401 , \11410 );
or \U$11433 ( \11614 , \11611 , \11612 , \11613 );
xor \U$11434 ( \11615 , \11610 , \11614 );
and \U$11435 ( \11616 , \11461 , \11465 );
and \U$11436 ( \11617 , \11465 , \11470 );
and \U$11437 ( \11618 , \11461 , \11470 );
or \U$11438 ( \11619 , \11616 , \11617 , \11618 );
and \U$11439 ( \11620 , \11445 , \11449 );
and \U$11440 ( \11621 , \11449 , \11454 );
and \U$11441 ( \11622 , \11445 , \11454 );
or \U$11442 ( \11623 , \11620 , \11621 , \11622 );
xor \U$11443 ( \11624 , \11619 , \11623 );
and \U$11444 ( \11625 , \11490 , \11494 );
and \U$11445 ( \11626 , \11494 , \11499 );
and \U$11446 ( \11627 , \11490 , \11499 );
or \U$11447 ( \11628 , \11625 , \11626 , \11627 );
xor \U$11448 ( \11629 , \11624 , \11628 );
xor \U$11449 ( \11630 , \11615 , \11629 );
and \U$11450 ( \11631 , \11372 , \11376 );
and \U$11451 ( \11632 , \11376 , \11381 );
and \U$11452 ( \11633 , \11372 , \11381 );
or \U$11453 ( \11634 , \11631 , \11632 , \11633 );
and \U$11454 ( \11635 , \11416 , \11420 );
and \U$11455 ( \11636 , \11420 , \11425 );
and \U$11456 ( \11637 , \11416 , \11425 );
or \U$11457 ( \11638 , \11635 , \11636 , \11637 );
xor \U$11458 ( \11639 , \11634 , \11638 );
and \U$11459 ( \11640 , \11430 , \11434 );
and \U$11460 ( \11641 , \11434 , \11439 );
and \U$11461 ( \11642 , \11430 , \11439 );
or \U$11462 ( \11643 , \11640 , \11641 , \11642 );
xor \U$11463 ( \11644 , \11639 , \11643 );
xor \U$11464 ( \11645 , \11630 , \11644 );
xor \U$11465 ( \11646 , \11601 , \11645 );
xor \U$11466 ( \11647 , \11592 , \11646 );
and \U$11467 ( \11648 , \11426 , \11440 );
and \U$11468 ( \11649 , \11440 , \11455 );
and \U$11469 ( \11650 , \11426 , \11455 );
or \U$11470 ( \11651 , \11648 , \11649 , \11650 );
and \U$11471 ( \11652 , \11471 , \11485 );
and \U$11472 ( \11653 , \11485 , \11500 );
and \U$11473 ( \11654 , \11471 , \11500 );
or \U$11474 ( \11655 , \11652 , \11653 , \11654 );
xor \U$11475 ( \11656 , \11651 , \11655 );
and \U$11476 ( \11657 , \11536 , \11540 );
and \U$11477 ( \11658 , \11540 , \11547 );
and \U$11478 ( \11659 , \11536 , \11547 );
or \U$11479 ( \11660 , \11657 , \11658 , \11659 );
xor \U$11480 ( \11661 , \11656 , \11660 );
and \U$11481 ( \11662 , \11475 , \11479 );
and \U$11482 ( \11663 , \11479 , \11484 );
and \U$11483 ( \11664 , \11475 , \11484 );
or \U$11484 ( \11665 , \11662 , \11663 , \11664 );
or \U$11485 ( \11666 , \11545 , \11546 );
xor \U$11486 ( \11667 , \11665 , \11666 );
and \U$11487 ( \11668 , \143 , \10408 );
and \U$11488 ( \11669 , \240 , \10116 );
nor \U$11489 ( \11670 , \11668 , \11669 );
xnor \U$11490 ( \11671 , \11670 , \10121 );
xor \U$11491 ( \11672 , \11667 , \11671 );
and \U$11492 ( \11673 , \134 , \10118 );
and \U$11493 ( \11674 , \307 , \7055 );
and \U$11494 ( \11675 , \412 , \6675 );
nor \U$11495 ( \11676 , \11674 , \11675 );
xnor \U$11496 ( \11677 , \11676 , \6680 );
and \U$11497 ( \11678 , \185 , \7489 );
and \U$11498 ( \11679 , \261 , \7137 );
nor \U$11499 ( \11680 , \11678 , \11679 );
xnor \U$11500 ( \11681 , \11680 , \7142 );
xor \U$11501 ( \11682 , \11677 , \11681 );
and \U$11502 ( \11683 , \197 , \8019 );
and \U$11503 ( \11684 , \178 , \7830 );
nor \U$11504 ( \11685 , \11683 , \11684 );
xnor \U$11505 ( \11686 , \11685 , \7713 );
xor \U$11506 ( \11687 , \11682 , \11686 );
xor \U$11507 ( \11688 , \11673 , \11687 );
and \U$11508 ( \11689 , \217 , \8540 );
and \U$11509 ( \11690 , \189 , \8292 );
nor \U$11510 ( \11691 , \11689 , \11690 );
xnor \U$11511 ( \11692 , \11691 , \8297 );
and \U$11512 ( \11693 , \232 , \9333 );
and \U$11513 ( \11694 , \209 , \9006 );
nor \U$11514 ( \11695 , \11693 , \11694 );
xnor \U$11515 ( \11696 , \11695 , \8848 );
xor \U$11516 ( \11697 , \11692 , \11696 );
and \U$11517 ( \11698 , \247 , \9765 );
and \U$11518 ( \11699 , \224 , \9644 );
nor \U$11519 ( \11700 , \11698 , \11699 );
xnor \U$11520 ( \11701 , \11700 , \9478 );
xor \U$11521 ( \11702 , \11697 , \11701 );
xor \U$11522 ( \11703 , \11688 , \11702 );
xor \U$11523 ( \11704 , \11672 , \11703 );
and \U$11524 ( \11705 , \3143 , \3103 );
and \U$11525 ( \11706 , \3395 , \2934 );
nor \U$11526 ( \11707 , \11705 , \11706 );
xnor \U$11527 ( \11708 , \11707 , \2839 );
and \U$11528 ( \11709 , \2826 , \3357 );
and \U$11529 ( \11710 , \3037 , \3255 );
nor \U$11530 ( \11711 , \11709 , \11710 );
xnor \U$11531 ( \11712 , \11711 , \3156 );
xor \U$11532 ( \11713 , \11708 , \11712 );
and \U$11533 ( \11714 , \2521 , \3813 );
and \U$11534 ( \11715 , \2757 , \3557 );
nor \U$11535 ( \11716 , \11714 , \11715 );
xnor \U$11536 ( \11717 , \11716 , \3562 );
xor \U$11537 ( \11718 , \11713 , \11717 );
and \U$11538 ( \11719 , \1484 , \5485 );
and \U$11539 ( \11720 , \1601 , \5275 );
nor \U$11540 ( \11721 , \11719 , \11720 );
xnor \U$11541 ( \11722 , \11721 , \5169 );
and \U$11542 ( \11723 , \1192 , \5996 );
and \U$11543 ( \11724 , \1333 , \5695 );
nor \U$11544 ( \11725 , \11723 , \11724 );
xnor \U$11545 ( \11726 , \11725 , \5687 );
xor \U$11546 ( \11727 , \11722 , \11726 );
and \U$11547 ( \11728 , \474 , \6401 );
and \U$11548 ( \11729 , \1147 , \6143 );
nor \U$11549 ( \11730 , \11728 , \11729 );
xnor \U$11550 ( \11731 , \11730 , \6148 );
xor \U$11551 ( \11732 , \11727 , \11731 );
xor \U$11552 ( \11733 , \11718 , \11732 );
and \U$11553 ( \11734 , \2182 , \4132 );
and \U$11554 ( \11735 , \2366 , \4012 );
nor \U$11555 ( \11736 , \11734 , \11735 );
xnor \U$11556 ( \11737 , \11736 , \3925 );
and \U$11557 ( \11738 , \1948 , \4581 );
and \U$11558 ( \11739 , \2090 , \4424 );
nor \U$11559 ( \11740 , \11738 , \11739 );
xnor \U$11560 ( \11741 , \11740 , \4377 );
xor \U$11561 ( \11742 , \11737 , \11741 );
and \U$11562 ( \11743 , \1684 , \5011 );
and \U$11563 ( \11744 , \1802 , \4878 );
nor \U$11564 ( \11745 , \11743 , \11744 );
xnor \U$11565 ( \11746 , \11745 , \4762 );
xor \U$11566 ( \11747 , \11742 , \11746 );
xor \U$11567 ( \11748 , \11733 , \11747 );
xor \U$11568 ( \11749 , \11704 , \11748 );
xor \U$11569 ( \11750 , \11661 , \11749 );
and \U$11570 ( \11751 , \11382 , \11396 );
and \U$11571 ( \11752 , \11396 , \11411 );
and \U$11572 ( \11753 , \11382 , \11411 );
or \U$11573 ( \11754 , \11751 , \11752 , \11753 );
and \U$11574 ( \11755 , \7231 , \296 );
and \U$11575 ( \11756 , \7556 , \168 );
nor \U$11576 ( \11757 , \11755 , \11756 );
xnor \U$11577 ( \11758 , \11757 , \173 );
and \U$11578 ( \11759 , \6790 , \438 );
and \U$11579 ( \11760 , \6945 , \336 );
nor \U$11580 ( \11761 , \11759 , \11760 );
xnor \U$11581 ( \11762 , \11761 , \320 );
xor \U$11582 ( \11763 , \11758 , \11762 );
and \U$11583 ( \11764 , \6281 , \1086 );
and \U$11584 ( \11765 , \6514 , \508 );
nor \U$11585 ( \11766 , \11764 , \11765 );
xnor \U$11586 ( \11767 , \11766 , \487 );
xor \U$11587 ( \11768 , \11763 , \11767 );
and \U$11588 ( \11769 , \4364 , \2121 );
and \U$11589 ( \11770 , \4654 , \2008 );
nor \U$11590 ( \11771 , \11769 , \11770 );
xnor \U$11591 ( \11772 , \11771 , \1961 );
and \U$11592 ( \11773 , \3912 , \2400 );
and \U$11593 ( \11774 , \4160 , \2246 );
nor \U$11594 ( \11775 , \11773 , \11774 );
xnor \U$11595 ( \11776 , \11775 , \2195 );
xor \U$11596 ( \11777 , \11772 , \11776 );
and \U$11597 ( \11778 , \3646 , \2669 );
and \U$11598 ( \11779 , \3736 , \2538 );
nor \U$11599 ( \11780 , \11778 , \11779 );
xnor \U$11600 ( \11781 , \11780 , \2534 );
xor \U$11601 ( \11782 , \11777 , \11781 );
xor \U$11602 ( \11783 , \11768 , \11782 );
and \U$11603 ( \11784 , \5674 , \1301 );
and \U$11604 ( \11785 , \6030 , \1246 );
nor \U$11605 ( \11786 , \11784 , \11785 );
xnor \U$11606 ( \11787 , \11786 , \1205 );
and \U$11607 ( \11788 , \5156 , \1578 );
and \U$11608 ( \11789 , \5469 , \1431 );
nor \U$11609 ( \11790 , \11788 , \11789 );
xnor \U$11610 ( \11791 , \11790 , \1436 );
xor \U$11611 ( \11792 , \11787 , \11791 );
and \U$11612 ( \11793 , \4749 , \1824 );
and \U$11613 ( \11794 , \4922 , \1739 );
nor \U$11614 ( \11795 , \11793 , \11794 );
xnor \U$11615 ( \11796 , \11795 , \1697 );
xor \U$11616 ( \11797 , \11792 , \11796 );
xor \U$11617 ( \11798 , \11783 , \11797 );
xor \U$11618 ( \11799 , \11754 , \11798 );
and \U$11619 ( \11800 , \8835 , \245 );
and \U$11620 ( \11801 , \9169 , \243 );
nor \U$11621 ( \11802 , \11800 , \11801 );
xnor \U$11622 ( \11803 , \11802 , \252 );
and \U$11623 ( \11804 , \8349 , \141 );
and \U$11624 ( \11805 , \8652 , \139 );
nor \U$11625 ( \11806 , \11804 , \11805 );
xnor \U$11626 ( \11807 , \11806 , \148 );
xor \U$11627 ( \11808 , \11803 , \11807 );
and \U$11628 ( \11809 , \7700 , \156 );
and \U$11629 ( \11810 , \8057 , \154 );
nor \U$11630 ( \11811 , \11809 , \11810 );
xnor \U$11631 ( \11812 , \11811 , \163 );
xor \U$11632 ( \11813 , \11808 , \11812 );
not \U$11633 ( \11814 , \202 );
and \U$11634 ( \11815 , \10206 , \215 );
and \U$11635 ( \11816 , \10584 , \213 );
nor \U$11636 ( \11817 , \11815 , \11816 );
xnor \U$11637 ( \11818 , \11817 , \222 );
xor \U$11638 ( \11819 , \11814 , \11818 );
and \U$11639 ( \11820 , \9465 , \230 );
and \U$11640 ( \11821 , \9897 , \228 );
nor \U$11641 ( \11822 , \11820 , \11821 );
xnor \U$11642 ( \11823 , \11822 , \237 );
xor \U$11643 ( \11824 , \11819 , \11823 );
xor \U$11644 ( \11825 , \11813 , \11824 );
xor \U$11645 ( \11826 , \11799 , \11825 );
xor \U$11646 ( \11827 , \11750 , \11826 );
xor \U$11647 ( \11828 , \11647 , \11827 );
xor \U$11648 ( \11829 , \11578 , \11828 );
xor \U$11649 ( \11830 , \11569 , \11829 );
and \U$11650 ( \11831 , \11297 , \11301 );
and \U$11651 ( \11832 , \11301 , \11306 );
and \U$11652 ( \11833 , \11297 , \11306 );
or \U$11653 ( \11834 , \11831 , \11832 , \11833 );
and \U$11654 ( \11835 , \11271 , \11275 );
and \U$11655 ( \11836 , \11275 , \11290 );
and \U$11656 ( \11837 , \11271 , \11290 );
or \U$11657 ( \11838 , \11835 , \11836 , \11837 );
xor \U$11658 ( \11839 , \11834 , \11838 );
and \U$11659 ( \11840 , \11368 , \11502 );
and \U$11660 ( \11841 , \11502 , \11549 );
and \U$11661 ( \11842 , \11368 , \11549 );
or \U$11662 ( \11843 , \11840 , \11841 , \11842 );
xor \U$11663 ( \11844 , \11839 , \11843 );
and \U$11664 ( \11845 , \11311 , \11315 );
and \U$11665 ( \11846 , \11315 , \11320 );
and \U$11666 ( \11847 , \11311 , \11320 );
or \U$11667 ( \11848 , \11845 , \11846 , \11847 );
and \U$11668 ( \11849 , \11333 , \11347 );
and \U$11669 ( \11850 , \11347 , \11550 );
and \U$11670 ( \11851 , \11333 , \11550 );
or \U$11671 ( \11852 , \11849 , \11850 , \11851 );
xor \U$11672 ( \11853 , \11848 , \11852 );
and \U$11673 ( \11854 , \11326 , \11330 );
and \U$11674 ( \11855 , \11330 , \11332 );
and \U$11675 ( \11856 , \11326 , \11332 );
or \U$11676 ( \11857 , \11854 , \11855 , \11856 );
and \U$11677 ( \11858 , \11337 , \11341 );
and \U$11678 ( \11859 , \11341 , \11346 );
and \U$11679 ( \11860 , \11337 , \11346 );
or \U$11680 ( \11861 , \11858 , \11859 , \11860 );
xor \U$11681 ( \11862 , \11857 , \11861 );
and \U$11682 ( \11863 , \11352 , \11353 );
and \U$11683 ( \11864 , \11353 , \11367 );
and \U$11684 ( \11865 , \11352 , \11367 );
or \U$11685 ( \11866 , \11863 , \11864 , \11865 );
xor \U$11686 ( \11867 , \11862 , \11866 );
xor \U$11687 ( \11868 , \11853 , \11867 );
xor \U$11688 ( \11869 , \11844 , \11868 );
xor \U$11689 ( \11870 , \11830 , \11869 );
and \U$11690 ( \11871 , \11252 , \11253 );
and \U$11691 ( \11872 , \11253 , \11553 );
and \U$11692 ( \11873 , \11252 , \11553 );
or \U$11693 ( \11874 , \11871 , \11872 , \11873 );
xor \U$11694 ( \11875 , \11870 , \11874 );
and \U$11695 ( \11876 , \11554 , \11558 );
and \U$11696 ( \11877 , \11559 , \11562 );
or \U$11697 ( \11878 , \11876 , \11877 );
xor \U$11698 ( \11879 , \11875 , \11878 );
buf g5515_GF_PartitionCandidate( \11880_nG5515 , \11879 );
buf \U$11699 ( \11881 , \11880_nG5515 );
and \U$11700 ( \11882 , \11573 , \11577 );
and \U$11701 ( \11883 , \11577 , \11828 );
and \U$11702 ( \11884 , \11573 , \11828 );
or \U$11703 ( \11885 , \11882 , \11883 , \11884 );
and \U$11704 ( \11886 , \11844 , \11868 );
xor \U$11705 ( \11887 , \11885 , \11886 );
and \U$11706 ( \11888 , \11848 , \11852 );
and \U$11707 ( \11889 , \11852 , \11867 );
and \U$11708 ( \11890 , \11848 , \11867 );
or \U$11709 ( \11891 , \11888 , \11889 , \11890 );
and \U$11710 ( \11892 , \11834 , \11838 );
and \U$11711 ( \11893 , \11838 , \11843 );
and \U$11712 ( \11894 , \11834 , \11843 );
or \U$11713 ( \11895 , \11892 , \11893 , \11894 );
and \U$11714 ( \11896 , \11592 , \11646 );
and \U$11715 ( \11897 , \11646 , \11827 );
and \U$11716 ( \11898 , \11592 , \11827 );
or \U$11717 ( \11899 , \11896 , \11897 , \11898 );
xor \U$11718 ( \11900 , \11895 , \11899 );
and \U$11719 ( \11901 , \11651 , \11655 );
and \U$11720 ( \11902 , \11655 , \11660 );
and \U$11721 ( \11903 , \11651 , \11660 );
or \U$11722 ( \11904 , \11901 , \11902 , \11903 );
and \U$11723 ( \11905 , \11582 , \11586 );
and \U$11724 ( \11906 , \11586 , \11591 );
and \U$11725 ( \11907 , \11582 , \11591 );
or \U$11726 ( \11908 , \11905 , \11906 , \11907 );
xor \U$11727 ( \11909 , \11904 , \11908 );
and \U$11728 ( \11910 , \11754 , \11798 );
and \U$11729 ( \11911 , \11798 , \11825 );
and \U$11730 ( \11912 , \11754 , \11825 );
or \U$11731 ( \11913 , \11910 , \11911 , \11912 );
xor \U$11732 ( \11914 , \11909 , \11913 );
xor \U$11733 ( \11915 , \11900 , \11914 );
xor \U$11734 ( \11916 , \11891 , \11915 );
and \U$11735 ( \11917 , \11857 , \11861 );
and \U$11736 ( \11918 , \11861 , \11866 );
and \U$11737 ( \11919 , \11857 , \11866 );
or \U$11738 ( \11920 , \11917 , \11918 , \11919 );
and \U$11739 ( \11921 , \11596 , \11600 );
and \U$11740 ( \11922 , \11600 , \11645 );
and \U$11741 ( \11923 , \11596 , \11645 );
or \U$11742 ( \11924 , \11921 , \11922 , \11923 );
xor \U$11743 ( \11925 , \11920 , \11924 );
and \U$11744 ( \11926 , \11661 , \11749 );
and \U$11745 ( \11927 , \11749 , \11826 );
and \U$11746 ( \11928 , \11661 , \11826 );
or \U$11747 ( \11929 , \11926 , \11927 , \11928 );
xor \U$11748 ( \11930 , \11925 , \11929 );
and \U$11749 ( \11931 , \11605 , \11609 );
and \U$11750 ( \11932 , \11609 , \11614 );
and \U$11751 ( \11933 , \11605 , \11614 );
or \U$11752 ( \11934 , \11931 , \11932 , \11933 );
and \U$11753 ( \11935 , \11619 , \11623 );
and \U$11754 ( \11936 , \11623 , \11628 );
and \U$11755 ( \11937 , \11619 , \11628 );
or \U$11756 ( \11938 , \11935 , \11936 , \11937 );
xor \U$11757 ( \11939 , \11934 , \11938 );
and \U$11758 ( \11940 , \11634 , \11638 );
and \U$11759 ( \11941 , \11638 , \11643 );
and \U$11760 ( \11942 , \11634 , \11643 );
or \U$11761 ( \11943 , \11940 , \11941 , \11942 );
xor \U$11762 ( \11944 , \11939 , \11943 );
and \U$11763 ( \11945 , \11615 , \11629 );
and \U$11764 ( \11946 , \11629 , \11644 );
and \U$11765 ( \11947 , \11615 , \11644 );
or \U$11766 ( \11948 , \11945 , \11946 , \11947 );
and \U$11767 ( \11949 , \11672 , \11703 );
and \U$11768 ( \11950 , \11703 , \11748 );
and \U$11769 ( \11951 , \11672 , \11748 );
or \U$11770 ( \11952 , \11949 , \11950 , \11951 );
xor \U$11771 ( \11953 , \11948 , \11952 );
and \U$11772 ( \11954 , \11708 , \11712 );
and \U$11773 ( \11955 , \11712 , \11717 );
and \U$11774 ( \11956 , \11708 , \11717 );
or \U$11775 ( \11957 , \11954 , \11955 , \11956 );
and \U$11776 ( \11958 , \11772 , \11776 );
and \U$11777 ( \11959 , \11776 , \11781 );
and \U$11778 ( \11960 , \11772 , \11781 );
or \U$11779 ( \11961 , \11958 , \11959 , \11960 );
xor \U$11780 ( \11962 , \11957 , \11961 );
and \U$11781 ( \11963 , \11787 , \11791 );
and \U$11782 ( \11964 , \11791 , \11796 );
and \U$11783 ( \11965 , \11787 , \11796 );
or \U$11784 ( \11966 , \11963 , \11964 , \11965 );
xor \U$11785 ( \11967 , \11962 , \11966 );
and \U$11786 ( \11968 , \11758 , \11762 );
and \U$11787 ( \11969 , \11762 , \11767 );
and \U$11788 ( \11970 , \11758 , \11767 );
or \U$11789 ( \11971 , \11968 , \11969 , \11970 );
and \U$11790 ( \11972 , \11803 , \11807 );
and \U$11791 ( \11973 , \11807 , \11812 );
and \U$11792 ( \11974 , \11803 , \11812 );
or \U$11793 ( \11975 , \11972 , \11973 , \11974 );
xor \U$11794 ( \11976 , \11971 , \11975 );
and \U$11795 ( \11977 , \11814 , \11818 );
and \U$11796 ( \11978 , \11818 , \11823 );
and \U$11797 ( \11979 , \11814 , \11823 );
or \U$11798 ( \11980 , \11977 , \11978 , \11979 );
xor \U$11799 ( \11981 , \11976 , \11980 );
xor \U$11800 ( \11982 , \11967 , \11981 );
and \U$11801 ( \11983 , \11677 , \11681 );
and \U$11802 ( \11984 , \11681 , \11686 );
and \U$11803 ( \11985 , \11677 , \11686 );
or \U$11804 ( \11986 , \11983 , \11984 , \11985 );
and \U$11805 ( \11987 , \11722 , \11726 );
and \U$11806 ( \11988 , \11726 , \11731 );
and \U$11807 ( \11989 , \11722 , \11731 );
or \U$11808 ( \11990 , \11987 , \11988 , \11989 );
xor \U$11809 ( \11991 , \11986 , \11990 );
and \U$11810 ( \11992 , \11737 , \11741 );
and \U$11811 ( \11993 , \11741 , \11746 );
and \U$11812 ( \11994 , \11737 , \11746 );
or \U$11813 ( \11995 , \11992 , \11993 , \11994 );
xor \U$11814 ( \11996 , \11991 , \11995 );
xor \U$11815 ( \11997 , \11982 , \11996 );
xor \U$11816 ( \11998 , \11953 , \11997 );
xor \U$11817 ( \11999 , \11944 , \11998 );
and \U$11818 ( \12000 , \11665 , \11666 );
and \U$11819 ( \12001 , \11666 , \11671 );
and \U$11820 ( \12002 , \11665 , \11671 );
or \U$11821 ( \12003 , \12000 , \12001 , \12002 );
and \U$11822 ( \12004 , \11673 , \11687 );
and \U$11823 ( \12005 , \11687 , \11702 );
and \U$11824 ( \12006 , \11673 , \11702 );
or \U$11825 ( \12007 , \12004 , \12005 , \12006 );
xor \U$11826 ( \12008 , \12003 , \12007 );
and \U$11827 ( \12009 , \11718 , \11732 );
and \U$11828 ( \12010 , \11732 , \11747 );
and \U$11829 ( \12011 , \11718 , \11747 );
or \U$11830 ( \12012 , \12009 , \12010 , \12011 );
xor \U$11831 ( \12013 , \12008 , \12012 );
and \U$11832 ( \12014 , \11768 , \11782 );
and \U$11833 ( \12015 , \11782 , \11797 );
and \U$11834 ( \12016 , \11768 , \11797 );
or \U$11835 ( \12017 , \12014 , \12015 , \12016 );
and \U$11836 ( \12018 , \11813 , \11824 );
xor \U$11837 ( \12019 , \12017 , \12018 );
and \U$11838 ( \12020 , \10584 , \215 );
not \U$11839 ( \12021 , \12020 );
xnor \U$11840 ( \12022 , \12021 , \222 );
and \U$11841 ( \12023 , \9897 , \230 );
and \U$11842 ( \12024 , \10206 , \228 );
nor \U$11843 ( \12025 , \12023 , \12024 );
xnor \U$11844 ( \12026 , \12025 , \237 );
xor \U$11845 ( \12027 , \12022 , \12026 );
and \U$11846 ( \12028 , \9169 , \245 );
and \U$11847 ( \12029 , \9465 , \243 );
nor \U$11848 ( \12030 , \12028 , \12029 );
xnor \U$11849 ( \12031 , \12030 , \252 );
xor \U$11850 ( \12032 , \12027 , \12031 );
and \U$11851 ( \12033 , \6945 , \438 );
and \U$11852 ( \12034 , \7231 , \336 );
nor \U$11853 ( \12035 , \12033 , \12034 );
xnor \U$11854 ( \12036 , \12035 , \320 );
and \U$11855 ( \12037 , \6514 , \1086 );
and \U$11856 ( \12038 , \6790 , \508 );
nor \U$11857 ( \12039 , \12037 , \12038 );
xnor \U$11858 ( \12040 , \12039 , \487 );
xor \U$11859 ( \12041 , \12036 , \12040 );
and \U$11860 ( \12042 , \6030 , \1301 );
and \U$11861 ( \12043 , \6281 , \1246 );
nor \U$11862 ( \12044 , \12042 , \12043 );
xnor \U$11863 ( \12045 , \12044 , \1205 );
xor \U$11864 ( \12046 , \12041 , \12045 );
xor \U$11865 ( \12047 , \12032 , \12046 );
and \U$11866 ( \12048 , \8652 , \141 );
and \U$11867 ( \12049 , \8835 , \139 );
nor \U$11868 ( \12050 , \12048 , \12049 );
xnor \U$11869 ( \12051 , \12050 , \148 );
and \U$11870 ( \12052 , \8057 , \156 );
and \U$11871 ( \12053 , \8349 , \154 );
nor \U$11872 ( \12054 , \12052 , \12053 );
xnor \U$11873 ( \12055 , \12054 , \163 );
xor \U$11874 ( \12056 , \12051 , \12055 );
and \U$11875 ( \12057 , \7556 , \296 );
and \U$11876 ( \12058 , \7700 , \168 );
nor \U$11877 ( \12059 , \12057 , \12058 );
xnor \U$11878 ( \12060 , \12059 , \173 );
xor \U$11879 ( \12061 , \12056 , \12060 );
xor \U$11880 ( \12062 , \12047 , \12061 );
xor \U$11881 ( \12063 , \12019 , \12062 );
xor \U$11882 ( \12064 , \12013 , \12063 );
and \U$11883 ( \12065 , \5469 , \1578 );
and \U$11884 ( \12066 , \5674 , \1431 );
nor \U$11885 ( \12067 , \12065 , \12066 );
xnor \U$11886 ( \12068 , \12067 , \1436 );
and \U$11887 ( \12069 , \4922 , \1824 );
and \U$11888 ( \12070 , \5156 , \1739 );
nor \U$11889 ( \12071 , \12069 , \12070 );
xnor \U$11890 ( \12072 , \12071 , \1697 );
xor \U$11891 ( \12073 , \12068 , \12072 );
and \U$11892 ( \12074 , \4654 , \2121 );
and \U$11893 ( \12075 , \4749 , \2008 );
nor \U$11894 ( \12076 , \12074 , \12075 );
xnor \U$11895 ( \12077 , \12076 , \1961 );
xor \U$11896 ( \12078 , \12073 , \12077 );
and \U$11897 ( \12079 , \3037 , \3357 );
and \U$11898 ( \12080 , \3143 , \3255 );
nor \U$11899 ( \12081 , \12079 , \12080 );
xnor \U$11900 ( \12082 , \12081 , \3156 );
and \U$11901 ( \12083 , \2757 , \3813 );
and \U$11902 ( \12084 , \2826 , \3557 );
nor \U$11903 ( \12085 , \12083 , \12084 );
xnor \U$11904 ( \12086 , \12085 , \3562 );
xor \U$11905 ( \12087 , \12082 , \12086 );
and \U$11906 ( \12088 , \2366 , \4132 );
and \U$11907 ( \12089 , \2521 , \4012 );
nor \U$11908 ( \12090 , \12088 , \12089 );
xnor \U$11909 ( \12091 , \12090 , \3925 );
xor \U$11910 ( \12092 , \12087 , \12091 );
xor \U$11911 ( \12093 , \12078 , \12092 );
and \U$11912 ( \12094 , \4160 , \2400 );
and \U$11913 ( \12095 , \4364 , \2246 );
nor \U$11914 ( \12096 , \12094 , \12095 );
xnor \U$11915 ( \12097 , \12096 , \2195 );
and \U$11916 ( \12098 , \3736 , \2669 );
and \U$11917 ( \12099 , \3912 , \2538 );
nor \U$11918 ( \12100 , \12098 , \12099 );
xnor \U$11919 ( \12101 , \12100 , \2534 );
xor \U$11920 ( \12102 , \12097 , \12101 );
and \U$11921 ( \12103 , \3395 , \3103 );
and \U$11922 ( \12104 , \3646 , \2934 );
nor \U$11923 ( \12105 , \12103 , \12104 );
xnor \U$11924 ( \12106 , \12105 , \2839 );
xor \U$11925 ( \12107 , \12102 , \12106 );
xor \U$11926 ( \12108 , \12093 , \12107 );
and \U$11927 ( \12109 , \1333 , \5996 );
and \U$11928 ( \12110 , \1484 , \5695 );
nor \U$11929 ( \12111 , \12109 , \12110 );
xnor \U$11930 ( \12112 , \12111 , \5687 );
and \U$11931 ( \12113 , \1147 , \6401 );
and \U$11932 ( \12114 , \1192 , \6143 );
nor \U$11933 ( \12115 , \12113 , \12114 );
xnor \U$11934 ( \12116 , \12115 , \6148 );
xor \U$11935 ( \12117 , \12112 , \12116 );
and \U$11936 ( \12118 , \412 , \7055 );
and \U$11937 ( \12119 , \474 , \6675 );
nor \U$11938 ( \12120 , \12118 , \12119 );
xnor \U$11939 ( \12121 , \12120 , \6680 );
xor \U$11940 ( \12122 , \12117 , \12121 );
and \U$11941 ( \12123 , \2090 , \4581 );
and \U$11942 ( \12124 , \2182 , \4424 );
nor \U$11943 ( \12125 , \12123 , \12124 );
xnor \U$11944 ( \12126 , \12125 , \4377 );
and \U$11945 ( \12127 , \1802 , \5011 );
and \U$11946 ( \12128 , \1948 , \4878 );
nor \U$11947 ( \12129 , \12127 , \12128 );
xnor \U$11948 ( \12130 , \12129 , \4762 );
xor \U$11949 ( \12131 , \12126 , \12130 );
and \U$11950 ( \12132 , \1601 , \5485 );
and \U$11951 ( \12133 , \1684 , \5275 );
nor \U$11952 ( \12134 , \12132 , \12133 );
xnor \U$11953 ( \12135 , \12134 , \5169 );
xor \U$11954 ( \12136 , \12131 , \12135 );
xor \U$11955 ( \12137 , \12122 , \12136 );
and \U$11956 ( \12138 , \261 , \7489 );
and \U$11957 ( \12139 , \307 , \7137 );
nor \U$11958 ( \12140 , \12138 , \12139 );
xnor \U$11959 ( \12141 , \12140 , \7142 );
and \U$11960 ( \12142 , \178 , \8019 );
and \U$11961 ( \12143 , \185 , \7830 );
nor \U$11962 ( \12144 , \12142 , \12143 );
xnor \U$11963 ( \12145 , \12144 , \7713 );
xor \U$11964 ( \12146 , \12141 , \12145 );
and \U$11965 ( \12147 , \189 , \8540 );
and \U$11966 ( \12148 , \197 , \8292 );
nor \U$11967 ( \12149 , \12147 , \12148 );
xnor \U$11968 ( \12150 , \12149 , \8297 );
xor \U$11969 ( \12151 , \12146 , \12150 );
xor \U$11970 ( \12152 , \12137 , \12151 );
xor \U$11971 ( \12153 , \12108 , \12152 );
and \U$11972 ( \12154 , \11692 , \11696 );
and \U$11973 ( \12155 , \11696 , \11701 );
and \U$11974 ( \12156 , \11692 , \11701 );
or \U$11975 ( \12157 , \12154 , \12155 , \12156 );
and \U$11976 ( \12158 , \209 , \9333 );
and \U$11977 ( \12159 , \217 , \9006 );
nor \U$11978 ( \12160 , \12158 , \12159 );
xnor \U$11979 ( \12161 , \12160 , \8848 );
and \U$11980 ( \12162 , \224 , \9765 );
and \U$11981 ( \12163 , \232 , \9644 );
nor \U$11982 ( \12164 , \12162 , \12163 );
xnor \U$11983 ( \12165 , \12164 , \9478 );
xor \U$11984 ( \12166 , \12161 , \12165 );
and \U$11985 ( \12167 , \240 , \10408 );
and \U$11986 ( \12168 , \247 , \10116 );
nor \U$11987 ( \12169 , \12167 , \12168 );
xnor \U$11988 ( \12170 , \12169 , \10121 );
xor \U$11989 ( \12171 , \12166 , \12170 );
xor \U$11990 ( \12172 , \12157 , \12171 );
and \U$11991 ( \12173 , \143 , \10118 );
not \U$11992 ( \12174 , \12173 );
xor \U$11993 ( \12175 , \12172 , \12174 );
xor \U$11994 ( \12176 , \12153 , \12175 );
xor \U$11995 ( \12177 , \12064 , \12176 );
xor \U$11996 ( \12178 , \11999 , \12177 );
xor \U$11997 ( \12179 , \11930 , \12178 );
xor \U$11998 ( \12180 , \11916 , \12179 );
xor \U$11999 ( \12181 , \11887 , \12180 );
and \U$12000 ( \12182 , \11569 , \11829 );
and \U$12001 ( \12183 , \11829 , \11869 );
and \U$12002 ( \12184 , \11569 , \11869 );
or \U$12003 ( \12185 , \12182 , \12183 , \12184 );
xor \U$12004 ( \12186 , \12181 , \12185 );
and \U$12005 ( \12187 , \11870 , \11874 );
and \U$12006 ( \12188 , \11875 , \11878 );
or \U$12007 ( \12189 , \12187 , \12188 );
xor \U$12008 ( \12190 , \12186 , \12189 );
buf g5513_GF_PartitionCandidate( \12191_nG5513 , \12190 );
buf \U$12009 ( \12192 , \12191_nG5513 );
and \U$12010 ( \12193 , \11891 , \11915 );
and \U$12011 ( \12194 , \11915 , \12179 );
and \U$12012 ( \12195 , \11891 , \12179 );
or \U$12013 ( \12196 , \12193 , \12194 , \12195 );
and \U$12014 ( \12197 , \11895 , \11899 );
and \U$12015 ( \12198 , \11899 , \11914 );
and \U$12016 ( \12199 , \11895 , \11914 );
or \U$12017 ( \12200 , \12197 , \12198 , \12199 );
and \U$12018 ( \12201 , \11930 , \12178 );
xor \U$12019 ( \12202 , \12200 , \12201 );
and \U$12020 ( \12203 , \11957 , \11961 );
and \U$12021 ( \12204 , \11961 , \11966 );
and \U$12022 ( \12205 , \11957 , \11966 );
or \U$12023 ( \12206 , \12203 , \12204 , \12205 );
and \U$12024 ( \12207 , \11971 , \11975 );
and \U$12025 ( \12208 , \11975 , \11980 );
and \U$12026 ( \12209 , \11971 , \11980 );
or \U$12027 ( \12210 , \12207 , \12208 , \12209 );
xor \U$12028 ( \12211 , \12206 , \12210 );
and \U$12029 ( \12212 , \11986 , \11990 );
and \U$12030 ( \12213 , \11990 , \11995 );
and \U$12031 ( \12214 , \11986 , \11995 );
or \U$12032 ( \12215 , \12212 , \12213 , \12214 );
xor \U$12033 ( \12216 , \12211 , \12215 );
and \U$12034 ( \12217 , \11967 , \11981 );
and \U$12035 ( \12218 , \11981 , \11996 );
and \U$12036 ( \12219 , \11967 , \11996 );
or \U$12037 ( \12220 , \12217 , \12218 , \12219 );
and \U$12038 ( \12221 , \12108 , \12152 );
and \U$12039 ( \12222 , \12152 , \12175 );
and \U$12040 ( \12223 , \12108 , \12175 );
or \U$12041 ( \12224 , \12221 , \12222 , \12223 );
xor \U$12042 ( \12225 , \12220 , \12224 );
and \U$12043 ( \12226 , \12112 , \12116 );
and \U$12044 ( \12227 , \12116 , \12121 );
and \U$12045 ( \12228 , \12112 , \12121 );
or \U$12046 ( \12229 , \12226 , \12227 , \12228 );
and \U$12047 ( \12230 , \12126 , \12130 );
and \U$12048 ( \12231 , \12130 , \12135 );
and \U$12049 ( \12232 , \12126 , \12135 );
or \U$12050 ( \12233 , \12230 , \12231 , \12232 );
xor \U$12051 ( \12234 , \12229 , \12233 );
and \U$12052 ( \12235 , \12141 , \12145 );
and \U$12053 ( \12236 , \12145 , \12150 );
and \U$12054 ( \12237 , \12141 , \12150 );
or \U$12055 ( \12238 , \12235 , \12236 , \12237 );
xor \U$12056 ( \12239 , \12234 , \12238 );
and \U$12057 ( \12240 , \12022 , \12026 );
and \U$12058 ( \12241 , \12026 , \12031 );
and \U$12059 ( \12242 , \12022 , \12031 );
or \U$12060 ( \12243 , \12240 , \12241 , \12242 );
and \U$12061 ( \12244 , \12036 , \12040 );
and \U$12062 ( \12245 , \12040 , \12045 );
and \U$12063 ( \12246 , \12036 , \12045 );
or \U$12064 ( \12247 , \12244 , \12245 , \12246 );
xor \U$12065 ( \12248 , \12243 , \12247 );
and \U$12066 ( \12249 , \12051 , \12055 );
and \U$12067 ( \12250 , \12055 , \12060 );
and \U$12068 ( \12251 , \12051 , \12060 );
or \U$12069 ( \12252 , \12249 , \12250 , \12251 );
xor \U$12070 ( \12253 , \12248 , \12252 );
xor \U$12071 ( \12254 , \12239 , \12253 );
and \U$12072 ( \12255 , \12068 , \12072 );
and \U$12073 ( \12256 , \12072 , \12077 );
and \U$12074 ( \12257 , \12068 , \12077 );
or \U$12075 ( \12258 , \12255 , \12256 , \12257 );
and \U$12076 ( \12259 , \12082 , \12086 );
and \U$12077 ( \12260 , \12086 , \12091 );
and \U$12078 ( \12261 , \12082 , \12091 );
or \U$12079 ( \12262 , \12259 , \12260 , \12261 );
xor \U$12080 ( \12263 , \12258 , \12262 );
and \U$12081 ( \12264 , \12097 , \12101 );
and \U$12082 ( \12265 , \12101 , \12106 );
and \U$12083 ( \12266 , \12097 , \12106 );
or \U$12084 ( \12267 , \12264 , \12265 , \12266 );
xor \U$12085 ( \12268 , \12263 , \12267 );
xor \U$12086 ( \12269 , \12254 , \12268 );
xor \U$12087 ( \12270 , \12225 , \12269 );
xor \U$12088 ( \12271 , \12216 , \12270 );
and \U$12089 ( \12272 , \12078 , \12092 );
and \U$12090 ( \12273 , \12092 , \12107 );
and \U$12091 ( \12274 , \12078 , \12107 );
or \U$12092 ( \12275 , \12272 , \12273 , \12274 );
and \U$12093 ( \12276 , \12122 , \12136 );
and \U$12094 ( \12277 , \12136 , \12151 );
and \U$12095 ( \12278 , \12122 , \12151 );
or \U$12096 ( \12279 , \12276 , \12277 , \12278 );
xor \U$12097 ( \12280 , \12275 , \12279 );
and \U$12098 ( \12281 , \12157 , \12171 );
and \U$12099 ( \12282 , \12171 , \12174 );
and \U$12100 ( \12283 , \12157 , \12174 );
or \U$12101 ( \12284 , \12281 , \12282 , \12283 );
xor \U$12102 ( \12285 , \12280 , \12284 );
and \U$12103 ( \12286 , \12161 , \12165 );
and \U$12104 ( \12287 , \12165 , \12170 );
and \U$12105 ( \12288 , \12161 , \12170 );
or \U$12106 ( \12289 , \12286 , \12287 , \12288 );
buf \U$12107 ( \12290 , \12173 );
xor \U$12108 ( \12291 , \12289 , \12290 );
and \U$12109 ( \12292 , \240 , \10118 );
xor \U$12110 ( \12293 , \12291 , \12292 );
and \U$12111 ( \12294 , \217 , \9333 );
and \U$12112 ( \12295 , \189 , \9006 );
nor \U$12113 ( \12296 , \12294 , \12295 );
xnor \U$12114 ( \12297 , \12296 , \8848 );
and \U$12115 ( \12298 , \232 , \9765 );
and \U$12116 ( \12299 , \209 , \9644 );
nor \U$12117 ( \12300 , \12298 , \12299 );
xnor \U$12118 ( \12301 , \12300 , \9478 );
xor \U$12119 ( \12302 , \12297 , \12301 );
and \U$12120 ( \12303 , \247 , \10408 );
and \U$12121 ( \12304 , \224 , \10116 );
nor \U$12122 ( \12305 , \12303 , \12304 );
xnor \U$12123 ( \12306 , \12305 , \10121 );
xor \U$12124 ( \12307 , \12302 , \12306 );
and \U$12125 ( \12308 , \307 , \7489 );
and \U$12126 ( \12309 , \412 , \7137 );
nor \U$12127 ( \12310 , \12308 , \12309 );
xnor \U$12128 ( \12311 , \12310 , \7142 );
and \U$12129 ( \12312 , \185 , \8019 );
and \U$12130 ( \12313 , \261 , \7830 );
nor \U$12131 ( \12314 , \12312 , \12313 );
xnor \U$12132 ( \12315 , \12314 , \7713 );
xor \U$12133 ( \12316 , \12311 , \12315 );
and \U$12134 ( \12317 , \197 , \8540 );
and \U$12135 ( \12318 , \178 , \8292 );
nor \U$12136 ( \12319 , \12317 , \12318 );
xnor \U$12137 ( \12320 , \12319 , \8297 );
xor \U$12138 ( \12321 , \12316 , \12320 );
xor \U$12139 ( \12322 , \12307 , \12321 );
and \U$12140 ( \12323 , \1484 , \5996 );
and \U$12141 ( \12324 , \1601 , \5695 );
nor \U$12142 ( \12325 , \12323 , \12324 );
xnor \U$12143 ( \12326 , \12325 , \5687 );
and \U$12144 ( \12327 , \1192 , \6401 );
and \U$12145 ( \12328 , \1333 , \6143 );
nor \U$12146 ( \12329 , \12327 , \12328 );
xnor \U$12147 ( \12330 , \12329 , \6148 );
xor \U$12148 ( \12331 , \12326 , \12330 );
and \U$12149 ( \12332 , \474 , \7055 );
and \U$12150 ( \12333 , \1147 , \6675 );
nor \U$12151 ( \12334 , \12332 , \12333 );
xnor \U$12152 ( \12335 , \12334 , \6680 );
xor \U$12153 ( \12336 , \12331 , \12335 );
xor \U$12154 ( \12337 , \12322 , \12336 );
xor \U$12155 ( \12338 , \12293 , \12337 );
and \U$12156 ( \12339 , \2182 , \4581 );
and \U$12157 ( \12340 , \2366 , \4424 );
nor \U$12158 ( \12341 , \12339 , \12340 );
xnor \U$12159 ( \12342 , \12341 , \4377 );
and \U$12160 ( \12343 , \1948 , \5011 );
and \U$12161 ( \12344 , \2090 , \4878 );
nor \U$12162 ( \12345 , \12343 , \12344 );
xnor \U$12163 ( \12346 , \12345 , \4762 );
xor \U$12164 ( \12347 , \12342 , \12346 );
and \U$12165 ( \12348 , \1684 , \5485 );
and \U$12166 ( \12349 , \1802 , \5275 );
nor \U$12167 ( \12350 , \12348 , \12349 );
xnor \U$12168 ( \12351 , \12350 , \5169 );
xor \U$12169 ( \12352 , \12347 , \12351 );
and \U$12170 ( \12353 , \4364 , \2400 );
and \U$12171 ( \12354 , \4654 , \2246 );
nor \U$12172 ( \12355 , \12353 , \12354 );
xnor \U$12173 ( \12356 , \12355 , \2195 );
and \U$12174 ( \12357 , \3912 , \2669 );
and \U$12175 ( \12358 , \4160 , \2538 );
nor \U$12176 ( \12359 , \12357 , \12358 );
xnor \U$12177 ( \12360 , \12359 , \2534 );
xor \U$12178 ( \12361 , \12356 , \12360 );
and \U$12179 ( \12362 , \3646 , \3103 );
and \U$12180 ( \12363 , \3736 , \2934 );
nor \U$12181 ( \12364 , \12362 , \12363 );
xnor \U$12182 ( \12365 , \12364 , \2839 );
xor \U$12183 ( \12366 , \12361 , \12365 );
xor \U$12184 ( \12367 , \12352 , \12366 );
and \U$12185 ( \12368 , \3143 , \3357 );
and \U$12186 ( \12369 , \3395 , \3255 );
nor \U$12187 ( \12370 , \12368 , \12369 );
xnor \U$12188 ( \12371 , \12370 , \3156 );
and \U$12189 ( \12372 , \2826 , \3813 );
and \U$12190 ( \12373 , \3037 , \3557 );
nor \U$12191 ( \12374 , \12372 , \12373 );
xnor \U$12192 ( \12375 , \12374 , \3562 );
xor \U$12193 ( \12376 , \12371 , \12375 );
and \U$12194 ( \12377 , \2521 , \4132 );
and \U$12195 ( \12378 , \2757 , \4012 );
nor \U$12196 ( \12379 , \12377 , \12378 );
xnor \U$12197 ( \12380 , \12379 , \3925 );
xor \U$12198 ( \12381 , \12376 , \12380 );
xor \U$12199 ( \12382 , \12367 , \12381 );
xor \U$12200 ( \12383 , \12338 , \12382 );
xor \U$12201 ( \12384 , \12285 , \12383 );
and \U$12202 ( \12385 , \12032 , \12046 );
and \U$12203 ( \12386 , \12046 , \12061 );
and \U$12204 ( \12387 , \12032 , \12061 );
or \U$12205 ( \12388 , \12385 , \12386 , \12387 );
not \U$12206 ( \12389 , \222 );
and \U$12207 ( \12390 , \10206 , \230 );
and \U$12208 ( \12391 , \10584 , \228 );
nor \U$12209 ( \12392 , \12390 , \12391 );
xnor \U$12210 ( \12393 , \12392 , \237 );
xor \U$12211 ( \12394 , \12389 , \12393 );
and \U$12212 ( \12395 , \9465 , \245 );
and \U$12213 ( \12396 , \9897 , \243 );
nor \U$12214 ( \12397 , \12395 , \12396 );
xnor \U$12215 ( \12398 , \12397 , \252 );
xor \U$12216 ( \12399 , \12394 , \12398 );
xor \U$12217 ( \12400 , \12388 , \12399 );
and \U$12218 ( \12401 , \7231 , \438 );
and \U$12219 ( \12402 , \7556 , \336 );
nor \U$12220 ( \12403 , \12401 , \12402 );
xnor \U$12221 ( \12404 , \12403 , \320 );
and \U$12222 ( \12405 , \6790 , \1086 );
and \U$12223 ( \12406 , \6945 , \508 );
nor \U$12224 ( \12407 , \12405 , \12406 );
xnor \U$12225 ( \12408 , \12407 , \487 );
xor \U$12226 ( \12409 , \12404 , \12408 );
and \U$12227 ( \12410 , \6281 , \1301 );
and \U$12228 ( \12411 , \6514 , \1246 );
nor \U$12229 ( \12412 , \12410 , \12411 );
xnor \U$12230 ( \12413 , \12412 , \1205 );
xor \U$12231 ( \12414 , \12409 , \12413 );
and \U$12232 ( \12415 , \8835 , \141 );
and \U$12233 ( \12416 , \9169 , \139 );
nor \U$12234 ( \12417 , \12415 , \12416 );
xnor \U$12235 ( \12418 , \12417 , \148 );
and \U$12236 ( \12419 , \8349 , \156 );
and \U$12237 ( \12420 , \8652 , \154 );
nor \U$12238 ( \12421 , \12419 , \12420 );
xnor \U$12239 ( \12422 , \12421 , \163 );
xor \U$12240 ( \12423 , \12418 , \12422 );
and \U$12241 ( \12424 , \7700 , \296 );
and \U$12242 ( \12425 , \8057 , \168 );
nor \U$12243 ( \12426 , \12424 , \12425 );
xnor \U$12244 ( \12427 , \12426 , \173 );
xor \U$12245 ( \12428 , \12423 , \12427 );
xor \U$12246 ( \12429 , \12414 , \12428 );
and \U$12247 ( \12430 , \5674 , \1578 );
and \U$12248 ( \12431 , \6030 , \1431 );
nor \U$12249 ( \12432 , \12430 , \12431 );
xnor \U$12250 ( \12433 , \12432 , \1436 );
and \U$12251 ( \12434 , \5156 , \1824 );
and \U$12252 ( \12435 , \5469 , \1739 );
nor \U$12253 ( \12436 , \12434 , \12435 );
xnor \U$12254 ( \12437 , \12436 , \1697 );
xor \U$12255 ( \12438 , \12433 , \12437 );
and \U$12256 ( \12439 , \4749 , \2121 );
and \U$12257 ( \12440 , \4922 , \2008 );
nor \U$12258 ( \12441 , \12439 , \12440 );
xnor \U$12259 ( \12442 , \12441 , \1961 );
xor \U$12260 ( \12443 , \12438 , \12442 );
xor \U$12261 ( \12444 , \12429 , \12443 );
xor \U$12262 ( \12445 , \12400 , \12444 );
xor \U$12263 ( \12446 , \12384 , \12445 );
xor \U$12264 ( \12447 , \12271 , \12446 );
xor \U$12265 ( \12448 , \12202 , \12447 );
xor \U$12266 ( \12449 , \12196 , \12448 );
and \U$12267 ( \12450 , \11904 , \11908 );
and \U$12268 ( \12451 , \11908 , \11913 );
and \U$12269 ( \12452 , \11904 , \11913 );
or \U$12270 ( \12453 , \12450 , \12451 , \12452 );
and \U$12271 ( \12454 , \11948 , \11952 );
and \U$12272 ( \12455 , \11952 , \11997 );
and \U$12273 ( \12456 , \11948 , \11997 );
or \U$12274 ( \12457 , \12454 , \12455 , \12456 );
xor \U$12275 ( \12458 , \12453 , \12457 );
and \U$12276 ( \12459 , \12013 , \12063 );
and \U$12277 ( \12460 , \12063 , \12176 );
and \U$12278 ( \12461 , \12013 , \12176 );
or \U$12279 ( \12462 , \12459 , \12460 , \12461 );
xor \U$12280 ( \12463 , \12458 , \12462 );
and \U$12281 ( \12464 , \11920 , \11924 );
and \U$12282 ( \12465 , \11924 , \11929 );
and \U$12283 ( \12466 , \11920 , \11929 );
or \U$12284 ( \12467 , \12464 , \12465 , \12466 );
and \U$12285 ( \12468 , \11944 , \11998 );
and \U$12286 ( \12469 , \11998 , \12177 );
and \U$12287 ( \12470 , \11944 , \12177 );
or \U$12288 ( \12471 , \12468 , \12469 , \12470 );
xor \U$12289 ( \12472 , \12467 , \12471 );
and \U$12290 ( \12473 , \11934 , \11938 );
and \U$12291 ( \12474 , \11938 , \11943 );
and \U$12292 ( \12475 , \11934 , \11943 );
or \U$12293 ( \12476 , \12473 , \12474 , \12475 );
and \U$12294 ( \12477 , \12003 , \12007 );
and \U$12295 ( \12478 , \12007 , \12012 );
and \U$12296 ( \12479 , \12003 , \12012 );
or \U$12297 ( \12480 , \12477 , \12478 , \12479 );
xor \U$12298 ( \12481 , \12476 , \12480 );
and \U$12299 ( \12482 , \12017 , \12018 );
and \U$12300 ( \12483 , \12018 , \12062 );
and \U$12301 ( \12484 , \12017 , \12062 );
or \U$12302 ( \12485 , \12482 , \12483 , \12484 );
xor \U$12303 ( \12486 , \12481 , \12485 );
xor \U$12304 ( \12487 , \12472 , \12486 );
xor \U$12305 ( \12488 , \12463 , \12487 );
xor \U$12306 ( \12489 , \12449 , \12488 );
and \U$12307 ( \12490 , \11885 , \11886 );
and \U$12308 ( \12491 , \11886 , \12180 );
and \U$12309 ( \12492 , \11885 , \12180 );
or \U$12310 ( \12493 , \12490 , \12491 , \12492 );
xor \U$12311 ( \12494 , \12489 , \12493 );
and \U$12312 ( \12495 , \12181 , \12185 );
and \U$12313 ( \12496 , \12186 , \12189 );
or \U$12314 ( \12497 , \12495 , \12496 );
xor \U$12315 ( \12498 , \12494 , \12497 );
buf g5511_GF_PartitionCandidate( \12499_nG5511 , \12498 );
buf \U$12316 ( \12500 , \12499_nG5511 );
and \U$12317 ( \12501 , \12200 , \12201 );
and \U$12318 ( \12502 , \12201 , \12447 );
and \U$12319 ( \12503 , \12200 , \12447 );
or \U$12320 ( \12504 , \12501 , \12502 , \12503 );
and \U$12321 ( \12505 , \12463 , \12487 );
xor \U$12322 ( \12506 , \12504 , \12505 );
and \U$12323 ( \12507 , \12467 , \12471 );
and \U$12324 ( \12508 , \12471 , \12486 );
and \U$12325 ( \12509 , \12467 , \12486 );
or \U$12326 ( \12510 , \12507 , \12508 , \12509 );
and \U$12327 ( \12511 , \12453 , \12457 );
and \U$12328 ( \12512 , \12457 , \12462 );
and \U$12329 ( \12513 , \12453 , \12462 );
or \U$12330 ( \12514 , \12511 , \12512 , \12513 );
and \U$12331 ( \12515 , \12216 , \12270 );
and \U$12332 ( \12516 , \12270 , \12446 );
and \U$12333 ( \12517 , \12216 , \12446 );
or \U$12334 ( \12518 , \12515 , \12516 , \12517 );
xor \U$12335 ( \12519 , \12514 , \12518 );
and \U$12336 ( \12520 , \12239 , \12253 );
and \U$12337 ( \12521 , \12253 , \12268 );
and \U$12338 ( \12522 , \12239 , \12268 );
or \U$12339 ( \12523 , \12520 , \12521 , \12522 );
and \U$12340 ( \12524 , \12293 , \12337 );
and \U$12341 ( \12525 , \12337 , \12382 );
and \U$12342 ( \12526 , \12293 , \12382 );
or \U$12343 ( \12527 , \12524 , \12525 , \12526 );
xor \U$12344 ( \12528 , \12523 , \12527 );
and \U$12345 ( \12529 , \12356 , \12360 );
and \U$12346 ( \12530 , \12360 , \12365 );
and \U$12347 ( \12531 , \12356 , \12365 );
or \U$12348 ( \12532 , \12529 , \12530 , \12531 );
and \U$12349 ( \12533 , \12371 , \12375 );
and \U$12350 ( \12534 , \12375 , \12380 );
and \U$12351 ( \12535 , \12371 , \12380 );
or \U$12352 ( \12536 , \12533 , \12534 , \12535 );
xor \U$12353 ( \12537 , \12532 , \12536 );
and \U$12354 ( \12538 , \12433 , \12437 );
and \U$12355 ( \12539 , \12437 , \12442 );
and \U$12356 ( \12540 , \12433 , \12442 );
or \U$12357 ( \12541 , \12538 , \12539 , \12540 );
xor \U$12358 ( \12542 , \12537 , \12541 );
xor \U$12359 ( \12543 , \12528 , \12542 );
xor \U$12360 ( \12544 , \12519 , \12543 );
xor \U$12361 ( \12545 , \12510 , \12544 );
and \U$12362 ( \12546 , \12206 , \12210 );
and \U$12363 ( \12547 , \12210 , \12215 );
and \U$12364 ( \12548 , \12206 , \12215 );
or \U$12365 ( \12549 , \12546 , \12547 , \12548 );
and \U$12366 ( \12550 , \12275 , \12279 );
and \U$12367 ( \12551 , \12279 , \12284 );
and \U$12368 ( \12552 , \12275 , \12284 );
or \U$12369 ( \12553 , \12550 , \12551 , \12552 );
xor \U$12370 ( \12554 , \12549 , \12553 );
and \U$12371 ( \12555 , \12388 , \12399 );
and \U$12372 ( \12556 , \12399 , \12444 );
and \U$12373 ( \12557 , \12388 , \12444 );
or \U$12374 ( \12558 , \12555 , \12556 , \12557 );
xor \U$12375 ( \12559 , \12554 , \12558 );
and \U$12376 ( \12560 , \12476 , \12480 );
and \U$12377 ( \12561 , \12480 , \12485 );
and \U$12378 ( \12562 , \12476 , \12485 );
or \U$12379 ( \12563 , \12560 , \12561 , \12562 );
and \U$12380 ( \12564 , \12220 , \12224 );
and \U$12381 ( \12565 , \12224 , \12269 );
and \U$12382 ( \12566 , \12220 , \12269 );
or \U$12383 ( \12567 , \12564 , \12565 , \12566 );
xor \U$12384 ( \12568 , \12563 , \12567 );
and \U$12385 ( \12569 , \12285 , \12383 );
and \U$12386 ( \12570 , \12383 , \12445 );
and \U$12387 ( \12571 , \12285 , \12445 );
or \U$12388 ( \12572 , \12569 , \12570 , \12571 );
xor \U$12389 ( \12573 , \12568 , \12572 );
xor \U$12390 ( \12574 , \12559 , \12573 );
and \U$12391 ( \12575 , \12229 , \12233 );
and \U$12392 ( \12576 , \12233 , \12238 );
and \U$12393 ( \12577 , \12229 , \12238 );
or \U$12394 ( \12578 , \12575 , \12576 , \12577 );
and \U$12395 ( \12579 , \12243 , \12247 );
and \U$12396 ( \12580 , \12247 , \12252 );
and \U$12397 ( \12581 , \12243 , \12252 );
or \U$12398 ( \12582 , \12579 , \12580 , \12581 );
xor \U$12399 ( \12583 , \12578 , \12582 );
and \U$12400 ( \12584 , \12258 , \12262 );
and \U$12401 ( \12585 , \12262 , \12267 );
and \U$12402 ( \12586 , \12258 , \12267 );
or \U$12403 ( \12587 , \12584 , \12585 , \12586 );
xor \U$12404 ( \12588 , \12583 , \12587 );
and \U$12405 ( \12589 , \12289 , \12290 );
and \U$12406 ( \12590 , \12290 , \12292 );
and \U$12407 ( \12591 , \12289 , \12292 );
or \U$12408 ( \12592 , \12589 , \12590 , \12591 );
and \U$12409 ( \12593 , \12307 , \12321 );
and \U$12410 ( \12594 , \12321 , \12336 );
and \U$12411 ( \12595 , \12307 , \12336 );
or \U$12412 ( \12596 , \12593 , \12594 , \12595 );
xor \U$12413 ( \12597 , \12592 , \12596 );
and \U$12414 ( \12598 , \12352 , \12366 );
and \U$12415 ( \12599 , \12366 , \12381 );
and \U$12416 ( \12600 , \12352 , \12381 );
or \U$12417 ( \12601 , \12598 , \12599 , \12600 );
xor \U$12418 ( \12602 , \12597 , \12601 );
xor \U$12419 ( \12603 , \12588 , \12602 );
and \U$12420 ( \12604 , \12389 , \12393 );
and \U$12421 ( \12605 , \12393 , \12398 );
and \U$12422 ( \12606 , \12389 , \12398 );
or \U$12423 ( \12607 , \12604 , \12605 , \12606 );
and \U$12424 ( \12608 , \12404 , \12408 );
and \U$12425 ( \12609 , \12408 , \12413 );
and \U$12426 ( \12610 , \12404 , \12413 );
or \U$12427 ( \12611 , \12608 , \12609 , \12610 );
xor \U$12428 ( \12612 , \12607 , \12611 );
and \U$12429 ( \12613 , \12418 , \12422 );
and \U$12430 ( \12614 , \12422 , \12427 );
and \U$12431 ( \12615 , \12418 , \12427 );
or \U$12432 ( \12616 , \12613 , \12614 , \12615 );
xor \U$12433 ( \12617 , \12612 , \12616 );
and \U$12434 ( \12618 , \12414 , \12428 );
and \U$12435 ( \12619 , \12428 , \12443 );
and \U$12436 ( \12620 , \12414 , \12443 );
or \U$12437 ( \12621 , \12618 , \12619 , \12620 );
and \U$12438 ( \12622 , \10584 , \230 );
not \U$12439 ( \12623 , \12622 );
xnor \U$12440 ( \12624 , \12623 , \237 );
and \U$12441 ( \12625 , \9897 , \245 );
and \U$12442 ( \12626 , \10206 , \243 );
nor \U$12443 ( \12627 , \12625 , \12626 );
xnor \U$12444 ( \12628 , \12627 , \252 );
xor \U$12445 ( \12629 , \12624 , \12628 );
and \U$12446 ( \12630 , \9169 , \141 );
and \U$12447 ( \12631 , \9465 , \139 );
nor \U$12448 ( \12632 , \12630 , \12631 );
xnor \U$12449 ( \12633 , \12632 , \148 );
xor \U$12450 ( \12634 , \12629 , \12633 );
and \U$12451 ( \12635 , \6945 , \1086 );
and \U$12452 ( \12636 , \7231 , \508 );
nor \U$12453 ( \12637 , \12635 , \12636 );
xnor \U$12454 ( \12638 , \12637 , \487 );
and \U$12455 ( \12639 , \6514 , \1301 );
and \U$12456 ( \12640 , \6790 , \1246 );
nor \U$12457 ( \12641 , \12639 , \12640 );
xnor \U$12458 ( \12642 , \12641 , \1205 );
xor \U$12459 ( \12643 , \12638 , \12642 );
and \U$12460 ( \12644 , \6030 , \1578 );
and \U$12461 ( \12645 , \6281 , \1431 );
nor \U$12462 ( \12646 , \12644 , \12645 );
xnor \U$12463 ( \12647 , \12646 , \1436 );
xor \U$12464 ( \12648 , \12643 , \12647 );
xor \U$12465 ( \12649 , \12634 , \12648 );
and \U$12466 ( \12650 , \8652 , \156 );
and \U$12467 ( \12651 , \8835 , \154 );
nor \U$12468 ( \12652 , \12650 , \12651 );
xnor \U$12469 ( \12653 , \12652 , \163 );
and \U$12470 ( \12654 , \8057 , \296 );
and \U$12471 ( \12655 , \8349 , \168 );
nor \U$12472 ( \12656 , \12654 , \12655 );
xnor \U$12473 ( \12657 , \12656 , \173 );
xor \U$12474 ( \12658 , \12653 , \12657 );
and \U$12475 ( \12659 , \7556 , \438 );
and \U$12476 ( \12660 , \7700 , \336 );
nor \U$12477 ( \12661 , \12659 , \12660 );
xnor \U$12478 ( \12662 , \12661 , \320 );
xor \U$12479 ( \12663 , \12658 , \12662 );
xor \U$12480 ( \12664 , \12649 , \12663 );
xor \U$12481 ( \12665 , \12621 , \12664 );
and \U$12482 ( \12666 , \3037 , \3813 );
and \U$12483 ( \12667 , \3143 , \3557 );
nor \U$12484 ( \12668 , \12666 , \12667 );
xnor \U$12485 ( \12669 , \12668 , \3562 );
and \U$12486 ( \12670 , \2757 , \4132 );
and \U$12487 ( \12671 , \2826 , \4012 );
nor \U$12488 ( \12672 , \12670 , \12671 );
xnor \U$12489 ( \12673 , \12672 , \3925 );
xor \U$12490 ( \12674 , \12669 , \12673 );
and \U$12491 ( \12675 , \2366 , \4581 );
and \U$12492 ( \12676 , \2521 , \4424 );
nor \U$12493 ( \12677 , \12675 , \12676 );
xnor \U$12494 ( \12678 , \12677 , \4377 );
xor \U$12495 ( \12679 , \12674 , \12678 );
and \U$12496 ( \12680 , \5469 , \1824 );
and \U$12497 ( \12681 , \5674 , \1739 );
nor \U$12498 ( \12682 , \12680 , \12681 );
xnor \U$12499 ( \12683 , \12682 , \1697 );
and \U$12500 ( \12684 , \4922 , \2121 );
and \U$12501 ( \12685 , \5156 , \2008 );
nor \U$12502 ( \12686 , \12684 , \12685 );
xnor \U$12503 ( \12687 , \12686 , \1961 );
xor \U$12504 ( \12688 , \12683 , \12687 );
and \U$12505 ( \12689 , \4654 , \2400 );
and \U$12506 ( \12690 , \4749 , \2246 );
nor \U$12507 ( \12691 , \12689 , \12690 );
xnor \U$12508 ( \12692 , \12691 , \2195 );
xor \U$12509 ( \12693 , \12688 , \12692 );
xor \U$12510 ( \12694 , \12679 , \12693 );
and \U$12511 ( \12695 , \4160 , \2669 );
and \U$12512 ( \12696 , \4364 , \2538 );
nor \U$12513 ( \12697 , \12695 , \12696 );
xnor \U$12514 ( \12698 , \12697 , \2534 );
and \U$12515 ( \12699 , \3736 , \3103 );
and \U$12516 ( \12700 , \3912 , \2934 );
nor \U$12517 ( \12701 , \12699 , \12700 );
xnor \U$12518 ( \12702 , \12701 , \2839 );
xor \U$12519 ( \12703 , \12698 , \12702 );
and \U$12520 ( \12704 , \3395 , \3357 );
and \U$12521 ( \12705 , \3646 , \3255 );
nor \U$12522 ( \12706 , \12704 , \12705 );
xnor \U$12523 ( \12707 , \12706 , \3156 );
xor \U$12524 ( \12708 , \12703 , \12707 );
xor \U$12525 ( \12709 , \12694 , \12708 );
xor \U$12526 ( \12710 , \12665 , \12709 );
xor \U$12527 ( \12711 , \12617 , \12710 );
and \U$12528 ( \12712 , \12311 , \12315 );
and \U$12529 ( \12713 , \12315 , \12320 );
and \U$12530 ( \12714 , \12311 , \12320 );
or \U$12531 ( \12715 , \12712 , \12713 , \12714 );
and \U$12532 ( \12716 , \12326 , \12330 );
and \U$12533 ( \12717 , \12330 , \12335 );
and \U$12534 ( \12718 , \12326 , \12335 );
or \U$12535 ( \12719 , \12716 , \12717 , \12718 );
xor \U$12536 ( \12720 , \12715 , \12719 );
and \U$12537 ( \12721 , \12342 , \12346 );
and \U$12538 ( \12722 , \12346 , \12351 );
and \U$12539 ( \12723 , \12342 , \12351 );
or \U$12540 ( \12724 , \12721 , \12722 , \12723 );
xor \U$12541 ( \12725 , \12720 , \12724 );
and \U$12542 ( \12726 , \261 , \8019 );
and \U$12543 ( \12727 , \307 , \7830 );
nor \U$12544 ( \12728 , \12726 , \12727 );
xnor \U$12545 ( \12729 , \12728 , \7713 );
and \U$12546 ( \12730 , \178 , \8540 );
and \U$12547 ( \12731 , \185 , \8292 );
nor \U$12548 ( \12732 , \12730 , \12731 );
xnor \U$12549 ( \12733 , \12732 , \8297 );
xor \U$12550 ( \12734 , \12729 , \12733 );
and \U$12551 ( \12735 , \189 , \9333 );
and \U$12552 ( \12736 , \197 , \9006 );
nor \U$12553 ( \12737 , \12735 , \12736 );
xnor \U$12554 ( \12738 , \12737 , \8848 );
xor \U$12555 ( \12739 , \12734 , \12738 );
and \U$12556 ( \12740 , \1333 , \6401 );
and \U$12557 ( \12741 , \1484 , \6143 );
nor \U$12558 ( \12742 , \12740 , \12741 );
xnor \U$12559 ( \12743 , \12742 , \6148 );
and \U$12560 ( \12744 , \1147 , \7055 );
and \U$12561 ( \12745 , \1192 , \6675 );
nor \U$12562 ( \12746 , \12744 , \12745 );
xnor \U$12563 ( \12747 , \12746 , \6680 );
xor \U$12564 ( \12748 , \12743 , \12747 );
and \U$12565 ( \12749 , \412 , \7489 );
and \U$12566 ( \12750 , \474 , \7137 );
nor \U$12567 ( \12751 , \12749 , \12750 );
xnor \U$12568 ( \12752 , \12751 , \7142 );
xor \U$12569 ( \12753 , \12748 , \12752 );
xor \U$12570 ( \12754 , \12739 , \12753 );
and \U$12571 ( \12755 , \2090 , \5011 );
and \U$12572 ( \12756 , \2182 , \4878 );
nor \U$12573 ( \12757 , \12755 , \12756 );
xnor \U$12574 ( \12758 , \12757 , \4762 );
and \U$12575 ( \12759 , \1802 , \5485 );
and \U$12576 ( \12760 , \1948 , \5275 );
nor \U$12577 ( \12761 , \12759 , \12760 );
xnor \U$12578 ( \12762 , \12761 , \5169 );
xor \U$12579 ( \12763 , \12758 , \12762 );
and \U$12580 ( \12764 , \1601 , \5996 );
and \U$12581 ( \12765 , \1684 , \5695 );
nor \U$12582 ( \12766 , \12764 , \12765 );
xnor \U$12583 ( \12767 , \12766 , \5687 );
xor \U$12584 ( \12768 , \12763 , \12767 );
xor \U$12585 ( \12769 , \12754 , \12768 );
xor \U$12586 ( \12770 , \12725 , \12769 );
and \U$12587 ( \12771 , \12297 , \12301 );
and \U$12588 ( \12772 , \12301 , \12306 );
and \U$12589 ( \12773 , \12297 , \12306 );
or \U$12590 ( \12774 , \12771 , \12772 , \12773 );
and \U$12591 ( \12775 , \209 , \9765 );
and \U$12592 ( \12776 , \217 , \9644 );
nor \U$12593 ( \12777 , \12775 , \12776 );
xnor \U$12594 ( \12778 , \12777 , \9478 );
and \U$12595 ( \12779 , \224 , \10408 );
and \U$12596 ( \12780 , \232 , \10116 );
nor \U$12597 ( \12781 , \12779 , \12780 );
xnor \U$12598 ( \12782 , \12781 , \10121 );
xor \U$12599 ( \12783 , \12778 , \12782 );
and \U$12600 ( \12784 , \247 , \10118 );
xor \U$12601 ( \12785 , \12783 , \12784 );
xnor \U$12602 ( \12786 , \12774 , \12785 );
xor \U$12603 ( \12787 , \12770 , \12786 );
xor \U$12604 ( \12788 , \12711 , \12787 );
xor \U$12605 ( \12789 , \12603 , \12788 );
xor \U$12606 ( \12790 , \12574 , \12789 );
xor \U$12607 ( \12791 , \12545 , \12790 );
xor \U$12608 ( \12792 , \12506 , \12791 );
and \U$12609 ( \12793 , \12196 , \12448 );
and \U$12610 ( \12794 , \12448 , \12488 );
and \U$12611 ( \12795 , \12196 , \12488 );
or \U$12612 ( \12796 , \12793 , \12794 , \12795 );
xor \U$12613 ( \12797 , \12792 , \12796 );
and \U$12614 ( \12798 , \12489 , \12493 );
and \U$12615 ( \12799 , \12494 , \12497 );
or \U$12616 ( \12800 , \12798 , \12799 );
xor \U$12617 ( \12801 , \12797 , \12800 );
buf g550f_GF_PartitionCandidate( \12802_nG550f , \12801 );
buf \U$12618 ( \12803 , \12802_nG550f );
and \U$12619 ( \12804 , \12510 , \12544 );
and \U$12620 ( \12805 , \12544 , \12790 );
and \U$12621 ( \12806 , \12510 , \12790 );
or \U$12622 ( \12807 , \12804 , \12805 , \12806 );
and \U$12623 ( \12808 , \12514 , \12518 );
and \U$12624 ( \12809 , \12518 , \12543 );
and \U$12625 ( \12810 , \12514 , \12543 );
or \U$12626 ( \12811 , \12808 , \12809 , \12810 );
and \U$12627 ( \12812 , \12559 , \12573 );
and \U$12628 ( \12813 , \12573 , \12789 );
and \U$12629 ( \12814 , \12559 , \12789 );
or \U$12630 ( \12815 , \12812 , \12813 , \12814 );
xor \U$12631 ( \12816 , \12811 , \12815 );
and \U$12632 ( \12817 , \12549 , \12553 );
and \U$12633 ( \12818 , \12553 , \12558 );
and \U$12634 ( \12819 , \12549 , \12558 );
or \U$12635 ( \12820 , \12817 , \12818 , \12819 );
and \U$12636 ( \12821 , \12523 , \12527 );
and \U$12637 ( \12822 , \12527 , \12542 );
and \U$12638 ( \12823 , \12523 , \12542 );
or \U$12639 ( \12824 , \12821 , \12822 , \12823 );
xor \U$12640 ( \12825 , \12820 , \12824 );
and \U$12641 ( \12826 , \12617 , \12710 );
and \U$12642 ( \12827 , \12710 , \12787 );
and \U$12643 ( \12828 , \12617 , \12787 );
or \U$12644 ( \12829 , \12826 , \12827 , \12828 );
xor \U$12645 ( \12830 , \12825 , \12829 );
xor \U$12646 ( \12831 , \12816 , \12830 );
xor \U$12647 ( \12832 , \12807 , \12831 );
and \U$12648 ( \12833 , \12563 , \12567 );
and \U$12649 ( \12834 , \12567 , \12572 );
and \U$12650 ( \12835 , \12563 , \12572 );
or \U$12651 ( \12836 , \12833 , \12834 , \12835 );
and \U$12652 ( \12837 , \12588 , \12602 );
and \U$12653 ( \12838 , \12602 , \12788 );
and \U$12654 ( \12839 , \12588 , \12788 );
or \U$12655 ( \12840 , \12837 , \12838 , \12839 );
xor \U$12656 ( \12841 , \12836 , \12840 );
and \U$12657 ( \12842 , \12578 , \12582 );
and \U$12658 ( \12843 , \12582 , \12587 );
and \U$12659 ( \12844 , \12578 , \12587 );
or \U$12660 ( \12845 , \12842 , \12843 , \12844 );
and \U$12661 ( \12846 , \12592 , \12596 );
and \U$12662 ( \12847 , \12596 , \12601 );
and \U$12663 ( \12848 , \12592 , \12601 );
or \U$12664 ( \12849 , \12846 , \12847 , \12848 );
xor \U$12665 ( \12850 , \12845 , \12849 );
and \U$12666 ( \12851 , \12621 , \12664 );
and \U$12667 ( \12852 , \12664 , \12709 );
and \U$12668 ( \12853 , \12621 , \12709 );
or \U$12669 ( \12854 , \12851 , \12852 , \12853 );
xor \U$12670 ( \12855 , \12850 , \12854 );
and \U$12671 ( \12856 , \12739 , \12753 );
and \U$12672 ( \12857 , \12753 , \12768 );
and \U$12673 ( \12858 , \12739 , \12768 );
or \U$12674 ( \12859 , \12856 , \12857 , \12858 );
and \U$12675 ( \12860 , \12679 , \12693 );
and \U$12676 ( \12861 , \12693 , \12708 );
and \U$12677 ( \12862 , \12679 , \12708 );
or \U$12678 ( \12863 , \12860 , \12861 , \12862 );
xor \U$12679 ( \12864 , \12859 , \12863 );
or \U$12680 ( \12865 , \12774 , \12785 );
xor \U$12681 ( \12866 , \12864 , \12865 );
and \U$12682 ( \12867 , \12607 , \12611 );
and \U$12683 ( \12868 , \12611 , \12616 );
and \U$12684 ( \12869 , \12607 , \12616 );
or \U$12685 ( \12870 , \12867 , \12868 , \12869 );
and \U$12686 ( \12871 , \12532 , \12536 );
and \U$12687 ( \12872 , \12536 , \12541 );
and \U$12688 ( \12873 , \12532 , \12541 );
or \U$12689 ( \12874 , \12871 , \12872 , \12873 );
xor \U$12690 ( \12875 , \12870 , \12874 );
and \U$12691 ( \12876 , \12715 , \12719 );
and \U$12692 ( \12877 , \12719 , \12724 );
and \U$12693 ( \12878 , \12715 , \12724 );
or \U$12694 ( \12879 , \12876 , \12877 , \12878 );
xor \U$12695 ( \12880 , \12875 , \12879 );
xor \U$12696 ( \12881 , \12866 , \12880 );
and \U$12697 ( \12882 , \12634 , \12648 );
and \U$12698 ( \12883 , \12648 , \12663 );
and \U$12699 ( \12884 , \12634 , \12663 );
or \U$12700 ( \12885 , \12882 , \12883 , \12884 );
and \U$12701 ( \12886 , \8835 , \156 );
and \U$12702 ( \12887 , \9169 , \154 );
nor \U$12703 ( \12888 , \12886 , \12887 );
xnor \U$12704 ( \12889 , \12888 , \163 );
and \U$12705 ( \12890 , \8349 , \296 );
and \U$12706 ( \12891 , \8652 , \168 );
nor \U$12707 ( \12892 , \12890 , \12891 );
xnor \U$12708 ( \12893 , \12892 , \173 );
xor \U$12709 ( \12894 , \12889 , \12893 );
and \U$12710 ( \12895 , \7700 , \438 );
and \U$12711 ( \12896 , \8057 , \336 );
nor \U$12712 ( \12897 , \12895 , \12896 );
xnor \U$12713 ( \12898 , \12897 , \320 );
xor \U$12714 ( \12899 , \12894 , \12898 );
xor \U$12715 ( \12900 , \12885 , \12899 );
not \U$12716 ( \12901 , \237 );
and \U$12717 ( \12902 , \10206 , \245 );
and \U$12718 ( \12903 , \10584 , \243 );
nor \U$12719 ( \12904 , \12902 , \12903 );
xnor \U$12720 ( \12905 , \12904 , \252 );
xor \U$12721 ( \12906 , \12901 , \12905 );
and \U$12722 ( \12907 , \9465 , \141 );
and \U$12723 ( \12908 , \9897 , \139 );
nor \U$12724 ( \12909 , \12907 , \12908 );
xnor \U$12725 ( \12910 , \12909 , \148 );
xor \U$12726 ( \12911 , \12906 , \12910 );
xor \U$12727 ( \12912 , \12900 , \12911 );
xor \U$12728 ( \12913 , \12881 , \12912 );
xor \U$12729 ( \12914 , \12855 , \12913 );
and \U$12730 ( \12915 , \12725 , \12769 );
and \U$12731 ( \12916 , \12769 , \12786 );
and \U$12732 ( \12917 , \12725 , \12786 );
or \U$12733 ( \12918 , \12915 , \12916 , \12917 );
and \U$12734 ( \12919 , \12669 , \12673 );
and \U$12735 ( \12920 , \12673 , \12678 );
and \U$12736 ( \12921 , \12669 , \12678 );
or \U$12737 ( \12922 , \12919 , \12920 , \12921 );
and \U$12738 ( \12923 , \12683 , \12687 );
and \U$12739 ( \12924 , \12687 , \12692 );
and \U$12740 ( \12925 , \12683 , \12692 );
or \U$12741 ( \12926 , \12923 , \12924 , \12925 );
xor \U$12742 ( \12927 , \12922 , \12926 );
and \U$12743 ( \12928 , \12698 , \12702 );
and \U$12744 ( \12929 , \12702 , \12707 );
and \U$12745 ( \12930 , \12698 , \12707 );
or \U$12746 ( \12931 , \12928 , \12929 , \12930 );
xor \U$12747 ( \12932 , \12927 , \12931 );
and \U$12748 ( \12933 , \12729 , \12733 );
and \U$12749 ( \12934 , \12733 , \12738 );
and \U$12750 ( \12935 , \12729 , \12738 );
or \U$12751 ( \12936 , \12933 , \12934 , \12935 );
and \U$12752 ( \12937 , \12743 , \12747 );
and \U$12753 ( \12938 , \12747 , \12752 );
and \U$12754 ( \12939 , \12743 , \12752 );
or \U$12755 ( \12940 , \12937 , \12938 , \12939 );
xor \U$12756 ( \12941 , \12936 , \12940 );
and \U$12757 ( \12942 , \12758 , \12762 );
and \U$12758 ( \12943 , \12762 , \12767 );
and \U$12759 ( \12944 , \12758 , \12767 );
or \U$12760 ( \12945 , \12942 , \12943 , \12944 );
xor \U$12761 ( \12946 , \12941 , \12945 );
xor \U$12762 ( \12947 , \12932 , \12946 );
and \U$12763 ( \12948 , \12624 , \12628 );
and \U$12764 ( \12949 , \12628 , \12633 );
and \U$12765 ( \12950 , \12624 , \12633 );
or \U$12766 ( \12951 , \12948 , \12949 , \12950 );
and \U$12767 ( \12952 , \12638 , \12642 );
and \U$12768 ( \12953 , \12642 , \12647 );
and \U$12769 ( \12954 , \12638 , \12647 );
or \U$12770 ( \12955 , \12952 , \12953 , \12954 );
xor \U$12771 ( \12956 , \12951 , \12955 );
and \U$12772 ( \12957 , \12653 , \12657 );
and \U$12773 ( \12958 , \12657 , \12662 );
and \U$12774 ( \12959 , \12653 , \12662 );
or \U$12775 ( \12960 , \12957 , \12958 , \12959 );
xor \U$12776 ( \12961 , \12956 , \12960 );
xor \U$12777 ( \12962 , \12947 , \12961 );
xor \U$12778 ( \12963 , \12918 , \12962 );
and \U$12779 ( \12964 , \7231 , \1086 );
and \U$12780 ( \12965 , \7556 , \508 );
nor \U$12781 ( \12966 , \12964 , \12965 );
xnor \U$12782 ( \12967 , \12966 , \487 );
and \U$12783 ( \12968 , \6790 , \1301 );
and \U$12784 ( \12969 , \6945 , \1246 );
nor \U$12785 ( \12970 , \12968 , \12969 );
xnor \U$12786 ( \12971 , \12970 , \1205 );
xor \U$12787 ( \12972 , \12967 , \12971 );
and \U$12788 ( \12973 , \6281 , \1578 );
and \U$12789 ( \12974 , \6514 , \1431 );
nor \U$12790 ( \12975 , \12973 , \12974 );
xnor \U$12791 ( \12976 , \12975 , \1436 );
xor \U$12792 ( \12977 , \12972 , \12976 );
and \U$12793 ( \12978 , \4364 , \2669 );
and \U$12794 ( \12979 , \4654 , \2538 );
nor \U$12795 ( \12980 , \12978 , \12979 );
xnor \U$12796 ( \12981 , \12980 , \2534 );
and \U$12797 ( \12982 , \3912 , \3103 );
and \U$12798 ( \12983 , \4160 , \2934 );
nor \U$12799 ( \12984 , \12982 , \12983 );
xnor \U$12800 ( \12985 , \12984 , \2839 );
xor \U$12801 ( \12986 , \12981 , \12985 );
and \U$12802 ( \12987 , \3646 , \3357 );
and \U$12803 ( \12988 , \3736 , \3255 );
nor \U$12804 ( \12989 , \12987 , \12988 );
xnor \U$12805 ( \12990 , \12989 , \3156 );
xor \U$12806 ( \12991 , \12986 , \12990 );
xor \U$12807 ( \12992 , \12977 , \12991 );
and \U$12808 ( \12993 , \5674 , \1824 );
and \U$12809 ( \12994 , \6030 , \1739 );
nor \U$12810 ( \12995 , \12993 , \12994 );
xnor \U$12811 ( \12996 , \12995 , \1697 );
and \U$12812 ( \12997 , \5156 , \2121 );
and \U$12813 ( \12998 , \5469 , \2008 );
nor \U$12814 ( \12999 , \12997 , \12998 );
xnor \U$12815 ( \13000 , \12999 , \1961 );
xor \U$12816 ( \13001 , \12996 , \13000 );
and \U$12817 ( \13002 , \4749 , \2400 );
and \U$12818 ( \13003 , \4922 , \2246 );
nor \U$12819 ( \13004 , \13002 , \13003 );
xnor \U$12820 ( \13005 , \13004 , \2195 );
xor \U$12821 ( \13006 , \13001 , \13005 );
xor \U$12822 ( \13007 , \12992 , \13006 );
and \U$12823 ( \13008 , \3143 , \3813 );
and \U$12824 ( \13009 , \3395 , \3557 );
nor \U$12825 ( \13010 , \13008 , \13009 );
xnor \U$12826 ( \13011 , \13010 , \3562 );
and \U$12827 ( \13012 , \2826 , \4132 );
and \U$12828 ( \13013 , \3037 , \4012 );
nor \U$12829 ( \13014 , \13012 , \13013 );
xnor \U$12830 ( \13015 , \13014 , \3925 );
xor \U$12831 ( \13016 , \13011 , \13015 );
and \U$12832 ( \13017 , \2521 , \4581 );
and \U$12833 ( \13018 , \2757 , \4424 );
nor \U$12834 ( \13019 , \13017 , \13018 );
xnor \U$12835 ( \13020 , \13019 , \4377 );
xor \U$12836 ( \13021 , \13016 , \13020 );
and \U$12837 ( \13022 , \1484 , \6401 );
and \U$12838 ( \13023 , \1601 , \6143 );
nor \U$12839 ( \13024 , \13022 , \13023 );
xnor \U$12840 ( \13025 , \13024 , \6148 );
and \U$12841 ( \13026 , \1192 , \7055 );
and \U$12842 ( \13027 , \1333 , \6675 );
nor \U$12843 ( \13028 , \13026 , \13027 );
xnor \U$12844 ( \13029 , \13028 , \6680 );
xor \U$12845 ( \13030 , \13025 , \13029 );
and \U$12846 ( \13031 , \474 , \7489 );
and \U$12847 ( \13032 , \1147 , \7137 );
nor \U$12848 ( \13033 , \13031 , \13032 );
xnor \U$12849 ( \13034 , \13033 , \7142 );
xor \U$12850 ( \13035 , \13030 , \13034 );
xor \U$12851 ( \13036 , \13021 , \13035 );
and \U$12852 ( \13037 , \2182 , \5011 );
and \U$12853 ( \13038 , \2366 , \4878 );
nor \U$12854 ( \13039 , \13037 , \13038 );
xnor \U$12855 ( \13040 , \13039 , \4762 );
and \U$12856 ( \13041 , \1948 , \5485 );
and \U$12857 ( \13042 , \2090 , \5275 );
nor \U$12858 ( \13043 , \13041 , \13042 );
xnor \U$12859 ( \13044 , \13043 , \5169 );
xor \U$12860 ( \13045 , \13040 , \13044 );
and \U$12861 ( \13046 , \1684 , \5996 );
and \U$12862 ( \13047 , \1802 , \5695 );
nor \U$12863 ( \13048 , \13046 , \13047 );
xnor \U$12864 ( \13049 , \13048 , \5687 );
xor \U$12865 ( \13050 , \13045 , \13049 );
xor \U$12866 ( \13051 , \13036 , \13050 );
xor \U$12867 ( \13052 , \13007 , \13051 );
and \U$12868 ( \13053 , \12778 , \12782 );
and \U$12869 ( \13054 , \12782 , \12784 );
and \U$12870 ( \13055 , \12778 , \12784 );
or \U$12871 ( \13056 , \13053 , \13054 , \13055 );
and \U$12872 ( \13057 , \217 , \9765 );
and \U$12873 ( \13058 , \189 , \9644 );
nor \U$12874 ( \13059 , \13057 , \13058 );
xnor \U$12875 ( \13060 , \13059 , \9478 );
and \U$12876 ( \13061 , \232 , \10408 );
and \U$12877 ( \13062 , \209 , \10116 );
nor \U$12878 ( \13063 , \13061 , \13062 );
xnor \U$12879 ( \13064 , \13063 , \10121 );
xor \U$12880 ( \13065 , \13060 , \13064 );
and \U$12881 ( \13066 , \224 , \10118 );
xor \U$12882 ( \13067 , \13065 , \13066 );
xor \U$12883 ( \13068 , \13056 , \13067 );
and \U$12884 ( \13069 , \307 , \8019 );
and \U$12885 ( \13070 , \412 , \7830 );
nor \U$12886 ( \13071 , \13069 , \13070 );
xnor \U$12887 ( \13072 , \13071 , \7713 );
and \U$12888 ( \13073 , \185 , \8540 );
and \U$12889 ( \13074 , \261 , \8292 );
nor \U$12890 ( \13075 , \13073 , \13074 );
xnor \U$12891 ( \13076 , \13075 , \8297 );
xor \U$12892 ( \13077 , \13072 , \13076 );
and \U$12893 ( \13078 , \197 , \9333 );
and \U$12894 ( \13079 , \178 , \9006 );
nor \U$12895 ( \13080 , \13078 , \13079 );
xnor \U$12896 ( \13081 , \13080 , \8848 );
xor \U$12897 ( \13082 , \13077 , \13081 );
xor \U$12898 ( \13083 , \13068 , \13082 );
xor \U$12899 ( \13084 , \13052 , \13083 );
xor \U$12900 ( \13085 , \12963 , \13084 );
xor \U$12901 ( \13086 , \12914 , \13085 );
xor \U$12902 ( \13087 , \12841 , \13086 );
xor \U$12903 ( \13088 , \12832 , \13087 );
and \U$12904 ( \13089 , \12504 , \12505 );
and \U$12905 ( \13090 , \12505 , \12791 );
and \U$12906 ( \13091 , \12504 , \12791 );
or \U$12907 ( \13092 , \13089 , \13090 , \13091 );
xor \U$12908 ( \13093 , \13088 , \13092 );
and \U$12909 ( \13094 , \12792 , \12796 );
and \U$12910 ( \13095 , \12797 , \12800 );
or \U$12911 ( \13096 , \13094 , \13095 );
xor \U$12912 ( \13097 , \13093 , \13096 );
buf g550d_GF_PartitionCandidate( \13098_nG550d , \13097 );
buf \U$12913 ( \13099 , \13098_nG550d );
and \U$12914 ( \13100 , \12811 , \12815 );
and \U$12915 ( \13101 , \12815 , \12830 );
and \U$12916 ( \13102 , \12811 , \12830 );
or \U$12917 ( \13103 , \13100 , \13101 , \13102 );
and \U$12918 ( \13104 , \12836 , \12840 );
and \U$12919 ( \13105 , \12840 , \13086 );
and \U$12920 ( \13106 , \12836 , \13086 );
or \U$12921 ( \13107 , \13104 , \13105 , \13106 );
and \U$12922 ( \13108 , \12820 , \12824 );
and \U$12923 ( \13109 , \12824 , \12829 );
and \U$12924 ( \13110 , \12820 , \12829 );
or \U$12925 ( \13111 , \13108 , \13109 , \13110 );
and \U$12926 ( \13112 , \12855 , \12913 );
and \U$12927 ( \13113 , \12913 , \13085 );
and \U$12928 ( \13114 , \12855 , \13085 );
or \U$12929 ( \13115 , \13112 , \13113 , \13114 );
xor \U$12930 ( \13116 , \13111 , \13115 );
and \U$12931 ( \13117 , \12932 , \12946 );
and \U$12932 ( \13118 , \12946 , \12961 );
and \U$12933 ( \13119 , \12932 , \12961 );
or \U$12934 ( \13120 , \13117 , \13118 , \13119 );
and \U$12935 ( \13121 , \13007 , \13051 );
and \U$12936 ( \13122 , \13051 , \13083 );
and \U$12937 ( \13123 , \13007 , \13083 );
or \U$12938 ( \13124 , \13121 , \13122 , \13123 );
xor \U$12939 ( \13125 , \13120 , \13124 );
and \U$12940 ( \13126 , \13011 , \13015 );
and \U$12941 ( \13127 , \13015 , \13020 );
and \U$12942 ( \13128 , \13011 , \13020 );
or \U$12943 ( \13129 , \13126 , \13127 , \13128 );
and \U$12944 ( \13130 , \12981 , \12985 );
and \U$12945 ( \13131 , \12985 , \12990 );
and \U$12946 ( \13132 , \12981 , \12990 );
or \U$12947 ( \13133 , \13130 , \13131 , \13132 );
xor \U$12948 ( \13134 , \13129 , \13133 );
and \U$12949 ( \13135 , \12996 , \13000 );
and \U$12950 ( \13136 , \13000 , \13005 );
and \U$12951 ( \13137 , \12996 , \13005 );
or \U$12952 ( \13138 , \13135 , \13136 , \13137 );
xor \U$12953 ( \13139 , \13134 , \13138 );
xor \U$12954 ( \13140 , \13125 , \13139 );
xor \U$12955 ( \13141 , \13116 , \13140 );
xor \U$12956 ( \13142 , \13107 , \13141 );
and \U$12957 ( \13143 , \12859 , \12863 );
and \U$12958 ( \13144 , \12863 , \12865 );
and \U$12959 ( \13145 , \12859 , \12865 );
or \U$12960 ( \13146 , \13143 , \13144 , \13145 );
and \U$12961 ( \13147 , \12870 , \12874 );
and \U$12962 ( \13148 , \12874 , \12879 );
and \U$12963 ( \13149 , \12870 , \12879 );
or \U$12964 ( \13150 , \13147 , \13148 , \13149 );
xor \U$12965 ( \13151 , \13146 , \13150 );
and \U$12966 ( \13152 , \12885 , \12899 );
and \U$12967 ( \13153 , \12899 , \12911 );
and \U$12968 ( \13154 , \12885 , \12911 );
or \U$12969 ( \13155 , \13152 , \13153 , \13154 );
xor \U$12970 ( \13156 , \13151 , \13155 );
and \U$12971 ( \13157 , \12845 , \12849 );
and \U$12972 ( \13158 , \12849 , \12854 );
and \U$12973 ( \13159 , \12845 , \12854 );
or \U$12974 ( \13160 , \13157 , \13158 , \13159 );
and \U$12975 ( \13161 , \12866 , \12880 );
and \U$12976 ( \13162 , \12880 , \12912 );
and \U$12977 ( \13163 , \12866 , \12912 );
or \U$12978 ( \13164 , \13161 , \13162 , \13163 );
xor \U$12979 ( \13165 , \13160 , \13164 );
and \U$12980 ( \13166 , \12918 , \12962 );
and \U$12981 ( \13167 , \12962 , \13084 );
and \U$12982 ( \13168 , \12918 , \13084 );
or \U$12983 ( \13169 , \13166 , \13167 , \13168 );
xor \U$12984 ( \13170 , \13165 , \13169 );
xor \U$12985 ( \13171 , \13156 , \13170 );
and \U$12986 ( \13172 , \12922 , \12926 );
and \U$12987 ( \13173 , \12926 , \12931 );
and \U$12988 ( \13174 , \12922 , \12931 );
or \U$12989 ( \13175 , \13172 , \13173 , \13174 );
and \U$12990 ( \13176 , \12936 , \12940 );
and \U$12991 ( \13177 , \12940 , \12945 );
and \U$12992 ( \13178 , \12936 , \12945 );
or \U$12993 ( \13179 , \13176 , \13177 , \13178 );
xor \U$12994 ( \13180 , \13175 , \13179 );
and \U$12995 ( \13181 , \12951 , \12955 );
and \U$12996 ( \13182 , \12955 , \12960 );
and \U$12997 ( \13183 , \12951 , \12960 );
or \U$12998 ( \13184 , \13181 , \13182 , \13183 );
xor \U$12999 ( \13185 , \13180 , \13184 );
and \U$13000 ( \13186 , \12977 , \12991 );
and \U$13001 ( \13187 , \12991 , \13006 );
and \U$13002 ( \13188 , \12977 , \13006 );
or \U$13003 ( \13189 , \13186 , \13187 , \13188 );
and \U$13004 ( \13190 , \13021 , \13035 );
and \U$13005 ( \13191 , \13035 , \13050 );
and \U$13006 ( \13192 , \13021 , \13050 );
or \U$13007 ( \13193 , \13190 , \13191 , \13192 );
xor \U$13008 ( \13194 , \13189 , \13193 );
and \U$13009 ( \13195 , \13056 , \13067 );
and \U$13010 ( \13196 , \13067 , \13082 );
and \U$13011 ( \13197 , \13056 , \13082 );
or \U$13012 ( \13198 , \13195 , \13196 , \13197 );
xor \U$13013 ( \13199 , \13194 , \13198 );
xor \U$13014 ( \13200 , \13185 , \13199 );
and \U$13015 ( \13201 , \12889 , \12893 );
and \U$13016 ( \13202 , \12893 , \12898 );
and \U$13017 ( \13203 , \12889 , \12898 );
or \U$13018 ( \13204 , \13201 , \13202 , \13203 );
and \U$13019 ( \13205 , \12901 , \12905 );
and \U$13020 ( \13206 , \12905 , \12910 );
and \U$13021 ( \13207 , \12901 , \12910 );
or \U$13022 ( \13208 , \13205 , \13206 , \13207 );
xor \U$13023 ( \13209 , \13204 , \13208 );
and \U$13024 ( \13210 , \12967 , \12971 );
and \U$13025 ( \13211 , \12971 , \12976 );
and \U$13026 ( \13212 , \12967 , \12976 );
or \U$13027 ( \13213 , \13210 , \13211 , \13212 );
xor \U$13028 ( \13214 , \13209 , \13213 );
and \U$13029 ( \13215 , \10584 , \245 );
not \U$13030 ( \13216 , \13215 );
xnor \U$13031 ( \13217 , \13216 , \252 );
and \U$13032 ( \13218 , \9897 , \141 );
and \U$13033 ( \13219 , \10206 , \139 );
nor \U$13034 ( \13220 , \13218 , \13219 );
xnor \U$13035 ( \13221 , \13220 , \148 );
xor \U$13036 ( \13222 , \13217 , \13221 );
and \U$13037 ( \13223 , \9169 , \156 );
and \U$13038 ( \13224 , \9465 , \154 );
nor \U$13039 ( \13225 , \13223 , \13224 );
xnor \U$13040 ( \13226 , \13225 , \163 );
xor \U$13041 ( \13227 , \13222 , \13226 );
and \U$13042 ( \13228 , \8652 , \296 );
and \U$13043 ( \13229 , \8835 , \168 );
nor \U$13044 ( \13230 , \13228 , \13229 );
xnor \U$13045 ( \13231 , \13230 , \173 );
and \U$13046 ( \13232 , \8057 , \438 );
and \U$13047 ( \13233 , \8349 , \336 );
nor \U$13048 ( \13234 , \13232 , \13233 );
xnor \U$13049 ( \13235 , \13234 , \320 );
xor \U$13050 ( \13236 , \13231 , \13235 );
and \U$13051 ( \13237 , \7556 , \1086 );
and \U$13052 ( \13238 , \7700 , \508 );
nor \U$13053 ( \13239 , \13237 , \13238 );
xnor \U$13054 ( \13240 , \13239 , \487 );
xor \U$13055 ( \13241 , \13236 , \13240 );
xor \U$13056 ( \13242 , \13227 , \13241 );
and \U$13057 ( \13243 , \4160 , \3103 );
and \U$13058 ( \13244 , \4364 , \2934 );
nor \U$13059 ( \13245 , \13243 , \13244 );
xnor \U$13060 ( \13246 , \13245 , \2839 );
and \U$13061 ( \13247 , \3736 , \3357 );
and \U$13062 ( \13248 , \3912 , \3255 );
nor \U$13063 ( \13249 , \13247 , \13248 );
xnor \U$13064 ( \13250 , \13249 , \3156 );
xor \U$13065 ( \13251 , \13246 , \13250 );
and \U$13066 ( \13252 , \3395 , \3813 );
and \U$13067 ( \13253 , \3646 , \3557 );
nor \U$13068 ( \13254 , \13252 , \13253 );
xnor \U$13069 ( \13255 , \13254 , \3562 );
xor \U$13070 ( \13256 , \13251 , \13255 );
and \U$13071 ( \13257 , \6945 , \1301 );
and \U$13072 ( \13258 , \7231 , \1246 );
nor \U$13073 ( \13259 , \13257 , \13258 );
xnor \U$13074 ( \13260 , \13259 , \1205 );
and \U$13075 ( \13261 , \6514 , \1578 );
and \U$13076 ( \13262 , \6790 , \1431 );
nor \U$13077 ( \13263 , \13261 , \13262 );
xnor \U$13078 ( \13264 , \13263 , \1436 );
xor \U$13079 ( \13265 , \13260 , \13264 );
and \U$13080 ( \13266 , \6030 , \1824 );
and \U$13081 ( \13267 , \6281 , \1739 );
nor \U$13082 ( \13268 , \13266 , \13267 );
xnor \U$13083 ( \13269 , \13268 , \1697 );
xor \U$13084 ( \13270 , \13265 , \13269 );
xor \U$13085 ( \13271 , \13256 , \13270 );
and \U$13086 ( \13272 , \5469 , \2121 );
and \U$13087 ( \13273 , \5674 , \2008 );
nor \U$13088 ( \13274 , \13272 , \13273 );
xnor \U$13089 ( \13275 , \13274 , \1961 );
and \U$13090 ( \13276 , \4922 , \2400 );
and \U$13091 ( \13277 , \5156 , \2246 );
nor \U$13092 ( \13278 , \13276 , \13277 );
xnor \U$13093 ( \13279 , \13278 , \2195 );
xor \U$13094 ( \13280 , \13275 , \13279 );
and \U$13095 ( \13281 , \4654 , \2669 );
and \U$13096 ( \13282 , \4749 , \2538 );
nor \U$13097 ( \13283 , \13281 , \13282 );
xnor \U$13098 ( \13284 , \13283 , \2534 );
xor \U$13099 ( \13285 , \13280 , \13284 );
xor \U$13100 ( \13286 , \13271 , \13285 );
xor \U$13101 ( \13287 , \13242 , \13286 );
xor \U$13102 ( \13288 , \13214 , \13287 );
and \U$13103 ( \13289 , \13025 , \13029 );
and \U$13104 ( \13290 , \13029 , \13034 );
and \U$13105 ( \13291 , \13025 , \13034 );
or \U$13106 ( \13292 , \13289 , \13290 , \13291 );
and \U$13107 ( \13293 , \13040 , \13044 );
and \U$13108 ( \13294 , \13044 , \13049 );
and \U$13109 ( \13295 , \13040 , \13049 );
or \U$13110 ( \13296 , \13293 , \13294 , \13295 );
xor \U$13111 ( \13297 , \13292 , \13296 );
and \U$13112 ( \13298 , \13072 , \13076 );
and \U$13113 ( \13299 , \13076 , \13081 );
and \U$13114 ( \13300 , \13072 , \13081 );
or \U$13115 ( \13301 , \13298 , \13299 , \13300 );
xor \U$13116 ( \13302 , \13297 , \13301 );
and \U$13117 ( \13303 , \3037 , \4132 );
and \U$13118 ( \13304 , \3143 , \4012 );
nor \U$13119 ( \13305 , \13303 , \13304 );
xnor \U$13120 ( \13306 , \13305 , \3925 );
and \U$13121 ( \13307 , \2757 , \4581 );
and \U$13122 ( \13308 , \2826 , \4424 );
nor \U$13123 ( \13309 , \13307 , \13308 );
xnor \U$13124 ( \13310 , \13309 , \4377 );
xor \U$13125 ( \13311 , \13306 , \13310 );
and \U$13126 ( \13312 , \2366 , \5011 );
and \U$13127 ( \13313 , \2521 , \4878 );
nor \U$13128 ( \13314 , \13312 , \13313 );
xnor \U$13129 ( \13315 , \13314 , \4762 );
xor \U$13130 ( \13316 , \13311 , \13315 );
and \U$13131 ( \13317 , \1333 , \7055 );
and \U$13132 ( \13318 , \1484 , \6675 );
nor \U$13133 ( \13319 , \13317 , \13318 );
xnor \U$13134 ( \13320 , \13319 , \6680 );
and \U$13135 ( \13321 , \1147 , \7489 );
and \U$13136 ( \13322 , \1192 , \7137 );
nor \U$13137 ( \13323 , \13321 , \13322 );
xnor \U$13138 ( \13324 , \13323 , \7142 );
xor \U$13139 ( \13325 , \13320 , \13324 );
and \U$13140 ( \13326 , \412 , \8019 );
and \U$13141 ( \13327 , \474 , \7830 );
nor \U$13142 ( \13328 , \13326 , \13327 );
xnor \U$13143 ( \13329 , \13328 , \7713 );
xor \U$13144 ( \13330 , \13325 , \13329 );
xor \U$13145 ( \13331 , \13316 , \13330 );
and \U$13146 ( \13332 , \2090 , \5485 );
and \U$13147 ( \13333 , \2182 , \5275 );
nor \U$13148 ( \13334 , \13332 , \13333 );
xnor \U$13149 ( \13335 , \13334 , \5169 );
and \U$13150 ( \13336 , \1802 , \5996 );
and \U$13151 ( \13337 , \1948 , \5695 );
nor \U$13152 ( \13338 , \13336 , \13337 );
xnor \U$13153 ( \13339 , \13338 , \5687 );
xor \U$13154 ( \13340 , \13335 , \13339 );
and \U$13155 ( \13341 , \1601 , \6401 );
and \U$13156 ( \13342 , \1684 , \6143 );
nor \U$13157 ( \13343 , \13341 , \13342 );
xnor \U$13158 ( \13344 , \13343 , \6148 );
xor \U$13159 ( \13345 , \13340 , \13344 );
xor \U$13160 ( \13346 , \13331 , \13345 );
xor \U$13161 ( \13347 , \13302 , \13346 );
and \U$13162 ( \13348 , \13060 , \13064 );
and \U$13163 ( \13349 , \13064 , \13066 );
and \U$13164 ( \13350 , \13060 , \13066 );
or \U$13165 ( \13351 , \13348 , \13349 , \13350 );
and \U$13166 ( \13352 , \261 , \8540 );
and \U$13167 ( \13353 , \307 , \8292 );
nor \U$13168 ( \13354 , \13352 , \13353 );
xnor \U$13169 ( \13355 , \13354 , \8297 );
and \U$13170 ( \13356 , \178 , \9333 );
and \U$13171 ( \13357 , \185 , \9006 );
nor \U$13172 ( \13358 , \13356 , \13357 );
xnor \U$13173 ( \13359 , \13358 , \8848 );
xor \U$13174 ( \13360 , \13355 , \13359 );
and \U$13175 ( \13361 , \189 , \9765 );
and \U$13176 ( \13362 , \197 , \9644 );
nor \U$13177 ( \13363 , \13361 , \13362 );
xnor \U$13178 ( \13364 , \13363 , \9478 );
xor \U$13179 ( \13365 , \13360 , \13364 );
xor \U$13180 ( \13366 , \13351 , \13365 );
and \U$13181 ( \13367 , \209 , \10408 );
and \U$13182 ( \13368 , \217 , \10116 );
nor \U$13183 ( \13369 , \13367 , \13368 );
xnor \U$13184 ( \13370 , \13369 , \10121 );
and \U$13185 ( \13371 , \232 , \10118 );
xnor \U$13186 ( \13372 , \13370 , \13371 );
xor \U$13187 ( \13373 , \13366 , \13372 );
xor \U$13188 ( \13374 , \13347 , \13373 );
xor \U$13189 ( \13375 , \13288 , \13374 );
xor \U$13190 ( \13376 , \13200 , \13375 );
xor \U$13191 ( \13377 , \13171 , \13376 );
xor \U$13192 ( \13378 , \13142 , \13377 );
xor \U$13193 ( \13379 , \13103 , \13378 );
and \U$13194 ( \13380 , \12807 , \12831 );
and \U$13195 ( \13381 , \12831 , \13087 );
and \U$13196 ( \13382 , \12807 , \13087 );
or \U$13197 ( \13383 , \13380 , \13381 , \13382 );
xor \U$13198 ( \13384 , \13379 , \13383 );
and \U$13199 ( \13385 , \13088 , \13092 );
and \U$13200 ( \13386 , \13093 , \13096 );
or \U$13201 ( \13387 , \13385 , \13386 );
xor \U$13202 ( \13388 , \13384 , \13387 );
buf g550b_GF_PartitionCandidate( \13389_nG550b , \13388 );
buf \U$13203 ( \13390 , \13389_nG550b );
and \U$13204 ( \13391 , \13107 , \13141 );
and \U$13205 ( \13392 , \13141 , \13377 );
and \U$13206 ( \13393 , \13107 , \13377 );
or \U$13207 ( \13394 , \13391 , \13392 , \13393 );
and \U$13208 ( \13395 , \13111 , \13115 );
and \U$13209 ( \13396 , \13115 , \13140 );
and \U$13210 ( \13397 , \13111 , \13140 );
or \U$13211 ( \13398 , \13395 , \13396 , \13397 );
and \U$13212 ( \13399 , \13156 , \13170 );
and \U$13213 ( \13400 , \13170 , \13376 );
and \U$13214 ( \13401 , \13156 , \13376 );
or \U$13215 ( \13402 , \13399 , \13400 , \13401 );
xor \U$13216 ( \13403 , \13398 , \13402 );
and \U$13217 ( \13404 , \13146 , \13150 );
and \U$13218 ( \13405 , \13150 , \13155 );
and \U$13219 ( \13406 , \13146 , \13155 );
or \U$13220 ( \13407 , \13404 , \13405 , \13406 );
and \U$13221 ( \13408 , \13120 , \13124 );
and \U$13222 ( \13409 , \13124 , \13139 );
and \U$13223 ( \13410 , \13120 , \13139 );
or \U$13224 ( \13411 , \13408 , \13409 , \13410 );
xor \U$13225 ( \13412 , \13407 , \13411 );
and \U$13226 ( \13413 , \13214 , \13287 );
and \U$13227 ( \13414 , \13287 , \13374 );
and \U$13228 ( \13415 , \13214 , \13374 );
or \U$13229 ( \13416 , \13413 , \13414 , \13415 );
xor \U$13230 ( \13417 , \13412 , \13416 );
xor \U$13231 ( \13418 , \13403 , \13417 );
xor \U$13232 ( \13419 , \13394 , \13418 );
and \U$13233 ( \13420 , \13160 , \13164 );
and \U$13234 ( \13421 , \13164 , \13169 );
and \U$13235 ( \13422 , \13160 , \13169 );
or \U$13236 ( \13423 , \13420 , \13421 , \13422 );
and \U$13237 ( \13424 , \13185 , \13199 );
and \U$13238 ( \13425 , \13199 , \13375 );
and \U$13239 ( \13426 , \13185 , \13375 );
or \U$13240 ( \13427 , \13424 , \13425 , \13426 );
xor \U$13241 ( \13428 , \13423 , \13427 );
and \U$13242 ( \13429 , \13175 , \13179 );
and \U$13243 ( \13430 , \13179 , \13184 );
and \U$13244 ( \13431 , \13175 , \13184 );
or \U$13245 ( \13432 , \13429 , \13430 , \13431 );
and \U$13246 ( \13433 , \13189 , \13193 );
and \U$13247 ( \13434 , \13193 , \13198 );
and \U$13248 ( \13435 , \13189 , \13198 );
or \U$13249 ( \13436 , \13433 , \13434 , \13435 );
xor \U$13250 ( \13437 , \13432 , \13436 );
and \U$13251 ( \13438 , \13227 , \13241 );
and \U$13252 ( \13439 , \13241 , \13286 );
and \U$13253 ( \13440 , \13227 , \13286 );
or \U$13254 ( \13441 , \13438 , \13439 , \13440 );
xor \U$13255 ( \13442 , \13437 , \13441 );
and \U$13256 ( \13443 , \13302 , \13346 );
and \U$13257 ( \13444 , \13346 , \13373 );
and \U$13258 ( \13445 , \13302 , \13373 );
or \U$13259 ( \13446 , \13443 , \13444 , \13445 );
and \U$13260 ( \13447 , \13260 , \13264 );
and \U$13261 ( \13448 , \13264 , \13269 );
and \U$13262 ( \13449 , \13260 , \13269 );
or \U$13263 ( \13450 , \13447 , \13448 , \13449 );
and \U$13264 ( \13451 , \13217 , \13221 );
and \U$13265 ( \13452 , \13221 , \13226 );
and \U$13266 ( \13453 , \13217 , \13226 );
or \U$13267 ( \13454 , \13451 , \13452 , \13453 );
xor \U$13268 ( \13455 , \13450 , \13454 );
and \U$13269 ( \13456 , \13231 , \13235 );
and \U$13270 ( \13457 , \13235 , \13240 );
and \U$13271 ( \13458 , \13231 , \13240 );
or \U$13272 ( \13459 , \13456 , \13457 , \13458 );
xor \U$13273 ( \13460 , \13455 , \13459 );
xor \U$13274 ( \13461 , \13446 , \13460 );
and \U$13275 ( \13462 , \13246 , \13250 );
and \U$13276 ( \13463 , \13250 , \13255 );
and \U$13277 ( \13464 , \13246 , \13255 );
or \U$13278 ( \13465 , \13462 , \13463 , \13464 );
and \U$13279 ( \13466 , \13306 , \13310 );
and \U$13280 ( \13467 , \13310 , \13315 );
and \U$13281 ( \13468 , \13306 , \13315 );
or \U$13282 ( \13469 , \13466 , \13467 , \13468 );
xor \U$13283 ( \13470 , \13465 , \13469 );
and \U$13284 ( \13471 , \13275 , \13279 );
and \U$13285 ( \13472 , \13279 , \13284 );
and \U$13286 ( \13473 , \13275 , \13284 );
or \U$13287 ( \13474 , \13471 , \13472 , \13473 );
xor \U$13288 ( \13475 , \13470 , \13474 );
and \U$13289 ( \13476 , \13320 , \13324 );
and \U$13290 ( \13477 , \13324 , \13329 );
and \U$13291 ( \13478 , \13320 , \13329 );
or \U$13292 ( \13479 , \13476 , \13477 , \13478 );
and \U$13293 ( \13480 , \13335 , \13339 );
and \U$13294 ( \13481 , \13339 , \13344 );
and \U$13295 ( \13482 , \13335 , \13344 );
or \U$13296 ( \13483 , \13480 , \13481 , \13482 );
xor \U$13297 ( \13484 , \13479 , \13483 );
and \U$13298 ( \13485 , \13355 , \13359 );
and \U$13299 ( \13486 , \13359 , \13364 );
and \U$13300 ( \13487 , \13355 , \13364 );
or \U$13301 ( \13488 , \13485 , \13486 , \13487 );
xor \U$13302 ( \13489 , \13484 , \13488 );
xor \U$13303 ( \13490 , \13475 , \13489 );
or \U$13304 ( \13491 , \13370 , \13371 );
and \U$13305 ( \13492 , \217 , \10408 );
and \U$13306 ( \13493 , \189 , \10116 );
nor \U$13307 ( \13494 , \13492 , \13493 );
xnor \U$13308 ( \13495 , \13494 , \10121 );
xor \U$13309 ( \13496 , \13491 , \13495 );
and \U$13310 ( \13497 , \209 , \10118 );
xor \U$13311 ( \13498 , \13496 , \13497 );
xor \U$13312 ( \13499 , \13490 , \13498 );
xor \U$13313 ( \13500 , \13461 , \13499 );
xor \U$13314 ( \13501 , \13442 , \13500 );
and \U$13315 ( \13502 , \13204 , \13208 );
and \U$13316 ( \13503 , \13208 , \13213 );
and \U$13317 ( \13504 , \13204 , \13213 );
or \U$13318 ( \13505 , \13502 , \13503 , \13504 );
and \U$13319 ( \13506 , \13129 , \13133 );
and \U$13320 ( \13507 , \13133 , \13138 );
and \U$13321 ( \13508 , \13129 , \13138 );
or \U$13322 ( \13509 , \13506 , \13507 , \13508 );
xor \U$13323 ( \13510 , \13505 , \13509 );
and \U$13324 ( \13511 , \13292 , \13296 );
and \U$13325 ( \13512 , \13296 , \13301 );
and \U$13326 ( \13513 , \13292 , \13301 );
or \U$13327 ( \13514 , \13511 , \13512 , \13513 );
xor \U$13328 ( \13515 , \13510 , \13514 );
and \U$13329 ( \13516 , \13256 , \13270 );
and \U$13330 ( \13517 , \13270 , \13285 );
and \U$13331 ( \13518 , \13256 , \13285 );
or \U$13332 ( \13519 , \13516 , \13517 , \13518 );
and \U$13333 ( \13520 , \13316 , \13330 );
and \U$13334 ( \13521 , \13330 , \13345 );
and \U$13335 ( \13522 , \13316 , \13345 );
or \U$13336 ( \13523 , \13520 , \13521 , \13522 );
xor \U$13337 ( \13524 , \13519 , \13523 );
and \U$13338 ( \13525 , \13351 , \13365 );
and \U$13339 ( \13526 , \13365 , \13372 );
and \U$13340 ( \13527 , \13351 , \13372 );
or \U$13341 ( \13528 , \13525 , \13526 , \13527 );
xor \U$13342 ( \13529 , \13524 , \13528 );
xor \U$13343 ( \13530 , \13515 , \13529 );
and \U$13344 ( \13531 , \1484 , \7055 );
and \U$13345 ( \13532 , \1601 , \6675 );
nor \U$13346 ( \13533 , \13531 , \13532 );
xnor \U$13347 ( \13534 , \13533 , \6680 );
and \U$13348 ( \13535 , \1192 , \7489 );
and \U$13349 ( \13536 , \1333 , \7137 );
nor \U$13350 ( \13537 , \13535 , \13536 );
xnor \U$13351 ( \13538 , \13537 , \7142 );
xor \U$13352 ( \13539 , \13534 , \13538 );
and \U$13353 ( \13540 , \474 , \8019 );
and \U$13354 ( \13541 , \1147 , \7830 );
nor \U$13355 ( \13542 , \13540 , \13541 );
xnor \U$13356 ( \13543 , \13542 , \7713 );
xor \U$13357 ( \13544 , \13539 , \13543 );
and \U$13358 ( \13545 , \307 , \8540 );
and \U$13359 ( \13546 , \412 , \8292 );
nor \U$13360 ( \13547 , \13545 , \13546 );
xnor \U$13361 ( \13548 , \13547 , \8297 );
and \U$13362 ( \13549 , \185 , \9333 );
and \U$13363 ( \13550 , \261 , \9006 );
nor \U$13364 ( \13551 , \13549 , \13550 );
xnor \U$13365 ( \13552 , \13551 , \8848 );
xor \U$13366 ( \13553 , \13548 , \13552 );
and \U$13367 ( \13554 , \197 , \9765 );
and \U$13368 ( \13555 , \178 , \9644 );
nor \U$13369 ( \13556 , \13554 , \13555 );
xnor \U$13370 ( \13557 , \13556 , \9478 );
xor \U$13371 ( \13558 , \13553 , \13557 );
xor \U$13372 ( \13559 , \13544 , \13558 );
and \U$13373 ( \13560 , \2182 , \5485 );
and \U$13374 ( \13561 , \2366 , \5275 );
nor \U$13375 ( \13562 , \13560 , \13561 );
xnor \U$13376 ( \13563 , \13562 , \5169 );
and \U$13377 ( \13564 , \1948 , \5996 );
and \U$13378 ( \13565 , \2090 , \5695 );
nor \U$13379 ( \13566 , \13564 , \13565 );
xnor \U$13380 ( \13567 , \13566 , \5687 );
xor \U$13381 ( \13568 , \13563 , \13567 );
and \U$13382 ( \13569 , \1684 , \6401 );
and \U$13383 ( \13570 , \1802 , \6143 );
nor \U$13384 ( \13571 , \13569 , \13570 );
xnor \U$13385 ( \13572 , \13571 , \6148 );
xor \U$13386 ( \13573 , \13568 , \13572 );
xor \U$13387 ( \13574 , \13559 , \13573 );
and \U$13388 ( \13575 , \3143 , \4132 );
and \U$13389 ( \13576 , \3395 , \4012 );
nor \U$13390 ( \13577 , \13575 , \13576 );
xnor \U$13391 ( \13578 , \13577 , \3925 );
and \U$13392 ( \13579 , \2826 , \4581 );
and \U$13393 ( \13580 , \3037 , \4424 );
nor \U$13394 ( \13581 , \13579 , \13580 );
xnor \U$13395 ( \13582 , \13581 , \4377 );
xor \U$13396 ( \13583 , \13578 , \13582 );
and \U$13397 ( \13584 , \2521 , \5011 );
and \U$13398 ( \13585 , \2757 , \4878 );
nor \U$13399 ( \13586 , \13584 , \13585 );
xnor \U$13400 ( \13587 , \13586 , \4762 );
xor \U$13401 ( \13588 , \13583 , \13587 );
and \U$13402 ( \13589 , \5674 , \2121 );
and \U$13403 ( \13590 , \6030 , \2008 );
nor \U$13404 ( \13591 , \13589 , \13590 );
xnor \U$13405 ( \13592 , \13591 , \1961 );
and \U$13406 ( \13593 , \5156 , \2400 );
and \U$13407 ( \13594 , \5469 , \2246 );
nor \U$13408 ( \13595 , \13593 , \13594 );
xnor \U$13409 ( \13596 , \13595 , \2195 );
xor \U$13410 ( \13597 , \13592 , \13596 );
and \U$13411 ( \13598 , \4749 , \2669 );
and \U$13412 ( \13599 , \4922 , \2538 );
nor \U$13413 ( \13600 , \13598 , \13599 );
xnor \U$13414 ( \13601 , \13600 , \2534 );
xor \U$13415 ( \13602 , \13597 , \13601 );
xor \U$13416 ( \13603 , \13588 , \13602 );
and \U$13417 ( \13604 , \4364 , \3103 );
and \U$13418 ( \13605 , \4654 , \2934 );
nor \U$13419 ( \13606 , \13604 , \13605 );
xnor \U$13420 ( \13607 , \13606 , \2839 );
and \U$13421 ( \13608 , \3912 , \3357 );
and \U$13422 ( \13609 , \4160 , \3255 );
nor \U$13423 ( \13610 , \13608 , \13609 );
xnor \U$13424 ( \13611 , \13610 , \3156 );
xor \U$13425 ( \13612 , \13607 , \13611 );
and \U$13426 ( \13613 , \3646 , \3813 );
and \U$13427 ( \13614 , \3736 , \3557 );
nor \U$13428 ( \13615 , \13613 , \13614 );
xnor \U$13429 ( \13616 , \13615 , \3562 );
xor \U$13430 ( \13617 , \13612 , \13616 );
xor \U$13431 ( \13618 , \13603 , \13617 );
xor \U$13432 ( \13619 , \13574 , \13618 );
and \U$13433 ( \13620 , \7231 , \1301 );
and \U$13434 ( \13621 , \7556 , \1246 );
nor \U$13435 ( \13622 , \13620 , \13621 );
xnor \U$13436 ( \13623 , \13622 , \1205 );
and \U$13437 ( \13624 , \6790 , \1578 );
and \U$13438 ( \13625 , \6945 , \1431 );
nor \U$13439 ( \13626 , \13624 , \13625 );
xnor \U$13440 ( \13627 , \13626 , \1436 );
xor \U$13441 ( \13628 , \13623 , \13627 );
and \U$13442 ( \13629 , \6281 , \1824 );
and \U$13443 ( \13630 , \6514 , \1739 );
nor \U$13444 ( \13631 , \13629 , \13630 );
xnor \U$13445 ( \13632 , \13631 , \1697 );
xor \U$13446 ( \13633 , \13628 , \13632 );
not \U$13447 ( \13634 , \252 );
and \U$13448 ( \13635 , \10206 , \141 );
and \U$13449 ( \13636 , \10584 , \139 );
nor \U$13450 ( \13637 , \13635 , \13636 );
xnor \U$13451 ( \13638 , \13637 , \148 );
xor \U$13452 ( \13639 , \13634 , \13638 );
and \U$13453 ( \13640 , \9465 , \156 );
and \U$13454 ( \13641 , \9897 , \154 );
nor \U$13455 ( \13642 , \13640 , \13641 );
xnor \U$13456 ( \13643 , \13642 , \163 );
xor \U$13457 ( \13644 , \13639 , \13643 );
xor \U$13458 ( \13645 , \13633 , \13644 );
and \U$13459 ( \13646 , \8835 , \296 );
and \U$13460 ( \13647 , \9169 , \168 );
nor \U$13461 ( \13648 , \13646 , \13647 );
xnor \U$13462 ( \13649 , \13648 , \173 );
and \U$13463 ( \13650 , \8349 , \438 );
and \U$13464 ( \13651 , \8652 , \336 );
nor \U$13465 ( \13652 , \13650 , \13651 );
xnor \U$13466 ( \13653 , \13652 , \320 );
xor \U$13467 ( \13654 , \13649 , \13653 );
and \U$13468 ( \13655 , \7700 , \1086 );
and \U$13469 ( \13656 , \8057 , \508 );
nor \U$13470 ( \13657 , \13655 , \13656 );
xnor \U$13471 ( \13658 , \13657 , \487 );
xor \U$13472 ( \13659 , \13654 , \13658 );
xor \U$13473 ( \13660 , \13645 , \13659 );
xor \U$13474 ( \13661 , \13619 , \13660 );
xor \U$13475 ( \13662 , \13530 , \13661 );
xor \U$13476 ( \13663 , \13501 , \13662 );
xor \U$13477 ( \13664 , \13428 , \13663 );
xor \U$13478 ( \13665 , \13419 , \13664 );
and \U$13479 ( \13666 , \13103 , \13378 );
xor \U$13480 ( \13667 , \13665 , \13666 );
and \U$13481 ( \13668 , \13379 , \13383 );
and \U$13482 ( \13669 , \13384 , \13387 );
or \U$13483 ( \13670 , \13668 , \13669 );
xor \U$13484 ( \13671 , \13667 , \13670 );
buf g5509_GF_PartitionCandidate( \13672_nG5509 , \13671 );
buf \U$13485 ( \13673 , \13672_nG5509 );
and \U$13486 ( \13674 , \13398 , \13402 );
and \U$13487 ( \13675 , \13402 , \13417 );
and \U$13488 ( \13676 , \13398 , \13417 );
or \U$13489 ( \13677 , \13674 , \13675 , \13676 );
and \U$13490 ( \13678 , \13423 , \13427 );
and \U$13491 ( \13679 , \13427 , \13663 );
and \U$13492 ( \13680 , \13423 , \13663 );
or \U$13493 ( \13681 , \13678 , \13679 , \13680 );
and \U$13494 ( \13682 , \13432 , \13436 );
and \U$13495 ( \13683 , \13436 , \13441 );
and \U$13496 ( \13684 , \13432 , \13441 );
or \U$13497 ( \13685 , \13682 , \13683 , \13684 );
and \U$13498 ( \13686 , \13446 , \13460 );
and \U$13499 ( \13687 , \13460 , \13499 );
and \U$13500 ( \13688 , \13446 , \13499 );
or \U$13501 ( \13689 , \13686 , \13687 , \13688 );
xor \U$13502 ( \13690 , \13685 , \13689 );
and \U$13503 ( \13691 , \13515 , \13529 );
and \U$13504 ( \13692 , \13529 , \13661 );
and \U$13505 ( \13693 , \13515 , \13661 );
or \U$13506 ( \13694 , \13691 , \13692 , \13693 );
xor \U$13507 ( \13695 , \13690 , \13694 );
xor \U$13508 ( \13696 , \13681 , \13695 );
and \U$13509 ( \13697 , \13407 , \13411 );
and \U$13510 ( \13698 , \13411 , \13416 );
and \U$13511 ( \13699 , \13407 , \13416 );
or \U$13512 ( \13700 , \13697 , \13698 , \13699 );
and \U$13513 ( \13701 , \13442 , \13500 );
and \U$13514 ( \13702 , \13500 , \13662 );
and \U$13515 ( \13703 , \13442 , \13662 );
or \U$13516 ( \13704 , \13701 , \13702 , \13703 );
xor \U$13517 ( \13705 , \13700 , \13704 );
and \U$13518 ( \13706 , \13505 , \13509 );
and \U$13519 ( \13707 , \13509 , \13514 );
and \U$13520 ( \13708 , \13505 , \13514 );
or \U$13521 ( \13709 , \13706 , \13707 , \13708 );
and \U$13522 ( \13710 , \13519 , \13523 );
and \U$13523 ( \13711 , \13523 , \13528 );
and \U$13524 ( \13712 , \13519 , \13528 );
or \U$13525 ( \13713 , \13710 , \13711 , \13712 );
xor \U$13526 ( \13714 , \13709 , \13713 );
and \U$13527 ( \13715 , \13574 , \13618 );
and \U$13528 ( \13716 , \13618 , \13660 );
and \U$13529 ( \13717 , \13574 , \13660 );
or \U$13530 ( \13718 , \13715 , \13716 , \13717 );
xor \U$13531 ( \13719 , \13714 , \13718 );
and \U$13532 ( \13720 , \13465 , \13469 );
and \U$13533 ( \13721 , \13469 , \13474 );
and \U$13534 ( \13722 , \13465 , \13474 );
or \U$13535 ( \13723 , \13720 , \13721 , \13722 );
and \U$13536 ( \13724 , \13479 , \13483 );
and \U$13537 ( \13725 , \13483 , \13488 );
and \U$13538 ( \13726 , \13479 , \13488 );
or \U$13539 ( \13727 , \13724 , \13725 , \13726 );
xor \U$13540 ( \13728 , \13723 , \13727 );
and \U$13541 ( \13729 , \13450 , \13454 );
and \U$13542 ( \13730 , \13454 , \13459 );
and \U$13543 ( \13731 , \13450 , \13459 );
or \U$13544 ( \13732 , \13729 , \13730 , \13731 );
xor \U$13545 ( \13733 , \13728 , \13732 );
and \U$13546 ( \13734 , \13491 , \13495 );
and \U$13547 ( \13735 , \13495 , \13497 );
and \U$13548 ( \13736 , \13491 , \13497 );
or \U$13549 ( \13737 , \13734 , \13735 , \13736 );
and \U$13550 ( \13738 , \13544 , \13558 );
and \U$13551 ( \13739 , \13558 , \13573 );
and \U$13552 ( \13740 , \13544 , \13573 );
or \U$13553 ( \13741 , \13738 , \13739 , \13740 );
xor \U$13554 ( \13742 , \13737 , \13741 );
and \U$13555 ( \13743 , \13588 , \13602 );
and \U$13556 ( \13744 , \13602 , \13617 );
and \U$13557 ( \13745 , \13588 , \13617 );
or \U$13558 ( \13746 , \13743 , \13744 , \13745 );
xor \U$13559 ( \13747 , \13742 , \13746 );
xor \U$13560 ( \13748 , \13733 , \13747 );
and \U$13561 ( \13749 , \13633 , \13644 );
and \U$13562 ( \13750 , \13644 , \13659 );
and \U$13563 ( \13751 , \13633 , \13659 );
or \U$13564 ( \13752 , \13749 , \13750 , \13751 );
and \U$13565 ( \13753 , \8652 , \438 );
and \U$13566 ( \13754 , \8835 , \336 );
nor \U$13567 ( \13755 , \13753 , \13754 );
xnor \U$13568 ( \13756 , \13755 , \320 );
and \U$13569 ( \13757 , \8057 , \1086 );
and \U$13570 ( \13758 , \8349 , \508 );
nor \U$13571 ( \13759 , \13757 , \13758 );
xnor \U$13572 ( \13760 , \13759 , \487 );
xor \U$13573 ( \13761 , \13756 , \13760 );
and \U$13574 ( \13762 , \7556 , \1301 );
and \U$13575 ( \13763 , \7700 , \1246 );
nor \U$13576 ( \13764 , \13762 , \13763 );
xnor \U$13577 ( \13765 , \13764 , \1205 );
xor \U$13578 ( \13766 , \13761 , \13765 );
xor \U$13579 ( \13767 , \13752 , \13766 );
and \U$13580 ( \13768 , \10584 , \141 );
not \U$13581 ( \13769 , \13768 );
xnor \U$13582 ( \13770 , \13769 , \148 );
and \U$13583 ( \13771 , \9897 , \156 );
and \U$13584 ( \13772 , \10206 , \154 );
nor \U$13585 ( \13773 , \13771 , \13772 );
xnor \U$13586 ( \13774 , \13773 , \163 );
xor \U$13587 ( \13775 , \13770 , \13774 );
and \U$13588 ( \13776 , \9169 , \296 );
and \U$13589 ( \13777 , \9465 , \168 );
nor \U$13590 ( \13778 , \13776 , \13777 );
xnor \U$13591 ( \13779 , \13778 , \173 );
xor \U$13592 ( \13780 , \13775 , \13779 );
xor \U$13593 ( \13781 , \13767 , \13780 );
xor \U$13594 ( \13782 , \13748 , \13781 );
xor \U$13595 ( \13783 , \13719 , \13782 );
and \U$13596 ( \13784 , \13475 , \13489 );
and \U$13597 ( \13785 , \13489 , \13498 );
and \U$13598 ( \13786 , \13475 , \13498 );
or \U$13599 ( \13787 , \13784 , \13785 , \13786 );
and \U$13600 ( \13788 , \13578 , \13582 );
and \U$13601 ( \13789 , \13582 , \13587 );
and \U$13602 ( \13790 , \13578 , \13587 );
or \U$13603 ( \13791 , \13788 , \13789 , \13790 );
and \U$13604 ( \13792 , \13592 , \13596 );
and \U$13605 ( \13793 , \13596 , \13601 );
and \U$13606 ( \13794 , \13592 , \13601 );
or \U$13607 ( \13795 , \13792 , \13793 , \13794 );
xor \U$13608 ( \13796 , \13791 , \13795 );
and \U$13609 ( \13797 , \13607 , \13611 );
and \U$13610 ( \13798 , \13611 , \13616 );
and \U$13611 ( \13799 , \13607 , \13616 );
or \U$13612 ( \13800 , \13797 , \13798 , \13799 );
xor \U$13613 ( \13801 , \13796 , \13800 );
and \U$13614 ( \13802 , \13623 , \13627 );
and \U$13615 ( \13803 , \13627 , \13632 );
and \U$13616 ( \13804 , \13623 , \13632 );
or \U$13617 ( \13805 , \13802 , \13803 , \13804 );
and \U$13618 ( \13806 , \13634 , \13638 );
and \U$13619 ( \13807 , \13638 , \13643 );
and \U$13620 ( \13808 , \13634 , \13643 );
or \U$13621 ( \13809 , \13806 , \13807 , \13808 );
xor \U$13622 ( \13810 , \13805 , \13809 );
and \U$13623 ( \13811 , \13649 , \13653 );
and \U$13624 ( \13812 , \13653 , \13658 );
and \U$13625 ( \13813 , \13649 , \13658 );
or \U$13626 ( \13814 , \13811 , \13812 , \13813 );
xor \U$13627 ( \13815 , \13810 , \13814 );
xor \U$13628 ( \13816 , \13801 , \13815 );
and \U$13629 ( \13817 , \13534 , \13538 );
and \U$13630 ( \13818 , \13538 , \13543 );
and \U$13631 ( \13819 , \13534 , \13543 );
or \U$13632 ( \13820 , \13817 , \13818 , \13819 );
and \U$13633 ( \13821 , \13548 , \13552 );
and \U$13634 ( \13822 , \13552 , \13557 );
and \U$13635 ( \13823 , \13548 , \13557 );
or \U$13636 ( \13824 , \13821 , \13822 , \13823 );
xor \U$13637 ( \13825 , \13820 , \13824 );
and \U$13638 ( \13826 , \13563 , \13567 );
and \U$13639 ( \13827 , \13567 , \13572 );
and \U$13640 ( \13828 , \13563 , \13572 );
or \U$13641 ( \13829 , \13826 , \13827 , \13828 );
xor \U$13642 ( \13830 , \13825 , \13829 );
xor \U$13643 ( \13831 , \13816 , \13830 );
xor \U$13644 ( \13832 , \13787 , \13831 );
and \U$13645 ( \13833 , \2090 , \5996 );
and \U$13646 ( \13834 , \2182 , \5695 );
nor \U$13647 ( \13835 , \13833 , \13834 );
xnor \U$13648 ( \13836 , \13835 , \5687 );
and \U$13649 ( \13837 , \1802 , \6401 );
and \U$13650 ( \13838 , \1948 , \6143 );
nor \U$13651 ( \13839 , \13837 , \13838 );
xnor \U$13652 ( \13840 , \13839 , \6148 );
xor \U$13653 ( \13841 , \13836 , \13840 );
and \U$13654 ( \13842 , \1601 , \7055 );
and \U$13655 ( \13843 , \1684 , \6675 );
nor \U$13656 ( \13844 , \13842 , \13843 );
xnor \U$13657 ( \13845 , \13844 , \6680 );
xor \U$13658 ( \13846 , \13841 , \13845 );
and \U$13659 ( \13847 , \3037 , \4581 );
and \U$13660 ( \13848 , \3143 , \4424 );
nor \U$13661 ( \13849 , \13847 , \13848 );
xnor \U$13662 ( \13850 , \13849 , \4377 );
and \U$13663 ( \13851 , \2757 , \5011 );
and \U$13664 ( \13852 , \2826 , \4878 );
nor \U$13665 ( \13853 , \13851 , \13852 );
xnor \U$13666 ( \13854 , \13853 , \4762 );
xor \U$13667 ( \13855 , \13850 , \13854 );
and \U$13668 ( \13856 , \2366 , \5485 );
and \U$13669 ( \13857 , \2521 , \5275 );
nor \U$13670 ( \13858 , \13856 , \13857 );
xnor \U$13671 ( \13859 , \13858 , \5169 );
xor \U$13672 ( \13860 , \13855 , \13859 );
xor \U$13673 ( \13861 , \13846 , \13860 );
and \U$13674 ( \13862 , \1333 , \7489 );
and \U$13675 ( \13863 , \1484 , \7137 );
nor \U$13676 ( \13864 , \13862 , \13863 );
xnor \U$13677 ( \13865 , \13864 , \7142 );
and \U$13678 ( \13866 , \1147 , \8019 );
and \U$13679 ( \13867 , \1192 , \7830 );
nor \U$13680 ( \13868 , \13866 , \13867 );
xnor \U$13681 ( \13869 , \13868 , \7713 );
xor \U$13682 ( \13870 , \13865 , \13869 );
and \U$13683 ( \13871 , \412 , \8540 );
and \U$13684 ( \13872 , \474 , \8292 );
nor \U$13685 ( \13873 , \13871 , \13872 );
xnor \U$13686 ( \13874 , \13873 , \8297 );
xor \U$13687 ( \13875 , \13870 , \13874 );
xor \U$13688 ( \13876 , \13861 , \13875 );
and \U$13689 ( \13877 , \6945 , \1578 );
and \U$13690 ( \13878 , \7231 , \1431 );
nor \U$13691 ( \13879 , \13877 , \13878 );
xnor \U$13692 ( \13880 , \13879 , \1436 );
and \U$13693 ( \13881 , \6514 , \1824 );
and \U$13694 ( \13882 , \6790 , \1739 );
nor \U$13695 ( \13883 , \13881 , \13882 );
xnor \U$13696 ( \13884 , \13883 , \1697 );
xor \U$13697 ( \13885 , \13880 , \13884 );
and \U$13698 ( \13886 , \6030 , \2121 );
and \U$13699 ( \13887 , \6281 , \2008 );
nor \U$13700 ( \13888 , \13886 , \13887 );
xnor \U$13701 ( \13889 , \13888 , \1961 );
xor \U$13702 ( \13890 , \13885 , \13889 );
and \U$13703 ( \13891 , \5469 , \2400 );
and \U$13704 ( \13892 , \5674 , \2246 );
nor \U$13705 ( \13893 , \13891 , \13892 );
xnor \U$13706 ( \13894 , \13893 , \2195 );
and \U$13707 ( \13895 , \4922 , \2669 );
and \U$13708 ( \13896 , \5156 , \2538 );
nor \U$13709 ( \13897 , \13895 , \13896 );
xnor \U$13710 ( \13898 , \13897 , \2534 );
xor \U$13711 ( \13899 , \13894 , \13898 );
and \U$13712 ( \13900 , \4654 , \3103 );
and \U$13713 ( \13901 , \4749 , \2934 );
nor \U$13714 ( \13902 , \13900 , \13901 );
xnor \U$13715 ( \13903 , \13902 , \2839 );
xor \U$13716 ( \13904 , \13899 , \13903 );
xor \U$13717 ( \13905 , \13890 , \13904 );
and \U$13718 ( \13906 , \4160 , \3357 );
and \U$13719 ( \13907 , \4364 , \3255 );
nor \U$13720 ( \13908 , \13906 , \13907 );
xnor \U$13721 ( \13909 , \13908 , \3156 );
and \U$13722 ( \13910 , \3736 , \3813 );
and \U$13723 ( \13911 , \3912 , \3557 );
nor \U$13724 ( \13912 , \13910 , \13911 );
xnor \U$13725 ( \13913 , \13912 , \3562 );
xor \U$13726 ( \13914 , \13909 , \13913 );
and \U$13727 ( \13915 , \3395 , \4132 );
and \U$13728 ( \13916 , \3646 , \4012 );
nor \U$13729 ( \13917 , \13915 , \13916 );
xnor \U$13730 ( \13918 , \13917 , \3925 );
xor \U$13731 ( \13919 , \13914 , \13918 );
xor \U$13732 ( \13920 , \13905 , \13919 );
xor \U$13733 ( \13921 , \13876 , \13920 );
and \U$13734 ( \13922 , \217 , \10118 );
and \U$13735 ( \13923 , \261 , \9333 );
and \U$13736 ( \13924 , \307 , \9006 );
nor \U$13737 ( \13925 , \13923 , \13924 );
xnor \U$13738 ( \13926 , \13925 , \8848 );
and \U$13739 ( \13927 , \178 , \9765 );
and \U$13740 ( \13928 , \185 , \9644 );
nor \U$13741 ( \13929 , \13927 , \13928 );
xnor \U$13742 ( \13930 , \13929 , \9478 );
xor \U$13743 ( \13931 , \13926 , \13930 );
and \U$13744 ( \13932 , \189 , \10408 );
and \U$13745 ( \13933 , \197 , \10116 );
nor \U$13746 ( \13934 , \13932 , \13933 );
xnor \U$13747 ( \13935 , \13934 , \10121 );
xor \U$13748 ( \13936 , \13931 , \13935 );
xnor \U$13749 ( \13937 , \13922 , \13936 );
xor \U$13750 ( \13938 , \13921 , \13937 );
xor \U$13751 ( \13939 , \13832 , \13938 );
xor \U$13752 ( \13940 , \13783 , \13939 );
xor \U$13753 ( \13941 , \13705 , \13940 );
xor \U$13754 ( \13942 , \13696 , \13941 );
xor \U$13755 ( \13943 , \13677 , \13942 );
and \U$13756 ( \13944 , \13394 , \13418 );
and \U$13757 ( \13945 , \13418 , \13664 );
and \U$13758 ( \13946 , \13394 , \13664 );
or \U$13759 ( \13947 , \13944 , \13945 , \13946 );
xor \U$13760 ( \13948 , \13943 , \13947 );
and \U$13761 ( \13949 , \13665 , \13666 );
and \U$13762 ( \13950 , \13667 , \13670 );
or \U$13763 ( \13951 , \13949 , \13950 );
xor \U$13764 ( \13952 , \13948 , \13951 );
buf g5507_GF_PartitionCandidate( \13953_nG5507 , \13952 );
buf \U$13765 ( \13954 , \13953_nG5507 );
and \U$13766 ( \13955 , \13681 , \13695 );
and \U$13767 ( \13956 , \13695 , \13941 );
and \U$13768 ( \13957 , \13681 , \13941 );
or \U$13769 ( \13958 , \13955 , \13956 , \13957 );
and \U$13770 ( \13959 , \13700 , \13704 );
and \U$13771 ( \13960 , \13704 , \13940 );
and \U$13772 ( \13961 , \13700 , \13940 );
or \U$13773 ( \13962 , \13959 , \13960 , \13961 );
and \U$13774 ( \13963 , \13685 , \13689 );
and \U$13775 ( \13964 , \13689 , \13694 );
and \U$13776 ( \13965 , \13685 , \13694 );
or \U$13777 ( \13966 , \13963 , \13964 , \13965 );
and \U$13778 ( \13967 , \13719 , \13782 );
and \U$13779 ( \13968 , \13782 , \13939 );
and \U$13780 ( \13969 , \13719 , \13939 );
or \U$13781 ( \13970 , \13967 , \13968 , \13969 );
xor \U$13782 ( \13971 , \13966 , \13970 );
and \U$13783 ( \13972 , \13723 , \13727 );
and \U$13784 ( \13973 , \13727 , \13732 );
and \U$13785 ( \13974 , \13723 , \13732 );
or \U$13786 ( \13975 , \13972 , \13973 , \13974 );
and \U$13787 ( \13976 , \13737 , \13741 );
and \U$13788 ( \13977 , \13741 , \13746 );
and \U$13789 ( \13978 , \13737 , \13746 );
or \U$13790 ( \13979 , \13976 , \13977 , \13978 );
xor \U$13791 ( \13980 , \13975 , \13979 );
and \U$13792 ( \13981 , \13752 , \13766 );
and \U$13793 ( \13982 , \13766 , \13780 );
and \U$13794 ( \13983 , \13752 , \13780 );
or \U$13795 ( \13984 , \13981 , \13982 , \13983 );
xor \U$13796 ( \13985 , \13980 , \13984 );
xor \U$13797 ( \13986 , \13971 , \13985 );
xor \U$13798 ( \13987 , \13962 , \13986 );
and \U$13799 ( \13988 , \13709 , \13713 );
and \U$13800 ( \13989 , \13713 , \13718 );
and \U$13801 ( \13990 , \13709 , \13718 );
or \U$13802 ( \13991 , \13988 , \13989 , \13990 );
and \U$13803 ( \13992 , \13733 , \13747 );
and \U$13804 ( \13993 , \13747 , \13781 );
and \U$13805 ( \13994 , \13733 , \13781 );
or \U$13806 ( \13995 , \13992 , \13993 , \13994 );
xor \U$13807 ( \13996 , \13991 , \13995 );
and \U$13808 ( \13997 , \13787 , \13831 );
and \U$13809 ( \13998 , \13831 , \13938 );
and \U$13810 ( \13999 , \13787 , \13938 );
or \U$13811 ( \14000 , \13997 , \13998 , \13999 );
xor \U$13812 ( \14001 , \13996 , \14000 );
and \U$13813 ( \14002 , \13791 , \13795 );
and \U$13814 ( \14003 , \13795 , \13800 );
and \U$13815 ( \14004 , \13791 , \13800 );
or \U$13816 ( \14005 , \14002 , \14003 , \14004 );
and \U$13817 ( \14006 , \13805 , \13809 );
and \U$13818 ( \14007 , \13809 , \13814 );
and \U$13819 ( \14008 , \13805 , \13814 );
or \U$13820 ( \14009 , \14006 , \14007 , \14008 );
xor \U$13821 ( \14010 , \14005 , \14009 );
and \U$13822 ( \14011 , \13820 , \13824 );
and \U$13823 ( \14012 , \13824 , \13829 );
and \U$13824 ( \14013 , \13820 , \13829 );
or \U$13825 ( \14014 , \14011 , \14012 , \14013 );
xor \U$13826 ( \14015 , \14010 , \14014 );
and \U$13827 ( \14016 , \13801 , \13815 );
and \U$13828 ( \14017 , \13815 , \13830 );
and \U$13829 ( \14018 , \13801 , \13830 );
or \U$13830 ( \14019 , \14016 , \14017 , \14018 );
and \U$13831 ( \14020 , \13876 , \13920 );
and \U$13832 ( \14021 , \13920 , \13937 );
and \U$13833 ( \14022 , \13876 , \13937 );
or \U$13834 ( \14023 , \14020 , \14021 , \14022 );
xor \U$13835 ( \14024 , \14019 , \14023 );
and \U$13836 ( \14025 , \13756 , \13760 );
and \U$13837 ( \14026 , \13760 , \13765 );
and \U$13838 ( \14027 , \13756 , \13765 );
or \U$13839 ( \14028 , \14025 , \14026 , \14027 );
and \U$13840 ( \14029 , \13880 , \13884 );
and \U$13841 ( \14030 , \13884 , \13889 );
and \U$13842 ( \14031 , \13880 , \13889 );
or \U$13843 ( \14032 , \14029 , \14030 , \14031 );
xor \U$13844 ( \14033 , \14028 , \14032 );
and \U$13845 ( \14034 , \13770 , \13774 );
and \U$13846 ( \14035 , \13774 , \13779 );
and \U$13847 ( \14036 , \13770 , \13779 );
or \U$13848 ( \14037 , \14034 , \14035 , \14036 );
xor \U$13849 ( \14038 , \14033 , \14037 );
xor \U$13850 ( \14039 , \14024 , \14038 );
xor \U$13851 ( \14040 , \14015 , \14039 );
and \U$13852 ( \14041 , \13846 , \13860 );
and \U$13853 ( \14042 , \13860 , \13875 );
and \U$13854 ( \14043 , \13846 , \13875 );
or \U$13855 ( \14044 , \14041 , \14042 , \14043 );
and \U$13856 ( \14045 , \13890 , \13904 );
and \U$13857 ( \14046 , \13904 , \13919 );
and \U$13858 ( \14047 , \13890 , \13919 );
or \U$13859 ( \14048 , \14045 , \14046 , \14047 );
xor \U$13860 ( \14049 , \14044 , \14048 );
or \U$13861 ( \14050 , \13922 , \13936 );
xor \U$13862 ( \14051 , \14049 , \14050 );
and \U$13863 ( \14052 , \13836 , \13840 );
and \U$13864 ( \14053 , \13840 , \13845 );
and \U$13865 ( \14054 , \13836 , \13845 );
or \U$13866 ( \14055 , \14052 , \14053 , \14054 );
and \U$13867 ( \14056 , \13926 , \13930 );
and \U$13868 ( \14057 , \13930 , \13935 );
and \U$13869 ( \14058 , \13926 , \13935 );
or \U$13870 ( \14059 , \14056 , \14057 , \14058 );
xor \U$13871 ( \14060 , \14055 , \14059 );
and \U$13872 ( \14061 , \13865 , \13869 );
and \U$13873 ( \14062 , \13869 , \13874 );
and \U$13874 ( \14063 , \13865 , \13874 );
or \U$13875 ( \14064 , \14061 , \14062 , \14063 );
xor \U$13876 ( \14065 , \14060 , \14064 );
and \U$13877 ( \14066 , \13850 , \13854 );
and \U$13878 ( \14067 , \13854 , \13859 );
and \U$13879 ( \14068 , \13850 , \13859 );
or \U$13880 ( \14069 , \14066 , \14067 , \14068 );
and \U$13881 ( \14070 , \13894 , \13898 );
and \U$13882 ( \14071 , \13898 , \13903 );
and \U$13883 ( \14072 , \13894 , \13903 );
or \U$13884 ( \14073 , \14070 , \14071 , \14072 );
xor \U$13885 ( \14074 , \14069 , \14073 );
and \U$13886 ( \14075 , \13909 , \13913 );
and \U$13887 ( \14076 , \13913 , \13918 );
and \U$13888 ( \14077 , \13909 , \13918 );
or \U$13889 ( \14078 , \14075 , \14076 , \14077 );
xor \U$13890 ( \14079 , \14074 , \14078 );
xor \U$13891 ( \14080 , \14065 , \14079 );
and \U$13892 ( \14081 , \189 , \10118 );
and \U$13893 ( \14082 , \1484 , \7489 );
and \U$13894 ( \14083 , \1601 , \7137 );
nor \U$13895 ( \14084 , \14082 , \14083 );
xnor \U$13896 ( \14085 , \14084 , \7142 );
and \U$13897 ( \14086 , \1192 , \8019 );
and \U$13898 ( \14087 , \1333 , \7830 );
nor \U$13899 ( \14088 , \14086 , \14087 );
xnor \U$13900 ( \14089 , \14088 , \7713 );
xor \U$13901 ( \14090 , \14085 , \14089 );
and \U$13902 ( \14091 , \474 , \8540 );
and \U$13903 ( \14092 , \1147 , \8292 );
nor \U$13904 ( \14093 , \14091 , \14092 );
xnor \U$13905 ( \14094 , \14093 , \8297 );
xor \U$13906 ( \14095 , \14090 , \14094 );
xor \U$13907 ( \14096 , \14081 , \14095 );
and \U$13908 ( \14097 , \307 , \9333 );
and \U$13909 ( \14098 , \412 , \9006 );
nor \U$13910 ( \14099 , \14097 , \14098 );
xnor \U$13911 ( \14100 , \14099 , \8848 );
and \U$13912 ( \14101 , \185 , \9765 );
and \U$13913 ( \14102 , \261 , \9644 );
nor \U$13914 ( \14103 , \14101 , \14102 );
xnor \U$13915 ( \14104 , \14103 , \9478 );
xor \U$13916 ( \14105 , \14100 , \14104 );
and \U$13917 ( \14106 , \197 , \10408 );
and \U$13918 ( \14107 , \178 , \10116 );
nor \U$13919 ( \14108 , \14106 , \14107 );
xnor \U$13920 ( \14109 , \14108 , \10121 );
xor \U$13921 ( \14110 , \14105 , \14109 );
xor \U$13922 ( \14111 , \14096 , \14110 );
xor \U$13923 ( \14112 , \14080 , \14111 );
xor \U$13924 ( \14113 , \14051 , \14112 );
not \U$13925 ( \14114 , \148 );
and \U$13926 ( \14115 , \10206 , \156 );
and \U$13927 ( \14116 , \10584 , \154 );
nor \U$13928 ( \14117 , \14115 , \14116 );
xnor \U$13929 ( \14118 , \14117 , \163 );
xor \U$13930 ( \14119 , \14114 , \14118 );
and \U$13931 ( \14120 , \9465 , \296 );
and \U$13932 ( \14121 , \9897 , \168 );
nor \U$13933 ( \14122 , \14120 , \14121 );
xnor \U$13934 ( \14123 , \14122 , \173 );
xor \U$13935 ( \14124 , \14119 , \14123 );
and \U$13936 ( \14125 , \8835 , \438 );
and \U$13937 ( \14126 , \9169 , \336 );
nor \U$13938 ( \14127 , \14125 , \14126 );
xnor \U$13939 ( \14128 , \14127 , \320 );
and \U$13940 ( \14129 , \8349 , \1086 );
and \U$13941 ( \14130 , \8652 , \508 );
nor \U$13942 ( \14131 , \14129 , \14130 );
xnor \U$13943 ( \14132 , \14131 , \487 );
xor \U$13944 ( \14133 , \14128 , \14132 );
and \U$13945 ( \14134 , \7700 , \1301 );
and \U$13946 ( \14135 , \8057 , \1246 );
nor \U$13947 ( \14136 , \14134 , \14135 );
xnor \U$13948 ( \14137 , \14136 , \1205 );
xor \U$13949 ( \14138 , \14133 , \14137 );
and \U$13950 ( \14139 , \5674 , \2400 );
and \U$13951 ( \14140 , \6030 , \2246 );
nor \U$13952 ( \14141 , \14139 , \14140 );
xnor \U$13953 ( \14142 , \14141 , \2195 );
and \U$13954 ( \14143 , \5156 , \2669 );
and \U$13955 ( \14144 , \5469 , \2538 );
nor \U$13956 ( \14145 , \14143 , \14144 );
xnor \U$13957 ( \14146 , \14145 , \2534 );
xor \U$13958 ( \14147 , \14142 , \14146 );
and \U$13959 ( \14148 , \4749 , \3103 );
and \U$13960 ( \14149 , \4922 , \2934 );
nor \U$13961 ( \14150 , \14148 , \14149 );
xnor \U$13962 ( \14151 , \14150 , \2839 );
xor \U$13963 ( \14152 , \14147 , \14151 );
xor \U$13964 ( \14153 , \14138 , \14152 );
and \U$13965 ( \14154 , \7231 , \1578 );
and \U$13966 ( \14155 , \7556 , \1431 );
nor \U$13967 ( \14156 , \14154 , \14155 );
xnor \U$13968 ( \14157 , \14156 , \1436 );
and \U$13969 ( \14158 , \6790 , \1824 );
and \U$13970 ( \14159 , \6945 , \1739 );
nor \U$13971 ( \14160 , \14158 , \14159 );
xnor \U$13972 ( \14161 , \14160 , \1697 );
xor \U$13973 ( \14162 , \14157 , \14161 );
and \U$13974 ( \14163 , \6281 , \2121 );
and \U$13975 ( \14164 , \6514 , \2008 );
nor \U$13976 ( \14165 , \14163 , \14164 );
xnor \U$13977 ( \14166 , \14165 , \1961 );
xor \U$13978 ( \14167 , \14162 , \14166 );
xor \U$13979 ( \14168 , \14153 , \14167 );
xor \U$13980 ( \14169 , \14124 , \14168 );
and \U$13981 ( \14170 , \2182 , \5996 );
and \U$13982 ( \14171 , \2366 , \5695 );
nor \U$13983 ( \14172 , \14170 , \14171 );
xnor \U$13984 ( \14173 , \14172 , \5687 );
and \U$13985 ( \14174 , \1948 , \6401 );
and \U$13986 ( \14175 , \2090 , \6143 );
nor \U$13987 ( \14176 , \14174 , \14175 );
xnor \U$13988 ( \14177 , \14176 , \6148 );
xor \U$13989 ( \14178 , \14173 , \14177 );
and \U$13990 ( \14179 , \1684 , \7055 );
and \U$13991 ( \14180 , \1802 , \6675 );
nor \U$13992 ( \14181 , \14179 , \14180 );
xnor \U$13993 ( \14182 , \14181 , \6680 );
xor \U$13994 ( \14183 , \14178 , \14182 );
and \U$13995 ( \14184 , \4364 , \3357 );
and \U$13996 ( \14185 , \4654 , \3255 );
nor \U$13997 ( \14186 , \14184 , \14185 );
xnor \U$13998 ( \14187 , \14186 , \3156 );
and \U$13999 ( \14188 , \3912 , \3813 );
and \U$14000 ( \14189 , \4160 , \3557 );
nor \U$14001 ( \14190 , \14188 , \14189 );
xnor \U$14002 ( \14191 , \14190 , \3562 );
xor \U$14003 ( \14192 , \14187 , \14191 );
and \U$14004 ( \14193 , \3646 , \4132 );
and \U$14005 ( \14194 , \3736 , \4012 );
nor \U$14006 ( \14195 , \14193 , \14194 );
xnor \U$14007 ( \14196 , \14195 , \3925 );
xor \U$14008 ( \14197 , \14192 , \14196 );
xor \U$14009 ( \14198 , \14183 , \14197 );
and \U$14010 ( \14199 , \3143 , \4581 );
and \U$14011 ( \14200 , \3395 , \4424 );
nor \U$14012 ( \14201 , \14199 , \14200 );
xnor \U$14013 ( \14202 , \14201 , \4377 );
and \U$14014 ( \14203 , \2826 , \5011 );
and \U$14015 ( \14204 , \3037 , \4878 );
nor \U$14016 ( \14205 , \14203 , \14204 );
xnor \U$14017 ( \14206 , \14205 , \4762 );
xor \U$14018 ( \14207 , \14202 , \14206 );
and \U$14019 ( \14208 , \2521 , \5485 );
and \U$14020 ( \14209 , \2757 , \5275 );
nor \U$14021 ( \14210 , \14208 , \14209 );
xnor \U$14022 ( \14211 , \14210 , \5169 );
xor \U$14023 ( \14212 , \14207 , \14211 );
xor \U$14024 ( \14213 , \14198 , \14212 );
xor \U$14025 ( \14214 , \14169 , \14213 );
xor \U$14026 ( \14215 , \14113 , \14214 );
xor \U$14027 ( \14216 , \14040 , \14215 );
xor \U$14028 ( \14217 , \14001 , \14216 );
xor \U$14029 ( \14218 , \13987 , \14217 );
xor \U$14030 ( \14219 , \13958 , \14218 );
and \U$14031 ( \14220 , \13677 , \13942 );
xor \U$14032 ( \14221 , \14219 , \14220 );
and \U$14033 ( \14222 , \13943 , \13947 );
and \U$14034 ( \14223 , \13948 , \13951 );
or \U$14035 ( \14224 , \14222 , \14223 );
xor \U$14036 ( \14225 , \14221 , \14224 );
buf g5505_GF_PartitionCandidate( \14226_nG5505 , \14225 );
buf \U$14037 ( \14227 , \14226_nG5505 );
and \U$14038 ( \14228 , \13962 , \13986 );
and \U$14039 ( \14229 , \13986 , \14217 );
and \U$14040 ( \14230 , \13962 , \14217 );
or \U$14041 ( \14231 , \14228 , \14229 , \14230 );
and \U$14042 ( \14232 , \13966 , \13970 );
and \U$14043 ( \14233 , \13970 , \13985 );
and \U$14044 ( \14234 , \13966 , \13985 );
or \U$14045 ( \14235 , \14232 , \14233 , \14234 );
and \U$14046 ( \14236 , \14001 , \14216 );
xor \U$14047 ( \14237 , \14235 , \14236 );
and \U$14048 ( \14238 , \13975 , \13979 );
and \U$14049 ( \14239 , \13979 , \13984 );
and \U$14050 ( \14240 , \13975 , \13984 );
or \U$14051 ( \14241 , \14238 , \14239 , \14240 );
and \U$14052 ( \14242 , \14019 , \14023 );
and \U$14053 ( \14243 , \14023 , \14038 );
and \U$14054 ( \14244 , \14019 , \14038 );
or \U$14055 ( \14245 , \14242 , \14243 , \14244 );
xor \U$14056 ( \14246 , \14241 , \14245 );
and \U$14057 ( \14247 , \14051 , \14112 );
and \U$14058 ( \14248 , \14112 , \14214 );
and \U$14059 ( \14249 , \14051 , \14214 );
or \U$14060 ( \14250 , \14247 , \14248 , \14249 );
xor \U$14061 ( \14251 , \14246 , \14250 );
xor \U$14062 ( \14252 , \14237 , \14251 );
xor \U$14063 ( \14253 , \14231 , \14252 );
and \U$14064 ( \14254 , \13991 , \13995 );
and \U$14065 ( \14255 , \13995 , \14000 );
and \U$14066 ( \14256 , \13991 , \14000 );
or \U$14067 ( \14257 , \14254 , \14255 , \14256 );
and \U$14068 ( \14258 , \14015 , \14039 );
and \U$14069 ( \14259 , \14039 , \14215 );
and \U$14070 ( \14260 , \14015 , \14215 );
or \U$14071 ( \14261 , \14258 , \14259 , \14260 );
xor \U$14072 ( \14262 , \14257 , \14261 );
and \U$14073 ( \14263 , \14005 , \14009 );
and \U$14074 ( \14264 , \14009 , \14014 );
and \U$14075 ( \14265 , \14005 , \14014 );
or \U$14076 ( \14266 , \14263 , \14264 , \14265 );
and \U$14077 ( \14267 , \14044 , \14048 );
and \U$14078 ( \14268 , \14048 , \14050 );
and \U$14079 ( \14269 , \14044 , \14050 );
or \U$14080 ( \14270 , \14267 , \14268 , \14269 );
xor \U$14081 ( \14271 , \14266 , \14270 );
and \U$14082 ( \14272 , \14124 , \14168 );
and \U$14083 ( \14273 , \14168 , \14213 );
and \U$14084 ( \14274 , \14124 , \14213 );
or \U$14085 ( \14275 , \14272 , \14273 , \14274 );
xor \U$14086 ( \14276 , \14271 , \14275 );
and \U$14087 ( \14277 , \14055 , \14059 );
and \U$14088 ( \14278 , \14059 , \14064 );
and \U$14089 ( \14279 , \14055 , \14064 );
or \U$14090 ( \14280 , \14277 , \14278 , \14279 );
and \U$14091 ( \14281 , \14028 , \14032 );
and \U$14092 ( \14282 , \14032 , \14037 );
and \U$14093 ( \14283 , \14028 , \14037 );
or \U$14094 ( \14284 , \14281 , \14282 , \14283 );
xor \U$14095 ( \14285 , \14280 , \14284 );
and \U$14096 ( \14286 , \14069 , \14073 );
and \U$14097 ( \14287 , \14073 , \14078 );
and \U$14098 ( \14288 , \14069 , \14078 );
or \U$14099 ( \14289 , \14286 , \14287 , \14288 );
xor \U$14100 ( \14290 , \14285 , \14289 );
and \U$14101 ( \14291 , \14138 , \14152 );
and \U$14102 ( \14292 , \14152 , \14167 );
and \U$14103 ( \14293 , \14138 , \14167 );
or \U$14104 ( \14294 , \14291 , \14292 , \14293 );
and \U$14105 ( \14295 , \14081 , \14095 );
and \U$14106 ( \14296 , \14095 , \14110 );
and \U$14107 ( \14297 , \14081 , \14110 );
or \U$14108 ( \14298 , \14295 , \14296 , \14297 );
xor \U$14109 ( \14299 , \14294 , \14298 );
and \U$14110 ( \14300 , \14183 , \14197 );
and \U$14111 ( \14301 , \14197 , \14212 );
and \U$14112 ( \14302 , \14183 , \14212 );
or \U$14113 ( \14303 , \14300 , \14301 , \14302 );
xor \U$14114 ( \14304 , \14299 , \14303 );
xor \U$14115 ( \14305 , \14290 , \14304 );
and \U$14116 ( \14306 , \10584 , \156 );
not \U$14117 ( \14307 , \14306 );
xnor \U$14118 ( \14308 , \14307 , \163 );
and \U$14119 ( \14309 , \9897 , \296 );
and \U$14120 ( \14310 , \10206 , \168 );
nor \U$14121 ( \14311 , \14309 , \14310 );
xnor \U$14122 ( \14312 , \14311 , \173 );
xor \U$14123 ( \14313 , \14308 , \14312 );
and \U$14124 ( \14314 , \9169 , \438 );
and \U$14125 ( \14315 , \9465 , \336 );
nor \U$14126 ( \14316 , \14314 , \14315 );
xnor \U$14127 ( \14317 , \14316 , \320 );
xor \U$14128 ( \14318 , \14313 , \14317 );
and \U$14129 ( \14319 , \8652 , \1086 );
and \U$14130 ( \14320 , \8835 , \508 );
nor \U$14131 ( \14321 , \14319 , \14320 );
xnor \U$14132 ( \14322 , \14321 , \487 );
and \U$14133 ( \14323 , \8057 , \1301 );
and \U$14134 ( \14324 , \8349 , \1246 );
nor \U$14135 ( \14325 , \14323 , \14324 );
xnor \U$14136 ( \14326 , \14325 , \1205 );
xor \U$14137 ( \14327 , \14322 , \14326 );
and \U$14138 ( \14328 , \7556 , \1578 );
and \U$14139 ( \14329 , \7700 , \1431 );
nor \U$14140 ( \14330 , \14328 , \14329 );
xnor \U$14141 ( \14331 , \14330 , \1436 );
xor \U$14142 ( \14332 , \14327 , \14331 );
and \U$14143 ( \14333 , \5469 , \2669 );
and \U$14144 ( \14334 , \5674 , \2538 );
nor \U$14145 ( \14335 , \14333 , \14334 );
xnor \U$14146 ( \14336 , \14335 , \2534 );
and \U$14147 ( \14337 , \4922 , \3103 );
and \U$14148 ( \14338 , \5156 , \2934 );
nor \U$14149 ( \14339 , \14337 , \14338 );
xnor \U$14150 ( \14340 , \14339 , \2839 );
xor \U$14151 ( \14341 , \14336 , \14340 );
and \U$14152 ( \14342 , \4654 , \3357 );
and \U$14153 ( \14343 , \4749 , \3255 );
nor \U$14154 ( \14344 , \14342 , \14343 );
xnor \U$14155 ( \14345 , \14344 , \3156 );
xor \U$14156 ( \14346 , \14341 , \14345 );
xor \U$14157 ( \14347 , \14332 , \14346 );
and \U$14158 ( \14348 , \6945 , \1824 );
and \U$14159 ( \14349 , \7231 , \1739 );
nor \U$14160 ( \14350 , \14348 , \14349 );
xnor \U$14161 ( \14351 , \14350 , \1697 );
and \U$14162 ( \14352 , \6514 , \2121 );
and \U$14163 ( \14353 , \6790 , \2008 );
nor \U$14164 ( \14354 , \14352 , \14353 );
xnor \U$14165 ( \14355 , \14354 , \1961 );
xor \U$14166 ( \14356 , \14351 , \14355 );
and \U$14167 ( \14357 , \6030 , \2400 );
and \U$14168 ( \14358 , \6281 , \2246 );
nor \U$14169 ( \14359 , \14357 , \14358 );
xnor \U$14170 ( \14360 , \14359 , \2195 );
xor \U$14171 ( \14361 , \14356 , \14360 );
xor \U$14172 ( \14362 , \14347 , \14361 );
xor \U$14173 ( \14363 , \14318 , \14362 );
and \U$14174 ( \14364 , \4160 , \3813 );
and \U$14175 ( \14365 , \4364 , \3557 );
nor \U$14176 ( \14366 , \14364 , \14365 );
xnor \U$14177 ( \14367 , \14366 , \3562 );
and \U$14178 ( \14368 , \3736 , \4132 );
and \U$14179 ( \14369 , \3912 , \4012 );
nor \U$14180 ( \14370 , \14368 , \14369 );
xnor \U$14181 ( \14371 , \14370 , \3925 );
xor \U$14182 ( \14372 , \14367 , \14371 );
and \U$14183 ( \14373 , \3395 , \4581 );
and \U$14184 ( \14374 , \3646 , \4424 );
nor \U$14185 ( \14375 , \14373 , \14374 );
xnor \U$14186 ( \14376 , \14375 , \4377 );
xor \U$14187 ( \14377 , \14372 , \14376 );
and \U$14188 ( \14378 , \2090 , \6401 );
and \U$14189 ( \14379 , \2182 , \6143 );
nor \U$14190 ( \14380 , \14378 , \14379 );
xnor \U$14191 ( \14381 , \14380 , \6148 );
and \U$14192 ( \14382 , \1802 , \7055 );
and \U$14193 ( \14383 , \1948 , \6675 );
nor \U$14194 ( \14384 , \14382 , \14383 );
xnor \U$14195 ( \14385 , \14384 , \6680 );
xor \U$14196 ( \14386 , \14381 , \14385 );
and \U$14197 ( \14387 , \1601 , \7489 );
and \U$14198 ( \14388 , \1684 , \7137 );
nor \U$14199 ( \14389 , \14387 , \14388 );
xnor \U$14200 ( \14390 , \14389 , \7142 );
xor \U$14201 ( \14391 , \14386 , \14390 );
xor \U$14202 ( \14392 , \14377 , \14391 );
and \U$14203 ( \14393 , \3037 , \5011 );
and \U$14204 ( \14394 , \3143 , \4878 );
nor \U$14205 ( \14395 , \14393 , \14394 );
xnor \U$14206 ( \14396 , \14395 , \4762 );
and \U$14207 ( \14397 , \2757 , \5485 );
and \U$14208 ( \14398 , \2826 , \5275 );
nor \U$14209 ( \14399 , \14397 , \14398 );
xnor \U$14210 ( \14400 , \14399 , \5169 );
xor \U$14211 ( \14401 , \14396 , \14400 );
and \U$14212 ( \14402 , \2366 , \5996 );
and \U$14213 ( \14403 , \2521 , \5695 );
nor \U$14214 ( \14404 , \14402 , \14403 );
xnor \U$14215 ( \14405 , \14404 , \5687 );
xor \U$14216 ( \14406 , \14401 , \14405 );
xor \U$14217 ( \14407 , \14392 , \14406 );
xor \U$14218 ( \14408 , \14363 , \14407 );
xor \U$14219 ( \14409 , \14305 , \14408 );
xor \U$14220 ( \14410 , \14276 , \14409 );
and \U$14221 ( \14411 , \14065 , \14079 );
and \U$14222 ( \14412 , \14079 , \14111 );
and \U$14223 ( \14413 , \14065 , \14111 );
or \U$14224 ( \14414 , \14411 , \14412 , \14413 );
and \U$14225 ( \14415 , \14128 , \14132 );
and \U$14226 ( \14416 , \14132 , \14137 );
and \U$14227 ( \14417 , \14128 , \14137 );
or \U$14228 ( \14418 , \14415 , \14416 , \14417 );
and \U$14229 ( \14419 , \14114 , \14118 );
and \U$14230 ( \14420 , \14118 , \14123 );
and \U$14231 ( \14421 , \14114 , \14123 );
or \U$14232 ( \14422 , \14419 , \14420 , \14421 );
xor \U$14233 ( \14423 , \14418 , \14422 );
and \U$14234 ( \14424 , \14157 , \14161 );
and \U$14235 ( \14425 , \14161 , \14166 );
and \U$14236 ( \14426 , \14157 , \14166 );
or \U$14237 ( \14427 , \14424 , \14425 , \14426 );
xor \U$14238 ( \14428 , \14423 , \14427 );
xor \U$14239 ( \14429 , \14414 , \14428 );
and \U$14240 ( \14430 , \14187 , \14191 );
and \U$14241 ( \14431 , \14191 , \14196 );
and \U$14242 ( \14432 , \14187 , \14196 );
or \U$14243 ( \14433 , \14430 , \14431 , \14432 );
and \U$14244 ( \14434 , \14142 , \14146 );
and \U$14245 ( \14435 , \14146 , \14151 );
and \U$14246 ( \14436 , \14142 , \14151 );
or \U$14247 ( \14437 , \14434 , \14435 , \14436 );
xor \U$14248 ( \14438 , \14433 , \14437 );
and \U$14249 ( \14439 , \14202 , \14206 );
and \U$14250 ( \14440 , \14206 , \14211 );
and \U$14251 ( \14441 , \14202 , \14211 );
or \U$14252 ( \14442 , \14439 , \14440 , \14441 );
xor \U$14253 ( \14443 , \14438 , \14442 );
and \U$14254 ( \14444 , \14173 , \14177 );
and \U$14255 ( \14445 , \14177 , \14182 );
and \U$14256 ( \14446 , \14173 , \14182 );
or \U$14257 ( \14447 , \14444 , \14445 , \14446 );
and \U$14258 ( \14448 , \14085 , \14089 );
and \U$14259 ( \14449 , \14089 , \14094 );
and \U$14260 ( \14450 , \14085 , \14094 );
or \U$14261 ( \14451 , \14448 , \14449 , \14450 );
xor \U$14262 ( \14452 , \14447 , \14451 );
and \U$14263 ( \14453 , \14100 , \14104 );
and \U$14264 ( \14454 , \14104 , \14109 );
and \U$14265 ( \14455 , \14100 , \14109 );
or \U$14266 ( \14456 , \14453 , \14454 , \14455 );
xor \U$14267 ( \14457 , \14452 , \14456 );
xor \U$14268 ( \14458 , \14443 , \14457 );
and \U$14269 ( \14459 , \261 , \9765 );
and \U$14270 ( \14460 , \307 , \9644 );
nor \U$14271 ( \14461 , \14459 , \14460 );
xnor \U$14272 ( \14462 , \14461 , \9478 );
and \U$14273 ( \14463 , \178 , \10408 );
and \U$14274 ( \14464 , \185 , \10116 );
nor \U$14275 ( \14465 , \14463 , \14464 );
xnor \U$14276 ( \14466 , \14465 , \10121 );
xor \U$14277 ( \14467 , \14462 , \14466 );
and \U$14278 ( \14468 , \197 , \10118 );
xor \U$14279 ( \14469 , \14467 , \14468 );
and \U$14280 ( \14470 , \1333 , \8019 );
and \U$14281 ( \14471 , \1484 , \7830 );
nor \U$14282 ( \14472 , \14470 , \14471 );
xnor \U$14283 ( \14473 , \14472 , \7713 );
and \U$14284 ( \14474 , \1147 , \8540 );
and \U$14285 ( \14475 , \1192 , \8292 );
nor \U$14286 ( \14476 , \14474 , \14475 );
xnor \U$14287 ( \14477 , \14476 , \8297 );
xor \U$14288 ( \14478 , \14473 , \14477 );
and \U$14289 ( \14479 , \412 , \9333 );
and \U$14290 ( \14480 , \474 , \9006 );
nor \U$14291 ( \14481 , \14479 , \14480 );
xnor \U$14292 ( \14482 , \14481 , \8848 );
xor \U$14293 ( \14483 , \14478 , \14482 );
xnor \U$14294 ( \14484 , \14469 , \14483 );
xor \U$14295 ( \14485 , \14458 , \14484 );
xor \U$14296 ( \14486 , \14429 , \14485 );
xor \U$14297 ( \14487 , \14410 , \14486 );
xor \U$14298 ( \14488 , \14262 , \14487 );
xor \U$14299 ( \14489 , \14253 , \14488 );
and \U$14300 ( \14490 , \13958 , \14218 );
xor \U$14301 ( \14491 , \14489 , \14490 );
and \U$14302 ( \14492 , \14219 , \14220 );
and \U$14303 ( \14493 , \14221 , \14224 );
or \U$14304 ( \14494 , \14492 , \14493 );
xor \U$14305 ( \14495 , \14491 , \14494 );
buf g5503_GF_PartitionCandidate( \14496_nG5503 , \14495 );
buf \U$14306 ( \14497 , \14496_nG5503 );
and \U$14307 ( \14498 , \14235 , \14236 );
and \U$14308 ( \14499 , \14236 , \14251 );
and \U$14309 ( \14500 , \14235 , \14251 );
or \U$14310 ( \14501 , \14498 , \14499 , \14500 );
and \U$14311 ( \14502 , \14257 , \14261 );
and \U$14312 ( \14503 , \14261 , \14487 );
and \U$14313 ( \14504 , \14257 , \14487 );
or \U$14314 ( \14505 , \14502 , \14503 , \14504 );
and \U$14315 ( \14506 , \14266 , \14270 );
and \U$14316 ( \14507 , \14270 , \14275 );
and \U$14317 ( \14508 , \14266 , \14275 );
or \U$14318 ( \14509 , \14506 , \14507 , \14508 );
and \U$14319 ( \14510 , \14290 , \14304 );
and \U$14320 ( \14511 , \14304 , \14408 );
and \U$14321 ( \14512 , \14290 , \14408 );
or \U$14322 ( \14513 , \14510 , \14511 , \14512 );
xor \U$14323 ( \14514 , \14509 , \14513 );
and \U$14324 ( \14515 , \14414 , \14428 );
and \U$14325 ( \14516 , \14428 , \14485 );
and \U$14326 ( \14517 , \14414 , \14485 );
or \U$14327 ( \14518 , \14515 , \14516 , \14517 );
xor \U$14328 ( \14519 , \14514 , \14518 );
xor \U$14329 ( \14520 , \14505 , \14519 );
and \U$14330 ( \14521 , \14241 , \14245 );
and \U$14331 ( \14522 , \14245 , \14250 );
and \U$14332 ( \14523 , \14241 , \14250 );
or \U$14333 ( \14524 , \14521 , \14522 , \14523 );
and \U$14334 ( \14525 , \14276 , \14409 );
and \U$14335 ( \14526 , \14409 , \14486 );
and \U$14336 ( \14527 , \14276 , \14486 );
or \U$14337 ( \14528 , \14525 , \14526 , \14527 );
xor \U$14338 ( \14529 , \14524 , \14528 );
and \U$14339 ( \14530 , \14280 , \14284 );
and \U$14340 ( \14531 , \14284 , \14289 );
and \U$14341 ( \14532 , \14280 , \14289 );
or \U$14342 ( \14533 , \14530 , \14531 , \14532 );
and \U$14343 ( \14534 , \14294 , \14298 );
and \U$14344 ( \14535 , \14298 , \14303 );
and \U$14345 ( \14536 , \14294 , \14303 );
or \U$14346 ( \14537 , \14534 , \14535 , \14536 );
xor \U$14347 ( \14538 , \14533 , \14537 );
and \U$14348 ( \14539 , \14318 , \14362 );
and \U$14349 ( \14540 , \14362 , \14407 );
and \U$14350 ( \14541 , \14318 , \14407 );
or \U$14351 ( \14542 , \14539 , \14540 , \14541 );
xor \U$14352 ( \14543 , \14538 , \14542 );
and \U$14353 ( \14544 , \14443 , \14457 );
and \U$14354 ( \14545 , \14457 , \14484 );
and \U$14355 ( \14546 , \14443 , \14484 );
or \U$14356 ( \14547 , \14544 , \14545 , \14546 );
and \U$14357 ( \14548 , \14381 , \14385 );
and \U$14358 ( \14549 , \14385 , \14390 );
and \U$14359 ( \14550 , \14381 , \14390 );
or \U$14360 ( \14551 , \14548 , \14549 , \14550 );
and \U$14361 ( \14552 , \14462 , \14466 );
and \U$14362 ( \14553 , \14466 , \14468 );
and \U$14363 ( \14554 , \14462 , \14468 );
or \U$14364 ( \14555 , \14552 , \14553 , \14554 );
xor \U$14365 ( \14556 , \14551 , \14555 );
and \U$14366 ( \14557 , \14473 , \14477 );
and \U$14367 ( \14558 , \14477 , \14482 );
and \U$14368 ( \14559 , \14473 , \14482 );
or \U$14369 ( \14560 , \14557 , \14558 , \14559 );
xor \U$14370 ( \14561 , \14556 , \14560 );
and \U$14371 ( \14562 , \14322 , \14326 );
and \U$14372 ( \14563 , \14326 , \14331 );
and \U$14373 ( \14564 , \14322 , \14331 );
or \U$14374 ( \14565 , \14562 , \14563 , \14564 );
and \U$14375 ( \14566 , \14351 , \14355 );
and \U$14376 ( \14567 , \14355 , \14360 );
and \U$14377 ( \14568 , \14351 , \14360 );
or \U$14378 ( \14569 , \14566 , \14567 , \14568 );
xor \U$14379 ( \14570 , \14565 , \14569 );
and \U$14380 ( \14571 , \14308 , \14312 );
and \U$14381 ( \14572 , \14312 , \14317 );
and \U$14382 ( \14573 , \14308 , \14317 );
or \U$14383 ( \14574 , \14571 , \14572 , \14573 );
xor \U$14384 ( \14575 , \14570 , \14574 );
xor \U$14385 ( \14576 , \14561 , \14575 );
and \U$14386 ( \14577 , \14336 , \14340 );
and \U$14387 ( \14578 , \14340 , \14345 );
and \U$14388 ( \14579 , \14336 , \14345 );
or \U$14389 ( \14580 , \14577 , \14578 , \14579 );
and \U$14390 ( \14581 , \14367 , \14371 );
and \U$14391 ( \14582 , \14371 , \14376 );
and \U$14392 ( \14583 , \14367 , \14376 );
or \U$14393 ( \14584 , \14581 , \14582 , \14583 );
xor \U$14394 ( \14585 , \14580 , \14584 );
and \U$14395 ( \14586 , \14396 , \14400 );
and \U$14396 ( \14587 , \14400 , \14405 );
and \U$14397 ( \14588 , \14396 , \14405 );
or \U$14398 ( \14589 , \14586 , \14587 , \14588 );
xor \U$14399 ( \14590 , \14585 , \14589 );
xor \U$14400 ( \14591 , \14576 , \14590 );
xor \U$14401 ( \14592 , \14547 , \14591 );
and \U$14402 ( \14593 , \307 , \9765 );
and \U$14403 ( \14594 , \412 , \9644 );
nor \U$14404 ( \14595 , \14593 , \14594 );
xnor \U$14405 ( \14596 , \14595 , \9478 );
and \U$14406 ( \14597 , \185 , \10408 );
and \U$14407 ( \14598 , \261 , \10116 );
nor \U$14408 ( \14599 , \14597 , \14598 );
xnor \U$14409 ( \14600 , \14599 , \10121 );
xor \U$14410 ( \14601 , \14596 , \14600 );
and \U$14411 ( \14602 , \178 , \10118 );
xor \U$14412 ( \14603 , \14601 , \14602 );
and \U$14413 ( \14604 , \2182 , \6401 );
and \U$14414 ( \14605 , \2366 , \6143 );
nor \U$14415 ( \14606 , \14604 , \14605 );
xnor \U$14416 ( \14607 , \14606 , \6148 );
and \U$14417 ( \14608 , \1948 , \7055 );
and \U$14418 ( \14609 , \2090 , \6675 );
nor \U$14419 ( \14610 , \14608 , \14609 );
xnor \U$14420 ( \14611 , \14610 , \6680 );
xor \U$14421 ( \14612 , \14607 , \14611 );
and \U$14422 ( \14613 , \1684 , \7489 );
and \U$14423 ( \14614 , \1802 , \7137 );
nor \U$14424 ( \14615 , \14613 , \14614 );
xnor \U$14425 ( \14616 , \14615 , \7142 );
xor \U$14426 ( \14617 , \14612 , \14616 );
xor \U$14427 ( \14618 , \14603 , \14617 );
and \U$14428 ( \14619 , \1484 , \8019 );
and \U$14429 ( \14620 , \1601 , \7830 );
nor \U$14430 ( \14621 , \14619 , \14620 );
xnor \U$14431 ( \14622 , \14621 , \7713 );
and \U$14432 ( \14623 , \1192 , \8540 );
and \U$14433 ( \14624 , \1333 , \8292 );
nor \U$14434 ( \14625 , \14623 , \14624 );
xnor \U$14435 ( \14626 , \14625 , \8297 );
xor \U$14436 ( \14627 , \14622 , \14626 );
and \U$14437 ( \14628 , \474 , \9333 );
and \U$14438 ( \14629 , \1147 , \9006 );
nor \U$14439 ( \14630 , \14628 , \14629 );
xnor \U$14440 ( \14631 , \14630 , \8848 );
xor \U$14441 ( \14632 , \14627 , \14631 );
xor \U$14442 ( \14633 , \14618 , \14632 );
and \U$14443 ( \14634 , \5674 , \2669 );
and \U$14444 ( \14635 , \6030 , \2538 );
nor \U$14445 ( \14636 , \14634 , \14635 );
xnor \U$14446 ( \14637 , \14636 , \2534 );
and \U$14447 ( \14638 , \5156 , \3103 );
and \U$14448 ( \14639 , \5469 , \2934 );
nor \U$14449 ( \14640 , \14638 , \14639 );
xnor \U$14450 ( \14641 , \14640 , \2839 );
xor \U$14451 ( \14642 , \14637 , \14641 );
and \U$14452 ( \14643 , \4749 , \3357 );
and \U$14453 ( \14644 , \4922 , \3255 );
nor \U$14454 ( \14645 , \14643 , \14644 );
xnor \U$14455 ( \14646 , \14645 , \3156 );
xor \U$14456 ( \14647 , \14642 , \14646 );
and \U$14457 ( \14648 , \4364 , \3813 );
and \U$14458 ( \14649 , \4654 , \3557 );
nor \U$14459 ( \14650 , \14648 , \14649 );
xnor \U$14460 ( \14651 , \14650 , \3562 );
and \U$14461 ( \14652 , \3912 , \4132 );
and \U$14462 ( \14653 , \4160 , \4012 );
nor \U$14463 ( \14654 , \14652 , \14653 );
xnor \U$14464 ( \14655 , \14654 , \3925 );
xor \U$14465 ( \14656 , \14651 , \14655 );
and \U$14466 ( \14657 , \3646 , \4581 );
and \U$14467 ( \14658 , \3736 , \4424 );
nor \U$14468 ( \14659 , \14657 , \14658 );
xnor \U$14469 ( \14660 , \14659 , \4377 );
xor \U$14470 ( \14661 , \14656 , \14660 );
xor \U$14471 ( \14662 , \14647 , \14661 );
and \U$14472 ( \14663 , \3143 , \5011 );
and \U$14473 ( \14664 , \3395 , \4878 );
nor \U$14474 ( \14665 , \14663 , \14664 );
xnor \U$14475 ( \14666 , \14665 , \4762 );
and \U$14476 ( \14667 , \2826 , \5485 );
and \U$14477 ( \14668 , \3037 , \5275 );
nor \U$14478 ( \14669 , \14667 , \14668 );
xnor \U$14479 ( \14670 , \14669 , \5169 );
xor \U$14480 ( \14671 , \14666 , \14670 );
and \U$14481 ( \14672 , \2521 , \5996 );
and \U$14482 ( \14673 , \2757 , \5695 );
nor \U$14483 ( \14674 , \14672 , \14673 );
xnor \U$14484 ( \14675 , \14674 , \5687 );
xor \U$14485 ( \14676 , \14671 , \14675 );
xor \U$14486 ( \14677 , \14662 , \14676 );
xor \U$14487 ( \14678 , \14633 , \14677 );
and \U$14488 ( \14679 , \8835 , \1086 );
and \U$14489 ( \14680 , \9169 , \508 );
nor \U$14490 ( \14681 , \14679 , \14680 );
xnor \U$14491 ( \14682 , \14681 , \487 );
and \U$14492 ( \14683 , \8349 , \1301 );
and \U$14493 ( \14684 , \8652 , \1246 );
nor \U$14494 ( \14685 , \14683 , \14684 );
xnor \U$14495 ( \14686 , \14685 , \1205 );
xor \U$14496 ( \14687 , \14682 , \14686 );
and \U$14497 ( \14688 , \7700 , \1578 );
and \U$14498 ( \14689 , \8057 , \1431 );
nor \U$14499 ( \14690 , \14688 , \14689 );
xnor \U$14500 ( \14691 , \14690 , \1436 );
xor \U$14501 ( \14692 , \14687 , \14691 );
and \U$14502 ( \14693 , \7231 , \1824 );
and \U$14503 ( \14694 , \7556 , \1739 );
nor \U$14504 ( \14695 , \14693 , \14694 );
xnor \U$14505 ( \14696 , \14695 , \1697 );
and \U$14506 ( \14697 , \6790 , \2121 );
and \U$14507 ( \14698 , \6945 , \2008 );
nor \U$14508 ( \14699 , \14697 , \14698 );
xnor \U$14509 ( \14700 , \14699 , \1961 );
xor \U$14510 ( \14701 , \14696 , \14700 );
and \U$14511 ( \14702 , \6281 , \2400 );
and \U$14512 ( \14703 , \6514 , \2246 );
nor \U$14513 ( \14704 , \14702 , \14703 );
xnor \U$14514 ( \14705 , \14704 , \2195 );
xor \U$14515 ( \14706 , \14701 , \14705 );
xor \U$14516 ( \14707 , \14692 , \14706 );
not \U$14517 ( \14708 , \163 );
and \U$14518 ( \14709 , \10206 , \296 );
and \U$14519 ( \14710 , \10584 , \168 );
nor \U$14520 ( \14711 , \14709 , \14710 );
xnor \U$14521 ( \14712 , \14711 , \173 );
xor \U$14522 ( \14713 , \14708 , \14712 );
and \U$14523 ( \14714 , \9465 , \438 );
and \U$14524 ( \14715 , \9897 , \336 );
nor \U$14525 ( \14716 , \14714 , \14715 );
xnor \U$14526 ( \14717 , \14716 , \320 );
xor \U$14527 ( \14718 , \14713 , \14717 );
xor \U$14528 ( \14719 , \14707 , \14718 );
xor \U$14529 ( \14720 , \14678 , \14719 );
xor \U$14530 ( \14721 , \14592 , \14720 );
xor \U$14531 ( \14722 , \14543 , \14721 );
and \U$14532 ( \14723 , \14332 , \14346 );
and \U$14533 ( \14724 , \14346 , \14361 );
and \U$14534 ( \14725 , \14332 , \14361 );
or \U$14535 ( \14726 , \14723 , \14724 , \14725 );
and \U$14536 ( \14727 , \14377 , \14391 );
and \U$14537 ( \14728 , \14391 , \14406 );
and \U$14538 ( \14729 , \14377 , \14406 );
or \U$14539 ( \14730 , \14727 , \14728 , \14729 );
xor \U$14540 ( \14731 , \14726 , \14730 );
or \U$14541 ( \14732 , \14469 , \14483 );
xor \U$14542 ( \14733 , \14731 , \14732 );
and \U$14543 ( \14734 , \14433 , \14437 );
and \U$14544 ( \14735 , \14437 , \14442 );
and \U$14545 ( \14736 , \14433 , \14442 );
or \U$14546 ( \14737 , \14734 , \14735 , \14736 );
and \U$14547 ( \14738 , \14418 , \14422 );
and \U$14548 ( \14739 , \14422 , \14427 );
and \U$14549 ( \14740 , \14418 , \14427 );
or \U$14550 ( \14741 , \14738 , \14739 , \14740 );
xor \U$14551 ( \14742 , \14737 , \14741 );
and \U$14552 ( \14743 , \14447 , \14451 );
and \U$14553 ( \14744 , \14451 , \14456 );
and \U$14554 ( \14745 , \14447 , \14456 );
or \U$14555 ( \14746 , \14743 , \14744 , \14745 );
xor \U$14556 ( \14747 , \14742 , \14746 );
xor \U$14557 ( \14748 , \14733 , \14747 );
xor \U$14558 ( \14749 , \14722 , \14748 );
xor \U$14559 ( \14750 , \14529 , \14749 );
xor \U$14560 ( \14751 , \14520 , \14750 );
xor \U$14561 ( \14752 , \14501 , \14751 );
and \U$14562 ( \14753 , \14231 , \14252 );
and \U$14563 ( \14754 , \14252 , \14488 );
and \U$14564 ( \14755 , \14231 , \14488 );
or \U$14565 ( \14756 , \14753 , \14754 , \14755 );
xor \U$14566 ( \14757 , \14752 , \14756 );
and \U$14567 ( \14758 , \14489 , \14490 );
and \U$14568 ( \14759 , \14491 , \14494 );
or \U$14569 ( \14760 , \14758 , \14759 );
xor \U$14570 ( \14761 , \14757 , \14760 );
buf g5501_GF_PartitionCandidate( \14762_nG5501 , \14761 );
buf \U$14571 ( \14763 , \14762_nG5501 );
and \U$14572 ( \14764 , \14505 , \14519 );
and \U$14573 ( \14765 , \14519 , \14750 );
and \U$14574 ( \14766 , \14505 , \14750 );
or \U$14575 ( \14767 , \14764 , \14765 , \14766 );
and \U$14576 ( \14768 , \14524 , \14528 );
and \U$14577 ( \14769 , \14528 , \14749 );
and \U$14578 ( \14770 , \14524 , \14749 );
or \U$14579 ( \14771 , \14768 , \14769 , \14770 );
and \U$14580 ( \14772 , \14533 , \14537 );
and \U$14581 ( \14773 , \14537 , \14542 );
and \U$14582 ( \14774 , \14533 , \14542 );
or \U$14583 ( \14775 , \14772 , \14773 , \14774 );
and \U$14584 ( \14776 , \14547 , \14591 );
and \U$14585 ( \14777 , \14591 , \14720 );
and \U$14586 ( \14778 , \14547 , \14720 );
or \U$14587 ( \14779 , \14776 , \14777 , \14778 );
xor \U$14588 ( \14780 , \14775 , \14779 );
and \U$14589 ( \14781 , \14733 , \14747 );
xor \U$14590 ( \14782 , \14780 , \14781 );
xor \U$14591 ( \14783 , \14771 , \14782 );
and \U$14592 ( \14784 , \14509 , \14513 );
and \U$14593 ( \14785 , \14513 , \14518 );
and \U$14594 ( \14786 , \14509 , \14518 );
or \U$14595 ( \14787 , \14784 , \14785 , \14786 );
and \U$14596 ( \14788 , \14543 , \14721 );
and \U$14597 ( \14789 , \14721 , \14748 );
and \U$14598 ( \14790 , \14543 , \14748 );
or \U$14599 ( \14791 , \14788 , \14789 , \14790 );
xor \U$14600 ( \14792 , \14787 , \14791 );
and \U$14601 ( \14793 , \14726 , \14730 );
and \U$14602 ( \14794 , \14730 , \14732 );
and \U$14603 ( \14795 , \14726 , \14732 );
or \U$14604 ( \14796 , \14793 , \14794 , \14795 );
and \U$14605 ( \14797 , \14737 , \14741 );
and \U$14606 ( \14798 , \14741 , \14746 );
and \U$14607 ( \14799 , \14737 , \14746 );
or \U$14608 ( \14800 , \14797 , \14798 , \14799 );
xor \U$14609 ( \14801 , \14796 , \14800 );
and \U$14610 ( \14802 , \14633 , \14677 );
and \U$14611 ( \14803 , \14677 , \14719 );
and \U$14612 ( \14804 , \14633 , \14719 );
or \U$14613 ( \14805 , \14802 , \14803 , \14804 );
xor \U$14614 ( \14806 , \14801 , \14805 );
and \U$14615 ( \14807 , \14561 , \14575 );
and \U$14616 ( \14808 , \14575 , \14590 );
and \U$14617 ( \14809 , \14561 , \14590 );
or \U$14618 ( \14810 , \14807 , \14808 , \14809 );
and \U$14619 ( \14811 , \14637 , \14641 );
and \U$14620 ( \14812 , \14641 , \14646 );
and \U$14621 ( \14813 , \14637 , \14646 );
or \U$14622 ( \14814 , \14811 , \14812 , \14813 );
and \U$14623 ( \14815 , \14651 , \14655 );
and \U$14624 ( \14816 , \14655 , \14660 );
and \U$14625 ( \14817 , \14651 , \14660 );
or \U$14626 ( \14818 , \14815 , \14816 , \14817 );
xor \U$14627 ( \14819 , \14814 , \14818 );
and \U$14628 ( \14820 , \14666 , \14670 );
and \U$14629 ( \14821 , \14670 , \14675 );
and \U$14630 ( \14822 , \14666 , \14675 );
or \U$14631 ( \14823 , \14820 , \14821 , \14822 );
xor \U$14632 ( \14824 , \14819 , \14823 );
and \U$14633 ( \14825 , \14682 , \14686 );
and \U$14634 ( \14826 , \14686 , \14691 );
and \U$14635 ( \14827 , \14682 , \14691 );
or \U$14636 ( \14828 , \14825 , \14826 , \14827 );
and \U$14637 ( \14829 , \14696 , \14700 );
and \U$14638 ( \14830 , \14700 , \14705 );
and \U$14639 ( \14831 , \14696 , \14705 );
or \U$14640 ( \14832 , \14829 , \14830 , \14831 );
xor \U$14641 ( \14833 , \14828 , \14832 );
and \U$14642 ( \14834 , \14708 , \14712 );
and \U$14643 ( \14835 , \14712 , \14717 );
and \U$14644 ( \14836 , \14708 , \14717 );
or \U$14645 ( \14837 , \14834 , \14835 , \14836 );
xor \U$14646 ( \14838 , \14833 , \14837 );
xor \U$14647 ( \14839 , \14824 , \14838 );
and \U$14648 ( \14840 , \14596 , \14600 );
and \U$14649 ( \14841 , \14600 , \14602 );
and \U$14650 ( \14842 , \14596 , \14602 );
or \U$14651 ( \14843 , \14840 , \14841 , \14842 );
and \U$14652 ( \14844 , \14607 , \14611 );
and \U$14653 ( \14845 , \14611 , \14616 );
and \U$14654 ( \14846 , \14607 , \14616 );
or \U$14655 ( \14847 , \14844 , \14845 , \14846 );
xor \U$14656 ( \14848 , \14843 , \14847 );
and \U$14657 ( \14849 , \14622 , \14626 );
and \U$14658 ( \14850 , \14626 , \14631 );
and \U$14659 ( \14851 , \14622 , \14631 );
or \U$14660 ( \14852 , \14849 , \14850 , \14851 );
xor \U$14661 ( \14853 , \14848 , \14852 );
xor \U$14662 ( \14854 , \14839 , \14853 );
xor \U$14663 ( \14855 , \14810 , \14854 );
and \U$14664 ( \14856 , \4160 , \4132 );
and \U$14665 ( \14857 , \4364 , \4012 );
nor \U$14666 ( \14858 , \14856 , \14857 );
xnor \U$14667 ( \14859 , \14858 , \3925 );
and \U$14668 ( \14860 , \3736 , \4581 );
and \U$14669 ( \14861 , \3912 , \4424 );
nor \U$14670 ( \14862 , \14860 , \14861 );
xnor \U$14671 ( \14863 , \14862 , \4377 );
xor \U$14672 ( \14864 , \14859 , \14863 );
and \U$14673 ( \14865 , \3395 , \5011 );
and \U$14674 ( \14866 , \3646 , \4878 );
nor \U$14675 ( \14867 , \14865 , \14866 );
xnor \U$14676 ( \14868 , \14867 , \4762 );
xor \U$14677 ( \14869 , \14864 , \14868 );
and \U$14678 ( \14870 , \3037 , \5485 );
and \U$14679 ( \14871 , \3143 , \5275 );
nor \U$14680 ( \14872 , \14870 , \14871 );
xnor \U$14681 ( \14873 , \14872 , \5169 );
and \U$14682 ( \14874 , \2757 , \5996 );
and \U$14683 ( \14875 , \2826 , \5695 );
nor \U$14684 ( \14876 , \14874 , \14875 );
xnor \U$14685 ( \14877 , \14876 , \5687 );
xor \U$14686 ( \14878 , \14873 , \14877 );
and \U$14687 ( \14879 , \2366 , \6401 );
and \U$14688 ( \14880 , \2521 , \6143 );
nor \U$14689 ( \14881 , \14879 , \14880 );
xnor \U$14690 ( \14882 , \14881 , \6148 );
xor \U$14691 ( \14883 , \14878 , \14882 );
xor \U$14692 ( \14884 , \14869 , \14883 );
and \U$14693 ( \14885 , \5469 , \3103 );
and \U$14694 ( \14886 , \5674 , \2934 );
nor \U$14695 ( \14887 , \14885 , \14886 );
xnor \U$14696 ( \14888 , \14887 , \2839 );
and \U$14697 ( \14889 , \4922 , \3357 );
and \U$14698 ( \14890 , \5156 , \3255 );
nor \U$14699 ( \14891 , \14889 , \14890 );
xnor \U$14700 ( \14892 , \14891 , \3156 );
xor \U$14701 ( \14893 , \14888 , \14892 );
and \U$14702 ( \14894 , \4654 , \3813 );
and \U$14703 ( \14895 , \4749 , \3557 );
nor \U$14704 ( \14896 , \14894 , \14895 );
xnor \U$14705 ( \14897 , \14896 , \3562 );
xor \U$14706 ( \14898 , \14893 , \14897 );
xor \U$14707 ( \14899 , \14884 , \14898 );
and \U$14708 ( \14900 , \6945 , \2121 );
and \U$14709 ( \14901 , \7231 , \2008 );
nor \U$14710 ( \14902 , \14900 , \14901 );
xnor \U$14711 ( \14903 , \14902 , \1961 );
and \U$14712 ( \14904 , \6514 , \2400 );
and \U$14713 ( \14905 , \6790 , \2246 );
nor \U$14714 ( \14906 , \14904 , \14905 );
xnor \U$14715 ( \14907 , \14906 , \2195 );
xor \U$14716 ( \14908 , \14903 , \14907 );
and \U$14717 ( \14909 , \6030 , \2669 );
and \U$14718 ( \14910 , \6281 , \2538 );
nor \U$14719 ( \14911 , \14909 , \14910 );
xnor \U$14720 ( \14912 , \14911 , \2534 );
xor \U$14721 ( \14913 , \14908 , \14912 );
and \U$14722 ( \14914 , \8652 , \1301 );
and \U$14723 ( \14915 , \8835 , \1246 );
nor \U$14724 ( \14916 , \14914 , \14915 );
xnor \U$14725 ( \14917 , \14916 , \1205 );
and \U$14726 ( \14918 , \8057 , \1578 );
and \U$14727 ( \14919 , \8349 , \1431 );
nor \U$14728 ( \14920 , \14918 , \14919 );
xnor \U$14729 ( \14921 , \14920 , \1436 );
xor \U$14730 ( \14922 , \14917 , \14921 );
and \U$14731 ( \14923 , \7556 , \1824 );
and \U$14732 ( \14924 , \7700 , \1739 );
nor \U$14733 ( \14925 , \14923 , \14924 );
xnor \U$14734 ( \14926 , \14925 , \1697 );
xor \U$14735 ( \14927 , \14922 , \14926 );
xor \U$14736 ( \14928 , \14913 , \14927 );
and \U$14737 ( \14929 , \10584 , \296 );
not \U$14738 ( \14930 , \14929 );
xnor \U$14739 ( \14931 , \14930 , \173 );
and \U$14740 ( \14932 , \9897 , \438 );
and \U$14741 ( \14933 , \10206 , \336 );
nor \U$14742 ( \14934 , \14932 , \14933 );
xnor \U$14743 ( \14935 , \14934 , \320 );
xor \U$14744 ( \14936 , \14931 , \14935 );
and \U$14745 ( \14937 , \9169 , \1086 );
and \U$14746 ( \14938 , \9465 , \508 );
nor \U$14747 ( \14939 , \14937 , \14938 );
xnor \U$14748 ( \14940 , \14939 , \487 );
xor \U$14749 ( \14941 , \14936 , \14940 );
xor \U$14750 ( \14942 , \14928 , \14941 );
xor \U$14751 ( \14943 , \14899 , \14942 );
and \U$14752 ( \14944 , \2090 , \7055 );
and \U$14753 ( \14945 , \2182 , \6675 );
nor \U$14754 ( \14946 , \14944 , \14945 );
xnor \U$14755 ( \14947 , \14946 , \6680 );
and \U$14756 ( \14948 , \1802 , \7489 );
and \U$14757 ( \14949 , \1948 , \7137 );
nor \U$14758 ( \14950 , \14948 , \14949 );
xnor \U$14759 ( \14951 , \14950 , \7142 );
xor \U$14760 ( \14952 , \14947 , \14951 );
and \U$14761 ( \14953 , \1601 , \8019 );
and \U$14762 ( \14954 , \1684 , \7830 );
nor \U$14763 ( \14955 , \14953 , \14954 );
xnor \U$14764 ( \14956 , \14955 , \7713 );
xor \U$14765 ( \14957 , \14952 , \14956 );
and \U$14766 ( \14958 , \1333 , \8540 );
and \U$14767 ( \14959 , \1484 , \8292 );
nor \U$14768 ( \14960 , \14958 , \14959 );
xnor \U$14769 ( \14961 , \14960 , \8297 );
and \U$14770 ( \14962 , \1147 , \9333 );
and \U$14771 ( \14963 , \1192 , \9006 );
nor \U$14772 ( \14964 , \14962 , \14963 );
xnor \U$14773 ( \14965 , \14964 , \8848 );
xor \U$14774 ( \14966 , \14961 , \14965 );
and \U$14775 ( \14967 , \412 , \9765 );
and \U$14776 ( \14968 , \474 , \9644 );
nor \U$14777 ( \14969 , \14967 , \14968 );
xnor \U$14778 ( \14970 , \14969 , \9478 );
xor \U$14779 ( \14971 , \14966 , \14970 );
xor \U$14780 ( \14972 , \14957 , \14971 );
and \U$14781 ( \14973 , \261 , \10408 );
and \U$14782 ( \14974 , \307 , \10116 );
nor \U$14783 ( \14975 , \14973 , \14974 );
xnor \U$14784 ( \14976 , \14975 , \10121 );
and \U$14785 ( \14977 , \185 , \10118 );
xnor \U$14786 ( \14978 , \14976 , \14977 );
xor \U$14787 ( \14979 , \14972 , \14978 );
xor \U$14788 ( \14980 , \14943 , \14979 );
xor \U$14789 ( \14981 , \14855 , \14980 );
xor \U$14790 ( \14982 , \14806 , \14981 );
and \U$14791 ( \14983 , \14551 , \14555 );
and \U$14792 ( \14984 , \14555 , \14560 );
and \U$14793 ( \14985 , \14551 , \14560 );
or \U$14794 ( \14986 , \14983 , \14984 , \14985 );
and \U$14795 ( \14987 , \14565 , \14569 );
and \U$14796 ( \14988 , \14569 , \14574 );
and \U$14797 ( \14989 , \14565 , \14574 );
or \U$14798 ( \14990 , \14987 , \14988 , \14989 );
xor \U$14799 ( \14991 , \14986 , \14990 );
and \U$14800 ( \14992 , \14580 , \14584 );
and \U$14801 ( \14993 , \14584 , \14589 );
and \U$14802 ( \14994 , \14580 , \14589 );
or \U$14803 ( \14995 , \14992 , \14993 , \14994 );
xor \U$14804 ( \14996 , \14991 , \14995 );
and \U$14805 ( \14997 , \14603 , \14617 );
and \U$14806 ( \14998 , \14617 , \14632 );
and \U$14807 ( \14999 , \14603 , \14632 );
or \U$14808 ( \15000 , \14997 , \14998 , \14999 );
and \U$14809 ( \15001 , \14647 , \14661 );
and \U$14810 ( \15002 , \14661 , \14676 );
and \U$14811 ( \15003 , \14647 , \14676 );
or \U$14812 ( \15004 , \15001 , \15002 , \15003 );
xor \U$14813 ( \15005 , \15000 , \15004 );
and \U$14814 ( \15006 , \14692 , \14706 );
and \U$14815 ( \15007 , \14706 , \14718 );
and \U$14816 ( \15008 , \14692 , \14718 );
or \U$14817 ( \15009 , \15006 , \15007 , \15008 );
xor \U$14818 ( \15010 , \15005 , \15009 );
xor \U$14819 ( \15011 , \14996 , \15010 );
xor \U$14820 ( \15012 , \14982 , \15011 );
xor \U$14821 ( \15013 , \14792 , \15012 );
xor \U$14822 ( \15014 , \14783 , \15013 );
xor \U$14823 ( \15015 , \14767 , \15014 );
and \U$14824 ( \15016 , \14501 , \14751 );
xor \U$14825 ( \15017 , \15015 , \15016 );
and \U$14826 ( \15018 , \14752 , \14756 );
and \U$14827 ( \15019 , \14757 , \14760 );
or \U$14828 ( \15020 , \15018 , \15019 );
xor \U$14829 ( \15021 , \15017 , \15020 );
buf g54ff_GF_PartitionCandidate( \15022_nG54ff , \15021 );
buf \U$14830 ( \15023 , \15022_nG54ff );
and \U$14831 ( \15024 , \14771 , \14782 );
and \U$14832 ( \15025 , \14782 , \15013 );
and \U$14833 ( \15026 , \14771 , \15013 );
or \U$14834 ( \15027 , \15024 , \15025 , \15026 );
and \U$14835 ( \15028 , \14787 , \14791 );
and \U$14836 ( \15029 , \14791 , \15012 );
and \U$14837 ( \15030 , \14787 , \15012 );
or \U$14838 ( \15031 , \15028 , \15029 , \15030 );
and \U$14839 ( \15032 , \14796 , \14800 );
and \U$14840 ( \15033 , \14800 , \14805 );
and \U$14841 ( \15034 , \14796 , \14805 );
or \U$14842 ( \15035 , \15032 , \15033 , \15034 );
and \U$14843 ( \15036 , \14810 , \14854 );
and \U$14844 ( \15037 , \14854 , \14980 );
and \U$14845 ( \15038 , \14810 , \14980 );
or \U$14846 ( \15039 , \15036 , \15037 , \15038 );
xor \U$14847 ( \15040 , \15035 , \15039 );
and \U$14848 ( \15041 , \14996 , \15010 );
xor \U$14849 ( \15042 , \15040 , \15041 );
xor \U$14850 ( \15043 , \15031 , \15042 );
and \U$14851 ( \15044 , \14775 , \14779 );
and \U$14852 ( \15045 , \14779 , \14781 );
and \U$14853 ( \15046 , \14775 , \14781 );
or \U$14854 ( \15047 , \15044 , \15045 , \15046 );
and \U$14855 ( \15048 , \14806 , \14981 );
and \U$14856 ( \15049 , \14981 , \15011 );
and \U$14857 ( \15050 , \14806 , \15011 );
or \U$14858 ( \15051 , \15048 , \15049 , \15050 );
xor \U$14859 ( \15052 , \15047 , \15051 );
and \U$14860 ( \15053 , \14986 , \14990 );
and \U$14861 ( \15054 , \14990 , \14995 );
and \U$14862 ( \15055 , \14986 , \14995 );
or \U$14863 ( \15056 , \15053 , \15054 , \15055 );
and \U$14864 ( \15057 , \15000 , \15004 );
and \U$14865 ( \15058 , \15004 , \15009 );
and \U$14866 ( \15059 , \15000 , \15009 );
or \U$14867 ( \15060 , \15057 , \15058 , \15059 );
xor \U$14868 ( \15061 , \15056 , \15060 );
and \U$14869 ( \15062 , \14899 , \14942 );
and \U$14870 ( \15063 , \14942 , \14979 );
and \U$14871 ( \15064 , \14899 , \14979 );
or \U$14872 ( \15065 , \15062 , \15063 , \15064 );
xor \U$14873 ( \15066 , \15061 , \15065 );
and \U$14874 ( \15067 , \14824 , \14838 );
and \U$14875 ( \15068 , \14838 , \14853 );
and \U$14876 ( \15069 , \14824 , \14853 );
or \U$14877 ( \15070 , \15067 , \15068 , \15069 );
and \U$14878 ( \15071 , \14947 , \14951 );
and \U$14879 ( \15072 , \14951 , \14956 );
and \U$14880 ( \15073 , \14947 , \14956 );
or \U$14881 ( \15074 , \15071 , \15072 , \15073 );
and \U$14882 ( \15075 , \14961 , \14965 );
and \U$14883 ( \15076 , \14965 , \14970 );
and \U$14884 ( \15077 , \14961 , \14970 );
or \U$14885 ( \15078 , \15075 , \15076 , \15077 );
xor \U$14886 ( \15079 , \15074 , \15078 );
or \U$14887 ( \15080 , \14976 , \14977 );
xor \U$14888 ( \15081 , \15079 , \15080 );
and \U$14889 ( \15082 , \14903 , \14907 );
and \U$14890 ( \15083 , \14907 , \14912 );
and \U$14891 ( \15084 , \14903 , \14912 );
or \U$14892 ( \15085 , \15082 , \15083 , \15084 );
and \U$14893 ( \15086 , \14917 , \14921 );
and \U$14894 ( \15087 , \14921 , \14926 );
and \U$14895 ( \15088 , \14917 , \14926 );
or \U$14896 ( \15089 , \15086 , \15087 , \15088 );
xor \U$14897 ( \15090 , \15085 , \15089 );
and \U$14898 ( \15091 , \14931 , \14935 );
and \U$14899 ( \15092 , \14935 , \14940 );
and \U$14900 ( \15093 , \14931 , \14940 );
or \U$14901 ( \15094 , \15091 , \15092 , \15093 );
xor \U$14902 ( \15095 , \15090 , \15094 );
xor \U$14903 ( \15096 , \15081 , \15095 );
and \U$14904 ( \15097 , \14859 , \14863 );
and \U$14905 ( \15098 , \14863 , \14868 );
and \U$14906 ( \15099 , \14859 , \14868 );
or \U$14907 ( \15100 , \15097 , \15098 , \15099 );
and \U$14908 ( \15101 , \14873 , \14877 );
and \U$14909 ( \15102 , \14877 , \14882 );
and \U$14910 ( \15103 , \14873 , \14882 );
or \U$14911 ( \15104 , \15101 , \15102 , \15103 );
xor \U$14912 ( \15105 , \15100 , \15104 );
and \U$14913 ( \15106 , \14888 , \14892 );
and \U$14914 ( \15107 , \14892 , \14897 );
and \U$14915 ( \15108 , \14888 , \14897 );
or \U$14916 ( \15109 , \15106 , \15107 , \15108 );
xor \U$14917 ( \15110 , \15105 , \15109 );
xor \U$14918 ( \15111 , \15096 , \15110 );
xor \U$14919 ( \15112 , \15070 , \15111 );
and \U$14920 ( \15113 , \5674 , \3103 );
and \U$14921 ( \15114 , \6030 , \2934 );
nor \U$14922 ( \15115 , \15113 , \15114 );
xnor \U$14923 ( \15116 , \15115 , \2839 );
and \U$14924 ( \15117 , \5156 , \3357 );
and \U$14925 ( \15118 , \5469 , \3255 );
nor \U$14926 ( \15119 , \15117 , \15118 );
xnor \U$14927 ( \15120 , \15119 , \3156 );
xor \U$14928 ( \15121 , \15116 , \15120 );
and \U$14929 ( \15122 , \4749 , \3813 );
and \U$14930 ( \15123 , \4922 , \3557 );
nor \U$14931 ( \15124 , \15122 , \15123 );
xnor \U$14932 ( \15125 , \15124 , \3562 );
xor \U$14933 ( \15126 , \15121 , \15125 );
and \U$14934 ( \15127 , \4364 , \4132 );
and \U$14935 ( \15128 , \4654 , \4012 );
nor \U$14936 ( \15129 , \15127 , \15128 );
xnor \U$14937 ( \15130 , \15129 , \3925 );
and \U$14938 ( \15131 , \3912 , \4581 );
and \U$14939 ( \15132 , \4160 , \4424 );
nor \U$14940 ( \15133 , \15131 , \15132 );
xnor \U$14941 ( \15134 , \15133 , \4377 );
xor \U$14942 ( \15135 , \15130 , \15134 );
and \U$14943 ( \15136 , \3646 , \5011 );
and \U$14944 ( \15137 , \3736 , \4878 );
nor \U$14945 ( \15138 , \15136 , \15137 );
xnor \U$14946 ( \15139 , \15138 , \4762 );
xor \U$14947 ( \15140 , \15135 , \15139 );
xor \U$14948 ( \15141 , \15126 , \15140 );
and \U$14949 ( \15142 , \3143 , \5485 );
and \U$14950 ( \15143 , \3395 , \5275 );
nor \U$14951 ( \15144 , \15142 , \15143 );
xnor \U$14952 ( \15145 , \15144 , \5169 );
and \U$14953 ( \15146 , \2826 , \5996 );
and \U$14954 ( \15147 , \3037 , \5695 );
nor \U$14955 ( \15148 , \15146 , \15147 );
xnor \U$14956 ( \15149 , \15148 , \5687 );
xor \U$14957 ( \15150 , \15145 , \15149 );
and \U$14958 ( \15151 , \2521 , \6401 );
and \U$14959 ( \15152 , \2757 , \6143 );
nor \U$14960 ( \15153 , \15151 , \15152 );
xnor \U$14961 ( \15154 , \15153 , \6148 );
xor \U$14962 ( \15155 , \15150 , \15154 );
xor \U$14963 ( \15156 , \15141 , \15155 );
and \U$14964 ( \15157 , \8835 , \1301 );
and \U$14965 ( \15158 , \9169 , \1246 );
nor \U$14966 ( \15159 , \15157 , \15158 );
xnor \U$14967 ( \15160 , \15159 , \1205 );
and \U$14968 ( \15161 , \8349 , \1578 );
and \U$14969 ( \15162 , \8652 , \1431 );
nor \U$14970 ( \15163 , \15161 , \15162 );
xnor \U$14971 ( \15164 , \15163 , \1436 );
xor \U$14972 ( \15165 , \15160 , \15164 );
and \U$14973 ( \15166 , \7700 , \1824 );
and \U$14974 ( \15167 , \8057 , \1739 );
nor \U$14975 ( \15168 , \15166 , \15167 );
xnor \U$14976 ( \15169 , \15168 , \1697 );
xor \U$14977 ( \15170 , \15165 , \15169 );
not \U$14978 ( \15171 , \173 );
and \U$14979 ( \15172 , \10206 , \438 );
and \U$14980 ( \15173 , \10584 , \336 );
nor \U$14981 ( \15174 , \15172 , \15173 );
xnor \U$14982 ( \15175 , \15174 , \320 );
xor \U$14983 ( \15176 , \15171 , \15175 );
and \U$14984 ( \15177 , \9465 , \1086 );
and \U$14985 ( \15178 , \9897 , \508 );
nor \U$14986 ( \15179 , \15177 , \15178 );
xnor \U$14987 ( \15180 , \15179 , \487 );
xor \U$14988 ( \15181 , \15176 , \15180 );
xor \U$14989 ( \15182 , \15170 , \15181 );
and \U$14990 ( \15183 , \7231 , \2121 );
and \U$14991 ( \15184 , \7556 , \2008 );
nor \U$14992 ( \15185 , \15183 , \15184 );
xnor \U$14993 ( \15186 , \15185 , \1961 );
and \U$14994 ( \15187 , \6790 , \2400 );
and \U$14995 ( \15188 , \6945 , \2246 );
nor \U$14996 ( \15189 , \15187 , \15188 );
xnor \U$14997 ( \15190 , \15189 , \2195 );
xor \U$14998 ( \15191 , \15186 , \15190 );
and \U$14999 ( \15192 , \6281 , \2669 );
and \U$15000 ( \15193 , \6514 , \2538 );
nor \U$15001 ( \15194 , \15192 , \15193 );
xnor \U$15002 ( \15195 , \15194 , \2534 );
xor \U$15003 ( \15196 , \15191 , \15195 );
xor \U$15004 ( \15197 , \15182 , \15196 );
xor \U$15005 ( \15198 , \15156 , \15197 );
and \U$15006 ( \15199 , \2182 , \7055 );
and \U$15007 ( \15200 , \2366 , \6675 );
nor \U$15008 ( \15201 , \15199 , \15200 );
xnor \U$15009 ( \15202 , \15201 , \6680 );
and \U$15010 ( \15203 , \1948 , \7489 );
and \U$15011 ( \15204 , \2090 , \7137 );
nor \U$15012 ( \15205 , \15203 , \15204 );
xnor \U$15013 ( \15206 , \15205 , \7142 );
xor \U$15014 ( \15207 , \15202 , \15206 );
and \U$15015 ( \15208 , \1684 , \8019 );
and \U$15016 ( \15209 , \1802 , \7830 );
nor \U$15017 ( \15210 , \15208 , \15209 );
xnor \U$15018 ( \15211 , \15210 , \7713 );
xor \U$15019 ( \15212 , \15207 , \15211 );
and \U$15020 ( \15213 , \1484 , \8540 );
and \U$15021 ( \15214 , \1601 , \8292 );
nor \U$15022 ( \15215 , \15213 , \15214 );
xnor \U$15023 ( \15216 , \15215 , \8297 );
and \U$15024 ( \15217 , \1192 , \9333 );
and \U$15025 ( \15218 , \1333 , \9006 );
nor \U$15026 ( \15219 , \15217 , \15218 );
xnor \U$15027 ( \15220 , \15219 , \8848 );
xor \U$15028 ( \15221 , \15216 , \15220 );
and \U$15029 ( \15222 , \474 , \9765 );
and \U$15030 ( \15223 , \1147 , \9644 );
nor \U$15031 ( \15224 , \15222 , \15223 );
xnor \U$15032 ( \15225 , \15224 , \9478 );
xor \U$15033 ( \15226 , \15221 , \15225 );
xor \U$15034 ( \15227 , \15212 , \15226 );
and \U$15035 ( \15228 , \307 , \10408 );
and \U$15036 ( \15229 , \412 , \10116 );
nor \U$15037 ( \15230 , \15228 , \15229 );
xnor \U$15038 ( \15231 , \15230 , \10121 );
and \U$15039 ( \15232 , \261 , \10118 );
xor \U$15040 ( \15233 , \15231 , \15232 );
xor \U$15041 ( \15234 , \15227 , \15233 );
xor \U$15042 ( \15235 , \15198 , \15234 );
xor \U$15043 ( \15236 , \15112 , \15235 );
xor \U$15044 ( \15237 , \15066 , \15236 );
and \U$15045 ( \15238 , \14814 , \14818 );
and \U$15046 ( \15239 , \14818 , \14823 );
and \U$15047 ( \15240 , \14814 , \14823 );
or \U$15048 ( \15241 , \15238 , \15239 , \15240 );
and \U$15049 ( \15242 , \14828 , \14832 );
and \U$15050 ( \15243 , \14832 , \14837 );
and \U$15051 ( \15244 , \14828 , \14837 );
or \U$15052 ( \15245 , \15242 , \15243 , \15244 );
xor \U$15053 ( \15246 , \15241 , \15245 );
and \U$15054 ( \15247 , \14843 , \14847 );
and \U$15055 ( \15248 , \14847 , \14852 );
and \U$15056 ( \15249 , \14843 , \14852 );
or \U$15057 ( \15250 , \15247 , \15248 , \15249 );
xor \U$15058 ( \15251 , \15246 , \15250 );
and \U$15059 ( \15252 , \14869 , \14883 );
and \U$15060 ( \15253 , \14883 , \14898 );
and \U$15061 ( \15254 , \14869 , \14898 );
or \U$15062 ( \15255 , \15252 , \15253 , \15254 );
and \U$15063 ( \15256 , \14913 , \14927 );
and \U$15064 ( \15257 , \14927 , \14941 );
and \U$15065 ( \15258 , \14913 , \14941 );
or \U$15066 ( \15259 , \15256 , \15257 , \15258 );
xor \U$15067 ( \15260 , \15255 , \15259 );
and \U$15068 ( \15261 , \14957 , \14971 );
and \U$15069 ( \15262 , \14971 , \14978 );
and \U$15070 ( \15263 , \14957 , \14978 );
or \U$15071 ( \15264 , \15261 , \15262 , \15263 );
xor \U$15072 ( \15265 , \15260 , \15264 );
xor \U$15073 ( \15266 , \15251 , \15265 );
xor \U$15074 ( \15267 , \15237 , \15266 );
xor \U$15075 ( \15268 , \15052 , \15267 );
xor \U$15076 ( \15269 , \15043 , \15268 );
xor \U$15077 ( \15270 , \15027 , \15269 );
and \U$15078 ( \15271 , \14767 , \15014 );
xor \U$15079 ( \15272 , \15270 , \15271 );
and \U$15080 ( \15273 , \15015 , \15016 );
and \U$15081 ( \15274 , \15017 , \15020 );
or \U$15082 ( \15275 , \15273 , \15274 );
xor \U$15083 ( \15276 , \15272 , \15275 );
buf g54fd_GF_PartitionCandidate( \15277_nG54fd , \15276 );
buf \U$15084 ( \15278 , \15277_nG54fd );
and \U$15085 ( \15279 , \15031 , \15042 );
and \U$15086 ( \15280 , \15042 , \15268 );
and \U$15087 ( \15281 , \15031 , \15268 );
or \U$15088 ( \15282 , \15279 , \15280 , \15281 );
and \U$15089 ( \15283 , \15047 , \15051 );
and \U$15090 ( \15284 , \15051 , \15267 );
and \U$15091 ( \15285 , \15047 , \15267 );
or \U$15092 ( \15286 , \15283 , \15284 , \15285 );
and \U$15093 ( \15287 , \15056 , \15060 );
and \U$15094 ( \15288 , \15060 , \15065 );
and \U$15095 ( \15289 , \15056 , \15065 );
or \U$15096 ( \15290 , \15287 , \15288 , \15289 );
and \U$15097 ( \15291 , \15070 , \15111 );
and \U$15098 ( \15292 , \15111 , \15235 );
and \U$15099 ( \15293 , \15070 , \15235 );
or \U$15100 ( \15294 , \15291 , \15292 , \15293 );
xor \U$15101 ( \15295 , \15290 , \15294 );
and \U$15102 ( \15296 , \15251 , \15265 );
xor \U$15103 ( \15297 , \15295 , \15296 );
xor \U$15104 ( \15298 , \15286 , \15297 );
and \U$15105 ( \15299 , \15035 , \15039 );
and \U$15106 ( \15300 , \15039 , \15041 );
and \U$15107 ( \15301 , \15035 , \15041 );
or \U$15108 ( \15302 , \15299 , \15300 , \15301 );
and \U$15109 ( \15303 , \15066 , \15236 );
and \U$15110 ( \15304 , \15236 , \15266 );
and \U$15111 ( \15305 , \15066 , \15266 );
or \U$15112 ( \15306 , \15303 , \15304 , \15305 );
xor \U$15113 ( \15307 , \15302 , \15306 );
and \U$15114 ( \15308 , \15241 , \15245 );
and \U$15115 ( \15309 , \15245 , \15250 );
and \U$15116 ( \15310 , \15241 , \15250 );
or \U$15117 ( \15311 , \15308 , \15309 , \15310 );
and \U$15118 ( \15312 , \15255 , \15259 );
and \U$15119 ( \15313 , \15259 , \15264 );
and \U$15120 ( \15314 , \15255 , \15264 );
or \U$15121 ( \15315 , \15312 , \15313 , \15314 );
xor \U$15122 ( \15316 , \15311 , \15315 );
and \U$15123 ( \15317 , \15156 , \15197 );
and \U$15124 ( \15318 , \15197 , \15234 );
and \U$15125 ( \15319 , \15156 , \15234 );
or \U$15126 ( \15320 , \15317 , \15318 , \15319 );
xor \U$15127 ( \15321 , \15316 , \15320 );
and \U$15128 ( \15322 , \15081 , \15095 );
and \U$15129 ( \15323 , \15095 , \15110 );
and \U$15130 ( \15324 , \15081 , \15110 );
or \U$15131 ( \15325 , \15322 , \15323 , \15324 );
and \U$15132 ( \15326 , \15160 , \15164 );
and \U$15133 ( \15327 , \15164 , \15169 );
and \U$15134 ( \15328 , \15160 , \15169 );
or \U$15135 ( \15329 , \15326 , \15327 , \15328 );
and \U$15136 ( \15330 , \15171 , \15175 );
and \U$15137 ( \15331 , \15175 , \15180 );
and \U$15138 ( \15332 , \15171 , \15180 );
or \U$15139 ( \15333 , \15330 , \15331 , \15332 );
xor \U$15140 ( \15334 , \15329 , \15333 );
and \U$15141 ( \15335 , \15186 , \15190 );
and \U$15142 ( \15336 , \15190 , \15195 );
and \U$15143 ( \15337 , \15186 , \15195 );
or \U$15144 ( \15338 , \15335 , \15336 , \15337 );
xor \U$15145 ( \15339 , \15334 , \15338 );
and \U$15146 ( \15340 , \15202 , \15206 );
and \U$15147 ( \15341 , \15206 , \15211 );
and \U$15148 ( \15342 , \15202 , \15211 );
or \U$15149 ( \15343 , \15340 , \15341 , \15342 );
and \U$15150 ( \15344 , \15216 , \15220 );
and \U$15151 ( \15345 , \15220 , \15225 );
and \U$15152 ( \15346 , \15216 , \15225 );
or \U$15153 ( \15347 , \15344 , \15345 , \15346 );
xor \U$15154 ( \15348 , \15343 , \15347 );
and \U$15155 ( \15349 , \15231 , \15232 );
xor \U$15156 ( \15350 , \15348 , \15349 );
xor \U$15157 ( \15351 , \15339 , \15350 );
and \U$15158 ( \15352 , \15116 , \15120 );
and \U$15159 ( \15353 , \15120 , \15125 );
and \U$15160 ( \15354 , \15116 , \15125 );
or \U$15161 ( \15355 , \15352 , \15353 , \15354 );
and \U$15162 ( \15356 , \15130 , \15134 );
and \U$15163 ( \15357 , \15134 , \15139 );
and \U$15164 ( \15358 , \15130 , \15139 );
or \U$15165 ( \15359 , \15356 , \15357 , \15358 );
xor \U$15166 ( \15360 , \15355 , \15359 );
and \U$15167 ( \15361 , \15145 , \15149 );
and \U$15168 ( \15362 , \15149 , \15154 );
and \U$15169 ( \15363 , \15145 , \15154 );
or \U$15170 ( \15364 , \15361 , \15362 , \15363 );
xor \U$15171 ( \15365 , \15360 , \15364 );
xor \U$15172 ( \15366 , \15351 , \15365 );
xor \U$15173 ( \15367 , \15325 , \15366 );
and \U$15174 ( \15368 , \4160 , \4581 );
and \U$15175 ( \15369 , \4364 , \4424 );
nor \U$15176 ( \15370 , \15368 , \15369 );
xnor \U$15177 ( \15371 , \15370 , \4377 );
and \U$15178 ( \15372 , \3736 , \5011 );
and \U$15179 ( \15373 , \3912 , \4878 );
nor \U$15180 ( \15374 , \15372 , \15373 );
xnor \U$15181 ( \15375 , \15374 , \4762 );
xor \U$15182 ( \15376 , \15371 , \15375 );
and \U$15183 ( \15377 , \3395 , \5485 );
and \U$15184 ( \15378 , \3646 , \5275 );
nor \U$15185 ( \15379 , \15377 , \15378 );
xnor \U$15186 ( \15380 , \15379 , \5169 );
xor \U$15187 ( \15381 , \15376 , \15380 );
and \U$15188 ( \15382 , \5469 , \3357 );
and \U$15189 ( \15383 , \5674 , \3255 );
nor \U$15190 ( \15384 , \15382 , \15383 );
xnor \U$15191 ( \15385 , \15384 , \3156 );
and \U$15192 ( \15386 , \4922 , \3813 );
and \U$15193 ( \15387 , \5156 , \3557 );
nor \U$15194 ( \15388 , \15386 , \15387 );
xnor \U$15195 ( \15389 , \15388 , \3562 );
xor \U$15196 ( \15390 , \15385 , \15389 );
and \U$15197 ( \15391 , \4654 , \4132 );
and \U$15198 ( \15392 , \4749 , \4012 );
nor \U$15199 ( \15393 , \15391 , \15392 );
xnor \U$15200 ( \15394 , \15393 , \3925 );
xor \U$15201 ( \15395 , \15390 , \15394 );
xor \U$15202 ( \15396 , \15381 , \15395 );
and \U$15203 ( \15397 , \3037 , \5996 );
and \U$15204 ( \15398 , \3143 , \5695 );
nor \U$15205 ( \15399 , \15397 , \15398 );
xnor \U$15206 ( \15400 , \15399 , \5687 );
and \U$15207 ( \15401 , \2757 , \6401 );
and \U$15208 ( \15402 , \2826 , \6143 );
nor \U$15209 ( \15403 , \15401 , \15402 );
xnor \U$15210 ( \15404 , \15403 , \6148 );
xor \U$15211 ( \15405 , \15400 , \15404 );
and \U$15212 ( \15406 , \2366 , \7055 );
and \U$15213 ( \15407 , \2521 , \6675 );
nor \U$15214 ( \15408 , \15406 , \15407 );
xnor \U$15215 ( \15409 , \15408 , \6680 );
xor \U$15216 ( \15410 , \15405 , \15409 );
xor \U$15217 ( \15411 , \15396 , \15410 );
and \U$15218 ( \15412 , \8652 , \1578 );
and \U$15219 ( \15413 , \8835 , \1431 );
nor \U$15220 ( \15414 , \15412 , \15413 );
xnor \U$15221 ( \15415 , \15414 , \1436 );
and \U$15222 ( \15416 , \8057 , \1824 );
and \U$15223 ( \15417 , \8349 , \1739 );
nor \U$15224 ( \15418 , \15416 , \15417 );
xnor \U$15225 ( \15419 , \15418 , \1697 );
xor \U$15226 ( \15420 , \15415 , \15419 );
and \U$15227 ( \15421 , \7556 , \2121 );
and \U$15228 ( \15422 , \7700 , \2008 );
nor \U$15229 ( \15423 , \15421 , \15422 );
xnor \U$15230 ( \15424 , \15423 , \1961 );
xor \U$15231 ( \15425 , \15420 , \15424 );
and \U$15232 ( \15426 , \10584 , \438 );
not \U$15233 ( \15427 , \15426 );
xnor \U$15234 ( \15428 , \15427 , \320 );
and \U$15235 ( \15429 , \9897 , \1086 );
and \U$15236 ( \15430 , \10206 , \508 );
nor \U$15237 ( \15431 , \15429 , \15430 );
xnor \U$15238 ( \15432 , \15431 , \487 );
xor \U$15239 ( \15433 , \15428 , \15432 );
and \U$15240 ( \15434 , \9169 , \1301 );
and \U$15241 ( \15435 , \9465 , \1246 );
nor \U$15242 ( \15436 , \15434 , \15435 );
xnor \U$15243 ( \15437 , \15436 , \1205 );
xor \U$15244 ( \15438 , \15433 , \15437 );
xor \U$15245 ( \15439 , \15425 , \15438 );
and \U$15246 ( \15440 , \6945 , \2400 );
and \U$15247 ( \15441 , \7231 , \2246 );
nor \U$15248 ( \15442 , \15440 , \15441 );
xnor \U$15249 ( \15443 , \15442 , \2195 );
and \U$15250 ( \15444 , \6514 , \2669 );
and \U$15251 ( \15445 , \6790 , \2538 );
nor \U$15252 ( \15446 , \15444 , \15445 );
xnor \U$15253 ( \15447 , \15446 , \2534 );
xor \U$15254 ( \15448 , \15443 , \15447 );
and \U$15255 ( \15449 , \6030 , \3103 );
and \U$15256 ( \15450 , \6281 , \2934 );
nor \U$15257 ( \15451 , \15449 , \15450 );
xnor \U$15258 ( \15452 , \15451 , \2839 );
xor \U$15259 ( \15453 , \15448 , \15452 );
xor \U$15260 ( \15454 , \15439 , \15453 );
xor \U$15261 ( \15455 , \15411 , \15454 );
and \U$15262 ( \15456 , \2090 , \7489 );
and \U$15263 ( \15457 , \2182 , \7137 );
nor \U$15264 ( \15458 , \15456 , \15457 );
xnor \U$15265 ( \15459 , \15458 , \7142 );
and \U$15266 ( \15460 , \1802 , \8019 );
and \U$15267 ( \15461 , \1948 , \7830 );
nor \U$15268 ( \15462 , \15460 , \15461 );
xnor \U$15269 ( \15463 , \15462 , \7713 );
xor \U$15270 ( \15464 , \15459 , \15463 );
and \U$15271 ( \15465 , \1601 , \8540 );
and \U$15272 ( \15466 , \1684 , \8292 );
nor \U$15273 ( \15467 , \15465 , \15466 );
xnor \U$15274 ( \15468 , \15467 , \8297 );
xor \U$15275 ( \15469 , \15464 , \15468 );
and \U$15276 ( \15470 , \1333 , \9333 );
and \U$15277 ( \15471 , \1484 , \9006 );
nor \U$15278 ( \15472 , \15470 , \15471 );
xnor \U$15279 ( \15473 , \15472 , \8848 );
and \U$15280 ( \15474 , \1147 , \9765 );
and \U$15281 ( \15475 , \1192 , \9644 );
nor \U$15282 ( \15476 , \15474 , \15475 );
xnor \U$15283 ( \15477 , \15476 , \9478 );
xor \U$15284 ( \15478 , \15473 , \15477 );
and \U$15285 ( \15479 , \412 , \10408 );
and \U$15286 ( \15480 , \474 , \10116 );
nor \U$15287 ( \15481 , \15479 , \15480 );
xnor \U$15288 ( \15482 , \15481 , \10121 );
xor \U$15289 ( \15483 , \15478 , \15482 );
xor \U$15290 ( \15484 , \15469 , \15483 );
and \U$15291 ( \15485 , \307 , \10118 );
not \U$15292 ( \15486 , \15485 );
xor \U$15293 ( \15487 , \15484 , \15486 );
xor \U$15294 ( \15488 , \15455 , \15487 );
xor \U$15295 ( \15489 , \15367 , \15488 );
xor \U$15296 ( \15490 , \15321 , \15489 );
and \U$15297 ( \15491 , \15126 , \15140 );
and \U$15298 ( \15492 , \15140 , \15155 );
and \U$15299 ( \15493 , \15126 , \15155 );
or \U$15300 ( \15494 , \15491 , \15492 , \15493 );
and \U$15301 ( \15495 , \15170 , \15181 );
and \U$15302 ( \15496 , \15181 , \15196 );
and \U$15303 ( \15497 , \15170 , \15196 );
or \U$15304 ( \15498 , \15495 , \15496 , \15497 );
xor \U$15305 ( \15499 , \15494 , \15498 );
and \U$15306 ( \15500 , \15212 , \15226 );
and \U$15307 ( \15501 , \15226 , \15233 );
and \U$15308 ( \15502 , \15212 , \15233 );
or \U$15309 ( \15503 , \15500 , \15501 , \15502 );
xor \U$15310 ( \15504 , \15499 , \15503 );
and \U$15311 ( \15505 , \15074 , \15078 );
and \U$15312 ( \15506 , \15078 , \15080 );
and \U$15313 ( \15507 , \15074 , \15080 );
or \U$15314 ( \15508 , \15505 , \15506 , \15507 );
and \U$15315 ( \15509 , \15085 , \15089 );
and \U$15316 ( \15510 , \15089 , \15094 );
and \U$15317 ( \15511 , \15085 , \15094 );
or \U$15318 ( \15512 , \15509 , \15510 , \15511 );
xor \U$15319 ( \15513 , \15508 , \15512 );
and \U$15320 ( \15514 , \15100 , \15104 );
and \U$15321 ( \15515 , \15104 , \15109 );
and \U$15322 ( \15516 , \15100 , \15109 );
or \U$15323 ( \15517 , \15514 , \15515 , \15516 );
xor \U$15324 ( \15518 , \15513 , \15517 );
xor \U$15325 ( \15519 , \15504 , \15518 );
xor \U$15326 ( \15520 , \15490 , \15519 );
xor \U$15327 ( \15521 , \15307 , \15520 );
xor \U$15328 ( \15522 , \15298 , \15521 );
xor \U$15329 ( \15523 , \15282 , \15522 );
and \U$15330 ( \15524 , \15027 , \15269 );
xor \U$15331 ( \15525 , \15523 , \15524 );
and \U$15332 ( \15526 , \15270 , \15271 );
and \U$15333 ( \15527 , \15272 , \15275 );
or \U$15334 ( \15528 , \15526 , \15527 );
xor \U$15335 ( \15529 , \15525 , \15528 );
buf g54fb_GF_PartitionCandidate( \15530_nG54fb , \15529 );
buf \U$15336 ( \15531 , \15530_nG54fb );
and \U$15337 ( \15532 , \15286 , \15297 );
and \U$15338 ( \15533 , \15297 , \15521 );
and \U$15339 ( \15534 , \15286 , \15521 );
or \U$15340 ( \15535 , \15532 , \15533 , \15534 );
and \U$15341 ( \15536 , \15302 , \15306 );
and \U$15342 ( \15537 , \15306 , \15520 );
and \U$15343 ( \15538 , \15302 , \15520 );
or \U$15344 ( \15539 , \15536 , \15537 , \15538 );
and \U$15345 ( \15540 , \15311 , \15315 );
and \U$15346 ( \15541 , \15315 , \15320 );
and \U$15347 ( \15542 , \15311 , \15320 );
or \U$15348 ( \15543 , \15540 , \15541 , \15542 );
and \U$15349 ( \15544 , \15325 , \15366 );
and \U$15350 ( \15545 , \15366 , \15488 );
and \U$15351 ( \15546 , \15325 , \15488 );
or \U$15352 ( \15547 , \15544 , \15545 , \15546 );
xor \U$15353 ( \15548 , \15543 , \15547 );
and \U$15354 ( \15549 , \15504 , \15518 );
xor \U$15355 ( \15550 , \15548 , \15549 );
xor \U$15356 ( \15551 , \15539 , \15550 );
and \U$15357 ( \15552 , \15290 , \15294 );
and \U$15358 ( \15553 , \15294 , \15296 );
and \U$15359 ( \15554 , \15290 , \15296 );
or \U$15360 ( \15555 , \15552 , \15553 , \15554 );
and \U$15361 ( \15556 , \15321 , \15489 );
and \U$15362 ( \15557 , \15489 , \15519 );
and \U$15363 ( \15558 , \15321 , \15519 );
or \U$15364 ( \15559 , \15556 , \15557 , \15558 );
xor \U$15365 ( \15560 , \15555 , \15559 );
and \U$15366 ( \15561 , \15494 , \15498 );
and \U$15367 ( \15562 , \15498 , \15503 );
and \U$15368 ( \15563 , \15494 , \15503 );
or \U$15369 ( \15564 , \15561 , \15562 , \15563 );
and \U$15370 ( \15565 , \15508 , \15512 );
and \U$15371 ( \15566 , \15512 , \15517 );
and \U$15372 ( \15567 , \15508 , \15517 );
or \U$15373 ( \15568 , \15565 , \15566 , \15567 );
xor \U$15374 ( \15569 , \15564 , \15568 );
and \U$15375 ( \15570 , \15411 , \15454 );
and \U$15376 ( \15571 , \15454 , \15487 );
and \U$15377 ( \15572 , \15411 , \15487 );
or \U$15378 ( \15573 , \15570 , \15571 , \15572 );
xor \U$15379 ( \15574 , \15569 , \15573 );
and \U$15380 ( \15575 , \15339 , \15350 );
and \U$15381 ( \15576 , \15350 , \15365 );
and \U$15382 ( \15577 , \15339 , \15365 );
or \U$15383 ( \15578 , \15575 , \15576 , \15577 );
and \U$15384 ( \15579 , \15459 , \15463 );
and \U$15385 ( \15580 , \15463 , \15468 );
and \U$15386 ( \15581 , \15459 , \15468 );
or \U$15387 ( \15582 , \15579 , \15580 , \15581 );
and \U$15388 ( \15583 , \15473 , \15477 );
and \U$15389 ( \15584 , \15477 , \15482 );
and \U$15390 ( \15585 , \15473 , \15482 );
or \U$15391 ( \15586 , \15583 , \15584 , \15585 );
xor \U$15392 ( \15587 , \15582 , \15586 );
buf \U$15393 ( \15588 , \15485 );
xor \U$15394 ( \15589 , \15587 , \15588 );
and \U$15395 ( \15590 , \15371 , \15375 );
and \U$15396 ( \15591 , \15375 , \15380 );
and \U$15397 ( \15592 , \15371 , \15380 );
or \U$15398 ( \15593 , \15590 , \15591 , \15592 );
and \U$15399 ( \15594 , \15385 , \15389 );
and \U$15400 ( \15595 , \15389 , \15394 );
and \U$15401 ( \15596 , \15385 , \15394 );
or \U$15402 ( \15597 , \15594 , \15595 , \15596 );
xor \U$15403 ( \15598 , \15593 , \15597 );
and \U$15404 ( \15599 , \15400 , \15404 );
and \U$15405 ( \15600 , \15404 , \15409 );
and \U$15406 ( \15601 , \15400 , \15409 );
or \U$15407 ( \15602 , \15599 , \15600 , \15601 );
xor \U$15408 ( \15603 , \15598 , \15602 );
xor \U$15409 ( \15604 , \15589 , \15603 );
and \U$15410 ( \15605 , \15415 , \15419 );
and \U$15411 ( \15606 , \15419 , \15424 );
and \U$15412 ( \15607 , \15415 , \15424 );
or \U$15413 ( \15608 , \15605 , \15606 , \15607 );
and \U$15414 ( \15609 , \15428 , \15432 );
and \U$15415 ( \15610 , \15432 , \15437 );
and \U$15416 ( \15611 , \15428 , \15437 );
or \U$15417 ( \15612 , \15609 , \15610 , \15611 );
xor \U$15418 ( \15613 , \15608 , \15612 );
and \U$15419 ( \15614 , \15443 , \15447 );
and \U$15420 ( \15615 , \15447 , \15452 );
and \U$15421 ( \15616 , \15443 , \15452 );
or \U$15422 ( \15617 , \15614 , \15615 , \15616 );
xor \U$15423 ( \15618 , \15613 , \15617 );
xor \U$15424 ( \15619 , \15604 , \15618 );
xor \U$15425 ( \15620 , \15578 , \15619 );
and \U$15426 ( \15621 , \8835 , \1578 );
and \U$15427 ( \15622 , \9169 , \1431 );
nor \U$15428 ( \15623 , \15621 , \15622 );
xnor \U$15429 ( \15624 , \15623 , \1436 );
and \U$15430 ( \15625 , \8349 , \1824 );
and \U$15431 ( \15626 , \8652 , \1739 );
nor \U$15432 ( \15627 , \15625 , \15626 );
xnor \U$15433 ( \15628 , \15627 , \1697 );
xor \U$15434 ( \15629 , \15624 , \15628 );
and \U$15435 ( \15630 , \7700 , \2121 );
and \U$15436 ( \15631 , \8057 , \2008 );
nor \U$15437 ( \15632 , \15630 , \15631 );
xnor \U$15438 ( \15633 , \15632 , \1961 );
xor \U$15439 ( \15634 , \15629 , \15633 );
not \U$15440 ( \15635 , \320 );
and \U$15441 ( \15636 , \10206 , \1086 );
and \U$15442 ( \15637 , \10584 , \508 );
nor \U$15443 ( \15638 , \15636 , \15637 );
xnor \U$15444 ( \15639 , \15638 , \487 );
xor \U$15445 ( \15640 , \15635 , \15639 );
and \U$15446 ( \15641 , \9465 , \1301 );
and \U$15447 ( \15642 , \9897 , \1246 );
nor \U$15448 ( \15643 , \15641 , \15642 );
xnor \U$15449 ( \15644 , \15643 , \1205 );
xor \U$15450 ( \15645 , \15640 , \15644 );
xor \U$15451 ( \15646 , \15634 , \15645 );
and \U$15452 ( \15647 , \7231 , \2400 );
and \U$15453 ( \15648 , \7556 , \2246 );
nor \U$15454 ( \15649 , \15647 , \15648 );
xnor \U$15455 ( \15650 , \15649 , \2195 );
and \U$15456 ( \15651 , \6790 , \2669 );
and \U$15457 ( \15652 , \6945 , \2538 );
nor \U$15458 ( \15653 , \15651 , \15652 );
xnor \U$15459 ( \15654 , \15653 , \2534 );
xor \U$15460 ( \15655 , \15650 , \15654 );
and \U$15461 ( \15656 , \6281 , \3103 );
and \U$15462 ( \15657 , \6514 , \2934 );
nor \U$15463 ( \15658 , \15656 , \15657 );
xnor \U$15464 ( \15659 , \15658 , \2839 );
xor \U$15465 ( \15660 , \15655 , \15659 );
xor \U$15466 ( \15661 , \15646 , \15660 );
and \U$15467 ( \15662 , \3143 , \5996 );
and \U$15468 ( \15663 , \3395 , \5695 );
nor \U$15469 ( \15664 , \15662 , \15663 );
xnor \U$15470 ( \15665 , \15664 , \5687 );
and \U$15471 ( \15666 , \2826 , \6401 );
and \U$15472 ( \15667 , \3037 , \6143 );
nor \U$15473 ( \15668 , \15666 , \15667 );
xnor \U$15474 ( \15669 , \15668 , \6148 );
xor \U$15475 ( \15670 , \15665 , \15669 );
and \U$15476 ( \15671 , \2521 , \7055 );
and \U$15477 ( \15672 , \2757 , \6675 );
nor \U$15478 ( \15673 , \15671 , \15672 );
xnor \U$15479 ( \15674 , \15673 , \6680 );
xor \U$15480 ( \15675 , \15670 , \15674 );
and \U$15481 ( \15676 , \4364 , \4581 );
and \U$15482 ( \15677 , \4654 , \4424 );
nor \U$15483 ( \15678 , \15676 , \15677 );
xnor \U$15484 ( \15679 , \15678 , \4377 );
and \U$15485 ( \15680 , \3912 , \5011 );
and \U$15486 ( \15681 , \4160 , \4878 );
nor \U$15487 ( \15682 , \15680 , \15681 );
xnor \U$15488 ( \15683 , \15682 , \4762 );
xor \U$15489 ( \15684 , \15679 , \15683 );
and \U$15490 ( \15685 , \3646 , \5485 );
and \U$15491 ( \15686 , \3736 , \5275 );
nor \U$15492 ( \15687 , \15685 , \15686 );
xnor \U$15493 ( \15688 , \15687 , \5169 );
xor \U$15494 ( \15689 , \15684 , \15688 );
xor \U$15495 ( \15690 , \15675 , \15689 );
and \U$15496 ( \15691 , \5674 , \3357 );
and \U$15497 ( \15692 , \6030 , \3255 );
nor \U$15498 ( \15693 , \15691 , \15692 );
xnor \U$15499 ( \15694 , \15693 , \3156 );
and \U$15500 ( \15695 , \5156 , \3813 );
and \U$15501 ( \15696 , \5469 , \3557 );
nor \U$15502 ( \15697 , \15695 , \15696 );
xnor \U$15503 ( \15698 , \15697 , \3562 );
xor \U$15504 ( \15699 , \15694 , \15698 );
and \U$15505 ( \15700 , \4749 , \4132 );
and \U$15506 ( \15701 , \4922 , \4012 );
nor \U$15507 ( \15702 , \15700 , \15701 );
xnor \U$15508 ( \15703 , \15702 , \3925 );
xor \U$15509 ( \15704 , \15699 , \15703 );
xor \U$15510 ( \15705 , \15690 , \15704 );
xor \U$15511 ( \15706 , \15661 , \15705 );
and \U$15512 ( \15707 , \412 , \10118 );
and \U$15513 ( \15708 , \2182 , \7489 );
and \U$15514 ( \15709 , \2366 , \7137 );
nor \U$15515 ( \15710 , \15708 , \15709 );
xnor \U$15516 ( \15711 , \15710 , \7142 );
and \U$15517 ( \15712 , \1948 , \8019 );
and \U$15518 ( \15713 , \2090 , \7830 );
nor \U$15519 ( \15714 , \15712 , \15713 );
xnor \U$15520 ( \15715 , \15714 , \7713 );
xor \U$15521 ( \15716 , \15711 , \15715 );
and \U$15522 ( \15717 , \1684 , \8540 );
and \U$15523 ( \15718 , \1802 , \8292 );
nor \U$15524 ( \15719 , \15717 , \15718 );
xnor \U$15525 ( \15720 , \15719 , \8297 );
xor \U$15526 ( \15721 , \15716 , \15720 );
xor \U$15527 ( \15722 , \15707 , \15721 );
and \U$15528 ( \15723 , \1484 , \9333 );
and \U$15529 ( \15724 , \1601 , \9006 );
nor \U$15530 ( \15725 , \15723 , \15724 );
xnor \U$15531 ( \15726 , \15725 , \8848 );
and \U$15532 ( \15727 , \1192 , \9765 );
and \U$15533 ( \15728 , \1333 , \9644 );
nor \U$15534 ( \15729 , \15727 , \15728 );
xnor \U$15535 ( \15730 , \15729 , \9478 );
xor \U$15536 ( \15731 , \15726 , \15730 );
and \U$15537 ( \15732 , \474 , \10408 );
and \U$15538 ( \15733 , \1147 , \10116 );
nor \U$15539 ( \15734 , \15732 , \15733 );
xnor \U$15540 ( \15735 , \15734 , \10121 );
xor \U$15541 ( \15736 , \15731 , \15735 );
xor \U$15542 ( \15737 , \15722 , \15736 );
xor \U$15543 ( \15738 , \15706 , \15737 );
xor \U$15544 ( \15739 , \15620 , \15738 );
xor \U$15545 ( \15740 , \15574 , \15739 );
and \U$15546 ( \15741 , \15381 , \15395 );
and \U$15547 ( \15742 , \15395 , \15410 );
and \U$15548 ( \15743 , \15381 , \15410 );
or \U$15549 ( \15744 , \15741 , \15742 , \15743 );
and \U$15550 ( \15745 , \15425 , \15438 );
and \U$15551 ( \15746 , \15438 , \15453 );
and \U$15552 ( \15747 , \15425 , \15453 );
or \U$15553 ( \15748 , \15745 , \15746 , \15747 );
xor \U$15554 ( \15749 , \15744 , \15748 );
and \U$15555 ( \15750 , \15469 , \15483 );
and \U$15556 ( \15751 , \15483 , \15486 );
and \U$15557 ( \15752 , \15469 , \15486 );
or \U$15558 ( \15753 , \15750 , \15751 , \15752 );
xor \U$15559 ( \15754 , \15749 , \15753 );
and \U$15560 ( \15755 , \15329 , \15333 );
and \U$15561 ( \15756 , \15333 , \15338 );
and \U$15562 ( \15757 , \15329 , \15338 );
or \U$15563 ( \15758 , \15755 , \15756 , \15757 );
and \U$15564 ( \15759 , \15343 , \15347 );
and \U$15565 ( \15760 , \15347 , \15349 );
and \U$15566 ( \15761 , \15343 , \15349 );
or \U$15567 ( \15762 , \15759 , \15760 , \15761 );
xor \U$15568 ( \15763 , \15758 , \15762 );
and \U$15569 ( \15764 , \15355 , \15359 );
and \U$15570 ( \15765 , \15359 , \15364 );
and \U$15571 ( \15766 , \15355 , \15364 );
or \U$15572 ( \15767 , \15764 , \15765 , \15766 );
xor \U$15573 ( \15768 , \15763 , \15767 );
xor \U$15574 ( \15769 , \15754 , \15768 );
xor \U$15575 ( \15770 , \15740 , \15769 );
xor \U$15576 ( \15771 , \15560 , \15770 );
xor \U$15577 ( \15772 , \15551 , \15771 );
xor \U$15578 ( \15773 , \15535 , \15772 );
and \U$15579 ( \15774 , \15282 , \15522 );
xor \U$15580 ( \15775 , \15773 , \15774 );
and \U$15581 ( \15776 , \15523 , \15524 );
and \U$15582 ( \15777 , \15525 , \15528 );
or \U$15583 ( \15778 , \15776 , \15777 );
xor \U$15584 ( \15779 , \15775 , \15778 );
buf g54f9_GF_PartitionCandidate( \15780_nG54f9 , \15779 );
buf \U$15585 ( \15781 , \15780_nG54f9 );
or \U$15586 ( \15782 , \1070 , \1171 , \1279 , \1390 , \1508 , \1629 , \1757 , \1888 , \2026 , \2167 , \2315 , \2466 , \2624 , \2785 , \2953 , \3124 , \3302 , \3483 , \3671 , \3862 , \4060 , \4261 , \4469 , \4680 , \4898 , \5118 , \5349 , \5580 , \5818 , \6059 , \6307 , \6558 , \6816 , \7077 , \7345 , \7616 , \7894 , \8175 , \8463 , \8754 , \9052 , \9353 , \9661 , \9972 , \10290 , \10611 , \10930 , \11248 , \11565 , \11881 , \12192 , \12500 , \12803 , \13099 , \13390 , \13673 , \13954 , \14227 , \14497 , \14763 , \15023 , \15278 , \15531 , \15781 );
and \U$15587 ( \15783 , \15539 , \15550 );
and \U$15588 ( \15784 , \15550 , \15771 );
and \U$15589 ( \15785 , \15539 , \15771 );
or \U$15590 ( \15786 , \15783 , \15784 , \15785 );
and \U$15591 ( \15787 , \15555 , \15559 );
and \U$15592 ( \15788 , \15559 , \15770 );
and \U$15593 ( \15789 , \15555 , \15770 );
or \U$15594 ( \15790 , \15787 , \15788 , \15789 );
and \U$15595 ( \15791 , \15564 , \15568 );
and \U$15596 ( \15792 , \15568 , \15573 );
and \U$15597 ( \15793 , \15564 , \15573 );
or \U$15598 ( \15794 , \15791 , \15792 , \15793 );
and \U$15599 ( \15795 , \15578 , \15619 );
and \U$15600 ( \15796 , \15619 , \15738 );
and \U$15601 ( \15797 , \15578 , \15738 );
or \U$15602 ( \15798 , \15795 , \15796 , \15797 );
xor \U$15603 ( \15799 , \15794 , \15798 );
and \U$15604 ( \15800 , \15754 , \15768 );
xor \U$15605 ( \15801 , \15799 , \15800 );
xor \U$15606 ( \15802 , \15790 , \15801 );
and \U$15607 ( \15803 , \15543 , \15547 );
and \U$15608 ( \15804 , \15547 , \15549 );
and \U$15609 ( \15805 , \15543 , \15549 );
or \U$15610 ( \15806 , \15803 , \15804 , \15805 );
and \U$15611 ( \15807 , \15574 , \15739 );
and \U$15612 ( \15808 , \15739 , \15769 );
and \U$15613 ( \15809 , \15574 , \15769 );
or \U$15614 ( \15810 , \15807 , \15808 , \15809 );
xor \U$15615 ( \15811 , \15806 , \15810 );
and \U$15616 ( \15812 , \15744 , \15748 );
and \U$15617 ( \15813 , \15748 , \15753 );
and \U$15618 ( \15814 , \15744 , \15753 );
or \U$15619 ( \15815 , \15812 , \15813 , \15814 );
and \U$15620 ( \15816 , \15758 , \15762 );
and \U$15621 ( \15817 , \15762 , \15767 );
and \U$15622 ( \15818 , \15758 , \15767 );
or \U$15623 ( \15819 , \15816 , \15817 , \15818 );
xor \U$15624 ( \15820 , \15815 , \15819 );
and \U$15625 ( \15821 , \15661 , \15705 );
and \U$15626 ( \15822 , \15705 , \15737 );
and \U$15627 ( \15823 , \15661 , \15737 );
or \U$15628 ( \15824 , \15821 , \15822 , \15823 );
xor \U$15629 ( \15825 , \15820 , \15824 );
and \U$15630 ( \15826 , \15589 , \15603 );
and \U$15631 ( \15827 , \15603 , \15618 );
and \U$15632 ( \15828 , \15589 , \15618 );
or \U$15633 ( \15829 , \15826 , \15827 , \15828 );
and \U$15634 ( \15830 , \15624 , \15628 );
and \U$15635 ( \15831 , \15628 , \15633 );
and \U$15636 ( \15832 , \15624 , \15633 );
or \U$15637 ( \15833 , \15830 , \15831 , \15832 );
and \U$15638 ( \15834 , \15635 , \15639 );
and \U$15639 ( \15835 , \15639 , \15644 );
and \U$15640 ( \15836 , \15635 , \15644 );
or \U$15641 ( \15837 , \15834 , \15835 , \15836 );
xor \U$15642 ( \15838 , \15833 , \15837 );
and \U$15643 ( \15839 , \15650 , \15654 );
and \U$15644 ( \15840 , \15654 , \15659 );
and \U$15645 ( \15841 , \15650 , \15659 );
or \U$15646 ( \15842 , \15839 , \15840 , \15841 );
xor \U$15647 ( \15843 , \15838 , \15842 );
and \U$15648 ( \15844 , \15665 , \15669 );
and \U$15649 ( \15845 , \15669 , \15674 );
and \U$15650 ( \15846 , \15665 , \15674 );
or \U$15651 ( \15847 , \15844 , \15845 , \15846 );
and \U$15652 ( \15848 , \15679 , \15683 );
and \U$15653 ( \15849 , \15683 , \15688 );
and \U$15654 ( \15850 , \15679 , \15688 );
or \U$15655 ( \15851 , \15848 , \15849 , \15850 );
xor \U$15656 ( \15852 , \15847 , \15851 );
and \U$15657 ( \15853 , \15694 , \15698 );
and \U$15658 ( \15854 , \15698 , \15703 );
and \U$15659 ( \15855 , \15694 , \15703 );
or \U$15660 ( \15856 , \15853 , \15854 , \15855 );
xor \U$15661 ( \15857 , \15852 , \15856 );
xor \U$15662 ( \15858 , \15843 , \15857 );
and \U$15663 ( \15859 , \15711 , \15715 );
and \U$15664 ( \15860 , \15715 , \15720 );
and \U$15665 ( \15861 , \15711 , \15720 );
or \U$15666 ( \15862 , \15859 , \15860 , \15861 );
and \U$15667 ( \15863 , \15726 , \15730 );
and \U$15668 ( \15864 , \15730 , \15735 );
and \U$15669 ( \15865 , \15726 , \15735 );
or \U$15670 ( \15866 , \15863 , \15864 , \15865 );
xnor \U$15671 ( \15867 , \15862 , \15866 );
xor \U$15672 ( \15868 , \15858 , \15867 );
xor \U$15673 ( \15869 , \15829 , \15868 );
and \U$15674 ( \15870 , \5469 , \3813 );
and \U$15675 ( \15871 , \5674 , \3557 );
nor \U$15676 ( \15872 , \15870 , \15871 );
xnor \U$15677 ( \15873 , \15872 , \3562 );
and \U$15678 ( \15874 , \4922 , \4132 );
and \U$15679 ( \15875 , \5156 , \4012 );
nor \U$15680 ( \15876 , \15874 , \15875 );
xnor \U$15681 ( \15877 , \15876 , \3925 );
xor \U$15682 ( \15878 , \15873 , \15877 );
and \U$15683 ( \15879 , \4654 , \4581 );
and \U$15684 ( \15880 , \4749 , \4424 );
nor \U$15685 ( \15881 , \15879 , \15880 );
xnor \U$15686 ( \15882 , \15881 , \4377 );
xor \U$15687 ( \15883 , \15878 , \15882 );
and \U$15688 ( \15884 , \4160 , \5011 );
and \U$15689 ( \15885 , \4364 , \4878 );
nor \U$15690 ( \15886 , \15884 , \15885 );
xnor \U$15691 ( \15887 , \15886 , \4762 );
and \U$15692 ( \15888 , \3736 , \5485 );
and \U$15693 ( \15889 , \3912 , \5275 );
nor \U$15694 ( \15890 , \15888 , \15889 );
xnor \U$15695 ( \15891 , \15890 , \5169 );
xor \U$15696 ( \15892 , \15887 , \15891 );
and \U$15697 ( \15893 , \3395 , \5996 );
and \U$15698 ( \15894 , \3646 , \5695 );
nor \U$15699 ( \15895 , \15893 , \15894 );
xnor \U$15700 ( \15896 , \15895 , \5687 );
xor \U$15701 ( \15897 , \15892 , \15896 );
xor \U$15702 ( \15898 , \15883 , \15897 );
and \U$15703 ( \15899 , \6945 , \2669 );
and \U$15704 ( \15900 , \7231 , \2538 );
nor \U$15705 ( \15901 , \15899 , \15900 );
xnor \U$15706 ( \15902 , \15901 , \2534 );
and \U$15707 ( \15903 , \6514 , \3103 );
and \U$15708 ( \15904 , \6790 , \2934 );
nor \U$15709 ( \15905 , \15903 , \15904 );
xnor \U$15710 ( \15906 , \15905 , \2839 );
xor \U$15711 ( \15907 , \15902 , \15906 );
and \U$15712 ( \15908 , \6030 , \3357 );
and \U$15713 ( \15909 , \6281 , \3255 );
nor \U$15714 ( \15910 , \15908 , \15909 );
xnor \U$15715 ( \15911 , \15910 , \3156 );
xor \U$15716 ( \15912 , \15907 , \15911 );
xor \U$15717 ( \15913 , \15898 , \15912 );
and \U$15718 ( \15914 , \3037 , \6401 );
and \U$15719 ( \15915 , \3143 , \6143 );
nor \U$15720 ( \15916 , \15914 , \15915 );
xnor \U$15721 ( \15917 , \15916 , \6148 );
and \U$15722 ( \15918 , \2757 , \7055 );
and \U$15723 ( \15919 , \2826 , \6675 );
nor \U$15724 ( \15920 , \15918 , \15919 );
xnor \U$15725 ( \15921 , \15920 , \6680 );
xor \U$15726 ( \15922 , \15917 , \15921 );
and \U$15727 ( \15923 , \2366 , \7489 );
and \U$15728 ( \15924 , \2521 , \7137 );
nor \U$15729 ( \15925 , \15923 , \15924 );
xnor \U$15730 ( \15926 , \15925 , \7142 );
xor \U$15731 ( \15927 , \15922 , \15926 );
and \U$15732 ( \15928 , \2090 , \8019 );
and \U$15733 ( \15929 , \2182 , \7830 );
nor \U$15734 ( \15930 , \15928 , \15929 );
xnor \U$15735 ( \15931 , \15930 , \7713 );
and \U$15736 ( \15932 , \1802 , \8540 );
and \U$15737 ( \15933 , \1948 , \8292 );
nor \U$15738 ( \15934 , \15932 , \15933 );
xnor \U$15739 ( \15935 , \15934 , \8297 );
xor \U$15740 ( \15936 , \15931 , \15935 );
and \U$15741 ( \15937 , \1601 , \9333 );
and \U$15742 ( \15938 , \1684 , \9006 );
nor \U$15743 ( \15939 , \15937 , \15938 );
xnor \U$15744 ( \15940 , \15939 , \8848 );
xor \U$15745 ( \15941 , \15936 , \15940 );
xor \U$15746 ( \15942 , \15927 , \15941 );
and \U$15747 ( \15943 , \1333 , \9765 );
and \U$15748 ( \15944 , \1484 , \9644 );
nor \U$15749 ( \15945 , \15943 , \15944 );
xnor \U$15750 ( \15946 , \15945 , \9478 );
and \U$15751 ( \15947 , \1147 , \10408 );
and \U$15752 ( \15948 , \1192 , \10116 );
nor \U$15753 ( \15949 , \15947 , \15948 );
xnor \U$15754 ( \15950 , \15949 , \10121 );
xor \U$15755 ( \15951 , \15946 , \15950 );
and \U$15756 ( \15952 , \474 , \10118 );
xor \U$15757 ( \15953 , \15951 , \15952 );
xor \U$15758 ( \15954 , \15942 , \15953 );
xor \U$15759 ( \15955 , \15913 , \15954 );
and \U$15760 ( \15956 , \10584 , \1086 );
not \U$15761 ( \15957 , \15956 );
xnor \U$15762 ( \15958 , \15957 , \487 );
and \U$15763 ( \15959 , \9897 , \1301 );
and \U$15764 ( \15960 , \10206 , \1246 );
nor \U$15765 ( \15961 , \15959 , \15960 );
xnor \U$15766 ( \15962 , \15961 , \1205 );
xor \U$15767 ( \15963 , \15958 , \15962 );
and \U$15768 ( \15964 , \9169 , \1578 );
and \U$15769 ( \15965 , \9465 , \1431 );
nor \U$15770 ( \15966 , \15964 , \15965 );
xnor \U$15771 ( \15967 , \15966 , \1436 );
xor \U$15772 ( \15968 , \15963 , \15967 );
and \U$15773 ( \15969 , \8652 , \1824 );
and \U$15774 ( \15970 , \8835 , \1739 );
nor \U$15775 ( \15971 , \15969 , \15970 );
xnor \U$15776 ( \15972 , \15971 , \1697 );
and \U$15777 ( \15973 , \8057 , \2121 );
and \U$15778 ( \15974 , \8349 , \2008 );
nor \U$15779 ( \15975 , \15973 , \15974 );
xnor \U$15780 ( \15976 , \15975 , \1961 );
xor \U$15781 ( \15977 , \15972 , \15976 );
and \U$15782 ( \15978 , \7556 , \2400 );
and \U$15783 ( \15979 , \7700 , \2246 );
nor \U$15784 ( \15980 , \15978 , \15979 );
xnor \U$15785 ( \15981 , \15980 , \2195 );
xor \U$15786 ( \15982 , \15977 , \15981 );
xor \U$15787 ( \15983 , \15968 , \15982 );
xor \U$15788 ( \15984 , \15955 , \15983 );
xor \U$15789 ( \15985 , \15869 , \15984 );
xor \U$15790 ( \15986 , \15825 , \15985 );
and \U$15791 ( \15987 , \15582 , \15586 );
and \U$15792 ( \15988 , \15586 , \15588 );
and \U$15793 ( \15989 , \15582 , \15588 );
or \U$15794 ( \15990 , \15987 , \15988 , \15989 );
and \U$15795 ( \15991 , \15593 , \15597 );
and \U$15796 ( \15992 , \15597 , \15602 );
and \U$15797 ( \15993 , \15593 , \15602 );
or \U$15798 ( \15994 , \15991 , \15992 , \15993 );
xor \U$15799 ( \15995 , \15990 , \15994 );
and \U$15800 ( \15996 , \15608 , \15612 );
and \U$15801 ( \15997 , \15612 , \15617 );
and \U$15802 ( \15998 , \15608 , \15617 );
or \U$15803 ( \15999 , \15996 , \15997 , \15998 );
xor \U$15804 ( \16000 , \15995 , \15999 );
and \U$15805 ( \16001 , \15634 , \15645 );
and \U$15806 ( \16002 , \15645 , \15660 );
and \U$15807 ( \16003 , \15634 , \15660 );
or \U$15808 ( \16004 , \16001 , \16002 , \16003 );
and \U$15809 ( \16005 , \15675 , \15689 );
and \U$15810 ( \16006 , \15689 , \15704 );
and \U$15811 ( \16007 , \15675 , \15704 );
or \U$15812 ( \16008 , \16005 , \16006 , \16007 );
xor \U$15813 ( \16009 , \16004 , \16008 );
and \U$15814 ( \16010 , \15707 , \15721 );
and \U$15815 ( \16011 , \15721 , \15736 );
and \U$15816 ( \16012 , \15707 , \15736 );
or \U$15817 ( \16013 , \16010 , \16011 , \16012 );
xor \U$15818 ( \16014 , \16009 , \16013 );
xor \U$15819 ( \16015 , \16000 , \16014 );
xor \U$15820 ( \16016 , \15986 , \16015 );
xor \U$15821 ( \16017 , \15811 , \16016 );
xor \U$15822 ( \16018 , \15802 , \16017 );
xor \U$15823 ( \16019 , \15786 , \16018 );
and \U$15824 ( \16020 , \15535 , \15772 );
xor \U$15825 ( \16021 , \16019 , \16020 );
and \U$15826 ( \16022 , \15773 , \15774 );
and \U$15827 ( \16023 , \15775 , \15778 );
or \U$15828 ( \16024 , \16022 , \16023 );
xor \U$15829 ( \16025 , \16021 , \16024 );
buf g54f7_GF_PartitionCandidate( \16026_nG54f7 , \16025 );
buf \U$15830 ( \16027 , \16026_nG54f7 );
and \U$15831 ( \16028 , \15790 , \15801 );
and \U$15832 ( \16029 , \15801 , \16017 );
and \U$15833 ( \16030 , \15790 , \16017 );
or \U$15834 ( \16031 , \16028 , \16029 , \16030 );
and \U$15835 ( \16032 , \15806 , \15810 );
and \U$15836 ( \16033 , \15810 , \16016 );
and \U$15837 ( \16034 , \15806 , \16016 );
or \U$15838 ( \16035 , \16032 , \16033 , \16034 );
and \U$15839 ( \16036 , \15815 , \15819 );
and \U$15840 ( \16037 , \15819 , \15824 );
and \U$15841 ( \16038 , \15815 , \15824 );
or \U$15842 ( \16039 , \16036 , \16037 , \16038 );
and \U$15843 ( \16040 , \15829 , \15868 );
and \U$15844 ( \16041 , \15868 , \15984 );
and \U$15845 ( \16042 , \15829 , \15984 );
or \U$15846 ( \16043 , \16040 , \16041 , \16042 );
xor \U$15847 ( \16044 , \16039 , \16043 );
and \U$15848 ( \16045 , \16000 , \16014 );
xor \U$15849 ( \16046 , \16044 , \16045 );
xor \U$15850 ( \16047 , \16035 , \16046 );
and \U$15851 ( \16048 , \15794 , \15798 );
and \U$15852 ( \16049 , \15798 , \15800 );
and \U$15853 ( \16050 , \15794 , \15800 );
or \U$15854 ( \16051 , \16048 , \16049 , \16050 );
and \U$15855 ( \16052 , \15825 , \15985 );
and \U$15856 ( \16053 , \15985 , \16015 );
and \U$15857 ( \16054 , \15825 , \16015 );
or \U$15858 ( \16055 , \16052 , \16053 , \16054 );
xor \U$15859 ( \16056 , \16051 , \16055 );
and \U$15860 ( \16057 , \15990 , \15994 );
and \U$15861 ( \16058 , \15994 , \15999 );
and \U$15862 ( \16059 , \15990 , \15999 );
or \U$15863 ( \16060 , \16057 , \16058 , \16059 );
and \U$15864 ( \16061 , \16004 , \16008 );
and \U$15865 ( \16062 , \16008 , \16013 );
and \U$15866 ( \16063 , \16004 , \16013 );
or \U$15867 ( \16064 , \16061 , \16062 , \16063 );
xor \U$15868 ( \16065 , \16060 , \16064 );
and \U$15869 ( \16066 , \15913 , \15954 );
and \U$15870 ( \16067 , \15954 , \15983 );
and \U$15871 ( \16068 , \15913 , \15983 );
or \U$15872 ( \16069 , \16066 , \16067 , \16068 );
xor \U$15873 ( \16070 , \16065 , \16069 );
and \U$15874 ( \16071 , \15843 , \15857 );
and \U$15875 ( \16072 , \15857 , \15867 );
and \U$15876 ( \16073 , \15843 , \15867 );
or \U$15877 ( \16074 , \16071 , \16072 , \16073 );
not \U$15878 ( \16075 , \487 );
and \U$15879 ( \16076 , \10206 , \1301 );
and \U$15880 ( \16077 , \10584 , \1246 );
nor \U$15881 ( \16078 , \16076 , \16077 );
xnor \U$15882 ( \16079 , \16078 , \1205 );
xor \U$15883 ( \16080 , \16075 , \16079 );
and \U$15884 ( \16081 , \9465 , \1578 );
and \U$15885 ( \16082 , \9897 , \1431 );
nor \U$15886 ( \16083 , \16081 , \16082 );
xnor \U$15887 ( \16084 , \16083 , \1436 );
xor \U$15888 ( \16085 , \16080 , \16084 );
and \U$15889 ( \16086 , \5674 , \3813 );
and \U$15890 ( \16087 , \6030 , \3557 );
nor \U$15891 ( \16088 , \16086 , \16087 );
xnor \U$15892 ( \16089 , \16088 , \3562 );
and \U$15893 ( \16090 , \5156 , \4132 );
and \U$15894 ( \16091 , \5469 , \4012 );
nor \U$15895 ( \16092 , \16090 , \16091 );
xnor \U$15896 ( \16093 , \16092 , \3925 );
xor \U$15897 ( \16094 , \16089 , \16093 );
and \U$15898 ( \16095 , \4749 , \4581 );
and \U$15899 ( \16096 , \4922 , \4424 );
nor \U$15900 ( \16097 , \16095 , \16096 );
xnor \U$15901 ( \16098 , \16097 , \4377 );
xor \U$15902 ( \16099 , \16094 , \16098 );
and \U$15903 ( \16100 , \8835 , \1824 );
and \U$15904 ( \16101 , \9169 , \1739 );
nor \U$15905 ( \16102 , \16100 , \16101 );
xnor \U$15906 ( \16103 , \16102 , \1697 );
and \U$15907 ( \16104 , \8349 , \2121 );
and \U$15908 ( \16105 , \8652 , \2008 );
nor \U$15909 ( \16106 , \16104 , \16105 );
xnor \U$15910 ( \16107 , \16106 , \1961 );
xor \U$15911 ( \16108 , \16103 , \16107 );
and \U$15912 ( \16109 , \7700 , \2400 );
and \U$15913 ( \16110 , \8057 , \2246 );
nor \U$15914 ( \16111 , \16109 , \16110 );
xnor \U$15915 ( \16112 , \16111 , \2195 );
xor \U$15916 ( \16113 , \16108 , \16112 );
xor \U$15917 ( \16114 , \16099 , \16113 );
and \U$15918 ( \16115 , \7231 , \2669 );
and \U$15919 ( \16116 , \7556 , \2538 );
nor \U$15920 ( \16117 , \16115 , \16116 );
xnor \U$15921 ( \16118 , \16117 , \2534 );
and \U$15922 ( \16119 , \6790 , \3103 );
and \U$15923 ( \16120 , \6945 , \2934 );
nor \U$15924 ( \16121 , \16119 , \16120 );
xnor \U$15925 ( \16122 , \16121 , \2839 );
xor \U$15926 ( \16123 , \16118 , \16122 );
and \U$15927 ( \16124 , \6281 , \3357 );
and \U$15928 ( \16125 , \6514 , \3255 );
nor \U$15929 ( \16126 , \16124 , \16125 );
xnor \U$15930 ( \16127 , \16126 , \3156 );
xor \U$15931 ( \16128 , \16123 , \16127 );
xor \U$15932 ( \16129 , \16114 , \16128 );
xor \U$15933 ( \16130 , \16085 , \16129 );
and \U$15934 ( \16131 , \4364 , \5011 );
and \U$15935 ( \16132 , \4654 , \4878 );
nor \U$15936 ( \16133 , \16131 , \16132 );
xnor \U$15937 ( \16134 , \16133 , \4762 );
and \U$15938 ( \16135 , \3912 , \5485 );
and \U$15939 ( \16136 , \4160 , \5275 );
nor \U$15940 ( \16137 , \16135 , \16136 );
xnor \U$15941 ( \16138 , \16137 , \5169 );
xor \U$15942 ( \16139 , \16134 , \16138 );
and \U$15943 ( \16140 , \3646 , \5996 );
and \U$15944 ( \16141 , \3736 , \5695 );
nor \U$15945 ( \16142 , \16140 , \16141 );
xnor \U$15946 ( \16143 , \16142 , \5687 );
xor \U$15947 ( \16144 , \16139 , \16143 );
and \U$15948 ( \16145 , \3143 , \6401 );
and \U$15949 ( \16146 , \3395 , \6143 );
nor \U$15950 ( \16147 , \16145 , \16146 );
xnor \U$15951 ( \16148 , \16147 , \6148 );
and \U$15952 ( \16149 , \2826 , \7055 );
and \U$15953 ( \16150 , \3037 , \6675 );
nor \U$15954 ( \16151 , \16149 , \16150 );
xnor \U$15955 ( \16152 , \16151 , \6680 );
xor \U$15956 ( \16153 , \16148 , \16152 );
and \U$15957 ( \16154 , \2521 , \7489 );
and \U$15958 ( \16155 , \2757 , \7137 );
nor \U$15959 ( \16156 , \16154 , \16155 );
xnor \U$15960 ( \16157 , \16156 , \7142 );
xor \U$15961 ( \16158 , \16153 , \16157 );
xor \U$15962 ( \16159 , \16144 , \16158 );
and \U$15963 ( \16160 , \2182 , \8019 );
and \U$15964 ( \16161 , \2366 , \7830 );
nor \U$15965 ( \16162 , \16160 , \16161 );
xnor \U$15966 ( \16163 , \16162 , \7713 );
and \U$15967 ( \16164 , \1948 , \8540 );
and \U$15968 ( \16165 , \2090 , \8292 );
nor \U$15969 ( \16166 , \16164 , \16165 );
xnor \U$15970 ( \16167 , \16166 , \8297 );
xor \U$15971 ( \16168 , \16163 , \16167 );
and \U$15972 ( \16169 , \1684 , \9333 );
and \U$15973 ( \16170 , \1802 , \9006 );
nor \U$15974 ( \16171 , \16169 , \16170 );
xnor \U$15975 ( \16172 , \16171 , \8848 );
xor \U$15976 ( \16173 , \16168 , \16172 );
xor \U$15977 ( \16174 , \16159 , \16173 );
xor \U$15978 ( \16175 , \16130 , \16174 );
xor \U$15979 ( \16176 , \16074 , \16175 );
and \U$15980 ( \16177 , \15958 , \15962 );
and \U$15981 ( \16178 , \15962 , \15967 );
and \U$15982 ( \16179 , \15958 , \15967 );
or \U$15983 ( \16180 , \16177 , \16178 , \16179 );
and \U$15984 ( \16181 , \15972 , \15976 );
and \U$15985 ( \16182 , \15976 , \15981 );
and \U$15986 ( \16183 , \15972 , \15981 );
or \U$15987 ( \16184 , \16181 , \16182 , \16183 );
xor \U$15988 ( \16185 , \16180 , \16184 );
and \U$15989 ( \16186 , \15902 , \15906 );
and \U$15990 ( \16187 , \15906 , \15911 );
and \U$15991 ( \16188 , \15902 , \15911 );
or \U$15992 ( \16189 , \16186 , \16187 , \16188 );
xor \U$15993 ( \16190 , \16185 , \16189 );
and \U$15994 ( \16191 , \15873 , \15877 );
and \U$15995 ( \16192 , \15877 , \15882 );
and \U$15996 ( \16193 , \15873 , \15882 );
or \U$15997 ( \16194 , \16191 , \16192 , \16193 );
and \U$15998 ( \16195 , \15887 , \15891 );
and \U$15999 ( \16196 , \15891 , \15896 );
and \U$16000 ( \16197 , \15887 , \15896 );
or \U$16001 ( \16198 , \16195 , \16196 , \16197 );
xor \U$16002 ( \16199 , \16194 , \16198 );
and \U$16003 ( \16200 , \15917 , \15921 );
and \U$16004 ( \16201 , \15921 , \15926 );
and \U$16005 ( \16202 , \15917 , \15926 );
or \U$16006 ( \16203 , \16200 , \16201 , \16202 );
xor \U$16007 ( \16204 , \16199 , \16203 );
xor \U$16008 ( \16205 , \16190 , \16204 );
and \U$16009 ( \16206 , \15931 , \15935 );
and \U$16010 ( \16207 , \15935 , \15940 );
and \U$16011 ( \16208 , \15931 , \15940 );
or \U$16012 ( \16209 , \16206 , \16207 , \16208 );
and \U$16013 ( \16210 , \15946 , \15950 );
and \U$16014 ( \16211 , \15950 , \15952 );
and \U$16015 ( \16212 , \15946 , \15952 );
or \U$16016 ( \16213 , \16210 , \16211 , \16212 );
xor \U$16017 ( \16214 , \16209 , \16213 );
and \U$16018 ( \16215 , \1484 , \9765 );
and \U$16019 ( \16216 , \1601 , \9644 );
nor \U$16020 ( \16217 , \16215 , \16216 );
xnor \U$16021 ( \16218 , \16217 , \9478 );
and \U$16022 ( \16219 , \1192 , \10408 );
and \U$16023 ( \16220 , \1333 , \10116 );
nor \U$16024 ( \16221 , \16219 , \16220 );
xnor \U$16025 ( \16222 , \16221 , \10121 );
xor \U$16026 ( \16223 , \16218 , \16222 );
and \U$16027 ( \16224 , \1147 , \10118 );
xor \U$16028 ( \16225 , \16223 , \16224 );
xor \U$16029 ( \16226 , \16214 , \16225 );
xor \U$16030 ( \16227 , \16205 , \16226 );
xor \U$16031 ( \16228 , \16176 , \16227 );
xor \U$16032 ( \16229 , \16070 , \16228 );
and \U$16033 ( \16230 , \15833 , \15837 );
and \U$16034 ( \16231 , \15837 , \15842 );
and \U$16035 ( \16232 , \15833 , \15842 );
or \U$16036 ( \16233 , \16230 , \16231 , \16232 );
and \U$16037 ( \16234 , \15847 , \15851 );
and \U$16038 ( \16235 , \15851 , \15856 );
and \U$16039 ( \16236 , \15847 , \15856 );
or \U$16040 ( \16237 , \16234 , \16235 , \16236 );
xor \U$16041 ( \16238 , \16233 , \16237 );
or \U$16042 ( \16239 , \15862 , \15866 );
xor \U$16043 ( \16240 , \16238 , \16239 );
and \U$16044 ( \16241 , \15883 , \15897 );
and \U$16045 ( \16242 , \15897 , \15912 );
and \U$16046 ( \16243 , \15883 , \15912 );
or \U$16047 ( \16244 , \16241 , \16242 , \16243 );
and \U$16048 ( \16245 , \15927 , \15941 );
and \U$16049 ( \16246 , \15941 , \15953 );
and \U$16050 ( \16247 , \15927 , \15953 );
or \U$16051 ( \16248 , \16245 , \16246 , \16247 );
xor \U$16052 ( \16249 , \16244 , \16248 );
and \U$16053 ( \16250 , \15968 , \15982 );
xor \U$16054 ( \16251 , \16249 , \16250 );
xor \U$16055 ( \16252 , \16240 , \16251 );
xor \U$16056 ( \16253 , \16229 , \16252 );
xor \U$16057 ( \16254 , \16056 , \16253 );
xor \U$16058 ( \16255 , \16047 , \16254 );
xor \U$16059 ( \16256 , \16031 , \16255 );
and \U$16060 ( \16257 , \15786 , \16018 );
xor \U$16061 ( \16258 , \16256 , \16257 );
and \U$16062 ( \16259 , \16019 , \16020 );
and \U$16063 ( \16260 , \16021 , \16024 );
or \U$16064 ( \16261 , \16259 , \16260 );
xor \U$16065 ( \16262 , \16258 , \16261 );
buf g54f5_GF_PartitionCandidate( \16263_nG54f5 , \16262 );
buf \U$16066 ( \16264 , \16263_nG54f5 );
and \U$16067 ( \16265 , \16035 , \16046 );
and \U$16068 ( \16266 , \16046 , \16254 );
and \U$16069 ( \16267 , \16035 , \16254 );
or \U$16070 ( \16268 , \16265 , \16266 , \16267 );
and \U$16071 ( \16269 , \16051 , \16055 );
and \U$16072 ( \16270 , \16055 , \16253 );
and \U$16073 ( \16271 , \16051 , \16253 );
or \U$16074 ( \16272 , \16269 , \16270 , \16271 );
and \U$16075 ( \16273 , \16060 , \16064 );
and \U$16076 ( \16274 , \16064 , \16069 );
and \U$16077 ( \16275 , \16060 , \16069 );
or \U$16078 ( \16276 , \16273 , \16274 , \16275 );
and \U$16079 ( \16277 , \16074 , \16175 );
and \U$16080 ( \16278 , \16175 , \16227 );
and \U$16081 ( \16279 , \16074 , \16227 );
or \U$16082 ( \16280 , \16277 , \16278 , \16279 );
xor \U$16083 ( \16281 , \16276 , \16280 );
and \U$16084 ( \16282 , \16240 , \16251 );
xor \U$16085 ( \16283 , \16281 , \16282 );
xor \U$16086 ( \16284 , \16272 , \16283 );
and \U$16087 ( \16285 , \16039 , \16043 );
and \U$16088 ( \16286 , \16043 , \16045 );
and \U$16089 ( \16287 , \16039 , \16045 );
or \U$16090 ( \16288 , \16285 , \16286 , \16287 );
and \U$16091 ( \16289 , \16070 , \16228 );
and \U$16092 ( \16290 , \16228 , \16252 );
and \U$16093 ( \16291 , \16070 , \16252 );
or \U$16094 ( \16292 , \16289 , \16290 , \16291 );
xor \U$16095 ( \16293 , \16288 , \16292 );
and \U$16096 ( \16294 , \16233 , \16237 );
and \U$16097 ( \16295 , \16237 , \16239 );
and \U$16098 ( \16296 , \16233 , \16239 );
or \U$16099 ( \16297 , \16294 , \16295 , \16296 );
and \U$16100 ( \16298 , \16244 , \16248 );
and \U$16101 ( \16299 , \16248 , \16250 );
and \U$16102 ( \16300 , \16244 , \16250 );
or \U$16103 ( \16301 , \16298 , \16299 , \16300 );
xor \U$16104 ( \16302 , \16297 , \16301 );
and \U$16105 ( \16303 , \16085 , \16129 );
and \U$16106 ( \16304 , \16129 , \16174 );
and \U$16107 ( \16305 , \16085 , \16174 );
or \U$16108 ( \16306 , \16303 , \16304 , \16305 );
xor \U$16109 ( \16307 , \16302 , \16306 );
and \U$16110 ( \16308 , \16190 , \16204 );
and \U$16111 ( \16309 , \16204 , \16226 );
and \U$16112 ( \16310 , \16190 , \16226 );
or \U$16113 ( \16311 , \16308 , \16309 , \16310 );
and \U$16114 ( \16312 , \16075 , \16079 );
and \U$16115 ( \16313 , \16079 , \16084 );
and \U$16116 ( \16314 , \16075 , \16084 );
or \U$16117 ( \16315 , \16312 , \16313 , \16314 );
and \U$16118 ( \16316 , \16103 , \16107 );
and \U$16119 ( \16317 , \16107 , \16112 );
and \U$16120 ( \16318 , \16103 , \16112 );
or \U$16121 ( \16319 , \16316 , \16317 , \16318 );
xor \U$16122 ( \16320 , \16315 , \16319 );
and \U$16123 ( \16321 , \16118 , \16122 );
and \U$16124 ( \16322 , \16122 , \16127 );
and \U$16125 ( \16323 , \16118 , \16127 );
or \U$16126 ( \16324 , \16321 , \16322 , \16323 );
xor \U$16127 ( \16325 , \16320 , \16324 );
xor \U$16128 ( \16326 , \16311 , \16325 );
and \U$16129 ( \16327 , \16089 , \16093 );
and \U$16130 ( \16328 , \16093 , \16098 );
and \U$16131 ( \16329 , \16089 , \16098 );
or \U$16132 ( \16330 , \16327 , \16328 , \16329 );
and \U$16133 ( \16331 , \16134 , \16138 );
and \U$16134 ( \16332 , \16138 , \16143 );
and \U$16135 ( \16333 , \16134 , \16143 );
or \U$16136 ( \16334 , \16331 , \16332 , \16333 );
xor \U$16137 ( \16335 , \16330 , \16334 );
and \U$16138 ( \16336 , \16148 , \16152 );
and \U$16139 ( \16337 , \16152 , \16157 );
and \U$16140 ( \16338 , \16148 , \16157 );
or \U$16141 ( \16339 , \16336 , \16337 , \16338 );
xor \U$16142 ( \16340 , \16335 , \16339 );
xor \U$16143 ( \16341 , \16326 , \16340 );
xor \U$16144 ( \16342 , \16307 , \16341 );
and \U$16145 ( \16343 , \16180 , \16184 );
and \U$16146 ( \16344 , \16184 , \16189 );
and \U$16147 ( \16345 , \16180 , \16189 );
or \U$16148 ( \16346 , \16343 , \16344 , \16345 );
and \U$16149 ( \16347 , \16194 , \16198 );
and \U$16150 ( \16348 , \16198 , \16203 );
and \U$16151 ( \16349 , \16194 , \16203 );
or \U$16152 ( \16350 , \16347 , \16348 , \16349 );
xor \U$16153 ( \16351 , \16346 , \16350 );
and \U$16154 ( \16352 , \16209 , \16213 );
and \U$16155 ( \16353 , \16213 , \16225 );
and \U$16156 ( \16354 , \16209 , \16225 );
or \U$16157 ( \16355 , \16352 , \16353 , \16354 );
xor \U$16158 ( \16356 , \16351 , \16355 );
and \U$16159 ( \16357 , \16099 , \16113 );
and \U$16160 ( \16358 , \16113 , \16128 );
and \U$16161 ( \16359 , \16099 , \16128 );
or \U$16162 ( \16360 , \16357 , \16358 , \16359 );
and \U$16163 ( \16361 , \16144 , \16158 );
and \U$16164 ( \16362 , \16158 , \16173 );
and \U$16165 ( \16363 , \16144 , \16173 );
or \U$16166 ( \16364 , \16361 , \16362 , \16363 );
xor \U$16167 ( \16365 , \16360 , \16364 );
and \U$16168 ( \16366 , \10584 , \1301 );
not \U$16169 ( \16367 , \16366 );
xnor \U$16170 ( \16368 , \16367 , \1205 );
and \U$16171 ( \16369 , \9897 , \1578 );
and \U$16172 ( \16370 , \10206 , \1431 );
nor \U$16173 ( \16371 , \16369 , \16370 );
xnor \U$16174 ( \16372 , \16371 , \1436 );
xor \U$16175 ( \16373 , \16368 , \16372 );
and \U$16176 ( \16374 , \9169 , \1824 );
and \U$16177 ( \16375 , \9465 , \1739 );
nor \U$16178 ( \16376 , \16374 , \16375 );
xnor \U$16179 ( \16377 , \16376 , \1697 );
xor \U$16180 ( \16378 , \16373 , \16377 );
xor \U$16181 ( \16379 , \16365 , \16378 );
xor \U$16182 ( \16380 , \16356 , \16379 );
and \U$16183 ( \16381 , \2090 , \8540 );
and \U$16184 ( \16382 , \2182 , \8292 );
nor \U$16185 ( \16383 , \16381 , \16382 );
xnor \U$16186 ( \16384 , \16383 , \8297 );
and \U$16187 ( \16385 , \1802 , \9333 );
and \U$16188 ( \16386 , \1948 , \9006 );
nor \U$16189 ( \16387 , \16385 , \16386 );
xnor \U$16190 ( \16388 , \16387 , \8848 );
xor \U$16191 ( \16389 , \16384 , \16388 );
and \U$16192 ( \16390 , \1601 , \9765 );
and \U$16193 ( \16391 , \1684 , \9644 );
nor \U$16194 ( \16392 , \16390 , \16391 );
xnor \U$16195 ( \16393 , \16392 , \9478 );
xor \U$16196 ( \16394 , \16389 , \16393 );
and \U$16197 ( \16395 , \4160 , \5485 );
and \U$16198 ( \16396 , \4364 , \5275 );
nor \U$16199 ( \16397 , \16395 , \16396 );
xnor \U$16200 ( \16398 , \16397 , \5169 );
and \U$16201 ( \16399 , \3736 , \5996 );
and \U$16202 ( \16400 , \3912 , \5695 );
nor \U$16203 ( \16401 , \16399 , \16400 );
xnor \U$16204 ( \16402 , \16401 , \5687 );
xor \U$16205 ( \16403 , \16398 , \16402 );
and \U$16206 ( \16404 , \3395 , \6401 );
and \U$16207 ( \16405 , \3646 , \6143 );
nor \U$16208 ( \16406 , \16404 , \16405 );
xnor \U$16209 ( \16407 , \16406 , \6148 );
xor \U$16210 ( \16408 , \16403 , \16407 );
xor \U$16211 ( \16409 , \16394 , \16408 );
and \U$16212 ( \16410 , \3037 , \7055 );
and \U$16213 ( \16411 , \3143 , \6675 );
nor \U$16214 ( \16412 , \16410 , \16411 );
xnor \U$16215 ( \16413 , \16412 , \6680 );
and \U$16216 ( \16414 , \2757 , \7489 );
and \U$16217 ( \16415 , \2826 , \7137 );
nor \U$16218 ( \16416 , \16414 , \16415 );
xnor \U$16219 ( \16417 , \16416 , \7142 );
xor \U$16220 ( \16418 , \16413 , \16417 );
and \U$16221 ( \16419 , \2366 , \8019 );
and \U$16222 ( \16420 , \2521 , \7830 );
nor \U$16223 ( \16421 , \16419 , \16420 );
xnor \U$16224 ( \16422 , \16421 , \7713 );
xor \U$16225 ( \16423 , \16418 , \16422 );
xor \U$16226 ( \16424 , \16409 , \16423 );
and \U$16227 ( \16425 , \5469 , \4132 );
and \U$16228 ( \16426 , \5674 , \4012 );
nor \U$16229 ( \16427 , \16425 , \16426 );
xnor \U$16230 ( \16428 , \16427 , \3925 );
and \U$16231 ( \16429 , \4922 , \4581 );
and \U$16232 ( \16430 , \5156 , \4424 );
nor \U$16233 ( \16431 , \16429 , \16430 );
xnor \U$16234 ( \16432 , \16431 , \4377 );
xor \U$16235 ( \16433 , \16428 , \16432 );
and \U$16236 ( \16434 , \4654 , \5011 );
and \U$16237 ( \16435 , \4749 , \4878 );
nor \U$16238 ( \16436 , \16434 , \16435 );
xnor \U$16239 ( \16437 , \16436 , \4762 );
xor \U$16240 ( \16438 , \16433 , \16437 );
and \U$16241 ( \16439 , \6945 , \3103 );
and \U$16242 ( \16440 , \7231 , \2934 );
nor \U$16243 ( \16441 , \16439 , \16440 );
xnor \U$16244 ( \16442 , \16441 , \2839 );
and \U$16245 ( \16443 , \6514 , \3357 );
and \U$16246 ( \16444 , \6790 , \3255 );
nor \U$16247 ( \16445 , \16443 , \16444 );
xnor \U$16248 ( \16446 , \16445 , \3156 );
xor \U$16249 ( \16447 , \16442 , \16446 );
and \U$16250 ( \16448 , \6030 , \3813 );
and \U$16251 ( \16449 , \6281 , \3557 );
nor \U$16252 ( \16450 , \16448 , \16449 );
xnor \U$16253 ( \16451 , \16450 , \3562 );
xor \U$16254 ( \16452 , \16447 , \16451 );
xor \U$16255 ( \16453 , \16438 , \16452 );
and \U$16256 ( \16454 , \8652 , \2121 );
and \U$16257 ( \16455 , \8835 , \2008 );
nor \U$16258 ( \16456 , \16454 , \16455 );
xnor \U$16259 ( \16457 , \16456 , \1961 );
and \U$16260 ( \16458 , \8057 , \2400 );
and \U$16261 ( \16459 , \8349 , \2246 );
nor \U$16262 ( \16460 , \16458 , \16459 );
xnor \U$16263 ( \16461 , \16460 , \2195 );
xor \U$16264 ( \16462 , \16457 , \16461 );
and \U$16265 ( \16463 , \7556 , \2669 );
and \U$16266 ( \16464 , \7700 , \2538 );
nor \U$16267 ( \16465 , \16463 , \16464 );
xnor \U$16268 ( \16466 , \16465 , \2534 );
xor \U$16269 ( \16467 , \16462 , \16466 );
xor \U$16270 ( \16468 , \16453 , \16467 );
xor \U$16271 ( \16469 , \16424 , \16468 );
and \U$16272 ( \16470 , \16218 , \16222 );
and \U$16273 ( \16471 , \16222 , \16224 );
and \U$16274 ( \16472 , \16218 , \16224 );
or \U$16275 ( \16473 , \16470 , \16471 , \16472 );
and \U$16276 ( \16474 , \16163 , \16167 );
and \U$16277 ( \16475 , \16167 , \16172 );
and \U$16278 ( \16476 , \16163 , \16172 );
or \U$16279 ( \16477 , \16474 , \16475 , \16476 );
xor \U$16280 ( \16478 , \16473 , \16477 );
and \U$16281 ( \16479 , \1333 , \10408 );
and \U$16282 ( \16480 , \1484 , \10116 );
nor \U$16283 ( \16481 , \16479 , \16480 );
xnor \U$16284 ( \16482 , \16481 , \10121 );
and \U$16285 ( \16483 , \1192 , \10118 );
xnor \U$16286 ( \16484 , \16482 , \16483 );
xor \U$16287 ( \16485 , \16478 , \16484 );
xor \U$16288 ( \16486 , \16469 , \16485 );
xor \U$16289 ( \16487 , \16380 , \16486 );
xor \U$16290 ( \16488 , \16342 , \16487 );
xor \U$16291 ( \16489 , \16293 , \16488 );
xor \U$16292 ( \16490 , \16284 , \16489 );
xor \U$16293 ( \16491 , \16268 , \16490 );
and \U$16294 ( \16492 , \16031 , \16255 );
xor \U$16295 ( \16493 , \16491 , \16492 );
and \U$16296 ( \16494 , \16256 , \16257 );
and \U$16297 ( \16495 , \16258 , \16261 );
or \U$16298 ( \16496 , \16494 , \16495 );
xor \U$16299 ( \16497 , \16493 , \16496 );
buf g54f3_GF_PartitionCandidate( \16498_nG54f3 , \16497 );
buf \U$16300 ( \16499 , \16498_nG54f3 );
and \U$16301 ( \16500 , \16272 , \16283 );
and \U$16302 ( \16501 , \16283 , \16489 );
and \U$16303 ( \16502 , \16272 , \16489 );
or \U$16304 ( \16503 , \16500 , \16501 , \16502 );
and \U$16305 ( \16504 , \16288 , \16292 );
and \U$16306 ( \16505 , \16292 , \16488 );
and \U$16307 ( \16506 , \16288 , \16488 );
or \U$16308 ( \16507 , \16504 , \16505 , \16506 );
and \U$16309 ( \16508 , \16297 , \16301 );
and \U$16310 ( \16509 , \16301 , \16306 );
and \U$16311 ( \16510 , \16297 , \16306 );
or \U$16312 ( \16511 , \16508 , \16509 , \16510 );
and \U$16313 ( \16512 , \16311 , \16325 );
and \U$16314 ( \16513 , \16325 , \16340 );
and \U$16315 ( \16514 , \16311 , \16340 );
or \U$16316 ( \16515 , \16512 , \16513 , \16514 );
xor \U$16317 ( \16516 , \16511 , \16515 );
and \U$16318 ( \16517 , \16356 , \16379 );
and \U$16319 ( \16518 , \16379 , \16486 );
and \U$16320 ( \16519 , \16356 , \16486 );
or \U$16321 ( \16520 , \16517 , \16518 , \16519 );
xor \U$16322 ( \16521 , \16516 , \16520 );
xor \U$16323 ( \16522 , \16507 , \16521 );
and \U$16324 ( \16523 , \16276 , \16280 );
and \U$16325 ( \16524 , \16280 , \16282 );
and \U$16326 ( \16525 , \16276 , \16282 );
or \U$16327 ( \16526 , \16523 , \16524 , \16525 );
and \U$16328 ( \16527 , \16307 , \16341 );
and \U$16329 ( \16528 , \16341 , \16487 );
and \U$16330 ( \16529 , \16307 , \16487 );
or \U$16331 ( \16530 , \16527 , \16528 , \16529 );
xor \U$16332 ( \16531 , \16526 , \16530 );
and \U$16333 ( \16532 , \16315 , \16319 );
and \U$16334 ( \16533 , \16319 , \16324 );
and \U$16335 ( \16534 , \16315 , \16324 );
or \U$16336 ( \16535 , \16532 , \16533 , \16534 );
and \U$16337 ( \16536 , \16330 , \16334 );
and \U$16338 ( \16537 , \16334 , \16339 );
and \U$16339 ( \16538 , \16330 , \16339 );
or \U$16340 ( \16539 , \16536 , \16537 , \16538 );
xor \U$16341 ( \16540 , \16535 , \16539 );
and \U$16342 ( \16541 , \16473 , \16477 );
and \U$16343 ( \16542 , \16477 , \16484 );
and \U$16344 ( \16543 , \16473 , \16484 );
or \U$16345 ( \16544 , \16541 , \16542 , \16543 );
xor \U$16346 ( \16545 , \16540 , \16544 );
and \U$16347 ( \16546 , \16346 , \16350 );
and \U$16348 ( \16547 , \16350 , \16355 );
and \U$16349 ( \16548 , \16346 , \16355 );
or \U$16350 ( \16549 , \16546 , \16547 , \16548 );
and \U$16351 ( \16550 , \16360 , \16364 );
and \U$16352 ( \16551 , \16364 , \16378 );
and \U$16353 ( \16552 , \16360 , \16378 );
or \U$16354 ( \16553 , \16550 , \16551 , \16552 );
xor \U$16355 ( \16554 , \16549 , \16553 );
and \U$16356 ( \16555 , \16424 , \16468 );
and \U$16357 ( \16556 , \16468 , \16485 );
and \U$16358 ( \16557 , \16424 , \16485 );
or \U$16359 ( \16558 , \16555 , \16556 , \16557 );
xor \U$16360 ( \16559 , \16554 , \16558 );
xor \U$16361 ( \16560 , \16545 , \16559 );
and \U$16362 ( \16561 , \16394 , \16408 );
and \U$16363 ( \16562 , \16408 , \16423 );
and \U$16364 ( \16563 , \16394 , \16423 );
or \U$16365 ( \16564 , \16561 , \16562 , \16563 );
and \U$16366 ( \16565 , \16438 , \16452 );
and \U$16367 ( \16566 , \16452 , \16467 );
and \U$16368 ( \16567 , \16438 , \16467 );
or \U$16369 ( \16568 , \16565 , \16566 , \16567 );
xor \U$16370 ( \16569 , \16564 , \16568 );
and \U$16371 ( \16570 , \8835 , \2121 );
and \U$16372 ( \16571 , \9169 , \2008 );
nor \U$16373 ( \16572 , \16570 , \16571 );
xnor \U$16374 ( \16573 , \16572 , \1961 );
and \U$16375 ( \16574 , \8349 , \2400 );
and \U$16376 ( \16575 , \8652 , \2246 );
nor \U$16377 ( \16576 , \16574 , \16575 );
xnor \U$16378 ( \16577 , \16576 , \2195 );
xor \U$16379 ( \16578 , \16573 , \16577 );
and \U$16380 ( \16579 , \7700 , \2669 );
and \U$16381 ( \16580 , \8057 , \2538 );
nor \U$16382 ( \16581 , \16579 , \16580 );
xnor \U$16383 ( \16582 , \16581 , \2534 );
xor \U$16384 ( \16583 , \16578 , \16582 );
xor \U$16385 ( \16584 , \16569 , \16583 );
and \U$16386 ( \16585 , \16368 , \16372 );
and \U$16387 ( \16586 , \16372 , \16377 );
and \U$16388 ( \16587 , \16368 , \16377 );
or \U$16389 ( \16588 , \16585 , \16586 , \16587 );
and \U$16390 ( \16589 , \16442 , \16446 );
and \U$16391 ( \16590 , \16446 , \16451 );
and \U$16392 ( \16591 , \16442 , \16451 );
or \U$16393 ( \16592 , \16589 , \16590 , \16591 );
xor \U$16394 ( \16593 , \16588 , \16592 );
and \U$16395 ( \16594 , \16457 , \16461 );
and \U$16396 ( \16595 , \16461 , \16466 );
and \U$16397 ( \16596 , \16457 , \16466 );
or \U$16398 ( \16597 , \16594 , \16595 , \16596 );
xor \U$16399 ( \16598 , \16593 , \16597 );
and \U$16400 ( \16599 , \16384 , \16388 );
and \U$16401 ( \16600 , \16388 , \16393 );
and \U$16402 ( \16601 , \16384 , \16393 );
or \U$16403 ( \16602 , \16599 , \16600 , \16601 );
or \U$16404 ( \16603 , \16482 , \16483 );
xor \U$16405 ( \16604 , \16602 , \16603 );
and \U$16406 ( \16605 , \1484 , \10408 );
and \U$16407 ( \16606 , \1601 , \10116 );
nor \U$16408 ( \16607 , \16605 , \16606 );
xnor \U$16409 ( \16608 , \16607 , \10121 );
xor \U$16410 ( \16609 , \16604 , \16608 );
xor \U$16411 ( \16610 , \16598 , \16609 );
and \U$16412 ( \16611 , \16428 , \16432 );
and \U$16413 ( \16612 , \16432 , \16437 );
and \U$16414 ( \16613 , \16428 , \16437 );
or \U$16415 ( \16614 , \16611 , \16612 , \16613 );
and \U$16416 ( \16615 , \16398 , \16402 );
and \U$16417 ( \16616 , \16402 , \16407 );
and \U$16418 ( \16617 , \16398 , \16407 );
or \U$16419 ( \16618 , \16615 , \16616 , \16617 );
xor \U$16420 ( \16619 , \16614 , \16618 );
and \U$16421 ( \16620 , \16413 , \16417 );
and \U$16422 ( \16621 , \16417 , \16422 );
and \U$16423 ( \16622 , \16413 , \16422 );
or \U$16424 ( \16623 , \16620 , \16621 , \16622 );
xor \U$16425 ( \16624 , \16619 , \16623 );
xor \U$16426 ( \16625 , \16610 , \16624 );
xor \U$16427 ( \16626 , \16584 , \16625 );
not \U$16428 ( \16627 , \1205 );
and \U$16429 ( \16628 , \10206 , \1578 );
and \U$16430 ( \16629 , \10584 , \1431 );
nor \U$16431 ( \16630 , \16628 , \16629 );
xnor \U$16432 ( \16631 , \16630 , \1436 );
xor \U$16433 ( \16632 , \16627 , \16631 );
and \U$16434 ( \16633 , \9465 , \1824 );
and \U$16435 ( \16634 , \9897 , \1739 );
nor \U$16436 ( \16635 , \16633 , \16634 );
xnor \U$16437 ( \16636 , \16635 , \1697 );
xor \U$16438 ( \16637 , \16632 , \16636 );
and \U$16439 ( \16638 , \1333 , \10118 );
and \U$16440 ( \16639 , \2182 , \8540 );
and \U$16441 ( \16640 , \2366 , \8292 );
nor \U$16442 ( \16641 , \16639 , \16640 );
xnor \U$16443 ( \16642 , \16641 , \8297 );
and \U$16444 ( \16643 , \1948 , \9333 );
and \U$16445 ( \16644 , \2090 , \9006 );
nor \U$16446 ( \16645 , \16643 , \16644 );
xnor \U$16447 ( \16646 , \16645 , \8848 );
xor \U$16448 ( \16647 , \16642 , \16646 );
and \U$16449 ( \16648 , \1684 , \9765 );
and \U$16450 ( \16649 , \1802 , \9644 );
nor \U$16451 ( \16650 , \16648 , \16649 );
xnor \U$16452 ( \16651 , \16650 , \9478 );
xor \U$16453 ( \16652 , \16647 , \16651 );
xor \U$16454 ( \16653 , \16638 , \16652 );
and \U$16455 ( \16654 , \3143 , \7055 );
and \U$16456 ( \16655 , \3395 , \6675 );
nor \U$16457 ( \16656 , \16654 , \16655 );
xnor \U$16458 ( \16657 , \16656 , \6680 );
and \U$16459 ( \16658 , \2826 , \7489 );
and \U$16460 ( \16659 , \3037 , \7137 );
nor \U$16461 ( \16660 , \16658 , \16659 );
xnor \U$16462 ( \16661 , \16660 , \7142 );
xor \U$16463 ( \16662 , \16657 , \16661 );
and \U$16464 ( \16663 , \2521 , \8019 );
and \U$16465 ( \16664 , \2757 , \7830 );
nor \U$16466 ( \16665 , \16663 , \16664 );
xnor \U$16467 ( \16666 , \16665 , \7713 );
xor \U$16468 ( \16667 , \16662 , \16666 );
xor \U$16469 ( \16668 , \16653 , \16667 );
xor \U$16470 ( \16669 , \16637 , \16668 );
and \U$16471 ( \16670 , \5674 , \4132 );
and \U$16472 ( \16671 , \6030 , \4012 );
nor \U$16473 ( \16672 , \16670 , \16671 );
xnor \U$16474 ( \16673 , \16672 , \3925 );
and \U$16475 ( \16674 , \5156 , \4581 );
and \U$16476 ( \16675 , \5469 , \4424 );
nor \U$16477 ( \16676 , \16674 , \16675 );
xnor \U$16478 ( \16677 , \16676 , \4377 );
xor \U$16479 ( \16678 , \16673 , \16677 );
and \U$16480 ( \16679 , \4749 , \5011 );
and \U$16481 ( \16680 , \4922 , \4878 );
nor \U$16482 ( \16681 , \16679 , \16680 );
xnor \U$16483 ( \16682 , \16681 , \4762 );
xor \U$16484 ( \16683 , \16678 , \16682 );
and \U$16485 ( \16684 , \7231 , \3103 );
and \U$16486 ( \16685 , \7556 , \2934 );
nor \U$16487 ( \16686 , \16684 , \16685 );
xnor \U$16488 ( \16687 , \16686 , \2839 );
and \U$16489 ( \16688 , \6790 , \3357 );
and \U$16490 ( \16689 , \6945 , \3255 );
nor \U$16491 ( \16690 , \16688 , \16689 );
xnor \U$16492 ( \16691 , \16690 , \3156 );
xor \U$16493 ( \16692 , \16687 , \16691 );
and \U$16494 ( \16693 , \6281 , \3813 );
and \U$16495 ( \16694 , \6514 , \3557 );
nor \U$16496 ( \16695 , \16693 , \16694 );
xnor \U$16497 ( \16696 , \16695 , \3562 );
xor \U$16498 ( \16697 , \16692 , \16696 );
xor \U$16499 ( \16698 , \16683 , \16697 );
and \U$16500 ( \16699 , \4364 , \5485 );
and \U$16501 ( \16700 , \4654 , \5275 );
nor \U$16502 ( \16701 , \16699 , \16700 );
xnor \U$16503 ( \16702 , \16701 , \5169 );
and \U$16504 ( \16703 , \3912 , \5996 );
and \U$16505 ( \16704 , \4160 , \5695 );
nor \U$16506 ( \16705 , \16703 , \16704 );
xnor \U$16507 ( \16706 , \16705 , \5687 );
xor \U$16508 ( \16707 , \16702 , \16706 );
and \U$16509 ( \16708 , \3646 , \6401 );
and \U$16510 ( \16709 , \3736 , \6143 );
nor \U$16511 ( \16710 , \16708 , \16709 );
xnor \U$16512 ( \16711 , \16710 , \6148 );
xor \U$16513 ( \16712 , \16707 , \16711 );
xor \U$16514 ( \16713 , \16698 , \16712 );
xor \U$16515 ( \16714 , \16669 , \16713 );
xor \U$16516 ( \16715 , \16626 , \16714 );
xor \U$16517 ( \16716 , \16560 , \16715 );
xor \U$16518 ( \16717 , \16531 , \16716 );
xor \U$16519 ( \16718 , \16522 , \16717 );
xor \U$16520 ( \16719 , \16503 , \16718 );
and \U$16521 ( \16720 , \16268 , \16490 );
xor \U$16522 ( \16721 , \16719 , \16720 );
and \U$16523 ( \16722 , \16491 , \16492 );
and \U$16524 ( \16723 , \16493 , \16496 );
or \U$16525 ( \16724 , \16722 , \16723 );
xor \U$16526 ( \16725 , \16721 , \16724 );
buf g54f1_GF_PartitionCandidate( \16726_nG54f1 , \16725 );
buf \U$16527 ( \16727 , \16726_nG54f1 );
and \U$16528 ( \16728 , \16507 , \16521 );
and \U$16529 ( \16729 , \16521 , \16717 );
and \U$16530 ( \16730 , \16507 , \16717 );
or \U$16531 ( \16731 , \16728 , \16729 , \16730 );
and \U$16532 ( \16732 , \16526 , \16530 );
and \U$16533 ( \16733 , \16530 , \16716 );
and \U$16534 ( \16734 , \16526 , \16716 );
or \U$16535 ( \16735 , \16732 , \16733 , \16734 );
and \U$16536 ( \16736 , \16549 , \16553 );
and \U$16537 ( \16737 , \16553 , \16558 );
and \U$16538 ( \16738 , \16549 , \16558 );
or \U$16539 ( \16739 , \16736 , \16737 , \16738 );
and \U$16540 ( \16740 , \16584 , \16625 );
and \U$16541 ( \16741 , \16625 , \16714 );
and \U$16542 ( \16742 , \16584 , \16714 );
or \U$16543 ( \16743 , \16740 , \16741 , \16742 );
xor \U$16544 ( \16744 , \16739 , \16743 );
and \U$16545 ( \16745 , \16638 , \16652 );
and \U$16546 ( \16746 , \16652 , \16667 );
and \U$16547 ( \16747 , \16638 , \16667 );
or \U$16548 ( \16748 , \16745 , \16746 , \16747 );
and \U$16549 ( \16749 , \16683 , \16697 );
and \U$16550 ( \16750 , \16697 , \16712 );
and \U$16551 ( \16751 , \16683 , \16712 );
or \U$16552 ( \16752 , \16749 , \16750 , \16751 );
xor \U$16553 ( \16753 , \16748 , \16752 );
and \U$16554 ( \16754 , \6945 , \3357 );
and \U$16555 ( \16755 , \7231 , \3255 );
nor \U$16556 ( \16756 , \16754 , \16755 );
xnor \U$16557 ( \16757 , \16756 , \3156 );
and \U$16558 ( \16758 , \6514 , \3813 );
and \U$16559 ( \16759 , \6790 , \3557 );
nor \U$16560 ( \16760 , \16758 , \16759 );
xnor \U$16561 ( \16761 , \16760 , \3562 );
xor \U$16562 ( \16762 , \16757 , \16761 );
and \U$16563 ( \16763 , \6030 , \4132 );
and \U$16564 ( \16764 , \6281 , \4012 );
nor \U$16565 ( \16765 , \16763 , \16764 );
xnor \U$16566 ( \16766 , \16765 , \3925 );
xor \U$16567 ( \16767 , \16762 , \16766 );
and \U$16568 ( \16768 , \10584 , \1578 );
not \U$16569 ( \16769 , \16768 );
xnor \U$16570 ( \16770 , \16769 , \1436 );
and \U$16571 ( \16771 , \9897 , \1824 );
and \U$16572 ( \16772 , \10206 , \1739 );
nor \U$16573 ( \16773 , \16771 , \16772 );
xnor \U$16574 ( \16774 , \16773 , \1697 );
xor \U$16575 ( \16775 , \16770 , \16774 );
and \U$16576 ( \16776 , \9169 , \2121 );
and \U$16577 ( \16777 , \9465 , \2008 );
nor \U$16578 ( \16778 , \16776 , \16777 );
xnor \U$16579 ( \16779 , \16778 , \1961 );
xor \U$16580 ( \16780 , \16775 , \16779 );
xor \U$16581 ( \16781 , \16767 , \16780 );
and \U$16582 ( \16782 , \8652 , \2400 );
and \U$16583 ( \16783 , \8835 , \2246 );
nor \U$16584 ( \16784 , \16782 , \16783 );
xnor \U$16585 ( \16785 , \16784 , \2195 );
and \U$16586 ( \16786 , \8057 , \2669 );
and \U$16587 ( \16787 , \8349 , \2538 );
nor \U$16588 ( \16788 , \16786 , \16787 );
xnor \U$16589 ( \16789 , \16788 , \2534 );
xor \U$16590 ( \16790 , \16785 , \16789 );
and \U$16591 ( \16791 , \7556 , \3103 );
and \U$16592 ( \16792 , \7700 , \2934 );
nor \U$16593 ( \16793 , \16791 , \16792 );
xnor \U$16594 ( \16794 , \16793 , \2839 );
xor \U$16595 ( \16795 , \16790 , \16794 );
xor \U$16596 ( \16796 , \16781 , \16795 );
xor \U$16597 ( \16797 , \16753 , \16796 );
xor \U$16598 ( \16798 , \16744 , \16797 );
xor \U$16599 ( \16799 , \16735 , \16798 );
and \U$16600 ( \16800 , \16511 , \16515 );
and \U$16601 ( \16801 , \16515 , \16520 );
and \U$16602 ( \16802 , \16511 , \16520 );
or \U$16603 ( \16803 , \16800 , \16801 , \16802 );
and \U$16604 ( \16804 , \16545 , \16559 );
and \U$16605 ( \16805 , \16559 , \16715 );
and \U$16606 ( \16806 , \16545 , \16715 );
or \U$16607 ( \16807 , \16804 , \16805 , \16806 );
xor \U$16608 ( \16808 , \16803 , \16807 );
and \U$16609 ( \16809 , \16588 , \16592 );
and \U$16610 ( \16810 , \16592 , \16597 );
and \U$16611 ( \16811 , \16588 , \16597 );
or \U$16612 ( \16812 , \16809 , \16810 , \16811 );
and \U$16613 ( \16813 , \16602 , \16603 );
and \U$16614 ( \16814 , \16603 , \16608 );
and \U$16615 ( \16815 , \16602 , \16608 );
or \U$16616 ( \16816 , \16813 , \16814 , \16815 );
xor \U$16617 ( \16817 , \16812 , \16816 );
and \U$16618 ( \16818 , \16614 , \16618 );
and \U$16619 ( \16819 , \16618 , \16623 );
and \U$16620 ( \16820 , \16614 , \16623 );
or \U$16621 ( \16821 , \16818 , \16819 , \16820 );
xor \U$16622 ( \16822 , \16817 , \16821 );
and \U$16623 ( \16823 , \16535 , \16539 );
and \U$16624 ( \16824 , \16539 , \16544 );
and \U$16625 ( \16825 , \16535 , \16544 );
or \U$16626 ( \16826 , \16823 , \16824 , \16825 );
and \U$16627 ( \16827 , \16564 , \16568 );
and \U$16628 ( \16828 , \16568 , \16583 );
and \U$16629 ( \16829 , \16564 , \16583 );
or \U$16630 ( \16830 , \16827 , \16828 , \16829 );
xor \U$16631 ( \16831 , \16826 , \16830 );
and \U$16632 ( \16832 , \16637 , \16668 );
and \U$16633 ( \16833 , \16668 , \16713 );
and \U$16634 ( \16834 , \16637 , \16713 );
or \U$16635 ( \16835 , \16832 , \16833 , \16834 );
xor \U$16636 ( \16836 , \16831 , \16835 );
xor \U$16637 ( \16837 , \16822 , \16836 );
and \U$16638 ( \16838 , \16598 , \16609 );
and \U$16639 ( \16839 , \16609 , \16624 );
and \U$16640 ( \16840 , \16598 , \16624 );
or \U$16641 ( \16841 , \16838 , \16839 , \16840 );
and \U$16642 ( \16842 , \16687 , \16691 );
and \U$16643 ( \16843 , \16691 , \16696 );
and \U$16644 ( \16844 , \16687 , \16696 );
or \U$16645 ( \16845 , \16842 , \16843 , \16844 );
and \U$16646 ( \16846 , \16627 , \16631 );
and \U$16647 ( \16847 , \16631 , \16636 );
and \U$16648 ( \16848 , \16627 , \16636 );
or \U$16649 ( \16849 , \16846 , \16847 , \16848 );
xor \U$16650 ( \16850 , \16845 , \16849 );
and \U$16651 ( \16851 , \16573 , \16577 );
and \U$16652 ( \16852 , \16577 , \16582 );
and \U$16653 ( \16853 , \16573 , \16582 );
or \U$16654 ( \16854 , \16851 , \16852 , \16853 );
xor \U$16655 ( \16855 , \16850 , \16854 );
xor \U$16656 ( \16856 , \16841 , \16855 );
and \U$16657 ( \16857 , \16673 , \16677 );
and \U$16658 ( \16858 , \16677 , \16682 );
and \U$16659 ( \16859 , \16673 , \16682 );
or \U$16660 ( \16860 , \16857 , \16858 , \16859 );
and \U$16661 ( \16861 , \16657 , \16661 );
and \U$16662 ( \16862 , \16661 , \16666 );
and \U$16663 ( \16863 , \16657 , \16666 );
or \U$16664 ( \16864 , \16861 , \16862 , \16863 );
xor \U$16665 ( \16865 , \16860 , \16864 );
and \U$16666 ( \16866 , \16702 , \16706 );
and \U$16667 ( \16867 , \16706 , \16711 );
and \U$16668 ( \16868 , \16702 , \16711 );
or \U$16669 ( \16869 , \16866 , \16867 , \16868 );
xor \U$16670 ( \16870 , \16865 , \16869 );
and \U$16671 ( \16871 , \3037 , \7489 );
and \U$16672 ( \16872 , \3143 , \7137 );
nor \U$16673 ( \16873 , \16871 , \16872 );
xnor \U$16674 ( \16874 , \16873 , \7142 );
and \U$16675 ( \16875 , \2757 , \8019 );
and \U$16676 ( \16876 , \2826 , \7830 );
nor \U$16677 ( \16877 , \16875 , \16876 );
xnor \U$16678 ( \16878 , \16877 , \7713 );
xor \U$16679 ( \16879 , \16874 , \16878 );
and \U$16680 ( \16880 , \2366 , \8540 );
and \U$16681 ( \16881 , \2521 , \8292 );
nor \U$16682 ( \16882 , \16880 , \16881 );
xnor \U$16683 ( \16883 , \16882 , \8297 );
xor \U$16684 ( \16884 , \16879 , \16883 );
and \U$16685 ( \16885 , \4160 , \5996 );
and \U$16686 ( \16886 , \4364 , \5695 );
nor \U$16687 ( \16887 , \16885 , \16886 );
xnor \U$16688 ( \16888 , \16887 , \5687 );
and \U$16689 ( \16889 , \3736 , \6401 );
and \U$16690 ( \16890 , \3912 , \6143 );
nor \U$16691 ( \16891 , \16889 , \16890 );
xnor \U$16692 ( \16892 , \16891 , \6148 );
xor \U$16693 ( \16893 , \16888 , \16892 );
and \U$16694 ( \16894 , \3395 , \7055 );
and \U$16695 ( \16895 , \3646 , \6675 );
nor \U$16696 ( \16896 , \16894 , \16895 );
xnor \U$16697 ( \16897 , \16896 , \6680 );
xor \U$16698 ( \16898 , \16893 , \16897 );
xor \U$16699 ( \16899 , \16884 , \16898 );
and \U$16700 ( \16900 , \5469 , \4581 );
and \U$16701 ( \16901 , \5674 , \4424 );
nor \U$16702 ( \16902 , \16900 , \16901 );
xnor \U$16703 ( \16903 , \16902 , \4377 );
and \U$16704 ( \16904 , \4922 , \5011 );
and \U$16705 ( \16905 , \5156 , \4878 );
nor \U$16706 ( \16906 , \16904 , \16905 );
xnor \U$16707 ( \16907 , \16906 , \4762 );
xor \U$16708 ( \16908 , \16903 , \16907 );
and \U$16709 ( \16909 , \4654 , \5485 );
and \U$16710 ( \16910 , \4749 , \5275 );
nor \U$16711 ( \16911 , \16909 , \16910 );
xnor \U$16712 ( \16912 , \16911 , \5169 );
xor \U$16713 ( \16913 , \16908 , \16912 );
xor \U$16714 ( \16914 , \16899 , \16913 );
xor \U$16715 ( \16915 , \16870 , \16914 );
and \U$16716 ( \16916 , \16642 , \16646 );
and \U$16717 ( \16917 , \16646 , \16651 );
and \U$16718 ( \16918 , \16642 , \16651 );
or \U$16719 ( \16919 , \16916 , \16917 , \16918 );
and \U$16720 ( \16920 , \2090 , \9333 );
and \U$16721 ( \16921 , \2182 , \9006 );
nor \U$16722 ( \16922 , \16920 , \16921 );
xnor \U$16723 ( \16923 , \16922 , \8848 );
and \U$16724 ( \16924 , \1802 , \9765 );
and \U$16725 ( \16925 , \1948 , \9644 );
nor \U$16726 ( \16926 , \16924 , \16925 );
xnor \U$16727 ( \16927 , \16926 , \9478 );
xor \U$16728 ( \16928 , \16923 , \16927 );
and \U$16729 ( \16929 , \1601 , \10408 );
and \U$16730 ( \16930 , \1684 , \10116 );
nor \U$16731 ( \16931 , \16929 , \16930 );
xnor \U$16732 ( \16932 , \16931 , \10121 );
xor \U$16733 ( \16933 , \16928 , \16932 );
xor \U$16734 ( \16934 , \16919 , \16933 );
and \U$16735 ( \16935 , \1484 , \10118 );
not \U$16736 ( \16936 , \16935 );
xor \U$16737 ( \16937 , \16934 , \16936 );
xor \U$16738 ( \16938 , \16915 , \16937 );
xor \U$16739 ( \16939 , \16856 , \16938 );
xor \U$16740 ( \16940 , \16837 , \16939 );
xor \U$16741 ( \16941 , \16808 , \16940 );
xor \U$16742 ( \16942 , \16799 , \16941 );
xor \U$16743 ( \16943 , \16731 , \16942 );
and \U$16744 ( \16944 , \16503 , \16718 );
xor \U$16745 ( \16945 , \16943 , \16944 );
and \U$16746 ( \16946 , \16719 , \16720 );
and \U$16747 ( \16947 , \16721 , \16724 );
or \U$16748 ( \16948 , \16946 , \16947 );
xor \U$16749 ( \16949 , \16945 , \16948 );
buf g54ef_GF_PartitionCandidate( \16950_nG54ef , \16949 );
buf \U$16750 ( \16951 , \16950_nG54ef );
and \U$16751 ( \16952 , \16735 , \16798 );
and \U$16752 ( \16953 , \16798 , \16941 );
and \U$16753 ( \16954 , \16735 , \16941 );
or \U$16754 ( \16955 , \16952 , \16953 , \16954 );
and \U$16755 ( \16956 , \16803 , \16807 );
and \U$16756 ( \16957 , \16807 , \16940 );
and \U$16757 ( \16958 , \16803 , \16940 );
or \U$16758 ( \16959 , \16956 , \16957 , \16958 );
and \U$16759 ( \16960 , \16826 , \16830 );
and \U$16760 ( \16961 , \16830 , \16835 );
and \U$16761 ( \16962 , \16826 , \16835 );
or \U$16762 ( \16963 , \16960 , \16961 , \16962 );
and \U$16763 ( \16964 , \16841 , \16855 );
and \U$16764 ( \16965 , \16855 , \16938 );
and \U$16765 ( \16966 , \16841 , \16938 );
or \U$16766 ( \16967 , \16964 , \16965 , \16966 );
xor \U$16767 ( \16968 , \16963 , \16967 );
and \U$16768 ( \16969 , \16884 , \16898 );
and \U$16769 ( \16970 , \16898 , \16913 );
and \U$16770 ( \16971 , \16884 , \16913 );
or \U$16771 ( \16972 , \16969 , \16970 , \16971 );
and \U$16772 ( \16973 , \16767 , \16780 );
and \U$16773 ( \16974 , \16780 , \16795 );
and \U$16774 ( \16975 , \16767 , \16795 );
or \U$16775 ( \16976 , \16973 , \16974 , \16975 );
xor \U$16776 ( \16977 , \16972 , \16976 );
not \U$16777 ( \16978 , \1436 );
and \U$16778 ( \16979 , \10206 , \1824 );
and \U$16779 ( \16980 , \10584 , \1739 );
nor \U$16780 ( \16981 , \16979 , \16980 );
xnor \U$16781 ( \16982 , \16981 , \1697 );
xor \U$16782 ( \16983 , \16978 , \16982 );
and \U$16783 ( \16984 , \9465 , \2121 );
and \U$16784 ( \16985 , \9897 , \2008 );
nor \U$16785 ( \16986 , \16984 , \16985 );
xnor \U$16786 ( \16987 , \16986 , \1961 );
xor \U$16787 ( \16988 , \16983 , \16987 );
xor \U$16788 ( \16989 , \16977 , \16988 );
xor \U$16789 ( \16990 , \16968 , \16989 );
xor \U$16790 ( \16991 , \16959 , \16990 );
and \U$16791 ( \16992 , \16739 , \16743 );
and \U$16792 ( \16993 , \16743 , \16797 );
and \U$16793 ( \16994 , \16739 , \16797 );
or \U$16794 ( \16995 , \16992 , \16993 , \16994 );
and \U$16795 ( \16996 , \16822 , \16836 );
and \U$16796 ( \16997 , \16836 , \16939 );
and \U$16797 ( \16998 , \16822 , \16939 );
or \U$16798 ( \16999 , \16996 , \16997 , \16998 );
xor \U$16799 ( \17000 , \16995 , \16999 );
and \U$16800 ( \17001 , \16845 , \16849 );
and \U$16801 ( \17002 , \16849 , \16854 );
and \U$16802 ( \17003 , \16845 , \16854 );
or \U$16803 ( \17004 , \17001 , \17002 , \17003 );
and \U$16804 ( \17005 , \16860 , \16864 );
and \U$16805 ( \17006 , \16864 , \16869 );
and \U$16806 ( \17007 , \16860 , \16869 );
or \U$16807 ( \17008 , \17005 , \17006 , \17007 );
xor \U$16808 ( \17009 , \17004 , \17008 );
and \U$16809 ( \17010 , \16919 , \16933 );
and \U$16810 ( \17011 , \16933 , \16936 );
and \U$16811 ( \17012 , \16919 , \16936 );
or \U$16812 ( \17013 , \17010 , \17011 , \17012 );
xor \U$16813 ( \17014 , \17009 , \17013 );
and \U$16814 ( \17015 , \16812 , \16816 );
and \U$16815 ( \17016 , \16816 , \16821 );
and \U$16816 ( \17017 , \16812 , \16821 );
or \U$16817 ( \17018 , \17015 , \17016 , \17017 );
and \U$16818 ( \17019 , \16748 , \16752 );
and \U$16819 ( \17020 , \16752 , \16796 );
and \U$16820 ( \17021 , \16748 , \16796 );
or \U$16821 ( \17022 , \17019 , \17020 , \17021 );
xor \U$16822 ( \17023 , \17018 , \17022 );
and \U$16823 ( \17024 , \16870 , \16914 );
and \U$16824 ( \17025 , \16914 , \16937 );
and \U$16825 ( \17026 , \16870 , \16937 );
or \U$16826 ( \17027 , \17024 , \17025 , \17026 );
xor \U$16827 ( \17028 , \17023 , \17027 );
xor \U$16828 ( \17029 , \17014 , \17028 );
and \U$16829 ( \17030 , \16757 , \16761 );
and \U$16830 ( \17031 , \16761 , \16766 );
and \U$16831 ( \17032 , \16757 , \16766 );
or \U$16832 ( \17033 , \17030 , \17031 , \17032 );
and \U$16833 ( \17034 , \16770 , \16774 );
and \U$16834 ( \17035 , \16774 , \16779 );
and \U$16835 ( \17036 , \16770 , \16779 );
or \U$16836 ( \17037 , \17034 , \17035 , \17036 );
xor \U$16837 ( \17038 , \17033 , \17037 );
and \U$16838 ( \17039 , \16785 , \16789 );
and \U$16839 ( \17040 , \16789 , \16794 );
and \U$16840 ( \17041 , \16785 , \16794 );
or \U$16841 ( \17042 , \17039 , \17040 , \17041 );
xor \U$16842 ( \17043 , \17038 , \17042 );
and \U$16843 ( \17044 , \16874 , \16878 );
and \U$16844 ( \17045 , \16878 , \16883 );
and \U$16845 ( \17046 , \16874 , \16883 );
or \U$16846 ( \17047 , \17044 , \17045 , \17046 );
and \U$16847 ( \17048 , \16888 , \16892 );
and \U$16848 ( \17049 , \16892 , \16897 );
and \U$16849 ( \17050 , \16888 , \16897 );
or \U$16850 ( \17051 , \17048 , \17049 , \17050 );
xor \U$16851 ( \17052 , \17047 , \17051 );
and \U$16852 ( \17053 , \16903 , \16907 );
and \U$16853 ( \17054 , \16907 , \16912 );
and \U$16854 ( \17055 , \16903 , \16912 );
or \U$16855 ( \17056 , \17053 , \17054 , \17055 );
xor \U$16856 ( \17057 , \17052 , \17056 );
xor \U$16857 ( \17058 , \17043 , \17057 );
and \U$16858 ( \17059 , \16923 , \16927 );
and \U$16859 ( \17060 , \16927 , \16932 );
and \U$16860 ( \17061 , \16923 , \16932 );
or \U$16861 ( \17062 , \17059 , \17060 , \17061 );
buf \U$16862 ( \17063 , \16935 );
xor \U$16863 ( \17064 , \17062 , \17063 );
and \U$16864 ( \17065 , \1601 , \10118 );
xor \U$16865 ( \17066 , \17064 , \17065 );
and \U$16866 ( \17067 , \3143 , \7489 );
and \U$16867 ( \17068 , \3395 , \7137 );
nor \U$16868 ( \17069 , \17067 , \17068 );
xnor \U$16869 ( \17070 , \17069 , \7142 );
and \U$16870 ( \17071 , \2826 , \8019 );
and \U$16871 ( \17072 , \3037 , \7830 );
nor \U$16872 ( \17073 , \17071 , \17072 );
xnor \U$16873 ( \17074 , \17073 , \7713 );
xor \U$16874 ( \17075 , \17070 , \17074 );
and \U$16875 ( \17076 , \2521 , \8540 );
and \U$16876 ( \17077 , \2757 , \8292 );
nor \U$16877 ( \17078 , \17076 , \17077 );
xnor \U$16878 ( \17079 , \17078 , \8297 );
xor \U$16879 ( \17080 , \17075 , \17079 );
and \U$16880 ( \17081 , \4364 , \5996 );
and \U$16881 ( \17082 , \4654 , \5695 );
nor \U$16882 ( \17083 , \17081 , \17082 );
xnor \U$16883 ( \17084 , \17083 , \5687 );
and \U$16884 ( \17085 , \3912 , \6401 );
and \U$16885 ( \17086 , \4160 , \6143 );
nor \U$16886 ( \17087 , \17085 , \17086 );
xnor \U$16887 ( \17088 , \17087 , \6148 );
xor \U$16888 ( \17089 , \17084 , \17088 );
and \U$16889 ( \17090 , \3646 , \7055 );
and \U$16890 ( \17091 , \3736 , \6675 );
nor \U$16891 ( \17092 , \17090 , \17091 );
xnor \U$16892 ( \17093 , \17092 , \6680 );
xor \U$16893 ( \17094 , \17089 , \17093 );
xor \U$16894 ( \17095 , \17080 , \17094 );
and \U$16895 ( \17096 , \2182 , \9333 );
and \U$16896 ( \17097 , \2366 , \9006 );
nor \U$16897 ( \17098 , \17096 , \17097 );
xnor \U$16898 ( \17099 , \17098 , \8848 );
and \U$16899 ( \17100 , \1948 , \9765 );
and \U$16900 ( \17101 , \2090 , \9644 );
nor \U$16901 ( \17102 , \17100 , \17101 );
xnor \U$16902 ( \17103 , \17102 , \9478 );
xor \U$16903 ( \17104 , \17099 , \17103 );
and \U$16904 ( \17105 , \1684 , \10408 );
and \U$16905 ( \17106 , \1802 , \10116 );
nor \U$16906 ( \17107 , \17105 , \17106 );
xnor \U$16907 ( \17108 , \17107 , \10121 );
xor \U$16908 ( \17109 , \17104 , \17108 );
xor \U$16909 ( \17110 , \17095 , \17109 );
xor \U$16910 ( \17111 , \17066 , \17110 );
and \U$16911 ( \17112 , \7231 , \3357 );
and \U$16912 ( \17113 , \7556 , \3255 );
nor \U$16913 ( \17114 , \17112 , \17113 );
xnor \U$16914 ( \17115 , \17114 , \3156 );
and \U$16915 ( \17116 , \6790 , \3813 );
and \U$16916 ( \17117 , \6945 , \3557 );
nor \U$16917 ( \17118 , \17116 , \17117 );
xnor \U$16918 ( \17119 , \17118 , \3562 );
xor \U$16919 ( \17120 , \17115 , \17119 );
and \U$16920 ( \17121 , \6281 , \4132 );
and \U$16921 ( \17122 , \6514 , \4012 );
nor \U$16922 ( \17123 , \17121 , \17122 );
xnor \U$16923 ( \17124 , \17123 , \3925 );
xor \U$16924 ( \17125 , \17120 , \17124 );
and \U$16925 ( \17126 , \5674 , \4581 );
and \U$16926 ( \17127 , \6030 , \4424 );
nor \U$16927 ( \17128 , \17126 , \17127 );
xnor \U$16928 ( \17129 , \17128 , \4377 );
and \U$16929 ( \17130 , \5156 , \5011 );
and \U$16930 ( \17131 , \5469 , \4878 );
nor \U$16931 ( \17132 , \17130 , \17131 );
xnor \U$16932 ( \17133 , \17132 , \4762 );
xor \U$16933 ( \17134 , \17129 , \17133 );
and \U$16934 ( \17135 , \4749 , \5485 );
and \U$16935 ( \17136 , \4922 , \5275 );
nor \U$16936 ( \17137 , \17135 , \17136 );
xnor \U$16937 ( \17138 , \17137 , \5169 );
xor \U$16938 ( \17139 , \17134 , \17138 );
xor \U$16939 ( \17140 , \17125 , \17139 );
and \U$16940 ( \17141 , \8835 , \2400 );
and \U$16941 ( \17142 , \9169 , \2246 );
nor \U$16942 ( \17143 , \17141 , \17142 );
xnor \U$16943 ( \17144 , \17143 , \2195 );
and \U$16944 ( \17145 , \8349 , \2669 );
and \U$16945 ( \17146 , \8652 , \2538 );
nor \U$16946 ( \17147 , \17145 , \17146 );
xnor \U$16947 ( \17148 , \17147 , \2534 );
xor \U$16948 ( \17149 , \17144 , \17148 );
and \U$16949 ( \17150 , \7700 , \3103 );
and \U$16950 ( \17151 , \8057 , \2934 );
nor \U$16951 ( \17152 , \17150 , \17151 );
xnor \U$16952 ( \17153 , \17152 , \2839 );
xor \U$16953 ( \17154 , \17149 , \17153 );
xor \U$16954 ( \17155 , \17140 , \17154 );
xor \U$16955 ( \17156 , \17111 , \17155 );
xor \U$16956 ( \17157 , \17058 , \17156 );
xor \U$16957 ( \17158 , \17029 , \17157 );
xor \U$16958 ( \17159 , \17000 , \17158 );
xor \U$16959 ( \17160 , \16991 , \17159 );
xor \U$16960 ( \17161 , \16955 , \17160 );
and \U$16961 ( \17162 , \16731 , \16942 );
xor \U$16962 ( \17163 , \17161 , \17162 );
and \U$16963 ( \17164 , \16943 , \16944 );
and \U$16964 ( \17165 , \16945 , \16948 );
or \U$16965 ( \17166 , \17164 , \17165 );
xor \U$16966 ( \17167 , \17163 , \17166 );
buf g54ed_GF_PartitionCandidate( \17168_nG54ed , \17167 );
buf \U$16967 ( \17169 , \17168_nG54ed );
and \U$16968 ( \17170 , \16959 , \16990 );
and \U$16969 ( \17171 , \16990 , \17159 );
and \U$16970 ( \17172 , \16959 , \17159 );
or \U$16971 ( \17173 , \17170 , \17171 , \17172 );
and \U$16972 ( \17174 , \16995 , \16999 );
and \U$16973 ( \17175 , \16999 , \17158 );
and \U$16974 ( \17176 , \16995 , \17158 );
or \U$16975 ( \17177 , \17174 , \17175 , \17176 );
and \U$16976 ( \17178 , \16963 , \16967 );
and \U$16977 ( \17179 , \16967 , \16989 );
and \U$16978 ( \17180 , \16963 , \16989 );
or \U$16979 ( \17181 , \17178 , \17179 , \17180 );
and \U$16980 ( \17182 , \17014 , \17028 );
and \U$16981 ( \17183 , \17028 , \17157 );
and \U$16982 ( \17184 , \17014 , \17157 );
or \U$16983 ( \17185 , \17182 , \17183 , \17184 );
xor \U$16984 ( \17186 , \17181 , \17185 );
and \U$16985 ( \17187 , \17115 , \17119 );
and \U$16986 ( \17188 , \17119 , \17124 );
and \U$16987 ( \17189 , \17115 , \17124 );
or \U$16988 ( \17190 , \17187 , \17188 , \17189 );
and \U$16989 ( \17191 , \16978 , \16982 );
and \U$16990 ( \17192 , \16982 , \16987 );
and \U$16991 ( \17193 , \16978 , \16987 );
or \U$16992 ( \17194 , \17191 , \17192 , \17193 );
xor \U$16993 ( \17195 , \17190 , \17194 );
and \U$16994 ( \17196 , \17144 , \17148 );
and \U$16995 ( \17197 , \17148 , \17153 );
and \U$16996 ( \17198 , \17144 , \17153 );
or \U$16997 ( \17199 , \17196 , \17197 , \17198 );
xor \U$16998 ( \17200 , \17195 , \17199 );
and \U$16999 ( \17201 , \17080 , \17094 );
and \U$17000 ( \17202 , \17094 , \17109 );
and \U$17001 ( \17203 , \17080 , \17109 );
or \U$17002 ( \17204 , \17201 , \17202 , \17203 );
and \U$17003 ( \17205 , \17125 , \17139 );
and \U$17004 ( \17206 , \17139 , \17154 );
and \U$17005 ( \17207 , \17125 , \17154 );
or \U$17006 ( \17208 , \17205 , \17206 , \17207 );
xor \U$17007 ( \17209 , \17204 , \17208 );
and \U$17008 ( \17210 , \10584 , \1824 );
not \U$17009 ( \17211 , \17210 );
xnor \U$17010 ( \17212 , \17211 , \1697 );
and \U$17011 ( \17213 , \9897 , \2121 );
and \U$17012 ( \17214 , \10206 , \2008 );
nor \U$17013 ( \17215 , \17213 , \17214 );
xnor \U$17014 ( \17216 , \17215 , \1961 );
xor \U$17015 ( \17217 , \17212 , \17216 );
and \U$17016 ( \17218 , \9169 , \2400 );
and \U$17017 ( \17219 , \9465 , \2246 );
nor \U$17018 ( \17220 , \17218 , \17219 );
xnor \U$17019 ( \17221 , \17220 , \2195 );
xor \U$17020 ( \17222 , \17217 , \17221 );
and \U$17021 ( \17223 , \8652 , \2669 );
and \U$17022 ( \17224 , \8835 , \2538 );
nor \U$17023 ( \17225 , \17223 , \17224 );
xnor \U$17024 ( \17226 , \17225 , \2534 );
and \U$17025 ( \17227 , \8057 , \3103 );
and \U$17026 ( \17228 , \8349 , \2934 );
nor \U$17027 ( \17229 , \17227 , \17228 );
xnor \U$17028 ( \17230 , \17229 , \2839 );
xor \U$17029 ( \17231 , \17226 , \17230 );
and \U$17030 ( \17232 , \7556 , \3357 );
and \U$17031 ( \17233 , \7700 , \3255 );
nor \U$17032 ( \17234 , \17232 , \17233 );
xnor \U$17033 ( \17235 , \17234 , \3156 );
xor \U$17034 ( \17236 , \17231 , \17235 );
xor \U$17035 ( \17237 , \17222 , \17236 );
and \U$17036 ( \17238 , \6945 , \3813 );
and \U$17037 ( \17239 , \7231 , \3557 );
nor \U$17038 ( \17240 , \17238 , \17239 );
xnor \U$17039 ( \17241 , \17240 , \3562 );
and \U$17040 ( \17242 , \6514 , \4132 );
and \U$17041 ( \17243 , \6790 , \4012 );
nor \U$17042 ( \17244 , \17242 , \17243 );
xnor \U$17043 ( \17245 , \17244 , \3925 );
xor \U$17044 ( \17246 , \17241 , \17245 );
and \U$17045 ( \17247 , \6030 , \4581 );
and \U$17046 ( \17248 , \6281 , \4424 );
nor \U$17047 ( \17249 , \17247 , \17248 );
xnor \U$17048 ( \17250 , \17249 , \4377 );
xor \U$17049 ( \17251 , \17246 , \17250 );
xor \U$17050 ( \17252 , \17237 , \17251 );
xor \U$17051 ( \17253 , \17209 , \17252 );
xor \U$17052 ( \17254 , \17200 , \17253 );
and \U$17053 ( \17255 , \17070 , \17074 );
and \U$17054 ( \17256 , \17074 , \17079 );
and \U$17055 ( \17257 , \17070 , \17079 );
or \U$17056 ( \17258 , \17255 , \17256 , \17257 );
and \U$17057 ( \17259 , \17129 , \17133 );
and \U$17058 ( \17260 , \17133 , \17138 );
and \U$17059 ( \17261 , \17129 , \17138 );
or \U$17060 ( \17262 , \17259 , \17260 , \17261 );
xor \U$17061 ( \17263 , \17258 , \17262 );
and \U$17062 ( \17264 , \17084 , \17088 );
and \U$17063 ( \17265 , \17088 , \17093 );
and \U$17064 ( \17266 , \17084 , \17093 );
or \U$17065 ( \17267 , \17264 , \17265 , \17266 );
xor \U$17066 ( \17268 , \17263 , \17267 );
and \U$17067 ( \17269 , \3037 , \8019 );
and \U$17068 ( \17270 , \3143 , \7830 );
nor \U$17069 ( \17271 , \17269 , \17270 );
xnor \U$17070 ( \17272 , \17271 , \7713 );
and \U$17071 ( \17273 , \2757 , \8540 );
and \U$17072 ( \17274 , \2826 , \8292 );
nor \U$17073 ( \17275 , \17273 , \17274 );
xnor \U$17074 ( \17276 , \17275 , \8297 );
xor \U$17075 ( \17277 , \17272 , \17276 );
and \U$17076 ( \17278 , \2366 , \9333 );
and \U$17077 ( \17279 , \2521 , \9006 );
nor \U$17078 ( \17280 , \17278 , \17279 );
xnor \U$17079 ( \17281 , \17280 , \8848 );
xor \U$17080 ( \17282 , \17277 , \17281 );
and \U$17081 ( \17283 , \5469 , \5011 );
and \U$17082 ( \17284 , \5674 , \4878 );
nor \U$17083 ( \17285 , \17283 , \17284 );
xnor \U$17084 ( \17286 , \17285 , \4762 );
and \U$17085 ( \17287 , \4922 , \5485 );
and \U$17086 ( \17288 , \5156 , \5275 );
nor \U$17087 ( \17289 , \17287 , \17288 );
xnor \U$17088 ( \17290 , \17289 , \5169 );
xor \U$17089 ( \17291 , \17286 , \17290 );
and \U$17090 ( \17292 , \4654 , \5996 );
and \U$17091 ( \17293 , \4749 , \5695 );
nor \U$17092 ( \17294 , \17292 , \17293 );
xnor \U$17093 ( \17295 , \17294 , \5687 );
xor \U$17094 ( \17296 , \17291 , \17295 );
xor \U$17095 ( \17297 , \17282 , \17296 );
and \U$17096 ( \17298 , \4160 , \6401 );
and \U$17097 ( \17299 , \4364 , \6143 );
nor \U$17098 ( \17300 , \17298 , \17299 );
xnor \U$17099 ( \17301 , \17300 , \6148 );
and \U$17100 ( \17302 , \3736 , \7055 );
and \U$17101 ( \17303 , \3912 , \6675 );
nor \U$17102 ( \17304 , \17302 , \17303 );
xnor \U$17103 ( \17305 , \17304 , \6680 );
xor \U$17104 ( \17306 , \17301 , \17305 );
and \U$17105 ( \17307 , \3395 , \7489 );
and \U$17106 ( \17308 , \3646 , \7137 );
nor \U$17107 ( \17309 , \17307 , \17308 );
xnor \U$17108 ( \17310 , \17309 , \7142 );
xor \U$17109 ( \17311 , \17306 , \17310 );
xor \U$17110 ( \17312 , \17297 , \17311 );
xor \U$17111 ( \17313 , \17268 , \17312 );
and \U$17112 ( \17314 , \17099 , \17103 );
and \U$17113 ( \17315 , \17103 , \17108 );
and \U$17114 ( \17316 , \17099 , \17108 );
or \U$17115 ( \17317 , \17314 , \17315 , \17316 );
and \U$17116 ( \17318 , \2090 , \9765 );
and \U$17117 ( \17319 , \2182 , \9644 );
nor \U$17118 ( \17320 , \17318 , \17319 );
xnor \U$17119 ( \17321 , \17320 , \9478 );
and \U$17120 ( \17322 , \1802 , \10408 );
and \U$17121 ( \17323 , \1948 , \10116 );
nor \U$17122 ( \17324 , \17322 , \17323 );
xnor \U$17123 ( \17325 , \17324 , \10121 );
xor \U$17124 ( \17326 , \17321 , \17325 );
and \U$17125 ( \17327 , \1684 , \10118 );
xor \U$17126 ( \17328 , \17326 , \17327 );
xnor \U$17127 ( \17329 , \17317 , \17328 );
xor \U$17128 ( \17330 , \17313 , \17329 );
xor \U$17129 ( \17331 , \17254 , \17330 );
xor \U$17130 ( \17332 , \17186 , \17331 );
xor \U$17131 ( \17333 , \17177 , \17332 );
and \U$17132 ( \17334 , \17004 , \17008 );
and \U$17133 ( \17335 , \17008 , \17013 );
and \U$17134 ( \17336 , \17004 , \17013 );
or \U$17135 ( \17337 , \17334 , \17335 , \17336 );
and \U$17136 ( \17338 , \16972 , \16976 );
and \U$17137 ( \17339 , \16976 , \16988 );
and \U$17138 ( \17340 , \16972 , \16988 );
or \U$17139 ( \17341 , \17338 , \17339 , \17340 );
xor \U$17140 ( \17342 , \17337 , \17341 );
and \U$17141 ( \17343 , \17066 , \17110 );
and \U$17142 ( \17344 , \17110 , \17155 );
and \U$17143 ( \17345 , \17066 , \17155 );
or \U$17144 ( \17346 , \17343 , \17344 , \17345 );
xor \U$17145 ( \17347 , \17342 , \17346 );
and \U$17146 ( \17348 , \17018 , \17022 );
and \U$17147 ( \17349 , \17022 , \17027 );
and \U$17148 ( \17350 , \17018 , \17027 );
or \U$17149 ( \17351 , \17348 , \17349 , \17350 );
and \U$17150 ( \17352 , \17043 , \17057 );
and \U$17151 ( \17353 , \17057 , \17156 );
and \U$17152 ( \17354 , \17043 , \17156 );
or \U$17153 ( \17355 , \17352 , \17353 , \17354 );
xor \U$17154 ( \17356 , \17351 , \17355 );
and \U$17155 ( \17357 , \17062 , \17063 );
and \U$17156 ( \17358 , \17063 , \17065 );
and \U$17157 ( \17359 , \17062 , \17065 );
or \U$17158 ( \17360 , \17357 , \17358 , \17359 );
and \U$17159 ( \17361 , \17033 , \17037 );
and \U$17160 ( \17362 , \17037 , \17042 );
and \U$17161 ( \17363 , \17033 , \17042 );
or \U$17162 ( \17364 , \17361 , \17362 , \17363 );
xor \U$17163 ( \17365 , \17360 , \17364 );
and \U$17164 ( \17366 , \17047 , \17051 );
and \U$17165 ( \17367 , \17051 , \17056 );
and \U$17166 ( \17368 , \17047 , \17056 );
or \U$17167 ( \17369 , \17366 , \17367 , \17368 );
xor \U$17168 ( \17370 , \17365 , \17369 );
xor \U$17169 ( \17371 , \17356 , \17370 );
xor \U$17170 ( \17372 , \17347 , \17371 );
xor \U$17171 ( \17373 , \17333 , \17372 );
xor \U$17172 ( \17374 , \17173 , \17373 );
and \U$17173 ( \17375 , \16955 , \17160 );
xor \U$17174 ( \17376 , \17374 , \17375 );
and \U$17175 ( \17377 , \17161 , \17162 );
and \U$17176 ( \17378 , \17163 , \17166 );
or \U$17177 ( \17379 , \17377 , \17378 );
xor \U$17178 ( \17380 , \17376 , \17379 );
buf g54eb_GF_PartitionCandidate( \17381_nG54eb , \17380 );
buf \U$17179 ( \17382 , \17381_nG54eb );
and \U$17180 ( \17383 , \17177 , \17332 );
and \U$17181 ( \17384 , \17332 , \17372 );
and \U$17182 ( \17385 , \17177 , \17372 );
or \U$17183 ( \17386 , \17383 , \17384 , \17385 );
and \U$17184 ( \17387 , \17181 , \17185 );
and \U$17185 ( \17388 , \17185 , \17331 );
and \U$17186 ( \17389 , \17181 , \17331 );
or \U$17187 ( \17390 , \17387 , \17388 , \17389 );
and \U$17188 ( \17391 , \17347 , \17371 );
xor \U$17189 ( \17392 , \17390 , \17391 );
and \U$17190 ( \17393 , \17351 , \17355 );
and \U$17191 ( \17394 , \17355 , \17370 );
and \U$17192 ( \17395 , \17351 , \17370 );
or \U$17193 ( \17396 , \17393 , \17394 , \17395 );
and \U$17194 ( \17397 , \17337 , \17341 );
and \U$17195 ( \17398 , \17341 , \17346 );
and \U$17196 ( \17399 , \17337 , \17346 );
or \U$17197 ( \17400 , \17397 , \17398 , \17399 );
and \U$17198 ( \17401 , \17200 , \17253 );
and \U$17199 ( \17402 , \17253 , \17330 );
and \U$17200 ( \17403 , \17200 , \17330 );
or \U$17201 ( \17404 , \17401 , \17402 , \17403 );
xor \U$17202 ( \17405 , \17400 , \17404 );
and \U$17203 ( \17406 , \17282 , \17296 );
and \U$17204 ( \17407 , \17296 , \17311 );
and \U$17205 ( \17408 , \17282 , \17311 );
or \U$17206 ( \17409 , \17406 , \17407 , \17408 );
and \U$17207 ( \17410 , \17222 , \17236 );
and \U$17208 ( \17411 , \17236 , \17251 );
and \U$17209 ( \17412 , \17222 , \17251 );
or \U$17210 ( \17413 , \17410 , \17411 , \17412 );
xor \U$17211 ( \17414 , \17409 , \17413 );
and \U$17212 ( \17415 , \8835 , \2669 );
and \U$17213 ( \17416 , \9169 , \2538 );
nor \U$17214 ( \17417 , \17415 , \17416 );
xnor \U$17215 ( \17418 , \17417 , \2534 );
and \U$17216 ( \17419 , \8349 , \3103 );
and \U$17217 ( \17420 , \8652 , \2934 );
nor \U$17218 ( \17421 , \17419 , \17420 );
xnor \U$17219 ( \17422 , \17421 , \2839 );
xor \U$17220 ( \17423 , \17418 , \17422 );
and \U$17221 ( \17424 , \7700 , \3357 );
and \U$17222 ( \17425 , \8057 , \3255 );
nor \U$17223 ( \17426 , \17424 , \17425 );
xnor \U$17224 ( \17427 , \17426 , \3156 );
xor \U$17225 ( \17428 , \17423 , \17427 );
xor \U$17226 ( \17429 , \17414 , \17428 );
xor \U$17227 ( \17430 , \17405 , \17429 );
xor \U$17228 ( \17431 , \17396 , \17430 );
and \U$17229 ( \17432 , \17190 , \17194 );
and \U$17230 ( \17433 , \17194 , \17199 );
and \U$17231 ( \17434 , \17190 , \17199 );
or \U$17232 ( \17435 , \17432 , \17433 , \17434 );
and \U$17233 ( \17436 , \17258 , \17262 );
and \U$17234 ( \17437 , \17262 , \17267 );
and \U$17235 ( \17438 , \17258 , \17267 );
or \U$17236 ( \17439 , \17436 , \17437 , \17438 );
xor \U$17237 ( \17440 , \17435 , \17439 );
or \U$17238 ( \17441 , \17317 , \17328 );
xor \U$17239 ( \17442 , \17440 , \17441 );
and \U$17240 ( \17443 , \17360 , \17364 );
and \U$17241 ( \17444 , \17364 , \17369 );
and \U$17242 ( \17445 , \17360 , \17369 );
or \U$17243 ( \17446 , \17443 , \17444 , \17445 );
and \U$17244 ( \17447 , \17204 , \17208 );
and \U$17245 ( \17448 , \17208 , \17252 );
and \U$17246 ( \17449 , \17204 , \17252 );
or \U$17247 ( \17450 , \17447 , \17448 , \17449 );
xor \U$17248 ( \17451 , \17446 , \17450 );
and \U$17249 ( \17452 , \17268 , \17312 );
and \U$17250 ( \17453 , \17312 , \17329 );
and \U$17251 ( \17454 , \17268 , \17329 );
or \U$17252 ( \17455 , \17452 , \17453 , \17454 );
xor \U$17253 ( \17456 , \17451 , \17455 );
xor \U$17254 ( \17457 , \17442 , \17456 );
and \U$17255 ( \17458 , \17212 , \17216 );
and \U$17256 ( \17459 , \17216 , \17221 );
and \U$17257 ( \17460 , \17212 , \17221 );
or \U$17258 ( \17461 , \17458 , \17459 , \17460 );
and \U$17259 ( \17462 , \17226 , \17230 );
and \U$17260 ( \17463 , \17230 , \17235 );
and \U$17261 ( \17464 , \17226 , \17235 );
or \U$17262 ( \17465 , \17462 , \17463 , \17464 );
xor \U$17263 ( \17466 , \17461 , \17465 );
and \U$17264 ( \17467 , \17241 , \17245 );
and \U$17265 ( \17468 , \17245 , \17250 );
and \U$17266 ( \17469 , \17241 , \17250 );
or \U$17267 ( \17470 , \17467 , \17468 , \17469 );
xor \U$17268 ( \17471 , \17466 , \17470 );
and \U$17269 ( \17472 , \17272 , \17276 );
and \U$17270 ( \17473 , \17276 , \17281 );
and \U$17271 ( \17474 , \17272 , \17281 );
or \U$17272 ( \17475 , \17472 , \17473 , \17474 );
and \U$17273 ( \17476 , \17286 , \17290 );
and \U$17274 ( \17477 , \17290 , \17295 );
and \U$17275 ( \17478 , \17286 , \17295 );
or \U$17276 ( \17479 , \17476 , \17477 , \17478 );
xor \U$17277 ( \17480 , \17475 , \17479 );
and \U$17278 ( \17481 , \17301 , \17305 );
and \U$17279 ( \17482 , \17305 , \17310 );
and \U$17280 ( \17483 , \17301 , \17310 );
or \U$17281 ( \17484 , \17481 , \17482 , \17483 );
xor \U$17282 ( \17485 , \17480 , \17484 );
xor \U$17283 ( \17486 , \17471 , \17485 );
not \U$17284 ( \17487 , \1697 );
and \U$17285 ( \17488 , \10206 , \2121 );
and \U$17286 ( \17489 , \10584 , \2008 );
nor \U$17287 ( \17490 , \17488 , \17489 );
xnor \U$17288 ( \17491 , \17490 , \1961 );
xor \U$17289 ( \17492 , \17487 , \17491 );
and \U$17290 ( \17493 , \9465 , \2400 );
and \U$17291 ( \17494 , \9897 , \2246 );
nor \U$17292 ( \17495 , \17493 , \17494 );
xnor \U$17293 ( \17496 , \17495 , \2195 );
xor \U$17294 ( \17497 , \17492 , \17496 );
and \U$17295 ( \17498 , \4364 , \6401 );
and \U$17296 ( \17499 , \4654 , \6143 );
nor \U$17297 ( \17500 , \17498 , \17499 );
xnor \U$17298 ( \17501 , \17500 , \6148 );
and \U$17299 ( \17502 , \3912 , \7055 );
and \U$17300 ( \17503 , \4160 , \6675 );
nor \U$17301 ( \17504 , \17502 , \17503 );
xnor \U$17302 ( \17505 , \17504 , \6680 );
xor \U$17303 ( \17506 , \17501 , \17505 );
and \U$17304 ( \17507 , \3646 , \7489 );
and \U$17305 ( \17508 , \3736 , \7137 );
nor \U$17306 ( \17509 , \17507 , \17508 );
xnor \U$17307 ( \17510 , \17509 , \7142 );
xor \U$17308 ( \17511 , \17506 , \17510 );
and \U$17309 ( \17512 , \5674 , \5011 );
and \U$17310 ( \17513 , \6030 , \4878 );
nor \U$17311 ( \17514 , \17512 , \17513 );
xnor \U$17312 ( \17515 , \17514 , \4762 );
and \U$17313 ( \17516 , \5156 , \5485 );
and \U$17314 ( \17517 , \5469 , \5275 );
nor \U$17315 ( \17518 , \17516 , \17517 );
xnor \U$17316 ( \17519 , \17518 , \5169 );
xor \U$17317 ( \17520 , \17515 , \17519 );
and \U$17318 ( \17521 , \4749 , \5996 );
and \U$17319 ( \17522 , \4922 , \5695 );
nor \U$17320 ( \17523 , \17521 , \17522 );
xnor \U$17321 ( \17524 , \17523 , \5687 );
xor \U$17322 ( \17525 , \17520 , \17524 );
xor \U$17323 ( \17526 , \17511 , \17525 );
and \U$17324 ( \17527 , \7231 , \3813 );
and \U$17325 ( \17528 , \7556 , \3557 );
nor \U$17326 ( \17529 , \17527 , \17528 );
xnor \U$17327 ( \17530 , \17529 , \3562 );
and \U$17328 ( \17531 , \6790 , \4132 );
and \U$17329 ( \17532 , \6945 , \4012 );
nor \U$17330 ( \17533 , \17531 , \17532 );
xnor \U$17331 ( \17534 , \17533 , \3925 );
xor \U$17332 ( \17535 , \17530 , \17534 );
and \U$17333 ( \17536 , \6281 , \4581 );
and \U$17334 ( \17537 , \6514 , \4424 );
nor \U$17335 ( \17538 , \17536 , \17537 );
xnor \U$17336 ( \17539 , \17538 , \4377 );
xor \U$17337 ( \17540 , \17535 , \17539 );
xor \U$17338 ( \17541 , \17526 , \17540 );
xor \U$17339 ( \17542 , \17497 , \17541 );
and \U$17340 ( \17543 , \17321 , \17325 );
and \U$17341 ( \17544 , \17325 , \17327 );
and \U$17342 ( \17545 , \17321 , \17327 );
or \U$17343 ( \17546 , \17543 , \17544 , \17545 );
and \U$17344 ( \17547 , \2182 , \9765 );
and \U$17345 ( \17548 , \2366 , \9644 );
nor \U$17346 ( \17549 , \17547 , \17548 );
xnor \U$17347 ( \17550 , \17549 , \9478 );
and \U$17348 ( \17551 , \1948 , \10408 );
and \U$17349 ( \17552 , \2090 , \10116 );
nor \U$17350 ( \17553 , \17551 , \17552 );
xnor \U$17351 ( \17554 , \17553 , \10121 );
xor \U$17352 ( \17555 , \17550 , \17554 );
and \U$17353 ( \17556 , \1802 , \10118 );
xor \U$17354 ( \17557 , \17555 , \17556 );
xor \U$17355 ( \17558 , \17546 , \17557 );
and \U$17356 ( \17559 , \3143 , \8019 );
and \U$17357 ( \17560 , \3395 , \7830 );
nor \U$17358 ( \17561 , \17559 , \17560 );
xnor \U$17359 ( \17562 , \17561 , \7713 );
and \U$17360 ( \17563 , \2826 , \8540 );
and \U$17361 ( \17564 , \3037 , \8292 );
nor \U$17362 ( \17565 , \17563 , \17564 );
xnor \U$17363 ( \17566 , \17565 , \8297 );
xor \U$17364 ( \17567 , \17562 , \17566 );
and \U$17365 ( \17568 , \2521 , \9333 );
and \U$17366 ( \17569 , \2757 , \9006 );
nor \U$17367 ( \17570 , \17568 , \17569 );
xnor \U$17368 ( \17571 , \17570 , \8848 );
xor \U$17369 ( \17572 , \17567 , \17571 );
xor \U$17370 ( \17573 , \17558 , \17572 );
xor \U$17371 ( \17574 , \17542 , \17573 );
xor \U$17372 ( \17575 , \17486 , \17574 );
xor \U$17373 ( \17576 , \17457 , \17575 );
xor \U$17374 ( \17577 , \17431 , \17576 );
xor \U$17375 ( \17578 , \17392 , \17577 );
xor \U$17376 ( \17579 , \17386 , \17578 );
and \U$17377 ( \17580 , \17173 , \17373 );
xor \U$17378 ( \17581 , \17579 , \17580 );
and \U$17379 ( \17582 , \17374 , \17375 );
and \U$17380 ( \17583 , \17376 , \17379 );
or \U$17381 ( \17584 , \17582 , \17583 );
xor \U$17382 ( \17585 , \17581 , \17584 );
buf g54e9_GF_PartitionCandidate( \17586_nG54e9 , \17585 );
buf \U$17383 ( \17587 , \17586_nG54e9 );
and \U$17384 ( \17588 , \17390 , \17391 );
and \U$17385 ( \17589 , \17391 , \17577 );
and \U$17386 ( \17590 , \17390 , \17577 );
or \U$17387 ( \17591 , \17588 , \17589 , \17590 );
and \U$17388 ( \17592 , \17396 , \17430 );
and \U$17389 ( \17593 , \17430 , \17576 );
and \U$17390 ( \17594 , \17396 , \17576 );
or \U$17391 ( \17595 , \17592 , \17593 , \17594 );
and \U$17392 ( \17596 , \17400 , \17404 );
and \U$17393 ( \17597 , \17404 , \17429 );
and \U$17394 ( \17598 , \17400 , \17429 );
or \U$17395 ( \17599 , \17596 , \17597 , \17598 );
and \U$17396 ( \17600 , \17442 , \17456 );
and \U$17397 ( \17601 , \17456 , \17575 );
and \U$17398 ( \17602 , \17442 , \17575 );
or \U$17399 ( \17603 , \17600 , \17601 , \17602 );
xor \U$17400 ( \17604 , \17599 , \17603 );
and \U$17401 ( \17605 , \17435 , \17439 );
and \U$17402 ( \17606 , \17439 , \17441 );
and \U$17403 ( \17607 , \17435 , \17441 );
or \U$17404 ( \17608 , \17605 , \17606 , \17607 );
and \U$17405 ( \17609 , \17409 , \17413 );
and \U$17406 ( \17610 , \17413 , \17428 );
and \U$17407 ( \17611 , \17409 , \17428 );
or \U$17408 ( \17612 , \17609 , \17610 , \17611 );
xor \U$17409 ( \17613 , \17608 , \17612 );
and \U$17410 ( \17614 , \17497 , \17541 );
and \U$17411 ( \17615 , \17541 , \17573 );
and \U$17412 ( \17616 , \17497 , \17573 );
or \U$17413 ( \17617 , \17614 , \17615 , \17616 );
xor \U$17414 ( \17618 , \17613 , \17617 );
xor \U$17415 ( \17619 , \17604 , \17618 );
xor \U$17416 ( \17620 , \17595 , \17619 );
and \U$17417 ( \17621 , \17446 , \17450 );
and \U$17418 ( \17622 , \17450 , \17455 );
and \U$17419 ( \17623 , \17446 , \17455 );
or \U$17420 ( \17624 , \17621 , \17622 , \17623 );
and \U$17421 ( \17625 , \17471 , \17485 );
and \U$17422 ( \17626 , \17485 , \17574 );
and \U$17423 ( \17627 , \17471 , \17574 );
or \U$17424 ( \17628 , \17625 , \17626 , \17627 );
xor \U$17425 ( \17629 , \17624 , \17628 );
and \U$17426 ( \17630 , \17461 , \17465 );
and \U$17427 ( \17631 , \17465 , \17470 );
and \U$17428 ( \17632 , \17461 , \17470 );
or \U$17429 ( \17633 , \17630 , \17631 , \17632 );
and \U$17430 ( \17634 , \17475 , \17479 );
and \U$17431 ( \17635 , \17479 , \17484 );
and \U$17432 ( \17636 , \17475 , \17484 );
or \U$17433 ( \17637 , \17634 , \17635 , \17636 );
xor \U$17434 ( \17638 , \17633 , \17637 );
and \U$17435 ( \17639 , \17546 , \17557 );
and \U$17436 ( \17640 , \17557 , \17572 );
and \U$17437 ( \17641 , \17546 , \17572 );
or \U$17438 ( \17642 , \17639 , \17640 , \17641 );
xor \U$17439 ( \17643 , \17638 , \17642 );
and \U$17440 ( \17644 , \17501 , \17505 );
and \U$17441 ( \17645 , \17505 , \17510 );
and \U$17442 ( \17646 , \17501 , \17510 );
or \U$17443 ( \17647 , \17644 , \17645 , \17646 );
and \U$17444 ( \17648 , \17515 , \17519 );
and \U$17445 ( \17649 , \17519 , \17524 );
and \U$17446 ( \17650 , \17515 , \17524 );
or \U$17447 ( \17651 , \17648 , \17649 , \17650 );
xor \U$17448 ( \17652 , \17647 , \17651 );
and \U$17449 ( \17653 , \17562 , \17566 );
and \U$17450 ( \17654 , \17566 , \17571 );
and \U$17451 ( \17655 , \17562 , \17571 );
or \U$17452 ( \17656 , \17653 , \17654 , \17655 );
xor \U$17453 ( \17657 , \17652 , \17656 );
and \U$17454 ( \17658 , \17487 , \17491 );
and \U$17455 ( \17659 , \17491 , \17496 );
and \U$17456 ( \17660 , \17487 , \17496 );
or \U$17457 ( \17661 , \17658 , \17659 , \17660 );
and \U$17458 ( \17662 , \17418 , \17422 );
and \U$17459 ( \17663 , \17422 , \17427 );
and \U$17460 ( \17664 , \17418 , \17427 );
or \U$17461 ( \17665 , \17662 , \17663 , \17664 );
xor \U$17462 ( \17666 , \17661 , \17665 );
and \U$17463 ( \17667 , \17530 , \17534 );
and \U$17464 ( \17668 , \17534 , \17539 );
and \U$17465 ( \17669 , \17530 , \17539 );
or \U$17466 ( \17670 , \17667 , \17668 , \17669 );
xor \U$17467 ( \17671 , \17666 , \17670 );
xor \U$17468 ( \17672 , \17657 , \17671 );
and \U$17469 ( \17673 , \17550 , \17554 );
and \U$17470 ( \17674 , \17554 , \17556 );
and \U$17471 ( \17675 , \17550 , \17556 );
or \U$17472 ( \17676 , \17673 , \17674 , \17675 );
and \U$17473 ( \17677 , \3037 , \8540 );
and \U$17474 ( \17678 , \3143 , \8292 );
nor \U$17475 ( \17679 , \17677 , \17678 );
xnor \U$17476 ( \17680 , \17679 , \8297 );
and \U$17477 ( \17681 , \2757 , \9333 );
and \U$17478 ( \17682 , \2826 , \9006 );
nor \U$17479 ( \17683 , \17681 , \17682 );
xnor \U$17480 ( \17684 , \17683 , \8848 );
xor \U$17481 ( \17685 , \17680 , \17684 );
and \U$17482 ( \17686 , \2366 , \9765 );
and \U$17483 ( \17687 , \2521 , \9644 );
nor \U$17484 ( \17688 , \17686 , \17687 );
xnor \U$17485 ( \17689 , \17688 , \9478 );
xor \U$17486 ( \17690 , \17685 , \17689 );
xor \U$17487 ( \17691 , \17676 , \17690 );
and \U$17488 ( \17692 , \2090 , \10408 );
and \U$17489 ( \17693 , \2182 , \10116 );
nor \U$17490 ( \17694 , \17692 , \17693 );
xnor \U$17491 ( \17695 , \17694 , \10121 );
and \U$17492 ( \17696 , \1948 , \10118 );
xnor \U$17493 ( \17697 , \17695 , \17696 );
xor \U$17494 ( \17698 , \17691 , \17697 );
xor \U$17495 ( \17699 , \17672 , \17698 );
xor \U$17496 ( \17700 , \17643 , \17699 );
and \U$17497 ( \17701 , \17511 , \17525 );
and \U$17498 ( \17702 , \17525 , \17540 );
and \U$17499 ( \17703 , \17511 , \17540 );
or \U$17500 ( \17704 , \17701 , \17702 , \17703 );
and \U$17501 ( \17705 , \5469 , \5485 );
and \U$17502 ( \17706 , \5674 , \5275 );
nor \U$17503 ( \17707 , \17705 , \17706 );
xnor \U$17504 ( \17708 , \17707 , \5169 );
and \U$17505 ( \17709 , \4922 , \5996 );
and \U$17506 ( \17710 , \5156 , \5695 );
nor \U$17507 ( \17711 , \17709 , \17710 );
xnor \U$17508 ( \17712 , \17711 , \5687 );
xor \U$17509 ( \17713 , \17708 , \17712 );
and \U$17510 ( \17714 , \4654 , \6401 );
and \U$17511 ( \17715 , \4749 , \6143 );
nor \U$17512 ( \17716 , \17714 , \17715 );
xnor \U$17513 ( \17717 , \17716 , \6148 );
xor \U$17514 ( \17718 , \17713 , \17717 );
and \U$17515 ( \17719 , \4160 , \7055 );
and \U$17516 ( \17720 , \4364 , \6675 );
nor \U$17517 ( \17721 , \17719 , \17720 );
xnor \U$17518 ( \17722 , \17721 , \6680 );
and \U$17519 ( \17723 , \3736 , \7489 );
and \U$17520 ( \17724 , \3912 , \7137 );
nor \U$17521 ( \17725 , \17723 , \17724 );
xnor \U$17522 ( \17726 , \17725 , \7142 );
xor \U$17523 ( \17727 , \17722 , \17726 );
and \U$17524 ( \17728 , \3395 , \8019 );
and \U$17525 ( \17729 , \3646 , \7830 );
nor \U$17526 ( \17730 , \17728 , \17729 );
xnor \U$17527 ( \17731 , \17730 , \7713 );
xor \U$17528 ( \17732 , \17727 , \17731 );
xor \U$17529 ( \17733 , \17718 , \17732 );
and \U$17530 ( \17734 , \6945 , \4132 );
and \U$17531 ( \17735 , \7231 , \4012 );
nor \U$17532 ( \17736 , \17734 , \17735 );
xnor \U$17533 ( \17737 , \17736 , \3925 );
and \U$17534 ( \17738 , \6514 , \4581 );
and \U$17535 ( \17739 , \6790 , \4424 );
nor \U$17536 ( \17740 , \17738 , \17739 );
xnor \U$17537 ( \17741 , \17740 , \4377 );
xor \U$17538 ( \17742 , \17737 , \17741 );
and \U$17539 ( \17743 , \6030 , \5011 );
and \U$17540 ( \17744 , \6281 , \4878 );
nor \U$17541 ( \17745 , \17743 , \17744 );
xnor \U$17542 ( \17746 , \17745 , \4762 );
xor \U$17543 ( \17747 , \17742 , \17746 );
xor \U$17544 ( \17748 , \17733 , \17747 );
xor \U$17545 ( \17749 , \17704 , \17748 );
and \U$17546 ( \17750 , \10584 , \2121 );
not \U$17547 ( \17751 , \17750 );
xnor \U$17548 ( \17752 , \17751 , \1961 );
and \U$17549 ( \17753 , \9897 , \2400 );
and \U$17550 ( \17754 , \10206 , \2246 );
nor \U$17551 ( \17755 , \17753 , \17754 );
xnor \U$17552 ( \17756 , \17755 , \2195 );
xor \U$17553 ( \17757 , \17752 , \17756 );
and \U$17554 ( \17758 , \9169 , \2669 );
and \U$17555 ( \17759 , \9465 , \2538 );
nor \U$17556 ( \17760 , \17758 , \17759 );
xnor \U$17557 ( \17761 , \17760 , \2534 );
xor \U$17558 ( \17762 , \17757 , \17761 );
and \U$17559 ( \17763 , \8652 , \3103 );
and \U$17560 ( \17764 , \8835 , \2934 );
nor \U$17561 ( \17765 , \17763 , \17764 );
xnor \U$17562 ( \17766 , \17765 , \2839 );
and \U$17563 ( \17767 , \8057 , \3357 );
and \U$17564 ( \17768 , \8349 , \3255 );
nor \U$17565 ( \17769 , \17767 , \17768 );
xnor \U$17566 ( \17770 , \17769 , \3156 );
xor \U$17567 ( \17771 , \17766 , \17770 );
and \U$17568 ( \17772 , \7556 , \3813 );
and \U$17569 ( \17773 , \7700 , \3557 );
nor \U$17570 ( \17774 , \17772 , \17773 );
xnor \U$17571 ( \17775 , \17774 , \3562 );
xor \U$17572 ( \17776 , \17771 , \17775 );
xor \U$17573 ( \17777 , \17762 , \17776 );
xor \U$17574 ( \17778 , \17749 , \17777 );
xor \U$17575 ( \17779 , \17700 , \17778 );
xor \U$17576 ( \17780 , \17629 , \17779 );
xor \U$17577 ( \17781 , \17620 , \17780 );
xor \U$17578 ( \17782 , \17591 , \17781 );
and \U$17579 ( \17783 , \17386 , \17578 );
xor \U$17580 ( \17784 , \17782 , \17783 );
and \U$17581 ( \17785 , \17579 , \17580 );
and \U$17582 ( \17786 , \17581 , \17584 );
or \U$17583 ( \17787 , \17785 , \17786 );
xor \U$17584 ( \17788 , \17784 , \17787 );
buf g54e7_GF_PartitionCandidate( \17789_nG54e7 , \17788 );
buf \U$17585 ( \17790 , \17789_nG54e7 );
and \U$17586 ( \17791 , \17599 , \17603 );
and \U$17587 ( \17792 , \17603 , \17618 );
and \U$17588 ( \17793 , \17599 , \17618 );
or \U$17589 ( \17794 , \17791 , \17792 , \17793 );
and \U$17590 ( \17795 , \17595 , \17619 );
and \U$17591 ( \17796 , \17619 , \17780 );
and \U$17592 ( \17797 , \17595 , \17780 );
or \U$17593 ( \17798 , \17795 , \17796 , \17797 );
xor \U$17594 ( \17799 , \17794 , \17798 );
and \U$17595 ( \17800 , \17624 , \17628 );
and \U$17596 ( \17801 , \17628 , \17779 );
and \U$17597 ( \17802 , \17624 , \17779 );
or \U$17598 ( \17803 , \17800 , \17801 , \17802 );
and \U$17599 ( \17804 , \17608 , \17612 );
and \U$17600 ( \17805 , \17612 , \17617 );
and \U$17601 ( \17806 , \17608 , \17617 );
or \U$17602 ( \17807 , \17804 , \17805 , \17806 );
and \U$17603 ( \17808 , \17643 , \17699 );
and \U$17604 ( \17809 , \17699 , \17778 );
and \U$17605 ( \17810 , \17643 , \17778 );
or \U$17606 ( \17811 , \17808 , \17809 , \17810 );
xor \U$17607 ( \17812 , \17807 , \17811 );
and \U$17608 ( \17813 , \17647 , \17651 );
and \U$17609 ( \17814 , \17651 , \17656 );
and \U$17610 ( \17815 , \17647 , \17656 );
or \U$17611 ( \17816 , \17813 , \17814 , \17815 );
and \U$17612 ( \17817 , \17661 , \17665 );
and \U$17613 ( \17818 , \17665 , \17670 );
and \U$17614 ( \17819 , \17661 , \17670 );
or \U$17615 ( \17820 , \17817 , \17818 , \17819 );
xor \U$17616 ( \17821 , \17816 , \17820 );
and \U$17617 ( \17822 , \17676 , \17690 );
and \U$17618 ( \17823 , \17690 , \17697 );
and \U$17619 ( \17824 , \17676 , \17697 );
or \U$17620 ( \17825 , \17822 , \17823 , \17824 );
xor \U$17621 ( \17826 , \17821 , \17825 );
xor \U$17622 ( \17827 , \17812 , \17826 );
xor \U$17623 ( \17828 , \17803 , \17827 );
and \U$17624 ( \17829 , \17633 , \17637 );
and \U$17625 ( \17830 , \17637 , \17642 );
and \U$17626 ( \17831 , \17633 , \17642 );
or \U$17627 ( \17832 , \17829 , \17830 , \17831 );
and \U$17628 ( \17833 , \17657 , \17671 );
and \U$17629 ( \17834 , \17671 , \17698 );
and \U$17630 ( \17835 , \17657 , \17698 );
or \U$17631 ( \17836 , \17833 , \17834 , \17835 );
xor \U$17632 ( \17837 , \17832 , \17836 );
and \U$17633 ( \17838 , \17704 , \17748 );
and \U$17634 ( \17839 , \17748 , \17777 );
and \U$17635 ( \17840 , \17704 , \17777 );
or \U$17636 ( \17841 , \17838 , \17839 , \17840 );
xor \U$17637 ( \17842 , \17837 , \17841 );
and \U$17638 ( \17843 , \17752 , \17756 );
and \U$17639 ( \17844 , \17756 , \17761 );
and \U$17640 ( \17845 , \17752 , \17761 );
or \U$17641 ( \17846 , \17843 , \17844 , \17845 );
and \U$17642 ( \17847 , \17766 , \17770 );
and \U$17643 ( \17848 , \17770 , \17775 );
and \U$17644 ( \17849 , \17766 , \17775 );
or \U$17645 ( \17850 , \17847 , \17848 , \17849 );
xor \U$17646 ( \17851 , \17846 , \17850 );
and \U$17647 ( \17852 , \17737 , \17741 );
and \U$17648 ( \17853 , \17741 , \17746 );
and \U$17649 ( \17854 , \17737 , \17746 );
or \U$17650 ( \17855 , \17852 , \17853 , \17854 );
xor \U$17651 ( \17856 , \17851 , \17855 );
and \U$17652 ( \17857 , \17718 , \17732 );
and \U$17653 ( \17858 , \17732 , \17747 );
and \U$17654 ( \17859 , \17718 , \17747 );
or \U$17655 ( \17860 , \17857 , \17858 , \17859 );
and \U$17656 ( \17861 , \17762 , \17776 );
xor \U$17657 ( \17862 , \17860 , \17861 );
not \U$17658 ( \17863 , \1961 );
and \U$17659 ( \17864 , \10206 , \2400 );
and \U$17660 ( \17865 , \10584 , \2246 );
nor \U$17661 ( \17866 , \17864 , \17865 );
xnor \U$17662 ( \17867 , \17866 , \2195 );
xor \U$17663 ( \17868 , \17863 , \17867 );
and \U$17664 ( \17869 , \9465 , \2669 );
and \U$17665 ( \17870 , \9897 , \2538 );
nor \U$17666 ( \17871 , \17869 , \17870 );
xnor \U$17667 ( \17872 , \17871 , \2534 );
xor \U$17668 ( \17873 , \17868 , \17872 );
and \U$17669 ( \17874 , \8835 , \3103 );
and \U$17670 ( \17875 , \9169 , \2934 );
nor \U$17671 ( \17876 , \17874 , \17875 );
xnor \U$17672 ( \17877 , \17876 , \2839 );
and \U$17673 ( \17878 , \8349 , \3357 );
and \U$17674 ( \17879 , \8652 , \3255 );
nor \U$17675 ( \17880 , \17878 , \17879 );
xnor \U$17676 ( \17881 , \17880 , \3156 );
xor \U$17677 ( \17882 , \17877 , \17881 );
and \U$17678 ( \17883 , \7700 , \3813 );
and \U$17679 ( \17884 , \8057 , \3557 );
nor \U$17680 ( \17885 , \17883 , \17884 );
xnor \U$17681 ( \17886 , \17885 , \3562 );
xor \U$17682 ( \17887 , \17882 , \17886 );
xor \U$17683 ( \17888 , \17873 , \17887 );
and \U$17684 ( \17889 , \7231 , \4132 );
and \U$17685 ( \17890 , \7556 , \4012 );
nor \U$17686 ( \17891 , \17889 , \17890 );
xnor \U$17687 ( \17892 , \17891 , \3925 );
and \U$17688 ( \17893 , \6790 , \4581 );
and \U$17689 ( \17894 , \6945 , \4424 );
nor \U$17690 ( \17895 , \17893 , \17894 );
xnor \U$17691 ( \17896 , \17895 , \4377 );
xor \U$17692 ( \17897 , \17892 , \17896 );
and \U$17693 ( \17898 , \6281 , \5011 );
and \U$17694 ( \17899 , \6514 , \4878 );
nor \U$17695 ( \17900 , \17898 , \17899 );
xnor \U$17696 ( \17901 , \17900 , \4762 );
xor \U$17697 ( \17902 , \17897 , \17901 );
xor \U$17698 ( \17903 , \17888 , \17902 );
xor \U$17699 ( \17904 , \17862 , \17903 );
xor \U$17700 ( \17905 , \17856 , \17904 );
and \U$17701 ( \17906 , \17708 , \17712 );
and \U$17702 ( \17907 , \17712 , \17717 );
and \U$17703 ( \17908 , \17708 , \17717 );
or \U$17704 ( \17909 , \17906 , \17907 , \17908 );
and \U$17705 ( \17910 , \17722 , \17726 );
and \U$17706 ( \17911 , \17726 , \17731 );
and \U$17707 ( \17912 , \17722 , \17731 );
or \U$17708 ( \17913 , \17910 , \17911 , \17912 );
xor \U$17709 ( \17914 , \17909 , \17913 );
and \U$17710 ( \17915 , \17680 , \17684 );
and \U$17711 ( \17916 , \17684 , \17689 );
and \U$17712 ( \17917 , \17680 , \17689 );
or \U$17713 ( \17918 , \17915 , \17916 , \17917 );
xor \U$17714 ( \17919 , \17914 , \17918 );
or \U$17715 ( \17920 , \17695 , \17696 );
and \U$17716 ( \17921 , \2182 , \10408 );
and \U$17717 ( \17922 , \2366 , \10116 );
nor \U$17718 ( \17923 , \17921 , \17922 );
xnor \U$17719 ( \17924 , \17923 , \10121 );
xor \U$17720 ( \17925 , \17920 , \17924 );
and \U$17721 ( \17926 , \2090 , \10118 );
xor \U$17722 ( \17927 , \17925 , \17926 );
xor \U$17723 ( \17928 , \17919 , \17927 );
and \U$17724 ( \17929 , \4364 , \7055 );
and \U$17725 ( \17930 , \4654 , \6675 );
nor \U$17726 ( \17931 , \17929 , \17930 );
xnor \U$17727 ( \17932 , \17931 , \6680 );
and \U$17728 ( \17933 , \3912 , \7489 );
and \U$17729 ( \17934 , \4160 , \7137 );
nor \U$17730 ( \17935 , \17933 , \17934 );
xnor \U$17731 ( \17936 , \17935 , \7142 );
xor \U$17732 ( \17937 , \17932 , \17936 );
and \U$17733 ( \17938 , \3646 , \8019 );
and \U$17734 ( \17939 , \3736 , \7830 );
nor \U$17735 ( \17940 , \17938 , \17939 );
xnor \U$17736 ( \17941 , \17940 , \7713 );
xor \U$17737 ( \17942 , \17937 , \17941 );
and \U$17738 ( \17943 , \5674 , \5485 );
and \U$17739 ( \17944 , \6030 , \5275 );
nor \U$17740 ( \17945 , \17943 , \17944 );
xnor \U$17741 ( \17946 , \17945 , \5169 );
and \U$17742 ( \17947 , \5156 , \5996 );
and \U$17743 ( \17948 , \5469 , \5695 );
nor \U$17744 ( \17949 , \17947 , \17948 );
xnor \U$17745 ( \17950 , \17949 , \5687 );
xor \U$17746 ( \17951 , \17946 , \17950 );
and \U$17747 ( \17952 , \4749 , \6401 );
and \U$17748 ( \17953 , \4922 , \6143 );
nor \U$17749 ( \17954 , \17952 , \17953 );
xnor \U$17750 ( \17955 , \17954 , \6148 );
xor \U$17751 ( \17956 , \17951 , \17955 );
xor \U$17752 ( \17957 , \17942 , \17956 );
and \U$17753 ( \17958 , \3143 , \8540 );
and \U$17754 ( \17959 , \3395 , \8292 );
nor \U$17755 ( \17960 , \17958 , \17959 );
xnor \U$17756 ( \17961 , \17960 , \8297 );
and \U$17757 ( \17962 , \2826 , \9333 );
and \U$17758 ( \17963 , \3037 , \9006 );
nor \U$17759 ( \17964 , \17962 , \17963 );
xnor \U$17760 ( \17965 , \17964 , \8848 );
xor \U$17761 ( \17966 , \17961 , \17965 );
and \U$17762 ( \17967 , \2521 , \9765 );
and \U$17763 ( \17968 , \2757 , \9644 );
nor \U$17764 ( \17969 , \17967 , \17968 );
xnor \U$17765 ( \17970 , \17969 , \9478 );
xor \U$17766 ( \17971 , \17966 , \17970 );
xor \U$17767 ( \17972 , \17957 , \17971 );
xor \U$17768 ( \17973 , \17928 , \17972 );
xor \U$17769 ( \17974 , \17905 , \17973 );
xor \U$17770 ( \17975 , \17842 , \17974 );
xor \U$17771 ( \17976 , \17828 , \17975 );
xor \U$17772 ( \17977 , \17799 , \17976 );
and \U$17773 ( \17978 , \17591 , \17781 );
xor \U$17774 ( \17979 , \17977 , \17978 );
and \U$17775 ( \17980 , \17782 , \17783 );
and \U$17776 ( \17981 , \17784 , \17787 );
or \U$17777 ( \17982 , \17980 , \17981 );
xor \U$17778 ( \17983 , \17979 , \17982 );
buf g54e5_GF_PartitionCandidate( \17984_nG54e5 , \17983 );
buf \U$17779 ( \17985 , \17984_nG54e5 );
and \U$17780 ( \17986 , \17803 , \17827 );
and \U$17781 ( \17987 , \17827 , \17975 );
and \U$17782 ( \17988 , \17803 , \17975 );
or \U$17783 ( \17989 , \17986 , \17987 , \17988 );
and \U$17784 ( \17990 , \17832 , \17836 );
and \U$17785 ( \17991 , \17836 , \17841 );
and \U$17786 ( \17992 , \17832 , \17841 );
or \U$17787 ( \17993 , \17990 , \17991 , \17992 );
and \U$17788 ( \17994 , \17856 , \17904 );
and \U$17789 ( \17995 , \17904 , \17973 );
and \U$17790 ( \17996 , \17856 , \17973 );
or \U$17791 ( \17997 , \17994 , \17995 , \17996 );
xor \U$17792 ( \17998 , \17993 , \17997 );
and \U$17793 ( \17999 , \17942 , \17956 );
and \U$17794 ( \18000 , \17956 , \17971 );
and \U$17795 ( \18001 , \17942 , \17971 );
or \U$17796 ( \18002 , \17999 , \18000 , \18001 );
and \U$17797 ( \18003 , \17873 , \17887 );
and \U$17798 ( \18004 , \17887 , \17902 );
and \U$17799 ( \18005 , \17873 , \17902 );
or \U$17800 ( \18006 , \18003 , \18004 , \18005 );
xor \U$17801 ( \18007 , \18002 , \18006 );
and \U$17802 ( \18008 , \8652 , \3357 );
and \U$17803 ( \18009 , \8835 , \3255 );
nor \U$17804 ( \18010 , \18008 , \18009 );
xnor \U$17805 ( \18011 , \18010 , \3156 );
and \U$17806 ( \18012 , \8057 , \3813 );
and \U$17807 ( \18013 , \8349 , \3557 );
nor \U$17808 ( \18014 , \18012 , \18013 );
xnor \U$17809 ( \18015 , \18014 , \3562 );
xor \U$17810 ( \18016 , \18011 , \18015 );
and \U$17811 ( \18017 , \7556 , \4132 );
and \U$17812 ( \18018 , \7700 , \4012 );
nor \U$17813 ( \18019 , \18017 , \18018 );
xnor \U$17814 ( \18020 , \18019 , \3925 );
xor \U$17815 ( \18021 , \18016 , \18020 );
xor \U$17816 ( \18022 , \18007 , \18021 );
xor \U$17817 ( \18023 , \17998 , \18022 );
xor \U$17818 ( \18024 , \17989 , \18023 );
and \U$17819 ( \18025 , \17807 , \17811 );
and \U$17820 ( \18026 , \17811 , \17826 );
and \U$17821 ( \18027 , \17807 , \17826 );
or \U$17822 ( \18028 , \18025 , \18026 , \18027 );
and \U$17823 ( \18029 , \17842 , \17974 );
xor \U$17824 ( \18030 , \18028 , \18029 );
and \U$17825 ( \18031 , \17909 , \17913 );
and \U$17826 ( \18032 , \17913 , \17918 );
and \U$17827 ( \18033 , \17909 , \17918 );
or \U$17828 ( \18034 , \18031 , \18032 , \18033 );
and \U$17829 ( \18035 , \17920 , \17924 );
and \U$17830 ( \18036 , \17924 , \17926 );
and \U$17831 ( \18037 , \17920 , \17926 );
or \U$17832 ( \18038 , \18035 , \18036 , \18037 );
xor \U$17833 ( \18039 , \18034 , \18038 );
and \U$17834 ( \18040 , \17846 , \17850 );
and \U$17835 ( \18041 , \17850 , \17855 );
and \U$17836 ( \18042 , \17846 , \17855 );
or \U$17837 ( \18043 , \18040 , \18041 , \18042 );
xor \U$17838 ( \18044 , \18039 , \18043 );
and \U$17839 ( \18045 , \17816 , \17820 );
and \U$17840 ( \18046 , \17820 , \17825 );
and \U$17841 ( \18047 , \17816 , \17825 );
or \U$17842 ( \18048 , \18045 , \18046 , \18047 );
and \U$17843 ( \18049 , \17860 , \17861 );
and \U$17844 ( \18050 , \17861 , \17903 );
and \U$17845 ( \18051 , \17860 , \17903 );
or \U$17846 ( \18052 , \18049 , \18050 , \18051 );
xor \U$17847 ( \18053 , \18048 , \18052 );
and \U$17848 ( \18054 , \17919 , \17927 );
and \U$17849 ( \18055 , \17927 , \17972 );
and \U$17850 ( \18056 , \17919 , \17972 );
or \U$17851 ( \18057 , \18054 , \18055 , \18056 );
xor \U$17852 ( \18058 , \18053 , \18057 );
xor \U$17853 ( \18059 , \18044 , \18058 );
and \U$17854 ( \18060 , \17863 , \17867 );
and \U$17855 ( \18061 , \17867 , \17872 );
and \U$17856 ( \18062 , \17863 , \17872 );
or \U$17857 ( \18063 , \18060 , \18061 , \18062 );
and \U$17858 ( \18064 , \17877 , \17881 );
and \U$17859 ( \18065 , \17881 , \17886 );
and \U$17860 ( \18066 , \17877 , \17886 );
or \U$17861 ( \18067 , \18064 , \18065 , \18066 );
xor \U$17862 ( \18068 , \18063 , \18067 );
and \U$17863 ( \18069 , \17892 , \17896 );
and \U$17864 ( \18070 , \17896 , \17901 );
and \U$17865 ( \18071 , \17892 , \17901 );
or \U$17866 ( \18072 , \18069 , \18070 , \18071 );
xor \U$17867 ( \18073 , \18068 , \18072 );
and \U$17868 ( \18074 , \17932 , \17936 );
and \U$17869 ( \18075 , \17936 , \17941 );
and \U$17870 ( \18076 , \17932 , \17941 );
or \U$17871 ( \18077 , \18074 , \18075 , \18076 );
and \U$17872 ( \18078 , \17946 , \17950 );
and \U$17873 ( \18079 , \17950 , \17955 );
and \U$17874 ( \18080 , \17946 , \17955 );
or \U$17875 ( \18081 , \18078 , \18079 , \18080 );
xor \U$17876 ( \18082 , \18077 , \18081 );
and \U$17877 ( \18083 , \17961 , \17965 );
and \U$17878 ( \18084 , \17965 , \17970 );
and \U$17879 ( \18085 , \17961 , \17970 );
or \U$17880 ( \18086 , \18083 , \18084 , \18085 );
xor \U$17881 ( \18087 , \18082 , \18086 );
xor \U$17882 ( \18088 , \18073 , \18087 );
and \U$17883 ( \18089 , \10584 , \2400 );
not \U$17884 ( \18090 , \18089 );
xnor \U$17885 ( \18091 , \18090 , \2195 );
and \U$17886 ( \18092 , \9897 , \2669 );
and \U$17887 ( \18093 , \10206 , \2538 );
nor \U$17888 ( \18094 , \18092 , \18093 );
xnor \U$17889 ( \18095 , \18094 , \2534 );
xor \U$17890 ( \18096 , \18091 , \18095 );
and \U$17891 ( \18097 , \9169 , \3103 );
and \U$17892 ( \18098 , \9465 , \2934 );
nor \U$17893 ( \18099 , \18097 , \18098 );
xnor \U$17894 ( \18100 , \18099 , \2839 );
xor \U$17895 ( \18101 , \18096 , \18100 );
and \U$17896 ( \18102 , \6945 , \4581 );
and \U$17897 ( \18103 , \7231 , \4424 );
nor \U$17898 ( \18104 , \18102 , \18103 );
xnor \U$17899 ( \18105 , \18104 , \4377 );
and \U$17900 ( \18106 , \6514 , \5011 );
and \U$17901 ( \18107 , \6790 , \4878 );
nor \U$17902 ( \18108 , \18106 , \18107 );
xnor \U$17903 ( \18109 , \18108 , \4762 );
xor \U$17904 ( \18110 , \18105 , \18109 );
and \U$17905 ( \18111 , \6030 , \5485 );
and \U$17906 ( \18112 , \6281 , \5275 );
nor \U$17907 ( \18113 , \18111 , \18112 );
xnor \U$17908 ( \18114 , \18113 , \5169 );
xor \U$17909 ( \18115 , \18110 , \18114 );
and \U$17910 ( \18116 , \5469 , \5996 );
and \U$17911 ( \18117 , \5674 , \5695 );
nor \U$17912 ( \18118 , \18116 , \18117 );
xnor \U$17913 ( \18119 , \18118 , \5687 );
and \U$17914 ( \18120 , \4922 , \6401 );
and \U$17915 ( \18121 , \5156 , \6143 );
nor \U$17916 ( \18122 , \18120 , \18121 );
xnor \U$17917 ( \18123 , \18122 , \6148 );
xor \U$17918 ( \18124 , \18119 , \18123 );
and \U$17919 ( \18125 , \4654 , \7055 );
and \U$17920 ( \18126 , \4749 , \6675 );
nor \U$17921 ( \18127 , \18125 , \18126 );
xnor \U$17922 ( \18128 , \18127 , \6680 );
xor \U$17923 ( \18129 , \18124 , \18128 );
xor \U$17924 ( \18130 , \18115 , \18129 );
and \U$17925 ( \18131 , \4160 , \7489 );
and \U$17926 ( \18132 , \4364 , \7137 );
nor \U$17927 ( \18133 , \18131 , \18132 );
xnor \U$17928 ( \18134 , \18133 , \7142 );
and \U$17929 ( \18135 , \3736 , \8019 );
and \U$17930 ( \18136 , \3912 , \7830 );
nor \U$17931 ( \18137 , \18135 , \18136 );
xnor \U$17932 ( \18138 , \18137 , \7713 );
xor \U$17933 ( \18139 , \18134 , \18138 );
and \U$17934 ( \18140 , \3395 , \8540 );
and \U$17935 ( \18141 , \3646 , \8292 );
nor \U$17936 ( \18142 , \18140 , \18141 );
xnor \U$17937 ( \18143 , \18142 , \8297 );
xor \U$17938 ( \18144 , \18139 , \18143 );
xor \U$17939 ( \18145 , \18130 , \18144 );
xor \U$17940 ( \18146 , \18101 , \18145 );
and \U$17941 ( \18147 , \2182 , \10118 );
and \U$17942 ( \18148 , \3037 , \9333 );
and \U$17943 ( \18149 , \3143 , \9006 );
nor \U$17944 ( \18150 , \18148 , \18149 );
xnor \U$17945 ( \18151 , \18150 , \8848 );
and \U$17946 ( \18152 , \2757 , \9765 );
and \U$17947 ( \18153 , \2826 , \9644 );
nor \U$17948 ( \18154 , \18152 , \18153 );
xnor \U$17949 ( \18155 , \18154 , \9478 );
xor \U$17950 ( \18156 , \18151 , \18155 );
and \U$17951 ( \18157 , \2366 , \10408 );
and \U$17952 ( \18158 , \2521 , \10116 );
nor \U$17953 ( \18159 , \18157 , \18158 );
xnor \U$17954 ( \18160 , \18159 , \10121 );
xor \U$17955 ( \18161 , \18156 , \18160 );
xnor \U$17956 ( \18162 , \18147 , \18161 );
xor \U$17957 ( \18163 , \18146 , \18162 );
xor \U$17958 ( \18164 , \18088 , \18163 );
xor \U$17959 ( \18165 , \18059 , \18164 );
xor \U$17960 ( \18166 , \18030 , \18165 );
xor \U$17961 ( \18167 , \18024 , \18166 );
and \U$17962 ( \18168 , \17794 , \17798 );
and \U$17963 ( \18169 , \17798 , \17976 );
and \U$17964 ( \18170 , \17794 , \17976 );
or \U$17965 ( \18171 , \18168 , \18169 , \18170 );
xor \U$17966 ( \18172 , \18167 , \18171 );
and \U$17967 ( \18173 , \17977 , \17978 );
and \U$17968 ( \18174 , \17979 , \17982 );
or \U$17969 ( \18175 , \18173 , \18174 );
xor \U$17970 ( \18176 , \18172 , \18175 );
buf g54e3_GF_PartitionCandidate( \18177_nG54e3 , \18176 );
buf \U$17971 ( \18178 , \18177_nG54e3 );
and \U$17972 ( \18179 , \18028 , \18029 );
and \U$17973 ( \18180 , \18029 , \18165 );
and \U$17974 ( \18181 , \18028 , \18165 );
or \U$17975 ( \18182 , \18179 , \18180 , \18181 );
and \U$17976 ( \18183 , \17993 , \17997 );
and \U$17977 ( \18184 , \17997 , \18022 );
and \U$17978 ( \18185 , \17993 , \18022 );
or \U$17979 ( \18186 , \18183 , \18184 , \18185 );
and \U$17980 ( \18187 , \18044 , \18058 );
and \U$17981 ( \18188 , \18058 , \18164 );
and \U$17982 ( \18189 , \18044 , \18164 );
or \U$17983 ( \18190 , \18187 , \18188 , \18189 );
xor \U$17984 ( \18191 , \18186 , \18190 );
and \U$17985 ( \18192 , \18034 , \18038 );
and \U$17986 ( \18193 , \18038 , \18043 );
and \U$17987 ( \18194 , \18034 , \18043 );
or \U$17988 ( \18195 , \18192 , \18193 , \18194 );
and \U$17989 ( \18196 , \18002 , \18006 );
and \U$17990 ( \18197 , \18006 , \18021 );
and \U$17991 ( \18198 , \18002 , \18021 );
or \U$17992 ( \18199 , \18196 , \18197 , \18198 );
xor \U$17993 ( \18200 , \18195 , \18199 );
and \U$17994 ( \18201 , \18101 , \18145 );
and \U$17995 ( \18202 , \18145 , \18162 );
and \U$17996 ( \18203 , \18101 , \18162 );
or \U$17997 ( \18204 , \18201 , \18202 , \18203 );
xor \U$17998 ( \18205 , \18200 , \18204 );
xor \U$17999 ( \18206 , \18191 , \18205 );
xor \U$18000 ( \18207 , \18182 , \18206 );
and \U$18001 ( \18208 , \18048 , \18052 );
and \U$18002 ( \18209 , \18052 , \18057 );
and \U$18003 ( \18210 , \18048 , \18057 );
or \U$18004 ( \18211 , \18208 , \18209 , \18210 );
and \U$18005 ( \18212 , \18073 , \18087 );
and \U$18006 ( \18213 , \18087 , \18163 );
and \U$18007 ( \18214 , \18073 , \18163 );
or \U$18008 ( \18215 , \18212 , \18213 , \18214 );
xor \U$18009 ( \18216 , \18211 , \18215 );
and \U$18010 ( \18217 , \18063 , \18067 );
and \U$18011 ( \18218 , \18067 , \18072 );
and \U$18012 ( \18219 , \18063 , \18072 );
or \U$18013 ( \18220 , \18217 , \18218 , \18219 );
and \U$18014 ( \18221 , \18077 , \18081 );
and \U$18015 ( \18222 , \18081 , \18086 );
and \U$18016 ( \18223 , \18077 , \18086 );
or \U$18017 ( \18224 , \18221 , \18222 , \18223 );
xor \U$18018 ( \18225 , \18220 , \18224 );
or \U$18019 ( \18226 , \18147 , \18161 );
xor \U$18020 ( \18227 , \18225 , \18226 );
and \U$18021 ( \18228 , \18115 , \18129 );
and \U$18022 ( \18229 , \18129 , \18144 );
and \U$18023 ( \18230 , \18115 , \18144 );
or \U$18024 ( \18231 , \18228 , \18229 , \18230 );
not \U$18025 ( \18232 , \2195 );
and \U$18026 ( \18233 , \10206 , \2669 );
and \U$18027 ( \18234 , \10584 , \2538 );
nor \U$18028 ( \18235 , \18233 , \18234 );
xnor \U$18029 ( \18236 , \18235 , \2534 );
xor \U$18030 ( \18237 , \18232 , \18236 );
and \U$18031 ( \18238 , \9465 , \3103 );
and \U$18032 ( \18239 , \9897 , \2934 );
nor \U$18033 ( \18240 , \18238 , \18239 );
xnor \U$18034 ( \18241 , \18240 , \2839 );
xor \U$18035 ( \18242 , \18237 , \18241 );
xor \U$18036 ( \18243 , \18231 , \18242 );
and \U$18037 ( \18244 , \7231 , \4581 );
and \U$18038 ( \18245 , \7556 , \4424 );
nor \U$18039 ( \18246 , \18244 , \18245 );
xnor \U$18040 ( \18247 , \18246 , \4377 );
and \U$18041 ( \18248 , \6790 , \5011 );
and \U$18042 ( \18249 , \6945 , \4878 );
nor \U$18043 ( \18250 , \18248 , \18249 );
xnor \U$18044 ( \18251 , \18250 , \4762 );
xor \U$18045 ( \18252 , \18247 , \18251 );
and \U$18046 ( \18253 , \6281 , \5485 );
and \U$18047 ( \18254 , \6514 , \5275 );
nor \U$18048 ( \18255 , \18253 , \18254 );
xnor \U$18049 ( \18256 , \18255 , \5169 );
xor \U$18050 ( \18257 , \18252 , \18256 );
and \U$18051 ( \18258 , \5674 , \5996 );
and \U$18052 ( \18259 , \6030 , \5695 );
nor \U$18053 ( \18260 , \18258 , \18259 );
xnor \U$18054 ( \18261 , \18260 , \5687 );
and \U$18055 ( \18262 , \5156 , \6401 );
and \U$18056 ( \18263 , \5469 , \6143 );
nor \U$18057 ( \18264 , \18262 , \18263 );
xnor \U$18058 ( \18265 , \18264 , \6148 );
xor \U$18059 ( \18266 , \18261 , \18265 );
and \U$18060 ( \18267 , \4749 , \7055 );
and \U$18061 ( \18268 , \4922 , \6675 );
nor \U$18062 ( \18269 , \18267 , \18268 );
xnor \U$18063 ( \18270 , \18269 , \6680 );
xor \U$18064 ( \18271 , \18266 , \18270 );
xor \U$18065 ( \18272 , \18257 , \18271 );
and \U$18066 ( \18273 , \8835 , \3357 );
and \U$18067 ( \18274 , \9169 , \3255 );
nor \U$18068 ( \18275 , \18273 , \18274 );
xnor \U$18069 ( \18276 , \18275 , \3156 );
and \U$18070 ( \18277 , \8349 , \3813 );
and \U$18071 ( \18278 , \8652 , \3557 );
nor \U$18072 ( \18279 , \18277 , \18278 );
xnor \U$18073 ( \18280 , \18279 , \3562 );
xor \U$18074 ( \18281 , \18276 , \18280 );
and \U$18075 ( \18282 , \7700 , \4132 );
and \U$18076 ( \18283 , \8057 , \4012 );
nor \U$18077 ( \18284 , \18282 , \18283 );
xnor \U$18078 ( \18285 , \18284 , \3925 );
xor \U$18079 ( \18286 , \18281 , \18285 );
xor \U$18080 ( \18287 , \18272 , \18286 );
xor \U$18081 ( \18288 , \18243 , \18287 );
xor \U$18082 ( \18289 , \18227 , \18288 );
and \U$18083 ( \18290 , \18105 , \18109 );
and \U$18084 ( \18291 , \18109 , \18114 );
and \U$18085 ( \18292 , \18105 , \18114 );
or \U$18086 ( \18293 , \18290 , \18291 , \18292 );
and \U$18087 ( \18294 , \18011 , \18015 );
and \U$18088 ( \18295 , \18015 , \18020 );
and \U$18089 ( \18296 , \18011 , \18020 );
or \U$18090 ( \18297 , \18294 , \18295 , \18296 );
xor \U$18091 ( \18298 , \18293 , \18297 );
and \U$18092 ( \18299 , \18091 , \18095 );
and \U$18093 ( \18300 , \18095 , \18100 );
and \U$18094 ( \18301 , \18091 , \18100 );
or \U$18095 ( \18302 , \18299 , \18300 , \18301 );
xor \U$18096 ( \18303 , \18298 , \18302 );
and \U$18097 ( \18304 , \18119 , \18123 );
and \U$18098 ( \18305 , \18123 , \18128 );
and \U$18099 ( \18306 , \18119 , \18128 );
or \U$18100 ( \18307 , \18304 , \18305 , \18306 );
and \U$18101 ( \18308 , \18151 , \18155 );
and \U$18102 ( \18309 , \18155 , \18160 );
and \U$18103 ( \18310 , \18151 , \18160 );
or \U$18104 ( \18311 , \18308 , \18309 , \18310 );
xor \U$18105 ( \18312 , \18307 , \18311 );
and \U$18106 ( \18313 , \18134 , \18138 );
and \U$18107 ( \18314 , \18138 , \18143 );
and \U$18108 ( \18315 , \18134 , \18143 );
or \U$18109 ( \18316 , \18313 , \18314 , \18315 );
xor \U$18110 ( \18317 , \18312 , \18316 );
xor \U$18111 ( \18318 , \18303 , \18317 );
and \U$18112 ( \18319 , \2366 , \10118 );
and \U$18113 ( \18320 , \3143 , \9333 );
and \U$18114 ( \18321 , \3395 , \9006 );
nor \U$18115 ( \18322 , \18320 , \18321 );
xnor \U$18116 ( \18323 , \18322 , \8848 );
and \U$18117 ( \18324 , \2826 , \9765 );
and \U$18118 ( \18325 , \3037 , \9644 );
nor \U$18119 ( \18326 , \18324 , \18325 );
xnor \U$18120 ( \18327 , \18326 , \9478 );
xor \U$18121 ( \18328 , \18323 , \18327 );
and \U$18122 ( \18329 , \2521 , \10408 );
and \U$18123 ( \18330 , \2757 , \10116 );
nor \U$18124 ( \18331 , \18329 , \18330 );
xnor \U$18125 ( \18332 , \18331 , \10121 );
xor \U$18126 ( \18333 , \18328 , \18332 );
xor \U$18127 ( \18334 , \18319 , \18333 );
and \U$18128 ( \18335 , \4364 , \7489 );
and \U$18129 ( \18336 , \4654 , \7137 );
nor \U$18130 ( \18337 , \18335 , \18336 );
xnor \U$18131 ( \18338 , \18337 , \7142 );
and \U$18132 ( \18339 , \3912 , \8019 );
and \U$18133 ( \18340 , \4160 , \7830 );
nor \U$18134 ( \18341 , \18339 , \18340 );
xnor \U$18135 ( \18342 , \18341 , \7713 );
xor \U$18136 ( \18343 , \18338 , \18342 );
and \U$18137 ( \18344 , \3646 , \8540 );
and \U$18138 ( \18345 , \3736 , \8292 );
nor \U$18139 ( \18346 , \18344 , \18345 );
xnor \U$18140 ( \18347 , \18346 , \8297 );
xor \U$18141 ( \18348 , \18343 , \18347 );
xor \U$18142 ( \18349 , \18334 , \18348 );
xor \U$18143 ( \18350 , \18318 , \18349 );
xor \U$18144 ( \18351 , \18289 , \18350 );
xor \U$18145 ( \18352 , \18216 , \18351 );
xor \U$18146 ( \18353 , \18207 , \18352 );
and \U$18147 ( \18354 , \17989 , \18023 );
and \U$18148 ( \18355 , \18023 , \18166 );
and \U$18149 ( \18356 , \17989 , \18166 );
or \U$18150 ( \18357 , \18354 , \18355 , \18356 );
xor \U$18151 ( \18358 , \18353 , \18357 );
and \U$18152 ( \18359 , \18167 , \18171 );
and \U$18153 ( \18360 , \18172 , \18175 );
or \U$18154 ( \18361 , \18359 , \18360 );
xor \U$18155 ( \18362 , \18358 , \18361 );
buf g54e1_GF_PartitionCandidate( \18363_nG54e1 , \18362 );
buf \U$18156 ( \18364 , \18363_nG54e1 );
and \U$18157 ( \18365 , \18186 , \18190 );
and \U$18158 ( \18366 , \18190 , \18205 );
and \U$18159 ( \18367 , \18186 , \18205 );
or \U$18160 ( \18368 , \18365 , \18366 , \18367 );
and \U$18161 ( \18369 , \18211 , \18215 );
and \U$18162 ( \18370 , \18215 , \18351 );
and \U$18163 ( \18371 , \18211 , \18351 );
or \U$18164 ( \18372 , \18369 , \18370 , \18371 );
and \U$18165 ( \18373 , \18220 , \18224 );
and \U$18166 ( \18374 , \18224 , \18226 );
and \U$18167 ( \18375 , \18220 , \18226 );
or \U$18168 ( \18376 , \18373 , \18374 , \18375 );
and \U$18169 ( \18377 , \18231 , \18242 );
and \U$18170 ( \18378 , \18242 , \18287 );
and \U$18171 ( \18379 , \18231 , \18287 );
or \U$18172 ( \18380 , \18377 , \18378 , \18379 );
xor \U$18173 ( \18381 , \18376 , \18380 );
and \U$18174 ( \18382 , \18303 , \18317 );
and \U$18175 ( \18383 , \18317 , \18349 );
and \U$18176 ( \18384 , \18303 , \18349 );
or \U$18177 ( \18385 , \18382 , \18383 , \18384 );
xor \U$18178 ( \18386 , \18381 , \18385 );
xor \U$18179 ( \18387 , \18372 , \18386 );
and \U$18180 ( \18388 , \18195 , \18199 );
and \U$18181 ( \18389 , \18199 , \18204 );
and \U$18182 ( \18390 , \18195 , \18204 );
or \U$18183 ( \18391 , \18388 , \18389 , \18390 );
and \U$18184 ( \18392 , \18227 , \18288 );
and \U$18185 ( \18393 , \18288 , \18350 );
and \U$18186 ( \18394 , \18227 , \18350 );
or \U$18187 ( \18395 , \18392 , \18393 , \18394 );
xor \U$18188 ( \18396 , \18391 , \18395 );
and \U$18189 ( \18397 , \18293 , \18297 );
and \U$18190 ( \18398 , \18297 , \18302 );
and \U$18191 ( \18399 , \18293 , \18302 );
or \U$18192 ( \18400 , \18397 , \18398 , \18399 );
and \U$18193 ( \18401 , \18307 , \18311 );
and \U$18194 ( \18402 , \18311 , \18316 );
and \U$18195 ( \18403 , \18307 , \18316 );
or \U$18196 ( \18404 , \18401 , \18402 , \18403 );
xor \U$18197 ( \18405 , \18400 , \18404 );
and \U$18198 ( \18406 , \18319 , \18333 );
and \U$18199 ( \18407 , \18333 , \18348 );
and \U$18200 ( \18408 , \18319 , \18348 );
or \U$18201 ( \18409 , \18406 , \18407 , \18408 );
xor \U$18202 ( \18410 , \18405 , \18409 );
and \U$18203 ( \18411 , \18257 , \18271 );
and \U$18204 ( \18412 , \18271 , \18286 );
and \U$18205 ( \18413 , \18257 , \18286 );
or \U$18206 ( \18414 , \18411 , \18412 , \18413 );
and \U$18207 ( \18415 , \10584 , \2669 );
not \U$18208 ( \18416 , \18415 );
xnor \U$18209 ( \18417 , \18416 , \2534 );
and \U$18210 ( \18418 , \9897 , \3103 );
and \U$18211 ( \18419 , \10206 , \2934 );
nor \U$18212 ( \18420 , \18418 , \18419 );
xnor \U$18213 ( \18421 , \18420 , \2839 );
xor \U$18214 ( \18422 , \18417 , \18421 );
and \U$18215 ( \18423 , \9169 , \3357 );
and \U$18216 ( \18424 , \9465 , \3255 );
nor \U$18217 ( \18425 , \18423 , \18424 );
xnor \U$18218 ( \18426 , \18425 , \3156 );
xor \U$18219 ( \18427 , \18422 , \18426 );
xor \U$18220 ( \18428 , \18414 , \18427 );
and \U$18221 ( \18429 , \8652 , \3813 );
and \U$18222 ( \18430 , \8835 , \3557 );
nor \U$18223 ( \18431 , \18429 , \18430 );
xnor \U$18224 ( \18432 , \18431 , \3562 );
and \U$18225 ( \18433 , \8057 , \4132 );
and \U$18226 ( \18434 , \8349 , \4012 );
nor \U$18227 ( \18435 , \18433 , \18434 );
xnor \U$18228 ( \18436 , \18435 , \3925 );
xor \U$18229 ( \18437 , \18432 , \18436 );
and \U$18230 ( \18438 , \7556 , \4581 );
and \U$18231 ( \18439 , \7700 , \4424 );
nor \U$18232 ( \18440 , \18438 , \18439 );
xnor \U$18233 ( \18441 , \18440 , \4377 );
xor \U$18234 ( \18442 , \18437 , \18441 );
and \U$18235 ( \18443 , \6945 , \5011 );
and \U$18236 ( \18444 , \7231 , \4878 );
nor \U$18237 ( \18445 , \18443 , \18444 );
xnor \U$18238 ( \18446 , \18445 , \4762 );
and \U$18239 ( \18447 , \6514 , \5485 );
and \U$18240 ( \18448 , \6790 , \5275 );
nor \U$18241 ( \18449 , \18447 , \18448 );
xnor \U$18242 ( \18450 , \18449 , \5169 );
xor \U$18243 ( \18451 , \18446 , \18450 );
and \U$18244 ( \18452 , \6030 , \5996 );
and \U$18245 ( \18453 , \6281 , \5695 );
nor \U$18246 ( \18454 , \18452 , \18453 );
xnor \U$18247 ( \18455 , \18454 , \5687 );
xor \U$18248 ( \18456 , \18451 , \18455 );
xor \U$18249 ( \18457 , \18442 , \18456 );
and \U$18250 ( \18458 , \5469 , \6401 );
and \U$18251 ( \18459 , \5674 , \6143 );
nor \U$18252 ( \18460 , \18458 , \18459 );
xnor \U$18253 ( \18461 , \18460 , \6148 );
and \U$18254 ( \18462 , \4922 , \7055 );
and \U$18255 ( \18463 , \5156 , \6675 );
nor \U$18256 ( \18464 , \18462 , \18463 );
xnor \U$18257 ( \18465 , \18464 , \6680 );
xor \U$18258 ( \18466 , \18461 , \18465 );
and \U$18259 ( \18467 , \4654 , \7489 );
and \U$18260 ( \18468 , \4749 , \7137 );
nor \U$18261 ( \18469 , \18467 , \18468 );
xnor \U$18262 ( \18470 , \18469 , \7142 );
xor \U$18263 ( \18471 , \18466 , \18470 );
xor \U$18264 ( \18472 , \18457 , \18471 );
xor \U$18265 ( \18473 , \18428 , \18472 );
xor \U$18266 ( \18474 , \18410 , \18473 );
and \U$18267 ( \18475 , \18247 , \18251 );
and \U$18268 ( \18476 , \18251 , \18256 );
and \U$18269 ( \18477 , \18247 , \18256 );
or \U$18270 ( \18478 , \18475 , \18476 , \18477 );
and \U$18271 ( \18479 , \18232 , \18236 );
and \U$18272 ( \18480 , \18236 , \18241 );
and \U$18273 ( \18481 , \18232 , \18241 );
or \U$18274 ( \18482 , \18479 , \18480 , \18481 );
xor \U$18275 ( \18483 , \18478 , \18482 );
and \U$18276 ( \18484 , \18276 , \18280 );
and \U$18277 ( \18485 , \18280 , \18285 );
and \U$18278 ( \18486 , \18276 , \18285 );
or \U$18279 ( \18487 , \18484 , \18485 , \18486 );
xor \U$18280 ( \18488 , \18483 , \18487 );
and \U$18281 ( \18489 , \18323 , \18327 );
and \U$18282 ( \18490 , \18327 , \18332 );
and \U$18283 ( \18491 , \18323 , \18332 );
or \U$18284 ( \18492 , \18489 , \18490 , \18491 );
and \U$18285 ( \18493 , \18261 , \18265 );
and \U$18286 ( \18494 , \18265 , \18270 );
and \U$18287 ( \18495 , \18261 , \18270 );
or \U$18288 ( \18496 , \18493 , \18494 , \18495 );
xor \U$18289 ( \18497 , \18492 , \18496 );
and \U$18290 ( \18498 , \18338 , \18342 );
and \U$18291 ( \18499 , \18342 , \18347 );
and \U$18292 ( \18500 , \18338 , \18347 );
or \U$18293 ( \18501 , \18498 , \18499 , \18500 );
xor \U$18294 ( \18502 , \18497 , \18501 );
xor \U$18295 ( \18503 , \18488 , \18502 );
and \U$18296 ( \18504 , \3037 , \9765 );
and \U$18297 ( \18505 , \3143 , \9644 );
nor \U$18298 ( \18506 , \18504 , \18505 );
xnor \U$18299 ( \18507 , \18506 , \9478 );
and \U$18300 ( \18508 , \2757 , \10408 );
and \U$18301 ( \18509 , \2826 , \10116 );
nor \U$18302 ( \18510 , \18508 , \18509 );
xnor \U$18303 ( \18511 , \18510 , \10121 );
xor \U$18304 ( \18512 , \18507 , \18511 );
and \U$18305 ( \18513 , \2521 , \10118 );
xor \U$18306 ( \18514 , \18512 , \18513 );
and \U$18307 ( \18515 , \4160 , \8019 );
and \U$18308 ( \18516 , \4364 , \7830 );
nor \U$18309 ( \18517 , \18515 , \18516 );
xnor \U$18310 ( \18518 , \18517 , \7713 );
and \U$18311 ( \18519 , \3736 , \8540 );
and \U$18312 ( \18520 , \3912 , \8292 );
nor \U$18313 ( \18521 , \18519 , \18520 );
xnor \U$18314 ( \18522 , \18521 , \8297 );
xor \U$18315 ( \18523 , \18518 , \18522 );
and \U$18316 ( \18524 , \3395 , \9333 );
and \U$18317 ( \18525 , \3646 , \9006 );
nor \U$18318 ( \18526 , \18524 , \18525 );
xnor \U$18319 ( \18527 , \18526 , \8848 );
xor \U$18320 ( \18528 , \18523 , \18527 );
xnor \U$18321 ( \18529 , \18514 , \18528 );
xor \U$18322 ( \18530 , \18503 , \18529 );
xor \U$18323 ( \18531 , \18474 , \18530 );
xor \U$18324 ( \18532 , \18396 , \18531 );
xor \U$18325 ( \18533 , \18387 , \18532 );
xor \U$18326 ( \18534 , \18368 , \18533 );
and \U$18327 ( \18535 , \18182 , \18206 );
and \U$18328 ( \18536 , \18206 , \18352 );
and \U$18329 ( \18537 , \18182 , \18352 );
or \U$18330 ( \18538 , \18535 , \18536 , \18537 );
xor \U$18331 ( \18539 , \18534 , \18538 );
and \U$18332 ( \18540 , \18353 , \18357 );
and \U$18333 ( \18541 , \18358 , \18361 );
or \U$18334 ( \18542 , \18540 , \18541 );
xor \U$18335 ( \18543 , \18539 , \18542 );
buf g54df_GF_PartitionCandidate( \18544_nG54df , \18543 );
buf \U$18336 ( \18545 , \18544_nG54df );
and \U$18337 ( \18546 , \18372 , \18386 );
and \U$18338 ( \18547 , \18386 , \18532 );
and \U$18339 ( \18548 , \18372 , \18532 );
or \U$18340 ( \18549 , \18546 , \18547 , \18548 );
and \U$18341 ( \18550 , \18391 , \18395 );
and \U$18342 ( \18551 , \18395 , \18531 );
and \U$18343 ( \18552 , \18391 , \18531 );
or \U$18344 ( \18553 , \18550 , \18551 , \18552 );
and \U$18345 ( \18554 , \18400 , \18404 );
and \U$18346 ( \18555 , \18404 , \18409 );
and \U$18347 ( \18556 , \18400 , \18409 );
or \U$18348 ( \18557 , \18554 , \18555 , \18556 );
and \U$18349 ( \18558 , \18414 , \18427 );
and \U$18350 ( \18559 , \18427 , \18472 );
and \U$18351 ( \18560 , \18414 , \18472 );
or \U$18352 ( \18561 , \18558 , \18559 , \18560 );
xor \U$18353 ( \18562 , \18557 , \18561 );
and \U$18354 ( \18563 , \18488 , \18502 );
and \U$18355 ( \18564 , \18502 , \18529 );
and \U$18356 ( \18565 , \18488 , \18529 );
or \U$18357 ( \18566 , \18563 , \18564 , \18565 );
xor \U$18358 ( \18567 , \18562 , \18566 );
xor \U$18359 ( \18568 , \18553 , \18567 );
and \U$18360 ( \18569 , \18376 , \18380 );
and \U$18361 ( \18570 , \18380 , \18385 );
and \U$18362 ( \18571 , \18376 , \18385 );
or \U$18363 ( \18572 , \18569 , \18570 , \18571 );
and \U$18364 ( \18573 , \18410 , \18473 );
and \U$18365 ( \18574 , \18473 , \18530 );
and \U$18366 ( \18575 , \18410 , \18530 );
or \U$18367 ( \18576 , \18573 , \18574 , \18575 );
xor \U$18368 ( \18577 , \18572 , \18576 );
and \U$18369 ( \18578 , \18478 , \18482 );
and \U$18370 ( \18579 , \18482 , \18487 );
and \U$18371 ( \18580 , \18478 , \18487 );
or \U$18372 ( \18581 , \18578 , \18579 , \18580 );
and \U$18373 ( \18582 , \18492 , \18496 );
and \U$18374 ( \18583 , \18496 , \18501 );
and \U$18375 ( \18584 , \18492 , \18501 );
or \U$18376 ( \18585 , \18582 , \18583 , \18584 );
xor \U$18377 ( \18586 , \18581 , \18585 );
or \U$18378 ( \18587 , \18514 , \18528 );
xor \U$18379 ( \18588 , \18586 , \18587 );
and \U$18380 ( \18589 , \18442 , \18456 );
and \U$18381 ( \18590 , \18456 , \18471 );
and \U$18382 ( \18591 , \18442 , \18471 );
or \U$18383 ( \18592 , \18589 , \18590 , \18591 );
and \U$18384 ( \18593 , \3143 , \9765 );
and \U$18385 ( \18594 , \3395 , \9644 );
nor \U$18386 ( \18595 , \18593 , \18594 );
xnor \U$18387 ( \18596 , \18595 , \9478 );
and \U$18388 ( \18597 , \2826 , \10408 );
and \U$18389 ( \18598 , \3037 , \10116 );
nor \U$18390 ( \18599 , \18597 , \18598 );
xnor \U$18391 ( \18600 , \18599 , \10121 );
xor \U$18392 ( \18601 , \18596 , \18600 );
and \U$18393 ( \18602 , \2757 , \10118 );
xor \U$18394 ( \18603 , \18601 , \18602 );
and \U$18395 ( \18604 , \4364 , \8019 );
and \U$18396 ( \18605 , \4654 , \7830 );
nor \U$18397 ( \18606 , \18604 , \18605 );
xnor \U$18398 ( \18607 , \18606 , \7713 );
and \U$18399 ( \18608 , \3912 , \8540 );
and \U$18400 ( \18609 , \4160 , \8292 );
nor \U$18401 ( \18610 , \18608 , \18609 );
xnor \U$18402 ( \18611 , \18610 , \8297 );
xor \U$18403 ( \18612 , \18607 , \18611 );
and \U$18404 ( \18613 , \3646 , \9333 );
and \U$18405 ( \18614 , \3736 , \9006 );
nor \U$18406 ( \18615 , \18613 , \18614 );
xnor \U$18407 ( \18616 , \18615 , \8848 );
xor \U$18408 ( \18617 , \18612 , \18616 );
xor \U$18409 ( \18618 , \18603 , \18617 );
and \U$18410 ( \18619 , \5674 , \6401 );
and \U$18411 ( \18620 , \6030 , \6143 );
nor \U$18412 ( \18621 , \18619 , \18620 );
xnor \U$18413 ( \18622 , \18621 , \6148 );
and \U$18414 ( \18623 , \5156 , \7055 );
and \U$18415 ( \18624 , \5469 , \6675 );
nor \U$18416 ( \18625 , \18623 , \18624 );
xnor \U$18417 ( \18626 , \18625 , \6680 );
xor \U$18418 ( \18627 , \18622 , \18626 );
and \U$18419 ( \18628 , \4749 , \7489 );
and \U$18420 ( \18629 , \4922 , \7137 );
nor \U$18421 ( \18630 , \18628 , \18629 );
xnor \U$18422 ( \18631 , \18630 , \7142 );
xor \U$18423 ( \18632 , \18627 , \18631 );
xor \U$18424 ( \18633 , \18618 , \18632 );
xor \U$18425 ( \18634 , \18592 , \18633 );
and \U$18426 ( \18635 , \8835 , \3813 );
and \U$18427 ( \18636 , \9169 , \3557 );
nor \U$18428 ( \18637 , \18635 , \18636 );
xnor \U$18429 ( \18638 , \18637 , \3562 );
and \U$18430 ( \18639 , \8349 , \4132 );
and \U$18431 ( \18640 , \8652 , \4012 );
nor \U$18432 ( \18641 , \18639 , \18640 );
xnor \U$18433 ( \18642 , \18641 , \3925 );
xor \U$18434 ( \18643 , \18638 , \18642 );
and \U$18435 ( \18644 , \7700 , \4581 );
and \U$18436 ( \18645 , \8057 , \4424 );
nor \U$18437 ( \18646 , \18644 , \18645 );
xnor \U$18438 ( \18647 , \18646 , \4377 );
xor \U$18439 ( \18648 , \18643 , \18647 );
and \U$18440 ( \18649 , \7231 , \5011 );
and \U$18441 ( \18650 , \7556 , \4878 );
nor \U$18442 ( \18651 , \18649 , \18650 );
xnor \U$18443 ( \18652 , \18651 , \4762 );
and \U$18444 ( \18653 , \6790 , \5485 );
and \U$18445 ( \18654 , \6945 , \5275 );
nor \U$18446 ( \18655 , \18653 , \18654 );
xnor \U$18447 ( \18656 , \18655 , \5169 );
xor \U$18448 ( \18657 , \18652 , \18656 );
and \U$18449 ( \18658 , \6281 , \5996 );
and \U$18450 ( \18659 , \6514 , \5695 );
nor \U$18451 ( \18660 , \18658 , \18659 );
xnor \U$18452 ( \18661 , \18660 , \5687 );
xor \U$18453 ( \18662 , \18657 , \18661 );
xor \U$18454 ( \18663 , \18648 , \18662 );
not \U$18455 ( \18664 , \2534 );
and \U$18456 ( \18665 , \10206 , \3103 );
and \U$18457 ( \18666 , \10584 , \2934 );
nor \U$18458 ( \18667 , \18665 , \18666 );
xnor \U$18459 ( \18668 , \18667 , \2839 );
xor \U$18460 ( \18669 , \18664 , \18668 );
and \U$18461 ( \18670 , \9465 , \3357 );
and \U$18462 ( \18671 , \9897 , \3255 );
nor \U$18463 ( \18672 , \18670 , \18671 );
xnor \U$18464 ( \18673 , \18672 , \3156 );
xor \U$18465 ( \18674 , \18669 , \18673 );
xor \U$18466 ( \18675 , \18663 , \18674 );
xor \U$18467 ( \18676 , \18634 , \18675 );
xor \U$18468 ( \18677 , \18588 , \18676 );
and \U$18469 ( \18678 , \18507 , \18511 );
and \U$18470 ( \18679 , \18511 , \18513 );
and \U$18471 ( \18680 , \18507 , \18513 );
or \U$18472 ( \18681 , \18678 , \18679 , \18680 );
and \U$18473 ( \18682 , \18518 , \18522 );
and \U$18474 ( \18683 , \18522 , \18527 );
and \U$18475 ( \18684 , \18518 , \18527 );
or \U$18476 ( \18685 , \18682 , \18683 , \18684 );
xor \U$18477 ( \18686 , \18681 , \18685 );
and \U$18478 ( \18687 , \18461 , \18465 );
and \U$18479 ( \18688 , \18465 , \18470 );
and \U$18480 ( \18689 , \18461 , \18470 );
or \U$18481 ( \18690 , \18687 , \18688 , \18689 );
xor \U$18482 ( \18691 , \18686 , \18690 );
and \U$18483 ( \18692 , \18432 , \18436 );
and \U$18484 ( \18693 , \18436 , \18441 );
and \U$18485 ( \18694 , \18432 , \18441 );
or \U$18486 ( \18695 , \18692 , \18693 , \18694 );
and \U$18487 ( \18696 , \18417 , \18421 );
and \U$18488 ( \18697 , \18421 , \18426 );
and \U$18489 ( \18698 , \18417 , \18426 );
or \U$18490 ( \18699 , \18696 , \18697 , \18698 );
xor \U$18491 ( \18700 , \18695 , \18699 );
and \U$18492 ( \18701 , \18446 , \18450 );
and \U$18493 ( \18702 , \18450 , \18455 );
and \U$18494 ( \18703 , \18446 , \18455 );
or \U$18495 ( \18704 , \18701 , \18702 , \18703 );
xor \U$18496 ( \18705 , \18700 , \18704 );
xor \U$18497 ( \18706 , \18691 , \18705 );
xor \U$18498 ( \18707 , \18677 , \18706 );
xor \U$18499 ( \18708 , \18577 , \18707 );
xor \U$18500 ( \18709 , \18568 , \18708 );
xor \U$18501 ( \18710 , \18549 , \18709 );
and \U$18502 ( \18711 , \18368 , \18533 );
xor \U$18503 ( \18712 , \18710 , \18711 );
and \U$18504 ( \18713 , \18534 , \18538 );
and \U$18505 ( \18714 , \18539 , \18542 );
or \U$18506 ( \18715 , \18713 , \18714 );
xor \U$18507 ( \18716 , \18712 , \18715 );
buf g54dd_GF_PartitionCandidate( \18717_nG54dd , \18716 );
buf \U$18508 ( \18718 , \18717_nG54dd );
and \U$18509 ( \18719 , \18553 , \18567 );
and \U$18510 ( \18720 , \18567 , \18708 );
and \U$18511 ( \18721 , \18553 , \18708 );
or \U$18512 ( \18722 , \18719 , \18720 , \18721 );
and \U$18513 ( \18723 , \18572 , \18576 );
and \U$18514 ( \18724 , \18576 , \18707 );
and \U$18515 ( \18725 , \18572 , \18707 );
or \U$18516 ( \18726 , \18723 , \18724 , \18725 );
and \U$18517 ( \18727 , \18581 , \18585 );
and \U$18518 ( \18728 , \18585 , \18587 );
and \U$18519 ( \18729 , \18581 , \18587 );
or \U$18520 ( \18730 , \18727 , \18728 , \18729 );
and \U$18521 ( \18731 , \18592 , \18633 );
and \U$18522 ( \18732 , \18633 , \18675 );
and \U$18523 ( \18733 , \18592 , \18675 );
or \U$18524 ( \18734 , \18731 , \18732 , \18733 );
xor \U$18525 ( \18735 , \18730 , \18734 );
and \U$18526 ( \18736 , \18691 , \18705 );
xor \U$18527 ( \18737 , \18735 , \18736 );
xor \U$18528 ( \18738 , \18726 , \18737 );
and \U$18529 ( \18739 , \18557 , \18561 );
and \U$18530 ( \18740 , \18561 , \18566 );
and \U$18531 ( \18741 , \18557 , \18566 );
or \U$18532 ( \18742 , \18739 , \18740 , \18741 );
and \U$18533 ( \18743 , \18588 , \18676 );
and \U$18534 ( \18744 , \18676 , \18706 );
and \U$18535 ( \18745 , \18588 , \18706 );
or \U$18536 ( \18746 , \18743 , \18744 , \18745 );
xor \U$18537 ( \18747 , \18742 , \18746 );
and \U$18538 ( \18748 , \18681 , \18685 );
and \U$18539 ( \18749 , \18685 , \18690 );
and \U$18540 ( \18750 , \18681 , \18690 );
or \U$18541 ( \18751 , \18748 , \18749 , \18750 );
and \U$18542 ( \18752 , \18695 , \18699 );
and \U$18543 ( \18753 , \18699 , \18704 );
and \U$18544 ( \18754 , \18695 , \18704 );
or \U$18545 ( \18755 , \18752 , \18753 , \18754 );
xor \U$18546 ( \18756 , \18751 , \18755 );
and \U$18547 ( \18757 , \18603 , \18617 );
and \U$18548 ( \18758 , \18617 , \18632 );
and \U$18549 ( \18759 , \18603 , \18632 );
or \U$18550 ( \18760 , \18757 , \18758 , \18759 );
xor \U$18551 ( \18761 , \18756 , \18760 );
and \U$18552 ( \18762 , \18648 , \18662 );
and \U$18553 ( \18763 , \18662 , \18674 );
and \U$18554 ( \18764 , \18648 , \18674 );
or \U$18555 ( \18765 , \18762 , \18763 , \18764 );
and \U$18556 ( \18766 , \10584 , \3103 );
not \U$18557 ( \18767 , \18766 );
xnor \U$18558 ( \18768 , \18767 , \2839 );
and \U$18559 ( \18769 , \9897 , \3357 );
and \U$18560 ( \18770 , \10206 , \3255 );
nor \U$18561 ( \18771 , \18769 , \18770 );
xnor \U$18562 ( \18772 , \18771 , \3156 );
xor \U$18563 ( \18773 , \18768 , \18772 );
and \U$18564 ( \18774 , \9169 , \3813 );
and \U$18565 ( \18775 , \9465 , \3557 );
nor \U$18566 ( \18776 , \18774 , \18775 );
xnor \U$18567 ( \18777 , \18776 , \3562 );
xor \U$18568 ( \18778 , \18773 , \18777 );
and \U$18569 ( \18779 , \6945 , \5485 );
and \U$18570 ( \18780 , \7231 , \5275 );
nor \U$18571 ( \18781 , \18779 , \18780 );
xnor \U$18572 ( \18782 , \18781 , \5169 );
and \U$18573 ( \18783 , \6514 , \5996 );
and \U$18574 ( \18784 , \6790 , \5695 );
nor \U$18575 ( \18785 , \18783 , \18784 );
xnor \U$18576 ( \18786 , \18785 , \5687 );
xor \U$18577 ( \18787 , \18782 , \18786 );
and \U$18578 ( \18788 , \6030 , \6401 );
and \U$18579 ( \18789 , \6281 , \6143 );
nor \U$18580 ( \18790 , \18788 , \18789 );
xnor \U$18581 ( \18791 , \18790 , \6148 );
xor \U$18582 ( \18792 , \18787 , \18791 );
xor \U$18583 ( \18793 , \18778 , \18792 );
and \U$18584 ( \18794 , \8652 , \4132 );
and \U$18585 ( \18795 , \8835 , \4012 );
nor \U$18586 ( \18796 , \18794 , \18795 );
xnor \U$18587 ( \18797 , \18796 , \3925 );
and \U$18588 ( \18798 , \8057 , \4581 );
and \U$18589 ( \18799 , \8349 , \4424 );
nor \U$18590 ( \18800 , \18798 , \18799 );
xnor \U$18591 ( \18801 , \18800 , \4377 );
xor \U$18592 ( \18802 , \18797 , \18801 );
and \U$18593 ( \18803 , \7556 , \5011 );
and \U$18594 ( \18804 , \7700 , \4878 );
nor \U$18595 ( \18805 , \18803 , \18804 );
xnor \U$18596 ( \18806 , \18805 , \4762 );
xor \U$18597 ( \18807 , \18802 , \18806 );
xor \U$18598 ( \18808 , \18793 , \18807 );
xor \U$18599 ( \18809 , \18765 , \18808 );
and \U$18600 ( \18810 , \4160 , \8540 );
and \U$18601 ( \18811 , \4364 , \8292 );
nor \U$18602 ( \18812 , \18810 , \18811 );
xnor \U$18603 ( \18813 , \18812 , \8297 );
and \U$18604 ( \18814 , \3736 , \9333 );
and \U$18605 ( \18815 , \3912 , \9006 );
nor \U$18606 ( \18816 , \18814 , \18815 );
xnor \U$18607 ( \18817 , \18816 , \8848 );
xor \U$18608 ( \18818 , \18813 , \18817 );
and \U$18609 ( \18819 , \3395 , \9765 );
and \U$18610 ( \18820 , \3646 , \9644 );
nor \U$18611 ( \18821 , \18819 , \18820 );
xnor \U$18612 ( \18822 , \18821 , \9478 );
xor \U$18613 ( \18823 , \18818 , \18822 );
and \U$18614 ( \18824 , \5469 , \7055 );
and \U$18615 ( \18825 , \5674 , \6675 );
nor \U$18616 ( \18826 , \18824 , \18825 );
xnor \U$18617 ( \18827 , \18826 , \6680 );
and \U$18618 ( \18828 , \4922 , \7489 );
and \U$18619 ( \18829 , \5156 , \7137 );
nor \U$18620 ( \18830 , \18828 , \18829 );
xnor \U$18621 ( \18831 , \18830 , \7142 );
xor \U$18622 ( \18832 , \18827 , \18831 );
and \U$18623 ( \18833 , \4654 , \8019 );
and \U$18624 ( \18834 , \4749 , \7830 );
nor \U$18625 ( \18835 , \18833 , \18834 );
xnor \U$18626 ( \18836 , \18835 , \7713 );
xor \U$18627 ( \18837 , \18832 , \18836 );
xor \U$18628 ( \18838 , \18823 , \18837 );
and \U$18629 ( \18839 , \3037 , \10408 );
and \U$18630 ( \18840 , \3143 , \10116 );
nor \U$18631 ( \18841 , \18839 , \18840 );
xnor \U$18632 ( \18842 , \18841 , \10121 );
and \U$18633 ( \18843 , \2826 , \10118 );
xnor \U$18634 ( \18844 , \18842 , \18843 );
xor \U$18635 ( \18845 , \18838 , \18844 );
xor \U$18636 ( \18846 , \18809 , \18845 );
xor \U$18637 ( \18847 , \18761 , \18846 );
and \U$18638 ( \18848 , \18638 , \18642 );
and \U$18639 ( \18849 , \18642 , \18647 );
and \U$18640 ( \18850 , \18638 , \18647 );
or \U$18641 ( \18851 , \18848 , \18849 , \18850 );
and \U$18642 ( \18852 , \18652 , \18656 );
and \U$18643 ( \18853 , \18656 , \18661 );
and \U$18644 ( \18854 , \18652 , \18661 );
or \U$18645 ( \18855 , \18852 , \18853 , \18854 );
xor \U$18646 ( \18856 , \18851 , \18855 );
and \U$18647 ( \18857 , \18664 , \18668 );
and \U$18648 ( \18858 , \18668 , \18673 );
and \U$18649 ( \18859 , \18664 , \18673 );
or \U$18650 ( \18860 , \18857 , \18858 , \18859 );
xor \U$18651 ( \18861 , \18856 , \18860 );
and \U$18652 ( \18862 , \18596 , \18600 );
and \U$18653 ( \18863 , \18600 , \18602 );
and \U$18654 ( \18864 , \18596 , \18602 );
or \U$18655 ( \18865 , \18862 , \18863 , \18864 );
and \U$18656 ( \18866 , \18607 , \18611 );
and \U$18657 ( \18867 , \18611 , \18616 );
and \U$18658 ( \18868 , \18607 , \18616 );
or \U$18659 ( \18869 , \18866 , \18867 , \18868 );
xor \U$18660 ( \18870 , \18865 , \18869 );
and \U$18661 ( \18871 , \18622 , \18626 );
and \U$18662 ( \18872 , \18626 , \18631 );
and \U$18663 ( \18873 , \18622 , \18631 );
or \U$18664 ( \18874 , \18871 , \18872 , \18873 );
xor \U$18665 ( \18875 , \18870 , \18874 );
xor \U$18666 ( \18876 , \18861 , \18875 );
xor \U$18667 ( \18877 , \18847 , \18876 );
xor \U$18668 ( \18878 , \18747 , \18877 );
xor \U$18669 ( \18879 , \18738 , \18878 );
xor \U$18670 ( \18880 , \18722 , \18879 );
and \U$18671 ( \18881 , \18549 , \18709 );
xor \U$18672 ( \18882 , \18880 , \18881 );
and \U$18673 ( \18883 , \18710 , \18711 );
and \U$18674 ( \18884 , \18712 , \18715 );
or \U$18675 ( \18885 , \18883 , \18884 );
xor \U$18676 ( \18886 , \18882 , \18885 );
buf g54db_GF_PartitionCandidate( \18887_nG54db , \18886 );
buf \U$18677 ( \18888 , \18887_nG54db );
and \U$18678 ( \18889 , \18726 , \18737 );
and \U$18679 ( \18890 , \18737 , \18878 );
and \U$18680 ( \18891 , \18726 , \18878 );
or \U$18681 ( \18892 , \18889 , \18890 , \18891 );
and \U$18682 ( \18893 , \18742 , \18746 );
and \U$18683 ( \18894 , \18746 , \18877 );
and \U$18684 ( \18895 , \18742 , \18877 );
or \U$18685 ( \18896 , \18893 , \18894 , \18895 );
and \U$18686 ( \18897 , \18751 , \18755 );
and \U$18687 ( \18898 , \18755 , \18760 );
and \U$18688 ( \18899 , \18751 , \18760 );
or \U$18689 ( \18900 , \18897 , \18898 , \18899 );
and \U$18690 ( \18901 , \18765 , \18808 );
and \U$18691 ( \18902 , \18808 , \18845 );
and \U$18692 ( \18903 , \18765 , \18845 );
or \U$18693 ( \18904 , \18901 , \18902 , \18903 );
xor \U$18694 ( \18905 , \18900 , \18904 );
and \U$18695 ( \18906 , \18861 , \18875 );
xor \U$18696 ( \18907 , \18905 , \18906 );
xor \U$18697 ( \18908 , \18896 , \18907 );
and \U$18698 ( \18909 , \18730 , \18734 );
and \U$18699 ( \18910 , \18734 , \18736 );
and \U$18700 ( \18911 , \18730 , \18736 );
or \U$18701 ( \18912 , \18909 , \18910 , \18911 );
and \U$18702 ( \18913 , \18761 , \18846 );
and \U$18703 ( \18914 , \18846 , \18876 );
and \U$18704 ( \18915 , \18761 , \18876 );
or \U$18705 ( \18916 , \18913 , \18914 , \18915 );
xor \U$18706 ( \18917 , \18912 , \18916 );
and \U$18707 ( \18918 , \18851 , \18855 );
and \U$18708 ( \18919 , \18855 , \18860 );
and \U$18709 ( \18920 , \18851 , \18860 );
or \U$18710 ( \18921 , \18918 , \18919 , \18920 );
and \U$18711 ( \18922 , \18865 , \18869 );
and \U$18712 ( \18923 , \18869 , \18874 );
and \U$18713 ( \18924 , \18865 , \18874 );
or \U$18714 ( \18925 , \18922 , \18923 , \18924 );
xor \U$18715 ( \18926 , \18921 , \18925 );
and \U$18716 ( \18927 , \18823 , \18837 );
and \U$18717 ( \18928 , \18837 , \18844 );
and \U$18718 ( \18929 , \18823 , \18844 );
or \U$18719 ( \18930 , \18927 , \18928 , \18929 );
xor \U$18720 ( \18931 , \18926 , \18930 );
and \U$18721 ( \18932 , \18778 , \18792 );
and \U$18722 ( \18933 , \18792 , \18807 );
and \U$18723 ( \18934 , \18778 , \18807 );
or \U$18724 ( \18935 , \18932 , \18933 , \18934 );
and \U$18725 ( \18936 , \7231 , \5485 );
and \U$18726 ( \18937 , \7556 , \5275 );
nor \U$18727 ( \18938 , \18936 , \18937 );
xnor \U$18728 ( \18939 , \18938 , \5169 );
and \U$18729 ( \18940 , \6790 , \5996 );
and \U$18730 ( \18941 , \6945 , \5695 );
nor \U$18731 ( \18942 , \18940 , \18941 );
xnor \U$18732 ( \18943 , \18942 , \5687 );
xor \U$18733 ( \18944 , \18939 , \18943 );
and \U$18734 ( \18945 , \6281 , \6401 );
and \U$18735 ( \18946 , \6514 , \6143 );
nor \U$18736 ( \18947 , \18945 , \18946 );
xnor \U$18737 ( \18948 , \18947 , \6148 );
xor \U$18738 ( \18949 , \18944 , \18948 );
not \U$18739 ( \18950 , \2839 );
and \U$18740 ( \18951 , \10206 , \3357 );
and \U$18741 ( \18952 , \10584 , \3255 );
nor \U$18742 ( \18953 , \18951 , \18952 );
xnor \U$18743 ( \18954 , \18953 , \3156 );
xor \U$18744 ( \18955 , \18950 , \18954 );
and \U$18745 ( \18956 , \9465 , \3813 );
and \U$18746 ( \18957 , \9897 , \3557 );
nor \U$18747 ( \18958 , \18956 , \18957 );
xnor \U$18748 ( \18959 , \18958 , \3562 );
xor \U$18749 ( \18960 , \18955 , \18959 );
xor \U$18750 ( \18961 , \18949 , \18960 );
and \U$18751 ( \18962 , \8835 , \4132 );
and \U$18752 ( \18963 , \9169 , \4012 );
nor \U$18753 ( \18964 , \18962 , \18963 );
xnor \U$18754 ( \18965 , \18964 , \3925 );
and \U$18755 ( \18966 , \8349 , \4581 );
and \U$18756 ( \18967 , \8652 , \4424 );
nor \U$18757 ( \18968 , \18966 , \18967 );
xnor \U$18758 ( \18969 , \18968 , \4377 );
xor \U$18759 ( \18970 , \18965 , \18969 );
and \U$18760 ( \18971 , \7700 , \5011 );
and \U$18761 ( \18972 , \8057 , \4878 );
nor \U$18762 ( \18973 , \18971 , \18972 );
xnor \U$18763 ( \18974 , \18973 , \4762 );
xor \U$18764 ( \18975 , \18970 , \18974 );
xor \U$18765 ( \18976 , \18961 , \18975 );
xor \U$18766 ( \18977 , \18935 , \18976 );
and \U$18767 ( \18978 , \4364 , \8540 );
and \U$18768 ( \18979 , \4654 , \8292 );
nor \U$18769 ( \18980 , \18978 , \18979 );
xnor \U$18770 ( \18981 , \18980 , \8297 );
and \U$18771 ( \18982 , \3912 , \9333 );
and \U$18772 ( \18983 , \4160 , \9006 );
nor \U$18773 ( \18984 , \18982 , \18983 );
xnor \U$18774 ( \18985 , \18984 , \8848 );
xor \U$18775 ( \18986 , \18981 , \18985 );
and \U$18776 ( \18987 , \3646 , \9765 );
and \U$18777 ( \18988 , \3736 , \9644 );
nor \U$18778 ( \18989 , \18987 , \18988 );
xnor \U$18779 ( \18990 , \18989 , \9478 );
xor \U$18780 ( \18991 , \18986 , \18990 );
and \U$18781 ( \18992 , \5674 , \7055 );
and \U$18782 ( \18993 , \6030 , \6675 );
nor \U$18783 ( \18994 , \18992 , \18993 );
xnor \U$18784 ( \18995 , \18994 , \6680 );
and \U$18785 ( \18996 , \5156 , \7489 );
and \U$18786 ( \18997 , \5469 , \7137 );
nor \U$18787 ( \18998 , \18996 , \18997 );
xnor \U$18788 ( \18999 , \18998 , \7142 );
xor \U$18789 ( \19000 , \18995 , \18999 );
and \U$18790 ( \19001 , \4749 , \8019 );
and \U$18791 ( \19002 , \4922 , \7830 );
nor \U$18792 ( \19003 , \19001 , \19002 );
xnor \U$18793 ( \19004 , \19003 , \7713 );
xor \U$18794 ( \19005 , \19000 , \19004 );
xor \U$18795 ( \19006 , \18991 , \19005 );
and \U$18796 ( \19007 , \3143 , \10408 );
and \U$18797 ( \19008 , \3395 , \10116 );
nor \U$18798 ( \19009 , \19007 , \19008 );
xnor \U$18799 ( \19010 , \19009 , \10121 );
and \U$18800 ( \19011 , \3037 , \10118 );
xor \U$18801 ( \19012 , \19010 , \19011 );
xor \U$18802 ( \19013 , \19006 , \19012 );
xor \U$18803 ( \19014 , \18977 , \19013 );
xor \U$18804 ( \19015 , \18931 , \19014 );
and \U$18805 ( \19016 , \18768 , \18772 );
and \U$18806 ( \19017 , \18772 , \18777 );
and \U$18807 ( \19018 , \18768 , \18777 );
or \U$18808 ( \19019 , \19016 , \19017 , \19018 );
and \U$18809 ( \19020 , \18782 , \18786 );
and \U$18810 ( \19021 , \18786 , \18791 );
and \U$18811 ( \19022 , \18782 , \18791 );
or \U$18812 ( \19023 , \19020 , \19021 , \19022 );
xor \U$18813 ( \19024 , \19019 , \19023 );
and \U$18814 ( \19025 , \18797 , \18801 );
and \U$18815 ( \19026 , \18801 , \18806 );
and \U$18816 ( \19027 , \18797 , \18806 );
or \U$18817 ( \19028 , \19025 , \19026 , \19027 );
xor \U$18818 ( \19029 , \19024 , \19028 );
and \U$18819 ( \19030 , \18813 , \18817 );
and \U$18820 ( \19031 , \18817 , \18822 );
and \U$18821 ( \19032 , \18813 , \18822 );
or \U$18822 ( \19033 , \19030 , \19031 , \19032 );
and \U$18823 ( \19034 , \18827 , \18831 );
and \U$18824 ( \19035 , \18831 , \18836 );
and \U$18825 ( \19036 , \18827 , \18836 );
or \U$18826 ( \19037 , \19034 , \19035 , \19036 );
xor \U$18827 ( \19038 , \19033 , \19037 );
or \U$18828 ( \19039 , \18842 , \18843 );
xor \U$18829 ( \19040 , \19038 , \19039 );
xor \U$18830 ( \19041 , \19029 , \19040 );
xor \U$18831 ( \19042 , \19015 , \19041 );
xor \U$18832 ( \19043 , \18917 , \19042 );
xor \U$18833 ( \19044 , \18908 , \19043 );
xor \U$18834 ( \19045 , \18892 , \19044 );
and \U$18835 ( \19046 , \18722 , \18879 );
xor \U$18836 ( \19047 , \19045 , \19046 );
and \U$18837 ( \19048 , \18880 , \18881 );
and \U$18838 ( \19049 , \18882 , \18885 );
or \U$18839 ( \19050 , \19048 , \19049 );
xor \U$18840 ( \19051 , \19047 , \19050 );
buf g54d9_GF_PartitionCandidate( \19052_nG54d9 , \19051 );
buf \U$18841 ( \19053 , \19052_nG54d9 );
and \U$18842 ( \19054 , \18896 , \18907 );
and \U$18843 ( \19055 , \18907 , \19043 );
and \U$18844 ( \19056 , \18896 , \19043 );
or \U$18845 ( \19057 , \19054 , \19055 , \19056 );
and \U$18846 ( \19058 , \18912 , \18916 );
and \U$18847 ( \19059 , \18916 , \19042 );
and \U$18848 ( \19060 , \18912 , \19042 );
or \U$18849 ( \19061 , \19058 , \19059 , \19060 );
and \U$18850 ( \19062 , \18921 , \18925 );
and \U$18851 ( \19063 , \18925 , \18930 );
and \U$18852 ( \19064 , \18921 , \18930 );
or \U$18853 ( \19065 , \19062 , \19063 , \19064 );
and \U$18854 ( \19066 , \18935 , \18976 );
and \U$18855 ( \19067 , \18976 , \19013 );
and \U$18856 ( \19068 , \18935 , \19013 );
or \U$18857 ( \19069 , \19066 , \19067 , \19068 );
xor \U$18858 ( \19070 , \19065 , \19069 );
and \U$18859 ( \19071 , \19029 , \19040 );
xor \U$18860 ( \19072 , \19070 , \19071 );
xor \U$18861 ( \19073 , \19061 , \19072 );
and \U$18862 ( \19074 , \18900 , \18904 );
and \U$18863 ( \19075 , \18904 , \18906 );
and \U$18864 ( \19076 , \18900 , \18906 );
or \U$18865 ( \19077 , \19074 , \19075 , \19076 );
and \U$18866 ( \19078 , \18931 , \19014 );
and \U$18867 ( \19079 , \19014 , \19041 );
and \U$18868 ( \19080 , \18931 , \19041 );
or \U$18869 ( \19081 , \19078 , \19079 , \19080 );
xor \U$18870 ( \19082 , \19077 , \19081 );
and \U$18871 ( \19083 , \19019 , \19023 );
and \U$18872 ( \19084 , \19023 , \19028 );
and \U$18873 ( \19085 , \19019 , \19028 );
or \U$18874 ( \19086 , \19083 , \19084 , \19085 );
and \U$18875 ( \19087 , \19033 , \19037 );
and \U$18876 ( \19088 , \19037 , \19039 );
and \U$18877 ( \19089 , \19033 , \19039 );
or \U$18878 ( \19090 , \19087 , \19088 , \19089 );
xor \U$18879 ( \19091 , \19086 , \19090 );
and \U$18880 ( \19092 , \18991 , \19005 );
and \U$18881 ( \19093 , \19005 , \19012 );
and \U$18882 ( \19094 , \18991 , \19012 );
or \U$18883 ( \19095 , \19092 , \19093 , \19094 );
xor \U$18884 ( \19096 , \19091 , \19095 );
and \U$18885 ( \19097 , \18949 , \18960 );
and \U$18886 ( \19098 , \18960 , \18975 );
and \U$18887 ( \19099 , \18949 , \18975 );
or \U$18888 ( \19100 , \19097 , \19098 , \19099 );
and \U$18889 ( \19101 , \8652 , \4581 );
and \U$18890 ( \19102 , \8835 , \4424 );
nor \U$18891 ( \19103 , \19101 , \19102 );
xnor \U$18892 ( \19104 , \19103 , \4377 );
and \U$18893 ( \19105 , \8057 , \5011 );
and \U$18894 ( \19106 , \8349 , \4878 );
nor \U$18895 ( \19107 , \19105 , \19106 );
xnor \U$18896 ( \19108 , \19107 , \4762 );
xor \U$18897 ( \19109 , \19104 , \19108 );
and \U$18898 ( \19110 , \7556 , \5485 );
and \U$18899 ( \19111 , \7700 , \5275 );
nor \U$18900 ( \19112 , \19110 , \19111 );
xnor \U$18901 ( \19113 , \19112 , \5169 );
xor \U$18902 ( \19114 , \19109 , \19113 );
and \U$18903 ( \19115 , \10584 , \3357 );
not \U$18904 ( \19116 , \19115 );
xnor \U$18905 ( \19117 , \19116 , \3156 );
and \U$18906 ( \19118 , \9897 , \3813 );
and \U$18907 ( \19119 , \10206 , \3557 );
nor \U$18908 ( \19120 , \19118 , \19119 );
xnor \U$18909 ( \19121 , \19120 , \3562 );
xor \U$18910 ( \19122 , \19117 , \19121 );
and \U$18911 ( \19123 , \9169 , \4132 );
and \U$18912 ( \19124 , \9465 , \4012 );
nor \U$18913 ( \19125 , \19123 , \19124 );
xnor \U$18914 ( \19126 , \19125 , \3925 );
xor \U$18915 ( \19127 , \19122 , \19126 );
xor \U$18916 ( \19128 , \19114 , \19127 );
and \U$18917 ( \19129 , \6945 , \5996 );
and \U$18918 ( \19130 , \7231 , \5695 );
nor \U$18919 ( \19131 , \19129 , \19130 );
xnor \U$18920 ( \19132 , \19131 , \5687 );
and \U$18921 ( \19133 , \6514 , \6401 );
and \U$18922 ( \19134 , \6790 , \6143 );
nor \U$18923 ( \19135 , \19133 , \19134 );
xnor \U$18924 ( \19136 , \19135 , \6148 );
xor \U$18925 ( \19137 , \19132 , \19136 );
and \U$18926 ( \19138 , \6030 , \7055 );
and \U$18927 ( \19139 , \6281 , \6675 );
nor \U$18928 ( \19140 , \19138 , \19139 );
xnor \U$18929 ( \19141 , \19140 , \6680 );
xor \U$18930 ( \19142 , \19137 , \19141 );
xor \U$18931 ( \19143 , \19128 , \19142 );
xor \U$18932 ( \19144 , \19100 , \19143 );
and \U$18933 ( \19145 , \4160 , \9333 );
and \U$18934 ( \19146 , \4364 , \9006 );
nor \U$18935 ( \19147 , \19145 , \19146 );
xnor \U$18936 ( \19148 , \19147 , \8848 );
and \U$18937 ( \19149 , \3736 , \9765 );
and \U$18938 ( \19150 , \3912 , \9644 );
nor \U$18939 ( \19151 , \19149 , \19150 );
xnor \U$18940 ( \19152 , \19151 , \9478 );
xor \U$18941 ( \19153 , \19148 , \19152 );
and \U$18942 ( \19154 , \3395 , \10408 );
and \U$18943 ( \19155 , \3646 , \10116 );
nor \U$18944 ( \19156 , \19154 , \19155 );
xnor \U$18945 ( \19157 , \19156 , \10121 );
xor \U$18946 ( \19158 , \19153 , \19157 );
and \U$18947 ( \19159 , \5469 , \7489 );
and \U$18948 ( \19160 , \5674 , \7137 );
nor \U$18949 ( \19161 , \19159 , \19160 );
xnor \U$18950 ( \19162 , \19161 , \7142 );
and \U$18951 ( \19163 , \4922 , \8019 );
and \U$18952 ( \19164 , \5156 , \7830 );
nor \U$18953 ( \19165 , \19163 , \19164 );
xnor \U$18954 ( \19166 , \19165 , \7713 );
xor \U$18955 ( \19167 , \19162 , \19166 );
and \U$18956 ( \19168 , \4654 , \8540 );
and \U$18957 ( \19169 , \4749 , \8292 );
nor \U$18958 ( \19170 , \19168 , \19169 );
xnor \U$18959 ( \19171 , \19170 , \8297 );
xor \U$18960 ( \19172 , \19167 , \19171 );
xor \U$18961 ( \19173 , \19158 , \19172 );
and \U$18962 ( \19174 , \3143 , \10118 );
not \U$18963 ( \19175 , \19174 );
xor \U$18964 ( \19176 , \19173 , \19175 );
xor \U$18965 ( \19177 , \19144 , \19176 );
xor \U$18966 ( \19178 , \19096 , \19177 );
and \U$18967 ( \19179 , \18939 , \18943 );
and \U$18968 ( \19180 , \18943 , \18948 );
and \U$18969 ( \19181 , \18939 , \18948 );
or \U$18970 ( \19182 , \19179 , \19180 , \19181 );
and \U$18971 ( \19183 , \18950 , \18954 );
and \U$18972 ( \19184 , \18954 , \18959 );
and \U$18973 ( \19185 , \18950 , \18959 );
or \U$18974 ( \19186 , \19183 , \19184 , \19185 );
xor \U$18975 ( \19187 , \19182 , \19186 );
and \U$18976 ( \19188 , \18965 , \18969 );
and \U$18977 ( \19189 , \18969 , \18974 );
and \U$18978 ( \19190 , \18965 , \18974 );
or \U$18979 ( \19191 , \19188 , \19189 , \19190 );
xor \U$18980 ( \19192 , \19187 , \19191 );
and \U$18981 ( \19193 , \18981 , \18985 );
and \U$18982 ( \19194 , \18985 , \18990 );
and \U$18983 ( \19195 , \18981 , \18990 );
or \U$18984 ( \19196 , \19193 , \19194 , \19195 );
and \U$18985 ( \19197 , \18995 , \18999 );
and \U$18986 ( \19198 , \18999 , \19004 );
and \U$18987 ( \19199 , \18995 , \19004 );
or \U$18988 ( \19200 , \19197 , \19198 , \19199 );
xor \U$18989 ( \19201 , \19196 , \19200 );
and \U$18990 ( \19202 , \19010 , \19011 );
xor \U$18991 ( \19203 , \19201 , \19202 );
xor \U$18992 ( \19204 , \19192 , \19203 );
xor \U$18993 ( \19205 , \19178 , \19204 );
xor \U$18994 ( \19206 , \19082 , \19205 );
xor \U$18995 ( \19207 , \19073 , \19206 );
xor \U$18996 ( \19208 , \19057 , \19207 );
and \U$18997 ( \19209 , \18892 , \19044 );
xor \U$18998 ( \19210 , \19208 , \19209 );
and \U$18999 ( \19211 , \19045 , \19046 );
and \U$19000 ( \19212 , \19047 , \19050 );
or \U$19001 ( \19213 , \19211 , \19212 );
xor \U$19002 ( \19214 , \19210 , \19213 );
buf g54d7_GF_PartitionCandidate( \19215_nG54d7 , \19214 );
buf \U$19003 ( \19216 , \19215_nG54d7 );
and \U$19004 ( \19217 , \19061 , \19072 );
and \U$19005 ( \19218 , \19072 , \19206 );
and \U$19006 ( \19219 , \19061 , \19206 );
or \U$19007 ( \19220 , \19217 , \19218 , \19219 );
and \U$19008 ( \19221 , \19077 , \19081 );
and \U$19009 ( \19222 , \19081 , \19205 );
and \U$19010 ( \19223 , \19077 , \19205 );
or \U$19011 ( \19224 , \19221 , \19222 , \19223 );
and \U$19012 ( \19225 , \19086 , \19090 );
and \U$19013 ( \19226 , \19090 , \19095 );
and \U$19014 ( \19227 , \19086 , \19095 );
or \U$19015 ( \19228 , \19225 , \19226 , \19227 );
and \U$19016 ( \19229 , \19100 , \19143 );
and \U$19017 ( \19230 , \19143 , \19176 );
and \U$19018 ( \19231 , \19100 , \19176 );
or \U$19019 ( \19232 , \19229 , \19230 , \19231 );
xor \U$19020 ( \19233 , \19228 , \19232 );
and \U$19021 ( \19234 , \19192 , \19203 );
xor \U$19022 ( \19235 , \19233 , \19234 );
xor \U$19023 ( \19236 , \19224 , \19235 );
and \U$19024 ( \19237 , \19065 , \19069 );
and \U$19025 ( \19238 , \19069 , \19071 );
and \U$19026 ( \19239 , \19065 , \19071 );
or \U$19027 ( \19240 , \19237 , \19238 , \19239 );
and \U$19028 ( \19241 , \19096 , \19177 );
and \U$19029 ( \19242 , \19177 , \19204 );
and \U$19030 ( \19243 , \19096 , \19204 );
or \U$19031 ( \19244 , \19241 , \19242 , \19243 );
xor \U$19032 ( \19245 , \19240 , \19244 );
and \U$19033 ( \19246 , \19182 , \19186 );
and \U$19034 ( \19247 , \19186 , \19191 );
and \U$19035 ( \19248 , \19182 , \19191 );
or \U$19036 ( \19249 , \19246 , \19247 , \19248 );
and \U$19037 ( \19250 , \19196 , \19200 );
and \U$19038 ( \19251 , \19200 , \19202 );
and \U$19039 ( \19252 , \19196 , \19202 );
or \U$19040 ( \19253 , \19250 , \19251 , \19252 );
xor \U$19041 ( \19254 , \19249 , \19253 );
and \U$19042 ( \19255 , \19158 , \19172 );
and \U$19043 ( \19256 , \19172 , \19175 );
and \U$19044 ( \19257 , \19158 , \19175 );
or \U$19045 ( \19258 , \19255 , \19256 , \19257 );
xor \U$19046 ( \19259 , \19254 , \19258 );
and \U$19047 ( \19260 , \19114 , \19127 );
and \U$19048 ( \19261 , \19127 , \19142 );
and \U$19049 ( \19262 , \19114 , \19142 );
or \U$19050 ( \19263 , \19260 , \19261 , \19262 );
and \U$19051 ( \19264 , \8835 , \4581 );
and \U$19052 ( \19265 , \9169 , \4424 );
nor \U$19053 ( \19266 , \19264 , \19265 );
xnor \U$19054 ( \19267 , \19266 , \4377 );
and \U$19055 ( \19268 , \8349 , \5011 );
and \U$19056 ( \19269 , \8652 , \4878 );
nor \U$19057 ( \19270 , \19268 , \19269 );
xnor \U$19058 ( \19271 , \19270 , \4762 );
xor \U$19059 ( \19272 , \19267 , \19271 );
and \U$19060 ( \19273 , \7700 , \5485 );
and \U$19061 ( \19274 , \8057 , \5275 );
nor \U$19062 ( \19275 , \19273 , \19274 );
xnor \U$19063 ( \19276 , \19275 , \5169 );
xor \U$19064 ( \19277 , \19272 , \19276 );
not \U$19065 ( \19278 , \3156 );
and \U$19066 ( \19279 , \10206 , \3813 );
and \U$19067 ( \19280 , \10584 , \3557 );
nor \U$19068 ( \19281 , \19279 , \19280 );
xnor \U$19069 ( \19282 , \19281 , \3562 );
xor \U$19070 ( \19283 , \19278 , \19282 );
and \U$19071 ( \19284 , \9465 , \4132 );
and \U$19072 ( \19285 , \9897 , \4012 );
nor \U$19073 ( \19286 , \19284 , \19285 );
xnor \U$19074 ( \19287 , \19286 , \3925 );
xor \U$19075 ( \19288 , \19283 , \19287 );
xor \U$19076 ( \19289 , \19277 , \19288 );
and \U$19077 ( \19290 , \7231 , \5996 );
and \U$19078 ( \19291 , \7556 , \5695 );
nor \U$19079 ( \19292 , \19290 , \19291 );
xnor \U$19080 ( \19293 , \19292 , \5687 );
and \U$19081 ( \19294 , \6790 , \6401 );
and \U$19082 ( \19295 , \6945 , \6143 );
nor \U$19083 ( \19296 , \19294 , \19295 );
xnor \U$19084 ( \19297 , \19296 , \6148 );
xor \U$19085 ( \19298 , \19293 , \19297 );
and \U$19086 ( \19299 , \6281 , \7055 );
and \U$19087 ( \19300 , \6514 , \6675 );
nor \U$19088 ( \19301 , \19299 , \19300 );
xnor \U$19089 ( \19302 , \19301 , \6680 );
xor \U$19090 ( \19303 , \19298 , \19302 );
xor \U$19091 ( \19304 , \19289 , \19303 );
xor \U$19092 ( \19305 , \19263 , \19304 );
and \U$19093 ( \19306 , \3395 , \10118 );
and \U$19094 ( \19307 , \4364 , \9333 );
and \U$19095 ( \19308 , \4654 , \9006 );
nor \U$19096 ( \19309 , \19307 , \19308 );
xnor \U$19097 ( \19310 , \19309 , \8848 );
and \U$19098 ( \19311 , \3912 , \9765 );
and \U$19099 ( \19312 , \4160 , \9644 );
nor \U$19100 ( \19313 , \19311 , \19312 );
xnor \U$19101 ( \19314 , \19313 , \9478 );
xor \U$19102 ( \19315 , \19310 , \19314 );
and \U$19103 ( \19316 , \3646 , \10408 );
and \U$19104 ( \19317 , \3736 , \10116 );
nor \U$19105 ( \19318 , \19316 , \19317 );
xnor \U$19106 ( \19319 , \19318 , \10121 );
xor \U$19107 ( \19320 , \19315 , \19319 );
xor \U$19108 ( \19321 , \19306 , \19320 );
and \U$19109 ( \19322 , \5674 , \7489 );
and \U$19110 ( \19323 , \6030 , \7137 );
nor \U$19111 ( \19324 , \19322 , \19323 );
xnor \U$19112 ( \19325 , \19324 , \7142 );
and \U$19113 ( \19326 , \5156 , \8019 );
and \U$19114 ( \19327 , \5469 , \7830 );
nor \U$19115 ( \19328 , \19326 , \19327 );
xnor \U$19116 ( \19329 , \19328 , \7713 );
xor \U$19117 ( \19330 , \19325 , \19329 );
and \U$19118 ( \19331 , \4749 , \8540 );
and \U$19119 ( \19332 , \4922 , \8292 );
nor \U$19120 ( \19333 , \19331 , \19332 );
xnor \U$19121 ( \19334 , \19333 , \8297 );
xor \U$19122 ( \19335 , \19330 , \19334 );
xor \U$19123 ( \19336 , \19321 , \19335 );
xor \U$19124 ( \19337 , \19305 , \19336 );
xor \U$19125 ( \19338 , \19259 , \19337 );
and \U$19126 ( \19339 , \19104 , \19108 );
and \U$19127 ( \19340 , \19108 , \19113 );
and \U$19128 ( \19341 , \19104 , \19113 );
or \U$19129 ( \19342 , \19339 , \19340 , \19341 );
and \U$19130 ( \19343 , \19117 , \19121 );
and \U$19131 ( \19344 , \19121 , \19126 );
and \U$19132 ( \19345 , \19117 , \19126 );
or \U$19133 ( \19346 , \19343 , \19344 , \19345 );
xor \U$19134 ( \19347 , \19342 , \19346 );
and \U$19135 ( \19348 , \19132 , \19136 );
and \U$19136 ( \19349 , \19136 , \19141 );
and \U$19137 ( \19350 , \19132 , \19141 );
or \U$19138 ( \19351 , \19348 , \19349 , \19350 );
xor \U$19139 ( \19352 , \19347 , \19351 );
and \U$19140 ( \19353 , \19148 , \19152 );
and \U$19141 ( \19354 , \19152 , \19157 );
and \U$19142 ( \19355 , \19148 , \19157 );
or \U$19143 ( \19356 , \19353 , \19354 , \19355 );
and \U$19144 ( \19357 , \19162 , \19166 );
and \U$19145 ( \19358 , \19166 , \19171 );
and \U$19146 ( \19359 , \19162 , \19171 );
or \U$19147 ( \19360 , \19357 , \19358 , \19359 );
xor \U$19148 ( \19361 , \19356 , \19360 );
buf \U$19149 ( \19362 , \19174 );
xor \U$19150 ( \19363 , \19361 , \19362 );
xor \U$19151 ( \19364 , \19352 , \19363 );
xor \U$19152 ( \19365 , \19338 , \19364 );
xor \U$19153 ( \19366 , \19245 , \19365 );
xor \U$19154 ( \19367 , \19236 , \19366 );
xor \U$19155 ( \19368 , \19220 , \19367 );
and \U$19156 ( \19369 , \19057 , \19207 );
xor \U$19157 ( \19370 , \19368 , \19369 );
and \U$19158 ( \19371 , \19208 , \19209 );
and \U$19159 ( \19372 , \19210 , \19213 );
or \U$19160 ( \19373 , \19371 , \19372 );
xor \U$19161 ( \19374 , \19370 , \19373 );
buf g54d5_GF_PartitionCandidate( \19375_nG54d5 , \19374 );
buf \U$19162 ( \19376 , \19375_nG54d5 );
and \U$19163 ( \19377 , \19224 , \19235 );
and \U$19164 ( \19378 , \19235 , \19366 );
and \U$19165 ( \19379 , \19224 , \19366 );
or \U$19166 ( \19380 , \19377 , \19378 , \19379 );
and \U$19167 ( \19381 , \19240 , \19244 );
and \U$19168 ( \19382 , \19244 , \19365 );
and \U$19169 ( \19383 , \19240 , \19365 );
or \U$19170 ( \19384 , \19381 , \19382 , \19383 );
and \U$19171 ( \19385 , \19249 , \19253 );
and \U$19172 ( \19386 , \19253 , \19258 );
and \U$19173 ( \19387 , \19249 , \19258 );
or \U$19174 ( \19388 , \19385 , \19386 , \19387 );
and \U$19175 ( \19389 , \19263 , \19304 );
and \U$19176 ( \19390 , \19304 , \19336 );
and \U$19177 ( \19391 , \19263 , \19336 );
or \U$19178 ( \19392 , \19389 , \19390 , \19391 );
xor \U$19179 ( \19393 , \19388 , \19392 );
and \U$19180 ( \19394 , \19352 , \19363 );
xor \U$19181 ( \19395 , \19393 , \19394 );
xor \U$19182 ( \19396 , \19384 , \19395 );
and \U$19183 ( \19397 , \19228 , \19232 );
and \U$19184 ( \19398 , \19232 , \19234 );
and \U$19185 ( \19399 , \19228 , \19234 );
or \U$19186 ( \19400 , \19397 , \19398 , \19399 );
and \U$19187 ( \19401 , \19259 , \19337 );
and \U$19188 ( \19402 , \19337 , \19364 );
and \U$19189 ( \19403 , \19259 , \19364 );
or \U$19190 ( \19404 , \19401 , \19402 , \19403 );
xor \U$19191 ( \19405 , \19400 , \19404 );
and \U$19192 ( \19406 , \19342 , \19346 );
and \U$19193 ( \19407 , \19346 , \19351 );
and \U$19194 ( \19408 , \19342 , \19351 );
or \U$19195 ( \19409 , \19406 , \19407 , \19408 );
and \U$19196 ( \19410 , \19356 , \19360 );
and \U$19197 ( \19411 , \19360 , \19362 );
and \U$19198 ( \19412 , \19356 , \19362 );
or \U$19199 ( \19413 , \19410 , \19411 , \19412 );
xor \U$19200 ( \19414 , \19409 , \19413 );
and \U$19201 ( \19415 , \19306 , \19320 );
and \U$19202 ( \19416 , \19320 , \19335 );
and \U$19203 ( \19417 , \19306 , \19335 );
or \U$19204 ( \19418 , \19415 , \19416 , \19417 );
xor \U$19205 ( \19419 , \19414 , \19418 );
and \U$19206 ( \19420 , \19277 , \19288 );
and \U$19207 ( \19421 , \19288 , \19303 );
and \U$19208 ( \19422 , \19277 , \19303 );
or \U$19209 ( \19423 , \19420 , \19421 , \19422 );
and \U$19210 ( \19424 , \10584 , \3813 );
not \U$19211 ( \19425 , \19424 );
xnor \U$19212 ( \19426 , \19425 , \3562 );
and \U$19213 ( \19427 , \9897 , \4132 );
and \U$19214 ( \19428 , \10206 , \4012 );
nor \U$19215 ( \19429 , \19427 , \19428 );
xnor \U$19216 ( \19430 , \19429 , \3925 );
xor \U$19217 ( \19431 , \19426 , \19430 );
and \U$19218 ( \19432 , \9169 , \4581 );
and \U$19219 ( \19433 , \9465 , \4424 );
nor \U$19220 ( \19434 , \19432 , \19433 );
xnor \U$19221 ( \19435 , \19434 , \4377 );
xor \U$19222 ( \19436 , \19431 , \19435 );
xor \U$19223 ( \19437 , \19423 , \19436 );
and \U$19224 ( \19438 , \8652 , \5011 );
and \U$19225 ( \19439 , \8835 , \4878 );
nor \U$19226 ( \19440 , \19438 , \19439 );
xnor \U$19227 ( \19441 , \19440 , \4762 );
and \U$19228 ( \19442 , \8057 , \5485 );
and \U$19229 ( \19443 , \8349 , \5275 );
nor \U$19230 ( \19444 , \19442 , \19443 );
xnor \U$19231 ( \19445 , \19444 , \5169 );
xor \U$19232 ( \19446 , \19441 , \19445 );
and \U$19233 ( \19447 , \7556 , \5996 );
and \U$19234 ( \19448 , \7700 , \5695 );
nor \U$19235 ( \19449 , \19447 , \19448 );
xnor \U$19236 ( \19450 , \19449 , \5687 );
xor \U$19237 ( \19451 , \19446 , \19450 );
xor \U$19238 ( \19452 , \19437 , \19451 );
xor \U$19239 ( \19453 , \19419 , \19452 );
and \U$19240 ( \19454 , \19267 , \19271 );
and \U$19241 ( \19455 , \19271 , \19276 );
and \U$19242 ( \19456 , \19267 , \19276 );
or \U$19243 ( \19457 , \19454 , \19455 , \19456 );
and \U$19244 ( \19458 , \19278 , \19282 );
and \U$19245 ( \19459 , \19282 , \19287 );
and \U$19246 ( \19460 , \19278 , \19287 );
or \U$19247 ( \19461 , \19458 , \19459 , \19460 );
xor \U$19248 ( \19462 , \19457 , \19461 );
and \U$19249 ( \19463 , \19293 , \19297 );
and \U$19250 ( \19464 , \19297 , \19302 );
and \U$19251 ( \19465 , \19293 , \19302 );
or \U$19252 ( \19466 , \19463 , \19464 , \19465 );
xor \U$19253 ( \19467 , \19462 , \19466 );
and \U$19254 ( \19468 , \5469 , \8019 );
and \U$19255 ( \19469 , \5674 , \7830 );
nor \U$19256 ( \19470 , \19468 , \19469 );
xnor \U$19257 ( \19471 , \19470 , \7713 );
and \U$19258 ( \19472 , \4922 , \8540 );
and \U$19259 ( \19473 , \5156 , \8292 );
nor \U$19260 ( \19474 , \19472 , \19473 );
xnor \U$19261 ( \19475 , \19474 , \8297 );
xor \U$19262 ( \19476 , \19471 , \19475 );
and \U$19263 ( \19477 , \4654 , \9333 );
and \U$19264 ( \19478 , \4749 , \9006 );
nor \U$19265 ( \19479 , \19477 , \19478 );
xnor \U$19266 ( \19480 , \19479 , \8848 );
xor \U$19267 ( \19481 , \19476 , \19480 );
and \U$19268 ( \19482 , \4160 , \9765 );
and \U$19269 ( \19483 , \4364 , \9644 );
nor \U$19270 ( \19484 , \19482 , \19483 );
xnor \U$19271 ( \19485 , \19484 , \9478 );
and \U$19272 ( \19486 , \3736 , \10408 );
and \U$19273 ( \19487 , \3912 , \10116 );
nor \U$19274 ( \19488 , \19486 , \19487 );
xnor \U$19275 ( \19489 , \19488 , \10121 );
xor \U$19276 ( \19490 , \19485 , \19489 );
and \U$19277 ( \19491 , \3646 , \10118 );
xor \U$19278 ( \19492 , \19490 , \19491 );
xor \U$19279 ( \19493 , \19481 , \19492 );
and \U$19280 ( \19494 , \6945 , \6401 );
and \U$19281 ( \19495 , \7231 , \6143 );
nor \U$19282 ( \19496 , \19494 , \19495 );
xnor \U$19283 ( \19497 , \19496 , \6148 );
and \U$19284 ( \19498 , \6514 , \7055 );
and \U$19285 ( \19499 , \6790 , \6675 );
nor \U$19286 ( \19500 , \19498 , \19499 );
xnor \U$19287 ( \19501 , \19500 , \6680 );
xor \U$19288 ( \19502 , \19497 , \19501 );
and \U$19289 ( \19503 , \6030 , \7489 );
and \U$19290 ( \19504 , \6281 , \7137 );
nor \U$19291 ( \19505 , \19503 , \19504 );
xnor \U$19292 ( \19506 , \19505 , \7142 );
xor \U$19293 ( \19507 , \19502 , \19506 );
xor \U$19294 ( \19508 , \19493 , \19507 );
xor \U$19295 ( \19509 , \19467 , \19508 );
and \U$19296 ( \19510 , \19310 , \19314 );
and \U$19297 ( \19511 , \19314 , \19319 );
and \U$19298 ( \19512 , \19310 , \19319 );
or \U$19299 ( \19513 , \19510 , \19511 , \19512 );
and \U$19300 ( \19514 , \19325 , \19329 );
and \U$19301 ( \19515 , \19329 , \19334 );
and \U$19302 ( \19516 , \19325 , \19334 );
or \U$19303 ( \19517 , \19514 , \19515 , \19516 );
xnor \U$19304 ( \19518 , \19513 , \19517 );
xor \U$19305 ( \19519 , \19509 , \19518 );
xor \U$19306 ( \19520 , \19453 , \19519 );
xor \U$19307 ( \19521 , \19405 , \19520 );
xor \U$19308 ( \19522 , \19396 , \19521 );
xor \U$19309 ( \19523 , \19380 , \19522 );
and \U$19310 ( \19524 , \19220 , \19367 );
xor \U$19311 ( \19525 , \19523 , \19524 );
and \U$19312 ( \19526 , \19368 , \19369 );
and \U$19313 ( \19527 , \19370 , \19373 );
or \U$19314 ( \19528 , \19526 , \19527 );
xor \U$19315 ( \19529 , \19525 , \19528 );
buf g54d3_GF_PartitionCandidate( \19530_nG54d3 , \19529 );
buf \U$19316 ( \19531 , \19530_nG54d3 );
and \U$19317 ( \19532 , \19384 , \19395 );
and \U$19318 ( \19533 , \19395 , \19521 );
and \U$19319 ( \19534 , \19384 , \19521 );
or \U$19320 ( \19535 , \19532 , \19533 , \19534 );
and \U$19321 ( \19536 , \19400 , \19404 );
and \U$19322 ( \19537 , \19404 , \19520 );
and \U$19323 ( \19538 , \19400 , \19520 );
or \U$19324 ( \19539 , \19536 , \19537 , \19538 );
and \U$19325 ( \19540 , \19409 , \19413 );
and \U$19326 ( \19541 , \19413 , \19418 );
and \U$19327 ( \19542 , \19409 , \19418 );
or \U$19328 ( \19543 , \19540 , \19541 , \19542 );
and \U$19329 ( \19544 , \19423 , \19436 );
and \U$19330 ( \19545 , \19436 , \19451 );
and \U$19331 ( \19546 , \19423 , \19451 );
or \U$19332 ( \19547 , \19544 , \19545 , \19546 );
xor \U$19333 ( \19548 , \19543 , \19547 );
and \U$19334 ( \19549 , \19467 , \19508 );
and \U$19335 ( \19550 , \19508 , \19518 );
and \U$19336 ( \19551 , \19467 , \19518 );
or \U$19337 ( \19552 , \19549 , \19550 , \19551 );
xor \U$19338 ( \19553 , \19548 , \19552 );
xor \U$19339 ( \19554 , \19539 , \19553 );
and \U$19340 ( \19555 , \19388 , \19392 );
and \U$19341 ( \19556 , \19392 , \19394 );
and \U$19342 ( \19557 , \19388 , \19394 );
or \U$19343 ( \19558 , \19555 , \19556 , \19557 );
and \U$19344 ( \19559 , \19419 , \19452 );
and \U$19345 ( \19560 , \19452 , \19519 );
and \U$19346 ( \19561 , \19419 , \19519 );
or \U$19347 ( \19562 , \19559 , \19560 , \19561 );
xor \U$19348 ( \19563 , \19558 , \19562 );
and \U$19349 ( \19564 , \19426 , \19430 );
and \U$19350 ( \19565 , \19430 , \19435 );
and \U$19351 ( \19566 , \19426 , \19435 );
or \U$19352 ( \19567 , \19564 , \19565 , \19566 );
and \U$19353 ( \19568 , \19441 , \19445 );
and \U$19354 ( \19569 , \19445 , \19450 );
and \U$19355 ( \19570 , \19441 , \19450 );
or \U$19356 ( \19571 , \19568 , \19569 , \19570 );
xor \U$19357 ( \19572 , \19567 , \19571 );
and \U$19358 ( \19573 , \19497 , \19501 );
and \U$19359 ( \19574 , \19501 , \19506 );
and \U$19360 ( \19575 , \19497 , \19506 );
or \U$19361 ( \19576 , \19573 , \19574 , \19575 );
xor \U$19362 ( \19577 , \19572 , \19576 );
and \U$19363 ( \19578 , \19457 , \19461 );
and \U$19364 ( \19579 , \19461 , \19466 );
and \U$19365 ( \19580 , \19457 , \19466 );
or \U$19366 ( \19581 , \19578 , \19579 , \19580 );
and \U$19367 ( \19582 , \19481 , \19492 );
and \U$19368 ( \19583 , \19492 , \19507 );
and \U$19369 ( \19584 , \19481 , \19507 );
or \U$19370 ( \19585 , \19582 , \19583 , \19584 );
xor \U$19371 ( \19586 , \19581 , \19585 );
or \U$19372 ( \19587 , \19513 , \19517 );
xor \U$19373 ( \19588 , \19586 , \19587 );
xor \U$19374 ( \19589 , \19577 , \19588 );
not \U$19375 ( \19590 , \3562 );
and \U$19376 ( \19591 , \10206 , \4132 );
and \U$19377 ( \19592 , \10584 , \4012 );
nor \U$19378 ( \19593 , \19591 , \19592 );
xnor \U$19379 ( \19594 , \19593 , \3925 );
xor \U$19380 ( \19595 , \19590 , \19594 );
and \U$19381 ( \19596 , \9465 , \4581 );
and \U$19382 ( \19597 , \9897 , \4424 );
nor \U$19383 ( \19598 , \19596 , \19597 );
xnor \U$19384 ( \19599 , \19598 , \4377 );
xor \U$19385 ( \19600 , \19595 , \19599 );
and \U$19386 ( \19601 , \19471 , \19475 );
and \U$19387 ( \19602 , \19475 , \19480 );
and \U$19388 ( \19603 , \19471 , \19480 );
or \U$19389 ( \19604 , \19601 , \19602 , \19603 );
and \U$19390 ( \19605 , \19485 , \19489 );
and \U$19391 ( \19606 , \19489 , \19491 );
and \U$19392 ( \19607 , \19485 , \19491 );
or \U$19393 ( \19608 , \19605 , \19606 , \19607 );
xor \U$19394 ( \19609 , \19604 , \19608 );
and \U$19395 ( \19610 , \4364 , \9765 );
and \U$19396 ( \19611 , \4654 , \9644 );
nor \U$19397 ( \19612 , \19610 , \19611 );
xnor \U$19398 ( \19613 , \19612 , \9478 );
and \U$19399 ( \19614 , \3912 , \10408 );
and \U$19400 ( \19615 , \4160 , \10116 );
nor \U$19401 ( \19616 , \19614 , \19615 );
xnor \U$19402 ( \19617 , \19616 , \10121 );
xor \U$19403 ( \19618 , \19613 , \19617 );
and \U$19404 ( \19619 , \3736 , \10118 );
xor \U$19405 ( \19620 , \19618 , \19619 );
xor \U$19406 ( \19621 , \19609 , \19620 );
xor \U$19407 ( \19622 , \19600 , \19621 );
and \U$19408 ( \19623 , \8835 , \5011 );
and \U$19409 ( \19624 , \9169 , \4878 );
nor \U$19410 ( \19625 , \19623 , \19624 );
xnor \U$19411 ( \19626 , \19625 , \4762 );
and \U$19412 ( \19627 , \8349 , \5485 );
and \U$19413 ( \19628 , \8652 , \5275 );
nor \U$19414 ( \19629 , \19627 , \19628 );
xnor \U$19415 ( \19630 , \19629 , \5169 );
xor \U$19416 ( \19631 , \19626 , \19630 );
and \U$19417 ( \19632 , \7700 , \5996 );
and \U$19418 ( \19633 , \8057 , \5695 );
nor \U$19419 ( \19634 , \19632 , \19633 );
xnor \U$19420 ( \19635 , \19634 , \5687 );
xor \U$19421 ( \19636 , \19631 , \19635 );
and \U$19422 ( \19637 , \5674 , \8019 );
and \U$19423 ( \19638 , \6030 , \7830 );
nor \U$19424 ( \19639 , \19637 , \19638 );
xnor \U$19425 ( \19640 , \19639 , \7713 );
and \U$19426 ( \19641 , \5156 , \8540 );
and \U$19427 ( \19642 , \5469 , \8292 );
nor \U$19428 ( \19643 , \19641 , \19642 );
xnor \U$19429 ( \19644 , \19643 , \8297 );
xor \U$19430 ( \19645 , \19640 , \19644 );
and \U$19431 ( \19646 , \4749 , \9333 );
and \U$19432 ( \19647 , \4922 , \9006 );
nor \U$19433 ( \19648 , \19646 , \19647 );
xnor \U$19434 ( \19649 , \19648 , \8848 );
xor \U$19435 ( \19650 , \19645 , \19649 );
xor \U$19436 ( \19651 , \19636 , \19650 );
and \U$19437 ( \19652 , \7231 , \6401 );
and \U$19438 ( \19653 , \7556 , \6143 );
nor \U$19439 ( \19654 , \19652 , \19653 );
xnor \U$19440 ( \19655 , \19654 , \6148 );
and \U$19441 ( \19656 , \6790 , \7055 );
and \U$19442 ( \19657 , \6945 , \6675 );
nor \U$19443 ( \19658 , \19656 , \19657 );
xnor \U$19444 ( \19659 , \19658 , \6680 );
xor \U$19445 ( \19660 , \19655 , \19659 );
and \U$19446 ( \19661 , \6281 , \7489 );
and \U$19447 ( \19662 , \6514 , \7137 );
nor \U$19448 ( \19663 , \19661 , \19662 );
xnor \U$19449 ( \19664 , \19663 , \7142 );
xor \U$19450 ( \19665 , \19660 , \19664 );
xor \U$19451 ( \19666 , \19651 , \19665 );
xor \U$19452 ( \19667 , \19622 , \19666 );
xor \U$19453 ( \19668 , \19589 , \19667 );
xor \U$19454 ( \19669 , \19563 , \19668 );
xor \U$19455 ( \19670 , \19554 , \19669 );
xor \U$19456 ( \19671 , \19535 , \19670 );
and \U$19457 ( \19672 , \19380 , \19522 );
xor \U$19458 ( \19673 , \19671 , \19672 );
and \U$19459 ( \19674 , \19523 , \19524 );
and \U$19460 ( \19675 , \19525 , \19528 );
or \U$19461 ( \19676 , \19674 , \19675 );
xor \U$19462 ( \19677 , \19673 , \19676 );
buf g54d1_GF_PartitionCandidate( \19678_nG54d1 , \19677 );
buf \U$19463 ( \19679 , \19678_nG54d1 );
and \U$19464 ( \19680 , \19539 , \19553 );
and \U$19465 ( \19681 , \19553 , \19669 );
and \U$19466 ( \19682 , \19539 , \19669 );
or \U$19467 ( \19683 , \19680 , \19681 , \19682 );
and \U$19468 ( \19684 , \19558 , \19562 );
and \U$19469 ( \19685 , \19562 , \19668 );
and \U$19470 ( \19686 , \19558 , \19668 );
or \U$19471 ( \19687 , \19684 , \19685 , \19686 );
and \U$19472 ( \19688 , \19543 , \19547 );
and \U$19473 ( \19689 , \19547 , \19552 );
and \U$19474 ( \19690 , \19543 , \19552 );
or \U$19475 ( \19691 , \19688 , \19689 , \19690 );
and \U$19476 ( \19692 , \19577 , \19588 );
and \U$19477 ( \19693 , \19588 , \19667 );
and \U$19478 ( \19694 , \19577 , \19667 );
or \U$19479 ( \19695 , \19692 , \19693 , \19694 );
xor \U$19480 ( \19696 , \19691 , \19695 );
and \U$19481 ( \19697 , \10584 , \4132 );
not \U$19482 ( \19698 , \19697 );
xnor \U$19483 ( \19699 , \19698 , \3925 );
and \U$19484 ( \19700 , \9897 , \4581 );
and \U$19485 ( \19701 , \10206 , \4424 );
nor \U$19486 ( \19702 , \19700 , \19701 );
xnor \U$19487 ( \19703 , \19702 , \4377 );
xor \U$19488 ( \19704 , \19699 , \19703 );
and \U$19489 ( \19705 , \9169 , \5011 );
and \U$19490 ( \19706 , \9465 , \4878 );
nor \U$19491 ( \19707 , \19705 , \19706 );
xnor \U$19492 ( \19708 , \19707 , \4762 );
xor \U$19493 ( \19709 , \19704 , \19708 );
and \U$19494 ( \19710 , \6945 , \7055 );
and \U$19495 ( \19711 , \7231 , \6675 );
nor \U$19496 ( \19712 , \19710 , \19711 );
xnor \U$19497 ( \19713 , \19712 , \6680 );
and \U$19498 ( \19714 , \6514 , \7489 );
and \U$19499 ( \19715 , \6790 , \7137 );
nor \U$19500 ( \19716 , \19714 , \19715 );
xnor \U$19501 ( \19717 , \19716 , \7142 );
xor \U$19502 ( \19718 , \19713 , \19717 );
and \U$19503 ( \19719 , \6030 , \8019 );
and \U$19504 ( \19720 , \6281 , \7830 );
nor \U$19505 ( \19721 , \19719 , \19720 );
xnor \U$19506 ( \19722 , \19721 , \7713 );
xor \U$19507 ( \19723 , \19718 , \19722 );
and \U$19508 ( \19724 , \8652 , \5485 );
and \U$19509 ( \19725 , \8835 , \5275 );
nor \U$19510 ( \19726 , \19724 , \19725 );
xnor \U$19511 ( \19727 , \19726 , \5169 );
and \U$19512 ( \19728 , \8057 , \5996 );
and \U$19513 ( \19729 , \8349 , \5695 );
nor \U$19514 ( \19730 , \19728 , \19729 );
xnor \U$19515 ( \19731 , \19730 , \5687 );
xor \U$19516 ( \19732 , \19727 , \19731 );
and \U$19517 ( \19733 , \7556 , \6401 );
and \U$19518 ( \19734 , \7700 , \6143 );
nor \U$19519 ( \19735 , \19733 , \19734 );
xnor \U$19520 ( \19736 , \19735 , \6148 );
xor \U$19521 ( \19737 , \19732 , \19736 );
xor \U$19522 ( \19738 , \19723 , \19737 );
and \U$19523 ( \19739 , \5469 , \8540 );
and \U$19524 ( \19740 , \5674 , \8292 );
nor \U$19525 ( \19741 , \19739 , \19740 );
xnor \U$19526 ( \19742 , \19741 , \8297 );
and \U$19527 ( \19743 , \4922 , \9333 );
and \U$19528 ( \19744 , \5156 , \9006 );
nor \U$19529 ( \19745 , \19743 , \19744 );
xnor \U$19530 ( \19746 , \19745 , \8848 );
xor \U$19531 ( \19747 , \19742 , \19746 );
and \U$19532 ( \19748 , \4654 , \9765 );
and \U$19533 ( \19749 , \4749 , \9644 );
nor \U$19534 ( \19750 , \19748 , \19749 );
xnor \U$19535 ( \19751 , \19750 , \9478 );
xor \U$19536 ( \19752 , \19747 , \19751 );
xor \U$19537 ( \19753 , \19738 , \19752 );
xor \U$19538 ( \19754 , \19709 , \19753 );
and \U$19539 ( \19755 , \19613 , \19617 );
and \U$19540 ( \19756 , \19617 , \19619 );
and \U$19541 ( \19757 , \19613 , \19619 );
or \U$19542 ( \19758 , \19755 , \19756 , \19757 );
and \U$19543 ( \19759 , \19640 , \19644 );
and \U$19544 ( \19760 , \19644 , \19649 );
and \U$19545 ( \19761 , \19640 , \19649 );
or \U$19546 ( \19762 , \19759 , \19760 , \19761 );
xor \U$19547 ( \19763 , \19758 , \19762 );
and \U$19548 ( \19764 , \4160 , \10408 );
and \U$19549 ( \19765 , \4364 , \10116 );
nor \U$19550 ( \19766 , \19764 , \19765 );
xnor \U$19551 ( \19767 , \19766 , \10121 );
and \U$19552 ( \19768 , \3912 , \10118 );
xnor \U$19553 ( \19769 , \19767 , \19768 );
xor \U$19554 ( \19770 , \19763 , \19769 );
xor \U$19555 ( \19771 , \19754 , \19770 );
xor \U$19556 ( \19772 , \19696 , \19771 );
xor \U$19557 ( \19773 , \19687 , \19772 );
and \U$19558 ( \19774 , \19567 , \19571 );
and \U$19559 ( \19775 , \19571 , \19576 );
and \U$19560 ( \19776 , \19567 , \19576 );
or \U$19561 ( \19777 , \19774 , \19775 , \19776 );
and \U$19562 ( \19778 , \19604 , \19608 );
and \U$19563 ( \19779 , \19608 , \19620 );
and \U$19564 ( \19780 , \19604 , \19620 );
or \U$19565 ( \19781 , \19778 , \19779 , \19780 );
xor \U$19566 ( \19782 , \19777 , \19781 );
and \U$19567 ( \19783 , \19636 , \19650 );
and \U$19568 ( \19784 , \19650 , \19665 );
and \U$19569 ( \19785 , \19636 , \19665 );
or \U$19570 ( \19786 , \19783 , \19784 , \19785 );
xor \U$19571 ( \19787 , \19782 , \19786 );
and \U$19572 ( \19788 , \19581 , \19585 );
and \U$19573 ( \19789 , \19585 , \19587 );
and \U$19574 ( \19790 , \19581 , \19587 );
or \U$19575 ( \19791 , \19788 , \19789 , \19790 );
and \U$19576 ( \19792 , \19600 , \19621 );
and \U$19577 ( \19793 , \19621 , \19666 );
and \U$19578 ( \19794 , \19600 , \19666 );
or \U$19579 ( \19795 , \19792 , \19793 , \19794 );
xor \U$19580 ( \19796 , \19791 , \19795 );
and \U$19581 ( \19797 , \19590 , \19594 );
and \U$19582 ( \19798 , \19594 , \19599 );
and \U$19583 ( \19799 , \19590 , \19599 );
or \U$19584 ( \19800 , \19797 , \19798 , \19799 );
and \U$19585 ( \19801 , \19626 , \19630 );
and \U$19586 ( \19802 , \19630 , \19635 );
and \U$19587 ( \19803 , \19626 , \19635 );
or \U$19588 ( \19804 , \19801 , \19802 , \19803 );
xor \U$19589 ( \19805 , \19800 , \19804 );
and \U$19590 ( \19806 , \19655 , \19659 );
and \U$19591 ( \19807 , \19659 , \19664 );
and \U$19592 ( \19808 , \19655 , \19664 );
or \U$19593 ( \19809 , \19806 , \19807 , \19808 );
xor \U$19594 ( \19810 , \19805 , \19809 );
xor \U$19595 ( \19811 , \19796 , \19810 );
xor \U$19596 ( \19812 , \19787 , \19811 );
xor \U$19597 ( \19813 , \19773 , \19812 );
xor \U$19598 ( \19814 , \19683 , \19813 );
and \U$19599 ( \19815 , \19535 , \19670 );
xor \U$19600 ( \19816 , \19814 , \19815 );
and \U$19601 ( \19817 , \19671 , \19672 );
and \U$19602 ( \19818 , \19673 , \19676 );
or \U$19603 ( \19819 , \19817 , \19818 );
xor \U$19604 ( \19820 , \19816 , \19819 );
buf g54cf_GF_PartitionCandidate( \19821_nG54cf , \19820 );
buf \U$19605 ( \19822 , \19821_nG54cf );
and \U$19606 ( \19823 , \19687 , \19772 );
and \U$19607 ( \19824 , \19772 , \19812 );
and \U$19608 ( \19825 , \19687 , \19812 );
or \U$19609 ( \19826 , \19823 , \19824 , \19825 );
and \U$19610 ( \19827 , \19691 , \19695 );
and \U$19611 ( \19828 , \19695 , \19771 );
and \U$19612 ( \19829 , \19691 , \19771 );
or \U$19613 ( \19830 , \19827 , \19828 , \19829 );
and \U$19614 ( \19831 , \19787 , \19811 );
xor \U$19615 ( \19832 , \19830 , \19831 );
and \U$19616 ( \19833 , \19791 , \19795 );
and \U$19617 ( \19834 , \19795 , \19810 );
and \U$19618 ( \19835 , \19791 , \19810 );
or \U$19619 ( \19836 , \19833 , \19834 , \19835 );
and \U$19620 ( \19837 , \19777 , \19781 );
and \U$19621 ( \19838 , \19781 , \19786 );
and \U$19622 ( \19839 , \19777 , \19786 );
or \U$19623 ( \19840 , \19837 , \19838 , \19839 );
and \U$19624 ( \19841 , \19709 , \19753 );
and \U$19625 ( \19842 , \19753 , \19770 );
and \U$19626 ( \19843 , \19709 , \19770 );
or \U$19627 ( \19844 , \19841 , \19842 , \19843 );
xor \U$19628 ( \19845 , \19840 , \19844 );
and \U$19629 ( \19846 , \19742 , \19746 );
and \U$19630 ( \19847 , \19746 , \19751 );
and \U$19631 ( \19848 , \19742 , \19751 );
or \U$19632 ( \19849 , \19846 , \19847 , \19848 );
or \U$19633 ( \19850 , \19767 , \19768 );
xor \U$19634 ( \19851 , \19849 , \19850 );
and \U$19635 ( \19852 , \4364 , \10408 );
and \U$19636 ( \19853 , \4654 , \10116 );
nor \U$19637 ( \19854 , \19852 , \19853 );
xnor \U$19638 ( \19855 , \19854 , \10121 );
xor \U$19639 ( \19856 , \19851 , \19855 );
xor \U$19640 ( \19857 , \19845 , \19856 );
xor \U$19641 ( \19858 , \19836 , \19857 );
and \U$19642 ( \19859 , \19713 , \19717 );
and \U$19643 ( \19860 , \19717 , \19722 );
and \U$19644 ( \19861 , \19713 , \19722 );
or \U$19645 ( \19862 , \19859 , \19860 , \19861 );
and \U$19646 ( \19863 , \19727 , \19731 );
and \U$19647 ( \19864 , \19731 , \19736 );
and \U$19648 ( \19865 , \19727 , \19736 );
or \U$19649 ( \19866 , \19863 , \19864 , \19865 );
xor \U$19650 ( \19867 , \19862 , \19866 );
and \U$19651 ( \19868 , \19699 , \19703 );
and \U$19652 ( \19869 , \19703 , \19708 );
and \U$19653 ( \19870 , \19699 , \19708 );
or \U$19654 ( \19871 , \19868 , \19869 , \19870 );
xor \U$19655 ( \19872 , \19867 , \19871 );
and \U$19656 ( \19873 , \19800 , \19804 );
and \U$19657 ( \19874 , \19804 , \19809 );
and \U$19658 ( \19875 , \19800 , \19809 );
or \U$19659 ( \19876 , \19873 , \19874 , \19875 );
and \U$19660 ( \19877 , \19723 , \19737 );
and \U$19661 ( \19878 , \19737 , \19752 );
and \U$19662 ( \19879 , \19723 , \19752 );
or \U$19663 ( \19880 , \19877 , \19878 , \19879 );
xor \U$19664 ( \19881 , \19876 , \19880 );
and \U$19665 ( \19882 , \19758 , \19762 );
and \U$19666 ( \19883 , \19762 , \19769 );
and \U$19667 ( \19884 , \19758 , \19769 );
or \U$19668 ( \19885 , \19882 , \19883 , \19884 );
xor \U$19669 ( \19886 , \19881 , \19885 );
xor \U$19670 ( \19887 , \19872 , \19886 );
and \U$19671 ( \19888 , \8835 , \5485 );
and \U$19672 ( \19889 , \9169 , \5275 );
nor \U$19673 ( \19890 , \19888 , \19889 );
xnor \U$19674 ( \19891 , \19890 , \5169 );
and \U$19675 ( \19892 , \8349 , \5996 );
and \U$19676 ( \19893 , \8652 , \5695 );
nor \U$19677 ( \19894 , \19892 , \19893 );
xnor \U$19678 ( \19895 , \19894 , \5687 );
xor \U$19679 ( \19896 , \19891 , \19895 );
and \U$19680 ( \19897 , \7700 , \6401 );
and \U$19681 ( \19898 , \8057 , \6143 );
nor \U$19682 ( \19899 , \19897 , \19898 );
xnor \U$19683 ( \19900 , \19899 , \6148 );
xor \U$19684 ( \19901 , \19896 , \19900 );
not \U$19685 ( \19902 , \3925 );
and \U$19686 ( \19903 , \10206 , \4581 );
and \U$19687 ( \19904 , \10584 , \4424 );
nor \U$19688 ( \19905 , \19903 , \19904 );
xnor \U$19689 ( \19906 , \19905 , \4377 );
xor \U$19690 ( \19907 , \19902 , \19906 );
and \U$19691 ( \19908 , \9465 , \5011 );
and \U$19692 ( \19909 , \9897 , \4878 );
nor \U$19693 ( \19910 , \19908 , \19909 );
xnor \U$19694 ( \19911 , \19910 , \4762 );
xor \U$19695 ( \19912 , \19907 , \19911 );
xor \U$19696 ( \19913 , \19901 , \19912 );
and \U$19697 ( \19914 , \4160 , \10118 );
and \U$19698 ( \19915 , \7231 , \7055 );
and \U$19699 ( \19916 , \7556 , \6675 );
nor \U$19700 ( \19917 , \19915 , \19916 );
xnor \U$19701 ( \19918 , \19917 , \6680 );
and \U$19702 ( \19919 , \6790 , \7489 );
and \U$19703 ( \19920 , \6945 , \7137 );
nor \U$19704 ( \19921 , \19919 , \19920 );
xnor \U$19705 ( \19922 , \19921 , \7142 );
xor \U$19706 ( \19923 , \19918 , \19922 );
and \U$19707 ( \19924 , \6281 , \8019 );
and \U$19708 ( \19925 , \6514 , \7830 );
nor \U$19709 ( \19926 , \19924 , \19925 );
xnor \U$19710 ( \19927 , \19926 , \7713 );
xor \U$19711 ( \19928 , \19923 , \19927 );
xor \U$19712 ( \19929 , \19914 , \19928 );
and \U$19713 ( \19930 , \5674 , \8540 );
and \U$19714 ( \19931 , \6030 , \8292 );
nor \U$19715 ( \19932 , \19930 , \19931 );
xnor \U$19716 ( \19933 , \19932 , \8297 );
and \U$19717 ( \19934 , \5156 , \9333 );
and \U$19718 ( \19935 , \5469 , \9006 );
nor \U$19719 ( \19936 , \19934 , \19935 );
xnor \U$19720 ( \19937 , \19936 , \8848 );
xor \U$19721 ( \19938 , \19933 , \19937 );
and \U$19722 ( \19939 , \4749 , \9765 );
and \U$19723 ( \19940 , \4922 , \9644 );
nor \U$19724 ( \19941 , \19939 , \19940 );
xnor \U$19725 ( \19942 , \19941 , \9478 );
xor \U$19726 ( \19943 , \19938 , \19942 );
xor \U$19727 ( \19944 , \19929 , \19943 );
xor \U$19728 ( \19945 , \19913 , \19944 );
xor \U$19729 ( \19946 , \19887 , \19945 );
xor \U$19730 ( \19947 , \19858 , \19946 );
xor \U$19731 ( \19948 , \19832 , \19947 );
xor \U$19732 ( \19949 , \19826 , \19948 );
and \U$19733 ( \19950 , \19683 , \19813 );
xor \U$19734 ( \19951 , \19949 , \19950 );
and \U$19735 ( \19952 , \19814 , \19815 );
and \U$19736 ( \19953 , \19816 , \19819 );
or \U$19737 ( \19954 , \19952 , \19953 );
xor \U$19738 ( \19955 , \19951 , \19954 );
buf g54cd_GF_PartitionCandidate( \19956_nG54cd , \19955 );
buf \U$19739 ( \19957 , \19956_nG54cd );
and \U$19740 ( \19958 , \19830 , \19831 );
and \U$19741 ( \19959 , \19831 , \19947 );
and \U$19742 ( \19960 , \19830 , \19947 );
or \U$19743 ( \19961 , \19958 , \19959 , \19960 );
and \U$19744 ( \19962 , \19836 , \19857 );
and \U$19745 ( \19963 , \19857 , \19946 );
and \U$19746 ( \19964 , \19836 , \19946 );
or \U$19747 ( \19965 , \19962 , \19963 , \19964 );
and \U$19748 ( \19966 , \19840 , \19844 );
and \U$19749 ( \19967 , \19844 , \19856 );
and \U$19750 ( \19968 , \19840 , \19856 );
or \U$19751 ( \19969 , \19966 , \19967 , \19968 );
and \U$19752 ( \19970 , \19872 , \19886 );
and \U$19753 ( \19971 , \19886 , \19945 );
and \U$19754 ( \19972 , \19872 , \19945 );
or \U$19755 ( \19973 , \19970 , \19971 , \19972 );
xor \U$19756 ( \19974 , \19969 , \19973 );
and \U$19757 ( \19975 , \19849 , \19850 );
and \U$19758 ( \19976 , \19850 , \19855 );
and \U$19759 ( \19977 , \19849 , \19855 );
or \U$19760 ( \19978 , \19975 , \19976 , \19977 );
and \U$19761 ( \19979 , \19862 , \19866 );
and \U$19762 ( \19980 , \19866 , \19871 );
and \U$19763 ( \19981 , \19862 , \19871 );
or \U$19764 ( \19982 , \19979 , \19980 , \19981 );
xor \U$19765 ( \19983 , \19978 , \19982 );
and \U$19766 ( \19984 , \19914 , \19928 );
and \U$19767 ( \19985 , \19928 , \19943 );
and \U$19768 ( \19986 , \19914 , \19943 );
or \U$19769 ( \19987 , \19984 , \19985 , \19986 );
xor \U$19770 ( \19988 , \19983 , \19987 );
xor \U$19771 ( \19989 , \19974 , \19988 );
xor \U$19772 ( \19990 , \19965 , \19989 );
and \U$19773 ( \19991 , \19876 , \19880 );
and \U$19774 ( \19992 , \19880 , \19885 );
and \U$19775 ( \19993 , \19876 , \19885 );
or \U$19776 ( \19994 , \19991 , \19992 , \19993 );
and \U$19777 ( \19995 , \19901 , \19912 );
and \U$19778 ( \19996 , \19912 , \19944 );
and \U$19779 ( \19997 , \19901 , \19944 );
or \U$19780 ( \19998 , \19995 , \19996 , \19997 );
xor \U$19781 ( \19999 , \19994 , \19998 );
and \U$19782 ( \20000 , \19918 , \19922 );
and \U$19783 ( \20001 , \19922 , \19927 );
and \U$19784 ( \20002 , \19918 , \19927 );
or \U$19785 ( \20003 , \20000 , \20001 , \20002 );
and \U$19786 ( \20004 , \19891 , \19895 );
and \U$19787 ( \20005 , \19895 , \19900 );
and \U$19788 ( \20006 , \19891 , \19900 );
or \U$19789 ( \20007 , \20004 , \20005 , \20006 );
xor \U$19790 ( \20008 , \20003 , \20007 );
and \U$19791 ( \20009 , \19902 , \19906 );
and \U$19792 ( \20010 , \19906 , \19911 );
and \U$19793 ( \20011 , \19902 , \19911 );
or \U$19794 ( \20012 , \20009 , \20010 , \20011 );
xor \U$19795 ( \20013 , \20008 , \20012 );
and \U$19796 ( \20014 , \8652 , \5996 );
and \U$19797 ( \20015 , \8835 , \5695 );
nor \U$19798 ( \20016 , \20014 , \20015 );
xnor \U$19799 ( \20017 , \20016 , \5687 );
and \U$19800 ( \20018 , \8057 , \6401 );
and \U$19801 ( \20019 , \8349 , \6143 );
nor \U$19802 ( \20020 , \20018 , \20019 );
xnor \U$19803 ( \20021 , \20020 , \6148 );
xor \U$19804 ( \20022 , \20017 , \20021 );
and \U$19805 ( \20023 , \7556 , \7055 );
and \U$19806 ( \20024 , \7700 , \6675 );
nor \U$19807 ( \20025 , \20023 , \20024 );
xnor \U$19808 ( \20026 , \20025 , \6680 );
xor \U$19809 ( \20027 , \20022 , \20026 );
and \U$19810 ( \20028 , \10584 , \4581 );
not \U$19811 ( \20029 , \20028 );
xnor \U$19812 ( \20030 , \20029 , \4377 );
and \U$19813 ( \20031 , \9897 , \5011 );
and \U$19814 ( \20032 , \10206 , \4878 );
nor \U$19815 ( \20033 , \20031 , \20032 );
xnor \U$19816 ( \20034 , \20033 , \4762 );
xor \U$19817 ( \20035 , \20030 , \20034 );
and \U$19818 ( \20036 , \9169 , \5485 );
and \U$19819 ( \20037 , \9465 , \5275 );
nor \U$19820 ( \20038 , \20036 , \20037 );
xnor \U$19821 ( \20039 , \20038 , \5169 );
xor \U$19822 ( \20040 , \20035 , \20039 );
xor \U$19823 ( \20041 , \20027 , \20040 );
and \U$19824 ( \20042 , \6945 , \7489 );
and \U$19825 ( \20043 , \7231 , \7137 );
nor \U$19826 ( \20044 , \20042 , \20043 );
xnor \U$19827 ( \20045 , \20044 , \7142 );
and \U$19828 ( \20046 , \6514 , \8019 );
and \U$19829 ( \20047 , \6790 , \7830 );
nor \U$19830 ( \20048 , \20046 , \20047 );
xnor \U$19831 ( \20049 , \20048 , \7713 );
xor \U$19832 ( \20050 , \20045 , \20049 );
and \U$19833 ( \20051 , \6030 , \8540 );
and \U$19834 ( \20052 , \6281 , \8292 );
nor \U$19835 ( \20053 , \20051 , \20052 );
xnor \U$19836 ( \20054 , \20053 , \8297 );
xor \U$19837 ( \20055 , \20050 , \20054 );
xor \U$19838 ( \20056 , \20041 , \20055 );
xor \U$19839 ( \20057 , \20013 , \20056 );
and \U$19840 ( \20058 , \19933 , \19937 );
and \U$19841 ( \20059 , \19937 , \19942 );
and \U$19842 ( \20060 , \19933 , \19942 );
or \U$19843 ( \20061 , \20058 , \20059 , \20060 );
and \U$19844 ( \20062 , \5469 , \9333 );
and \U$19845 ( \20063 , \5674 , \9006 );
nor \U$19846 ( \20064 , \20062 , \20063 );
xnor \U$19847 ( \20065 , \20064 , \8848 );
and \U$19848 ( \20066 , \4922 , \9765 );
and \U$19849 ( \20067 , \5156 , \9644 );
nor \U$19850 ( \20068 , \20066 , \20067 );
xnor \U$19851 ( \20069 , \20068 , \9478 );
xor \U$19852 ( \20070 , \20065 , \20069 );
and \U$19853 ( \20071 , \4654 , \10408 );
and \U$19854 ( \20072 , \4749 , \10116 );
nor \U$19855 ( \20073 , \20071 , \20072 );
xnor \U$19856 ( \20074 , \20073 , \10121 );
xor \U$19857 ( \20075 , \20070 , \20074 );
xor \U$19858 ( \20076 , \20061 , \20075 );
and \U$19859 ( \20077 , \4364 , \10118 );
not \U$19860 ( \20078 , \20077 );
xor \U$19861 ( \20079 , \20076 , \20078 );
xor \U$19862 ( \20080 , \20057 , \20079 );
xor \U$19863 ( \20081 , \19999 , \20080 );
xor \U$19864 ( \20082 , \19990 , \20081 );
xor \U$19865 ( \20083 , \19961 , \20082 );
and \U$19866 ( \20084 , \19826 , \19948 );
xor \U$19867 ( \20085 , \20083 , \20084 );
and \U$19868 ( \20086 , \19949 , \19950 );
and \U$19869 ( \20087 , \19951 , \19954 );
or \U$19870 ( \20088 , \20086 , \20087 );
xor \U$19871 ( \20089 , \20085 , \20088 );
buf g54cb_GF_PartitionCandidate( \20090_nG54cb , \20089 );
buf \U$19872 ( \20091 , \20090_nG54cb );
and \U$19873 ( \20092 , \19969 , \19973 );
and \U$19874 ( \20093 , \19973 , \19988 );
and \U$19875 ( \20094 , \19969 , \19988 );
or \U$19876 ( \20095 , \20092 , \20093 , \20094 );
and \U$19877 ( \20096 , \19965 , \19989 );
and \U$19878 ( \20097 , \19989 , \20081 );
and \U$19879 ( \20098 , \19965 , \20081 );
or \U$19880 ( \20099 , \20096 , \20097 , \20098 );
xor \U$19881 ( \20100 , \20095 , \20099 );
and \U$19882 ( \20101 , \19994 , \19998 );
and \U$19883 ( \20102 , \19998 , \20080 );
and \U$19884 ( \20103 , \19994 , \20080 );
or \U$19885 ( \20104 , \20101 , \20102 , \20103 );
and \U$19886 ( \20105 , \19978 , \19982 );
and \U$19887 ( \20106 , \19982 , \19987 );
and \U$19888 ( \20107 , \19978 , \19987 );
or \U$19889 ( \20108 , \20105 , \20106 , \20107 );
and \U$19890 ( \20109 , \20013 , \20056 );
and \U$19891 ( \20110 , \20056 , \20079 );
and \U$19892 ( \20111 , \20013 , \20079 );
or \U$19893 ( \20112 , \20109 , \20110 , \20111 );
xor \U$19894 ( \20113 , \20108 , \20112 );
and \U$19895 ( \20114 , \20017 , \20021 );
and \U$19896 ( \20115 , \20021 , \20026 );
and \U$19897 ( \20116 , \20017 , \20026 );
or \U$19898 ( \20117 , \20114 , \20115 , \20116 );
and \U$19899 ( \20118 , \20030 , \20034 );
and \U$19900 ( \20119 , \20034 , \20039 );
and \U$19901 ( \20120 , \20030 , \20039 );
or \U$19902 ( \20121 , \20118 , \20119 , \20120 );
xor \U$19903 ( \20122 , \20117 , \20121 );
and \U$19904 ( \20123 , \20045 , \20049 );
and \U$19905 ( \20124 , \20049 , \20054 );
and \U$19906 ( \20125 , \20045 , \20054 );
or \U$19907 ( \20126 , \20123 , \20124 , \20125 );
xor \U$19908 ( \20127 , \20122 , \20126 );
xor \U$19909 ( \20128 , \20113 , \20127 );
xor \U$19910 ( \20129 , \20104 , \20128 );
and \U$19911 ( \20130 , \20003 , \20007 );
and \U$19912 ( \20131 , \20007 , \20012 );
and \U$19913 ( \20132 , \20003 , \20012 );
or \U$19914 ( \20133 , \20130 , \20131 , \20132 );
and \U$19915 ( \20134 , \20027 , \20040 );
and \U$19916 ( \20135 , \20040 , \20055 );
and \U$19917 ( \20136 , \20027 , \20055 );
or \U$19918 ( \20137 , \20134 , \20135 , \20136 );
xor \U$19919 ( \20138 , \20133 , \20137 );
and \U$19920 ( \20139 , \20061 , \20075 );
and \U$19921 ( \20140 , \20075 , \20078 );
and \U$19922 ( \20141 , \20061 , \20078 );
or \U$19923 ( \20142 , \20139 , \20140 , \20141 );
xor \U$19924 ( \20143 , \20138 , \20142 );
not \U$19925 ( \20144 , \4377 );
and \U$19926 ( \20145 , \10206 , \5011 );
and \U$19927 ( \20146 , \10584 , \4878 );
nor \U$19928 ( \20147 , \20145 , \20146 );
xnor \U$19929 ( \20148 , \20147 , \4762 );
xor \U$19930 ( \20149 , \20144 , \20148 );
and \U$19931 ( \20150 , \9465 , \5485 );
and \U$19932 ( \20151 , \9897 , \5275 );
nor \U$19933 ( \20152 , \20150 , \20151 );
xnor \U$19934 ( \20153 , \20152 , \5169 );
xor \U$19935 ( \20154 , \20149 , \20153 );
and \U$19936 ( \20155 , \20065 , \20069 );
and \U$19937 ( \20156 , \20069 , \20074 );
and \U$19938 ( \20157 , \20065 , \20074 );
or \U$19939 ( \20158 , \20155 , \20156 , \20157 );
buf \U$19940 ( \20159 , \20077 );
xor \U$19941 ( \20160 , \20158 , \20159 );
and \U$19942 ( \20161 , \4654 , \10118 );
xor \U$19943 ( \20162 , \20160 , \20161 );
xor \U$19944 ( \20163 , \20154 , \20162 );
and \U$19945 ( \20164 , \8835 , \5996 );
and \U$19946 ( \20165 , \9169 , \5695 );
nor \U$19947 ( \20166 , \20164 , \20165 );
xnor \U$19948 ( \20167 , \20166 , \5687 );
and \U$19949 ( \20168 , \8349 , \6401 );
and \U$19950 ( \20169 , \8652 , \6143 );
nor \U$19951 ( \20170 , \20168 , \20169 );
xnor \U$19952 ( \20171 , \20170 , \6148 );
xor \U$19953 ( \20172 , \20167 , \20171 );
and \U$19954 ( \20173 , \7700 , \7055 );
and \U$19955 ( \20174 , \8057 , \6675 );
nor \U$19956 ( \20175 , \20173 , \20174 );
xnor \U$19957 ( \20176 , \20175 , \6680 );
xor \U$19958 ( \20177 , \20172 , \20176 );
and \U$19959 ( \20178 , \5674 , \9333 );
and \U$19960 ( \20179 , \6030 , \9006 );
nor \U$19961 ( \20180 , \20178 , \20179 );
xnor \U$19962 ( \20181 , \20180 , \8848 );
and \U$19963 ( \20182 , \5156 , \9765 );
and \U$19964 ( \20183 , \5469 , \9644 );
nor \U$19965 ( \20184 , \20182 , \20183 );
xnor \U$19966 ( \20185 , \20184 , \9478 );
xor \U$19967 ( \20186 , \20181 , \20185 );
and \U$19968 ( \20187 , \4749 , \10408 );
and \U$19969 ( \20188 , \4922 , \10116 );
nor \U$19970 ( \20189 , \20187 , \20188 );
xnor \U$19971 ( \20190 , \20189 , \10121 );
xor \U$19972 ( \20191 , \20186 , \20190 );
xor \U$19973 ( \20192 , \20177 , \20191 );
and \U$19974 ( \20193 , \7231 , \7489 );
and \U$19975 ( \20194 , \7556 , \7137 );
nor \U$19976 ( \20195 , \20193 , \20194 );
xnor \U$19977 ( \20196 , \20195 , \7142 );
and \U$19978 ( \20197 , \6790 , \8019 );
and \U$19979 ( \20198 , \6945 , \7830 );
nor \U$19980 ( \20199 , \20197 , \20198 );
xnor \U$19981 ( \20200 , \20199 , \7713 );
xor \U$19982 ( \20201 , \20196 , \20200 );
and \U$19983 ( \20202 , \6281 , \8540 );
and \U$19984 ( \20203 , \6514 , \8292 );
nor \U$19985 ( \20204 , \20202 , \20203 );
xnor \U$19986 ( \20205 , \20204 , \8297 );
xor \U$19987 ( \20206 , \20201 , \20205 );
xor \U$19988 ( \20207 , \20192 , \20206 );
xor \U$19989 ( \20208 , \20163 , \20207 );
xor \U$19990 ( \20209 , \20143 , \20208 );
xor \U$19991 ( \20210 , \20129 , \20209 );
xor \U$19992 ( \20211 , \20100 , \20210 );
and \U$19993 ( \20212 , \19961 , \20082 );
xor \U$19994 ( \20213 , \20211 , \20212 );
and \U$19995 ( \20214 , \20083 , \20084 );
and \U$19996 ( \20215 , \20085 , \20088 );
or \U$19997 ( \20216 , \20214 , \20215 );
xor \U$19998 ( \20217 , \20213 , \20216 );
buf g54c9_GF_PartitionCandidate( \20218_nG54c9 , \20217 );
buf \U$19999 ( \20219 , \20218_nG54c9 );
and \U$20000 ( \20220 , \20104 , \20128 );
and \U$20001 ( \20221 , \20128 , \20209 );
and \U$20002 ( \20222 , \20104 , \20209 );
or \U$20003 ( \20223 , \20220 , \20221 , \20222 );
and \U$20004 ( \20224 , \20108 , \20112 );
and \U$20005 ( \20225 , \20112 , \20127 );
and \U$20006 ( \20226 , \20108 , \20127 );
or \U$20007 ( \20227 , \20224 , \20225 , \20226 );
and \U$20008 ( \20228 , \20143 , \20208 );
xor \U$20009 ( \20229 , \20227 , \20228 );
and \U$20010 ( \20230 , \20158 , \20159 );
and \U$20011 ( \20231 , \20159 , \20161 );
and \U$20012 ( \20232 , \20158 , \20161 );
or \U$20013 ( \20233 , \20230 , \20231 , \20232 );
and \U$20014 ( \20234 , \20117 , \20121 );
and \U$20015 ( \20235 , \20121 , \20126 );
and \U$20016 ( \20236 , \20117 , \20126 );
or \U$20017 ( \20237 , \20234 , \20235 , \20236 );
xor \U$20018 ( \20238 , \20233 , \20237 );
and \U$20019 ( \20239 , \20177 , \20191 );
and \U$20020 ( \20240 , \20191 , \20206 );
and \U$20021 ( \20241 , \20177 , \20206 );
or \U$20022 ( \20242 , \20239 , \20240 , \20241 );
xor \U$20023 ( \20243 , \20238 , \20242 );
xor \U$20024 ( \20244 , \20229 , \20243 );
xor \U$20025 ( \20245 , \20223 , \20244 );
and \U$20026 ( \20246 , \20133 , \20137 );
and \U$20027 ( \20247 , \20137 , \20142 );
and \U$20028 ( \20248 , \20133 , \20142 );
or \U$20029 ( \20249 , \20246 , \20247 , \20248 );
and \U$20030 ( \20250 , \20154 , \20162 );
and \U$20031 ( \20251 , \20162 , \20207 );
and \U$20032 ( \20252 , \20154 , \20207 );
or \U$20033 ( \20253 , \20250 , \20251 , \20252 );
xor \U$20034 ( \20254 , \20249 , \20253 );
and \U$20035 ( \20255 , \20144 , \20148 );
and \U$20036 ( \20256 , \20148 , \20153 );
and \U$20037 ( \20257 , \20144 , \20153 );
or \U$20038 ( \20258 , \20255 , \20256 , \20257 );
and \U$20039 ( \20259 , \20167 , \20171 );
and \U$20040 ( \20260 , \20171 , \20176 );
and \U$20041 ( \20261 , \20167 , \20176 );
or \U$20042 ( \20262 , \20259 , \20260 , \20261 );
xor \U$20043 ( \20263 , \20258 , \20262 );
and \U$20044 ( \20264 , \20196 , \20200 );
and \U$20045 ( \20265 , \20200 , \20205 );
and \U$20046 ( \20266 , \20196 , \20205 );
or \U$20047 ( \20267 , \20264 , \20265 , \20266 );
xor \U$20048 ( \20268 , \20263 , \20267 );
and \U$20049 ( \20269 , \10584 , \5011 );
not \U$20050 ( \20270 , \20269 );
xnor \U$20051 ( \20271 , \20270 , \4762 );
and \U$20052 ( \20272 , \9897 , \5485 );
and \U$20053 ( \20273 , \10206 , \5275 );
nor \U$20054 ( \20274 , \20272 , \20273 );
xnor \U$20055 ( \20275 , \20274 , \5169 );
xor \U$20056 ( \20276 , \20271 , \20275 );
and \U$20057 ( \20277 , \9169 , \5996 );
and \U$20058 ( \20278 , \9465 , \5695 );
nor \U$20059 ( \20279 , \20277 , \20278 );
xnor \U$20060 ( \20280 , \20279 , \5687 );
xor \U$20061 ( \20281 , \20276 , \20280 );
and \U$20062 ( \20282 , \6945 , \8019 );
and \U$20063 ( \20283 , \7231 , \7830 );
nor \U$20064 ( \20284 , \20282 , \20283 );
xnor \U$20065 ( \20285 , \20284 , \7713 );
and \U$20066 ( \20286 , \6514 , \8540 );
and \U$20067 ( \20287 , \6790 , \8292 );
nor \U$20068 ( \20288 , \20286 , \20287 );
xnor \U$20069 ( \20289 , \20288 , \8297 );
xor \U$20070 ( \20290 , \20285 , \20289 );
and \U$20071 ( \20291 , \6030 , \9333 );
and \U$20072 ( \20292 , \6281 , \9006 );
nor \U$20073 ( \20293 , \20291 , \20292 );
xnor \U$20074 ( \20294 , \20293 , \8848 );
xor \U$20075 ( \20295 , \20290 , \20294 );
xor \U$20076 ( \20296 , \20281 , \20295 );
and \U$20077 ( \20297 , \8652 , \6401 );
and \U$20078 ( \20298 , \8835 , \6143 );
nor \U$20079 ( \20299 , \20297 , \20298 );
xnor \U$20080 ( \20300 , \20299 , \6148 );
and \U$20081 ( \20301 , \8057 , \7055 );
and \U$20082 ( \20302 , \8349 , \6675 );
nor \U$20083 ( \20303 , \20301 , \20302 );
xnor \U$20084 ( \20304 , \20303 , \6680 );
xor \U$20085 ( \20305 , \20300 , \20304 );
and \U$20086 ( \20306 , \7556 , \7489 );
and \U$20087 ( \20307 , \7700 , \7137 );
nor \U$20088 ( \20308 , \20306 , \20307 );
xnor \U$20089 ( \20309 , \20308 , \7142 );
xor \U$20090 ( \20310 , \20305 , \20309 );
xor \U$20091 ( \20311 , \20296 , \20310 );
xor \U$20092 ( \20312 , \20268 , \20311 );
and \U$20093 ( \20313 , \20181 , \20185 );
and \U$20094 ( \20314 , \20185 , \20190 );
and \U$20095 ( \20315 , \20181 , \20190 );
or \U$20096 ( \20316 , \20313 , \20314 , \20315 );
and \U$20097 ( \20317 , \5469 , \9765 );
and \U$20098 ( \20318 , \5674 , \9644 );
nor \U$20099 ( \20319 , \20317 , \20318 );
xnor \U$20100 ( \20320 , \20319 , \9478 );
and \U$20101 ( \20321 , \4922 , \10408 );
and \U$20102 ( \20322 , \5156 , \10116 );
nor \U$20103 ( \20323 , \20321 , \20322 );
xnor \U$20104 ( \20324 , \20323 , \10121 );
xor \U$20105 ( \20325 , \20320 , \20324 );
and \U$20106 ( \20326 , \4749 , \10118 );
xor \U$20107 ( \20327 , \20325 , \20326 );
xnor \U$20108 ( \20328 , \20316 , \20327 );
xor \U$20109 ( \20329 , \20312 , \20328 );
xor \U$20110 ( \20330 , \20254 , \20329 );
xor \U$20111 ( \20331 , \20245 , \20330 );
and \U$20112 ( \20332 , \20095 , \20099 );
and \U$20113 ( \20333 , \20099 , \20210 );
and \U$20114 ( \20334 , \20095 , \20210 );
or \U$20115 ( \20335 , \20332 , \20333 , \20334 );
xor \U$20116 ( \20336 , \20331 , \20335 );
and \U$20117 ( \20337 , \20211 , \20212 );
and \U$20118 ( \20338 , \20213 , \20216 );
or \U$20119 ( \20339 , \20337 , \20338 );
xor \U$20120 ( \20340 , \20336 , \20339 );
buf g54c7_GF_PartitionCandidate( \20341_nG54c7 , \20340 );
buf \U$20121 ( \20342 , \20341_nG54c7 );
and \U$20122 ( \20343 , \20227 , \20228 );
and \U$20123 ( \20344 , \20228 , \20243 );
and \U$20124 ( \20345 , \20227 , \20243 );
or \U$20125 ( \20346 , \20343 , \20344 , \20345 );
and \U$20126 ( \20347 , \20249 , \20253 );
and \U$20127 ( \20348 , \20253 , \20329 );
and \U$20128 ( \20349 , \20249 , \20329 );
or \U$20129 ( \20350 , \20347 , \20348 , \20349 );
and \U$20130 ( \20351 , \20258 , \20262 );
and \U$20131 ( \20352 , \20262 , \20267 );
and \U$20132 ( \20353 , \20258 , \20267 );
or \U$20133 ( \20354 , \20351 , \20352 , \20353 );
and \U$20134 ( \20355 , \20281 , \20295 );
and \U$20135 ( \20356 , \20295 , \20310 );
and \U$20136 ( \20357 , \20281 , \20310 );
or \U$20137 ( \20358 , \20355 , \20356 , \20357 );
xor \U$20138 ( \20359 , \20354 , \20358 );
or \U$20139 ( \20360 , \20316 , \20327 );
xor \U$20140 ( \20361 , \20359 , \20360 );
xor \U$20141 ( \20362 , \20350 , \20361 );
and \U$20142 ( \20363 , \20233 , \20237 );
and \U$20143 ( \20364 , \20237 , \20242 );
and \U$20144 ( \20365 , \20233 , \20242 );
or \U$20145 ( \20366 , \20363 , \20364 , \20365 );
and \U$20146 ( \20367 , \20268 , \20311 );
and \U$20147 ( \20368 , \20311 , \20328 );
and \U$20148 ( \20369 , \20268 , \20328 );
or \U$20149 ( \20370 , \20367 , \20368 , \20369 );
xor \U$20150 ( \20371 , \20366 , \20370 );
and \U$20151 ( \20372 , \20271 , \20275 );
and \U$20152 ( \20373 , \20275 , \20280 );
and \U$20153 ( \20374 , \20271 , \20280 );
or \U$20154 ( \20375 , \20372 , \20373 , \20374 );
and \U$20155 ( \20376 , \20285 , \20289 );
and \U$20156 ( \20377 , \20289 , \20294 );
and \U$20157 ( \20378 , \20285 , \20294 );
or \U$20158 ( \20379 , \20376 , \20377 , \20378 );
xor \U$20159 ( \20380 , \20375 , \20379 );
and \U$20160 ( \20381 , \20300 , \20304 );
and \U$20161 ( \20382 , \20304 , \20309 );
and \U$20162 ( \20383 , \20300 , \20309 );
or \U$20163 ( \20384 , \20381 , \20382 , \20383 );
xor \U$20164 ( \20385 , \20380 , \20384 );
and \U$20165 ( \20386 , \20320 , \20324 );
and \U$20166 ( \20387 , \20324 , \20326 );
and \U$20167 ( \20388 , \20320 , \20326 );
or \U$20168 ( \20389 , \20386 , \20387 , \20388 );
and \U$20169 ( \20390 , \5674 , \9765 );
and \U$20170 ( \20391 , \6030 , \9644 );
nor \U$20171 ( \20392 , \20390 , \20391 );
xnor \U$20172 ( \20393 , \20392 , \9478 );
and \U$20173 ( \20394 , \5156 , \10408 );
and \U$20174 ( \20395 , \5469 , \10116 );
nor \U$20175 ( \20396 , \20394 , \20395 );
xnor \U$20176 ( \20397 , \20396 , \10121 );
xor \U$20177 ( \20398 , \20393 , \20397 );
and \U$20178 ( \20399 , \4922 , \10118 );
xor \U$20179 ( \20400 , \20398 , \20399 );
xor \U$20180 ( \20401 , \20389 , \20400 );
and \U$20181 ( \20402 , \7231 , \8019 );
and \U$20182 ( \20403 , \7556 , \7830 );
nor \U$20183 ( \20404 , \20402 , \20403 );
xnor \U$20184 ( \20405 , \20404 , \7713 );
and \U$20185 ( \20406 , \6790 , \8540 );
and \U$20186 ( \20407 , \6945 , \8292 );
nor \U$20187 ( \20408 , \20406 , \20407 );
xnor \U$20188 ( \20409 , \20408 , \8297 );
xor \U$20189 ( \20410 , \20405 , \20409 );
and \U$20190 ( \20411 , \6281 , \9333 );
and \U$20191 ( \20412 , \6514 , \9006 );
nor \U$20192 ( \20413 , \20411 , \20412 );
xnor \U$20193 ( \20414 , \20413 , \8848 );
xor \U$20194 ( \20415 , \20410 , \20414 );
xor \U$20195 ( \20416 , \20401 , \20415 );
xor \U$20196 ( \20417 , \20385 , \20416 );
not \U$20197 ( \20418 , \4762 );
and \U$20198 ( \20419 , \10206 , \5485 );
and \U$20199 ( \20420 , \10584 , \5275 );
nor \U$20200 ( \20421 , \20419 , \20420 );
xnor \U$20201 ( \20422 , \20421 , \5169 );
xor \U$20202 ( \20423 , \20418 , \20422 );
and \U$20203 ( \20424 , \9465 , \5996 );
and \U$20204 ( \20425 , \9897 , \5695 );
nor \U$20205 ( \20426 , \20424 , \20425 );
xnor \U$20206 ( \20427 , \20426 , \5687 );
xor \U$20207 ( \20428 , \20423 , \20427 );
and \U$20208 ( \20429 , \8835 , \6401 );
and \U$20209 ( \20430 , \9169 , \6143 );
nor \U$20210 ( \20431 , \20429 , \20430 );
xnor \U$20211 ( \20432 , \20431 , \6148 );
and \U$20212 ( \20433 , \8349 , \7055 );
and \U$20213 ( \20434 , \8652 , \6675 );
nor \U$20214 ( \20435 , \20433 , \20434 );
xnor \U$20215 ( \20436 , \20435 , \6680 );
xor \U$20216 ( \20437 , \20432 , \20436 );
and \U$20217 ( \20438 , \7700 , \7489 );
and \U$20218 ( \20439 , \8057 , \7137 );
nor \U$20219 ( \20440 , \20438 , \20439 );
xnor \U$20220 ( \20441 , \20440 , \7142 );
xor \U$20221 ( \20442 , \20437 , \20441 );
xor \U$20222 ( \20443 , \20428 , \20442 );
xor \U$20223 ( \20444 , \20417 , \20443 );
xor \U$20224 ( \20445 , \20371 , \20444 );
xor \U$20225 ( \20446 , \20362 , \20445 );
xor \U$20226 ( \20447 , \20346 , \20446 );
and \U$20227 ( \20448 , \20223 , \20244 );
and \U$20228 ( \20449 , \20244 , \20330 );
and \U$20229 ( \20450 , \20223 , \20330 );
or \U$20230 ( \20451 , \20448 , \20449 , \20450 );
xor \U$20231 ( \20452 , \20447 , \20451 );
and \U$20232 ( \20453 , \20331 , \20335 );
and \U$20233 ( \20454 , \20336 , \20339 );
or \U$20234 ( \20455 , \20453 , \20454 );
xor \U$20235 ( \20456 , \20452 , \20455 );
buf g54c5_GF_PartitionCandidate( \20457_nG54c5 , \20456 );
buf \U$20236 ( \20458 , \20457_nG54c5 );
and \U$20237 ( \20459 , \20350 , \20361 );
and \U$20238 ( \20460 , \20361 , \20445 );
and \U$20239 ( \20461 , \20350 , \20445 );
or \U$20240 ( \20462 , \20459 , \20460 , \20461 );
and \U$20241 ( \20463 , \20366 , \20370 );
and \U$20242 ( \20464 , \20370 , \20444 );
and \U$20243 ( \20465 , \20366 , \20444 );
or \U$20244 ( \20466 , \20463 , \20464 , \20465 );
and \U$20245 ( \20467 , \20375 , \20379 );
and \U$20246 ( \20468 , \20379 , \20384 );
and \U$20247 ( \20469 , \20375 , \20384 );
or \U$20248 ( \20470 , \20467 , \20468 , \20469 );
and \U$20249 ( \20471 , \20389 , \20400 );
and \U$20250 ( \20472 , \20400 , \20415 );
and \U$20251 ( \20473 , \20389 , \20415 );
or \U$20252 ( \20474 , \20471 , \20472 , \20473 );
xor \U$20253 ( \20475 , \20470 , \20474 );
and \U$20254 ( \20476 , \20428 , \20442 );
xor \U$20255 ( \20477 , \20475 , \20476 );
xor \U$20256 ( \20478 , \20466 , \20477 );
and \U$20257 ( \20479 , \20354 , \20358 );
and \U$20258 ( \20480 , \20358 , \20360 );
and \U$20259 ( \20481 , \20354 , \20360 );
or \U$20260 ( \20482 , \20479 , \20480 , \20481 );
and \U$20261 ( \20483 , \20385 , \20416 );
and \U$20262 ( \20484 , \20416 , \20443 );
and \U$20263 ( \20485 , \20385 , \20443 );
or \U$20264 ( \20486 , \20483 , \20484 , \20485 );
xor \U$20265 ( \20487 , \20482 , \20486 );
and \U$20266 ( \20488 , \20418 , \20422 );
and \U$20267 ( \20489 , \20422 , \20427 );
and \U$20268 ( \20490 , \20418 , \20427 );
or \U$20269 ( \20491 , \20488 , \20489 , \20490 );
and \U$20270 ( \20492 , \20405 , \20409 );
and \U$20271 ( \20493 , \20409 , \20414 );
and \U$20272 ( \20494 , \20405 , \20414 );
or \U$20273 ( \20495 , \20492 , \20493 , \20494 );
xor \U$20274 ( \20496 , \20491 , \20495 );
and \U$20275 ( \20497 , \20432 , \20436 );
and \U$20276 ( \20498 , \20436 , \20441 );
and \U$20277 ( \20499 , \20432 , \20441 );
or \U$20278 ( \20500 , \20497 , \20498 , \20499 );
xor \U$20279 ( \20501 , \20496 , \20500 );
and \U$20280 ( \20502 , \20393 , \20397 );
and \U$20281 ( \20503 , \20397 , \20399 );
and \U$20282 ( \20504 , \20393 , \20399 );
or \U$20283 ( \20505 , \20502 , \20503 , \20504 );
and \U$20284 ( \20506 , \6945 , \8540 );
and \U$20285 ( \20507 , \7231 , \8292 );
nor \U$20286 ( \20508 , \20506 , \20507 );
xnor \U$20287 ( \20509 , \20508 , \8297 );
and \U$20288 ( \20510 , \6514 , \9333 );
and \U$20289 ( \20511 , \6790 , \9006 );
nor \U$20290 ( \20512 , \20510 , \20511 );
xnor \U$20291 ( \20513 , \20512 , \8848 );
xor \U$20292 ( \20514 , \20509 , \20513 );
and \U$20293 ( \20515 , \6030 , \9765 );
and \U$20294 ( \20516 , \6281 , \9644 );
nor \U$20295 ( \20517 , \20515 , \20516 );
xnor \U$20296 ( \20518 , \20517 , \9478 );
xor \U$20297 ( \20519 , \20514 , \20518 );
xor \U$20298 ( \20520 , \20505 , \20519 );
and \U$20299 ( \20521 , \5469 , \10408 );
and \U$20300 ( \20522 , \5674 , \10116 );
nor \U$20301 ( \20523 , \20521 , \20522 );
xnor \U$20302 ( \20524 , \20523 , \10121 );
and \U$20303 ( \20525 , \5156 , \10118 );
xnor \U$20304 ( \20526 , \20524 , \20525 );
xor \U$20305 ( \20527 , \20520 , \20526 );
xor \U$20306 ( \20528 , \20501 , \20527 );
and \U$20307 ( \20529 , \8652 , \7055 );
and \U$20308 ( \20530 , \8835 , \6675 );
nor \U$20309 ( \20531 , \20529 , \20530 );
xnor \U$20310 ( \20532 , \20531 , \6680 );
and \U$20311 ( \20533 , \8057 , \7489 );
and \U$20312 ( \20534 , \8349 , \7137 );
nor \U$20313 ( \20535 , \20533 , \20534 );
xnor \U$20314 ( \20536 , \20535 , \7142 );
xor \U$20315 ( \20537 , \20532 , \20536 );
and \U$20316 ( \20538 , \7556 , \8019 );
and \U$20317 ( \20539 , \7700 , \7830 );
nor \U$20318 ( \20540 , \20538 , \20539 );
xnor \U$20319 ( \20541 , \20540 , \7713 );
xor \U$20320 ( \20542 , \20537 , \20541 );
and \U$20321 ( \20543 , \10584 , \5485 );
not \U$20322 ( \20544 , \20543 );
xnor \U$20323 ( \20545 , \20544 , \5169 );
and \U$20324 ( \20546 , \9897 , \5996 );
and \U$20325 ( \20547 , \10206 , \5695 );
nor \U$20326 ( \20548 , \20546 , \20547 );
xnor \U$20327 ( \20549 , \20548 , \5687 );
xor \U$20328 ( \20550 , \20545 , \20549 );
and \U$20329 ( \20551 , \9169 , \6401 );
and \U$20330 ( \20552 , \9465 , \6143 );
nor \U$20331 ( \20553 , \20551 , \20552 );
xnor \U$20332 ( \20554 , \20553 , \6148 );
xor \U$20333 ( \20555 , \20550 , \20554 );
xor \U$20334 ( \20556 , \20542 , \20555 );
xor \U$20335 ( \20557 , \20528 , \20556 );
xor \U$20336 ( \20558 , \20487 , \20557 );
xor \U$20337 ( \20559 , \20478 , \20558 );
xor \U$20338 ( \20560 , \20462 , \20559 );
and \U$20339 ( \20561 , \20346 , \20446 );
xor \U$20340 ( \20562 , \20560 , \20561 );
and \U$20341 ( \20563 , \20447 , \20451 );
and \U$20342 ( \20564 , \20452 , \20455 );
or \U$20343 ( \20565 , \20563 , \20564 );
xor \U$20344 ( \20566 , \20562 , \20565 );
buf g54c3_GF_PartitionCandidate( \20567_nG54c3 , \20566 );
buf \U$20345 ( \20568 , \20567_nG54c3 );
and \U$20346 ( \20569 , \20466 , \20477 );
and \U$20347 ( \20570 , \20477 , \20558 );
and \U$20348 ( \20571 , \20466 , \20558 );
or \U$20349 ( \20572 , \20569 , \20570 , \20571 );
and \U$20350 ( \20573 , \20482 , \20486 );
and \U$20351 ( \20574 , \20486 , \20557 );
and \U$20352 ( \20575 , \20482 , \20557 );
or \U$20353 ( \20576 , \20573 , \20574 , \20575 );
and \U$20354 ( \20577 , \20491 , \20495 );
and \U$20355 ( \20578 , \20495 , \20500 );
and \U$20356 ( \20579 , \20491 , \20500 );
or \U$20357 ( \20580 , \20577 , \20578 , \20579 );
and \U$20358 ( \20581 , \20505 , \20519 );
and \U$20359 ( \20582 , \20519 , \20526 );
and \U$20360 ( \20583 , \20505 , \20526 );
or \U$20361 ( \20584 , \20581 , \20582 , \20583 );
xor \U$20362 ( \20585 , \20580 , \20584 );
and \U$20363 ( \20586 , \20542 , \20555 );
xor \U$20364 ( \20587 , \20585 , \20586 );
xor \U$20365 ( \20588 , \20576 , \20587 );
and \U$20366 ( \20589 , \20470 , \20474 );
and \U$20367 ( \20590 , \20474 , \20476 );
and \U$20368 ( \20591 , \20470 , \20476 );
or \U$20369 ( \20592 , \20589 , \20590 , \20591 );
and \U$20370 ( \20593 , \20501 , \20527 );
and \U$20371 ( \20594 , \20527 , \20556 );
and \U$20372 ( \20595 , \20501 , \20556 );
or \U$20373 ( \20596 , \20593 , \20594 , \20595 );
xor \U$20374 ( \20597 , \20592 , \20596 );
and \U$20375 ( \20598 , \20509 , \20513 );
and \U$20376 ( \20599 , \20513 , \20518 );
and \U$20377 ( \20600 , \20509 , \20518 );
or \U$20378 ( \20601 , \20598 , \20599 , \20600 );
and \U$20379 ( \20602 , \20532 , \20536 );
and \U$20380 ( \20603 , \20536 , \20541 );
and \U$20381 ( \20604 , \20532 , \20541 );
or \U$20382 ( \20605 , \20602 , \20603 , \20604 );
xor \U$20383 ( \20606 , \20601 , \20605 );
and \U$20384 ( \20607 , \20545 , \20549 );
and \U$20385 ( \20608 , \20549 , \20554 );
and \U$20386 ( \20609 , \20545 , \20554 );
or \U$20387 ( \20610 , \20607 , \20608 , \20609 );
xor \U$20388 ( \20611 , \20606 , \20610 );
or \U$20389 ( \20612 , \20524 , \20525 );
and \U$20390 ( \20613 , \5674 , \10408 );
and \U$20391 ( \20614 , \6030 , \10116 );
nor \U$20392 ( \20615 , \20613 , \20614 );
xnor \U$20393 ( \20616 , \20615 , \10121 );
xor \U$20394 ( \20617 , \20612 , \20616 );
and \U$20395 ( \20618 , \5469 , \10118 );
xor \U$20396 ( \20619 , \20617 , \20618 );
xor \U$20397 ( \20620 , \20611 , \20619 );
not \U$20398 ( \20621 , \5169 );
and \U$20399 ( \20622 , \10206 , \5996 );
and \U$20400 ( \20623 , \10584 , \5695 );
nor \U$20401 ( \20624 , \20622 , \20623 );
xnor \U$20402 ( \20625 , \20624 , \5687 );
xor \U$20403 ( \20626 , \20621 , \20625 );
and \U$20404 ( \20627 , \9465 , \6401 );
and \U$20405 ( \20628 , \9897 , \6143 );
nor \U$20406 ( \20629 , \20627 , \20628 );
xnor \U$20407 ( \20630 , \20629 , \6148 );
xor \U$20408 ( \20631 , \20626 , \20630 );
and \U$20409 ( \20632 , \8835 , \7055 );
and \U$20410 ( \20633 , \9169 , \6675 );
nor \U$20411 ( \20634 , \20632 , \20633 );
xnor \U$20412 ( \20635 , \20634 , \6680 );
and \U$20413 ( \20636 , \8349 , \7489 );
and \U$20414 ( \20637 , \8652 , \7137 );
nor \U$20415 ( \20638 , \20636 , \20637 );
xnor \U$20416 ( \20639 , \20638 , \7142 );
xor \U$20417 ( \20640 , \20635 , \20639 );
and \U$20418 ( \20641 , \7700 , \8019 );
and \U$20419 ( \20642 , \8057 , \7830 );
nor \U$20420 ( \20643 , \20641 , \20642 );
xnor \U$20421 ( \20644 , \20643 , \7713 );
xor \U$20422 ( \20645 , \20640 , \20644 );
xor \U$20423 ( \20646 , \20631 , \20645 );
and \U$20424 ( \20647 , \7231 , \8540 );
and \U$20425 ( \20648 , \7556 , \8292 );
nor \U$20426 ( \20649 , \20647 , \20648 );
xnor \U$20427 ( \20650 , \20649 , \8297 );
and \U$20428 ( \20651 , \6790 , \9333 );
and \U$20429 ( \20652 , \6945 , \9006 );
nor \U$20430 ( \20653 , \20651 , \20652 );
xnor \U$20431 ( \20654 , \20653 , \8848 );
xor \U$20432 ( \20655 , \20650 , \20654 );
and \U$20433 ( \20656 , \6281 , \9765 );
and \U$20434 ( \20657 , \6514 , \9644 );
nor \U$20435 ( \20658 , \20656 , \20657 );
xnor \U$20436 ( \20659 , \20658 , \9478 );
xor \U$20437 ( \20660 , \20655 , \20659 );
xor \U$20438 ( \20661 , \20646 , \20660 );
xor \U$20439 ( \20662 , \20620 , \20661 );
xor \U$20440 ( \20663 , \20597 , \20662 );
xor \U$20441 ( \20664 , \20588 , \20663 );
xor \U$20442 ( \20665 , \20572 , \20664 );
and \U$20443 ( \20666 , \20462 , \20559 );
xor \U$20444 ( \20667 , \20665 , \20666 );
and \U$20445 ( \20668 , \20560 , \20561 );
and \U$20446 ( \20669 , \20562 , \20565 );
or \U$20447 ( \20670 , \20668 , \20669 );
xor \U$20448 ( \20671 , \20667 , \20670 );
buf g54c1_GF_PartitionCandidate( \20672_nG54c1 , \20671 );
buf \U$20449 ( \20673 , \20672_nG54c1 );
and \U$20450 ( \20674 , \20576 , \20587 );
and \U$20451 ( \20675 , \20587 , \20663 );
and \U$20452 ( \20676 , \20576 , \20663 );
or \U$20453 ( \20677 , \20674 , \20675 , \20676 );
and \U$20454 ( \20678 , \20592 , \20596 );
and \U$20455 ( \20679 , \20596 , \20662 );
and \U$20456 ( \20680 , \20592 , \20662 );
or \U$20457 ( \20681 , \20678 , \20679 , \20680 );
and \U$20458 ( \20682 , \20601 , \20605 );
and \U$20459 ( \20683 , \20605 , \20610 );
and \U$20460 ( \20684 , \20601 , \20610 );
or \U$20461 ( \20685 , \20682 , \20683 , \20684 );
and \U$20462 ( \20686 , \20612 , \20616 );
and \U$20463 ( \20687 , \20616 , \20618 );
and \U$20464 ( \20688 , \20612 , \20618 );
or \U$20465 ( \20689 , \20686 , \20687 , \20688 );
xor \U$20466 ( \20690 , \20685 , \20689 );
and \U$20467 ( \20691 , \20631 , \20645 );
and \U$20468 ( \20692 , \20645 , \20660 );
and \U$20469 ( \20693 , \20631 , \20660 );
or \U$20470 ( \20694 , \20691 , \20692 , \20693 );
xor \U$20471 ( \20695 , \20690 , \20694 );
xor \U$20472 ( \20696 , \20681 , \20695 );
and \U$20473 ( \20697 , \20580 , \20584 );
and \U$20474 ( \20698 , \20584 , \20586 );
and \U$20475 ( \20699 , \20580 , \20586 );
or \U$20476 ( \20700 , \20697 , \20698 , \20699 );
and \U$20477 ( \20701 , \20611 , \20619 );
and \U$20478 ( \20702 , \20619 , \20661 );
and \U$20479 ( \20703 , \20611 , \20661 );
or \U$20480 ( \20704 , \20701 , \20702 , \20703 );
xor \U$20481 ( \20705 , \20700 , \20704 );
and \U$20482 ( \20706 , \20621 , \20625 );
and \U$20483 ( \20707 , \20625 , \20630 );
and \U$20484 ( \20708 , \20621 , \20630 );
or \U$20485 ( \20709 , \20706 , \20707 , \20708 );
and \U$20486 ( \20710 , \20635 , \20639 );
and \U$20487 ( \20711 , \20639 , \20644 );
and \U$20488 ( \20712 , \20635 , \20644 );
or \U$20489 ( \20713 , \20710 , \20711 , \20712 );
xor \U$20490 ( \20714 , \20709 , \20713 );
and \U$20491 ( \20715 , \20650 , \20654 );
and \U$20492 ( \20716 , \20654 , \20659 );
and \U$20493 ( \20717 , \20650 , \20659 );
or \U$20494 ( \20718 , \20715 , \20716 , \20717 );
xor \U$20495 ( \20719 , \20714 , \20718 );
and \U$20496 ( \20720 , \5674 , \10118 );
and \U$20497 ( \20721 , \6945 , \9333 );
and \U$20498 ( \20722 , \7231 , \9006 );
nor \U$20499 ( \20723 , \20721 , \20722 );
xnor \U$20500 ( \20724 , \20723 , \8848 );
and \U$20501 ( \20725 , \6514 , \9765 );
and \U$20502 ( \20726 , \6790 , \9644 );
nor \U$20503 ( \20727 , \20725 , \20726 );
xnor \U$20504 ( \20728 , \20727 , \9478 );
xor \U$20505 ( \20729 , \20724 , \20728 );
and \U$20506 ( \20730 , \6030 , \10408 );
and \U$20507 ( \20731 , \6281 , \10116 );
nor \U$20508 ( \20732 , \20730 , \20731 );
xnor \U$20509 ( \20733 , \20732 , \10121 );
xor \U$20510 ( \20734 , \20729 , \20733 );
xnor \U$20511 ( \20735 , \20720 , \20734 );
xor \U$20512 ( \20736 , \20719 , \20735 );
and \U$20513 ( \20737 , \8652 , \7489 );
and \U$20514 ( \20738 , \8835 , \7137 );
nor \U$20515 ( \20739 , \20737 , \20738 );
xnor \U$20516 ( \20740 , \20739 , \7142 );
and \U$20517 ( \20741 , \8057 , \8019 );
and \U$20518 ( \20742 , \8349 , \7830 );
nor \U$20519 ( \20743 , \20741 , \20742 );
xnor \U$20520 ( \20744 , \20743 , \7713 );
xor \U$20521 ( \20745 , \20740 , \20744 );
and \U$20522 ( \20746 , \7556 , \8540 );
and \U$20523 ( \20747 , \7700 , \8292 );
nor \U$20524 ( \20748 , \20746 , \20747 );
xnor \U$20525 ( \20749 , \20748 , \8297 );
xor \U$20526 ( \20750 , \20745 , \20749 );
and \U$20527 ( \20751 , \10584 , \5996 );
not \U$20528 ( \20752 , \20751 );
xnor \U$20529 ( \20753 , \20752 , \5687 );
and \U$20530 ( \20754 , \9897 , \6401 );
and \U$20531 ( \20755 , \10206 , \6143 );
nor \U$20532 ( \20756 , \20754 , \20755 );
xnor \U$20533 ( \20757 , \20756 , \6148 );
xor \U$20534 ( \20758 , \20753 , \20757 );
and \U$20535 ( \20759 , \9169 , \7055 );
and \U$20536 ( \20760 , \9465 , \6675 );
nor \U$20537 ( \20761 , \20759 , \20760 );
xnor \U$20538 ( \20762 , \20761 , \6680 );
xor \U$20539 ( \20763 , \20758 , \20762 );
xor \U$20540 ( \20764 , \20750 , \20763 );
xor \U$20541 ( \20765 , \20736 , \20764 );
xor \U$20542 ( \20766 , \20705 , \20765 );
xor \U$20543 ( \20767 , \20696 , \20766 );
xor \U$20544 ( \20768 , \20677 , \20767 );
and \U$20545 ( \20769 , \20572 , \20664 );
xor \U$20546 ( \20770 , \20768 , \20769 );
and \U$20547 ( \20771 , \20665 , \20666 );
and \U$20548 ( \20772 , \20667 , \20670 );
or \U$20549 ( \20773 , \20771 , \20772 );
xor \U$20550 ( \20774 , \20770 , \20773 );
buf g54bf_GF_PartitionCandidate( \20775_nG54bf , \20774 );
buf \U$20551 ( \20776 , \20775_nG54bf );
and \U$20552 ( \20777 , \20681 , \20695 );
and \U$20553 ( \20778 , \20695 , \20766 );
and \U$20554 ( \20779 , \20681 , \20766 );
or \U$20555 ( \20780 , \20777 , \20778 , \20779 );
and \U$20556 ( \20781 , \20700 , \20704 );
and \U$20557 ( \20782 , \20704 , \20765 );
and \U$20558 ( \20783 , \20700 , \20765 );
or \U$20559 ( \20784 , \20781 , \20782 , \20783 );
and \U$20560 ( \20785 , \20709 , \20713 );
and \U$20561 ( \20786 , \20713 , \20718 );
and \U$20562 ( \20787 , \20709 , \20718 );
or \U$20563 ( \20788 , \20785 , \20786 , \20787 );
or \U$20564 ( \20789 , \20720 , \20734 );
xor \U$20565 ( \20790 , \20788 , \20789 );
and \U$20566 ( \20791 , \20750 , \20763 );
xor \U$20567 ( \20792 , \20790 , \20791 );
xor \U$20568 ( \20793 , \20784 , \20792 );
and \U$20569 ( \20794 , \20685 , \20689 );
and \U$20570 ( \20795 , \20689 , \20694 );
and \U$20571 ( \20796 , \20685 , \20694 );
or \U$20572 ( \20797 , \20794 , \20795 , \20796 );
and \U$20573 ( \20798 , \20719 , \20735 );
and \U$20574 ( \20799 , \20735 , \20764 );
and \U$20575 ( \20800 , \20719 , \20764 );
or \U$20576 ( \20801 , \20798 , \20799 , \20800 );
xor \U$20577 ( \20802 , \20797 , \20801 );
not \U$20578 ( \20803 , \5687 );
and \U$20579 ( \20804 , \10206 , \6401 );
and \U$20580 ( \20805 , \10584 , \6143 );
nor \U$20581 ( \20806 , \20804 , \20805 );
xnor \U$20582 ( \20807 , \20806 , \6148 );
xor \U$20583 ( \20808 , \20803 , \20807 );
and \U$20584 ( \20809 , \9465 , \7055 );
and \U$20585 ( \20810 , \9897 , \6675 );
nor \U$20586 ( \20811 , \20809 , \20810 );
xnor \U$20587 ( \20812 , \20811 , \6680 );
xor \U$20588 ( \20813 , \20808 , \20812 );
and \U$20589 ( \20814 , \20740 , \20744 );
and \U$20590 ( \20815 , \20744 , \20749 );
and \U$20591 ( \20816 , \20740 , \20749 );
or \U$20592 ( \20817 , \20814 , \20815 , \20816 );
and \U$20593 ( \20818 , \20753 , \20757 );
and \U$20594 ( \20819 , \20757 , \20762 );
and \U$20595 ( \20820 , \20753 , \20762 );
or \U$20596 ( \20821 , \20818 , \20819 , \20820 );
xor \U$20597 ( \20822 , \20817 , \20821 );
and \U$20598 ( \20823 , \20724 , \20728 );
and \U$20599 ( \20824 , \20728 , \20733 );
and \U$20600 ( \20825 , \20724 , \20733 );
or \U$20601 ( \20826 , \20823 , \20824 , \20825 );
xor \U$20602 ( \20827 , \20822 , \20826 );
xor \U$20603 ( \20828 , \20813 , \20827 );
and \U$20604 ( \20829 , \6030 , \10118 );
and \U$20605 ( \20830 , \8835 , \7489 );
and \U$20606 ( \20831 , \9169 , \7137 );
nor \U$20607 ( \20832 , \20830 , \20831 );
xnor \U$20608 ( \20833 , \20832 , \7142 );
and \U$20609 ( \20834 , \8349 , \8019 );
and \U$20610 ( \20835 , \8652 , \7830 );
nor \U$20611 ( \20836 , \20834 , \20835 );
xnor \U$20612 ( \20837 , \20836 , \7713 );
xor \U$20613 ( \20838 , \20833 , \20837 );
and \U$20614 ( \20839 , \7700 , \8540 );
and \U$20615 ( \20840 , \8057 , \8292 );
nor \U$20616 ( \20841 , \20839 , \20840 );
xnor \U$20617 ( \20842 , \20841 , \8297 );
xor \U$20618 ( \20843 , \20838 , \20842 );
xor \U$20619 ( \20844 , \20829 , \20843 );
and \U$20620 ( \20845 , \7231 , \9333 );
and \U$20621 ( \20846 , \7556 , \9006 );
nor \U$20622 ( \20847 , \20845 , \20846 );
xnor \U$20623 ( \20848 , \20847 , \8848 );
and \U$20624 ( \20849 , \6790 , \9765 );
and \U$20625 ( \20850 , \6945 , \9644 );
nor \U$20626 ( \20851 , \20849 , \20850 );
xnor \U$20627 ( \20852 , \20851 , \9478 );
xor \U$20628 ( \20853 , \20848 , \20852 );
and \U$20629 ( \20854 , \6281 , \10408 );
and \U$20630 ( \20855 , \6514 , \10116 );
nor \U$20631 ( \20856 , \20854 , \20855 );
xnor \U$20632 ( \20857 , \20856 , \10121 );
xor \U$20633 ( \20858 , \20853 , \20857 );
xor \U$20634 ( \20859 , \20844 , \20858 );
xor \U$20635 ( \20860 , \20828 , \20859 );
xor \U$20636 ( \20861 , \20802 , \20860 );
xor \U$20637 ( \20862 , \20793 , \20861 );
xor \U$20638 ( \20863 , \20780 , \20862 );
and \U$20639 ( \20864 , \20677 , \20767 );
xor \U$20640 ( \20865 , \20863 , \20864 );
and \U$20641 ( \20866 , \20768 , \20769 );
and \U$20642 ( \20867 , \20770 , \20773 );
or \U$20643 ( \20868 , \20866 , \20867 );
xor \U$20644 ( \20869 , \20865 , \20868 );
buf g54bd_GF_PartitionCandidate( \20870_nG54bd , \20869 );
buf \U$20645 ( \20871 , \20870_nG54bd );
and \U$20646 ( \20872 , \20784 , \20792 );
and \U$20647 ( \20873 , \20792 , \20861 );
and \U$20648 ( \20874 , \20784 , \20861 );
or \U$20649 ( \20875 , \20872 , \20873 , \20874 );
and \U$20650 ( \20876 , \20797 , \20801 );
and \U$20651 ( \20877 , \20801 , \20860 );
and \U$20652 ( \20878 , \20797 , \20860 );
or \U$20653 ( \20879 , \20876 , \20877 , \20878 );
and \U$20654 ( \20880 , \20788 , \20789 );
and \U$20655 ( \20881 , \20789 , \20791 );
and \U$20656 ( \20882 , \20788 , \20791 );
or \U$20657 ( \20883 , \20880 , \20881 , \20882 );
and \U$20658 ( \20884 , \20813 , \20827 );
and \U$20659 ( \20885 , \20827 , \20859 );
and \U$20660 ( \20886 , \20813 , \20859 );
or \U$20661 ( \20887 , \20884 , \20885 , \20886 );
xor \U$20662 ( \20888 , \20883 , \20887 );
and \U$20663 ( \20889 , \6945 , \9765 );
and \U$20664 ( \20890 , \7231 , \9644 );
nor \U$20665 ( \20891 , \20889 , \20890 );
xnor \U$20666 ( \20892 , \20891 , \9478 );
and \U$20667 ( \20893 , \6514 , \10408 );
and \U$20668 ( \20894 , \6790 , \10116 );
nor \U$20669 ( \20895 , \20893 , \20894 );
xnor \U$20670 ( \20896 , \20895 , \10121 );
xor \U$20671 ( \20897 , \20892 , \20896 );
and \U$20672 ( \20898 , \6281 , \10118 );
xor \U$20673 ( \20899 , \20897 , \20898 );
and \U$20674 ( \20900 , \8652 , \8019 );
and \U$20675 ( \20901 , \8835 , \7830 );
nor \U$20676 ( \20902 , \20900 , \20901 );
xnor \U$20677 ( \20903 , \20902 , \7713 );
and \U$20678 ( \20904 , \8057 , \8540 );
and \U$20679 ( \20905 , \8349 , \8292 );
nor \U$20680 ( \20906 , \20904 , \20905 );
xnor \U$20681 ( \20907 , \20906 , \8297 );
xor \U$20682 ( \20908 , \20903 , \20907 );
and \U$20683 ( \20909 , \7556 , \9333 );
and \U$20684 ( \20910 , \7700 , \9006 );
nor \U$20685 ( \20911 , \20909 , \20910 );
xnor \U$20686 ( \20912 , \20911 , \8848 );
xor \U$20687 ( \20913 , \20908 , \20912 );
xnor \U$20688 ( \20914 , \20899 , \20913 );
xor \U$20689 ( \20915 , \20888 , \20914 );
xor \U$20690 ( \20916 , \20879 , \20915 );
and \U$20691 ( \20917 , \20833 , \20837 );
and \U$20692 ( \20918 , \20837 , \20842 );
and \U$20693 ( \20919 , \20833 , \20842 );
or \U$20694 ( \20920 , \20917 , \20918 , \20919 );
and \U$20695 ( \20921 , \20803 , \20807 );
and \U$20696 ( \20922 , \20807 , \20812 );
and \U$20697 ( \20923 , \20803 , \20812 );
or \U$20698 ( \20924 , \20921 , \20922 , \20923 );
xor \U$20699 ( \20925 , \20920 , \20924 );
and \U$20700 ( \20926 , \20848 , \20852 );
and \U$20701 ( \20927 , \20852 , \20857 );
and \U$20702 ( \20928 , \20848 , \20857 );
or \U$20703 ( \20929 , \20926 , \20927 , \20928 );
xor \U$20704 ( \20930 , \20925 , \20929 );
and \U$20705 ( \20931 , \20817 , \20821 );
and \U$20706 ( \20932 , \20821 , \20826 );
and \U$20707 ( \20933 , \20817 , \20826 );
or \U$20708 ( \20934 , \20931 , \20932 , \20933 );
and \U$20709 ( \20935 , \20829 , \20843 );
and \U$20710 ( \20936 , \20843 , \20858 );
and \U$20711 ( \20937 , \20829 , \20858 );
or \U$20712 ( \20938 , \20935 , \20936 , \20937 );
xor \U$20713 ( \20939 , \20934 , \20938 );
and \U$20714 ( \20940 , \10584 , \6401 );
not \U$20715 ( \20941 , \20940 );
xnor \U$20716 ( \20942 , \20941 , \6148 );
and \U$20717 ( \20943 , \9897 , \7055 );
and \U$20718 ( \20944 , \10206 , \6675 );
nor \U$20719 ( \20945 , \20943 , \20944 );
xnor \U$20720 ( \20946 , \20945 , \6680 );
xor \U$20721 ( \20947 , \20942 , \20946 );
and \U$20722 ( \20948 , \9169 , \7489 );
and \U$20723 ( \20949 , \9465 , \7137 );
nor \U$20724 ( \20950 , \20948 , \20949 );
xnor \U$20725 ( \20951 , \20950 , \7142 );
xor \U$20726 ( \20952 , \20947 , \20951 );
xor \U$20727 ( \20953 , \20939 , \20952 );
xor \U$20728 ( \20954 , \20930 , \20953 );
xor \U$20729 ( \20955 , \20916 , \20954 );
xor \U$20730 ( \20956 , \20875 , \20955 );
and \U$20731 ( \20957 , \20780 , \20862 );
xor \U$20732 ( \20958 , \20956 , \20957 );
and \U$20733 ( \20959 , \20863 , \20864 );
and \U$20734 ( \20960 , \20865 , \20868 );
or \U$20735 ( \20961 , \20959 , \20960 );
xor \U$20736 ( \20962 , \20958 , \20961 );
buf g54bb_GF_PartitionCandidate( \20963_nG54bb , \20962 );
buf \U$20737 ( \20964 , \20963_nG54bb );
and \U$20738 ( \20965 , \20879 , \20915 );
and \U$20739 ( \20966 , \20915 , \20954 );
and \U$20740 ( \20967 , \20879 , \20954 );
or \U$20741 ( \20968 , \20965 , \20966 , \20967 );
and \U$20742 ( \20969 , \20883 , \20887 );
and \U$20743 ( \20970 , \20887 , \20914 );
and \U$20744 ( \20971 , \20883 , \20914 );
or \U$20745 ( \20972 , \20969 , \20970 , \20971 );
and \U$20746 ( \20973 , \20930 , \20953 );
xor \U$20747 ( \20974 , \20972 , \20973 );
and \U$20748 ( \20975 , \20934 , \20938 );
and \U$20749 ( \20976 , \20938 , \20952 );
and \U$20750 ( \20977 , \20934 , \20952 );
or \U$20751 ( \20978 , \20975 , \20976 , \20977 );
and \U$20752 ( \20979 , \20892 , \20896 );
and \U$20753 ( \20980 , \20896 , \20898 );
and \U$20754 ( \20981 , \20892 , \20898 );
or \U$20755 ( \20982 , \20979 , \20980 , \20981 );
and \U$20756 ( \20983 , \20942 , \20946 );
and \U$20757 ( \20984 , \20946 , \20951 );
and \U$20758 ( \20985 , \20942 , \20951 );
or \U$20759 ( \20986 , \20983 , \20984 , \20985 );
xor \U$20760 ( \20987 , \20982 , \20986 );
and \U$20761 ( \20988 , \20903 , \20907 );
and \U$20762 ( \20989 , \20907 , \20912 );
and \U$20763 ( \20990 , \20903 , \20912 );
or \U$20764 ( \20991 , \20988 , \20989 , \20990 );
xor \U$20765 ( \20992 , \20987 , \20991 );
xor \U$20766 ( \20993 , \20978 , \20992 );
and \U$20767 ( \20994 , \20920 , \20924 );
and \U$20768 ( \20995 , \20924 , \20929 );
and \U$20769 ( \20996 , \20920 , \20929 );
or \U$20770 ( \20997 , \20994 , \20995 , \20996 );
or \U$20771 ( \20998 , \20899 , \20913 );
xor \U$20772 ( \20999 , \20997 , \20998 );
not \U$20773 ( \21000 , \6148 );
and \U$20774 ( \21001 , \10206 , \7055 );
and \U$20775 ( \21002 , \10584 , \6675 );
nor \U$20776 ( \21003 , \21001 , \21002 );
xnor \U$20777 ( \21004 , \21003 , \6680 );
xor \U$20778 ( \21005 , \21000 , \21004 );
and \U$20779 ( \21006 , \9465 , \7489 );
and \U$20780 ( \21007 , \9897 , \7137 );
nor \U$20781 ( \21008 , \21006 , \21007 );
xnor \U$20782 ( \21009 , \21008 , \7142 );
xor \U$20783 ( \21010 , \21005 , \21009 );
and \U$20784 ( \21011 , \7231 , \9765 );
and \U$20785 ( \21012 , \7556 , \9644 );
nor \U$20786 ( \21013 , \21011 , \21012 );
xnor \U$20787 ( \21014 , \21013 , \9478 );
and \U$20788 ( \21015 , \6790 , \10408 );
and \U$20789 ( \21016 , \6945 , \10116 );
nor \U$20790 ( \21017 , \21015 , \21016 );
xnor \U$20791 ( \21018 , \21017 , \10121 );
xor \U$20792 ( \21019 , \21014 , \21018 );
and \U$20793 ( \21020 , \6514 , \10118 );
xor \U$20794 ( \21021 , \21019 , \21020 );
xor \U$20795 ( \21022 , \21010 , \21021 );
and \U$20796 ( \21023 , \8835 , \8019 );
and \U$20797 ( \21024 , \9169 , \7830 );
nor \U$20798 ( \21025 , \21023 , \21024 );
xnor \U$20799 ( \21026 , \21025 , \7713 );
and \U$20800 ( \21027 , \8349 , \8540 );
and \U$20801 ( \21028 , \8652 , \8292 );
nor \U$20802 ( \21029 , \21027 , \21028 );
xnor \U$20803 ( \21030 , \21029 , \8297 );
xor \U$20804 ( \21031 , \21026 , \21030 );
and \U$20805 ( \21032 , \7700 , \9333 );
and \U$20806 ( \21033 , \8057 , \9006 );
nor \U$20807 ( \21034 , \21032 , \21033 );
xnor \U$20808 ( \21035 , \21034 , \8848 );
xor \U$20809 ( \21036 , \21031 , \21035 );
xor \U$20810 ( \21037 , \21022 , \21036 );
xor \U$20811 ( \21038 , \20999 , \21037 );
xor \U$20812 ( \21039 , \20993 , \21038 );
xor \U$20813 ( \21040 , \20974 , \21039 );
xor \U$20814 ( \21041 , \20968 , \21040 );
and \U$20815 ( \21042 , \20875 , \20955 );
xor \U$20816 ( \21043 , \21041 , \21042 );
and \U$20817 ( \21044 , \20956 , \20957 );
and \U$20818 ( \21045 , \20958 , \20961 );
or \U$20819 ( \21046 , \21044 , \21045 );
xor \U$20820 ( \21047 , \21043 , \21046 );
buf g54b9_GF_PartitionCandidate( \21048_nG54b9 , \21047 );
buf \U$20821 ( \21049 , \21048_nG54b9 );
and \U$20822 ( \21050 , \20978 , \20992 );
and \U$20823 ( \21051 , \20992 , \21038 );
and \U$20824 ( \21052 , \20978 , \21038 );
or \U$20825 ( \21053 , \21050 , \21051 , \21052 );
and \U$20826 ( \21054 , \20972 , \20973 );
and \U$20827 ( \21055 , \20973 , \21039 );
and \U$20828 ( \21056 , \20972 , \21039 );
or \U$20829 ( \21057 , \21054 , \21055 , \21056 );
xor \U$20830 ( \21058 , \21053 , \21057 );
and \U$20831 ( \21059 , \20997 , \20998 );
and \U$20832 ( \21060 , \20998 , \21037 );
and \U$20833 ( \21061 , \20997 , \21037 );
or \U$20834 ( \21062 , \21059 , \21060 , \21061 );
and \U$20835 ( \21063 , \21000 , \21004 );
and \U$20836 ( \21064 , \21004 , \21009 );
and \U$20837 ( \21065 , \21000 , \21009 );
or \U$20838 ( \21066 , \21063 , \21064 , \21065 );
and \U$20839 ( \21067 , \21014 , \21018 );
and \U$20840 ( \21068 , \21018 , \21020 );
and \U$20841 ( \21069 , \21014 , \21020 );
or \U$20842 ( \21070 , \21067 , \21068 , \21069 );
xor \U$20843 ( \21071 , \21066 , \21070 );
and \U$20844 ( \21072 , \21026 , \21030 );
and \U$20845 ( \21073 , \21030 , \21035 );
and \U$20846 ( \21074 , \21026 , \21035 );
or \U$20847 ( \21075 , \21072 , \21073 , \21074 );
xor \U$20848 ( \21076 , \21071 , \21075 );
xor \U$20849 ( \21077 , \21062 , \21076 );
and \U$20850 ( \21078 , \20982 , \20986 );
and \U$20851 ( \21079 , \20986 , \20991 );
and \U$20852 ( \21080 , \20982 , \20991 );
or \U$20853 ( \21081 , \21078 , \21079 , \21080 );
and \U$20854 ( \21082 , \21010 , \21021 );
and \U$20855 ( \21083 , \21021 , \21036 );
and \U$20856 ( \21084 , \21010 , \21036 );
or \U$20857 ( \21085 , \21082 , \21083 , \21084 );
xor \U$20858 ( \21086 , \21081 , \21085 );
and \U$20859 ( \21087 , \10584 , \7055 );
not \U$20860 ( \21088 , \21087 );
xnor \U$20861 ( \21089 , \21088 , \6680 );
and \U$20862 ( \21090 , \9897 , \7489 );
and \U$20863 ( \21091 , \10206 , \7137 );
nor \U$20864 ( \21092 , \21090 , \21091 );
xnor \U$20865 ( \21093 , \21092 , \7142 );
xor \U$20866 ( \21094 , \21089 , \21093 );
and \U$20867 ( \21095 , \9169 , \8019 );
and \U$20868 ( \21096 , \9465 , \7830 );
nor \U$20869 ( \21097 , \21095 , \21096 );
xnor \U$20870 ( \21098 , \21097 , \7713 );
xor \U$20871 ( \21099 , \21094 , \21098 );
and \U$20872 ( \21100 , \8652 , \8540 );
and \U$20873 ( \21101 , \8835 , \8292 );
nor \U$20874 ( \21102 , \21100 , \21101 );
xnor \U$20875 ( \21103 , \21102 , \8297 );
and \U$20876 ( \21104 , \8057 , \9333 );
and \U$20877 ( \21105 , \8349 , \9006 );
nor \U$20878 ( \21106 , \21104 , \21105 );
xnor \U$20879 ( \21107 , \21106 , \8848 );
xor \U$20880 ( \21108 , \21103 , \21107 );
and \U$20881 ( \21109 , \7556 , \9765 );
and \U$20882 ( \21110 , \7700 , \9644 );
nor \U$20883 ( \21111 , \21109 , \21110 );
xnor \U$20884 ( \21112 , \21111 , \9478 );
xor \U$20885 ( \21113 , \21108 , \21112 );
xor \U$20886 ( \21114 , \21099 , \21113 );
and \U$20887 ( \21115 , \6945 , \10408 );
and \U$20888 ( \21116 , \7231 , \10116 );
nor \U$20889 ( \21117 , \21115 , \21116 );
xnor \U$20890 ( \21118 , \21117 , \10121 );
and \U$20891 ( \21119 , \6790 , \10118 );
xnor \U$20892 ( \21120 , \21118 , \21119 );
xor \U$20893 ( \21121 , \21114 , \21120 );
xor \U$20894 ( \21122 , \21086 , \21121 );
xor \U$20895 ( \21123 , \21077 , \21122 );
xor \U$20896 ( \21124 , \21058 , \21123 );
and \U$20897 ( \21125 , \20968 , \21040 );
xor \U$20898 ( \21126 , \21124 , \21125 );
and \U$20899 ( \21127 , \21041 , \21042 );
and \U$20900 ( \21128 , \21043 , \21046 );
or \U$20901 ( \21129 , \21127 , \21128 );
xor \U$20902 ( \21130 , \21126 , \21129 );
buf g54b7_GF_PartitionCandidate( \21131_nG54b7 , \21130 );
buf \U$20903 ( \21132 , \21131_nG54b7 );
and \U$20904 ( \21133 , \21062 , \21076 );
and \U$20905 ( \21134 , \21076 , \21122 );
and \U$20906 ( \21135 , \21062 , \21122 );
or \U$20907 ( \21136 , \21133 , \21134 , \21135 );
and \U$20908 ( \21137 , \21081 , \21085 );
and \U$20909 ( \21138 , \21085 , \21121 );
and \U$20910 ( \21139 , \21081 , \21121 );
or \U$20911 ( \21140 , \21137 , \21138 , \21139 );
and \U$20912 ( \21141 , \21089 , \21093 );
and \U$20913 ( \21142 , \21093 , \21098 );
and \U$20914 ( \21143 , \21089 , \21098 );
or \U$20915 ( \21144 , \21141 , \21142 , \21143 );
and \U$20916 ( \21145 , \21103 , \21107 );
and \U$20917 ( \21146 , \21107 , \21112 );
and \U$20918 ( \21147 , \21103 , \21112 );
or \U$20919 ( \21148 , \21145 , \21146 , \21147 );
xor \U$20920 ( \21149 , \21144 , \21148 );
or \U$20921 ( \21150 , \21118 , \21119 );
xor \U$20922 ( \21151 , \21149 , \21150 );
xor \U$20923 ( \21152 , \21140 , \21151 );
and \U$20924 ( \21153 , \21066 , \21070 );
and \U$20925 ( \21154 , \21070 , \21075 );
and \U$20926 ( \21155 , \21066 , \21075 );
or \U$20927 ( \21156 , \21153 , \21154 , \21155 );
and \U$20928 ( \21157 , \21099 , \21113 );
and \U$20929 ( \21158 , \21113 , \21120 );
and \U$20930 ( \21159 , \21099 , \21120 );
or \U$20931 ( \21160 , \21157 , \21158 , \21159 );
xor \U$20932 ( \21161 , \21156 , \21160 );
not \U$20933 ( \21162 , \6680 );
and \U$20934 ( \21163 , \10206 , \7489 );
and \U$20935 ( \21164 , \10584 , \7137 );
nor \U$20936 ( \21165 , \21163 , \21164 );
xnor \U$20937 ( \21166 , \21165 , \7142 );
xor \U$20938 ( \21167 , \21162 , \21166 );
and \U$20939 ( \21168 , \9465 , \8019 );
and \U$20940 ( \21169 , \9897 , \7830 );
nor \U$20941 ( \21170 , \21168 , \21169 );
xnor \U$20942 ( \21171 , \21170 , \7713 );
xor \U$20943 ( \21172 , \21167 , \21171 );
and \U$20944 ( \21173 , \8835 , \8540 );
and \U$20945 ( \21174 , \9169 , \8292 );
nor \U$20946 ( \21175 , \21173 , \21174 );
xnor \U$20947 ( \21176 , \21175 , \8297 );
and \U$20948 ( \21177 , \8349 , \9333 );
and \U$20949 ( \21178 , \8652 , \9006 );
nor \U$20950 ( \21179 , \21177 , \21178 );
xnor \U$20951 ( \21180 , \21179 , \8848 );
xor \U$20952 ( \21181 , \21176 , \21180 );
and \U$20953 ( \21182 , \7700 , \9765 );
and \U$20954 ( \21183 , \8057 , \9644 );
nor \U$20955 ( \21184 , \21182 , \21183 );
xnor \U$20956 ( \21185 , \21184 , \9478 );
xor \U$20957 ( \21186 , \21181 , \21185 );
xor \U$20958 ( \21187 , \21172 , \21186 );
and \U$20959 ( \21188 , \7231 , \10408 );
and \U$20960 ( \21189 , \7556 , \10116 );
nor \U$20961 ( \21190 , \21188 , \21189 );
xnor \U$20962 ( \21191 , \21190 , \10121 );
and \U$20963 ( \21192 , \6945 , \10118 );
xor \U$20964 ( \21193 , \21191 , \21192 );
xor \U$20965 ( \21194 , \21187 , \21193 );
xor \U$20966 ( \21195 , \21161 , \21194 );
xor \U$20967 ( \21196 , \21152 , \21195 );
xor \U$20968 ( \21197 , \21136 , \21196 );
and \U$20969 ( \21198 , \21053 , \21057 );
and \U$20970 ( \21199 , \21057 , \21123 );
and \U$20971 ( \21200 , \21053 , \21123 );
or \U$20972 ( \21201 , \21198 , \21199 , \21200 );
xor \U$20973 ( \21202 , \21197 , \21201 );
and \U$20974 ( \21203 , \21124 , \21125 );
and \U$20975 ( \21204 , \21126 , \21129 );
or \U$20976 ( \21205 , \21203 , \21204 );
xor \U$20977 ( \21206 , \21202 , \21205 );
buf g54b5_GF_PartitionCandidate( \21207_nG54b5 , \21206 );
buf \U$20978 ( \21208 , \21207_nG54b5 );
and \U$20979 ( \21209 , \21140 , \21151 );
and \U$20980 ( \21210 , \21151 , \21195 );
and \U$20981 ( \21211 , \21140 , \21195 );
or \U$20982 ( \21212 , \21209 , \21210 , \21211 );
and \U$20983 ( \21213 , \21156 , \21160 );
and \U$20984 ( \21214 , \21160 , \21194 );
and \U$20985 ( \21215 , \21156 , \21194 );
or \U$20986 ( \21216 , \21213 , \21214 , \21215 );
and \U$20987 ( \21217 , \21162 , \21166 );
and \U$20988 ( \21218 , \21166 , \21171 );
and \U$20989 ( \21219 , \21162 , \21171 );
or \U$20990 ( \21220 , \21217 , \21218 , \21219 );
and \U$20991 ( \21221 , \21176 , \21180 );
and \U$20992 ( \21222 , \21180 , \21185 );
and \U$20993 ( \21223 , \21176 , \21185 );
or \U$20994 ( \21224 , \21221 , \21222 , \21223 );
xor \U$20995 ( \21225 , \21220 , \21224 );
and \U$20996 ( \21226 , \21191 , \21192 );
xor \U$20997 ( \21227 , \21225 , \21226 );
xor \U$20998 ( \21228 , \21216 , \21227 );
and \U$20999 ( \21229 , \21144 , \21148 );
and \U$21000 ( \21230 , \21148 , \21150 );
and \U$21001 ( \21231 , \21144 , \21150 );
or \U$21002 ( \21232 , \21229 , \21230 , \21231 );
and \U$21003 ( \21233 , \21172 , \21186 );
and \U$21004 ( \21234 , \21186 , \21193 );
and \U$21005 ( \21235 , \21172 , \21193 );
or \U$21006 ( \21236 , \21233 , \21234 , \21235 );
xor \U$21007 ( \21237 , \21232 , \21236 );
and \U$21008 ( \21238 , \8652 , \9333 );
and \U$21009 ( \21239 , \8835 , \9006 );
nor \U$21010 ( \21240 , \21238 , \21239 );
xnor \U$21011 ( \21241 , \21240 , \8848 );
and \U$21012 ( \21242 , \8057 , \9765 );
and \U$21013 ( \21243 , \8349 , \9644 );
nor \U$21014 ( \21244 , \21242 , \21243 );
xnor \U$21015 ( \21245 , \21244 , \9478 );
xor \U$21016 ( \21246 , \21241 , \21245 );
and \U$21017 ( \21247 , \7556 , \10408 );
and \U$21018 ( \21248 , \7700 , \10116 );
nor \U$21019 ( \21249 , \21247 , \21248 );
xnor \U$21020 ( \21250 , \21249 , \10121 );
xor \U$21021 ( \21251 , \21246 , \21250 );
and \U$21022 ( \21252 , \10584 , \7489 );
not \U$21023 ( \21253 , \21252 );
xnor \U$21024 ( \21254 , \21253 , \7142 );
and \U$21025 ( \21255 , \9897 , \8019 );
and \U$21026 ( \21256 , \10206 , \7830 );
nor \U$21027 ( \21257 , \21255 , \21256 );
xnor \U$21028 ( \21258 , \21257 , \7713 );
xor \U$21029 ( \21259 , \21254 , \21258 );
and \U$21030 ( \21260 , \9169 , \8540 );
and \U$21031 ( \21261 , \9465 , \8292 );
nor \U$21032 ( \21262 , \21260 , \21261 );
xnor \U$21033 ( \21263 , \21262 , \8297 );
xor \U$21034 ( \21264 , \21259 , \21263 );
xor \U$21035 ( \21265 , \21251 , \21264 );
and \U$21036 ( \21266 , \7231 , \10118 );
not \U$21037 ( \21267 , \21266 );
xor \U$21038 ( \21268 , \21265 , \21267 );
xor \U$21039 ( \21269 , \21237 , \21268 );
xor \U$21040 ( \21270 , \21228 , \21269 );
xor \U$21041 ( \21271 , \21212 , \21270 );
and \U$21042 ( \21272 , \21136 , \21196 );
xor \U$21043 ( \21273 , \21271 , \21272 );
and \U$21044 ( \21274 , \21197 , \21201 );
and \U$21045 ( \21275 , \21202 , \21205 );
or \U$21046 ( \21276 , \21274 , \21275 );
xor \U$21047 ( \21277 , \21273 , \21276 );
buf g54b3_GF_PartitionCandidate( \21278_nG54b3 , \21277 );
buf \U$21048 ( \21279 , \21278_nG54b3 );
and \U$21049 ( \21280 , \21216 , \21227 );
and \U$21050 ( \21281 , \21227 , \21269 );
and \U$21051 ( \21282 , \21216 , \21269 );
or \U$21052 ( \21283 , \21280 , \21281 , \21282 );
and \U$21053 ( \21284 , \21232 , \21236 );
and \U$21054 ( \21285 , \21236 , \21268 );
and \U$21055 ( \21286 , \21232 , \21268 );
or \U$21056 ( \21287 , \21284 , \21285 , \21286 );
and \U$21057 ( \21288 , \21241 , \21245 );
and \U$21058 ( \21289 , \21245 , \21250 );
and \U$21059 ( \21290 , \21241 , \21250 );
or \U$21060 ( \21291 , \21288 , \21289 , \21290 );
and \U$21061 ( \21292 , \21254 , \21258 );
and \U$21062 ( \21293 , \21258 , \21263 );
and \U$21063 ( \21294 , \21254 , \21263 );
or \U$21064 ( \21295 , \21292 , \21293 , \21294 );
xor \U$21065 ( \21296 , \21291 , \21295 );
buf \U$21066 ( \21297 , \21266 );
xor \U$21067 ( \21298 , \21296 , \21297 );
xor \U$21068 ( \21299 , \21287 , \21298 );
and \U$21069 ( \21300 , \21220 , \21224 );
and \U$21070 ( \21301 , \21224 , \21226 );
and \U$21071 ( \21302 , \21220 , \21226 );
or \U$21072 ( \21303 , \21300 , \21301 , \21302 );
and \U$21073 ( \21304 , \21251 , \21264 );
and \U$21074 ( \21305 , \21264 , \21267 );
and \U$21075 ( \21306 , \21251 , \21267 );
or \U$21076 ( \21307 , \21304 , \21305 , \21306 );
xor \U$21077 ( \21308 , \21303 , \21307 );
and \U$21078 ( \21309 , \7556 , \10118 );
and \U$21079 ( \21310 , \8835 , \9333 );
and \U$21080 ( \21311 , \9169 , \9006 );
nor \U$21081 ( \21312 , \21310 , \21311 );
xnor \U$21082 ( \21313 , \21312 , \8848 );
and \U$21083 ( \21314 , \8349 , \9765 );
and \U$21084 ( \21315 , \8652 , \9644 );
nor \U$21085 ( \21316 , \21314 , \21315 );
xnor \U$21086 ( \21317 , \21316 , \9478 );
xor \U$21087 ( \21318 , \21313 , \21317 );
and \U$21088 ( \21319 , \7700 , \10408 );
and \U$21089 ( \21320 , \8057 , \10116 );
nor \U$21090 ( \21321 , \21319 , \21320 );
xnor \U$21091 ( \21322 , \21321 , \10121 );
xor \U$21092 ( \21323 , \21318 , \21322 );
xor \U$21093 ( \21324 , \21309 , \21323 );
not \U$21094 ( \21325 , \7142 );
and \U$21095 ( \21326 , \10206 , \8019 );
and \U$21096 ( \21327 , \10584 , \7830 );
nor \U$21097 ( \21328 , \21326 , \21327 );
xnor \U$21098 ( \21329 , \21328 , \7713 );
xor \U$21099 ( \21330 , \21325 , \21329 );
and \U$21100 ( \21331 , \9465 , \8540 );
and \U$21101 ( \21332 , \9897 , \8292 );
nor \U$21102 ( \21333 , \21331 , \21332 );
xnor \U$21103 ( \21334 , \21333 , \8297 );
xor \U$21104 ( \21335 , \21330 , \21334 );
xor \U$21105 ( \21336 , \21324 , \21335 );
xor \U$21106 ( \21337 , \21308 , \21336 );
xor \U$21107 ( \21338 , \21299 , \21337 );
xor \U$21108 ( \21339 , \21283 , \21338 );
and \U$21109 ( \21340 , \21212 , \21270 );
xor \U$21110 ( \21341 , \21339 , \21340 );
and \U$21111 ( \21342 , \21271 , \21272 );
and \U$21112 ( \21343 , \21273 , \21276 );
or \U$21113 ( \21344 , \21342 , \21343 );
xor \U$21114 ( \21345 , \21341 , \21344 );
buf g54b1_GF_PartitionCandidate( \21346_nG54b1 , \21345 );
buf \U$21115 ( \21347 , \21346_nG54b1 );
and \U$21116 ( \21348 , \21287 , \21298 );
and \U$21117 ( \21349 , \21298 , \21337 );
and \U$21118 ( \21350 , \21287 , \21337 );
or \U$21119 ( \21351 , \21348 , \21349 , \21350 );
and \U$21120 ( \21352 , \21303 , \21307 );
and \U$21121 ( \21353 , \21307 , \21336 );
and \U$21122 ( \21354 , \21303 , \21336 );
or \U$21123 ( \21355 , \21352 , \21353 , \21354 );
and \U$21124 ( \21356 , \21291 , \21295 );
and \U$21125 ( \21357 , \21295 , \21297 );
and \U$21126 ( \21358 , \21291 , \21297 );
or \U$21127 ( \21359 , \21356 , \21357 , \21358 );
and \U$21128 ( \21360 , \21309 , \21323 );
and \U$21129 ( \21361 , \21323 , \21335 );
and \U$21130 ( \21362 , \21309 , \21335 );
or \U$21131 ( \21363 , \21360 , \21361 , \21362 );
xor \U$21132 ( \21364 , \21359 , \21363 );
and \U$21133 ( \21365 , \8652 , \9765 );
and \U$21134 ( \21366 , \8835 , \9644 );
nor \U$21135 ( \21367 , \21365 , \21366 );
xnor \U$21136 ( \21368 , \21367 , \9478 );
and \U$21137 ( \21369 , \8057 , \10408 );
and \U$21138 ( \21370 , \8349 , \10116 );
nor \U$21139 ( \21371 , \21369 , \21370 );
xnor \U$21140 ( \21372 , \21371 , \10121 );
xor \U$21141 ( \21373 , \21368 , \21372 );
and \U$21142 ( \21374 , \7700 , \10118 );
xor \U$21143 ( \21375 , \21373 , \21374 );
xor \U$21144 ( \21376 , \21364 , \21375 );
xor \U$21145 ( \21377 , \21355 , \21376 );
and \U$21146 ( \21378 , \10584 , \8019 );
not \U$21147 ( \21379 , \21378 );
xnor \U$21148 ( \21380 , \21379 , \7713 );
and \U$21149 ( \21381 , \9897 , \8540 );
and \U$21150 ( \21382 , \10206 , \8292 );
nor \U$21151 ( \21383 , \21381 , \21382 );
xnor \U$21152 ( \21384 , \21383 , \8297 );
xor \U$21153 ( \21385 , \21380 , \21384 );
and \U$21154 ( \21386 , \9169 , \9333 );
and \U$21155 ( \21387 , \9465 , \9006 );
nor \U$21156 ( \21388 , \21386 , \21387 );
xnor \U$21157 ( \21389 , \21388 , \8848 );
xor \U$21158 ( \21390 , \21385 , \21389 );
and \U$21159 ( \21391 , \21313 , \21317 );
and \U$21160 ( \21392 , \21317 , \21322 );
and \U$21161 ( \21393 , \21313 , \21322 );
or \U$21162 ( \21394 , \21391 , \21392 , \21393 );
and \U$21163 ( \21395 , \21325 , \21329 );
and \U$21164 ( \21396 , \21329 , \21334 );
and \U$21165 ( \21397 , \21325 , \21334 );
or \U$21166 ( \21398 , \21395 , \21396 , \21397 );
xnor \U$21167 ( \21399 , \21394 , \21398 );
xor \U$21168 ( \21400 , \21390 , \21399 );
xor \U$21169 ( \21401 , \21377 , \21400 );
xor \U$21170 ( \21402 , \21351 , \21401 );
and \U$21171 ( \21403 , \21283 , \21338 );
xor \U$21172 ( \21404 , \21402 , \21403 );
and \U$21173 ( \21405 , \21339 , \21340 );
and \U$21174 ( \21406 , \21341 , \21344 );
or \U$21175 ( \21407 , \21405 , \21406 );
xor \U$21176 ( \21408 , \21404 , \21407 );
buf g54af_GF_PartitionCandidate( \21409_nG54af , \21408 );
buf \U$21177 ( \21410 , \21409_nG54af );
and \U$21178 ( \21411 , \21355 , \21376 );
and \U$21179 ( \21412 , \21376 , \21400 );
and \U$21180 ( \21413 , \21355 , \21400 );
or \U$21181 ( \21414 , \21411 , \21412 , \21413 );
and \U$21182 ( \21415 , \21359 , \21363 );
and \U$21183 ( \21416 , \21363 , \21375 );
and \U$21184 ( \21417 , \21359 , \21375 );
or \U$21185 ( \21418 , \21415 , \21416 , \21417 );
and \U$21186 ( \21419 , \21390 , \21399 );
xor \U$21187 ( \21420 , \21418 , \21419 );
or \U$21188 ( \21421 , \21394 , \21398 );
not \U$21189 ( \21422 , \7713 );
and \U$21190 ( \21423 , \10206 , \8540 );
and \U$21191 ( \21424 , \10584 , \8292 );
nor \U$21192 ( \21425 , \21423 , \21424 );
xnor \U$21193 ( \21426 , \21425 , \8297 );
xor \U$21194 ( \21427 , \21422 , \21426 );
and \U$21195 ( \21428 , \9465 , \9333 );
and \U$21196 ( \21429 , \9897 , \9006 );
nor \U$21197 ( \21430 , \21428 , \21429 );
xnor \U$21198 ( \21431 , \21430 , \8848 );
xor \U$21199 ( \21432 , \21427 , \21431 );
xor \U$21200 ( \21433 , \21421 , \21432 );
and \U$21201 ( \21434 , \21380 , \21384 );
and \U$21202 ( \21435 , \21384 , \21389 );
and \U$21203 ( \21436 , \21380 , \21389 );
or \U$21204 ( \21437 , \21434 , \21435 , \21436 );
and \U$21205 ( \21438 , \21368 , \21372 );
and \U$21206 ( \21439 , \21372 , \21374 );
and \U$21207 ( \21440 , \21368 , \21374 );
or \U$21208 ( \21441 , \21438 , \21439 , \21440 );
xor \U$21209 ( \21442 , \21437 , \21441 );
and \U$21210 ( \21443 , \8835 , \9765 );
and \U$21211 ( \21444 , \9169 , \9644 );
nor \U$21212 ( \21445 , \21443 , \21444 );
xnor \U$21213 ( \21446 , \21445 , \9478 );
and \U$21214 ( \21447 , \8349 , \10408 );
and \U$21215 ( \21448 , \8652 , \10116 );
nor \U$21216 ( \21449 , \21447 , \21448 );
xnor \U$21217 ( \21450 , \21449 , \10121 );
xor \U$21218 ( \21451 , \21446 , \21450 );
and \U$21219 ( \21452 , \8057 , \10118 );
xor \U$21220 ( \21453 , \21451 , \21452 );
xor \U$21221 ( \21454 , \21442 , \21453 );
xor \U$21222 ( \21455 , \21433 , \21454 );
xor \U$21223 ( \21456 , \21420 , \21455 );
xor \U$21224 ( \21457 , \21414 , \21456 );
and \U$21225 ( \21458 , \21351 , \21401 );
xor \U$21226 ( \21459 , \21457 , \21458 );
and \U$21227 ( \21460 , \21402 , \21403 );
and \U$21228 ( \21461 , \21404 , \21407 );
or \U$21229 ( \21462 , \21460 , \21461 );
xor \U$21230 ( \21463 , \21459 , \21462 );
buf g54ad_GF_PartitionCandidate( \21464_nG54ad , \21463 );
buf \U$21231 ( \21465 , \21464_nG54ad );
and \U$21232 ( \21466 , \21421 , \21432 );
and \U$21233 ( \21467 , \21432 , \21454 );
and \U$21234 ( \21468 , \21421 , \21454 );
or \U$21235 ( \21469 , \21466 , \21467 , \21468 );
and \U$21236 ( \21470 , \21418 , \21419 );
and \U$21237 ( \21471 , \21419 , \21455 );
and \U$21238 ( \21472 , \21418 , \21455 );
or \U$21239 ( \21473 , \21470 , \21471 , \21472 );
xor \U$21240 ( \21474 , \21469 , \21473 );
and \U$21241 ( \21475 , \21437 , \21441 );
and \U$21242 ( \21476 , \21441 , \21453 );
and \U$21243 ( \21477 , \21437 , \21453 );
or \U$21244 ( \21478 , \21475 , \21476 , \21477 );
and \U$21245 ( \21479 , \10584 , \8540 );
not \U$21246 ( \21480 , \21479 );
xnor \U$21247 ( \21481 , \21480 , \8297 );
and \U$21248 ( \21482 , \9897 , \9333 );
and \U$21249 ( \21483 , \10206 , \9006 );
nor \U$21250 ( \21484 , \21482 , \21483 );
xnor \U$21251 ( \21485 , \21484 , \8848 );
xor \U$21252 ( \21486 , \21481 , \21485 );
and \U$21253 ( \21487 , \9169 , \9765 );
and \U$21254 ( \21488 , \9465 , \9644 );
nor \U$21255 ( \21489 , \21487 , \21488 );
xnor \U$21256 ( \21490 , \21489 , \9478 );
xor \U$21257 ( \21491 , \21486 , \21490 );
xor \U$21258 ( \21492 , \21478 , \21491 );
and \U$21259 ( \21493 , \21422 , \21426 );
and \U$21260 ( \21494 , \21426 , \21431 );
and \U$21261 ( \21495 , \21422 , \21431 );
or \U$21262 ( \21496 , \21493 , \21494 , \21495 );
and \U$21263 ( \21497 , \21446 , \21450 );
and \U$21264 ( \21498 , \21450 , \21452 );
and \U$21265 ( \21499 , \21446 , \21452 );
or \U$21266 ( \21500 , \21497 , \21498 , \21499 );
xor \U$21267 ( \21501 , \21496 , \21500 );
and \U$21268 ( \21502 , \8652 , \10408 );
and \U$21269 ( \21503 , \8835 , \10116 );
nor \U$21270 ( \21504 , \21502 , \21503 );
xnor \U$21271 ( \21505 , \21504 , \10121 );
and \U$21272 ( \21506 , \8349 , \10118 );
xnor \U$21273 ( \21507 , \21505 , \21506 );
xor \U$21274 ( \21508 , \21501 , \21507 );
xor \U$21275 ( \21509 , \21492 , \21508 );
xor \U$21276 ( \21510 , \21474 , \21509 );
and \U$21277 ( \21511 , \21414 , \21456 );
xor \U$21278 ( \21512 , \21510 , \21511 );
and \U$21279 ( \21513 , \21457 , \21458 );
and \U$21280 ( \21514 , \21459 , \21462 );
or \U$21281 ( \21515 , \21513 , \21514 );
xor \U$21282 ( \21516 , \21512 , \21515 );
buf g54ab_GF_PartitionCandidate( \21517_nG54ab , \21516 );
buf \U$21283 ( \21518 , \21517_nG54ab );
and \U$21284 ( \21519 , \21478 , \21491 );
and \U$21285 ( \21520 , \21491 , \21508 );
and \U$21286 ( \21521 , \21478 , \21508 );
or \U$21287 ( \21522 , \21519 , \21520 , \21521 );
and \U$21288 ( \21523 , \21496 , \21500 );
and \U$21289 ( \21524 , \21500 , \21507 );
and \U$21290 ( \21525 , \21496 , \21507 );
or \U$21291 ( \21526 , \21523 , \21524 , \21525 );
and \U$21292 ( \21527 , \21481 , \21485 );
and \U$21293 ( \21528 , \21485 , \21490 );
and \U$21294 ( \21529 , \21481 , \21490 );
or \U$21295 ( \21530 , \21527 , \21528 , \21529 );
or \U$21296 ( \21531 , \21505 , \21506 );
xor \U$21297 ( \21532 , \21530 , \21531 );
and \U$21298 ( \21533 , \8835 , \10408 );
and \U$21299 ( \21534 , \9169 , \10116 );
nor \U$21300 ( \21535 , \21533 , \21534 );
xnor \U$21301 ( \21536 , \21535 , \10121 );
xor \U$21302 ( \21537 , \21532 , \21536 );
xor \U$21303 ( \21538 , \21526 , \21537 );
and \U$21304 ( \21539 , \8652 , \10118 );
not \U$21305 ( \21540 , \8297 );
and \U$21306 ( \21541 , \10206 , \9333 );
and \U$21307 ( \21542 , \10584 , \9006 );
nor \U$21308 ( \21543 , \21541 , \21542 );
xnor \U$21309 ( \21544 , \21543 , \8848 );
xor \U$21310 ( \21545 , \21540 , \21544 );
and \U$21311 ( \21546 , \9465 , \9765 );
and \U$21312 ( \21547 , \9897 , \9644 );
nor \U$21313 ( \21548 , \21546 , \21547 );
xnor \U$21314 ( \21549 , \21548 , \9478 );
xor \U$21315 ( \21550 , \21545 , \21549 );
xor \U$21316 ( \21551 , \21539 , \21550 );
xor \U$21317 ( \21552 , \21538 , \21551 );
xor \U$21318 ( \21553 , \21522 , \21552 );
and \U$21319 ( \21554 , \21469 , \21473 );
and \U$21320 ( \21555 , \21473 , \21509 );
and \U$21321 ( \21556 , \21469 , \21509 );
or \U$21322 ( \21557 , \21554 , \21555 , \21556 );
xor \U$21323 ( \21558 , \21553 , \21557 );
and \U$21324 ( \21559 , \21510 , \21511 );
and \U$21325 ( \21560 , \21512 , \21515 );
or \U$21326 ( \21561 , \21559 , \21560 );
xor \U$21327 ( \21562 , \21558 , \21561 );
buf g54a9_GF_PartitionCandidate( \21563_nG54a9 , \21562 );
buf \U$21328 ( \21564 , \21563_nG54a9 );
and \U$21329 ( \21565 , \21526 , \21537 );
and \U$21330 ( \21566 , \21537 , \21551 );
and \U$21331 ( \21567 , \21526 , \21551 );
or \U$21332 ( \21568 , \21565 , \21566 , \21567 );
and \U$21333 ( \21569 , \21530 , \21531 );
and \U$21334 ( \21570 , \21531 , \21536 );
and \U$21335 ( \21571 , \21530 , \21536 );
or \U$21336 ( \21572 , \21569 , \21570 , \21571 );
and \U$21337 ( \21573 , \21539 , \21550 );
xor \U$21338 ( \21574 , \21572 , \21573 );
and \U$21339 ( \21575 , \21540 , \21544 );
and \U$21340 ( \21576 , \21544 , \21549 );
and \U$21341 ( \21577 , \21540 , \21549 );
or \U$21342 ( \21578 , \21575 , \21576 , \21577 );
and \U$21343 ( \21579 , \10584 , \9333 );
not \U$21344 ( \21580 , \21579 );
xnor \U$21345 ( \21581 , \21580 , \8848 );
and \U$21346 ( \21582 , \9897 , \9765 );
and \U$21347 ( \21583 , \10206 , \9644 );
nor \U$21348 ( \21584 , \21582 , \21583 );
xnor \U$21349 ( \21585 , \21584 , \9478 );
xor \U$21350 ( \21586 , \21581 , \21585 );
and \U$21351 ( \21587 , \9169 , \10408 );
and \U$21352 ( \21588 , \9465 , \10116 );
nor \U$21353 ( \21589 , \21587 , \21588 );
xnor \U$21354 ( \21590 , \21589 , \10121 );
xor \U$21355 ( \21591 , \21586 , \21590 );
xor \U$21356 ( \21592 , \21578 , \21591 );
and \U$21357 ( \21593 , \8835 , \10118 );
not \U$21358 ( \21594 , \21593 );
xor \U$21359 ( \21595 , \21592 , \21594 );
xor \U$21360 ( \21596 , \21574 , \21595 );
xor \U$21361 ( \21597 , \21568 , \21596 );
and \U$21362 ( \21598 , \21522 , \21552 );
xor \U$21363 ( \21599 , \21597 , \21598 );
and \U$21364 ( \21600 , \21553 , \21557 );
and \U$21365 ( \21601 , \21558 , \21561 );
or \U$21366 ( \21602 , \21600 , \21601 );
xor \U$21367 ( \21603 , \21599 , \21602 );
buf g54a7_GF_PartitionCandidate( \21604_nG54a7 , \21603 );
buf \U$21368 ( \21605 , \21604_nG54a7 );
and \U$21369 ( \21606 , \21572 , \21573 );
and \U$21370 ( \21607 , \21573 , \21595 );
and \U$21371 ( \21608 , \21572 , \21595 );
or \U$21372 ( \21609 , \21606 , \21607 , \21608 );
and \U$21373 ( \21610 , \21578 , \21591 );
and \U$21374 ( \21611 , \21591 , \21594 );
and \U$21375 ( \21612 , \21578 , \21594 );
or \U$21376 ( \21613 , \21610 , \21611 , \21612 );
not \U$21377 ( \21614 , \8848 );
and \U$21378 ( \21615 , \10206 , \9765 );
and \U$21379 ( \21616 , \10584 , \9644 );
nor \U$21380 ( \21617 , \21615 , \21616 );
xnor \U$21381 ( \21618 , \21617 , \9478 );
xor \U$21382 ( \21619 , \21614 , \21618 );
and \U$21383 ( \21620 , \9465 , \10408 );
and \U$21384 ( \21621 , \9897 , \10116 );
nor \U$21385 ( \21622 , \21620 , \21621 );
xnor \U$21386 ( \21623 , \21622 , \10121 );
xor \U$21387 ( \21624 , \21619 , \21623 );
xor \U$21388 ( \21625 , \21613 , \21624 );
and \U$21389 ( \21626 , \21581 , \21585 );
and \U$21390 ( \21627 , \21585 , \21590 );
and \U$21391 ( \21628 , \21581 , \21590 );
or \U$21392 ( \21629 , \21626 , \21627 , \21628 );
buf \U$21393 ( \21630 , \21593 );
xor \U$21394 ( \21631 , \21629 , \21630 );
and \U$21395 ( \21632 , \9169 , \10118 );
xor \U$21396 ( \21633 , \21631 , \21632 );
xor \U$21397 ( \21634 , \21625 , \21633 );
xor \U$21398 ( \21635 , \21609 , \21634 );
and \U$21399 ( \21636 , \21568 , \21596 );
xor \U$21400 ( \21637 , \21635 , \21636 );
and \U$21401 ( \21638 , \21597 , \21598 );
and \U$21402 ( \21639 , \21599 , \21602 );
or \U$21403 ( \21640 , \21638 , \21639 );
xor \U$21404 ( \21641 , \21637 , \21640 );
buf g54a5_GF_PartitionCandidate( \21642_nG54a5 , \21641 );
buf \U$21405 ( \21643 , \21642_nG54a5 );
and \U$21406 ( \21644 , \21629 , \21630 );
and \U$21407 ( \21645 , \21630 , \21632 );
and \U$21408 ( \21646 , \21629 , \21632 );
or \U$21409 ( \21647 , \21644 , \21645 , \21646 );
and \U$21410 ( \21648 , \21613 , \21624 );
and \U$21411 ( \21649 , \21624 , \21633 );
and \U$21412 ( \21650 , \21613 , \21633 );
or \U$21413 ( \21651 , \21648 , \21649 , \21650 );
xor \U$21414 ( \21652 , \21647 , \21651 );
and \U$21415 ( \21653 , \21614 , \21618 );
and \U$21416 ( \21654 , \21618 , \21623 );
and \U$21417 ( \21655 , \21614 , \21623 );
or \U$21418 ( \21656 , \21653 , \21654 , \21655 );
and \U$21419 ( \21657 , \10584 , \9765 );
not \U$21420 ( \21658 , \21657 );
xnor \U$21421 ( \21659 , \21658 , \9478 );
and \U$21422 ( \21660 , \9897 , \10408 );
and \U$21423 ( \21661 , \10206 , \10116 );
nor \U$21424 ( \21662 , \21660 , \21661 );
xnor \U$21425 ( \21663 , \21662 , \10121 );
xor \U$21426 ( \21664 , \21659 , \21663 );
and \U$21427 ( \21665 , \9465 , \10118 );
xor \U$21428 ( \21666 , \21664 , \21665 );
xnor \U$21429 ( \21667 , \21656 , \21666 );
xor \U$21430 ( \21668 , \21652 , \21667 );
and \U$21431 ( \21669 , \21609 , \21634 );
xor \U$21432 ( \21670 , \21668 , \21669 );
and \U$21433 ( \21671 , \21635 , \21636 );
and \U$21434 ( \21672 , \21637 , \21640 );
or \U$21435 ( \21673 , \21671 , \21672 );
xor \U$21436 ( \21674 , \21670 , \21673 );
buf g54a3_GF_PartitionCandidate( \21675_nG54a3 , \21674 );
buf \U$21437 ( \21676 , \21675_nG54a3 );
and \U$21438 ( \21677 , \21659 , \21663 );
and \U$21439 ( \21678 , \21663 , \21665 );
and \U$21440 ( \21679 , \21659 , \21665 );
or \U$21441 ( \21680 , \21677 , \21678 , \21679 );
or \U$21442 ( \21681 , \21656 , \21666 );
xor \U$21443 ( \21682 , \21680 , \21681 );
not \U$21444 ( \21683 , \9478 );
and \U$21445 ( \21684 , \10206 , \10408 );
and \U$21446 ( \21685 , \10584 , \10116 );
nor \U$21447 ( \21686 , \21684 , \21685 );
xnor \U$21448 ( \21687 , \21686 , \10121 );
xor \U$21449 ( \21688 , \21683 , \21687 );
and \U$21450 ( \21689 , \9897 , \10118 );
xor \U$21451 ( \21690 , \21688 , \21689 );
xor \U$21452 ( \21691 , \21682 , \21690 );
and \U$21453 ( \21692 , \21647 , \21651 );
and \U$21454 ( \21693 , \21651 , \21667 );
and \U$21455 ( \21694 , \21647 , \21667 );
or \U$21456 ( \21695 , \21692 , \21693 , \21694 );
xor \U$21457 ( \21696 , \21691 , \21695 );
and \U$21458 ( \21697 , \21668 , \21669 );
and \U$21459 ( \21698 , \21670 , \21673 );
or \U$21460 ( \21699 , \21697 , \21698 );
xor \U$21461 ( \21700 , \21696 , \21699 );
buf g54a1_GF_PartitionCandidate( \21701_nG54a1 , \21700 );
buf \U$21462 ( \21702 , \21701_nG54a1 );
and \U$21463 ( \21703 , \21683 , \21687 );
and \U$21464 ( \21704 , \21687 , \21689 );
and \U$21465 ( \21705 , \21683 , \21689 );
or \U$21466 ( \21706 , \21703 , \21704 , \21705 );
and \U$21467 ( \21707 , \10584 , \10408 );
not \U$21468 ( \21708 , \21707 );
xnor \U$21469 ( \21709 , \21708 , \10121 );
and \U$21470 ( \21710 , \10206 , \10118 );
xnor \U$21471 ( \21711 , \21709 , \21710 );
xor \U$21472 ( \21712 , \21706 , \21711 );
and \U$21473 ( \21713 , \21680 , \21681 );
and \U$21474 ( \21714 , \21681 , \21690 );
and \U$21475 ( \21715 , \21680 , \21690 );
or \U$21476 ( \21716 , \21713 , \21714 , \21715 );
xor \U$21477 ( \21717 , \21712 , \21716 );
and \U$21478 ( \21718 , \21691 , \21695 );
and \U$21479 ( \21719 , \21696 , \21699 );
or \U$21480 ( \21720 , \21718 , \21719 );
xor \U$21481 ( \21721 , \21717 , \21720 );
buf g549f_GF_PartitionCandidate( \21722_nG549f , \21721 );
buf \U$21482 ( \21723 , \21722_nG549f );
or \U$21483 ( \21724 , \21709 , \21710 );
not \U$21484 ( \21725 , \10121 );
xor \U$21485 ( \21726 , \21724 , \21725 );
and \U$21486 ( \21727 , \10584 , \10118 );
xor \U$21487 ( \21728 , \21726 , \21727 );
and \U$21488 ( \21729 , \21706 , \21711 );
xor \U$21489 ( \21730 , \21728 , \21729 );
and \U$21490 ( \21731 , \21712 , \21716 );
and \U$21491 ( \21732 , \21717 , \21720 );
or \U$21492 ( \21733 , \21731 , \21732 );
xor \U$21493 ( \21734 , \21730 , \21733 );
buf g549d_GF_PartitionCandidate( \21735_nG549d , \21734 );
buf \U$21494 ( \21736 , \21735_nG549d );
xor \U$21495 ( \21737 , \649 , \1063 );
buf g557b_GF_PartitionCandidate( \21738_nG557b , \21737 );
buf \U$21496 ( \21739 , \21738_nG557b );
xor \U$21497 ( \21740 , \594 , \1065 );
buf g5579_GF_PartitionCandidate( \21741_nG5579 , \21740 );
buf \U$21498 ( \21742 , \21741_nG5579 );
xor \U$21499 ( \21743 , \865 , \1055 );
buf g5583_GF_PartitionCandidate( \21744_nG5583 , \21743 );
buf \U$21500 ( \21745 , \21744_nG5583 );
xor \U$21501 ( \21746 , \812 , \1057 );
buf g5581_GF_PartitionCandidate( \21747_nG5581 , \21746 );
buf \U$21502 ( \21748 , \21747_nG5581 );
xor \U$21503 ( \21749 , \773 , \1059 );
buf g557f_GF_PartitionCandidate( \21750_nG557f , \21749 );
buf \U$21504 ( \21751 , \21750_nG557f );
xor \U$21505 ( \21752 , \720 , \1061 );
buf g557d_GF_PartitionCandidate( \21753_nG557d , \21752 );
buf \U$21506 ( \21754 , \21753_nG557d );
xor \U$21507 ( \21755 , \907 , \1051 );
buf g5587_GF_PartitionCandidate( \21756_nG5587 , \21755 );
buf \U$21508 ( \21757 , \21756_nG5587 );
xor \U$21509 ( \21758 , \873 , \1053 );
buf g5585_GF_PartitionCandidate( \21759_nG5585 , \21758 );
buf \U$21510 ( \21760 , \21759_nG5585 );
xor \U$21511 ( \21761 , \941 , \1049 );
buf g5589_GF_PartitionCandidate( \21762_nG5589 , \21761 );
buf \U$21512 ( \21763 , \21762_nG5589 );
xor \U$21513 ( \21764 , \949 , \1047 );
buf g558b_GF_PartitionCandidate( \21765_nG558b , \21764 );
buf \U$21514 ( \21766 , \21765_nG558b );
xor \U$21515 ( \21767 , \994 , \1043 );
buf g558f_GF_PartitionCandidate( \21768_nG558f , \21767 );
buf \U$21516 ( \21769 , \21768_nG558f );
xor \U$21517 ( \21770 , \975 , \1045 );
buf g558d_GF_PartitionCandidate( \21771_nG558d , \21770 );
buf \U$21518 ( \21772 , \21771_nG558d );
xor \U$21519 ( \21773 , \1031 , \1034 );
buf g5599_GF_PartitionCandidate( \21774_nG5599 , \21773 );
buf \U$21520 ( \21775 , \21774_nG5599 );
xor \U$21521 ( \21776 , \1027 , \1035 );
buf g5597_GF_PartitionCandidate( \21777_nG5597 , \21776 );
buf \U$21522 ( \21778 , \21777_nG5597 );
xor \U$21523 ( \21779 , \1022 , \1037 );
buf g5595_GF_PartitionCandidate( \21780_nG5595 , \21779 );
buf \U$21524 ( \21781 , \21780_nG5595 );
xor \U$21525 ( \21782 , \1014 , \1039 );
buf g5593_GF_PartitionCandidate( \21783_nG5593 , \21782 );
buf \U$21526 ( \21784 , \21783_nG5593 );
xor \U$21527 ( \21785 , \1002 , \1041 );
buf g5591_GF_PartitionCandidate( \21786_nG5591 , \21785 );
buf \U$21528 ( \21787 , \21786_nG5591 );
xor \U$21529 ( \21788 , \1033 , \179 );
buf g559b_GF_PartitionCandidate( \21789_nG559b , \21788 );
buf \U$21530 ( \21790 , \21789_nG559b );
and \U$21531 ( \21791 , \21775 , \21778 , \21781 , \21784 , \21787 , \21790 );
or \U$21532 ( \21792 , \21769 , \21772 , \21791 );
and \U$21533 ( \21793 , \21766 , \21792 );
or \U$21534 ( \21794 , \21763 , \21793 );
and \U$21535 ( \21795 , \21757 , \21760 , \21794 );
or \U$21536 ( \21796 , \21745 , \21748 , \21751 , \21754 , \21795 );
and \U$21537 ( \21797 , \21739 , \21742 , \21796 );
or \U$21538 ( \21798 , \16027 , \16264 , \16499 , \16727 , \16951 , \17169 , \17382 , \17587 , \17790 , \17985 , \18178 , \18364 , \18545 , \18718 , \18888 , \19053 , \19216 , \19376 , \19531 , \19679 , \19822 , \19957 , \20091 , \20219 , \20342 , \20458 , \20568 , \20673 , \20776 , \20871 , \20964 , \21049 , \21132 , \21208 , \21279 , \21347 , \21410 , \21465 , \21518 , \21564 , \21605 , \21643 , \21676 , \21702 , \21723 , \21736 , \21797 );
or \U$21539 ( \21799 , \15782 , \21798 );
buf \U$21540 ( \21800 , \21799 );
buf \U$21541 ( \21801 , \1069_nG5577 );
buf \U$21542 ( \21802 , \1170_nG5575 );
buf \U$21543 ( \21803 , \1278_nG5573 );
buf \U$21544 ( \21804 , \1389_nG5571 );
buf \U$21545 ( \21805 , \1507_nG556f );
buf \U$21546 ( \21806 , \1628_nG556d );
buf \U$21547 ( \21807 , \1756_nG556b );
buf \U$21548 ( \21808 , \1887_nG5569 );
buf \U$21549 ( \21809 , \2025_nG5567 );
buf \U$21550 ( \21810 , \2166_nG5565 );
buf \U$21551 ( \21811 , \2314_nG5563 );
buf \U$21552 ( \21812 , \2465_nG5561 );
buf \U$21553 ( \21813 , \2623_nG555f );
buf \U$21554 ( \21814 , \2784_nG555d );
buf \U$21555 ( \21815 , \2952_nG555b );
buf \U$21556 ( \21816 , \3123_nG5559 );
buf \U$21557 ( \21817 , \3301_nG5557 );
buf \U$21558 ( \21818 , \3482_nG5555 );
buf \U$21559 ( \21819 , \3670_nG5553 );
buf \U$21560 ( \21820 , \3861_nG5551 );
buf \U$21561 ( \21821 , \4059_nG554f );
buf \U$21562 ( \21822 , \4260_nG554d );
buf \U$21563 ( \21823 , \4468_nG554b );
buf \U$21564 ( \21824 , \4679_nG5549 );
buf \U$21565 ( \21825 , \4897_nG5547 );
buf \U$21566 ( \21826 , \5117_nG5545 );
buf \U$21567 ( \21827 , \5348_nG5543 );
buf \U$21568 ( \21828 , \5579_nG5541 );
buf \U$21569 ( \21829 , \5817_nG553f );
buf \U$21570 ( \21830 , \6058_nG553d );
buf \U$21571 ( \21831 , \6306_nG553b );
buf \U$21572 ( \21832 , \6557_nG5539 );
buf \U$21573 ( \21833 , \6815_nG5537 );
buf \U$21574 ( \21834 , \7076_nG5535 );
buf \U$21575 ( \21835 , \7344_nG5533 );
buf \U$21576 ( \21836 , \7615_nG5531 );
buf \U$21577 ( \21837 , \7893_nG552f );
buf \U$21578 ( \21838 , \8174_nG552d );
buf \U$21579 ( \21839 , \8462_nG552b );
buf \U$21580 ( \21840 , \8753_nG5529 );
buf \U$21581 ( \21841 , \9051_nG5527 );
buf \U$21582 ( \21842 , \9352_nG5525 );
buf \U$21583 ( \21843 , \9660_nG5523 );
buf \U$21584 ( \21844 , \9971_nG5521 );
buf \U$21585 ( \21845 , \10289_nG551f );
buf \U$21586 ( \21846 , \10610_nG551d );
buf \U$21587 ( \21847 , \10929_nG551b );
buf \U$21588 ( \21848 , \11247_nG5519 );
buf \U$21589 ( \21849 , \11564_nG5517 );
buf \U$21590 ( \21850 , \11880_nG5515 );
buf \U$21591 ( \21851 , \12191_nG5513 );
buf \U$21592 ( \21852 , \12499_nG5511 );
buf \U$21593 ( \21853 , \12802_nG550f );
buf \U$21594 ( \21854 , \13098_nG550d );
buf \U$21595 ( \21855 , \13389_nG550b );
buf \U$21596 ( \21856 , \13672_nG5509 );
buf \U$21597 ( \21857 , \13953_nG5507 );
buf \U$21598 ( \21858 , \14226_nG5505 );
buf \U$21599 ( \21859 , \14496_nG5503 );
buf \U$21600 ( \21860 , \14762_nG5501 );
buf \U$21601 ( \21861 , \15022_nG54ff );
buf \U$21602 ( \21862 , \15277_nG54fd );
buf \U$21603 ( \21863 , \15530_nG54fb );
buf \U$21604 ( \21864 , \15780_nG54f9 );
or \U$21605 ( \21865 , \21801 , \21802 , \21803 , \21804 , \21805 , \21806 , \21807 , \21808 , \21809 , \21810 , \21811 , \21812 , \21813 , \21814 , \21815 , \21816 , \21817 , \21818 , \21819 , \21820 , \21821 , \21822 , \21823 , \21824 , \21825 , \21826 , \21827 , \21828 , \21829 , \21830 , \21831 , \21832 , \21833 , \21834 , \21835 , \21836 , \21837 , \21838 , \21839 , \21840 , \21841 , \21842 , \21843 , \21844 , \21845 , \21846 , \21847 , \21848 , \21849 , \21850 , \21851 , \21852 , \21853 , \21854 , \21855 , \21856 , \21857 , \21858 , \21859 , \21860 , \21861 , \21862 , \21863 , \21864 );
buf \U$21606 ( \21866 , \16026_nG54f7 );
buf \U$21607 ( \21867 , \16263_nG54f5 );
buf \U$21608 ( \21868 , \16498_nG54f3 );
buf \U$21609 ( \21869 , \16726_nG54f1 );
buf \U$21610 ( \21870 , \16950_nG54ef );
buf \U$21611 ( \21871 , \17168_nG54ed );
buf \U$21612 ( \21872 , \17381_nG54eb );
buf \U$21613 ( \21873 , \17586_nG54e9 );
buf \U$21614 ( \21874 , \17789_nG54e7 );
buf \U$21615 ( \21875 , \17984_nG54e5 );
buf \U$21616 ( \21876 , \18177_nG54e3 );
buf \U$21617 ( \21877 , \18363_nG54e1 );
buf \U$21618 ( \21878 , \18544_nG54df );
buf \U$21619 ( \21879 , \18717_nG54dd );
buf \U$21620 ( \21880 , \18887_nG54db );
buf \U$21621 ( \21881 , \19052_nG54d9 );
buf \U$21622 ( \21882 , \19215_nG54d7 );
buf \U$21623 ( \21883 , \19375_nG54d5 );
buf \U$21624 ( \21884 , \19530_nG54d3 );
buf \U$21625 ( \21885 , \19678_nG54d1 );
buf \U$21626 ( \21886 , \19821_nG54cf );
buf \U$21627 ( \21887 , \19956_nG54cd );
buf \U$21628 ( \21888 , \20090_nG54cb );
buf \U$21629 ( \21889 , \20218_nG54c9 );
buf \U$21630 ( \21890 , \20341_nG54c7 );
buf \U$21631 ( \21891 , \20457_nG54c5 );
buf \U$21632 ( \21892 , \20567_nG54c3 );
buf \U$21633 ( \21893 , \20672_nG54c1 );
buf \U$21634 ( \21894 , \20775_nG54bf );
buf \U$21635 ( \21895 , \20870_nG54bd );
buf \U$21636 ( \21896 , \20963_nG54bb );
buf \U$21637 ( \21897 , \21048_nG54b9 );
buf \U$21638 ( \21898 , \21131_nG54b7 );
buf \U$21639 ( \21899 , \21207_nG54b5 );
buf \U$21640 ( \21900 , \21278_nG54b3 );
buf \U$21641 ( \21901 , \21346_nG54b1 );
buf \U$21642 ( \21902 , \21409_nG54af );
buf \U$21643 ( \21903 , \21464_nG54ad );
buf \U$21644 ( \21904 , \21517_nG54ab );
buf \U$21645 ( \21905 , \21563_nG54a9 );
buf \U$21646 ( \21906 , \21604_nG54a7 );
buf \U$21647 ( \21907 , \21642_nG54a5 );
buf \U$21648 ( \21908 , \21675_nG54a3 );
buf \U$21649 ( \21909 , \21701_nG54a1 );
buf \U$21650 ( \21910 , \21722_nG549f );
buf \U$21651 ( \21911 , \21735_nG549d );
buf \U$21652 ( \21912 , \21738_nG557b );
buf \U$21653 ( \21913 , \21741_nG5579 );
buf \U$21654 ( \21914 , \21750_nG557f );
buf \U$21655 ( \21915 , \21753_nG557d );
buf \U$21656 ( \21916 , \21759_nG5585 );
buf \U$21657 ( \21917 , \21744_nG5583 );
buf \U$21658 ( \21918 , \21747_nG5581 );
buf \U$21659 ( \21919 , \21765_nG558b );
buf \U$21660 ( \21920 , \21762_nG5589 );
buf \U$21661 ( \21921 , \21756_nG5587 );
buf \U$21662 ( \21922 , \21771_nG558d );
buf \U$21663 ( \21923 , \21768_nG558f );
buf \U$21664 ( \21924 , \21786_nG5591 );
buf \U$21665 ( \21925 , \21780_nG5595 );
buf \U$21666 ( \21926 , \21783_nG5593 );
buf \U$21667 ( \21927 , \21789_nG559b );
buf \U$21668 ( \21928 , \21774_nG5599 );
buf \U$21669 ( \21929 , \21777_nG5597 );
and \U$21670 ( \21930 , \21927 , \21928 , \21929 );
or \U$21671 ( \21931 , \21925 , \21926 , \21930 );
and \U$21672 ( \21932 , \21924 , \21931 );
or \U$21673 ( \21933 , \21923 , \21932 );
and \U$21674 ( \21934 , \21922 , \21933 );
or \U$21675 ( \21935 , \21919 , \21920 , \21921 , \21934 );
and \U$21676 ( \21936 , \21916 , \21917 , \21918 , \21935 );
or \U$21677 ( \21937 , \21914 , \21915 , \21936 );
and \U$21678 ( \21938 , \21912 , \21913 , \21937 );
or \U$21679 ( \21939 , \21866 , \21867 , \21868 , \21869 , \21870 , \21871 , \21872 , \21873 , \21874 , \21875 , \21876 , \21877 , \21878 , \21879 , \21880 , \21881 , \21882 , \21883 , \21884 , \21885 , \21886 , \21887 , \21888 , \21889 , \21890 , \21891 , \21892 , \21893 , \21894 , \21895 , \21896 , \21897 , \21898 , \21899 , \21900 , \21901 , \21902 , \21903 , \21904 , \21905 , \21906 , \21907 , \21908 , \21909 , \21910 , \21911 , \21938 );
nor \U$21680 ( \21940 , \21865 , \21939 );
buf \U$21681 ( \21941 , \21940 );
and \U$21682 ( \21942 , \21800 , \21941 );
not \U$21683 ( \21943 , \21942 );
_DC g56b6 ( \21944_nG56b6 , 1'b0 , \21943 );
buf \U$21684 ( \21945 , \21944_nG56b6 );
endmodule

