//
// Conformal-LEC Version 20.10-d131 (29-Jun-2020)
//
module top(RIc0d85f0_34,RIc0d9478_65,RIc0d9658_69,RIc0d8398_29,RIc0d96d0_70,RIc0d9748_71,RIc0d8320_28,RIc0da288_95,RIc0d7768_3,
        RIc0da300_96,RIc0da378_97,RIc0d76f0_2,RIc0d9b08_79,RIc0d7ee8_19,RIc0d9b80_80,RIc0d9bf8_81,RIc0d7e70_18,RIc0d7a38_9,RIc0d9fb8_89,
        RIc0da030_90,RIc0da0a8_91,RIc0d79c0_8,RIc0d7858_5,RIc0da198_93,RIc0da210_94,RIc0d77e0_4,RIc0d7948_7,RIc0da120_92,RIc0d78d0_6,
        RIc0d7d08_15,RIc0d9ce8_83,RIc0d9d60_84,RIc0d9dd8_85,RIc0d7c90_14,RIc0d9f40_88,RIc0d9ec8_87,RIc0d7b28_11,RIc0d7ab0_10,RIc0d8578_33,
        RIc0d8410_30,RIc0d9568_67,RIc0d95e0_68,RIc0da3f0_98,RIc0da468_99,RIc0d98b0_74,RIc0d9928_75,RIc0d9838_73,RIc0d8140_24,RIc0d80c8_23,
        RIc0d82a8_27,RIc0d9e50_86,RIc0d7ba0_12,RIc0d7678_1,RIc0d7c18_13,RIc0d7df8_17,RIc0d7d80_16,RIc0d9c70_82,RIc0d8050_22,RIc0d99a0_76,
        RIc0d9a18_77,RIc0d7fd8_21,RIc0d7f60_20,RIc0d9a90_78,RIc0d8500_32,RIc0d94f0_66,RIc0d8488_31,RIc0d8230_26,RIc0d97c0_72,RIc0d81b8_25,
        RIc0d8668_35,RIc0da4e0_100,RIc0da558_101,RIc0d86e0_36,RIc0d8758_37,RIc0da5d0_102,RIc0da648_103,RIc0d87d0_38,RIc0d8848_39,RIc0da6c0_104,
        RIc0da738_105,RIc0d8b90_46,RIc0d8b18_45,RIc0dabe8_115,RIc0dac60_116,RIc0dacd8_117,RIc0da828_107,RIc0da8a0_108,RIc0da918_109,RIc0d8d70_50,
        RIc0d8cf8_49,RIc0daaf8_113,RIc0dab70_114,RIc0d9040_56,RIc0d8fc8_55,RIc0d9220_60,RIc0d91a8_59,RIc0d8aa0_44,RIc0d8a28_43,RIc0daa08_111,
        RIc0daa80_112,RIc0d89b0_42,RIc0d8938_41,RIc0db188_127,RIc0db200_128,RIc0d9130_58,RIc0d90b8_57,RIc0da7b0_106,RIc0d8e60_52,RIc0d8de8_51,
        RIc0d9400_64,RIc0d9388_63,RIc0dafa8_123,RIc0db020_124,RIc0db098_125,RIc0dad50_118,RIc0dadc8_119,RIc0daeb8_121,RIc0daf30_122,RIc0dae40_120,
        RIc0d8c80_48,RIc0d8c08_47,RIc0d9310_62,RIc0d9298_61,RIc0d8f50_54,RIc0d8ed8_53,RIc0da990_110,RIc0db110_126,RIc0d88c0_40,R_81_84446b8,
        R_82_8444760,R_83_8444808,R_84_84448b0,R_85_8444958,R_86_8444a00,R_87_9bec6f8,R_88_9bec7a0,R_89_9bec848,R_8a_9bec8f0,R_8b_9bec998,
        R_8c_9beca40,R_8d_9becae8,R_8e_9becb90,R_8f_9becc38,R_90_9becce0,R_91_9becd88,R_92_9bece30,R_93_9beced8,R_94_9becf80,R_95_9bed028,
        R_96_9bed0d0,R_97_9bed178,R_98_9bed220,R_99_9bed2c8,R_9a_9bed370,R_9b_9bed418,R_9c_9bed4c0,R_9d_9bed568,R_9e_9bed610,R_9f_9bed6b8,
        R_a0_9bed760,R_a1_9bed808,R_a2_9bed8b0,R_a3_9bed958,R_a4_9beda00,R_a5_9bedaa8,R_a6_9bedb50,R_a7_9bedbf8,R_a8_9bedca0,R_a9_9bedd48,
        R_aa_9beddf0,R_ab_9bede98,R_ac_9bedf40,R_ad_9bedfe8,R_ae_9bee090,R_af_9bee138,R_b0_9bee1e0,R_b1_9bee288,R_b2_9bee330,R_b3_9bee3d8,
        R_b4_9bee480,R_b5_9bee528,R_b6_9bee5d0,R_b7_9bee678,R_b8_9bee720,R_b9_9bee7c8,R_ba_9bee870,R_bb_9bee918,R_bc_9bee9c0,R_bd_9beea68,
        R_be_9beeb10,R_bf_9beebb8,R_c0_9beec60,R_c1_9beed08,R_c2_9beedb0,R_c3_9beee58,R_c4_9beef00,R_c5_9beefa8,R_c6_9bef050,R_c7_9bef0f8,
        R_c8_9bef1a0,R_c9_9bef248,R_ca_9bef2f0,R_cb_9bef398,R_cc_9bef440,R_cd_9bef4e8,R_ce_9bef590,R_cf_9bef638,R_d0_9bef6e0,R_d1_9bef788,
        R_d2_9bef830,R_d3_9bef8d8,R_d4_9bef980,R_d5_9befa28,R_d6_9befad0,R_d7_9befb78,R_d8_9befc20,R_d9_9befcc8,R_da_9befd70,R_db_9befe18,
        R_dc_9befec0,R_dd_9beff68,R_de_9bf0010,R_df_9bf00b8,R_e0_9bf0160,R_e1_9bf0208,R_e2_9bf02b0,R_e3_9bf0358,R_e4_9bf0400,R_e5_9bf04a8,
        R_e6_9bf0550,R_e7_9bf05f8,R_e8_9bf06a0,R_e9_9bf0748,R_ea_9bf07f0,R_eb_9bf0898,R_ec_9bf0940,R_ed_9bf09e8,R_ee_9bf0a90,R_ef_9bf0b38,
        R_f0_9bf0be0,R_f1_9bf0c88,R_f2_9bf0d30,R_f3_9bf0dd8);
input RIc0d85f0_34,RIc0d9478_65,RIc0d9658_69,RIc0d8398_29,RIc0d96d0_70,RIc0d9748_71,RIc0d8320_28,RIc0da288_95,RIc0d7768_3,
        RIc0da300_96,RIc0da378_97,RIc0d76f0_2,RIc0d9b08_79,RIc0d7ee8_19,RIc0d9b80_80,RIc0d9bf8_81,RIc0d7e70_18,RIc0d7a38_9,RIc0d9fb8_89,
        RIc0da030_90,RIc0da0a8_91,RIc0d79c0_8,RIc0d7858_5,RIc0da198_93,RIc0da210_94,RIc0d77e0_4,RIc0d7948_7,RIc0da120_92,RIc0d78d0_6,
        RIc0d7d08_15,RIc0d9ce8_83,RIc0d9d60_84,RIc0d9dd8_85,RIc0d7c90_14,RIc0d9f40_88,RIc0d9ec8_87,RIc0d7b28_11,RIc0d7ab0_10,RIc0d8578_33,
        RIc0d8410_30,RIc0d9568_67,RIc0d95e0_68,RIc0da3f0_98,RIc0da468_99,RIc0d98b0_74,RIc0d9928_75,RIc0d9838_73,RIc0d8140_24,RIc0d80c8_23,
        RIc0d82a8_27,RIc0d9e50_86,RIc0d7ba0_12,RIc0d7678_1,RIc0d7c18_13,RIc0d7df8_17,RIc0d7d80_16,RIc0d9c70_82,RIc0d8050_22,RIc0d99a0_76,
        RIc0d9a18_77,RIc0d7fd8_21,RIc0d7f60_20,RIc0d9a90_78,RIc0d8500_32,RIc0d94f0_66,RIc0d8488_31,RIc0d8230_26,RIc0d97c0_72,RIc0d81b8_25,
        RIc0d8668_35,RIc0da4e0_100,RIc0da558_101,RIc0d86e0_36,RIc0d8758_37,RIc0da5d0_102,RIc0da648_103,RIc0d87d0_38,RIc0d8848_39,RIc0da6c0_104,
        RIc0da738_105,RIc0d8b90_46,RIc0d8b18_45,RIc0dabe8_115,RIc0dac60_116,RIc0dacd8_117,RIc0da828_107,RIc0da8a0_108,RIc0da918_109,RIc0d8d70_50,
        RIc0d8cf8_49,RIc0daaf8_113,RIc0dab70_114,RIc0d9040_56,RIc0d8fc8_55,RIc0d9220_60,RIc0d91a8_59,RIc0d8aa0_44,RIc0d8a28_43,RIc0daa08_111,
        RIc0daa80_112,RIc0d89b0_42,RIc0d8938_41,RIc0db188_127,RIc0db200_128,RIc0d9130_58,RIc0d90b8_57,RIc0da7b0_106,RIc0d8e60_52,RIc0d8de8_51,
        RIc0d9400_64,RIc0d9388_63,RIc0dafa8_123,RIc0db020_124,RIc0db098_125,RIc0dad50_118,RIc0dadc8_119,RIc0daeb8_121,RIc0daf30_122,RIc0dae40_120,
        RIc0d8c80_48,RIc0d8c08_47,RIc0d9310_62,RIc0d9298_61,RIc0d8f50_54,RIc0d8ed8_53,RIc0da990_110,RIc0db110_126,RIc0d88c0_40;
output R_81_84446b8,R_82_8444760,R_83_8444808,R_84_84448b0,R_85_8444958,R_86_8444a00,R_87_9bec6f8,R_88_9bec7a0,R_89_9bec848,
        R_8a_9bec8f0,R_8b_9bec998,R_8c_9beca40,R_8d_9becae8,R_8e_9becb90,R_8f_9becc38,R_90_9becce0,R_91_9becd88,R_92_9bece30,R_93_9beced8,
        R_94_9becf80,R_95_9bed028,R_96_9bed0d0,R_97_9bed178,R_98_9bed220,R_99_9bed2c8,R_9a_9bed370,R_9b_9bed418,R_9c_9bed4c0,R_9d_9bed568,
        R_9e_9bed610,R_9f_9bed6b8,R_a0_9bed760,R_a1_9bed808,R_a2_9bed8b0,R_a3_9bed958,R_a4_9beda00,R_a5_9bedaa8,R_a6_9bedb50,R_a7_9bedbf8,
        R_a8_9bedca0,R_a9_9bedd48,R_aa_9beddf0,R_ab_9bede98,R_ac_9bedf40,R_ad_9bedfe8,R_ae_9bee090,R_af_9bee138,R_b0_9bee1e0,R_b1_9bee288,
        R_b2_9bee330,R_b3_9bee3d8,R_b4_9bee480,R_b5_9bee528,R_b6_9bee5d0,R_b7_9bee678,R_b8_9bee720,R_b9_9bee7c8,R_ba_9bee870,R_bb_9bee918,
        R_bc_9bee9c0,R_bd_9beea68,R_be_9beeb10,R_bf_9beebb8,R_c0_9beec60,R_c1_9beed08,R_c2_9beedb0,R_c3_9beee58,R_c4_9beef00,R_c5_9beefa8,
        R_c6_9bef050,R_c7_9bef0f8,R_c8_9bef1a0,R_c9_9bef248,R_ca_9bef2f0,R_cb_9bef398,R_cc_9bef440,R_cd_9bef4e8,R_ce_9bef590,R_cf_9bef638,
        R_d0_9bef6e0,R_d1_9bef788,R_d2_9bef830,R_d3_9bef8d8,R_d4_9bef980,R_d5_9befa28,R_d6_9befad0,R_d7_9befb78,R_d8_9befc20,R_d9_9befcc8,
        R_da_9befd70,R_db_9befe18,R_dc_9befec0,R_dd_9beff68,R_de_9bf0010,R_df_9bf00b8,R_e0_9bf0160,R_e1_9bf0208,R_e2_9bf02b0,R_e3_9bf0358,
        R_e4_9bf0400,R_e5_9bf04a8,R_e6_9bf0550,R_e7_9bf05f8,R_e8_9bf06a0,R_e9_9bf0748,R_ea_9bf07f0,R_eb_9bf0898,R_ec_9bf0940,R_ed_9bf09e8,
        R_ee_9bf0a90,R_ef_9bf0b38,R_f0_9bf0be0,R_f1_9bf0c88,R_f2_9bf0d30,R_f3_9bf0dd8;

wire \244_ZERO , \245_ONE , \246 , \247 , \248 , \249 , \250 , \251 , \252 ,
         \253 , \254 , \255 , \256 , \257 , \258 , \259 , \260 , \261 , \262 ,
         \263 , \264 , \265 , \266 , \267 , \268 , \269 , \270 , \271 , \272 ,
         \273 , \274 , \275 , \276 , \277 , \278 , \279 , \280 , \281 , \282 ,
         \283 , \284 , \285 , \286 , \287 , \288 , \289 , \290 , \291 , \292 ,
         \293 , \294 , \295 , \296 , \297 , \298 , \299 , \300 , \301 , \302 ,
         \303 , \304 , \305 , \306 , \307 , \308 , \309 , \310 , \311 , \312 ,
         \313 , \314 , \315 , \316 , \317 , \318 , \319 , \320 , \321 , \322 ,
         \323 , \324 , \325 , \326 , \327 , \328 , \329 , \330 , \331 , \332 ,
         \333 , \334 , \335 , \336 , \337 , \338 , \339 , \340 , \341 , \342 ,
         \343 , \344 , \345 , \346 , \347 , \348 , \349 , \350 , \351 , \352 ,
         \353 , \354 , \355 , \356 , \357 , \358 , \359 , \360 , \361 , \362 ,
         \363 , \364 , \365 , \366 , \367 , \368 , \369 , \370 , \371 , \372 ,
         \373 , \374 , \375 , \376 , \377 , \378 , \379 , \380 , \381 , \382 ,
         \383 , \384 , \385 , \386 , \387 , \388 , \389 , \390 , \391 , \392 ,
         \393 , \394 , \395 , \396 , \397 , \398 , \399 , \400 , \401 , \402 ,
         \403 , \404 , \405 , \406 , \407 , \408 , \409 , \410 , \411 , \412 ,
         \413 , \414 , \415 , \416 , \417 , \418 , \419 , \420 , \421 , \422 ,
         \423 , \424 , \425 , \426 , \427 , \428 , \429 , \430 , \431 , \432 ,
         \433 , \434 , \435 , \436 , \437 , \438 , \439 , \440 , \441 , \442 ,
         \443 , \444 , \445 , \446 , \447 , \448 , \449 , \450 , \451 , \452 ,
         \453 , \454 , \455 , \456 , \457 , \458 , \459 , \460 , \461 , \462 ,
         \463 , \464 , \465 , \466 , \467 , \468 , \469 , \470 , \471 , \472 ,
         \473 , \474 , \475 , \476 , \477 , \478 , \479 , \480 , \481 , \482 ,
         \483 , \484 , \485 , \486 , \487 , \488 , \489 , \490 , \491 , \492 ,
         \493 , \494 , \495 , \496 , \497 , \498 , \499 , \500 , \501 , \502 ,
         \503 , \504 , \505 , \506 , \507 , \508 , \509 , \510 , \511 , \512 ,
         \513 , \514 , \515 , \516 , \517 , \518 , \519 , \520 , \521 , \522 ,
         \523 , \524 , \525 , \526 , \527 , \528 , \529 , \530 , \531 , \532 ,
         \533 , \534 , \535 , \536 , \537 , \538 , \539 , \540 , \541 , \542 ,
         \543 , \544 , \545 , \546 , \547 , \548 , \549 , \550 , \551 , \552 ,
         \553 , \554 , \555 , \556 , \557 , \558 , \559 , \560 , \561 , \562 ,
         \563 , \564 , \565 , \566 , \567 , \568 , \569 , \570 , \571 , \572 ,
         \573 , \574 , \575 , \576 , \577 , \578 , \579 , \580 , \581 , \582 ,
         \583 , \584 , \585 , \586 , \587 , \588 , \589 , \590 , \591 , \592 ,
         \593 , \594 , \595 , \596 , \597 , \598 , \599 , \600 , \601 , \602 ,
         \603 , \604 , \605 , \606 , \607 , \608 , \609 , \610 , \611 , \612 ,
         \613 , \614 , \615 , \616 , \617 , \618 , \619 , \620 , \621 , \622 ,
         \623 , \624 , \625 , \626 , \627 , \628 , \629 , \630 , \631 , \632 ,
         \633 , \634 , \635 , \636 , \637 , \638 , \639 , \640 , \641 , \642 ,
         \643 , \644 , \645 , \646 , \647 , \648 , \649 , \650 , \651 , \652 ,
         \653 , \654 , \655 , \656 , \657 , \658 , \659 , \660 , \661 , \662 ,
         \663 , \664 , \665 , \666 , \667 , \668 , \669 , \670 , \671 , \672 ,
         \673 , \674 , \675 , \676 , \677 , \678 , \679 , \680 , \681 , \682 ,
         \683 , \684 , \685 , \686 , \687 , \688 , \689 , \690 , \691 , \692 ,
         \693 , \694 , \695 , \696 , \697 , \698 , \699 , \700 , \701 , \702 ,
         \703 , \704 , \705 , \706 , \707 , \708 , \709 , \710 , \711 , \712 ,
         \713 , \714 , \715 , \716 , \717 , \718 , \719 , \720 , \721 , \722 ,
         \723 , \724 , \725 , \726 , \727 , \728 , \729 , \730 , \731 , \732 ,
         \733 , \734 , \735 , \736 , \737 , \738 , \739 , \740 , \741 , \742 ,
         \743 , \744 , \745 , \746 , \747 , \748 , \749 , \750 , \751 , \752 ,
         \753 , \754 , \755 , \756 , \757 , \758 , \759 , \760 , \761 , \762 ,
         \763 , \764 , \765 , \766 , \767 , \768 , \769 , \770 , \771 , \772 ,
         \773 , \774 , \775 , \776 , \777 , \778 , \779 , \780 , \781 , \782 ,
         \783 , \784 , \785 , \786 , \787 , \788 , \789 , \790 , \791 , \792 ,
         \793 , \794 , \795 , \796 , \797 , \798 , \799 , \800 , \801 , \802 ,
         \803 , \804 , \805 , \806 , \807 , \808 , \809 , \810 , \811 , \812 ,
         \813 , \814 , \815 , \816 , \817 , \818 , \819 , \820 , \821 , \822 ,
         \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 , \831 , \832 ,
         \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 , \841 , \842 ,
         \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 , \851 , \852 ,
         \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 , \861 , \862 ,
         \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 , \871 , \872 ,
         \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 , \881 , \882 ,
         \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 , \891 , \892 ,
         \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 , \901 , \902 ,
         \903 , \904 , \905 , \906 , \907 , \908 , \909 , \910 , \911 , \912 ,
         \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 , \921 , \922 ,
         \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 , \931 , \932 ,
         \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 ,
         \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 , \951 , \952 ,
         \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 , \961 , \962 ,
         \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 ,
         \973 , \974 , \975 , \976 , \977 , \978 , \979 , \980 , \981 , \982 ,
         \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 ,
         \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 ,
         \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 ,
         \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 ,
         \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 ,
         \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 ,
         \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 ,
         \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 ,
         \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 ,
         \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 ,
         \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 ,
         \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 ,
         \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 ,
         \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 ,
         \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 ,
         \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 ,
         \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 ,
         \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 ,
         \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 ,
         \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 ,
         \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 ,
         \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 ,
         \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 ,
         \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 ,
         \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 ,
         \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 ,
         \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 ,
         \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 ,
         \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 ,
         \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 ,
         \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 ,
         \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 ,
         \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 ,
         \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 ,
         \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 ,
         \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 ,
         \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 ,
         \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 ,
         \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 ,
         \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 ,
         \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 ,
         \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 ,
         \1403 , \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 ,
         \1413 , \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 ,
         \1423 , \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 ,
         \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 ,
         \1443 , \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 ,
         \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 ,
         \1463 , \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 ,
         \1473 , \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 ,
         \1483 , \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 ,
         \1493 , \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 ,
         \1503 , \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 ,
         \1513 , \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 ,
         \1523 , \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 ,
         \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 ,
         \1543 , \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 ,
         \1553 , \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 ,
         \1563 , \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 ,
         \1573 , \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 ,
         \1583 , \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 ,
         \1593 , \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 ,
         \1603 , \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 ,
         \1613 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 ,
         \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 ,
         \1633 , \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 ,
         \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 ,
         \1653 , \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 ,
         \1663 , \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 ,
         \1673 , \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 ,
         \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 ,
         \1693 , \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 ,
         \1703 , \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 ,
         \1713 , \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 ,
         \1723 , \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 ,
         \1733 , \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 ,
         \1743 , \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 ,
         \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 ,
         \1763 , \1764 , \1765 , \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 ,
         \1773 , \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 ,
         \1783 , \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 ,
         \1793 , \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 ,
         \1803 , \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 ,
         \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 ,
         \1823 , \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 ,
         \1833 , \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 ,
         \1843 , \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 ,
         \1853 , \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 ,
         \1863 , \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 ,
         \1873 , \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 ,
         \1883 , \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 ,
         \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 ,
         \1903 , \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 ,
         \1913 , \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 ,
         \1923 , \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 ,
         \1933 , \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 ,
         \1943 , \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 ,
         \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 ,
         \1963 , \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 ,
         \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 ,
         \1983 , \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 ,
         \1993 , \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 ,
         \2003 , \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 ,
         \2013 , \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 ,
         \2023 , \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 ,
         \2033 , \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 ,
         \2043 , \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 ,
         \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 ,
         \2063 , \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 ,
         \2073 , \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 ,
         \2083 , \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 ,
         \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 ,
         \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 ,
         \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 ,
         \2123 , \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 ,
         \2133 , \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 ,
         \2143 , \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 ,
         \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 ,
         \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 ,
         \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 ,
         \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 ,
         \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 ,
         \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 ,
         \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 ,
         \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 ,
         \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 ,
         \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 ,
         \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 ,
         \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 ,
         \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 ,
         \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 ,
         \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 ,
         \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 ,
         \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 ,
         \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 ,
         \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 ,
         \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 ,
         \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 ,
         \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 ,
         \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 ,
         \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 ,
         \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 ,
         \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 ,
         \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 ,
         \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 ,
         \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 ,
         \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 ,
         \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 ,
         \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 ,
         \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 ,
         \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 ,
         \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 ,
         \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 ,
         \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 ,
         \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 ,
         \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 ,
         \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 ,
         \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 ,
         \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 ,
         \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 ,
         \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 ,
         \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 ,
         \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 ,
         \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 ,
         \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 ,
         \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 ,
         \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 ,
         \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 ,
         \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 ,
         \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 ,
         \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 ,
         \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 ,
         \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 ,
         \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 ,
         \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 ,
         \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 ,
         \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 ,
         \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 ,
         \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 ,
         \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 ,
         \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 ,
         \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 ,
         \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 ,
         \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 ,
         \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 ,
         \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 ,
         \2843 , \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 ,
         \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 ,
         \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 ,
         \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 ,
         \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 ,
         \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 ,
         \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 ,
         \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 ,
         \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 ,
         \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 ,
         \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 ,
         \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 ,
         \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 ,
         \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 ,
         \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 ,
         \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 ,
         \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 ,
         \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 ,
         \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 ,
         \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 ,
         \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 ,
         \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 ,
         \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 ,
         \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 ,
         \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 ,
         \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 ,
         \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 ,
         \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 ,
         \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 ,
         \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 ,
         \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 ,
         \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 ,
         \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 ,
         \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 ,
         \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 ,
         \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 ,
         \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 ,
         \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 ,
         \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 ,
         \3233 , \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 ,
         \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 ,
         \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 ,
         \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 ,
         \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 ,
         \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 ,
         \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 ,
         \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 ,
         \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 ,
         \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 ,
         \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 ,
         \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 ,
         \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 ,
         \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 ,
         \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 ,
         \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 ,
         \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 ,
         \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 ,
         \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 ,
         \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 ,
         \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 ,
         \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 ,
         \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 ,
         \3463 , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 ,
         \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 ,
         \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 ,
         \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 ,
         \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 ,
         \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 ,
         \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 ,
         \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 ,
         \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 ,
         \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 ,
         \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 ,
         \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 ,
         \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 ,
         \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 ,
         \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 ,
         \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 ,
         \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 ,
         \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 ,
         \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 ,
         \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 ,
         \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 ,
         \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 ,
         \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 ,
         \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 ,
         \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 ,
         \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 ,
         \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 ,
         \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 ,
         \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 ,
         \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 ,
         \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 ,
         \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 ,
         \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 ,
         \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 ,
         \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 ,
         \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 ,
         \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 ,
         \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 ,
         \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 ,
         \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 ,
         \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 ,
         \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 ,
         \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 ,
         \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 ,
         \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 ,
         \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 ,
         \3923 , \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 ,
         \3933 , \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 ,
         \3943 , \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 ,
         \3953 , \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 ,
         \3963 , \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 ,
         \3973 , \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 ,
         \3983 , \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 ,
         \3993 , \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 ,
         \4003 , \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 ,
         \4013 , \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 ,
         \4023 , \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 ,
         \4033 , \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 ,
         \4043 , \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 ,
         \4053 , \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 ,
         \4063 , \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 ,
         \4073 , \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 ,
         \4083 , \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 ,
         \4093 , \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 ,
         \4103 , \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 ,
         \4113 , \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 ,
         \4123 , \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 ,
         \4133 , \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 ,
         \4143 , \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 ,
         \4153 , \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 ,
         \4163 , \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 ,
         \4173 , \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 ,
         \4183 , \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 ,
         \4193 , \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 ,
         \4203 , \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 ,
         \4213 , \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 ,
         \4223 , \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 ,
         \4233 , \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 ,
         \4243 , \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 ,
         \4253 , \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 ,
         \4263 , \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 ,
         \4273 , \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 ,
         \4283 , \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 ,
         \4293 , \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 ,
         \4303 , \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 ,
         \4313 , \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 ,
         \4323 , \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 ,
         \4333 , \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 ,
         \4343 , \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 ,
         \4353 , \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 ,
         \4363 , \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 ,
         \4373 , \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 ,
         \4383 , \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 ,
         \4393 , \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 ,
         \4403 , \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 ,
         \4413 , \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 ,
         \4423 , \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 ,
         \4433 , \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 ,
         \4443 , \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 ,
         \4453 , \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 ,
         \4463 , \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 ,
         \4473 , \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 ,
         \4483 , \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 ,
         \4493 , \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 ,
         \4503 , \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 ,
         \4513 , \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 ,
         \4523 , \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 ,
         \4533 , \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 ,
         \4543 , \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 ,
         \4553 , \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 ,
         \4563 , \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 ,
         \4573 , \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 ,
         \4583 , \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 ,
         \4593 , \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 ,
         \4603 , \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 ,
         \4613 , \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 ,
         \4623 , \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 ,
         \4633 , \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 ,
         \4643 , \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 ,
         \4653 , \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 ,
         \4663 , \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 ,
         \4673 , \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 ,
         \4683 , \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 ,
         \4693 , \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 ,
         \4703 , \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 ,
         \4713 , \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 ,
         \4723 , \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 ,
         \4733 , \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 ,
         \4743 , \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 ,
         \4753 , \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 ,
         \4763 , \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 ,
         \4773 , \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 ,
         \4783 , \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 ,
         \4793 , \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 ,
         \4803 , \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 ,
         \4813 , \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 ,
         \4823 , \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 ,
         \4833 , \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 ,
         \4843 , \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 ,
         \4853 , \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 ,
         \4863 , \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 ,
         \4873 , \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 ,
         \4883 , \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 ,
         \4893 , \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 ,
         \4903 , \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 ,
         \4913 , \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 ,
         \4923 , \4924 , \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 ,
         \4933 , \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 ,
         \4943 , \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 ,
         \4953 , \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 ,
         \4963 , \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 ,
         \4973 , \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 ,
         \4983 , \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 ,
         \4993 , \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 ,
         \5003 , \5004 , \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 ,
         \5013 , \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 ,
         \5023 , \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 ,
         \5033 , \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 ,
         \5043 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 ,
         \5053 , \5054 , \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 ,
         \5063 , \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 ,
         \5073 , \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 ,
         \5083 , \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 ,
         \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 ,
         \5103 , \5104 , \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 ,
         \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 ,
         \5123 , \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 ,
         \5133 , \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 ,
         \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 ,
         \5153 , \5154 , \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 ,
         \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 ,
         \5173 , \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 ,
         \5183 , \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 ,
         \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 ,
         \5203 , \5204 , \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 ,
         \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 ,
         \5223 , \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 ,
         \5233 , \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 ,
         \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 ,
         \5253 , \5254 , \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 ,
         \5263 , \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 ,
         \5273 , \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 ,
         \5283 , \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 ,
         \5293 , \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 ,
         \5303 , \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 ,
         \5313 , \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 ,
         \5323 , \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 ,
         \5333 , \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 ,
         \5343 , \5344 , \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 ,
         \5353 , \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 ,
         \5363 , \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 ,
         \5373 , \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 ,
         \5383 , \5384 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 ,
         \5393 , \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 ,
         \5403 , \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 ,
         \5413 , \5414 , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 ,
         \5423 , \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 ,
         \5433 , \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 ,
         \5443 , \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 ,
         \5453 , \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 ,
         \5463 , \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 ,
         \5473 , \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 ,
         \5483 , \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 ,
         \5493 , \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 ,
         \5503 , \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 ,
         \5513 , \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 ,
         \5523 , \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 ,
         \5533 , \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 ,
         \5543 , \5544 , \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 ,
         \5553 , \5554 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 ,
         \5563 , \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 ,
         \5573 , \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 ,
         \5583 , \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 ,
         \5593 , \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 ,
         \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 ,
         \5613 , \5614 , \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 ,
         \5623 , \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 ,
         \5633 , \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 ,
         \5643 , \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 ,
         \5653 , \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 ,
         \5663 , \5664 , \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 ,
         \5673 , \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 ,
         \5683 , \5684 , \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 ,
         \5693 , \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 ,
         \5703 , \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 ,
         \5713 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 ,
         \5723 , \5724 , \5725 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 , \5732 ,
         \5733 , \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 ,
         \5743 , \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 ,
         \5753 , \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 ,
         \5763 , \5764 , \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 ,
         \5773 , \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 ,
         \5783 , \5784 , \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 ,
         \5793 , \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 , \5802 ,
         \5803 , \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 ,
         \5813 , \5814 , \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821 , \5822 ,
         \5823 , \5824 , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 ,
         \5833 , \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 ,
         \5843 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 ,
         \5853 , \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 ,
         \5863 , \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 ,
         \5873 , \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 ,
         \5883 , \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 ,
         \5893 , \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 ,
         \5903 , \5904 , \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 ,
         \5913 , \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 ,
         \5923 , \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 ,
         \5933 , \5934 , \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 ,
         \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 ,
         \5953 , \5954 , \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 ,
         \5963 , \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 ,
         \5973 , \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 ,
         \5983 , \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 ,
         \5993 , \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 ,
         \6003 , \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 ,
         \6013 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 ,
         \6023 , \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 ,
         \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 ,
         \6043 , \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 ,
         \6053 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 ,
         \6063 , \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 ,
         \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 ,
         \6083 , \6084 , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 ,
         \6093 , \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 ,
         \6103 , \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 ,
         \6113 , \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 ,
         \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 ,
         \6133 , \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 ,
         \6143 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 ,
         \6153 , \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 ,
         \6163 , \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 ,
         \6173 , \6174 , \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 ,
         \6183 , \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 ,
         \6193 , \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 ,
         \6203 , \6204 , \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 ,
         \6213 , \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 ,
         \6223 , \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 ,
         \6233 , \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 ,
         \6243 , \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 ,
         \6253 , \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 ,
         \6263 , \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 ,
         \6273 , \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 ,
         \6283 , \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 ,
         \6293 , \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 ,
         \6303 , \6304 , \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 ,
         \6313 , \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 ,
         \6323 , \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 ,
         \6333 , \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 ,
         \6343 , \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 ,
         \6353 , \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 ,
         \6363 , \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 ,
         \6373 , \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 ,
         \6383 , \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 ,
         \6393 , \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 ,
         \6403 , \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 ,
         \6413 , \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 ,
         \6423 , \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 ,
         \6433 , \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 ,
         \6443 , \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 ,
         \6453 , \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 ,
         \6463 , \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 ,
         \6473 , \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 ,
         \6483 , \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 ,
         \6493 , \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 ,
         \6503 , \6504 , \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 ,
         \6513 , \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 ,
         \6523 , \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 ,
         \6533 , \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 ,
         \6543 , \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 ,
         \6553 , \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 ,
         \6563 , \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 ,
         \6573 , \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 ,
         \6583 , \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 ,
         \6593 , \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 ,
         \6603 , \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 ,
         \6613 , \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 ,
         \6623 , \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 ,
         \6633 , \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 ,
         \6643 , \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 ,
         \6653 , \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 ,
         \6663 , \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 ,
         \6673 , \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 ,
         \6683 , \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 ,
         \6693 , \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 ,
         \6703 , \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 ,
         \6713 , \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 ,
         \6723 , \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 ,
         \6733 , \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 ,
         \6743 , \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 ,
         \6753 , \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 ,
         \6763 , \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 ,
         \6773 , \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 ,
         \6783 , \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 ,
         \6793 , \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 ,
         \6803 , \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 ,
         \6813 , \6814 , \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 ,
         \6823 , \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 ,
         \6833 , \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 ,
         \6843 , \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 ,
         \6853 , \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 ,
         \6863 , \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 ,
         \6873 , \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 ,
         \6883 , \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 ,
         \6893 , \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 ,
         \6903 , \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 ,
         \6913 , \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 ,
         \6923 , \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 ,
         \6933 , \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 ,
         \6943 , \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 ,
         \6953 , \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 ,
         \6963 , \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 ,
         \6973 , \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 ,
         \6983 , \6984 , \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 ,
         \6993 , \6994 , \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 ,
         \7003 , \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 ,
         \7013 , \7014 , \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 ,
         \7023 , \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 ,
         \7033 , \7034 , \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 ,
         \7043 , \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 ,
         \7053 , \7054 , \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 ,
         \7063 , \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 ,
         \7073 , \7074 , \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 ,
         \7083 , \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 ,
         \7093 , \7094 , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 ,
         \7103 , \7104 , \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 ,
         \7113 , \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 ,
         \7123 , \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132 ,
         \7133 , \7134 , \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 ,
         \7143 , \7144 , \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 , \7152 ,
         \7153 , \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 ,
         \7163 , \7164 , \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172 ,
         \7173 , \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 ,
         \7183 , \7184 , \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 ,
         \7193 , \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 ,
         \7203 , \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 ,
         \7213 , \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222 ,
         \7223 , \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232 ,
         \7233 , \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242 ,
         \7243 , \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252 ,
         \7253 , \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262 ,
         \7263 , \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272 ,
         \7273 , \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 , \7282 ,
         \7283 , \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 ,
         \7293 , \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 ,
         \7303 , \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 ,
         \7313 , \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 , \7322 ,
         \7323 , \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 ,
         \7333 , \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 ,
         \7343 , \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 , \7352 ,
         \7353 , \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 ,
         \7363 , \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 ,
         \7373 , \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 , \7382 ,
         \7383 , \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 ,
         \7393 , \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 ,
         \7403 , \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 ,
         \7413 , \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 ,
         \7423 , \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 , \7432 ,
         \7433 , \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 , \7442 ,
         \7443 , \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 , \7452 ,
         \7453 , \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 , \7462 ,
         \7463 , \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 , \7472 ,
         \7473 , \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 , \7482 ,
         \7483 , \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 , \7492 ,
         \7493 , \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 , \7502 ,
         \7503 , \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 , \7512 ,
         \7513 , \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 , \7522 ,
         \7523 , \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 , \7532 ,
         \7533 , \7534 , \7535 , \7536 , \7537 , \7538 , \7539 , \7540 , \7541 , \7542 ,
         \7543 , \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 , \7552 ,
         \7553 , \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 , \7562 ,
         \7563 , \7564 , \7565 , \7566 , \7567 , \7568 , \7569 , \7570 , \7571 , \7572 ,
         \7573 , \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 , \7582 ,
         \7583 , \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 , \7592 ,
         \7593 , \7594 , \7595 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 , \7602 ,
         \7603 , \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 , \7612 ,
         \7613 , \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 , \7621 , \7622 ,
         \7623 , \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 , \7632 ,
         \7633 , \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 , \7642 ,
         \7643 , \7644 , \7645 , \7646 , \7647 , \7648 , \7649 , \7650 , \7651 , \7652 ,
         \7653 , \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 , \7662 ,
         \7663 , \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 , \7672 ,
         \7673 , \7674 , \7675 , \7676 , \7677 , \7678 , \7679 , \7680 , \7681 , \7682 ,
         \7683 , \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 , \7692 ,
         \7693 , \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 , \7702 ,
         \7703 , \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 , \7712 ,
         \7713 , \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 , \7722 ,
         \7723 , \7724 , \7725 , \7726 , \7727 , \7728 , \7729 , \7730 , \7731 , \7732 ,
         \7733 , \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 , \7742 ,
         \7743 , \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 , \7752 ,
         \7753 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 , \7762 ,
         \7763 , \7764 , \7765 , \7766 , \7767 , \7768 , \7769 , \7770 , \7771 , \7772 ,
         \7773 , \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 , \7782 ,
         \7783 , \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791 , \7792 ,
         \7793 , \7794 , \7795 , \7796 , \7797 , \7798 , \7799 , \7800 , \7801 , \7802 ,
         \7803 , \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 , \7811 , \7812 ,
         \7813 , \7814 , \7815 , \7816 , \7817 , \7818 , \7819 , \7820 , \7821 , \7822 ,
         \7823 , \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 , \7832 ,
         \7833 , \7834 , \7835 , \7836 , \7837 , \7838 , \7839 , \7840 , \7841 , \7842 ,
         \7843 , \7844 , \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 , \7852 ,
         \7853 , \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 , \7862 ,
         \7863 , \7864 , \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 , \7872 ,
         \7873 , \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 ,
         \7883 , \7884 , \7885 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891 , \7892 ,
         \7893 , \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 ,
         \7903 , \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 ,
         \7913 , \7914 , \7915 , \7916 , \7917 , \7918 , \7919 , \7920 , \7921 , \7922 ,
         \7923 , \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 ,
         \7933 , \7934 , \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 , \7942 ,
         \7943 , \7944 , \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 , \7952 ,
         \7953 , \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 ,
         \7963 , \7964 , \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 , \7972 ,
         \7973 , \7974 , \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 ,
         \7983 , \7984 , \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 , \7992 ,
         \7993 , \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 , \8002 ,
         \8003 , \8004 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 ,
         \8013 , \8014 , \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 , \8022 ,
         \8023 , \8024 , \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 , \8032 ,
         \8033 , \8034 , \8035 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 , \8042 ,
         \8043 , \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 ,
         \8053 , \8054 , \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 , \8062 ,
         \8063 , \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 , \8072 ,
         \8073 , \8074 , \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 , \8082 ,
         \8083 , \8084 , \8085 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 , \8092 ,
         \8093 , \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 ,
         \8103 , \8104 , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 , \8112 ,
         \8113 , \8114 , \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 , \8122 ,
         \8123 , \8124 , \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 , \8132 ,
         \8133 , \8134 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 , \8142 ,
         \8143 , \8144 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 , \8152 ,
         \8153 , \8154 , \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 , \8162 ,
         \8163 , \8164 , \8165 , \8166 , \8167 , \8168 , \8169 , \8170 , \8171 , \8172 ,
         \8173 , \8174 , \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 , \8182 ,
         \8183 , \8184 , \8185 , \8186 , \8187 , \8188 , \8189 , \8190 , \8191 , \8192 ,
         \8193 , \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 , \8202 ,
         \8203 , \8204 , \8205 , \8206 , \8207 , \8208 , \8209 , \8210 , \8211 , \8212 ,
         \8213 , \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 , \8222 ,
         \8223 , \8224 , \8225 , \8226 , \8227 , \8228 , \8229 , \8230 , \8231 , \8232 ,
         \8233 , \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 , \8242 ,
         \8243 , \8244 , \8245 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 , \8252 ,
         \8253 , \8254 , \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 , \8262 ,
         \8263 , \8264 , \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271 , \8272 ,
         \8273 , \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 , \8282 ,
         \8283 , \8284 , \8285 , \8286 , \8287 , \8288 , \8289 , \8290 , \8291 , \8292 ,
         \8293 , \8294 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 , \8302 ,
         \8303 , \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 , \8312 ,
         \8313 , \8314 , \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 , \8322 ,
         \8323 , \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 , \8332 ,
         \8333 , \8334 , \8335 , \8336 , \8337 , \8338 , \8339 , \8340 , \8341 , \8342 ,
         \8343 , \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 , \8352 ,
         \8353 , \8354 , \8355 , \8356 , \8357 , \8358 , \8359 , \8360 , \8361 , \8362 ,
         \8363 , \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 , \8372 ,
         \8373 , \8374 , \8375 , \8376 , \8377 , \8378 , \8379 , \8380 , \8381 , \8382 ,
         \8383 , \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 , \8392 ,
         \8393 , \8394 , \8395 , \8396 , \8397 , \8398 , \8399 , \8400 , \8401 , \8402 ,
         \8403 , \8404 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 , \8412 ,
         \8413 , \8414 , \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 , \8422 ,
         \8423 , \8424 , \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 , \8432 ,
         \8433 , \8434 , \8435 , \8436 , \8437 , \8438 , \8439 , \8440 , \8441 , \8442 ,
         \8443 , \8444 , \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 , \8452 ,
         \8453 , \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 , \8462 ,
         \8463 , \8464 , \8465 , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 , \8472 ,
         \8473 , \8474 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 , \8482 ,
         \8483 , \8484 , \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 , \8492 ,
         \8493 , \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 , \8502 ,
         \8503 , \8504 , \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511 , \8512 ,
         \8513 , \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 , \8522 ,
         \8523 , \8524 , \8525 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 , \8532 ,
         \8533 , \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 , \8542 ,
         \8543 , \8544 , \8545 , \8546 , \8547 , \8548 , \8549 , \8550 , \8551 , \8552 ,
         \8553 , \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 , \8562 ,
         \8563 , \8564 , \8565 , \8566 , \8567 , \8568 , \8569 , \8570 , \8571 , \8572 ,
         \8573 , \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 , \8582 ,
         \8583 , \8584 , \8585 , \8586 , \8587 , \8588 , \8589 , \8590 , \8591 , \8592 ,
         \8593 , \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 ,
         \8603 , \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 , \8612 ,
         \8613 , \8614 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 , \8622 ,
         \8623 , \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 , \8632 ,
         \8633 , \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 ,
         \8643 , \8644 , \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 ,
         \8653 , \8654 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 ,
         \8663 , \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 , \8672 ,
         \8673 , \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 , \8682 ,
         \8683 , \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 ,
         \8693 , \8694 , \8695 , \8696 , \8697 , \8698 , \8699 , \8700 , \8701 , \8702 ,
         \8703 , \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 ,
         \8713 , \8714 , \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 , \8722 ,
         \8723 , \8724 , \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 , \8732 ,
         \8733 , \8734 , \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 , \8742 ,
         \8743 , \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 , \8752 ,
         \8753 , \8754 , \8755 , \8756 , \8757 , \8758 , \8759 , \8760 , \8761 , \8762 ,
         \8763 , \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 , \8772 ,
         \8773 , \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 , \8782 ,
         \8783 , \8784 , \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 , \8792 ,
         \8793 , \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 , \8802 ,
         \8803 , \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 , \8812 ,
         \8813 , \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 , \8822 ,
         \8823 , \8824 , \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 , \8832 ,
         \8833 , \8834 , \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 , \8842 ,
         \8843 , \8844 , \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 , \8852 ,
         \8853 , \8854 , \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 , \8862 ,
         \8863 , \8864 , \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 , \8872 ,
         \8873 , \8874 , \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 , \8882 ,
         \8883 , \8884 , \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 , \8892 ,
         \8893 , \8894 , \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 , \8902 ,
         \8903 , \8904 , \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 , \8912 ,
         \8913 , \8914 , \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 , \8922 ,
         \8923 , \8924 , \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 , \8932 ,
         \8933 , \8934 , \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 , \8942 ,
         \8943 , \8944 , \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 , \8952 ,
         \8953 , \8954 , \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 , \8962 ,
         \8963 , \8964 , \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 , \8972 ,
         \8973 , \8974 , \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 , \8982 ,
         \8983 , \8984 , \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 , \8992 ,
         \8993 , \8994 , \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 , \9002 ,
         \9003 , \9004 , \9005 , \9006 , \9007 , \9008 , \9009 , \9010 , \9011 , \9012 ,
         \9013 , \9014 , \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 , \9022 ,
         \9023 , \9024 , \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 , \9032 ,
         \9033 , \9034 , \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 , \9042 ,
         \9043 , \9044 , \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 , \9052 ,
         \9053 , \9054 , \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 , \9062 ,
         \9063 , \9064 , \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 , \9072 ,
         \9073 , \9074 , \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 , \9082 ,
         \9083 , \9084 , \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 , \9092 ,
         \9093 , \9094 , \9095 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 , \9102 ,
         \9103 , \9104 , \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 , \9112 ,
         \9113 , \9114 , \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 , \9122 ,
         \9123 , \9124 , \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 , \9132 ,
         \9133 , \9134 , \9135 , \9136 , \9137 , \9138 , \9139 , \9140 , \9141 , \9142 ,
         \9143 , \9144 , \9145 , \9146 , \9147 , \9148 , \9149 , \9150 , \9151 , \9152 ,
         \9153 , \9154 , \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 , \9162 ,
         \9163 , \9164 , \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 , \9172 ,
         \9173 , \9174 , \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 , \9182 ,
         \9183 , \9184 , \9185 , \9186 , \9187 , \9188 , \9189 , \9190 , \9191 , \9192 ,
         \9193 , \9194 , \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 , \9202 ,
         \9203 , \9204 , \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 , \9212 ,
         \9213 , \9214 , \9215 , \9216 , \9217 , \9218 , \9219 , \9220 , \9221 , \9222 ,
         \9223 , \9224 , \9225 , \9226 , \9227 , \9228 , \9229 , \9230 , \9231 , \9232 ,
         \9233 , \9234 , \9235 , \9236 , \9237 , \9238 , \9239 , \9240 , \9241 , \9242 ,
         \9243 , \9244 , \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 , \9252 ,
         \9253 , \9254 , \9255 , \9256 , \9257 , \9258 , \9259 , \9260 , \9261 , \9262 ,
         \9263 , \9264 , \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 , \9272 ,
         \9273 , \9274 , \9275 , \9276 , \9277 , \9278 , \9279 , \9280 , \9281 , \9282 ,
         \9283 , \9284 , \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 , \9292 ,
         \9293 , \9294 , \9295 , \9296 , \9297 , \9298 , \9299 , \9300 , \9301 , \9302 ,
         \9303 , \9304 , \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 , \9312 ,
         \9313 , \9314 , \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 , \9322 ,
         \9323 , \9324 , \9325 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 , \9332 ,
         \9333 , \9334 , \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 , \9342 ,
         \9343 , \9344 , \9345 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 , \9352 ,
         \9353 , \9354 , \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 , \9362 ,
         \9363 , \9364 , \9365 , \9366 , \9367 , \9368 , \9369 , \9370 , \9371 , \9372 ,
         \9373 , \9374 , \9375 , \9376 , \9377 , \9378 , \9379 , \9380 , \9381 , \9382 ,
         \9383 , \9384 , \9385 , \9386 , \9387 , \9388 , \9389 , \9390 , \9391 , \9392 ,
         \9393 , \9394 , \9395 , \9396 , \9397 , \9398 , \9399 , \9400 , \9401 , \9402 ,
         \9403 , \9404 , \9405 , \9406 , \9407 , \9408 , \9409 , \9410 , \9411 , \9412 ,
         \9413 , \9414 , \9415 , \9416 , \9417 , \9418 , \9419 , \9420 , \9421 , \9422 ,
         \9423 , \9424 , \9425 , \9426 , \9427 , \9428 , \9429 , \9430 , \9431 , \9432 ,
         \9433 , \9434 , \9435 , \9436 , \9437 , \9438 , \9439 , \9440 , \9441 , \9442 ,
         \9443 , \9444 , \9445 , \9446 , \9447 , \9448 , \9449 , \9450 , \9451 , \9452 ,
         \9453 , \9454 , \9455 , \9456 , \9457 , \9458 , \9459 , \9460 , \9461 , \9462 ,
         \9463 , \9464 , \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471 , \9472 ,
         \9473 , \9474 , \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 , \9482 ,
         \9483 , \9484 , \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491 , \9492 ,
         \9493 , \9494 , \9495 , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 , \9502 ,
         \9503 , \9504 , \9505 , \9506 , \9507 , \9508 , \9509 , \9510 , \9511 , \9512 ,
         \9513 , \9514 , \9515 , \9516 , \9517 , \9518 , \9519 , \9520 , \9521 , \9522 ,
         \9523 , \9524 , \9525 , \9526 , \9527 , \9528 , \9529 , \9530 , \9531 , \9532 ,
         \9533 , \9534 , \9535 , \9536 , \9537 , \9538 , \9539 , \9540 , \9541 , \9542 ,
         \9543 , \9544 , \9545 , \9546 , \9547 , \9548 , \9549 , \9550 , \9551 , \9552 ,
         \9553 , \9554 , \9555 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 , \9562 ,
         \9563 , \9564 , \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 , \9572 ,
         \9573 , \9574 , \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 , \9582 ,
         \9583 , \9584 , \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 , \9592 ,
         \9593 , \9594 , \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 , \9602 ,
         \9603 , \9604 , \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 , \9612 ,
         \9613 , \9614 , \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 , \9622 ,
         \9623 , \9624 , \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 ,
         \9633 , \9634 , \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 ,
         \9643 , \9644 , \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 ,
         \9653 , \9654 , \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 ,
         \9663 , \9664 , \9665 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 , \9672 ,
         \9673 , \9674 , \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 ,
         \9683 , \9684 , \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 ,
         \9693 , \9694 , \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 , \9702 ,
         \9703 , \9704 , \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 ,
         \9713 , \9714 , \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 ,
         \9723 , \9724 , \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 ,
         \9733 , \9734 , \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 ,
         \9743 , \9744 , \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 ,
         \9753 , \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 ,
         \9763 , \9764 , \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 ,
         \9773 , \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 ,
         \9783 , \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 ,
         \9793 , \9794 , \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 ,
         \9803 , \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 ,
         \9813 , \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 ,
         \9823 , \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 ,
         \9833 , \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 ,
         \9843 , \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 ,
         \9853 , \9854 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 ,
         \9863 , \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 ,
         \9873 , \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 ,
         \9883 , \9884 , \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 ,
         \9893 , \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 ,
         \9903 , \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 ,
         \9913 , \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 ,
         \9923 , \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 ,
         \9933 , \9934 , \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 ,
         \9943 , \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 ,
         \9953 , \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 ,
         \9963 , \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 ,
         \9973 , \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 ,
         \9983 , \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 ,
         \9993 , \9994 , \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 ,
         \10003 , \10004 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 ,
         \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 ,
         \10023 , \10024 , \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 ,
         \10033 , \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 ,
         \10043 , \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 ,
         \10053 , \10054 , \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 , \10062 ,
         \10063 , \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 ,
         \10073 , \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 ,
         \10083 , \10084 , \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 ,
         \10093 , \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 ,
         \10103 , \10104 , \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 ,
         \10113 , \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 ,
         \10123 , \10124 , \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 , \10132 ,
         \10133 , \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 ,
         \10143 , \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 ,
         \10153 , \10154 , \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 ,
         \10163 , \10164 , \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 ,
         \10173 , \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 ,
         \10183 , \10184 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 ,
         \10193 , \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 ,
         \10203 , \10204 , \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 , \10212 ,
         \10213 , \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 ,
         \10223 , \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 ,
         \10233 , \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 ,
         \10243 , \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 ,
         \10253 , \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 , \10262 ,
         \10263 , \10264 , \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 ,
         \10273 , \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 ,
         \10283 , \10284 , \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 , \10292 ,
         \10293 , \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 ,
         \10303 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 ,
         \10313 , \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 ,
         \10323 , \10324 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 ,
         \10333 , \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 ,
         \10343 , \10344 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 ,
         \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 ,
         \10363 , \10364 , \10365 , \10366 , \10367 , \10368 , \10369 , \10370 , \10371 , \10372 ,
         \10373 , \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 ,
         \10383 , \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 ,
         \10393 , \10394 , \10395 , \10396 , \10397 , \10398 , \10399 , \10400 , \10401 , \10402 ,
         \10403 , \10404 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 ,
         \10413 , \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 , \10422 ,
         \10423 , \10424 , \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 ,
         \10433 , \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 ,
         \10443 , \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 ,
         \10453 , \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 ,
         \10463 , \10464 , \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 ,
         \10473 , \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 ,
         \10483 , \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 ,
         \10493 , \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 ,
         \10503 , \10504 , \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 ,
         \10513 , \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 ,
         \10523 , \10524 , \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 , \10532 ,
         \10533 , \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 ,
         \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 ,
         \10553 , \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 ,
         \10563 , \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 ,
         \10573 , \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 ,
         \10583 , \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 ,
         \10593 , \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 ,
         \10603 , \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 , \10612 ,
         \10613 , \10614 , \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 , \10622 ,
         \10623 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 ,
         \10633 , \10634 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 ,
         \10643 , \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 ,
         \10653 , \10654 , \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 ,
         \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 ,
         \10673 , \10674 , \10675 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 , \10682 ,
         \10683 , \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 ,
         \10693 , \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 , \10702 ,
         \10703 , \10704 , \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 , \10712 ,
         \10713 , \10714 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 ,
         \10723 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 ,
         \10733 , \10734 , \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 , \10742 ,
         \10743 , \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 ,
         \10753 , \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 ,
         \10763 , \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 ,
         \10773 , \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 ,
         \10783 , \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 ,
         \10793 , \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 , \10802 ,
         \10803 , \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 ,
         \10813 , \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 ,
         \10823 , \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 ,
         \10833 , \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 ,
         \10843 , \10844 , \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 ,
         \10853 , \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 ,
         \10863 , \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 ,
         \10873 , \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 ,
         \10883 , \10884 , \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 ,
         \10893 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 ,
         \10903 , \10904 , \10905 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 , \10912 ,
         \10913 , \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 ,
         \10923 , \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 , \10932 ,
         \10933 , \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 , \10942 ,
         \10943 , \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 ,
         \10953 , \10954 , \10955 , \10956 , \10957 , \10958 , \10959 , \10960 , \10961 , \10962 ,
         \10963 , \10964 , \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 , \10972 ,
         \10973 , \10974 , \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 , \10982 ,
         \10983 , \10984 , \10985 , \10986 , \10987 , \10988 , \10989 , \10990 , \10991 , \10992 ,
         \10993 , \10994 , \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 , \11002 ,
         \11003 , \11004 , \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 , \11012 ,
         \11013 , \11014 , \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 , \11022 ,
         \11023 , \11024 , \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 , \11032 ,
         \11033 , \11034 , \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 , \11042 ,
         \11043 , \11044 , \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 , \11052 ,
         \11053 , \11054 , \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 , \11062 ,
         \11063 , \11064 , \11065 , \11066 , \11067 , \11068 , \11069 , \11070 , \11071 , \11072 ,
         \11073 , \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 ,
         \11083 , \11084 , \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 , \11092 ,
         \11093 , \11094 , \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 , \11102 ,
         \11103 , \11104 , \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 , \11112 ,
         \11113 , \11114 , \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 , \11122 ,
         \11123 , \11124 , \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 , \11132 ,
         \11133 , \11134 , \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 , \11142 ,
         \11143 , \11144 , \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 , \11152 ,
         \11153 , \11154 , \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 , \11162 ,
         \11163 , \11164 , \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 , \11172 ,
         \11173 , \11174 , \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 , \11182 ,
         \11183 , \11184 , \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 , \11192 ,
         \11193 , \11194 , \11195 , \11196 , \11197 , \11198 , \11199 , \11200 , \11201 , \11202 ,
         \11203 , \11204 , \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 , \11212 ,
         \11213 , \11214 , \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 , \11222 ,
         \11223 , \11224 , \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 , \11232 ,
         \11233 , \11234 , \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 , \11242 ,
         \11243 , \11244 , \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 , \11252 ,
         \11253 , \11254 , \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 , \11262 ,
         \11263 , \11264 , \11265 , \11266 , \11267 , \11268 , \11269 , \11270 , \11271 , \11272 ,
         \11273 , \11274 , \11275 , \11276 , \11277 , \11278 , \11279 , \11280 , \11281 , \11282 ,
         \11283 , \11284 , \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 , \11292 ,
         \11293 , \11294 , \11295 , \11296 , \11297 , \11298 , \11299 , \11300 , \11301 , \11302 ,
         \11303 , \11304 , \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 , \11312 ,
         \11313 , \11314 , \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 , \11322 ,
         \11323 , \11324 , \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 , \11332 ,
         \11333 , \11334 , \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 , \11342 ,
         \11343 , \11344 , \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 , \11352 ,
         \11353 , \11354 , \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 , \11362 ,
         \11363 , \11364 , \11365 , \11366 , \11367 , \11368 , \11369 , \11370 , \11371 , \11372 ,
         \11373 , \11374 , \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 , \11382 ,
         \11383 , \11384 , \11385 , \11386 , \11387 , \11388 , \11389 , \11390 , \11391 , \11392 ,
         \11393 , \11394 , \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 , \11402 ,
         \11403 , \11404 , \11405 , \11406 , \11407 , \11408 , \11409 , \11410 , \11411 , \11412 ,
         \11413 , \11414 , \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 , \11422 ,
         \11423 , \11424 , \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 , \11432 ,
         \11433 , \11434 , \11435 , \11436 , \11437 , \11438 , \11439 , \11440 , \11441 , \11442 ,
         \11443 , \11444 , \11445 , \11446 , \11447 , \11448 , \11449 , \11450 , \11451 , \11452 ,
         \11453 , \11454 , \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 , \11462 ,
         \11463 , \11464 , \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 , \11472 ,
         \11473 , \11474 , \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 , \11482 ,
         \11483 , \11484 , \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 , \11492 ,
         \11493 , \11494 , \11495 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 , \11502 ,
         \11503 , \11504 , \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 , \11512 ,
         \11513 , \11514 , \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 , \11522 ,
         \11523 , \11524 , \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 , \11532 ,
         \11533 , \11534 , \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 , \11542 ,
         \11543 , \11544 , \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 , \11552 ,
         \11553 , \11554 , \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 , \11562 ,
         \11563 , \11564 , \11565 , \11566 , \11567 , \11568 , \11569 , \11570 , \11571 , \11572 ,
         \11573 , \11574 , \11575 , \11576 , \11577 , \11578 , \11579 , \11580 , \11581 , \11582 ,
         \11583 , \11584 , \11585 , \11586 , \11587 , \11588 , \11589 , \11590 , \11591 , \11592 ,
         \11593 , \11594 , \11595 , \11596 , \11597 , \11598 , \11599 , \11600 , \11601 , \11602 ,
         \11603 , \11604 , \11605 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 , \11612 ,
         \11613 , \11614 , \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 , \11622 ,
         \11623 , \11624 , \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 , \11632 ,
         \11633 , \11634 , \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 , \11642 ,
         \11643 , \11644 , \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 , \11652 ,
         \11653 , \11654 , \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661 , \11662 ,
         \11663 , \11664 , \11665 , \11666 , \11667 , \11668 , \11669 , \11670 , \11671 , \11672 ,
         \11673 , \11674 , \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 , \11682 ,
         \11683 , \11684 , \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 , \11692 ,
         \11693 , \11694 , \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 , \11702 ,
         \11703 , \11704 , \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 , \11712 ,
         \11713 , \11714 , \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 , \11722 ,
         \11723 , \11724 , \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 , \11732 ,
         \11733 , \11734 , \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 , \11742 ,
         \11743 , \11744 , \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 , \11752 ,
         \11753 , \11754 , \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 , \11762 ,
         \11763 , \11764 , \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 , \11772 ,
         \11773 , \11774 , \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 , \11782 ,
         \11783 , \11784 , \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 , \11792 ,
         \11793 , \11794 , \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 , \11802 ,
         \11803 , \11804 , \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 , \11812 ,
         \11813 , \11814 , \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 , \11822 ,
         \11823 , \11824 , \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 , \11832 ,
         \11833 , \11834 , \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 , \11842 ,
         \11843 , \11844 , \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 , \11852 ,
         \11853 , \11854 , \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 , \11862 ,
         \11863 , \11864 , \11865 , \11866 , \11867 , \11868 , \11869 , \11870 , \11871 , \11872 ,
         \11873 , \11874 , \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 , \11882 ,
         \11883 , \11884 , \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 , \11892 ,
         \11893 , \11894 , \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 , \11902 ,
         \11903 , \11904 , \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 , \11912 ,
         \11913 , \11914 , \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 , \11922 ,
         \11923 , \11924 , \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 , \11932 ,
         \11933 , \11934 , \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 , \11942 ,
         \11943 , \11944 , \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 , \11952 ,
         \11953 , \11954 , \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 , \11962 ,
         \11963 , \11964 , \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 , \11972 ,
         \11973 , \11974 , \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 , \11982 ,
         \11983 , \11984 , \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 , \11992 ,
         \11993 , \11994 , \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 , \12002 ,
         \12003 , \12004 , \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 , \12012 ,
         \12013 , \12014 , \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 , \12022 ,
         \12023 , \12024 , \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 , \12032 ,
         \12033 , \12034 , \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 , \12042 ,
         \12043 , \12044 , \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 , \12052 ,
         \12053 , \12054 , \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 , \12062 ,
         \12063 , \12064 , \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 , \12072 ,
         \12073 , \12074 , \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 , \12082 ,
         \12083 , \12084 , \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 , \12092 ,
         \12093 , \12094 , \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 , \12102 ,
         \12103 , \12104 , \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 , \12112 ,
         \12113 , \12114 , \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 , \12122 ,
         \12123 , \12124 , \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 , \12132 ,
         \12133 , \12134 , \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 , \12142 ,
         \12143 , \12144 , \12145 , \12146 , \12147 , \12148 , \12149 , \12150 , \12151 , \12152 ,
         \12153 , \12154 , \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 , \12162 ,
         \12163 , \12164 , \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 , \12172 ,
         \12173 , \12174 , \12175 , \12176 , \12177 , \12178 , \12179 , \12180 , \12181 , \12182 ,
         \12183 , \12184 , \12185 , \12186 , \12187 , \12188 , \12189 , \12190 , \12191 , \12192 ,
         \12193 , \12194 , \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 , \12202 ,
         \12203 , \12204 , \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 , \12212 ,
         \12213 , \12214 , \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 , \12222 ,
         \12223 , \12224 , \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 , \12232 ,
         \12233 , \12234 , \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 , \12242 ,
         \12243 , \12244 , \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 , \12252 ,
         \12253 , \12254 , \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 , \12262 ,
         \12263 , \12264 , \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 , \12272 ,
         \12273 , \12274 , \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 , \12282 ,
         \12283 , \12284 , \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 , \12292 ,
         \12293 , \12294 , \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 , \12302 ,
         \12303 , \12304 , \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 , \12312 ,
         \12313 , \12314 , \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 , \12322 ,
         \12323 , \12324 , \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 , \12332 ,
         \12333 , \12334 , \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 , \12342 ,
         \12343 , \12344 , \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 , \12352 ,
         \12353 , \12354 , \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 , \12362 ,
         \12363 , \12364 , \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 , \12372 ,
         \12373 , \12374 , \12375 , \12376 , \12377 , \12378 , \12379 , \12380 , \12381 , \12382 ,
         \12383 , \12384 , \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 , \12392 ,
         \12393 , \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 ,
         \12403 , \12404 , \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 , \12412 ,
         \12413 , \12414 , \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 , \12422 ,
         \12423 , \12424 , \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 , \12432 ,
         \12433 , \12434 , \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 , \12442 ,
         \12443 , \12444 , \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 , \12452 ,
         \12453 , \12454 , \12455 , \12456 , \12457 , \12458 , \12459 , \12460 , \12461 , \12462 ,
         \12463 , \12464 , \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 , \12472 ,
         \12473 , \12474 , \12475 , \12476 , \12477 , \12478 , \12479 , \12480 , \12481 , \12482 ,
         \12483 , \12484 , \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 , \12492 ,
         \12493 , \12494 , \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 , \12502 ,
         \12503 , \12504 , \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 , \12512 ,
         \12513 , \12514 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 ,
         \12523 , \12524 , \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 , \12532 ,
         \12533 , \12534 , \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 , \12542 ,
         \12543 , \12544 , \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 , \12552 ,
         \12553 , \12554 , \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 , \12562 ,
         \12563 , \12564 , \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 , \12572 ,
         \12573 , \12574 , \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 ,
         \12583 , \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 ,
         \12593 , \12594 , \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 , \12602 ,
         \12603 , \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 , \12612 ,
         \12613 , \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 , \12622 ,
         \12623 , \12624 , \12625 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 ,
         \12633 , \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 ,
         \12643 , \12644 , \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 , \12652 ,
         \12653 , \12654 , \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 , \12662 ,
         \12663 , \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 ,
         \12673 , \12674 , \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 ,
         \12683 , \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 ,
         \12693 , \12694 , \12695 , \12696 , \12697 , \12698 , \12699 , \12700 , \12701 , \12702 ,
         \12703 , \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 ,
         \12713 , \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 , \12722 ,
         \12723 , \12724 , \12725 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 ,
         \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 ,
         \12743 , \12744 , \12745 , \12746 , \12747 , \12748 , \12749 , \12750 , \12751 , \12752 ,
         \12753 , \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 ,
         \12763 , \12764 , \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 , \12772 ,
         \12773 , \12774 , \12775 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 , \12782 ,
         \12783 , \12784 , \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 , \12792 ,
         \12793 , \12794 , \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801 , \12802 ,
         \12803 , \12804 , \12805 , \12806 , \12807 , \12808 , \12809 , \12810 , \12811 , \12812 ,
         \12813 , \12814 , \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 , \12822 ,
         \12823 , \12824 , \12825 , \12826 , \12827 , \12828 , \12829 , \12830 , \12831 , \12832 ,
         \12833 , \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 ,
         \12843 , \12844 , \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851 , \12852 ,
         \12853 , \12854 , \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 , \12862 ,
         \12863 , \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 ,
         \12873 , \12874 , \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 ,
         \12883 , \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 ,
         \12893 , \12894 , \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 , \12902 ,
         \12903 , \12904 , \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 , \12912 ,
         \12913 , \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 ,
         \12923 , \12924 , \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 ,
         \12933 , \12934 , \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 , \12942 ,
         \12943 , \12944 , \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 , \12952 ,
         \12953 , \12954 , \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 ,
         \12963 , \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 ,
         \12973 , \12974 , \12975 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 , \12982 ,
         \12983 , \12984 , \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 ,
         \12993 , \12994 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 ,
         \13003 , \13004 , \13005 , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 , \13012 ,
         \13013 , \13014 , \13015 , \13016 , \13017 , \13018 , \13019 , \13020 , \13021 , \13022 ,
         \13023 , \13024 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 ,
         \13033 , \13034 , \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 , \13042 ,
         \13043 , \13044 , \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 , \13052 ,
         \13053 , \13054 , \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 , \13062 ,
         \13063 , \13064 , \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 , \13072 ,
         \13073 , \13074 , \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 , \13082 ,
         \13083 , \13084 , \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 , \13092 ,
         \13093 , \13094 , \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 , \13102 ,
         \13103 , \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 ,
         \13113 , \13114 , \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 ,
         \13123 , \13124 , \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 ,
         \13133 , \13134 , \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 , \13142 ,
         \13143 , \13144 , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 ,
         \13153 , \13154 , \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 ,
         \13163 , \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 , \13172 ,
         \13173 , \13174 , \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 , \13182 ,
         \13183 , \13184 , \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 , \13192 ,
         \13193 , \13194 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 ,
         \13203 , \13204 , \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 , \13212 ,
         \13213 , \13214 , \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 , \13222 ,
         \13223 , \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 ,
         \13233 , \13234 , \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 , \13242 ,
         \13243 , \13244 , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 , \13252 ,
         \13253 , \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 ,
         \13263 , \13264 , \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 , \13272 ,
         \13273 , \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 ,
         \13283 , \13284 , \13285 , \13286 , \13287 , \13288 , \13289 , \13290 , \13291 , \13292 ,
         \13293 , \13294 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 ,
         \13303 , \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 , \13312 ,
         \13313 , \13314 , \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 , \13322 ,
         \13323 , \13324 , \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 , \13332 ,
         \13333 , \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 ,
         \13343 , \13344 , \13345 , \13346 , \13347 , \13348 , \13349 , \13350 , \13351 , \13352 ,
         \13353 , \13354 , \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 , \13362 ,
         \13363 , \13364 , \13365 , \13366 , \13367 , \13368 , \13369 , \13370 , \13371 , \13372 ,
         \13373 , \13374 , \13375 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 , \13382 ,
         \13383 , \13384 , \13385 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 , \13392 ,
         \13393 , \13394 , \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 ,
         \13403 , \13404 , \13405 , \13406 , \13407 , \13408 , \13409 , \13410 , \13411 , \13412 ,
         \13413 , \13414 , \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 ,
         \13423 , \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 , \13432 ,
         \13433 , \13434 , \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 , \13442 ,
         \13443 , \13444 , \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 , \13452 ,
         \13453 , \13454 , \13455 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 ,
         \13463 , \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 ,
         \13473 , \13474 , \13475 , \13476 , \13477 , \13478 , \13479 , \13480 , \13481 , \13482 ,
         \13483 , \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 ,
         \13493 , \13494 , \13495 , \13496 , \13497 , \13498 , \13499 , \13500 , \13501 , \13502 ,
         \13503 , \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 ,
         \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 , \13522 ,
         \13523 , \13524 , \13525 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 , \13532 ,
         \13533 , \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 , \13542 ,
         \13543 , \13544 , \13545 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 , \13552 ,
         \13553 , \13554 , \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 , \13562 ,
         \13563 , \13564 , \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 ,
         \13573 , \13574 , \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 , \13582 ,
         \13583 , \13584 , \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 , \13592 ,
         \13593 , \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 , \13602 ,
         \13603 , \13604 , \13605 , \13606 , \13607 , \13608 , \13609 , \13610 , \13611 , \13612 ,
         \13613 , \13614 , \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 , \13622 ,
         \13623 , \13624 , \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 , \13632 ,
         \13633 , \13634 , \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 , \13642 ,
         \13643 , \13644 , \13645 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 , \13652 ,
         \13653 , \13654 , \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 , \13662 ,
         \13663 , \13664 , \13665 , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 , \13672 ,
         \13673 , \13674 , \13675 , \13676 , \13677 , \13678 , \13679 , \13680 , \13681 , \13682 ,
         \13683 , \13684 , \13685 , \13686 , \13687 , \13688 , \13689 , \13690 , \13691 , \13692 ,
         \13693 , \13694 , \13695 , \13696 , \13697 , \13698 , \13699 , \13700 , \13701 , \13702 ,
         \13703 , \13704 , \13705 , \13706 , \13707 , \13708 , \13709 , \13710 , \13711 , \13712 ,
         \13713 , \13714 , \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 , \13722 ,
         \13723 , \13724 , \13725 , \13726 , \13727 , \13728 , \13729 , \13730 , \13731 , \13732 ,
         \13733 , \13734 , \13735 , \13736 , \13737 , \13738 , \13739 , \13740 , \13741 , \13742 ,
         \13743 , \13744 , \13745 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 , \13752 ,
         \13753 , \13754 , \13755 , \13756 , \13757 , \13758 , \13759 , \13760 , \13761 , \13762 ,
         \13763 , \13764 , \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 , \13772 ,
         \13773 , \13774 , \13775 , \13776 , \13777 , \13778 , \13779 , \13780 , \13781 , \13782 ,
         \13783 , \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 ,
         \13793 , \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 , \13802 ,
         \13803 , \13804 , \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 , \13812 ,
         \13813 , \13814 , \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 , \13822 ,
         \13823 , \13824 , \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 , \13832 ,
         \13833 , \13834 , \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 ,
         \13843 , \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 , \13852 ,
         \13853 , \13854 , \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 , \13862 ,
         \13863 , \13864 , \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 , \13872 ,
         \13873 , \13874 , \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 , \13882 ,
         \13883 , \13884 , \13885 , \13886 , \13887 , \13888 , \13889 , \13890 , \13891 , \13892 ,
         \13893 , \13894 , \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 , \13902 ,
         \13903 , \13904 , \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 , \13912 ,
         \13913 , \13914 , \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 , \13922 ,
         \13923 , \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 ,
         \13933 , \13934 , \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 , \13942 ,
         \13943 , \13944 , \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 , \13952 ,
         \13953 , \13954 , \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 , \13962 ,
         \13963 , \13964 , \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 , \13972 ,
         \13973 , \13974 , \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 , \13982 ,
         \13983 , \13984 , \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 , \13992 ,
         \13993 , \13994 , \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 , \14002 ,
         \14003 , \14004 , \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 , \14012 ,
         \14013 , \14014 , \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 , \14022 ,
         \14023 , \14024 , \14025 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 , \14032 ,
         \14033 , \14034 , \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 , \14042 ,
         \14043 , \14044 , \14045 , \14046 , \14047 , \14048 , \14049 , \14050 , \14051 , \14052 ,
         \14053 , \14054 , \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 , \14062 ,
         \14063 , \14064 , \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 , \14072 ,
         \14073 , \14074 , \14075 , \14076 , \14077 , \14078 , \14079 , \14080 , \14081 , \14082 ,
         \14083 , \14084 , \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 , \14092 ,
         \14093 , \14094 , \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 , \14102 ,
         \14103 , \14104 , \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 , \14112 ,
         \14113 , \14114 , \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 , \14122 ,
         \14123 , \14124 , \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 , \14132 ,
         \14133 , \14134 , \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 , \14142 ,
         \14143 , \14144 , \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 , \14152 ,
         \14153 , \14154 , \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 , \14162 ,
         \14163 , \14164 , \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 , \14172 ,
         \14173 , \14174 , \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 , \14182 ,
         \14183 , \14184 , \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 , \14192 ,
         \14193 , \14194 , \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 , \14202 ,
         \14203 , \14204 , \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 , \14212 ,
         \14213 , \14214 , \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 , \14222 ,
         \14223 , \14224 , \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 , \14232 ,
         \14233 , \14234 , \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 , \14242 ,
         \14243 , \14244 , \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 , \14252 ,
         \14253 , \14254 , \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 , \14262 ,
         \14263 , \14264 , \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 , \14272 ,
         \14273 , \14274 , \14275 , \14276 , \14277 , \14278 , \14279 , \14280 , \14281 , \14282 ,
         \14283 , \14284 , \14285 , \14286 , \14287 , \14288 , \14289 , \14290 , \14291 , \14292 ,
         \14293 , \14294 , \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 , \14302 ,
         \14303 , \14304 , \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 , \14312 ,
         \14313 , \14314 , \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 , \14322 ,
         \14323 , \14324 , \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 , \14332 ,
         \14333 , \14334 , \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 , \14342 ,
         \14343 , \14344 , \14345 , \14346 , \14347 , \14348 , \14349 , \14350 , \14351 , \14352 ,
         \14353 , \14354 , \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 , \14362 ,
         \14363 , \14364 , \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 , \14372 ,
         \14373 , \14374 , \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 , \14382 ,
         \14383 , \14384 , \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 , \14392 ,
         \14393 , \14394 , \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 , \14402 ,
         \14403 , \14404 , \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 , \14412 ,
         \14413 , \14414 , \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 , \14422 ,
         \14423 , \14424 , \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 , \14432 ,
         \14433 , \14434 , \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 , \14442 ,
         \14443 , \14444 , \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 , \14452 ,
         \14453 , \14454 , \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 , \14462 ,
         \14463 , \14464 , \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 , \14472 ,
         \14473 , \14474 , \14475 , \14476 , \14477 , \14478 , \14479 , \14480 , \14481 , \14482 ,
         \14483 , \14484 , \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 , \14492 ,
         \14493 , \14494 , \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 , \14502 ,
         \14503 , \14504 , \14505 , \14506 , \14507 , \14508 , \14509 , \14510 , \14511 , \14512 ,
         \14513 , \14514 , \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 , \14522 ,
         \14523 , \14524 , \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 , \14532 ,
         \14533 , \14534 , \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 , \14542 ,
         \14543 , \14544 , \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 , \14552 ,
         \14553 , \14554 , \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 , \14562 ,
         \14563 , \14564 , \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 , \14572 ,
         \14573 , \14574 , \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 , \14582 ,
         \14583 , \14584 , \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 , \14592 ,
         \14593 , \14594 , \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 , \14602 ,
         \14603 , \14604 , \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 , \14612 ,
         \14613 , \14614 , \14615 , \14616 , \14617 , \14618 , \14619 , \14620 , \14621 , \14622 ,
         \14623 , \14624 , \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 , \14632 ,
         \14633 , \14634 , \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 , \14642 ,
         \14643 , \14644 , \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 , \14652 ,
         \14653 , \14654 , \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 , \14662 ,
         \14663 , \14664 , \14665 , \14666 , \14667 , \14668 , \14669 , \14670 , \14671 , \14672 ,
         \14673 , \14674 , \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 , \14682 ,
         \14683 , \14684 , \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 , \14692 ,
         \14693 , \14694 , \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 , \14702 ,
         \14703 , \14704 , \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 , \14712 ,
         \14713 , \14714 , \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 , \14722 ,
         \14723 , \14724 , \14725 , \14726 , \14727 , \14728 , \14729 , \14730 , \14731 , \14732 ,
         \14733 , \14734 , \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 , \14742 ,
         \14743 , \14744 , \14745 , \14746 , \14747 , \14748 , \14749 , \14750 , \14751 , \14752 ,
         \14753 , \14754 , \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 , \14762 ,
         \14763 , \14764 , \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 , \14772 ,
         \14773 , \14774 , \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 , \14782 ,
         \14783 , \14784 , \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14791 , \14792 ,
         \14793 , \14794 , \14795 , \14796 , \14797 , \14798 , \14799 , \14800 , \14801 , \14802 ,
         \14803 , \14804 , \14805 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 , \14812 ,
         \14813 , \14814 , \14815 , \14816 , \14817 , \14818 , \14819 , \14820 , \14821 , \14822 ,
         \14823 , \14824 , \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831 , \14832 ,
         \14833 , \14834 , \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 , \14842 ,
         \14843 , \14844 , \14845 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 , \14852 ,
         \14853 , \14854 , \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 , \14862 ,
         \14863 , \14864 , \14865 , \14866 , \14867 , \14868 , \14869 , \14870 , \14871 , \14872 ,
         \14873 , \14874 , \14875 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 , \14882 ,
         \14883 , \14884 , \14885 , \14886 , \14887 , \14888 , \14889 , \14890 , \14891 , \14892 ,
         \14893 , \14894 , \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 , \14902 ,
         \14903 , \14904 , \14905 , \14906 , \14907 , \14908 , \14909 , \14910 , \14911 , \14912 ,
         \14913 , \14914 , \14915 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 , \14922 ,
         \14923 , \14924 , \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 , \14932 ,
         \14933 , \14934 , \14935 , \14936 , \14937 , \14938 , \14939 , \14940 , \14941 , \14942 ,
         \14943 , \14944 , \14945 , \14946 , \14947 , \14948 , \14949 , \14950 , \14951 , \14952 ,
         \14953 , \14954 , \14955 , \14956 , \14957 , \14958 , \14959 , \14960 , \14961 , \14962 ,
         \14963 , \14964 , \14965 , \14966 , \14967 , \14968 , \14969 , \14970 , \14971 , \14972 ,
         \14973 , \14974 , \14975 , \14976 , \14977 , \14978 , \14979 , \14980 , \14981 , \14982 ,
         \14983 , \14984 , \14985 , \14986 , \14987 , \14988 , \14989 , \14990 , \14991 , \14992 ,
         \14993 , \14994 , \14995 , \14996 , \14997 , \14998 , \14999 , \15000 , \15001 , \15002 ,
         \15003 , \15004 , \15005 , \15006 , \15007 , \15008 , \15009 , \15010 , \15011 , \15012 ,
         \15013 , \15014 , \15015 , \15016 , \15017 , \15018 , \15019 , \15020 , \15021 , \15022 ,
         \15023 , \15024 , \15025 , \15026 , \15027 , \15028 , \15029 , \15030 , \15031 , \15032 ,
         \15033 , \15034 , \15035 , \15036 , \15037 , \15038 , \15039 , \15040 , \15041 , \15042 ,
         \15043 , \15044 , \15045 , \15046 , \15047 , \15048 , \15049 , \15050 , \15051 , \15052 ,
         \15053 , \15054 , \15055 , \15056 , \15057 , \15058 , \15059 , \15060 , \15061 , \15062 ,
         \15063 , \15064 , \15065 , \15066 , \15067 , \15068 , \15069 , \15070 , \15071 , \15072 ,
         \15073 , \15074 , \15075 , \15076 , \15077 , \15078 , \15079 , \15080 , \15081 , \15082 ,
         \15083 , \15084 , \15085 , \15086 , \15087 , \15088 , \15089 , \15090 , \15091 , \15092 ,
         \15093 , \15094 , \15095 , \15096 , \15097 , \15098 , \15099 , \15100 , \15101 , \15102 ,
         \15103 , \15104 , \15105 , \15106 , \15107 , \15108 , \15109 , \15110 , \15111 , \15112 ,
         \15113 , \15114 , \15115 , \15116 , \15117 , \15118 , \15119 , \15120 , \15121 , \15122 ,
         \15123 , \15124 , \15125 , \15126 , \15127 , \15128 , \15129 , \15130 , \15131 , \15132 ,
         \15133 , \15134 , \15135 , \15136 , \15137 , \15138 , \15139 , \15140 , \15141 , \15142 ,
         \15143 , \15144 , \15145 , \15146 , \15147 , \15148 , \15149 , \15150 , \15151 , \15152 ,
         \15153 , \15154 , \15155 , \15156 , \15157 , \15158 , \15159 , \15160 , \15161 , \15162 ,
         \15163 , \15164 , \15165 , \15166 , \15167 , \15168 , \15169 , \15170 , \15171 , \15172 ,
         \15173 , \15174 , \15175 , \15176 , \15177 , \15178 , \15179 , \15180 , \15181 , \15182 ,
         \15183 , \15184 , \15185 , \15186 , \15187 , \15188 , \15189 , \15190 , \15191 , \15192 ,
         \15193 , \15194 , \15195 , \15196 , \15197 , \15198 , \15199 , \15200 , \15201 , \15202 ,
         \15203 , \15204 , \15205 , \15206 , \15207 , \15208 , \15209 , \15210 , \15211 , \15212 ,
         \15213 , \15214 , \15215 , \15216 , \15217 , \15218 , \15219 , \15220 , \15221 , \15222 ,
         \15223 , \15224 , \15225 , \15226 , \15227 , \15228 , \15229 , \15230 , \15231 , \15232 ,
         \15233 , \15234 , \15235 , \15236 , \15237 , \15238 , \15239 , \15240 , \15241 , \15242 ,
         \15243 , \15244 , \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 , \15252 ,
         \15253 , \15254 , \15255 , \15256 , \15257 , \15258 , \15259 , \15260 , \15261 , \15262 ,
         \15263 , \15264 , \15265 , \15266 , \15267 , \15268 , \15269 , \15270 , \15271 , \15272 ,
         \15273 , \15274 , \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 , \15282 ,
         \15283 , \15284 , \15285 , \15286 , \15287 , \15288 , \15289 , \15290 , \15291 , \15292 ,
         \15293 , \15294 , \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 , \15302 ,
         \15303 , \15304 , \15305 , \15306 , \15307 , \15308 , \15309 , \15310 , \15311 , \15312 ,
         \15313 , \15314 , \15315 , \15316 , \15317 , \15318 , \15319 , \15320 , \15321 , \15322 ,
         \15323 , \15324 , \15325 , \15326 , \15327 , \15328 , \15329 , \15330 , \15331 , \15332 ,
         \15333 , \15334 , \15335 , \15336 , \15337 , \15338 , \15339 , \15340 , \15341 , \15342 ,
         \15343 , \15344 , \15345 , \15346 , \15347 , \15348 , \15349 , \15350 , \15351 , \15352 ,
         \15353 , \15354 , \15355 , \15356 , \15357 , \15358 , \15359 , \15360 , \15361 , \15362 ,
         \15363 , \15364 , \15365 , \15366 , \15367 , \15368 , \15369 , \15370 , \15371 , \15372 ,
         \15373 , \15374 , \15375 , \15376 , \15377 , \15378 , \15379 , \15380 , \15381 , \15382 ,
         \15383 , \15384 , \15385 , \15386 , \15387 , \15388 , \15389 , \15390 , \15391 , \15392 ,
         \15393 , \15394 , \15395 , \15396 , \15397 , \15398 , \15399 , \15400 , \15401 , \15402 ,
         \15403 , \15404 , \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411 , \15412 ,
         \15413 , \15414 , \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 , \15422 ,
         \15423 , \15424 , \15425 , \15426 , \15427 , \15428 , \15429 , \15430 , \15431 , \15432 ,
         \15433 , \15434 , \15435 , \15436 , \15437 , \15438 , \15439 , \15440 , \15441 , \15442 ,
         \15443 , \15444 , \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 , \15452 ,
         \15453 , \15454 , \15455 , \15456 , \15457 , \15458 , \15459 , \15460 , \15461 , \15462 ,
         \15463 , \15464 , \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15471 , \15472 ,
         \15473 , \15474 , \15475 , \15476 , \15477 , \15478 , \15479 , \15480 , \15481 , \15482 ,
         \15483 , \15484 , \15485 , \15486 , \15487 , \15488 , \15489 , \15490 , \15491 , \15492 ,
         \15493 , \15494 , \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 , \15502 ,
         \15503 , \15504 , \15505 , \15506 , \15507 , \15508 , \15509 , \15510 , \15511 , \15512 ,
         \15513 , \15514 , \15515 , \15516 , \15517 , \15518 , \15519 , \15520 , \15521 , \15522 ,
         \15523 , \15524 , \15525 , \15526 , \15527 , \15528 , \15529 , \15530 , \15531 , \15532 ,
         \15533 , \15534 , \15535 , \15536 , \15537 , \15538 , \15539 , \15540 , \15541 , \15542 ,
         \15543 , \15544 , \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 , \15552 ,
         \15553 , \15554 , \15555 , \15556 , \15557 , \15558 , \15559 , \15560 , \15561 , \15562 ,
         \15563 , \15564 , \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 , \15572 ,
         \15573 , \15574 , \15575 , \15576 , \15577 , \15578 , \15579 , \15580 , \15581 , \15582 ,
         \15583 , \15584 , \15585 , \15586 , \15587 , \15588 , \15589 , \15590 , \15591 , \15592 ,
         \15593 , \15594 , \15595 , \15596 , \15597 , \15598 , \15599 , \15600 , \15601 , \15602 ,
         \15603 , \15604 , \15605 , \15606 , \15607 , \15608 , \15609 , \15610 , \15611 , \15612 ,
         \15613 , \15614 , \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 , \15622 ,
         \15623 , \15624 , \15625 , \15626 , \15627 , \15628 , \15629 , \15630 , \15631 , \15632 ,
         \15633 , \15634 , \15635 , \15636 , \15637 , \15638 , \15639 , \15640 , \15641 , \15642 ,
         \15643 , \15644 , \15645 , \15646 , \15647 , \15648 , \15649 , \15650 , \15651 , \15652 ,
         \15653 , \15654 , \15655 , \15656 , \15657 , \15658 , \15659 , \15660 , \15661 , \15662 ,
         \15663 , \15664 , \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 , \15672 ,
         \15673 , \15674 , \15675 , \15676 , \15677 , \15678 , \15679 , \15680 , \15681 , \15682 ,
         \15683 , \15684 , \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 , \15692 ,
         \15693 , \15694 , \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 , \15702 ,
         \15703 , \15704 , \15705 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 , \15712 ,
         \15713 , \15714 , \15715 , \15716 , \15717 , \15718 , \15719 , \15720 , \15721 , \15722 ,
         \15723 , \15724 , \15725 , \15726 , \15727 , \15728 , \15729 , \15730 , \15731 , \15732 ,
         \15733 , \15734 , \15735 , \15736 , \15737 , \15738 , \15739 , \15740 , \15741 , \15742 ,
         \15743 , \15744 , \15745 , \15746 , \15747 , \15748 , \15749 , \15750 , \15751 , \15752 ,
         \15753 , \15754 , \15755 , \15756 , \15757 , \15758 , \15759 , \15760 , \15761 , \15762 ,
         \15763 , \15764 , \15765 , \15766 , \15767 , \15768 , \15769 , \15770 , \15771 , \15772 ,
         \15773 , \15774 , \15775 , \15776 , \15777 , \15778 , \15779 , \15780 , \15781 , \15782 ,
         \15783 , \15784 , \15785 , \15786 , \15787 , \15788 , \15789 , \15790 , \15791 , \15792 ,
         \15793 , \15794 , \15795 , \15796 , \15797 , \15798 , \15799 , \15800 , \15801 , \15802 ,
         \15803 , \15804 , \15805 , \15806 , \15807 , \15808 , \15809 , \15810 , \15811 , \15812 ,
         \15813 , \15814 , \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , \15821 , \15822 ,
         \15823 , \15824 , \15825 , \15826 , \15827 , \15828 , \15829 , \15830 , \15831 , \15832 ,
         \15833 , \15834 , \15835 , \15836 , \15837 , \15838 , \15839 , \15840 , \15841 , \15842 ,
         \15843 , \15844 , \15845 , \15846 , \15847 , \15848 , \15849 , \15850 , \15851 , \15852 ,
         \15853 , \15854 , \15855 , \15856 , \15857 , \15858 , \15859 , \15860 , \15861 , \15862 ,
         \15863 , \15864 , \15865 , \15866 , \15867 , \15868 , \15869 , \15870 , \15871 , \15872 ,
         \15873 , \15874 , \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 , \15882 ,
         \15883 , \15884 , \15885 , \15886 , \15887 , \15888 , \15889 , \15890 , \15891 , \15892 ,
         \15893 , \15894 , \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 , \15902 ,
         \15903 , \15904 , \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 , \15912 ,
         \15913 , \15914 , \15915 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 , \15922 ,
         \15923 , \15924 , \15925 , \15926 , \15927 , \15928 , \15929 , \15930 , \15931 , \15932 ,
         \15933 , \15934 , \15935 , \15936 , \15937 , \15938 , \15939 , \15940 , \15941 , \15942 ,
         \15943 , \15944 , \15945 , \15946 , \15947 , \15948 , \15949 , \15950 , \15951 , \15952 ,
         \15953 , \15954 , \15955 , \15956 , \15957 , \15958 , \15959 , \15960 , \15961 , \15962 ,
         \15963 , \15964 , \15965 , \15966 , \15967 , \15968 , \15969 , \15970 , \15971 , \15972 ,
         \15973 , \15974 , \15975 , \15976 , \15977 , \15978 , \15979 , \15980 , \15981 , \15982 ,
         \15983 , \15984 , \15985 , \15986 , \15987 , \15988 , \15989 , \15990 , \15991 , \15992 ,
         \15993 , \15994 , \15995 , \15996 , \15997 , \15998 , \15999 , \16000 , \16001 , \16002 ,
         \16003 , \16004 , \16005 , \16006 , \16007 , \16008 , \16009 , \16010 , \16011 , \16012 ,
         \16013 , \16014 , \16015 , \16016 , \16017 , \16018 , \16019 , \16020 , \16021 , \16022 ,
         \16023 , \16024 , \16025 , \16026 , \16027 , \16028 , \16029 , \16030 , \16031 , \16032 ,
         \16033 , \16034 , \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 , \16042 ,
         \16043 , \16044 , \16045 , \16046 , \16047 , \16048 , \16049 , \16050 , \16051 , \16052 ,
         \16053 , \16054 , \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 , \16062 ,
         \16063 , \16064 , \16065 , \16066 , \16067 , \16068 , \16069 , \16070 , \16071 , \16072 ,
         \16073 , \16074 , \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 , \16082 ,
         \16083 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 , \16092 ,
         \16093 , \16094 , \16095 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 , \16102 ,
         \16103 , \16104 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 , \16112 ,
         \16113 , \16114 , \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 , \16122 ,
         \16123 , \16124 , \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 , \16132 ,
         \16133 , \16134 , \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 , \16142 ,
         \16143 , \16144 , \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 , \16152 ,
         \16153 , \16154 , \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 , \16162 ,
         \16163 , \16164 , \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 , \16172 ,
         \16173 , \16174 , \16175 , \16176 , \16177 , \16178 , \16179 , \16180 , \16181 , \16182 ,
         \16183 , \16184 , \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 , \16192 ,
         \16193 , \16194 , \16195 , \16196 , \16197 , \16198 , \16199 , \16200 , \16201 , \16202 ,
         \16203 , \16204 , \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 , \16212 ,
         \16213 , \16214 , \16215 , \16216 , \16217 , \16218 , \16219 , \16220 , \16221 , \16222 ,
         \16223 , \16224 , \16225 , \16226 , \16227 , \16228 , \16229 , \16230 , \16231 , \16232 ,
         \16233 , \16234 , \16235 , \16236 , \16237 , \16238 , \16239 , \16240 , \16241 , \16242 ,
         \16243 , \16244 , \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 , \16252 ,
         \16253 , \16254 , \16255 , \16256 , \16257 , \16258 , \16259 , \16260 , \16261 , \16262 ,
         \16263 , \16264 , \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 , \16272 ,
         \16273 , \16274 , \16275 , \16276 , \16277 , \16278 , \16279 , \16280 , \16281 , \16282 ,
         \16283 , \16284 , \16285 , \16286 , \16287 , \16288 , \16289 , \16290 , \16291 , \16292 ,
         \16293 , \16294 , \16295 , \16296 , \16297 , \16298 , \16299 , \16300 , \16301 , \16302 ,
         \16303 , \16304 , \16305 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 , \16312 ,
         \16313 , \16314 , \16315 , \16316 , \16317 , \16318 , \16319 , \16320 , \16321 , \16322 ,
         \16323 , \16324 , \16325 , \16326 , \16327 , \16328 , \16329 , \16330 , \16331 , \16332 ,
         \16333 , \16334 , \16335 , \16336 , \16337 , \16338 , \16339 , \16340 , \16341 , \16342 ,
         \16343 , \16344 , \16345 , \16346 , \16347 , \16348 , \16349 , \16350 , \16351 , \16352 ,
         \16353 , \16354 , \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 , \16362 ,
         \16363 , \16364 , \16365 , \16366 , \16367 , \16368 , \16369 , \16370 , \16371 , \16372 ,
         \16373 , \16374 , \16375 , \16376 , \16377 , \16378 , \16379 , \16380 , \16381 , \16382 ,
         \16383 , \16384 , \16385 , \16386 , \16387 , \16388 , \16389 , \16390 , \16391 , \16392 ,
         \16393 , \16394 , \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 , \16402 ,
         \16403 , \16404 , \16405 , \16406 , \16407 , \16408 , \16409 , \16410 , \16411 , \16412 ,
         \16413 , \16414 , \16415 , \16416 , \16417 , \16418 , \16419 , \16420 , \16421 , \16422 ,
         \16423 , \16424 , \16425 , \16426 , \16427 , \16428 , \16429 , \16430 , \16431 , \16432 ,
         \16433 , \16434 , \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 , \16442 ,
         \16443 , \16444 , \16445 , \16446 , \16447 , \16448 , \16449 , \16450 , \16451 , \16452 ,
         \16453 , \16454 , \16455 , \16456 , \16457 , \16458 , \16459 , \16460 , \16461 , \16462 ,
         \16463 , \16464 , \16465 , \16466 , \16467 , \16468 , \16469 , \16470 , \16471 , \16472 ,
         \16473 , \16474 , \16475 , \16476 , \16477 , \16478 , \16479 , \16480 , \16481 , \16482 ,
         \16483 , \16484 , \16485 , \16486 , \16487 , \16488 , \16489 , \16490 , \16491 , \16492 ,
         \16493 , \16494 , \16495 , \16496 , \16497 , \16498 , \16499 , \16500 , \16501 , \16502 ,
         \16503 , \16504 , \16505 , \16506 , \16507 , \16508 , \16509 , \16510 , \16511 , \16512 ,
         \16513 , \16514 , \16515 , \16516 , \16517 , \16518 , \16519 , \16520 , \16521 , \16522 ,
         \16523 , \16524 , \16525 , \16526 , \16527 , \16528 , \16529 , \16530 , \16531 , \16532 ,
         \16533 , \16534 , \16535 , \16536 , \16537 , \16538 , \16539 , \16540 , \16541 , \16542 ,
         \16543 , \16544 , \16545 , \16546 , \16547 , \16548 , \16549 , \16550 , \16551 , \16552 ,
         \16553 , \16554 , \16555 , \16556 , \16557 , \16558 , \16559 , \16560 , \16561 , \16562 ,
         \16563 , \16564 , \16565 , \16566 , \16567 , \16568 , \16569 , \16570 , \16571 , \16572 ,
         \16573 , \16574 , \16575 , \16576 , \16577 , \16578 , \16579 , \16580 , \16581 , \16582 ,
         \16583 , \16584 , \16585 , \16586 , \16587 , \16588 , \16589 , \16590 , \16591 , \16592 ,
         \16593 , \16594 , \16595 , \16596 , \16597 , \16598 , \16599 , \16600 , \16601 , \16602 ,
         \16603 , \16604 , \16605 , \16606 , \16607 , \16608 , \16609 , \16610 , \16611 , \16612 ,
         \16613 , \16614 , \16615 , \16616 , \16617 , \16618 , \16619 , \16620 , \16621 , \16622 ,
         \16623 , \16624 , \16625 , \16626 , \16627 , \16628 , \16629 , \16630 , \16631 , \16632 ,
         \16633 , \16634 , \16635 , \16636 , \16637 , \16638 , \16639 , \16640 , \16641 , \16642 ,
         \16643 , \16644 , \16645 , \16646 , \16647 , \16648 , \16649 , \16650 , \16651 , \16652 ,
         \16653 , \16654 , \16655 , \16656 , \16657 , \16658 , \16659 , \16660 , \16661 , \16662 ,
         \16663 , \16664 , \16665 , \16666 , \16667 , \16668 , \16669 , \16670 , \16671 , \16672 ,
         \16673 , \16674 , \16675 , \16676 , \16677 , \16678 , \16679 , \16680 , \16681 , \16682 ,
         \16683 , \16684 , \16685 , \16686 , \16687 , \16688 , \16689 , \16690 , \16691 , \16692 ,
         \16693 , \16694 , \16695 , \16696 , \16697 , \16698 , \16699 , \16700 , \16701 , \16702 ,
         \16703 , \16704 , \16705 , \16706 , \16707 , \16708 , \16709 , \16710 , \16711 , \16712 ,
         \16713 , \16714 , \16715 , \16716 , \16717 , \16718 , \16719 , \16720 , \16721 , \16722 ,
         \16723 , \16724 , \16725 , \16726 , \16727 , \16728 , \16729 , \16730 , \16731 , \16732 ,
         \16733 , \16734 , \16735 , \16736 , \16737 , \16738 , \16739 , \16740 , \16741 , \16742 ,
         \16743 , \16744 , \16745 , \16746 , \16747 , \16748 , \16749 , \16750 , \16751 , \16752 ,
         \16753 , \16754 , \16755 , \16756 , \16757 , \16758 , \16759 , \16760 , \16761 , \16762 ,
         \16763 , \16764 , \16765 , \16766 , \16767 , \16768 , \16769 , \16770 , \16771 , \16772 ,
         \16773 , \16774 , \16775 , \16776 , \16777 , \16778 , \16779 , \16780 , \16781 , \16782 ,
         \16783 , \16784 , \16785 , \16786 , \16787 , \16788 , \16789 , \16790 , \16791 , \16792 ,
         \16793 , \16794 , \16795 , \16796 , \16797 , \16798 , \16799 , \16800 , \16801 , \16802 ,
         \16803 , \16804 , \16805 , \16806 , \16807 , \16808 , \16809 , \16810 , \16811 , \16812 ,
         \16813 , \16814 , \16815 , \16816 , \16817 , \16818 , \16819 , \16820 , \16821 , \16822 ,
         \16823 , \16824 , \16825 , \16826 , \16827 , \16828 , \16829 , \16830 , \16831 , \16832 ,
         \16833 , \16834 , \16835 , \16836 , \16837 , \16838 , \16839 , \16840 , \16841 , \16842 ,
         \16843 , \16844 , \16845 , \16846 , \16847 , \16848 , \16849 , \16850 , \16851 , \16852 ,
         \16853 , \16854 , \16855 , \16856 , \16857 , \16858 , \16859 , \16860 , \16861 , \16862 ,
         \16863 , \16864 , \16865 , \16866 , \16867 , \16868 , \16869 , \16870 , \16871 , \16872 ,
         \16873 , \16874 , \16875 , \16876 , \16877 , \16878 , \16879 , \16880 , \16881 , \16882 ,
         \16883 , \16884 , \16885 , \16886 , \16887 , \16888 , \16889 , \16890 , \16891 , \16892 ,
         \16893 , \16894 , \16895 , \16896 , \16897 , \16898 , \16899 , \16900 , \16901 , \16902 ,
         \16903 , \16904 , \16905 , \16906 , \16907 , \16908 , \16909 , \16910 , \16911 , \16912 ,
         \16913 , \16914 , \16915 , \16916 , \16917 , \16918 , \16919 , \16920 , \16921 , \16922 ,
         \16923 , \16924 , \16925 , \16926 , \16927 , \16928 , \16929 , \16930 , \16931 , \16932 ,
         \16933 , \16934 , \16935 , \16936 , \16937 , \16938 , \16939 , \16940 , \16941 , \16942 ,
         \16943 , \16944 , \16945 , \16946 , \16947 , \16948 , \16949 , \16950 , \16951 , \16952 ,
         \16953 , \16954 , \16955 , \16956 , \16957 , \16958 , \16959 , \16960 , \16961 , \16962 ,
         \16963 , \16964 , \16965 , \16966 , \16967 , \16968 , \16969 , \16970 , \16971 , \16972 ,
         \16973 , \16974 , \16975 , \16976 , \16977 , \16978 , \16979 , \16980 , \16981 , \16982 ,
         \16983 , \16984 , \16985 , \16986 , \16987 , \16988 , \16989 , \16990 , \16991 , \16992 ,
         \16993 , \16994 , \16995 , \16996 , \16997 , \16998 , \16999 , \17000 , \17001 , \17002 ,
         \17003 , \17004 , \17005 , \17006 , \17007 , \17008 , \17009 , \17010 , \17011 , \17012 ,
         \17013 , \17014 , \17015 , \17016 , \17017 , \17018 , \17019 , \17020 , \17021 , \17022 ,
         \17023 , \17024 , \17025 , \17026 , \17027 , \17028 , \17029 , \17030 , \17031 , \17032 ,
         \17033 , \17034 , \17035 , \17036 , \17037 , \17038 , \17039 , \17040 , \17041 , \17042 ,
         \17043 , \17044 , \17045 , \17046 , \17047 , \17048 , \17049 , \17050 , \17051 , \17052 ,
         \17053 , \17054 , \17055 , \17056 , \17057 , \17058 , \17059 , \17060 , \17061 , \17062 ,
         \17063 , \17064 , \17065 , \17066 , \17067 , \17068 , \17069 , \17070 , \17071 , \17072 ,
         \17073 , \17074 , \17075 , \17076 , \17077 , \17078 , \17079 , \17080 , \17081 , \17082 ,
         \17083 , \17084 , \17085 , \17086 , \17087 , \17088 , \17089 , \17090 , \17091 , \17092 ,
         \17093 , \17094 , \17095 , \17096 , \17097 , \17098 , \17099 , \17100 , \17101 , \17102 ,
         \17103 , \17104 , \17105 , \17106 , \17107 , \17108 , \17109 , \17110 , \17111 , \17112 ,
         \17113 , \17114 , \17115 , \17116 , \17117 , \17118 , \17119 , \17120 , \17121 , \17122 ,
         \17123 , \17124 , \17125 , \17126 , \17127 , \17128 , \17129 , \17130 , \17131 , \17132 ,
         \17133 , \17134 , \17135 , \17136 , \17137 , \17138 , \17139 , \17140 , \17141 , \17142 ,
         \17143 , \17144 , \17145 , \17146 , \17147 , \17148 , \17149 , \17150 , \17151 , \17152 ,
         \17153 , \17154 , \17155 , \17156 , \17157 , \17158 , \17159 , \17160 , \17161 , \17162 ,
         \17163 , \17164 , \17165 , \17166 , \17167 , \17168 , \17169 , \17170 , \17171 , \17172 ,
         \17173 , \17174 , \17175 , \17176 , \17177 , \17178 , \17179 , \17180 , \17181 , \17182 ,
         \17183 , \17184 , \17185 , \17186 , \17187 , \17188 , \17189 , \17190 , \17191 , \17192 ,
         \17193 , \17194 , \17195 , \17196 , \17197 , \17198 , \17199 , \17200 , \17201 , \17202 ,
         \17203 , \17204 , \17205 , \17206 , \17207 , \17208 , \17209 , \17210 , \17211 , \17212 ,
         \17213 , \17214 , \17215 , \17216 , \17217 , \17218 , \17219 , \17220 , \17221 , \17222 ,
         \17223 , \17224 , \17225 , \17226 , \17227 , \17228 , \17229 , \17230 , \17231 , \17232 ,
         \17233 , \17234 , \17235 , \17236 , \17237 , \17238 , \17239 , \17240 , \17241 , \17242 ,
         \17243 , \17244 , \17245 , \17246 , \17247 , \17248 , \17249 , \17250 , \17251 , \17252 ,
         \17253 , \17254 , \17255 , \17256 , \17257 , \17258 , \17259 , \17260 , \17261 , \17262 ,
         \17263 , \17264 , \17265 , \17266 , \17267 , \17268 , \17269 , \17270 , \17271 , \17272 ,
         \17273 , \17274 , \17275 , \17276 , \17277 , \17278 , \17279 , \17280 , \17281 , \17282 ,
         \17283 , \17284 , \17285 , \17286 , \17287 , \17288 , \17289 , \17290 , \17291 , \17292 ,
         \17293 , \17294 , \17295 , \17296 , \17297 , \17298 , \17299 , \17300 , \17301 , \17302 ,
         \17303 , \17304 , \17305 , \17306 , \17307 , \17308 , \17309 , \17310 , \17311 , \17312 ,
         \17313 , \17314 , \17315 , \17316 , \17317 , \17318 , \17319 , \17320 , \17321 , \17322 ,
         \17323 , \17324 , \17325 , \17326 , \17327 , \17328 , \17329 , \17330 , \17331 , \17332 ,
         \17333 , \17334 , \17335 , \17336 , \17337 , \17338 , \17339 , \17340 , \17341 , \17342 ,
         \17343 , \17344 , \17345 , \17346 , \17347 , \17348 , \17349 , \17350 , \17351 , \17352 ,
         \17353 , \17354 , \17355 , \17356 , \17357 , \17358 , \17359 , \17360 , \17361 , \17362 ,
         \17363 , \17364 , \17365 , \17366 , \17367 , \17368 , \17369 , \17370 , \17371 , \17372 ,
         \17373 , \17374 , \17375 , \17376 , \17377 , \17378 , \17379 , \17380 , \17381 , \17382 ,
         \17383 , \17384 , \17385 , \17386 , \17387 , \17388 , \17389 , \17390 , \17391 , \17392 ,
         \17393 , \17394 , \17395 , \17396 , \17397 , \17398 , \17399 , \17400 , \17401 , \17402 ,
         \17403 , \17404 , \17405 , \17406 , \17407 , \17408 , \17409 , \17410 , \17411 , \17412 ,
         \17413 , \17414 , \17415 , \17416 , \17417 , \17418 , \17419 , \17420 , \17421 , \17422 ,
         \17423 , \17424 , \17425 , \17426 , \17427 , \17428 , \17429 , \17430 , \17431 , \17432 ,
         \17433 , \17434 , \17435 , \17436 , \17437 , \17438 , \17439 , \17440 , \17441 , \17442 ,
         \17443 , \17444 , \17445 , \17446 , \17447 , \17448 , \17449 , \17450 , \17451 , \17452 ,
         \17453 , \17454 , \17455 , \17456 , \17457 , \17458 , \17459 , \17460 , \17461 , \17462 ,
         \17463 , \17464 , \17465 , \17466 , \17467 , \17468 , \17469 , \17470 , \17471 , \17472 ,
         \17473 , \17474 , \17475 , \17476 , \17477 , \17478 , \17479 , \17480 , \17481 , \17482 ,
         \17483 , \17484 , \17485 , \17486 , \17487 , \17488 , \17489 , \17490 , \17491 , \17492 ,
         \17493 , \17494 , \17495 , \17496 , \17497 , \17498 , \17499 , \17500 , \17501 , \17502 ,
         \17503 , \17504 , \17505 , \17506 , \17507 , \17508 , \17509 , \17510 , \17511 , \17512 ,
         \17513 , \17514 , \17515 , \17516 , \17517 , \17518 , \17519 , \17520 , \17521 , \17522 ,
         \17523 , \17524 , \17525 , \17526 , \17527 , \17528 , \17529 , \17530 , \17531 , \17532 ,
         \17533 , \17534 , \17535 , \17536 , \17537 , \17538 , \17539 , \17540 , \17541 , \17542 ,
         \17543 , \17544 , \17545 , \17546 , \17547 , \17548 , \17549 , \17550 , \17551 , \17552 ,
         \17553 , \17554 , \17555 , \17556 , \17557 , \17558 , \17559 , \17560 , \17561 , \17562 ,
         \17563 , \17564 , \17565 , \17566 , \17567 , \17568 , \17569 , \17570 , \17571 , \17572 ,
         \17573 , \17574 , \17575 , \17576 , \17577 , \17578 , \17579 , \17580 , \17581 , \17582 ,
         \17583 , \17584 , \17585 , \17586 , \17587 , \17588 , \17589 , \17590 , \17591 , \17592 ,
         \17593 , \17594 , \17595 , \17596 , \17597 , \17598 , \17599 , \17600 , \17601 , \17602 ,
         \17603 , \17604 , \17605 , \17606 , \17607 , \17608 , \17609 , \17610 , \17611 , \17612 ,
         \17613 , \17614 , \17615 , \17616 , \17617 , \17618 , \17619 , \17620 , \17621 , \17622 ,
         \17623 , \17624 , \17625 , \17626 , \17627 , \17628 , \17629 , \17630 , \17631 , \17632 ,
         \17633 , \17634 , \17635 , \17636 , \17637 , \17638 , \17639 , \17640 , \17641 , \17642 ,
         \17643 , \17644 , \17645 , \17646 , \17647 , \17648 , \17649 , \17650 , \17651 , \17652 ,
         \17653 , \17654 , \17655 , \17656 , \17657 , \17658 , \17659 , \17660 , \17661 , \17662 ,
         \17663 , \17664 , \17665 , \17666 , \17667 , \17668 , \17669 , \17670 , \17671 , \17672 ,
         \17673 , \17674 , \17675 , \17676 , \17677 , \17678 , \17679 , \17680 , \17681 , \17682 ,
         \17683 , \17684 , \17685 , \17686 , \17687 , \17688 , \17689 , \17690 , \17691 , \17692 ,
         \17693 , \17694 , \17695 , \17696 , \17697 , \17698 , \17699 , \17700 , \17701 , \17702 ,
         \17703 , \17704 , \17705 , \17706 , \17707 , \17708 , \17709 , \17710 , \17711 , \17712 ,
         \17713 , \17714 , \17715 , \17716 , \17717 , \17718 , \17719 , \17720 , \17721 , \17722 ,
         \17723 , \17724 , \17725 , \17726 , \17727 , \17728 , \17729 , \17730 , \17731 , \17732 ,
         \17733 , \17734 , \17735 , \17736 , \17737 , \17738 , \17739 , \17740 , \17741 , \17742 ,
         \17743 , \17744 , \17745 , \17746 , \17747 , \17748 , \17749 , \17750 , \17751 , \17752 ,
         \17753 , \17754 , \17755 , \17756 , \17757 , \17758 , \17759 , \17760 , \17761 , \17762 ,
         \17763 , \17764 , \17765 , \17766 , \17767 , \17768 , \17769 , \17770 , \17771 , \17772 ,
         \17773 , \17774 , \17775 , \17776 , \17777 , \17778 , \17779 , \17780 , \17781 , \17782 ,
         \17783 , \17784 , \17785 , \17786 , \17787 , \17788 , \17789 , \17790 , \17791 , \17792 ,
         \17793 , \17794 , \17795 , \17796 , \17797 , \17798 , \17799 , \17800 , \17801 , \17802 ,
         \17803 , \17804 , \17805 , \17806 , \17807 , \17808 , \17809 , \17810 , \17811 , \17812 ,
         \17813 , \17814 , \17815 , \17816 , \17817 , \17818 , \17819 , \17820 , \17821 , \17822 ,
         \17823 , \17824 , \17825 , \17826 , \17827 , \17828 , \17829 , \17830 , \17831 , \17832 ,
         \17833 , \17834 , \17835 , \17836 , \17837 , \17838 , \17839 , \17840 , \17841 , \17842 ,
         \17843 , \17844 , \17845 , \17846 , \17847 , \17848 , \17849 , \17850 , \17851 , \17852 ,
         \17853 , \17854 , \17855 , \17856 , \17857 , \17858 , \17859 , \17860 , \17861 , \17862 ,
         \17863 , \17864 , \17865 , \17866 , \17867 , \17868 , \17869 , \17870 , \17871 , \17872 ,
         \17873 , \17874 , \17875 , \17876 , \17877 , \17878 , \17879 , \17880 , \17881 , \17882 ,
         \17883 , \17884 , \17885 , \17886 , \17887 , \17888 , \17889 , \17890 , \17891 , \17892 ,
         \17893 , \17894 , \17895 , \17896 , \17897 , \17898 , \17899 , \17900 , \17901 , \17902 ,
         \17903 , \17904 , \17905 , \17906 , \17907 , \17908 , \17909 , \17910 , \17911 , \17912 ,
         \17913 , \17914 , \17915 , \17916 , \17917 , \17918 , \17919 , \17920 , \17921 , \17922 ,
         \17923 , \17924 , \17925 , \17926 , \17927 , \17928 , \17929 , \17930 , \17931 , \17932 ,
         \17933 , \17934 , \17935 , \17936 , \17937 , \17938 , \17939 , \17940 , \17941 , \17942 ,
         \17943 , \17944 , \17945 , \17946 , \17947 , \17948 , \17949 , \17950 , \17951 , \17952 ,
         \17953 , \17954 , \17955 , \17956 , \17957 , \17958 , \17959 , \17960 , \17961 , \17962 ,
         \17963 , \17964 , \17965 , \17966 , \17967 , \17968 , \17969 , \17970 , \17971 , \17972 ,
         \17973 , \17974 , \17975 , \17976 , \17977 , \17978 , \17979 , \17980 , \17981 , \17982 ,
         \17983 , \17984 , \17985 , \17986 , \17987 , \17988 , \17989 , \17990 , \17991 , \17992 ,
         \17993 , \17994 , \17995 , \17996 , \17997 , \17998 , \17999 , \18000 , \18001 , \18002 ,
         \18003 , \18004 , \18005 , \18006 , \18007 , \18008 , \18009 , \18010 , \18011 , \18012 ,
         \18013 , \18014 , \18015 , \18016 , \18017 , \18018 , \18019 , \18020 , \18021 , \18022 ,
         \18023 , \18024 , \18025 , \18026 , \18027 , \18028 , \18029 , \18030 , \18031 , \18032 ,
         \18033 , \18034 , \18035 , \18036 , \18037 , \18038 , \18039 , \18040 , \18041 , \18042 ,
         \18043 , \18044 , \18045 , \18046 , \18047 , \18048 , \18049 , \18050 , \18051 , \18052 ,
         \18053 , \18054 , \18055 , \18056 , \18057 , \18058 , \18059 , \18060 , \18061 , \18062 ,
         \18063 , \18064 , \18065 , \18066 , \18067 , \18068 , \18069 , \18070 , \18071 , \18072 ,
         \18073 , \18074 , \18075 , \18076 , \18077 , \18078 , \18079 , \18080 , \18081 , \18082 ,
         \18083 , \18084 , \18085 , \18086 , \18087 , \18088 , \18089 , \18090 , \18091 , \18092 ,
         \18093 , \18094 , \18095 , \18096 , \18097 , \18098 , \18099 , \18100 , \18101 , \18102 ,
         \18103 , \18104 , \18105 , \18106 , \18107 , \18108 , \18109 , \18110 , \18111 , \18112 ,
         \18113 , \18114 , \18115 , \18116 , \18117 , \18118 , \18119 , \18120 , \18121 , \18122 ,
         \18123 , \18124 , \18125 , \18126 , \18127 , \18128 , \18129 , \18130 , \18131 , \18132 ,
         \18133 , \18134 , \18135 , \18136 , \18137 , \18138 , \18139 , \18140 , \18141 , \18142 ,
         \18143 , \18144 , \18145 , \18146 , \18147 , \18148 , \18149 , \18150 , \18151 , \18152 ,
         \18153 , \18154 , \18155 , \18156 , \18157 , \18158 , \18159 , \18160 , \18161 , \18162 ,
         \18163 , \18164 , \18165 , \18166 , \18167 , \18168 , \18169 , \18170 , \18171 , \18172 ,
         \18173 , \18174 , \18175 , \18176 , \18177 , \18178 , \18179 , \18180 , \18181 , \18182 ,
         \18183 , \18184 , \18185 , \18186 , \18187 , \18188 , \18189 , \18190 , \18191 , \18192 ,
         \18193 , \18194 , \18195 , \18196 , \18197 , \18198 , \18199 , \18200 , \18201 , \18202 ,
         \18203 , \18204 , \18205 , \18206 , \18207 , \18208 , \18209 , \18210 , \18211 , \18212 ,
         \18213 , \18214 , \18215 , \18216 , \18217 , \18218 , \18219 , \18220 , \18221 , \18222 ,
         \18223 , \18224 , \18225 , \18226 , \18227 , \18228 , \18229 , \18230 , \18231 , \18232 ,
         \18233 , \18234 , \18235 , \18236 , \18237 , \18238 , \18239 , \18240 , \18241 , \18242 ,
         \18243 , \18244 , \18245 , \18246 , \18247 , \18248 , \18249 , \18250 , \18251 , \18252 ,
         \18253 , \18254 , \18255 , \18256 , \18257 , \18258 , \18259 , \18260 , \18261 , \18262 ,
         \18263 , \18264 , \18265 , \18266 , \18267 , \18268 , \18269 , \18270 , \18271 , \18272 ,
         \18273 , \18274 , \18275 , \18276 , \18277 , \18278 , \18279 , \18280 , \18281 , \18282 ,
         \18283 , \18284 , \18285 , \18286 , \18287 , \18288 , \18289 , \18290 , \18291 , \18292 ,
         \18293 , \18294 , \18295 , \18296 , \18297 , \18298 , \18299 , \18300 , \18301 , \18302 ,
         \18303 , \18304 , \18305 , \18306 , \18307 , \18308 , \18309 , \18310 , \18311 , \18312 ,
         \18313 , \18314 , \18315 , \18316 , \18317 , \18318 , \18319 , \18320 , \18321 , \18322 ,
         \18323 , \18324 , \18325 , \18326 , \18327 , \18328 , \18329 , \18330 , \18331 , \18332 ,
         \18333 , \18334 , \18335 , \18336 , \18337 , \18338 , \18339 , \18340 , \18341 , \18342 ,
         \18343 , \18344 , \18345 , \18346 , \18347 , \18348 , \18349 , \18350 , \18351 , \18352 ,
         \18353 , \18354 , \18355 , \18356 , \18357 , \18358 , \18359 , \18360 , \18361 , \18362 ,
         \18363 , \18364 , \18365 , \18366 , \18367 , \18368 , \18369 , \18370 , \18371 , \18372 ,
         \18373 , \18374 , \18375 , \18376 , \18377 , \18378 , \18379 , \18380 , \18381 , \18382 ,
         \18383 , \18384 , \18385 , \18386 , \18387 , \18388 , \18389 , \18390 , \18391 , \18392 ,
         \18393 , \18394 , \18395 , \18396 , \18397 , \18398 , \18399 , \18400 , \18401 , \18402 ,
         \18403 , \18404 , \18405 , \18406 , \18407 , \18408 , \18409 , \18410 , \18411 , \18412 ,
         \18413 , \18414 , \18415 , \18416 , \18417 , \18418 , \18419 , \18420 , \18421 , \18422 ,
         \18423 , \18424 , \18425 , \18426 , \18427 , \18428 , \18429 , \18430 , \18431 , \18432 ,
         \18433 , \18434 , \18435 , \18436 , \18437 , \18438 , \18439 , \18440 , \18441 , \18442 ,
         \18443 , \18444 , \18445 , \18446 , \18447 , \18448 , \18449 , \18450 , \18451 , \18452 ,
         \18453 , \18454 , \18455 , \18456 , \18457 , \18458 , \18459 , \18460 , \18461 , \18462 ,
         \18463 , \18464 , \18465 , \18466 , \18467 , \18468 , \18469 , \18470 , \18471 , \18472 ,
         \18473 , \18474 , \18475 , \18476 , \18477 , \18478 , \18479 , \18480 , \18481 , \18482 ,
         \18483 , \18484 , \18485 , \18486 , \18487 , \18488 , \18489 , \18490 , \18491 , \18492 ,
         \18493 , \18494 , \18495 , \18496 , \18497 , \18498 , \18499 , \18500 , \18501 , \18502 ,
         \18503 , \18504 , \18505 , \18506 , \18507 , \18508 , \18509 , \18510 , \18511 , \18512 ,
         \18513 , \18514 , \18515 , \18516 , \18517 , \18518 , \18519 , \18520 , \18521 , \18522 ,
         \18523 , \18524 , \18525 , \18526 , \18527 , \18528 , \18529 , \18530 , \18531 , \18532 ,
         \18533 , \18534 , \18535 , \18536 , \18537 , \18538 , \18539 , \18540 , \18541 , \18542 ,
         \18543 , \18544 , \18545 , \18546 , \18547 , \18548 , \18549 , \18550 , \18551 , \18552 ,
         \18553 , \18554 , \18555 , \18556 , \18557 , \18558 , \18559 , \18560 , \18561 , \18562 ,
         \18563 , \18564 , \18565 , \18566 , \18567 , \18568 , \18569 , \18570 , \18571 , \18572 ,
         \18573 , \18574 , \18575 , \18576 , \18577 , \18578 , \18579 , \18580 , \18581 , \18582 ,
         \18583 , \18584 , \18585 , \18586 , \18587 , \18588 , \18589 , \18590 , \18591 , \18592 ,
         \18593 , \18594 , \18595 , \18596 , \18597 , \18598 , \18599 , \18600 , \18601 , \18602 ,
         \18603 , \18604 , \18605 , \18606 , \18607 , \18608 , \18609 , \18610 , \18611 , \18612 ,
         \18613 , \18614 , \18615 , \18616 , \18617 , \18618 , \18619 , \18620 , \18621 , \18622 ,
         \18623 , \18624 , \18625 , \18626 , \18627 , \18628 , \18629 , \18630 , \18631 , \18632 ,
         \18633 , \18634 , \18635 , \18636 , \18637 , \18638 , \18639 , \18640 , \18641 , \18642 ,
         \18643 , \18644 , \18645 , \18646 , \18647 , \18648 , \18649 , \18650 , \18651 , \18652 ,
         \18653 , \18654 , \18655 , \18656 , \18657 , \18658 , \18659 , \18660 , \18661 , \18662 ,
         \18663 , \18664 , \18665 , \18666 , \18667 , \18668 , \18669 , \18670 , \18671 , \18672 ,
         \18673 , \18674 , \18675 , \18676 , \18677 , \18678 , \18679 , \18680 , \18681 , \18682 ,
         \18683 , \18684 , \18685 , \18686 , \18687 , \18688 , \18689 , \18690 , \18691 , \18692 ,
         \18693 , \18694 , \18695 , \18696 , \18697 , \18698 , \18699 , \18700 , \18701 , \18702 ,
         \18703 , \18704 , \18705 , \18706 , \18707 , \18708 , \18709 , \18710 , \18711 , \18712 ,
         \18713 , \18714 , \18715 , \18716 , \18717 , \18718 , \18719 , \18720 , \18721 , \18722 ,
         \18723 , \18724 , \18725 , \18726 , \18727 , \18728 , \18729 , \18730 , \18731 , \18732 ,
         \18733 , \18734 , \18735 , \18736 , \18737 , \18738 , \18739 , \18740 , \18741 , \18742 ,
         \18743 , \18744 , \18745 , \18746 , \18747 , \18748 , \18749 , \18750 , \18751 , \18752 ,
         \18753 , \18754 , \18755 , \18756 , \18757 , \18758 , \18759 , \18760 , \18761 , \18762 ,
         \18763 , \18764 , \18765 , \18766 , \18767 , \18768 , \18769 , \18770 , \18771 , \18772 ,
         \18773 , \18774 , \18775 , \18776 , \18777 , \18778 , \18779 , \18780 , \18781 , \18782 ,
         \18783 , \18784 , \18785 , \18786 , \18787 , \18788 , \18789 , \18790 , \18791 , \18792 ,
         \18793 , \18794 , \18795 , \18796 , \18797 , \18798 , \18799 , \18800 , \18801 , \18802 ,
         \18803 , \18804 , \18805 , \18806 , \18807 , \18808 , \18809 , \18810 , \18811 , \18812 ,
         \18813 , \18814 , \18815 , \18816 , \18817 , \18818 , \18819 , \18820 , \18821 , \18822 ,
         \18823 , \18824 , \18825 , \18826 , \18827 , \18828 , \18829 , \18830 , \18831 , \18832 ,
         \18833 , \18834 , \18835 , \18836 , \18837 , \18838 , \18839 , \18840 , \18841 , \18842 ,
         \18843 , \18844 , \18845 , \18846 , \18847 , \18848 , \18849 , \18850 , \18851 , \18852 ,
         \18853 , \18854 , \18855 , \18856 , \18857 , \18858 , \18859 , \18860 , \18861 , \18862 ,
         \18863 , \18864 , \18865 , \18866 , \18867 , \18868 , \18869 , \18870 , \18871 , \18872 ,
         \18873 , \18874 , \18875 , \18876 , \18877 , \18878 , \18879 , \18880 , \18881 , \18882 ,
         \18883 , \18884 , \18885 , \18886 , \18887 , \18888 , \18889 , \18890 , \18891 , \18892 ,
         \18893 , \18894 , \18895 , \18896 , \18897 , \18898 , \18899 , \18900 , \18901 , \18902 ,
         \18903 , \18904 , \18905 , \18906 , \18907 , \18908 , \18909 , \18910 , \18911 , \18912 ,
         \18913 , \18914 , \18915 , \18916 , \18917 , \18918 , \18919 , \18920 , \18921 , \18922 ,
         \18923 , \18924 , \18925 , \18926 , \18927 , \18928 , \18929 , \18930 , \18931 , \18932 ,
         \18933 , \18934 , \18935 , \18936 , \18937 , \18938 , \18939 , \18940 , \18941 , \18942 ,
         \18943 , \18944 , \18945 , \18946 , \18947 , \18948 , \18949 , \18950 , \18951 , \18952 ,
         \18953 , \18954 , \18955 , \18956 , \18957 , \18958 , \18959 , \18960 , \18961 , \18962 ,
         \18963 , \18964 , \18965 , \18966 , \18967 , \18968 , \18969 , \18970 , \18971 , \18972 ,
         \18973 , \18974 , \18975 , \18976 , \18977 , \18978 , \18979 , \18980 , \18981 , \18982 ,
         \18983 , \18984 , \18985 , \18986 , \18987 , \18988 , \18989 , \18990 , \18991 , \18992 ,
         \18993 , \18994 , \18995 , \18996 , \18997 , \18998 , \18999 , \19000 , \19001 , \19002 ,
         \19003 , \19004 , \19005 , \19006 , \19007 , \19008 , \19009 , \19010 , \19011 , \19012 ,
         \19013 , \19014 , \19015 , \19016 , \19017 , \19018 , \19019 , \19020 , \19021 , \19022 ,
         \19023 , \19024 , \19025 , \19026 , \19027 , \19028 , \19029 , \19030 , \19031 , \19032 ,
         \19033 , \19034 , \19035 , \19036 , \19037 , \19038 , \19039 , \19040 , \19041 , \19042 ,
         \19043 , \19044 , \19045 , \19046 , \19047 , \19048 , \19049 , \19050 , \19051 , \19052 ,
         \19053 , \19054 , \19055 , \19056 , \19057 , \19058 , \19059 , \19060 , \19061 , \19062 ,
         \19063 , \19064 , \19065 , \19066 , \19067 , \19068 , \19069 , \19070 , \19071 , \19072 ,
         \19073 , \19074 , \19075 , \19076 , \19077 , \19078 , \19079 , \19080 , \19081 , \19082 ,
         \19083 , \19084 , \19085 , \19086 , \19087 , \19088 , \19089 , \19090 , \19091 , \19092 ,
         \19093 , \19094 , \19095 , \19096 , \19097 , \19098 , \19099 , \19100 , \19101 , \19102 ,
         \19103 , \19104 , \19105 , \19106 , \19107 , \19108 , \19109 , \19110 , \19111 , \19112 ,
         \19113 , \19114 , \19115 , \19116 , \19117 , \19118 , \19119 , \19120 , \19121 , \19122 ,
         \19123 , \19124 , \19125 , \19126 , \19127 , \19128 , \19129 , \19130 , \19131 , \19132 ,
         \19133 , \19134 , \19135 , \19136 , \19137 , \19138 , \19139 , \19140 , \19141 , \19142 ,
         \19143 , \19144 , \19145 , \19146 , \19147 , \19148 , \19149 , \19150 , \19151 , \19152 ,
         \19153 , \19154 , \19155 , \19156 , \19157 , \19158 , \19159 , \19160 , \19161 , \19162 ,
         \19163 , \19164 , \19165 , \19166 , \19167 , \19168 , \19169 , \19170 , \19171 , \19172 ,
         \19173 , \19174 , \19175 , \19176 , \19177 , \19178 , \19179 , \19180 , \19181 , \19182 ,
         \19183 , \19184 , \19185 , \19186 , \19187 , \19188 , \19189 , \19190 , \19191 , \19192 ,
         \19193 , \19194 , \19195 , \19196 , \19197 , \19198 , \19199 , \19200 , \19201 , \19202 ,
         \19203 , \19204 , \19205 , \19206 , \19207 , \19208 , \19209 , \19210 , \19211 , \19212 ,
         \19213 , \19214 , \19215 , \19216 , \19217 , \19218 , \19219 , \19220 , \19221 , \19222 ,
         \19223 , \19224 , \19225 , \19226 , \19227 , \19228 , \19229 , \19230 , \19231 , \19232 ,
         \19233 , \19234 , \19235 , \19236 , \19237 , \19238 , \19239 , \19240 , \19241 , \19242 ,
         \19243 , \19244 , \19245 , \19246 , \19247 , \19248 , \19249 , \19250 , \19251 , \19252 ,
         \19253 , \19254 , \19255 , \19256 , \19257 , \19258 , \19259 , \19260 , \19261 , \19262 ,
         \19263 , \19264 , \19265 , \19266 , \19267 , \19268 , \19269 , \19270 , \19271 , \19272 ,
         \19273 , \19274 , \19275 , \19276 , \19277 , \19278 , \19279 , \19280 , \19281 , \19282 ,
         \19283 , \19284 , \19285 , \19286 , \19287 , \19288 , \19289 , \19290 , \19291 , \19292 ,
         \19293 , \19294 , \19295 , \19296 , \19297 , \19298 , \19299 , \19300 , \19301 , \19302 ,
         \19303 , \19304 , \19305 , \19306 , \19307 , \19308 , \19309 , \19310 , \19311 , \19312 ,
         \19313 , \19314 , \19315 , \19316 , \19317 , \19318 , \19319 , \19320 , \19321 , \19322 ,
         \19323 , \19324 , \19325 , \19326 , \19327 , \19328 , \19329 , \19330 , \19331 , \19332 ,
         \19333 , \19334 , \19335 , \19336 , \19337 , \19338 , \19339 , \19340 , \19341 , \19342 ,
         \19343 , \19344 , \19345 , \19346 , \19347 , \19348 , \19349 , \19350 , \19351 , \19352 ,
         \19353 , \19354 , \19355 , \19356 , \19357 , \19358 , \19359 , \19360 , \19361 , \19362 ,
         \19363 , \19364 , \19365 , \19366 , \19367 , \19368 , \19369 , \19370 , \19371 , \19372 ,
         \19373 , \19374 , \19375 , \19376 , \19377 , \19378 , \19379 , \19380 , \19381 , \19382 ,
         \19383 , \19384 , \19385 , \19386 , \19387 , \19388 , \19389 , \19390 , \19391 , \19392 ,
         \19393 , \19394 , \19395 , \19396 , \19397 , \19398 , \19399 , \19400 , \19401 , \19402 ,
         \19403 , \19404 , \19405 , \19406 , \19407 , \19408 , \19409 , \19410 , \19411 , \19412 ,
         \19413 , \19414 , \19415 , \19416 , \19417 , \19418 , \19419 , \19420 , \19421 , \19422 ,
         \19423 , \19424 , \19425 , \19426 , \19427 , \19428 , \19429 , \19430 , \19431 , \19432 ,
         \19433 , \19434 , \19435 , \19436 , \19437 , \19438 , \19439 , \19440 , \19441 , \19442 ,
         \19443 , \19444 , \19445 , \19446 , \19447 , \19448 , \19449 , \19450 , \19451 , \19452 ,
         \19453 , \19454 , \19455 , \19456 , \19457 , \19458 , \19459 , \19460 , \19461 , \19462 ,
         \19463 , \19464 , \19465 , \19466 , \19467 , \19468 , \19469 , \19470 , \19471 , \19472 ,
         \19473 , \19474 , \19475 , \19476 , \19477 , \19478 , \19479 , \19480 , \19481 , \19482 ,
         \19483 , \19484 , \19485 , \19486 , \19487 , \19488 , \19489 , \19490 , \19491 , \19492 ,
         \19493 , \19494 , \19495 , \19496 , \19497 , \19498 , \19499 , \19500 , \19501 , \19502 ,
         \19503 , \19504 , \19505 , \19506 , \19507 , \19508 , \19509 , \19510 , \19511 , \19512 ,
         \19513 , \19514 , \19515 , \19516 , \19517 , \19518 , \19519 , \19520 , \19521 , \19522 ,
         \19523 , \19524 , \19525 , \19526 , \19527 , \19528 , \19529 , \19530 , \19531 , \19532 ,
         \19533 , \19534 , \19535 , \19536 , \19537 , \19538 , \19539 , \19540 , \19541 , \19542 ,
         \19543 , \19544 , \19545 , \19546 , \19547 , \19548 , \19549 , \19550 , \19551 , \19552 ,
         \19553 , \19554 , \19555 , \19556 , \19557 , \19558 , \19559 , \19560 , \19561 , \19562 ,
         \19563 , \19564 , \19565 , \19566 , \19567 , \19568 , \19569 , \19570 , \19571 , \19572 ,
         \19573 , \19574 , \19575 , \19576 , \19577 , \19578 , \19579 , \19580 , \19581 , \19582 ,
         \19583 , \19584 , \19585 , \19586 , \19587 , \19588 , \19589 , \19590 , \19591 , \19592 ,
         \19593 , \19594 , \19595 , \19596 , \19597 , \19598 , \19599 , \19600 , \19601 , \19602 ,
         \19603 , \19604 , \19605 , \19606 , \19607 , \19608 , \19609 , \19610 , \19611 , \19612 ,
         \19613 , \19614 , \19615 , \19616 , \19617 , \19618 , \19619 , \19620 , \19621 , \19622 ,
         \19623 , \19624 , \19625 , \19626 , \19627 , \19628 , \19629 , \19630 , \19631 , \19632 ,
         \19633 , \19634 , \19635 , \19636 , \19637 , \19638 , \19639 , \19640 , \19641 , \19642 ,
         \19643 , \19644 , \19645 , \19646 , \19647 , \19648 , \19649 , \19650 , \19651 , \19652 ,
         \19653 , \19654 , \19655 , \19656 , \19657 , \19658 , \19659 , \19660 , \19661 , \19662 ,
         \19663 , \19664 , \19665 , \19666 , \19667 , \19668 , \19669 , \19670 , \19671 , \19672 ,
         \19673 , \19674 , \19675 , \19676 , \19677 , \19678 , \19679 , \19680 , \19681 , \19682 ,
         \19683 , \19684 , \19685 , \19686 , \19687 , \19688 , \19689 , \19690 , \19691 , \19692 ,
         \19693 , \19694 , \19695 , \19696 , \19697 , \19698 , \19699 , \19700 , \19701 , \19702 ,
         \19703 , \19704 , \19705 , \19706 , \19707 , \19708 , \19709 , \19710 , \19711 , \19712 ,
         \19713 , \19714 , \19715 , \19716 , \19717 , \19718 , \19719 , \19720 , \19721 , \19722 ,
         \19723 , \19724 , \19725 , \19726 , \19727 , \19728 , \19729 , \19730 , \19731 , \19732 ,
         \19733 , \19734 , \19735 , \19736 , \19737 , \19738 , \19739 , \19740 , \19741 , \19742 ,
         \19743 , \19744 , \19745 , \19746 , \19747 , \19748 , \19749 , \19750 , \19751 , \19752 ,
         \19753 , \19754 , \19755 , \19756 , \19757 , \19758 , \19759 , \19760 , \19761 , \19762 ,
         \19763 , \19764 , \19765 , \19766 , \19767 , \19768 , \19769 , \19770 , \19771 , \19772 ,
         \19773 , \19774 , \19775 , \19776 , \19777 , \19778 , \19779 , \19780 , \19781 , \19782 ,
         \19783 , \19784 , \19785 , \19786 , \19787 , \19788 , \19789 , \19790 , \19791 , \19792 ,
         \19793 , \19794 , \19795 , \19796 , \19797 , \19798 , \19799 , \19800 , \19801 , \19802 ,
         \19803 , \19804 , \19805 , \19806 , \19807 , \19808 , \19809 , \19810 , \19811 , \19812 ,
         \19813 , \19814 , \19815 , \19816 , \19817 , \19818 , \19819 , \19820 , \19821 , \19822 ,
         \19823 , \19824 , \19825 , \19826 , \19827 , \19828 , \19829 , \19830 , \19831 , \19832 ,
         \19833 , \19834 , \19835 , \19836 , \19837 , \19838 , \19839 , \19840 , \19841 , \19842 ,
         \19843 , \19844 , \19845 , \19846 , \19847 , \19848 , \19849 , \19850 , \19851 , \19852 ,
         \19853 , \19854 , \19855 , \19856 , \19857 , \19858 , \19859 , \19860 , \19861 , \19862 ,
         \19863 , \19864 , \19865 , \19866 , \19867 , \19868 , \19869 , \19870 , \19871 , \19872 ,
         \19873 , \19874 , \19875 , \19876 , \19877 , \19878 , \19879 , \19880 , \19881 , \19882 ,
         \19883 , \19884 , \19885 , \19886 , \19887 , \19888 , \19889 , \19890 , \19891 , \19892 ,
         \19893 , \19894 , \19895 , \19896 , \19897 , \19898 , \19899 , \19900 , \19901 , \19902 ,
         \19903 , \19904 , \19905 , \19906 , \19907 , \19908 , \19909 , \19910 , \19911 , \19912 ,
         \19913 , \19914 , \19915 , \19916 , \19917 , \19918 , \19919 , \19920 , \19921 , \19922 ,
         \19923 , \19924 , \19925 , \19926 , \19927 , \19928 , \19929 , \19930 , \19931 , \19932 ,
         \19933 , \19934 , \19935 , \19936 , \19937 , \19938 , \19939 , \19940 , \19941 , \19942 ,
         \19943 , \19944 , \19945 , \19946 , \19947 , \19948 , \19949 , \19950 , \19951 , \19952 ,
         \19953 , \19954 , \19955 , \19956 , \19957 , \19958 , \19959 , \19960 , \19961 , \19962 ,
         \19963 , \19964 , \19965 , \19966 , \19967 , \19968 , \19969 , \19970 , \19971 , \19972 ,
         \19973 , \19974 , \19975 , \19976 , \19977 , \19978 , \19979 , \19980 , \19981 , \19982 ,
         \19983 , \19984 , \19985 , \19986 , \19987 , \19988 , \19989 , \19990 , \19991 , \19992 ,
         \19993 , \19994 , \19995 , \19996 , \19997 , \19998 , \19999 , \20000 , \20001 , \20002 ,
         \20003 , \20004 , \20005 , \20006 , \20007 , \20008 , \20009 , \20010 , \20011 , \20012 ,
         \20013 , \20014 , \20015 , \20016 , \20017 , \20018 , \20019 , \20020 , \20021 , \20022 ,
         \20023 , \20024 , \20025 , \20026 , \20027 , \20028 , \20029 , \20030 , \20031 , \20032 ,
         \20033 , \20034 , \20035 , \20036 , \20037 , \20038 , \20039 , \20040 , \20041 , \20042 ,
         \20043 , \20044 , \20045 , \20046 , \20047 , \20048 , \20049 , \20050 , \20051 , \20052 ,
         \20053 , \20054 , \20055 , \20056 , \20057 , \20058 , \20059 , \20060 , \20061 , \20062 ,
         \20063 , \20064 , \20065 , \20066 , \20067 , \20068 , \20069 , \20070 , \20071 , \20072 ,
         \20073 , \20074 , \20075 , \20076 , \20077 , \20078 , \20079 , \20080 , \20081 , \20082 ,
         \20083 , \20084 , \20085 , \20086 , \20087 , \20088 , \20089 , \20090 , \20091 , \20092 ,
         \20093 , \20094 , \20095 , \20096 , \20097 , \20098 , \20099 , \20100 , \20101 , \20102 ,
         \20103 , \20104 , \20105 , \20106 , \20107 , \20108 , \20109 , \20110 , \20111 , \20112 ,
         \20113 , \20114 , \20115 , \20116 , \20117 , \20118 , \20119 , \20120 , \20121 , \20122 ,
         \20123 , \20124 , \20125 , \20126 , \20127 , \20128 , \20129 , \20130 , \20131 , \20132 ,
         \20133 , \20134 , \20135 , \20136 , \20137 , \20138 , \20139 , \20140 , \20141 , \20142 ,
         \20143 , \20144 , \20145 , \20146 , \20147 , \20148 , \20149 , \20150 , \20151 , \20152 ,
         \20153 , \20154 , \20155 , \20156 , \20157 , \20158 , \20159 , \20160 , \20161 , \20162 ,
         \20163 , \20164 , \20165 , \20166 , \20167 , \20168 , \20169 , \20170 , \20171 , \20172 ,
         \20173 , \20174 , \20175 , \20176 , \20177 , \20178 , \20179 , \20180 , \20181 , \20182 ,
         \20183 , \20184 , \20185 , \20186 , \20187 , \20188 , \20189 , \20190 , \20191 , \20192 ,
         \20193 , \20194 , \20195 , \20196 , \20197 , \20198 , \20199 , \20200 , \20201 , \20202 ,
         \20203 , \20204 , \20205 , \20206 , \20207 , \20208 , \20209 , \20210 , \20211 , \20212 ,
         \20213 , \20214 , \20215 , \20216 , \20217 , \20218 , \20219 , \20220 , \20221 , \20222 ,
         \20223 , \20224 , \20225 , \20226 , \20227 , \20228 , \20229 , \20230 , \20231 , \20232 ,
         \20233 , \20234 , \20235 , \20236 , \20237 , \20238 , \20239 , \20240 , \20241 , \20242 ,
         \20243 , \20244 , \20245 , \20246 , \20247 , \20248 , \20249 , \20250 , \20251 , \20252 ,
         \20253 , \20254 , \20255 , \20256 , \20257 , \20258 , \20259 , \20260 , \20261 , \20262 ,
         \20263 , \20264 , \20265 , \20266 , \20267 , \20268 , \20269 , \20270 , \20271 , \20272 ,
         \20273 , \20274 , \20275 , \20276 , \20277 , \20278 , \20279 , \20280 , \20281 , \20282 ,
         \20283 , \20284 , \20285 , \20286 , \20287 , \20288 , \20289 , \20290 , \20291 , \20292 ,
         \20293 , \20294 , \20295 , \20296 , \20297 , \20298 , \20299 , \20300 , \20301 , \20302 ,
         \20303 , \20304 , \20305 , \20306 , \20307 , \20308 , \20309 , \20310 , \20311 , \20312 ,
         \20313 , \20314 , \20315 , \20316 , \20317 , \20318 , \20319 , \20320 , \20321 , \20322 ,
         \20323 , \20324 , \20325 , \20326 , \20327 , \20328 , \20329 , \20330 , \20331 , \20332 ,
         \20333 , \20334 , \20335 , \20336 , \20337 , \20338 , \20339 , \20340 , \20341 , \20342 ,
         \20343 , \20344 , \20345 , \20346 , \20347 , \20348 , \20349 , \20350 , \20351 , \20352 ,
         \20353 , \20354 , \20355 , \20356 , \20357 , \20358 , \20359 , \20360 , \20361 , \20362 ,
         \20363 , \20364 , \20365 , \20366 , \20367 , \20368 , \20369 , \20370 , \20371 , \20372 ,
         \20373 , \20374 , \20375 , \20376 , \20377 , \20378 , \20379 , \20380 , \20381 , \20382 ,
         \20383 , \20384 , \20385 , \20386 , \20387 , \20388 , \20389 , \20390 , \20391 , \20392 ,
         \20393 , \20394 , \20395 , \20396 , \20397 , \20398 , \20399 , \20400 , \20401 , \20402 ,
         \20403 , \20404 , \20405 , \20406 , \20407 , \20408 , \20409 , \20410 , \20411 , \20412 ,
         \20413 , \20414 , \20415 , \20416 , \20417 , \20418 , \20419 , \20420 , \20421 , \20422 ,
         \20423 , \20424 , \20425 , \20426 , \20427 , \20428 , \20429 , \20430 , \20431 , \20432 ,
         \20433 , \20434 , \20435 , \20436 , \20437 , \20438 , \20439 , \20440 , \20441 , \20442 ,
         \20443 , \20444 , \20445 , \20446 , \20447 , \20448 , \20449 , \20450 , \20451 , \20452 ,
         \20453 , \20454 , \20455 , \20456 , \20457 , \20458 , \20459 , \20460 , \20461 , \20462 ,
         \20463 , \20464 , \20465 , \20466 , \20467 , \20468 , \20469 , \20470 , \20471 , \20472 ,
         \20473 , \20474 , \20475 , \20476 , \20477 , \20478 , \20479 , \20480 , \20481 , \20482 ,
         \20483 , \20484 , \20485 , \20486 , \20487 , \20488 , \20489 , \20490 , \20491 , \20492 ,
         \20493 , \20494 , \20495 , \20496 , \20497 , \20498 , \20499 , \20500 , \20501 , \20502 ,
         \20503 , \20504 , \20505 , \20506 , \20507 , \20508 , \20509 , \20510 , \20511 , \20512 ,
         \20513 , \20514 , \20515 , \20516 , \20517 , \20518 , \20519 , \20520 , \20521 , \20522 ,
         \20523 , \20524 , \20525 , \20526 , \20527 , \20528 , \20529 , \20530 , \20531 , \20532 ,
         \20533 , \20534 , \20535 , \20536 , \20537 , \20538 , \20539 , \20540 , \20541 , \20542 ,
         \20543 , \20544 , \20545 , \20546 , \20547 , \20548 , \20549 , \20550 , \20551 , \20552 ,
         \20553 , \20554 , \20555 , \20556 , \20557 , \20558 , \20559 , \20560 , \20561 , \20562 ,
         \20563 , \20564 , \20565 , \20566 , \20567 , \20568 , \20569 , \20570 , \20571 , \20572 ,
         \20573 , \20574 , \20575 , \20576 , \20577 , \20578 , \20579 , \20580 , \20581 , \20582 ,
         \20583 , \20584 , \20585 , \20586 , \20587 , \20588 , \20589 , \20590 , \20591 , \20592 ,
         \20593 , \20594 , \20595 , \20596 , \20597 , \20598 , \20599 , \20600 , \20601 , \20602 ,
         \20603 , \20604 , \20605 , \20606 , \20607 , \20608 , \20609 , \20610 , \20611 , \20612 ,
         \20613 , \20614 , \20615 , \20616 , \20617 , \20618 , \20619 , \20620 , \20621 , \20622 ,
         \20623 , \20624 , \20625 , \20626 , \20627 , \20628 , \20629 , \20630 , \20631 , \20632 ,
         \20633 , \20634 , \20635 , \20636 , \20637 , \20638 , \20639 , \20640 , \20641 , \20642 ,
         \20643 , \20644 , \20645 , \20646 , \20647 , \20648 , \20649 , \20650 , \20651 , \20652 ,
         \20653 , \20654 , \20655 , \20656 , \20657 , \20658 , \20659 , \20660 , \20661 , \20662 ,
         \20663 , \20664 , \20665 , \20666 , \20667 , \20668 , \20669 , \20670 , \20671 , \20672 ,
         \20673 , \20674 , \20675 , \20676 , \20677 , \20678 , \20679 , \20680 , \20681 , \20682 ,
         \20683 , \20684 , \20685 , \20686 , \20687 , \20688 , \20689 , \20690 , \20691 , \20692 ,
         \20693 , \20694 , \20695 , \20696 , \20697 , \20698 , \20699 , \20700 , \20701 , \20702 ,
         \20703 , \20704 , \20705 , \20706 , \20707 , \20708 , \20709 , \20710 , \20711 , \20712 ,
         \20713 , \20714 , \20715 , \20716 , \20717 , \20718 , \20719 , \20720 , \20721 , \20722 ,
         \20723 , \20724 , \20725 , \20726 , \20727 , \20728 , \20729 , \20730 , \20731 , \20732 ,
         \20733 , \20734 , \20735 , \20736 , \20737 , \20738 , \20739 , \20740 , \20741 , \20742 ,
         \20743 , \20744 , \20745 , \20746 , \20747 , \20748 , \20749 , \20750 , \20751 , \20752 ,
         \20753 , \20754 , \20755 , \20756 , \20757 , \20758 , \20759 , \20760 , \20761 , \20762 ,
         \20763 , \20764 , \20765 , \20766 , \20767 , \20768 , \20769 , \20770 , \20771 , \20772 ,
         \20773 , \20774 , \20775 , \20776 , \20777 , \20778 , \20779 , \20780 , \20781 , \20782 ,
         \20783 , \20784 , \20785 , \20786 , \20787 , \20788 , \20789 , \20790 , \20791 , \20792 ,
         \20793 , \20794 , \20795 , \20796 , \20797 , \20798 , \20799 , \20800 , \20801 , \20802 ,
         \20803 , \20804 , \20805 , \20806 , \20807 , \20808 , \20809 , \20810 , \20811 , \20812 ,
         \20813 , \20814 , \20815 , \20816 , \20817 , \20818 , \20819 , \20820 , \20821 , \20822 ,
         \20823 , \20824 , \20825 , \20826 , \20827 , \20828 , \20829 , \20830 , \20831 , \20832 ,
         \20833 , \20834 , \20835 , \20836 , \20837 , \20838 , \20839 , \20840 , \20841 , \20842 ,
         \20843 , \20844 , \20845 , \20846 , \20847 , \20848 , \20849 , \20850 , \20851 , \20852 ,
         \20853 , \20854 , \20855 , \20856 , \20857 , \20858 , \20859 , \20860 , \20861 , \20862 ,
         \20863 , \20864 , \20865 , \20866 , \20867 , \20868 , \20869 , \20870 , \20871 , \20872 ,
         \20873 , \20874 , \20875 , \20876 , \20877 , \20878 , \20879 , \20880 , \20881 , \20882 ,
         \20883 , \20884 , \20885 , \20886 , \20887 , \20888 , \20889 , \20890 , \20891 , \20892 ,
         \20893 , \20894 , \20895 , \20896 , \20897 , \20898 , \20899 , \20900 , \20901 , \20902 ,
         \20903 , \20904 , \20905 , \20906 , \20907 , \20908 , \20909 , \20910 , \20911 , \20912 ,
         \20913 , \20914 , \20915 , \20916 , \20917 , \20918 , \20919 , \20920 , \20921 , \20922 ,
         \20923 , \20924 , \20925 , \20926 , \20927 , \20928 , \20929 , \20930 , \20931 , \20932 ,
         \20933 , \20934 , \20935 , \20936 , \20937 , \20938 , \20939 , \20940 , \20941 , \20942 ,
         \20943 , \20944 , \20945 , \20946 , \20947 , \20948 , \20949 , \20950 , \20951 , \20952 ,
         \20953 , \20954 , \20955 , \20956 , \20957 , \20958 , \20959 , \20960 , \20961 , \20962 ,
         \20963 , \20964 , \20965 , \20966 , \20967 , \20968 , \20969 , \20970 , \20971 , \20972 ,
         \20973 , \20974 , \20975 , \20976 , \20977 , \20978 , \20979 , \20980 , \20981 , \20982 ,
         \20983 , \20984 , \20985 , \20986 , \20987 , \20988 , \20989 , \20990 , \20991 , \20992 ,
         \20993 , \20994 , \20995 , \20996 , \20997 , \20998 , \20999 , \21000 , \21001 , \21002 ,
         \21003 , \21004 , \21005 , \21006 , \21007 , \21008 , \21009 , \21010 , \21011 , \21012 ,
         \21013 , \21014 , \21015 , \21016 , \21017 , \21018 , \21019 , \21020 , \21021 , \21022 ,
         \21023 , \21024 , \21025 , \21026 , \21027 , \21028 , \21029 , \21030 , \21031 , \21032 ,
         \21033 , \21034 , \21035 , \21036 , \21037 , \21038 , \21039 , \21040 , \21041 , \21042 ,
         \21043 , \21044 , \21045 , \21046 , \21047 , \21048 , \21049 , \21050 , \21051 , \21052 ,
         \21053 , \21054 , \21055 , \21056 , \21057 , \21058 , \21059 , \21060 , \21061 , \21062 ,
         \21063 , \21064 , \21065 , \21066 , \21067 , \21068 , \21069 , \21070 , \21071 , \21072 ,
         \21073 , \21074 , \21075 , \21076 , \21077 , \21078 , \21079 , \21080 , \21081 , \21082 ,
         \21083 , \21084 , \21085 , \21086 , \21087 , \21088 , \21089 , \21090 , \21091 , \21092 ,
         \21093 , \21094 , \21095 , \21096 , \21097 , \21098 , \21099 , \21100 , \21101 , \21102 ,
         \21103 , \21104 , \21105 , \21106 , \21107 , \21108 , \21109 , \21110 , \21111 , \21112 ,
         \21113 , \21114 , \21115 , \21116 , \21117 , \21118 , \21119 , \21120 , \21121 , \21122 ,
         \21123 , \21124 , \21125 , \21126 , \21127 , \21128 , \21129 , \21130 , \21131 , \21132 ,
         \21133 , \21134 , \21135 , \21136 , \21137 , \21138 , \21139 , \21140 , \21141 , \21142 ,
         \21143 , \21144 , \21145 , \21146 , \21147 , \21148 , \21149 , \21150 , \21151 , \21152 ,
         \21153 , \21154 , \21155 , \21156 , \21157 , \21158 , \21159 , \21160 , \21161 , \21162 ,
         \21163 , \21164 , \21165 , \21166 , \21167 , \21168 , \21169 , \21170 , \21171 , \21172 ,
         \21173 , \21174 , \21175 , \21176 , \21177 , \21178 , \21179 , \21180 , \21181 , \21182 ,
         \21183 , \21184 , \21185 , \21186 , \21187 , \21188 , \21189 , \21190 , \21191 , \21192 ,
         \21193 , \21194 , \21195 , \21196 , \21197 , \21198 , \21199 , \21200 , \21201 , \21202 ,
         \21203 , \21204 , \21205 , \21206 , \21207 , \21208 , \21209 , \21210 , \21211 , \21212 ,
         \21213 , \21214 , \21215 , \21216 , \21217 , \21218 , \21219 , \21220 , \21221 , \21222 ,
         \21223 , \21224 , \21225 , \21226 , \21227 , \21228 , \21229 , \21230 , \21231 , \21232 ,
         \21233 , \21234 , \21235 , \21236 , \21237 , \21238 , \21239 , \21240 , \21241 , \21242 ,
         \21243 , \21244 , \21245 , \21246 , \21247 , \21248 , \21249 , \21250 , \21251 , \21252 ,
         \21253 , \21254 , \21255 , \21256 , \21257 , \21258 , \21259 , \21260 , \21261 , \21262 ,
         \21263 , \21264 , \21265 , \21266 , \21267 , \21268 , \21269 , \21270 , \21271 , \21272 ,
         \21273 , \21274 , \21275 , \21276 , \21277 , \21278 , \21279 , \21280 , \21281 , \21282 ,
         \21283 , \21284 , \21285 , \21286 , \21287 , \21288 , \21289 , \21290 , \21291 , \21292 ,
         \21293 , \21294 , \21295 , \21296 , \21297 , \21298 , \21299 , \21300 , \21301 , \21302 ,
         \21303 , \21304 , \21305 , \21306 , \21307 , \21308 , \21309 , \21310 , \21311 , \21312 ,
         \21313 , \21314 , \21315 , \21316 , \21317 , \21318 , \21319 , \21320 , \21321 , \21322 ,
         \21323 , \21324 , \21325 , \21326 , \21327 , \21328 , \21329 , \21330 , \21331 , \21332 ,
         \21333 , \21334 , \21335 , \21336 , \21337 , \21338 , \21339 , \21340 , \21341 , \21342 ,
         \21343 , \21344 , \21345 , \21346 , \21347 , \21348 , \21349 , \21350 , \21351 , \21352 ,
         \21353 , \21354 , \21355 , \21356 , \21357 , \21358 , \21359 , \21360 , \21361 , \21362 ,
         \21363 , \21364 , \21365 , \21366 , \21367 , \21368 , \21369 , \21370 , \21371 , \21372 ,
         \21373 , \21374 , \21375 , \21376 , \21377 , \21378 , \21379 , \21380 , \21381 , \21382 ,
         \21383 , \21384 , \21385 , \21386 , \21387 , \21388 , \21389 , \21390 , \21391 , \21392 ,
         \21393 , \21394 , \21395 , \21396 , \21397 , \21398 , \21399 , \21400 , \21401 , \21402 ,
         \21403 , \21404 , \21405 , \21406 , \21407 , \21408 , \21409 , \21410 , \21411 , \21412 ,
         \21413 , \21414 , \21415 , \21416 , \21417 , \21418 , \21419 , \21420 , \21421 , \21422 ,
         \21423 , \21424 , \21425 , \21426 , \21427 , \21428 , \21429 , \21430 , \21431 , \21432 ,
         \21433 , \21434 , \21435 , \21436 , \21437 , \21438 , \21439 , \21440 , \21441 , \21442 ,
         \21443 , \21444 , \21445 , \21446 , \21447 , \21448 , \21449 , \21450 , \21451 , \21452 ,
         \21453 , \21454 , \21455 , \21456 , \21457 , \21458 , \21459 , \21460 , \21461 , \21462 ,
         \21463 , \21464 , \21465 , \21466 , \21467 , \21468 , \21469 , \21470 , \21471 , \21472 ,
         \21473 , \21474 , \21475 , \21476 , \21477 , \21478 , \21479 , \21480 , \21481 , \21482 ,
         \21483 , \21484 , \21485 , \21486 , \21487 , \21488 , \21489 , \21490 , \21491 , \21492 ,
         \21493 , \21494 , \21495 , \21496 , \21497 , \21498 , \21499 , \21500 , \21501 , \21502 ,
         \21503 , \21504 , \21505 , \21506 , \21507 , \21508 , \21509 , \21510 , \21511 , \21512 ,
         \21513 , \21514 , \21515 , \21516 , \21517 , \21518 , \21519 , \21520 , \21521 , \21522 ,
         \21523 , \21524 , \21525 , \21526 , \21527 , \21528 , \21529 , \21530 , \21531 , \21532 ,
         \21533 , \21534 , \21535 , \21536 , \21537 , \21538 , \21539 , \21540 , \21541 , \21542 ,
         \21543 , \21544 , \21545 , \21546 , \21547 , \21548 , \21549 , \21550 , \21551 , \21552 ,
         \21553 , \21554 , \21555 , \21556 , \21557 , \21558 , \21559 , \21560 , \21561 , \21562 ,
         \21563 , \21564 , \21565 , \21566 , \21567 , \21568 , \21569 , \21570 , \21571 , \21572 ,
         \21573 , \21574 , \21575 , \21576 , \21577 , \21578 , \21579 , \21580 , \21581 , \21582 ,
         \21583 , \21584 , \21585 , \21586 , \21587 , \21588 , \21589 , \21590 , \21591 , \21592 ,
         \21593 , \21594 , \21595 , \21596 , \21597 , \21598 , \21599 , \21600 , \21601 , \21602 ,
         \21603 , \21604 , \21605 , \21606 , \21607 , \21608 , \21609 , \21610 , \21611 , \21612 ,
         \21613 , \21614 , \21615 , \21616 , \21617 , \21618 , \21619 , \21620 , \21621 , \21622 ,
         \21623 , \21624 , \21625 , \21626 , \21627 , \21628 , \21629 , \21630 , \21631 , \21632 ,
         \21633 , \21634 , \21635 , \21636 , \21637 , \21638 , \21639 , \21640 , \21641 , \21642 ,
         \21643 , \21644 , \21645 , \21646 , \21647 , \21648 , \21649 , \21650 , \21651 , \21652 ,
         \21653 , \21654 , \21655 , \21656 , \21657 , \21658 , \21659 , \21660 , \21661 , \21662 ,
         \21663 , \21664 , \21665 , \21666 , \21667 , \21668 , \21669 , \21670 , \21671 , \21672 ,
         \21673 , \21674 , \21675 , \21676 , \21677 , \21678 , \21679 , \21680 , \21681 , \21682 ,
         \21683 , \21684 , \21685 , \21686 , \21687 , \21688 , \21689 , \21690 , \21691 , \21692 ,
         \21693 , \21694 , \21695 , \21696 , \21697 , \21698 , \21699 , \21700 , \21701 , \21702 ,
         \21703 , \21704 , \21705 , \21706 , \21707 , \21708 , \21709 , \21710 , \21711 , \21712 ,
         \21713 , \21714 , \21715 , \21716 , \21717 , \21718 , \21719 , \21720 , \21721 , \21722 ,
         \21723 , \21724 , \21725 , \21726 , \21727 , \21728 , \21729 , \21730 , \21731 , \21732 ,
         \21733 , \21734 , \21735 , \21736 , \21737 , \21738 , \21739 , \21740 , \21741 , \21742 ,
         \21743 , \21744 , \21745 , \21746 , \21747 , \21748 , \21749 , \21750 , \21751 , \21752 ,
         \21753 , \21754 , \21755 , \21756 , \21757 , \21758 , \21759 , \21760 , \21761 , \21762 ,
         \21763 , \21764 , \21765 , \21766 , \21767 , \21768 , \21769 , \21770 , \21771 , \21772 ,
         \21773 , \21774 , \21775 , \21776 , \21777 , \21778 , \21779 , \21780 , \21781 , \21782 ,
         \21783 , \21784 , \21785 , \21786 , \21787 , \21788 , \21789 , \21790 , \21791 , \21792 ,
         \21793 , \21794 , \21795 , \21796 , \21797 , \21798 , \21799 , \21800 , \21801 , \21802 ,
         \21803 , \21804 , \21805 , \21806 , \21807 , \21808 , \21809 , \21810 , \21811 , \21812 ,
         \21813 , \21814 , \21815 , \21816 , \21817 , \21818 , \21819 , \21820 , \21821 , \21822 ,
         \21823 , \21824 , \21825 , \21826 , \21827 , \21828 , \21829 , \21830 , \21831 , \21832 ,
         \21833 , \21834 , \21835 , \21836 , \21837 , \21838 , \21839 , \21840 , \21841 , \21842 ,
         \21843 , \21844 , \21845 , \21846 , \21847 , \21848 , \21849 , \21850 , \21851 , \21852 ,
         \21853 , \21854 , \21855 , \21856 , \21857 , \21858 , \21859 , \21860 , \21861 , \21862 ,
         \21863 , \21864 , \21865 , \21866 , \21867 , \21868 , \21869 , \21870 , \21871 , \21872 ,
         \21873 , \21874 , \21875 , \21876 , \21877 , \21878 , \21879 , \21880 , \21881 , \21882 ,
         \21883 , \21884 , \21885 , \21886 , \21887 , \21888 , \21889 , \21890 , \21891 , \21892 ,
         \21893 , \21894 , \21895 , \21896 , \21897 , \21898 , \21899 , \21900 , \21901 , \21902 ,
         \21903 , \21904 , \21905 , \21906 , \21907 , \21908 , \21909 , \21910 , \21911 , \21912 ,
         \21913 , \21914 , \21915 , \21916 , \21917 , \21918 , \21919 , \21920 , \21921 , \21922 ,
         \21923 , \21924 , \21925 , \21926 , \21927 , \21928 , \21929 , \21930 , \21931 , \21932 ,
         \21933 , \21934 , \21935 , \21936 , \21937 , \21938 , \21939 , \21940 , \21941 , \21942 ,
         \21943 , \21944 , \21945 , \21946 , \21947 , \21948 , \21949 , \21950 , \21951 , \21952 ,
         \21953 , \21954 , \21955 , \21956 , \21957 , \21958 , \21959 , \21960 , \21961 , \21962 ,
         \21963 , \21964 , \21965 , \21966 , \21967 , \21968 , \21969 , \21970 , \21971 , \21972 ,
         \21973 , \21974 , \21975 , \21976 , \21977 , \21978 , \21979 , \21980 , \21981 , \21982 ,
         \21983 , \21984 , \21985 , \21986 , \21987 , \21988 , \21989 , \21990 , \21991 , \21992 ,
         \21993 , \21994 , \21995 , \21996 , \21997 , \21998 , \21999 , \22000 , \22001 , \22002 ,
         \22003 , \22004 , \22005 , \22006 , \22007 , \22008 , \22009 , \22010 , \22011 , \22012 ,
         \22013 , \22014 , \22015 , \22016 , \22017 , \22018 , \22019 , \22020 , \22021 , \22022 ,
         \22023 , \22024 , \22025 , \22026 , \22027 , \22028 , \22029 , \22030 , \22031 , \22032 ,
         \22033 , \22034 , \22035 , \22036 , \22037 , \22038 , \22039 , \22040 , \22041 , \22042 ,
         \22043 , \22044 , \22045 , \22046 , \22047 , \22048 , \22049 , \22050 , \22051 , \22052 ,
         \22053 , \22054 , \22055 , \22056 , \22057 , \22058 , \22059 , \22060 , \22061 , \22062 ,
         \22063 , \22064 , \22065 , \22066 , \22067 , \22068 , \22069 , \22070 , \22071 , \22072 ,
         \22073 , \22074 , \22075 , \22076 , \22077 , \22078 , \22079 , \22080 , \22081 , \22082 ,
         \22083 , \22084 , \22085 , \22086 , \22087 , \22088 , \22089 , \22090 , \22091 , \22092 ,
         \22093 , \22094 , \22095 , \22096 , \22097 , \22098 , \22099 , \22100 , \22101 , \22102 ,
         \22103 , \22104 , \22105 , \22106 , \22107 , \22108 , \22109 , \22110 , \22111 , \22112 ,
         \22113 , \22114 , \22115 , \22116 , \22117 , \22118 , \22119 , \22120 , \22121 , \22122 ,
         \22123 , \22124 , \22125 , \22126 , \22127 , \22128 , \22129 , \22130 , \22131 , \22132 ,
         \22133 , \22134 , \22135 , \22136 , \22137 , \22138 , \22139 , \22140 , \22141 , \22142 ,
         \22143 , \22144 , \22145 , \22146 , \22147 , \22148 , \22149 , \22150 , \22151 , \22152 ,
         \22153 , \22154 , \22155 , \22156 , \22157 , \22158 , \22159 , \22160 , \22161 , \22162 ,
         \22163 , \22164 , \22165 , \22166 , \22167 , \22168 , \22169 , \22170 , \22171 , \22172 ,
         \22173 , \22174 , \22175 , \22176 , \22177 , \22178 , \22179 , \22180 , \22181 , \22182 ,
         \22183 , \22184 , \22185 , \22186 , \22187 , \22188 , \22189 , \22190 , \22191 , \22192 ,
         \22193 , \22194 , \22195 , \22196 , \22197 , \22198 , \22199 , \22200 , \22201 , \22202 ,
         \22203 , \22204 , \22205 , \22206 , \22207 , \22208 , \22209 , \22210 , \22211 , \22212 ,
         \22213 , \22214 , \22215 , \22216 , \22217 , \22218 , \22219 , \22220 , \22221 , \22222 ,
         \22223 , \22224 , \22225 , \22226 , \22227 , \22228 , \22229 , \22230 , \22231 , \22232 ,
         \22233 , \22234 , \22235 , \22236 , \22237 , \22238 , \22239 , \22240 , \22241 , \22242 ,
         \22243 , \22244 , \22245 , \22246 , \22247 , \22248 , \22249 , \22250 , \22251 , \22252 ,
         \22253 , \22254 , \22255 , \22256 , \22257 , \22258 , \22259 , \22260 , \22261 , \22262 ,
         \22263 , \22264 , \22265 , \22266 , \22267 , \22268 , \22269 , \22270 , \22271 , \22272 ,
         \22273 , \22274 , \22275 , \22276 , \22277 , \22278 , \22279 , \22280 , \22281 , \22282 ,
         \22283 , \22284 , \22285 , \22286 , \22287 , \22288 , \22289 , \22290 , \22291 , \22292 ,
         \22293 , \22294 , \22295 , \22296 , \22297 , \22298 , \22299 , \22300 , \22301 , \22302 ,
         \22303 , \22304 , \22305 , \22306 , \22307 , \22308 , \22309 , \22310 , \22311 , \22312 ,
         \22313 , \22314 , \22315 , \22316 , \22317 , \22318 , \22319 , \22320 , \22321 , \22322 ,
         \22323 , \22324 , \22325 , \22326 , \22327 , \22328 , \22329 , \22330 , \22331 , \22332 ,
         \22333 , \22334 , \22335 , \22336 , \22337 , \22338 , \22339 , \22340 , \22341 , \22342 ,
         \22343 , \22344 , \22345 , \22346 , \22347 , \22348 , \22349 , \22350 , \22351 , \22352 ,
         \22353 , \22354 , \22355 , \22356 , \22357 , \22358 , \22359 , \22360 , \22361 , \22362 ,
         \22363 , \22364 , \22365 , \22366 , \22367 , \22368 , \22369 , \22370 , \22371 , \22372 ,
         \22373 , \22374 , \22375 , \22376 , \22377 , \22378 , \22379 , \22380 , \22381 , \22382 ,
         \22383 , \22384 , \22385 , \22386 , \22387 , \22388 , \22389 , \22390 , \22391 , \22392 ,
         \22393 , \22394 , \22395 , \22396 , \22397 , \22398 , \22399 , \22400 , \22401 , \22402 ,
         \22403 , \22404 , \22405 , \22406 , \22407 , \22408 , \22409 , \22410 , \22411 , \22412 ,
         \22413 , \22414 , \22415 , \22416 , \22417 , \22418 , \22419 , \22420 , \22421 , \22422 ,
         \22423 , \22424 , \22425 , \22426 , \22427 , \22428 , \22429 , \22430 , \22431 , \22432 ,
         \22433 , \22434 , \22435 , \22436 , \22437 , \22438 , \22439 , \22440 , \22441 , \22442 ,
         \22443 , \22444 , \22445 , \22446 , \22447 , \22448 , \22449 , \22450 , \22451 , \22452 ,
         \22453 , \22454 , \22455 , \22456 , \22457 , \22458 , \22459 , \22460 , \22461 , \22462 ,
         \22463 , \22464 , \22465 , \22466 , \22467 , \22468 , \22469 , \22470 , \22471 , \22472 ,
         \22473 , \22474 , \22475 , \22476 , \22477 , \22478 , \22479 , \22480 , \22481 , \22482 ,
         \22483 , \22484 , \22485 , \22486 , \22487 , \22488 , \22489 , \22490 , \22491 , \22492 ,
         \22493 , \22494 , \22495 , \22496 , \22497 , \22498 , \22499 , \22500 , \22501 , \22502 ,
         \22503 , \22504 , \22505 , \22506 , \22507 , \22508 , \22509 , \22510 , \22511 , \22512 ,
         \22513 , \22514 , \22515 , \22516 , \22517 , \22518 , \22519 , \22520 , \22521 , \22522 ,
         \22523 , \22524 , \22525 , \22526 , \22527 , \22528 , \22529 , \22530 , \22531 , \22532 ,
         \22533 , \22534 , \22535 , \22536 , \22537 , \22538 , \22539 , \22540 , \22541 , \22542 ,
         \22543 , \22544 , \22545 , \22546 , \22547 , \22548 , \22549 , \22550 , \22551 , \22552 ,
         \22553 , \22554 , \22555 , \22556 , \22557 , \22558 , \22559 , \22560 , \22561 , \22562 ,
         \22563 , \22564 , \22565 , \22566 , \22567 , \22568 , \22569 , \22570 , \22571 , \22572 ,
         \22573 , \22574 , \22575 , \22576 , \22577 , \22578 , \22579 , \22580 , \22581 , \22582 ,
         \22583 , \22584 , \22585 , \22586 , \22587 , \22588 , \22589 , \22590 , \22591 , \22592 ,
         \22593 , \22594 , \22595 , \22596 , \22597 , \22598 , \22599 , \22600 , \22601 , \22602 ,
         \22603 , \22604 , \22605 , \22606 , \22607 , \22608 , \22609 , \22610 , \22611 , \22612 ,
         \22613 , \22614 , \22615 , \22616 , \22617 , \22618 , \22619 , \22620 , \22621 , \22622 ,
         \22623 , \22624 , \22625 , \22626 , \22627 , \22628 , \22629 , \22630 , \22631 , \22632 ,
         \22633 , \22634 , \22635 , \22636 , \22637 , \22638 , \22639 , \22640 , \22641 , \22642 ,
         \22643 , \22644 , \22645 , \22646 , \22647 , \22648 , \22649 , \22650 , \22651 , \22652 ,
         \22653 , \22654 , \22655 , \22656 , \22657 , \22658 , \22659 , \22660 , \22661 , \22662 ,
         \22663 , \22664 , \22665 , \22666 , \22667 , \22668 , \22669 , \22670 , \22671 , \22672 ,
         \22673 , \22674 , \22675 , \22676 , \22677 , \22678 , \22679 , \22680 , \22681 , \22682 ,
         \22683 , \22684 , \22685 , \22686 , \22687 , \22688 , \22689 , \22690 , \22691 , \22692 ,
         \22693 , \22694 , \22695 , \22696 , \22697 , \22698 , \22699 , \22700 , \22701 , \22702 ,
         \22703 , \22704 , \22705 , \22706 , \22707 , \22708 , \22709 , \22710 , \22711 , \22712 ,
         \22713 , \22714 , \22715 , \22716 , \22717 , \22718 , \22719 , \22720 , \22721 , \22722 ,
         \22723 , \22724 , \22725 , \22726 , \22727 , \22728 , \22729 , \22730 , \22731 , \22732 ,
         \22733 , \22734 , \22735 , \22736 , \22737 , \22738 , \22739 , \22740 , \22741 , \22742 ,
         \22743 , \22744 , \22745 , \22746 , \22747 , \22748 , \22749 , \22750 , \22751 , \22752 ,
         \22753 , \22754 , \22755 , \22756 , \22757 , \22758 , \22759 , \22760 , \22761 , \22762 ,
         \22763 , \22764 , \22765 , \22766 , \22767 , \22768 , \22769 , \22770 , \22771 , \22772 ,
         \22773 , \22774 , \22775 , \22776 , \22777 , \22778 , \22779 , \22780 , \22781 , \22782 ,
         \22783 , \22784 , \22785 , \22786 , \22787 , \22788 , \22789 , \22790 , \22791 , \22792 ,
         \22793 , \22794 , \22795 , \22796 , \22797 , \22798 , \22799 , \22800 , \22801 , \22802 ,
         \22803 , \22804 , \22805 , \22806 , \22807 , \22808 , \22809 , \22810 , \22811 , \22812 ,
         \22813 , \22814 , \22815 , \22816 , \22817 , \22818 , \22819 , \22820 , \22821 , \22822 ,
         \22823 , \22824 , \22825 , \22826 , \22827 , \22828 , \22829 , \22830 , \22831 , \22832 ,
         \22833 , \22834 , \22835 , \22836 , \22837 , \22838 , \22839 , \22840 , \22841 , \22842 ,
         \22843 , \22844 , \22845 , \22846 , \22847 , \22848 , \22849 , \22850 , \22851 , \22852 ,
         \22853 , \22854 , \22855 , \22856 , \22857 , \22858 , \22859 , \22860 , \22861 , \22862 ,
         \22863 , \22864 , \22865 , \22866 , \22867 , \22868 , \22869 , \22870 , \22871 , \22872 ,
         \22873 , \22874 , \22875 , \22876 , \22877 , \22878 , \22879 , \22880 , \22881 , \22882 ,
         \22883 , \22884 , \22885 , \22886 , \22887 , \22888 , \22889 , \22890 , \22891 , \22892 ,
         \22893 , \22894 , \22895 , \22896 , \22897 , \22898 , \22899 , \22900 , \22901 , \22902 ,
         \22903 , \22904 , \22905 , \22906 , \22907 , \22908 , \22909 , \22910 , \22911 , \22912 ,
         \22913 , \22914 , \22915 , \22916 , \22917 , \22918 , \22919 , \22920 , \22921 , \22922 ,
         \22923 , \22924 , \22925 , \22926 , \22927 , \22928 , \22929 , \22930 , \22931 , \22932 ,
         \22933 , \22934 , \22935 , \22936 , \22937 , \22938 , \22939 , \22940 , \22941 , \22942 ,
         \22943 , \22944 , \22945 , \22946 , \22947 , \22948 , \22949 , \22950 , \22951 , \22952 ,
         \22953 , \22954 , \22955 , \22956 , \22957 , \22958 , \22959 , \22960 , \22961 , \22962 ,
         \22963 , \22964 , \22965 , \22966 , \22967 , \22968 , \22969 , \22970 , \22971 , \22972 ,
         \22973 , \22974 , \22975 , \22976 , \22977 , \22978 , \22979 , \22980 , \22981 , \22982 ,
         \22983 , \22984 , \22985 , \22986 , \22987 , \22988 , \22989 , \22990 , \22991 , \22992 ,
         \22993 , \22994 , \22995 , \22996 , \22997 , \22998 , \22999 , \23000 , \23001 , \23002 ,
         \23003 , \23004 , \23005 , \23006 , \23007 , \23008 , \23009 , \23010 , \23011 , \23012 ,
         \23013 , \23014 , \23015 , \23016 , \23017 , \23018 , \23019 , \23020 , \23021 , \23022 ,
         \23023 , \23024 , \23025 , \23026 , \23027 , \23028 , \23029 , \23030 , \23031 , \23032 ,
         \23033 , \23034 , \23035 , \23036 , \23037 , \23038 , \23039 , \23040 , \23041 , \23042 ,
         \23043 , \23044 , \23045 , \23046 , \23047 , \23048 , \23049 , \23050 , \23051 , \23052 ,
         \23053 , \23054 , \23055 , \23056 , \23057 , \23058 , \23059 , \23060 , \23061 , \23062 ,
         \23063 , \23064 , \23065 , \23066 , \23067 , \23068 , \23069 , \23070 , \23071 , \23072 ,
         \23073 , \23074 , \23075 , \23076 , \23077 , \23078 , \23079 , \23080 , \23081 , \23082 ,
         \23083 , \23084 , \23085 , \23086 , \23087 , \23088 , \23089 , \23090 , \23091 , \23092 ,
         \23093 , \23094 , \23095 , \23096 , \23097 , \23098 , \23099 , \23100 , \23101 , \23102 ,
         \23103 , \23104 , \23105 , \23106 , \23107 , \23108 , \23109 , \23110 , \23111 , \23112 ,
         \23113 , \23114 , \23115 , \23116 , \23117 , \23118 , \23119 , \23120 , \23121 , \23122 ,
         \23123 , \23124 , \23125 , \23126 , \23127 , \23128 , \23129 , \23130 , \23131 , \23132 ,
         \23133 , \23134 , \23135 , \23136 , \23137 , \23138 , \23139 , \23140 , \23141 , \23142 ,
         \23143 , \23144 , \23145 , \23146 , \23147 , \23148 , \23149 , \23150 , \23151 , \23152 ,
         \23153 , \23154 , \23155 , \23156 , \23157 , \23158 , \23159 , \23160 , \23161 , \23162 ,
         \23163 , \23164 , \23165 , \23166 , \23167 , \23168 , \23169 , \23170 , \23171 , \23172 ,
         \23173 , \23174 , \23175 , \23176 , \23177 , \23178 , \23179 , \23180 , \23181 , \23182 ,
         \23183 , \23184 , \23185 , \23186 , \23187 , \23188 , \23189 , \23190 , \23191 , \23192 ,
         \23193 , \23194 , \23195 , \23196 , \23197 , \23198 , \23199 , \23200 , \23201 , \23202 ,
         \23203 , \23204 , \23205 , \23206 , \23207 , \23208 , \23209 , \23210 , \23211 , \23212 ,
         \23213 , \23214 , \23215 , \23216 , \23217 , \23218 , \23219 , \23220 , \23221 , \23222 ,
         \23223 , \23224 , \23225 , \23226 , \23227 , \23228 , \23229 , \23230 , \23231 , \23232 ,
         \23233 , \23234 , \23235 , \23236 , \23237 , \23238 , \23239 , \23240 , \23241 , \23242 ,
         \23243 , \23244 , \23245 , \23246 , \23247 , \23248 , \23249 , \23250 , \23251 , \23252 ,
         \23253 , \23254 , \23255 , \23256 , \23257 , \23258 , \23259 , \23260 , \23261 , \23262 ,
         \23263 , \23264 , \23265 , \23266 , \23267 , \23268 , \23269 , \23270 , \23271 , \23272 ,
         \23273 , \23274 , \23275 , \23276 , \23277 , \23278 , \23279 , \23280 , \23281 , \23282 ,
         \23283 , \23284 , \23285 , \23286 , \23287 , \23288 , \23289 , \23290 , \23291 , \23292 ,
         \23293 , \23294 , \23295 , \23296 , \23297 , \23298 , \23299 , \23300 , \23301 , \23302 ,
         \23303 , \23304 , \23305 , \23306 , \23307 , \23308 , \23309 , \23310 , \23311 , \23312 ,
         \23313 , \23314 , \23315 , \23316 , \23317 , \23318 , \23319 , \23320 , \23321 , \23322 ,
         \23323 , \23324 , \23325 , \23326 , \23327 , \23328 , \23329 , \23330 , \23331 , \23332 ,
         \23333 , \23334 , \23335 , \23336 , \23337 , \23338 , \23339 , \23340 , \23341 , \23342 ,
         \23343 , \23344 , \23345 , \23346 , \23347 , \23348 , \23349 , \23350 , \23351 , \23352 ,
         \23353 , \23354 , \23355 , \23356 , \23357 , \23358 , \23359 , \23360 , \23361 , \23362 ,
         \23363 , \23364 , \23365 , \23366 , \23367 , \23368 , \23369 , \23370 , \23371 , \23372 ,
         \23373 , \23374 , \23375 , \23376 , \23377 , \23378 , \23379 , \23380 , \23381 , \23382 ,
         \23383 , \23384 , \23385 , \23386 , \23387 , \23388 , \23389 , \23390 , \23391 , \23392 ,
         \23393 , \23394 , \23395 , \23396 , \23397 , \23398 , \23399 , \23400 , \23401 , \23402 ,
         \23403 , \23404 , \23405 , \23406 , \23407 , \23408 , \23409 , \23410 , \23411 , \23412 ,
         \23413 , \23414 , \23415 , \23416 , \23417 , \23418 , \23419 , \23420 , \23421 , \23422 ,
         \23423 , \23424 , \23425 , \23426 , \23427 , \23428 , \23429 , \23430 , \23431 , \23432 ,
         \23433 , \23434 , \23435 , \23436 , \23437 , \23438 , \23439 , \23440 , \23441 , \23442 ,
         \23443 , \23444 , \23445 , \23446 , \23447 , \23448 , \23449 , \23450 , \23451 , \23452 ,
         \23453 , \23454 , \23455 , \23456 , \23457 , \23458 , \23459 , \23460 , \23461 , \23462 ,
         \23463 , \23464 , \23465 , \23466 , \23467 , \23468 , \23469 , \23470 , \23471 , \23472 ,
         \23473 , \23474 , \23475 , \23476 , \23477 , \23478 , \23479 , \23480 , \23481 , \23482 ,
         \23483 , \23484 , \23485 , \23486 , \23487 , \23488 , \23489 , \23490 , \23491 , \23492 ,
         \23493 , \23494 , \23495 , \23496 , \23497 , \23498 , \23499 , \23500 , \23501 , \23502 ,
         \23503 , \23504 , \23505 , \23506 , \23507 , \23508 , \23509 , \23510 , \23511 , \23512 ,
         \23513 , \23514 , \23515 , \23516 , \23517 , \23518 , \23519 , \23520 , \23521 , \23522 ,
         \23523 , \23524 , \23525 , \23526 , \23527 , \23528 , \23529 , \23530 , \23531 , \23532 ,
         \23533 , \23534 , \23535 , \23536 , \23537 , \23538 , \23539 , \23540 , \23541 , \23542 ,
         \23543 , \23544 , \23545 , \23546 , \23547 , \23548 , \23549 , \23550 , \23551 , \23552 ,
         \23553 , \23554 , \23555 , \23556 , \23557 , \23558 , \23559 , \23560 , \23561 , \23562 ,
         \23563 , \23564 , \23565 , \23566 , \23567 , \23568 , \23569 , \23570 , \23571 , \23572 ,
         \23573 , \23574 , \23575 , \23576 , \23577 , \23578 , \23579 , \23580 , \23581 , \23582 ,
         \23583 , \23584 , \23585 , \23586 , \23587 , \23588 , \23589 , \23590 , \23591 , \23592 ,
         \23593 , \23594 , \23595 , \23596 , \23597 , \23598 , \23599 , \23600 , \23601 , \23602 ,
         \23603 , \23604 , \23605 , \23606 , \23607 , \23608 , \23609 , \23610 , \23611 , \23612 ,
         \23613 , \23614 , \23615 , \23616 , \23617 , \23618 , \23619 , \23620 , \23621 , \23622 ,
         \23623 , \23624 , \23625 , \23626 , \23627 , \23628 , \23629 , \23630 , \23631 , \23632 ,
         \23633 , \23634 , \23635 , \23636 , \23637 , \23638 , \23639 , \23640 , \23641 , \23642 ,
         \23643 , \23644 , \23645 , \23646 , \23647 , \23648 , \23649 , \23650 , \23651 , \23652 ,
         \23653 , \23654 , \23655 , \23656 , \23657 , \23658 , \23659 , \23660 , \23661 , \23662 ,
         \23663 , \23664 , \23665 , \23666 , \23667 , \23668 , \23669 , \23670 , \23671 , \23672 ,
         \23673 , \23674 , \23675 , \23676 , \23677 , \23678 , \23679 , \23680 , \23681 , \23682 ,
         \23683 , \23684 , \23685 , \23686 , \23687 , \23688 , \23689 , \23690 , \23691 , \23692 ,
         \23693 , \23694 , \23695 , \23696 , \23697 , \23698 , \23699 , \23700 , \23701 , \23702 ,
         \23703 , \23704 , \23705 , \23706 , \23707 , \23708 , \23709 , \23710 , \23711 , \23712 ,
         \23713 , \23714 , \23715 , \23716 , \23717 , \23718 , \23719 , \23720 , \23721 , \23722 ,
         \23723 , \23724 , \23725 , \23726 , \23727 , \23728 , \23729 , \23730 , \23731 , \23732 ,
         \23733 , \23734 , \23735 , \23736 , \23737 , \23738 , \23739 , \23740 , \23741 , \23742 ,
         \23743 , \23744 , \23745 , \23746 , \23747 , \23748 , \23749 , \23750 , \23751 , \23752 ,
         \23753 , \23754 , \23755 , \23756 , \23757 , \23758 , \23759 , \23760 , \23761 , \23762 ,
         \23763 , \23764 , \23765 , \23766 , \23767 , \23768 , \23769 , \23770 , \23771 , \23772 ,
         \23773 , \23774 , \23775 , \23776 , \23777 , \23778 , \23779 , \23780 , \23781 , \23782 ,
         \23783 , \23784 , \23785 , \23786 , \23787 , \23788 , \23789 , \23790 , \23791 , \23792 ,
         \23793 , \23794 , \23795 , \23796 , \23797 , \23798 , \23799 , \23800 , \23801 , \23802 ,
         \23803 , \23804 , \23805 , \23806 , \23807 , \23808 , \23809 , \23810 , \23811 , \23812 ,
         \23813 , \23814 , \23815 , \23816 , \23817 , \23818 , \23819 , \23820 , \23821 , \23822 ,
         \23823 , \23824 , \23825 , \23826 , \23827 , \23828 , \23829 , \23830 , \23831 , \23832 ,
         \23833 , \23834 , \23835 , \23836 , \23837 , \23838 , \23839 , \23840 , \23841 , \23842 ,
         \23843 , \23844 , \23845 , \23846 , \23847 , \23848 , \23849 , \23850 , \23851 , \23852 ,
         \23853 , \23854 , \23855 , \23856 , \23857 , \23858 , \23859 , \23860 , \23861 , \23862 ,
         \23863 , \23864 , \23865 , \23866 , \23867 , \23868 , \23869 , \23870 , \23871 , \23872 ,
         \23873 , \23874 , \23875 , \23876 , \23877 , \23878 , \23879 , \23880 , \23881 , \23882 ,
         \23883 , \23884 , \23885 , \23886 , \23887 , \23888 , \23889 , \23890 , \23891 , \23892 ,
         \23893 , \23894 , \23895 , \23896 , \23897 , \23898 , \23899 , \23900 , \23901 , \23902 ,
         \23903 , \23904 , \23905 , \23906 , \23907 , \23908 , \23909 , \23910 , \23911 , \23912 ,
         \23913 , \23914 , \23915 , \23916 , \23917 , \23918 , \23919 , \23920 , \23921 , \23922 ,
         \23923 , \23924 , \23925 , \23926 , \23927 , \23928 , \23929 , \23930 , \23931 , \23932 ,
         \23933 , \23934 , \23935 , \23936 , \23937 , \23938 , \23939 , \23940 , \23941 , \23942 ,
         \23943 , \23944 , \23945 , \23946 , \23947 , \23948 , \23949 , \23950 , \23951 , \23952 ,
         \23953 , \23954 , \23955 , \23956 , \23957 , \23958 , \23959 , \23960 , \23961 , \23962 ,
         \23963 , \23964 , \23965 , \23966 , \23967 , \23968 , \23969 , \23970 , \23971 , \23972 ,
         \23973 , \23974 , \23975 , \23976 , \23977 , \23978 , \23979 , \23980 , \23981 , \23982 ,
         \23983 , \23984 , \23985 , \23986 , \23987 , \23988 , \23989 , \23990 , \23991 , \23992 ,
         \23993 , \23994 , \23995 , \23996 , \23997 , \23998 , \23999 , \24000 , \24001 , \24002 ,
         \24003 , \24004 , \24005 , \24006 , \24007 , \24008 , \24009 , \24010 , \24011 , \24012 ,
         \24013 , \24014 , \24015 , \24016 , \24017 , \24018 , \24019 , \24020 , \24021 , \24022 ,
         \24023 , \24024 , \24025 , \24026 , \24027 , \24028 , \24029 , \24030 , \24031 , \24032 ,
         \24033 , \24034 , \24035 , \24036 , \24037 , \24038 , \24039 , \24040 , \24041 , \24042 ,
         \24043 , \24044 , \24045 , \24046 , \24047 , \24048 , \24049 , \24050 , \24051 , \24052 ,
         \24053 , \24054 , \24055 , \24056 , \24057 , \24058 , \24059 , \24060 , \24061 , \24062 ,
         \24063 , \24064 , \24065 , \24066 , \24067 , \24068 , \24069 , \24070 , \24071 , \24072 ,
         \24073 , \24074 , \24075 , \24076 , \24077 , \24078 , \24079 , \24080 , \24081 , \24082 ,
         \24083 , \24084 , \24085 , \24086 , \24087 , \24088 , \24089 , \24090 , \24091 , \24092 ,
         \24093 , \24094 , \24095 , \24096 , \24097 , \24098 , \24099 , \24100 , \24101 , \24102 ,
         \24103 , \24104 , \24105 , \24106 , \24107 , \24108 , \24109 , \24110 , \24111 , \24112 ,
         \24113 , \24114 , \24115 , \24116 , \24117 , \24118 , \24119 , \24120 , \24121 , \24122 ,
         \24123 , \24124 , \24125 , \24126 , \24127 , \24128 , \24129 , \24130 , \24131 , \24132 ,
         \24133 , \24134 , \24135 , \24136 , \24137 , \24138 , \24139 , \24140 , \24141 , \24142 ,
         \24143 , \24144 , \24145 , \24146 , \24147 , \24148 , \24149 , \24150 , \24151 , \24152 ,
         \24153 , \24154 , \24155 , \24156 , \24157 , \24158 , \24159 , \24160 , \24161 , \24162 ,
         \24163 , \24164 , \24165 , \24166 , \24167 , \24168 , \24169 , \24170 , \24171 , \24172 ,
         \24173 , \24174 , \24175 , \24176 , \24177 , \24178 , \24179 , \24180 , \24181 , \24182 ,
         \24183 , \24184 , \24185 , \24186 , \24187 , \24188 , \24189 , \24190 , \24191 , \24192 ,
         \24193 , \24194 , \24195 , \24196 , \24197 , \24198 , \24199 , \24200 , \24201 , \24202 ,
         \24203 , \24204 , \24205 , \24206 , \24207 , \24208 , \24209 , \24210 , \24211 , \24212 ,
         \24213 , \24214 , \24215 , \24216 , \24217 , \24218 , \24219 , \24220 , \24221 , \24222 ,
         \24223 , \24224 , \24225 , \24226 , \24227 , \24228 , \24229 , \24230 , \24231 , \24232 ,
         \24233 , \24234 , \24235 , \24236 , \24237 , \24238 , \24239 , \24240 , \24241 , \24242 ,
         \24243 , \24244 , \24245 , \24246 , \24247 , \24248 , \24249 , \24250 , \24251 , \24252 ,
         \24253 , \24254 , \24255 , \24256 , \24257 , \24258 , \24259 , \24260 , \24261 , \24262 ,
         \24263 , \24264 , \24265 , \24266 , \24267 , \24268 , \24269 , \24270 , \24271 , \24272 ,
         \24273 , \24274 , \24275 , \24276 , \24277 , \24278 , \24279 , \24280 , \24281 , \24282 ,
         \24283 , \24284 , \24285 , \24286 , \24287 , \24288 , \24289 , \24290 , \24291 , \24292 ,
         \24293 , \24294 , \24295 , \24296 , \24297 , \24298 , \24299 , \24300 , \24301 , \24302 ,
         \24303 , \24304 , \24305 , \24306 , \24307 , \24308 , \24309 , \24310 , \24311 , \24312 ,
         \24313 , \24314 , \24315 , \24316 , \24317 , \24318 , \24319 , \24320 , \24321 , \24322 ,
         \24323 , \24324 , \24325 , \24326 , \24327 , \24328 , \24329 , \24330 , \24331 , \24332 ,
         \24333 , \24334 , \24335 , \24336 , \24337 , \24338 , \24339 , \24340 , \24341 , \24342 ,
         \24343 , \24344 , \24345 , \24346 , \24347 , \24348 , \24349 , \24350 , \24351 , \24352 ,
         \24353 , \24354 , \24355 , \24356 , \24357 , \24358 , \24359 , \24360 , \24361 , \24362 ,
         \24363 , \24364 , \24365 , \24366 , \24367 , \24368 , \24369 , \24370 , \24371 , \24372 ,
         \24373 , \24374 , \24375 , \24376 , \24377 , \24378 , \24379 , \24380 , \24381 , \24382 ,
         \24383 , \24384 , \24385 , \24386 , \24387 , \24388 , \24389 , \24390 , \24391 , \24392 ,
         \24393 , \24394 , \24395 , \24396 , \24397 , \24398 , \24399 , \24400 , \24401 , \24402 ,
         \24403 , \24404 , \24405 , \24406 , \24407 , \24408 , \24409 , \24410 , \24411 , \24412 ,
         \24413 , \24414 , \24415 , \24416 , \24417 , \24418 , \24419 , \24420 , \24421 , \24422 ,
         \24423 , \24424 , \24425 , \24426 , \24427 , \24428 , \24429 , \24430 , \24431 , \24432 ,
         \24433 , \24434 , \24435 , \24436 , \24437 , \24438 , \24439 , \24440 , \24441 , \24442 ,
         \24443 , \24444 , \24445 , \24446 , \24447 , \24448 , \24449 , \24450 , \24451 , \24452 ,
         \24453 , \24454 , \24455 , \24456 , \24457 , \24458 , \24459 , \24460 , \24461 , \24462 ,
         \24463 , \24464 , \24465 , \24466 , \24467 , \24468 , \24469 , \24470 , \24471 , \24472 ,
         \24473 , \24474 , \24475 , \24476 , \24477 , \24478 , \24479 , \24480 , \24481 , \24482 ,
         \24483 , \24484 , \24485 , \24486 , \24487 , \24488 , \24489 , \24490 , \24491 , \24492 ,
         \24493 , \24494 , \24495 , \24496 , \24497 , \24498 , \24499 , \24500 , \24501 , \24502 ,
         \24503 , \24504 , \24505 , \24506 , \24507 , \24508 , \24509 , \24510 , \24511 , \24512 ,
         \24513 , \24514 , \24515 , \24516 , \24517 , \24518 , \24519 , \24520 , \24521 , \24522 ,
         \24523 , \24524 , \24525 , \24526 , \24527 , \24528 , \24529 , \24530 , \24531 , \24532 ,
         \24533 , \24534 , \24535 , \24536 , \24537 , \24538 , \24539 , \24540 , \24541 , \24542 ,
         \24543 , \24544 , \24545 , \24546 , \24547 , \24548 , \24549 , \24550 , \24551 , \24552 ,
         \24553 , \24554 , \24555 , \24556 , \24557 , \24558 , \24559 , \24560 , \24561 , \24562 ,
         \24563 , \24564 , \24565 , \24566 , \24567 , \24568 , \24569 , \24570 , \24571 , \24572 ,
         \24573 , \24574 , \24575 , \24576 , \24577 , \24578 , \24579 , \24580 , \24581 , \24582 ,
         \24583 , \24584 , \24585 , \24586 , \24587 , \24588 , \24589 , \24590 , \24591 , \24592 ,
         \24593 , \24594 , \24595 , \24596 , \24597 , \24598 , \24599 , \24600 , \24601 , \24602 ,
         \24603 , \24604 , \24605 , \24606 , \24607 , \24608 , \24609 , \24610 , \24611 , \24612 ,
         \24613 , \24614 , \24615 , \24616 , \24617 , \24618 , \24619 , \24620 , \24621 , \24622 ,
         \24623 , \24624 , \24625 , \24626 , \24627 , \24628 , \24629 , \24630 , \24631 , \24632 ,
         \24633 , \24634 , \24635 , \24636 , \24637 , \24638 , \24639 , \24640 , \24641 , \24642 ,
         \24643 , \24644 , \24645 , \24646 , \24647 , \24648 , \24649 , \24650 , \24651 , \24652 ,
         \24653 , \24654 , \24655 , \24656 , \24657 , \24658 , \24659 , \24660 , \24661 , \24662 ,
         \24663 , \24664 , \24665 , \24666 , \24667 , \24668 , \24669 , \24670 , \24671 , \24672 ,
         \24673 , \24674 , \24675 , \24676 , \24677 , \24678 , \24679 , \24680 , \24681 , \24682 ,
         \24683 , \24684 , \24685 , \24686 , \24687 , \24688 , \24689 , \24690 , \24691 , \24692 ,
         \24693 , \24694 , \24695 , \24696 , \24697 , \24698 , \24699 , \24700 , \24701 , \24702 ,
         \24703 , \24704 , \24705 , \24706 , \24707 , \24708 , \24709 , \24710 , \24711 , \24712 ,
         \24713 , \24714 , \24715 , \24716 , \24717 , \24718 , \24719 , \24720 , \24721 , \24722 ,
         \24723 , \24724 , \24725 , \24726 , \24727 , \24728 , \24729 , \24730 , \24731 , \24732 ,
         \24733 , \24734 , \24735 , \24736 , \24737 , \24738 , \24739 , \24740 , \24741 , \24742 ,
         \24743 , \24744 , \24745 , \24746 , \24747 , \24748 , \24749 , \24750 , \24751 , \24752 ,
         \24753 , \24754 , \24755 , \24756 , \24757 , \24758 , \24759 , \24760 , \24761 , \24762 ,
         \24763 , \24764 , \24765 , \24766 , \24767 , \24768 , \24769 , \24770 , \24771 , \24772 ,
         \24773 , \24774 , \24775 , \24776 , \24777 , \24778 , \24779 , \24780 , \24781 , \24782 ,
         \24783 , \24784 , \24785 , \24786 , \24787 , \24788 , \24789 , \24790 , \24791 , \24792 ,
         \24793 , \24794 , \24795 , \24796 , \24797 , \24798 , \24799 , \24800 , \24801 , \24802 ,
         \24803 , \24804 , \24805 , \24806 , \24807 , \24808 , \24809 , \24810 , \24811 , \24812 ,
         \24813 , \24814 , \24815 , \24816 , \24817 , \24818 , \24819 , \24820 , \24821 , \24822 ,
         \24823 , \24824 , \24825 , \24826 , \24827 , \24828 , \24829 , \24830 , \24831 , \24832 ,
         \24833 , \24834 , \24835 , \24836 , \24837 , \24838 , \24839 , \24840 , \24841 , \24842 ,
         \24843 , \24844 , \24845 , \24846 , \24847 , \24848 , \24849 , \24850 , \24851 , \24852 ,
         \24853 , \24854 , \24855 , \24856 , \24857 , \24858 , \24859 , \24860 , \24861 , \24862 ,
         \24863 , \24864 , \24865 , \24866 , \24867 , \24868 , \24869 , \24870 , \24871 , \24872 ,
         \24873 , \24874 , \24875 , \24876 , \24877 , \24878 , \24879 , \24880 , \24881 , \24882 ,
         \24883 , \24884 , \24885 , \24886 , \24887 , \24888 , \24889 , \24890 , \24891 , \24892 ,
         \24893 , \24894 , \24895 , \24896 , \24897 , \24898 , \24899 , \24900 , \24901 , \24902 ,
         \24903 , \24904 , \24905 , \24906 , \24907 , \24908 , \24909 , \24910 , \24911 , \24912 ,
         \24913 , \24914 , \24915 , \24916 , \24917 , \24918 , \24919 , \24920 , \24921 , \24922 ,
         \24923 , \24924 , \24925 , \24926 , \24927 , \24928 , \24929 , \24930 , \24931 , \24932 ,
         \24933 , \24934 , \24935 , \24936 , \24937 , \24938 , \24939 , \24940 , \24941 , \24942 ,
         \24943 , \24944 , \24945 , \24946 , \24947 , \24948 , \24949 , \24950 , \24951 , \24952 ,
         \24953 , \24954 , \24955 , \24956 , \24957 , \24958 , \24959 , \24960 , \24961 , \24962 ,
         \24963 , \24964 , \24965 , \24966 , \24967 , \24968 , \24969 , \24970 , \24971 , \24972 ,
         \24973 , \24974 , \24975 , \24976 , \24977 , \24978 , \24979 , \24980 , \24981 , \24982 ,
         \24983 , \24984 , \24985 , \24986 , \24987 , \24988 , \24989 , \24990 , \24991 , \24992 ,
         \24993 , \24994 , \24995 , \24996 , \24997 , \24998 , \24999 , \25000 , \25001 , \25002 ,
         \25003 , \25004 , \25005 , \25006 , \25007 , \25008 , \25009 , \25010 , \25011 , \25012 ,
         \25013 , \25014 , \25015 , \25016 , \25017 , \25018 , \25019 , \25020 , \25021 , \25022 ,
         \25023 , \25024 , \25025 , \25026 , \25027 , \25028 , \25029 , \25030 , \25031 , \25032 ,
         \25033 , \25034 , \25035 , \25036 , \25037 , \25038 , \25039 , \25040 , \25041 , \25042 ,
         \25043 , \25044 , \25045 , \25046 , \25047 , \25048 , \25049 , \25050 , \25051 , \25052 ,
         \25053 , \25054 , \25055 , \25056 , \25057 , \25058 , \25059 , \25060 , \25061 , \25062 ,
         \25063 , \25064 , \25065 , \25066 , \25067 , \25068 , \25069 , \25070 , \25071 , \25072 ,
         \25073 , \25074 , \25075 , \25076 , \25077 , \25078 , \25079 , \25080 , \25081 , \25082 ,
         \25083 , \25084 , \25085 , \25086 , \25087 , \25088 , \25089 , \25090 , \25091 , \25092 ,
         \25093 , \25094 , \25095 , \25096 , \25097 , \25098 , \25099 , \25100 , \25101 , \25102 ,
         \25103 , \25104 , \25105 , \25106 , \25107 , \25108 , \25109 , \25110 , \25111 , \25112 ,
         \25113 , \25114 , \25115 , \25116 , \25117 , \25118 , \25119 , \25120 , \25121 , \25122 ,
         \25123 , \25124 , \25125 , \25126 , \25127 , \25128 , \25129 , \25130 , \25131 , \25132 ,
         \25133 , \25134 , \25135 , \25136 , \25137 , \25138 , \25139 , \25140 , \25141 , \25142 ,
         \25143 , \25144 , \25145 , \25146 , \25147 , \25148 , \25149 , \25150 , \25151 , \25152 ,
         \25153 , \25154 , \25155 , \25156 , \25157 , \25158 , \25159 , \25160 , \25161 , \25162 ,
         \25163 , \25164 , \25165 , \25166 , \25167 , \25168 , \25169 , \25170 , \25171 , \25172 ,
         \25173 , \25174 , \25175 , \25176 , \25177 , \25178 , \25179 , \25180 , \25181 , \25182 ,
         \25183 , \25184 , \25185 , \25186 , \25187 , \25188 , \25189 , \25190 , \25191 , \25192 ,
         \25193 , \25194 , \25195 , \25196 , \25197 , \25198 , \25199 , \25200 , \25201 , \25202 ,
         \25203 , \25204 , \25205 , \25206 , \25207 , \25208 , \25209 , \25210 , \25211 , \25212 ,
         \25213 , \25214 , \25215 , \25216 , \25217 , \25218 , \25219 , \25220 , \25221 , \25222 ,
         \25223 , \25224 , \25225 , \25226 , \25227 , \25228 , \25229 , \25230 , \25231 , \25232 ,
         \25233 , \25234 , \25235 , \25236 , \25237 , \25238 , \25239 , \25240 , \25241 , \25242 ,
         \25243 , \25244 , \25245 , \25246 , \25247 , \25248 , \25249 , \25250 , \25251 , \25252 ,
         \25253 , \25254 , \25255 , \25256 , \25257 , \25258 , \25259 , \25260 , \25261 , \25262 ,
         \25263 , \25264 , \25265 , \25266 , \25267 , \25268 , \25269 , \25270 , \25271 , \25272 ,
         \25273 , \25274 , \25275 , \25276 , \25277 , \25278 , \25279 , \25280 , \25281 , \25282 ,
         \25283 , \25284 , \25285 , \25286 , \25287 , \25288 , \25289 , \25290 , \25291 , \25292 ,
         \25293 , \25294 , \25295 , \25296 , \25297 , \25298 , \25299 , \25300 , \25301 , \25302 ,
         \25303 , \25304 , \25305 , \25306 , \25307 , \25308 , \25309 , \25310 , \25311 , \25312 ,
         \25313 , \25314 , \25315 , \25316 , \25317 , \25318 , \25319 , \25320 , \25321 , \25322 ,
         \25323 , \25324 , \25325 , \25326 , \25327 , \25328 , \25329 , \25330 , \25331 , \25332 ,
         \25333 , \25334 , \25335 , \25336 , \25337 , \25338 , \25339 , \25340 , \25341 , \25342 ,
         \25343 , \25344 , \25345 , \25346 , \25347 , \25348 , \25349 , \25350 , \25351 , \25352 ,
         \25353 , \25354 , \25355 , \25356 , \25357 , \25358 , \25359 , \25360 , \25361 , \25362 ,
         \25363 , \25364 , \25365 , \25366 , \25367 , \25368 , \25369 , \25370 , \25371 , \25372 ,
         \25373 , \25374 , \25375 , \25376 , \25377 , \25378 , \25379 , \25380 , \25381 , \25382 ,
         \25383 , \25384 , \25385 , \25386 , \25387 , \25388 , \25389 , \25390 , \25391 , \25392 ,
         \25393 , \25394 , \25395 , \25396 , \25397 , \25398 , \25399 , \25400 , \25401 , \25402 ,
         \25403 , \25404 , \25405 , \25406 , \25407 , \25408 , \25409 , \25410 , \25411 , \25412 ,
         \25413 , \25414 , \25415 , \25416 , \25417 , \25418 , \25419 , \25420 , \25421 , \25422 ,
         \25423 , \25424 , \25425 , \25426 , \25427 , \25428 , \25429 , \25430 , \25431 , \25432 ,
         \25433 , \25434 , \25435 , \25436 , \25437 , \25438 , \25439 , \25440 , \25441 , \25442 ,
         \25443 , \25444 , \25445 , \25446 , \25447 , \25448 , \25449 , \25450 , \25451 , \25452 ,
         \25453 , \25454 , \25455 , \25456 , \25457 , \25458 , \25459 , \25460 , \25461 , \25462 ,
         \25463 , \25464 , \25465 , \25466 , \25467 , \25468 , \25469 , \25470 , \25471 , \25472 ,
         \25473 , \25474 , \25475 , \25476 , \25477 , \25478 , \25479 , \25480 , \25481 , \25482 ,
         \25483 , \25484 , \25485 , \25486 , \25487 , \25488 , \25489 , \25490 , \25491 , \25492 ,
         \25493 , \25494 , \25495 , \25496 , \25497 , \25498 , \25499 , \25500 , \25501 , \25502 ,
         \25503 , \25504 , \25505 , \25506 , \25507 , \25508 , \25509 , \25510 , \25511 , \25512 ,
         \25513 , \25514 , \25515 , \25516 , \25517 , \25518 , \25519 , \25520 , \25521 , \25522 ,
         \25523 , \25524 , \25525 , \25526 , \25527 , \25528 , \25529 , \25530 , \25531 , \25532 ,
         \25533 , \25534 , \25535 , \25536 , \25537 , \25538 , \25539 , \25540 , \25541 , \25542 ,
         \25543 , \25544 , \25545 , \25546 , \25547 , \25548 , \25549 , \25550 , \25551 , \25552 ,
         \25553 , \25554 , \25555 , \25556 , \25557 , \25558 , \25559 , \25560 , \25561 , \25562 ,
         \25563 , \25564 , \25565 , \25566 , \25567 , \25568 , \25569 , \25570 , \25571 , \25572 ,
         \25573 , \25574 , \25575 , \25576 , \25577 , \25578 , \25579 , \25580 , \25581 , \25582 ,
         \25583 , \25584 , \25585 , \25586 , \25587 , \25588 , \25589 , \25590 , \25591 , \25592 ,
         \25593 , \25594 , \25595 , \25596 , \25597 , \25598 , \25599 , \25600 , \25601 , \25602 ,
         \25603 , \25604 , \25605 , \25606 , \25607 , \25608 , \25609 , \25610 , \25611 , \25612 ,
         \25613 , \25614 , \25615 , \25616 , \25617 , \25618 , \25619 , \25620 , \25621 , \25622 ,
         \25623 , \25624 , \25625 , \25626 , \25627 , \25628 , \25629 , \25630 , \25631 , \25632 ,
         \25633 , \25634 , \25635 , \25636 , \25637 , \25638 , \25639 , \25640 , \25641 , \25642 ,
         \25643 , \25644 , \25645 , \25646 , \25647 , \25648 , \25649 , \25650 , \25651 , \25652 ,
         \25653 , \25654 , \25655 , \25656 , \25657 , \25658 , \25659 , \25660 , \25661 , \25662 ,
         \25663 , \25664 , \25665 , \25666 , \25667 , \25668 , \25669 , \25670 , \25671 , \25672 ,
         \25673 , \25674 , \25675 , \25676 , \25677 , \25678 , \25679 , \25680 , \25681 , \25682 ,
         \25683 , \25684 , \25685 , \25686 , \25687 , \25688 , \25689 , \25690 , \25691 , \25692 ,
         \25693 , \25694 , \25695 , \25696 , \25697 , \25698 , \25699 , \25700 , \25701 , \25702 ,
         \25703 , \25704 , \25705 , \25706 , \25707 , \25708 , \25709 , \25710 , \25711 , \25712 ,
         \25713 , \25714 , \25715 , \25716 , \25717 , \25718 , \25719 , \25720 , \25721 , \25722 ,
         \25723 , \25724 , \25725 , \25726 , \25727 , \25728 , \25729 , \25730 , \25731 , \25732 ,
         \25733 , \25734 , \25735 , \25736 , \25737 , \25738 , \25739 , \25740 , \25741 , \25742 ,
         \25743 , \25744 , \25745 , \25746 , \25747 , \25748 , \25749 , \25750 , \25751 , \25752 ,
         \25753 , \25754 , \25755 , \25756 , \25757 , \25758 , \25759 , \25760 , \25761 , \25762 ,
         \25763 , \25764 , \25765 , \25766 , \25767 , \25768 , \25769 , \25770 , \25771 , \25772 ,
         \25773 , \25774 , \25775 , \25776 , \25777 , \25778 , \25779 , \25780 , \25781 , \25782 ,
         \25783 , \25784 , \25785 , \25786 , \25787 , \25788 , \25789 , \25790 , \25791 , \25792 ,
         \25793 , \25794 , \25795 , \25796 , \25797 , \25798 , \25799 , \25800 , \25801 , \25802 ,
         \25803 , \25804 , \25805 , \25806 , \25807 , \25808 , \25809 , \25810 , \25811 , \25812 ,
         \25813 , \25814 , \25815 , \25816 , \25817 , \25818 , \25819 , \25820 , \25821 , \25822 ,
         \25823 , \25824 , \25825 , \25826 , \25827 , \25828 , \25829 , \25830 , \25831 , \25832 ,
         \25833 , \25834 , \25835 , \25836 , \25837 , \25838 , \25839 , \25840 , \25841 , \25842 ,
         \25843 , \25844 , \25845 , \25846 , \25847 , \25848 , \25849 , \25850 , \25851 , \25852 ,
         \25853 , \25854 , \25855 , \25856 , \25857 , \25858 , \25859 , \25860 , \25861 , \25862 ,
         \25863 , \25864 , \25865 , \25866 , \25867 , \25868 , \25869 , \25870 , \25871 , \25872 ,
         \25873 , \25874 , \25875 , \25876 , \25877 , \25878 , \25879 , \25880 , \25881 , \25882 ,
         \25883 , \25884 , \25885 , \25886 , \25887 , \25888 , \25889 , \25890 , \25891 , \25892 ,
         \25893 , \25894 , \25895 , \25896 , \25897 , \25898 , \25899 , \25900 , \25901 , \25902 ,
         \25903 , \25904 , \25905 , \25906 , \25907 , \25908 , \25909 , \25910 , \25911 , \25912 ,
         \25913 , \25914 , \25915 , \25916 , \25917 , \25918 , \25919 , \25920 , \25921 , \25922 ,
         \25923 , \25924 , \25925 , \25926 , \25927 , \25928 , \25929 , \25930 , \25931 , \25932 ,
         \25933 , \25934 , \25935 , \25936 , \25937 , \25938 , \25939 , \25940 , \25941 , \25942 ,
         \25943 , \25944 , \25945 , \25946 , \25947 , \25948 , \25949 , \25950 , \25951 , \25952 ,
         \25953 , \25954 , \25955 , \25956 , \25957 , \25958 , \25959 , \25960 , \25961 , \25962 ,
         \25963 , \25964 , \25965 , \25966 , \25967 , \25968 , \25969 , \25970 , \25971 , \25972 ,
         \25973 , \25974 , \25975 , \25976 , \25977 , \25978 , \25979 , \25980 , \25981 , \25982 ,
         \25983 , \25984 , \25985 , \25986 , \25987 , \25988 , \25989 , \25990 , \25991 , \25992 ,
         \25993 , \25994 , \25995 , \25996 , \25997 , \25998 , \25999 , \26000 , \26001 , \26002 ,
         \26003 , \26004 , \26005 , \26006 , \26007 , \26008 , \26009 , \26010 , \26011 , \26012 ,
         \26013 , \26014 , \26015 , \26016 , \26017 , \26018 , \26019 , \26020 , \26021 , \26022 ,
         \26023 , \26024 , \26025 , \26026 , \26027 , \26028 , \26029 , \26030 , \26031 , \26032 ,
         \26033 , \26034 , \26035 , \26036 , \26037 , \26038 , \26039 , \26040 , \26041 , \26042 ,
         \26043 , \26044 , \26045 , \26046 , \26047 , \26048 , \26049 , \26050 , \26051 , \26052 ,
         \26053 , \26054 , \26055 , \26056 , \26057 , \26058 , \26059 , \26060 , \26061 , \26062 ,
         \26063 , \26064 , \26065 , \26066 , \26067 , \26068 , \26069 , \26070 , \26071 , \26072 ,
         \26073 , \26074 , \26075 , \26076 , \26077 , \26078 , \26079 , \26080 , \26081 , \26082 ,
         \26083 , \26084 , \26085 , \26086 , \26087 , \26088 , \26089 , \26090 , \26091 , \26092 ,
         \26093 , \26094 , \26095 , \26096 , \26097 , \26098 , \26099 , \26100 , \26101 , \26102 ,
         \26103 , \26104 , \26105 , \26106 , \26107 , \26108 , \26109 , \26110 , \26111 , \26112 ,
         \26113 , \26114 , \26115 , \26116 , \26117 , \26118 , \26119 , \26120 , \26121 , \26122 ,
         \26123 , \26124 , \26125 , \26126 , \26127 , \26128 , \26129 , \26130 , \26131 , \26132 ,
         \26133 , \26134 , \26135 , \26136 , \26137 , \26138 , \26139 , \26140 , \26141 , \26142 ,
         \26143 , \26144 , \26145 , \26146 , \26147 , \26148 , \26149 , \26150 , \26151 , \26152 ,
         \26153 , \26154 , \26155 , \26156 , \26157 , \26158 , \26159 , \26160 , \26161 , \26162 ,
         \26163 , \26164 , \26165 , \26166 , \26167 , \26168 , \26169 , \26170 , \26171 , \26172 ,
         \26173 , \26174 , \26175 , \26176 , \26177 , \26178 , \26179 , \26180 , \26181 , \26182 ,
         \26183 , \26184 , \26185 , \26186 , \26187 , \26188 , \26189 , \26190 , \26191 , \26192 ,
         \26193 , \26194 , \26195 , \26196 , \26197 , \26198 , \26199 , \26200 , \26201 , \26202 ,
         \26203 , \26204 , \26205 , \26206 , \26207 , \26208 , \26209 , \26210 , \26211 , \26212 ,
         \26213 , \26214 , \26215 , \26216 , \26217 , \26218 , \26219 , \26220 , \26221 , \26222 ,
         \26223 , \26224 , \26225 , \26226 , \26227 , \26228 , \26229 , \26230 , \26231 , \26232 ,
         \26233 , \26234 , \26235 , \26236 , \26237 , \26238 , \26239 , \26240 , \26241 , \26242 ,
         \26243 , \26244 , \26245 , \26246 , \26247 , \26248 , \26249 , \26250 , \26251 , \26252 ,
         \26253 , \26254 , \26255 , \26256 , \26257 , \26258 , \26259 , \26260 , \26261 , \26262 ,
         \26263 , \26264 , \26265 , \26266 , \26267 , \26268 , \26269 , \26270 , \26271 , \26272 ,
         \26273 , \26274 , \26275 , \26276 , \26277 , \26278 , \26279 , \26280 , \26281 , \26282 ,
         \26283 , \26284 , \26285 , \26286 , \26287 , \26288 , \26289 , \26290 , \26291 , \26292 ,
         \26293 , \26294 , \26295 , \26296 , \26297 , \26298 , \26299 , \26300 , \26301 , \26302 ,
         \26303 , \26304 , \26305 , \26306 , \26307 , \26308 , \26309 , \26310 , \26311 , \26312 ,
         \26313 , \26314 , \26315 , \26316 , \26317 , \26318 , \26319 , \26320 , \26321 , \26322 ,
         \26323 , \26324 , \26325 , \26326 , \26327 , \26328 , \26329 , \26330 , \26331 , \26332 ,
         \26333 , \26334 , \26335 , \26336 , \26337 , \26338 , \26339 , \26340 , \26341 , \26342 ,
         \26343 , \26344 , \26345 , \26346 , \26347 , \26348 , \26349 , \26350 , \26351 , \26352 ,
         \26353 , \26354 , \26355 , \26356 , \26357 , \26358 , \26359 , \26360 , \26361 , \26362 ,
         \26363 , \26364 , \26365 , \26366 , \26367 , \26368 , \26369 , \26370 , \26371 , \26372 ,
         \26373 , \26374 , \26375 , \26376 , \26377 , \26378 , \26379 , \26380 , \26381 , \26382 ,
         \26383 , \26384 , \26385 , \26386 , \26387 , \26388 , \26389 , \26390 , \26391 , \26392 ,
         \26393 , \26394 , \26395 , \26396 , \26397 , \26398 , \26399 , \26400 , \26401 , \26402 ,
         \26403 , \26404 , \26405 , \26406 , \26407 , \26408 , \26409 , \26410 , \26411 , \26412 ,
         \26413 , \26414 , \26415 , \26416 , \26417 , \26418 , \26419 , \26420 , \26421 , \26422 ,
         \26423 , \26424 , \26425 , \26426 , \26427 , \26428 , \26429 , \26430 , \26431 , \26432 ,
         \26433 , \26434 , \26435 , \26436 , \26437 , \26438 , \26439 , \26440 , \26441 , \26442 ,
         \26443 , \26444 , \26445 , \26446 , \26447 , \26448 , \26449 , \26450 , \26451 , \26452 ,
         \26453 , \26454 , \26455 , \26456 , \26457 , \26458 , \26459 , \26460 , \26461 , \26462 ,
         \26463 , \26464 , \26465 , \26466 , \26467 , \26468 , \26469 , \26470 , \26471 , \26472 ,
         \26473 , \26474 , \26475 , \26476 , \26477 , \26478 , \26479 , \26480 , \26481 , \26482 ,
         \26483 , \26484 , \26485 , \26486 , \26487 , \26488 , \26489 , \26490 , \26491 , \26492 ,
         \26493 , \26494 , \26495 , \26496 , \26497 , \26498 , \26499 , \26500 , \26501 , \26502 ,
         \26503 , \26504 , \26505 , \26506 , \26507 , \26508 , \26509 , \26510 , \26511 , \26512 ,
         \26513 , \26514 , \26515 , \26516 , \26517 , \26518 , \26519 , \26520 , \26521 , \26522 ,
         \26523 , \26524 , \26525 , \26526 , \26527 , \26528 , \26529 , \26530 , \26531 , \26532 ,
         \26533 , \26534 , \26535 , \26536 , \26537 , \26538 , \26539 , \26540 , \26541 , \26542 ,
         \26543 , \26544 , \26545 , \26546 , \26547 , \26548 , \26549 , \26550 , \26551 , \26552 ,
         \26553 , \26554 , \26555 , \26556 , \26557 , \26558 , \26559 , \26560 , \26561 , \26562 ,
         \26563 , \26564 , \26565 , \26566 , \26567 , \26568 , \26569 , \26570 , \26571 , \26572 ,
         \26573 , \26574 , \26575 , \26576 , \26577 , \26578 , \26579 , \26580 , \26581 , \26582 ,
         \26583 , \26584 , \26585 , \26586 , \26587 , \26588 , \26589 , \26590 , \26591 , \26592 ,
         \26593 , \26594 , \26595 , \26596 , \26597 , \26598 , \26599 , \26600 , \26601 , \26602 ,
         \26603 , \26604 , \26605 , \26606 , \26607 , \26608 , \26609 , \26610 , \26611 , \26612 ,
         \26613 , \26614 , \26615 , \26616 , \26617 , \26618 , \26619 , \26620 , \26621 , \26622 ,
         \26623 , \26624 , \26625 , \26626 , \26627 , \26628 , \26629 , \26630 , \26631 , \26632 ,
         \26633 , \26634 , \26635 , \26636 , \26637 , \26638 , \26639 , \26640 , \26641 , \26642 ,
         \26643 , \26644 , \26645 , \26646 , \26647 , \26648 , \26649 , \26650 , \26651 , \26652 ,
         \26653 , \26654 , \26655 , \26656 , \26657 , \26658 , \26659 , \26660 , \26661 , \26662 ,
         \26663 , \26664 , \26665 , \26666 , \26667 , \26668 , \26669 , \26670 , \26671 , \26672 ,
         \26673 , \26674 , \26675 , \26676 , \26677 , \26678 , \26679 , \26680 , \26681 , \26682 ,
         \26683 , \26684 , \26685 , \26686 , \26687 , \26688 , \26689 , \26690 , \26691 , \26692 ,
         \26693 , \26694 , \26695 , \26696 , \26697 , \26698 , \26699 , \26700 , \26701 , \26702 ,
         \26703 , \26704 , \26705 , \26706 , \26707 , \26708 , \26709 , \26710 , \26711 , \26712 ,
         \26713 , \26714 , \26715 , \26716 , \26717 , \26718 , \26719 , \26720 , \26721 , \26722 ,
         \26723 , \26724 , \26725 , \26726 , \26727 , \26728 , \26729 , \26730 , \26731 , \26732 ,
         \26733 , \26734 , \26735 , \26736 , \26737 , \26738 , \26739 , \26740 , \26741 , \26742 ,
         \26743 , \26744 , \26745 , \26746 , \26747 , \26748 , \26749 , \26750 , \26751 , \26752 ,
         \26753 , \26754 , \26755 , \26756 , \26757 , \26758 , \26759 , \26760 , \26761 , \26762 ,
         \26763 , \26764 , \26765 , \26766 , \26767 , \26768 , \26769 , \26770 , \26771 , \26772 ,
         \26773 , \26774 , \26775 , \26776 , \26777 , \26778 , \26779 , \26780 , \26781 , \26782 ,
         \26783 , \26784 , \26785 , \26786 , \26787 , \26788 , \26789 , \26790 , \26791 , \26792 ,
         \26793 , \26794 , \26795 , \26796 , \26797 , \26798 , \26799 , \26800 , \26801 , \26802 ,
         \26803 , \26804 , \26805 , \26806 , \26807 , \26808 , \26809 , \26810 , \26811 , \26812 ,
         \26813 , \26814 , \26815 , \26816 , \26817 , \26818 , \26819 , \26820 , \26821 , \26822 ,
         \26823 , \26824 , \26825 , \26826 , \26827 , \26828 , \26829 , \26830 , \26831 , \26832 ,
         \26833 , \26834 , \26835 , \26836 , \26837 , \26838 , \26839 , \26840 , \26841 , \26842 ,
         \26843 , \26844 , \26845 , \26846 , \26847 , \26848 , \26849 , \26850 , \26851 , \26852 ,
         \26853 , \26854 , \26855 , \26856 , \26857 , \26858 , \26859 , \26860 , \26861 , \26862 ,
         \26863 , \26864 , \26865 , \26866 , \26867 , \26868 , \26869 , \26870 , \26871 , \26872 ,
         \26873 , \26874 , \26875 , \26876 , \26877 , \26878 , \26879 , \26880 , \26881 , \26882 ,
         \26883 , \26884 , \26885 , \26886 , \26887 , \26888 , \26889 , \26890 , \26891 , \26892 ,
         \26893 , \26894 , \26895 , \26896 , \26897 , \26898 , \26899 , \26900 , \26901 , \26902 ,
         \26903 , \26904 , \26905 , \26906 , \26907 , \26908 , \26909 , \26910 , \26911 , \26912 ,
         \26913 , \26914 , \26915 , \26916 , \26917 , \26918 , \26919 , \26920 , \26921 , \26922 ,
         \26923 , \26924 , \26925 , \26926 , \26927 , \26928 , \26929 , \26930 , \26931 , \26932 ,
         \26933 , \26934 , \26935 , \26936 , \26937 , \26938 , \26939 , \26940 , \26941 , \26942 ,
         \26943 , \26944 , \26945 , \26946 , \26947 , \26948 , \26949 , \26950 , \26951 , \26952 ,
         \26953 , \26954 , \26955 , \26956 , \26957 , \26958 , \26959 , \26960 , \26961 , \26962 ,
         \26963 , \26964 , \26965 , \26966 , \26967 , \26968 , \26969 , \26970 , \26971 , \26972 ,
         \26973 , \26974 , \26975 , \26976 , \26977 , \26978 , \26979 , \26980 , \26981 , \26982 ,
         \26983 , \26984 , \26985 , \26986 , \26987 , \26988 , \26989 , \26990 , \26991 , \26992 ,
         \26993 , \26994 , \26995 , \26996 , \26997 , \26998 , \26999 , \27000 , \27001 , \27002 ,
         \27003 , \27004 , \27005 , \27006 , \27007 , \27008 , \27009 , \27010 , \27011 , \27012 ,
         \27013 , \27014 , \27015 , \27016 , \27017 , \27018 , \27019 , \27020 , \27021 , \27022 ,
         \27023 , \27024 , \27025 , \27026 , \27027 , \27028 , \27029 , \27030 , \27031 , \27032 ,
         \27033 , \27034 , \27035 , \27036 , \27037 , \27038 , \27039 , \27040 , \27041 , \27042 ,
         \27043 , \27044 , \27045 , \27046 , \27047 , \27048 , \27049 , \27050 , \27051 , \27052 ,
         \27053 , \27054 , \27055 , \27056 , \27057 , \27058 , \27059 , \27060 , \27061 , \27062 ,
         \27063 , \27064 , \27065 , \27066 , \27067 , \27068 , \27069 , \27070 , \27071 , \27072 ,
         \27073 , \27074 , \27075 , \27076 , \27077 , \27078 , \27079 , \27080 , \27081 , \27082 ,
         \27083 , \27084 , \27085 , \27086 , \27087 , \27088 , \27089 , \27090 , \27091 , \27092 ,
         \27093 , \27094 , \27095 , \27096 , \27097 , \27098 , \27099 , \27100 , \27101 , \27102 ,
         \27103 , \27104 , \27105 , \27106 , \27107 , \27108 , \27109 , \27110 , \27111 , \27112 ,
         \27113 , \27114 , \27115 , \27116 , \27117 , \27118 , \27119 , \27120 , \27121 , \27122 ,
         \27123 , \27124 , \27125 , \27126 , \27127 , \27128 , \27129 , \27130 , \27131 , \27132 ,
         \27133 , \27134 , \27135 , \27136 , \27137 , \27138 , \27139 , \27140 , \27141 , \27142 ,
         \27143 , \27144 , \27145 , \27146 , \27147 , \27148 , \27149 , \27150 , \27151 , \27152 ,
         \27153 , \27154 , \27155 , \27156 , \27157 , \27158 , \27159 , \27160 , \27161 , \27162 ,
         \27163 , \27164 , \27165 , \27166 , \27167 , \27168 , \27169 , \27170 , \27171 , \27172 ,
         \27173 , \27174 , \27175 , \27176 , \27177 , \27178 , \27179 , \27180 , \27181 , \27182 ,
         \27183 , \27184 , \27185 , \27186 , \27187 , \27188 , \27189 , \27190 , \27191 , \27192 ,
         \27193 , \27194 , \27195 , \27196 , \27197 , \27198 , \27199 , \27200 , \27201 , \27202 ,
         \27203 , \27204 , \27205 , \27206 , \27207 , \27208 , \27209 , \27210 , \27211 , \27212 ,
         \27213 , \27214 , \27215 , \27216 , \27217 , \27218 , \27219 , \27220 , \27221 , \27222 ,
         \27223 , \27224 , \27225 , \27226 , \27227 , \27228 , \27229 , \27230 , \27231 , \27232 ,
         \27233 , \27234 , \27235 , \27236 , \27237 , \27238 , \27239 , \27240 , \27241 , \27242 ,
         \27243 , \27244 , \27245 , \27246 , \27247 , \27248 , \27249 , \27250 , \27251 , \27252 ,
         \27253 , \27254 , \27255 , \27256 , \27257 , \27258 , \27259 , \27260 , \27261 , \27262 ,
         \27263 , \27264 , \27265 , \27266 , \27267 , \27268 , \27269 , \27270 , \27271 , \27272 ,
         \27273 , \27274 , \27275 , \27276 , \27277 , \27278 , \27279 , \27280 , \27281 , \27282 ,
         \27283 , \27284 , \27285 , \27286 , \27287 , \27288 , \27289 , \27290 , \27291 , \27292 ,
         \27293 , \27294 , \27295 , \27296 , \27297 , \27298 , \27299 , \27300 , \27301 , \27302 ,
         \27303 , \27304 , \27305 , \27306 , \27307 , \27308 , \27309 , \27310 , \27311 , \27312 ,
         \27313 , \27314 , \27315 , \27316 , \27317 , \27318 , \27319 , \27320 , \27321 , \27322 ,
         \27323 , \27324 , \27325 , \27326 , \27327 , \27328 , \27329 , \27330 , \27331 , \27332 ,
         \27333 , \27334 , \27335 , \27336 , \27337 , \27338 , \27339 , \27340 , \27341 , \27342 ,
         \27343 , \27344 , \27345 , \27346 , \27347 , \27348 , \27349 , \27350 , \27351 , \27352 ,
         \27353 , \27354 , \27355 , \27356 , \27357 , \27358 , \27359 , \27360 , \27361 , \27362 ,
         \27363 , \27364 , \27365 , \27366 , \27367 , \27368 , \27369 , \27370 , \27371 , \27372 ,
         \27373 , \27374 , \27375 , \27376 , \27377 , \27378 , \27379 , \27380 , \27381 , \27382 ,
         \27383 , \27384 , \27385 , \27386 , \27387 , \27388 , \27389 , \27390 , \27391 , \27392 ,
         \27393 , \27394 , \27395 , \27396 , \27397 , \27398 , \27399 , \27400 , \27401 , \27402 ,
         \27403 , \27404 , \27405 , \27406 , \27407 , \27408 , \27409 , \27410 , \27411 , \27412 ,
         \27413 , \27414 , \27415 , \27416 , \27417 , \27418 , \27419 , \27420 , \27421 , \27422 ,
         \27423 , \27424 , \27425 , \27426 , \27427 , \27428 , \27429 , \27430 , \27431 , \27432 ,
         \27433 , \27434 , \27435 , \27436 , \27437 , \27438 , \27439 , \27440 , \27441 , \27442 ,
         \27443 , \27444 , \27445 , \27446 , \27447 , \27448 , \27449 , \27450 , \27451 , \27452 ,
         \27453 , \27454 , \27455 , \27456 , \27457 , \27458 , \27459 , \27460 , \27461 , \27462 ,
         \27463 , \27464 , \27465 , \27466 , \27467 , \27468 , \27469 , \27470 , \27471 , \27472 ,
         \27473 , \27474 , \27475 , \27476 , \27477 , \27478 , \27479 , \27480 , \27481 , \27482 ,
         \27483 , \27484 , \27485 , \27486 , \27487 , \27488 , \27489 , \27490 , \27491 , \27492 ,
         \27493 , \27494 , \27495 , \27496 , \27497 , \27498 , \27499 , \27500 , \27501 , \27502 ,
         \27503 , \27504 , \27505 , \27506 , \27507 , \27508 , \27509 , \27510 , \27511 , \27512 ,
         \27513 , \27514 , \27515 , \27516 , \27517 , \27518 , \27519 , \27520 , \27521 , \27522 ,
         \27523 , \27524 , \27525 , \27526 , \27527 , \27528 , \27529 , \27530 , \27531 , \27532 ,
         \27533 , \27534 , \27535 , \27536 , \27537 , \27538 , \27539 , \27540 , \27541 , \27542 ,
         \27543 , \27544 , \27545 , \27546 , \27547 , \27548 , \27549 , \27550 , \27551 , \27552 ,
         \27553 , \27554 , \27555 , \27556 , \27557 , \27558 , \27559 , \27560 , \27561 , \27562 ,
         \27563 , \27564 , \27565 , \27566 , \27567 , \27568 , \27569 , \27570 , \27571 , \27572 ,
         \27573 , \27574 , \27575 , \27576 , \27577 , \27578 , \27579 , \27580 , \27581 , \27582 ,
         \27583 , \27584 , \27585 , \27586 , \27587 , \27588 , \27589 , \27590 , \27591 , \27592 ,
         \27593 , \27594 , \27595 , \27596 , \27597 , \27598 , \27599 , \27600 , \27601 , \27602 ,
         \27603 , \27604 , \27605 , \27606 , \27607 , \27608 , \27609 , \27610 , \27611 , \27612 ,
         \27613 , \27614 , \27615 , \27616 , \27617 , \27618 , \27619 , \27620 , \27621 , \27622 ,
         \27623 , \27624 , \27625 , \27626 , \27627 , \27628 , \27629 , \27630 , \27631 , \27632 ,
         \27633 , \27634 , \27635 , \27636 , \27637 , \27638 , \27639 , \27640 , \27641 , \27642 ,
         \27643 , \27644 , \27645 , \27646 , \27647 , \27648 , \27649 , \27650 , \27651 , \27652 ,
         \27653 , \27654 , \27655 , \27656 , \27657 , \27658 , \27659 , \27660 , \27661 , \27662 ,
         \27663 , \27664 , \27665 , \27666 , \27667 , \27668 , \27669 , \27670 , \27671 , \27672 ,
         \27673 , \27674 , \27675 , \27676 , \27677 , \27678 , \27679 , \27680 , \27681 , \27682 ,
         \27683 , \27684 , \27685 , \27686 , \27687 , \27688 , \27689 , \27690 , \27691 , \27692 ,
         \27693 , \27694 , \27695 , \27696 , \27697 , \27698 , \27699 , \27700 , \27701 , \27702 ,
         \27703 , \27704 , \27705 , \27706 , \27707 , \27708 , \27709 , \27710 , \27711 , \27712 ,
         \27713 , \27714 , \27715 , \27716 , \27717 , \27718 , \27719 , \27720 , \27721 , \27722 ,
         \27723 , \27724 , \27725 , \27726 , \27727 , \27728 , \27729 , \27730 , \27731 , \27732 ,
         \27733 , \27734 , \27735 , \27736 , \27737 , \27738 , \27739 , \27740 , \27741 , \27742 ,
         \27743 , \27744 , \27745 , \27746 , \27747 , \27748 , \27749 , \27750 , \27751 , \27752 ,
         \27753 , \27754 , \27755 , \27756 , \27757 , \27758 , \27759 , \27760 , \27761 , \27762 ,
         \27763 , \27764 , \27765 , \27766 , \27767 , \27768 , \27769 , \27770 , \27771 , \27772 ,
         \27773 , \27774 , \27775 , \27776 , \27777 , \27778 , \27779 , \27780 , \27781 , \27782 ,
         \27783 , \27784 , \27785 , \27786 , \27787 , \27788 , \27789 , \27790 , \27791 , \27792 ,
         \27793 , \27794 , \27795 , \27796 , \27797 , \27798 , \27799 , \27800 , \27801 , \27802 ,
         \27803 , \27804 , \27805 , \27806 , \27807 , \27808 , \27809 , \27810 , \27811 , \27812 ,
         \27813 , \27814 , \27815 , \27816 , \27817 , \27818 , \27819 , \27820 , \27821 , \27822 ,
         \27823 , \27824 , \27825 , \27826 , \27827 , \27828 , \27829 , \27830 , \27831 , \27832 ,
         \27833 , \27834 , \27835 , \27836 , \27837 , \27838 , \27839 , \27840 , \27841 , \27842 ,
         \27843 , \27844 , \27845 , \27846 , \27847 , \27848 , \27849 , \27850 , \27851 , \27852 ,
         \27853 , \27854 , \27855 , \27856 , \27857 , \27858 , \27859 , \27860 , \27861 , \27862 ,
         \27863 , \27864 , \27865 , \27866 , \27867 , \27868 , \27869 , \27870 , \27871 , \27872 ,
         \27873 , \27874 , \27875 , \27876 , \27877 , \27878 , \27879 , \27880 , \27881 , \27882 ,
         \27883 , \27884 , \27885 , \27886 , \27887 , \27888 , \27889 , \27890 , \27891 , \27892 ,
         \27893 , \27894 , \27895 , \27896 , \27897 , \27898 , \27899 , \27900 , \27901 , \27902 ,
         \27903 , \27904 , \27905 , \27906 , \27907 , \27908 , \27909 , \27910 , \27911 , \27912 ,
         \27913 , \27914 , \27915 , \27916 , \27917 , \27918 , \27919 , \27920 , \27921 , \27922 ,
         \27923 , \27924 , \27925 , \27926 , \27927 , \27928 , \27929 , \27930 , \27931 , \27932 ,
         \27933 , \27934 , \27935 , \27936 , \27937 , \27938 , \27939 , \27940 , \27941 , \27942 ,
         \27943 , \27944 , \27945 , \27946 , \27947 , \27948 , \27949 , \27950 , \27951 , \27952 ,
         \27953 , \27954 , \27955 , \27956 , \27957 , \27958 , \27959 , \27960 , \27961 , \27962 ,
         \27963 , \27964 , \27965 , \27966 , \27967 , \27968 , \27969 , \27970 , \27971 , \27972 ,
         \27973 , \27974 , \27975 , \27976 , \27977 , \27978 , \27979 , \27980 , \27981 , \27982 ,
         \27983 , \27984 , \27985 , \27986 , \27987 , \27988 , \27989 , \27990 , \27991 , \27992 ,
         \27993 , \27994 , \27995 , \27996 , \27997 , \27998 , \27999 , \28000 , \28001 , \28002 ,
         \28003 , \28004 , \28005 , \28006 , \28007 , \28008 , \28009 , \28010 , \28011 , \28012 ,
         \28013 , \28014 , \28015 , \28016 , \28017 , \28018 , \28019 , \28020 , \28021 , \28022 ,
         \28023 , \28024 , \28025 , \28026 , \28027 , \28028 , \28029 , \28030 , \28031 , \28032 ,
         \28033 , \28034 , \28035 , \28036 , \28037 , \28038 , \28039 , \28040 , \28041 , \28042 ,
         \28043 , \28044 , \28045 , \28046 , \28047 , \28048 , \28049 , \28050 , \28051 , \28052 ,
         \28053 , \28054 , \28055 , \28056 , \28057 , \28058 , \28059 , \28060 , \28061 , \28062 ,
         \28063 , \28064 , \28065 , \28066 , \28067 , \28068 , \28069 , \28070 , \28071 , \28072 ,
         \28073 , \28074 , \28075 , \28076 , \28077 , \28078 , \28079 , \28080 , \28081 , \28082 ,
         \28083 , \28084 , \28085 , \28086 , \28087 , \28088 , \28089 , \28090 , \28091 , \28092 ,
         \28093 , \28094 , \28095 , \28096 , \28097 , \28098 , \28099 , \28100 , \28101 , \28102 ,
         \28103 , \28104 , \28105 , \28106 , \28107 , \28108 , \28109 , \28110 , \28111 , \28112 ,
         \28113 , \28114 , \28115 , \28116 , \28117 , \28118 , \28119 , \28120 , \28121 , \28122 ,
         \28123 , \28124 , \28125 , \28126 , \28127 , \28128 , \28129 , \28130 , \28131 , \28132 ,
         \28133 , \28134 , \28135 , \28136 , \28137 , \28138 , \28139 , \28140 , \28141 , \28142 ,
         \28143 , \28144 , \28145 , \28146 , \28147 , \28148 , \28149 , \28150 , \28151 , \28152 ,
         \28153 , \28154 , \28155 , \28156 , \28157 , \28158 , \28159 , \28160 , \28161 , \28162 ,
         \28163 , \28164 , \28165 , \28166 , \28167 , \28168 , \28169 , \28170 , \28171 , \28172 ,
         \28173 , \28174 , \28175 , \28176 , \28177 , \28178 , \28179 , \28180 , \28181 , \28182 ,
         \28183 , \28184 , \28185 , \28186 , \28187 , \28188 , \28189 , \28190 , \28191 , \28192 ,
         \28193 , \28194 , \28195 , \28196 , \28197 , \28198 , \28199 , \28200 , \28201 , \28202 ,
         \28203 , \28204 , \28205 , \28206 , \28207 , \28208 , \28209 , \28210 , \28211 , \28212 ,
         \28213 , \28214 , \28215 , \28216 , \28217 , \28218 , \28219 , \28220 , \28221 , \28222 ,
         \28223 , \28224 , \28225 , \28226 , \28227 , \28228 , \28229 , \28230 , \28231 , \28232 ,
         \28233 , \28234 , \28235 , \28236 , \28237 , \28238 , \28239 , \28240 , \28241 , \28242 ,
         \28243 , \28244 , \28245 , \28246 , \28247 , \28248 , \28249 , \28250 , \28251 , \28252 ,
         \28253 , \28254 , \28255 , \28256 , \28257 , \28258 , \28259 , \28260 , \28261 , \28262 ,
         \28263 , \28264 , \28265 , \28266 , \28267 , \28268 , \28269 , \28270 , \28271 , \28272 ,
         \28273 , \28274 , \28275 , \28276 , \28277 , \28278 , \28279 , \28280 , \28281 , \28282 ,
         \28283 , \28284 , \28285 , \28286 , \28287 , \28288 , \28289 , \28290 , \28291 , \28292 ,
         \28293 , \28294 , \28295 , \28296 , \28297 , \28298 , \28299 , \28300 , \28301 , \28302 ,
         \28303 , \28304 , \28305 , \28306 , \28307 , \28308 , \28309 , \28310 , \28311 , \28312 ,
         \28313 , \28314 , \28315 , \28316 , \28317 , \28318 , \28319 , \28320 , \28321 , \28322 ,
         \28323 , \28324 , \28325 , \28326 , \28327 , \28328 , \28329 , \28330 , \28331 , \28332 ,
         \28333 , \28334 , \28335 , \28336 , \28337 , \28338 , \28339 , \28340 , \28341 , \28342 ,
         \28343 , \28344 , \28345 , \28346 , \28347 , \28348 , \28349 , \28350 , \28351 , \28352 ,
         \28353 , \28354 , \28355 , \28356 , \28357 , \28358 , \28359 , \28360 , \28361 , \28362 ,
         \28363 , \28364 , \28365 , \28366 , \28367 , \28368 , \28369 , \28370 , \28371 , \28372 ,
         \28373 , \28374 , \28375 , \28376 , \28377 , \28378 , \28379 , \28380 , \28381 , \28382 ,
         \28383 , \28384 , \28385 , \28386 , \28387 , \28388 , \28389 , \28390 , \28391 , \28392 ,
         \28393 , \28394 , \28395 , \28396 , \28397 , \28398 , \28399 , \28400 , \28401 , \28402 ,
         \28403 , \28404 , \28405 , \28406 , \28407 , \28408 , \28409 , \28410 , \28411 , \28412 ,
         \28413 , \28414 , \28415 , \28416 , \28417 , \28418 , \28419 , \28420 , \28421 , \28422 ,
         \28423 , \28424 , \28425 , \28426 , \28427 , \28428 , \28429 , \28430 , \28431 , \28432 ,
         \28433 , \28434 , \28435 , \28436 , \28437 , \28438 , \28439 , \28440 , \28441 , \28442 ,
         \28443 , \28444 , \28445 , \28446 , \28447 , \28448 , \28449 , \28450 , \28451 , \28452 ,
         \28453 , \28454 , \28455 , \28456 , \28457 , \28458 , \28459 , \28460 , \28461 , \28462 ,
         \28463 , \28464 , \28465 , \28466 , \28467 , \28468 , \28469 , \28470 , \28471 , \28472 ,
         \28473 , \28474 , \28475 , \28476 , \28477 , \28478 , \28479 , \28480 , \28481 , \28482 ,
         \28483 , \28484 , \28485 , \28486 , \28487 , \28488 , \28489 , \28490 , \28491 , \28492 ,
         \28493 , \28494 , \28495 , \28496 , \28497 , \28498 , \28499 , \28500 , \28501 , \28502 ,
         \28503 , \28504 , \28505 , \28506 , \28507 , \28508 , \28509 , \28510 , \28511 , \28512 ,
         \28513 , \28514 , \28515 , \28516 , \28517 , \28518 , \28519 , \28520 , \28521 , \28522 ,
         \28523 , \28524 , \28525 , \28526 , \28527 , \28528 , \28529 , \28530 , \28531 , \28532 ,
         \28533 , \28534 , \28535 , \28536 , \28537 , \28538 , \28539 , \28540 , \28541 , \28542 ,
         \28543 , \28544 , \28545 , \28546 , \28547 , \28548 , \28549 , \28550 , \28551 , \28552 ,
         \28553 , \28554 , \28555 , \28556 , \28557 , \28558 , \28559 , \28560 , \28561 , \28562 ,
         \28563 , \28564 , \28565 , \28566 , \28567 , \28568 , \28569 , \28570 , \28571 , \28572 ,
         \28573 , \28574 , \28575 , \28576 , \28577 , \28578 , \28579 , \28580 , \28581 , \28582 ,
         \28583 , \28584 , \28585 , \28586 , \28587 , \28588 , \28589 , \28590 , \28591 , \28592 ,
         \28593 , \28594 , \28595 , \28596 , \28597 , \28598 , \28599 , \28600 , \28601 , \28602 ,
         \28603 , \28604 , \28605 , \28606 , \28607 , \28608 , \28609 , \28610 , \28611 , \28612 ,
         \28613 , \28614 , \28615 , \28616 , \28617 , \28618 , \28619 , \28620 , \28621 , \28622 ,
         \28623 , \28624 , \28625 , \28626 , \28627 , \28628 , \28629 , \28630 , \28631 , \28632 ,
         \28633 , \28634 , \28635 , \28636 , \28637 , \28638 , \28639 , \28640 , \28641 , \28642 ,
         \28643 , \28644 , \28645 , \28646 , \28647 , \28648 , \28649 , \28650 , \28651 , \28652 ,
         \28653 , \28654 , \28655 , \28656 , \28657 , \28658 , \28659 , \28660 , \28661 , \28662 ,
         \28663 , \28664 , \28665 , \28666 , \28667 , \28668 , \28669 , \28670 , \28671 , \28672 ,
         \28673 , \28674 , \28675 , \28676 , \28677 , \28678 , \28679 , \28680 , \28681 , \28682 ,
         \28683 , \28684 , \28685 , \28686 , \28687 , \28688 , \28689 , \28690 , \28691 , \28692 ,
         \28693 , \28694 , \28695 , \28696 , \28697 , \28698 , \28699 , \28700 , \28701 , \28702 ,
         \28703 , \28704 , \28705 , \28706 , \28707 , \28708 , \28709 , \28710 , \28711 , \28712 ,
         \28713 , \28714 , \28715 , \28716 , \28717 , \28718 , \28719 , \28720 , \28721 , \28722 ,
         \28723 , \28724 , \28725 , \28726 , \28727 , \28728 , \28729 , \28730 , \28731 , \28732 ,
         \28733 , \28734 , \28735 , \28736 , \28737 , \28738 , \28739 , \28740 , \28741 , \28742 ,
         \28743 , \28744 , \28745 , \28746 , \28747 , \28748 , \28749 , \28750 , \28751 , \28752 ,
         \28753 , \28754 , \28755 , \28756 , \28757 , \28758 , \28759 , \28760 , \28761 , \28762 ,
         \28763 , \28764 , \28765 , \28766 , \28767 , \28768 , \28769 , \28770 , \28771 , \28772 ,
         \28773 , \28774 , \28775 , \28776 , \28777 , \28778 , \28779 , \28780 , \28781 , \28782 ,
         \28783 , \28784 , \28785 , \28786 , \28787 , \28788 , \28789 , \28790 , \28791 , \28792 ,
         \28793 , \28794 , \28795 , \28796 , \28797 , \28798 , \28799 , \28800 , \28801 , \28802 ,
         \28803 , \28804 , \28805 , \28806 , \28807 , \28808 , \28809 , \28810 , \28811 , \28812 ,
         \28813 , \28814 , \28815 , \28816 , \28817 , \28818 , \28819 , \28820 , \28821 , \28822 ,
         \28823 , \28824 , \28825 , \28826 , \28827 , \28828 , \28829 , \28830 , \28831 , \28832 ,
         \28833 , \28834 , \28835 , \28836 , \28837 , \28838 , \28839 , \28840 , \28841 , \28842 ,
         \28843 , \28844 , \28845 , \28846 , \28847 , \28848 , \28849 , \28850 , \28851 , \28852 ,
         \28853 , \28854 , \28855 , \28856 , \28857 , \28858 , \28859 , \28860 , \28861 , \28862 ,
         \28863 , \28864 , \28865 , \28866 , \28867 , \28868 , \28869 , \28870 , \28871 , \28872 ,
         \28873 , \28874 , \28875 , \28876 , \28877 , \28878 , \28879 , \28880 , \28881 , \28882 ,
         \28883 , \28884 , \28885 , \28886 , \28887 , \28888 , \28889 , \28890 , \28891 , \28892 ,
         \28893 , \28894 , \28895 , \28896 , \28897 , \28898 , \28899 , \28900 , \28901 , \28902 ,
         \28903 , \28904 , \28905 , \28906 , \28907 , \28908 , \28909 , \28910 , \28911 , \28912 ,
         \28913 , \28914 , \28915 , \28916 , \28917 , \28918 , \28919 , \28920 , \28921 , \28922 ,
         \28923 , \28924 , \28925 , \28926 , \28927 , \28928 , \28929 , \28930 , \28931 , \28932 ,
         \28933 , \28934 , \28935 , \28936 , \28937 , \28938 , \28939 , \28940 , \28941 , \28942 ,
         \28943 , \28944 , \28945 , \28946 , \28947 , \28948 , \28949 , \28950 , \28951 , \28952 ,
         \28953 , \28954 , \28955 , \28956 , \28957 , \28958 , \28959 , \28960 , \28961 , \28962 ,
         \28963 , \28964 , \28965 , \28966 , \28967 , \28968 , \28969 , \28970 , \28971 , \28972 ,
         \28973 , \28974 , \28975 , \28976 , \28977 , \28978 , \28979 , \28980 , \28981 , \28982 ,
         \28983 , \28984 , \28985 , \28986 , \28987 , \28988 , \28989 , \28990 , \28991 , \28992 ,
         \28993 , \28994 , \28995 , \28996 , \28997 , \28998 , \28999 , \29000 , \29001 , \29002 ,
         \29003 , \29004 , \29005 , \29006 , \29007 , \29008 , \29009 , \29010 , \29011 , \29012 ,
         \29013 , \29014 , \29015 , \29016 , \29017 , \29018 , \29019 , \29020 , \29021 , \29022 ,
         \29023 , \29024 , \29025 , \29026 , \29027 , \29028 , \29029 , \29030 , \29031 , \29032 ,
         \29033 , \29034 , \29035 , \29036 , \29037 , \29038 , \29039 , \29040 , \29041 , \29042 ,
         \29043 , \29044 , \29045 , \29046 , \29047 , \29048 , \29049 , \29050 , \29051 , \29052 ,
         \29053 , \29054 , \29055 , \29056 , \29057 , \29058 , \29059 , \29060 , \29061 , \29062 ,
         \29063 , \29064 , \29065 , \29066 , \29067 , \29068 , \29069 , \29070 , \29071 , \29072 ,
         \29073 , \29074 , \29075 , \29076 , \29077 , \29078 , \29079 , \29080 , \29081 , \29082 ,
         \29083 , \29084 , \29085 , \29086 , \29087 , \29088 , \29089 , \29090 , \29091 , \29092 ,
         \29093 , \29094 , \29095 , \29096 , \29097 , \29098 , \29099 , \29100 , \29101 , \29102 ,
         \29103 , \29104 , \29105 , \29106 , \29107 , \29108 , \29109 , \29110 , \29111 , \29112 ,
         \29113 , \29114 , \29115 , \29116 , \29117 , \29118 , \29119 , \29120 , \29121 , \29122 ,
         \29123 , \29124 , \29125 , \29126 , \29127 , \29128 , \29129 , \29130 , \29131 , \29132 ,
         \29133 , \29134 , \29135 , \29136 , \29137 , \29138 , \29139 , \29140 , \29141 , \29142 ,
         \29143 , \29144 , \29145 , \29146 , \29147 , \29148 , \29149 , \29150 , \29151 , \29152 ,
         \29153 , \29154 , \29155 , \29156 , \29157 , \29158 , \29159 , \29160 , \29161 , \29162 ,
         \29163 , \29164 , \29165 , \29166 , \29167 , \29168 , \29169 , \29170 , \29171 , \29172 ,
         \29173 , \29174 , \29175 , \29176 , \29177 , \29178 , \29179 , \29180 , \29181 , \29182 ,
         \29183 , \29184 , \29185 , \29186 , \29187 , \29188 , \29189 , \29190 , \29191 , \29192 ,
         \29193 , \29194 , \29195 , \29196 , \29197 , \29198 , \29199 , \29200 , \29201 , \29202 ,
         \29203 , \29204 , \29205 , \29206 , \29207 , \29208 , \29209 , \29210 , \29211 , \29212 ,
         \29213 , \29214 , \29215 , \29216 , \29217 , \29218 , \29219 , \29220 , \29221 , \29222 ,
         \29223 , \29224 , \29225 , \29226 , \29227 , \29228 , \29229 , \29230 , \29231 , \29232 ,
         \29233 , \29234 , \29235 , \29236 , \29237 , \29238 , \29239 , \29240 , \29241 , \29242 ,
         \29243 , \29244 , \29245 , \29246 , \29247 , \29248 , \29249 , \29250 , \29251 , \29252 ,
         \29253 , \29254 , \29255 , \29256 , \29257 , \29258 , \29259 , \29260 , \29261 , \29262 ,
         \29263 , \29264 , \29265 , \29266 , \29267 , \29268 , \29269 , \29270 , \29271 , \29272 ,
         \29273 , \29274 , \29275 , \29276 , \29277 , \29278 , \29279 , \29280 , \29281 , \29282 ,
         \29283 , \29284 , \29285 , \29286 , \29287 , \29288 , \29289 , \29290 , \29291 , \29292 ,
         \29293 , \29294 , \29295 , \29296 , \29297 , \29298 , \29299 , \29300 , \29301 , \29302 ,
         \29303 , \29304 , \29305 , \29306 , \29307 , \29308 , \29309 , \29310 , \29311 , \29312 ,
         \29313 , \29314 , \29315 , \29316 , \29317 , \29318 , \29319 , \29320 , \29321 , \29322 ,
         \29323 , \29324 , \29325 , \29326 , \29327 , \29328 , \29329 , \29330 , \29331 , \29332 ,
         \29333 , \29334 , \29335 , \29336 , \29337 , \29338 , \29339 , \29340 , \29341 , \29342 ,
         \29343 , \29344 , \29345 , \29346 , \29347 , \29348 , \29349 , \29350 , \29351 , \29352 ,
         \29353 , \29354 , \29355 , \29356 , \29357 , \29358 , \29359 , \29360 , \29361 , \29362 ,
         \29363 , \29364 , \29365 , \29366 , \29367 , \29368 , \29369 , \29370 , \29371 , \29372 ,
         \29373 , \29374 , \29375 , \29376 , \29377 , \29378 , \29379 , \29380 , \29381 , \29382 ,
         \29383 , \29384 , \29385 , \29386 , \29387 , \29388 , \29389 , \29390 , \29391 , \29392 ,
         \29393 , \29394 , \29395 , \29396 , \29397 , \29398 , \29399 , \29400 , \29401 , \29402 ,
         \29403 , \29404 , \29405 , \29406 , \29407 , \29408 , \29409 , \29410 , \29411 , \29412 ,
         \29413 , \29414 , \29415 , \29416 , \29417 , \29418 , \29419 , \29420 , \29421 , \29422 ,
         \29423 , \29424 , \29425 , \29426 , \29427 , \29428 , \29429 , \29430 , \29431 , \29432 ,
         \29433 , \29434 , \29435 , \29436 , \29437 , \29438 , \29439 , \29440 , \29441 , \29442 ,
         \29443 , \29444 , \29445 , \29446 , \29447 , \29448 , \29449 , \29450 , \29451 , \29452 ,
         \29453 , \29454 , \29455 , \29456 , \29457 , \29458 , \29459 , \29460 , \29461 , \29462 ,
         \29463 , \29464 , \29465 , \29466 , \29467 , \29468 , \29469 , \29470 , \29471 , \29472 ,
         \29473 , \29474 , \29475 , \29476 , \29477 , \29478 , \29479 , \29480 , \29481 , \29482 ,
         \29483 , \29484 , \29485 , \29486 , \29487 , \29488 , \29489 , \29490 , \29491 , \29492 ,
         \29493 , \29494 , \29495 , \29496 , \29497 , \29498 , \29499 , \29500 , \29501 , \29502 ,
         \29503 , \29504 , \29505 , \29506 , \29507 , \29508 , \29509 , \29510 , \29511 , \29512 ,
         \29513 , \29514 , \29515 , \29516 , \29517 , \29518 , \29519 , \29520 , \29521 , \29522 ,
         \29523 , \29524 , \29525 , \29526 , \29527 , \29528 , \29529 , \29530 , \29531 , \29532 ,
         \29533 , \29534 , \29535 , \29536 , \29537 , \29538 , \29539 , \29540 , \29541 , \29542 ,
         \29543 , \29544 , \29545 , \29546 , \29547 , \29548 , \29549 , \29550 , \29551 , \29552 ,
         \29553 , \29554 , \29555 , \29556 , \29557 , \29558 , \29559 , \29560 , \29561 , \29562 ,
         \29563 , \29564 , \29565 , \29566 , \29567 , \29568 , \29569 , \29570 , \29571 , \29572 ,
         \29573 , \29574 , \29575 , \29576 , \29577 , \29578 , \29579 , \29580 , \29581 , \29582 ,
         \29583 , \29584 , \29585 , \29586 , \29587 , \29588 , \29589 , \29590 , \29591 , \29592 ,
         \29593 , \29594 , \29595 , \29596 , \29597 , \29598 , \29599 , \29600 , \29601 , \29602 ,
         \29603 , \29604 , \29605 , \29606 , \29607 , \29608 , \29609 , \29610 , \29611 , \29612 ,
         \29613 , \29614 , \29615 , \29616 , \29617 , \29618 , \29619 , \29620 , \29621 , \29622 ,
         \29623 , \29624 , \29625 , \29626 , \29627 , \29628 , \29629 , \29630 , \29631 , \29632 ,
         \29633 , \29634 , \29635 , \29636 , \29637 , \29638 , \29639 , \29640 , \29641 , \29642 ,
         \29643 , \29644 , \29645 , \29646 , \29647 , \29648 , \29649 , \29650 , \29651 , \29652 ,
         \29653 , \29654 , \29655 , \29656 , \29657 , \29658 , \29659 , \29660 , \29661 , \29662 ,
         \29663 , \29664 , \29665 , \29666 , \29667 , \29668 , \29669 , \29670 , \29671 , \29672 ,
         \29673 , \29674 , \29675 , \29676 , \29677 , \29678 , \29679 , \29680 , \29681 , \29682 ,
         \29683 , \29684 , \29685 , \29686 , \29687 , \29688 , \29689 , \29690 , \29691 , \29692 ,
         \29693 , \29694 , \29695 , \29696 , \29697 , \29698 , \29699 , \29700 , \29701 , \29702 ,
         \29703 , \29704 , \29705 , \29706 , \29707 , \29708 , \29709 , \29710 , \29711 , \29712 ,
         \29713 , \29714 , \29715 , \29716 , \29717 , \29718 , \29719 , \29720 , \29721 , \29722 ,
         \29723 , \29724 , \29725 , \29726 , \29727 , \29728 , \29729 , \29730 , \29731 , \29732 ,
         \29733 , \29734 , \29735 , \29736 , \29737 , \29738 , \29739 , \29740 , \29741 , \29742 ,
         \29743 , \29744 , \29745 , \29746 , \29747 , \29748 , \29749 , \29750 , \29751 , \29752 ,
         \29753 , \29754 , \29755 , \29756 , \29757 , \29758 , \29759 , \29760 , \29761 , \29762 ,
         \29763 , \29764 , \29765 , \29766 , \29767 , \29768 , \29769 , \29770 , \29771 , \29772 ,
         \29773 , \29774 , \29775 , \29776 , \29777 , \29778 , \29779 , \29780 , \29781 , \29782 ,
         \29783 , \29784 , \29785 , \29786 , \29787 , \29788 , \29789 , \29790 , \29791 , \29792 ,
         \29793 , \29794 , \29795 , \29796 , \29797 , \29798 , \29799 , \29800 , \29801 , \29802 ,
         \29803 , \29804 , \29805 , \29806 , \29807 , \29808 , \29809 , \29810 , \29811 , \29812 ,
         \29813 , \29814 , \29815 , \29816 , \29817 , \29818 , \29819 , \29820 , \29821 , \29822 ,
         \29823 , \29824 , \29825 , \29826 , \29827 , \29828 , \29829 , \29830 , \29831 , \29832 ,
         \29833 , \29834 , \29835 , \29836 , \29837 , \29838 , \29839 , \29840 , \29841 , \29842 ,
         \29843 , \29844 , \29845 , \29846 , \29847 , \29848 , \29849 , \29850 , \29851 , \29852 ,
         \29853 , \29854 , \29855 , \29856 , \29857 , \29858 , \29859 , \29860 , \29861 , \29862 ,
         \29863 , \29864 , \29865 , \29866 , \29867 , \29868 , \29869 , \29870 , \29871 , \29872 ,
         \29873 , \29874 , \29875 , \29876 , \29877 , \29878 , \29879 , \29880 , \29881 , \29882 ,
         \29883 , \29884 , \29885 , \29886 , \29887 , \29888 , \29889 , \29890 , \29891 , \29892 ,
         \29893 , \29894 , \29895 , \29896 , \29897 , \29898 , \29899 , \29900 , \29901 , \29902 ,
         \29903 , \29904 , \29905 , \29906 , \29907 , \29908 , \29909 , \29910 , \29911 , \29912 ,
         \29913 , \29914 , \29915 , \29916 , \29917 , \29918 , \29919 , \29920 , \29921 , \29922 ,
         \29923 , \29924 , \29925 , \29926 , \29927 , \29928 , \29929 , \29930 , \29931 , \29932 ,
         \29933 , \29934 , \29935 , \29936 , \29937 , \29938 , \29939 , \29940 , \29941 , \29942 ,
         \29943 , \29944 , \29945 , \29946 , \29947 , \29948 , \29949 , \29950 , \29951 , \29952 ,
         \29953 , \29954 , \29955 , \29956 , \29957 , \29958 , \29959 , \29960 , \29961 , \29962 ,
         \29963 , \29964 , \29965 , \29966 , \29967 , \29968 , \29969 , \29970 , \29971 , \29972 ,
         \29973 , \29974 , \29975 , \29976 , \29977 , \29978 , \29979 , \29980 , \29981 , \29982 ,
         \29983 , \29984 , \29985 , \29986 , \29987 , \29988 , \29989 , \29990 , \29991 , \29992 ,
         \29993 , \29994 , \29995 , \29996 , \29997 , \29998 , \29999 , \30000 , \30001 , \30002 ,
         \30003 , \30004 , \30005 , \30006 , \30007 , \30008 , \30009 , \30010 , \30011 , \30012 ,
         \30013 , \30014 , \30015 , \30016 , \30017 , \30018 , \30019 , \30020 , \30021 , \30022 ,
         \30023 , \30024 , \30025 , \30026 , \30027 , \30028 , \30029 , \30030 , \30031 , \30032 ,
         \30033 , \30034 , \30035 , \30036 , \30037 , \30038 , \30039 , \30040 , \30041 , \30042 ,
         \30043 , \30044 , \30045 , \30046 , \30047 , \30048 , \30049 , \30050 , \30051 , \30052 ,
         \30053 , \30054 , \30055 , \30056 , \30057 , \30058 , \30059 , \30060 , \30061 , \30062 ,
         \30063 , \30064 , \30065 , \30066 , \30067 , \30068 , \30069 , \30070 , \30071 , \30072 ,
         \30073 , \30074 , \30075 , \30076 , \30077 , \30078 , \30079 , \30080 , \30081 , \30082 ,
         \30083 , \30084 , \30085 , \30086 , \30087 , \30088 , \30089 , \30090 , \30091 , \30092 ,
         \30093 , \30094 , \30095 , \30096 , \30097 , \30098 , \30099 , \30100 , \30101 , \30102 ,
         \30103 , \30104 , \30105 , \30106 , \30107 , \30108 , \30109 , \30110 , \30111 , \30112 ,
         \30113 , \30114 , \30115 , \30116 , \30117 , \30118 , \30119 , \30120 , \30121 , \30122 ,
         \30123 , \30124 , \30125 , \30126 , \30127 , \30128 , \30129 , \30130 , \30131 , \30132 ,
         \30133 , \30134 , \30135 , \30136 , \30137 , \30138 , \30139 , \30140 , \30141 , \30142 ,
         \30143 , \30144 , \30145 , \30146 , \30147 , \30148 , \30149 , \30150 , \30151 , \30152 ,
         \30153 , \30154 , \30155 , \30156 , \30157 , \30158 , \30159 , \30160 , \30161 , \30162 ,
         \30163 , \30164 , \30165 , \30166 , \30167 , \30168 , \30169 , \30170 , \30171 , \30172 ,
         \30173 , \30174 , \30175 , \30176 , \30177 , \30178 , \30179 , \30180 , \30181 , \30182 ,
         \30183 , \30184 , \30185 , \30186 , \30187 , \30188 , \30189 , \30190 , \30191 , \30192 ,
         \30193 , \30194 , \30195 , \30196 , \30197 , \30198 , \30199 , \30200 , \30201 , \30202 ,
         \30203 , \30204 , \30205 , \30206 , \30207 , \30208 , \30209 , \30210 , \30211 , \30212 ,
         \30213 , \30214 , \30215 , \30216 , \30217 , \30218 , \30219 , \30220 , \30221 , \30222 ,
         \30223 , \30224 , \30225 , \30226 , \30227 , \30228 , \30229 , \30230 , \30231 , \30232 ,
         \30233 , \30234 , \30235 , \30236 , \30237 , \30238 , \30239 , \30240 , \30241 , \30242 ,
         \30243 , \30244 , \30245 , \30246 , \30247 , \30248 , \30249 , \30250 , \30251 , \30252 ,
         \30253 , \30254 , \30255 , \30256 , \30257 , \30258 , \30259 , \30260 , \30261 , \30262 ,
         \30263 , \30264 , \30265 , \30266 , \30267 , \30268 , \30269 , \30270 , \30271 , \30272 ,
         \30273 , \30274 , \30275 , \30276 , \30277 , \30278 , \30279 , \30280 , \30281 , \30282 ,
         \30283 , \30284 , \30285 , \30286 , \30287 , \30288 , \30289 , \30290 , \30291 , \30292 ,
         \30293 , \30294 , \30295 , \30296 , \30297 , \30298 , \30299 , \30300 , \30301 , \30302 ,
         \30303 , \30304 , \30305 , \30306 , \30307 , \30308 , \30309 , \30310 , \30311 , \30312 ,
         \30313 , \30314 , \30315 , \30316 , \30317 , \30318 , \30319 , \30320 , \30321 , \30322 ,
         \30323 , \30324 , \30325 , \30326 , \30327 , \30328 , \30329 , \30330 , \30331 , \30332 ,
         \30333 , \30334 , \30335 , \30336 , \30337 , \30338 , \30339 , \30340 , \30341 , \30342 ,
         \30343 , \30344 , \30345 , \30346 , \30347 , \30348 , \30349 , \30350 , \30351 , \30352 ,
         \30353 , \30354 , \30355 , \30356 , \30357 , \30358 , \30359 , \30360 , \30361 , \30362 ,
         \30363 , \30364 , \30365 , \30366 , \30367 , \30368 , \30369 , \30370 , \30371 , \30372 ,
         \30373 , \30374 , \30375 , \30376 , \30377 , \30378 , \30379 , \30380 , \30381 , \30382 ,
         \30383 , \30384 , \30385 , \30386 , \30387 , \30388 , \30389 , \30390 , \30391 , \30392 ,
         \30393 , \30394 , \30395 , \30396 , \30397 , \30398 , \30399 , \30400 , \30401 , \30402 ,
         \30403 , \30404 , \30405 , \30406 , \30407 , \30408 , \30409 , \30410 , \30411 , \30412 ,
         \30413 , \30414 , \30415 , \30416 , \30417 , \30418 , \30419 , \30420 , \30421 , \30422 ,
         \30423 , \30424 , \30425 , \30426 , \30427 , \30428 , \30429 , \30430 , \30431 , \30432 ,
         \30433 , \30434 , \30435 , \30436 , \30437 , \30438 , \30439 , \30440 , \30441 , \30442 ,
         \30443 , \30444 , \30445 , \30446 , \30447 , \30448 , \30449 , \30450 , \30451 , \30452 ,
         \30453 , \30454 , \30455 , \30456 , \30457 , \30458 , \30459 , \30460 , \30461 , \30462 ,
         \30463 , \30464 , \30465 , \30466 , \30467 , \30468 , \30469 , \30470 , \30471 , \30472 ,
         \30473 , \30474 , \30475 , \30476 , \30477 , \30478 , \30479 , \30480 , \30481 , \30482 ,
         \30483 , \30484 , \30485 , \30486 , \30487 , \30488 , \30489 , \30490 , \30491 , \30492 ,
         \30493 , \30494 , \30495 , \30496 , \30497 , \30498 , \30499 , \30500 , \30501 , \30502 ,
         \30503 , \30504 , \30505 , \30506 , \30507 , \30508 , \30509 , \30510 , \30511 , \30512 ,
         \30513 , \30514 , \30515 , \30516 , \30517 , \30518 , \30519 , \30520 , \30521 , \30522 ,
         \30523 , \30524 , \30525 , \30526 , \30527 , \30528 , \30529 , \30530 , \30531 , \30532 ,
         \30533 , \30534 , \30535 , \30536 , \30537 , \30538 , \30539 , \30540 , \30541 , \30542 ,
         \30543 , \30544 , \30545 , \30546 , \30547 , \30548 , \30549 , \30550 , \30551 , \30552 ,
         \30553 , \30554 , \30555 , \30556 , \30557 , \30558 , \30559 , \30560 , \30561 , \30562 ,
         \30563 , \30564 , \30565 , \30566 , \30567 , \30568 , \30569 , \30570 , \30571 , \30572 ,
         \30573 , \30574 , \30575 , \30576 , \30577 , \30578 , \30579 , \30580 , \30581 , \30582 ,
         \30583 , \30584 , \30585 , \30586 , \30587 , \30588 , \30589 , \30590 , \30591 , \30592 ,
         \30593 , \30594 , \30595 , \30596 , \30597 , \30598 , \30599 , \30600 , \30601 , \30602 ,
         \30603 , \30604 , \30605 , \30606 , \30607 , \30608 , \30609 , \30610 , \30611 , \30612 ,
         \30613 , \30614 , \30615 , \30616 , \30617 , \30618 , \30619 , \30620 , \30621 , \30622 ,
         \30623 , \30624 , \30625 , \30626 , \30627 , \30628 , \30629 , \30630 , \30631 , \30632 ,
         \30633 , \30634 , \30635 , \30636 , \30637 , \30638 , \30639 , \30640 , \30641 , \30642 ,
         \30643 , \30644 , \30645 , \30646 , \30647 , \30648 , \30649 , \30650 , \30651 , \30652 ,
         \30653 , \30654 , \30655 , \30656 , \30657 , \30658 , \30659 , \30660 , \30661 , \30662 ,
         \30663 , \30664 , \30665 , \30666 , \30667 , \30668 , \30669 , \30670 , \30671 , \30672 ,
         \30673 , \30674 , \30675 , \30676 , \30677 , \30678 , \30679 , \30680 , \30681 , \30682 ,
         \30683 , \30684 , \30685 , \30686 , \30687 , \30688 , \30689 , \30690 , \30691 , \30692 ,
         \30693 , \30694 , \30695 , \30696 , \30697 , \30698 , \30699 , \30700 , \30701 , \30702 ,
         \30703 , \30704 , \30705 , \30706 , \30707 , \30708 , \30709 , \30710 , \30711 , \30712 ,
         \30713 , \30714 , \30715 , \30716 , \30717 , \30718 , \30719 , \30720 , \30721 , \30722 ,
         \30723 , \30724 , \30725 , \30726 , \30727 , \30728 , \30729 , \30730 , \30731 , \30732 ,
         \30733 , \30734 , \30735 , \30736 , \30737 , \30738 , \30739 , \30740 , \30741 , \30742 ,
         \30743 , \30744 , \30745 , \30746 , \30747 , \30748 , \30749 , \30750 , \30751 , \30752 ,
         \30753 , \30754 , \30755 , \30756 , \30757 , \30758 , \30759 , \30760 , \30761 , \30762 ,
         \30763 , \30764 , \30765 , \30766 , \30767 , \30768 , \30769 , \30770 , \30771 , \30772 ,
         \30773 , \30774 , \30775 , \30776 , \30777 , \30778 , \30779 , \30780 , \30781 , \30782 ,
         \30783 , \30784 , \30785 , \30786 , \30787 , \30788 , \30789 , \30790 , \30791 , \30792 ,
         \30793 , \30794 , \30795 , \30796 , \30797 , \30798 , \30799 , \30800 , \30801 , \30802 ,
         \30803 , \30804 , \30805 , \30806 , \30807 , \30808 , \30809 , \30810 , \30811 , \30812 ,
         \30813 , \30814 , \30815 , \30816 , \30817 , \30818 , \30819 , \30820 , \30821 , \30822 ,
         \30823 , \30824 , \30825 , \30826 , \30827 , \30828 , \30829 , \30830 , \30831 , \30832 ,
         \30833 , \30834 , \30835 , \30836 , \30837 , \30838 , \30839 , \30840 , \30841 , \30842 ,
         \30843 , \30844 , \30845 , \30846 , \30847 , \30848 , \30849 , \30850 , \30851 , \30852 ,
         \30853 , \30854 , \30855 , \30856 , \30857 , \30858 , \30859 , \30860 , \30861 , \30862 ,
         \30863 , \30864 , \30865 , \30866 , \30867 , \30868 , \30869 , \30870 , \30871 , \30872 ,
         \30873 , \30874 , \30875 , \30876 , \30877 , \30878 , \30879 , \30880 , \30881 , \30882 ,
         \30883 , \30884 , \30885 , \30886 , \30887 , \30888 , \30889 , \30890 , \30891 , \30892 ,
         \30893 , \30894 , \30895 , \30896 , \30897 , \30898 , \30899 , \30900 , \30901 , \30902 ,
         \30903 , \30904 , \30905 , \30906 , \30907 , \30908 , \30909 , \30910 , \30911 , \30912 ,
         \30913 , \30914 , \30915 , \30916 , \30917 , \30918 , \30919 , \30920 , \30921 , \30922 ,
         \30923 , \30924 , \30925 , \30926 , \30927 , \30928 , \30929 , \30930 , \30931 , \30932 ,
         \30933 , \30934 , \30935 , \30936 , \30937 , \30938 , \30939 , \30940 , \30941 , \30942 ,
         \30943 , \30944 , \30945 , \30946 , \30947 , \30948 , \30949 , \30950 , \30951 , \30952 ,
         \30953 , \30954 , \30955 , \30956 , \30957 , \30958 , \30959 , \30960 , \30961 , \30962 ,
         \30963 , \30964 , \30965 , \30966 , \30967 , \30968 , \30969 , \30970 , \30971 , \30972 ,
         \30973 , \30974 , \30975 , \30976 , \30977 , \30978 , \30979 , \30980 , \30981 , \30982 ,
         \30983 , \30984 , \30985 , \30986 , \30987 , \30988 , \30989 , \30990 , \30991 , \30992 ,
         \30993 , \30994 , \30995 , \30996 , \30997 , \30998 , \30999 , \31000 , \31001 , \31002 ,
         \31003 , \31004 , \31005 , \31006 , \31007 , \31008 , \31009 , \31010 , \31011 , \31012 ,
         \31013 , \31014 , \31015 , \31016 , \31017 , \31018 , \31019 , \31020 , \31021 , \31022 ,
         \31023 , \31024 , \31025 , \31026 , \31027 , \31028 , \31029 , \31030 , \31031 , \31032 ,
         \31033 , \31034 , \31035 , \31036 , \31037 , \31038 , \31039 , \31040 , \31041 , \31042 ,
         \31043 , \31044 , \31045 , \31046 , \31047 , \31048 , \31049 , \31050 , \31051 , \31052 ,
         \31053 , \31054 , \31055 , \31056 , \31057 , \31058 , \31059 , \31060 , \31061 , \31062 ,
         \31063 , \31064 , \31065 , \31066 , \31067 , \31068 , \31069 , \31070 , \31071 , \31072 ,
         \31073 , \31074 , \31075 , \31076 , \31077 , \31078 , \31079 , \31080 , \31081 , \31082 ,
         \31083 , \31084 , \31085 , \31086 , \31087 , \31088 , \31089 , \31090 , \31091 , \31092 ,
         \31093 , \31094 , \31095 , \31096 , \31097 , \31098 , \31099 , \31100 , \31101 , \31102 ,
         \31103 , \31104 , \31105 , \31106 , \31107 , \31108 , \31109 , \31110 , \31111 , \31112 ,
         \31113 , \31114 , \31115 , \31116 , \31117 , \31118 , \31119 , \31120 , \31121 , \31122 ,
         \31123 , \31124 , \31125 , \31126 , \31127 , \31128 , \31129 , \31130 , \31131 , \31132 ,
         \31133 , \31134 , \31135 , \31136 , \31137 , \31138 , \31139 , \31140 , \31141 , \31142 ,
         \31143 , \31144 , \31145 , \31146 , \31147 , \31148 , \31149 , \31150 , \31151 , \31152 ,
         \31153 , \31154 , \31155 , \31156 , \31157 , \31158 , \31159 , \31160 , \31161 , \31162 ,
         \31163 , \31164 , \31165 , \31166 , \31167 , \31168 , \31169 , \31170 , \31171 , \31172 ,
         \31173 , \31174 , \31175 , \31176 , \31177 , \31178 , \31179 , \31180 , \31181 , \31182 ,
         \31183 , \31184 , \31185 , \31186 , \31187 , \31188 , \31189 , \31190 , \31191 , \31192 ,
         \31193 , \31194 , \31195 , \31196 , \31197 , \31198 , \31199 , \31200 , \31201 , \31202 ,
         \31203 , \31204 , \31205 , \31206 , \31207 , \31208 , \31209 , \31210 , \31211 , \31212 ,
         \31213 , \31214 , \31215 , \31216 , \31217 , \31218 , \31219 , \31220 , \31221 , \31222 ,
         \31223 , \31224 , \31225 , \31226 , \31227 , \31228 , \31229 , \31230 , \31231 , \31232 ,
         \31233 , \31234 , \31235 , \31236 , \31237 , \31238 , \31239 , \31240 , \31241 , \31242 ,
         \31243 , \31244 , \31245 , \31246 , \31247 , \31248 , \31249 , \31250 , \31251 , \31252 ,
         \31253 , \31254 , \31255 , \31256 , \31257 , \31258 , \31259 , \31260 , \31261 , \31262 ,
         \31263 , \31264 , \31265 , \31266 , \31267 , \31268 , \31269 , \31270 , \31271 , \31272 ,
         \31273 , \31274 , \31275 , \31276 , \31277 , \31278 , \31279 , \31280 , \31281 , \31282 ,
         \31283 , \31284 , \31285 , \31286 , \31287 , \31288 , \31289 , \31290 , \31291 , \31292 ,
         \31293 , \31294 , \31295 , \31296 , \31297 , \31298 , \31299 , \31300 , \31301 , \31302 ,
         \31303 , \31304 , \31305 , \31306 , \31307 , \31308 , \31309 , \31310 , \31311 , \31312 ,
         \31313 , \31314 , \31315 , \31316 , \31317 , \31318 , \31319 , \31320 , \31321 , \31322 ,
         \31323 , \31324 , \31325 , \31326 , \31327 , \31328 , \31329 , \31330 , \31331 , \31332 ,
         \31333 , \31334 , \31335 , \31336 , \31337 , \31338 , \31339 , \31340 , \31341 , \31342 ,
         \31343 , \31344 , \31345 , \31346 , \31347 , \31348 , \31349 , \31350 , \31351 , \31352 ,
         \31353 , \31354 , \31355 , \31356 , \31357 , \31358 , \31359 , \31360 , \31361 , \31362 ,
         \31363 , \31364 , \31365 , \31366 , \31367 , \31368 , \31369 , \31370 , \31371 , \31372 ,
         \31373 , \31374 , \31375 , \31376 , \31377 , \31378 , \31379 , \31380 , \31381 , \31382 ,
         \31383 , \31384 , \31385 , \31386 , \31387 , \31388 , \31389 , \31390 , \31391 , \31392 ,
         \31393 , \31394 , \31395 , \31396 , \31397 , \31398 , \31399 , \31400 , \31401 , \31402 ,
         \31403 , \31404 , \31405 , \31406 , \31407 , \31408 , \31409 , \31410 , \31411 , \31412 ,
         \31413 , \31414 , \31415 , \31416 , \31417 , \31418 , \31419 , \31420 , \31421 , \31422 ,
         \31423 , \31424 , \31425 , \31426 , \31427 , \31428 , \31429 , \31430 , \31431 , \31432 ,
         \31433 , \31434 , \31435 , \31436 , \31437 , \31438 , \31439 , \31440 , \31441 , \31442 ,
         \31443 , \31444 , \31445 , \31446 , \31447 , \31448 , \31449 , \31450 , \31451 , \31452 ,
         \31453 , \31454 , \31455 , \31456 , \31457 , \31458 , \31459 , \31460 , \31461 , \31462 ,
         \31463 , \31464 , \31465 , \31466 , \31467 , \31468 , \31469 , \31470 , \31471 , \31472 ,
         \31473 , \31474 , \31475 , \31476 , \31477 , \31478 , \31479 , \31480 , \31481 , \31482 ,
         \31483 , \31484 , \31485 , \31486 , \31487 , \31488 , \31489 , \31490 , \31491 , \31492 ,
         \31493 , \31494 , \31495 , \31496 , \31497 , \31498 , \31499 , \31500 , \31501 , \31502 ,
         \31503 , \31504 , \31505 , \31506 , \31507 , \31508 , \31509 , \31510 , \31511 , \31512 ,
         \31513 , \31514 , \31515 , \31516 , \31517 , \31518 , \31519 , \31520 , \31521 , \31522 ,
         \31523 , \31524 , \31525 , \31526 , \31527 , \31528 , \31529 , \31530 , \31531 , \31532 ,
         \31533 , \31534 , \31535 , \31536 , \31537 , \31538 , \31539 , \31540 , \31541 , \31542 ,
         \31543 , \31544 , \31545 , \31546 , \31547 , \31548 , \31549 , \31550 , \31551 , \31552 ,
         \31553 , \31554 , \31555 , \31556 , \31557 , \31558 , \31559 , \31560 , \31561 , \31562 ,
         \31563 , \31564 , \31565 , \31566 , \31567 , \31568 , \31569 , \31570 , \31571 , \31572 ,
         \31573 , \31574 , \31575 , \31576 , \31577 , \31578 , \31579 , \31580 , \31581 , \31582 ,
         \31583 , \31584 , \31585 , \31586 , \31587 , \31588 , \31589 , \31590 , \31591 , \31592 ,
         \31593 , \31594 , \31595 , \31596 , \31597 , \31598 , \31599 , \31600 , \31601 , \31602 ,
         \31603 , \31604 , \31605 , \31606 , \31607 , \31608 , \31609 , \31610 , \31611 , \31612 ,
         \31613 , \31614 , \31615 , \31616 , \31617 , \31618 , \31619 , \31620 , \31621 , \31622 ,
         \31623 , \31624 , \31625 , \31626 , \31627 , \31628 , \31629 , \31630 , \31631 , \31632 ,
         \31633 , \31634 , \31635 , \31636 , \31637 , \31638 , \31639 , \31640 , \31641 , \31642 ,
         \31643 , \31644 , \31645 , \31646 , \31647 , \31648 , \31649 , \31650 , \31651 , \31652 ,
         \31653 , \31654 , \31655 , \31656 , \31657 , \31658 , \31659 , \31660 , \31661 , \31662 ,
         \31663 , \31664 , \31665 , \31666 , \31667 , \31668 , \31669 , \31670 , \31671 , \31672 ,
         \31673 , \31674 , \31675 , \31676 , \31677 , \31678 , \31679 , \31680 , \31681 , \31682 ,
         \31683 , \31684 , \31685 , \31686 , \31687 , \31688 , \31689 , \31690 , \31691 , \31692 ,
         \31693 , \31694 , \31695 , \31696 , \31697 , \31698 , \31699 , \31700 , \31701 , \31702 ,
         \31703 , \31704 , \31705 , \31706 , \31707 , \31708 , \31709 , \31710 , \31711 , \31712 ,
         \31713 , \31714 , \31715 , \31716 , \31717 , \31718 , \31719 , \31720 , \31721 , \31722 ,
         \31723 , \31724 , \31725 , \31726 , \31727 , \31728 , \31729 , \31730 , \31731 , \31732 ,
         \31733 , \31734 , \31735 , \31736 , \31737 , \31738 , \31739 , \31740 , \31741 , \31742 ,
         \31743 , \31744 , \31745 , \31746 , \31747 , \31748 , \31749 , \31750 , \31751 , \31752 ,
         \31753 , \31754 , \31755 , \31756 , \31757 , \31758 , \31759 , \31760 , \31761 , \31762 ,
         \31763 , \31764 , \31765 , \31766 , \31767 , \31768 , \31769 , \31770 , \31771 , \31772 ,
         \31773 , \31774 , \31775 , \31776 , \31777 , \31778 , \31779 , \31780 , \31781 , \31782 ,
         \31783 , \31784 , \31785 , \31786 , \31787 , \31788 , \31789 , \31790 , \31791 , \31792 ,
         \31793 , \31794 , \31795 , \31796 , \31797 , \31798 , \31799 , \31800 , \31801 , \31802 ,
         \31803 , \31804 , \31805 , \31806 , \31807 , \31808 , \31809 , \31810 , \31811 , \31812 ,
         \31813 , \31814 , \31815 , \31816 , \31817 , \31818 , \31819 , \31820 , \31821 , \31822 ,
         \31823 , \31824 , \31825 , \31826 , \31827 , \31828 , \31829 , \31830 , \31831 , \31832 ,
         \31833 , \31834 , \31835 , \31836 , \31837 , \31838 , \31839 , \31840 , \31841 , \31842 ,
         \31843 , \31844 , \31845 , \31846 , \31847 , \31848 , \31849 , \31850 , \31851 , \31852 ,
         \31853 , \31854 , \31855 , \31856 , \31857 , \31858 , \31859 , \31860 , \31861 , \31862 ,
         \31863 , \31864 , \31865 , \31866 , \31867 , \31868 , \31869 , \31870 , \31871 , \31872 ,
         \31873 , \31874 , \31875 , \31876 , \31877 , \31878 , \31879 , \31880 , \31881 , \31882 ,
         \31883 , \31884 , \31885 , \31886 , \31887 , \31888 , \31889 , \31890 , \31891 , \31892 ,
         \31893 , \31894 , \31895 , \31896 , \31897 , \31898 , \31899 , \31900 , \31901 , \31902 ,
         \31903 , \31904 , \31905 , \31906 , \31907 , \31908 , \31909 , \31910 , \31911 , \31912 ,
         \31913 , \31914 , \31915 , \31916 , \31917 , \31918 , \31919 , \31920 , \31921 , \31922 ,
         \31923 , \31924 , \31925 , \31926 , \31927 , \31928 , \31929 , \31930 , \31931 , \31932 ,
         \31933 , \31934 , \31935 , \31936 , \31937 , \31938 , \31939 , \31940 , \31941 , \31942 ,
         \31943 , \31944 , \31945 , \31946 , \31947 , \31948 , \31949 , \31950 , \31951 , \31952 ,
         \31953 , \31954 , \31955 , \31956 , \31957 , \31958 , \31959 , \31960 , \31961 , \31962 ,
         \31963 , \31964 , \31965 , \31966 , \31967 , \31968 , \31969 , \31970 , \31971 , \31972 ,
         \31973 , \31974 , \31975 , \31976 , \31977 , \31978 , \31979 , \31980 , \31981 , \31982 ,
         \31983 , \31984 , \31985 , \31986 , \31987 , \31988 , \31989 , \31990 , \31991 , \31992 ,
         \31993 , \31994 , \31995 , \31996 , \31997 , \31998 , \31999 , \32000 , \32001 , \32002 ,
         \32003 , \32004 , \32005 , \32006 , \32007 , \32008 , \32009 , \32010 , \32011 , \32012 ,
         \32013 , \32014 , \32015 , \32016 , \32017 , \32018 , \32019 , \32020 , \32021 , \32022 ,
         \32023 , \32024 , \32025 , \32026 , \32027 , \32028 , \32029 , \32030 , \32031 , \32032 ,
         \32033 , \32034 , \32035 , \32036 , \32037 , \32038 , \32039 , \32040 , \32041 , \32042 ,
         \32043 , \32044 , \32045 , \32046 , \32047 , \32048 , \32049 , \32050 , \32051 , \32052 ,
         \32053 , \32054 , \32055 , \32056 , \32057 , \32058 , \32059 , \32060 , \32061 , \32062 ,
         \32063 , \32064 , \32065 , \32066 , \32067 , \32068 , \32069 , \32070 , \32071 , \32072 ,
         \32073 , \32074 , \32075 , \32076 , \32077 , \32078 , \32079 , \32080 , \32081 , \32082 ,
         \32083 , \32084 , \32085 , \32086 , \32087 , \32088 , \32089 , \32090 , \32091 , \32092 ,
         \32093 , \32094 , \32095 , \32096 , \32097 , \32098 , \32099 , \32100 , \32101 , \32102 ,
         \32103 , \32104 , \32105 , \32106 , \32107 , \32108 , \32109 , \32110 , \32111 , \32112 ,
         \32113 , \32114 , \32115 , \32116 , \32117 , \32118 , \32119 , \32120 , \32121 , \32122 ,
         \32123 , \32124 , \32125 , \32126 , \32127 , \32128 , \32129 , \32130 , \32131 , \32132 ,
         \32133 , \32134 , \32135 , \32136 , \32137 , \32138 , \32139 , \32140 , \32141 , \32142 ,
         \32143 , \32144 , \32145 , \32146 , \32147 , \32148 , \32149 , \32150 , \32151 , \32152 ,
         \32153 , \32154 , \32155 , \32156 , \32157 , \32158 , \32159 , \32160 , \32161 , \32162 ,
         \32163 , \32164 , \32165 , \32166 , \32167 , \32168 , \32169 , \32170 , \32171 , \32172 ,
         \32173 , \32174 , \32175 , \32176 , \32177 , \32178 , \32179 , \32180 , \32181 , \32182 ,
         \32183 , \32184 , \32185 , \32186 , \32187 , \32188 , \32189 , \32190 , \32191 , \32192 ,
         \32193 , \32194 , \32195 , \32196 , \32197 , \32198 , \32199 , \32200 , \32201 , \32202 ,
         \32203 , \32204 , \32205 , \32206 , \32207 , \32208 , \32209 , \32210 , \32211 , \32212 ,
         \32213 , \32214 , \32215 , \32216 , \32217 , \32218 , \32219 , \32220 , \32221 , \32222 ,
         \32223 , \32224 , \32225 , \32226 , \32227 , \32228 , \32229 , \32230 , \32231 , \32232 ,
         \32233 , \32234 , \32235 , \32236 , \32237 , \32238 , \32239 , \32240 , \32241 , \32242 ,
         \32243 , \32244 , \32245 , \32246 , \32247 , \32248 , \32249 , \32250 , \32251 , \32252 ,
         \32253 , \32254 , \32255 , \32256 , \32257 , \32258 , \32259 , \32260 , \32261 , \32262 ,
         \32263 , \32264 , \32265 , \32266 , \32267 , \32268 , \32269 , \32270 , \32271 , \32272 ,
         \32273 , \32274 , \32275 , \32276 , \32277 , \32278 , \32279 , \32280 , \32281 , \32282 ,
         \32283 , \32284 , \32285 , \32286 , \32287 , \32288 , \32289 , \32290 , \32291 , \32292 ,
         \32293 , \32294 , \32295 , \32296 , \32297 , \32298 , \32299 , \32300 , \32301 , \32302 ,
         \32303 , \32304 , \32305 , \32306 , \32307 , \32308 , \32309 , \32310 , \32311 , \32312 ,
         \32313 , \32314 , \32315 , \32316 , \32317 , \32318 , \32319 , \32320 , \32321 , \32322 ,
         \32323 , \32324 , \32325 , \32326 , \32327 , \32328 , \32329 , \32330 , \32331 , \32332 ,
         \32333 , \32334 , \32335 , \32336 , \32337 , \32338 , \32339 , \32340 , \32341 , \32342 ,
         \32343 , \32344 , \32345 , \32346 , \32347 , \32348 , \32349 , \32350 , \32351 , \32352 ,
         \32353 , \32354 , \32355 , \32356 , \32357 , \32358 , \32359 , \32360 , \32361 , \32362 ,
         \32363 , \32364 , \32365 , \32366 , \32367 , \32368 , \32369 , \32370 , \32371 , \32372 ,
         \32373 , \32374 , \32375 , \32376 , \32377 , \32378 , \32379 , \32380 , \32381 , \32382 ,
         \32383 , \32384 , \32385 , \32386 , \32387 , \32388 , \32389 , \32390 , \32391 , \32392 ,
         \32393 , \32394 , \32395 , \32396 , \32397 , \32398 , \32399 , \32400 , \32401 , \32402 ,
         \32403 , \32404 , \32405 , \32406 , \32407 , \32408 , \32409 , \32410 , \32411 , \32412 ,
         \32413 , \32414 , \32415 , \32416 , \32417 , \32418 , \32419 , \32420 , \32421 , \32422 ,
         \32423 , \32424 , \32425 , \32426 , \32427 , \32428 , \32429 , \32430 , \32431 , \32432 ,
         \32433 , \32434 , \32435 , \32436 , \32437 , \32438 , \32439 , \32440 , \32441 , \32442 ,
         \32443 , \32444 , \32445 , \32446 , \32447 , \32448 , \32449 , \32450 , \32451 , \32452 ,
         \32453 , \32454 , \32455 , \32456 , \32457 , \32458 , \32459 , \32460 , \32461 , \32462 ,
         \32463 , \32464 , \32465 , \32466 , \32467 , \32468 , \32469 , \32470 , \32471 , \32472 ,
         \32473 , \32474 , \32475 , \32476 , \32477 , \32478 , \32479 , \32480 , \32481 , \32482 ,
         \32483 , \32484 , \32485 , \32486 , \32487 , \32488 , \32489 , \32490 , \32491 , \32492 ,
         \32493 , \32494 , \32495 , \32496 , \32497 , \32498 , \32499 , \32500 , \32501 , \32502 ,
         \32503 , \32504 , \32505 , \32506 , \32507 , \32508 , \32509 , \32510 , \32511 , \32512 ,
         \32513 , \32514 , \32515 , \32516 , \32517 , \32518 , \32519 , \32520 , \32521 , \32522 ,
         \32523 , \32524 , \32525 , \32526 , \32527 , \32528 , \32529 , \32530 , \32531 , \32532 ,
         \32533 , \32534 , \32535 , \32536 , \32537 , \32538 , \32539 , \32540 , \32541 , \32542 ,
         \32543 , \32544 , \32545 , \32546 , \32547 , \32548 , \32549 , \32550 , \32551 , \32552 ,
         \32553 , \32554 , \32555 , \32556 , \32557 , \32558 , \32559 , \32560 , \32561 , \32562 ,
         \32563 , \32564 , \32565 , \32566 , \32567 , \32568 , \32569 , \32570 , \32571 , \32572 ,
         \32573 , \32574 , \32575 , \32576 , \32577 , \32578 , \32579 , \32580 , \32581 , \32582 ,
         \32583 , \32584 , \32585 , \32586 , \32587 , \32588 , \32589 , \32590 , \32591 , \32592 ,
         \32593 , \32594 , \32595 , \32596 , \32597 , \32598 , \32599 , \32600 , \32601 , \32602 ,
         \32603 , \32604 , \32605 , \32606 , \32607 , \32608 , \32609 , \32610 , \32611 , \32612 ,
         \32613 , \32614 , \32615 , \32616 , \32617 , \32618 , \32619 , \32620 , \32621 , \32622 ,
         \32623 , \32624 , \32625 , \32626 , \32627 , \32628 , \32629 , \32630 , \32631 , \32632 ,
         \32633 , \32634 , \32635 , \32636 , \32637 , \32638 , \32639 , \32640 , \32641 , \32642 ,
         \32643 , \32644 , \32645 , \32646 , \32647 , \32648 , \32649 , \32650 , \32651 , \32652 ,
         \32653 , \32654 , \32655 , \32656 , \32657 , \32658 , \32659 , \32660 , \32661 , \32662 ,
         \32663 , \32664 , \32665 , \32666 , \32667 , \32668 , \32669 , \32670 , \32671 , \32672 ,
         \32673 , \32674 , \32675 , \32676 , \32677 , \32678 , \32679 , \32680 , \32681 , \32682 ,
         \32683 , \32684 , \32685 , \32686 , \32687 , \32688 , \32689 , \32690 , \32691 , \32692 ,
         \32693 , \32694 , \32695 , \32696 , \32697 , \32698 , \32699 , \32700 , \32701 , \32702 ,
         \32703 , \32704 , \32705 , \32706 , \32707 , \32708 , \32709 , \32710 , \32711 , \32712 ,
         \32713 , \32714 , \32715 , \32716 , \32717 , \32718 , \32719 , \32720 , \32721 , \32722 ,
         \32723 , \32724 , \32725 , \32726 , \32727 , \32728 , \32729 , \32730 , \32731 , \32732 ,
         \32733 , \32734 , \32735 , \32736 , \32737 , \32738 , \32739 , \32740 , \32741 , \32742 ,
         \32743 , \32744 , \32745 , \32746 , \32747 , \32748 , \32749 , \32750 , \32751 , \32752 ,
         \32753 , \32754 , \32755 , \32756 , \32757 , \32758 , \32759 , \32760 , \32761 , \32762 ,
         \32763 , \32764 , \32765 , \32766 , \32767 , \32768 , \32769 , \32770 , \32771 , \32772 ,
         \32773 , \32774 , \32775 , \32776 , \32777 , \32778 , \32779 , \32780 , \32781 , \32782 ,
         \32783 , \32784 , \32785 , \32786 , \32787 , \32788 , \32789 , \32790 , \32791 , \32792 ,
         \32793 , \32794 , \32795 , \32796 , \32797 , \32798 , \32799 , \32800 , \32801 , \32802 ,
         \32803 , \32804 , \32805 , \32806 , \32807 , \32808 , \32809 , \32810 , \32811 , \32812 ,
         \32813 , \32814 , \32815 , \32816 , \32817 , \32818 , \32819 , \32820 , \32821 , \32822 ,
         \32823 , \32824 , \32825 , \32826 , \32827 , \32828 , \32829 , \32830 , \32831 , \32832 ,
         \32833 , \32834 , \32835 , \32836 , \32837 , \32838 , \32839 , \32840 , \32841 , \32842 ,
         \32843 , \32844 , \32845 , \32846 , \32847 , \32848 , \32849 , \32850 , \32851 , \32852 ,
         \32853 , \32854 , \32855 , \32856 , \32857 , \32858 , \32859 , \32860 , \32861 , \32862 ,
         \32863 , \32864 , \32865 , \32866 , \32867 , \32868 , \32869 , \32870 , \32871 , \32872 ,
         \32873 , \32874 , \32875 , \32876 , \32877 , \32878 , \32879 , \32880 , \32881 , \32882 ,
         \32883 , \32884 , \32885 , \32886 , \32887 , \32888 , \32889 , \32890 , \32891 , \32892 ,
         \32893 , \32894 , \32895 , \32896 , \32897 , \32898 , \32899 , \32900 , \32901 , \32902 ,
         \32903 , \32904 , \32905 , \32906 , \32907 , \32908 , \32909 , \32910 , \32911 , \32912 ,
         \32913 , \32914 , \32915 , \32916 , \32917 , \32918 , \32919 , \32920 , \32921 , \32922 ,
         \32923 , \32924 , \32925 , \32926 , \32927 , \32928 , \32929 , \32930 , \32931 , \32932 ,
         \32933 , \32934 , \32935 , \32936 , \32937 , \32938 , \32939 , \32940 , \32941 , \32942 ,
         \32943 , \32944 , \32945 , \32946 , \32947 , \32948 , \32949 , \32950 , \32951 , \32952 ,
         \32953 , \32954 , \32955 , \32956 , \32957 , \32958 , \32959 , \32960 , \32961 , \32962 ,
         \32963 , \32964 , \32965 , \32966 , \32967 , \32968 , \32969 , \32970 , \32971 , \32972 ,
         \32973 , \32974 , \32975 , \32976 , \32977 , \32978 , \32979 , \32980 , \32981 , \32982 ,
         \32983 , \32984 , \32985 , \32986 , \32987 , \32988 , \32989 , \32990 , \32991 , \32992 ,
         \32993 , \32994 , \32995 , \32996 , \32997 , \32998 , \32999 , \33000 , \33001 , \33002 ,
         \33003 , \33004 , \33005 , \33006 , \33007 , \33008 , \33009 , \33010 , \33011 , \33012 ,
         \33013 , \33014 , \33015 , \33016 , \33017 , \33018 , \33019 , \33020 , \33021 , \33022 ,
         \33023 , \33024 , \33025 , \33026 , \33027 , \33028 , \33029 , \33030 , \33031 , \33032 ,
         \33033 , \33034 , \33035 , \33036 , \33037 , \33038 , \33039 , \33040 , \33041 , \33042 ,
         \33043 , \33044 , \33045 , \33046 , \33047 , \33048 , \33049 , \33050 , \33051 , \33052 ,
         \33053 , \33054 , \33055 , \33056 , \33057 , \33058 , \33059 , \33060 , \33061 , \33062 ,
         \33063 , \33064 , \33065 , \33066 , \33067 , \33068 , \33069 , \33070 , \33071 , \33072 ,
         \33073 , \33074 , \33075 , \33076 , \33077 , \33078 , \33079 , \33080 , \33081 , \33082 ,
         \33083 , \33084 , \33085 , \33086 , \33087 , \33088 , \33089 , \33090 , \33091 , \33092 ,
         \33093 , \33094 , \33095 , \33096 , \33097 , \33098 , \33099 , \33100 , \33101 , \33102 ,
         \33103 , \33104 , \33105 , \33106 , \33107 , \33108 , \33109 , \33110 , \33111 , \33112 ,
         \33113 , \33114 , \33115 , \33116 , \33117 , \33118 , \33119 , \33120 , \33121 , \33122 ,
         \33123 , \33124 , \33125 , \33126 , \33127 , \33128 , \33129 , \33130 , \33131 , \33132 ,
         \33133 , \33134 , \33135 , \33136 , \33137 , \33138 , \33139 , \33140 , \33141 , \33142 ,
         \33143 , \33144 , \33145 , \33146 , \33147 , \33148 , \33149 , \33150 , \33151 , \33152 ,
         \33153 , \33154 , \33155 , \33156 , \33157 , \33158 , \33159 , \33160 , \33161 , \33162 ,
         \33163 , \33164 , \33165 , \33166 , \33167 , \33168 , \33169 , \33170 , \33171 , \33172 ,
         \33173 , \33174 , \33175 , \33176 , \33177 , \33178 , \33179 , \33180 , \33181 , \33182 ,
         \33183 , \33184 , \33185 , \33186 , \33187 , \33188 , \33189 , \33190 , \33191 , \33192 ,
         \33193 , \33194 , \33195 , \33196 , \33197 , \33198 , \33199 , \33200 , \33201 , \33202 ,
         \33203 , \33204 , \33205 , \33206 , \33207 , \33208 , \33209 , \33210 , \33211 , \33212 ,
         \33213 , \33214 , \33215 , \33216 , \33217 , \33218 , \33219 , \33220 , \33221 , \33222 ,
         \33223 , \33224 , \33225 , \33226 , \33227 , \33228 , \33229 , \33230 , \33231 , \33232 ,
         \33233 , \33234 , \33235 , \33236 , \33237 , \33238 , \33239 , \33240 , \33241 , \33242 ,
         \33243 , \33244 , \33245 , \33246 , \33247 , \33248 , \33249 , \33250 , \33251 , \33252 ,
         \33253 , \33254 , \33255 , \33256 , \33257 , \33258 , \33259 , \33260 , \33261 , \33262 ,
         \33263 , \33264 , \33265 , \33266 , \33267 , \33268 , \33269 , \33270 , \33271 , \33272 ,
         \33273 , \33274 , \33275 , \33276 , \33277 , \33278 , \33279 , \33280 , \33281 , \33282 ,
         \33283 , \33284 , \33285 , \33286 , \33287 , \33288 , \33289 , \33290 , \33291 , \33292 ,
         \33293 , \33294 , \33295 , \33296 , \33297 , \33298 , \33299 , \33300 , \33301 , \33302 ,
         \33303 , \33304 , \33305 , \33306 , \33307 , \33308 , \33309 , \33310 , \33311 , \33312 ,
         \33313 , \33314 , \33315 , \33316 , \33317 , \33318 , \33319 , \33320 , \33321 , \33322 ,
         \33323 , \33324 , \33325 , \33326 , \33327 , \33328 , \33329 , \33330 , \33331 , \33332 ,
         \33333 , \33334 , \33335 , \33336 , \33337 , \33338 , \33339 , \33340 , \33341 , \33342 ,
         \33343 , \33344 , \33345 , \33346 , \33347 , \33348 , \33349 , \33350 , \33351 , \33352 ,
         \33353 , \33354 , \33355 , \33356 , \33357 , \33358 , \33359 , \33360 , \33361 , \33362 ,
         \33363 , \33364 , \33365 , \33366 , \33367 , \33368 , \33369 , \33370 , \33371 , \33372 ,
         \33373 , \33374 , \33375 , \33376 , \33377 , \33378 , \33379 , \33380 , \33381 , \33382 ,
         \33383 , \33384 , \33385 , \33386 , \33387 , \33388 , \33389 , \33390 , \33391 , \33392 ,
         \33393 , \33394 , \33395 , \33396 , \33397 , \33398 , \33399 , \33400 , \33401 , \33402 ,
         \33403 , \33404 , \33405 , \33406 , \33407 , \33408 , \33409 , \33410 , \33411 , \33412 ,
         \33413 , \33414 , \33415 , \33416 , \33417 , \33418 , \33419 , \33420 , \33421 , \33422 ,
         \33423 , \33424 , \33425 , \33426 , \33427 , \33428 , \33429 , \33430 , \33431 , \33432 ,
         \33433 , \33434 , \33435 , \33436 , \33437 , \33438 , \33439 , \33440 , \33441 , \33442 ,
         \33443 , \33444 , \33445 , \33446 , \33447 , \33448 , \33449 , \33450 , \33451 , \33452 ,
         \33453 , \33454 , \33455 , \33456 , \33457 , \33458 , \33459 , \33460 , \33461 , \33462 ,
         \33463 , \33464 , \33465 , \33466 , \33467 , \33468 , \33469 , \33470 , \33471 , \33472 ,
         \33473 , \33474 , \33475 , \33476 , \33477 , \33478 , \33479 , \33480 , \33481 , \33482 ,
         \33483 , \33484 , \33485 , \33486 , \33487 , \33488 , \33489 , \33490 , \33491 , \33492 ,
         \33493 , \33494 , \33495 , \33496 , \33497 , \33498 , \33499 , \33500 , \33501 , \33502 ,
         \33503 , \33504 , \33505 , \33506 , \33507 , \33508 , \33509 , \33510 , \33511 , \33512 ,
         \33513 , \33514 , \33515 , \33516 , \33517 , \33518 , \33519 , \33520 , \33521 , \33522 ,
         \33523 , \33524 , \33525 , \33526 , \33527 , \33528 , \33529 , \33530 , \33531 , \33532 ,
         \33533 , \33534 , \33535 , \33536 , \33537 , \33538 , \33539 , \33540 , \33541 , \33542 ,
         \33543 , \33544 , \33545 , \33546 , \33547 , \33548 , \33549 , \33550 , \33551 , \33552 ,
         \33553 , \33554 , \33555 , \33556 , \33557 , \33558 , \33559 , \33560 , \33561 , \33562 ,
         \33563 , \33564 , \33565 , \33566 , \33567 , \33568 , \33569 , \33570 , \33571 , \33572 ,
         \33573 , \33574 , \33575 , \33576 , \33577 , \33578 , \33579 , \33580 , \33581 , \33582 ,
         \33583 , \33584 , \33585 , \33586 , \33587 , \33588 , \33589 , \33590 , \33591 , \33592 ,
         \33593 , \33594 , \33595 , \33596 , \33597 , \33598 , \33599 , \33600 , \33601 , \33602 ,
         \33603 , \33604 , \33605 , \33606 , \33607 , \33608 , \33609 , \33610 , \33611 , \33612 ,
         \33613 , \33614 , \33615 , \33616 , \33617 , \33618 , \33619 , \33620 , \33621 , \33622 ,
         \33623 , \33624 , \33625 , \33626 , \33627 , \33628 , \33629 , \33630 , \33631 , \33632 ,
         \33633 , \33634 , \33635 , \33636 , \33637 , \33638 , \33639 , \33640 , \33641 , \33642 ,
         \33643 , \33644 , \33645 , \33646 , \33647 , \33648 , \33649 , \33650 , \33651 , \33652 ,
         \33653 , \33654 , \33655 , \33656 , \33657 , \33658 , \33659 , \33660 , \33661 , \33662 ,
         \33663 , \33664 , \33665 , \33666 , \33667 , \33668 , \33669 , \33670 , \33671 , \33672 ,
         \33673 , \33674 , \33675 , \33676 , \33677 , \33678 , \33679 , \33680 , \33681 , \33682 ,
         \33683 , \33684 , \33685 , \33686 , \33687 , \33688 , \33689 , \33690 , \33691 , \33692 ,
         \33693 , \33694 , \33695 , \33696 , \33697 , \33698 , \33699 , \33700 , \33701 , \33702 ,
         \33703 , \33704 , \33705 , \33706 , \33707 , \33708 , \33709 , \33710 , \33711 , \33712 ,
         \33713 , \33714 , \33715 , \33716 , \33717 , \33718 , \33719 , \33720 , \33721 , \33722 ,
         \33723 , \33724 , \33725 , \33726 , \33727 , \33728 , \33729 , \33730 , \33731 , \33732 ,
         \33733 , \33734 , \33735 , \33736 , \33737 , \33738 , \33739 , \33740 , \33741 , \33742 ,
         \33743 , \33744 , \33745 , \33746 , \33747 , \33748 , \33749 , \33750 , \33751 , \33752 ,
         \33753 , \33754 , \33755 , \33756 , \33757 , \33758 , \33759 , \33760 , \33761 , \33762 ,
         \33763 , \33764 , \33765 , \33766 , \33767 , \33768 , \33769 , \33770 , \33771 , \33772 ,
         \33773 , \33774 , \33775 , \33776 , \33777 , \33778 , \33779 , \33780 , \33781 , \33782 ,
         \33783 , \33784 , \33785 , \33786 , \33787 , \33788 , \33789 , \33790 , \33791 , \33792 ,
         \33793 , \33794 , \33795 , \33796 , \33797 , \33798 , \33799 , \33800 , \33801 , \33802 ,
         \33803 , \33804 , \33805 , \33806 , \33807 , \33808 , \33809 , \33810 , \33811 , \33812 ,
         \33813 , \33814 , \33815 , \33816 , \33817 , \33818 , \33819 , \33820 , \33821 , \33822 ,
         \33823 , \33824 , \33825 , \33826 , \33827 , \33828 , \33829 , \33830 , \33831 , \33832 ,
         \33833 , \33834 , \33835 , \33836 , \33837 , \33838 , \33839 , \33840 , \33841 , \33842 ,
         \33843 , \33844 , \33845 , \33846 , \33847 , \33848 , \33849 , \33850 , \33851 , \33852 ,
         \33853 , \33854 , \33855 , \33856 , \33857 , \33858 , \33859 , \33860 , \33861 , \33862 ,
         \33863 , \33864 , \33865 , \33866 , \33867 , \33868 , \33869 , \33870 , \33871 , \33872 ,
         \33873 , \33874 , \33875 , \33876 , \33877 , \33878 , \33879 , \33880 , \33881 , \33882 ,
         \33883 , \33884 , \33885 , \33886 , \33887 , \33888 , \33889 , \33890 , \33891 , \33892 ,
         \33893 , \33894 , \33895 , \33896 , \33897 , \33898 , \33899 , \33900 , \33901 , \33902 ,
         \33903 , \33904 , \33905 , \33906 , \33907 , \33908 , \33909 , \33910 , \33911 , \33912 ,
         \33913 , \33914 , \33915 , \33916 , \33917 , \33918 , \33919 , \33920 , \33921 , \33922 ,
         \33923 , \33924 , \33925 , \33926 , \33927 , \33928 , \33929 , \33930 , \33931 , \33932 ,
         \33933 , \33934 , \33935 , \33936 , \33937 , \33938 , \33939 , \33940 , \33941 , \33942 ,
         \33943 , \33944 , \33945 , \33946 , \33947 , \33948 , \33949 , \33950 , \33951 , \33952 ,
         \33953 , \33954 , \33955 , \33956 , \33957 , \33958 , \33959 , \33960 , \33961 , \33962 ,
         \33963 , \33964 , \33965 , \33966 , \33967 , \33968 , \33969 , \33970 , \33971 , \33972 ,
         \33973 , \33974 , \33975 , \33976 , \33977 , \33978 , \33979 , \33980 , \33981 , \33982 ,
         \33983 , \33984 , \33985 , \33986 , \33987 , \33988 , \33989 , \33990 , \33991 , \33992 ,
         \33993 , \33994 , \33995 , \33996 , \33997 , \33998 , \33999 , \34000 , \34001 , \34002 ,
         \34003 , \34004 , \34005 , \34006 , \34007 , \34008 , \34009 , \34010 , \34011 , \34012 ,
         \34013 , \34014 , \34015 , \34016 , \34017 , \34018 , \34019 , \34020 , \34021 , \34022 ,
         \34023 , \34024 , \34025 , \34026 , \34027 , \34028 , \34029 , \34030 , \34031 , \34032 ,
         \34033 , \34034 , \34035 , \34036 , \34037 , \34038 , \34039 , \34040 , \34041 , \34042 ,
         \34043 , \34044 , \34045 , \34046 , \34047 , \34048 , \34049 , \34050 , \34051 , \34052 ,
         \34053 , \34054 , \34055 , \34056 , \34057 , \34058 , \34059 , \34060 , \34061 , \34062 ,
         \34063 , \34064 , \34065 , \34066 , \34067 , \34068 , \34069 , \34070 , \34071 , \34072 ,
         \34073 , \34074 , \34075 , \34076 , \34077 , \34078 , \34079 , \34080 , \34081 , \34082 ,
         \34083 , \34084 , \34085 , \34086 , \34087 , \34088 , \34089 , \34090 , \34091 , \34092 ,
         \34093 , \34094 , \34095 , \34096 , \34097 , \34098 , \34099 , \34100 , \34101 , \34102 ,
         \34103 , \34104 , \34105 , \34106 , \34107 , \34108 , \34109 , \34110 , \34111 , \34112 ,
         \34113 , \34114 , \34115 , \34116 , \34117 , \34118 , \34119 , \34120 , \34121 , \34122 ,
         \34123 , \34124 , \34125 , \34126 , \34127 , \34128 , \34129 , \34130 , \34131 , \34132 ,
         \34133 , \34134 , \34135 , \34136 , \34137 , \34138 , \34139 , \34140 , \34141 , \34142 ,
         \34143 , \34144 , \34145 , \34146 , \34147 , \34148 , \34149 , \34150 , \34151 , \34152 ,
         \34153 , \34154 , \34155 , \34156 , \34157 , \34158 , \34159 , \34160 , \34161 , \34162 ,
         \34163 , \34164 , \34165 , \34166 , \34167 , \34168 , \34169 , \34170 , \34171 , \34172 ,
         \34173 , \34174 , \34175 , \34176 , \34177 , \34178 , \34179 , \34180 , \34181 , \34182 ,
         \34183 , \34184 , \34185 , \34186 , \34187 , \34188 , \34189 , \34190 , \34191 , \34192 ,
         \34193 , \34194 , \34195 , \34196 , \34197 , \34198 , \34199 , \34200 , \34201 , \34202 ,
         \34203 , \34204 , \34205 , \34206 , \34207 , \34208 , \34209 , \34210 , \34211 , \34212 ,
         \34213 , \34214 , \34215 , \34216 , \34217 , \34218 , \34219 , \34220 , \34221 , \34222 ,
         \34223 , \34224 , \34225 , \34226 , \34227 , \34228 , \34229 , \34230 , \34231 , \34232 ,
         \34233 , \34234 , \34235 , \34236 , \34237 , \34238 , \34239 , \34240 , \34241 , \34242 ,
         \34243 , \34244 , \34245 , \34246 , \34247 , \34248 , \34249 , \34250 , \34251 , \34252 ,
         \34253 , \34254 , \34255 , \34256 , \34257 , \34258 , \34259 , \34260 , \34261 , \34262 ,
         \34263 , \34264 , \34265 , \34266 , \34267 , \34268 , \34269 , \34270 , \34271 , \34272 ,
         \34273 , \34274 , \34275 , \34276 , \34277 , \34278 , \34279 , \34280 , \34281 , \34282 ,
         \34283 , \34284 , \34285 , \34286 , \34287 , \34288 , \34289 , \34290 , \34291 , \34292 ,
         \34293 , \34294 , \34295 , \34296 , \34297 , \34298 , \34299 , \34300 , \34301 , \34302 ,
         \34303 , \34304 , \34305 , \34306 , \34307 , \34308 , \34309 , \34310 , \34311 , \34312 ,
         \34313 , \34314 , \34315 , \34316 , \34317 , \34318 , \34319 , \34320 , \34321 , \34322 ,
         \34323 , \34324 , \34325 , \34326 , \34327 , \34328 , \34329 , \34330 , \34331 , \34332 ,
         \34333 , \34334 , \34335 , \34336 , \34337 , \34338 , \34339 , \34340 , \34341 , \34342 ,
         \34343 , \34344 , \34345 , \34346 , \34347 , \34348 , \34349 , \34350 , \34351 , \34352 ,
         \34353 , \34354 , \34355 , \34356 , \34357 , \34358 , \34359 , \34360 , \34361 , \34362 ,
         \34363 , \34364 , \34365 , \34366 , \34367 , \34368 , \34369 , \34370 , \34371 , \34372 ,
         \34373 , \34374 , \34375 , \34376 , \34377 , \34378 , \34379 , \34380 , \34381 , \34382 ,
         \34383 , \34384 , \34385 , \34386 , \34387 , \34388 , \34389 , \34390 , \34391 , \34392 ,
         \34393 , \34394 , \34395 , \34396 , \34397 , \34398 , \34399 , \34400 , \34401 , \34402 ,
         \34403 , \34404 , \34405 , \34406 , \34407 , \34408 , \34409 , \34410 , \34411 , \34412 ,
         \34413 , \34414 , \34415 , \34416 , \34417 , \34418 , \34419 , \34420 , \34421 , \34422 ,
         \34423 , \34424 , \34425 , \34426 , \34427 , \34428 , \34429 , \34430 , \34431 , \34432 ,
         \34433 , \34434 , \34435 , \34436 , \34437 , \34438 , \34439 , \34440 , \34441 , \34442 ,
         \34443 , \34444 , \34445 , \34446 , \34447 , \34448 , \34449 , \34450 , \34451 , \34452 ,
         \34453 , \34454 , \34455 , \34456 , \34457 , \34458 , \34459 , \34460 , \34461 , \34462 ,
         \34463 , \34464 , \34465 , \34466 , \34467 , \34468 , \34469 , \34470 , \34471 , \34472 ,
         \34473 , \34474 , \34475 , \34476 , \34477 , \34478 , \34479 , \34480 , \34481 , \34482 ,
         \34483 , \34484 , \34485 , \34486 , \34487 , \34488 , \34489 , \34490 , \34491 , \34492 ,
         \34493 , \34494 , \34495 , \34496 , \34497 , \34498 , \34499 , \34500 , \34501 , \34502 ,
         \34503 , \34504 , \34505 , \34506 , \34507 , \34508 , \34509 , \34510 , \34511 , \34512 ,
         \34513 , \34514 , \34515 , \34516 , \34517 , \34518 , \34519 , \34520 , \34521 , \34522 ,
         \34523 , \34524 , \34525 , \34526 , \34527 , \34528 , \34529 , \34530 , \34531 , \34532 ,
         \34533 , \34534 , \34535 , \34536 , \34537 , \34538 , \34539 , \34540 , \34541 , \34542 ,
         \34543 , \34544 , \34545 , \34546 , \34547 , \34548 , \34549 , \34550 , \34551 , \34552 ,
         \34553 , \34554 , \34555 , \34556 , \34557 , \34558 , \34559 , \34560 , \34561 , \34562 ,
         \34563 , \34564 , \34565 , \34566 , \34567 , \34568 , \34569 , \34570 , \34571 , \34572 ,
         \34573 , \34574 , \34575 , \34576 , \34577 , \34578 , \34579 , \34580 , \34581 , \34582 ,
         \34583 , \34584 , \34585 , \34586 , \34587 , \34588 , \34589 , \34590 , \34591 , \34592 ,
         \34593 , \34594 , \34595 , \34596 , \34597 , \34598 , \34599 , \34600 , \34601 , \34602 ,
         \34603 , \34604 , \34605 , \34606 , \34607 , \34608 , \34609 , \34610 , \34611 , \34612 ,
         \34613 , \34614 , \34615 , \34616 , \34617 , \34618 , \34619 , \34620 , \34621 , \34622 ,
         \34623 , \34624 , \34625 , \34626 , \34627 , \34628 , \34629 , \34630 , \34631 , \34632 ,
         \34633 , \34634 , \34635 , \34636 , \34637 , \34638 , \34639 , \34640 , \34641 , \34642 ,
         \34643 , \34644 , \34645 , \34646 , \34647 , \34648 , \34649 , \34650 , \34651 , \34652 ,
         \34653 , \34654 , \34655 , \34656 , \34657 , \34658 , \34659 , \34660 , \34661 , \34662 ,
         \34663 , \34664 , \34665 , \34666 , \34667 , \34668 , \34669 , \34670 , \34671 , \34672 ,
         \34673 , \34674 , \34675 , \34676 , \34677 , \34678 , \34679 , \34680 , \34681 , \34682 ,
         \34683 , \34684 , \34685 , \34686 , \34687 , \34688 , \34689 , \34690 , \34691 , \34692 ,
         \34693 , \34694 , \34695 , \34696 , \34697 , \34698 , \34699 , \34700 , \34701 , \34702 ,
         \34703 , \34704 , \34705 , \34706 , \34707 , \34708 , \34709 , \34710 , \34711 , \34712 ,
         \34713 , \34714 , \34715 , \34716 , \34717 , \34718 , \34719 , \34720 , \34721 , \34722 ,
         \34723 , \34724 , \34725 , \34726 , \34727 , \34728 , \34729 , \34730 , \34731 , \34732 ,
         \34733 , \34734 , \34735 , \34736 , \34737 , \34738 , \34739 , \34740 , \34741 , \34742 ,
         \34743 , \34744 , \34745 , \34746 , \34747 , \34748 , \34749 , \34750 , \34751 , \34752 ,
         \34753 , \34754 , \34755 , \34756 , \34757 , \34758 , \34759 , \34760 , \34761 , \34762 ,
         \34763 , \34764 , \34765 , \34766 , \34767 , \34768 , \34769 , \34770 , \34771 , \34772 ,
         \34773 , \34774 , \34775 , \34776 , \34777 , \34778 , \34779 , \34780 , \34781 , \34782 ,
         \34783 , \34784 , \34785 , \34786 , \34787 , \34788 , \34789 , \34790 , \34791 , \34792 ,
         \34793 , \34794 , \34795 , \34796 , \34797 , \34798 , \34799 , \34800 , \34801 , \34802 ,
         \34803 , \34804 , \34805 , \34806 , \34807 , \34808 , \34809 , \34810 , \34811 , \34812 ,
         \34813 , \34814 , \34815 , \34816 , \34817 , \34818 , \34819 , \34820 , \34821 , \34822 ,
         \34823 , \34824 , \34825 , \34826 , \34827 , \34828 , \34829 , \34830 , \34831 , \34832 ,
         \34833 , \34834 , \34835 , \34836 , \34837 , \34838 , \34839 , \34840 , \34841 , \34842 ,
         \34843 , \34844 , \34845 , \34846 , \34847 , \34848 , \34849 , \34850 , \34851 , \34852 ,
         \34853 , \34854 , \34855 , \34856 , \34857 , \34858 , \34859 , \34860 , \34861 , \34862 ,
         \34863 , \34864 , \34865 , \34866 , \34867 , \34868 , \34869 , \34870 , \34871 , \34872 ,
         \34873 , \34874 , \34875 , \34876 , \34877 , \34878 , \34879 , \34880 , \34881 , \34882 ,
         \34883 , \34884 , \34885 , \34886 , \34887 , \34888 , \34889 , \34890 , \34891 , \34892 ,
         \34893 , \34894 , \34895 , \34896 , \34897 , \34898 , \34899 , \34900 , \34901 , \34902 ,
         \34903 , \34904 , \34905 , \34906 , \34907 , \34908 , \34909 , \34910 , \34911 , \34912 ,
         \34913 , \34914 , \34915 , \34916 , \34917 , \34918 , \34919 , \34920 , \34921 , \34922 ,
         \34923 , \34924 , \34925 , \34926 , \34927 , \34928 , \34929 , \34930 , \34931 , \34932 ,
         \34933 , \34934 , \34935 , \34936 , \34937 , \34938 , \34939 , \34940 , \34941 , \34942 ,
         \34943 , \34944 , \34945 , \34946 , \34947 , \34948 , \34949 , \34950 , \34951 , \34952 ,
         \34953 , \34954 , \34955 , \34956 , \34957 , \34958 , \34959 , \34960 , \34961 , \34962 ,
         \34963 , \34964 , \34965 , \34966 , \34967 , \34968 , \34969 , \34970 , \34971 , \34972 ,
         \34973 , \34974 , \34975 , \34976 , \34977 , \34978 , \34979 , \34980 , \34981 , \34982 ,
         \34983 , \34984 , \34985 , \34986 , \34987 , \34988 , \34989 , \34990 , \34991 , \34992 ,
         \34993 , \34994 , \34995 , \34996 , \34997 , \34998 , \34999 , \35000 , \35001 , \35002 ,
         \35003 , \35004 , \35005 , \35006 , \35007 , \35008 , \35009 , \35010 , \35011 , \35012 ,
         \35013 , \35014 , \35015 , \35016 , \35017 , \35018 , \35019 , \35020 , \35021 , \35022 ,
         \35023 , \35024 , \35025 , \35026 , \35027 , \35028 , \35029 , \35030 , \35031 , \35032 ,
         \35033 , \35034 , \35035 , \35036 , \35037 , \35038 , \35039 , \35040 , \35041 , \35042 ,
         \35043 , \35044 , \35045 , \35046 , \35047 , \35048 , \35049 , \35050 , \35051 , \35052 ,
         \35053 , \35054 , \35055 , \35056 , \35057 , \35058 , \35059 , \35060 , \35061 , \35062 ,
         \35063 , \35064 , \35065 , \35066 , \35067 , \35068 , \35069 , \35070 , \35071 , \35072 ,
         \35073 , \35074 , \35075 , \35076 , \35077 , \35078 , \35079 , \35080 , \35081 , \35082 ,
         \35083 , \35084 , \35085 , \35086 , \35087 , \35088 , \35089 , \35090 , \35091 , \35092 ,
         \35093 , \35094 , \35095 , \35096 , \35097 , \35098 , \35099 , \35100 , \35101 , \35102 ,
         \35103 , \35104 , \35105 , \35106 , \35107 , \35108 , \35109 , \35110 , \35111 , \35112 ,
         \35113 , \35114 , \35115 , \35116 , \35117 , \35118 , \35119 , \35120 , \35121 , \35122 ,
         \35123 , \35124 , \35125 , \35126 , \35127 , \35128 , \35129 , \35130 , \35131 , \35132 ,
         \35133 , \35134 , \35135 , \35136 , \35137 , \35138 , \35139 , \35140 , \35141 , \35142 ,
         \35143 , \35144 , \35145 , \35146 , \35147 , \35148 , \35149 , \35150 , \35151 , \35152 ,
         \35153 , \35154 , \35155 , \35156 , \35157 , \35158 , \35159 , \35160 , \35161 , \35162 ,
         \35163 , \35164 , \35165 , \35166 , \35167 , \35168 , \35169 , \35170 , \35171 , \35172 ,
         \35173 , \35174 , \35175 , \35176 , \35177 , \35178 , \35179 , \35180 , \35181 , \35182 ,
         \35183 , \35184 , \35185 , \35186 , \35187 , \35188 , \35189 , \35190 , \35191 , \35192 ,
         \35193 , \35194 , \35195 , \35196 , \35197 , \35198 , \35199 , \35200 , \35201 , \35202 ,
         \35203 , \35204 , \35205 , \35206 , \35207 , \35208 , \35209 , \35210 , \35211 , \35212 ,
         \35213 , \35214 , \35215 , \35216 , \35217 , \35218 , \35219 , \35220 , \35221 , \35222 ,
         \35223 , \35224 , \35225 , \35226 , \35227 , \35228 , \35229 , \35230 , \35231 , \35232 ,
         \35233 , \35234 , \35235 , \35236 , \35237 , \35238 , \35239 , \35240 , \35241 , \35242 ,
         \35243 , \35244 , \35245 , \35246 , \35247 , \35248 , \35249 , \35250 , \35251 , \35252 ,
         \35253 , \35254 , \35255 , \35256 , \35257 , \35258 , \35259 , \35260 , \35261 , \35262 ,
         \35263 , \35264 , \35265 , \35266 , \35267 , \35268 , \35269 , \35270 , \35271 , \35272 ,
         \35273 , \35274 , \35275 , \35276 , \35277 , \35278 , \35279 , \35280 , \35281 , \35282 ,
         \35283 , \35284 , \35285 , \35286 , \35287 , \35288 , \35289 , \35290 , \35291 , \35292 ,
         \35293 , \35294 , \35295 , \35296 , \35297 , \35298 , \35299 , \35300 , \35301 , \35302 ,
         \35303 , \35304 , \35305 , \35306 , \35307 , \35308 , \35309 , \35310 , \35311 , \35312 ,
         \35313 , \35314 , \35315 , \35316 , \35317 , \35318 , \35319 , \35320 , \35321 , \35322 ,
         \35323 , \35324 , \35325 , \35326 , \35327 , \35328 , \35329 , \35330 , \35331 , \35332 ,
         \35333 , \35334 , \35335 , \35336 , \35337 , \35338 , \35339 , \35340 , \35341 , \35342 ,
         \35343 , \35344 , \35345 , \35346 , \35347 , \35348 , \35349 , \35350 , \35351 , \35352 ,
         \35353 , \35354 , \35355 , \35356 , \35357 , \35358 , \35359 , \35360 , \35361 , \35362 ,
         \35363 , \35364 , \35365 , \35366 , \35367 , \35368 , \35369 , \35370 , \35371 , \35372 ,
         \35373 , \35374 , \35375 , \35376 , \35377 , \35378 , \35379 , \35380 , \35381 , \35382 ,
         \35383 , \35384 , \35385 , \35386 , \35387 , \35388 , \35389 , \35390 , \35391 , \35392 ,
         \35393 , \35394 , \35395 , \35396 , \35397 , \35398 , \35399 , \35400 , \35401 , \35402 ,
         \35403 , \35404 , \35405 , \35406 , \35407 , \35408 , \35409 , \35410 , \35411 , \35412 ,
         \35413 , \35414 , \35415 , \35416 , \35417 , \35418 , \35419 , \35420 , \35421 , \35422 ,
         \35423 , \35424 , \35425 , \35426 , \35427 , \35428 , \35429 , \35430 , \35431 , \35432 ,
         \35433 , \35434 , \35435 , \35436 , \35437 , \35438 , \35439 , \35440 , \35441 , \35442 ,
         \35443 , \35444 , \35445 , \35446 , \35447 , \35448 , \35449 , \35450 , \35451 , \35452 ,
         \35453 , \35454 , \35455 , \35456 , \35457 , \35458 , \35459 , \35460 , \35461 , \35462 ,
         \35463 , \35464 , \35465 , \35466 , \35467 , \35468 , \35469 , \35470 , \35471 , \35472 ,
         \35473 , \35474 , \35475 , \35476 , \35477 , \35478 , \35479 , \35480 , \35481 , \35482 ,
         \35483 , \35484 , \35485 , \35486 , \35487 , \35488 , \35489 , \35490 , \35491 , \35492 ,
         \35493 , \35494 , \35495 , \35496 , \35497 , \35498 , \35499 , \35500 , \35501 , \35502 ,
         \35503 , \35504 , \35505 , \35506 , \35507 , \35508 , \35509 , \35510 , \35511 , \35512 ,
         \35513 , \35514 , \35515 , \35516 , \35517 , \35518 , \35519 , \35520 , \35521 , \35522 ,
         \35523 , \35524 , \35525 , \35526 , \35527 , \35528 , \35529 , \35530 , \35531 , \35532 ,
         \35533 , \35534 , \35535 , \35536 , \35537 , \35538 , \35539 , \35540 , \35541 , \35542 ,
         \35543 , \35544 , \35545 , \35546 , \35547 , \35548 , \35549 , \35550 , \35551 , \35552 ,
         \35553 , \35554 , \35555 , \35556 , \35557 , \35558 , \35559 , \35560 , \35561 , \35562 ,
         \35563 , \35564 , \35565 , \35566 , \35567 , \35568 , \35569 , \35570 , \35571 , \35572 ,
         \35573 , \35574 , \35575 , \35576 , \35577 , \35578 , \35579 , \35580 , \35581 , \35582 ,
         \35583 , \35584 , \35585 , \35586 , \35587 , \35588 , \35589 , \35590 , \35591 , \35592 ,
         \35593 , \35594 , \35595 , \35596 , \35597 , \35598 , \35599 , \35600 , \35601 , \35602 ,
         \35603 , \35604 , \35605 , \35606 , \35607 , \35608 , \35609 , \35610 , \35611 , \35612 ,
         \35613 , \35614 , \35615 , \35616 , \35617 , \35618 , \35619 , \35620 , \35621 , \35622 ,
         \35623 , \35624 , \35625 , \35626 , \35627 , \35628 , \35629 , \35630 , \35631 , \35632 ,
         \35633 , \35634 , \35635 , \35636 , \35637 , \35638 , \35639 , \35640 , \35641 , \35642 ,
         \35643 , \35644 , \35645 , \35646 , \35647 , \35648 , \35649 , \35650 , \35651 , \35652 ,
         \35653 , \35654 , \35655 , \35656 , \35657 , \35658 , \35659 , \35660 , \35661 , \35662 ,
         \35663 , \35664 , \35665 , \35666 , \35667 , \35668 , \35669 , \35670 , \35671 , \35672 ,
         \35673 , \35674 , \35675 , \35676 , \35677 , \35678 , \35679 , \35680 , \35681 , \35682 ,
         \35683 , \35684 , \35685 , \35686 , \35687 , \35688 , \35689 , \35690 , \35691 , \35692 ,
         \35693 , \35694 , \35695 , \35696 , \35697 , \35698 , \35699 , \35700 , \35701 , \35702 ,
         \35703 , \35704 , \35705 , \35706 , \35707 , \35708 , \35709 , \35710 , \35711 , \35712 ,
         \35713 , \35714 , \35715 , \35716 , \35717 , \35718 , \35719 , \35720 , \35721 , \35722 ,
         \35723 , \35724 , \35725 , \35726 , \35727 , \35728 , \35729 , \35730 , \35731 , \35732 ,
         \35733 , \35734 , \35735 , \35736 , \35737 , \35738 , \35739 , \35740 , \35741 , \35742 ,
         \35743 , \35744 , \35745 , \35746 , \35747 , \35748 , \35749 , \35750 , \35751 , \35752 ,
         \35753 , \35754 , \35755 , \35756 , \35757 , \35758 , \35759 , \35760 , \35761 , \35762 ,
         \35763 , \35764 , \35765 , \35766 , \35767 , \35768 , \35769 , \35770 , \35771 , \35772 ,
         \35773 , \35774 , \35775 , \35776 , \35777 , \35778 , \35779 , \35780 , \35781 , \35782 ,
         \35783 , \35784 , \35785 , \35786 , \35787 , \35788 , \35789 , \35790 , \35791 , \35792 ,
         \35793 , \35794 , \35795 , \35796 , \35797 , \35798 , \35799 , \35800 , \35801 , \35802 ,
         \35803 , \35804 , \35805 , \35806 , \35807 , \35808 , \35809 , \35810 , \35811 , \35812 ,
         \35813 , \35814 , \35815 , \35816 , \35817 , \35818 , \35819 , \35820 , \35821 , \35822 ,
         \35823 , \35824 , \35825 , \35826 , \35827 , \35828 , \35829 , \35830 , \35831 , \35832 ,
         \35833 , \35834 , \35835 , \35836 , \35837 , \35838 , \35839 , \35840 , \35841 , \35842 ,
         \35843 , \35844 , \35845 , \35846 , \35847 , \35848 , \35849 , \35850 , \35851 , \35852 ,
         \35853 , \35854 , \35855 , \35856 , \35857 , \35858 , \35859 , \35860 , \35861 , \35862 ,
         \35863 , \35864 , \35865 , \35866 , \35867 , \35868 , \35869 , \35870 , \35871 , \35872 ,
         \35873 , \35874 , \35875 , \35876 , \35877 , \35878 , \35879 , \35880 , \35881 , \35882 ,
         \35883 , \35884 , \35885 , \35886 , \35887 , \35888 , \35889 , \35890 , \35891 , \35892 ,
         \35893 , \35894 , \35895 , \35896 , \35897 , \35898 , \35899 , \35900 , \35901 , \35902 ,
         \35903 , \35904 , \35905 , \35906 , \35907 , \35908 , \35909 , \35910 , \35911 , \35912 ,
         \35913 , \35914 , \35915 , \35916 , \35917 , \35918 , \35919 , \35920 , \35921 , \35922 ,
         \35923 , \35924 , \35925 , \35926 , \35927 , \35928 , \35929 , \35930 , \35931 , \35932 ,
         \35933 , \35934 , \35935 , \35936 , \35937 , \35938 , \35939 , \35940 , \35941 , \35942 ,
         \35943 , \35944 , \35945 , \35946 , \35947 , \35948 , \35949 , \35950 , \35951 , \35952 ,
         \35953 , \35954 , \35955 , \35956 , \35957 , \35958 , \35959 , \35960 , \35961 , \35962 ,
         \35963 , \35964 , \35965 , \35966 , \35967 , \35968 , \35969 , \35970 , \35971 , \35972 ,
         \35973 , \35974 , \35975 , \35976 , \35977 , \35978 , \35979 , \35980 , \35981 , \35982 ,
         \35983 , \35984 , \35985 , \35986 , \35987 , \35988 , \35989 , \35990 , \35991 , \35992 ,
         \35993 , \35994 , \35995 , \35996 , \35997 , \35998 , \35999 , \36000 , \36001 , \36002 ,
         \36003 , \36004 , \36005 , \36006 , \36007 , \36008 , \36009 , \36010 , \36011 , \36012 ,
         \36013 , \36014 , \36015 , \36016 , \36017 , \36018 , \36019 , \36020 , \36021 , \36022 ,
         \36023 , \36024 , \36025 , \36026 , \36027 , \36028 , \36029 , \36030 , \36031 , \36032 ,
         \36033 , \36034 , \36035 , \36036 , \36037 , \36038 , \36039 , \36040 , \36041 , \36042 ,
         \36043 , \36044 , \36045 , \36046 , \36047 , \36048 , \36049 , \36050 , \36051 , \36052 ,
         \36053 , \36054 , \36055 , \36056 , \36057 , \36058 , \36059 , \36060 , \36061 , \36062 ,
         \36063 , \36064 , \36065 , \36066 , \36067 , \36068 , \36069 , \36070 , \36071 , \36072 ,
         \36073 , \36074 , \36075 , \36076 , \36077 , \36078 , \36079 , \36080 , \36081 , \36082 ,
         \36083 , \36084 , \36085 , \36086 , \36087 , \36088 , \36089 , \36090 , \36091 , \36092 ,
         \36093 , \36094 , \36095 , \36096 , \36097 , \36098 , \36099 , \36100 , \36101 , \36102 ,
         \36103 , \36104 , \36105 , \36106 , \36107 , \36108 , \36109 , \36110 , \36111 , \36112 ,
         \36113 , \36114 , \36115 , \36116 , \36117 , \36118 , \36119 , \36120 , \36121 , \36122 ,
         \36123 , \36124 , \36125 , \36126 , \36127 , \36128 , \36129 , \36130 , \36131 , \36132 ,
         \36133 , \36134 , \36135 , \36136 , \36137 , \36138 , \36139 , \36140 , \36141 , \36142 ,
         \36143 , \36144 , \36145 , \36146 , \36147 , \36148 , \36149 , \36150 , \36151 , \36152 ,
         \36153 , \36154 , \36155 , \36156 , \36157 , \36158 , \36159 , \36160 , \36161 , \36162 ,
         \36163 , \36164 , \36165 , \36166 , \36167 , \36168 , \36169 , \36170 , \36171 , \36172 ,
         \36173 , \36174 , \36175 , \36176 , \36177 , \36178 , \36179 , \36180 , \36181 , \36182 ,
         \36183 , \36184 , \36185 , \36186 , \36187 , \36188 , \36189 , \36190 , \36191 , \36192 ,
         \36193 , \36194 , \36195 , \36196 , \36197 , \36198 , \36199 , \36200 , \36201 , \36202 ,
         \36203 , \36204 , \36205 , \36206 , \36207 , \36208 , \36209 , \36210 , \36211 , \36212 ,
         \36213 , \36214 , \36215 , \36216 , \36217 , \36218 , \36219 , \36220 , \36221 , \36222 ,
         \36223 , \36224 , \36225 , \36226 , \36227 , \36228 , \36229 , \36230 , \36231 , \36232 ,
         \36233 , \36234 , \36235 , \36236 , \36237 , \36238 , \36239 , \36240 , \36241 , \36242 ,
         \36243 , \36244 , \36245 , \36246 , \36247 , \36248 , \36249 , \36250 , \36251 , \36252 ,
         \36253 , \36254 , \36255 , \36256 , \36257 , \36258 , \36259 , \36260 , \36261 , \36262 ,
         \36263 , \36264 , \36265 , \36266 , \36267 , \36268 , \36269 , \36270 , \36271 , \36272 ,
         \36273 , \36274 , \36275 , \36276 , \36277 , \36278 , \36279 , \36280 , \36281 , \36282 ,
         \36283 , \36284 , \36285 , \36286 , \36287 , \36288 , \36289 , \36290 , \36291 , \36292 ,
         \36293 , \36294 , \36295 , \36296 , \36297 , \36298 , \36299 , \36300 , \36301 , \36302 ,
         \36303 , \36304 , \36305 , \36306 , \36307 , \36308 , \36309 , \36310 , \36311 , \36312 ,
         \36313 , \36314 , \36315 , \36316 , \36317 , \36318 , \36319 , \36320 , \36321 , \36322 ,
         \36323 , \36324 , \36325 , \36326 , \36327 , \36328 , \36329 , \36330 , \36331 , \36332 ,
         \36333 , \36334 , \36335 , \36336 , \36337 , \36338 , \36339 , \36340 , \36341 , \36342 ,
         \36343 , \36344 , \36345 , \36346 , \36347 , \36348 , \36349 , \36350 , \36351 , \36352 ,
         \36353 , \36354 , \36355 , \36356 , \36357 , \36358 , \36359 , \36360 , \36361 , \36362 ,
         \36363 , \36364 , \36365 , \36366 , \36367 , \36368 , \36369 , \36370 , \36371 , \36372 ,
         \36373 , \36374 , \36375 , \36376 , \36377 , \36378 , \36379 , \36380 , \36381 , \36382 ,
         \36383 , \36384 , \36385 , \36386 , \36387 , \36388 , \36389 , \36390 , \36391 , \36392 ,
         \36393 , \36394 , \36395 , \36396 , \36397 , \36398 , \36399 , \36400 , \36401 , \36402 ,
         \36403 , \36404 , \36405 , \36406 , \36407 , \36408 , \36409 , \36410 , \36411 , \36412 ,
         \36413 , \36414 , \36415 , \36416 , \36417 , \36418 , \36419 , \36420 , \36421 , \36422 ,
         \36423 , \36424 , \36425 , \36426 , \36427 , \36428 , \36429 , \36430 , \36431 , \36432 ,
         \36433 , \36434 , \36435 , \36436 , \36437 , \36438 , \36439 , \36440 , \36441 , \36442 ,
         \36443 , \36444 , \36445 , \36446 , \36447 , \36448 , \36449 , \36450 , \36451 , \36452 ,
         \36453 , \36454 , \36455 , \36456 , \36457 , \36458 , \36459 , \36460 , \36461 , \36462 ,
         \36463 , \36464 , \36465 , \36466 , \36467 , \36468 , \36469 , \36470 , \36471 , \36472 ,
         \36473 , \36474 , \36475 , \36476 , \36477 , \36478 , \36479 , \36480 , \36481 , \36482 ,
         \36483 , \36484 , \36485 , \36486 , \36487 , \36488 , \36489 , \36490 , \36491 , \36492 ,
         \36493 , \36494 , \36495 , \36496 , \36497 , \36498 , \36499 , \36500 , \36501 , \36502 ,
         \36503 , \36504 , \36505 , \36506 , \36507 , \36508 , \36509 , \36510 , \36511 , \36512 ,
         \36513 , \36514 , \36515 , \36516 , \36517 , \36518 , \36519 , \36520 , \36521 , \36522 ,
         \36523 , \36524 , \36525 , \36526 , \36527 , \36528 , \36529 , \36530 , \36531 , \36532 ,
         \36533 , \36534 , \36535 , \36536 , \36537 , \36538 , \36539 , \36540 , \36541 , \36542 ,
         \36543 , \36544 , \36545 , \36546 , \36547 , \36548 , \36549 , \36550 , \36551 , \36552 ,
         \36553 , \36554 , \36555 , \36556 , \36557 , \36558 , \36559 , \36560 , \36561 , \36562 ,
         \36563 , \36564 , \36565 , \36566 , \36567 , \36568 , \36569 , \36570 , \36571 , \36572 ,
         \36573 , \36574 , \36575 , \36576 , \36577 , \36578 , \36579 , \36580 , \36581 , \36582 ,
         \36583 , \36584 , \36585 , \36586 , \36587 , \36588 , \36589 , \36590 , \36591 , \36592 ,
         \36593 , \36594 , \36595 , \36596 , \36597 , \36598 , \36599 , \36600 , \36601 , \36602 ,
         \36603 , \36604 , \36605 , \36606 , \36607 , \36608 , \36609 , \36610 , \36611 , \36612 ,
         \36613 , \36614 , \36615 , \36616 , \36617 , \36618 , \36619 , \36620 , \36621 , \36622 ,
         \36623 , \36624 , \36625 , \36626 , \36627 , \36628 , \36629 , \36630 , \36631 , \36632 ,
         \36633 , \36634 , \36635 , \36636 , \36637 , \36638 , \36639 , \36640 , \36641 , \36642 ,
         \36643 , \36644 , \36645 , \36646 , \36647 , \36648 , \36649 , \36650 , \36651 , \36652 ,
         \36653 , \36654 , \36655 , \36656 , \36657 , \36658 , \36659 , \36660 , \36661 , \36662 ,
         \36663 , \36664 , \36665 , \36666 , \36667 , \36668 , \36669 , \36670 , \36671 , \36672 ,
         \36673 , \36674 , \36675 , \36676 , \36677 , \36678 , \36679 , \36680 , \36681 , \36682 ,
         \36683 , \36684 , \36685 , \36686 , \36687 , \36688 , \36689 , \36690 , \36691 , \36692 ,
         \36693 , \36694 , \36695 , \36696 , \36697 , \36698 , \36699 , \36700 , \36701 , \36702 ,
         \36703 , \36704 , \36705 , \36706 , \36707 , \36708 , \36709 , \36710 , \36711 , \36712 ,
         \36713 , \36714 , \36715 , \36716 , \36717 , \36718 , \36719 , \36720 , \36721 , \36722 ,
         \36723 , \36724 , \36725 , \36726 , \36727 , \36728 , \36729 , \36730 , \36731 , \36732 ,
         \36733 , \36734 , \36735 , \36736 , \36737 , \36738 , \36739 , \36740 , \36741 , \36742 ,
         \36743 , \36744 , \36745 , \36746 , \36747 , \36748 , \36749 , \36750 , \36751 , \36752 ,
         \36753 , \36754 , \36755 , \36756 , \36757 , \36758 , \36759 , \36760 , \36761 , \36762 ,
         \36763 , \36764 , \36765 , \36766 , \36767 , \36768 , \36769 , \36770 , \36771 , \36772 ,
         \36773 , \36774 , \36775 , \36776 , \36777 , \36778 , \36779 , \36780 , \36781 , \36782 ,
         \36783 , \36784 , \36785 , \36786 , \36787 , \36788 , \36789 , \36790 , \36791 , \36792 ,
         \36793 , \36794 , \36795 , \36796 , \36797 , \36798 , \36799 , \36800 , \36801 , \36802 ,
         \36803 , \36804 , \36805 , \36806 , \36807 , \36808 , \36809 , \36810 , \36811 , \36812 ,
         \36813 , \36814 , \36815 , \36816 , \36817 , \36818 , \36819 , \36820 , \36821 , \36822 ,
         \36823 , \36824 , \36825 , \36826 , \36827 , \36828 , \36829 , \36830 , \36831 , \36832 ,
         \36833 , \36834 , \36835 , \36836 , \36837 , \36838 , \36839 , \36840 , \36841 , \36842 ,
         \36843 , \36844 , \36845 , \36846 , \36847 , \36848 , \36849 , \36850 , \36851 , \36852 ,
         \36853 , \36854 , \36855 , \36856 , \36857 , \36858 , \36859 , \36860 , \36861 , \36862 ,
         \36863 , \36864 , \36865 , \36866 , \36867 , \36868 , \36869 , \36870 , \36871 , \36872 ,
         \36873 , \36874 , \36875 , \36876 , \36877 , \36878 , \36879 , \36880 , \36881 , \36882 ,
         \36883 , \36884 , \36885 , \36886 , \36887 , \36888 , \36889 , \36890 , \36891 , \36892 ,
         \36893 , \36894 , \36895 , \36896 , \36897 , \36898 , \36899 , \36900 , \36901 , \36902 ,
         \36903 , \36904 , \36905 , \36906 , \36907 , \36908 , \36909 , \36910 , \36911 , \36912 ,
         \36913 , \36914 , \36915 , \36916 , \36917 , \36918 , \36919 , \36920 , \36921 , \36922 ,
         \36923 , \36924 , \36925 , \36926 , \36927 , \36928 , \36929 , \36930 , \36931 , \36932 ,
         \36933 , \36934 , \36935 , \36936 , \36937 , \36938 , \36939 , \36940 , \36941 , \36942 ,
         \36943 , \36944 , \36945 , \36946 , \36947 , \36948 , \36949 , \36950 , \36951 , \36952 ,
         \36953 , \36954 , \36955 , \36956 , \36957 , \36958 , \36959 , \36960 , \36961 , \36962 ,
         \36963 , \36964 , \36965 , \36966 , \36967 , \36968 , \36969 , \36970 , \36971 , \36972 ,
         \36973 , \36974 , \36975 , \36976 , \36977 , \36978 , \36979 , \36980 , \36981 , \36982 ,
         \36983 , \36984 , \36985 , \36986 , \36987 , \36988 , \36989 , \36990 , \36991 , \36992 ,
         \36993 , \36994 , \36995 , \36996 , \36997 , \36998 , \36999 , \37000 , \37001 , \37002 ,
         \37003 , \37004 , \37005 , \37006 , \37007 , \37008 , \37009 , \37010 , \37011 , \37012 ,
         \37013 , \37014 , \37015 , \37016 , \37017 , \37018 , \37019 , \37020 , \37021 , \37022 ,
         \37023 , \37024 , \37025 , \37026 , \37027 , \37028 , \37029 , \37030 , \37031 , \37032 ,
         \37033 , \37034 , \37035 , \37036 , \37037 , \37038 , \37039 , \37040 , \37041 , \37042 ,
         \37043 , \37044 , \37045 , \37046 , \37047 , \37048 , \37049 , \37050 , \37051 , \37052 ,
         \37053 , \37054 , \37055 , \37056 , \37057 , \37058 , \37059 , \37060 , \37061 , \37062 ,
         \37063 , \37064 , \37065 , \37066 , \37067 , \37068 , \37069 , \37070 , \37071 , \37072 ,
         \37073 , \37074 , \37075 , \37076 , \37077 , \37078 , \37079 , \37080 , \37081 , \37082 ,
         \37083 , \37084 , \37085 , \37086 , \37087 , \37088 , \37089 , \37090 , \37091 , \37092 ,
         \37093 , \37094 , \37095 , \37096 , \37097 , \37098 , \37099 , \37100 , \37101 , \37102 ,
         \37103 , \37104 , \37105 , \37106 , \37107 , \37108 , \37109 , \37110 , \37111 , \37112 ,
         \37113 , \37114 , \37115 , \37116 , \37117 , \37118 , \37119 , \37120 , \37121 , \37122 ,
         \37123 , \37124 , \37125 , \37126 , \37127 , \37128 , \37129 , \37130 , \37131 , \37132 ,
         \37133 , \37134 , \37135 , \37136 , \37137 , \37138 , \37139 , \37140 , \37141 , \37142 ,
         \37143 , \37144 , \37145 , \37146 , \37147 , \37148 , \37149 , \37150 , \37151 , \37152 ,
         \37153 , \37154 , \37155 , \37156 , \37157 , \37158 , \37159 , \37160 , \37161 , \37162 ,
         \37163 , \37164 , \37165 , \37166 , \37167 , \37168 , \37169 , \37170 , \37171 , \37172 ,
         \37173 , \37174 , \37175 , \37176 , \37177 , \37178 , \37179 , \37180 , \37181 , \37182 ,
         \37183 , \37184 , \37185 , \37186 , \37187 , \37188 , \37189 , \37190 , \37191 , \37192 ,
         \37193 , \37194 , \37195 , \37196 , \37197 , \37198 , \37199 , \37200 , \37201 , \37202 ,
         \37203 , \37204 , \37205 , \37206 , \37207 , \37208 , \37209 , \37210 , \37211 , \37212 ,
         \37213 , \37214 , \37215 , \37216 , \37217 , \37218 , \37219 , \37220 , \37221 , \37222 ,
         \37223 , \37224 , \37225 , \37226 , \37227 , \37228 , \37229 , \37230 , \37231 , \37232 ,
         \37233 , \37234 , \37235 , \37236 , \37237 , \37238 , \37239 , \37240 , \37241 , \37242 ,
         \37243 , \37244 , \37245 , \37246 , \37247 , \37248 , \37249 , \37250 , \37251 , \37252 ,
         \37253 , \37254 , \37255 , \37256 , \37257 , \37258 , \37259 , \37260 , \37261 , \37262 ,
         \37263 , \37264 , \37265 , \37266 , \37267 , \37268 , \37269 , \37270 , \37271 , \37272 ,
         \37273 , \37274 , \37275 , \37276 , \37277 , \37278 , \37279 , \37280 , \37281 , \37282 ,
         \37283 , \37284 , \37285 , \37286 , \37287 , \37288 , \37289 , \37290 , \37291 , \37292 ,
         \37293 , \37294 , \37295 , \37296 , \37297 , \37298 , \37299 , \37300 , \37301 , \37302 ,
         \37303 , \37304 , \37305 , \37306 , \37307 , \37308 , \37309 , \37310 , \37311 , \37312 ,
         \37313 , \37314 , \37315 , \37316 , \37317 , \37318 , \37319 , \37320 , \37321 , \37322 ,
         \37323 , \37324 , \37325 , \37326 , \37327 , \37328 , \37329 , \37330 , \37331 , \37332 ,
         \37333 , \37334 , \37335 , \37336 , \37337 , \37338 , \37339 , \37340 , \37341 , \37342 ,
         \37343 , \37344 , \37345 , \37346 , \37347 , \37348 , \37349 , \37350 , \37351 , \37352 ,
         \37353 , \37354 , \37355 , \37356 , \37357 , \37358 , \37359 , \37360 , \37361 , \37362 ,
         \37363 , \37364 , \37365 , \37366 , \37367 , \37368 , \37369 , \37370 , \37371 , \37372 ,
         \37373 , \37374 , \37375 , \37376 , \37377 , \37378 , \37379 , \37380 , \37381 , \37382 ,
         \37383 , \37384 , \37385 , \37386 , \37387 , \37388 , \37389 , \37390 , \37391 , \37392 ,
         \37393 , \37394 , \37395 , \37396 , \37397 , \37398 , \37399 , \37400 , \37401 , \37402 ,
         \37403 , \37404 , \37405 , \37406 , \37407 , \37408 , \37409 , \37410 , \37411 , \37412 ,
         \37413 , \37414 , \37415 , \37416 , \37417 , \37418 , \37419 , \37420 , \37421 , \37422 ,
         \37423 , \37424 , \37425 , \37426 , \37427 , \37428 , \37429 , \37430 , \37431 , \37432 ,
         \37433 , \37434 , \37435 , \37436 , \37437 , \37438 , \37439 , \37440 , \37441 , \37442 ,
         \37443 , \37444 , \37445 , \37446 , \37447 , \37448 , \37449 , \37450 , \37451 , \37452 ,
         \37453 , \37454 , \37455 , \37456 , \37457 , \37458 , \37459 , \37460 , \37461 , \37462 ,
         \37463 , \37464 , \37465 , \37466 , \37467 , \37468 , \37469 , \37470 , \37471 , \37472 ,
         \37473 , \37474 , \37475 , \37476 , \37477 , \37478 , \37479 , \37480 , \37481 , \37482 ,
         \37483 , \37484 , \37485 , \37486 , \37487 , \37488 , \37489 , \37490 , \37491 , \37492 ,
         \37493 , \37494 , \37495 , \37496 , \37497 , \37498 , \37499 , \37500 , \37501 , \37502 ,
         \37503 , \37504 , \37505 , \37506 , \37507 , \37508 , \37509 , \37510 , \37511 , \37512 ,
         \37513 , \37514 , \37515 , \37516 , \37517 , \37518 , \37519 , \37520 , \37521 , \37522 ,
         \37523 , \37524 , \37525 , \37526 , \37527 , \37528 , \37529 , \37530 , \37531 , \37532 ,
         \37533 , \37534 , \37535 , \37536 , \37537 , \37538 , \37539 , \37540 , \37541 , \37542 ,
         \37543 , \37544 , \37545 , \37546 , \37547 , \37548 , \37549 , \37550 , \37551 , \37552 ,
         \37553 , \37554 , \37555 , \37556 , \37557 , \37558 , \37559 , \37560 , \37561 , \37562 ,
         \37563 , \37564 , \37565 , \37566 , \37567 , \37568 , \37569 , \37570 , \37571 , \37572 ,
         \37573 , \37574 , \37575 , \37576 , \37577 , \37578 , \37579 , \37580 , \37581 , \37582 ,
         \37583 , \37584 , \37585 , \37586 , \37587 , \37588 , \37589 , \37590 , \37591 , \37592 ,
         \37593 , \37594 , \37595 , \37596 , \37597 , \37598 , \37599 , \37600 , \37601 , \37602 ,
         \37603 , \37604 , \37605 , \37606 , \37607 , \37608 , \37609 , \37610 , \37611 , \37612 ,
         \37613 , \37614 , \37615 , \37616 , \37617 , \37618 , \37619 , \37620 , \37621 , \37622 ,
         \37623 , \37624 , \37625 , \37626 , \37627 , \37628 , \37629 , \37630 , \37631 , \37632 ,
         \37633 , \37634 , \37635 , \37636 , \37637 , \37638 , \37639 , \37640 , \37641 , \37642 ,
         \37643 , \37644 , \37645 , \37646 , \37647 , \37648 , \37649 , \37650 , \37651 , \37652 ,
         \37653 , \37654 , \37655 , \37656 , \37657 , \37658 , \37659 , \37660 , \37661 , \37662 ,
         \37663 , \37664 , \37665 , \37666 , \37667 , \37668 , \37669 , \37670 , \37671 , \37672 ,
         \37673 , \37674 , \37675 , \37676 , \37677 , \37678 , \37679 , \37680 , \37681 , \37682 ,
         \37683 , \37684 , \37685 , \37686 , \37687 , \37688 , \37689 , \37690 , \37691 , \37692 ,
         \37693 , \37694 , \37695 , \37696 , \37697 , \37698 , \37699 , \37700 , \37701 , \37702 ,
         \37703 , \37704 , \37705 , \37706 , \37707 , \37708 , \37709 , \37710 , \37711 , \37712 ,
         \37713 , \37714 , \37715 , \37716 , \37717 , \37718 , \37719 , \37720 , \37721 , \37722 ,
         \37723 , \37724 , \37725 , \37726 , \37727 , \37728 , \37729 , \37730 , \37731 , \37732 ,
         \37733 , \37734 , \37735 , \37736 , \37737 , \37738 , \37739 , \37740 , \37741 , \37742 ,
         \37743 , \37744 , \37745 , \37746 , \37747 , \37748 , \37749 , \37750 , \37751 , \37752 ,
         \37753 , \37754 , \37755 , \37756 , \37757 , \37758 , \37759 , \37760 , \37761 , \37762 ,
         \37763 , \37764 , \37765 , \37766 , \37767 , \37768 , \37769 , \37770 , \37771 , \37772 ,
         \37773 , \37774 , \37775 , \37776 , \37777 , \37778 , \37779 , \37780 , \37781 , \37782 ,
         \37783 , \37784 , \37785 , \37786 , \37787 , \37788 , \37789 , \37790 , \37791 , \37792 ,
         \37793 , \37794 , \37795 , \37796 , \37797 , \37798 , \37799 , \37800 , \37801 , \37802 ,
         \37803 , \37804 , \37805 , \37806 , \37807 , \37808 , \37809 , \37810 , \37811 , \37812 ,
         \37813 , \37814 , \37815 , \37816 , \37817 , \37818 , \37819 , \37820 , \37821 , \37822 ,
         \37823 , \37824 , \37825 , \37826 , \37827 , \37828 , \37829 , \37830 , \37831 , \37832 ,
         \37833 , \37834 , \37835 , \37836 , \37837 , \37838 , \37839 , \37840 , \37841 , \37842 ,
         \37843 , \37844 , \37845 , \37846 , \37847 , \37848 , \37849 , \37850 , \37851 , \37852 ,
         \37853 , \37854 , \37855 , \37856 , \37857 , \37858 , \37859 , \37860 , \37861 , \37862 ,
         \37863 , \37864 , \37865 , \37866 , \37867 , \37868 , \37869 , \37870 , \37871 , \37872 ,
         \37873 , \37874 , \37875 , \37876 , \37877 , \37878 , \37879 , \37880 , \37881 , \37882 ,
         \37883 , \37884 , \37885 , \37886 , \37887 , \37888 , \37889 , \37890 , \37891 , \37892 ,
         \37893 , \37894 , \37895 , \37896 , \37897 , \37898 , \37899 , \37900 , \37901 , \37902 ,
         \37903 , \37904 , \37905 , \37906 , \37907 , \37908 , \37909 , \37910 , \37911 , \37912 ,
         \37913 , \37914 , \37915 , \37916 , \37917 , \37918 , \37919 , \37920 , \37921 , \37922 ,
         \37923 , \37924 , \37925 , \37926 , \37927 , \37928 , \37929 , \37930 , \37931 , \37932 ,
         \37933 , \37934 , \37935 , \37936 , \37937 , \37938 , \37939 , \37940 , \37941 , \37942 ,
         \37943 , \37944 , \37945 , \37946 , \37947 , \37948 , \37949 , \37950 , \37951 , \37952 ,
         \37953 , \37954 , \37955 , \37956 , \37957 , \37958 , \37959 , \37960 , \37961 , \37962 ,
         \37963 , \37964 , \37965 , \37966 , \37967 , \37968 , \37969 , \37970 , \37971 , \37972 ,
         \37973 , \37974 , \37975 , \37976 , \37977 , \37978 , \37979 , \37980 , \37981 , \37982 ,
         \37983 , \37984 , \37985 , \37986 , \37987 , \37988 , \37989 , \37990 , \37991 , \37992 ,
         \37993 , \37994 , \37995 , \37996 , \37997 , \37998 , \37999 , \38000 , \38001 , \38002 ,
         \38003 , \38004 , \38005 , \38006 , \38007 , \38008 , \38009 , \38010 , \38011 , \38012 ,
         \38013 , \38014 , \38015 , \38016 , \38017 , \38018 , \38019 , \38020 , \38021 , \38022 ,
         \38023 , \38024 , \38025 , \38026 , \38027 , \38028 , \38029 , \38030 , \38031 , \38032 ,
         \38033 , \38034 , \38035 , \38036 , \38037 , \38038 , \38039 , \38040 , \38041 , \38042 ,
         \38043 , \38044 , \38045 , \38046 , \38047 , \38048 , \38049 , \38050 , \38051 , \38052 ,
         \38053 , \38054 , \38055 , \38056 , \38057 , \38058 , \38059 , \38060 , \38061 , \38062 ,
         \38063 , \38064 , \38065 , \38066 , \38067 , \38068 , \38069 , \38070 , \38071 , \38072 ,
         \38073 , \38074 , \38075 , \38076 , \38077 , \38078 , \38079 , \38080 , \38081 , \38082 ,
         \38083 , \38084 , \38085 , \38086 , \38087 , \38088 , \38089 , \38090 , \38091 , \38092 ,
         \38093 , \38094 , \38095 , \38096 , \38097 , \38098 , \38099 , \38100 , \38101 , \38102 ,
         \38103 , \38104 , \38105 , \38106 , \38107 , \38108 , \38109 , \38110 , \38111 , \38112 ,
         \38113 , \38114 , \38115 , \38116 , \38117 , \38118 , \38119 , \38120 , \38121 , \38122 ,
         \38123 , \38124 , \38125 , \38126 , \38127 , \38128 , \38129 , \38130 , \38131 , \38132 ,
         \38133 , \38134 , \38135 , \38136 , \38137 , \38138 , \38139 , \38140 , \38141 , \38142 ,
         \38143 , \38144 , \38145 , \38146 , \38147 , \38148 , \38149 , \38150 , \38151 , \38152 ,
         \38153 , \38154 , \38155 , \38156 , \38157 , \38158 , \38159 , \38160 , \38161 , \38162 ,
         \38163 , \38164 , \38165 , \38166 , \38167 , \38168 , \38169 , \38170 , \38171 , \38172 ,
         \38173 , \38174 , \38175 , \38176 , \38177 , \38178 , \38179 , \38180 , \38181 , \38182 ,
         \38183 , \38184 , \38185 , \38186 , \38187 , \38188 , \38189 , \38190 , \38191 , \38192 ,
         \38193 , \38194 , \38195 , \38196 , \38197 , \38198 , \38199 , \38200 , \38201 , \38202 ,
         \38203 , \38204 , \38205 , \38206 , \38207 , \38208 , \38209 , \38210 , \38211 , \38212 ,
         \38213 , \38214 , \38215 , \38216 , \38217 , \38218 , \38219 , \38220 , \38221 , \38222 ,
         \38223 , \38224 , \38225 , \38226 , \38227 , \38228 , \38229 , \38230 , \38231 , \38232 ,
         \38233 , \38234 , \38235 , \38236 , \38237 , \38238 , \38239 , \38240 , \38241 , \38242 ,
         \38243 , \38244 , \38245 , \38246 , \38247 , \38248 , \38249 , \38250 , \38251 , \38252 ,
         \38253 , \38254 , \38255 , \38256 , \38257 , \38258 , \38259 , \38260 , \38261 , \38262 ,
         \38263 , \38264 , \38265 , \38266 , \38267 , \38268 , \38269 , \38270 , \38271 , \38272 ,
         \38273 , \38274 , \38275 , \38276 , \38277 , \38278 , \38279 , \38280 , \38281 , \38282 ,
         \38283 , \38284 , \38285 , \38286 , \38287 , \38288 , \38289 , \38290 , \38291 , \38292 ,
         \38293 , \38294 , \38295 , \38296 , \38297 , \38298 , \38299 , \38300 , \38301 , \38302 ,
         \38303 , \38304 , \38305 , \38306 , \38307 , \38308 , \38309 , \38310 , \38311 , \38312 ,
         \38313 , \38314 , \38315 , \38316 , \38317 , \38318 , \38319 , \38320 , \38321 , \38322 ,
         \38323 , \38324 , \38325 , \38326 , \38327 , \38328 , \38329 , \38330 , \38331 , \38332 ,
         \38333 , \38334 , \38335 , \38336 , \38337 , \38338 , \38339 , \38340 , \38341 , \38342 ,
         \38343 , \38344 , \38345 , \38346 , \38347 , \38348 , \38349 , \38350 , \38351 , \38352 ,
         \38353 , \38354 , \38355 , \38356 , \38357 , \38358 , \38359 , \38360 , \38361 , \38362 ,
         \38363 , \38364 , \38365 , \38366 , \38367 , \38368 , \38369 , \38370 , \38371 , \38372 ,
         \38373 , \38374 , \38375 , \38376 , \38377 , \38378 , \38379 , \38380 , \38381 , \38382 ,
         \38383 , \38384 , \38385 , \38386 , \38387 , \38388 , \38389 , \38390 , \38391 , \38392 ,
         \38393 , \38394 , \38395 , \38396 , \38397 , \38398 , \38399 , \38400 , \38401 , \38402 ,
         \38403 , \38404 , \38405 , \38406 , \38407 , \38408 , \38409 , \38410 , \38411 , \38412 ,
         \38413 , \38414 , \38415 , \38416 , \38417 , \38418 , \38419 , \38420 , \38421 , \38422 ,
         \38423 , \38424 , \38425 , \38426 , \38427 , \38428 , \38429 , \38430 , \38431 , \38432 ,
         \38433 , \38434 , \38435 , \38436 , \38437 , \38438 , \38439 , \38440 , \38441 , \38442 ,
         \38443 , \38444 , \38445 , \38446 , \38447 , \38448 , \38449 , \38450 , \38451 , \38452 ,
         \38453 , \38454 , \38455 , \38456 , \38457 , \38458 , \38459 , \38460 , \38461 , \38462 ,
         \38463 , \38464 , \38465 , \38466 , \38467 , \38468 , \38469 , \38470 , \38471 , \38472 ,
         \38473 , \38474 , \38475 , \38476 , \38477 , \38478 , \38479 , \38480 , \38481 , \38482 ,
         \38483 , \38484 , \38485 , \38486 , \38487 , \38488 , \38489 , \38490 , \38491 , \38492 ,
         \38493 , \38494 , \38495 , \38496 , \38497 , \38498 , \38499 , \38500 , \38501 , \38502 ,
         \38503 , \38504 , \38505 , \38506 , \38507 , \38508 , \38509 , \38510 , \38511 , \38512 ,
         \38513 , \38514 , \38515 , \38516 , \38517 , \38518 , \38519 , \38520 , \38521 , \38522 ,
         \38523 , \38524 , \38525 , \38526 , \38527 , \38528 , \38529 , \38530 , \38531 , \38532 ,
         \38533 , \38534 , \38535 , \38536 , \38537 , \38538 , \38539 , \38540 , \38541 , \38542 ,
         \38543 , \38544 , \38545 , \38546 , \38547 , \38548 , \38549 , \38550 , \38551 , \38552 ,
         \38553 , \38554 , \38555 , \38556 , \38557 , \38558 , \38559 , \38560 , \38561 , \38562 ,
         \38563 , \38564 , \38565 , \38566 , \38567 , \38568 , \38569 , \38570 , \38571 , \38572 ,
         \38573 , \38574 , \38575 , \38576 , \38577 , \38578 , \38579 , \38580 , \38581 , \38582 ,
         \38583 , \38584 , \38585 , \38586 , \38587 , \38588 , \38589 , \38590 , \38591 , \38592 ,
         \38593 , \38594 , \38595 , \38596 , \38597 , \38598 , \38599 , \38600 , \38601 , \38602 ,
         \38603 , \38604 , \38605 , \38606 , \38607 , \38608 , \38609 , \38610 , \38611 , \38612 ,
         \38613 , \38614 , \38615 , \38616 , \38617 , \38618 , \38619 , \38620 , \38621 , \38622 ,
         \38623 , \38624 , \38625 , \38626 , \38627 , \38628 , \38629 , \38630 , \38631 , \38632 ,
         \38633 , \38634 , \38635 , \38636 , \38637 , \38638 , \38639 , \38640 , \38641 , \38642 ,
         \38643 , \38644 , \38645 , \38646 , \38647 , \38648 , \38649 , \38650 , \38651 , \38652 ,
         \38653 , \38654 , \38655 , \38656 , \38657 , \38658 , \38659 , \38660 , \38661 , \38662 ,
         \38663 , \38664 , \38665 , \38666 , \38667 , \38668 , \38669 , \38670 , \38671 , \38672 ,
         \38673 , \38674 , \38675 , \38676 , \38677 , \38678 , \38679 , \38680 , \38681 , \38682 ,
         \38683 , \38684 , \38685 , \38686 , \38687 , \38688 , \38689 , \38690 , \38691 , \38692 ,
         \38693 , \38694 , \38695 , \38696 , \38697 , \38698 , \38699 , \38700 , \38701 , \38702 ,
         \38703 , \38704 , \38705 , \38706 , \38707 , \38708 , \38709 , \38710 , \38711 , \38712 ,
         \38713 , \38714 , \38715 , \38716 , \38717 , \38718 , \38719 , \38720 , \38721 , \38722 ,
         \38723 , \38724 , \38725 , \38726 , \38727 , \38728 , \38729 , \38730 , \38731 , \38732 ,
         \38733 , \38734 , \38735 , \38736 , \38737 , \38738 , \38739 , \38740 , \38741 , \38742 ,
         \38743 , \38744 , \38745 , \38746 , \38747 , \38748 , \38749 , \38750 , \38751 , \38752 ,
         \38753 , \38754 , \38755 , \38756 , \38757 , \38758 , \38759 , \38760 , \38761 , \38762 ,
         \38763 , \38764 , \38765 , \38766 , \38767 , \38768 , \38769 , \38770 , \38771 , \38772 ,
         \38773 , \38774 , \38775 , \38776 , \38777 , \38778 , \38779 , \38780 , \38781 , \38782 ,
         \38783 , \38784 , \38785 , \38786 , \38787 , \38788 , \38789 , \38790 , \38791 , \38792 ,
         \38793 , \38794 , \38795 , \38796 , \38797 , \38798 , \38799 , \38800 , \38801 , \38802 ,
         \38803 , \38804 , \38805 , \38806 , \38807 , \38808 , \38809 , \38810 , \38811 , \38812 ,
         \38813 , \38814 , \38815 , \38816 , \38817 , \38818 , \38819 , \38820 , \38821 , \38822 ,
         \38823 , \38824 , \38825 , \38826 , \38827 , \38828 , \38829 , \38830 , \38831 , \38832 ,
         \38833 , \38834 , \38835 , \38836 , \38837 , \38838 , \38839 , \38840 , \38841 , \38842 ,
         \38843 , \38844 , \38845 , \38846 , \38847 , \38848 , \38849 , \38850 , \38851 , \38852 ,
         \38853 , \38854 , \38855 , \38856 , \38857 , \38858 , \38859 , \38860 , \38861 , \38862 ,
         \38863 , \38864 , \38865 , \38866 , \38867 , \38868 , \38869 , \38870 , \38871 , \38872 ,
         \38873 , \38874 , \38875 , \38876 , \38877 , \38878 , \38879 , \38880 , \38881 , \38882 ,
         \38883 , \38884 , \38885 , \38886 , \38887 , \38888 , \38889 , \38890 , \38891 , \38892 ,
         \38893 , \38894 , \38895 , \38896 , \38897 , \38898 , \38899 , \38900 , \38901 , \38902 ,
         \38903 , \38904 , \38905 , \38906 , \38907 , \38908 , \38909 , \38910 , \38911 , \38912 ,
         \38913 , \38914 , \38915 , \38916 , \38917 , \38918 , \38919 , \38920 , \38921 , \38922 ,
         \38923 , \38924 , \38925 , \38926 , \38927 , \38928 , \38929 , \38930 , \38931 , \38932 ,
         \38933 , \38934 , \38935 , \38936 , \38937 , \38938 , \38939 , \38940 , \38941 , \38942 ,
         \38943 , \38944 , \38945 , \38946 , \38947 , \38948 , \38949 , \38950 , \38951 , \38952 ,
         \38953 , \38954 , \38955 , \38956 , \38957 , \38958 , \38959 , \38960 , \38961 , \38962 ,
         \38963 , \38964 , \38965 , \38966 , \38967 , \38968 , \38969 , \38970 , \38971 , \38972 ,
         \38973 , \38974 , \38975 , \38976 , \38977 , \38978 , \38979 , \38980 , \38981 , \38982 ,
         \38983 , \38984 , \38985 , \38986 , \38987 , \38988 , \38989 , \38990 , \38991 , \38992 ,
         \38993 , \38994 , \38995 , \38996 , \38997 , \38998 , \38999 , \39000 , \39001 , \39002 ,
         \39003 , \39004 , \39005 , \39006 , \39007 , \39008 , \39009 , \39010 , \39011 , \39012 ,
         \39013 , \39014 , \39015 , \39016 , \39017 , \39018 , \39019 , \39020 , \39021 , \39022 ,
         \39023 , \39024 , \39025 , \39026 , \39027 , \39028 , \39029 , \39030 , \39031 , \39032 ,
         \39033 , \39034 , \39035 , \39036 , \39037 , \39038 , \39039 , \39040 , \39041 , \39042 ,
         \39043 , \39044 , \39045 , \39046 , \39047 , \39048 , \39049 , \39050 , \39051 , \39052 ,
         \39053 , \39054 , \39055 , \39056 , \39057 , \39058 , \39059 , \39060 , \39061 , \39062 ,
         \39063 , \39064 , \39065 , \39066 , \39067 , \39068 , \39069 , \39070 , \39071 , \39072 ,
         \39073 , \39074 , \39075 , \39076 , \39077 , \39078 , \39079 , \39080 , \39081 , \39082 ,
         \39083 , \39084 , \39085 , \39086 , \39087 , \39088 , \39089 , \39090 , \39091 , \39092 ,
         \39093 , \39094 , \39095 , \39096 , \39097 , \39098 , \39099 , \39100 , \39101 , \39102 ,
         \39103 , \39104 , \39105 , \39106 , \39107 , \39108 , \39109 , \39110 , \39111 , \39112 ,
         \39113 , \39114 , \39115 , \39116 , \39117 , \39118 , \39119 , \39120 , \39121 , \39122 ,
         \39123 , \39124 , \39125 , \39126 , \39127 , \39128 , \39129 , \39130 , \39131 , \39132 ,
         \39133 , \39134 , \39135 , \39136 , \39137 , \39138 , \39139 , \39140 , \39141 , \39142 ,
         \39143 , \39144 , \39145 , \39146 , \39147 , \39148 , \39149 , \39150 , \39151 , \39152 ,
         \39153 , \39154 , \39155 , \39156 , \39157 , \39158 , \39159 , \39160 , \39161 , \39162 ,
         \39163 , \39164 , \39165 , \39166 , \39167 , \39168 , \39169 , \39170 , \39171 , \39172 ,
         \39173 , \39174 , \39175 , \39176 , \39177 , \39178 , \39179 , \39180 , \39181 , \39182 ,
         \39183 , \39184 , \39185 , \39186 , \39187 , \39188 , \39189 , \39190 , \39191 , \39192 ,
         \39193 , \39194 , \39195 , \39196 , \39197 , \39198 , \39199 , \39200 , \39201 , \39202 ,
         \39203 , \39204 , \39205 , \39206 , \39207 , \39208 , \39209 , \39210 , \39211 , \39212 ,
         \39213 , \39214 , \39215 , \39216 , \39217 , \39218 , \39219 , \39220 , \39221 , \39222 ,
         \39223 , \39224 , \39225 , \39226 , \39227 , \39228 , \39229 , \39230 , \39231 , \39232 ,
         \39233 , \39234 , \39235 , \39236 , \39237 , \39238 , \39239 , \39240 , \39241 , \39242 ,
         \39243 , \39244 , \39245 , \39246 , \39247 , \39248 , \39249 , \39250 , \39251 , \39252 ,
         \39253 , \39254 , \39255 , \39256 , \39257 , \39258 , \39259 , \39260 , \39261 , \39262 ,
         \39263 , \39264 , \39265 , \39266 , \39267 , \39268 , \39269 , \39270 , \39271 , \39272 ,
         \39273 , \39274 , \39275 , \39276 , \39277 , \39278 , \39279 , \39280 , \39281 , \39282 ,
         \39283 , \39284 , \39285 , \39286 , \39287 , \39288 , \39289 , \39290 , \39291 , \39292 ,
         \39293 , \39294 , \39295 , \39296 , \39297 , \39298 , \39299 , \39300 , \39301 , \39302 ,
         \39303 , \39304 , \39305 , \39306 , \39307 , \39308 , \39309 , \39310 , \39311 , \39312 ,
         \39313 , \39314 , \39315 , \39316 , \39317 , \39318 , \39319 , \39320 , \39321 , \39322 ,
         \39323 , \39324 , \39325 , \39326 , \39327 , \39328 , \39329 , \39330 , \39331 , \39332 ,
         \39333 , \39334 , \39335 , \39336 , \39337 , \39338 , \39339 , \39340 , \39341 , \39342 ,
         \39343 , \39344 , \39345 , \39346 , \39347 , \39348 , \39349 , \39350 , \39351 , \39352 ,
         \39353 , \39354 , \39355 , \39356 , \39357 , \39358 , \39359 , \39360 , \39361 , \39362 ,
         \39363 , \39364 , \39365 , \39366 , \39367 , \39368 , \39369 , \39370 , \39371 , \39372 ,
         \39373 , \39374 , \39375 , \39376 , \39377 , \39378 , \39379 , \39380 , \39381 , \39382 ,
         \39383 , \39384 , \39385 , \39386 , \39387 , \39388 , \39389 , \39390 , \39391 , \39392 ,
         \39393 , \39394 , \39395 , \39396 , \39397 , \39398 , \39399 , \39400 , \39401 , \39402 ,
         \39403 , \39404 , \39405 , \39406 , \39407 , \39408 , \39409 , \39410 , \39411 , \39412 ,
         \39413 , \39414 , \39415 , \39416 , \39417 , \39418 , \39419 , \39420 , \39421 , \39422 ,
         \39423 , \39424 , \39425 , \39426 , \39427 , \39428 , \39429 , \39430 , \39431 , \39432 ,
         \39433 , \39434 , \39435 , \39436 , \39437 , \39438 , \39439 , \39440 , \39441 , \39442 ,
         \39443 , \39444 , \39445 , \39446 , \39447 , \39448 , \39449 , \39450 , \39451 , \39452 ,
         \39453 , \39454 , \39455 , \39456 , \39457 , \39458 , \39459 , \39460 , \39461 , \39462 ,
         \39463 , \39464 , \39465 , \39466 , \39467 , \39468 , \39469 , \39470 , \39471 , \39472 ,
         \39473 , \39474 , \39475 , \39476 , \39477 , \39478 , \39479 , \39480 , \39481 , \39482 ,
         \39483 , \39484 , \39485 , \39486 , \39487 , \39488 , \39489 , \39490 , \39491 , \39492 ,
         \39493 , \39494 , \39495 , \39496 , \39497 , \39498 , \39499 , \39500 , \39501 , \39502 ,
         \39503 , \39504 , \39505 , \39506 , \39507 , \39508 , \39509 , \39510 , \39511 , \39512 ,
         \39513 , \39514 , \39515 , \39516 , \39517 , \39518 , \39519 , \39520 , \39521 , \39522 ,
         \39523 , \39524 , \39525 , \39526 , \39527 , \39528 , \39529 , \39530 , \39531 , \39532 ,
         \39533 , \39534 , \39535 , \39536 , \39537 , \39538 , \39539 , \39540 , \39541 , \39542 ,
         \39543 , \39544 , \39545 , \39546 , \39547 , \39548 , \39549 , \39550 , \39551 , \39552 ,
         \39553 , \39554 , \39555 , \39556 , \39557 , \39558 , \39559 , \39560 , \39561 , \39562 ,
         \39563 , \39564 , \39565 , \39566 , \39567 , \39568 , \39569 , \39570 , \39571 , \39572 ,
         \39573 , \39574 , \39575 , \39576 , \39577 , \39578 , \39579 , \39580 , \39581 , \39582 ,
         \39583 , \39584 , \39585 , \39586 , \39587 , \39588 , \39589 , \39590 , \39591 , \39592 ,
         \39593 , \39594 , \39595 , \39596 , \39597 , \39598 , \39599 , \39600 , \39601 , \39602 ,
         \39603 , \39604 , \39605 , \39606 , \39607 , \39608 , \39609 , \39610 , \39611 , \39612 ,
         \39613 , \39614 , \39615 , \39616 , \39617 , \39618 , \39619 , \39620 , \39621 , \39622 ,
         \39623 , \39624 , \39625 , \39626 , \39627 , \39628 , \39629 , \39630 , \39631 , \39632 ,
         \39633 , \39634 , \39635 , \39636 , \39637 , \39638 , \39639 , \39640 , \39641 , \39642 ,
         \39643 , \39644 , \39645 , \39646 , \39647 , \39648 , \39649 , \39650 , \39651 , \39652 ,
         \39653 , \39654 , \39655 , \39656 , \39657 , \39658 , \39659 , \39660 , \39661 , \39662 ,
         \39663 , \39664 , \39665 , \39666 , \39667 , \39668 , \39669 , \39670 , \39671 , \39672 ,
         \39673 , \39674 , \39675 , \39676 , \39677 , \39678 , \39679 , \39680 , \39681 , \39682 ,
         \39683 , \39684 , \39685 , \39686 , \39687 , \39688 , \39689 , \39690 , \39691 , \39692 ,
         \39693 , \39694 , \39695 , \39696 , \39697 , \39698 , \39699 , \39700 , \39701 , \39702 ,
         \39703 , \39704 , \39705 , \39706 , \39707 , \39708 , \39709 , \39710 , \39711 , \39712 ,
         \39713 , \39714 , \39715 , \39716 , \39717 , \39718 , \39719 , \39720 , \39721 , \39722 ,
         \39723 , \39724 , \39725 , \39726 , \39727 , \39728 , \39729 , \39730 , \39731 , \39732 ,
         \39733 , \39734 , \39735 , \39736 , \39737 , \39738 , \39739 , \39740 , \39741 , \39742 ,
         \39743 , \39744 , \39745 , \39746 , \39747 , \39748 , \39749 , \39750 , \39751 , \39752 ,
         \39753 , \39754 , \39755 , \39756 , \39757 , \39758 , \39759 , \39760 , \39761 , \39762 ,
         \39763 , \39764 , \39765 , \39766 , \39767 , \39768 , \39769 , \39770 , \39771 , \39772 ,
         \39773 , \39774 , \39775 , \39776 , \39777 , \39778 , \39779 , \39780 , \39781 , \39782 ,
         \39783 , \39784 , \39785 , \39786 , \39787 , \39788 , \39789 , \39790 , \39791 , \39792 ,
         \39793 , \39794 , \39795 , \39796 , \39797 , \39798 , \39799 , \39800 , \39801 , \39802 ,
         \39803 , \39804 , \39805 , \39806 , \39807 , \39808 , \39809 , \39810 , \39811 , \39812 ,
         \39813 , \39814 , \39815 , \39816 , \39817 , \39818 , \39819 , \39820 , \39821 , \39822 ,
         \39823 , \39824 , \39825 , \39826 , \39827 , \39828 , \39829 , \39830 , \39831 , \39832 ,
         \39833 , \39834 , \39835 , \39836 , \39837 , \39838 , \39839 , \39840 , \39841 , \39842 ,
         \39843 , \39844 , \39845 , \39846 , \39847 , \39848 , \39849 , \39850 , \39851 , \39852 ,
         \39853 , \39854 , \39855 , \39856 , \39857 , \39858 , \39859 , \39860 , \39861 , \39862 ,
         \39863 , \39864 , \39865 , \39866 , \39867 , \39868 , \39869 , \39870 , \39871 , \39872 ,
         \39873 , \39874 , \39875 , \39876 , \39877 , \39878 , \39879 , \39880 , \39881 , \39882 ,
         \39883 , \39884 , \39885 , \39886 , \39887 , \39888 , \39889 , \39890 , \39891 , \39892 ,
         \39893 , \39894 , \39895 , \39896 , \39897 , \39898 , \39899 , \39900 , \39901 , \39902 ,
         \39903 , \39904 , \39905 , \39906 , \39907 , \39908 , \39909 , \39910 , \39911 , \39912 ,
         \39913 , \39914 , \39915 , \39916 , \39917 , \39918 , \39919 , \39920 , \39921 , \39922 ,
         \39923 , \39924 , \39925 , \39926 , \39927 , \39928 , \39929 , \39930 , \39931 , \39932 ,
         \39933 , \39934 , \39935 , \39936 , \39937 , \39938 , \39939 , \39940 , \39941 , \39942 ,
         \39943 , \39944 , \39945 , \39946 , \39947 , \39948 , \39949 , \39950 , \39951 , \39952 ,
         \39953 , \39954 , \39955 , \39956 , \39957 , \39958 , \39959 , \39960 , \39961 , \39962 ,
         \39963 , \39964 , \39965 , \39966 , \39967 , \39968 , \39969 , \39970 , \39971 , \39972 ,
         \39973 , \39974 , \39975 , \39976 , \39977 , \39978 , \39979 , \39980 , \39981 , \39982 ,
         \39983 , \39984 , \39985 , \39986 , \39987 , \39988 , \39989 , \39990 , \39991 , \39992 ,
         \39993 , \39994 , \39995 , \39996 , \39997 , \39998 , \39999 , \40000 , \40001 , \40002 ,
         \40003 , \40004 , \40005 , \40006 , \40007 , \40008 , \40009 , \40010 , \40011 , \40012 ,
         \40013 , \40014 , \40015 , \40016 , \40017 , \40018 , \40019 , \40020 , \40021 , \40022 ,
         \40023 , \40024 , \40025 , \40026 , \40027 , \40028 , \40029 , \40030 , \40031 , \40032 ,
         \40033 , \40034 , \40035 , \40036 , \40037 , \40038 , \40039 , \40040 , \40041 , \40042 ,
         \40043 , \40044 , \40045 , \40046 , \40047 , \40048 , \40049 , \40050 , \40051 , \40052 ,
         \40053 , \40054 , \40055 , \40056 , \40057 , \40058 , \40059 , \40060 , \40061 , \40062 ,
         \40063 , \40064 , \40065 , \40066 , \40067 , \40068 , \40069 , \40070 , \40071 , \40072 ,
         \40073 , \40074 , \40075 , \40076 , \40077 , \40078 , \40079 , \40080 , \40081 , \40082 ,
         \40083 , \40084 , \40085 , \40086 , \40087 , \40088 , \40089 , \40090 , \40091 , \40092 ,
         \40093 , \40094 , \40095 , \40096 , \40097 , \40098 , \40099 , \40100 , \40101 , \40102 ,
         \40103 , \40104 , \40105 , \40106 , \40107 , \40108 , \40109 , \40110 , \40111 , \40112 ,
         \40113 , \40114 , \40115 , \40116 , \40117 , \40118 , \40119 , \40120 , \40121 , \40122 ,
         \40123 , \40124 , \40125 , \40126 , \40127 , \40128 , \40129 , \40130 , \40131 , \40132 ,
         \40133 , \40134 , \40135 , \40136 , \40137 , \40138 , \40139 , \40140 , \40141 , \40142 ,
         \40143 , \40144 , \40145 , \40146 , \40147 , \40148 , \40149 , \40150 , \40151 , \40152 ,
         \40153 , \40154 , \40155 , \40156 , \40157 , \40158 , \40159 , \40160 , \40161 , \40162 ,
         \40163 , \40164 , \40165 , \40166 , \40167 , \40168 , \40169 , \40170 , \40171 , \40172 ,
         \40173 , \40174 , \40175 , \40176 , \40177 , \40178 , \40179 , \40180 , \40181 , \40182 ,
         \40183 , \40184 , \40185 , \40186 , \40187 , \40188 , \40189 , \40190 , \40191 , \40192 ,
         \40193 , \40194 , \40195 , \40196 , \40197 , \40198 , \40199 , \40200 , \40201 , \40202 ,
         \40203 , \40204 , \40205 , \40206 , \40207 , \40208 , \40209 , \40210 , \40211 , \40212 ,
         \40213 , \40214 , \40215 , \40216 , \40217 , \40218 , \40219 , \40220 , \40221 , \40222 ,
         \40223 , \40224 , \40225 , \40226 , \40227 , \40228 , \40229 , \40230 , \40231 , \40232 ,
         \40233 , \40234 , \40235 , \40236 , \40237 , \40238 , \40239 , \40240 , \40241 , \40242 ,
         \40243 , \40244 , \40245 , \40246 , \40247 , \40248 , \40249 , \40250 , \40251 , \40252 ,
         \40253 , \40254 , \40255 , \40256 , \40257 , \40258 , \40259 , \40260 , \40261 , \40262 ,
         \40263 , \40264 , \40265 , \40266 , \40267 , \40268 , \40269 , \40270 , \40271 , \40272 ,
         \40273 , \40274 , \40275 , \40276 , \40277 , \40278 , \40279 , \40280 , \40281 , \40282 ,
         \40283 , \40284 , \40285 , \40286 , \40287 , \40288 , \40289 , \40290 , \40291 , \40292 ,
         \40293 , \40294 , \40295 , \40296 , \40297 , \40298 , \40299 , \40300 , \40301 , \40302 ,
         \40303 , \40304 , \40305 , \40306 , \40307 , \40308 , \40309 , \40310 , \40311 , \40312 ,
         \40313 , \40314 , \40315 , \40316 , \40317 , \40318 , \40319 , \40320 , \40321 , \40322 ,
         \40323 , \40324 , \40325 , \40326 , \40327 , \40328 , \40329 , \40330 , \40331 , \40332 ,
         \40333 , \40334 , \40335 , \40336 , \40337 , \40338 , \40339 , \40340 , \40341 , \40342 ,
         \40343 , \40344 , \40345 , \40346 , \40347 , \40348 , \40349 , \40350 , \40351 , \40352 ,
         \40353 , \40354 , \40355 , \40356 , \40357 , \40358 , \40359 , \40360 , \40361 , \40362 ,
         \40363 , \40364 , \40365 , \40366 , \40367 , \40368 , \40369 , \40370 , \40371 , \40372 ,
         \40373 , \40374 , \40375 , \40376 , \40377 , \40378 , \40379 , \40380 , \40381 , \40382 ,
         \40383 , \40384 , \40385 , \40386 , \40387 , \40388 , \40389 , \40390 , \40391 , \40392 ,
         \40393 , \40394 , \40395 , \40396 , \40397 , \40398 , \40399 , \40400 , \40401 , \40402 ,
         \40403 , \40404 , \40405 , \40406 , \40407 , \40408 , \40409 , \40410 , \40411 , \40412 ,
         \40413 , \40414 , \40415 , \40416 , \40417 , \40418 , \40419 , \40420 , \40421 , \40422 ,
         \40423 , \40424 , \40425 , \40426 , \40427 , \40428 , \40429 , \40430 , \40431 , \40432 ,
         \40433 , \40434 , \40435 , \40436 , \40437 , \40438 , \40439 , \40440 , \40441 , \40442 ,
         \40443 , \40444 , \40445 , \40446 , \40447 , \40448 , \40449 , \40450 , \40451 , \40452 ,
         \40453 , \40454 , \40455 , \40456 , \40457 , \40458 , \40459 , \40460 , \40461 , \40462 ,
         \40463 , \40464 , \40465 , \40466 , \40467 , \40468 , \40469 , \40470 , \40471 , \40472 ,
         \40473 , \40474 , \40475 , \40476 , \40477 , \40478 , \40479 , \40480 , \40481 , \40482 ,
         \40483 , \40484 , \40485 , \40486 , \40487 , \40488 , \40489 , \40490 , \40491 , \40492 ,
         \40493 , \40494 , \40495 , \40496 , \40497 , \40498 , \40499 , \40500 , \40501 , \40502 ,
         \40503 , \40504 , \40505 , \40506 , \40507 , \40508 , \40509 , \40510 , \40511 , \40512 ,
         \40513 , \40514 , \40515 , \40516 , \40517 , \40518 , \40519 , \40520 , \40521 , \40522 ,
         \40523 , \40524 , \40525 , \40526 , \40527 , \40528 , \40529 , \40530 , \40531 , \40532 ,
         \40533 , \40534 , \40535 , \40536 , \40537 , \40538 , \40539 , \40540 , \40541 , \40542 ,
         \40543 , \40544 , \40545 , \40546 , \40547 , \40548 , \40549 , \40550 , \40551 , \40552 ,
         \40553 , \40554 , \40555 , \40556 , \40557 , \40558 , \40559 , \40560 , \40561 , \40562 ,
         \40563 , \40564 , \40565 , \40566 , \40567 , \40568 , \40569 , \40570 , \40571 , \40572 ,
         \40573 , \40574 , \40575 , \40576 , \40577 , \40578 , \40579 , \40580 , \40581 , \40582 ,
         \40583 , \40584 , \40585 , \40586 , \40587 , \40588 , \40589 , \40590 , \40591 , \40592 ,
         \40593 , \40594 , \40595 , \40596 , \40597 , \40598 , \40599 , \40600 , \40601 , \40602 ,
         \40603 , \40604 , \40605 , \40606 , \40607 , \40608 , \40609 , \40610 , \40611 , \40612 ,
         \40613 , \40614 , \40615 , \40616 , \40617 , \40618 , \40619 , \40620 , \40621 , \40622 ,
         \40623 , \40624 , \40625 , \40626 , \40627 , \40628 , \40629 , \40630 , \40631 , \40632 ,
         \40633 , \40634 , \40635 , \40636 , \40637 , \40638 , \40639 , \40640 , \40641 , \40642 ,
         \40643 , \40644 , \40645 , \40646 , \40647 , \40648 , \40649 , \40650 , \40651 , \40652 ,
         \40653 , \40654 , \40655 , \40656 , \40657 , \40658 , \40659 , \40660 , \40661 , \40662 ,
         \40663 , \40664 , \40665 , \40666 , \40667 , \40668 , \40669 , \40670 , \40671 , \40672 ,
         \40673 , \40674 , \40675 , \40676 , \40677 , \40678 , \40679 , \40680 , \40681 , \40682 ,
         \40683 , \40684 , \40685 , \40686 , \40687 , \40688 , \40689 , \40690 , \40691 , \40692 ,
         \40693 , \40694 , \40695 , \40696 , \40697 , \40698 , \40699 , \40700 , \40701 , \40702 ,
         \40703 , \40704 , \40705 , \40706 , \40707 , \40708 , \40709 , \40710 , \40711 , \40712 ,
         \40713 , \40714 , \40715 , \40716 , \40717 , \40718 , \40719 , \40720 , \40721 , \40722 ,
         \40723 , \40724 , \40725 , \40726 , \40727 , \40728 , \40729 , \40730 , \40731 , \40732 ,
         \40733 , \40734 , \40735 , \40736 , \40737 , \40738 , \40739 , \40740 , \40741 , \40742 ,
         \40743 , \40744 , \40745 , \40746 , \40747 , \40748 , \40749 , \40750 , \40751 , \40752 ,
         \40753 , \40754 , \40755 , \40756 , \40757 , \40758 , \40759 , \40760 , \40761 , \40762 ,
         \40763 , \40764 , \40765 , \40766 , \40767 , \40768 , \40769 , \40770 , \40771 , \40772 ,
         \40773 , \40774 , \40775 , \40776 , \40777 , \40778 , \40779 , \40780 , \40781 , \40782 ,
         \40783 , \40784 , \40785 , \40786 , \40787 , \40788 , \40789 , \40790 , \40791 , \40792 ,
         \40793 , \40794 , \40795 , \40796 , \40797 , \40798 , \40799 , \40800 , \40801 , \40802 ,
         \40803 , \40804 , \40805 , \40806 , \40807 , \40808 , \40809 , \40810 , \40811 , \40812 ,
         \40813 , \40814 , \40815 , \40816 , \40817 , \40818 , \40819 , \40820 , \40821 , \40822 ,
         \40823 , \40824 , \40825 , \40826 , \40827 , \40828 , \40829 , \40830 , \40831 , \40832 ,
         \40833 , \40834 , \40835 , \40836 , \40837 , \40838 , \40839 , \40840 , \40841 , \40842 ,
         \40843 , \40844 , \40845 , \40846 , \40847 , \40848 , \40849 , \40850 , \40851 , \40852 ,
         \40853 , \40854 , \40855 , \40856 , \40857 , \40858 , \40859 , \40860 , \40861 , \40862 ,
         \40863 , \40864 , \40865 , \40866 , \40867 , \40868 , \40869 , \40870 , \40871 , \40872 ,
         \40873 , \40874 , \40875 , \40876 , \40877 , \40878 , \40879 , \40880 , \40881 , \40882 ,
         \40883 , \40884 , \40885 , \40886 , \40887 , \40888 , \40889 , \40890 , \40891 , \40892 ,
         \40893 , \40894 , \40895 , \40896 , \40897 , \40898 , \40899 , \40900 , \40901 , \40902 ,
         \40903 , \40904 , \40905 , \40906 , \40907 , \40908 , \40909 , \40910 , \40911 , \40912 ,
         \40913 , \40914 , \40915 , \40916 , \40917 , \40918 , \40919 , \40920 , \40921 , \40922 ,
         \40923 , \40924 , \40925 , \40926 , \40927 , \40928 , \40929 , \40930 , \40931 , \40932 ,
         \40933 , \40934 , \40935 , \40936 , \40937 , \40938 , \40939 , \40940 , \40941 , \40942 ,
         \40943 , \40944 , \40945 , \40946 , \40947 , \40948 , \40949 , \40950 , \40951 , \40952 ,
         \40953 , \40954 , \40955 , \40956 , \40957 , \40958 , \40959 , \40960 , \40961 , \40962 ,
         \40963 , \40964 , \40965 , \40966 , \40967 , \40968 , \40969 , \40970 , \40971 , \40972 ,
         \40973 , \40974 , \40975 , \40976 , \40977 , \40978 , \40979 , \40980 , \40981 , \40982 ,
         \40983 , \40984 , \40985 , \40986 , \40987 , \40988 , \40989 , \40990 , \40991 , \40992 ,
         \40993 , \40994 , \40995 , \40996 , \40997 , \40998 , \40999 , \41000 , \41001 , \41002 ,
         \41003 , \41004 , \41005 , \41006 , \41007 , \41008 , \41009 , \41010 , \41011 , \41012 ,
         \41013 , \41014 , \41015 , \41016 , \41017 , \41018 , \41019 , \41020 , \41021 , \41022 ,
         \41023 , \41024 , \41025 , \41026 , \41027 , \41028 , \41029 , \41030 , \41031 , \41032 ,
         \41033 , \41034 , \41035 , \41036 , \41037 , \41038 , \41039 , \41040 , \41041 , \41042 ,
         \41043 , \41044 , \41045 , \41046 , \41047 , \41048 , \41049 , \41050 , \41051 , \41052 ,
         \41053 , \41054 , \41055 , \41056 , \41057 , \41058 , \41059 , \41060 , \41061 , \41062 ,
         \41063 , \41064 , \41065 , \41066 , \41067 , \41068 , \41069 , \41070 , \41071 , \41072 ,
         \41073 , \41074 , \41075 , \41076 , \41077 , \41078 , \41079 , \41080 , \41081 , \41082 ,
         \41083 , \41084 , \41085 , \41086 , \41087 , \41088 , \41089 , \41090 , \41091 , \41092 ,
         \41093 , \41094 , \41095 , \41096 , \41097 , \41098 , \41099 , \41100 , \41101 , \41102 ,
         \41103 , \41104 , \41105 , \41106 , \41107 , \41108 , \41109 , \41110 , \41111 , \41112 ,
         \41113 , \41114 , \41115 , \41116 , \41117 , \41118 , \41119 , \41120 , \41121 , \41122 ,
         \41123 , \41124 , \41125 , \41126 , \41127 , \41128 , \41129 , \41130 , \41131 , \41132 ,
         \41133 , \41134 , \41135 , \41136 , \41137 , \41138 , \41139 , \41140 , \41141 , \41142 ,
         \41143 , \41144 , \41145 , \41146 , \41147 , \41148 , \41149 , \41150 , \41151 , \41152 ,
         \41153 , \41154 , \41155 , \41156 , \41157 , \41158 , \41159 , \41160 , \41161 , \41162 ,
         \41163 , \41164 , \41165 , \41166 , \41167 , \41168 , \41169 , \41170 , \41171 , \41172 ,
         \41173 , \41174 , \41175 , \41176 , \41177 , \41178 , \41179 , \41180 , \41181 , \41182 ,
         \41183 , \41184 , \41185 , \41186 , \41187 , \41188 , \41189 , \41190 , \41191 , \41192 ,
         \41193 , \41194 , \41195 , \41196 , \41197 , \41198 , \41199 , \41200 , \41201 , \41202 ,
         \41203 , \41204 , \41205 , \41206 , \41207 , \41208 , \41209 , \41210 , \41211 , \41212 ,
         \41213 , \41214 , \41215 , \41216 , \41217 , \41218 , \41219 , \41220 , \41221 , \41222 ,
         \41223 , \41224 , \41225 , \41226 , \41227 , \41228 , \41229 , \41230 , \41231 , \41232 ,
         \41233 , \41234 , \41235 , \41236 , \41237 , \41238 , \41239 , \41240 , \41241 , \41242 ,
         \41243 , \41244 , \41245 , \41246 , \41247 , \41248 , \41249 , \41250 , \41251 , \41252 ,
         \41253 , \41254 , \41255 , \41256 , \41257 , \41258 , \41259 , \41260 , \41261 , \41262 ,
         \41263 , \41264 , \41265 , \41266 , \41267 , \41268 , \41269 , \41270 , \41271 , \41272 ,
         \41273 , \41274 , \41275 , \41276 , \41277 , \41278 , \41279 , \41280 , \41281 , \41282 ,
         \41283 , \41284 , \41285 , \41286 , \41287 , \41288 , \41289 , \41290 , \41291 , \41292 ,
         \41293 , \41294 , \41295 , \41296 , \41297 , \41298 , \41299 , \41300 , \41301 , \41302 ,
         \41303 , \41304 , \41305 , \41306 , \41307 , \41308 , \41309 , \41310 , \41311 , \41312 ,
         \41313 , \41314 , \41315 , \41316 , \41317 , \41318 , \41319 , \41320 , \41321 , \41322 ,
         \41323 , \41324 , \41325 , \41326 , \41327 , \41328 , \41329 , \41330 , \41331 , \41332 ,
         \41333 , \41334 , \41335 , \41336 , \41337 , \41338 , \41339 , \41340 , \41341 , \41342 ,
         \41343 , \41344 , \41345 , \41346 , \41347 , \41348 , \41349 , \41350 , \41351 , \41352 ,
         \41353 , \41354 , \41355 , \41356 , \41357 , \41358 , \41359 , \41360 , \41361 , \41362 ,
         \41363 , \41364 , \41365 , \41366 , \41367 , \41368 , \41369 , \41370 , \41371 , \41372 ,
         \41373 , \41374 , \41375 , \41376 , \41377 , \41378 , \41379 , \41380 , \41381 , \41382 ,
         \41383 , \41384 , \41385 , \41386 , \41387 , \41388 , \41389 , \41390 , \41391 , \41392 ,
         \41393 , \41394 , \41395 , \41396 , \41397 , \41398 , \41399 , \41400 , \41401 , \41402 ,
         \41403 , \41404 , \41405 , \41406 , \41407 , \41408 , \41409 , \41410 , \41411 , \41412 ,
         \41413 , \41414 , \41415 , \41416 , \41417 , \41418 , \41419 , \41420 , \41421 , \41422 ,
         \41423 , \41424 , \41425 , \41426 , \41427 , \41428 , \41429 , \41430 , \41431 , \41432 ,
         \41433 , \41434 , \41435 , \41436 , \41437 , \41438 , \41439 , \41440 , \41441 , \41442 ,
         \41443 , \41444 , \41445 , \41446 , \41447 , \41448 , \41449 , \41450 , \41451 , \41452 ,
         \41453 , \41454 , \41455 , \41456 , \41457 , \41458 , \41459 , \41460 , \41461 , \41462 ,
         \41463 , \41464 , \41465 , \41466 , \41467 , \41468 , \41469 , \41470 , \41471 , \41472 ,
         \41473 , \41474 , \41475 , \41476 , \41477 , \41478 , \41479 , \41480 , \41481 , \41482 ,
         \41483 , \41484 , \41485 , \41486 , \41487 , \41488 , \41489 , \41490 , \41491 , \41492 ,
         \41493 , \41494 , \41495 , \41496 , \41497 , \41498 , \41499 , \41500 , \41501 , \41502 ,
         \41503 , \41504 , \41505 , \41506 , \41507 , \41508 , \41509 , \41510 , \41511 , \41512 ,
         \41513 , \41514 , \41515 , \41516 , \41517 , \41518 , \41519 , \41520 , \41521 , \41522 ,
         \41523 , \41524 , \41525 , \41526 , \41527 , \41528 , \41529 , \41530 , \41531 , \41532 ,
         \41533 , \41534 , \41535 , \41536 , \41537 , \41538 , \41539 , \41540 , \41541 , \41542 ,
         \41543 , \41544 , \41545 , \41546 , \41547 , \41548 , \41549 , \41550 , \41551 , \41552 ,
         \41553 , \41554 , \41555 , \41556 , \41557 , \41558 , \41559 , \41560 , \41561 , \41562 ,
         \41563 , \41564 , \41565 , \41566 , \41567 , \41568 , \41569 , \41570 , \41571 , \41572 ,
         \41573 , \41574 , \41575 , \41576 , \41577 , \41578 , \41579 , \41580 , \41581 , \41582 ,
         \41583 , \41584 , \41585 , \41586 , \41587 , \41588 , \41589 , \41590 , \41591 , \41592 ,
         \41593 , \41594 , \41595 , \41596 , \41597 , \41598 , \41599 , \41600 , \41601 , \41602 ,
         \41603 , \41604 , \41605 , \41606 , \41607 , \41608 , \41609 , \41610 , \41611 , \41612 ,
         \41613 , \41614 , \41615 , \41616 , \41617 , \41618 , \41619 , \41620 , \41621 , \41622 ,
         \41623 , \41624 , \41625 , \41626 , \41627 , \41628 , \41629 , \41630 , \41631 , \41632 ,
         \41633 , \41634 , \41635 , \41636 , \41637 , \41638 , \41639 , \41640 , \41641 , \41642 ,
         \41643 , \41644 , \41645 , \41646 , \41647 , \41648 , \41649 , \41650 , \41651 , \41652 ,
         \41653 , \41654 , \41655 , \41656 , \41657 , \41658 , \41659 , \41660 , \41661 , \41662 ,
         \41663 , \41664 , \41665 , \41666 , \41667 , \41668 , \41669 , \41670 , \41671 , \41672 ,
         \41673 , \41674 , \41675 , \41676 , \41677 , \41678 , \41679 , \41680 , \41681 , \41682 ,
         \41683 , \41684 , \41685 , \41686 , \41687 , \41688 , \41689 , \41690 , \41691 , \41692 ,
         \41693 , \41694 , \41695 , \41696 , \41697 , \41698 , \41699 , \41700 , \41701 , \41702 ,
         \41703 , \41704 , \41705 , \41706 , \41707 , \41708 , \41709 , \41710 , \41711 , \41712 ,
         \41713 , \41714 , \41715 , \41716 , \41717 , \41718 , \41719 , \41720 , \41721 , \41722 ,
         \41723 , \41724 , \41725 , \41726 , \41727 , \41728 , \41729 , \41730 , \41731 , \41732 ,
         \41733 , \41734 , \41735 , \41736 , \41737 , \41738 , \41739 , \41740 , \41741 , \41742 ,
         \41743 , \41744 , \41745 , \41746 , \41747 , \41748 , \41749 , \41750 , \41751 , \41752 ,
         \41753 , \41754 , \41755 , \41756 , \41757 , \41758 , \41759 , \41760 , \41761 , \41762 ,
         \41763 , \41764 , \41765 , \41766 , \41767 , \41768 , \41769 , \41770 , \41771 , \41772 ,
         \41773 , \41774 , \41775 , \41776 , \41777 , \41778 , \41779 , \41780 , \41781 , \41782 ,
         \41783 , \41784 , \41785 , \41786 , \41787 , \41788 , \41789 , \41790 , \41791 , \41792 ,
         \41793 , \41794 , \41795 , \41796 , \41797 , \41798 , \41799 , \41800 , \41801 , \41802 ,
         \41803 , \41804 , \41805 , \41806 , \41807 , \41808 , \41809 , \41810 , \41811 , \41812 ,
         \41813 , \41814 , \41815 , \41816 , \41817 , \41818 , \41819 , \41820 , \41821 , \41822 ,
         \41823 , \41824 , \41825 , \41826 , \41827 , \41828 , \41829 , \41830 , \41831 , \41832 ,
         \41833 , \41834 , \41835 , \41836 , \41837 , \41838 , \41839 , \41840 , \41841 , \41842 ,
         \41843 , \41844 , \41845 , \41846 , \41847 , \41848 , \41849 , \41850 , \41851 , \41852 ,
         \41853 , \41854 , \41855 , \41856 , \41857 , \41858 , \41859 , \41860 , \41861 , \41862 ,
         \41863 , \41864 , \41865 , \41866 , \41867 , \41868 , \41869 , \41870 , \41871 , \41872 ,
         \41873 , \41874 , \41875 , \41876 , \41877 , \41878 , \41879 , \41880 , \41881 , \41882 ,
         \41883 , \41884 , \41885 , \41886 , \41887 , \41888 , \41889 , \41890 , \41891 , \41892 ,
         \41893 , \41894 , \41895 , \41896 , \41897 , \41898 , \41899 , \41900 , \41901 , \41902 ,
         \41903 , \41904 , \41905 , \41906 , \41907 , \41908 , \41909 , \41910 , \41911 , \41912 ,
         \41913 , \41914 , \41915 , \41916 , \41917 , \41918 , \41919 , \41920 , \41921 , \41922 ,
         \41923 , \41924 , \41925 , \41926 , \41927 , \41928 , \41929 , \41930 , \41931 , \41932 ,
         \41933 , \41934 , \41935 , \41936 , \41937 , \41938 , \41939 , \41940 , \41941 , \41942 ,
         \41943 , \41944 , \41945 , \41946 , \41947 , \41948 , \41949 , \41950 , \41951 , \41952 ,
         \41953 , \41954 , \41955 , \41956 , \41957 , \41958 , \41959 , \41960 , \41961 , \41962 ,
         \41963 , \41964 , \41965 , \41966 , \41967 , \41968 , \41969 , \41970 , \41971 , \41972 ,
         \41973 , \41974 , \41975 , \41976 , \41977 , \41978 , \41979 , \41980 , \41981 , \41982 ,
         \41983 , \41984 , \41985 , \41986 , \41987 , \41988 , \41989 , \41990 , \41991 , \41992 ,
         \41993 , \41994 , \41995 , \41996 , \41997 , \41998 , \41999 , \42000 , \42001 , \42002 ,
         \42003 , \42004 , \42005 , \42006 , \42007 , \42008 , \42009 , \42010 , \42011 , \42012 ,
         \42013 , \42014 , \42015 , \42016 , \42017 , \42018 , \42019 , \42020 , \42021 , \42022 ,
         \42023 , \42024 , \42025 , \42026 , \42027 , \42028 , \42029 , \42030 , \42031 , \42032 ,
         \42033 , \42034 , \42035 , \42036 , \42037 , \42038 , \42039 , \42040 , \42041 , \42042 ,
         \42043 , \42044 , \42045 , \42046 , \42047 , \42048 , \42049 , \42050 , \42051 , \42052 ,
         \42053 , \42054 , \42055 , \42056 , \42057 , \42058 , \42059 , \42060 , \42061 , \42062 ,
         \42063 , \42064 , \42065 , \42066 , \42067 , \42068 , \42069 , \42070 , \42071 , \42072 ,
         \42073 , \42074 , \42075 , \42076 , \42077 , \42078 , \42079 , \42080 , \42081 , \42082 ,
         \42083 , \42084 , \42085 , \42086 , \42087 , \42088 , \42089 , \42090 , \42091 , \42092 ,
         \42093 , \42094 , \42095 , \42096 , \42097 , \42098 , \42099 , \42100 , \42101 , \42102 ,
         \42103 , \42104 , \42105 , \42106 , \42107 , \42108 , \42109 , \42110 , \42111 , \42112 ,
         \42113 , \42114 , \42115 , \42116 , \42117 , \42118 , \42119 , \42120 , \42121 , \42122 ,
         \42123 , \42124 , \42125 , \42126 , \42127 , \42128 , \42129 , \42130 , \42131 , \42132 ,
         \42133 , \42134 , \42135 , \42136 , \42137 , \42138 , \42139 , \42140 , \42141 , \42142 ,
         \42143 , \42144 , \42145 , \42146 , \42147 , \42148 , \42149 , \42150 , \42151 , \42152 ,
         \42153 , \42154 , \42155 , \42156 , \42157 , \42158 , \42159 , \42160 , \42161 , \42162 ,
         \42163 , \42164 , \42165 , \42166 , \42167 , \42168 , \42169 , \42170 , \42171 , \42172 ,
         \42173 , \42174 , \42175 , \42176 , \42177 , \42178 , \42179 , \42180 , \42181 , \42182 ,
         \42183 , \42184 , \42185 , \42186 , \42187 , \42188 , \42189 , \42190 , \42191 , \42192 ,
         \42193 , \42194 , \42195 , \42196 , \42197 , \42198 , \42199 , \42200 , \42201 , \42202 ,
         \42203 , \42204 , \42205 , \42206 , \42207 , \42208 , \42209 , \42210 , \42211 , \42212 ,
         \42213 , \42214 , \42215 , \42216 , \42217 , \42218 , \42219 , \42220 , \42221 , \42222 ,
         \42223 , \42224 , \42225 , \42226 , \42227 , \42228 , \42229 , \42230 , \42231 , \42232 ,
         \42233 , \42234 , \42235 , \42236 , \42237 , \42238 , \42239 , \42240 , \42241 , \42242 ,
         \42243 , \42244 , \42245 , \42246 , \42247 , \42248 , \42249 , \42250 , \42251 , \42252 ,
         \42253 , \42254 , \42255 , \42256 , \42257 , \42258 , \42259 , \42260 , \42261 , \42262 ,
         \42263 , \42264 , \42265 , \42266 , \42267 , \42268 , \42269 , \42270 , \42271 , \42272 ,
         \42273 , \42274 , \42275 , \42276 , \42277 , \42278 , \42279 , \42280 , \42281 , \42282 ,
         \42283 , \42284 , \42285 , \42286 , \42287 , \42288 , \42289 , \42290 , \42291 , \42292 ,
         \42293 , \42294 , \42295 , \42296 , \42297 , \42298 , \42299 , \42300 , \42301 , \42302 ,
         \42303 , \42304 , \42305 , \42306 , \42307 , \42308 , \42309 , \42310 , \42311 , \42312 ,
         \42313 , \42314 , \42315 , \42316 , \42317 , \42318 , \42319 , \42320 , \42321 , \42322 ,
         \42323 , \42324 , \42325 , \42326 , \42327 , \42328 , \42329 , \42330 , \42331 , \42332 ,
         \42333 , \42334 , \42335 , \42336 , \42337 , \42338 , \42339 , \42340 , \42341 , \42342 ,
         \42343 , \42344 , \42345 , \42346 , \42347 , \42348 , \42349 , \42350 , \42351 , \42352 ,
         \42353 , \42354 , \42355 , \42356 , \42357 , \42358 , \42359 , \42360 , \42361 , \42362 ,
         \42363 , \42364 , \42365 , \42366 , \42367 , \42368 , \42369 , \42370 , \42371 , \42372 ,
         \42373 , \42374 , \42375 , \42376 , \42377 , \42378 , \42379 , \42380 , \42381 , \42382 ,
         \42383 , \42384 , \42385 , \42386 , \42387 , \42388 , \42389 , \42390 , \42391 , \42392 ,
         \42393 , \42394 , \42395 , \42396 , \42397 , \42398 , \42399 , \42400 , \42401 , \42402 ,
         \42403 , \42404 , \42405 , \42406 , \42407 , \42408 , \42409 , \42410 , \42411 , \42412 ,
         \42413 , \42414 , \42415 , \42416 , \42417 , \42418 , \42419 , \42420 , \42421 , \42422 ,
         \42423 , \42424 , \42425 , \42426 , \42427 , \42428 , \42429 , \42430 , \42431 , \42432 ,
         \42433 , \42434 , \42435 , \42436 , \42437 , \42438 , \42439 , \42440 , \42441 , \42442 ,
         \42443 , \42444 , \42445 , \42446 , \42447 , \42448 , \42449 , \42450 , \42451 , \42452 ,
         \42453 , \42454 , \42455 , \42456 , \42457 , \42458 , \42459 , \42460 , \42461 , \42462 ,
         \42463 , \42464 , \42465 , \42466 , \42467 , \42468 , \42469 , \42470 , \42471 , \42472 ,
         \42473 , \42474 , \42475 , \42476 , \42477 , \42478 , \42479 , \42480 , \42481 , \42482 ,
         \42483 , \42484 , \42485 , \42486 , \42487 , \42488 , \42489 , \42490 , \42491 , \42492 ,
         \42493 , \42494 , \42495 , \42496 , \42497 , \42498 , \42499 , \42500 , \42501 , \42502 ,
         \42503 , \42504 , \42505 , \42506 , \42507 , \42508 , \42509 , \42510 , \42511 , \42512 ,
         \42513 , \42514 , \42515 , \42516 , \42517 , \42518 , \42519 , \42520 , \42521 , \42522 ,
         \42523 , \42524 , \42525 , \42526 , \42527 , \42528 , \42529 , \42530 , \42531 , \42532 ,
         \42533 , \42534 , \42535 , \42536 , \42537 , \42538 , \42539 , \42540 , \42541 , \42542 ,
         \42543 , \42544 , \42545 , \42546 , \42547 , \42548 , \42549 , \42550 , \42551 , \42552 ,
         \42553 , \42554 , \42555 , \42556 , \42557 , \42558 , \42559 , \42560 , \42561 , \42562 ,
         \42563 , \42564 , \42565 , \42566 , \42567 , \42568 , \42569 , \42570 , \42571 , \42572 ,
         \42573 , \42574 , \42575 , \42576 , \42577 , \42578 , \42579 , \42580 , \42581 , \42582 ,
         \42583 , \42584 , \42585 , \42586 , \42587 , \42588 , \42589 , \42590 , \42591 , \42592 ,
         \42593 , \42594 , \42595 , \42596 , \42597 , \42598 , \42599 , \42600 , \42601 , \42602 ,
         \42603 , \42604 , \42605 , \42606 , \42607 , \42608 , \42609 , \42610 , \42611 , \42612 ,
         \42613 , \42614 , \42615 , \42616 , \42617 , \42618 , \42619 , \42620 , \42621 , \42622 ,
         \42623 , \42624 , \42625 , \42626 , \42627 , \42628 , \42629 , \42630 , \42631 , \42632 ,
         \42633 , \42634 , \42635 , \42636 , \42637 , \42638 , \42639 , \42640 , \42641 , \42642 ,
         \42643 , \42644 , \42645 , \42646 , \42647 , \42648 , \42649 , \42650 , \42651 , \42652 ,
         \42653 , \42654 , \42655 , \42656 , \42657 , \42658 , \42659 , \42660 , \42661 , \42662 ,
         \42663 , \42664 , \42665 , \42666 , \42667 , \42668 , \42669 , \42670 , \42671 , \42672 ,
         \42673 , \42674 , \42675 , \42676 , \42677 , \42678 , \42679 , \42680 , \42681 , \42682 ,
         \42683 , \42684 , \42685 , \42686 , \42687 , \42688 , \42689 , \42690 , \42691 , \42692 ,
         \42693 , \42694 , \42695 , \42696 , \42697 , \42698 , \42699 , \42700 , \42701 , \42702 ,
         \42703 , \42704 , \42705 , \42706 , \42707 , \42708 , \42709 , \42710 , \42711 , \42712 ,
         \42713 , \42714 , \42715 , \42716 , \42717 , \42718 , \42719 , \42720 , \42721 , \42722 ,
         \42723 , \42724 , \42725 , \42726 , \42727 , \42728 , \42729 , \42730 , \42731 , \42732 ,
         \42733 , \42734 , \42735 , \42736 , \42737 , \42738 , \42739 , \42740 , \42741 , \42742 ,
         \42743 , \42744 , \42745 , \42746 , \42747 , \42748 , \42749 , \42750 , \42751 , \42752 ,
         \42753 , \42754 , \42755 , \42756 , \42757 , \42758 , \42759 , \42760 , \42761 , \42762 ,
         \42763 , \42764 , \42765 , \42766 , \42767 , \42768 , \42769 , \42770 , \42771 , \42772 ,
         \42773 , \42774 , \42775 , \42776 , \42777 , \42778 , \42779 , \42780 , \42781 , \42782 ,
         \42783 , \42784 , \42785 , \42786 , \42787 , \42788 , \42789 , \42790 , \42791 , \42792 ,
         \42793 , \42794 , \42795 , \42796 , \42797 , \42798 , \42799 , \42800 , \42801 , \42802 ,
         \42803 , \42804 , \42805 , \42806 , \42807 , \42808 , \42809 , \42810 , \42811 , \42812 ,
         \42813 , \42814 , \42815 , \42816 , \42817 , \42818 , \42819 , \42820 , \42821 , \42822 ,
         \42823 , \42824 , \42825 , \42826 , \42827 , \42828 , \42829 , \42830 , \42831 , \42832 ,
         \42833 , \42834 , \42835 , \42836 , \42837 , \42838 , \42839 , \42840 , \42841 , \42842 ,
         \42843 , \42844 , \42845 , \42846 , \42847 , \42848 , \42849 , \42850 , \42851 , \42852 ,
         \42853 , \42854 , \42855 , \42856 , \42857 , \42858 , \42859 , \42860 , \42861 , \42862 ,
         \42863 , \42864 , \42865 , \42866 , \42867 , \42868 , \42869 , \42870 , \42871 , \42872 ,
         \42873 , \42874 , \42875 , \42876 , \42877 , \42878 , \42879 , \42880 , \42881 , \42882 ,
         \42883 , \42884 , \42885 , \42886 , \42887 , \42888 , \42889 , \42890 , \42891 , \42892 ,
         \42893 , \42894 , \42895 , \42896 , \42897 , \42898 , \42899 , \42900 , \42901 , \42902 ,
         \42903 , \42904 , \42905 , \42906 , \42907 , \42908 , \42909 , \42910 , \42911 , \42912 ,
         \42913 , \42914 , \42915 , \42916 , \42917 , \42918 , \42919 , \42920 , \42921 , \42922 ,
         \42923 , \42924 , \42925 , \42926 , \42927 , \42928 , \42929 , \42930 , \42931 , \42932 ,
         \42933 , \42934 , \42935 , \42936 , \42937 , \42938 , \42939 , \42940 , \42941 , \42942 ,
         \42943 , \42944 , \42945 , \42946 , \42947 , \42948 , \42949 , \42950 , \42951 , \42952 ,
         \42953 , \42954 , \42955 , \42956 , \42957 , \42958 , \42959 , \42960 , \42961 , \42962 ,
         \42963 , \42964 , \42965 , \42966 , \42967 , \42968 , \42969 , \42970 , \42971 , \42972 ,
         \42973 , \42974 , \42975 , \42976 , \42977 , \42978 , \42979 , \42980 , \42981 , \42982 ,
         \42983 , \42984 , \42985 , \42986 , \42987 , \42988 , \42989 , \42990 , \42991 , \42992 ,
         \42993 , \42994 , \42995 , \42996 , \42997 , \42998 , \42999 , \43000 , \43001 , \43002 ,
         \43003 , \43004 , \43005 , \43006 , \43007 , \43008 , \43009 , \43010 , \43011 , \43012 ,
         \43013 , \43014 , \43015 , \43016 , \43017 , \43018 , \43019 , \43020 , \43021 , \43022 ,
         \43023 , \43024 , \43025 , \43026 , \43027 , \43028 , \43029 , \43030 , \43031 , \43032 ,
         \43033 , \43034 , \43035 , \43036 , \43037 , \43038 , \43039 , \43040 , \43041 , \43042 ,
         \43043 , \43044 , \43045 , \43046 , \43047 , \43048 , \43049 , \43050 , \43051 , \43052 ,
         \43053 , \43054 , \43055 , \43056 , \43057 , \43058 , \43059 , \43060 , \43061 , \43062 ,
         \43063 , \43064 , \43065 , \43066 , \43067 , \43068 , \43069 , \43070 , \43071 , \43072 ,
         \43073 , \43074 , \43075 , \43076 , \43077 , \43078 , \43079 , \43080 , \43081 , \43082 ,
         \43083 , \43084 , \43085 , \43086 , \43087 , \43088 , \43089 , \43090 , \43091 , \43092 ,
         \43093 , \43094 , \43095 , \43096 , \43097 , \43098 , \43099 , \43100 , \43101 , \43102 ,
         \43103 , \43104 , \43105 , \43106 , \43107 , \43108 , \43109 , \43110 , \43111 , \43112 ,
         \43113 , \43114 , \43115 , \43116 , \43117 , \43118 , \43119 , \43120 , \43121 , \43122 ,
         \43123 , \43124 , \43125 , \43126 , \43127 , \43128 , \43129 , \43130 , \43131 , \43132 ,
         \43133 , \43134 , \43135 , \43136 , \43137 , \43138 , \43139 , \43140 , \43141 , \43142 ,
         \43143 , \43144 , \43145 , \43146 , \43147 , \43148 , \43149 , \43150 , \43151 , \43152 ,
         \43153 , \43154 , \43155 , \43156 , \43157 , \43158 , \43159 , \43160 , \43161 , \43162 ,
         \43163 , \43164 , \43165 , \43166 , \43167 , \43168 , \43169 , \43170 , \43171 , \43172 ,
         \43173 , \43174 , \43175 , \43176 , \43177 , \43178 , \43179 , \43180 , \43181 , \43182 ,
         \43183 , \43184 , \43185 , \43186 , \43187 , \43188 , \43189 , \43190 , \43191 , \43192 ,
         \43193 , \43194 , \43195 , \43196 , \43197 , \43198 , \43199 , \43200 , \43201 , \43202 ,
         \43203 , \43204 , \43205 , \43206 , \43207 , \43208 , \43209 , \43210 , \43211 , \43212 ,
         \43213 , \43214 , \43215 , \43216 , \43217 , \43218 , \43219 , \43220 , \43221 , \43222 ,
         \43223 , \43224 , \43225 , \43226 , \43227 , \43228 , \43229 , \43230 , \43231 , \43232 ,
         \43233 , \43234 , \43235 , \43236 , \43237 , \43238 , \43239 , \43240 , \43241 , \43242 ,
         \43243 , \43244 , \43245 , \43246 , \43247 , \43248 , \43249 , \43250 , \43251 , \43252 ,
         \43253 , \43254 , \43255 , \43256 , \43257 , \43258 , \43259 , \43260 , \43261 , \43262 ,
         \43263 , \43264 , \43265 , \43266 , \43267 , \43268 , \43269 , \43270 , \43271 , \43272 ,
         \43273 , \43274 , \43275 , \43276 , \43277 , \43278 , \43279 , \43280 , \43281 , \43282 ,
         \43283 , \43284 , \43285 , \43286 , \43287 , \43288 , \43289 , \43290 , \43291 , \43292 ,
         \43293 , \43294 , \43295 , \43296 , \43297 , \43298 , \43299 , \43300 , \43301 , \43302 ,
         \43303 , \43304 , \43305 , \43306 , \43307 , \43308 , \43309 , \43310 , \43311 , \43312 ,
         \43313 , \43314 , \43315 , \43316 , \43317 , \43318 , \43319 , \43320 , \43321 , \43322 ,
         \43323 , \43324 , \43325 , \43326 , \43327 , \43328 , \43329 , \43330 , \43331 , \43332 ,
         \43333 , \43334 , \43335 , \43336 , \43337 , \43338 , \43339 , \43340 , \43341 , \43342 ,
         \43343 , \43344 , \43345 , \43346 , \43347 , \43348 , \43349 , \43350 , \43351 , \43352 ,
         \43353 , \43354 , \43355 , \43356 , \43357 , \43358 , \43359 , \43360 , \43361 , \43362 ,
         \43363 , \43364 , \43365 , \43366 , \43367 , \43368 , \43369 , \43370 , \43371 , \43372 ,
         \43373 , \43374 , \43375 , \43376 , \43377 , \43378 , \43379 , \43380 , \43381 , \43382 ,
         \43383 , \43384 , \43385 , \43386 , \43387 , \43388 , \43389 , \43390 , \43391 , \43392 ,
         \43393 , \43394 , \43395 , \43396 , \43397 , \43398 , \43399 , \43400 , \43401 , \43402 ,
         \43403 , \43404 , \43405 , \43406 , \43407 , \43408 , \43409 , \43410 , \43411 , \43412 ,
         \43413 , \43414 , \43415 , \43416 , \43417 , \43418 , \43419 , \43420 , \43421 , \43422 ,
         \43423 , \43424 , \43425 , \43426 , \43427 , \43428 , \43429 , \43430 , \43431 , \43432 ,
         \43433 , \43434 , \43435 , \43436 , \43437 , \43438 , \43439 , \43440 , \43441 , \43442 ,
         \43443 , \43444 , \43445 , \43446 , \43447 , \43448 , \43449 , \43450 , \43451 , \43452 ,
         \43453 , \43454 , \43455 , \43456 , \43457 , \43458 , \43459 , \43460 , \43461 , \43462 ,
         \43463 , \43464 , \43465 , \43466 , \43467 , \43468 , \43469 , \43470 , \43471 , \43472 ,
         \43473 , \43474 , \43475 , \43476 , \43477 , \43478 , \43479 , \43480 , \43481 , \43482 ,
         \43483 , \43484 , \43485 , \43486 , \43487 , \43488 , \43489 , \43490 , \43491 , \43492 ,
         \43493 , \43494 , \43495 , \43496 , \43497 , \43498 , \43499 , \43500 , \43501 , \43502 ,
         \43503 , \43504 , \43505 , \43506 , \43507 , \43508 , \43509 , \43510 , \43511 , \43512 ,
         \43513 , \43514 , \43515 , \43516 , \43517 , \43518 , \43519 , \43520 , \43521 , \43522 ,
         \43523 , \43524 , \43525 , \43526 , \43527 , \43528 , \43529 , \43530 , \43531 , \43532 ,
         \43533 , \43534 , \43535 , \43536 , \43537 , \43538 , \43539 , \43540 , \43541 , \43542 ,
         \43543 , \43544 , \43545 , \43546 , \43547 , \43548 , \43549 , \43550 , \43551 , \43552 ,
         \43553 , \43554 , \43555 , \43556 , \43557 , \43558 , \43559 , \43560 , \43561 , \43562 ,
         \43563 , \43564 , \43565 , \43566 , \43567 , \43568 , \43569 , \43570 , \43571 , \43572 ,
         \43573 , \43574 , \43575 , \43576 , \43577 , \43578 , \43579 , \43580 , \43581 , \43582 ,
         \43583 , \43584 , \43585 , \43586 , \43587 , \43588 , \43589 , \43590 , \43591 , \43592 ,
         \43593 , \43594 , \43595 , \43596 , \43597 , \43598 , \43599 , \43600 , \43601 , \43602 ,
         \43603 , \43604 , \43605 , \43606 , \43607 , \43608 , \43609 , \43610 , \43611 , \43612 ,
         \43613 , \43614 , \43615 , \43616 , \43617 , \43618 , \43619 , \43620 , \43621 , \43622 ,
         \43623 , \43624 , \43625 , \43626 , \43627 , \43628 , \43629 , \43630 , \43631 , \43632 ,
         \43633 , \43634 , \43635 , \43636 , \43637 , \43638 , \43639 , \43640 , \43641 , \43642 ,
         \43643 , \43644 , \43645 , \43646 , \43647 , \43648 , \43649 , \43650 , \43651 , \43652 ,
         \43653 , \43654 , \43655 , \43656 , \43657 , \43658 , \43659 , \43660 , \43661 , \43662 ,
         \43663 , \43664 , \43665 , \43666 , \43667 , \43668 , \43669 , \43670 , \43671 , \43672 ,
         \43673 , \43674 , \43675 , \43676 , \43677 , \43678 , \43679 , \43680 , \43681 , \43682 ,
         \43683 , \43684 , \43685 , \43686 , \43687 , \43688 , \43689 , \43690 , \43691 , \43692 ,
         \43693 , \43694 , \43695 , \43696 , \43697 , \43698 , \43699 , \43700 , \43701 , \43702 ,
         \43703 , \43704 , \43705 , \43706 , \43707 , \43708 , \43709 , \43710 , \43711 , \43712 ,
         \43713 , \43714 , \43715 , \43716 , \43717 , \43718 , \43719 , \43720 , \43721 , \43722 ,
         \43723 , \43724 , \43725 , \43726 , \43727 , \43728 , \43729 , \43730 , \43731 , \43732 ,
         \43733 , \43734 , \43735 , \43736 , \43737 , \43738 , \43739 , \43740 , \43741 , \43742 ,
         \43743 , \43744 , \43745 , \43746 , \43747 , \43748 , \43749 , \43750 , \43751 , \43752 ,
         \43753 , \43754 , \43755 , \43756 , \43757 , \43758 , \43759 , \43760 , \43761 , \43762 ,
         \43763 , \43764 , \43765 , \43766 , \43767 , \43768 , \43769 , \43770 , \43771 , \43772 ,
         \43773 , \43774 , \43775 , \43776 , \43777 , \43778 , \43779 , \43780 , \43781 , \43782 ,
         \43783 , \43784 , \43785 , \43786 , \43787 , \43788 , \43789 , \43790 , \43791 , \43792 ,
         \43793 , \43794 , \43795 , \43796 , \43797 , \43798 , \43799 , \43800 , \43801 , \43802 ,
         \43803 , \43804 , \43805 , \43806 , \43807 , \43808 , \43809 , \43810 , \43811 , \43812 ,
         \43813 , \43814 , \43815 , \43816 , \43817 , \43818 , \43819 , \43820 , \43821 , \43822 ,
         \43823 , \43824 , \43825 , \43826 , \43827 , \43828 , \43829 , \43830 , \43831 , \43832 ,
         \43833 , \43834 , \43835 , \43836 , \43837 , \43838 , \43839 , \43840 , \43841 , \43842 ,
         \43843 , \43844 , \43845 , \43846 , \43847 , \43848 , \43849 , \43850 , \43851 , \43852 ,
         \43853 , \43854 , \43855 , \43856 , \43857 , \43858 , \43859 , \43860 , \43861 , \43862 ,
         \43863 , \43864 , \43865 , \43866 , \43867 , \43868 , \43869 , \43870 , \43871 , \43872 ,
         \43873 , \43874 , \43875 , \43876 , \43877 , \43878 , \43879 , \43880 , \43881 , \43882 ,
         \43883 , \43884 , \43885 , \43886 , \43887 , \43888 , \43889 , \43890 , \43891 , \43892 ,
         \43893 , \43894 , \43895 , \43896 , \43897 , \43898 , \43899 , \43900 , \43901 , \43902 ,
         \43903 , \43904 , \43905 , \43906 , \43907 , \43908 , \43909 , \43910 , \43911 , \43912 ,
         \43913 , \43914 , \43915 , \43916 , \43917 , \43918 , \43919 , \43920 , \43921 , \43922 ,
         \43923 , \43924 , \43925 , \43926 , \43927 , \43928 , \43929 , \43930 , \43931 , \43932 ,
         \43933 , \43934 , \43935 , \43936 , \43937 , \43938 , \43939 , \43940 , \43941 , \43942 ,
         \43943 , \43944 , \43945 , \43946 , \43947 , \43948 , \43949 , \43950 , \43951 , \43952 ,
         \43953 , \43954 , \43955 , \43956 , \43957 , \43958 , \43959 , \43960 , \43961 , \43962 ,
         \43963 , \43964 , \43965 , \43966 , \43967 , \43968 , \43969 , \43970 , \43971 , \43972 ,
         \43973 , \43974 , \43975 , \43976 , \43977 , \43978 , \43979 , \43980 , \43981 , \43982 ,
         \43983 , \43984 , \43985 , \43986 , \43987 , \43988 , \43989 , \43990 , \43991 , \43992 ,
         \43993 , \43994 , \43995 , \43996 , \43997 , \43998 , \43999 , \44000 , \44001 , \44002 ,
         \44003 , \44004 , \44005 , \44006 , \44007 , \44008 , \44009 , \44010 , \44011 , \44012 ,
         \44013 , \44014 , \44015 , \44016 , \44017 , \44018 , \44019 , \44020 , \44021 , \44022 ,
         \44023 , \44024 , \44025 , \44026 , \44027 , \44028 , \44029 , \44030 , \44031 , \44032 ,
         \44033 , \44034 , \44035 , \44036 , \44037 , \44038 , \44039 , \44040 , \44041 , \44042 ,
         \44043 , \44044 , \44045 , \44046 , \44047 , \44048 , \44049 , \44050 , \44051 , \44052 ,
         \44053 , \44054 , \44055 , \44056 , \44057 , \44058 , \44059 , \44060 , \44061 , \44062 ,
         \44063 , \44064 , \44065 , \44066 , \44067 , \44068 , \44069 , \44070 , \44071 , \44072 ,
         \44073 , \44074 , \44075 , \44076 , \44077 , \44078 , \44079 , \44080 , \44081 , \44082 ,
         \44083 , \44084 , \44085 , \44086 , \44087 , \44088 , \44089 , \44090 , \44091 , \44092 ,
         \44093 , \44094 , \44095 , \44096 , \44097 , \44098 , \44099 , \44100 , \44101 , \44102 ,
         \44103 , \44104 , \44105 , \44106 , \44107 , \44108 , \44109 , \44110 , \44111 , \44112 ,
         \44113 , \44114 , \44115 , \44116 , \44117 , \44118 , \44119 , \44120 , \44121 , \44122 ,
         \44123 , \44124 , \44125 , \44126 , \44127 , \44128 , \44129 , \44130 , \44131 , \44132 ,
         \44133 , \44134 , \44135 , \44136 , \44137 , \44138 , \44139 , \44140 , \44141 , \44142 ,
         \44143 , \44144 , \44145 , \44146 , \44147 , \44148 , \44149 , \44150 , \44151 , \44152 ,
         \44153 , \44154 , \44155 , \44156 , \44157 , \44158 , \44159 , \44160 , \44161 , \44162 ,
         \44163 , \44164 , \44165 , \44166 , \44167 , \44168 , \44169 , \44170 , \44171 , \44172 ,
         \44173 , \44174 , \44175 , \44176 , \44177 , \44178 , \44179 , \44180 , \44181 , \44182 ,
         \44183 , \44184 , \44185 , \44186 , \44187 , \44188 , \44189 , \44190 , \44191 , \44192 ,
         \44193 , \44194 , \44195 , \44196 , \44197 , \44198 , \44199 , \44200 , \44201 , \44202 ,
         \44203 , \44204 , \44205 , \44206 , \44207 , \44208 , \44209 , \44210 , \44211 , \44212 ,
         \44213 , \44214 , \44215 , \44216 , \44217 , \44218 , \44219 , \44220 , \44221 , \44222 ,
         \44223 , \44224 , \44225 , \44226 , \44227 , \44228 , \44229 , \44230 , \44231 , \44232 ,
         \44233 , \44234 , \44235 , \44236 , \44237 , \44238 , \44239 , \44240 , \44241 , \44242 ,
         \44243 , \44244 , \44245 , \44246 , \44247 , \44248 , \44249 , \44250 , \44251 , \44252 ,
         \44253 , \44254 , \44255 , \44256 , \44257 , \44258 , \44259 , \44260 , \44261 , \44262 ,
         \44263 , \44264 , \44265 , \44266 , \44267 , \44268 , \44269 , \44270 , \44271 , \44272 ,
         \44273 , \44274 , \44275 , \44276 , \44277 , \44278 , \44279 , \44280 , \44281 , \44282 ,
         \44283 , \44284 , \44285 , \44286 , \44287 , \44288 , \44289 , \44290 , \44291 , \44292 ,
         \44293 , \44294 , \44295 , \44296 , \44297 , \44298 , \44299 , \44300 , \44301 , \44302 ,
         \44303 , \44304 , \44305 , \44306 , \44307 , \44308 , \44309 , \44310 , \44311 , \44312 ,
         \44313 , \44314 , \44315 , \44316 , \44317 , \44318 , \44319 , \44320 , \44321 , \44322 ,
         \44323 , \44324 , \44325 , \44326 , \44327 , \44328 , \44329 , \44330 , \44331 , \44332 ,
         \44333 , \44334 , \44335 , \44336 , \44337 , \44338 , \44339 , \44340 , \44341 , \44342 ,
         \44343 , \44344 , \44345 , \44346 , \44347 , \44348 , \44349 , \44350 , \44351 , \44352 ,
         \44353 , \44354 , \44355 , \44356 , \44357 , \44358 , \44359 , \44360 , \44361 , \44362 ,
         \44363 , \44364 , \44365 , \44366 , \44367 , \44368 , \44369 , \44370 , \44371 , \44372 ,
         \44373 , \44374 , \44375 , \44376 , \44377 , \44378 , \44379 , \44380 , \44381 , \44382 ,
         \44383 , \44384 , \44385 , \44386 , \44387 , \44388 , \44389 , \44390 , \44391 , \44392 ,
         \44393 , \44394 , \44395 , \44396 , \44397 , \44398 , \44399 , \44400 , \44401 , \44402 ,
         \44403 , \44404 , \44405 , \44406 , \44407 , \44408 , \44409 , \44410 , \44411 , \44412 ,
         \44413 , \44414 , \44415 , \44416 , \44417 , \44418 , \44419 , \44420 , \44421 , \44422 ,
         \44423 , \44424 , \44425 , \44426 , \44427 , \44428 , \44429 , \44430 , \44431 , \44432 ,
         \44433 , \44434 , \44435 , \44436 , \44437 , \44438 , \44439 , \44440 , \44441 , \44442 ,
         \44443 , \44444 , \44445 , \44446 , \44447 , \44448 , \44449 , \44450 , \44451 , \44452 ,
         \44453 , \44454 , \44455 , \44456 , \44457 , \44458 , \44459 , \44460 , \44461 , \44462 ,
         \44463 , \44464 , \44465 , \44466 , \44467 , \44468 , \44469 , \44470 , \44471 , \44472 ,
         \44473 , \44474 , \44475 , \44476 , \44477 , \44478 , \44479 , \44480 , \44481 , \44482 ,
         \44483 , \44484 , \44485 , \44486 , \44487 , \44488 , \44489 , \44490 , \44491 , \44492 ,
         \44493 , \44494 , \44495 , \44496 , \44497 , \44498 , \44499 , \44500 , \44501 , \44502 ,
         \44503 , \44504 , \44505 , \44506 , \44507 , \44508 , \44509 , \44510 , \44511 , \44512 ,
         \44513 , \44514 , \44515 , \44516 , \44517 , \44518 , \44519 , \44520 , \44521 , \44522 ,
         \44523 , \44524 , \44525 , \44526 , \44527 , \44528 , \44529 , \44530 , \44531 , \44532 ,
         \44533 , \44534 , \44535 , \44536 , \44537 , \44538 , \44539 , \44540 , \44541 , \44542 ,
         \44543 , \44544 , \44545 , \44546 , \44547 , \44548 , \44549 , \44550 , \44551 , \44552 ,
         \44553 , \44554 , \44555 , \44556 , \44557 , \44558 , \44559 , \44560 , \44561 , \44562 ,
         \44563 , \44564 , \44565 , \44566 , \44567 , \44568 , \44569 , \44570 , \44571 , \44572 ,
         \44573 , \44574 , \44575 , \44576 , \44577 , \44578 , \44579 , \44580 , \44581 , \44582 ,
         \44583 , \44584 , \44585 , \44586 , \44587 , \44588 , \44589 , \44590 , \44591 , \44592 ,
         \44593 , \44594 , \44595 , \44596 , \44597 , \44598 , \44599 , \44600 , \44601 , \44602 ,
         \44603 , \44604 , \44605 , \44606 , \44607 , \44608 , \44609 , \44610 , \44611 , \44612 ,
         \44613 , \44614 , \44615 , \44616 , \44617 , \44618 , \44619 , \44620 , \44621 , \44622 ,
         \44623 , \44624 , \44625 , \44626 , \44627 , \44628 , \44629 , \44630 , \44631 , \44632 ,
         \44633 , \44634 , \44635 , \44636 , \44637 , \44638 , \44639 , \44640 , \44641 , \44642 ,
         \44643 , \44644 , \44645 , \44646 , \44647 , \44648 , \44649 , \44650 , \44651 , \44652 ,
         \44653 , \44654 , \44655 , \44656 , \44657 , \44658 , \44659 , \44660 , \44661 , \44662 ,
         \44663 , \44664 , \44665 , \44666 , \44667 , \44668 , \44669 , \44670 , \44671 , \44672 ,
         \44673 , \44674 , \44675 , \44676 , \44677 , \44678 , \44679 , \44680 , \44681 , \44682 ,
         \44683 , \44684 , \44685 , \44686 , \44687 , \44688 , \44689 , \44690 , \44691 , \44692 ,
         \44693 , \44694 , \44695 , \44696 , \44697 , \44698 , \44699 , \44700 , \44701 , \44702 ,
         \44703 , \44704 , \44705 , \44706 , \44707 , \44708 , \44709 , \44710 , \44711 , \44712 ,
         \44713 , \44714 , \44715 , \44716 , \44717 , \44718 , \44719 , \44720 , \44721 , \44722 ,
         \44723 , \44724 , \44725 , \44726 , \44727 , \44728 , \44729 , \44730 , \44731 , \44732 ,
         \44733 , \44734 , \44735 , \44736 , \44737 , \44738 , \44739 , \44740 , \44741 , \44742 ,
         \44743 , \44744 , \44745 , \44746 , \44747 , \44748 , \44749 , \44750 , \44751 , \44752 ,
         \44753 , \44754 , \44755 , \44756 , \44757 , \44758 , \44759 , \44760 , \44761 , \44762 ,
         \44763 , \44764 , \44765 , \44766 , \44767 , \44768 , \44769 , \44770 , \44771 , \44772 ,
         \44773 , \44774 , \44775 , \44776 , \44777 , \44778 , \44779 , \44780 , \44781 , \44782 ,
         \44783 , \44784 , \44785 , \44786 , \44787 , \44788 , \44789 , \44790 , \44791 , \44792 ,
         \44793 , \44794 , \44795 , \44796 , \44797 , \44798 , \44799 , \44800 , \44801 , \44802 ,
         \44803 , \44804 , \44805 , \44806 , \44807 , \44808 , \44809 , \44810 , \44811 , \44812 ,
         \44813 , \44814 , \44815 , \44816 , \44817 , \44818 , \44819 , \44820 , \44821 , \44822 ,
         \44823 , \44824 , \44825 , \44826 , \44827 , \44828 , \44829 , \44830 , \44831 , \44832 ,
         \44833 , \44834 , \44835 , \44836 , \44837 , \44838 , \44839 , \44840 , \44841 , \44842 ,
         \44843 , \44844 , \44845 , \44846 , \44847 , \44848 , \44849 , \44850 , \44851 , \44852 ,
         \44853 , \44854 , \44855 , \44856 , \44857 , \44858 , \44859 , \44860 , \44861 , \44862 ,
         \44863 , \44864 , \44865 , \44866 , \44867 , \44868 , \44869 , \44870 , \44871 , \44872 ,
         \44873 , \44874 , \44875 , \44876 , \44877 , \44878 , \44879 , \44880 , \44881 , \44882 ,
         \44883 , \44884 , \44885 , \44886 , \44887 , \44888 , \44889 , \44890 , \44891 , \44892 ,
         \44893 , \44894 , \44895 , \44896 , \44897 , \44898 , \44899 , \44900 , \44901 , \44902 ,
         \44903 , \44904 , \44905 , \44906 , \44907 , \44908 , \44909 , \44910 , \44911 , \44912 ,
         \44913 , \44914 , \44915 , \44916 , \44917 , \44918 , \44919 , \44920 , \44921 , \44922 ,
         \44923 , \44924 , \44925 , \44926 , \44927 , \44928 , \44929 , \44930 , \44931 , \44932 ,
         \44933 , \44934 , \44935 , \44936 , \44937 , \44938 , \44939 , \44940 , \44941 , \44942 ,
         \44943 , \44944 , \44945 , \44946 , \44947 , \44948 , \44949 , \44950 , \44951 , \44952 ,
         \44953 , \44954 , \44955 , \44956 , \44957 , \44958 , \44959 , \44960 , \44961 , \44962 ,
         \44963 , \44964 , \44965 , \44966 , \44967 , \44968 , \44969 , \44970 , \44971 , \44972 ,
         \44973 , \44974 , \44975 , \44976 , \44977 , \44978 , \44979 , \44980 , \44981 , \44982 ,
         \44983 , \44984 , \44985 , \44986 , \44987 , \44988 , \44989 , \44990 , \44991 , \44992 ,
         \44993 , \44994 , \44995 , \44996 , \44997 , \44998 , \44999 , \45000 , \45001 , \45002 ,
         \45003 , \45004 , \45005 , \45006 , \45007 , \45008 , \45009 , \45010 , \45011 , \45012 ,
         \45013 , \45014 , \45015 , \45016 , \45017 , \45018 , \45019 , \45020 , \45021 , \45022 ,
         \45023 , \45024 , \45025 , \45026 , \45027 , \45028 , \45029 , \45030 , \45031 , \45032 ,
         \45033 , \45034 , \45035 , \45036 , \45037 , \45038 , \45039 , \45040 , \45041 , \45042 ,
         \45043 , \45044 , \45045 , \45046 , \45047 , \45048 , \45049 , \45050 , \45051 , \45052 ,
         \45053 , \45054 , \45055 , \45056 , \45057 , \45058 , \45059 , \45060 , \45061 , \45062 ,
         \45063 , \45064 , \45065 , \45066 , \45067 , \45068 , \45069 , \45070 , \45071 , \45072 ,
         \45073 , \45074 , \45075 , \45076 , \45077 , \45078 , \45079 , \45080 , \45081 , \45082 ,
         \45083 , \45084 , \45085 , \45086 , \45087 , \45088 , \45089 , \45090 , \45091 , \45092 ,
         \45093 , \45094 , \45095 , \45096 , \45097 , \45098 , \45099 , \45100 , \45101 , \45102 ,
         \45103 , \45104 , \45105 , \45106 , \45107 , \45108 , \45109 , \45110 , \45111 , \45112 ,
         \45113 , \45114 , \45115 , \45116 , \45117 , \45118 , \45119 , \45120 , \45121 , \45122 ,
         \45123 , \45124 , \45125 , \45126 , \45127 , \45128 , \45129 , \45130 , \45131 , \45132 ,
         \45133 , \45134 , \45135 , \45136 , \45137 , \45138 , \45139 , \45140 , \45141 , \45142 ,
         \45143 , \45144 , \45145 , \45146 , \45147 , \45148 , \45149 , \45150 , \45151 , \45152 ,
         \45153 , \45154 , \45155 , \45156 , \45157 , \45158 , \45159 , \45160 , \45161 , \45162 ,
         \45163 , \45164 , \45165 , \45166 , \45167 , \45168 , \45169 , \45170 , \45171 , \45172 ,
         \45173 , \45174 , \45175 , \45176 , \45177 , \45178 , \45179 , \45180 , \45181 , \45182 ,
         \45183 , \45184 , \45185 , \45186 , \45187 , \45188 , \45189 , \45190 , \45191 , \45192 ,
         \45193 , \45194 , \45195 , \45196 , \45197 , \45198 , \45199 , \45200 , \45201 , \45202 ,
         \45203 , \45204 , \45205 , \45206 , \45207 , \45208 , \45209 , \45210 , \45211 , \45212 ,
         \45213 , \45214 , \45215 , \45216 , \45217 , \45218 , \45219 , \45220 , \45221 , \45222 ,
         \45223 , \45224 , \45225 , \45226 , \45227 , \45228 , \45229 , \45230 , \45231 , \45232 ,
         \45233 , \45234 , \45235 , \45236 , \45237 , \45238 , \45239 , \45240 , \45241 , \45242 ,
         \45243 , \45244 , \45245 , \45246 , \45247 , \45248 , \45249 , \45250 , \45251 , \45252 ,
         \45253 , \45254 , \45255 , \45256 , \45257 , \45258 , \45259 , \45260 , \45261 , \45262 ,
         \45263 , \45264 , \45265 , \45266 , \45267 , \45268 , \45269 , \45270 , \45271 , \45272 ,
         \45273 , \45274 , \45275 , \45276 , \45277 , \45278 , \45279 , \45280 , \45281 , \45282 ,
         \45283 , \45284 , \45285 , \45286 , \45287 , \45288 , \45289 , \45290 , \45291 , \45292 ,
         \45293 , \45294 , \45295 , \45296 , \45297 , \45298 , \45299 , \45300 , \45301 , \45302 ,
         \45303 , \45304 , \45305 , \45306 , \45307 , \45308 , \45309 , \45310 , \45311 , \45312 ,
         \45313 , \45314 , \45315 , \45316 , \45317 , \45318 , \45319 , \45320 , \45321 , \45322 ,
         \45323 , \45324 , \45325 , \45326 , \45327 , \45328 , \45329 , \45330 , \45331 , \45332 ,
         \45333 , \45334 , \45335 , \45336 , \45337 , \45338 , \45339 , \45340 , \45341 , \45342 ,
         \45343 , \45344 , \45345 , \45346 , \45347 , \45348 , \45349 , \45350 , \45351 , \45352 ,
         \45353 , \45354 , \45355 , \45356 , \45357 , \45358 , \45359 , \45360 , \45361 , \45362 ,
         \45363 , \45364 , \45365 , \45366 , \45367 , \45368 , \45369 , \45370 , \45371 , \45372 ,
         \45373 , \45374 , \45375 , \45376 , \45377 , \45378 , \45379 , \45380 , \45381 , \45382 ,
         \45383 , \45384 , \45385 , \45386 , \45387 , \45388 , \45389 , \45390 , \45391 , \45392 ,
         \45393 , \45394 , \45395 , \45396 , \45397 , \45398 , \45399 , \45400 , \45401 , \45402 ,
         \45403 , \45404 , \45405 , \45406 , \45407 , \45408 , \45409 , \45410 , \45411 , \45412 ,
         \45413 , \45414 , \45415 , \45416 , \45417 , \45418 , \45419 , \45420 , \45421 , \45422 ,
         \45423 , \45424 , \45425 , \45426 , \45427 , \45428 , \45429 , \45430 , \45431 , \45432 ,
         \45433 , \45434 , \45435 , \45436 , \45437 , \45438 , \45439 , \45440 , \45441 , \45442 ,
         \45443 , \45444 , \45445 , \45446 , \45447 , \45448 , \45449 , \45450 , \45451 , \45452 ,
         \45453 , \45454 , \45455 , \45456 , \45457 , \45458 , \45459 , \45460 , \45461 , \45462 ,
         \45463 , \45464 , \45465 , \45466 , \45467 , \45468 , \45469 , \45470 , \45471 , \45472 ,
         \45473 , \45474 , \45475 , \45476 , \45477 , \45478 , \45479 , \45480 , \45481 , \45482 ,
         \45483 , \45484 , \45485 , \45486 , \45487 , \45488 , \45489 , \45490 , \45491 , \45492 ,
         \45493 , \45494 , \45495 , \45496 , \45497 , \45498 , \45499 , \45500 , \45501 , \45502 ,
         \45503 , \45504 , \45505 , \45506 , \45507 , \45508 , \45509 , \45510 , \45511 , \45512 ,
         \45513 , \45514 , \45515 , \45516 , \45517 , \45518 , \45519 , \45520 , \45521 , \45522 ,
         \45523 , \45524 , \45525 , \45526 , \45527 , \45528 , \45529 , \45530 , \45531 , \45532 ,
         \45533 , \45534 , \45535 , \45536 , \45537 , \45538 , \45539 , \45540 , \45541 , \45542 ,
         \45543 , \45544 , \45545 , \45546 , \45547 , \45548 , \45549 , \45550 , \45551 , \45552 ,
         \45553 , \45554 , \45555 , \45556 , \45557 , \45558 , \45559 , \45560 , \45561 , \45562 ,
         \45563 , \45564 , \45565 , \45566 , \45567 , \45568 , \45569 , \45570 , \45571 , \45572 ,
         \45573 , \45574 , \45575 , \45576 , \45577 , \45578 , \45579 , \45580 , \45581 , \45582 ,
         \45583 , \45584 , \45585 , \45586 , \45587 , \45588 , \45589 , \45590 , \45591 , \45592 ,
         \45593 , \45594 , \45595 , \45596 , \45597 , \45598 , \45599 , \45600 , \45601 , \45602 ,
         \45603 , \45604 , \45605 , \45606 , \45607 , \45608 , \45609 , \45610 , \45611 , \45612 ,
         \45613 , \45614 , \45615 , \45616 , \45617 , \45618 , \45619 , \45620 , \45621 , \45622 ,
         \45623 , \45624 , \45625 , \45626 , \45627 , \45628 , \45629 , \45630 , \45631 , \45632 ,
         \45633 , \45634 , \45635 , \45636 , \45637 , \45638 , \45639 , \45640 , \45641 , \45642 ,
         \45643 , \45644 , \45645 , \45646 , \45647 , \45648 , \45649 , \45650 , \45651 , \45652 ,
         \45653 , \45654 , \45655 , \45656 , \45657 , \45658 , \45659 , \45660 , \45661 , \45662 ,
         \45663 , \45664 , \45665 , \45666 , \45667 , \45668 , \45669 , \45670 , \45671 , \45672 ,
         \45673 , \45674 , \45675 , \45676 , \45677 , \45678 , \45679 , \45680 , \45681 , \45682 ,
         \45683 , \45684 , \45685 , \45686 , \45687 , \45688 , \45689 , \45690 , \45691 , \45692 ,
         \45693 , \45694 , \45695 , \45696 , \45697 , \45698 , \45699 , \45700 , \45701 , \45702 ,
         \45703 , \45704 , \45705 , \45706 , \45707 , \45708 , \45709 , \45710 , \45711 , \45712 ,
         \45713 , \45714 , \45715 , \45716 , \45717 , \45718 , \45719 , \45720 , \45721 , \45722 ,
         \45723 , \45724 , \45725 , \45726 , \45727 , \45728 , \45729 , \45730 , \45731 , \45732 ,
         \45733 , \45734 , \45735 , \45736 , \45737 , \45738 , \45739 , \45740 , \45741 , \45742 ,
         \45743 , \45744 , \45745 , \45746 , \45747 , \45748 , \45749 , \45750 , \45751 , \45752 ,
         \45753 , \45754 , \45755 , \45756 , \45757 , \45758 , \45759 , \45760 , \45761 , \45762 ,
         \45763 , \45764 , \45765 , \45766 , \45767 , \45768 , \45769 , \45770 , \45771 , \45772 ,
         \45773 , \45774 , \45775 , \45776 , \45777 , \45778 , \45779 , \45780 , \45781 , \45782 ,
         \45783 , \45784 , \45785 , \45786 , \45787 , \45788 , \45789 , \45790 , \45791 , \45792 ,
         \45793 , \45794 , \45795 , \45796 , \45797 , \45798 , \45799 , \45800 , \45801 , \45802 ,
         \45803 , \45804 , \45805 , \45806 , \45807 , \45808 , \45809 , \45810 , \45811 , \45812 ,
         \45813 , \45814 , \45815 , \45816 , \45817 , \45818 , \45819 , \45820 , \45821 , \45822 ,
         \45823 , \45824 , \45825 , \45826 , \45827 , \45828 , \45829 , \45830 , \45831 , \45832 ,
         \45833 , \45834 , \45835 , \45836 , \45837 , \45838 , \45839 , \45840 , \45841 , \45842 ,
         \45843 , \45844 , \45845 , \45846 , \45847 , \45848 , \45849 , \45850 , \45851 , \45852 ,
         \45853 , \45854 , \45855 , \45856 , \45857 , \45858 , \45859 , \45860 , \45861 , \45862 ,
         \45863 , \45864 , \45865 , \45866 , \45867 , \45868 , \45869 , \45870 , \45871 , \45872 ,
         \45873 , \45874 , \45875 , \45876 , \45877 , \45878 , \45879 , \45880 , \45881 , \45882 ,
         \45883 , \45884 , \45885 , \45886 , \45887 , \45888 , \45889 , \45890 , \45891 , \45892 ,
         \45893 , \45894 , \45895 , \45896 , \45897 , \45898 , \45899 , \45900 , \45901 , \45902 ,
         \45903 , \45904 , \45905 , \45906 , \45907 , \45908 , \45909 , \45910 , \45911 , \45912 ,
         \45913 , \45914 , \45915 , \45916 , \45917 , \45918 , \45919 , \45920 , \45921 , \45922 ,
         \45923 , \45924 , \45925 , \45926 , \45927 , \45928 , \45929 , \45930 , \45931 , \45932 ,
         \45933 , \45934 , \45935 , \45936 , \45937 , \45938 , \45939 , \45940 , \45941 , \45942 ,
         \45943 , \45944 , \45945 , \45946 , \45947 , \45948 , \45949 , \45950 , \45951 , \45952 ,
         \45953 , \45954 , \45955 , \45956 , \45957 , \45958 , \45959 , \45960 , \45961 , \45962 ,
         \45963 , \45964 , \45965 , \45966 , \45967 , \45968 , \45969 , \45970 , \45971 , \45972 ,
         \45973 , \45974 , \45975 , \45976 , \45977 , \45978 , \45979 , \45980 , \45981 , \45982 ,
         \45983 , \45984 , \45985 , \45986 , \45987 , \45988 , \45989 , \45990 , \45991 , \45992 ,
         \45993 , \45994 , \45995 , \45996 , \45997 , \45998 , \45999 , \46000 , \46001 , \46002 ,
         \46003 , \46004 , \46005 , \46006 , \46007 , \46008 , \46009 , \46010 , \46011 , \46012 ,
         \46013 , \46014 , \46015 , \46016 , \46017 , \46018 , \46019 , \46020 , \46021 , \46022 ,
         \46023 , \46024 , \46025 , \46026 , \46027 , \46028 , \46029 , \46030 , \46031 , \46032 ,
         \46033 , \46034 , \46035 , \46036 , \46037 , \46038 , \46039 , \46040 , \46041 , \46042 ,
         \46043 , \46044 , \46045 , \46046 , \46047 , \46048 , \46049 , \46050 , \46051 , \46052 ,
         \46053 , \46054 , \46055 , \46056 , \46057 , \46058 , \46059 , \46060 , \46061 , \46062 ,
         \46063 , \46064 , \46065 , \46066 , \46067 , \46068 , \46069 , \46070 , \46071 , \46072 ,
         \46073 , \46074 , \46075 , \46076 , \46077 , \46078 , \46079 , \46080 , \46081 , \46082 ,
         \46083 , \46084 , \46085 , \46086 , \46087 , \46088 , \46089 , \46090 , \46091 , \46092 ,
         \46093 , \46094 , \46095 , \46096 , \46097 , \46098 , \46099 , \46100 , \46101 , \46102 ,
         \46103 , \46104 , \46105 , \46106 , \46107 , \46108 , \46109 , \46110 , \46111 , \46112 ,
         \46113 , \46114 , \46115 , \46116 , \46117 , \46118 , \46119 , \46120 , \46121 , \46122 ,
         \46123 , \46124 , \46125 , \46126 , \46127 , \46128 , \46129 , \46130 , \46131 , \46132 ,
         \46133 , \46134 , \46135 , \46136 , \46137 , \46138 , \46139 , \46140 , \46141 , \46142 ,
         \46143 , \46144 , \46145 , \46146 , \46147 , \46148 , \46149 , \46150 , \46151 , \46152 ,
         \46153 , \46154 , \46155 , \46156 , \46157 , \46158 , \46159 , \46160 , \46161 , \46162 ,
         \46163 , \46164 , \46165 , \46166 , \46167 , \46168 , \46169 , \46170 , \46171 , \46172 ,
         \46173 , \46174 , \46175 , \46176 , \46177 , \46178 , \46179 , \46180 , \46181 , \46182 ,
         \46183 , \46184 , \46185 , \46186 , \46187 , \46188 , \46189 , \46190 , \46191 , \46192 ,
         \46193 , \46194 , \46195 , \46196 , \46197 , \46198 , \46199 , \46200 , \46201 , \46202 ,
         \46203 , \46204 , \46205 , \46206 , \46207 , \46208 , \46209 , \46210 , \46211 , \46212 ,
         \46213 , \46214 , \46215 , \46216 , \46217 , \46218 , \46219 , \46220 , \46221 , \46222 ,
         \46223 , \46224 , \46225 , \46226 , \46227 , \46228 , \46229 , \46230 , \46231 , \46232 ,
         \46233 , \46234 , \46235 , \46236 , \46237 , \46238 , \46239 , \46240 , \46241 , \46242 ,
         \46243 , \46244 , \46245 , \46246 , \46247 , \46248 , \46249 , \46250 , \46251 , \46252 ,
         \46253 , \46254 , \46255 , \46256 , \46257 , \46258 , \46259 , \46260 , \46261 , \46262 ,
         \46263 , \46264 , \46265 , \46266 , \46267 , \46268 , \46269 , \46270 , \46271 , \46272 ,
         \46273 , \46274 , \46275 , \46276 , \46277 , \46278 , \46279 , \46280 , \46281 , \46282 ,
         \46283 , \46284 , \46285 , \46286 , \46287 , \46288 , \46289 , \46290 , \46291 , \46292 ,
         \46293 , \46294 , \46295 , \46296 , \46297 , \46298 , \46299 , \46300 , \46301 , \46302 ,
         \46303 , \46304 , \46305 , \46306 , \46307 , \46308 , \46309 , \46310 , \46311 , \46312 ,
         \46313 , \46314 , \46315 , \46316 , \46317 , \46318 , \46319 , \46320 , \46321 , \46322 ,
         \46323 , \46324 , \46325 , \46326 , \46327 , \46328 , \46329 , \46330 , \46331 , \46332 ,
         \46333 , \46334 , \46335 , \46336 , \46337 , \46338 , \46339 , \46340 , \46341 , \46342 ,
         \46343 , \46344 , \46345 , \46346 , \46347 , \46348 , \46349 , \46350 , \46351 , \46352 ,
         \46353 , \46354 , \46355 , \46356 , \46357 , \46358 , \46359 , \46360 , \46361 , \46362 ,
         \46363 , \46364 , \46365 , \46366 , \46367 , \46368 , \46369 , \46370 , \46371 , \46372 ,
         \46373 , \46374 , \46375 , \46376 , \46377 , \46378 , \46379 , \46380 , \46381 , \46382 ,
         \46383 , \46384 , \46385 , \46386 , \46387 , \46388 , \46389 , \46390 , \46391 , \46392 ,
         \46393 , \46394 , \46395 , \46396 , \46397 , \46398 , \46399 , \46400 , \46401 , \46402 ,
         \46403 , \46404 , \46405 , \46406 , \46407 , \46408 , \46409 , \46410 , \46411 , \46412 ,
         \46413 , \46414 , \46415 , \46416 , \46417 , \46418 , \46419 , \46420 , \46421 , \46422 ,
         \46423 , \46424 , \46425 , \46426 , \46427 , \46428 , \46429 , \46430 , \46431 , \46432 ,
         \46433 , \46434 , \46435 , \46436 , \46437 , \46438 , \46439 , \46440 , \46441 , \46442 ,
         \46443 , \46444 , \46445 , \46446 , \46447 , \46448 , \46449 , \46450 , \46451 , \46452 ,
         \46453 , \46454 , \46455 , \46456 , \46457 , \46458 , \46459 , \46460 , \46461 , \46462 ,
         \46463 , \46464 , \46465 , \46466 , \46467 , \46468 , \46469 , \46470 , \46471 , \46472 ,
         \46473 , \46474 , \46475 , \46476 , \46477 , \46478 , \46479 , \46480 , \46481 , \46482 ,
         \46483 , \46484 , \46485 , \46486 , \46487 , \46488 , \46489 , \46490 , \46491 , \46492 ,
         \46493 , \46494 , \46495 , \46496 , \46497 , \46498 , \46499 , \46500 , \46501 , \46502 ,
         \46503 , \46504 , \46505 , \46506 , \46507 , \46508 , \46509 , \46510 , \46511 , \46512 ,
         \46513 , \46514 , \46515 , \46516 , \46517 , \46518 , \46519 , \46520 , \46521 , \46522 ,
         \46523 , \46524 , \46525 , \46526 , \46527 , \46528 , \46529 , \46530 , \46531 , \46532 ,
         \46533 , \46534 , \46535 , \46536 , \46537 , \46538 , \46539 , \46540 , \46541 , \46542 ,
         \46543 , \46544 , \46545 , \46546 , \46547 , \46548 , \46549 , \46550 , \46551 , \46552 ,
         \46553 , \46554 , \46555 , \46556 , \46557 , \46558 , \46559 , \46560 , \46561 , \46562 ,
         \46563 , \46564 , \46565 , \46566 , \46567 , \46568 , \46569 , \46570 , \46571 , \46572 ,
         \46573 , \46574 , \46575 , \46576 , \46577 , \46578 , \46579 , \46580 , \46581 , \46582 ,
         \46583 , \46584 , \46585 , \46586 , \46587 , \46588 , \46589 , \46590 , \46591 , \46592 ,
         \46593 , \46594 , \46595 , \46596 , \46597 , \46598 , \46599 , \46600 , \46601 , \46602 ,
         \46603 , \46604 , \46605 , \46606 , \46607 , \46608 , \46609 , \46610 , \46611 , \46612 ,
         \46613 , \46614 , \46615 , \46616 , \46617 , \46618 , \46619 , \46620 , \46621 , \46622 ,
         \46623 , \46624 , \46625 , \46626 , \46627 , \46628 , \46629 , \46630 , \46631 , \46632 ,
         \46633 , \46634 , \46635 , \46636 , \46637 , \46638 , \46639 , \46640 , \46641 , \46642 ,
         \46643 , \46644 , \46645 , \46646 , \46647 , \46648 , \46649 , \46650 , \46651 , \46652 ,
         \46653 , \46654 , \46655 , \46656 , \46657 , \46658 , \46659 , \46660 , \46661 , \46662 ,
         \46663 , \46664 , \46665 , \46666 , \46667 , \46668 , \46669 , \46670 , \46671 , \46672 ,
         \46673 , \46674 , \46675 , \46676 , \46677 , \46678 , \46679 , \46680 , \46681 , \46682 ,
         \46683 , \46684 , \46685 , \46686 , \46687 , \46688 , \46689 , \46690 , \46691 , \46692 ,
         \46693 , \46694 , \46695 , \46696 , \46697 , \46698 , \46699 , \46700 , \46701 , \46702 ,
         \46703 , \46704 , \46705 , \46706 , \46707 , \46708 , \46709 , \46710 , \46711 , \46712 ,
         \46713 , \46714 , \46715 , \46716 , \46717 , \46718 , \46719 , \46720 , \46721 , \46722 ,
         \46723 , \46724 , \46725 , \46726 , \46727 , \46728 , \46729 , \46730 , \46731 , \46732 ,
         \46733 , \46734 , \46735 , \46736 , \46737 , \46738 , \46739 , \46740 , \46741 , \46742 ,
         \46743 , \46744 , \46745 , \46746 , \46747 , \46748 , \46749 , \46750 , \46751 , \46752 ,
         \46753 , \46754 , \46755 , \46756 , \46757 , \46758 , \46759 , \46760 , \46761 , \46762 ,
         \46763 , \46764 , \46765 , \46766 , \46767 , \46768 , \46769 , \46770 , \46771 , \46772 ,
         \46773 , \46774 , \46775 , \46776 , \46777 , \46778 , \46779 , \46780 , \46781 , \46782 ,
         \46783 , \46784 , \46785 , \46786 , \46787 , \46788 , \46789 , \46790 , \46791 , \46792 ,
         \46793 , \46794 , \46795 , \46796 , \46797 , \46798 , \46799 , \46800 , \46801 , \46802 ,
         \46803 , \46804 , \46805 , \46806 , \46807 , \46808 , \46809 , \46810 , \46811 , \46812 ,
         \46813 , \46814 , \46815 , \46816 , \46817 , \46818 , \46819 , \46820 , \46821 , \46822 ,
         \46823 , \46824 , \46825 , \46826 , \46827 , \46828 , \46829 , \46830 , \46831 , \46832 ,
         \46833 , \46834 , \46835 , \46836 , \46837 , \46838 , \46839 , \46840 , \46841 , \46842 ,
         \46843 , \46844 , \46845 , \46846 , \46847 , \46848 , \46849 , \46850 , \46851 , \46852 ,
         \46853 , \46854 , \46855 , \46856 , \46857 , \46858 , \46859 , \46860 , \46861 , \46862 ,
         \46863 , \46864 , \46865 , \46866 , \46867 , \46868 , \46869 , \46870 , \46871 , \46872 ,
         \46873 , \46874 , \46875 , \46876 , \46877 , \46878 , \46879 , \46880 , \46881 , \46882 ,
         \46883 , \46884 , \46885 , \46886 , \46887 , \46888 , \46889 , \46890 , \46891 , \46892 ,
         \46893 , \46894 , \46895 , \46896 , \46897 , \46898 , \46899 , \46900 , \46901 , \46902 ,
         \46903 , \46904 , \46905 , \46906 , \46907 , \46908 , \46909 , \46910 , \46911 , \46912 ,
         \46913 , \46914 , \46915 , \46916 , \46917 , \46918 , \46919 , \46920 , \46921 , \46922 ,
         \46923 , \46924 , \46925 , \46926 , \46927 , \46928 , \46929 , \46930 , \46931 , \46932 ,
         \46933 , \46934 , \46935 , \46936 , \46937 , \46938 , \46939 , \46940 , \46941 , \46942 ,
         \46943 , \46944 , \46945 , \46946 , \46947 , \46948 , \46949 , \46950 , \46951 , \46952 ,
         \46953 , \46954 , \46955 , \46956 , \46957 , \46958 , \46959 , \46960 , \46961 , \46962 ,
         \46963 , \46964 , \46965 , \46966 , \46967 , \46968 , \46969 , \46970 , \46971 , \46972 ,
         \46973 , \46974 , \46975 , \46976 , \46977 , \46978 , \46979 , \46980 , \46981 , \46982 ,
         \46983 , \46984 , \46985 , \46986 , \46987 , \46988 , \46989 , \46990 , \46991 , \46992 ,
         \46993 , \46994 , \46995 , \46996 , \46997 , \46998 , \46999 , \47000 , \47001 , \47002 ,
         \47003 , \47004 , \47005 , \47006 , \47007 , \47008 , \47009 , \47010 , \47011 , \47012 ,
         \47013 , \47014 , \47015 , \47016 , \47017 , \47018 , \47019 , \47020 , \47021 , \47022 ,
         \47023 , \47024 , \47025 , \47026 , \47027 , \47028 , \47029 , \47030 , \47031 , \47032 ,
         \47033 , \47034 , \47035 , \47036 , \47037 , \47038 , \47039 , \47040 , \47041 , \47042 ,
         \47043 , \47044 , \47045 , \47046 , \47047 , \47048 , \47049 , \47050 , \47051 , \47052 ,
         \47053 , \47054 , \47055 , \47056 , \47057 , \47058 , \47059 , \47060 , \47061 , \47062 ,
         \47063 , \47064 , \47065 , \47066 , \47067 , \47068 , \47069 , \47070 , \47071 , \47072 ,
         \47073 , \47074 , \47075 , \47076 , \47077 , \47078 , \47079 , \47080 , \47081 , \47082 ,
         \47083 , \47084 , \47085 , \47086 , \47087 , \47088 , \47089 , \47090 , \47091 , \47092 ,
         \47093 , \47094 , \47095 , \47096 , \47097 , \47098 , \47099 , \47100 , \47101 , \47102 ,
         \47103 , \47104 , \47105 , \47106 , \47107 , \47108 , \47109 , \47110 , \47111 , \47112 ,
         \47113 , \47114 , \47115 , \47116 , \47117 , \47118 , \47119 , \47120 , \47121 , \47122 ,
         \47123 , \47124 , \47125 , \47126 , \47127 , \47128 , \47129 , \47130 , \47131 , \47132 ,
         \47133 , \47134 , \47135 , \47136 , \47137 , \47138 , \47139 , \47140 , \47141 , \47142 ,
         \47143 , \47144 , \47145 , \47146 , \47147 , \47148 , \47149 , \47150 , \47151 , \47152 ,
         \47153 , \47154 , \47155 , \47156 , \47157 , \47158 , \47159 , \47160 , \47161 , \47162 ,
         \47163 , \47164 , \47165 , \47166 , \47167 , \47168 , \47169 , \47170 , \47171 , \47172 ,
         \47173 , \47174 , \47175 , \47176 , \47177 , \47178 , \47179 , \47180 , \47181 , \47182 ,
         \47183 , \47184 , \47185 , \47186 , \47187 , \47188 , \47189 , \47190 , \47191 , \47192 ,
         \47193 , \47194 , \47195 , \47196 , \47197 , \47198 , \47199 , \47200 , \47201 , \47202 ,
         \47203 , \47204 , \47205 , \47206 , \47207 , \47208 , \47209 , \47210 , \47211 , \47212 ,
         \47213 , \47214 , \47215 , \47216 , \47217 , \47218 , \47219 , \47220 , \47221 , \47222 ,
         \47223 , \47224 , \47225 , \47226 , \47227 , \47228 , \47229 , \47230 , \47231 , \47232 ,
         \47233 , \47234 , \47235 , \47236 , \47237 , \47238 , \47239 , \47240 , \47241 , \47242 ,
         \47243 , \47244 , \47245 , \47246 , \47247 , \47248 , \47249 , \47250 , \47251 , \47252 ,
         \47253 , \47254 , \47255 , \47256 , \47257 , \47258 , \47259 , \47260 , \47261 , \47262 ,
         \47263 , \47264 , \47265 , \47266 , \47267 , \47268 , \47269 , \47270 , \47271 , \47272 ,
         \47273 , \47274 , \47275 , \47276 , \47277 , \47278 , \47279 , \47280 , \47281 , \47282 ,
         \47283 , \47284 , \47285 , \47286 , \47287 , \47288 , \47289 , \47290 , \47291 , \47292 ,
         \47293 , \47294 , \47295 , \47296 , \47297 , \47298 , \47299 , \47300 , \47301 , \47302 ,
         \47303 , \47304 , \47305 , \47306 , \47307 , \47308 , \47309 , \47310 , \47311 , \47312 ,
         \47313 , \47314 , \47315 , \47316 , \47317 , \47318 , \47319 , \47320 , \47321 , \47322 ,
         \47323 , \47324 , \47325 , \47326 , \47327 , \47328 , \47329 , \47330 , \47331 , \47332 ,
         \47333 , \47334 , \47335 , \47336 , \47337 , \47338 , \47339 , \47340 , \47341 , \47342 ,
         \47343 , \47344 , \47345 , \47346 , \47347 , \47348 , \47349 , \47350 , \47351 , \47352 ,
         \47353 , \47354 , \47355 , \47356 , \47357 , \47358 , \47359 , \47360 , \47361 , \47362 ,
         \47363 , \47364 , \47365 , \47366 , \47367 , \47368 , \47369 , \47370 , \47371 , \47372 ,
         \47373 , \47374 , \47375 , \47376 , \47377 , \47378 , \47379 , \47380 , \47381 , \47382 ,
         \47383 , \47384 , \47385 , \47386 , \47387 , \47388 , \47389 , \47390 , \47391 , \47392 ,
         \47393 , \47394 , \47395 , \47396 , \47397 , \47398 , \47399 , \47400 , \47401 , \47402 ,
         \47403 , \47404 , \47405 , \47406 , \47407 , \47408 , \47409 , \47410 , \47411 , \47412 ,
         \47413 , \47414 , \47415 , \47416 , \47417 , \47418 , \47419 , \47420 , \47421 , \47422 ,
         \47423 , \47424 , \47425 , \47426 , \47427 , \47428 , \47429 , \47430 , \47431 , \47432 ,
         \47433 , \47434 , \47435 , \47436 , \47437 , \47438 , \47439 , \47440 , \47441 , \47442 ,
         \47443 , \47444 , \47445 , \47446 , \47447 , \47448 , \47449 , \47450 , \47451 , \47452 ,
         \47453 , \47454 , \47455 , \47456 , \47457 , \47458 , \47459 , \47460 , \47461 , \47462 ,
         \47463 , \47464 , \47465 , \47466 , \47467 , \47468 , \47469 , \47470 , \47471 , \47472 ,
         \47473 , \47474 , \47475 , \47476 , \47477 , \47478 , \47479 , \47480 , \47481 , \47482 ,
         \47483 , \47484 , \47485 , \47486 , \47487 , \47488 , \47489 , \47490 , \47491 , \47492 ,
         \47493 , \47494 , \47495 , \47496 , \47497 , \47498 , \47499 , \47500 , \47501 , \47502 ,
         \47503 , \47504 , \47505 , \47506 , \47507 , \47508 , \47509 , \47510 , \47511 , \47512 ,
         \47513 , \47514 , \47515 , \47516 , \47517 , \47518 , \47519 , \47520 , \47521 , \47522 ,
         \47523 , \47524 , \47525 , \47526 , \47527 , \47528 , \47529 , \47530 , \47531 , \47532 ,
         \47533 , \47534 , \47535 , \47536 , \47537 , \47538 , \47539 , \47540 , \47541 , \47542 ,
         \47543 , \47544 , \47545 , \47546 , \47547 , \47548 , \47549 , \47550 , \47551 , \47552 ,
         \47553 , \47554 , \47555 , \47556 , \47557 , \47558 , \47559 , \47560 , \47561 , \47562 ,
         \47563 , \47564 , \47565 , \47566 , \47567 , \47568 , \47569 , \47570 , \47571 , \47572 ,
         \47573 , \47574 , \47575 , \47576 , \47577 , \47578 , \47579 , \47580 , \47581 , \47582 ,
         \47583 , \47584 , \47585 , \47586 , \47587 , \47588 , \47589 , \47590 , \47591 , \47592 ,
         \47593 , \47594 , \47595 , \47596 , \47597 , \47598 , \47599 , \47600 , \47601 , \47602 ,
         \47603 , \47604 , \47605 , \47606 , \47607 , \47608 , \47609 , \47610 , \47611 , \47612 ,
         \47613 , \47614 , \47615 , \47616 , \47617 , \47618 , \47619 , \47620 , \47621 , \47622 ,
         \47623 , \47624 , \47625 , \47626 , \47627 , \47628 , \47629 , \47630 , \47631 , \47632 ,
         \47633 , \47634 , \47635 , \47636 , \47637 , \47638 , \47639 , \47640 , \47641 , \47642 ,
         \47643 , \47644 , \47645 , \47646 , \47647 , \47648 , \47649 , \47650 , \47651 , \47652 ,
         \47653 , \47654 , \47655 , \47656 , \47657 , \47658 , \47659 , \47660 , \47661 , \47662 ,
         \47663 , \47664 , \47665 , \47666 , \47667 , \47668 , \47669 , \47670 , \47671 , \47672 ,
         \47673 , \47674 , \47675 , \47676 , \47677 , \47678 , \47679 , \47680 , \47681 , \47682 ,
         \47683 , \47684 , \47685 , \47686 , \47687 , \47688 , \47689 , \47690 , \47691 , \47692 ,
         \47693 , \47694 , \47695 , \47696 , \47697 , \47698 , \47699 , \47700 , \47701 , \47702 ,
         \47703 , \47704 , \47705 , \47706 , \47707 , \47708 , \47709 , \47710 , \47711 , \47712 ,
         \47713 , \47714 , \47715 , \47716 , \47717 , \47718 , \47719 , \47720 , \47721 , \47722 ,
         \47723 , \47724 , \47725 , \47726 , \47727 , \47728 , \47729 , \47730 , \47731 , \47732 ,
         \47733 , \47734 , \47735 , \47736 , \47737 , \47738 , \47739 , \47740 , \47741 , \47742 ,
         \47743 , \47744 , \47745 , \47746 , \47747 , \47748 , \47749 , \47750 , \47751 , \47752 ,
         \47753 , \47754 , \47755 , \47756 , \47757 , \47758 , \47759 , \47760 , \47761 , \47762 ,
         \47763 , \47764 , \47765 , \47766 , \47767 , \47768 , \47769 , \47770 , \47771 , \47772 ,
         \47773 , \47774 , \47775 , \47776 , \47777 , \47778 , \47779 , \47780 , \47781 , \47782 ,
         \47783 , \47784 , \47785 , \47786 , \47787 , \47788 , \47789 , \47790 , \47791 , \47792 ,
         \47793 , \47794 , \47795 , \47796 , \47797 , \47798 , \47799 , \47800 , \47801 , \47802 ,
         \47803 , \47804 , \47805 , \47806 , \47807 , \47808 , \47809 , \47810 , \47811 , \47812 ,
         \47813 , \47814 , \47815 , \47816 , \47817 , \47818 , \47819 , \47820 , \47821 , \47822 ,
         \47823 , \47824 , \47825 , \47826 , \47827 , \47828 , \47829 , \47830 , \47831 , \47832 ,
         \47833 , \47834 , \47835 , \47836 , \47837 , \47838 , \47839 , \47840 , \47841 , \47842 ,
         \47843 , \47844 , \47845 , \47846 , \47847 , \47848 , \47849 , \47850 , \47851 , \47852 ,
         \47853 , \47854 , \47855 , \47856 , \47857 , \47858 , \47859 , \47860 , \47861 , \47862 ,
         \47863 , \47864 , \47865 , \47866 , \47867 , \47868 , \47869 , \47870 , \47871 , \47872 ,
         \47873 , \47874 , \47875 , \47876 , \47877 , \47878 , \47879 , \47880 , \47881 , \47882 ,
         \47883 , \47884 , \47885 , \47886 , \47887 , \47888 , \47889 , \47890 , \47891 , \47892 ,
         \47893 , \47894 , \47895 , \47896 , \47897 , \47898 , \47899 , \47900 , \47901 , \47902 ,
         \47903 , \47904 , \47905 , \47906 , \47907 , \47908 , \47909 , \47910 , \47911 , \47912 ,
         \47913 , \47914 , \47915 , \47916 , \47917 , \47918 , \47919 , \47920 , \47921 , \47922 ,
         \47923 , \47924 , \47925 , \47926 , \47927 , \47928 , \47929 , \47930 , \47931 , \47932 ,
         \47933 , \47934 , \47935 , \47936 , \47937 , \47938 , \47939 , \47940 , \47941 , \47942 ,
         \47943 , \47944 , \47945 , \47946 , \47947 , \47948 , \47949 , \47950 , \47951 , \47952 ,
         \47953 , \47954 , \47955 , \47956 , \47957 , \47958 , \47959 , \47960 , \47961 , \47962 ,
         \47963 , \47964 , \47965 , \47966 , \47967 , \47968 , \47969 , \47970 , \47971 , \47972 ,
         \47973 , \47974 , \47975 , \47976 , \47977 , \47978 , \47979 , \47980 , \47981 , \47982 ,
         \47983 , \47984 , \47985 , \47986 , \47987 , \47988 , \47989 , \47990 , \47991 , \47992 ,
         \47993 , \47994 , \47995 , \47996 , \47997 , \47998 , \47999 , \48000 , \48001 , \48002 ,
         \48003 , \48004 , \48005 , \48006 , \48007 , \48008 , \48009 , \48010 , \48011 , \48012 ,
         \48013 , \48014 , \48015 , \48016 , \48017 , \48018 , \48019 , \48020 , \48021 , \48022 ,
         \48023 , \48024 , \48025 , \48026 , \48027 , \48028 , \48029 , \48030 , \48031 , \48032 ,
         \48033 , \48034 , \48035 , \48036 , \48037 , \48038 , \48039 , \48040 , \48041 , \48042 ,
         \48043 , \48044 , \48045 , \48046 , \48047 , \48048 , \48049 , \48050 , \48051 , \48052 ,
         \48053 , \48054 , \48055 , \48056 , \48057 , \48058 , \48059 , \48060 , \48061 , \48062 ,
         \48063 , \48064 , \48065 , \48066 , \48067 , \48068 , \48069 , \48070 , \48071 , \48072 ,
         \48073 , \48074 , \48075 , \48076 , \48077 , \48078 , \48079 , \48080 , \48081 , \48082 ,
         \48083 , \48084 , \48085 , \48086 , \48087 , \48088 , \48089 , \48090 , \48091 , \48092 ,
         \48093 , \48094 , \48095 , \48096 , \48097 , \48098 , \48099 , \48100 , \48101 , \48102 ,
         \48103 , \48104 , \48105 , \48106 , \48107 , \48108 , \48109 , \48110 , \48111 , \48112 ,
         \48113 , \48114 , \48115 , \48116 , \48117 , \48118 , \48119 , \48120 , \48121 , \48122 ,
         \48123 , \48124 , \48125 , \48126 , \48127 , \48128 , \48129 , \48130 , \48131 , \48132 ,
         \48133 , \48134 , \48135 , \48136 , \48137 , \48138 , \48139 , \48140 , \48141 , \48142 ,
         \48143 , \48144 , \48145 , \48146 , \48147 , \48148 , \48149 , \48150 , \48151 , \48152 ,
         \48153 , \48154 , \48155 , \48156 , \48157 , \48158 , \48159 , \48160 , \48161 , \48162 ,
         \48163 , \48164 , \48165 , \48166 , \48167 , \48168 , \48169 , \48170 , \48171 , \48172 ,
         \48173 , \48174 , \48175 , \48176 , \48177 , \48178 , \48179 , \48180 , \48181 , \48182 ,
         \48183 , \48184 , \48185 , \48186 , \48187 , \48188 , \48189 , \48190 , \48191 , \48192 ,
         \48193 , \48194 , \48195 , \48196 , \48197 , \48198 , \48199 , \48200 , \48201 , \48202 ,
         \48203 , \48204 , \48205 , \48206 , \48207 , \48208 , \48209 , \48210 , \48211 , \48212 ,
         \48213 , \48214 , \48215 , \48216 , \48217 , \48218 , \48219 , \48220 , \48221 , \48222 ,
         \48223 , \48224 , \48225 , \48226 , \48227 , \48228 , \48229 , \48230 , \48231 , \48232 ,
         \48233 , \48234 , \48235 , \48236 , \48237 , \48238 , \48239 , \48240 , \48241 , \48242 ,
         \48243 , \48244 , \48245 , \48246 , \48247 , \48248 , \48249 , \48250 , \48251 , \48252 ,
         \48253 , \48254 , \48255 , \48256 , \48257 , \48258 , \48259 , \48260 , \48261 , \48262 ,
         \48263 , \48264 , \48265 , \48266 , \48267 , \48268 , \48269 , \48270 , \48271 , \48272 ,
         \48273 , \48274 , \48275 , \48276 , \48277 , \48278 , \48279 , \48280 , \48281 , \48282 ,
         \48283 , \48284 , \48285 , \48286 , \48287 , \48288 , \48289 , \48290 , \48291 , \48292 ,
         \48293 , \48294 , \48295 , \48296 , \48297 , \48298 , \48299 , \48300 , \48301 , \48302 ,
         \48303 , \48304 , \48305 , \48306 , \48307 , \48308 , \48309 , \48310 , \48311 , \48312 ,
         \48313 , \48314 , \48315 , \48316 , \48317 , \48318 , \48319 , \48320 , \48321 , \48322 ,
         \48323 , \48324 , \48325 , \48326 , \48327 , \48328 , \48329 , \48330 , \48331 , \48332 ,
         \48333 , \48334 , \48335 , \48336 , \48337 , \48338 , \48339 , \48340 , \48341 , \48342 ,
         \48343 , \48344 , \48345 , \48346 , \48347 , \48348 , \48349 , \48350 , \48351 , \48352 ,
         \48353 , \48354 , \48355 , \48356 , \48357 , \48358 , \48359 , \48360 , \48361 , \48362 ,
         \48363 , \48364 , \48365 , \48366 , \48367 , \48368 , \48369 , \48370 , \48371 , \48372 ,
         \48373 , \48374 , \48375 , \48376 , \48377 , \48378 , \48379 , \48380 , \48381 , \48382 ,
         \48383 , \48384 , \48385 , \48386 , \48387 , \48388 , \48389 , \48390 , \48391 , \48392 ,
         \48393 , \48394 , \48395 , \48396 , \48397 , \48398 , \48399 , \48400 , \48401 , \48402 ,
         \48403 , \48404 , \48405 , \48406 , \48407 , \48408 , \48409 , \48410 , \48411 , \48412 ,
         \48413 , \48414 , \48415 , \48416 , \48417 , \48418 , \48419 , \48420 , \48421 , \48422 ,
         \48423 , \48424 , \48425 , \48426 , \48427 , \48428 , \48429 , \48430 , \48431 , \48432 ,
         \48433 , \48434 , \48435 , \48436 , \48437 , \48438 , \48439 , \48440 , \48441 , \48442 ,
         \48443 , \48444 , \48445 , \48446 , \48447 , \48448 , \48449 , \48450 , \48451 , \48452 ,
         \48453 , \48454 , \48455 , \48456 , \48457 , \48458 , \48459 , \48460 , \48461 , \48462 ,
         \48463 , \48464 , \48465 , \48466 , \48467 , \48468 , \48469 , \48470 , \48471 , \48472 ,
         \48473 , \48474 , \48475 , \48476 , \48477 , \48478 , \48479 , \48480 , \48481 , \48482 ,
         \48483 , \48484 , \48485 , \48486 , \48487 , \48488 , \48489 , \48490 , \48491 , \48492 ,
         \48493 , \48494 , \48495 , \48496 , \48497 , \48498 , \48499 , \48500 , \48501 , \48502 ,
         \48503 , \48504 , \48505 , \48506 , \48507 , \48508 , \48509 , \48510 , \48511 , \48512 ,
         \48513 , \48514 , \48515 , \48516 , \48517 , \48518 , \48519 , \48520 , \48521 , \48522 ,
         \48523 , \48524 , \48525 , \48526 , \48527 , \48528 , \48529 , \48530 , \48531 , \48532 ,
         \48533 , \48534 , \48535 , \48536 , \48537 , \48538 , \48539 , \48540 , \48541 , \48542 ,
         \48543 , \48544 , \48545 , \48546 , \48547 , \48548 , \48549 , \48550 , \48551 , \48552 ,
         \48553 , \48554 , \48555 , \48556 , \48557 , \48558 , \48559 , \48560 , \48561 , \48562 ,
         \48563 , \48564 , \48565 , \48566 , \48567 , \48568 , \48569 , \48570 , \48571 , \48572 ,
         \48573 , \48574 , \48575 , \48576 , \48577 , \48578 , \48579 , \48580 , \48581 , \48582 ,
         \48583 , \48584 , \48585 , \48586 , \48587 , \48588 , \48589 , \48590 , \48591 , \48592 ,
         \48593 , \48594 , \48595 , \48596 , \48597 , \48598 , \48599 , \48600 , \48601 , \48602 ,
         \48603 , \48604 , \48605 , \48606 , \48607 , \48608 , \48609 , \48610 , \48611 , \48612 ,
         \48613 , \48614 , \48615 , \48616 , \48617 , \48618 , \48619 , \48620 , \48621 , \48622 ,
         \48623 , \48624 , \48625 , \48626 , \48627 , \48628 , \48629 , \48630 , \48631 , \48632 ,
         \48633 , \48634 , \48635 , \48636 , \48637 , \48638 , \48639 , \48640 , \48641 , \48642 ,
         \48643 , \48644 , \48645 , \48646 , \48647 , \48648 , \48649 , \48650 , \48651 , \48652 ,
         \48653 , \48654 , \48655 , \48656 , \48657 , \48658 , \48659 , \48660 , \48661 , \48662 ,
         \48663 , \48664 , \48665 , \48666 , \48667 , \48668 , \48669 , \48670 , \48671 , \48672 ,
         \48673 , \48674 , \48675 , \48676 , \48677 , \48678 , \48679 , \48680 , \48681 , \48682 ,
         \48683 , \48684 , \48685 , \48686 , \48687 , \48688 , \48689 , \48690 , \48691 , \48692 ,
         \48693 , \48694 , \48695 , \48696 , \48697 , \48698 , \48699 , \48700 , \48701 , \48702 ,
         \48703 , \48704 , \48705 , \48706 , \48707 , \48708 , \48709 , \48710 , \48711 , \48712 ,
         \48713 , \48714 , \48715 , \48716 , \48717 , \48718 , \48719 , \48720 , \48721 , \48722 ,
         \48723 , \48724 , \48725 , \48726 , \48727 , \48728 , \48729 , \48730 , \48731 , \48732 ,
         \48733 , \48734 , \48735 , \48736 , \48737 , \48738 , \48739 , \48740 , \48741 , \48742 ,
         \48743 , \48744 , \48745 , \48746 , \48747 , \48748 , \48749 , \48750 , \48751 , \48752 ,
         \48753 , \48754 , \48755 , \48756 , \48757 , \48758 , \48759 , \48760 , \48761 , \48762 ,
         \48763 , \48764 , \48765 , \48766 , \48767 , \48768 , \48769 , \48770 , \48771 , \48772 ,
         \48773 , \48774 , \48775 , \48776 , \48777 , \48778 , \48779 , \48780 , \48781 , \48782 ,
         \48783 , \48784 , \48785 , \48786 , \48787 , \48788 , \48789 , \48790 , \48791 , \48792 ,
         \48793 , \48794 , \48795 , \48796 , \48797 , \48798 , \48799 , \48800 , \48801 , \48802 ,
         \48803 , \48804 , \48805 , \48806 , \48807 , \48808 , \48809 , \48810 , \48811 , \48812 ,
         \48813 , \48814 , \48815 , \48816 , \48817 , \48818 , \48819 , \48820 , \48821 , \48822 ,
         \48823 , \48824 , \48825 , \48826 , \48827 , \48828 , \48829 , \48830 , \48831 , \48832 ,
         \48833 , \48834 , \48835 , \48836 , \48837 , \48838 , \48839 , \48840 , \48841 , \48842 ,
         \48843 , \48844 , \48845 , \48846 , \48847 , \48848 , \48849 , \48850 , \48851 , \48852 ,
         \48853 , \48854 , \48855 , \48856 , \48857 , \48858 , \48859 , \48860 , \48861 , \48862 ,
         \48863 , \48864 , \48865 , \48866 , \48867 , \48868 , \48869 , \48870 , \48871 , \48872 ,
         \48873 , \48874 , \48875 , \48876 , \48877 , \48878 , \48879 , \48880 , \48881 , \48882 ,
         \48883 , \48884 , \48885 , \48886 , \48887 , \48888 , \48889 , \48890 , \48891 , \48892 ,
         \48893 , \48894 , \48895 , \48896 , \48897 , \48898 , \48899 , \48900 , \48901 , \48902 ,
         \48903 , \48904 , \48905 , \48906 , \48907 , \48908 , \48909 , \48910 , \48911 , \48912 ,
         \48913 , \48914 , \48915 , \48916 , \48917 , \48918 , \48919 , \48920 , \48921 , \48922 ,
         \48923 , \48924 , \48925 , \48926 , \48927 , \48928 , \48929 , \48930 , \48931 , \48932 ,
         \48933 , \48934 , \48935 , \48936 , \48937 , \48938 , \48939 , \48940 , \48941 , \48942 ,
         \48943 , \48944 , \48945 , \48946 , \48947 , \48948 , \48949 , \48950 , \48951 , \48952 ,
         \48953 , \48954 , \48955 , \48956 , \48957 , \48958 , \48959 , \48960 , \48961 , \48962 ,
         \48963 , \48964 , \48965 , \48966 , \48967 , \48968 , \48969 , \48970 , \48971 , \48972 ,
         \48973 , \48974 , \48975 , \48976 , \48977 , \48978 , \48979 , \48980 , \48981 , \48982 ,
         \48983 , \48984 , \48985 , \48986 , \48987 , \48988 , \48989 , \48990 , \48991 , \48992 ,
         \48993 , \48994 , \48995 , \48996 , \48997 , \48998 , \48999 , \49000 , \49001 , \49002 ,
         \49003 , \49004 , \49005 , \49006 , \49007 , \49008 , \49009 , \49010 , \49011 , \49012 ,
         \49013 , \49014 , \49015 , \49016 , \49017 , \49018 , \49019 , \49020 , \49021 , \49022 ,
         \49023 , \49024 , \49025 , \49026 , \49027 , \49028 , \49029 , \49030 , \49031 , \49032 ,
         \49033 , \49034 , \49035 , \49036 , \49037 , \49038 , \49039 , \49040 , \49041 , \49042 ,
         \49043 , \49044 , \49045 , \49046 , \49047 , \49048 , \49049 , \49050 , \49051 , \49052 ,
         \49053 , \49054 , \49055 , \49056 , \49057 , \49058 , \49059 , \49060 , \49061 , \49062 ,
         \49063 , \49064 , \49065 , \49066 , \49067 , \49068 , \49069 , \49070 , \49071 , \49072 ,
         \49073 , \49074 , \49075 , \49076 , \49077 , \49078 , \49079 , \49080 , \49081 , \49082 ,
         \49083 , \49084 , \49085 , \49086 , \49087 , \49088 , \49089 , \49090 , \49091 , \49092 ,
         \49093 , \49094 , \49095 , \49096 , \49097 , \49098 , \49099 , \49100 , \49101 , \49102 ,
         \49103 , \49104 , \49105 , \49106 , \49107 , \49108 , \49109 , \49110 , \49111 , \49112 ,
         \49113 , \49114 , \49115 , \49116 , \49117 , \49118 , \49119 , \49120 , \49121 , \49122 ,
         \49123 , \49124 , \49125 , \49126 , \49127 , \49128 , \49129 , \49130 , \49131 , \49132 ,
         \49133 , \49134 , \49135 , \49136 , \49137 , \49138 , \49139 , \49140 , \49141 , \49142 ,
         \49143 , \49144 , \49145 , \49146 , \49147 , \49148 , \49149 , \49150 , \49151 , \49152 ,
         \49153 , \49154 , \49155 , \49156 , \49157 , \49158 , \49159 , \49160 , \49161 , \49162 ,
         \49163 , \49164 , \49165 , \49166 , \49167 , \49168 , \49169 , \49170 , \49171 , \49172 ,
         \49173 , \49174 , \49175 , \49176 , \49177 , \49178 , \49179 , \49180 , \49181 , \49182 ,
         \49183 , \49184 , \49185 , \49186 , \49187 , \49188 , \49189 , \49190 , \49191 , \49192 ,
         \49193 , \49194 , \49195 , \49196 , \49197 , \49198 , \49199 , \49200 , \49201 , \49202 ,
         \49203 , \49204 , \49205 , \49206 , \49207 , \49208 , \49209 , \49210 , \49211 , \49212 ,
         \49213 , \49214 , \49215 , \49216 , \49217 , \49218 , \49219 , \49220 , \49221 , \49222 ,
         \49223 , \49224 , \49225 , \49226 , \49227 , \49228 , \49229 , \49230 , \49231 , \49232 ,
         \49233 , \49234 , \49235 , \49236 , \49237 , \49238 , \49239 , \49240 , \49241 , \49242 ,
         \49243 , \49244 , \49245 , \49246 , \49247 , \49248 , \49249 , \49250 , \49251 , \49252 ,
         \49253 , \49254 , \49255 , \49256 , \49257 , \49258 , \49259 , \49260 , \49261 , \49262 ,
         \49263 , \49264 , \49265 , \49266 , \49267 , \49268 , \49269 , \49270 , \49271 , \49272 ,
         \49273 , \49274 , \49275 , \49276 , \49277 , \49278 , \49279 , \49280 , \49281 , \49282 ,
         \49283 , \49284 , \49285 , \49286 , \49287 , \49288 , \49289 , \49290 , \49291 , \49292 ,
         \49293 , \49294 , \49295 , \49296 , \49297 , \49298 , \49299 , \49300 , \49301 , \49302 ,
         \49303 , \49304 , \49305 , \49306 , \49307 , \49308 , \49309 , \49310 , \49311 , \49312 ,
         \49313 , \49314 , \49315 , \49316 , \49317 , \49318 , \49319 , \49320 , \49321 , \49322 ,
         \49323 , \49324 , \49325 , \49326 , \49327 , \49328 , \49329 , \49330 , \49331 , \49332 ,
         \49333 , \49334 , \49335 , \49336 , \49337 , \49338 , \49339 , \49340 , \49341 , \49342 ,
         \49343 , \49344 , \49345 , \49346 , \49347 , \49348 , \49349 , \49350 , \49351 , \49352 ,
         \49353 , \49354 , \49355 , \49356 , \49357 , \49358 , \49359 , \49360 , \49361 , \49362 ,
         \49363 , \49364 , \49365 , \49366 , \49367 , \49368 , \49369 , \49370 , \49371 , \49372 ,
         \49373 , \49374 , \49375 , \49376 , \49377 , \49378 , \49379 , \49380 , \49381 , \49382 ,
         \49383 , \49384 , \49385 , \49386 , \49387 , \49388 , \49389 , \49390 , \49391 , \49392 ,
         \49393 , \49394 , \49395 , \49396 , \49397 , \49398 , \49399 , \49400 , \49401 , \49402 ,
         \49403 , \49404 , \49405 , \49406 , \49407 , \49408 , \49409 , \49410 , \49411 , \49412 ,
         \49413 , \49414 , \49415 , \49416 , \49417 , \49418 , \49419 , \49420 , \49421 , \49422 ,
         \49423 , \49424 , \49425 , \49426 , \49427 , \49428 , \49429 , \49430 , \49431 , \49432 ,
         \49433 , \49434 , \49435 , \49436 , \49437 , \49438 , \49439 , \49440 , \49441 , \49442 ,
         \49443 , \49444 , \49445 , \49446 , \49447 , \49448 , \49449 , \49450 , \49451 , \49452 ,
         \49453 , \49454 , \49455 , \49456 , \49457 , \49458 , \49459 , \49460 , \49461 , \49462 ,
         \49463 , \49464 , \49465 , \49466 , \49467 , \49468 , \49469 , \49470 , \49471 , \49472 ,
         \49473 , \49474 , \49475 , \49476 , \49477 , \49478 , \49479 , \49480 , \49481 , \49482 ,
         \49483 , \49484 , \49485 , \49486 , \49487 , \49488 , \49489 , \49490 , \49491 , \49492 ,
         \49493 , \49494 , \49495 , \49496 , \49497 , \49498 , \49499 , \49500 , \49501 , \49502 ,
         \49503 , \49504 , \49505 , \49506 , \49507 , \49508 , \49509 , \49510 , \49511 , \49512 ,
         \49513 , \49514 , \49515 , \49516 , \49517 , \49518 , \49519 , \49520 , \49521 , \49522 ,
         \49523 , \49524 , \49525 , \49526 , \49527 , \49528 , \49529 , \49530 , \49531 , \49532 ,
         \49533 , \49534 , \49535 , \49536 , \49537 , \49538 , \49539 , \49540 , \49541 , \49542 ,
         \49543 , \49544 , \49545 , \49546 , \49547 , \49548 , \49549 , \49550 , \49551 , \49552 ,
         \49553 , \49554 , \49555 , \49556 , \49557 , \49558 , \49559 , \49560 , \49561 , \49562 ,
         \49563 , \49564 , \49565 , \49566 , \49567 , \49568 , \49569 , \49570 , \49571 , \49572 ,
         \49573 , \49574 , \49575 , \49576 , \49577 , \49578 , \49579 , \49580 , \49581 , \49582 ,
         \49583 , \49584 , \49585 , \49586 , \49587 , \49588 , \49589 , \49590 , \49591 , \49592 ,
         \49593 , \49594 , \49595 , \49596 , \49597 , \49598 , \49599 , \49600 , \49601 , \49602 ,
         \49603 , \49604 , \49605 , \49606 , \49607 , \49608 , \49609 , \49610 , \49611 , \49612 ,
         \49613 , \49614 , \49615 , \49616 , \49617 , \49618 , \49619 , \49620 , \49621 , \49622 ,
         \49623 , \49624 , \49625 , \49626 , \49627 , \49628 , \49629 , \49630 , \49631 , \49632 ,
         \49633 , \49634 , \49635 , \49636 , \49637 , \49638 , \49639 , \49640 , \49641 , \49642 ,
         \49643 , \49644 , \49645 , \49646 , \49647 , \49648 , \49649 , \49650 , \49651 , \49652 ,
         \49653 , \49654 , \49655 , \49656 , \49657 , \49658 , \49659 , \49660 , \49661 , \49662 ,
         \49663 , \49664 , \49665 , \49666 , \49667 , \49668 , \49669 , \49670 , \49671 , \49672 ,
         \49673 , \49674 , \49675 , \49676 , \49677 , \49678 , \49679 , \49680 , \49681 , \49682 ,
         \49683 , \49684 , \49685 , \49686 , \49687 , \49688 , \49689 , \49690 , \49691 , \49692 ,
         \49693 , \49694 , \49695 , \49696 , \49697 , \49698 , \49699 , \49700 , \49701 , \49702 ,
         \49703 , \49704 , \49705 , \49706 , \49707 , \49708 , \49709 , \49710 , \49711 , \49712 ,
         \49713 , \49714 , \49715 , \49716 , \49717 , \49718 , \49719 , \49720 , \49721 , \49722 ,
         \49723 , \49724 , \49725 , \49726 , \49727 , \49728 , \49729 , \49730 , \49731 , \49732 ,
         \49733 , \49734 , \49735 , \49736 , \49737 , \49738 , \49739 , \49740 , \49741 , \49742 ,
         \49743 , \49744 , \49745 , \49746 , \49747 , \49748 , \49749 , \49750 , \49751 , \49752 ,
         \49753 , \49754 , \49755 , \49756 , \49757 , \49758 , \49759 , \49760 , \49761 , \49762 ,
         \49763 , \49764 , \49765 , \49766 , \49767 , \49768 , \49769 , \49770 , \49771 , \49772 ,
         \49773 , \49774 , \49775 , \49776 , \49777 , \49778 , \49779 , \49780 , \49781 , \49782 ,
         \49783 , \49784 , \49785 , \49786 , \49787 , \49788 , \49789 , \49790 , \49791 , \49792 ,
         \49793 , \49794 , \49795 , \49796 , \49797 , \49798 , \49799 , \49800 , \49801 , \49802 ,
         \49803 , \49804 , \49805 , \49806 , \49807 , \49808 , \49809 , \49810 , \49811 , \49812 ,
         \49813 , \49814 , \49815 , \49816 , \49817 , \49818 , \49819 , \49820 , \49821 , \49822 ,
         \49823 , \49824 , \49825 , \49826 , \49827 , \49828 , \49829 , \49830 , \49831 , \49832 ,
         \49833 , \49834 , \49835 , \49836 , \49837 , \49838 , \49839 , \49840 , \49841 , \49842 ,
         \49843 , \49844 , \49845 , \49846 , \49847 , \49848 , \49849 , \49850 , \49851 , \49852 ,
         \49853 , \49854 , \49855 , \49856 , \49857 , \49858 , \49859 , \49860 , \49861 , \49862 ,
         \49863 , \49864 , \49865 , \49866 , \49867 , \49868 , \49869 , \49870 , \49871 , \49872 ,
         \49873 , \49874 , \49875 , \49876 , \49877 , \49878 , \49879 , \49880 , \49881 , \49882 ,
         \49883 , \49884 , \49885 , \49886 , \49887 , \49888 , \49889 , \49890 , \49891 , \49892 ,
         \49893 , \49894 , \49895 , \49896 , \49897 , \49898 , \49899 , \49900 , \49901 , \49902 ,
         \49903 , \49904 , \49905 , \49906 , \49907 , \49908 , \49909 , \49910 , \49911 , \49912 ,
         \49913 , \49914 , \49915 , \49916 , \49917 , \49918 , \49919 , \49920 , \49921 , \49922 ,
         \49923 , \49924 , \49925 , \49926 , \49927 , \49928 , \49929 , \49930 , \49931 , \49932 ,
         \49933 , \49934 , \49935 , \49936 , \49937 , \49938 , \49939 , \49940 , \49941 , \49942 ,
         \49943 , \49944 , \49945 , \49946 , \49947 , \49948 , \49949 , \49950 , \49951 , \49952 ,
         \49953 , \49954 , \49955 , \49956 , \49957 , \49958 , \49959 , \49960 , \49961 , \49962 ,
         \49963 , \49964 , \49965 , \49966 , \49967 , \49968 , \49969 , \49970 , \49971 , \49972 ,
         \49973 , \49974 , \49975 , \49976 , \49977 , \49978 , \49979 , \49980 , \49981 , \49982 ,
         \49983 , \49984 , \49985 , \49986 , \49987 , \49988 , \49989 , \49990 , \49991 , \49992 ,
         \49993 , \49994 , \49995 , \49996 , \49997 , \49998 , \49999 , \50000 , \50001 , \50002 ,
         \50003 , \50004 , \50005 , \50006 , \50007 , \50008 , \50009 , \50010 , \50011 , \50012 ,
         \50013 , \50014 , \50015 , \50016 , \50017 , \50018 , \50019 , \50020 , \50021 , \50022 ,
         \50023 , \50024 , \50025 , \50026 , \50027 , \50028 , \50029 , \50030 , \50031 , \50032 ,
         \50033 , \50034 , \50035 , \50036 , \50037 , \50038 , \50039 , \50040 , \50041 , \50042 ,
         \50043 , \50044 , \50045 , \50046 , \50047 , \50048 , \50049 , \50050 , \50051 , \50052 ,
         \50053 , \50054 , \50055 , \50056 , \50057 , \50058 , \50059 , \50060 , \50061 , \50062 ,
         \50063 , \50064 , \50065 , \50066 , \50067 , \50068 , \50069 , \50070 , \50071 , \50072 ,
         \50073 , \50074 , \50075 , \50076 , \50077 , \50078 , \50079 , \50080 , \50081 , \50082 ,
         \50083 , \50084 , \50085 , \50086 , \50087 , \50088 , \50089 , \50090 , \50091 , \50092 ,
         \50093 , \50094 , \50095 , \50096 , \50097 , \50098 , \50099 , \50100 , \50101 , \50102 ,
         \50103 , \50104 , \50105 , \50106 , \50107 , \50108 , \50109 , \50110 , \50111 , \50112 ,
         \50113 , \50114 , \50115 , \50116 , \50117 , \50118 , \50119 , \50120 , \50121 , \50122 ,
         \50123 , \50124 , \50125 , \50126 , \50127 , \50128 , \50129 , \50130 , \50131 , \50132 ,
         \50133 , \50134 , \50135 , \50136 , \50137 , \50138 , \50139 , \50140 , \50141 , \50142 ,
         \50143 , \50144 , \50145 , \50146 , \50147 , \50148 , \50149 , \50150 , \50151 , \50152 ,
         \50153 , \50154 , \50155 , \50156 , \50157 , \50158 , \50159 , \50160 , \50161 , \50162 ,
         \50163 , \50164 , \50165 , \50166 , \50167 , \50168 , \50169 , \50170 , \50171 , \50172 ,
         \50173 , \50174 , \50175 , \50176 , \50177 , \50178 , \50179 , \50180 , \50181 , \50182 ,
         \50183 , \50184 , \50185 , \50186 , \50187 , \50188 , \50189 , \50190 , \50191 , \50192 ,
         \50193 , \50194 , \50195 , \50196 , \50197 , \50198 , \50199 , \50200 , \50201 , \50202 ,
         \50203 , \50204 , \50205 , \50206 , \50207 , \50208 , \50209 , \50210 , \50211 , \50212 ,
         \50213 , \50214 , \50215 , \50216 , \50217 , \50218 , \50219 , \50220 , \50221 , \50222 ,
         \50223 , \50224 , \50225 , \50226 , \50227 , \50228 , \50229 , \50230 , \50231 , \50232 ,
         \50233 , \50234 , \50235 , \50236 , \50237 , \50238 , \50239 , \50240 , \50241 , \50242 ,
         \50243 , \50244 , \50245 , \50246 , \50247 , \50248 , \50249 , \50250 , \50251 , \50252 ,
         \50253 , \50254 , \50255 , \50256 , \50257 , \50258 , \50259 , \50260 , \50261 , \50262 ,
         \50263 , \50264 , \50265 , \50266 , \50267 , \50268 , \50269 , \50270 , \50271 , \50272 ,
         \50273 , \50274 , \50275 , \50276 , \50277 , \50278 , \50279 , \50280 , \50281 , \50282 ,
         \50283 , \50284 , \50285 , \50286 , \50287 , \50288 , \50289 , \50290 , \50291 , \50292 ,
         \50293 , \50294 , \50295 , \50296 , \50297 , \50298 , \50299 , \50300 , \50301 , \50302 ,
         \50303 , \50304 , \50305 , \50306 , \50307 , \50308 , \50309 , \50310 , \50311 , \50312 ,
         \50313 , \50314 , \50315 , \50316 , \50317 , \50318 , \50319 , \50320 , \50321 , \50322 ,
         \50323 , \50324 , \50325 , \50326 , \50327 , \50328 , \50329 , \50330 , \50331 , \50332 ,
         \50333 , \50334 , \50335 , \50336 , \50337 , \50338 , \50339 , \50340 , \50341 , \50342 ,
         \50343 , \50344 , \50345 , \50346 , \50347 , \50348 , \50349 , \50350 , \50351 , \50352 ,
         \50353 , \50354 , \50355 , \50356 , \50357 , \50358 , \50359 , \50360 , \50361 , \50362 ,
         \50363 , \50364 , \50365 , \50366 , \50367 , \50368 , \50369 , \50370 , \50371 , \50372 ,
         \50373 , \50374 , \50375 , \50376 , \50377 , \50378 , \50379 , \50380 , \50381 , \50382 ,
         \50383 , \50384 , \50385 , \50386 , \50387 , \50388 , \50389 , \50390 , \50391 , \50392 ,
         \50393 , \50394 , \50395 , \50396 , \50397 , \50398 , \50399 , \50400 , \50401 , \50402 ,
         \50403 , \50404 , \50405 , \50406 , \50407 , \50408 , \50409 , \50410 , \50411 , \50412 ,
         \50413 , \50414 , \50415 , \50416 , \50417 , \50418 , \50419 , \50420 , \50421 , \50422 ,
         \50423 , \50424 , \50425 , \50426 , \50427 , \50428 , \50429 , \50430 , \50431 , \50432 ,
         \50433 , \50434 , \50435 , \50436 , \50437 , \50438 , \50439 , \50440 , \50441 , \50442 ,
         \50443 , \50444 , \50445 , \50446 , \50447 , \50448 , \50449 , \50450 , \50451 , \50452 ,
         \50453 , \50454 , \50455 , \50456 , \50457 , \50458 , \50459 , \50460 , \50461 , \50462 ,
         \50463 , \50464 , \50465 , \50466 , \50467 , \50468 , \50469 , \50470 , \50471 , \50472 ,
         \50473 , \50474 , \50475 , \50476 , \50477 , \50478 , \50479 , \50480 , \50481 , \50482 ,
         \50483 , \50484 , \50485 , \50486 , \50487 , \50488 , \50489 , \50490 , \50491 , \50492 ,
         \50493 , \50494 , \50495 , \50496 , \50497 , \50498 , \50499 , \50500 , \50501 , \50502 ,
         \50503 , \50504 , \50505 , \50506 , \50507 , \50508 , \50509 , \50510 , \50511 , \50512 ,
         \50513 , \50514 , \50515 , \50516 , \50517 , \50518 , \50519 , \50520 , \50521 , \50522 ,
         \50523 , \50524 , \50525 , \50526 , \50527 , \50528 , \50529 , \50530 , \50531 , \50532 ,
         \50533 , \50534 , \50535 , \50536 , \50537 , \50538 , \50539 , \50540 , \50541 , \50542 ,
         \50543 , \50544 , \50545 , \50546 , \50547 , \50548 , \50549 , \50550 , \50551 , \50552 ,
         \50553 , \50554 , \50555 , \50556 , \50557 , \50558 , \50559 , \50560 , \50561 , \50562 ,
         \50563 , \50564 , \50565 , \50566 , \50567 , \50568 , \50569 , \50570 , \50571 , \50572 ,
         \50573 , \50574 , \50575 , \50576 , \50577 , \50578 , \50579 , \50580 , \50581 , \50582 ,
         \50583 , \50584 , \50585 , \50586 , \50587 , \50588 , \50589 , \50590 , \50591 , \50592 ,
         \50593 , \50594 , \50595 , \50596 , \50597 , \50598 , \50599 , \50600 , \50601 , \50602 ,
         \50603 , \50604 , \50605 , \50606 , \50607 , \50608 , \50609 , \50610 , \50611 , \50612 ,
         \50613 , \50614 , \50615 , \50616 , \50617 , \50618 , \50619 , \50620 , \50621 , \50622 ,
         \50623 , \50624 , \50625 , \50626 , \50627 , \50628 , \50629 , \50630 , \50631 , \50632 ,
         \50633 , \50634 , \50635 , \50636 , \50637 , \50638 , \50639 , \50640 , \50641 , \50642 ,
         \50643 , \50644 , \50645 , \50646 , \50647 , \50648 , \50649 , \50650 , \50651 , \50652 ,
         \50653 , \50654 , \50655 , \50656 , \50657 , \50658 , \50659 , \50660 , \50661 , \50662 ,
         \50663 , \50664 , \50665 , \50666 , \50667 , \50668 , \50669 , \50670 , \50671 , \50672 ,
         \50673 , \50674 , \50675 , \50676 , \50677 , \50678 , \50679 , \50680 , \50681 , \50682 ,
         \50683 , \50684 , \50685 , \50686 , \50687 , \50688 , \50689 , \50690 , \50691 , \50692 ,
         \50693 , \50694 , \50695 , \50696 , \50697 , \50698 , \50699 , \50700 , \50701 , \50702 ,
         \50703 , \50704 , \50705 , \50706 , \50707 , \50708 , \50709 , \50710 , \50711 , \50712 ,
         \50713 , \50714 , \50715 , \50716 , \50717 , \50718 , \50719 , \50720 , \50721 , \50722 ,
         \50723 , \50724 , \50725 , \50726 , \50727 , \50728 , \50729 , \50730 , \50731 , \50732 ,
         \50733 , \50734 , \50735 , \50736 , \50737 , \50738 , \50739 , \50740 , \50741 , \50742 ,
         \50743 , \50744 , \50745 , \50746 , \50747 , \50748 , \50749 , \50750 , \50751 , \50752 ,
         \50753 , \50754 , \50755 , \50756 , \50757 , \50758 , \50759 , \50760 , \50761 , \50762 ,
         \50763 , \50764 , \50765 , \50766 , \50767 , \50768 , \50769 , \50770 , \50771 , \50772 ,
         \50773 , \50774 , \50775 , \50776 , \50777 , \50778 , \50779 , \50780 , \50781 , \50782 ,
         \50783 , \50784 , \50785 , \50786 , \50787 , \50788 , \50789 , \50790 , \50791 , \50792 ,
         \50793 , \50794 , \50795 , \50796 , \50797 , \50798 , \50799 , \50800 , \50801 , \50802 ,
         \50803 , \50804 , \50805 , \50806 , \50807 , \50808 , \50809 , \50810 , \50811 , \50812 ,
         \50813 , \50814 , \50815 , \50816 , \50817 , \50818 , \50819 , \50820 , \50821 , \50822 ,
         \50823 , \50824 , \50825 , \50826 , \50827 , \50828 , \50829 , \50830 , \50831 , \50832 ,
         \50833 , \50834 , \50835 , \50836 , \50837 , \50838 , \50839 , \50840 , \50841 , \50842 ,
         \50843 , \50844 , \50845 , \50846 , \50847 , \50848 , \50849 , \50850 , \50851 , \50852 ,
         \50853 , \50854 , \50855 , \50856 , \50857 , \50858 , \50859 , \50860 , \50861 , \50862 ,
         \50863 , \50864 , \50865 , \50866 , \50867 , \50868 , \50869 , \50870 , \50871 , \50872 ,
         \50873 , \50874 , \50875 , \50876 , \50877 , \50878 , \50879 , \50880 , \50881 , \50882 ,
         \50883 , \50884 , \50885 , \50886 , \50887 , \50888 , \50889 , \50890 , \50891 , \50892 ,
         \50893 , \50894 , \50895 , \50896 , \50897 , \50898 , \50899 , \50900 , \50901 , \50902 ,
         \50903 , \50904 , \50905 , \50906 , \50907 , \50908 , \50909 , \50910 , \50911 , \50912 ,
         \50913 , \50914 , \50915 , \50916 , \50917 , \50918 , \50919 , \50920 , \50921 , \50922 ,
         \50923 , \50924 , \50925 , \50926 , \50927 , \50928 , \50929 , \50930 , \50931 , \50932 ,
         \50933 , \50934 , \50935 , \50936 , \50937 , \50938 , \50939 , \50940 , \50941 , \50942 ,
         \50943 , \50944 , \50945 , \50946 , \50947 , \50948 , \50949 , \50950 , \50951 , \50952 ,
         \50953 , \50954 , \50955 , \50956 , \50957 , \50958 , \50959 , \50960 , \50961 , \50962 ,
         \50963 , \50964 , \50965 , \50966 , \50967 , \50968 , \50969 , \50970 , \50971 , \50972 ,
         \50973 , \50974 , \50975 , \50976 , \50977 , \50978 , \50979 , \50980 , \50981 , \50982 ,
         \50983 , \50984 , \50985 , \50986 , \50987 , \50988 , \50989 , \50990 , \50991 , \50992 ,
         \50993 , \50994 , \50995 , \50996 , \50997 , \50998 , \50999 , \51000 , \51001 , \51002 ,
         \51003 , \51004 , \51005 , \51006 , \51007 , \51008 , \51009 , \51010 , \51011 , \51012 ,
         \51013 , \51014 , \51015 , \51016 , \51017 , \51018 , \51019 , \51020 , \51021 , \51022 ,
         \51023 , \51024 , \51025 , \51026 , \51027 , \51028 , \51029 , \51030 , \51031 , \51032 ,
         \51033 , \51034 , \51035 , \51036 , \51037 , \51038 , \51039 , \51040 , \51041 , \51042 ,
         \51043 , \51044 , \51045 , \51046 , \51047 , \51048 , \51049 , \51050 , \51051 , \51052 ,
         \51053 , \51054 , \51055 , \51056 , \51057 , \51058 , \51059 , \51060 , \51061 , \51062 ,
         \51063 , \51064 , \51065 , \51066 , \51067 , \51068 , \51069 , \51070 , \51071 , \51072 ,
         \51073 , \51074 , \51075 , \51076 , \51077 , \51078 , \51079 , \51080 , \51081 , \51082 ,
         \51083 , \51084 , \51085 , \51086 , \51087 , \51088 , \51089 , \51090 , \51091 , \51092 ,
         \51093 , \51094 , \51095 , \51096 , \51097 , \51098 , \51099 , \51100 , \51101 , \51102 ,
         \51103 , \51104 , \51105 , \51106 , \51107 , \51108 , \51109 , \51110 , \51111 , \51112 ,
         \51113 , \51114 , \51115 , \51116 , \51117 , \51118 , \51119 , \51120 , \51121 , \51122 ,
         \51123 , \51124 , \51125 , \51126 , \51127 , \51128 , \51129 , \51130 , \51131 , \51132 ,
         \51133 , \51134 , \51135 , \51136 , \51137 , \51138 , \51139 , \51140 , \51141 , \51142 ,
         \51143 , \51144 , \51145 , \51146 , \51147 , \51148 , \51149 , \51150 , \51151 , \51152 ,
         \51153 , \51154 , \51155 , \51156 , \51157 , \51158 , \51159 , \51160 , \51161 , \51162 ,
         \51163 , \51164 , \51165 , \51166 , \51167 , \51168 , \51169 , \51170 , \51171 , \51172 ,
         \51173 , \51174 , \51175 , \51176 , \51177 , \51178 , \51179 , \51180 , \51181 , \51182 ,
         \51183 , \51184 , \51185 , \51186 , \51187 , \51188 , \51189 , \51190 , \51191 , \51192 ,
         \51193 , \51194 , \51195 , \51196 , \51197 , \51198 , \51199 , \51200 , \51201 , \51202 ,
         \51203 , \51204 , \51205 , \51206 , \51207 , \51208 , \51209 , \51210 , \51211 , \51212 ,
         \51213 , \51214 , \51215 , \51216 , \51217 , \51218 , \51219 , \51220 , \51221 , \51222 ,
         \51223 , \51224 , \51225 , \51226 , \51227 , \51228 , \51229 , \51230 , \51231 , \51232 ,
         \51233 , \51234 , \51235 , \51236 , \51237 , \51238 , \51239 , \51240 , \51241 , \51242 ,
         \51243 , \51244 , \51245 , \51246 , \51247 , \51248 , \51249 , \51250 , \51251 , \51252 ,
         \51253 , \51254 , \51255 , \51256 , \51257 , \51258 , \51259 , \51260 , \51261 , \51262 ,
         \51263 , \51264 , \51265 , \51266 , \51267 , \51268 , \51269 , \51270 , \51271 , \51272 ,
         \51273 , \51274 , \51275 , \51276 , \51277 , \51278 , \51279 , \51280 , \51281 , \51282 ,
         \51283 , \51284 , \51285 , \51286 , \51287 , \51288 , \51289 , \51290 , \51291 , \51292 ,
         \51293 , \51294 , \51295 , \51296 , \51297 , \51298 , \51299 , \51300 , \51301 , \51302 ,
         \51303 , \51304 , \51305 , \51306 , \51307 , \51308 , \51309 , \51310 , \51311 , \51312 ,
         \51313 , \51314 , \51315 , \51316 , \51317 , \51318 , \51319 , \51320 , \51321 , \51322 ,
         \51323 , \51324 , \51325 , \51326 , \51327 , \51328 , \51329 , \51330 , \51331 , \51332 ,
         \51333 , \51334 , \51335 , \51336 , \51337 , \51338 , \51339 , \51340 , \51341 , \51342 ,
         \51343 , \51344 , \51345 , \51346 , \51347 , \51348 , \51349 , \51350 , \51351 , \51352 ,
         \51353 , \51354 , \51355 , \51356 , \51357 , \51358 , \51359 , \51360 , \51361 , \51362 ,
         \51363 , \51364 , \51365 , \51366 , \51367 , \51368 , \51369 , \51370 , \51371 , \51372 ,
         \51373 , \51374 , \51375 , \51376 , \51377 , \51378 , \51379 , \51380 , \51381 , \51382 ,
         \51383 , \51384 , \51385 , \51386 , \51387 , \51388 , \51389 , \51390 , \51391 , \51392 ,
         \51393 , \51394 , \51395 , \51396 , \51397 , \51398 , \51399 , \51400 , \51401 , \51402 ,
         \51403 , \51404 , \51405 , \51406 , \51407 , \51408 , \51409 , \51410 , \51411 , \51412 ,
         \51413 , \51414 , \51415 , \51416 , \51417 , \51418 , \51419 , \51420 , \51421 , \51422 ,
         \51423 , \51424 , \51425 , \51426 , \51427 , \51428 , \51429 , \51430 , \51431 , \51432 ,
         \51433 , \51434 , \51435 , \51436 , \51437 , \51438 , \51439 , \51440 , \51441 , \51442 ,
         \51443 , \51444 , \51445 , \51446 , \51447 , \51448 , \51449 , \51450 , \51451 , \51452 ,
         \51453 , \51454 , \51455 , \51456 , \51457 , \51458 , \51459 , \51460 , \51461 , \51462 ,
         \51463 , \51464 , \51465 , \51466 , \51467 , \51468 , \51469 , \51470 , \51471 , \51472 ,
         \51473 , \51474 , \51475 , \51476 , \51477 , \51478 , \51479 , \51480 , \51481 , \51482 ,
         \51483 , \51484 , \51485 , \51486 , \51487 , \51488 , \51489 , \51490 , \51491 , \51492 ,
         \51493 , \51494 , \51495 , \51496 , \51497 , \51498 , \51499 , \51500 , \51501 , \51502 ,
         \51503 , \51504 , \51505 , \51506 , \51507 , \51508 , \51509 , \51510 , \51511 , \51512 ,
         \51513 , \51514 , \51515 , \51516 , \51517 , \51518 , \51519 , \51520 , \51521 , \51522 ,
         \51523 , \51524 , \51525 , \51526 , \51527 , \51528 , \51529 , \51530 , \51531 , \51532 ,
         \51533 , \51534 , \51535 , \51536 , \51537 , \51538 , \51539 , \51540 , \51541 , \51542 ,
         \51543 , \51544 , \51545 , \51546 , \51547 , \51548 , \51549 , \51550 , \51551 , \51552 ,
         \51553 , \51554 , \51555 , \51556 , \51557 , \51558 , \51559 , \51560 , \51561 , \51562 ,
         \51563 , \51564 , \51565 , \51566 , \51567 , \51568 , \51569 , \51570 , \51571 , \51572 ,
         \51573 , \51574 , \51575 , \51576 , \51577 , \51578 , \51579 , \51580 , \51581 , \51582 ,
         \51583 , \51584 , \51585 , \51586 , \51587 , \51588 , \51589 , \51590 , \51591 , \51592 ,
         \51593 , \51594 , \51595 , \51596 , \51597 , \51598 , \51599 , \51600 , \51601 , \51602 ,
         \51603 , \51604 , \51605 , \51606 , \51607 , \51608 , \51609 , \51610 , \51611 , \51612 ,
         \51613 , \51614 , \51615 , \51616 , \51617 , \51618 , \51619 , \51620 , \51621 , \51622 ,
         \51623 , \51624 , \51625 , \51626 , \51627 , \51628 , \51629 , \51630 , \51631 , \51632 ,
         \51633 , \51634 , \51635 , \51636 , \51637 , \51638 , \51639 , \51640 , \51641 , \51642 ,
         \51643 , \51644 , \51645 , \51646 , \51647 , \51648 , \51649 , \51650 , \51651 , \51652 ,
         \51653 , \51654 , \51655 , \51656 , \51657 , \51658 , \51659 , \51660 , \51661 , \51662 ,
         \51663 , \51664 , \51665 , \51666 , \51667 , \51668 , \51669 , \51670 , \51671 , \51672 ,
         \51673 , \51674 , \51675 , \51676 , \51677 , \51678 , \51679 , \51680 , \51681 , \51682 ,
         \51683 , \51684 , \51685 , \51686 , \51687 , \51688 , \51689 , \51690 , \51691 , \51692 ,
         \51693 , \51694 , \51695 , \51696 , \51697 , \51698 , \51699 , \51700 , \51701 , \51702 ,
         \51703 , \51704 , \51705 , \51706 , \51707 , \51708 , \51709 , \51710 , \51711 , \51712 ,
         \51713 , \51714 , \51715 , \51716 , \51717 , \51718 , \51719 , \51720 , \51721 , \51722 ,
         \51723 , \51724 , \51725 , \51726 , \51727 , \51728 , \51729 , \51730 , \51731 , \51732 ,
         \51733 , \51734 , \51735 , \51736 , \51737 , \51738 , \51739 , \51740 , \51741 , \51742 ,
         \51743 , \51744 , \51745 , \51746 , \51747 , \51748 , \51749 , \51750 , \51751 , \51752 ,
         \51753 , \51754 , \51755 , \51756 , \51757 , \51758 , \51759 , \51760 , \51761 , \51762 ,
         \51763 , \51764 , \51765 , \51766 , \51767 , \51768 , \51769 , \51770 , \51771 , \51772 ,
         \51773 , \51774 , \51775 , \51776 , \51777 , \51778 , \51779 , \51780 , \51781 , \51782 ,
         \51783 , \51784 , \51785 , \51786 , \51787 , \51788 , \51789 , \51790 , \51791 , \51792 ,
         \51793 , \51794 , \51795 , \51796 , \51797 , \51798 , \51799 , \51800 , \51801 , \51802 ,
         \51803 , \51804 , \51805 , \51806 , \51807 , \51808 , \51809 , \51810 , \51811 , \51812 ,
         \51813 , \51814 , \51815 , \51816 , \51817 , \51818 , \51819 , \51820 , \51821 , \51822 ,
         \51823 , \51824 , \51825 , \51826 , \51827 , \51828 , \51829 , \51830 , \51831 , \51832 ,
         \51833 , \51834 , \51835 , \51836 , \51837 , \51838 , \51839 , \51840 , \51841 , \51842 ,
         \51843 , \51844 , \51845 , \51846 , \51847 , \51848 , \51849 , \51850 , \51851 , \51852 ,
         \51853 , \51854 , \51855 , \51856 , \51857 , \51858 , \51859 , \51860 , \51861 , \51862 ,
         \51863 , \51864 , \51865 , \51866 , \51867 , \51868 , \51869 , \51870 , \51871 , \51872 ,
         \51873 , \51874 , \51875 , \51876 , \51877 , \51878 , \51879 , \51880 , \51881 , \51882 ,
         \51883 , \51884 , \51885 , \51886 , \51887 , \51888 , \51889 , \51890 , \51891 , \51892 ,
         \51893 , \51894 , \51895 , \51896 , \51897 , \51898 , \51899 , \51900 , \51901 , \51902 ,
         \51903 , \51904 , \51905 , \51906 , \51907 , \51908 , \51909 , \51910 , \51911 , \51912 ,
         \51913 , \51914 , \51915 , \51916 , \51917 , \51918 , \51919 , \51920 , \51921 , \51922 ,
         \51923 , \51924 , \51925 , \51926 , \51927 , \51928 , \51929 , \51930 , \51931 , \51932 ,
         \51933 , \51934 , \51935 , \51936 , \51937 , \51938 , \51939 , \51940 , \51941 , \51942 ,
         \51943 , \51944 , \51945 , \51946 , \51947 , \51948 , \51949 , \51950 , \51951 , \51952 ,
         \51953 , \51954 , \51955 , \51956 , \51957 , \51958 , \51959 , \51960 , \51961 , \51962 ,
         \51963 , \51964 , \51965 , \51966 , \51967 , \51968 , \51969 , \51970 , \51971 , \51972 ,
         \51973 , \51974 , \51975 , \51976 , \51977 , \51978 , \51979 , \51980 , \51981 , \51982 ,
         \51983 , \51984 , \51985 , \51986 , \51987 , \51988 , \51989 , \51990 , \51991 , \51992 ,
         \51993 , \51994 , \51995 , \51996 , \51997 , \51998 , \51999 , \52000 , \52001 , \52002 ,
         \52003 , \52004 , \52005 , \52006 , \52007 , \52008 , \52009 , \52010 , \52011 , \52012 ,
         \52013 , \52014 , \52015 , \52016 , \52017 , \52018 , \52019 , \52020 , \52021 , \52022 ,
         \52023 , \52024 , \52025 , \52026 , \52027 , \52028 , \52029 , \52030 , \52031 , \52032 ,
         \52033 , \52034 , \52035 , \52036 , \52037 , \52038 , \52039 , \52040 , \52041 , \52042 ,
         \52043 , \52044 , \52045 , \52046 , \52047 , \52048 , \52049 , \52050 , \52051 , \52052 ,
         \52053 , \52054 , \52055 , \52056 , \52057 , \52058 , \52059 , \52060 , \52061 , \52062 ,
         \52063 , \52064 , \52065 , \52066 , \52067 , \52068 , \52069 , \52070 , \52071 , \52072 ,
         \52073 , \52074 , \52075 , \52076 , \52077 , \52078 , \52079 , \52080 , \52081 , \52082 ,
         \52083 , \52084 , \52085 , \52086 , \52087 , \52088 , \52089 , \52090 , \52091 , \52092 ,
         \52093 , \52094 , \52095 , \52096 , \52097 , \52098 , \52099 , \52100 , \52101 , \52102 ,
         \52103 , \52104 , \52105 , \52106 , \52107 , \52108 , \52109 , \52110 , \52111 , \52112 ,
         \52113 , \52114 , \52115 , \52116 , \52117 , \52118 , \52119 , \52120 , \52121 , \52122 ,
         \52123 , \52124 , \52125 , \52126 , \52127 , \52128 , \52129 , \52130 , \52131 , \52132 ,
         \52133 , \52134 , \52135 , \52136 , \52137 , \52138 , \52139 , \52140 , \52141 , \52142 ,
         \52143 , \52144 , \52145 , \52146 , \52147 , \52148 , \52149 , \52150 , \52151 , \52152 ,
         \52153 , \52154 , \52155 , \52156 , \52157 , \52158 , \52159 , \52160 , \52161 , \52162 ,
         \52163 , \52164 , \52165 , \52166 , \52167 , \52168 , \52169 , \52170 , \52171 , \52172 ,
         \52173 , \52174 , \52175 , \52176 , \52177 , \52178 , \52179 , \52180 , \52181 , \52182 ,
         \52183 , \52184 , \52185 , \52186 , \52187 , \52188 , \52189 , \52190 , \52191 , \52192 ,
         \52193 , \52194 , \52195 , \52196 , \52197 , \52198 , \52199 , \52200 , \52201 , \52202 ,
         \52203 , \52204 , \52205 , \52206 , \52207 , \52208 , \52209 , \52210 , \52211 , \52212 ,
         \52213 , \52214 , \52215 , \52216 , \52217 , \52218 , \52219 , \52220 , \52221 , \52222 ,
         \52223 , \52224 , \52225 , \52226 , \52227 , \52228 , \52229 , \52230 , \52231 , \52232 ,
         \52233 , \52234 , \52235 , \52236 , \52237 , \52238 , \52239 , \52240 , \52241 , \52242 ,
         \52243 , \52244 , \52245 , \52246 , \52247 , \52248 , \52249 , \52250 , \52251 , \52252 ,
         \52253 , \52254 , \52255 , \52256 , \52257 , \52258 , \52259 , \52260 , \52261 , \52262 ,
         \52263 , \52264 , \52265 , \52266 , \52267 , \52268 , \52269 , \52270 , \52271 , \52272 ,
         \52273 , \52274 , \52275 , \52276 , \52277 , \52278 , \52279 , \52280 , \52281 , \52282 ,
         \52283 , \52284 , \52285 , \52286 , \52287 , \52288 , \52289 , \52290 , \52291 , \52292 ,
         \52293 , \52294 , \52295 , \52296 , \52297 , \52298 , \52299 , \52300 , \52301 , \52302 ,
         \52303 , \52304 , \52305 , \52306 , \52307 , \52308 , \52309 , \52310 , \52311 , \52312 ,
         \52313 , \52314 , \52315 , \52316 , \52317 , \52318 , \52319 , \52320 , \52321 , \52322 ,
         \52323 , \52324 , \52325 , \52326 , \52327 , \52328 , \52329 , \52330 , \52331 , \52332 ,
         \52333 , \52334 , \52335 , \52336 , \52337 , \52338 , \52339 , \52340 , \52341 , \52342 ,
         \52343 , \52344 , \52345 , \52346 , \52347 , \52348 , \52349 , \52350 , \52351 , \52352 ,
         \52353 , \52354 , \52355 , \52356 , \52357 , \52358 , \52359 , \52360 , \52361 , \52362 ,
         \52363 , \52364 , \52365 , \52366 , \52367 , \52368 , \52369 , \52370 , \52371 , \52372 ,
         \52373 , \52374 , \52375 , \52376 , \52377 , \52378 , \52379 , \52380 , \52381 , \52382 ,
         \52383 , \52384 , \52385 , \52386 , \52387 , \52388 , \52389 , \52390 , \52391 , \52392 ,
         \52393 , \52394 , \52395 , \52396 , \52397 , \52398 , \52399 , \52400 , \52401 , \52402 ,
         \52403 , \52404 , \52405 , \52406 , \52407 , \52408 , \52409 , \52410 , \52411 , \52412 ,
         \52413 , \52414 , \52415 , \52416 , \52417 , \52418 , \52419 , \52420 , \52421 , \52422 ,
         \52423 , \52424 , \52425 , \52426 , \52427 , \52428 , \52429 , \52430 , \52431 , \52432 ,
         \52433 , \52434 , \52435 , \52436 , \52437 , \52438 , \52439 , \52440 , \52441 , \52442 ,
         \52443 , \52444 , \52445 , \52446 , \52447 , \52448 , \52449 , \52450 , \52451 , \52452 ,
         \52453 , \52454 , \52455 , \52456 , \52457 , \52458 , \52459 , \52460 , \52461 , \52462 ,
         \52463 , \52464 , \52465 , \52466 , \52467 , \52468 , \52469 , \52470 , \52471 , \52472 ,
         \52473 , \52474 , \52475 , \52476 , \52477 , \52478 , \52479 , \52480 , \52481 , \52482 ,
         \52483 , \52484 , \52485 , \52486 , \52487 , \52488 , \52489 , \52490 , \52491 , \52492 ,
         \52493 , \52494 , \52495 , \52496 , \52497 , \52498 , \52499 , \52500 , \52501 , \52502 ,
         \52503 , \52504 , \52505 , \52506 , \52507 , \52508 , \52509 , \52510 , \52511 , \52512 ,
         \52513 , \52514 , \52515 , \52516 , \52517 , \52518 , \52519 , \52520 , \52521 , \52522 ,
         \52523 , \52524 , \52525 , \52526 , \52527 , \52528 , \52529 , \52530 , \52531 , \52532 ,
         \52533 , \52534 , \52535 , \52536 , \52537 , \52538 , \52539 , \52540 , \52541 , \52542 ,
         \52543 , \52544 , \52545 , \52546 , \52547 , \52548 , \52549 , \52550 , \52551 , \52552 ,
         \52553 , \52554 , \52555 , \52556 , \52557 , \52558 , \52559 , \52560 , \52561 , \52562 ,
         \52563 , \52564 , \52565 , \52566 , \52567 , \52568 , \52569 , \52570 , \52571 , \52572 ,
         \52573 , \52574 , \52575 , \52576 , \52577 , \52578 , \52579 , \52580 , \52581 , \52582 ,
         \52583 , \52584 , \52585 , \52586 , \52587 , \52588 , \52589 , \52590 , \52591 , \52592 ,
         \52593 , \52594 , \52595 , \52596 , \52597 , \52598 , \52599 , \52600 , \52601 , \52602 ,
         \52603 , \52604 , \52605 , \52606 , \52607 , \52608 , \52609 , \52610 , \52611 , \52612 ,
         \52613 , \52614 , \52615 , \52616 , \52617 , \52618 , \52619 , \52620 , \52621 , \52622 ,
         \52623 , \52624 , \52625 , \52626 , \52627 , \52628 , \52629 , \52630 , \52631 , \52632 ,
         \52633 , \52634 , \52635 , \52636 , \52637 , \52638 , \52639 , \52640 , \52641 , \52642 ,
         \52643 , \52644 , \52645 , \52646 , \52647 , \52648 , \52649 , \52650 , \52651 , \52652 ,
         \52653 , \52654 , \52655 , \52656 , \52657 , \52658 , \52659 , \52660 , \52661 , \52662 ,
         \52663 , \52664 , \52665 , \52666 , \52667 , \52668 , \52669 , \52670 , \52671 , \52672 ,
         \52673 , \52674 , \52675 , \52676 , \52677 , \52678 , \52679 , \52680 , \52681 , \52682 ,
         \52683 , \52684 , \52685 , \52686 , \52687 , \52688 , \52689 , \52690 , \52691 , \52692 ,
         \52693 , \52694 , \52695 , \52696 , \52697 , \52698 , \52699 , \52700 , \52701 , \52702 ,
         \52703 , \52704 , \52705 , \52706 , \52707 , \52708 , \52709 , \52710 , \52711 , \52712 ,
         \52713 , \52714 , \52715 , \52716 , \52717 , \52718 , \52719 , \52720 , \52721 , \52722 ,
         \52723 , \52724 , \52725 , \52726 , \52727 , \52728 , \52729 , \52730 , \52731 , \52732 ,
         \52733 , \52734 , \52735 , \52736 , \52737 , \52738 , \52739 , \52740 , \52741 , \52742 ,
         \52743 , \52744 , \52745 , \52746 , \52747 , \52748 , \52749 , \52750 , \52751 , \52752 ,
         \52753 , \52754 , \52755 , \52756 , \52757 , \52758 , \52759 , \52760 , \52761 , \52762 ,
         \52763 , \52764 , \52765 , \52766 , \52767 , \52768 , \52769 , \52770 , \52771 , \52772 ,
         \52773 , \52774 , \52775 , \52776 , \52777 , \52778 , \52779 , \52780 , \52781 , \52782 ,
         \52783 , \52784 , \52785 , \52786 , \52787 , \52788 , \52789 , \52790 , \52791 , \52792 ,
         \52793 , \52794 , \52795 , \52796 , \52797 , \52798 , \52799 , \52800 , \52801 , \52802 ,
         \52803 , \52804 , \52805 , \52806 , \52807 , \52808 , \52809 , \52810 , \52811 , \52812 ,
         \52813 , \52814 , \52815 , \52816 , \52817 , \52818 , \52819 , \52820 , \52821 , \52822 ,
         \52823 , \52824 , \52825 , \52826 , \52827 , \52828 , \52829 , \52830 , \52831 , \52832 ,
         \52833 , \52834 , \52835 , \52836 , \52837 , \52838 , \52839 , \52840 , \52841 , \52842 ,
         \52843 , \52844 , \52845 , \52846 , \52847 , \52848 , \52849 , \52850 , \52851 , \52852 ,
         \52853 , \52854 , \52855 , \52856 , \52857 , \52858 , \52859 , \52860 , \52861 , \52862 ,
         \52863 , \52864 , \52865 , \52866 , \52867 , \52868 , \52869 , \52870 , \52871 , \52872 ,
         \52873 , \52874 , \52875 , \52876 , \52877 , \52878 , \52879 , \52880 , \52881 , \52882 ,
         \52883 , \52884 , \52885 , \52886 , \52887 , \52888 , \52889 , \52890 , \52891 , \52892 ,
         \52893 , \52894 , \52895 , \52896 , \52897 , \52898 , \52899 , \52900 , \52901 , \52902 ,
         \52903 , \52904 , \52905 , \52906 , \52907 , \52908 , \52909 , \52910 , \52911 , \52912 ,
         \52913 , \52914 , \52915 , \52916 , \52917 , \52918 , \52919 , \52920 , \52921 , \52922 ,
         \52923 , \52924 , \52925 , \52926 , \52927 , \52928 , \52929 , \52930 , \52931 , \52932 ,
         \52933 , \52934 , \52935 , \52936 , \52937 , \52938 , \52939 , \52940 , \52941 , \52942 ,
         \52943 , \52944 , \52945 , \52946 , \52947 , \52948 , \52949 , \52950 , \52951 , \52952 ,
         \52953 , \52954 , \52955 , \52956 , \52957 , \52958 , \52959 , \52960 , \52961 , \52962 ,
         \52963 , \52964 , \52965 , \52966 , \52967 , \52968 , \52969 , \52970 , \52971 , \52972 ,
         \52973 , \52974 , \52975 , \52976 , \52977 , \52978 , \52979 , \52980 , \52981 , \52982 ,
         \52983 , \52984 , \52985 , \52986 , \52987 , \52988 , \52989 , \52990 , \52991 , \52992 ,
         \52993 , \52994 , \52995 , \52996 , \52997 , \52998 , \52999 , \53000 , \53001 , \53002 ,
         \53003 , \53004 , \53005 , \53006 , \53007 , \53008 , \53009 , \53010 , \53011 , \53012 ,
         \53013 , \53014 , \53015 , \53016 , \53017 , \53018 , \53019 , \53020 , \53021 , \53022 ,
         \53023 , \53024 , \53025 , \53026 , \53027 , \53028 , \53029 , \53030 , \53031 , \53032 ,
         \53033 , \53034 , \53035 , \53036 , \53037 , \53038 , \53039 , \53040 , \53041 , \53042 ,
         \53043 , \53044 , \53045 , \53046 , \53047 , \53048 , \53049 , \53050 , \53051 , \53052 ,
         \53053 , \53054 , \53055 , \53056 , \53057 , \53058 , \53059 , \53060 , \53061 , \53062 ,
         \53063 , \53064 , \53065 , \53066 , \53067 , \53068 , \53069 , \53070 , \53071 , \53072 ,
         \53073 , \53074 , \53075 , \53076 , \53077 , \53078 , \53079 , \53080 , \53081 , \53082 ,
         \53083 , \53084 , \53085 , \53086 , \53087 , \53088 , \53089 , \53090 , \53091 , \53092 ,
         \53093 , \53094 , \53095 , \53096 , \53097 , \53098 , \53099 , \53100 , \53101 , \53102 ,
         \53103 , \53104 , \53105 , \53106 , \53107 , \53108 , \53109 , \53110 , \53111 , \53112 ,
         \53113 , \53114 , \53115 , \53116 , \53117 , \53118 , \53119 , \53120 , \53121 , \53122 ,
         \53123 , \53124 , \53125 , \53126 , \53127 , \53128 , \53129 , \53130 , \53131 , \53132 ,
         \53133 , \53134 , \53135 , \53136 , \53137 , \53138 , \53139 , \53140 , \53141 , \53142 ,
         \53143 , \53144 , \53145 , \53146 , \53147 , \53148 , \53149 , \53150 , \53151 , \53152 ,
         \53153 , \53154 , \53155 , \53156 , \53157 , \53158 , \53159 , \53160 , \53161 , \53162 ,
         \53163 , \53164 , \53165 , \53166 , \53167 , \53168 , \53169 , \53170 , \53171 , \53172 ,
         \53173 , \53174 , \53175 , \53176 , \53177 , \53178 , \53179 , \53180 , \53181 , \53182 ,
         \53183 , \53184 , \53185 , \53186 , \53187 , \53188 , \53189 , \53190 , \53191 , \53192 ,
         \53193 , \53194 , \53195 , \53196 , \53197 , \53198 , \53199 , \53200 , \53201 , \53202 ,
         \53203 , \53204 , \53205 , \53206 , \53207 , \53208 , \53209 , \53210 , \53211 , \53212 ,
         \53213 , \53214 , \53215 , \53216 , \53217 , \53218 , \53219 , \53220 , \53221 , \53222 ,
         \53223 , \53224 , \53225 , \53226 , \53227 , \53228 , \53229 , \53230 , \53231 , \53232 ,
         \53233 , \53234 , \53235 , \53236 , \53237 , \53238 , \53239 , \53240 , \53241 , \53242 ,
         \53243 , \53244 , \53245 , \53246 , \53247 , \53248 , \53249 , \53250 , \53251 , \53252 ,
         \53253 , \53254 , \53255 , \53256 , \53257 , \53258 , \53259 , \53260 , \53261 , \53262 ,
         \53263 , \53264 , \53265 , \53266 , \53267 , \53268 , \53269 , \53270 , \53271 , \53272 ,
         \53273 , \53274 , \53275 , \53276 , \53277 , \53278 , \53279 , \53280 , \53281 , \53282 ,
         \53283 , \53284 , \53285 , \53286 , \53287 , \53288 , \53289 , \53290 , \53291 , \53292 ,
         \53293 , \53294 , \53295 , \53296 , \53297 , \53298 , \53299 , \53300 , \53301 , \53302 ,
         \53303 , \53304 , \53305 , \53306 , \53307 , \53308 , \53309 , \53310 , \53311 , \53312 ,
         \53313 , \53314 , \53315 , \53316 , \53317 , \53318 , \53319 , \53320 , \53321 , \53322 ,
         \53323 , \53324 , \53325 , \53326 , \53327 , \53328 , \53329 , \53330 , \53331 , \53332 ,
         \53333 , \53334 , \53335 , \53336 , \53337 , \53338 , \53339 , \53340 , \53341 , \53342 ,
         \53343 , \53344 , \53345 , \53346 , \53347 , \53348 , \53349 , \53350 , \53351 , \53352 ,
         \53353 , \53354 , \53355 , \53356 , \53357 , \53358 , \53359 , \53360 , \53361 , \53362 ,
         \53363 , \53364 , \53365 , \53366 , \53367 , \53368 , \53369 , \53370 , \53371 , \53372 ,
         \53373 , \53374 , \53375 , \53376 , \53377 , \53378 , \53379 , \53380 , \53381 , \53382 ,
         \53383 , \53384 , \53385 , \53386 , \53387 , \53388 , \53389 , \53390 , \53391 , \53392 ,
         \53393 , \53394 , \53395 , \53396 , \53397 , \53398 , \53399 , \53400 , \53401 , \53402 ,
         \53403 , \53404 , \53405 , \53406 , \53407 , \53408 , \53409 , \53410 , \53411 , \53412 ,
         \53413 , \53414 , \53415 , \53416 , \53417 , \53418 , \53419 , \53420 , \53421 , \53422 ,
         \53423 , \53424 , \53425 , \53426 , \53427 , \53428 , \53429 , \53430 , \53431 , \53432 ,
         \53433 , \53434 , \53435 , \53436 , \53437 , \53438 , \53439 , \53440 , \53441 , \53442 ,
         \53443 , \53444 , \53445 , \53446 , \53447 , \53448 , \53449 , \53450 , \53451 , \53452 ,
         \53453 , \53454 , \53455 , \53456 , \53457 , \53458 , \53459 , \53460 , \53461 , \53462 ,
         \53463 , \53464 , \53465 , \53466 , \53467 , \53468 , \53469 , \53470 , \53471 , \53472 ,
         \53473 , \53474 , \53475 , \53476 , \53477 , \53478 , \53479 , \53480 , \53481 , \53482 ,
         \53483 , \53484 , \53485 , \53486 , \53487 , \53488 , \53489 , \53490 , \53491 , \53492 ,
         \53493 , \53494 , \53495 , \53496 , \53497 , \53498 , \53499 , \53500 , \53501 , \53502 ,
         \53503 , \53504 , \53505 , \53506 , \53507 , \53508 , \53509 , \53510 , \53511 , \53512 ,
         \53513 , \53514 , \53515 , \53516 , \53517 , \53518 , \53519 , \53520 , \53521 , \53522 ,
         \53523 , \53524 , \53525 , \53526 , \53527 , \53528 , \53529 , \53530 , \53531 , \53532 ,
         \53533 , \53534 , \53535 , \53536 , \53537 , \53538 , \53539 , \53540 , \53541 , \53542 ,
         \53543 , \53544 , \53545 , \53546 , \53547 , \53548 , \53549 , \53550 , \53551 , \53552 ,
         \53553 , \53554 , \53555 , \53556 , \53557 , \53558 , \53559 , \53560 , \53561 , \53562 ,
         \53563 , \53564 , \53565 , \53566 , \53567 , \53568 , \53569 , \53570 , \53571 , \53572 ,
         \53573 , \53574 , \53575 , \53576 , \53577 , \53578 , \53579 , \53580 , \53581 , \53582 ,
         \53583 , \53584 , \53585 , \53586 , \53587 , \53588 , \53589 , \53590 , \53591 , \53592 ,
         \53593 , \53594 , \53595 , \53596 , \53597 , \53598 , \53599 , \53600 , \53601 , \53602 ,
         \53603 , \53604 , \53605 , \53606 , \53607 , \53608 , \53609 , \53610 , \53611 , \53612 ,
         \53613 , \53614 , \53615 , \53616 , \53617 , \53618 , \53619 , \53620 , \53621 , \53622 ,
         \53623 , \53624 , \53625 , \53626 , \53627 , \53628 , \53629 , \53630 , \53631 , \53632 ,
         \53633 , \53634 , \53635 , \53636 , \53637 , \53638 , \53639 , \53640 , \53641 , \53642 ,
         \53643 , \53644 , \53645 , \53646 , \53647 , \53648 , \53649 , \53650 , \53651 , \53652 ,
         \53653 , \53654 , \53655 , \53656 , \53657 , \53658 , \53659 , \53660 , \53661 , \53662 ,
         \53663 , \53664 , \53665 , \53666 , \53667 , \53668 , \53669 , \53670 , \53671 , \53672 ,
         \53673 , \53674 , \53675 , \53676 , \53677 , \53678 , \53679 , \53680 , \53681 , \53682 ,
         \53683 , \53684 , \53685 , \53686 , \53687 , \53688 , \53689 , \53690 , \53691 , \53692 ,
         \53693 , \53694 , \53695 , \53696 , \53697 , \53698 , \53699 , \53700 , \53701 , \53702 ,
         \53703 , \53704 , \53705 , \53706 , \53707 , \53708 , \53709 , \53710 , \53711 , \53712 ,
         \53713 , \53714 , \53715 , \53716 , \53717 , \53718 , \53719 , \53720 , \53721 , \53722 ,
         \53723 , \53724 , \53725 , \53726 , \53727 , \53728 , \53729 , \53730 , \53731 , \53732 ,
         \53733 , \53734 , \53735 , \53736 , \53737 , \53738 , \53739 , \53740 , \53741 , \53742 ,
         \53743 , \53744 , \53745 , \53746 , \53747 , \53748 , \53749 , \53750 , \53751 , \53752 ,
         \53753 , \53754 , \53755 , \53756 , \53757 , \53758 , \53759 , \53760 , \53761 , \53762 ,
         \53763 , \53764 , \53765 , \53766 , \53767 , \53768 , \53769 , \53770 , \53771 , \53772 ,
         \53773 , \53774 , \53775 , \53776 , \53777 , \53778 , \53779 , \53780 , \53781 , \53782 ,
         \53783 , \53784 , \53785 , \53786 , \53787 , \53788 , \53789 , \53790 , \53791 , \53792 ,
         \53793 , \53794 , \53795 , \53796 , \53797 , \53798 , \53799 , \53800 , \53801 , \53802 ,
         \53803 , \53804 , \53805 , \53806 , \53807 , \53808 , \53809 , \53810 , \53811 , \53812 ,
         \53813 , \53814 , \53815 , \53816 , \53817 , \53818 , \53819 , \53820 , \53821 , \53822 ,
         \53823 , \53824 , \53825 , \53826 , \53827 , \53828 , \53829 , \53830 , \53831 , \53832 ,
         \53833 , \53834 , \53835 , \53836 , \53837 , \53838 , \53839 , \53840 , \53841 , \53842 ,
         \53843 , \53844 , \53845 , \53846 , \53847 , \53848 , \53849 , \53850 , \53851 , \53852 ,
         \53853 , \53854 , \53855 , \53856 , \53857 , \53858 , \53859 , \53860 , \53861 , \53862 ,
         \53863 , \53864 , \53865 , \53866 , \53867 , \53868 , \53869 , \53870 , \53871 , \53872 ,
         \53873 , \53874 , \53875 , \53876 , \53877 , \53878 , \53879 , \53880 , \53881 , \53882 ,
         \53883 , \53884 , \53885 , \53886 , \53887 , \53888 , \53889 , \53890 , \53891 , \53892 ,
         \53893 , \53894 , \53895 , \53896 , \53897 , \53898 , \53899 , \53900 , \53901 , \53902 ,
         \53903 , \53904 , \53905 , \53906 , \53907 , \53908 , \53909 , \53910 , \53911 , \53912 ,
         \53913 , \53914 , \53915 , \53916 , \53917 , \53918 , \53919 , \53920 , \53921 , \53922 ,
         \53923 , \53924 , \53925 , \53926 , \53927 , \53928 , \53929 , \53930 , \53931 , \53932 ,
         \53933 , \53934 , \53935 , \53936 , \53937 , \53938 , \53939 , \53940 , \53941 , \53942 ,
         \53943 , \53944 , \53945 , \53946 , \53947 , \53948 , \53949 , \53950 , \53951 , \53952 ,
         \53953 , \53954 , \53955 , \53956 , \53957 , \53958 , \53959 , \53960 , \53961 , \53962 ,
         \53963 , \53964 , \53965 , \53966 , \53967 , \53968 , \53969 , \53970 , \53971 , \53972 ,
         \53973 , \53974 , \53975 , \53976 , \53977 , \53978 , \53979 , \53980 , \53981 , \53982 ,
         \53983 , \53984 , \53985 , \53986 , \53987 , \53988 , \53989 , \53990 , \53991 , \53992 ,
         \53993 , \53994 , \53995 , \53996 , \53997 , \53998 , \53999 , \54000 , \54001 , \54002 ,
         \54003 , \54004 , \54005 , \54006 , \54007 , \54008 , \54009 , \54010 , \54011 , \54012 ,
         \54013 , \54014 , \54015 , \54016 , \54017 , \54018 , \54019 , \54020 , \54021 , \54022 ,
         \54023 , \54024 , \54025 , \54026 , \54027 , \54028 , \54029 , \54030 , \54031 , \54032 ,
         \54033 , \54034 , \54035 , \54036 , \54037 , \54038 , \54039 , \54040 , \54041 , \54042 ,
         \54043 , \54044 , \54045 , \54046 , \54047 , \54048 , \54049 , \54050 , \54051 , \54052 ,
         \54053 , \54054 , \54055 , \54056 , \54057 , \54058 , \54059 , \54060 , \54061 , \54062 ,
         \54063 , \54064 , \54065 , \54066 , \54067 , \54068 , \54069 , \54070 , \54071 , \54072 ,
         \54073 , \54074 , \54075 , \54076 , \54077 , \54078 , \54079 , \54080 , \54081 , \54082 ,
         \54083 , \54084 , \54085 , \54086 , \54087 , \54088 , \54089 , \54090 , \54091 , \54092 ,
         \54093 , \54094 , \54095 , \54096 , \54097 , \54098 , \54099 , \54100 , \54101 , \54102 ,
         \54103 , \54104 , \54105 , \54106 , \54107 , \54108 , \54109 , \54110 , \54111 , \54112 ,
         \54113 , \54114 , \54115 , \54116 , \54117 , \54118 , \54119 , \54120 , \54121 , \54122 ,
         \54123 , \54124 , \54125 , \54126 , \54127 , \54128 , \54129 , \54130 , \54131 , \54132 ,
         \54133 , \54134 , \54135 , \54136 , \54137 , \54138 , \54139 , \54140 , \54141 , \54142 ,
         \54143 , \54144 , \54145 , \54146 , \54147 , \54148 , \54149 , \54150 , \54151 , \54152 ,
         \54153 , \54154 , \54155 , \54156 , \54157 , \54158 , \54159 , \54160 , \54161 , \54162 ,
         \54163 , \54164 , \54165 , \54166 , \54167 , \54168 , \54169 , \54170 , \54171 , \54172 ,
         \54173 , \54174 , \54175 , \54176 , \54177 , \54178 , \54179 , \54180 , \54181 , \54182 ,
         \54183 , \54184 , \54185 , \54186 , \54187 , \54188 , \54189 , \54190 , \54191 , \54192 ,
         \54193 , \54194 , \54195 , \54196 , \54197 , \54198 , \54199 , \54200 , \54201 , \54202 ,
         \54203 , \54204 , \54205 , \54206 , \54207 , \54208 , \54209 , \54210 , \54211 , \54212 ,
         \54213 , \54214 , \54215 , \54216 , \54217 , \54218 , \54219 , \54220 , \54221 , \54222 ,
         \54223 , \54224 , \54225 , \54226 , \54227 , \54228 , \54229 , \54230 , \54231 , \54232 ,
         \54233 , \54234 , \54235 , \54236 , \54237 , \54238 , \54239 , \54240 , \54241 , \54242 ,
         \54243 , \54244 , \54245 , \54246 , \54247 , \54248 , \54249 , \54250 , \54251 , \54252 ,
         \54253 , \54254 , \54255 , \54256 , \54257 , \54258 , \54259 , \54260 , \54261 , \54262 ,
         \54263 , \54264 , \54265 , \54266 , \54267 , \54268 , \54269 , \54270 , \54271 , \54272 ,
         \54273 , \54274 , \54275 , \54276 , \54277 , \54278 , \54279 , \54280 , \54281 , \54282 ,
         \54283 , \54284 , \54285 , \54286 , \54287 , \54288 , \54289 , \54290 , \54291 , \54292 ,
         \54293 , \54294 , \54295 , \54296 , \54297 , \54298 , \54299 , \54300 , \54301 , \54302 ,
         \54303 , \54304 , \54305 , \54306 , \54307 , \54308 , \54309 , \54310 , \54311 , \54312 ,
         \54313 , \54314 , \54315 , \54316 , \54317 , \54318 , \54319 , \54320 , \54321 , \54322 ,
         \54323 , \54324 , \54325 , \54326 , \54327 , \54328 , \54329 , \54330 , \54331 , \54332 ,
         \54333 , \54334 , \54335 , \54336 , \54337 , \54338 , \54339 , \54340 , \54341 , \54342 ,
         \54343 , \54344 , \54345 , \54346 , \54347 , \54348 , \54349 , \54350 , \54351 , \54352 ,
         \54353 , \54354 , \54355 , \54356 , \54357 , \54358 , \54359 , \54360 , \54361 , \54362 ,
         \54363 , \54364 , \54365 , \54366 , \54367 , \54368 , \54369 , \54370 , \54371 , \54372 ,
         \54373 , \54374 , \54375 , \54376 , \54377 , \54378 , \54379 , \54380 , \54381 , \54382 ,
         \54383 , \54384 , \54385 , \54386 , \54387 , \54388 , \54389 , \54390 , \54391 , \54392 ,
         \54393 , \54394 , \54395 , \54396 , \54397 , \54398 , \54399 , \54400 , \54401 , \54402 ,
         \54403 , \54404 , \54405 , \54406 , \54407 , \54408 , \54409 , \54410 , \54411 , \54412 ,
         \54413 , \54414 , \54415 , \54416 , \54417 , \54418 , \54419 , \54420 , \54421 , \54422 ,
         \54423 , \54424 , \54425 , \54426 , \54427 , \54428 , \54429 , \54430 , \54431 , \54432 ,
         \54433 , \54434 , \54435 , \54436 , \54437 , \54438 , \54439 , \54440 , \54441 , \54442 ,
         \54443 , \54444 , \54445 , \54446 , \54447 , \54448 , \54449 , \54450 , \54451 , \54452 ,
         \54453 , \54454 , \54455 , \54456 , \54457 , \54458 , \54459 , \54460 , \54461 , \54462 ,
         \54463 , \54464 , \54465 , \54466 , \54467 , \54468 , \54469 , \54470 , \54471 , \54472 ,
         \54473 , \54474 , \54475 , \54476 , \54477 , \54478 , \54479 , \54480 , \54481 , \54482 ,
         \54483 , \54484 , \54485 , \54486 , \54487 , \54488 , \54489 , \54490 , \54491 , \54492 ,
         \54493 , \54494 , \54495 , \54496 , \54497 , \54498 , \54499 , \54500 , \54501 , \54502 ,
         \54503 , \54504 , \54505 , \54506 , \54507 , \54508 , \54509 , \54510 , \54511 , \54512 ,
         \54513 , \54514 , \54515 , \54516 , \54517 , \54518 , \54519 , \54520 , \54521 , \54522 ,
         \54523 , \54524 , \54525 , \54526 , \54527 , \54528 , \54529 , \54530 , \54531 , \54532 ,
         \54533 , \54534 , \54535 , \54536 , \54537 , \54538 , \54539 , \54540 , \54541 , \54542 ,
         \54543 , \54544 , \54545 , \54546 , \54547 , \54548 , \54549 , \54550 , \54551 , \54552 ,
         \54553 , \54554 , \54555 , \54556 , \54557 , \54558 , \54559 , \54560 , \54561 , \54562 ,
         \54563 , \54564 , \54565 , \54566 , \54567 , \54568 , \54569 , \54570 , \54571 , \54572 ,
         \54573 , \54574 , \54575 , \54576 , \54577 , \54578 , \54579 , \54580 , \54581 , \54582 ,
         \54583 , \54584 , \54585 , \54586 , \54587 , \54588 , \54589 , \54590 , \54591 , \54592 ,
         \54593 , \54594 , \54595 , \54596 , \54597 , \54598 , \54599 , \54600 , \54601 , \54602 ,
         \54603 , \54604 , \54605 , \54606 , \54607 , \54608 , \54609 , \54610 , \54611 , \54612 ,
         \54613 , \54614 , \54615 , \54616 , \54617 , \54618 , \54619 , \54620 , \54621 , \54622 ,
         \54623 , \54624 , \54625 , \54626 , \54627 , \54628 , \54629 , \54630 , \54631 , \54632 ,
         \54633 , \54634 , \54635 , \54636 , \54637 , \54638 , \54639 , \54640 , \54641 , \54642 ,
         \54643 , \54644 , \54645 , \54646 , \54647 , \54648 , \54649 , \54650 , \54651 , \54652 ,
         \54653 , \54654 , \54655 , \54656 , \54657 , \54658 , \54659 , \54660 , \54661 , \54662 ,
         \54663 , \54664 , \54665 , \54666 , \54667 , \54668 , \54669 , \54670 , \54671 , \54672 ,
         \54673 , \54674 , \54675 , \54676 , \54677 , \54678 , \54679 , \54680 , \54681 , \54682 ,
         \54683 , \54684 , \54685 , \54686 , \54687 , \54688 , \54689 , \54690 , \54691 , \54692 ,
         \54693 , \54694 , \54695 , \54696 , \54697 , \54698 , \54699 , \54700 , \54701 , \54702 ,
         \54703 , \54704 , \54705 , \54706 , \54707 , \54708 , \54709 , \54710 , \54711 , \54712 ,
         \54713 , \54714 , \54715 , \54716 , \54717 , \54718 , \54719 , \54720 , \54721 , \54722 ,
         \54723 , \54724 , \54725 , \54726 , \54727 , \54728 , \54729 , \54730 , \54731 , \54732 ,
         \54733 , \54734 , \54735 , \54736 , \54737 , \54738 , \54739 , \54740 , \54741 , \54742 ,
         \54743 , \54744 , \54745 , \54746 , \54747 , \54748 , \54749 , \54750 , \54751 , \54752 ,
         \54753 , \54754 , \54755 , \54756 , \54757 , \54758 , \54759 , \54760 , \54761 , \54762 ,
         \54763 , \54764 , \54765 , \54766 , \54767 , \54768 , \54769 , \54770 , \54771 , \54772 ,
         \54773 , \54774 , \54775 , \54776 , \54777 , \54778 , \54779 , \54780 , \54781 , \54782 ,
         \54783 , \54784 , \54785 , \54786 , \54787 , \54788 , \54789 , \54790 , \54791 , \54792 ,
         \54793 , \54794 , \54795 , \54796 , \54797 , \54798 , \54799 , \54800 , \54801 , \54802 ,
         \54803 , \54804 , \54805 , \54806 , \54807 , \54808 , \54809 , \54810 , \54811 , \54812 ,
         \54813 , \54814 , \54815 , \54816 , \54817 , \54818 , \54819 , \54820 , \54821 , \54822 ,
         \54823 , \54824 , \54825 , \54826 , \54827 , \54828 , \54829 , \54830 , \54831 , \54832 ,
         \54833 , \54834 , \54835 , \54836 , \54837 , \54838 , \54839 , \54840 , \54841 , \54842 ,
         \54843 , \54844 , \54845 , \54846 , \54847 , \54848 , \54849 , \54850 , \54851 , \54852 ,
         \54853 , \54854 , \54855 , \54856 , \54857 , \54858 , \54859 , \54860 , \54861 , \54862 ,
         \54863 , \54864 , \54865 , \54866 , \54867 , \54868 , \54869 , \54870 , \54871 , \54872 ,
         \54873 , \54874 , \54875 , \54876 , \54877 , \54878 , \54879 , \54880 , \54881 , \54882 ,
         \54883 , \54884 , \54885 , \54886 , \54887 , \54888 , \54889 , \54890 , \54891 , \54892 ,
         \54893 , \54894 , \54895 , \54896 , \54897 , \54898 , \54899 , \54900 , \54901 , \54902 ,
         \54903 , \54904 , \54905 , \54906 , \54907 , \54908 , \54909 , \54910 , \54911 , \54912 ,
         \54913 , \54914 , \54915 , \54916 , \54917 , \54918 , \54919 , \54920 , \54921 , \54922 ,
         \54923 , \54924 , \54925 , \54926 , \54927 , \54928 , \54929 , \54930 , \54931 , \54932 ,
         \54933 , \54934 , \54935 , \54936 , \54937 , \54938 , \54939 , \54940 , \54941 , \54942 ,
         \54943 , \54944 , \54945 , \54946 , \54947 , \54948 , \54949 , \54950 , \54951 , \54952 ,
         \54953 , \54954 , \54955 , \54956 , \54957 , \54958 , \54959 , \54960 , \54961 , \54962 ,
         \54963 , \54964 , \54965 , \54966 , \54967 , \54968 , \54969 , \54970 , \54971 , \54972 ,
         \54973 , \54974 , \54975 , \54976 , \54977 , \54978 , \54979 , \54980 , \54981 , \54982 ,
         \54983 , \54984 , \54985 , \54986 , \54987 , \54988 , \54989 , \54990 , \54991 , \54992 ,
         \54993 , \54994 , \54995 , \54996 , \54997 , \54998 , \54999 , \55000 , \55001 , \55002 ,
         \55003 , \55004 , \55005 , \55006 , \55007 , \55008 , \55009 , \55010 , \55011 , \55012 ,
         \55013 , \55014 , \55015 , \55016 , \55017 , \55018 , \55019 , \55020 , \55021 , \55022 ,
         \55023 , \55024 , \55025 , \55026 , \55027 , \55028 , \55029 , \55030 , \55031 , \55032 ,
         \55033 , \55034 , \55035 , \55036 , \55037 , \55038 , \55039 , \55040 , \55041 , \55042 ,
         \55043 , \55044 , \55045 , \55046 , \55047 , \55048 , \55049 , \55050 , \55051 , \55052 ,
         \55053 , \55054 , \55055 , \55056 , \55057 , \55058 , \55059 , \55060 , \55061 , \55062 ,
         \55063 , \55064 , \55065 , \55066 , \55067 , \55068 , \55069 , \55070 , \55071 , \55072 ,
         \55073 , \55074 , \55075 , \55076 , \55077 , \55078 , \55079 , \55080 , \55081 , \55082 ,
         \55083 , \55084 , \55085 , \55086 , \55087 , \55088 , \55089 , \55090 , \55091 , \55092 ,
         \55093 , \55094 , \55095 , \55096 , \55097 , \55098 , \55099 , \55100 , \55101 , \55102 ,
         \55103 , \55104 , \55105 , \55106 , \55107 , \55108 , \55109 , \55110 , \55111 , \55112 ,
         \55113 , \55114 , \55115 , \55116 , \55117 , \55118 , \55119 , \55120 , \55121 , \55122 ,
         \55123 , \55124 , \55125 , \55126 , \55127 , \55128 , \55129 , \55130 , \55131 , \55132 ,
         \55133 , \55134 , \55135 , \55136 , \55137 , \55138 , \55139 , \55140 , \55141 , \55142 ,
         \55143 , \55144 , \55145 , \55146 , \55147 , \55148 , \55149 , \55150 , \55151 , \55152 ,
         \55153 , \55154 , \55155 , \55156 , \55157 , \55158 , \55159 , \55160 , \55161 , \55162 ,
         \55163 , \55164 , \55165 , \55166 , \55167 , \55168 , \55169 , \55170 , \55171 , \55172 ,
         \55173 , \55174 , \55175 , \55176 , \55177 , \55178 , \55179 , \55180 , \55181 , \55182 ,
         \55183 , \55184 , \55185 , \55186 , \55187 , \55188 , \55189 , \55190 , \55191 , \55192 ,
         \55193 , \55194 , \55195 , \55196 , \55197 , \55198 , \55199 , \55200 , \55201 , \55202 ,
         \55203 , \55204 , \55205 , \55206 , \55207 , \55208 , \55209 , \55210 , \55211 , \55212 ,
         \55213 , \55214 , \55215 , \55216 , \55217 , \55218 , \55219 , \55220 , \55221 , \55222 ,
         \55223 , \55224 , \55225 , \55226 , \55227 , \55228 , \55229 , \55230 , \55231 , \55232 ,
         \55233 , \55234 , \55235 , \55236 , \55237 , \55238 , \55239 , \55240 , \55241 , \55242 ,
         \55243 , \55244 , \55245 , \55246 , \55247 , \55248 , \55249 , \55250 , \55251 , \55252 ,
         \55253 , \55254 , \55255 , \55256 , \55257 , \55258 , \55259 , \55260 , \55261 , \55262 ,
         \55263 , \55264 , \55265 , \55266 , \55267 , \55268 , \55269 , \55270 , \55271 , \55272 ,
         \55273 , \55274 , \55275 , \55276 , \55277 , \55278 , \55279 , \55280 , \55281 , \55282 ,
         \55283 , \55284 , \55285 , \55286 , \55287 , \55288 , \55289 , \55290 , \55291 , \55292 ,
         \55293 , \55294 , \55295 , \55296 , \55297 , \55298 , \55299 , \55300 , \55301 , \55302 ,
         \55303 , \55304 , \55305 , \55306 , \55307 , \55308 , \55309 , \55310 , \55311 , \55312 ,
         \55313 , \55314 , \55315 , \55316 , \55317 , \55318 , \55319 , \55320 , \55321 , \55322 ,
         \55323 , \55324 , \55325 , \55326 , \55327 , \55328 , \55329 , \55330 , \55331 , \55332 ,
         \55333 , \55334 , \55335 , \55336 , \55337 , \55338 , \55339 , \55340 , \55341 , \55342 ,
         \55343 , \55344 , \55345 , \55346 , \55347 , \55348 , \55349 , \55350 , \55351 , \55352 ,
         \55353 , \55354 , \55355 , \55356 , \55357 , \55358 , \55359 , \55360 , \55361 , \55362 ,
         \55363 , \55364 , \55365 , \55366 , \55367 , \55368 , \55369 , \55370 , \55371 , \55372 ,
         \55373 , \55374 , \55375 , \55376 , \55377 , \55378 , \55379 , \55380 , \55381 , \55382 ,
         \55383 , \55384 , \55385 , \55386 , \55387 , \55388 , \55389 , \55390 , \55391 , \55392 ,
         \55393 , \55394 , \55395 , \55396 , \55397 , \55398 , \55399 , \55400 , \55401 , \55402 ,
         \55403 , \55404 , \55405 , \55406 , \55407 , \55408 , \55409 , \55410 , \55411 , \55412 ,
         \55413 , \55414 , \55415 , \55416 , \55417 , \55418 , \55419 , \55420 , \55421 , \55422 ,
         \55423 , \55424 , \55425 , \55426 , \55427 , \55428 , \55429 , \55430 , \55431 , \55432 ,
         \55433 , \55434 , \55435 , \55436 , \55437 , \55438 , \55439 , \55440 , \55441 , \55442 ,
         \55443 , \55444 , \55445 , \55446 , \55447 , \55448 , \55449 , \55450 , \55451 , \55452 ,
         \55453 , \55454 , \55455 , \55456 , \55457 , \55458 , \55459 , \55460 , \55461 , \55462 ,
         \55463 , \55464 , \55465 , \55466 , \55467 , \55468 , \55469 , \55470 , \55471 , \55472 ,
         \55473 , \55474 , \55475 , \55476 , \55477 , \55478 , \55479 , \55480 , \55481 , \55482 ,
         \55483 , \55484 , \55485 , \55486 , \55487 , \55488 , \55489 , \55490 , \55491 , \55492 ,
         \55493 , \55494 , \55495 , \55496 , \55497 , \55498 , \55499 , \55500 , \55501 , \55502 ,
         \55503 , \55504 , \55505 , \55506 , \55507 , \55508 , \55509 , \55510 , \55511 , \55512 ,
         \55513 , \55514 , \55515 , \55516 , \55517 , \55518 , \55519 , \55520 , \55521 , \55522 ,
         \55523 , \55524 , \55525 , \55526 , \55527 , \55528 , \55529 , \55530 , \55531 , \55532 ,
         \55533 , \55534 , \55535 , \55536 , \55537 , \55538 , \55539 , \55540 , \55541 , \55542 ,
         \55543 , \55544 , \55545 , \55546 , \55547 , \55548 , \55549 , \55550 , \55551 , \55552 ,
         \55553 , \55554 , \55555 , \55556 , \55557 , \55558 , \55559 , \55560 , \55561 , \55562 ,
         \55563 , \55564 , \55565 , \55566 , \55567 , \55568 , \55569 , \55570 , \55571 , \55572 ,
         \55573 , \55574 , \55575 , \55576 , \55577 , \55578 , \55579 , \55580 , \55581 , \55582 ,
         \55583 , \55584 , \55585 , \55586 , \55587 , \55588 , \55589 , \55590 , \55591 , \55592 ,
         \55593 , \55594 , \55595 , \55596 , \55597 , \55598 , \55599 , \55600 , \55601 , \55602 ,
         \55603 , \55604 , \55605 , \55606 , \55607 , \55608 , \55609 , \55610 , \55611 , \55612 ,
         \55613 , \55614 , \55615 , \55616 , \55617 , \55618 , \55619 , \55620 , \55621 , \55622 ,
         \55623 , \55624 , \55625 , \55626 , \55627 , \55628 , \55629 , \55630 , \55631 , \55632 ,
         \55633 , \55634 , \55635 , \55636 , \55637 , \55638 , \55639 , \55640 , \55641 , \55642 ,
         \55643 , \55644 , \55645 , \55646 , \55647 , \55648 , \55649 , \55650 , \55651 , \55652 ,
         \55653 , \55654 , \55655 , \55656 , \55657 , \55658 , \55659 , \55660 , \55661 , \55662 ,
         \55663 , \55664 , \55665 , \55666 , \55667 , \55668 , \55669 , \55670 , \55671 , \55672 ,
         \55673 , \55674 , \55675 , \55676 , \55677 , \55678 , \55679 , \55680 , \55681 , \55682 ,
         \55683 , \55684 , \55685 , \55686 , \55687 , \55688 , \55689 , \55690 , \55691 , \55692 ,
         \55693 , \55694 , \55695 , \55696 , \55697 , \55698 , \55699 , \55700 , \55701 , \55702 ,
         \55703 , \55704 , \55705 , \55706 , \55707 , \55708 , \55709 , \55710 , \55711 , \55712 ,
         \55713 , \55714 , \55715 , \55716 , \55717 , \55718 , \55719 , \55720 , \55721 , \55722 ,
         \55723 , \55724 , \55725 , \55726 , \55727 , \55728 , \55729 , \55730 , \55731 , \55732 ,
         \55733 , \55734 , \55735 , \55736 , \55737 , \55738 , \55739 , \55740 , \55741 , \55742 ,
         \55743 , \55744 , \55745 , \55746 , \55747 , \55748 , \55749 , \55750 , \55751 , \55752 ,
         \55753 , \55754 , \55755 , \55756 , \55757 , \55758 , \55759 , \55760 , \55761 , \55762 ,
         \55763 , \55764 , \55765 , \55766 , \55767 , \55768 , \55769 , \55770 , \55771 , \55772 ,
         \55773 , \55774 , \55775 , \55776 , \55777 , \55778 , \55779 , \55780 , \55781 , \55782 ,
         \55783 , \55784 , \55785 , \55786 , \55787 , \55788 , \55789 , \55790 , \55791 , \55792 ,
         \55793 , \55794 , \55795 , \55796 , \55797 , \55798 , \55799 , \55800 , \55801 , \55802 ,
         \55803 , \55804 , \55805 , \55806 , \55807 , \55808 , \55809 , \55810 , \55811 , \55812 ,
         \55813 , \55814 , \55815 , \55816 , \55817 , \55818 , \55819 , \55820 , \55821 , \55822 ,
         \55823 , \55824 , \55825 , \55826 , \55827 , \55828 , \55829 , \55830 , \55831 , \55832 ,
         \55833 , \55834 , \55835 , \55836 , \55837 , \55838 , \55839 , \55840 , \55841 , \55842 ,
         \55843 , \55844 , \55845 , \55846 , \55847 , \55848 , \55849 , \55850 , \55851 , \55852 ,
         \55853 , \55854 , \55855 , \55856 , \55857 , \55858 , \55859 , \55860 , \55861 , \55862 ,
         \55863 , \55864 , \55865 , \55866 , \55867 , \55868 , \55869 , \55870 , \55871 , \55872 ,
         \55873 , \55874 , \55875 , \55876 , \55877 , \55878 , \55879 , \55880 , \55881 , \55882 ,
         \55883 , \55884 , \55885 , \55886 , \55887 , \55888 , \55889 , \55890 , \55891 , \55892 ,
         \55893 , \55894 , \55895 , \55896 , \55897 , \55898 , \55899 , \55900 , \55901 , \55902 ,
         \55903 , \55904 , \55905 , \55906 , \55907 , \55908 , \55909 , \55910 , \55911 , \55912 ,
         \55913 , \55914 , \55915 , \55916 , \55917 , \55918 , \55919 , \55920 , \55921 , \55922 ,
         \55923 , \55924 , \55925 , \55926 , \55927 , \55928 , \55929 , \55930 , \55931 , \55932 ,
         \55933 , \55934 , \55935 , \55936 , \55937 , \55938 , \55939 , \55940 , \55941 , \55942 ,
         \55943 , \55944 , \55945 , \55946 , \55947 , \55948 , \55949 , \55950 , \55951 , \55952 ,
         \55953 , \55954 , \55955 , \55956 , \55957 , \55958 , \55959 , \55960 , \55961 , \55962 ,
         \55963 , \55964 , \55965 , \55966 , \55967 , \55968 , \55969 , \55970 , \55971 , \55972 ,
         \55973 , \55974 , \55975 , \55976 , \55977 , \55978 , \55979 , \55980 , \55981 , \55982 ,
         \55983 , \55984 , \55985 , \55986 , \55987 , \55988 , \55989 , \55990 , \55991 , \55992 ,
         \55993 , \55994 , \55995 , \55996 , \55997 , \55998 , \55999 , \56000 , \56001 , \56002 ,
         \56003 , \56004 , \56005 , \56006 , \56007 , \56008 , \56009 , \56010 , \56011 , \56012 ,
         \56013 , \56014 , \56015 , \56016 , \56017 , \56018 , \56019 , \56020 , \56021 , \56022 ,
         \56023 , \56024 , \56025 , \56026 , \56027 , \56028 , \56029 , \56030 , \56031 , \56032 ,
         \56033 , \56034 , \56035 , \56036 , \56037 , \56038 , \56039 , \56040 , \56041 , \56042 ,
         \56043 , \56044 , \56045 , \56046 , \56047 , \56048 , \56049 , \56050 , \56051 , \56052 ,
         \56053 , \56054 , \56055 , \56056 , \56057 , \56058 , \56059 , \56060 , \56061 , \56062 ,
         \56063 , \56064 , \56065 , \56066 , \56067 , \56068 , \56069 , \56070 , \56071 , \56072 ,
         \56073 , \56074 , \56075 , \56076 , \56077 , \56078 , \56079 , \56080 , \56081 , \56082 ,
         \56083 , \56084 , \56085 , \56086 , \56087 , \56088 , \56089 , \56090 , \56091 , \56092 ,
         \56093 , \56094 , \56095 , \56096 , \56097 , \56098 , \56099 , \56100 , \56101 , \56102 ,
         \56103 , \56104 , \56105 , \56106 , \56107 , \56108 , \56109 , \56110 , \56111 , \56112 ,
         \56113 , \56114 , \56115 , \56116 , \56117 , \56118 , \56119 , \56120 , \56121 , \56122 ,
         \56123 , \56124 , \56125 , \56126 , \56127 , \56128 , \56129 , \56130 , \56131 , \56132 ,
         \56133 , \56134 , \56135 , \56136 , \56137 , \56138 , \56139 , \56140 , \56141 , \56142 ,
         \56143 , \56144 , \56145 , \56146 , \56147 , \56148 , \56149 , \56150 , \56151 , \56152 ,
         \56153 , \56154 , \56155 , \56156 , \56157 , \56158 , \56159 , \56160 , \56161 , \56162 ,
         \56163 , \56164 , \56165 , \56166 , \56167 , \56168 , \56169 , \56170 , \56171 , \56172 ,
         \56173 , \56174 , \56175 , \56176 , \56177 , \56178 , \56179 , \56180 , \56181 , \56182 ,
         \56183 , \56184 , \56185 , \56186 , \56187 , \56188 , \56189 , \56190 , \56191 , \56192 ,
         \56193 , \56194 , \56195 , \56196 , \56197 , \56198 , \56199 , \56200 , \56201 , \56202 ,
         \56203 , \56204 , \56205 , \56206 , \56207 , \56208 , \56209 , \56210 , \56211 , \56212 ,
         \56213 , \56214 , \56215 , \56216 , \56217 , \56218 , \56219 , \56220 , \56221 , \56222 ,
         \56223 , \56224 , \56225 , \56226 , \56227 , \56228 , \56229 , \56230 , \56231 , \56232 ,
         \56233 , \56234 , \56235 , \56236 , \56237 , \56238 , \56239 , \56240 , \56241 , \56242 ,
         \56243 , \56244 , \56245 , \56246 , \56247 , \56248 , \56249 , \56250 , \56251 , \56252 ,
         \56253 , \56254 , \56255 , \56256 , \56257 , \56258 , \56259 , \56260 , \56261 , \56262 ,
         \56263 , \56264 , \56265 , \56266 , \56267 , \56268 , \56269 , \56270 , \56271 , \56272 ,
         \56273 , \56274 , \56275 , \56276 , \56277 , \56278 , \56279 , \56280 , \56281 , \56282 ,
         \56283 , \56284 , \56285 , \56286 , \56287 , \56288 , \56289 , \56290 , \56291 , \56292 ,
         \56293 , \56294 , \56295 , \56296 , \56297 , \56298 , \56299 , \56300 , \56301 , \56302 ,
         \56303 , \56304 , \56305 , \56306 , \56307 , \56308 , \56309 , \56310 , \56311 , \56312 ,
         \56313 , \56314 , \56315 , \56316 , \56317 , \56318 , \56319 , \56320 , \56321 , \56322 ,
         \56323 , \56324 , \56325 , \56326 , \56327 , \56328 , \56329 , \56330 , \56331 , \56332 ,
         \56333 , \56334 , \56335 , \56336 , \56337 , \56338 , \56339 , \56340 , \56341 , \56342 ,
         \56343 , \56344 , \56345 , \56346 , \56347 , \56348 , \56349 , \56350 , \56351 , \56352 ,
         \56353 , \56354 , \56355 , \56356 , \56357 , \56358 , \56359 , \56360 , \56361 , \56362 ,
         \56363 , \56364 , \56365 , \56366 , \56367 , \56368 , \56369 , \56370 , \56371 , \56372 ,
         \56373 , \56374 , \56375 , \56376 , \56377 , \56378 , \56379 , \56380 , \56381 , \56382 ,
         \56383 , \56384 , \56385 , \56386 , \56387 , \56388 , \56389 , \56390 , \56391 , \56392 ,
         \56393 , \56394 , \56395 , \56396 , \56397 , \56398 , \56399 , \56400 , \56401 , \56402 ,
         \56403 , \56404 , \56405 , \56406 , \56407 , \56408 , \56409 , \56410 , \56411 , \56412 ,
         \56413 , \56414 , \56415 , \56416 , \56417 , \56418 , \56419 , \56420 , \56421 , \56422 ,
         \56423 , \56424 , \56425 , \56426 , \56427 , \56428 , \56429 , \56430 , \56431 , \56432 ,
         \56433 , \56434 , \56435 , \56436 , \56437 , \56438 , \56439 , \56440 , \56441 , \56442 ,
         \56443 , \56444 , \56445 , \56446 , \56447 , \56448 , \56449 , \56450 , \56451 , \56452 ,
         \56453 , \56454 , \56455 , \56456 , \56457 , \56458 , \56459 , \56460 , \56461 , \56462 ,
         \56463 , \56464 , \56465 , \56466 , \56467 , \56468 , \56469 , \56470 , \56471 , \56472 ,
         \56473 , \56474 , \56475 , \56476 , \56477 , \56478 , \56479 , \56480 , \56481 , \56482 ,
         \56483 , \56484 , \56485 , \56486 , \56487 , \56488 , \56489 , \56490 , \56491 , \56492 ,
         \56493 , \56494 , \56495 , \56496 , \56497 , \56498 , \56499 , \56500 , \56501 , \56502 ,
         \56503 , \56504 , \56505 , \56506 , \56507 , \56508 , \56509 , \56510 , \56511 , \56512 ,
         \56513 , \56514 , \56515 , \56516 , \56517 , \56518 , \56519 , \56520 , \56521 , \56522 ,
         \56523 , \56524 , \56525 , \56526 , \56527 , \56528 , \56529 , \56530 , \56531 , \56532 ,
         \56533 , \56534 , \56535 , \56536 , \56537 , \56538 , \56539 , \56540 , \56541 , \56542 ,
         \56543 , \56544 , \56545 , \56546 , \56547 , \56548 , \56549 , \56550 , \56551 , \56552 ,
         \56553 , \56554 , \56555 , \56556 , \56557 , \56558 , \56559 , \56560 , \56561 , \56562 ,
         \56563 , \56564 , \56565 , \56566 , \56567 , \56568 , \56569 , \56570 , \56571 , \56572 ,
         \56573 , \56574 , \56575 , \56576 , \56577 , \56578 , \56579 , \56580 , \56581 , \56582 ,
         \56583 , \56584 , \56585 , \56586 , \56587 , \56588 , \56589 , \56590 , \56591 , \56592 ,
         \56593 , \56594 , \56595 , \56596 , \56597 , \56598 , \56599 , \56600 , \56601 , \56602 ,
         \56603 , \56604 , \56605 , \56606 , \56607 , \56608 , \56609 , \56610 , \56611 , \56612 ,
         \56613 , \56614 , \56615 , \56616 , \56617 , \56618 , \56619 , \56620 , \56621 , \56622 ,
         \56623 , \56624 , \56625 , \56626 , \56627 , \56628 , \56629 , \56630 , \56631 , \56632 ,
         \56633 , \56634 , \56635 , \56636 , \56637 , \56638 , \56639 , \56640 , \56641 , \56642 ,
         \56643 , \56644 , \56645 , \56646 , \56647 , \56648 , \56649 , \56650 , \56651 , \56652 ,
         \56653 , \56654 , \56655 , \56656 , \56657 , \56658 , \56659 , \56660 , \56661 , \56662 ,
         \56663 , \56664 , \56665 , \56666 , \56667 , \56668 , \56669 , \56670 , \56671 , \56672 ,
         \56673 , \56674 , \56675 , \56676 , \56677 , \56678 , \56679 , \56680 , \56681 , \56682 ,
         \56683 , \56684 , \56685 , \56686 , \56687 , \56688 , \56689 , \56690 , \56691 , \56692 ,
         \56693 , \56694 , \56695 , \56696 , \56697 , \56698 , \56699 , \56700 , \56701 , \56702 ,
         \56703 , \56704 , \56705 , \56706 , \56707 , \56708 , \56709 , \56710 , \56711 , \56712 ,
         \56713 , \56714 , \56715 , \56716 , \56717 , \56718 , \56719 , \56720 , \56721 , \56722 ,
         \56723 , \56724 , \56725 , \56726 , \56727 , \56728 , \56729 , \56730 , \56731 , \56732 ,
         \56733 , \56734 , \56735 , \56736 , \56737 , \56738 , \56739 , \56740 , \56741 , \56742 ,
         \56743 , \56744 , \56745 , \56746 , \56747 , \56748 , \56749 , \56750 , \56751 , \56752 ,
         \56753 , \56754 , \56755 , \56756 , \56757 , \56758 , \56759 , \56760 , \56761 , \56762 ,
         \56763 , \56764 , \56765 , \56766 , \56767 , \56768 , \56769 , \56770 , \56771 , \56772 ,
         \56773 , \56774 , \56775 , \56776 , \56777 , \56778 , \56779 , \56780 , \56781 , \56782 ,
         \56783 , \56784 , \56785 , \56786 , \56787 , \56788 , \56789 , \56790 , \56791 , \56792 ,
         \56793 , \56794 , \56795 , \56796 , \56797 , \56798 , \56799 , \56800 , \56801 , \56802 ,
         \56803 , \56804 , \56805 , \56806 , \56807 , \56808 , \56809 , \56810 , \56811 , \56812 ,
         \56813 , \56814 , \56815 , \56816 , \56817 , \56818 , \56819 , \56820 , \56821 , \56822 ,
         \56823 , \56824 , \56825 , \56826 , \56827 , \56828 , \56829 , \56830 , \56831 , \56832 ,
         \56833 , \56834 , \56835 , \56836 , \56837 , \56838 , \56839 , \56840 , \56841 , \56842 ,
         \56843 , \56844 , \56845 , \56846 , \56847 , \56848 , \56849 , \56850 , \56851 , \56852 ,
         \56853 , \56854 , \56855 , \56856 , \56857 , \56858 , \56859 , \56860 , \56861 , \56862 ,
         \56863 , \56864 , \56865 , \56866 , \56867 , \56868 , \56869 , \56870 , \56871 , \56872 ,
         \56873 , \56874 , \56875 , \56876 , \56877 , \56878 , \56879 , \56880 , \56881 , \56882 ,
         \56883 , \56884 , \56885 , \56886 , \56887 , \56888 , \56889 , \56890 , \56891 , \56892 ,
         \56893 , \56894 , \56895 , \56896 , \56897 , \56898 , \56899 , \56900 , \56901 , \56902 ,
         \56903 , \56904 , \56905 , \56906 , \56907 , \56908 , \56909 , \56910 , \56911 , \56912 ,
         \56913 , \56914 , \56915 , \56916 , \56917 , \56918 , \56919 , \56920 , \56921 , \56922 ,
         \56923 , \56924 , \56925 , \56926 , \56927 , \56928 , \56929 , \56930 , \56931 , \56932 ,
         \56933 , \56934 , \56935 , \56936 , \56937 , \56938 , \56939 , \56940 , \56941 , \56942 ,
         \56943 , \56944 , \56945 , \56946 , \56947 , \56948 , \56949 , \56950 , \56951 , \56952 ,
         \56953 , \56954 , \56955 , \56956 , \56957 , \56958 , \56959 , \56960 , \56961 , \56962 ,
         \56963 , \56964 , \56965 , \56966 , \56967 , \56968 , \56969 , \56970 , \56971 , \56972 ,
         \56973 , \56974 , \56975 , \56976 , \56977 , \56978 , \56979 , \56980 , \56981 , \56982 ,
         \56983 , \56984 , \56985 , \56986 , \56987 , \56988 , \56989 , \56990 , \56991 , \56992 ,
         \56993 , \56994 , \56995 , \56996 , \56997 , \56998 , \56999 , \57000 , \57001 , \57002 ,
         \57003 , \57004 , \57005 , \57006 , \57007 , \57008 , \57009 , \57010 , \57011 , \57012 ,
         \57013 , \57014 , \57015 , \57016 , \57017 , \57018 , \57019 , \57020 , \57021 , \57022 ,
         \57023 , \57024 , \57025 , \57026 , \57027 , \57028 , \57029 , \57030 , \57031 , \57032 ,
         \57033 , \57034 , \57035 , \57036 , \57037 , \57038 , \57039 , \57040 , \57041 , \57042 ,
         \57043 , \57044 , \57045 , \57046 , \57047 , \57048 , \57049 , \57050 , \57051 , \57052 ,
         \57053 , \57054 , \57055 , \57056 , \57057 , \57058 , \57059 , \57060 , \57061 , \57062 ,
         \57063 , \57064 , \57065 , \57066 , \57067 , \57068 , \57069 , \57070 , \57071 , \57072 ,
         \57073 , \57074 , \57075 , \57076 , \57077 , \57078 , \57079 , \57080 , \57081 , \57082 ,
         \57083 , \57084 , \57085 , \57086 , \57087 , \57088 , \57089 , \57090 , \57091 , \57092 ,
         \57093 , \57094 , \57095 , \57096 , \57097 , \57098 , \57099 , \57100 , \57101 , \57102 ,
         \57103 , \57104 , \57105 , \57106 , \57107 , \57108 , \57109 , \57110 , \57111 , \57112 ,
         \57113 , \57114 , \57115 , \57116 , \57117 , \57118 , \57119 , \57120 , \57121 , \57122 ,
         \57123 , \57124 , \57125 , \57126 , \57127 , \57128 , \57129 , \57130 , \57131 , \57132 ,
         \57133 , \57134 , \57135 , \57136 , \57137 , \57138 , \57139 , \57140 , \57141 , \57142 ,
         \57143 , \57144 , \57145 , \57146 , \57147 , \57148 , \57149 , \57150 , \57151 , \57152 ,
         \57153 , \57154 , \57155 , \57156 , \57157 , \57158 , \57159 , \57160 , \57161 , \57162 ,
         \57163 , \57164 , \57165 , \57166 , \57167 , \57168 , \57169 , \57170 , \57171 , \57172 ,
         \57173 , \57174 , \57175 , \57176 , \57177 , \57178 , \57179 , \57180 , \57181 , \57182 ,
         \57183 , \57184 , \57185 , \57186 , \57187 , \57188 , \57189 , \57190 , \57191 , \57192 ,
         \57193 , \57194 , \57195 , \57196 , \57197 , \57198 , \57199 , \57200 , \57201 , \57202 ,
         \57203 , \57204 , \57205 , \57206 , \57207 , \57208 , \57209 , \57210 , \57211 , \57212 ,
         \57213 , \57214 , \57215 , \57216 , \57217 , \57218 , \57219 , \57220 , \57221 , \57222 ,
         \57223 , \57224 , \57225 , \57226 , \57227 , \57228 , \57229 , \57230 , \57231 , \57232 ,
         \57233 , \57234 , \57235 , \57236 , \57237 , \57238 , \57239 , \57240 , \57241 , \57242 ,
         \57243 , \57244 , \57245 , \57246 , \57247 , \57248 , \57249 , \57250 , \57251 , \57252 ,
         \57253 , \57254 , \57255 , \57256 , \57257 , \57258 , \57259 , \57260 , \57261 , \57262 ,
         \57263 , \57264 , \57265 , \57266 , \57267 , \57268 , \57269 , \57270 , \57271 , \57272 ,
         \57273 , \57274 , \57275 , \57276 , \57277 , \57278 , \57279 , \57280 , \57281 , \57282 ,
         \57283 , \57284 , \57285 , \57286 , \57287 , \57288 , \57289 , \57290 , \57291 , \57292 ,
         \57293 , \57294 , \57295 , \57296 , \57297 , \57298 , \57299 , \57300 , \57301 , \57302 ,
         \57303 , \57304 , \57305 , \57306 , \57307 , \57308 , \57309 , \57310 , \57311 , \57312 ,
         \57313 , \57314 , \57315 , \57316 , \57317 , \57318 , \57319 , \57320 , \57321 , \57322 ,
         \57323 , \57324 , \57325 , \57326 , \57327 , \57328 , \57329 , \57330 , \57331 , \57332 ,
         \57333 , \57334 , \57335 , \57336 , \57337 , \57338 , \57339 , \57340 , \57341 , \57342 ,
         \57343 , \57344 , \57345 , \57346 , \57347 , \57348 , \57349 , \57350 , \57351 , \57352 ,
         \57353 , \57354 , \57355 , \57356 , \57357 , \57358 , \57359 , \57360 , \57361 , \57362 ,
         \57363 , \57364 , \57365 , \57366 , \57367 , \57368 , \57369 , \57370 , \57371 , \57372 ,
         \57373 , \57374 , \57375 , \57376 , \57377 , \57378 , \57379 , \57380 , \57381 , \57382 ,
         \57383 , \57384 , \57385 , \57386 , \57387 , \57388 , \57389 , \57390 , \57391 , \57392 ,
         \57393 , \57394 , \57395 , \57396 , \57397 , \57398 , \57399 , \57400 , \57401 , \57402 ,
         \57403 , \57404 , \57405 , \57406 , \57407 , \57408 , \57409 , \57410 , \57411 , \57412 ,
         \57413 , \57414 , \57415 , \57416 , \57417 , \57418 , \57419 , \57420 , \57421 , \57422 ,
         \57423 , \57424 , \57425 , \57426 , \57427 , \57428 , \57429 , \57430 , \57431 , \57432 ,
         \57433 , \57434 , \57435 , \57436 , \57437 , \57438 , \57439 , \57440 , \57441 , \57442 ,
         \57443 , \57444 , \57445 , \57446 , \57447 , \57448 , \57449 , \57450 , \57451 , \57452 ,
         \57453 , \57454 , \57455 , \57456 , \57457 , \57458 , \57459 , \57460 , \57461 , \57462 ,
         \57463 , \57464 , \57465 , \57466 , \57467 , \57468 , \57469 , \57470 , \57471 , \57472 ,
         \57473 , \57474 , \57475 , \57476 , \57477 , \57478 , \57479 , \57480 , \57481 , \57482 ,
         \57483 , \57484 , \57485 , \57486 , \57487 , \57488 , \57489 , \57490 , \57491 , \57492 ,
         \57493 , \57494 , \57495 , \57496 , \57497 , \57498 , \57499 , \57500 , \57501 , \57502 ,
         \57503 , \57504 , \57505 , \57506 , \57507 , \57508 , \57509 , \57510 , \57511 , \57512 ,
         \57513 , \57514 , \57515 , \57516 , \57517 , \57518 , \57519 , \57520 , \57521 , \57522 ,
         \57523 , \57524 , \57525 , \57526 , \57527 , \57528 , \57529 , \57530 , \57531 , \57532 ,
         \57533 , \57534 , \57535 , \57536 , \57537 , \57538 , \57539 , \57540 , \57541 , \57542 ,
         \57543 , \57544 , \57545 , \57546 , \57547 , \57548 , \57549 , \57550 , \57551 , \57552 ,
         \57553 , \57554 , \57555 , \57556 , \57557 , \57558 , \57559 , \57560 , \57561 , \57562 ,
         \57563 , \57564 , \57565 , \57566 , \57567 , \57568 , \57569 , \57570 , \57571 , \57572 ,
         \57573 , \57574 , \57575 , \57576 , \57577 , \57578 , \57579 , \57580 , \57581 , \57582 ,
         \57583 , \57584 , \57585 , \57586 , \57587 , \57588 , \57589 , \57590 , \57591 , \57592 ,
         \57593 , \57594 , \57595 , \57596 , \57597 , \57598 , \57599 , \57600 , \57601 , \57602 ,
         \57603 , \57604 , \57605 , \57606 , \57607 , \57608 , \57609 , \57610 , \57611 , \57612 ,
         \57613 , \57614 , \57615 , \57616 , \57617 , \57618 , \57619 , \57620 , \57621 , \57622 ,
         \57623 , \57624 , \57625 , \57626 , \57627 , \57628 , \57629 , \57630 , \57631 , \57632 ,
         \57633 , \57634 , \57635 , \57636 , \57637 , \57638 , \57639 , \57640 , \57641 , \57642 ,
         \57643 , \57644 , \57645 , \57646 , \57647 , \57648 , \57649 , \57650 , \57651 , \57652 ,
         \57653 , \57654 , \57655 , \57656 , \57657 , \57658 , \57659 , \57660 , \57661 , \57662 ,
         \57663 , \57664 , \57665 , \57666 , \57667 , \57668 , \57669 , \57670 , \57671 , \57672 ,
         \57673 , \57674 , \57675 , \57676 , \57677 , \57678 , \57679 , \57680 , \57681 , \57682 ,
         \57683 , \57684 , \57685 , \57686 , \57687 , \57688 , \57689 , \57690 , \57691 , \57692 ,
         \57693 , \57694 , \57695 , \57696 , \57697 , \57698 , \57699 , \57700 , \57701 , \57702 ,
         \57703 , \57704 , \57705 , \57706 , \57707 , \57708 , \57709 , \57710 , \57711 , \57712 ,
         \57713 , \57714 , \57715 , \57716 , \57717 , \57718 , \57719 , \57720 , \57721 , \57722 ,
         \57723 , \57724 , \57725 , \57726 , \57727 , \57728 , \57729 , \57730 , \57731 , \57732 ,
         \57733 , \57734 , \57735 , \57736 , \57737 , \57738 , \57739 , \57740 , \57741 , \57742 ,
         \57743 , \57744 , \57745 , \57746 , \57747 , \57748 , \57749 , \57750 , \57751 , \57752 ,
         \57753 , \57754 , \57755 , \57756 , \57757 , \57758 , \57759 , \57760 , \57761 , \57762 ,
         \57763 , \57764 , \57765 , \57766 , \57767 , \57768 , \57769 , \57770 , \57771 , \57772 ,
         \57773 , \57774 , \57775 , \57776 , \57777 , \57778 , \57779 , \57780 , \57781 , \57782 ,
         \57783 , \57784 , \57785 , \57786 , \57787 , \57788 , \57789 , \57790 , \57791 , \57792 ,
         \57793 , \57794 , \57795 , \57796 , \57797 , \57798 , \57799 , \57800 , \57801 , \57802 ,
         \57803 , \57804 , \57805 , \57806 , \57807 , \57808 , \57809 , \57810 , \57811 , \57812 ,
         \57813 , \57814 , \57815 , \57816 , \57817 , \57818 , \57819 , \57820 , \57821 , \57822 ,
         \57823 , \57824 , \57825 , \57826 , \57827 , \57828 , \57829 , \57830 , \57831 , \57832 ,
         \57833 , \57834 , \57835 , \57836 , \57837 , \57838 , \57839 , \57840 , \57841 , \57842 ,
         \57843 , \57844 , \57845 , \57846 , \57847 , \57848 , \57849 , \57850 , \57851 , \57852 ,
         \57853 , \57854 , \57855 , \57856 , \57857 , \57858 , \57859 , \57860 , \57861 , \57862 ,
         \57863 , \57864 , \57865 , \57866 , \57867 , \57868 , \57869 , \57870 , \57871 , \57872 ,
         \57873 , \57874 , \57875 , \57876 , \57877 , \57878 , \57879 , \57880 , \57881 , \57882 ,
         \57883 , \57884 , \57885 , \57886 , \57887 , \57888 , \57889 , \57890 , \57891 , \57892 ,
         \57893 , \57894 , \57895 , \57896 , \57897 , \57898 , \57899 , \57900 , \57901 , \57902 ,
         \57903 , \57904 , \57905 , \57906 , \57907 , \57908 , \57909 , \57910 , \57911 , \57912 ,
         \57913 , \57914 , \57915 , \57916 , \57917 , \57918 , \57919 , \57920 , \57921 , \57922 ,
         \57923 , \57924 , \57925 , \57926 , \57927 , \57928 , \57929 , \57930 , \57931 , \57932 ,
         \57933 , \57934 , \57935 , \57936 , \57937 , \57938 , \57939 , \57940 , \57941 , \57942 ,
         \57943 , \57944 , \57945 , \57946 , \57947 , \57948 , \57949 , \57950 , \57951 , \57952 ,
         \57953 , \57954 , \57955 , \57956 , \57957 , \57958 , \57959 , \57960 , \57961 , \57962 ,
         \57963 , \57964 , \57965 , \57966 , \57967 , \57968 , \57969 , \57970 , \57971 , \57972 ,
         \57973 , \57974 , \57975 , \57976 , \57977 , \57978 , \57979 , \57980 , \57981 , \57982 ,
         \57983 , \57984 , \57985 , \57986 , \57987 , \57988 , \57989 , \57990 , \57991 , \57992 ,
         \57993 , \57994 , \57995 , \57996 , \57997 , \57998 , \57999 , \58000 , \58001 , \58002 ,
         \58003 , \58004 , \58005 , \58006 , \58007 , \58008 , \58009 , \58010 , \58011 , \58012 ,
         \58013 , \58014 , \58015 , \58016 , \58017 , \58018 , \58019 , \58020 , \58021 , \58022 ,
         \58023 , \58024 , \58025 , \58026 , \58027 , \58028 , \58029 , \58030 , \58031 , \58032 ,
         \58033 , \58034 , \58035 , \58036 , \58037 , \58038 , \58039 , \58040 , \58041 , \58042 ,
         \58043 , \58044 , \58045 , \58046 , \58047 , \58048 , \58049 , \58050 , \58051 , \58052 ,
         \58053 , \58054 , \58055 , \58056 , \58057 , \58058 , \58059 , \58060 , \58061 , \58062 ,
         \58063 , \58064 , \58065 , \58066 , \58067 , \58068 , \58069 , \58070 , \58071 , \58072 ,
         \58073 , \58074 , \58075 , \58076 , \58077 , \58078 , \58079 , \58080 , \58081 , \58082 ,
         \58083 , \58084 , \58085 , \58086 , \58087 , \58088 , \58089 , \58090 , \58091 , \58092 ,
         \58093 , \58094 , \58095 , \58096 , \58097 , \58098 , \58099 , \58100 , \58101 , \58102 ,
         \58103 , \58104 , \58105 , \58106 , \58107 , \58108 , \58109 , \58110 , \58111 , \58112 ,
         \58113 , \58114 , \58115 , \58116 , \58117 , \58118 , \58119 , \58120 , \58121 , \58122 ,
         \58123 , \58124 , \58125 , \58126 , \58127 , \58128 , \58129 , \58130 , \58131 , \58132 ,
         \58133 , \58134 , \58135 , \58136 , \58137 , \58138 , \58139 , \58140 , \58141 , \58142 ,
         \58143 , \58144 , \58145 , \58146 , \58147 , \58148 , \58149 , \58150 , \58151 , \58152 ,
         \58153 , \58154 , \58155 , \58156 , \58157 , \58158 , \58159 , \58160 , \58161 , \58162 ,
         \58163 , \58164 , \58165 , \58166 , \58167 , \58168 , \58169 , \58170 , \58171 , \58172 ,
         \58173 , \58174 , \58175 , \58176 , \58177 , \58178 , \58179 , \58180 , \58181 , \58182 ,
         \58183 , \58184 , \58185 , \58186 , \58187 , \58188 , \58189 , \58190 , \58191 , \58192 ,
         \58193 , \58194 , \58195 , \58196 , \58197 , \58198 , \58199 , \58200 , \58201 , \58202 ,
         \58203 , \58204 , \58205 , \58206 , \58207 , \58208 , \58209 , \58210 , \58211 , \58212 ,
         \58213 , \58214 , \58215 , \58216 , \58217 , \58218 , \58219 , \58220 , \58221 , \58222 ,
         \58223 , \58224 , \58225 , \58226 , \58227 , \58228 , \58229 , \58230 , \58231 , \58232 ,
         \58233 , \58234 , \58235 , \58236 , \58237 , \58238 , \58239 , \58240 , \58241 , \58242 ,
         \58243 , \58244 , \58245 , \58246 , \58247 , \58248 , \58249 , \58250 , \58251 , \58252 ,
         \58253 , \58254 , \58255 , \58256 , \58257 , \58258 , \58259 , \58260 , \58261 , \58262 ,
         \58263 , \58264 , \58265 , \58266 , \58267 , \58268 , \58269 , \58270 , \58271 , \58272 ,
         \58273 , \58274 , \58275 , \58276 , \58277 , \58278 , \58279 , \58280 , \58281 , \58282 ,
         \58283 , \58284 , \58285 , \58286 , \58287 , \58288 , \58289 , \58290 , \58291 , \58292 ,
         \58293 , \58294 , \58295 , \58296 , \58297 , \58298 , \58299 , \58300 , \58301 , \58302 ,
         \58303 , \58304 , \58305 , \58306 , \58307 , \58308 , \58309 , \58310 , \58311 , \58312 ,
         \58313 , \58314 , \58315 , \58316 , \58317 , \58318 , \58319 , \58320 , \58321 , \58322 ,
         \58323 , \58324 , \58325 , \58326 , \58327 , \58328 , \58329 , \58330 , \58331 , \58332 ,
         \58333 , \58334 , \58335 , \58336 , \58337 , \58338 , \58339 , \58340 , \58341 , \58342 ,
         \58343 , \58344 , \58345 , \58346 , \58347 , \58348 , \58349 , \58350 , \58351 , \58352 ,
         \58353 , \58354 , \58355 , \58356 , \58357 , \58358 , \58359 , \58360 , \58361 , \58362 ,
         \58363 , \58364 , \58365 , \58366 , \58367 , \58368 , \58369 , \58370 , \58371 , \58372 ,
         \58373 , \58374 , \58375 , \58376 , \58377 , \58378 , \58379 , \58380 , \58381 , \58382 ,
         \58383 , \58384 , \58385 , \58386 , \58387 , \58388 , \58389 , \58390 , \58391 , \58392 ,
         \58393 , \58394 , \58395 , \58396 , \58397 , \58398 , \58399 , \58400 , \58401 , \58402 ,
         \58403 , \58404 , \58405 , \58406 , \58407 , \58408 , \58409 , \58410 , \58411 , \58412 ,
         \58413 , \58414 , \58415 , \58416 , \58417 , \58418 , \58419 , \58420 , \58421 , \58422 ,
         \58423 , \58424 , \58425 , \58426 , \58427 , \58428 , \58429 , \58430 , \58431 , \58432 ,
         \58433 , \58434 , \58435 , \58436 , \58437 , \58438 , \58439 , \58440 , \58441 , \58442 ,
         \58443 , \58444 , \58445 , \58446 , \58447 , \58448 , \58449 , \58450 , \58451 , \58452 ,
         \58453 , \58454 , \58455 , \58456 , \58457 , \58458 , \58459 , \58460 , \58461 , \58462 ,
         \58463 , \58464 , \58465 , \58466 , \58467 , \58468 , \58469 , \58470 , \58471 , \58472 ,
         \58473 , \58474 , \58475 , \58476 , \58477 , \58478 , \58479 , \58480 , \58481 , \58482 ,
         \58483 , \58484 , \58485 , \58486 , \58487 , \58488 , \58489 , \58490 , \58491 , \58492 ,
         \58493 , \58494 , \58495 , \58496 , \58497 , \58498 , \58499 , \58500 , \58501 , \58502 ,
         \58503 , \58504 , \58505 , \58506 , \58507 , \58508 , \58509 , \58510 , \58511 , \58512 ,
         \58513 , \58514 , \58515 , \58516 , \58517 , \58518 , \58519 , \58520 , \58521 , \58522 ,
         \58523 , \58524 , \58525 , \58526 , \58527 , \58528 , \58529 , \58530 , \58531 , \58532 ,
         \58533 , \58534 , \58535 , \58536 , \58537 , \58538 , \58539 , \58540 , \58541 , \58542 ,
         \58543 , \58544 , \58545 , \58546 , \58547 , \58548 , \58549 , \58550 , \58551 , \58552 ,
         \58553 , \58554 , \58555 , \58556 , \58557 , \58558 , \58559 , \58560 , \58561 , \58562 ,
         \58563 , \58564 , \58565 , \58566 , \58567 , \58568 , \58569 , \58570 , \58571 , \58572 ,
         \58573 , \58574 , \58575 , \58576 , \58577 , \58578 , \58579 , \58580 , \58581 , \58582 ,
         \58583 , \58584 , \58585 , \58586 , \58587 , \58588 , \58589 , \58590 , \58591 , \58592 ,
         \58593 , \58594 , \58595 , \58596 , \58597 , \58598 , \58599 , \58600 , \58601 , \58602 ,
         \58603 , \58604 , \58605 , \58606 , \58607 , \58608 , \58609 , \58610 , \58611 , \58612 ,
         \58613 , \58614 , \58615 , \58616 , \58617 , \58618 , \58619 , \58620 , \58621 , \58622 ,
         \58623 , \58624 , \58625 , \58626 , \58627 , \58628 , \58629 , \58630 , \58631 , \58632 ,
         \58633 , \58634 , \58635 , \58636 , \58637 , \58638 , \58639 , \58640 , \58641 , \58642 ,
         \58643 , \58644 , \58645 , \58646 , \58647 , \58648 , \58649 , \58650 , \58651 , \58652 ,
         \58653 , \58654 , \58655 , \58656 , \58657 , \58658 , \58659 , \58660 , \58661 , \58662 ,
         \58663 , \58664 , \58665 , \58666 , \58667 , \58668 , \58669 , \58670 , \58671 , \58672 ,
         \58673 , \58674 , \58675 , \58676 , \58677 , \58678 , \58679 , \58680 , \58681 , \58682 ,
         \58683 , \58684 , \58685 , \58686 , \58687 , \58688 , \58689 , \58690 , \58691 , \58692 ,
         \58693 , \58694 , \58695 , \58696 , \58697 , \58698 , \58699 , \58700 , \58701 , \58702 ,
         \58703 , \58704 , \58705 , \58706 , \58707 , \58708 , \58709 , \58710 , \58711 , \58712 ,
         \58713 , \58714 , \58715 , \58716 , \58717 , \58718 , \58719 , \58720 , \58721 , \58722 ,
         \58723 , \58724 , \58725 , \58726 , \58727 , \58728 , \58729 , \58730 , \58731 , \58732 ,
         \58733 , \58734 , \58735 , \58736 , \58737 , \58738 , \58739 , \58740 , \58741 , \58742 ,
         \58743 , \58744 , \58745 , \58746 , \58747 , \58748 , \58749 , \58750 , \58751 , \58752 ,
         \58753 , \58754 , \58755 , \58756 , \58757 , \58758 , \58759 , \58760 , \58761 , \58762 ,
         \58763 , \58764 , \58765 , \58766 , \58767 , \58768 , \58769 , \58770 , \58771 , \58772 ,
         \58773 , \58774 , \58775 , \58776 , \58777 , \58778 , \58779 , \58780 , \58781 , \58782 ,
         \58783 , \58784 , \58785 , \58786 , \58787 , \58788 , \58789 , \58790 , \58791 , \58792 ,
         \58793 , \58794 , \58795 , \58796 , \58797 , \58798 , \58799 , \58800 , \58801 , \58802 ,
         \58803 , \58804 , \58805 , \58806 , \58807 , \58808 , \58809 , \58810 , \58811 , \58812 ,
         \58813 , \58814 , \58815 , \58816 , \58817 , \58818 , \58819 , \58820 , \58821 , \58822 ,
         \58823 , \58824 , \58825 , \58826 , \58827 , \58828 , \58829 , \58830 , \58831 , \58832 ,
         \58833 , \58834 , \58835 , \58836 , \58837 , \58838 , \58839 , \58840 , \58841 , \58842 ,
         \58843 , \58844 , \58845 , \58846 , \58847 , \58848 , \58849 , \58850 , \58851 , \58852 ,
         \58853 , \58854 , \58855 , \58856 , \58857 , \58858 , \58859 , \58860 , \58861 , \58862 ,
         \58863 , \58864 , \58865 , \58866 , \58867 , \58868 , \58869 , \58870 , \58871 , \58872 ,
         \58873 , \58874 , \58875 , \58876 , \58877 , \58878 , \58879 , \58880 , \58881 , \58882 ,
         \58883 , \58884 , \58885 , \58886 , \58887 , \58888 , \58889 , \58890 , \58891 , \58892 ,
         \58893 , \58894 , \58895 , \58896 , \58897 , \58898 , \58899 , \58900 , \58901 , \58902 ,
         \58903 , \58904 , \58905 , \58906 , \58907 , \58908 , \58909 , \58910 , \58911 , \58912 ,
         \58913 , \58914 , \58915 , \58916 , \58917 , \58918 , \58919 , \58920 , \58921 , \58922 ,
         \58923 , \58924 , \58925 , \58926 , \58927 , \58928 , \58929 , \58930 , \58931 , \58932 ,
         \58933 , \58934 , \58935 , \58936 , \58937 , \58938 , \58939 , \58940 , \58941 , \58942 ,
         \58943 , \58944 , \58945 , \58946 , \58947 , \58948 , \58949 , \58950 , \58951 , \58952 ,
         \58953 , \58954 , \58955 , \58956 , \58957 , \58958 , \58959 , \58960 , \58961 , \58962 ,
         \58963 , \58964 , \58965 , \58966 , \58967 , \58968 , \58969 , \58970 , \58971 , \58972 ,
         \58973 , \58974 , \58975 , \58976 , \58977 , \58978 , \58979 , \58980 , \58981 , \58982 ,
         \58983 , \58984 , \58985 , \58986 , \58987 , \58988 , \58989 , \58990 , \58991 , \58992 ,
         \58993 , \58994 , \58995 , \58996 , \58997 , \58998 , \58999 , \59000 , \59001 , \59002 ,
         \59003 , \59004 , \59005 , \59006 , \59007 , \59008 , \59009 , \59010 , \59011 , \59012 ,
         \59013 , \59014 , \59015 , \59016 , \59017 , \59018 , \59019 , \59020 , \59021 , \59022 ,
         \59023 , \59024 , \59025 , \59026 , \59027 , \59028 , \59029 , \59030 , \59031 , \59032 ,
         \59033 , \59034 , \59035 , \59036 , \59037 , \59038 , \59039 , \59040 , \59041 , \59042 ,
         \59043 , \59044 , \59045 , \59046 , \59047 , \59048 , \59049 , \59050 , \59051 , \59052 ,
         \59053 , \59054 , \59055 , \59056 , \59057 , \59058 , \59059 , \59060 , \59061 , \59062 ,
         \59063 , \59064 , \59065 , \59066 , \59067 , \59068 , \59069 , \59070 , \59071 , \59072 ,
         \59073 , \59074 , \59075 , \59076 , \59077 , \59078 , \59079 , \59080 , \59081 , \59082 ,
         \59083 , \59084 , \59085 , \59086 , \59087 , \59088 , \59089 , \59090 , \59091 , \59092 ,
         \59093 , \59094 , \59095 , \59096 , \59097 , \59098 , \59099 , \59100 , \59101 , \59102 ,
         \59103 , \59104 , \59105 , \59106 , \59107 , \59108 , \59109 , \59110 , \59111 , \59112 ,
         \59113 , \59114 , \59115 , \59116 , \59117 , \59118 , \59119 , \59120 , \59121 , \59122 ,
         \59123 , \59124 , \59125 , \59126 , \59127 , \59128 , \59129 , \59130 , \59131 , \59132 ,
         \59133 , \59134 , \59135 , \59136 , \59137 , \59138 , \59139 , \59140 , \59141 , \59142 ,
         \59143 , \59144 , \59145 , \59146 , \59147 , \59148 , \59149 , \59150 , \59151 , \59152 ,
         \59153 , \59154 , \59155 , \59156 , \59157 , \59158 , \59159 , \59160 , \59161 , \59162 ,
         \59163 , \59164 , \59165 , \59166 , \59167 , \59168 , \59169 , \59170 , \59171 , \59172 ,
         \59173 , \59174 , \59175 , \59176 , \59177 , \59178 , \59179 , \59180 , \59181 , \59182 ,
         \59183 , \59184 , \59185 , \59186 , \59187 , \59188 , \59189 , \59190 , \59191 , \59192 ,
         \59193 , \59194 , \59195 , \59196 , \59197 , \59198 , \59199 , \59200 , \59201 , \59202 ,
         \59203 , \59204 , \59205 , \59206 , \59207 , \59208 , \59209 , \59210 , \59211 , \59212 ,
         \59213 , \59214 , \59215 , \59216 , \59217 , \59218 , \59219 , \59220 , \59221 , \59222 ,
         \59223 , \59224 , \59225 , \59226 , \59227 , \59228 , \59229 , \59230 , \59231 , \59232 ,
         \59233 , \59234 , \59235 , \59236 , \59237 , \59238 , \59239 , \59240 , \59241 , \59242 ,
         \59243 , \59244 , \59245 , \59246 , \59247 , \59248 , \59249 , \59250 , \59251 , \59252 ,
         \59253 , \59254 , \59255 , \59256 , \59257 , \59258 , \59259 , \59260 , \59261 , \59262 ,
         \59263 , \59264 , \59265 , \59266 , \59267 , \59268 , \59269 , \59270 , \59271 , \59272 ,
         \59273 , \59274 , \59275 , \59276 , \59277 , \59278 , \59279 , \59280 , \59281 , \59282 ,
         \59283 , \59284 , \59285 , \59286 , \59287 , \59288 , \59289 , \59290 , \59291 , \59292 ,
         \59293 , \59294 , \59295 , \59296 , \59297 , \59298 , \59299 , \59300 , \59301 , \59302 ,
         \59303 , \59304 , \59305 , \59306 , \59307 , \59308 , \59309 , \59310 , \59311 , \59312 ,
         \59313 , \59314 , \59315 , \59316 , \59317 , \59318 , \59319 , \59320 , \59321 , \59322 ,
         \59323 , \59324 , \59325 , \59326 , \59327 , \59328 , \59329 , \59330 , \59331 , \59332 ,
         \59333 , \59334 , \59335 , \59336 , \59337 , \59338 , \59339 , \59340 , \59341 , \59342 ,
         \59343 , \59344 , \59345 , \59346 , \59347 , \59348 , \59349 , \59350 , \59351 , \59352 ,
         \59353 , \59354 , \59355 , \59356 , \59357 , \59358 , \59359 , \59360 , \59361 , \59362 ,
         \59363 , \59364 , \59365 , \59366 , \59367 , \59368 , \59369 , \59370 , \59371 , \59372 ,
         \59373 , \59374 , \59375 , \59376 , \59377 , \59378 , \59379 , \59380 , \59381 , \59382 ,
         \59383 , \59384 , \59385 , \59386 , \59387 , \59388 , \59389 , \59390 , \59391 , \59392 ,
         \59393 , \59394 , \59395 , \59396 , \59397 , \59398 , \59399 , \59400 , \59401 , \59402 ,
         \59403 , \59404 , \59405 , \59406 , \59407 , \59408 , \59409 , \59410 , \59411 , \59412 ,
         \59413 , \59414 , \59415 , \59416 , \59417 , \59418 , \59419 , \59420 , \59421 , \59422 ,
         \59423 , \59424 , \59425 , \59426 , \59427 , \59428 , \59429 , \59430 , \59431 , \59432 ,
         \59433 , \59434 , \59435 , \59436 , \59437 , \59438 , \59439 , \59440 , \59441 , \59442 ,
         \59443 , \59444 , \59445 , \59446 , \59447 , \59448 , \59449 , \59450 , \59451 , \59452 ,
         \59453 , \59454 , \59455 , \59456 , \59457 , \59458 , \59459 , \59460 , \59461 , \59462 ,
         \59463 , \59464 , \59465 , \59466 , \59467 , \59468 , \59469 , \59470 , \59471 , \59472 ,
         \59473 , \59474 , \59475 , \59476 , \59477 , \59478 , \59479 , \59480 , \59481 , \59482 ,
         \59483 , \59484 , \59485 , \59486 , \59487 , \59488 , \59489 , \59490 , \59491 , \59492 ,
         \59493 , \59494 , \59495 , \59496 , \59497 , \59498 , \59499 , \59500 , \59501 , \59502 ,
         \59503 , \59504 , \59505 , \59506 , \59507 , \59508 , \59509 , \59510 , \59511 , \59512 ,
         \59513 , \59514 , \59515 , \59516 , \59517 , \59518 , \59519 , \59520 , \59521 , \59522 ,
         \59523 , \59524 , \59525 , \59526 , \59527 , \59528 , \59529 , \59530 , \59531 , \59532 ,
         \59533 , \59534 , \59535 , \59536 , \59537 , \59538 , \59539 , \59540 , \59541 , \59542 ,
         \59543 , \59544 , \59545 , \59546 , \59547 , \59548 , \59549 , \59550 , \59551 , \59552 ,
         \59553 , \59554 , \59555 , \59556 , \59557 , \59558 , \59559 , \59560 , \59561 , \59562 ,
         \59563 , \59564 , \59565 , \59566 , \59567 , \59568 , \59569 , \59570 , \59571 , \59572 ,
         \59573 , \59574 , \59575 , \59576 , \59577 , \59578 , \59579 , \59580 , \59581 , \59582 ,
         \59583 , \59584 , \59585 , \59586 , \59587 , \59588 , \59589 , \59590 , \59591 , \59592 ,
         \59593 , \59594 , \59595 , \59596 , \59597 , \59598 , \59599 , \59600 , \59601 , \59602 ,
         \59603 , \59604 , \59605 , \59606 , \59607 , \59608 , \59609 , \59610 , \59611 , \59612 ,
         \59613 , \59614 , \59615 , \59616 , \59617 , \59618 , \59619 , \59620 , \59621 , \59622 ,
         \59623 , \59624 , \59625 , \59626 , \59627 , \59628 , \59629 , \59630 , \59631 , \59632 ,
         \59633 , \59634 , \59635 , \59636 , \59637 , \59638 , \59639 , \59640 , \59641 , \59642 ,
         \59643 , \59644 , \59645 , \59646 , \59647 , \59648 , \59649 , \59650 , \59651 , \59652 ,
         \59653 , \59654 , \59655 , \59656 , \59657 , \59658 , \59659 , \59660 , \59661 , \59662 ,
         \59663 , \59664 , \59665 , \59666 , \59667 , \59668 , \59669 , \59670 , \59671 , \59672 ,
         \59673 , \59674 , \59675 , \59676 , \59677 , \59678 , \59679 , \59680 , \59681 , \59682 ,
         \59683 , \59684 , \59685 , \59686 , \59687 , \59688 , \59689 , \59690 , \59691 , \59692 ,
         \59693 , \59694 , \59695 , \59696 , \59697 , \59698 , \59699 , \59700 , \59701 , \59702 ,
         \59703 , \59704 , \59705 , \59706 , \59707 , \59708 , \59709 , \59710 , \59711 , \59712 ,
         \59713 , \59714 , \59715 , \59716 , \59717 , \59718 , \59719 , \59720 , \59721 , \59722 ,
         \59723 , \59724 , \59725 , \59726 , \59727 , \59728 , \59729 , \59730 , \59731 , \59732 ,
         \59733 , \59734 , \59735 , \59736 , \59737 , \59738 , \59739 , \59740 , \59741 , \59742 ,
         \59743 , \59744 , \59745 , \59746 , \59747 , \59748 , \59749 , \59750 , \59751 , \59752 ,
         \59753 , \59754 , \59755 , \59756 , \59757 , \59758 , \59759 , \59760 , \59761 , \59762 ,
         \59763 , \59764 , \59765 , \59766 , \59767 , \59768 , \59769 , \59770 , \59771 , \59772 ,
         \59773 , \59774 , \59775 , \59776 , \59777 , \59778 , \59779 , \59780 , \59781 , \59782 ,
         \59783 , \59784 , \59785 , \59786 , \59787 , \59788 , \59789 , \59790 , \59791 , \59792 ,
         \59793 , \59794 , \59795 , \59796 , \59797 , \59798 , \59799 , \59800 , \59801 , \59802 ,
         \59803 , \59804 , \59805 , \59806 , \59807 , \59808 , \59809 , \59810 , \59811 , \59812 ,
         \59813 , \59814 , \59815 , \59816 , \59817 , \59818 , \59819 , \59820 , \59821 , \59822 ,
         \59823 , \59824 , \59825 , \59826 , \59827 , \59828 , \59829 , \59830 , \59831 , \59832 ,
         \59833 , \59834 , \59835 , \59836 , \59837 , \59838 , \59839 , \59840 , \59841 , \59842 ,
         \59843 , \59844 , \59845 , \59846 , \59847 , \59848 , \59849 , \59850 , \59851 , \59852 ,
         \59853 , \59854 , \59855 , \59856 , \59857 , \59858 , \59859 , \59860 , \59861 , \59862 ,
         \59863 , \59864 , \59865 , \59866 , \59867 , \59868 , \59869 , \59870 , \59871 , \59872 ,
         \59873 , \59874 , \59875 , \59876 , \59877 , \59878 , \59879 , \59880 , \59881 , \59882 ,
         \59883 , \59884 , \59885 , \59886 , \59887 , \59888 , \59889 , \59890 , \59891 , \59892 ,
         \59893 , \59894 , \59895 , \59896 , \59897 , \59898 , \59899 , \59900 , \59901 , \59902 ,
         \59903 , \59904 , \59905 , \59906 , \59907 , \59908 , \59909 , \59910 , \59911 , \59912 ,
         \59913 , \59914 , \59915 , \59916 , \59917 , \59918 , \59919 , \59920 , \59921 , \59922 ,
         \59923 , \59924 , \59925 , \59926 , \59927 , \59928 , \59929 , \59930 , \59931 , \59932 ,
         \59933 , \59934 , \59935 , \59936 , \59937 , \59938 , \59939 , \59940 , \59941 , \59942 ,
         \59943 , \59944 , \59945 , \59946 , \59947 , \59948 , \59949 , \59950 , \59951 , \59952 ,
         \59953 , \59954 , \59955 , \59956 , \59957 , \59958 , \59959 , \59960 , \59961 , \59962 ,
         \59963 , \59964 , \59965 , \59966 , \59967 , \59968 , \59969 , \59970 , \59971 , \59972 ,
         \59973 , \59974 , \59975 , \59976 , \59977 , \59978 , \59979 , \59980 , \59981 , \59982 ,
         \59983 , \59984 , \59985 , \59986 , \59987 , \59988 , \59989 , \59990 , \59991 , \59992 ,
         \59993 , \59994 , \59995 , \59996 , \59997 , \59998 , \59999 , \60000 , \60001 , \60002 ,
         \60003 , \60004 , \60005 , \60006 , \60007 , \60008 , \60009 , \60010 , \60011 , \60012 ,
         \60013 , \60014 , \60015 , \60016 , \60017 , \60018 , \60019 , \60020 , \60021 , \60022 ,
         \60023 , \60024 , \60025 , \60026 , \60027 , \60028 , \60029 , \60030 , \60031 , \60032 ,
         \60033 , \60034 , \60035 , \60036 , \60037 , \60038 , \60039 , \60040 , \60041 , \60042 ,
         \60043 , \60044 , \60045 , \60046 , \60047 , \60048 , \60049 , \60050 , \60051 , \60052 ,
         \60053 , \60054 , \60055 , \60056 , \60057 , \60058 , \60059 , \60060 , \60061 , \60062 ,
         \60063 , \60064 , \60065 , \60066 , \60067 , \60068 , \60069 , \60070 , \60071 , \60072 ,
         \60073 , \60074 , \60075 , \60076 , \60077 , \60078 , \60079 , \60080 , \60081 , \60082 ,
         \60083 , \60084 , \60085 , \60086 , \60087 , \60088 , \60089 , \60090 , \60091 , \60092 ,
         \60093 , \60094 , \60095 , \60096 , \60097 , \60098 , \60099 , \60100 , \60101 , \60102 ,
         \60103 , \60104 , \60105 , \60106 , \60107 , \60108 , \60109 , \60110 , \60111 , \60112 ,
         \60113 , \60114 , \60115 , \60116 , \60117 , \60118 , \60119 , \60120 , \60121 , \60122 ,
         \60123 , \60124 , \60125 , \60126 , \60127 , \60128 , \60129 , \60130 , \60131 , \60132 ,
         \60133 , \60134 , \60135 , \60136 , \60137 , \60138 , \60139 , \60140 , \60141 , \60142 ,
         \60143 , \60144 , \60145 , \60146 , \60147 , \60148 , \60149 , \60150 , \60151 , \60152 ,
         \60153 , \60154 , \60155 , \60156 , \60157 , \60158 , \60159 , \60160 , \60161 , \60162 ,
         \60163 , \60164 , \60165 , \60166 , \60167 , \60168 , \60169 , \60170 , \60171 , \60172 ,
         \60173 , \60174 , \60175 , \60176 , \60177 , \60178 , \60179 , \60180 , \60181 , \60182 ,
         \60183 , \60184 , \60185 , \60186 , \60187 , \60188 , \60189 , \60190 , \60191 , \60192 ,
         \60193 , \60194 , \60195 , \60196 , \60197 , \60198 , \60199 , \60200 , \60201 , \60202 ,
         \60203 , \60204 , \60205 , \60206 , \60207 , \60208 , \60209 , \60210 , \60211 , \60212 ,
         \60213 , \60214 , \60215 , \60216 , \60217 , \60218 , \60219 , \60220 , \60221 , \60222 ,
         \60223 , \60224 , \60225 , \60226 , \60227 , \60228 , \60229 , \60230 , \60231 , \60232 ,
         \60233 , \60234 , \60235 , \60236 , \60237 , \60238 , \60239 , \60240 , \60241 , \60242 ,
         \60243 , \60244 , \60245 , \60246 , \60247 , \60248 , \60249 , \60250 , \60251 , \60252 ,
         \60253 , \60254 , \60255 , \60256 , \60257 , \60258 , \60259 , \60260 , \60261 , \60262 ,
         \60263 , \60264 , \60265 , \60266 , \60267 , \60268 , \60269 , \60270 , \60271 , \60272 ,
         \60273 , \60274 , \60275 , \60276 , \60277 , \60278 , \60279 , \60280 , \60281 , \60282 ,
         \60283 , \60284 , \60285 , \60286 , \60287 , \60288 , \60289 , \60290 , \60291 , \60292 ,
         \60293 , \60294 , \60295 , \60296 , \60297 , \60298 , \60299 , \60300 , \60301 , \60302 ,
         \60303 , \60304 , \60305 , \60306 , \60307 , \60308 , \60309 , \60310 , \60311 , \60312 ,
         \60313 , \60314 , \60315 , \60316 , \60317 , \60318 , \60319 , \60320 , \60321 , \60322 ,
         \60323 , \60324 , \60325 , \60326 , \60327 , \60328 , \60329 , \60330 , \60331 , \60332 ,
         \60333 , \60334 , \60335 , \60336 , \60337 , \60338 , \60339 , \60340 , \60341 , \60342 ,
         \60343 , \60344 , \60345 , \60346 , \60347 , \60348 , \60349 , \60350 , \60351 , \60352 ,
         \60353 , \60354 , \60355 , \60356 , \60357 , \60358 , \60359 , \60360 , \60361 , \60362 ,
         \60363 , \60364 , \60365 , \60366 , \60367 , \60368 , \60369 , \60370 , \60371 , \60372 ,
         \60373 , \60374 , \60375 , \60376 , \60377 , \60378 , \60379 , \60380 , \60381 , \60382 ,
         \60383 , \60384 , \60385 , \60386 , \60387 , \60388 , \60389 , \60390 , \60391 , \60392 ,
         \60393 , \60394 , \60395 , \60396 , \60397 , \60398 , \60399 , \60400 , \60401 , \60402 ,
         \60403 , \60404 , \60405 , \60406 , \60407 , \60408 , \60409 , \60410 , \60411 , \60412 ,
         \60413 , \60414 , \60415 , \60416 , \60417 , \60418 , \60419 , \60420 , \60421 , \60422 ,
         \60423 , \60424 , \60425 , \60426 , \60427 , \60428 , \60429 , \60430 , \60431 , \60432 ,
         \60433 , \60434 , \60435 , \60436 , \60437 , \60438 , \60439 , \60440 , \60441 , \60442 ,
         \60443 , \60444 , \60445 , \60446 , \60447 , \60448 , \60449 , \60450 , \60451 , \60452 ,
         \60453 , \60454 , \60455 , \60456 , \60457 , \60458 , \60459 , \60460 , \60461 , \60462 ,
         \60463 , \60464 , \60465 , \60466 , \60467 , \60468 , \60469 , \60470 , \60471 , \60472 ,
         \60473 , \60474 , \60475 , \60476 , \60477 , \60478 , \60479 , \60480 , \60481 , \60482 ,
         \60483 , \60484 , \60485 , \60486 , \60487 , \60488 , \60489 , \60490 , \60491 , \60492 ,
         \60493 , \60494 , \60495 , \60496 , \60497 , \60498 , \60499 , \60500 , \60501 , \60502 ,
         \60503 , \60504 , \60505 , \60506 , \60507 , \60508 , \60509 , \60510 , \60511 , \60512 ,
         \60513 , \60514 , \60515 , \60516 , \60517 , \60518 , \60519 , \60520 , \60521 , \60522 ,
         \60523 , \60524 , \60525 , \60526 , \60527 , \60528 , \60529 , \60530 , \60531 , \60532 ,
         \60533 , \60534 , \60535 , \60536 , \60537 , \60538 , \60539 , \60540 , \60541 , \60542 ,
         \60543 , \60544 , \60545 , \60546 , \60547 , \60548 , \60549 , \60550 , \60551 , \60552 ,
         \60553 , \60554 , \60555 , \60556 , \60557 , \60558 , \60559 , \60560 , \60561 , \60562 ,
         \60563 , \60564 , \60565 , \60566 , \60567 , \60568 , \60569 , \60570 , \60571 , \60572 ,
         \60573 , \60574 , \60575 , \60576 , \60577 , \60578 , \60579 , \60580 , \60581 , \60582 ,
         \60583 , \60584 , \60585 , \60586 , \60587 , \60588 , \60589 , \60590 , \60591 , \60592 ,
         \60593 , \60594 , \60595 , \60596 , \60597 , \60598 , \60599 , \60600 , \60601 , \60602 ,
         \60603 , \60604 , \60605 , \60606 , \60607 , \60608 , \60609 , \60610 , \60611 , \60612 ,
         \60613 , \60614 , \60615 , \60616 , \60617 , \60618 , \60619 , \60620 , \60621 , \60622 ,
         \60623 , \60624 , \60625 , \60626 , \60627 , \60628 , \60629 , \60630 , \60631 , \60632 ,
         \60633 , \60634 , \60635 , \60636 , \60637 , \60638 , \60639 , \60640 , \60641 , \60642 ,
         \60643 , \60644 , \60645 , \60646 , \60647 , \60648 , \60649 , \60650 , \60651 , \60652 ,
         \60653 , \60654 , \60655 , \60656 , \60657 , \60658 , \60659 , \60660 , \60661 , \60662 ,
         \60663 , \60664 , \60665 , \60666 , \60667 , \60668 , \60669 , \60670 , \60671 , \60672 ,
         \60673 , \60674 , \60675 , \60676 , \60677 , \60678 , \60679 , \60680 , \60681 , \60682 ,
         \60683 , \60684 , \60685 , \60686 , \60687 , \60688 , \60689 , \60690 , \60691 , \60692 ,
         \60693 , \60694 , \60695 , \60696 , \60697 , \60698 , \60699 , \60700 , \60701 , \60702 ,
         \60703 , \60704 , \60705 , \60706 , \60707 , \60708 , \60709 , \60710 , \60711 , \60712 ,
         \60713 , \60714 , \60715 , \60716 , \60717 , \60718 , \60719 , \60720 , \60721 , \60722 ,
         \60723 , \60724 , \60725 , \60726 , \60727 , \60728 , \60729 , \60730 , \60731 , \60732 ,
         \60733 , \60734 , \60735 , \60736 , \60737 , \60738 , \60739 , \60740 , \60741 , \60742 ,
         \60743 , \60744 , \60745 , \60746 , \60747 , \60748 , \60749 , \60750 , \60751 , \60752 ,
         \60753 , \60754 , \60755 , \60756 , \60757 , \60758 , \60759 , \60760 , \60761 , \60762 ,
         \60763 , \60764 , \60765 , \60766 , \60767 , \60768 , \60769 , \60770 , \60771 , \60772 ,
         \60773 , \60774 , \60775 , \60776 , \60777 , \60778 , \60779 , \60780 , \60781 , \60782 ,
         \60783 , \60784 , \60785 , \60786 , \60787 , \60788 , \60789 , \60790 , \60791 , \60792 ,
         \60793 , \60794 , \60795 , \60796 , \60797 , \60798 , \60799 , \60800 , \60801 , \60802 ,
         \60803 , \60804 , \60805 , \60806 , \60807 , \60808 , \60809 , \60810 , \60811 , \60812 ,
         \60813 , \60814 , \60815 , \60816 , \60817 , \60818 , \60819 , \60820 , \60821 , \60822 ,
         \60823 , \60824 , \60825 , \60826 , \60827 , \60828 , \60829 , \60830 , \60831 , \60832 ,
         \60833 , \60834 , \60835 , \60836 , \60837 , \60838 , \60839 , \60840 , \60841 , \60842 ,
         \60843 , \60844 , \60845 , \60846 , \60847 , \60848 , \60849 , \60850 , \60851 , \60852 ,
         \60853 , \60854 , \60855 , \60856 , \60857 , \60858 , \60859 , \60860 , \60861 , \60862 ,
         \60863 , \60864 , \60865 , \60866 , \60867 , \60868 , \60869 , \60870 , \60871 , \60872 ,
         \60873 , \60874 , \60875 , \60876 , \60877 , \60878 , \60879 , \60880 , \60881 , \60882 ,
         \60883 , \60884 , \60885 , \60886 , \60887 , \60888 , \60889 , \60890 , \60891 , \60892 ,
         \60893 , \60894 , \60895 , \60896 , \60897 , \60898 , \60899 , \60900 , \60901 , \60902 ,
         \60903 , \60904 , \60905 , \60906 , \60907 , \60908 , \60909 , \60910 , \60911 , \60912 ,
         \60913 , \60914 , \60915 , \60916 , \60917 , \60918 , \60919 , \60920 , \60921 , \60922 ,
         \60923 , \60924 , \60925 , \60926 , \60927 , \60928 , \60929 , \60930 , \60931 , \60932 ,
         \60933 , \60934 , \60935 , \60936 , \60937 , \60938 , \60939 , \60940 , \60941 , \60942 ,
         \60943 , \60944 , \60945 , \60946 , \60947 , \60948 , \60949 , \60950 , \60951 , \60952 ,
         \60953 , \60954 , \60955 , \60956 , \60957 , \60958 , \60959 , \60960 , \60961 , \60962 ,
         \60963 , \60964 , \60965 , \60966 , \60967 , \60968 , \60969 , \60970 , \60971 , \60972 ,
         \60973 , \60974 , \60975 , \60976 , \60977 , \60978 , \60979 , \60980 , \60981 , \60982 ,
         \60983 , \60984 , \60985 , \60986 , \60987 , \60988 , \60989 , \60990 , \60991 , \60992 ,
         \60993 , \60994 , \60995 , \60996 , \60997 , \60998 , \60999 , \61000 , \61001 , \61002 ,
         \61003 , \61004 , \61005 , \61006 , \61007 , \61008 , \61009 , \61010 , \61011 , \61012 ,
         \61013 , \61014 , \61015 , \61016 , \61017 , \61018 , \61019 , \61020 , \61021 , \61022 ,
         \61023 , \61024 , \61025 , \61026 , \61027 , \61028 , \61029 , \61030 , \61031 , \61032 ,
         \61033 , \61034 , \61035 , \61036 , \61037 , \61038 , \61039 , \61040 , \61041 , \61042 ,
         \61043 , \61044 , \61045 , \61046 , \61047 , \61048 , \61049 , \61050 , \61051 , \61052 ,
         \61053 , \61054 , \61055 , \61056 , \61057 , \61058 , \61059 , \61060 , \61061 , \61062 ,
         \61063 , \61064 , \61065 , \61066 , \61067 , \61068 , \61069 , \61070 , \61071 , \61072 ,
         \61073 , \61074 , \61075 , \61076 , \61077 , \61078 , \61079 , \61080 , \61081 , \61082 ,
         \61083 , \61084 , \61085 , \61086 , \61087 , \61088 , \61089 , \61090 , \61091 , \61092 ,
         \61093 , \61094 , \61095 , \61096 , \61097 , \61098 , \61099 , \61100 , \61101 , \61102 ,
         \61103 , \61104 , \61105 , \61106 , \61107 , \61108 , \61109 , \61110 , \61111 , \61112 ,
         \61113 , \61114 , \61115 , \61116 , \61117 , \61118 , \61119 , \61120 , \61121 , \61122 ,
         \61123 , \61124 , \61125 , \61126 , \61127 , \61128 , \61129 , \61130 , \61131 , \61132 ,
         \61133 , \61134 , \61135 , \61136 , \61137 , \61138 , \61139 , \61140 , \61141 , \61142 ,
         \61143 , \61144 , \61145 , \61146 , \61147 , \61148 , \61149 , \61150 , \61151 , \61152 ,
         \61153 , \61154 , \61155 , \61156 , \61157 , \61158 , \61159 , \61160 , \61161 , \61162 ,
         \61163 , \61164 , \61165 , \61166 , \61167 , \61168 , \61169 , \61170 , \61171 , \61172 ,
         \61173 , \61174 , \61175 , \61176 , \61177 , \61178 , \61179 , \61180 , \61181 , \61182 ,
         \61183 , \61184 , \61185 , \61186 , \61187 , \61188 , \61189 , \61190 , \61191 , \61192 ,
         \61193 , \61194 , \61195 , \61196 , \61197 , \61198 , \61199 , \61200 , \61201 , \61202 ,
         \61203 , \61204 , \61205 , \61206 , \61207 , \61208 , \61209 , \61210 , \61211 , \61212 ,
         \61213 , \61214 , \61215 , \61216 , \61217 , \61218 , \61219 , \61220 , \61221 , \61222 ,
         \61223 , \61224 , \61225 , \61226 , \61227 , \61228 , \61229 , \61230 , \61231 , \61232 ,
         \61233 , \61234 , \61235 , \61236 , \61237 , \61238 , \61239 , \61240 , \61241 , \61242 ,
         \61243 , \61244 , \61245 , \61246 , \61247 , \61248 , \61249 , \61250 , \61251 , \61252 ,
         \61253 , \61254 , \61255 , \61256 , \61257 , \61258 , \61259 , \61260 , \61261 , \61262 ,
         \61263 , \61264 , \61265 , \61266 , \61267 , \61268 , \61269 , \61270 , \61271 , \61272 ,
         \61273 , \61274 , \61275 , \61276 , \61277 , \61278 , \61279 , \61280 , \61281 , \61282 ,
         \61283 , \61284 , \61285 , \61286 , \61287 , \61288 , \61289 , \61290 , \61291 , \61292 ,
         \61293 , \61294 , \61295 , \61296 , \61297 , \61298 , \61299 , \61300 , \61301 , \61302 ,
         \61303 , \61304 , \61305 , \61306 , \61307 , \61308 , \61309 , \61310 , \61311 , \61312 ,
         \61313 , \61314 , \61315 , \61316 , \61317 , \61318 , \61319 , \61320 , \61321 , \61322 ,
         \61323 , \61324 , \61325 , \61326 , \61327 , \61328 , \61329 , \61330 , \61331 , \61332 ,
         \61333 , \61334 , \61335 , \61336 , \61337 , \61338 , \61339 , \61340 , \61341 , \61342 ,
         \61343 , \61344 , \61345 , \61346 , \61347 , \61348 , \61349 , \61350 , \61351 , \61352 ,
         \61353 , \61354 , \61355 , \61356 , \61357 , \61358 , \61359 , \61360 , \61361 , \61362 ,
         \61363 , \61364 , \61365 , \61366 , \61367 , \61368 , \61369 , \61370 , \61371 , \61372 ,
         \61373 , \61374 , \61375 , \61376 , \61377 , \61378 , \61379 , \61380 , \61381 , \61382 ,
         \61383 , \61384 , \61385 , \61386 , \61387 , \61388 , \61389 , \61390 , \61391 , \61392 ,
         \61393 , \61394 , \61395 , \61396 , \61397 , \61398 , \61399 , \61400 , \61401 , \61402 ,
         \61403 , \61404 , \61405 , \61406 , \61407 , \61408 , \61409 , \61410 , \61411 , \61412 ,
         \61413 , \61414 , \61415 , \61416 , \61417 , \61418 , \61419 , \61420 , \61421 , \61422 ,
         \61423 , \61424 , \61425 , \61426 , \61427 , \61428 , \61429 , \61430 , \61431 , \61432 ,
         \61433 , \61434 , \61435 , \61436 , \61437 , \61438 , \61439 , \61440 , \61441 , \61442 ,
         \61443 , \61444 , \61445 , \61446 , \61447 , \61448 , \61449 , \61450 , \61451 , \61452 ,
         \61453 , \61454 , \61455 , \61456 , \61457 , \61458 , \61459 , \61460 , \61461 , \61462 ,
         \61463 , \61464 , \61465 , \61466 , \61467 , \61468 , \61469 , \61470 , \61471 , \61472 ,
         \61473 , \61474 , \61475 , \61476 , \61477 , \61478 , \61479 , \61480 , \61481 , \61482 ,
         \61483 , \61484 , \61485 , \61486 , \61487 , \61488 , \61489 , \61490 , \61491 , \61492 ,
         \61493 , \61494 , \61495 , \61496 , \61497 , \61498 , \61499 , \61500 , \61501 , \61502 ,
         \61503 , \61504 , \61505 , \61506 , \61507 , \61508 , \61509 , \61510 , \61511 , \61512 ,
         \61513 , \61514 , \61515 , \61516 , \61517 , \61518 , \61519 , \61520 , \61521 , \61522 ,
         \61523 , \61524 , \61525 , \61526 , \61527 , \61528 , \61529 , \61530 , \61531 , \61532 ,
         \61533 , \61534 , \61535 , \61536 , \61537 , \61538 , \61539 , \61540 , \61541 , \61542 ,
         \61543 , \61544 , \61545 , \61546 , \61547 , \61548 , \61549 , \61550 , \61551 , \61552 ,
         \61553 , \61554 , \61555 , \61556 , \61557 , \61558 , \61559 , \61560 , \61561 , \61562 ,
         \61563 , \61564 , \61565 , \61566 , \61567 , \61568 , \61569 , \61570 , \61571 , \61572 ,
         \61573 , \61574 , \61575 , \61576 , \61577 , \61578 , \61579 , \61580 , \61581 , \61582 ,
         \61583 , \61584 , \61585 , \61586 , \61587 , \61588 , \61589 , \61590 , \61591 , \61592 ,
         \61593 , \61594 , \61595 , \61596 , \61597 , \61598 , \61599 , \61600 , \61601 , \61602 ,
         \61603 , \61604 , \61605 , \61606 , \61607 , \61608 , \61609 , \61610 , \61611 , \61612 ,
         \61613 , \61614 , \61615 , \61616 , \61617 , \61618 , \61619 , \61620 , \61621 , \61622 ,
         \61623 , \61624 , \61625 , \61626 , \61627 , \61628 , \61629 , \61630 , \61631 , \61632 ,
         \61633 , \61634 , \61635 , \61636 , \61637 , \61638 , \61639 , \61640 , \61641 , \61642 ,
         \61643 , \61644 , \61645 , \61646 , \61647 , \61648 , \61649 , \61650 , \61651 , \61652 ,
         \61653 , \61654 , \61655 , \61656 , \61657 , \61658 , \61659 , \61660 , \61661 , \61662 ,
         \61663 , \61664 , \61665 , \61666 , \61667 , \61668 , \61669 , \61670 , \61671 , \61672 ,
         \61673 , \61674 , \61675 , \61676 , \61677 , \61678 , \61679 , \61680 , \61681 , \61682 ,
         \61683 , \61684 , \61685 , \61686 , \61687 , \61688 , \61689 , \61690 , \61691 , \61692 ,
         \61693 , \61694 , \61695 , \61696 , \61697 , \61698 , \61699 , \61700 , \61701 , \61702 ,
         \61703 , \61704 , \61705 , \61706 , \61707 , \61708 , \61709 , \61710 , \61711 , \61712 ,
         \61713 , \61714 , \61715 , \61716 , \61717 , \61718 , \61719 , \61720 , \61721 , \61722 ,
         \61723 , \61724 , \61725 , \61726 , \61727 , \61728 , \61729 , \61730 , \61731 , \61732 ,
         \61733 , \61734 , \61735 , \61736 , \61737 , \61738 , \61739 , \61740 , \61741 , \61742 ,
         \61743 , \61744 , \61745 , \61746 , \61747 , \61748 , \61749 , \61750 , \61751 , \61752 ,
         \61753 , \61754 , \61755 , \61756 , \61757 , \61758 , \61759 , \61760 , \61761 , \61762 ,
         \61763 , \61764 , \61765 , \61766 , \61767 , \61768 , \61769 , \61770 , \61771 , \61772 ,
         \61773 , \61774 , \61775 , \61776 , \61777 , \61778 , \61779 , \61780 , \61781 , \61782 ,
         \61783 , \61784 , \61785 , \61786 , \61787 , \61788 , \61789 , \61790 , \61791 , \61792 ,
         \61793 , \61794 , \61795 , \61796 , \61797 , \61798 , \61799 , \61800 , \61801 , \61802 ,
         \61803 , \61804 , \61805 , \61806 , \61807 , \61808 , \61809 , \61810 , \61811 , \61812 ,
         \61813 , \61814 , \61815 , \61816 , \61817 , \61818 , \61819 , \61820 , \61821 , \61822 ,
         \61823 , \61824 , \61825 , \61826 , \61827 , \61828 , \61829 , \61830 , \61831 , \61832 ,
         \61833 , \61834 , \61835 , \61836 , \61837 , \61838 , \61839 , \61840 , \61841 , \61842 ,
         \61843 , \61844 , \61845 , \61846 , \61847 , \61848 , \61849 , \61850 , \61851 , \61852 ,
         \61853 , \61854 , \61855 , \61856 , \61857 , \61858 , \61859 , \61860 , \61861 , \61862 ,
         \61863 , \61864 , \61865 , \61866 , \61867 , \61868 , \61869 , \61870 , \61871 , \61872 ,
         \61873 , \61874 , \61875 , \61876 , \61877 , \61878 , \61879 , \61880 , \61881 , \61882 ,
         \61883 , \61884 , \61885 , \61886 , \61887 , \61888 , \61889 , \61890 , \61891 , \61892 ,
         \61893 , \61894 , \61895 , \61896 , \61897 , \61898 , \61899 , \61900 , \61901 , \61902 ,
         \61903 , \61904 , \61905 , \61906 , \61907 , \61908 , \61909 , \61910 , \61911 , \61912 ,
         \61913 , \61914 , \61915 , \61916 , \61917 , \61918 , \61919 , \61920 , \61921 , \61922 ,
         \61923 , \61924 , \61925 , \61926 , \61927 , \61928 , \61929 , \61930 , \61931 , \61932 ,
         \61933 , \61934 , \61935 , \61936 , \61937 , \61938 , \61939 , \61940 , \61941 , \61942 ,
         \61943 , \61944 , \61945 , \61946 , \61947 , \61948 , \61949 , \61950 , \61951 , \61952 ,
         \61953 , \61954 , \61955 , \61956 , \61957 , \61958 , \61959 , \61960 , \61961 , \61962 ,
         \61963 , \61964 , \61965 , \61966 , \61967 , \61968 , \61969 , \61970 , \61971 , \61972 ,
         \61973 , \61974 , \61975 , \61976 , \61977 , \61978 , \61979 , \61980 , \61981 , \61982 ,
         \61983 , \61984 , \61985 , \61986 , \61987 , \61988 , \61989 , \61990 , \61991 , \61992 ,
         \61993 , \61994 , \61995 , \61996 , \61997 , \61998 , \61999 , \62000 , \62001 , \62002 ,
         \62003 , \62004 , \62005 , \62006 , \62007 , \62008 , \62009 , \62010 , \62011 , \62012 ,
         \62013 , \62014 , \62015 , \62016 , \62017 , \62018 , \62019 , \62020 , \62021 , \62022 ,
         \62023 , \62024 , \62025 , \62026 , \62027 , \62028 , \62029 , \62030 , \62031 , \62032 ,
         \62033 , \62034 , \62035 , \62036 , \62037 , \62038 , \62039 , \62040 , \62041 , \62042 ,
         \62043 , \62044 , \62045 , \62046 , \62047 , \62048 , \62049 , \62050 , \62051 , \62052 ,
         \62053 , \62054 , \62055 , \62056 , \62057 , \62058 , \62059 , \62060 , \62061 , \62062 ,
         \62063 , \62064 , \62065 , \62066 , \62067 , \62068 , \62069 , \62070 , \62071 , \62072 ,
         \62073 , \62074 , \62075 , \62076 , \62077 , \62078 , \62079 , \62080 , \62081 , \62082 ,
         \62083 , \62084 , \62085 , \62086 , \62087 , \62088 , \62089 , \62090 , \62091 , \62092 ,
         \62093 , \62094 , \62095 , \62096 , \62097 , \62098 , \62099 , \62100 , \62101 , \62102 ,
         \62103 , \62104 , \62105 , \62106 , \62107 , \62108 , \62109 , \62110 , \62111 , \62112 ,
         \62113 , \62114 , \62115 , \62116 , \62117 , \62118 , \62119 , \62120 , \62121 , \62122 ,
         \62123 , \62124 , \62125 , \62126 , \62127 , \62128 , \62129 , \62130 , \62131 , \62132 ,
         \62133 , \62134 , \62135 , \62136 , \62137 , \62138 , \62139 , \62140 , \62141 , \62142 ,
         \62143 , \62144 , \62145 , \62146 , \62147 , \62148 , \62149 , \62150 , \62151 , \62152 ,
         \62153 , \62154 , \62155 , \62156 , \62157 , \62158 , \62159 , \62160 , \62161 , \62162 ,
         \62163 , \62164 , \62165 , \62166 , \62167 , \62168 , \62169 , \62170 , \62171 , \62172 ,
         \62173 , \62174 , \62175 , \62176 , \62177 , \62178 , \62179 , \62180 , \62181 , \62182 ,
         \62183 , \62184 , \62185 , \62186 , \62187 , \62188 , \62189 , \62190 , \62191 , \62192 ,
         \62193 , \62194 , \62195 , \62196 , \62197 , \62198 , \62199 , \62200 , \62201 , \62202 ,
         \62203 , \62204 , \62205 , \62206 , \62207 , \62208 , \62209 , \62210 , \62211 , \62212 ,
         \62213 , \62214 , \62215 , \62216 , \62217 , \62218 , \62219 , \62220 , \62221 , \62222 ,
         \62223 , \62224 , \62225 , \62226 , \62227 , \62228 , \62229 , \62230 , \62231 , \62232 ,
         \62233 , \62234 , \62235 , \62236 , \62237 , \62238 , \62239 , \62240 , \62241 , \62242 ,
         \62243 , \62244 , \62245 , \62246 , \62247 , \62248 , \62249 , \62250 , \62251 , \62252 ,
         \62253 , \62254 , \62255 , \62256 , \62257 , \62258 , \62259 , \62260 , \62261 , \62262 ,
         \62263 , \62264 , \62265 , \62266 , \62267 , \62268 , \62269 , \62270 , \62271 , \62272 ,
         \62273 , \62274 , \62275 , \62276 , \62277 , \62278 , \62279 , \62280 , \62281 , \62282 ,
         \62283 , \62284 , \62285 , \62286 , \62287 , \62288 , \62289 , \62290 , \62291 , \62292 ,
         \62293 , \62294 , \62295 , \62296 , \62297 , \62298 , \62299 , \62300 , \62301 , \62302 ,
         \62303 , \62304 , \62305 , \62306 , \62307 , \62308 , \62309 , \62310 , \62311 , \62312 ,
         \62313 , \62314 , \62315 , \62316 , \62317 , \62318 , \62319 , \62320 , \62321 , \62322 ,
         \62323 , \62324 , \62325 , \62326 , \62327 , \62328 , \62329 , \62330 , \62331 , \62332 ,
         \62333 , \62334 , \62335 , \62336 , \62337 , \62338 , \62339 , \62340 , \62341 , \62342 ,
         \62343 , \62344 , \62345 , \62346 , \62347 , \62348 , \62349 , \62350 , \62351 , \62352 ,
         \62353 , \62354 , \62355 , \62356 , \62357 , \62358 , \62359 , \62360 , \62361 , \62362 ,
         \62363 , \62364 , \62365 , \62366 , \62367 , \62368 , \62369 , \62370 , \62371 , \62372 ,
         \62373 , \62374 , \62375 , \62376 , \62377 , \62378 , \62379 , \62380 , \62381 , \62382 ,
         \62383 , \62384 , \62385 , \62386 , \62387 , \62388 , \62389 , \62390 , \62391 , \62392 ,
         \62393 , \62394 , \62395 , \62396 , \62397 , \62398 , \62399 , \62400 , \62401 , \62402 ,
         \62403 , \62404 , \62405 , \62406 , \62407 , \62408 , \62409 , \62410 , \62411 , \62412 ,
         \62413 , \62414 , \62415 , \62416 , \62417 , \62418 , \62419 , \62420 , \62421 , \62422 ,
         \62423 , \62424 , \62425 , \62426 , \62427 , \62428 , \62429 , \62430 , \62431 , \62432 ,
         \62433 , \62434 , \62435 , \62436 , \62437 , \62438 , \62439 , \62440 , \62441 , \62442 ,
         \62443 , \62444 , \62445 , \62446 , \62447 , \62448 , \62449 , \62450 , \62451 , \62452 ,
         \62453 , \62454 , \62455 , \62456 , \62457 , \62458 , \62459 , \62460 , \62461 , \62462 ,
         \62463 , \62464 , \62465 , \62466 , \62467 , \62468 , \62469 , \62470 , \62471 , \62472 ,
         \62473 , \62474 , \62475 , \62476 , \62477 , \62478 , \62479 , \62480 , \62481 , \62482 ,
         \62483 , \62484 , \62485 , \62486 , \62487 , \62488 , \62489 , \62490 , \62491 , \62492 ,
         \62493 , \62494 , \62495 , \62496 , \62497 , \62498 , \62499 , \62500 , \62501 , \62502 ,
         \62503 , \62504 , \62505 , \62506 , \62507 , \62508 , \62509 , \62510 , \62511 , \62512 ,
         \62513 , \62514 , \62515 , \62516 , \62517 , \62518 , \62519 , \62520 , \62521 , \62522 ,
         \62523 , \62524 , \62525 , \62526 , \62527 , \62528 , \62529 , \62530 , \62531 , \62532 ,
         \62533 , \62534 , \62535 , \62536 , \62537 , \62538 , \62539 , \62540 , \62541 , \62542 ,
         \62543 , \62544 , \62545 , \62546 , \62547 , \62548 , \62549 , \62550 , \62551 , \62552 ,
         \62553 , \62554 , \62555 , \62556 , \62557 , \62558 , \62559 , \62560 , \62561 , \62562 ,
         \62563 , \62564 , \62565 , \62566 , \62567 , \62568 , \62569 , \62570 , \62571 , \62572 ,
         \62573 , \62574 , \62575 , \62576 , \62577 , \62578 , \62579 , \62580 , \62581 , \62582 ,
         \62583 , \62584 , \62585 , \62586 , \62587 , \62588 , \62589 , \62590 , \62591 , \62592 ,
         \62593 , \62594 , \62595 , \62596 , \62597 , \62598 , \62599 , \62600 , \62601 , \62602 ,
         \62603 , \62604 , \62605 , \62606 , \62607 , \62608 , \62609 , \62610 , \62611 , \62612 ,
         \62613 , \62614 , \62615 , \62616 , \62617 , \62618 , \62619 , \62620 , \62621 , \62622 ,
         \62623 , \62624 , \62625 , \62626 , \62627 , \62628 , \62629 , \62630 , \62631 , \62632 ,
         \62633 , \62634 , \62635 , \62636 , \62637 , \62638 , \62639 , \62640 , \62641 , \62642 ,
         \62643 , \62644 , \62645 , \62646 , \62647 , \62648 , \62649 , \62650 , \62651 , \62652 ,
         \62653 , \62654 , \62655 , \62656 , \62657 , \62658 , \62659 , \62660 , \62661 , \62662 ,
         \62663 , \62664 , \62665 , \62666 , \62667 , \62668 , \62669 , \62670 , \62671 , \62672 ,
         \62673 , \62674 , \62675 , \62676 , \62677 , \62678 , \62679 , \62680 , \62681 , \62682 ,
         \62683 , \62684 , \62685 , \62686 , \62687 , \62688 , \62689 , \62690 , \62691 , \62692 ,
         \62693 , \62694 , \62695 , \62696 , \62697 , \62698 , \62699 , \62700 , \62701 , \62702 ,
         \62703 , \62704 , \62705 , \62706 , \62707 , \62708 , \62709 , \62710 , \62711 , \62712 ,
         \62713 , \62714 , \62715 , \62716 , \62717 , \62718 , \62719 , \62720 , \62721 , \62722 ,
         \62723 , \62724 , \62725 , \62726 , \62727 , \62728 , \62729 , \62730 , \62731 , \62732 ,
         \62733 , \62734 , \62735 , \62736 , \62737 , \62738 , \62739 , \62740 , \62741 , \62742 ,
         \62743 , \62744 , \62745 , \62746 , \62747 , \62748 , \62749 , \62750 , \62751 , \62752 ,
         \62753 , \62754 , \62755 , \62756 , \62757 , \62758 , \62759 , \62760 , \62761 , \62762 ,
         \62763 , \62764 , \62765 , \62766 , \62767 , \62768 , \62769 , \62770 , \62771 , \62772 ,
         \62773 , \62774 , \62775 , \62776 , \62777 , \62778 , \62779 , \62780 , \62781 , \62782 ,
         \62783 , \62784 , \62785 , \62786 , \62787 , \62788 , \62789 , \62790 , \62791 , \62792 ,
         \62793 , \62794 , \62795 , \62796 , \62797 , \62798 , \62799 , \62800 , \62801 , \62802 ,
         \62803 , \62804 , \62805 , \62806 , \62807 , \62808 , \62809 , \62810 , \62811 , \62812 ,
         \62813 , \62814 , \62815 , \62816 , \62817 , \62818 , \62819 , \62820 , \62821 , \62822 ,
         \62823 , \62824 , \62825 , \62826 , \62827 , \62828 , \62829 , \62830 , \62831 , \62832 ,
         \62833 , \62834 , \62835 , \62836 , \62837 , \62838 , \62839 , \62840 , \62841 , \62842 ,
         \62843 , \62844 , \62845 , \62846 , \62847 , \62848 , \62849 , \62850 , \62851 , \62852 ,
         \62853 , \62854 , \62855 , \62856 , \62857 , \62858 , \62859 , \62860 , \62861 , \62862 ,
         \62863 , \62864 , \62865 , \62866 , \62867 , \62868 , \62869 , \62870 , \62871 , \62872 ,
         \62873 , \62874 , \62875 , \62876 , \62877 , \62878 , \62879 , \62880 , \62881 , \62882 ,
         \62883 , \62884 , \62885 , \62886 , \62887 , \62888 , \62889 , \62890 , \62891 , \62892 ,
         \62893 , \62894 , \62895 , \62896 , \62897 , \62898 , \62899 , \62900 , \62901 , \62902 ,
         \62903 , \62904 , \62905 , \62906 , \62907 , \62908 , \62909 , \62910 , \62911 , \62912 ,
         \62913 , \62914 , \62915 , \62916 , \62917 , \62918 , \62919 , \62920 , \62921 , \62922 ,
         \62923 , \62924 , \62925 , \62926 , \62927 , \62928 , \62929 , \62930 , \62931 , \62932 ,
         \62933 , \62934 , \62935 , \62936 , \62937 , \62938 , \62939 , \62940 , \62941 , \62942 ,
         \62943 , \62944 , \62945 , \62946 , \62947 , \62948 , \62949 , \62950 , \62951 , \62952 ,
         \62953 , \62954 , \62955 , \62956 , \62957 , \62958 , \62959 , \62960 , \62961 , \62962 ,
         \62963 , \62964 , \62965 , \62966 , \62967 , \62968 , \62969 , \62970 , \62971 , \62972 ,
         \62973 , \62974 , \62975 , \62976 , \62977 , \62978 , \62979 , \62980 , \62981 , \62982 ,
         \62983 , \62984 , \62985 , \62986 , \62987 , \62988 , \62989 , \62990 , \62991 , \62992 ,
         \62993 , \62994 , \62995 , \62996 , \62997 , \62998 , \62999 , \63000 , \63001 , \63002 ,
         \63003 , \63004 , \63005 , \63006 , \63007 , \63008 , \63009 , \63010 , \63011 , \63012 ,
         \63013 , \63014 , \63015 , \63016 , \63017 , \63018 , \63019 , \63020 , \63021 , \63022 ,
         \63023 , \63024 , \63025 , \63026 , \63027 , \63028 , \63029 , \63030 , \63031 , \63032 ,
         \63033 , \63034 , \63035 , \63036 , \63037 , \63038 , \63039 , \63040 , \63041 , \63042 ,
         \63043 , \63044 , \63045 , \63046 , \63047 , \63048 , \63049 , \63050 , \63051 , \63052 ,
         \63053 , \63054 , \63055 , \63056 , \63057 , \63058 , \63059 , \63060 , \63061 , \63062 ,
         \63063 , \63064 , \63065 , \63066 , \63067 , \63068 , \63069 , \63070 , \63071 , \63072 ,
         \63073 , \63074 , \63075 , \63076 , \63077 , \63078 , \63079 , \63080 , \63081 , \63082 ,
         \63083 , \63084 , \63085 , \63086 , \63087 , \63088 , \63089 , \63090 , \63091 , \63092 ,
         \63093 , \63094 , \63095 , \63096 , \63097 , \63098 , \63099 , \63100 , \63101 , \63102 ,
         \63103 , \63104 , \63105 , \63106 , \63107 , \63108 , \63109 , \63110 , \63111 , \63112 ,
         \63113 , \63114 , \63115 , \63116 , \63117 , \63118 , \63119 , \63120 , \63121 , \63122 ,
         \63123 , \63124 , \63125 , \63126 , \63127 , \63128 , \63129 , \63130 , \63131 , \63132 ,
         \63133 , \63134 , \63135 , \63136 , \63137 , \63138 , \63139 , \63140 , \63141 , \63142 ,
         \63143 , \63144 , \63145 , \63146 , \63147 , \63148 , \63149 , \63150 , \63151 , \63152 ,
         \63153 , \63154 , \63155 , \63156 , \63157 , \63158 , \63159 , \63160 , \63161 , \63162 ,
         \63163 , \63164 , \63165 , \63166 , \63167 , \63168 , \63169 , \63170 , \63171 , \63172 ,
         \63173 , \63174 , \63175 , \63176 , \63177 , \63178 , \63179 , \63180 , \63181 , \63182 ,
         \63183 , \63184 , \63185 , \63186 , \63187 , \63188 , \63189 , \63190 , \63191 , \63192 ,
         \63193 , \63194 , \63195 , \63196 , \63197 , \63198 , \63199 , \63200 , \63201 , \63202 ,
         \63203 , \63204 , \63205 , \63206 , \63207 , \63208 , \63209 , \63210 , \63211 , \63212 ,
         \63213 , \63214 , \63215 , \63216 , \63217 , \63218 , \63219 , \63220 , \63221 , \63222 ,
         \63223 , \63224 , \63225 , \63226 , \63227 , \63228 , \63229 , \63230 , \63231 , \63232 ,
         \63233 , \63234 , \63235 , \63236 , \63237 , \63238 , \63239 , \63240 , \63241 , \63242 ,
         \63243 , \63244 , \63245 , \63246 , \63247 , \63248 , \63249 , \63250 , \63251 , \63252 ,
         \63253 , \63254 , \63255 , \63256 , \63257 , \63258 , \63259 , \63260 , \63261 , \63262 ,
         \63263 , \63264 , \63265 , \63266 , \63267 , \63268 , \63269 , \63270 , \63271 , \63272 ,
         \63273 , \63274 , \63275 , \63276 , \63277 , \63278 , \63279 , \63280 , \63281 , \63282 ,
         \63283 , \63284 , \63285 , \63286 , \63287 , \63288 , \63289 , \63290 , \63291 , \63292 ,
         \63293 , \63294 , \63295 , \63296 , \63297 , \63298 , \63299 , \63300 , \63301 , \63302 ,
         \63303 , \63304 , \63305 , \63306 , \63307 , \63308 , \63309 , \63310 , \63311 , \63312 ,
         \63313 , \63314 , \63315 , \63316 , \63317 , \63318 , \63319 , \63320 , \63321 , \63322 ,
         \63323 , \63324 , \63325 , \63326 , \63327 , \63328 , \63329 , \63330 , \63331 , \63332 ,
         \63333 , \63334 , \63335 , \63336 , \63337 , \63338 , \63339 , \63340 , \63341 , \63342 ,
         \63343 , \63344 , \63345 , \63346 , \63347 , \63348 , \63349 , \63350 , \63351 , \63352 ,
         \63353 , \63354 , \63355 , \63356 , \63357 , \63358 , \63359 , \63360 , \63361 , \63362 ,
         \63363 , \63364 , \63365 , \63366 , \63367 , \63368 , \63369 , \63370 , \63371 , \63372 ,
         \63373 , \63374 , \63375 , \63376 , \63377 , \63378 , \63379 , \63380 , \63381 , \63382 ,
         \63383 , \63384 , \63385 , \63386 , \63387 , \63388 , \63389 , \63390 , \63391 , \63392 ,
         \63393 , \63394 , \63395 , \63396 , \63397 , \63398 , \63399 , \63400 , \63401 , \63402 ,
         \63403 , \63404 , \63405 , \63406 , \63407 , \63408 , \63409 , \63410 , \63411 , \63412 ,
         \63413 , \63414 , \63415 , \63416 , \63417 , \63418 , \63419 , \63420 , \63421 , \63422 ,
         \63423 , \63424 , \63425 , \63426 , \63427 , \63428 , \63429 , \63430 , \63431 , \63432 ,
         \63433 , \63434 , \63435 , \63436 , \63437 , \63438 , \63439 , \63440 , \63441 , \63442 ,
         \63443 , \63444 , \63445 , \63446 , \63447 , \63448 , \63449 , \63450 , \63451 , \63452 ,
         \63453 , \63454 , \63455 , \63456 , \63457 , \63458 , \63459 , \63460 , \63461 , \63462 ,
         \63463 , \63464 , \63465 , \63466 , \63467 , \63468 , \63469 , \63470 , \63471 , \63472 ,
         \63473 , \63474 , \63475 , \63476 , \63477 , \63478 , \63479 , \63480 , \63481 , \63482 ,
         \63483 , \63484 , \63485 , \63486 , \63487 , \63488 , \63489 , \63490 , \63491 , \63492 ,
         \63493 , \63494 , \63495 , \63496 , \63497 , \63498 , \63499 , \63500 , \63501 , \63502 ,
         \63503 , \63504 , \63505 , \63506 , \63507 , \63508 , \63509 , \63510 , \63511 , \63512 ,
         \63513 , \63514 , \63515 , \63516 , \63517 , \63518 , \63519 , \63520 , \63521 , \63522 ,
         \63523 , \63524 , \63525 , \63526 , \63527 , \63528 , \63529 , \63530 , \63531 , \63532 ,
         \63533 , \63534 , \63535 , \63536 , \63537 , \63538 , \63539 , \63540 , \63541 , \63542 ,
         \63543 , \63544 , \63545 , \63546 , \63547 , \63548 , \63549 , \63550 , \63551 , \63552 ,
         \63553 , \63554 , \63555 , \63556 , \63557 , \63558 , \63559 , \63560 , \63561 , \63562 ,
         \63563 , \63564 , \63565 , \63566 , \63567 , \63568 , \63569 , \63570 , \63571 , \63572 ,
         \63573 , \63574 , \63575 , \63576 , \63577 , \63578 , \63579 , \63580 , \63581 , \63582 ,
         \63583 , \63584 , \63585 , \63586 , \63587 , \63588 , \63589 , \63590 , \63591 , \63592 ,
         \63593 , \63594 , \63595 , \63596 , \63597 , \63598 , \63599 , \63600 , \63601 , \63602 ,
         \63603 , \63604 , \63605 , \63606 , \63607 , \63608 , \63609 , \63610 , \63611 , \63612 ,
         \63613 , \63614 , \63615 , \63616 , \63617 , \63618 , \63619 , \63620 , \63621 , \63622 ,
         \63623 , \63624 , \63625 , \63626 , \63627 , \63628 , \63629 , \63630 , \63631 , \63632 ,
         \63633 , \63634 , \63635 , \63636 , \63637 , \63638 , \63639 , \63640 , \63641 , \63642 ,
         \63643 , \63644 , \63645 , \63646 , \63647 , \63648 , \63649 , \63650 , \63651 , \63652 ,
         \63653 , \63654 , \63655 , \63656 , \63657 , \63658 , \63659 , \63660 , \63661 , \63662 ,
         \63663 , \63664 , \63665 , \63666 , \63667 , \63668 , \63669 , \63670 , \63671 , \63672 ,
         \63673 , \63674 , \63675 , \63676 , \63677 , \63678 , \63679 , \63680 , \63681 , \63682 ,
         \63683 , \63684 , \63685 , \63686 , \63687 , \63688 , \63689 , \63690 , \63691 , \63692 ,
         \63693 , \63694 , \63695 , \63696 , \63697 , \63698 , \63699 , \63700 , \63701 , \63702 ,
         \63703 , \63704 , \63705 , \63706 , \63707 , \63708 , \63709 , \63710 , \63711 , \63712 ,
         \63713 , \63714 , \63715 , \63716 , \63717 , \63718 , \63719 , \63720 , \63721 , \63722 ,
         \63723 , \63724 , \63725 , \63726 , \63727 , \63728 , \63729 , \63730 , \63731 , \63732 ,
         \63733 , \63734 , \63735 , \63736 , \63737 , \63738 , \63739 , \63740 , \63741 , \63742 ,
         \63743 , \63744 , \63745 , \63746 , \63747 , \63748 , \63749 , \63750 , \63751 , \63752 ,
         \63753 , \63754 , \63755 , \63756 , \63757 , \63758 , \63759 , \63760 , \63761 , \63762 ,
         \63763 , \63764 , \63765 , \63766 , \63767 , \63768 , \63769 , \63770 , \63771 , \63772 ,
         \63773 , \63774 , \63775 , \63776 , \63777 , \63778 , \63779 , \63780 , \63781 , \63782 ,
         \63783 , \63784 , \63785 , \63786 , \63787 , \63788 , \63789 , \63790 , \63791 , \63792 ,
         \63793 , \63794 , \63795 , \63796 , \63797 , \63798 , \63799 , \63800 , \63801 , \63802 ,
         \63803 , \63804 , \63805 , \63806 , \63807 , \63808 , \63809 , \63810 , \63811 , \63812 ,
         \63813 , \63814 , \63815 , \63816 , \63817 , \63818 , \63819 , \63820 , \63821 , \63822 ,
         \63823 , \63824 , \63825 , \63826 , \63827 , \63828 , \63829 , \63830 , \63831 , \63832 ,
         \63833 , \63834 , \63835 , \63836 , \63837 , \63838 , \63839 , \63840 , \63841 , \63842 ,
         \63843 , \63844 , \63845 , \63846 , \63847 , \63848 , \63849 , \63850 , \63851 , \63852 ,
         \63853 , \63854 , \63855 , \63856 , \63857 , \63858 , \63859 , \63860 , \63861 , \63862 ,
         \63863 , \63864 , \63865 , \63866 , \63867 , \63868 , \63869 , \63870 , \63871 , \63872 ,
         \63873 , \63874 , \63875 , \63876 , \63877 , \63878 , \63879 , \63880 , \63881 , \63882 ,
         \63883 , \63884 , \63885 , \63886 , \63887 , \63888 , \63889 , \63890 , \63891 , \63892 ,
         \63893 , \63894 , \63895 , \63896 , \63897 , \63898 , \63899 , \63900 , \63901 , \63902 ,
         \63903 , \63904 , \63905 , \63906 , \63907 , \63908 , \63909 , \63910 , \63911 , \63912 ,
         \63913 , \63914 , \63915 , \63916 , \63917 , \63918 , \63919 , \63920 , \63921 , \63922 ,
         \63923 , \63924 , \63925 , \63926 , \63927 , \63928 , \63929 , \63930 , \63931 , \63932 ,
         \63933 , \63934 , \63935 , \63936 , \63937 , \63938 , \63939 , \63940 , \63941 , \63942 ,
         \63943 , \63944 , \63945 , \63946 , \63947 , \63948 , \63949 , \63950 , \63951 , \63952 ,
         \63953 , \63954 , \63955 , \63956 , \63957 , \63958 , \63959 , \63960 , \63961 , \63962 ,
         \63963 , \63964 , \63965 , \63966 , \63967 , \63968 , \63969 , \63970 , \63971 , \63972 ,
         \63973 , \63974 , \63975 , \63976 , \63977 , \63978 , \63979 , \63980 , \63981 , \63982 ,
         \63983 , \63984 , \63985 , \63986 , \63987 , \63988 , \63989 , \63990 , \63991 , \63992 ,
         \63993 , \63994 , \63995 , \63996 , \63997 , \63998 , \63999 , \64000 , \64001 , \64002 ,
         \64003 , \64004 , \64005 , \64006 , \64007 , \64008 , \64009 , \64010 , \64011 , \64012 ,
         \64013 , \64014 , \64015 , \64016 , \64017 , \64018 , \64019 , \64020 , \64021 , \64022 ,
         \64023 , \64024 , \64025 , \64026 , \64027 , \64028 , \64029 , \64030 , \64031 , \64032 ,
         \64033 , \64034 , \64035 , \64036 , \64037 , \64038 , \64039 , \64040 , \64041 , \64042 ,
         \64043 , \64044 , \64045 , \64046 , \64047 , \64048 , \64049 , \64050 , \64051 , \64052 ,
         \64053 , \64054 , \64055 , \64056 , \64057 , \64058 , \64059 , \64060 , \64061 , \64062 ,
         \64063 , \64064 , \64065 , \64066 , \64067 , \64068 , \64069 , \64070 , \64071 , \64072 ,
         \64073 , \64074 , \64075 , \64076 , \64077 , \64078 , \64079 , \64080 , \64081 , \64082 ,
         \64083 , \64084 , \64085 , \64086 , \64087 , \64088 , \64089 , \64090 , \64091 , \64092 ,
         \64093 , \64094 , \64095 , \64096 , \64097 , \64098 , \64099 , \64100 , \64101 , \64102 ,
         \64103 , \64104 , \64105 , \64106 , \64107 , \64108 , \64109 , \64110 , \64111 , \64112 ,
         \64113 , \64114 , \64115 , \64116 , \64117 , \64118 , \64119 , \64120 , \64121 , \64122 ,
         \64123 , \64124 , \64125 , \64126 , \64127 , \64128 , \64129 , \64130 , \64131 , \64132 ,
         \64133 , \64134 , \64135 , \64136 , \64137 , \64138 , \64139 , \64140 , \64141 , \64142 ,
         \64143 , \64144 , \64145 , \64146 , \64147 , \64148 , \64149 , \64150 , \64151 , \64152 ,
         \64153 , \64154 , \64155 , \64156 , \64157 , \64158 , \64159 , \64160 , \64161 , \64162 ,
         \64163 , \64164 , \64165 , \64166 , \64167 , \64168 , \64169 , \64170 , \64171 , \64172 ,
         \64173 , \64174 , \64175 , \64176 , \64177 , \64178 , \64179 , \64180 , \64181 , \64182 ,
         \64183 , \64184 , \64185 , \64186 , \64187 , \64188 , \64189 , \64190 , \64191 , \64192 ,
         \64193 , \64194 , \64195 , \64196 , \64197 , \64198 , \64199 , \64200 , \64201 , \64202 ,
         \64203 , \64204 , \64205 , \64206 , \64207 , \64208 , \64209 , \64210 , \64211 , \64212 ,
         \64213 , \64214 , \64215 , \64216 , \64217 , \64218 , \64219 , \64220 , \64221 , \64222 ,
         \64223 , \64224 , \64225 , \64226 , \64227 , \64228 , \64229 , \64230 , \64231 , \64232 ,
         \64233 , \64234 , \64235 , \64236 , \64237 , \64238 , \64239 , \64240 , \64241 , \64242 ,
         \64243 , \64244 , \64245 , \64246 , \64247 , \64248 , \64249 , \64250 , \64251 , \64252 ,
         \64253 , \64254 , \64255 , \64256 , \64257 , \64258 , \64259 , \64260 , \64261 , \64262 ,
         \64263 , \64264 , \64265 , \64266 , \64267 , \64268 , \64269 , \64270 , \64271 , \64272 ,
         \64273 , \64274 , \64275 , \64276 , \64277 , \64278 , \64279 , \64280 , \64281 , \64282 ,
         \64283 , \64284 , \64285 , \64286 , \64287 , \64288 , \64289 , \64290 , \64291 , \64292 ,
         \64293 , \64294 , \64295 , \64296 , \64297 , \64298 , \64299 , \64300 , \64301 , \64302 ,
         \64303 , \64304 , \64305 , \64306 , \64307 , \64308 , \64309 , \64310 , \64311 , \64312 ,
         \64313 , \64314 , \64315 , \64316 , \64317 , \64318 , \64319 , \64320 , \64321 , \64322 ,
         \64323 , \64324 , \64325 , \64326 , \64327 , \64328 , \64329 , \64330 , \64331 , \64332 ,
         \64333 , \64334 , \64335 , \64336 , \64337 , \64338 , \64339 , \64340 , \64341 , \64342 ,
         \64343 , \64344 , \64345 , \64346 , \64347 , \64348 , \64349 , \64350 , \64351 , \64352 ,
         \64353 , \64354 , \64355 , \64356 , \64357 , \64358 , \64359 , \64360 , \64361 , \64362 ,
         \64363 , \64364 , \64365 , \64366 , \64367 , \64368 , \64369 , \64370 , \64371 , \64372 ,
         \64373 , \64374 , \64375 , \64376 , \64377 , \64378 , \64379 , \64380 , \64381 , \64382 ,
         \64383 , \64384 , \64385 , \64386 , \64387 , \64388 , \64389 , \64390 , \64391 , \64392 ,
         \64393 , \64394 , \64395 , \64396 , \64397 , \64398 , \64399 , \64400 , \64401 , \64402 ,
         \64403 , \64404 , \64405 , \64406 , \64407 , \64408 , \64409 , \64410 , \64411 , \64412 ,
         \64413 , \64414 , \64415 , \64416 , \64417 , \64418 , \64419 , \64420 , \64421 , \64422 ,
         \64423 , \64424 , \64425 , \64426 , \64427 , \64428 , \64429 , \64430 , \64431 , \64432 ,
         \64433 , \64434 , \64435 , \64436 , \64437 , \64438 , \64439 , \64440 , \64441 , \64442 ,
         \64443 , \64444 , \64445 , \64446 , \64447 , \64448 , \64449 , \64450 , \64451 , \64452 ,
         \64453 , \64454 , \64455 , \64456 , \64457 , \64458 , \64459 , \64460 , \64461 , \64462 ,
         \64463 , \64464 , \64465 , \64466 , \64467 , \64468 , \64469 , \64470 , \64471 , \64472 ,
         \64473 , \64474 , \64475 , \64476 , \64477 , \64478 , \64479 , \64480 , \64481 , \64482 ,
         \64483 , \64484 , \64485 , \64486 , \64487 , \64488 , \64489 , \64490 , \64491 , \64492 ,
         \64493 , \64494 , \64495 , \64496 , \64497 , \64498 , \64499 , \64500 , \64501 , \64502 ,
         \64503 , \64504 , \64505 , \64506 , \64507 , \64508 , \64509 , \64510 , \64511 , \64512 ,
         \64513 , \64514 , \64515 , \64516 , \64517 , \64518 , \64519 , \64520 , \64521 , \64522 ,
         \64523 , \64524 , \64525 , \64526 , \64527 , \64528 , \64529 , \64530 , \64531 , \64532 ,
         \64533 , \64534 , \64535 , \64536 , \64537 , \64538 , \64539 , \64540 , \64541 , \64542 ,
         \64543 , \64544 , \64545 , \64546 , \64547 , \64548 , \64549 , \64550 , \64551 , \64552 ,
         \64553 , \64554 , \64555 , \64556 , \64557 , \64558 , \64559 , \64560 , \64561 , \64562 ,
         \64563 , \64564 , \64565 , \64566 , \64567 , \64568 , \64569 , \64570 , \64571 , \64572 ,
         \64573 , \64574 , \64575 , \64576 , \64577 , \64578 , \64579 , \64580 , \64581 , \64582 ,
         \64583 , \64584 , \64585 , \64586 , \64587 , \64588 , \64589 , \64590 , \64591 , \64592 ,
         \64593 , \64594 , \64595 , \64596 , \64597 , \64598 , \64599 , \64600 , \64601 , \64602 ,
         \64603 , \64604 , \64605 , \64606 , \64607 , \64608 , \64609 , \64610 , \64611 , \64612 ,
         \64613 , \64614 , \64615 , \64616 , \64617 , \64618 , \64619 , \64620 , \64621 , \64622 ,
         \64623 , \64624 , \64625 , \64626 , \64627 , \64628 , \64629 , \64630 , \64631 , \64632 ,
         \64633 , \64634 , \64635 , \64636 , \64637 , \64638 , \64639 , \64640 , \64641 , \64642 ,
         \64643 , \64644 , \64645 , \64646 , \64647 , \64648 , \64649 , \64650 , \64651 , \64652 ,
         \64653 , \64654 , \64655 , \64656 , \64657 , \64658 , \64659 , \64660 , \64661 , \64662 ,
         \64663 , \64664 , \64665 , \64666 , \64667 , \64668 , \64669 , \64670 , \64671 , \64672 ,
         \64673 , \64674 , \64675 , \64676 , \64677 , \64678 , \64679 , \64680 , \64681 , \64682 ,
         \64683 , \64684 , \64685 , \64686 , \64687 , \64688 , \64689 , \64690 , \64691 , \64692 ,
         \64693 , \64694 , \64695 , \64696 , \64697 , \64698 , \64699 , \64700 , \64701 , \64702 ,
         \64703 , \64704 , \64705 , \64706 , \64707 , \64708 , \64709 , \64710 , \64711 , \64712 ,
         \64713 , \64714 , \64715 , \64716 , \64717 , \64718 , \64719 , \64720 , \64721 , \64722 ,
         \64723 , \64724 , \64725 , \64726 , \64727 , \64728 , \64729 , \64730 , \64731 , \64732 ,
         \64733 , \64734 , \64735 , \64736 , \64737 , \64738 , \64739 , \64740 , \64741 , \64742 ,
         \64743 , \64744 , \64745 , \64746 , \64747 , \64748 , \64749 , \64750 , \64751 , \64752 ,
         \64753 , \64754 , \64755 , \64756 , \64757 , \64758 , \64759 , \64760 , \64761 , \64762 ,
         \64763 , \64764 , \64765 , \64766 , \64767 , \64768 , \64769 , \64770 , \64771 , \64772 ,
         \64773 , \64774 , \64775 , \64776 , \64777 , \64778 , \64779 , \64780 , \64781 , \64782 ,
         \64783 , \64784 , \64785 , \64786 , \64787 , \64788 , \64789 , \64790 , \64791 , \64792 ,
         \64793 , \64794 , \64795 , \64796 , \64797 , \64798 , \64799 , \64800 , \64801 , \64802 ,
         \64803 , \64804 , \64805 , \64806 , \64807 , \64808 , \64809 , \64810 , \64811 , \64812 ,
         \64813 , \64814 , \64815 , \64816 , \64817 , \64818 , \64819 , \64820 , \64821 , \64822 ,
         \64823 , \64824 , \64825 , \64826 , \64827 , \64828 , \64829 , \64830 , \64831 , \64832 ,
         \64833 , \64834 , \64835 , \64836 , \64837 , \64838 , \64839 , \64840 , \64841 , \64842 ,
         \64843 , \64844 , \64845 , \64846 , \64847 , \64848 , \64849 , \64850 , \64851 , \64852 ,
         \64853 , \64854 , \64855 , \64856 , \64857 , \64858 , \64859 , \64860 , \64861 , \64862 ,
         \64863 , \64864 , \64865 , \64866 , \64867 , \64868 , \64869 , \64870 , \64871 , \64872 ,
         \64873 , \64874 , \64875 , \64876 , \64877 , \64878 , \64879 , \64880 , \64881 , \64882 ,
         \64883 , \64884 , \64885 , \64886 , \64887 , \64888 , \64889 , \64890 , \64891 , \64892 ,
         \64893 , \64894 , \64895 , \64896 , \64897 , \64898 , \64899 , \64900 , \64901 , \64902 ,
         \64903 , \64904 , \64905 , \64906 , \64907 , \64908 , \64909 , \64910 , \64911 , \64912 ,
         \64913 , \64914 , \64915 , \64916 , \64917 , \64918 , \64919 , \64920 , \64921 , \64922 ,
         \64923 , \64924 , \64925 , \64926 , \64927 , \64928 , \64929 , \64930 , \64931 , \64932 ,
         \64933 , \64934 , \64935 , \64936 , \64937 , \64938 , \64939 , \64940 , \64941 , \64942 ,
         \64943 , \64944 , \64945 , \64946 , \64947 , \64948 , \64949 , \64950 , \64951 , \64952 ,
         \64953 , \64954 , \64955 , \64956 , \64957 , \64958 , \64959 , \64960 , \64961 , \64962 ,
         \64963 , \64964 , \64965 , \64966 , \64967 , \64968 , \64969 , \64970 , \64971 , \64972 ,
         \64973 , \64974 , \64975 , \64976 , \64977 , \64978 , \64979 , \64980 , \64981 , \64982 ,
         \64983 , \64984 , \64985 , \64986 , \64987 , \64988 , \64989 , \64990 , \64991 , \64992 ,
         \64993 , \64994 , \64995 , \64996 , \64997 , \64998 , \64999 , \65000 , \65001 , \65002 ,
         \65003 , \65004 , \65005 , \65006 , \65007 , \65008 , \65009 , \65010 , \65011 , \65012 ,
         \65013 , \65014 , \65015 , \65016 , \65017 , \65018 , \65019 , \65020 , \65021 , \65022 ,
         \65023 , \65024 , \65025 , \65026 , \65027 , \65028 , \65029 , \65030 , \65031 , \65032 ,
         \65033 , \65034 , \65035 , \65036 , \65037 , \65038 , \65039 , \65040 , \65041 , \65042 ,
         \65043 , \65044 , \65045 , \65046 , \65047 , \65048 , \65049 , \65050 , \65051 , \65052 ,
         \65053 , \65054 , \65055 , \65056 , \65057 , \65058 , \65059 , \65060 , \65061 , \65062 ,
         \65063 , \65064 , \65065 , \65066 , \65067 , \65068 , \65069 , \65070 , \65071 , \65072 ,
         \65073 , \65074 , \65075 , \65076 , \65077 , \65078 , \65079 , \65080 , \65081 , \65082 ,
         \65083 , \65084 , \65085 , \65086 , \65087 , \65088 , \65089 , \65090 , \65091 , \65092 ,
         \65093 , \65094 , \65095 , \65096 , \65097 , \65098 , \65099 , \65100 , \65101 , \65102 ,
         \65103 , \65104 , \65105 , \65106 , \65107 , \65108 , \65109 , \65110 , \65111 , \65112 ,
         \65113 , \65114 , \65115 , \65116 , \65117 , \65118 , \65119 , \65120 , \65121 , \65122 ,
         \65123 , \65124 , \65125 , \65126 , \65127 , \65128 , \65129 , \65130 , \65131 , \65132 ,
         \65133 , \65134 , \65135 , \65136 , \65137 , \65138 , \65139 , \65140 , \65141 , \65142 ,
         \65143 , \65144 , \65145 , \65146 , \65147 , \65148 , \65149 , \65150 , \65151 , \65152 ,
         \65153 , \65154 , \65155 , \65156 , \65157 , \65158 , \65159 , \65160 , \65161 , \65162 ,
         \65163 , \65164 , \65165 , \65166 , \65167 , \65168 , \65169 , \65170 , \65171 , \65172 ,
         \65173 , \65174 , \65175 , \65176 , \65177 , \65178 , \65179 , \65180 , \65181 , \65182 ,
         \65183 , \65184 , \65185 , \65186 , \65187 , \65188 , \65189 , \65190 , \65191 , \65192 ,
         \65193 , \65194 , \65195 , \65196 , \65197 , \65198 , \65199 , \65200 , \65201 , \65202 ,
         \65203 , \65204 , \65205 , \65206 , \65207 , \65208 , \65209 , \65210 , \65211 , \65212 ,
         \65213 , \65214 , \65215 , \65216 , \65217 , \65218 , \65219 , \65220 , \65221 , \65222 ,
         \65223 , \65224 , \65225 , \65226 , \65227 , \65228 , \65229 , \65230 , \65231 , \65232 ,
         \65233 , \65234 , \65235 , \65236 , \65237 , \65238 , \65239 , \65240 , \65241 , \65242 ,
         \65243 , \65244 , \65245 , \65246 , \65247 , \65248 , \65249 , \65250 , \65251 , \65252 ,
         \65253 , \65254 , \65255 , \65256 , \65257 , \65258 , \65259 , \65260 , \65261 , \65262 ,
         \65263 , \65264 , \65265 , \65266 , \65267 , \65268 , \65269 , \65270 , \65271 , \65272 ,
         \65273 , \65274 , \65275 , \65276 , \65277 , \65278 , \65279 , \65280 , \65281 , \65282 ,
         \65283 , \65284 , \65285 , \65286 , \65287 , \65288 , \65289 , \65290 , \65291 , \65292 ,
         \65293 , \65294 , \65295 , \65296 , \65297 , \65298 , \65299 , \65300 , \65301 , \65302 ,
         \65303 , \65304 , \65305 , \65306 , \65307 , \65308 , \65309 , \65310 , \65311 , \65312 ,
         \65313 , \65314 , \65315 , \65316 , \65317 , \65318 , \65319 , \65320 , \65321 , \65322 ,
         \65323 , \65324 , \65325 , \65326 , \65327 , \65328 , \65329 , \65330 , \65331 , \65332 ,
         \65333 , \65334 , \65335 , \65336 , \65337 , \65338 , \65339 , \65340 , \65341 , \65342 ,
         \65343 , \65344 , \65345 , \65346 , \65347 , \65348 , \65349 , \65350 , \65351 , \65352 ,
         \65353 , \65354 , \65355 , \65356 , \65357 , \65358 , \65359 , \65360 , \65361 , \65362 ,
         \65363 , \65364 , \65365 , \65366 , \65367 , \65368 , \65369 , \65370 , \65371 , \65372 ,
         \65373 , \65374 , \65375 , \65376 , \65377 , \65378 , \65379 , \65380 , \65381 , \65382 ,
         \65383 , \65384 , \65385 , \65386 , \65387 , \65388 , \65389 , \65390 , \65391 , \65392 ,
         \65393 , \65394 , \65395 , \65396 , \65397 , \65398 , \65399 , \65400 , \65401 , \65402 ,
         \65403 , \65404 , \65405 , \65406 , \65407 , \65408 , \65409 , \65410 , \65411 , \65412 ,
         \65413 , \65414 , \65415 , \65416 , \65417 , \65418 , \65419 , \65420 , \65421 , \65422 ,
         \65423 , \65424 , \65425 , \65426 , \65427 , \65428 , \65429 , \65430 , \65431 , \65432 ,
         \65433 , \65434 , \65435 , \65436 , \65437 , \65438 , \65439 , \65440 , \65441 , \65442 ,
         \65443 , \65444 , \65445 , \65446 , \65447 , \65448 , \65449 , \65450 , \65451 , \65452 ,
         \65453 , \65454 , \65455 , \65456 , \65457 , \65458 , \65459 , \65460 , \65461 , \65462 ,
         \65463 , \65464 , \65465 , \65466 , \65467 , \65468 , \65469 , \65470 , \65471 , \65472 ,
         \65473 , \65474 , \65475 , \65476 , \65477 , \65478 , \65479 , \65480 , \65481 , \65482 ,
         \65483 , \65484 , \65485 , \65486 , \65487 , \65488 , \65489 , \65490 , \65491 , \65492 ,
         \65493 , \65494 , \65495 , \65496 , \65497 , \65498 , \65499 , \65500 , \65501 , \65502 ,
         \65503 , \65504 , \65505 , \65506 , \65507 , \65508 , \65509 , \65510 , \65511 , \65512 ,
         \65513 , \65514 , \65515 , \65516 , \65517 , \65518 , \65519 , \65520 , \65521 , \65522 ,
         \65523 , \65524 , \65525 , \65526 , \65527 , \65528 , \65529 , \65530 , \65531 , \65532 ,
         \65533 , \65534 , \65535 , \65536 , \65537 , \65538 , \65539 , \65540 , \65541 , \65542 ,
         \65543 , \65544 , \65545 , \65546 , \65547 , \65548 , \65549 , \65550 , \65551 , \65552 ,
         \65553 , \65554 , \65555 , \65556 , \65557 , \65558 , \65559 , \65560 , \65561 , \65562 ,
         \65563 , \65564 , \65565 , \65566 , \65567 , \65568 , \65569 , \65570 , \65571 , \65572 ,
         \65573 , \65574 , \65575 , \65576 , \65577 , \65578 , \65579 , \65580 , \65581 , \65582 ,
         \65583 , \65584 , \65585 , \65586 , \65587 , \65588 , \65589 , \65590 , \65591 , \65592 ,
         \65593 , \65594 , \65595 , \65596 , \65597 , \65598 , \65599 , \65600 , \65601 , \65602 ,
         \65603 , \65604 , \65605 , \65606 , \65607 , \65608 , \65609 , \65610 , \65611 , \65612 ,
         \65613 , \65614 , \65615 , \65616 , \65617 , \65618 , \65619 , \65620 , \65621 , \65622 ,
         \65623 , \65624 , \65625 , \65626 , \65627 , \65628 , \65629 , \65630 , \65631 , \65632 ,
         \65633 , \65634 , \65635 , \65636 , \65637 , \65638 , \65639 , \65640 , \65641 , \65642 ,
         \65643 , \65644 , \65645 , \65646 , \65647 , \65648 , \65649 , \65650 , \65651 , \65652 ,
         \65653 , \65654 , \65655 , \65656 , \65657 , \65658 , \65659 , \65660 , \65661 , \65662 ,
         \65663 , \65664 , \65665 , \65666 , \65667 , \65668 , \65669 , \65670 , \65671 , \65672 ,
         \65673 , \65674 , \65675 , \65676 , \65677 , \65678 , \65679 , \65680 , \65681 , \65682 ,
         \65683 , \65684 , \65685 , \65686 , \65687 , \65688 , \65689 , \65690 , \65691 , \65692 ,
         \65693 , \65694 , \65695 , \65696 , \65697 , \65698 , \65699 , \65700 , \65701 , \65702 ,
         \65703 , \65704 , \65705 , \65706 , \65707 , \65708 , \65709 , \65710 , \65711 , \65712 ,
         \65713 , \65714 , \65715 , \65716 , \65717 , \65718 , \65719 , \65720 , \65721 , \65722 ,
         \65723 , \65724 , \65725 , \65726 , \65727 , \65728 , \65729 , \65730 , \65731 , \65732 ,
         \65733 , \65734 , \65735 , \65736 , \65737 , \65738 , \65739 , \65740 , \65741 , \65742 ,
         \65743 , \65744 , \65745 , \65746 , \65747 , \65748 , \65749 , \65750 , \65751 , \65752 ,
         \65753 , \65754 , \65755 , \65756 , \65757 , \65758 , \65759 , \65760 , \65761 , \65762 ,
         \65763 , \65764 , \65765 , \65766 , \65767 , \65768 , \65769 , \65770 , \65771 , \65772 ,
         \65773 , \65774 , \65775 , \65776 , \65777 , \65778 , \65779 , \65780 , \65781 , \65782 ,
         \65783 , \65784 , \65785 , \65786 , \65787 , \65788 , \65789 , \65790 , \65791 , \65792 ,
         \65793 , \65794 , \65795 , \65796 , \65797 , \65798 , \65799 , \65800 , \65801 , \65802 ,
         \65803 , \65804 , \65805 , \65806 , \65807 , \65808 , \65809 , \65810 , \65811 , \65812 ,
         \65813 , \65814 , \65815 , \65816 , \65817 , \65818 , \65819 , \65820 , \65821 , \65822 ,
         \65823 , \65824 , \65825 , \65826 , \65827 , \65828 , \65829 , \65830 , \65831 , \65832 ,
         \65833 , \65834 , \65835 , \65836 , \65837 , \65838 , \65839 , \65840 , \65841 , \65842 ,
         \65843 , \65844 , \65845 , \65846 , \65847 , \65848 , \65849 , \65850 , \65851 , \65852 ,
         \65853 , \65854 , \65855 , \65856 , \65857 , \65858 , \65859 , \65860 , \65861 , \65862 ,
         \65863 , \65864 , \65865 , \65866 , \65867 , \65868 , \65869 , \65870 , \65871 , \65872 ,
         \65873 , \65874 , \65875 , \65876 , \65877 , \65878 , \65879 , \65880 , \65881 , \65882 ,
         \65883 , \65884 , \65885 , \65886 , \65887 , \65888 , \65889 , \65890 , \65891 , \65892 ,
         \65893 , \65894 , \65895 , \65896 , \65897 , \65898 , \65899 , \65900 , \65901 , \65902 ,
         \65903 , \65904 , \65905 , \65906 , \65907 , \65908 , \65909 , \65910 , \65911 , \65912 ,
         \65913 , \65914 , \65915 , \65916 , \65917 , \65918 , \65919 , \65920 , \65921 , \65922 ,
         \65923 , \65924 , \65925 , \65926 , \65927 , \65928 , \65929 , \65930 , \65931 , \65932 ,
         \65933 , \65934 , \65935 , \65936 , \65937 , \65938 , \65939 , \65940 , \65941 , \65942 ,
         \65943 , \65944 , \65945 , \65946 , \65947 , \65948 , \65949 , \65950 , \65951 , \65952 ,
         \65953 , \65954 , \65955 , \65956 , \65957 , \65958 , \65959 , \65960 , \65961 , \65962 ,
         \65963 , \65964 , \65965 , \65966 , \65967 , \65968 , \65969 , \65970 , \65971 , \65972 ,
         \65973 , \65974 , \65975 , \65976 , \65977 , \65978 , \65979 , \65980 , \65981 , \65982 ,
         \65983 , \65984 , \65985 , \65986 , \65987 , \65988 , \65989 , \65990 , \65991 , \65992 ,
         \65993 , \65994 , \65995 , \65996 , \65997 , \65998 , \65999 , \66000 , \66001 , \66002 ,
         \66003 , \66004 , \66005 , \66006 , \66007 , \66008 , \66009 , \66010 , \66011 , \66012 ,
         \66013 , \66014 , \66015 , \66016 , \66017 , \66018 , \66019 , \66020 , \66021 , \66022 ,
         \66023 , \66024 , \66025 , \66026 , \66027 , \66028 , \66029 , \66030 , \66031 , \66032 ,
         \66033 , \66034 , \66035 , \66036 , \66037 , \66038 , \66039 , \66040 , \66041 , \66042 ,
         \66043 , \66044 , \66045 , \66046 , \66047 , \66048 , \66049 , \66050 , \66051 , \66052 ,
         \66053 , \66054 , \66055 , \66056 , \66057 , \66058 , \66059 , \66060 , \66061 , \66062 ,
         \66063 , \66064 , \66065 , \66066 , \66067 , \66068 , \66069 , \66070 , \66071 , \66072 ,
         \66073 , \66074 , \66075 , \66076 , \66077 , \66078 , \66079 , \66080 , \66081 , \66082 ,
         \66083 , \66084 , \66085 , \66086 , \66087 , \66088 , \66089 , \66090 , \66091 , \66092 ,
         \66093 , \66094 , \66095 , \66096 , \66097 , \66098 , \66099 , \66100 , \66101 , \66102 ,
         \66103 , \66104 , \66105 , \66106 , \66107 , \66108 , \66109 , \66110 , \66111 , \66112 ,
         \66113 , \66114 , \66115 , \66116 , \66117 , \66118 , \66119 , \66120 , \66121 , \66122 ,
         \66123 , \66124 , \66125 , \66126 , \66127 , \66128 , \66129 , \66130 , \66131 , \66132 ,
         \66133 , \66134 , \66135 , \66136 , \66137 , \66138 , \66139 , \66140 , \66141 , \66142 ,
         \66143 , \66144 , \66145 , \66146 , \66147 , \66148 , \66149 , \66150 , \66151 , \66152 ,
         \66153 , \66154 , \66155 , \66156 , \66157 , \66158 , \66159 , \66160 , \66161 , \66162 ,
         \66163 , \66164 , \66165 , \66166 , \66167 , \66168 , \66169 , \66170 , \66171 , \66172 ,
         \66173 , \66174 , \66175 , \66176 , \66177 , \66178 , \66179 , \66180 , \66181 , \66182 ,
         \66183 , \66184 , \66185 , \66186 , \66187 , \66188 , \66189 , \66190 , \66191 , \66192 ,
         \66193 , \66194 , \66195 , \66196 , \66197 , \66198 , \66199 , \66200 , \66201 , \66202 ,
         \66203 , \66204 , \66205 , \66206 , \66207 , \66208 , \66209 , \66210 , \66211 , \66212 ,
         \66213 , \66214 , \66215 , \66216 , \66217 , \66218 , \66219 , \66220 , \66221 , \66222 ,
         \66223 , \66224 , \66225 , \66226 , \66227 , \66228 , \66229 , \66230 , \66231 , \66232 ,
         \66233 , \66234 , \66235 , \66236 , \66237 , \66238 , \66239 , \66240 , \66241 , \66242 ,
         \66243 , \66244 , \66245 , \66246 , \66247 , \66248 , \66249 , \66250 , \66251 , \66252 ,
         \66253 , \66254 , \66255 , \66256 , \66257 , \66258 , \66259 , \66260 , \66261 , \66262 ,
         \66263 , \66264 , \66265 , \66266 , \66267 , \66268 , \66269 , \66270 , \66271 , \66272 ,
         \66273 , \66274 , \66275 , \66276 , \66277 , \66278 , \66279 , \66280 , \66281 , \66282 ,
         \66283 , \66284 , \66285 , \66286 , \66287 , \66288 , \66289 , \66290 , \66291 , \66292 ,
         \66293 , \66294 , \66295 , \66296 , \66297 , \66298 , \66299 , \66300 , \66301 , \66302 ,
         \66303 , \66304 , \66305 , \66306 , \66307 , \66308 , \66309 , \66310 , \66311 , \66312 ,
         \66313 , \66314 , \66315 , \66316 , \66317 , \66318 , \66319 , \66320 , \66321 , \66322 ,
         \66323 , \66324 , \66325 , \66326 , \66327 , \66328 , \66329 , \66330 , \66331 , \66332 ,
         \66333 , \66334 , \66335 , \66336 , \66337 , \66338 , \66339 , \66340 , \66341 , \66342 ,
         \66343 , \66344 , \66345 , \66346 , \66347 , \66348 , \66349 , \66350 , \66351 , \66352 ,
         \66353 , \66354 , \66355 , \66356 , \66357 , \66358 , \66359 , \66360 , \66361 , \66362 ,
         \66363 , \66364 , \66365 , \66366 , \66367 , \66368 , \66369 , \66370 , \66371 , \66372 ,
         \66373 , \66374 , \66375 , \66376 , \66377 , \66378 , \66379 , \66380 , \66381 , \66382 ,
         \66383 , \66384 , \66385 , \66386 , \66387 , \66388 , \66389 , \66390 , \66391 , \66392 ,
         \66393 , \66394 , \66395 , \66396 , \66397 , \66398 , \66399 , \66400 , \66401 , \66402 ,
         \66403 , \66404 , \66405 , \66406 , \66407 , \66408 , \66409 , \66410 , \66411 , \66412 ,
         \66413 , \66414 , \66415 , \66416 , \66417 , \66418 , \66419 , \66420 , \66421 , \66422 ,
         \66423 , \66424 , \66425 , \66426 , \66427 , \66428 , \66429 , \66430 , \66431 , \66432 ,
         \66433 , \66434 , \66435 , \66436 , \66437 , \66438 , \66439 , \66440 , \66441 , \66442 ,
         \66443 , \66444 , \66445 , \66446 , \66447 , \66448 , \66449 , \66450 , \66451 , \66452 ,
         \66453 , \66454 , \66455 , \66456 , \66457 , \66458 , \66459 , \66460 , \66461 , \66462 ,
         \66463 , \66464 , \66465 , \66466 , \66467 , \66468 , \66469 , \66470 , \66471 , \66472 ,
         \66473 , \66474 , \66475 , \66476 , \66477 , \66478 , \66479 , \66480 , \66481 , \66482 ,
         \66483 , \66484 , \66485 , \66486 , \66487 , \66488 , \66489 , \66490 , \66491 , \66492 ,
         \66493 , \66494 , \66495 , \66496 , \66497 , \66498 , \66499 , \66500 , \66501 , \66502 ,
         \66503 , \66504 , \66505 , \66506 , \66507 , \66508 , \66509 , \66510 , \66511 , \66512 ,
         \66513 , \66514 , \66515 , \66516 , \66517 , \66518 , \66519 , \66520 , \66521 , \66522 ,
         \66523 , \66524 , \66525 , \66526 , \66527 , \66528 , \66529 , \66530 , \66531 , \66532 ,
         \66533 , \66534 , \66535 , \66536 , \66537 , \66538 , \66539 , \66540 , \66541 , \66542 ,
         \66543 , \66544 , \66545 , \66546 , \66547 , \66548 , \66549 , \66550 , \66551 , \66552 ,
         \66553 , \66554 , \66555 , \66556 , \66557 , \66558 , \66559 , \66560 , \66561 , \66562 ,
         \66563 , \66564 , \66565 , \66566 , \66567 , \66568 , \66569 , \66570 , \66571 , \66572 ,
         \66573 , \66574 , \66575 , \66576 , \66577 , \66578 , \66579 , \66580 , \66581 , \66582 ,
         \66583 , \66584 , \66585 , \66586 , \66587 , \66588 , \66589 , \66590 , \66591 , \66592 ,
         \66593 , \66594 , \66595 , \66596 , \66597 , \66598 , \66599 , \66600 , \66601 , \66602 ,
         \66603 , \66604 , \66605 , \66606 , \66607 , \66608 , \66609 , \66610 , \66611 , \66612 ,
         \66613 , \66614 , \66615 , \66616 , \66617 , \66618 , \66619 , \66620 , \66621 , \66622 ,
         \66623 , \66624 , \66625 , \66626 , \66627 , \66628 , \66629 , \66630 , \66631 , \66632 ,
         \66633 , \66634 , \66635 , \66636 , \66637 , \66638 , \66639 , \66640 , \66641 , \66642 ,
         \66643 , \66644 , \66645 , \66646 , \66647 , \66648 , \66649 , \66650 , \66651 , \66652 ,
         \66653 , \66654 , \66655 , \66656 , \66657 , \66658 , \66659 , \66660 , \66661 , \66662 ,
         \66663 , \66664 , \66665 , \66666 , \66667 , \66668 , \66669 , \66670 , \66671 , \66672 ,
         \66673 , \66674 , \66675 , \66676 , \66677 , \66678 , \66679 , \66680 , \66681 , \66682 ,
         \66683 , \66684 , \66685 , \66686 , \66687 , \66688 , \66689 , \66690 , \66691 , \66692 ,
         \66693 , \66694 , \66695 , \66696 , \66697 , \66698 , \66699 , \66700 , \66701 , \66702 ,
         \66703 , \66704 , \66705 , \66706 , \66707 , \66708 , \66709 , \66710 , \66711 , \66712 ,
         \66713 , \66714 , \66715 , \66716 , \66717 , \66718 , \66719 , \66720 , \66721 , \66722 ,
         \66723 , \66724 , \66725 , \66726 , \66727 , \66728 , \66729 , \66730 , \66731 , \66732 ,
         \66733 , \66734 , \66735 , \66736 , \66737 , \66738 , \66739 , \66740 , \66741 , \66742 ,
         \66743 , \66744 , \66745 , \66746 , \66747 , \66748 , \66749 , \66750 , \66751 , \66752 ,
         \66753 , \66754 , \66755 , \66756 , \66757 , \66758 , \66759 , \66760 , \66761 , \66762 ,
         \66763 , \66764 , \66765 , \66766 , \66767 , \66768 , \66769 , \66770 , \66771 , \66772 ,
         \66773 , \66774 , \66775 , \66776 , \66777 , \66778 , \66779 , \66780 , \66781 , \66782 ,
         \66783 , \66784 , \66785 , \66786 , \66787 , \66788 , \66789 , \66790 , \66791 , \66792 ,
         \66793 , \66794 , \66795 , \66796 , \66797 , \66798 , \66799 , \66800 , \66801 , \66802 ,
         \66803 , \66804 , \66805 , \66806 , \66807 , \66808 , \66809 , \66810 , \66811 , \66812 ,
         \66813 , \66814 , \66815 , \66816 , \66817 , \66818 , \66819 , \66820 , \66821 , \66822 ,
         \66823 , \66824 , \66825 , \66826 , \66827 , \66828 , \66829 , \66830 , \66831 , \66832 ,
         \66833 , \66834 , \66835 , \66836 , \66837 , \66838 , \66839 , \66840 , \66841 , \66842 ,
         \66843 , \66844 , \66845 , \66846 , \66847 , \66848 , \66849 , \66850 , \66851 , \66852 ,
         \66853 , \66854 , \66855 , \66856 , \66857 , \66858 , \66859 , \66860 , \66861 , \66862 ,
         \66863 , \66864 , \66865 , \66866 , \66867 , \66868 , \66869 , \66870 , \66871 , \66872 ,
         \66873 , \66874 , \66875 , \66876 , \66877 , \66878 , \66879 , \66880 , \66881 , \66882 ,
         \66883 , \66884 , \66885 , \66886 , \66887 , \66888 , \66889 , \66890 , \66891 , \66892 ,
         \66893 , \66894 , \66895 , \66896 , \66897 , \66898 , \66899 , \66900 , \66901 , \66902 ,
         \66903 , \66904 , \66905 , \66906 , \66907 , \66908 , \66909 , \66910 , \66911 , \66912 ,
         \66913 , \66914 , \66915 , \66916 , \66917 , \66918 , \66919 , \66920 , \66921 , \66922 ,
         \66923 , \66924 , \66925 , \66926 , \66927 , \66928 , \66929 , \66930 , \66931 , \66932 ,
         \66933 , \66934 , \66935 , \66936 , \66937 , \66938 , \66939 , \66940 , \66941 , \66942 ,
         \66943 , \66944 , \66945 , \66946 , \66947 , \66948 , \66949 , \66950 , \66951 , \66952 ,
         \66953 , \66954 , \66955 , \66956 , \66957 , \66958 , \66959 , \66960 , \66961 , \66962 ,
         \66963 , \66964 , \66965 , \66966 , \66967 , \66968 , \66969 , \66970 , \66971 , \66972 ,
         \66973 , \66974 , \66975 , \66976 , \66977 , \66978 , \66979 , \66980 , \66981 , \66982 ,
         \66983 , \66984 , \66985 , \66986 , \66987 , \66988 , \66989 , \66990 , \66991 , \66992 ,
         \66993 , \66994 , \66995 , \66996 , \66997 , \66998 , \66999 , \67000 , \67001 , \67002 ,
         \67003 , \67004 , \67005 , \67006 , \67007 , \67008 , \67009 , \67010 , \67011 , \67012 ,
         \67013 , \67014 , \67015 , \67016 , \67017 , \67018 , \67019 , \67020 , \67021 , \67022 ,
         \67023 , \67024 , \67025 , \67026 , \67027 , \67028 , \67029 , \67030 , \67031 , \67032 ,
         \67033 , \67034 , \67035 , \67036 , \67037 , \67038 , \67039 , \67040 , \67041 , \67042 ,
         \67043 , \67044 , \67045 , \67046 , \67047 , \67048 , \67049 , \67050 , \67051 , \67052 ,
         \67053 , \67054 , \67055 , \67056 , \67057 , \67058 , \67059 , \67060 , \67061 , \67062 ,
         \67063 , \67064 , \67065 , \67066 , \67067 , \67068 , \67069 , \67070 , \67071 , \67072 ,
         \67073 , \67074 , \67075 , \67076 , \67077 , \67078 , \67079 , \67080 , \67081 , \67082 ,
         \67083 , \67084 , \67085 , \67086 , \67087 , \67088 , \67089 , \67090 , \67091 , \67092 ,
         \67093 , \67094 , \67095 , \67096 , \67097 , \67098 , \67099 , \67100 , \67101 , \67102 ,
         \67103 , \67104 , \67105 , \67106 , \67107 , \67108 , \67109 , \67110 , \67111 , \67112 ,
         \67113 , \67114 , \67115 , \67116 , \67117 , \67118 , \67119 , \67120 , \67121 , \67122 ,
         \67123 , \67124 , \67125 , \67126 , \67127 , \67128 , \67129 , \67130 , \67131 , \67132 ,
         \67133 , \67134 , \67135 , \67136 , \67137 , \67138 , \67139 , \67140 , \67141 , \67142 ,
         \67143 , \67144 , \67145 , \67146 , \67147 , \67148 , \67149 , \67150 , \67151 , \67152 ,
         \67153 , \67154 , \67155 , \67156 , \67157 , \67158 , \67159 , \67160 , \67161 , \67162 ,
         \67163 , \67164 , \67165 , \67166 , \67167 , \67168 , \67169 , \67170 , \67171 , \67172 ,
         \67173 , \67174 , \67175 , \67176 , \67177 , \67178 , \67179 , \67180 , \67181 , \67182 ,
         \67183 , \67184 , \67185 , \67186 , \67187 , \67188 , \67189 , \67190 , \67191 , \67192 ,
         \67193 , \67194 , \67195 , \67196 , \67197 , \67198 , \67199 , \67200 , \67201 , \67202 ,
         \67203 , \67204 , \67205 , \67206 , \67207 , \67208 , \67209 , \67210 , \67211 , \67212 ,
         \67213 , \67214 , \67215 , \67216 , \67217 , \67218 , \67219 , \67220 , \67221 , \67222 ,
         \67223 , \67224 , \67225 , \67226 , \67227 , \67228 , \67229 , \67230 , \67231 , \67232 ,
         \67233 , \67234 , \67235 , \67236 , \67237 , \67238 , \67239 , \67240 , \67241 , \67242 ,
         \67243 , \67244 , \67245 , \67246 , \67247 , \67248 , \67249 , \67250 , \67251 , \67252 ,
         \67253 , \67254 , \67255 , \67256 , \67257 , \67258 , \67259 , \67260 , \67261 , \67262 ,
         \67263 , \67264 , \67265 , \67266 , \67267 , \67268 , \67269 , \67270 , \67271 , \67272 ,
         \67273 , \67274 , \67275 , \67276 , \67277 , \67278 , \67279 , \67280 , \67281 , \67282 ,
         \67283 , \67284 , \67285 , \67286 , \67287 , \67288 , \67289 , \67290 , \67291 , \67292 ,
         \67293 , \67294 , \67295 , \67296 , \67297 , \67298 , \67299 , \67300 , \67301 , \67302 ,
         \67303 , \67304 , \67305 , \67306 , \67307 , \67308 , \67309 , \67310 , \67311 , \67312 ,
         \67313 , \67314 , \67315 , \67316 , \67317 , \67318 , \67319 , \67320 , \67321 , \67322 ,
         \67323 , \67324 , \67325 , \67326 , \67327 , \67328 , \67329 , \67330 , \67331 , \67332 ,
         \67333 , \67334 , \67335 , \67336 , \67337 , \67338 , \67339 , \67340 , \67341 , \67342 ,
         \67343 , \67344 , \67345 , \67346 , \67347 , \67348 , \67349 , \67350 , \67351 , \67352 ,
         \67353 , \67354 , \67355 , \67356 , \67357 , \67358 , \67359 , \67360 , \67361 , \67362 ,
         \67363 , \67364 , \67365 , \67366 , \67367 , \67368 , \67369 , \67370 , \67371 , \67372 ,
         \67373 , \67374 , \67375 , \67376 , \67377 , \67378 , \67379 , \67380 , \67381 , \67382 ,
         \67383 , \67384 , \67385 , \67386 , \67387 , \67388 , \67389 , \67390 , \67391 , \67392 ,
         \67393 , \67394 , \67395 , \67396 , \67397 , \67398 , \67399 , \67400 , \67401 , \67402 ,
         \67403 , \67404 , \67405 , \67406 , \67407 , \67408 , \67409 , \67410 , \67411 , \67412 ,
         \67413 , \67414 , \67415 , \67416 , \67417 , \67418 , \67419 , \67420 , \67421 , \67422 ,
         \67423 , \67424 , \67425 , \67426 , \67427 , \67428 , \67429 , \67430 , \67431 , \67432 ,
         \67433 , \67434 , \67435 , \67436 , \67437 , \67438 , \67439 , \67440 , \67441 , \67442 ,
         \67443 , \67444 , \67445 , \67446 , \67447 , \67448 , \67449 , \67450 , \67451 , \67452 ,
         \67453 , \67454 , \67455 , \67456 , \67457 , \67458 , \67459 , \67460 , \67461 , \67462 ,
         \67463 , \67464 , \67465 , \67466 , \67467 , \67468 , \67469 , \67470 , \67471 , \67472 ,
         \67473 , \67474 , \67475 , \67476 , \67477 , \67478 , \67479 , \67480 , \67481 , \67482 ,
         \67483 , \67484 , \67485 , \67486 , \67487 , \67488 , \67489 , \67490 , \67491 , \67492 ,
         \67493 , \67494 , \67495 , \67496 , \67497 , \67498 , \67499 , \67500 , \67501 , \67502 ,
         \67503 , \67504 , \67505 , \67506 , \67507 , \67508 , \67509 , \67510 , \67511 , \67512 ,
         \67513 , \67514 , \67515 , \67516 , \67517 , \67518 , \67519 , \67520 , \67521 , \67522 ,
         \67523 , \67524 , \67525 , \67526 , \67527 , \67528 , \67529 , \67530 , \67531 , \67532 ,
         \67533 , \67534 , \67535 , \67536 , \67537 , \67538 , \67539 , \67540 , \67541 , \67542 ,
         \67543 , \67544 , \67545 , \67546 , \67547 , \67548 , \67549 , \67550 , \67551 , \67552 ,
         \67553 , \67554 , \67555 , \67556 , \67557 , \67558 , \67559 , \67560 , \67561 , \67562 ,
         \67563 , \67564 , \67565 , \67566 , \67567 , \67568 , \67569 , \67570 , \67571 , \67572 ,
         \67573 , \67574 , \67575 , \67576 , \67577 , \67578 , \67579 , \67580 , \67581 , \67582 ,
         \67583 , \67584 , \67585 , \67586 , \67587 , \67588 , \67589 , \67590 , \67591 , \67592 ,
         \67593 , \67594 , \67595 , \67596 , \67597 , \67598 , \67599 , \67600 , \67601 , \67602 ,
         \67603 , \67604 , \67605 , \67606 , \67607 , \67608 , \67609 , \67610 , \67611 , \67612 ,
         \67613 , \67614 , \67615 , \67616 , \67617 , \67618 , \67619 , \67620 , \67621 , \67622 ,
         \67623 , \67624 , \67625 , \67626 , \67627 , \67628 , \67629 , \67630 , \67631 , \67632 ,
         \67633 , \67634 , \67635 , \67636 , \67637 , \67638 , \67639 , \67640 , \67641 , \67642 ,
         \67643 , \67644 , \67645 , \67646 , \67647 , \67648 , \67649 , \67650 , \67651 , \67652 ,
         \67653 , \67654 , \67655 , \67656 , \67657 , \67658 , \67659 , \67660 , \67661 , \67662 ,
         \67663 , \67664 , \67665 , \67666 , \67667 , \67668 , \67669 , \67670 , \67671 , \67672 ,
         \67673 , \67674 , \67675 , \67676 , \67677 , \67678 , \67679 , \67680 , \67681 , \67682 ,
         \67683 , \67684 , \67685 , \67686 , \67687 , \67688 , \67689 , \67690 , \67691 , \67692 ,
         \67693 , \67694 , \67695 , \67696 , \67697 , \67698 , \67699 , \67700 , \67701 , \67702 ,
         \67703 , \67704 , \67705 , \67706 , \67707 , \67708 , \67709 , \67710 , \67711 , \67712 ,
         \67713 , \67714 , \67715 , \67716 , \67717 , \67718 , \67719 , \67720 , \67721 , \67722 ,
         \67723 , \67724 , \67725 , \67726 , \67727 , \67728 , \67729 , \67730 , \67731 , \67732 ,
         \67733 , \67734 , \67735 , \67736 , \67737 , \67738 , \67739 , \67740 , \67741 , \67742 ,
         \67743 , \67744 , \67745 , \67746 , \67747 , \67748 , \67749 , \67750 , \67751 , \67752 ,
         \67753 , \67754 , \67755 , \67756 , \67757 , \67758 , \67759 , \67760 , \67761 , \67762 ,
         \67763 , \67764 , \67765 , \67766 , \67767 , \67768 , \67769 , \67770 , \67771 , \67772 ,
         \67773 , \67774 , \67775 , \67776 , \67777 , \67778 , \67779 , \67780 , \67781 , \67782 ,
         \67783 , \67784 , \67785 , \67786 , \67787 , \67788 , \67789 , \67790 , \67791 , \67792 ,
         \67793 , \67794 , \67795 , \67796 , \67797 , \67798 , \67799 , \67800 , \67801 , \67802 ,
         \67803 , \67804 , \67805 , \67806 , \67807 , \67808 , \67809 , \67810 , \67811 , \67812 ,
         \67813 , \67814 , \67815 , \67816 , \67817 , \67818 , \67819 , \67820 , \67821 , \67822 ,
         \67823 , \67824 , \67825 , \67826 , \67827 , \67828 , \67829 , \67830 , \67831 , \67832 ,
         \67833 , \67834 , \67835 , \67836 , \67837 , \67838 , \67839 , \67840 , \67841 , \67842 ,
         \67843 , \67844 , \67845 , \67846 , \67847 , \67848 , \67849 , \67850 , \67851 , \67852 ,
         \67853 , \67854 , \67855 , \67856 , \67857 , \67858 , \67859 , \67860 , \67861 , \67862 ,
         \67863 , \67864 , \67865 , \67866 , \67867 , \67868 , \67869 , \67870 , \67871 , \67872 ,
         \67873 , \67874 , \67875 , \67876 , \67877 , \67878 , \67879 , \67880 , \67881 , \67882 ,
         \67883 , \67884 , \67885 , \67886 , \67887 , \67888 , \67889 , \67890 , \67891 , \67892 ,
         \67893 , \67894 , \67895 , \67896 , \67897 , \67898 , \67899 , \67900 , \67901 , \67902 ,
         \67903 , \67904 , \67905 , \67906 , \67907 , \67908 , \67909 , \67910 , \67911 , \67912 ,
         \67913 , \67914 , \67915 , \67916 , \67917 , \67918 , \67919 , \67920 , \67921 , \67922 ,
         \67923 , \67924 , \67925 , \67926 , \67927 , \67928 , \67929 , \67930 , \67931 , \67932 ,
         \67933 , \67934 , \67935 , \67936 , \67937 , \67938 , \67939 , \67940 , \67941 , \67942 ,
         \67943 , \67944 , \67945 , \67946 , \67947 , \67948 , \67949 , \67950 , \67951 , \67952 ,
         \67953 , \67954 , \67955 , \67956 , \67957 , \67958 , \67959 , \67960 , \67961 , \67962 ,
         \67963 , \67964 , \67965 , \67966 , \67967 , \67968 , \67969 , \67970 , \67971 , \67972 ,
         \67973 , \67974 , \67975 , \67976 , \67977 , \67978 , \67979 , \67980 , \67981 , \67982 ,
         \67983 , \67984 , \67985 , \67986 , \67987 , \67988 , \67989 , \67990 , \67991 , \67992 ,
         \67993 , \67994 , \67995 , \67996 , \67997 , \67998 , \67999 , \68000 , \68001 , \68002 ,
         \68003 , \68004 , \68005 , \68006 , \68007 , \68008 , \68009 , \68010 , \68011 , \68012 ,
         \68013 , \68014 , \68015 , \68016 , \68017 , \68018 , \68019 , \68020 , \68021 , \68022 ,
         \68023 , \68024 , \68025 , \68026 , \68027 , \68028 , \68029 , \68030 , \68031 , \68032 ,
         \68033 , \68034 , \68035 , \68036 , \68037 , \68038 , \68039 , \68040 , \68041 , \68042 ,
         \68043 , \68044 , \68045 , \68046 , \68047 , \68048 , \68049 , \68050 , \68051 , \68052 ,
         \68053 , \68054 , \68055 , \68056 , \68057 , \68058 , \68059 , \68060 , \68061 , \68062 ,
         \68063 , \68064 , \68065 , \68066 , \68067 , \68068 , \68069 , \68070 , \68071 , \68072 ,
         \68073 , \68074 , \68075 , \68076 , \68077 , \68078 , \68079 , \68080 , \68081 , \68082 ,
         \68083 , \68084 , \68085 , \68086 , \68087 , \68088 , \68089 , \68090 , \68091 , \68092 ,
         \68093 , \68094 , \68095 , \68096 , \68097 , \68098 , \68099 , \68100 , \68101 , \68102 ,
         \68103 , \68104 , \68105 , \68106 , \68107 , \68108 , \68109 , \68110 , \68111 , \68112 ,
         \68113 , \68114 , \68115 , \68116 , \68117 , \68118 , \68119 , \68120 , \68121 , \68122 ,
         \68123 , \68124 , \68125 , \68126 , \68127 , \68128 , \68129 , \68130 , \68131 , \68132 ,
         \68133 , \68134 , \68135 , \68136 , \68137 , \68138 , \68139 , \68140 , \68141 , \68142 ,
         \68143 , \68144 , \68145 , \68146 , \68147 , \68148 , \68149 , \68150 , \68151 , \68152 ,
         \68153 , \68154 , \68155 , \68156 , \68157 , \68158 , \68159 , \68160 , \68161 , \68162 ,
         \68163 , \68164 , \68165 , \68166 , \68167 , \68168 , \68169 , \68170 , \68171 , \68172 ,
         \68173 , \68174 , \68175 , \68176 , \68177 , \68178 , \68179 , \68180 , \68181 , \68182 ,
         \68183 , \68184 , \68185 , \68186 , \68187 , \68188 , \68189 , \68190 , \68191 , \68192 ,
         \68193 , \68194 , \68195 , \68196 , \68197 , \68198 , \68199 , \68200 , \68201 , \68202 ,
         \68203 , \68204 , \68205 , \68206 , \68207 , \68208 , \68209 , \68210 , \68211 , \68212 ,
         \68213 , \68214 , \68215 , \68216 , \68217 , \68218 , \68219 , \68220 , \68221 , \68222 ,
         \68223 , \68224 , \68225 , \68226 , \68227 , \68228 , \68229 , \68230 , \68231 , \68232 ,
         \68233 , \68234 , \68235 , \68236 , \68237 , \68238 , \68239 , \68240 , \68241 , \68242 ,
         \68243 , \68244 , \68245 , \68246 , \68247 , \68248 , \68249 , \68250 , \68251 , \68252 ,
         \68253 , \68254 , \68255 , \68256 , \68257 , \68258 , \68259 , \68260 , \68261 , \68262 ,
         \68263 , \68264 , \68265 , \68266 , \68267 , \68268 , \68269 , \68270 , \68271 , \68272 ,
         \68273 , \68274 , \68275 , \68276 , \68277 , \68278 , \68279 , \68280 , \68281 , \68282 ,
         \68283 , \68284 , \68285 , \68286 , \68287 , \68288 , \68289 , \68290 , \68291 , \68292 ,
         \68293 , \68294 , \68295 , \68296 , \68297 , \68298 , \68299 , \68300 , \68301 , \68302 ,
         \68303 , \68304 , \68305 , \68306 , \68307 , \68308 , \68309 , \68310 , \68311 , \68312 ,
         \68313 , \68314 , \68315 , \68316 , \68317 , \68318 , \68319 , \68320 , \68321 , \68322 ,
         \68323 , \68324 , \68325 , \68326 , \68327 , \68328 , \68329 , \68330 , \68331 , \68332 ,
         \68333 , \68334 , \68335 , \68336 , \68337 , \68338 , \68339 , \68340 , \68341 , \68342 ,
         \68343 , \68344 , \68345 , \68346 , \68347 , \68348 , \68349 , \68350 , \68351 , \68352 ,
         \68353 , \68354 , \68355 , \68356 , \68357 , \68358 , \68359 , \68360 , \68361 , \68362 ,
         \68363 , \68364 , \68365 , \68366 , \68367 , \68368 , \68369 , \68370 , \68371 , \68372 ,
         \68373 , \68374 , \68375 , \68376 , \68377 , \68378 , \68379 , \68380 , \68381 , \68382 ,
         \68383 , \68384 , \68385 , \68386 , \68387 , \68388 , \68389 , \68390 , \68391 , \68392 ,
         \68393 , \68394 , \68395 , \68396 , \68397 , \68398 , \68399 , \68400 , \68401 , \68402 ,
         \68403 , \68404 , \68405 , \68406 , \68407 , \68408 , \68409 , \68410 , \68411 , \68412 ,
         \68413 , \68414 , \68415 , \68416 , \68417 , \68418 , \68419 , \68420 , \68421 , \68422 ,
         \68423 , \68424 , \68425 , \68426 , \68427 , \68428 , \68429 , \68430 , \68431 , \68432 ,
         \68433 , \68434 , \68435 , \68436 , \68437 , \68438 , \68439 , \68440 , \68441 , \68442 ,
         \68443 , \68444 , \68445 , \68446 , \68447 , \68448 , \68449 , \68450 , \68451 , \68452 ,
         \68453 , \68454 , \68455 , \68456 , \68457 , \68458 , \68459 , \68460 , \68461 , \68462 ,
         \68463 , \68464 , \68465 , \68466 , \68467 , \68468 , \68469 , \68470 , \68471 , \68472 ,
         \68473 , \68474 , \68475 , \68476 , \68477 , \68478 , \68479 , \68480 , \68481 , \68482 ,
         \68483 , \68484 , \68485 , \68486 , \68487 , \68488 , \68489 , \68490 , \68491 , \68492 ,
         \68493 , \68494 , \68495 , \68496 , \68497 , \68498 , \68499 , \68500 , \68501 , \68502 ,
         \68503 , \68504 , \68505 , \68506 , \68507 , \68508 , \68509 , \68510 , \68511 , \68512 ,
         \68513 , \68514 , \68515 , \68516 , \68517 , \68518 , \68519 , \68520 , \68521 , \68522 ,
         \68523 , \68524 , \68525 , \68526 , \68527 , \68528 , \68529 , \68530 , \68531 , \68532 ,
         \68533 , \68534 , \68535 , \68536 , \68537 , \68538 , \68539 , \68540 , \68541 , \68542 ,
         \68543 , \68544 , \68545 , \68546 , \68547 , \68548 , \68549 , \68550 , \68551 , \68552 ,
         \68553 , \68554 , \68555 , \68556 , \68557 , \68558 , \68559 , \68560 , \68561 , \68562 ,
         \68563 , \68564 , \68565 , \68566 , \68567 , \68568 , \68569 , \68570 , \68571 , \68572 ,
         \68573 , \68574 , \68575 , \68576 , \68577 , \68578 , \68579 , \68580 , \68581 , \68582 ,
         \68583 , \68584 , \68585 , \68586 , \68587 , \68588 , \68589 , \68590 , \68591 , \68592 ,
         \68593 , \68594 , \68595 , \68596 , \68597 , \68598 , \68599 , \68600 , \68601 , \68602 ,
         \68603 , \68604 , \68605 , \68606 , \68607 , \68608 , \68609 , \68610 , \68611 , \68612 ,
         \68613 , \68614 , \68615 , \68616 , \68617 , \68618 , \68619 , \68620 , \68621 , \68622 ,
         \68623 , \68624 , \68625 , \68626 , \68627 , \68628 , \68629 , \68630 , \68631 , \68632 ,
         \68633 , \68634 , \68635 , \68636 , \68637 , \68638 , \68639 , \68640 , \68641 , \68642 ,
         \68643 , \68644 , \68645 , \68646 , \68647 , \68648 , \68649 , \68650 , \68651 , \68652 ,
         \68653 , \68654 , \68655 , \68656 , \68657 , \68658 , \68659 , \68660 , \68661 , \68662 ,
         \68663 , \68664 , \68665 , \68666 , \68667 , \68668 , \68669 , \68670 , \68671 , \68672 ,
         \68673 , \68674 , \68675 , \68676 , \68677 , \68678 , \68679 , \68680 , \68681 , \68682 ,
         \68683 , \68684 , \68685 , \68686 , \68687 , \68688 , \68689 , \68690 , \68691 , \68692 ,
         \68693 , \68694 , \68695 , \68696 , \68697 , \68698 , \68699 , \68700 , \68701 , \68702 ,
         \68703 , \68704 , \68705 , \68706 , \68707 , \68708 , \68709 , \68710 , \68711 , \68712 ,
         \68713 , \68714 , \68715 , \68716 , \68717 , \68718 , \68719 , \68720 , \68721 , \68722 ,
         \68723 , \68724 , \68725 , \68726 , \68727 , \68728 , \68729 , \68730 , \68731 , \68732 ,
         \68733 , \68734 , \68735 , \68736 , \68737 , \68738 , \68739 , \68740 , \68741 , \68742 ,
         \68743 , \68744 , \68745 , \68746 , \68747 , \68748 , \68749 , \68750 , \68751 , \68752 ,
         \68753 , \68754 , \68755 , \68756 , \68757 , \68758 , \68759 , \68760 , \68761 , \68762 ,
         \68763 , \68764 , \68765 , \68766 , \68767 , \68768 , \68769 , \68770 , \68771 , \68772 ,
         \68773 , \68774 , \68775 , \68776 , \68777 , \68778 , \68779 , \68780 , \68781 , \68782 ,
         \68783 , \68784 , \68785 , \68786 , \68787 , \68788 , \68789 , \68790 , \68791 , \68792 ,
         \68793 , \68794 , \68795 , \68796 , \68797 , \68798 , \68799 , \68800 , \68801 , \68802 ,
         \68803 , \68804 , \68805 , \68806 , \68807 , \68808 , \68809 , \68810 , \68811 , \68812 ,
         \68813 , \68814 , \68815 , \68816 , \68817 , \68818 , \68819 , \68820 , \68821 , \68822 ,
         \68823 , \68824 , \68825 , \68826 , \68827 , \68828 , \68829 , \68830 , \68831 , \68832 ,
         \68833 , \68834 , \68835 , \68836 , \68837 , \68838 , \68839 , \68840 , \68841 , \68842 ,
         \68843 , \68844 , \68845 , \68846 , \68847 , \68848 , \68849 , \68850 , \68851 , \68852 ,
         \68853 , \68854 , \68855 , \68856 , \68857 , \68858 , \68859 , \68860 , \68861 , \68862 ,
         \68863 , \68864 , \68865 , \68866 , \68867 , \68868 , \68869 , \68870 , \68871 , \68872 ,
         \68873 , \68874 , \68875 , \68876 , \68877 , \68878 , \68879 , \68880 , \68881 , \68882 ,
         \68883 , \68884 , \68885 , \68886 , \68887 , \68888 , \68889 , \68890 , \68891 , \68892 ,
         \68893 , \68894 , \68895 , \68896 , \68897 , \68898 , \68899 , \68900 , \68901 , \68902 ,
         \68903 , \68904 , \68905 , \68906 , \68907 , \68908 , \68909 , \68910 , \68911 , \68912 ,
         \68913 , \68914 , \68915 , \68916 , \68917 , \68918 , \68919 , \68920 , \68921 , \68922 ,
         \68923 , \68924 , \68925 , \68926 , \68927 , \68928 , \68929 , \68930 , \68931 , \68932 ,
         \68933 , \68934 , \68935 , \68936 , \68937 , \68938 , \68939 , \68940 , \68941 , \68942 ,
         \68943 , \68944 , \68945 , \68946 , \68947 , \68948 , \68949 , \68950 , \68951 , \68952 ,
         \68953 , \68954 , \68955 , \68956 , \68957 , \68958 , \68959 , \68960 , \68961 , \68962 ,
         \68963 , \68964 , \68965 , \68966 , \68967 , \68968 , \68969 , \68970 , \68971 , \68972 ,
         \68973 , \68974 , \68975 , \68976 , \68977 , \68978 , \68979 , \68980 , \68981 , \68982 ,
         \68983 , \68984 , \68985 , \68986 , \68987 , \68988 , \68989 , \68990 , \68991 , \68992 ,
         \68993 , \68994 , \68995 , \68996 , \68997 , \68998 , \68999 , \69000 , \69001 , \69002 ,
         \69003 , \69004 , \69005 , \69006 , \69007 , \69008 , \69009 , \69010 , \69011 , \69012 ,
         \69013 , \69014 , \69015 , \69016 , \69017 , \69018 , \69019 , \69020 , \69021 , \69022 ,
         \69023 , \69024 , \69025 , \69026 , \69027 , \69028 , \69029 , \69030 , \69031 , \69032 ,
         \69033 , \69034 , \69035 , \69036 , \69037 , \69038 , \69039 , \69040 , \69041 , \69042 ,
         \69043 , \69044 , \69045 , \69046 , \69047 , \69048 , \69049 , \69050 , \69051 , \69052 ,
         \69053 , \69054 , \69055 , \69056 , \69057 , \69058 , \69059 , \69060 , \69061 , \69062 ,
         \69063 , \69064 , \69065 , \69066 , \69067 , \69068 , \69069 , \69070 , \69071 , \69072 ,
         \69073 , \69074 , \69075 , \69076 , \69077 , \69078 , \69079 , \69080 , \69081 , \69082 ,
         \69083 , \69084 , \69085 , \69086 , \69087 , \69088 , \69089 , \69090 , \69091 , \69092 ,
         \69093 , \69094 , \69095 , \69096 , \69097 , \69098 , \69099 , \69100 , \69101 , \69102 ,
         \69103 , \69104 , \69105 , \69106 , \69107 , \69108 , \69109 , \69110 , \69111 , \69112 ,
         \69113 , \69114 , \69115 , \69116 , \69117 , \69118 , \69119 , \69120 , \69121 , \69122 ,
         \69123 , \69124 , \69125 , \69126 , \69127 , \69128 , \69129 , \69130 , \69131 , \69132 ,
         \69133 , \69134 , \69135 , \69136 , \69137 , \69138 , \69139 , \69140 , \69141 , \69142 ,
         \69143 , \69144 , \69145 , \69146 , \69147 , \69148 , \69149 , \69150 , \69151 , \69152 ,
         \69153 , \69154 , \69155 , \69156 , \69157 , \69158 , \69159 , \69160 , \69161 , \69162 ,
         \69163 , \69164 , \69165 , \69166 , \69167 , \69168 , \69169 , \69170 , \69171 , \69172 ,
         \69173 , \69174 , \69175 , \69176 , \69177 , \69178 , \69179 , \69180 , \69181 , \69182 ,
         \69183 , \69184 , \69185 , \69186 , \69187 , \69188 , \69189 , \69190 , \69191 , \69192 ,
         \69193 , \69194 , \69195 , \69196 , \69197 , \69198 , \69199 , \69200 , \69201 , \69202 ,
         \69203 , \69204 , \69205 , \69206 , \69207 , \69208 , \69209 , \69210 , \69211 , \69212 ,
         \69213 , \69214 , \69215 , \69216 , \69217 , \69218 , \69219 , \69220 , \69221 , \69222 ,
         \69223 , \69224 , \69225 , \69226 , \69227 , \69228 , \69229 , \69230 , \69231 , \69232 ,
         \69233 , \69234 , \69235 , \69236 , \69237 , \69238 , \69239 , \69240 , \69241 , \69242 ,
         \69243 , \69244 , \69245 , \69246 , \69247 , \69248 , \69249 , \69250 , \69251 , \69252 ,
         \69253 , \69254 , \69255 , \69256 , \69257 , \69258 , \69259 , \69260 , \69261 , \69262 ,
         \69263 , \69264 , \69265 , \69266 , \69267 , \69268 , \69269 , \69270 , \69271 , \69272 ,
         \69273 , \69274 , \69275 , \69276 , \69277 , \69278 , \69279 , \69280 , \69281 , \69282 ,
         \69283 , \69284 , \69285 , \69286 , \69287 , \69288 , \69289 , \69290 , \69291 , \69292 ,
         \69293 , \69294 , \69295 , \69296 , \69297 , \69298 , \69299 , \69300 , \69301 , \69302 ,
         \69303 , \69304 , \69305 , \69306 , \69307 , \69308 , \69309 , \69310 , \69311 , \69312 ,
         \69313 , \69314 , \69315 , \69316 , \69317 , \69318 , \69319 , \69320 , \69321 , \69322 ,
         \69323 , \69324 , \69325 , \69326 , \69327 , \69328 , \69329 , \69330 , \69331 , \69332 ,
         \69333 , \69334 , \69335 , \69336 , \69337 , \69338 , \69339 , \69340 , \69341 , \69342 ,
         \69343 , \69344 , \69345 , \69346 , \69347 , \69348 , \69349 , \69350 , \69351 , \69352 ,
         \69353 , \69354 , \69355 , \69356 , \69357 , \69358 , \69359 , \69360 , \69361 , \69362 ,
         \69363 , \69364 , \69365 , \69366 , \69367 , \69368 , \69369 , \69370 , \69371 , \69372 ,
         \69373 , \69374 , \69375 , \69376 , \69377 , \69378 , \69379 , \69380 , \69381 , \69382 ,
         \69383 , \69384 , \69385 , \69386 , \69387 , \69388 , \69389 , \69390 , \69391 , \69392 ,
         \69393 , \69394 , \69395 , \69396 , \69397 , \69398 , \69399 , \69400 , \69401 , \69402 ,
         \69403 , \69404 , \69405 , \69406 , \69407 , \69408 , \69409 , \69410 , \69411 , \69412 ,
         \69413 , \69414 , \69415 , \69416 , \69417 , \69418 , \69419 , \69420 , \69421 , \69422 ,
         \69423 , \69424 , \69425 , \69426 , \69427 , \69428 , \69429 , \69430 , \69431 , \69432 ,
         \69433 , \69434 , \69435 , \69436 , \69437 , \69438 , \69439 , \69440 , \69441 , \69442 ,
         \69443 , \69444 , \69445 , \69446 , \69447 , \69448 , \69449 , \69450 , \69451 , \69452 ,
         \69453 , \69454 , \69455 , \69456 , \69457 , \69458 , \69459 , \69460 , \69461 , \69462 ,
         \69463 , \69464 , \69465 , \69466 , \69467 , \69468 , \69469 , \69470 , \69471 , \69472 ,
         \69473 , \69474 , \69475 , \69476 , \69477 , \69478 , \69479 , \69480 , \69481 , \69482 ,
         \69483 , \69484 , \69485 , \69486 , \69487 , \69488 , \69489 , \69490 , \69491 , \69492 ,
         \69493 , \69494 , \69495 , \69496 , \69497 , \69498 , \69499 , \69500 , \69501 , \69502 ,
         \69503 , \69504 , \69505 , \69506 , \69507 , \69508 , \69509 , \69510 , \69511 , \69512 ,
         \69513 , \69514 , \69515 , \69516 , \69517 , \69518 , \69519 , \69520 , \69521 , \69522 ,
         \69523 , \69524 , \69525 , \69526 , \69527 , \69528 , \69529 , \69530 , \69531 , \69532 ,
         \69533 , \69534 , \69535 , \69536 , \69537 , \69538 , \69539 , \69540 , \69541 , \69542 ,
         \69543 , \69544 , \69545 , \69546 , \69547 , \69548 , \69549 , \69550 , \69551 , \69552 ,
         \69553 , \69554 , \69555 , \69556 , \69557 , \69558 , \69559 , \69560 , \69561 , \69562 ,
         \69563 , \69564 , \69565 , \69566 , \69567 , \69568 , \69569 , \69570 , \69571 , \69572 ,
         \69573 , \69574 , \69575 , \69576 , \69577 , \69578 , \69579 , \69580 , \69581 , \69582 ,
         \69583 , \69584 , \69585 , \69586 , \69587 , \69588 , \69589 , \69590 , \69591 , \69592 ,
         \69593 , \69594 , \69595 , \69596 , \69597 , \69598 , \69599 , \69600 , \69601 , \69602 ,
         \69603 , \69604 , \69605 , \69606 , \69607 , \69608 , \69609 , \69610 , \69611 , \69612 ,
         \69613 , \69614 , \69615 , \69616 , \69617 , \69618 , \69619 , \69620 , \69621 , \69622 ,
         \69623 , \69624 , \69625 , \69626 , \69627 , \69628 , \69629 , \69630 , \69631 , \69632 ,
         \69633 , \69634 , \69635 , \69636 , \69637 , \69638 , \69639 , \69640 , \69641 , \69642 ,
         \69643 , \69644 , \69645 , \69646 , \69647 , \69648 , \69649 , \69650 , \69651 , \69652 ,
         \69653 , \69654 , \69655 , \69656 , \69657 , \69658 , \69659 , \69660 , \69661 , \69662 ,
         \69663 , \69664 , \69665 , \69666 , \69667 , \69668 , \69669 , \69670 , \69671 , \69672 ,
         \69673 , \69674 , \69675 , \69676 , \69677 , \69678 , \69679 , \69680 , \69681 , \69682 ,
         \69683 , \69684 , \69685 , \69686 , \69687 , \69688 , \69689 , \69690 , \69691 , \69692 ,
         \69693 , \69694 , \69695 , \69696 , \69697 , \69698 , \69699 , \69700 , \69701 , \69702 ,
         \69703 , \69704 , \69705 , \69706 , \69707 , \69708 , \69709 , \69710 , \69711 , \69712 ,
         \69713 , \69714 , \69715 , \69716 , \69717 , \69718 , \69719 , \69720 , \69721 , \69722 ,
         \69723 , \69724 , \69725 , \69726 , \69727 , \69728 , \69729 , \69730 , \69731 , \69732 ,
         \69733 , \69734 , \69735 , \69736 , \69737 , \69738 , \69739 , \69740 , \69741 , \69742 ,
         \69743 , \69744 , \69745 , \69746 , \69747 , \69748 , \69749 , \69750 , \69751 , \69752 ,
         \69753 , \69754 , \69755 , \69756 , \69757 , \69758 , \69759 , \69760 , \69761 , \69762 ,
         \69763 , \69764 , \69765 , \69766 , \69767 , \69768 , \69769 , \69770 , \69771 , \69772 ,
         \69773 , \69774 , \69775 , \69776 , \69777 , \69778 , \69779 , \69780 , \69781 , \69782 ,
         \69783 , \69784 , \69785 , \69786 , \69787 , \69788 , \69789 , \69790 , \69791 , \69792 ,
         \69793 , \69794 , \69795 , \69796 , \69797 , \69798 , \69799 , \69800 , \69801 , \69802 ,
         \69803 , \69804 , \69805 , \69806 , \69807 , \69808 , \69809 , \69810 , \69811 , \69812 ,
         \69813 , \69814 , \69815 , \69816 , \69817 , \69818 , \69819 , \69820 , \69821 , \69822 ,
         \69823 , \69824 , \69825 , \69826 , \69827 , \69828 , \69829 , \69830 , \69831 , \69832 ,
         \69833 , \69834 , \69835 , \69836 , \69837 , \69838 , \69839 , \69840 , \69841 , \69842 ,
         \69843 , \69844 , \69845 , \69846 , \69847 , \69848 , \69849 , \69850 , \69851 , \69852 ,
         \69853 , \69854 , \69855 , \69856 , \69857 , \69858 , \69859 , \69860 , \69861 , \69862 ,
         \69863 , \69864 , \69865 , \69866 , \69867 , \69868 , \69869 , \69870 , \69871 , \69872 ,
         \69873 , \69874 , \69875 , \69876 , \69877 , \69878 , \69879 , \69880 , \69881 , \69882 ,
         \69883 , \69884 , \69885 , \69886 , \69887 , \69888 , \69889 , \69890 , \69891 , \69892 ,
         \69893 , \69894 , \69895 , \69896 , \69897 , \69898 , \69899 , \69900 , \69901 , \69902 ,
         \69903 , \69904 , \69905 , \69906 , \69907 , \69908 , \69909 , \69910 , \69911 , \69912 ,
         \69913 , \69914 , \69915 , \69916 , \69917 , \69918 , \69919 , \69920 , \69921 , \69922 ,
         \69923 , \69924 , \69925 , \69926 , \69927 , \69928 , \69929 , \69930 , \69931 , \69932 ,
         \69933 , \69934 , \69935 , \69936 , \69937 , \69938 , \69939 , \69940 , \69941 , \69942 ,
         \69943 , \69944 , \69945 , \69946 , \69947 , \69948 , \69949 , \69950 , \69951 , \69952 ,
         \69953 , \69954 , \69955 , \69956 , \69957 , \69958 , \69959 , \69960 , \69961 , \69962 ,
         \69963 , \69964 , \69965 , \69966 , \69967 , \69968 , \69969 , \69970 , \69971 , \69972 ,
         \69973 , \69974 , \69975 , \69976 , \69977 , \69978 , \69979 , \69980 , \69981 , \69982 ,
         \69983 , \69984 , \69985 , \69986 , \69987 , \69988 , \69989 , \69990 , \69991 , \69992 ,
         \69993 , \69994 , \69995 , \69996 , \69997 , \69998 , \69999 , \70000 , \70001 , \70002 ,
         \70003 , \70004 , \70005 , \70006 , \70007 , \70008 , \70009 , \70010 , \70011 , \70012 ,
         \70013 , \70014 , \70015 , \70016 , \70017 , \70018 , \70019 , \70020 , \70021 , \70022 ,
         \70023 , \70024 , \70025 , \70026 , \70027 , \70028 , \70029 , \70030 , \70031 , \70032 ,
         \70033 , \70034 , \70035 , \70036 , \70037 , \70038 , \70039 , \70040 , \70041 , \70042 ,
         \70043 , \70044 , \70045 , \70046 , \70047 , \70048 , \70049 , \70050 , \70051 , \70052 ,
         \70053 , \70054 , \70055 , \70056 , \70057 , \70058 , \70059 , \70060 , \70061 , \70062 ,
         \70063 , \70064 , \70065 , \70066 , \70067 , \70068 , \70069 , \70070 , \70071 , \70072 ,
         \70073 , \70074 , \70075 , \70076 , \70077 , \70078 , \70079 , \70080 , \70081 , \70082 ,
         \70083 , \70084 , \70085 , \70086 , \70087 , \70088 , \70089 , \70090 , \70091 , \70092 ,
         \70093 , \70094 , \70095 , \70096 , \70097 , \70098 , \70099 , \70100 , \70101 , \70102 ,
         \70103 , \70104 , \70105 , \70106 , \70107 , \70108 , \70109 , \70110 , \70111 , \70112 ,
         \70113 , \70114 , \70115 , \70116 , \70117 , \70118 , \70119 , \70120 , \70121 , \70122 ,
         \70123 , \70124 , \70125 , \70126 , \70127 , \70128 , \70129 , \70130 , \70131 , \70132 ,
         \70133 , \70134 , \70135 , \70136 , \70137 , \70138 , \70139 , \70140 , \70141 , \70142 ,
         \70143 , \70144 , \70145 , \70146 , \70147 , \70148 , \70149 , \70150 , \70151 , \70152 ,
         \70153 , \70154 , \70155 , \70156 , \70157 , \70158 , \70159 , \70160 , \70161 , \70162 ,
         \70163 , \70164 , \70165 , \70166 , \70167 , \70168 , \70169 , \70170 , \70171 , \70172 ,
         \70173 , \70174 , \70175 , \70176 , \70177 , \70178 , \70179 , \70180 , \70181 , \70182 ,
         \70183 , \70184 , \70185 , \70186 , \70187 , \70188 , \70189 , \70190 , \70191 , \70192 ,
         \70193 , \70194 , \70195 , \70196 , \70197 , \70198 , \70199 , \70200 , \70201 , \70202 ,
         \70203 , \70204 , \70205 , \70206 , \70207 , \70208 , \70209 , \70210 , \70211 , \70212 ,
         \70213 , \70214 , \70215 , \70216 , \70217 , \70218 , \70219 , \70220 , \70221 , \70222 ,
         \70223 , \70224 , \70225 , \70226 , \70227 , \70228 , \70229 , \70230 , \70231 , \70232 ,
         \70233 , \70234 , \70235 , \70236 , \70237 , \70238 , \70239 , \70240 , \70241 , \70242 ,
         \70243 , \70244 , \70245 , \70246 , \70247 , \70248 , \70249 , \70250 , \70251 , \70252 ,
         \70253 , \70254 , \70255 , \70256 , \70257 , \70258 , \70259 , \70260 , \70261 , \70262 ,
         \70263 , \70264 , \70265 , \70266 , \70267 , \70268 , \70269 , \70270 , \70271 , \70272 ,
         \70273 , \70274 , \70275 , \70276 , \70277 , \70278 , \70279 , \70280 , \70281 , \70282 ,
         \70283 , \70284 , \70285 , \70286 , \70287 , \70288 , \70289 , \70290 , \70291 , \70292 ,
         \70293 , \70294 , \70295 , \70296 , \70297 , \70298 , \70299 , \70300 , \70301 , \70302 ,
         \70303 , \70304 , \70305 , \70306 , \70307 , \70308 , \70309 , \70310 , \70311 , \70312 ,
         \70313 , \70314 , \70315 , \70316 , \70317 , \70318 , \70319 , \70320 , \70321 , \70322 ,
         \70323 , \70324 , \70325 , \70326 , \70327 , \70328 , \70329 , \70330 , \70331 , \70332 ,
         \70333 , \70334 , \70335 , \70336 , \70337 , \70338 , \70339 , \70340 , \70341 , \70342 ,
         \70343 , \70344 , \70345 , \70346 , \70347 , \70348 , \70349 , \70350 , \70351 , \70352 ,
         \70353 , \70354 , \70355 , \70356 , \70357 , \70358 , \70359 , \70360 , \70361 , \70362 ,
         \70363 , \70364 , \70365 , \70366 , \70367 , \70368 , \70369 , \70370 , \70371 , \70372 ,
         \70373 , \70374 , \70375 , \70376 , \70377 , \70378 , \70379 , \70380 , \70381 , \70382 ,
         \70383 , \70384 , \70385 , \70386 , \70387 , \70388 , \70389 , \70390 , \70391 , \70392 ,
         \70393 , \70394 , \70395 , \70396 , \70397 , \70398 , \70399 , \70400 , \70401 , \70402 ,
         \70403 , \70404 , \70405 , \70406 , \70407 , \70408 , \70409 , \70410 , \70411 , \70412 ,
         \70413 , \70414 , \70415 , \70416 , \70417 , \70418 , \70419 , \70420 , \70421 , \70422 ,
         \70423 , \70424 , \70425 , \70426 , \70427 , \70428 , \70429 , \70430 , \70431 , \70432 ,
         \70433 , \70434 , \70435 , \70436 , \70437 , \70438 , \70439 , \70440 , \70441 , \70442 ,
         \70443 , \70444 , \70445 , \70446 , \70447 , \70448 , \70449 , \70450 , \70451 , \70452 ,
         \70453 , \70454 , \70455 , \70456 , \70457 , \70458 , \70459 , \70460 , \70461 , \70462 ,
         \70463 , \70464 , \70465 , \70466 , \70467 , \70468 , \70469 , \70470 , \70471 , \70472 ,
         \70473 , \70474 , \70475 , \70476 , \70477 , \70478 , \70479 , \70480 , \70481 , \70482 ,
         \70483 , \70484 , \70485 , \70486 , \70487 , \70488 , \70489 , \70490 , \70491 , \70492 ,
         \70493 , \70494 , \70495 , \70496 , \70497 , \70498 , \70499 , \70500 , \70501 , \70502 ,
         \70503 , \70504 , \70505 , \70506 , \70507 , \70508 , \70509 , \70510 , \70511 , \70512 ,
         \70513 , \70514 , \70515 , \70516 , \70517 , \70518 , \70519 , \70520 , \70521 , \70522 ,
         \70523 , \70524 , \70525 , \70526 , \70527 , \70528 , \70529 , \70530 , \70531 , \70532 ,
         \70533 , \70534 , \70535 , \70536 , \70537 , \70538 , \70539 , \70540 , \70541 , \70542 ,
         \70543 , \70544 , \70545 , \70546 , \70547 , \70548 , \70549 , \70550 , \70551 , \70552 ,
         \70553 , \70554 , \70555 , \70556 , \70557 , \70558 , \70559 , \70560 , \70561 , \70562 ,
         \70563 , \70564 , \70565 , \70566 , \70567 , \70568 , \70569 , \70570 , \70571 , \70572 ,
         \70573 , \70574 , \70575 , \70576 , \70577 , \70578 , \70579 , \70580 , \70581 , \70582 ,
         \70583 , \70584 , \70585 , \70586 , \70587 , \70588 , \70589 , \70590 , \70591 , \70592 ,
         \70593 , \70594 , \70595 , \70596 , \70597 , \70598 , \70599 , \70600 , \70601 , \70602 ,
         \70603 , \70604 , \70605 , \70606 , \70607 , \70608 , \70609 , \70610 , \70611 , \70612 ,
         \70613 , \70614 , \70615 , \70616 , \70617 , \70618 , \70619 , \70620 , \70621 , \70622 ,
         \70623 , \70624 , \70625 , \70626 , \70627 , \70628 , \70629 , \70630 , \70631 , \70632 ,
         \70633 , \70634 , \70635 , \70636 , \70637 , \70638 , \70639 , \70640 , \70641 , \70642 ,
         \70643 , \70644 , \70645 , \70646 , \70647 , \70648 , \70649 , \70650 , \70651 , \70652 ,
         \70653 , \70654 , \70655 , \70656 , \70657 , \70658 , \70659 , \70660 , \70661 , \70662 ,
         \70663 , \70664 , \70665 , \70666 , \70667 , \70668 , \70669 , \70670 , \70671 , \70672 ,
         \70673 , \70674 , \70675 , \70676 , \70677 , \70678 , \70679 , \70680 , \70681 , \70682 ,
         \70683 , \70684 , \70685 , \70686 , \70687 , \70688 , \70689 , \70690 , \70691 , \70692 ,
         \70693 , \70694 , \70695 , \70696 , \70697 , \70698 , \70699 , \70700 , \70701 , \70702 ,
         \70703 , \70704 , \70705 , \70706 , \70707 , \70708 , \70709 , \70710 , \70711 , \70712 ,
         \70713 , \70714 , \70715 , \70716 , \70717 , \70718 , \70719 , \70720 , \70721 , \70722 ,
         \70723 , \70724 , \70725 , \70726 , \70727 , \70728 , \70729 , \70730 , \70731 , \70732 ,
         \70733 , \70734 , \70735 , \70736 , \70737 , \70738 , \70739 , \70740 , \70741 , \70742 ,
         \70743 , \70744 , \70745 , \70746 , \70747 , \70748 , \70749 , \70750 , \70751 , \70752 ,
         \70753 , \70754 , \70755 , \70756 , \70757 , \70758 , \70759 , \70760 , \70761 , \70762 ,
         \70763 , \70764 , \70765 , \70766 , \70767 , \70768 , \70769 , \70770 , \70771 , \70772 ,
         \70773 , \70774 , \70775 , \70776 , \70777 , \70778 , \70779 , \70780 , \70781 , \70782 ,
         \70783 , \70784 , \70785 , \70786 , \70787 , \70788 , \70789 , \70790 , \70791 , \70792 ,
         \70793 , \70794 , \70795 , \70796 , \70797 , \70798 , \70799 , \70800 , \70801 , \70802 ,
         \70803 , \70804 , \70805 , \70806 , \70807 , \70808 , \70809 , \70810 , \70811 , \70812 ,
         \70813 , \70814 , \70815 , \70816 , \70817 , \70818 , \70819 , \70820 , \70821 , \70822 ,
         \70823 , \70824 , \70825 , \70826 , \70827 , \70828 , \70829 , \70830 , \70831 , \70832 ,
         \70833 , \70834 , \70835 , \70836 , \70837 , \70838 , \70839 , \70840 , \70841 , \70842 ,
         \70843 , \70844 , \70845 , \70846 , \70847 , \70848 , \70849 , \70850 , \70851 , \70852 ,
         \70853 , \70854 , \70855 , \70856 , \70857 , \70858 , \70859 , \70860 , \70861 , \70862 ,
         \70863 , \70864 , \70865 , \70866 , \70867 , \70868 , \70869 , \70870 , \70871 , \70872 ,
         \70873 , \70874 , \70875 , \70876 , \70877 , \70878 , \70879 , \70880 , \70881 , \70882 ,
         \70883 , \70884 , \70885 , \70886 , \70887 , \70888 , \70889 , \70890 , \70891 , \70892 ,
         \70893 , \70894 , \70895 , \70896 , \70897 , \70898 , \70899 , \70900 , \70901 , \70902 ,
         \70903 , \70904 , \70905 , \70906 , \70907 , \70908 , \70909 , \70910 , \70911 , \70912 ,
         \70913 , \70914 , \70915 , \70916 , \70917 , \70918 , \70919 , \70920 , \70921 , \70922 ,
         \70923 , \70924 , \70925 , \70926 , \70927 , \70928 , \70929 , \70930 , \70931 , \70932 ,
         \70933 , \70934 , \70935 , \70936 , \70937 , \70938 , \70939 , \70940 , \70941 , \70942 ,
         \70943 , \70944 , \70945 , \70946 , \70947 , \70948 , \70949 , \70950 , \70951 , \70952 ,
         \70953 , \70954 , \70955 , \70956 , \70957 , \70958 , \70959 , \70960 , \70961 , \70962 ,
         \70963 , \70964 , \70965 , \70966 , \70967 , \70968 , \70969 , \70970 , \70971 , \70972 ,
         \70973 , \70974 , \70975 , \70976 , \70977 , \70978 , \70979 , \70980 , \70981 , \70982 ,
         \70983 , \70984 , \70985 , \70986 , \70987 , \70988 , \70989 , \70990 , \70991 , \70992 ,
         \70993 , \70994 , \70995 , \70996 , \70997 , \70998 , \70999 , \71000 , \71001 , \71002 ,
         \71003 , \71004 , \71005 , \71006 , \71007 , \71008 , \71009 , \71010 , \71011 , \71012 ,
         \71013 , \71014 , \71015 , \71016 , \71017 , \71018 , \71019 , \71020 , \71021 , \71022 ,
         \71023 , \71024 , \71025 , \71026 , \71027 , \71028 , \71029 , \71030 , \71031 , \71032 ,
         \71033 , \71034 , \71035 , \71036 , \71037 , \71038 , \71039 , \71040 , \71041 , \71042 ,
         \71043 , \71044 , \71045 , \71046 , \71047 , \71048 , \71049 , \71050 , \71051 , \71052 ,
         \71053 , \71054 , \71055 , \71056 , \71057 , \71058 , \71059 , \71060 , \71061 , \71062 ,
         \71063 , \71064 , \71065 , \71066 , \71067 , \71068 , \71069 , \71070 , \71071 , \71072 ,
         \71073 , \71074 , \71075 , \71076 , \71077 , \71078 , \71079 , \71080 , \71081 , \71082 ,
         \71083 , \71084 , \71085 , \71086 , \71087 , \71088 , \71089 , \71090 , \71091 , \71092 ,
         \71093 , \71094 , \71095 , \71096 , \71097 , \71098 , \71099 , \71100 , \71101 , \71102 ,
         \71103 , \71104 , \71105 , \71106 , \71107 , \71108 , \71109 , \71110 , \71111 , \71112 ,
         \71113 , \71114 , \71115 , \71116 , \71117 , \71118 , \71119 , \71120 , \71121 , \71122 ,
         \71123 , \71124 , \71125 , \71126 , \71127 , \71128 , \71129 , \71130 , \71131 , \71132 ,
         \71133 , \71134 , \71135 , \71136 , \71137 , \71138 , \71139 , \71140 , \71141 , \71142 ,
         \71143 , \71144 , \71145 , \71146 , \71147 , \71148 , \71149 , \71150 , \71151 , \71152 ,
         \71153 , \71154 , \71155 , \71156 , \71157 , \71158 , \71159 , \71160 , \71161 , \71162 ,
         \71163 , \71164 , \71165 , \71166 , \71167 , \71168 , \71169 , \71170 , \71171 , \71172 ,
         \71173 , \71174 , \71175 , \71176 , \71177 , \71178 , \71179 , \71180 , \71181 , \71182 ,
         \71183 , \71184 , \71185 , \71186 , \71187 , \71188 , \71189 , \71190 , \71191 , \71192 ,
         \71193 , \71194 , \71195 , \71196 , \71197 , \71198 , \71199 , \71200 , \71201 , \71202 ,
         \71203 , \71204 , \71205 , \71206 , \71207 , \71208 , \71209 , \71210 , \71211 , \71212 ,
         \71213 , \71214 , \71215 , \71216 , \71217 , \71218 , \71219 , \71220 , \71221 , \71222 ,
         \71223 , \71224 , \71225 , \71226 , \71227 , \71228 , \71229 , \71230 , \71231 , \71232 ,
         \71233 , \71234 , \71235 , \71236 , \71237 , \71238 , \71239 , \71240 , \71241 , \71242 ,
         \71243 , \71244 , \71245 , \71246 , \71247 , \71248 , \71249 , \71250 , \71251 , \71252 ,
         \71253 , \71254 , \71255 , \71256 , \71257 , \71258 , \71259 , \71260 , \71261 , \71262 ,
         \71263 , \71264 , \71265 , \71266 , \71267 , \71268 , \71269 , \71270 , \71271 , \71272 ,
         \71273 , \71274 , \71275 , \71276 , \71277 , \71278 , \71279 , \71280 , \71281 , \71282 ,
         \71283 , \71284 , \71285 , \71286 , \71287 , \71288 , \71289 , \71290 , \71291 , \71292 ,
         \71293 , \71294 , \71295 , \71296 , \71297 , \71298 , \71299 , \71300 , \71301 , \71302 ,
         \71303 , \71304 , \71305 , \71306 , \71307 , \71308 , \71309 , \71310 , \71311 , \71312 ,
         \71313 , \71314 , \71315 , \71316 , \71317 , \71318 , \71319 , \71320 , \71321 , \71322 ,
         \71323 , \71324 , \71325 , \71326 , \71327 , \71328 , \71329 , \71330 , \71331 , \71332 ,
         \71333 , \71334 , \71335 , \71336 , \71337 , \71338 , \71339 , \71340 , \71341 , \71342 ,
         \71343 , \71344 , \71345 , \71346 , \71347 , \71348 , \71349 , \71350 , \71351 , \71352 ,
         \71353 , \71354 , \71355 , \71356 , \71357 , \71358 , \71359 , \71360 , \71361 , \71362 ,
         \71363 , \71364 , \71365 , \71366 , \71367 , \71368 , \71369 , \71370 , \71371 , \71372 ,
         \71373 , \71374 , \71375 , \71376 , \71377 , \71378 , \71379 , \71380 , \71381 , \71382 ,
         \71383 , \71384 , \71385 , \71386 , \71387 , \71388 , \71389 , \71390 , \71391 , \71392 ,
         \71393 , \71394 , \71395 , \71396 , \71397 , \71398 , \71399 , \71400 , \71401 , \71402 ,
         \71403 , \71404 , \71405 , \71406 , \71407 , \71408 , \71409 , \71410 , \71411 , \71412 ,
         \71413 , \71414 , \71415 , \71416 , \71417 , \71418 , \71419 , \71420 , \71421 , \71422 ,
         \71423 , \71424 , \71425 , \71426 , \71427 , \71428 , \71429 , \71430 , \71431 , \71432 ,
         \71433 , \71434 , \71435 , \71436 , \71437 , \71438 , \71439 , \71440 , \71441 , \71442 ,
         \71443 , \71444 , \71445 , \71446 , \71447 , \71448 , \71449 , \71450 , \71451 , \71452 ,
         \71453 , \71454 , \71455 , \71456 , \71457 , \71458 , \71459 , \71460 , \71461 , \71462 ,
         \71463 , \71464 , \71465 , \71466 , \71467 , \71468 , \71469 , \71470 , \71471 , \71472 ,
         \71473 , \71474 , \71475 , \71476 , \71477 , \71478 , \71479 , \71480 , \71481 , \71482 ,
         \71483 , \71484 , \71485 , \71486 , \71487 , \71488 , \71489 , \71490 , \71491 , \71492 ,
         \71493 , \71494 , \71495 , \71496 , \71497 , \71498 , \71499 , \71500 , \71501 , \71502 ,
         \71503 , \71504 , \71505 , \71506 , \71507 , \71508 , \71509 , \71510 , \71511 , \71512 ,
         \71513 , \71514 , \71515 , \71516 , \71517 , \71518 , \71519 , \71520 , \71521 , \71522 ,
         \71523 , \71524 , \71525 , \71526 , \71527 , \71528 , \71529 , \71530 , \71531 , \71532 ,
         \71533 , \71534 , \71535 , \71536 , \71537 , \71538 , \71539 , \71540 , \71541 , \71542 ,
         \71543 , \71544 , \71545 , \71546 , \71547 , \71548 , \71549 , \71550 , \71551 , \71552 ,
         \71553 , \71554 , \71555 , \71556 , \71557 , \71558 , \71559 , \71560 , \71561 , \71562 ,
         \71563 , \71564 , \71565 , \71566 , \71567 , \71568 , \71569 , \71570 , \71571 , \71572 ,
         \71573 , \71574 , \71575 , \71576 , \71577 , \71578 , \71579 , \71580 , \71581 , \71582 ,
         \71583 , \71584 , \71585 , \71586 , \71587 , \71588 , \71589 , \71590 , \71591 , \71592 ,
         \71593 , \71594 , \71595 , \71596 , \71597 , \71598 , \71599 , \71600 , \71601 , \71602 ,
         \71603 , \71604 , \71605 , \71606 , \71607 , \71608 , \71609 , \71610 , \71611 , \71612 ,
         \71613 , \71614 , \71615 , \71616 , \71617 , \71618 , \71619 , \71620 , \71621 , \71622 ,
         \71623 , \71624 , \71625 , \71626 , \71627 , \71628 , \71629 , \71630 , \71631 , \71632 ,
         \71633 , \71634 , \71635 , \71636 , \71637 , \71638 , \71639 , \71640 , \71641 , \71642 ,
         \71643 , \71644 , \71645 , \71646 , \71647 , \71648 , \71649 , \71650 , \71651 , \71652 ,
         \71653 , \71654 , \71655 , \71656 , \71657 , \71658 , \71659 , \71660 , \71661 , \71662 ,
         \71663 , \71664 , \71665 , \71666 , \71667 , \71668 , \71669 , \71670 , \71671 , \71672 ,
         \71673 , \71674 , \71675 , \71676 , \71677 , \71678 , \71679 , \71680 , \71681 , \71682 ,
         \71683 , \71684 , \71685 , \71686 , \71687 , \71688 , \71689 , \71690 , \71691 , \71692 ,
         \71693 , \71694 , \71695 , \71696 , \71697 , \71698 , \71699 , \71700 , \71701 , \71702 ,
         \71703 , \71704 , \71705 , \71706 , \71707 , \71708 , \71709 , \71710 , \71711 , \71712 ,
         \71713 , \71714 , \71715 , \71716 , \71717 , \71718 , \71719 , \71720 , \71721 , \71722 ,
         \71723 , \71724 , \71725 , \71726 , \71727 , \71728 , \71729 , \71730 , \71731 , \71732 ,
         \71733 , \71734 , \71735 , \71736 , \71737 , \71738 , \71739 , \71740 , \71741 , \71742 ,
         \71743 , \71744 , \71745 , \71746 , \71747 , \71748 , \71749 , \71750 , \71751 , \71752 ,
         \71753 , \71754 , \71755 , \71756 , \71757 , \71758 , \71759 , \71760 , \71761 , \71762 ,
         \71763 , \71764 , \71765 , \71766 , \71767 , \71768 , \71769 , \71770 , \71771 , \71772 ,
         \71773 , \71774 , \71775 , \71776 , \71777 , \71778 , \71779 , \71780 , \71781 , \71782 ,
         \71783 , \71784 , \71785 , \71786 , \71787 , \71788 , \71789 , \71790 , \71791 , \71792 ,
         \71793 , \71794 , \71795 , \71796 , \71797 , \71798 , \71799 , \71800 , \71801 , \71802 ,
         \71803 , \71804 , \71805 , \71806 , \71807 , \71808 , \71809 , \71810 , \71811 , \71812 ,
         \71813 , \71814 , \71815 , \71816 , \71817 , \71818 , \71819 , \71820 , \71821 , \71822 ,
         \71823 , \71824 , \71825 , \71826 , \71827 , \71828 , \71829 , \71830 , \71831 , \71832 ,
         \71833 , \71834 , \71835 , \71836 , \71837 , \71838 , \71839 , \71840 , \71841 , \71842 ,
         \71843 , \71844 , \71845 , \71846 , \71847 , \71848 , \71849 , \71850 , \71851 , \71852 ,
         \71853 , \71854 , \71855 , \71856 , \71857 , \71858 , \71859 , \71860 , \71861 , \71862 ,
         \71863 , \71864 , \71865 , \71866 , \71867 , \71868 , \71869 , \71870 , \71871 , \71872 ,
         \71873 , \71874 , \71875 , \71876 , \71877 , \71878 , \71879 , \71880 , \71881 , \71882 ,
         \71883 , \71884 , \71885 , \71886 , \71887 , \71888 , \71889 , \71890 , \71891 , \71892 ,
         \71893 , \71894 , \71895 , \71896 , \71897 , \71898 , \71899 , \71900 , \71901 , \71902 ,
         \71903 , \71904 , \71905 , \71906 , \71907 , \71908 , \71909 , \71910 , \71911 , \71912 ,
         \71913 , \71914 , \71915 , \71916 , \71917 , \71918 , \71919 , \71920 , \71921 , \71922 ,
         \71923 , \71924 , \71925 , \71926 , \71927 , \71928 , \71929 , \71930 , \71931 , \71932 ,
         \71933 , \71934 , \71935 , \71936 , \71937 , \71938 , \71939 , \71940 , \71941 , \71942 ,
         \71943 , \71944 , \71945 , \71946 , \71947 , \71948 , \71949 , \71950 , \71951 , \71952 ,
         \71953 , \71954 , \71955 , \71956 , \71957 , \71958 , \71959 , \71960 , \71961 , \71962 ,
         \71963 , \71964 , \71965 , \71966 , \71967 , \71968 , \71969 , \71970 , \71971 , \71972 ,
         \71973 , \71974 , \71975 , \71976 , \71977 , \71978 , \71979 , \71980 , \71981 , \71982 ,
         \71983 , \71984 , \71985 , \71986 , \71987 , \71988 , \71989 , \71990 , \71991 , \71992 ,
         \71993 , \71994 , \71995 , \71996 , \71997 , \71998 , \71999 , \72000 , \72001 , \72002 ,
         \72003 , \72004 , \72005 , \72006 , \72007 , \72008 , \72009 , \72010 , \72011 , \72012 ,
         \72013 , \72014 , \72015 , \72016 , \72017 , \72018 , \72019 , \72020 , \72021 , \72022 ,
         \72023 , \72024 , \72025 , \72026 , \72027 , \72028 , \72029 , \72030 , \72031 , \72032 ,
         \72033 , \72034 , \72035 , \72036 , \72037 , \72038 , \72039 , \72040 , \72041 , \72042 ,
         \72043 , \72044 , \72045 , \72046 , \72047 , \72048 , \72049 , \72050 , \72051 , \72052 ,
         \72053 , \72054 , \72055 , \72056 , \72057 , \72058 , \72059 , \72060 , \72061 , \72062 ,
         \72063 , \72064 , \72065 , \72066 , \72067 , \72068 , \72069 , \72070 , \72071 , \72072 ,
         \72073 , \72074 , \72075 , \72076 , \72077 , \72078 , \72079 , \72080 , \72081 , \72082 ,
         \72083 , \72084 , \72085 , \72086 , \72087 , \72088 , \72089 , \72090 , \72091 , \72092 ,
         \72093 , \72094 , \72095 , \72096 , \72097 , \72098 , \72099 , \72100 , \72101 , \72102 ,
         \72103 , \72104 , \72105 , \72106 , \72107 , \72108 , \72109 , \72110 , \72111 , \72112 ,
         \72113 , \72114 , \72115 , \72116 , \72117 , \72118 , \72119 , \72120 , \72121 , \72122 ,
         \72123 , \72124 , \72125 , \72126 , \72127 , \72128 , \72129 , \72130 , \72131 , \72132 ,
         \72133 , \72134 , \72135 , \72136 , \72137 , \72138 , \72139 , \72140 , \72141 , \72142 ,
         \72143 , \72144 , \72145 , \72146 , \72147 , \72148 , \72149 , \72150 , \72151 , \72152 ,
         \72153 , \72154 , \72155 , \72156 , \72157 , \72158 , \72159 , \72160 , \72161 , \72162 ,
         \72163 , \72164 , \72165 , \72166 , \72167 , \72168 , \72169 , \72170 , \72171 , \72172 ,
         \72173 , \72174 , \72175 , \72176 , \72177 , \72178 , \72179 , \72180 , \72181 , \72182 ,
         \72183 , \72184 , \72185 , \72186 , \72187 , \72188 , \72189 , \72190 , \72191 , \72192 ,
         \72193 , \72194 , \72195 , \72196 , \72197 , \72198 , \72199 , \72200 , \72201 , \72202 ,
         \72203 , \72204 , \72205 , \72206 , \72207 , \72208 , \72209 , \72210 , \72211 , \72212 ,
         \72213 , \72214 , \72215 , \72216 , \72217 , \72218 , \72219 , \72220 , \72221 , \72222 ,
         \72223 , \72224 , \72225 , \72226 , \72227 , \72228 , \72229 , \72230 , \72231 , \72232 ,
         \72233 , \72234 , \72235 , \72236 , \72237 , \72238 , \72239 , \72240 , \72241 , \72242 ,
         \72243 , \72244 , \72245 , \72246 , \72247 , \72248 , \72249 , \72250 , \72251 , \72252 ,
         \72253 , \72254 , \72255 , \72256 , \72257 , \72258 , \72259 , \72260 , \72261 , \72262 ,
         \72263 , \72264 , \72265 , \72266 , \72267 , \72268 , \72269 , \72270 , \72271 , \72272 ,
         \72273 , \72274 , \72275 , \72276 , \72277 , \72278 , \72279 , \72280 , \72281 , \72282 ,
         \72283 , \72284 , \72285 , \72286 , \72287 , \72288 , \72289 , \72290 , \72291 , \72292 ,
         \72293 , \72294 , \72295 , \72296 , \72297 , \72298 , \72299 , \72300 , \72301 , \72302 ,
         \72303 , \72304 , \72305 , \72306 , \72307 , \72308 , \72309 , \72310 , \72311 , \72312 ,
         \72313 , \72314 , \72315 , \72316 , \72317 , \72318 , \72319 , \72320 , \72321 , \72322 ,
         \72323 , \72324 , \72325 , \72326 , \72327 , \72328 , \72329 , \72330 , \72331 , \72332 ,
         \72333 , \72334 , \72335 , \72336 , \72337 , \72338 , \72339 , \72340 , \72341 , \72342 ,
         \72343 , \72344 , \72345 , \72346 , \72347 , \72348 , \72349 , \72350 , \72351 , \72352 ,
         \72353 , \72354 , \72355 , \72356 , \72357 , \72358 , \72359 , \72360 , \72361 , \72362 ,
         \72363 , \72364 , \72365 , \72366 , \72367 , \72368 , \72369 , \72370 , \72371 , \72372 ,
         \72373 , \72374 , \72375 , \72376 , \72377 , \72378 , \72379 , \72380 , \72381 , \72382 ,
         \72383 , \72384 , \72385 , \72386 , \72387 , \72388 , \72389 , \72390 , \72391 , \72392 ,
         \72393 , \72394 , \72395 , \72396 , \72397 , \72398 , \72399 , \72400 , \72401 , \72402 ,
         \72403 , \72404 , \72405 , \72406 , \72407 , \72408 , \72409 , \72410 , \72411 , \72412 ,
         \72413 , \72414 , \72415 , \72416 , \72417 , \72418 , \72419 , \72420 , \72421 , \72422 ,
         \72423 , \72424 , \72425 , \72426 , \72427 , \72428 , \72429 , \72430 , \72431 , \72432 ,
         \72433 , \72434 , \72435 , \72436 , \72437 , \72438 , \72439 , \72440 , \72441 , \72442 ,
         \72443 , \72444 , \72445 , \72446 , \72447 , \72448 , \72449 , \72450 , \72451 , \72452 ,
         \72453 , \72454 , \72455 , \72456 , \72457 , \72458 , \72459 , \72460 , \72461 , \72462 ,
         \72463 , \72464 , \72465 , \72466 , \72467 , \72468 , \72469 , \72470 , \72471 , \72472 ,
         \72473 , \72474 , \72475 , \72476 , \72477 , \72478 , \72479 , \72480 , \72481 , \72482 ,
         \72483 , \72484 , \72485 , \72486 , \72487 , \72488 , \72489 , \72490 , \72491 , \72492 ,
         \72493 , \72494 , \72495 , \72496 , \72497 , \72498 , \72499 , \72500 , \72501 , \72502 ,
         \72503 , \72504 , \72505 , \72506 , \72507 , \72508 , \72509 , \72510 , \72511 , \72512 ,
         \72513 , \72514 , \72515 , \72516 , \72517 , \72518 , \72519 , \72520 , \72521 , \72522 ,
         \72523 , \72524 , \72525 , \72526 , \72527 , \72528 , \72529 , \72530 , \72531 , \72532 ,
         \72533 , \72534 , \72535 , \72536 , \72537 , \72538 , \72539 , \72540 , \72541 , \72542 ,
         \72543 , \72544 , \72545 , \72546 , \72547 , \72548 , \72549 , \72550 , \72551 , \72552 ,
         \72553 , \72554 , \72555 , \72556 , \72557 , \72558 , \72559 , \72560 , \72561 , \72562 ,
         \72563 , \72564 , \72565 , \72566 , \72567 , \72568 , \72569 , \72570 , \72571 , \72572 ,
         \72573 , \72574 , \72575 , \72576 , \72577 , \72578 , \72579 , \72580 , \72581 , \72582 ,
         \72583 , \72584 , \72585 , \72586 , \72587 , \72588 , \72589 , \72590 , \72591 , \72592 ,
         \72593 , \72594 , \72595 , \72596 , \72597 , \72598 , \72599 , \72600 , \72601 , \72602 ,
         \72603 , \72604 , \72605 , \72606 , \72607 , \72608 , \72609 , \72610 , \72611 , \72612 ,
         \72613 , \72614 , \72615 , \72616 , \72617 , \72618 , \72619 , \72620 , \72621 , \72622 ,
         \72623 , \72624 , \72625 , \72626 , \72627 , \72628 , \72629 , \72630 , \72631 , \72632 ,
         \72633 , \72634 , \72635 , \72636 , \72637 , \72638 , \72639 , \72640 , \72641 , \72642 ,
         \72643 , \72644 , \72645 , \72646 , \72647 , \72648 , \72649 , \72650 , \72651 , \72652 ,
         \72653 , \72654 , \72655 , \72656 , \72657 , \72658 , \72659 , \72660 , \72661 , \72662 ,
         \72663 , \72664 , \72665 , \72666 , \72667 , \72668 , \72669 , \72670 , \72671 , \72672 ,
         \72673 , \72674 , \72675 , \72676 , \72677 , \72678 , \72679 , \72680 , \72681 , \72682 ,
         \72683 , \72684 , \72685 , \72686 , \72687 , \72688 , \72689 , \72690 , \72691 , \72692 ,
         \72693 , \72694 , \72695 , \72696 , \72697 , \72698 , \72699 , \72700 , \72701 , \72702 ,
         \72703 , \72704 , \72705 , \72706 , \72707 , \72708 , \72709 , \72710 , \72711 , \72712 ,
         \72713 , \72714 , \72715 , \72716 , \72717 , \72718 , \72719 , \72720 , \72721 , \72722 ,
         \72723 , \72724 , \72725 , \72726 , \72727 , \72728 , \72729 , \72730 , \72731 , \72732 ,
         \72733 , \72734 , \72735 , \72736 , \72737 , \72738 , \72739 , \72740 , \72741 , \72742 ,
         \72743 , \72744 , \72745 , \72746 , \72747 , \72748 , \72749 , \72750 , \72751 , \72752 ,
         \72753 , \72754 , \72755 , \72756 , \72757 , \72758 , \72759 , \72760 , \72761 , \72762 ,
         \72763 , \72764 , \72765 , \72766 , \72767 , \72768 , \72769 , \72770 , \72771 , \72772 ,
         \72773 , \72774 , \72775 , \72776 , \72777 , \72778 , \72779 , \72780 , \72781 , \72782 ,
         \72783 , \72784 , \72785 , \72786 , \72787 , \72788 , \72789 , \72790 , \72791 , \72792 ,
         \72793 , \72794 , \72795 , \72796 , \72797 , \72798 , \72799 , \72800 , \72801 , \72802 ,
         \72803 , \72804 , \72805 , \72806 , \72807 , \72808 , \72809 , \72810 , \72811 , \72812 ,
         \72813 , \72814 , \72815 , \72816 , \72817 , \72818 , \72819 , \72820 , \72821 , \72822 ,
         \72823 , \72824 , \72825 , \72826 , \72827 , \72828 , \72829 , \72830 , \72831 , \72832 ,
         \72833 , \72834 , \72835 , \72836 , \72837 , \72838 , \72839 , \72840 , \72841 , \72842 ,
         \72843 , \72844 , \72845 , \72846 , \72847 , \72848 , \72849 , \72850 , \72851 , \72852 ,
         \72853 , \72854 , \72855 , \72856 , \72857 , \72858 , \72859 , \72860 , \72861 , \72862 ,
         \72863 , \72864 , \72865 , \72866 , \72867 , \72868 , \72869 , \72870 , \72871 , \72872 ,
         \72873 , \72874 , \72875 , \72876 , \72877 , \72878 , \72879 , \72880 , \72881 , \72882 ,
         \72883 , \72884 , \72885 , \72886 , \72887 , \72888 , \72889 , \72890 , \72891 , \72892 ,
         \72893 , \72894 , \72895 , \72896 , \72897 , \72898 , \72899 , \72900 , \72901 , \72902 ,
         \72903 , \72904 , \72905 , \72906 , \72907 , \72908 , \72909 , \72910 , \72911 , \72912 ,
         \72913 , \72914 , \72915 , \72916 , \72917 , \72918 , \72919 , \72920 , \72921 , \72922 ,
         \72923 , \72924 , \72925 , \72926 , \72927 , \72928 , \72929 , \72930 , \72931 , \72932 ,
         \72933 , \72934 , \72935 , \72936 , \72937 , \72938 , \72939 , \72940 , \72941 , \72942 ,
         \72943 , \72944 , \72945 , \72946 , \72947 , \72948 , \72949 , \72950 , \72951 , \72952 ,
         \72953 , \72954 , \72955 , \72956 , \72957 , \72958 , \72959 , \72960 , \72961 , \72962 ,
         \72963 , \72964 , \72965 , \72966 , \72967 , \72968 , \72969 , \72970 , \72971 , \72972 ,
         \72973 , \72974 , \72975 , \72976 , \72977 , \72978 , \72979 , \72980 , \72981 , \72982 ,
         \72983 , \72984 , \72985 , \72986 , \72987 , \72988 , \72989 , \72990 , \72991 , \72992 ,
         \72993 , \72994 , \72995 , \72996 , \72997 , \72998 , \72999 , \73000 , \73001 , \73002 ,
         \73003 , \73004 , \73005 , \73006 , \73007 , \73008 , \73009 , \73010 , \73011 , \73012 ,
         \73013 , \73014 , \73015 , \73016 , \73017 , \73018 , \73019 , \73020 , \73021 , \73022 ,
         \73023 , \73024 , \73025 , \73026 , \73027 , \73028 , \73029 , \73030 , \73031 , \73032 ,
         \73033 , \73034 , \73035 , \73036 , \73037 , \73038 , \73039 , \73040 , \73041 , \73042 ,
         \73043 , \73044 , \73045 , \73046 , \73047 , \73048 , \73049 , \73050 , \73051 , \73052 ,
         \73053 , \73054 , \73055 , \73056 , \73057 , \73058 , \73059 , \73060 , \73061 , \73062 ,
         \73063 , \73064 , \73065 , \73066 , \73067 , \73068 , \73069 , \73070 , \73071 , \73072 ,
         \73073 , \73074 , \73075 , \73076 , \73077 , \73078 , \73079 , \73080 , \73081 , \73082 ,
         \73083 , \73084 , \73085 , \73086 , \73087 , \73088 , \73089 , \73090 , \73091 , \73092 ,
         \73093 , \73094 , \73095 , \73096 , \73097 , \73098 , \73099 , \73100 , \73101 , \73102 ,
         \73103 , \73104 , \73105 , \73106 , \73107 , \73108 , \73109 , \73110 , \73111 , \73112 ,
         \73113 , \73114 , \73115 , \73116 , \73117 , \73118 , \73119 , \73120 , \73121 , \73122 ,
         \73123 , \73124 , \73125 , \73126 , \73127 , \73128 , \73129 , \73130 , \73131 , \73132 ,
         \73133 , \73134 , \73135 , \73136 , \73137 , \73138 , \73139 , \73140 , \73141 , \73142 ,
         \73143 , \73144 , \73145 , \73146 , \73147 , \73148 , \73149 , \73150 , \73151 , \73152 ,
         \73153 , \73154 , \73155 , \73156 , \73157 , \73158 , \73159 , \73160 , \73161 , \73162 ,
         \73163 , \73164 , \73165 , \73166 , \73167 , \73168 , \73169 , \73170 , \73171 , \73172 ,
         \73173 , \73174 , \73175 , \73176 , \73177 , \73178 , \73179 , \73180 , \73181 , \73182 ,
         \73183 , \73184 , \73185 , \73186 , \73187 , \73188 , \73189 , \73190 , \73191 , \73192 ,
         \73193 , \73194 , \73195 , \73196 , \73197 , \73198 , \73199 , \73200 , \73201 , \73202 ,
         \73203 , \73204 , \73205 , \73206 , \73207 , \73208 , \73209 , \73210 , \73211 , \73212 ,
         \73213 , \73214 , \73215 , \73216 , \73217 , \73218 , \73219 , \73220 , \73221 , \73222 ,
         \73223 , \73224 , \73225 , \73226 , \73227 , \73228 , \73229 , \73230 , \73231 , \73232 ,
         \73233 , \73234 , \73235 , \73236 , \73237 , \73238 , \73239 , \73240 , \73241 , \73242 ,
         \73243 , \73244 , \73245 , \73246 , \73247 , \73248 , \73249 , \73250 , \73251 , \73252 ,
         \73253 , \73254 , \73255 , \73256 , \73257 , \73258 , \73259 , \73260 , \73261 , \73262 ,
         \73263 , \73264 , \73265 , \73266 , \73267 , \73268 , \73269 , \73270 , \73271 , \73272 ,
         \73273 , \73274 , \73275 , \73276 , \73277 , \73278 , \73279 , \73280 , \73281 , \73282 ,
         \73283 , \73284 , \73285 , \73286 , \73287 , \73288 , \73289 , \73290 , \73291 , \73292 ,
         \73293 , \73294 , \73295 , \73296 , \73297 , \73298 , \73299 , \73300 , \73301 , \73302 ,
         \73303 , \73304 , \73305 , \73306 , \73307 , \73308 , \73309 , \73310 , \73311 , \73312 ,
         \73313 , \73314 , \73315 , \73316 , \73317 , \73318 , \73319 , \73320 , \73321 , \73322 ,
         \73323 , \73324 , \73325 , \73326 , \73327 , \73328 , \73329 , \73330 , \73331 , \73332 ,
         \73333 , \73334 , \73335 , \73336 , \73337 , \73338 , \73339 , \73340 , \73341 , \73342 ,
         \73343 , \73344 , \73345 , \73346 , \73347 , \73348 , \73349 , \73350 , \73351 , \73352 ,
         \73353 , \73354 , \73355 , \73356 , \73357 , \73358 , \73359 , \73360 , \73361 , \73362 ,
         \73363 , \73364 , \73365 , \73366 , \73367 , \73368 , \73369 , \73370 , \73371 , \73372 ,
         \73373 , \73374 , \73375 , \73376 , \73377 , \73378 , \73379 , \73380 , \73381 , \73382 ,
         \73383 , \73384 , \73385 , \73386 , \73387 , \73388 , \73389 , \73390 , \73391 , \73392 ,
         \73393 , \73394 , \73395 , \73396 , \73397 , \73398 , \73399 , \73400 , \73401 , \73402 ,
         \73403 , \73404 , \73405 , \73406 , \73407 , \73408 , \73409 , \73410 , \73411 , \73412 ,
         \73413 , \73414 , \73415 , \73416 , \73417 , \73418 , \73419 , \73420 , \73421 , \73422 ,
         \73423 , \73424 , \73425 , \73426 , \73427 , \73428 , \73429 , \73430 , \73431 , \73432 ,
         \73433 , \73434 , \73435 , \73436 , \73437 , \73438 , \73439 , \73440 , \73441 , \73442 ,
         \73443 , \73444 , \73445 , \73446 , \73447 , \73448 , \73449 , \73450 , \73451 , \73452 ,
         \73453 , \73454 , \73455 , \73456 , \73457 , \73458 , \73459 , \73460 , \73461 , \73462 ,
         \73463 , \73464 , \73465 , \73466 , \73467 , \73468 , \73469 , \73470 , \73471 , \73472 ,
         \73473 , \73474 , \73475 , \73476 , \73477 , \73478 , \73479 , \73480 , \73481 , \73482 ,
         \73483 , \73484 , \73485 , \73486 , \73487 , \73488 , \73489 , \73490 , \73491 , \73492 ,
         \73493 , \73494 , \73495 , \73496 , \73497 , \73498 , \73499 , \73500 , \73501 , \73502 ,
         \73503 , \73504 , \73505 , \73506 , \73507 , \73508 , \73509 , \73510 , \73511 , \73512 ,
         \73513 , \73514 , \73515 , \73516 , \73517 , \73518 , \73519 , \73520 , \73521 , \73522 ,
         \73523 , \73524 , \73525 , \73526 , \73527 , \73528 , \73529 , \73530 , \73531 , \73532 ,
         \73533 , \73534 , \73535 , \73536 , \73537 , \73538 , \73539 , \73540 , \73541 , \73542 ,
         \73543 , \73544 , \73545 , \73546 , \73547 , \73548 , \73549 , \73550 , \73551 , \73552 ,
         \73553 , \73554 , \73555 , \73556 , \73557 , \73558 , \73559 , \73560 , \73561 , \73562 ,
         \73563 , \73564 , \73565 , \73566 , \73567 , \73568 , \73569 , \73570 , \73571 , \73572 ,
         \73573 , \73574 , \73575 , \73576 , \73577 , \73578 , \73579 , \73580 , \73581 , \73582 ,
         \73583 , \73584 , \73585 , \73586 , \73587 , \73588 , \73589 , \73590 , \73591 , \73592 ,
         \73593 , \73594 , \73595 , \73596 , \73597 , \73598 , \73599 , \73600 , \73601 , \73602 ,
         \73603 , \73604 , \73605 , \73606 , \73607 , \73608 , \73609 , \73610 , \73611 , \73612 ,
         \73613 , \73614 , \73615 , \73616 , \73617 , \73618 , \73619 , \73620 , \73621 , \73622 ,
         \73623 , \73624 , \73625 , \73626 , \73627 , \73628 , \73629 , \73630 , \73631 , \73632 ,
         \73633 , \73634 , \73635 , \73636 , \73637 , \73638 , \73639 , \73640 , \73641 , \73642 ,
         \73643 , \73644 , \73645 , \73646 , \73647 , \73648 , \73649 , \73650 , \73651 , \73652 ,
         \73653 , \73654 , \73655 , \73656 , \73657 , \73658 , \73659 , \73660 , \73661 , \73662 ,
         \73663 , \73664 , \73665 , \73666 , \73667 , \73668 , \73669 , \73670 , \73671 , \73672 ,
         \73673 , \73674 , \73675 , \73676 , \73677 , \73678 , \73679 , \73680 , \73681 , \73682 ,
         \73683 , \73684 , \73685 , \73686 , \73687 , \73688 , \73689 , \73690 , \73691 , \73692 ,
         \73693 , \73694 , \73695 , \73696 , \73697 , \73698 , \73699 , \73700 , \73701 , \73702 ,
         \73703 , \73704 , \73705 , \73706 , \73707 , \73708 , \73709 , \73710 , \73711 , \73712 ,
         \73713 , \73714 , \73715 , \73716 , \73717 , \73718 , \73719 , \73720 , \73721 , \73722 ,
         \73723 , \73724 , \73725 , \73726 , \73727 , \73728 , \73729 , \73730 , \73731 , \73732 ,
         \73733 , \73734 , \73735 , \73736 , \73737 , \73738 , \73739 , \73740 , \73741 , \73742 ,
         \73743 , \73744 , \73745 , \73746 , \73747 , \73748 , \73749 , \73750 , \73751 , \73752 ,
         \73753 , \73754 , \73755 , \73756 , \73757 , \73758 , \73759 , \73760 , \73761 , \73762 ,
         \73763 , \73764 , \73765 , \73766 , \73767 , \73768 , \73769 , \73770 , \73771 , \73772 ,
         \73773 , \73774 , \73775 , \73776 , \73777 , \73778 , \73779 , \73780 , \73781 , \73782 ,
         \73783 , \73784 , \73785 , \73786 , \73787 , \73788 , \73789 , \73790 , \73791 , \73792 ,
         \73793 , \73794 , \73795 , \73796 , \73797 , \73798 , \73799 , \73800 , \73801 , \73802 ,
         \73803 , \73804 , \73805 , \73806 , \73807 , \73808 , \73809 , \73810 , \73811 , \73812 ,
         \73813 , \73814 , \73815 , \73816 , \73817 , \73818 , \73819 , \73820 , \73821 , \73822 ,
         \73823 , \73824 , \73825 , \73826 , \73827 , \73828 , \73829 , \73830 , \73831 , \73832 ,
         \73833 , \73834 , \73835 , \73836 , \73837 , \73838 , \73839 , \73840 , \73841 , \73842 ,
         \73843 , \73844 , \73845 , \73846 , \73847 , \73848 , \73849 , \73850 , \73851 , \73852 ,
         \73853 , \73854 , \73855 , \73856 , \73857 , \73858 , \73859 , \73860 , \73861 , \73862 ,
         \73863 , \73864 , \73865 , \73866 , \73867 , \73868 , \73869 , \73870 , \73871 , \73872 ,
         \73873 , \73874 , \73875 , \73876 , \73877 , \73878 , \73879 , \73880 , \73881 , \73882 ,
         \73883 , \73884 , \73885 , \73886 , \73887 , \73888 , \73889 , \73890 , \73891 , \73892 ,
         \73893 , \73894 , \73895 , \73896 , \73897 , \73898 , \73899 , \73900 , \73901 , \73902 ,
         \73903 , \73904 , \73905 , \73906 , \73907 , \73908 , \73909 , \73910 , \73911 , \73912 ,
         \73913 , \73914 , \73915 , \73916 , \73917 , \73918 , \73919 , \73920 , \73921 , \73922 ,
         \73923 , \73924 , \73925 , \73926 , \73927 , \73928 , \73929 , \73930 , \73931 , \73932 ,
         \73933 , \73934 , \73935 , \73936 , \73937 , \73938 , \73939 , \73940 , \73941 , \73942 ,
         \73943 , \73944 , \73945 , \73946 , \73947 , \73948 , \73949 , \73950 , \73951 , \73952 ,
         \73953 , \73954 , \73955 , \73956 , \73957 , \73958 , \73959 , \73960 , \73961 , \73962 ,
         \73963 , \73964 , \73965 , \73966 , \73967 , \73968 , \73969 , \73970 , \73971 , \73972 ,
         \73973 , \73974 , \73975 , \73976 , \73977 , \73978 , \73979 , \73980 , \73981 , \73982 ,
         \73983 , \73984 , \73985 , \73986 , \73987 , \73988 , \73989 , \73990 , \73991 , \73992 ,
         \73993 , \73994 , \73995 , \73996 , \73997 , \73998 , \73999 , \74000 , \74001 , \74002 ,
         \74003 , \74004 , \74005 , \74006 , \74007 , \74008 , \74009 , \74010 , \74011 , \74012 ,
         \74013 , \74014 , \74015 , \74016 , \74017 , \74018 , \74019 , \74020 , \74021 , \74022 ,
         \74023 , \74024 , \74025 , \74026 , \74027 , \74028 , \74029 , \74030 , \74031 , \74032 ,
         \74033 , \74034 , \74035 , \74036 , \74037 , \74038 , \74039 , \74040 , \74041 , \74042 ,
         \74043 , \74044 , \74045 , \74046 , \74047 , \74048 , \74049 , \74050 , \74051 , \74052 ,
         \74053 , \74054 , \74055 , \74056 , \74057 , \74058 , \74059 , \74060 , \74061 , \74062 ,
         \74063 , \74064 , \74065 , \74066 , \74067 , \74068 , \74069 , \74070 , \74071 , \74072 ,
         \74073 , \74074 , \74075 , \74076 , \74077 , \74078 , \74079 , \74080 , \74081 , \74082 ,
         \74083 , \74084 , \74085 , \74086 , \74087 , \74088 , \74089 , \74090 , \74091 , \74092 ,
         \74093 , \74094 , \74095 , \74096 , \74097 , \74098 , \74099 , \74100 , \74101 , \74102 ,
         \74103 , \74104 , \74105 , \74106 , \74107 , \74108 , \74109 , \74110 , \74111 , \74112 ,
         \74113 , \74114 , \74115 , \74116 , \74117 , \74118 , \74119 , \74120 , \74121 , \74122 ,
         \74123 , \74124 , \74125 , \74126 , \74127 , \74128 , \74129 , \74130 , \74131 , \74132 ,
         \74133 , \74134 , \74135 , \74136 , \74137 , \74138 , \74139 , \74140 , \74141 , \74142 ,
         \74143 , \74144 , \74145 , \74146 , \74147 , \74148 , \74149 , \74150 , \74151 , \74152 ,
         \74153 , \74154 , \74155 , \74156 , \74157 , \74158 , \74159 , \74160 , \74161 , \74162 ,
         \74163 , \74164 , \74165 , \74166 , \74167 , \74168 , \74169 , \74170 , \74171 , \74172 ,
         \74173 , \74174 , \74175 , \74176 , \74177 , \74178 , \74179 , \74180 , \74181 , \74182 ,
         \74183 , \74184 , \74185 , \74186 , \74187 , \74188 , \74189 , \74190 , \74191 , \74192 ,
         \74193 , \74194 , \74195 , \74196 , \74197 , \74198 , \74199 , \74200 , \74201 , \74202 ,
         \74203 , \74204 , \74205 , \74206 , \74207 , \74208 , \74209 , \74210 , \74211 , \74212 ,
         \74213 , \74214 , \74215 , \74216 , \74217 , \74218 , \74219 , \74220 , \74221 , \74222 ,
         \74223 , \74224 , \74225 , \74226 , \74227 , \74228 , \74229 , \74230 , \74231 , \74232 ,
         \74233 , \74234 , \74235 , \74236 , \74237 , \74238 , \74239 , \74240 , \74241 , \74242 ,
         \74243 , \74244 , \74245 , \74246 , \74247 , \74248 , \74249 , \74250 , \74251 , \74252 ,
         \74253 , \74254 , \74255 , \74256 , \74257 , \74258 , \74259 , \74260 , \74261 , \74262 ,
         \74263 , \74264 , \74265 , \74266 , \74267 , \74268 , \74269 , \74270 , \74271 , \74272 ,
         \74273 , \74274 , \74275 , \74276 , \74277 , \74278 , \74279 , \74280 , \74281 , \74282 ,
         \74283 , \74284 , \74285 , \74286 , \74287 , \74288 , \74289 , \74290 , \74291 , \74292 ,
         \74293 , \74294 , \74295 , \74296 , \74297 , \74298 , \74299 , \74300 , \74301 , \74302 ,
         \74303 , \74304 , \74305 , \74306 , \74307 , \74308 , \74309 , \74310 , \74311 , \74312 ,
         \74313 , \74314 , \74315 , \74316 , \74317 , \74318 , \74319 , \74320 , \74321 , \74322 ,
         \74323 , \74324 , \74325 , \74326 , \74327 , \74328 , \74329 , \74330 , \74331 , \74332 ,
         \74333 , \74334 , \74335 , \74336 , \74337 , \74338 , \74339 , \74340 , \74341 , \74342 ,
         \74343 , \74344 , \74345 , \74346 , \74347 , \74348 , \74349 , \74350 , \74351 , \74352 ,
         \74353 , \74354 , \74355 , \74356 , \74357 , \74358 , \74359 , \74360 , \74361 , \74362 ,
         \74363 , \74364 , \74365 , \74366 , \74367 , \74368 , \74369 , \74370 , \74371 , \74372 ,
         \74373 , \74374 , \74375 , \74376 , \74377 , \74378 , \74379 , \74380 , \74381 , \74382 ,
         \74383 , \74384 , \74385 , \74386 , \74387 , \74388 , \74389 , \74390 , \74391 , \74392 ,
         \74393 , \74394 , \74395 , \74396 , \74397 , \74398 , \74399 , \74400 , \74401 , \74402 ,
         \74403 , \74404 , \74405 , \74406 , \74407 , \74408 , \74409 , \74410 , \74411 , \74412 ,
         \74413 , \74414 , \74415 , \74416 , \74417 , \74418 , \74419 , \74420 , \74421 , \74422 ,
         \74423 , \74424 , \74425 , \74426 , \74427 , \74428 , \74429 , \74430 , \74431 , \74432 ,
         \74433 , \74434 , \74435 , \74436 , \74437 , \74438 , \74439 , \74440 , \74441 , \74442 ,
         \74443 , \74444 , \74445 , \74446 , \74447 , \74448 , \74449 , \74450 , \74451 , \74452 ,
         \74453 , \74454 , \74455 , \74456 , \74457 , \74458 , \74459 , \74460 , \74461 , \74462 ,
         \74463 , \74464 , \74465 , \74466 , \74467 , \74468 , \74469 , \74470 , \74471 , \74472 ,
         \74473 , \74474 , \74475 , \74476 , \74477 , \74478 , \74479 , \74480 , \74481 , \74482 ,
         \74483 , \74484 , \74485 , \74486 , \74487 , \74488 , \74489 , \74490 , \74491 , \74492 ,
         \74493 , \74494 , \74495 , \74496 , \74497 , \74498 , \74499 , \74500 , \74501 , \74502 ,
         \74503 , \74504 , \74505 , \74506 , \74507 , \74508 , \74509 , \74510 , \74511 , \74512 ,
         \74513 , \74514 , \74515 , \74516 , \74517 , \74518 , \74519 , \74520 , \74521 , \74522 ,
         \74523 , \74524 , \74525 , \74526 , \74527 , \74528 , \74529 , \74530 , \74531 , \74532 ,
         \74533 , \74534 , \74535 , \74536 , \74537 , \74538 , \74539 , \74540 , \74541 , \74542 ,
         \74543 , \74544 , \74545 , \74546 , \74547 , \74548 , \74549 , \74550 , \74551 , \74552 ,
         \74553 , \74554 , \74555 , \74556 , \74557 , \74558 , \74559 , \74560 , \74561 , \74562 ,
         \74563 , \74564 , \74565 , \74566 , \74567 , \74568 , \74569 , \74570 , \74571 , \74572 ,
         \74573 , \74574 , \74575 , \74576 , \74577 , \74578 , \74579 , \74580 , \74581 , \74582 ,
         \74583 , \74584 , \74585 , \74586 , \74587 , \74588 , \74589 , \74590 , \74591 , \74592 ,
         \74593 , \74594 , \74595 , \74596 , \74597 , \74598 , \74599 , \74600 , \74601 , \74602 ,
         \74603 , \74604 , \74605 , \74606 , \74607 , \74608 , \74609 , \74610 , \74611 , \74612 ,
         \74613 , \74614 , \74615 , \74616 , \74617 , \74618 , \74619 , \74620 , \74621 , \74622 ,
         \74623 , \74624 , \74625 , \74626 , \74627 , \74628 , \74629 , \74630 , \74631 , \74632 ,
         \74633 , \74634 , \74635 , \74636 , \74637 , \74638 , \74639 , \74640 , \74641 , \74642 ,
         \74643 , \74644 , \74645 , \74646 , \74647 , \74648 , \74649 , \74650 , \74651 , \74652 ,
         \74653 , \74654 , \74655 , \74656 , \74657 , \74658 , \74659 , \74660 , \74661 , \74662 ,
         \74663 , \74664 , \74665 , \74666 , \74667 , \74668 , \74669 , \74670 , \74671 , \74672 ,
         \74673 , \74674 , \74675 , \74676 , \74677 , \74678 , \74679 , \74680 , \74681 , \74682 ,
         \74683 , \74684 , \74685 , \74686 , \74687 , \74688 , \74689 , \74690 , \74691 , \74692 ,
         \74693 , \74694 , \74695 , \74696 , \74697 , \74698 , \74699 , \74700 , \74701 , \74702 ,
         \74703 , \74704 , \74705 , \74706 , \74707 , \74708 , \74709 , \74710 , \74711 , \74712 ,
         \74713 , \74714 , \74715 , \74716 , \74717 , \74718 , \74719 , \74720 , \74721 , \74722 ,
         \74723 , \74724 , \74725 , \74726 , \74727 , \74728 , \74729 , \74730 , \74731 , \74732 ,
         \74733 , \74734 , \74735 , \74736 , \74737 , \74738 , \74739 , \74740 , \74741 , \74742 ,
         \74743 , \74744 , \74745 , \74746 , \74747 , \74748 , \74749 , \74750 , \74751 , \74752 ,
         \74753 , \74754 , \74755 , \74756 , \74757 , \74758 , \74759 , \74760 , \74761 , \74762 ,
         \74763 , \74764 , \74765 , \74766 , \74767 , \74768 , \74769 , \74770 , \74771 , \74772 ,
         \74773 , \74774 , \74775 , \74776 , \74777 , \74778 , \74779 , \74780 , \74781 , \74782 ,
         \74783 , \74784 , \74785 , \74786 , \74787 , \74788 , \74789 , \74790 , \74791 , \74792 ,
         \74793 , \74794 , \74795 , \74796 , \74797 , \74798 , \74799 , \74800 , \74801 , \74802 ,
         \74803 , \74804 , \74805 , \74806 , \74807 , \74808 , \74809 , \74810 , \74811 , \74812 ,
         \74813 , \74814 , \74815 , \74816 , \74817 , \74818 , \74819 , \74820 , \74821 , \74822 ,
         \74823 , \74824 , \74825 , \74826 , \74827 , \74828 , \74829 , \74830 , \74831 , \74832 ,
         \74833 , \74834 , \74835 , \74836 , \74837 , \74838 , \74839 , \74840 , \74841 , \74842 ,
         \74843 , \74844 , \74845 , \74846 , \74847 , \74848 , \74849 , \74850 , \74851 , \74852 ,
         \74853 , \74854 , \74855 , \74856 , \74857 , \74858 , \74859 , \74860 , \74861 , \74862 ,
         \74863 , \74864 , \74865 , \74866 , \74867 , \74868 , \74869 , \74870 , \74871 , \74872 ,
         \74873 , \74874 , \74875 , \74876 , \74877 , \74878 , \74879 , \74880 , \74881 , \74882 ,
         \74883 , \74884 , \74885 , \74886 , \74887 , \74888 , \74889 , \74890 , \74891 , \74892 ,
         \74893 , \74894 , \74895 , \74896 , \74897 , \74898 , \74899 , \74900 , \74901 , \74902 ,
         \74903 , \74904 , \74905 , \74906 , \74907 , \74908 , \74909 , \74910 , \74911 , \74912 ,
         \74913 , \74914 , \74915 , \74916 , \74917 , \74918 , \74919 , \74920 , \74921 , \74922 ,
         \74923 , \74924 , \74925 , \74926 , \74927 , \74928 , \74929 , \74930 , \74931 , \74932 ,
         \74933 , \74934 , \74935 , \74936 , \74937 , \74938 , \74939 , \74940 , \74941 , \74942 ,
         \74943 , \74944 , \74945 , \74946 , \74947 , \74948 , \74949 , \74950 , \74951 , \74952 ,
         \74953 , \74954 , \74955 , \74956 , \74957 , \74958 , \74959 , \74960 , \74961 , \74962 ,
         \74963 , \74964 , \74965 , \74966 , \74967 , \74968 , \74969 , \74970 , \74971 , \74972 ,
         \74973 , \74974 , \74975 , \74976 , \74977 , \74978 , \74979 , \74980 , \74981 , \74982 ,
         \74983 , \74984 , \74985 , \74986 , \74987 , \74988 , \74989 , \74990 , \74991 , \74992 ,
         \74993 , \74994 , \74995 , \74996 , \74997 , \74998 , \74999 , \75000 , \75001 , \75002 ,
         \75003 , \75004 , \75005 , \75006 , \75007 , \75008 , \75009 , \75010 , \75011 , \75012 ,
         \75013 , \75014 , \75015 , \75016 , \75017 , \75018 , \75019 , \75020 , \75021 , \75022 ,
         \75023 , \75024 , \75025 , \75026 , \75027 , \75028 , \75029 , \75030 , \75031 , \75032 ,
         \75033 , \75034 , \75035 , \75036 , \75037 , \75038 , \75039 , \75040 , \75041 , \75042 ,
         \75043 , \75044 , \75045 , \75046 , \75047 , \75048 , \75049 , \75050 , \75051 , \75052 ,
         \75053 , \75054 , \75055 , \75056 , \75057 , \75058 , \75059 , \75060 , \75061 , \75062 ,
         \75063 , \75064 , \75065 , \75066 , \75067 , \75068 , \75069 , \75070 , \75071 , \75072 ,
         \75073 , \75074 , \75075 , \75076 , \75077 , \75078 , \75079 , \75080 , \75081 , \75082 ,
         \75083 , \75084 , \75085 , \75086 , \75087 , \75088 , \75089 , \75090 , \75091 , \75092 ,
         \75093 , \75094 , \75095 , \75096 , \75097 , \75098 , \75099 , \75100 , \75101 , \75102 ,
         \75103 , \75104 , \75105 , \75106 , \75107 , \75108 , \75109 , \75110 , \75111 , \75112 ,
         \75113 , \75114 , \75115 , \75116 , \75117 , \75118 , \75119 , \75120 , \75121 , \75122 ,
         \75123 , \75124 , \75125 , \75126 , \75127 , \75128 , \75129 , \75130 , \75131 , \75132 ,
         \75133 , \75134 , \75135 , \75136 , \75137 , \75138 , \75139 , \75140 , \75141 , \75142 ,
         \75143 , \75144 , \75145 , \75146 , \75147 , \75148 , \75149 , \75150 , \75151 , \75152 ,
         \75153 , \75154 , \75155 , \75156 , \75157 , \75158 , \75159 , \75160 , \75161 , \75162 ,
         \75163 , \75164 , \75165 , \75166 , \75167 , \75168 , \75169 , \75170 , \75171 , \75172 ,
         \75173 , \75174 , \75175 , \75176 , \75177 , \75178 , \75179 , \75180 , \75181 , \75182 ,
         \75183 , \75184 , \75185 , \75186 , \75187 , \75188 , \75189 , \75190 , \75191 , \75192 ,
         \75193 , \75194 , \75195 , \75196 , \75197 , \75198 , \75199 , \75200 , \75201 , \75202 ,
         \75203 , \75204 , \75205 , \75206 , \75207 , \75208 , \75209 , \75210 , \75211 , \75212 ,
         \75213 , \75214 , \75215 , \75216 , \75217 , \75218 , \75219 , \75220 , \75221 , \75222 ,
         \75223 , \75224 , \75225 , \75226 , \75227 , \75228 , \75229 , \75230 , \75231 , \75232 ,
         \75233 , \75234 , \75235 , \75236 , \75237 , \75238 , \75239 , \75240 , \75241 , \75242 ,
         \75243 , \75244 , \75245 , \75246 , \75247 , \75248 , \75249 , \75250 , \75251 , \75252 ,
         \75253 , \75254 , \75255 , \75256 , \75257 , \75258 , \75259 , \75260 , \75261 , \75262 ,
         \75263 , \75264 , \75265 , \75266 , \75267 , \75268 , \75269 , \75270 , \75271 , \75272 ,
         \75273 , \75274 , \75275 , \75276 , \75277 , \75278 , \75279 , \75280 , \75281 , \75282 ,
         \75283 , \75284 , \75285 , \75286 , \75287 , \75288 , \75289 , \75290 , \75291 , \75292 ,
         \75293 , \75294 , \75295 , \75296 , \75297 , \75298 , \75299 , \75300 , \75301 , \75302 ,
         \75303 , \75304 , \75305 , \75306 , \75307 , \75308 , \75309 , \75310 , \75311 , \75312 ,
         \75313 , \75314 , \75315 , \75316 , \75317 , \75318 , \75319 , \75320 , \75321 , \75322 ,
         \75323 , \75324 , \75325 , \75326 , \75327 , \75328 , \75329 , \75330 , \75331 , \75332 ,
         \75333 , \75334 , \75335 , \75336 , \75337 , \75338 , \75339 , \75340 , \75341 , \75342 ,
         \75343 , \75344 , \75345 , \75346 , \75347 , \75348 , \75349 , \75350 , \75351 , \75352 ,
         \75353 , \75354 , \75355 , \75356 , \75357 , \75358 , \75359 , \75360 , \75361 , \75362 ,
         \75363 , \75364 , \75365 , \75366 , \75367 , \75368 , \75369 , \75370 , \75371 , \75372 ,
         \75373 , \75374 , \75375 , \75376 , \75377 , \75378 , \75379 , \75380 , \75381 , \75382 ,
         \75383 , \75384 , \75385 , \75386 , \75387 , \75388 , \75389 , \75390 , \75391 , \75392 ,
         \75393 , \75394 , \75395 , \75396 , \75397 , \75398 , \75399 , \75400 , \75401 , \75402 ,
         \75403 , \75404 , \75405 , \75406 , \75407 , \75408 , \75409 , \75410 , \75411 , \75412 ,
         \75413 , \75414 , \75415 , \75416 , \75417 , \75418 , \75419 , \75420 , \75421 , \75422 ,
         \75423 , \75424 , \75425 , \75426 , \75427 , \75428 , \75429 , \75430 , \75431 , \75432 ,
         \75433 , \75434 , \75435 , \75436 , \75437 , \75438 , \75439 , \75440 , \75441 , \75442 ,
         \75443 , \75444 , \75445 , \75446 , \75447 , \75448 , \75449 , \75450 , \75451 , \75452 ,
         \75453 , \75454 , \75455 , \75456 , \75457 , \75458 , \75459 , \75460 , \75461 , \75462 ,
         \75463 , \75464 , \75465 , \75466 , \75467 , \75468 , \75469 , \75470 , \75471 , \75472 ,
         \75473 , \75474 , \75475 , \75476 , \75477 , \75478 , \75479 , \75480 , \75481 , \75482 ,
         \75483 , \75484 , \75485 , \75486 , \75487 , \75488 , \75489 , \75490 , \75491 , \75492 ,
         \75493 , \75494 , \75495 , \75496 , \75497 , \75498 , \75499 , \75500 , \75501 , \75502 ,
         \75503 , \75504 , \75505 , \75506 , \75507 , \75508 , \75509 , \75510 , \75511 , \75512 ,
         \75513 , \75514 , \75515 , \75516 , \75517 , \75518 , \75519 , \75520 , \75521 , \75522 ,
         \75523 , \75524 , \75525 , \75526 , \75527 , \75528 , \75529 , \75530 , \75531 , \75532 ,
         \75533 , \75534 , \75535 , \75536 , \75537 , \75538 , \75539 , \75540 , \75541 , \75542 ,
         \75543 , \75544 , \75545 , \75546 , \75547 , \75548 , \75549 , \75550 , \75551 , \75552 ,
         \75553 , \75554 , \75555 , \75556 , \75557 , \75558 , \75559 , \75560 , \75561 , \75562 ,
         \75563 , \75564 , \75565 , \75566 , \75567 , \75568 , \75569 , \75570 , \75571 , \75572 ,
         \75573 , \75574 , \75575 , \75576 , \75577 , \75578 , \75579 , \75580 , \75581 , \75582 ,
         \75583 , \75584 , \75585 , \75586 , \75587 , \75588 , \75589 , \75590 , \75591 , \75592 ,
         \75593 , \75594 , \75595 , \75596 , \75597 , \75598 , \75599 , \75600 , \75601 , \75602 ,
         \75603 , \75604 , \75605 , \75606 , \75607 , \75608 , \75609 , \75610 , \75611 , \75612 ,
         \75613 , \75614 , \75615 , \75616 , \75617 , \75618 , \75619 , \75620 , \75621 , \75622 ,
         \75623 , \75624 , \75625 , \75626 , \75627 , \75628 , \75629 , \75630 , \75631 , \75632 ,
         \75633 , \75634 , \75635 , \75636 , \75637 , \75638 , \75639 , \75640 , \75641 , \75642 ,
         \75643 , \75644 , \75645 , \75646 , \75647 , \75648 , \75649 , \75650 , \75651 , \75652 ,
         \75653 , \75654 , \75655 , \75656 , \75657 , \75658 , \75659 , \75660 , \75661 , \75662 ,
         \75663 , \75664 , \75665 , \75666 , \75667 , \75668 , \75669 , \75670 , \75671 , \75672 ,
         \75673 , \75674 , \75675 , \75676 , \75677 , \75678 , \75679 , \75680 , \75681 , \75682 ,
         \75683 , \75684 , \75685 , \75686 , \75687 , \75688 , \75689 , \75690 , \75691 , \75692 ,
         \75693 , \75694 , \75695 , \75696 , \75697 , \75698 , \75699 , \75700 , \75701 , \75702 ,
         \75703 , \75704 , \75705 , \75706 , \75707 , \75708 , \75709 , \75710 , \75711 , \75712 ,
         \75713 , \75714 , \75715 , \75716 , \75717 , \75718 , \75719 , \75720 , \75721 , \75722 ,
         \75723 , \75724 , \75725 , \75726 , \75727 , \75728 , \75729 , \75730 , \75731 , \75732 ,
         \75733 , \75734 , \75735 , \75736 , \75737 , \75738 , \75739 , \75740 , \75741 , \75742 ,
         \75743 , \75744 , \75745 , \75746 , \75747 , \75748 , \75749 , \75750 , \75751 , \75752 ,
         \75753 , \75754 , \75755 , \75756 , \75757 , \75758 , \75759 , \75760 , \75761 , \75762 ,
         \75763 , \75764 , \75765 , \75766 , \75767 , \75768 , \75769 , \75770 , \75771 , \75772 ,
         \75773 , \75774 , \75775 , \75776 , \75777 , \75778 , \75779 , \75780 , \75781 , \75782 ,
         \75783 , \75784 , \75785 , \75786 , \75787 , \75788 , \75789 , \75790 , \75791 , \75792 ,
         \75793 , \75794 , \75795 , \75796 , \75797 , \75798 , \75799 , \75800 , \75801 , \75802 ,
         \75803 , \75804 , \75805 , \75806 , \75807 , \75808 , \75809 , \75810 , \75811 , \75812 ,
         \75813 , \75814 , \75815 , \75816 , \75817 , \75818 , \75819 , \75820 , \75821 , \75822 ,
         \75823 , \75824 , \75825 , \75826 , \75827 , \75828 , \75829 , \75830 , \75831 , \75832 ,
         \75833 , \75834 , \75835 , \75836 , \75837 , \75838 , \75839 , \75840 , \75841 , \75842 ,
         \75843 , \75844 , \75845 , \75846 , \75847 , \75848 , \75849 , \75850 , \75851 , \75852 ,
         \75853 , \75854 , \75855 , \75856 , \75857 , \75858 , \75859 , \75860 , \75861 , \75862 ,
         \75863 , \75864 , \75865 , \75866 , \75867 , \75868 , \75869 , \75870 , \75871 , \75872 ,
         \75873 , \75874 , \75875 , \75876 , \75877 , \75878 , \75879 , \75880 , \75881 , \75882 ,
         \75883 , \75884 , \75885 , \75886 , \75887 , \75888 , \75889 , \75890 , \75891 , \75892 ,
         \75893 , \75894 , \75895 , \75896 , \75897 , \75898 , \75899 , \75900 , \75901 , \75902 ,
         \75903 , \75904 , \75905 , \75906 , \75907 , \75908 , \75909 , \75910 , \75911 , \75912 ,
         \75913 , \75914 , \75915 , \75916 , \75917 , \75918 , \75919 , \75920 , \75921 , \75922 ,
         \75923 , \75924 , \75925 , \75926 , \75927 , \75928 , \75929 , \75930 , \75931 , \75932 ,
         \75933 , \75934 , \75935 , \75936 , \75937 , \75938 , \75939 , \75940 , \75941 , \75942 ,
         \75943 , \75944 , \75945 , \75946 , \75947 , \75948 , \75949 , \75950 , \75951 , \75952 ,
         \75953 , \75954 , \75955 , \75956 , \75957 , \75958 , \75959 , \75960 , \75961 , \75962 ,
         \75963 , \75964 , \75965 , \75966 , \75967 , \75968 , \75969 , \75970 , \75971 , \75972 ,
         \75973 , \75974 , \75975 , \75976 , \75977 , \75978 , \75979 , \75980 , \75981 , \75982 ,
         \75983 , \75984 , \75985 , \75986 , \75987 , \75988 , \75989 , \75990 , \75991 , \75992 ,
         \75993 , \75994 , \75995 , \75996 , \75997 , \75998 , \75999 , \76000 , \76001 , \76002 ,
         \76003 , \76004 , \76005 , \76006 , \76007 , \76008 , \76009 , \76010 , \76011 , \76012 ,
         \76013 , \76014 , \76015 , \76016 , \76017 , \76018 , \76019 , \76020 , \76021 , \76022 ,
         \76023 , \76024 , \76025 , \76026 , \76027 , \76028 , \76029 , \76030 , \76031 , \76032 ,
         \76033 , \76034 , \76035 , \76036 , \76037 , \76038 , \76039 , \76040 , \76041 , \76042 ,
         \76043 , \76044 , \76045 , \76046 , \76047 , \76048 , \76049 , \76050 , \76051 , \76052 ,
         \76053 , \76054 , \76055 , \76056 , \76057 , \76058 , \76059 , \76060 , \76061 , \76062 ,
         \76063 , \76064 , \76065 , \76066 , \76067 , \76068 , \76069 , \76070 , \76071 , \76072 ,
         \76073 , \76074 , \76075 , \76076 , \76077 , \76078 , \76079 , \76080 , \76081 , \76082 ,
         \76083 , \76084 , \76085 , \76086 , \76087 , \76088 , \76089 , \76090 , \76091 , \76092 ,
         \76093 , \76094 , \76095 , \76096 , \76097 , \76098 , \76099 , \76100 , \76101 , \76102 ,
         \76103 , \76104 , \76105 , \76106 , \76107 , \76108 , \76109 , \76110 , \76111 , \76112 ,
         \76113 , \76114 , \76115 , \76116 , \76117 , \76118 , \76119 , \76120 , \76121 , \76122 ,
         \76123 , \76124 , \76125 , \76126 , \76127 , \76128 , \76129 , \76130 , \76131 , \76132 ,
         \76133 , \76134 , \76135 , \76136 , \76137 , \76138 , \76139 , \76140 , \76141 , \76142 ,
         \76143 , \76144 , \76145 , \76146 , \76147 , \76148 , \76149 , \76150 , \76151 , \76152 ,
         \76153 , \76154 , \76155 , \76156 , \76157 , \76158 , \76159 , \76160 , \76161 , \76162 ,
         \76163 , \76164 , \76165 , \76166 , \76167 , \76168 , \76169 , \76170 , \76171 , \76172 ,
         \76173 , \76174 , \76175 , \76176 , \76177 , \76178 , \76179 , \76180 , \76181 , \76182 ,
         \76183 , \76184 , \76185 , \76186 , \76187 , \76188 , \76189 , \76190 , \76191 , \76192 ,
         \76193 , \76194 , \76195 , \76196 , \76197 , \76198 , \76199 , \76200 , \76201 , \76202 ,
         \76203 , \76204 , \76205 , \76206 , \76207 , \76208 , \76209 , \76210 , \76211 , \76212 ,
         \76213 , \76214 , \76215 , \76216 , \76217 , \76218 , \76219 , \76220 , \76221 , \76222 ,
         \76223 , \76224 , \76225 , \76226 , \76227 , \76228 , \76229 , \76230 , \76231 , \76232 ,
         \76233 , \76234 , \76235 , \76236 , \76237 , \76238 , \76239 , \76240 , \76241 , \76242 ,
         \76243 , \76244 , \76245 , \76246 , \76247 , \76248 , \76249 , \76250 , \76251 , \76252 ,
         \76253 , \76254 , \76255 , \76256 , \76257 , \76258 , \76259 , \76260 , \76261 , \76262 ,
         \76263 , \76264 , \76265 , \76266 , \76267 , \76268 , \76269 , \76270 , \76271 , \76272 ,
         \76273 , \76274 , \76275 , \76276 , \76277 , \76278 , \76279 , \76280 , \76281 , \76282 ,
         \76283 , \76284 , \76285 , \76286 , \76287 , \76288 , \76289 , \76290 , \76291 , \76292 ,
         \76293 , \76294 , \76295 , \76296 , \76297 , \76298 , \76299 , \76300 , \76301 , \76302 ,
         \76303 , \76304 , \76305 , \76306 , \76307 , \76308 , \76309 , \76310 , \76311 , \76312 ,
         \76313 , \76314 , \76315 , \76316 , \76317 , \76318 , \76319 , \76320 , \76321 , \76322 ,
         \76323 , \76324 , \76325 , \76326 , \76327 , \76328 , \76329 , \76330 , \76331 , \76332 ,
         \76333 , \76334 , \76335 , \76336 , \76337 , \76338 , \76339 , \76340 , \76341 , \76342 ,
         \76343 , \76344 , \76345 , \76346 , \76347 , \76348 , \76349 , \76350 , \76351 , \76352 ,
         \76353 , \76354 , \76355 , \76356 , \76357 , \76358 , \76359 , \76360 , \76361 , \76362 ,
         \76363 , \76364 , \76365 , \76366 , \76367 , \76368 , \76369 , \76370 , \76371 , \76372 ,
         \76373 , \76374 , \76375 , \76376 , \76377 , \76378 , \76379 , \76380 , \76381 , \76382 ,
         \76383 , \76384 , \76385 , \76386 , \76387 , \76388 , \76389 , \76390 , \76391 , \76392 ,
         \76393 , \76394 , \76395 , \76396 , \76397 , \76398 , \76399 , \76400 , \76401 , \76402 ,
         \76403 , \76404 , \76405 , \76406 , \76407 , \76408 , \76409 , \76410 , \76411 , \76412 ,
         \76413 , \76414 , \76415 , \76416 , \76417 , \76418 , \76419 , \76420 , \76421 , \76422 ,
         \76423 , \76424 , \76425 , \76426 , \76427 , \76428 , \76429 , \76430 , \76431 , \76432 ,
         \76433 , \76434 , \76435 , \76436 , \76437 , \76438 , \76439 , \76440 , \76441 , \76442 ,
         \76443 , \76444 , \76445 , \76446 , \76447 , \76448 , \76449 , \76450 , \76451 , \76452 ,
         \76453 , \76454 , \76455 , \76456 , \76457 , \76458 , \76459 , \76460 , \76461 , \76462 ,
         \76463 , \76464 , \76465 , \76466 , \76467 , \76468 , \76469 , \76470 , \76471 , \76472 ,
         \76473 , \76474 , \76475 , \76476 , \76477 , \76478 , \76479 , \76480 , \76481 , \76482 ;
buf \U$labaj7679 ( R_81_84446b8, \73053 );
buf \U$labaj7680 ( R_82_8444760, \73126 );
buf \U$labaj7681 ( R_83_8444808, \73169 );
buf \U$labaj7682 ( R_84_84448b0, \73204 );
buf \U$labaj7683 ( R_85_8444958, \73245 );
buf \U$labaj7684 ( R_86_8444a00, \73280 );
buf \U$labaj7685 ( R_87_9bec6f8, \73318 );
buf \U$labaj7686 ( R_88_9bec7a0, \73345 );
buf \U$labaj7687 ( R_89_9bec848, \73386 );
buf \U$labaj7688 ( R_8a_9bec8f0, \73447 );
buf \U$labaj7689 ( R_8b_9bec998, \73474 );
buf \U$labaj7690 ( R_8c_9beca40, \73490 );
buf \U$labaj7691 ( R_8d_9becae8, \73542 );
buf \U$labaj7692 ( R_8e_9becb90, \73569 );
buf \U$labaj7693 ( R_8f_9becc38, \73610 );
buf \U$labaj7694 ( R_90_9becce0, \73634 );
buf \U$labaj7695 ( R_91_9becd88, \73702 );
buf \U$labaj7696 ( R_92_9bece30, \73745 );
buf \U$labaj7697 ( R_93_9beced8, \73782 );
buf \U$labaj7698 ( R_94_9becf80, \73809 );
buf \U$labaj7699 ( R_95_9bed028, \73858 );
buf \U$labaj7700 ( R_96_9bed0d0, \73882 );
buf \U$labaj7701 ( R_97_9bed178, \73910 );
buf \U$labaj7702 ( R_98_9bed220, \73935 );
buf \U$labaj7703 ( R_99_9bed2c8, \73986 );
buf \U$labaj7704 ( R_9a_9bed370, \74010 );
buf \U$labaj7705 ( R_9b_9bed418, \74044 );
buf \U$labaj7706 ( R_9c_9bed4c0, \74072 );
buf \U$labaj7707 ( R_9d_9bed568, \74102 );
buf \U$labaj7708 ( R_9e_9bed610, \74132 );
buf \U$labaj7709 ( R_9f_9bed6b8, \74156 );
buf \U$labaj7710 ( R_a0_9bed760, \74172 );
buf \U$labaj7711 ( R_a1_9bed808, \74273 );
buf \U$labaj7712 ( R_a2_9bed8b0, \74315 );
buf \U$labaj7713 ( R_a3_9bed958, \74352 );
buf \U$labaj7714 ( R_a4_9beda00, \74379 );
buf \U$labaj7715 ( R_a5_9bedaa8, \74430 );
buf \U$labaj7716 ( R_a6_9bedb50, \74457 );
buf \U$labaj7717 ( R_a7_9bedbf8, \74491 );
buf \U$labaj7718 ( R_a8_9bedca0, \74518 );
buf \U$labaj7719 ( R_a9_9bedd48, \74579 );
buf \U$labaj7720 ( R_aa_9beddf0, \74600 );
buf \U$labaj7721 ( R_ab_9bede98, \74636 );
buf \U$labaj7722 ( R_ac_9bedf40, \74651 );
buf \U$labaj7723 ( R_ad_9bedfe8, \74678 );
buf \U$labaj7724 ( R_ae_9bee090, \74705 );
buf \U$labaj7725 ( R_af_9bee138, \74729 );
buf \U$labaj7726 ( R_b0_9bee1e0, \74747 );
buf \U$labaj7727 ( R_b1_9bee288, \74826 );
buf \U$labaj7728 ( R_b2_9bee330, \74857 );
buf \U$labaj7729 ( R_b3_9bee3d8, \74887 );
buf \U$labaj7730 ( R_b4_9bee480, \74915 );
buf \U$labaj7731 ( R_b5_9bee528, \74942 );
buf \U$labaj7732 ( R_b6_9bee5d0, \74977 );
buf \U$labaj7733 ( R_b7_9bee678, \75001 );
buf \U$labaj7734 ( R_b8_9bee720, \75016 );
buf \U$labaj7735 ( R_b9_9bee7c8, \75075 );
buf \U$labaj7736 ( R_ba_9bee870, \75102 );
buf \U$labaj7737 ( R_bb_9bee918, \75129 );
buf \U$labaj7738 ( R_bc_9bee9c0, \75144 );
buf \U$labaj7739 ( R_bd_9beea68, \75190 );
buf \U$labaj7740 ( R_be_9beeb10, \75205 );
buf \U$labaj7741 ( R_bf_9beebb8, \75229 );
buf \U$labaj7742 ( R_c0_9beec60, \75239 );
buf \U$labaj7743 ( R_c1_9beed08, \75296 );
buf \U$labaj7744 ( R_c2_9beedb0, \75328 );
buf \U$labaj7745 ( R_c3_9beee58, \75352 );
buf \U$labaj7746 ( R_c4_9beef00, \75367 );
buf \U$labaj7747 ( R_c5_9beefa8, \75407 );
buf \U$labaj7748 ( R_c6_9bef050, \75422 );
buf \U$labaj7749 ( R_c7_9bef0f8, \75446 );
buf \U$labaj7750 ( R_c8_9bef1a0, \75461 );
buf \U$labaj7751 ( R_c9_9bef248, \75506 );
buf \U$labaj7752 ( R_ca_9bef2f0, \75521 );
buf \U$labaj7753 ( R_cb_9bef398, \75545 );
buf \U$labaj7754 ( R_cc_9bef440, \75560 );
buf \U$labaj7755 ( R_cd_9bef4e8, \75603 );
buf \U$labaj7756 ( R_ce_9bef590, \75618 );
buf \U$labaj7757 ( R_cf_9bef638, \75642 );
buf \U$labaj7758 ( R_d0_9bef6e0, \75657 );
buf \U$labaj7759 ( R_d1_9bef788, \75709 );
buf \U$labaj7760 ( R_d2_9bef830, \75724 );
buf \U$labaj7761 ( R_d3_9bef8d8, \75749 );
buf \U$labaj7762 ( R_d4_9bef980, \75764 );
buf \U$labaj7763 ( R_d5_9befa28, \75804 );
buf \U$labaj7764 ( R_d6_9befad0, \75819 );
buf \U$labaj7765 ( R_d7_9befb78, \75846 );
buf \U$labaj7766 ( R_d8_9befc20, \75861 );
buf \U$labaj7767 ( R_d9_9befcc8, \75904 );
buf \U$labaj7768 ( R_da_9befd70, \75919 );
buf \U$labaj7769 ( R_db_9befe18, \75946 );
buf \U$labaj7770 ( R_dc_9befec0, \75961 );
buf \U$labaj7771 ( R_dd_9beff68, \75993 );
buf \U$labaj7772 ( R_de_9bf0010, \76008 );
buf \U$labaj7773 ( R_df_9bf00b8, \76032 );
buf \U$labaj7774 ( R_e0_9bf0160, \76048 );
buf \U$labaj7775 ( R_e1_9bf0208, \76101 );
buf \U$labaj7776 ( R_e2_9bf02b0, \76116 );
buf \U$labaj7777 ( R_e3_9bf0358, \76140 );
buf \U$labaj7778 ( R_e4_9bf0400, \76155 );
buf \U$labaj7779 ( R_e5_9bf04a8, \76195 );
buf \U$labaj7780 ( R_e6_9bf0550, \76210 );
buf \U$labaj7781 ( R_e7_9bf05f8, \76238 );
buf \U$labaj7782 ( R_e8_9bf06a0, \76254 );
buf \U$labaj7783 ( R_e9_9bf0748, \76285 );
buf \U$labaj7784 ( R_ea_9bf07f0, \76300 );
buf \U$labaj7785 ( R_eb_9bf0898, \76317 );
buf \U$labaj7786 ( R_ec_9bf0940, \76326 );
buf \U$labaj7787 ( R_ed_9bf09e8, \76354 );
buf \U$labaj7788 ( R_ee_9bf0a90, \76369 );
buf \U$labaj7789 ( R_ef_9bf0b38, \76392 );
buf \U$labaj7790 ( R_f0_9bf0be0, \76407 );
buf \U$labaj7791 ( R_f1_9bf0c88, \76441 );
buf \U$labaj7792 ( R_f2_9bf0d30, \76456 );
buf \U$labaj7793 ( R_f3_9bf0dd8, \76482 );
buf \U$1 ( \246 , RIc0d85f0_34);
buf \U$2 ( \247 , RIc0d9478_65);
and \U$3 ( \248 , \246 , \247 );
buf \U$4 ( \249 , \248 );
buf \U$5 ( \250 , \249 );
xnor \U$6 ( \251 , RIc0d9658_69, RIc0d8398_29);
buf \U$7 ( \252 , \251 );
not \U$8 ( \253 , \252 );
buf \U$9 ( \254 , \253 );
buf \U$10 ( \255 , \254 );
not \U$11 ( \256 , \255 );
buf \U$12 ( \257 , RIc0d96d0_70);
buf \U$13 ( \258 , RIc0d9748_71);
and \U$14 ( \259 , \257 , \258 );
not \U$15 ( \260 , \257 );
buf \U$16 ( \261 , RIc0d9748_71);
not \U$17 ( \262 , \261 );
buf \U$18 ( \263 , \262 );
buf \U$19 ( \264 , \263 );
and \U$20 ( \265 , \260 , \264 );
nor \U$21 ( \266 , \259 , \265 );
buf \U$22 ( \267 , \266 );
buf \U$23 ( \268 , \267 );
not \U$24 ( \269 , \268 );
buf \U$25 ( \270 , \269 );
buf \U$26 ( \271 , \270 );
xor \U$27 ( \272 , RIc0d96d0_70, RIc0d9658_69);
buf \U$28 ( \273 , \272 );
nand \U$29 ( \274 , \271 , \273 );
buf \U$30 ( \275 , \274 );
buf \U$31 ( \276 , \275 );
not \U$32 ( \277 , \276 );
buf \U$33 ( \278 , \277 );
buf \U$36 ( \279 , \278 );
buf \U$37 ( \280 , \279 );
not \U$38 ( \281 , \280 );
or \U$39 ( \282 , \256 , \281 );
buf \U$42 ( \283 , \267 );
buf \U$45 ( \284 , \283 );
buf \U$46 ( \285 , \284 );
buf \U$47 ( \286 , RIc0d9658_69);
buf \U$48 ( \287 , RIc0d8320_28);
xor \U$49 ( \288 , \286 , \287 );
buf \U$50 ( \289 , \288 );
buf \U$51 ( \290 , \289 );
nand \U$52 ( \291 , \285 , \290 );
buf \U$53 ( \292 , \291 );
buf \U$54 ( \293 , \292 );
nand \U$55 ( \294 , \282 , \293 );
buf \U$56 ( \295 , \294 );
buf \U$57 ( \296 , \295 );
xor \U$58 ( \297 , \250 , \296 );
buf \U$59 ( \298 , RIc0da288_95);
buf \U$60 ( \299 , RIc0d7768_3);
and \U$61 ( \300 , \298 , \299 );
not \U$62 ( \301 , \298 );
buf \U$63 ( \302 , RIc0d7768_3);
not \U$64 ( \303 , \302 );
buf \U$65 ( \304 , \303 );
buf \U$66 ( \305 , \304 );
and \U$67 ( \306 , \301 , \305 );
nor \U$68 ( \307 , \300 , \306 );
buf \U$69 ( \308 , \307 );
buf \U$70 ( \309 , \308 );
not \U$71 ( \310 , \309 );
buf \U$72 ( \311 , RIc0da288_95);
buf \U$73 ( \312 , RIc0da300_96);
xor \U$74 ( \313 , \311 , \312 );
buf \U$75 ( \314 , \313 );
buf \U$76 ( \315 , \314 );
buf \U$77 ( \316 , RIc0da300_96);
not \U$78 ( \317 , \316 );
buf \U$79 ( \318 , RIc0da378_97);
nand \U$80 ( \319 , \317 , \318 );
buf \U$81 ( \320 , \319 );
buf \U$82 ( \321 , \320 );
buf \U$83 ( \322 , RIc0da378_97);
not \U$84 ( \323 , \322 );
buf \U$85 ( \324 , RIc0da300_96);
nand \U$86 ( \325 , \323 , \324 );
buf \U$87 ( \326 , \325 );
buf \U$88 ( \327 , \326 );
and \U$89 ( \328 , \315 , \321 , \327 );
buf \U$90 ( \329 , \328 );
buf \U$93 ( \330 , \329 );
buf \U$94 ( \331 , \330 );
not \U$95 ( \332 , \331 );
buf \U$96 ( \333 , \332 );
buf \U$97 ( \334 , \333 );
not \U$98 ( \335 , \334 );
buf \U$99 ( \336 , \335 );
buf \U$100 ( \337 , \336 );
not \U$101 ( \338 , \337 );
or \U$102 ( \339 , \310 , \338 );
buf \U$103 ( \340 , RIc0da300_96);
buf \U$104 ( \341 , RIc0da378_97);
xor \U$105 ( \342 , \340 , \341 );
buf \U$106 ( \343 , \342 );
buf \U$109 ( \344 , \343 );
buf \U$110 ( \345 , \344 );
buf \U$111 ( \346 , RIc0da288_95);
buf \U$112 ( \347 , RIc0d76f0_2);
and \U$113 ( \348 , \346 , \347 );
not \U$114 ( \349 , \346 );
buf \U$115 ( \350 , RIc0d76f0_2);
not \U$116 ( \351 , \350 );
buf \U$117 ( \352 , \351 );
buf \U$118 ( \353 , \352 );
and \U$119 ( \354 , \349 , \353 );
nor \U$120 ( \355 , \348 , \354 );
buf \U$121 ( \356 , \355 );
buf \U$122 ( \357 , \356 );
nand \U$123 ( \358 , \345 , \357 );
buf \U$124 ( \359 , \358 );
buf \U$125 ( \360 , \359 );
nand \U$126 ( \361 , \339 , \360 );
buf \U$127 ( \362 , \361 );
buf \U$128 ( \363 , \362 );
xor \U$129 ( \364 , \297 , \363 );
buf \U$130 ( \365 , \364 );
buf \U$131 ( \366 , \365 );
buf \U$132 ( \367 , RIc0d9b08_79);
buf \U$133 ( \368 , RIc0d7ee8_19);
xor \U$134 ( \369 , \367 , \368 );
buf \U$135 ( \370 , \369 );
buf \U$136 ( \371 , \370 );
not \U$137 ( \372 , \371 );
buf \U$138 ( \373 , RIc0d9b80_80);
not \U$139 ( \374 , \373 );
buf \U$140 ( \375 , RIc0d9b08_79);
nand \U$141 ( \376 , \374 , \375 );
buf \U$142 ( \377 , \376 );
not \U$143 ( \378 , \377 );
buf \U$144 ( \379 , RIc0d9b08_79);
not \U$145 ( \380 , \379 );
buf \U$146 ( \381 , RIc0d9b80_80);
nand \U$147 ( \382 , \380 , \381 );
buf \U$148 ( \383 , \382 );
not \U$149 ( \384 , \383 );
or \U$150 ( \385 , \378 , \384 );
buf \U$151 ( \386 , RIc0d9b80_80);
buf \U$152 ( \387 , RIc0d9bf8_81);
xor \U$153 ( \388 , \386 , \387 );
buf \U$154 ( \389 , \388 );
not \U$155 ( \390 , \389 );
nand \U$156 ( \391 , \385 , \390 );
buf \U$157 ( \392 , \391 );
buf \U$159 ( \393 , \392 );
buf \U$160 ( \394 , \393 );
not \U$161 ( \395 , \394 );
buf \U$162 ( \396 , \395 );
buf \U$165 ( \397 , \396 );
buf \U$166 ( \398 , \397 );
not \U$167 ( \399 , \398 );
or \U$168 ( \400 , \372 , \399 );
buf \U$169 ( \401 , \389 );
buf \U$170 ( \402 , \401 );
buf \U$171 ( \403 , \402 );
buf \U$172 ( \404 , \403 );
buf \U$173 ( \405 , RIc0d7e70_18);
buf \U$174 ( \406 , RIc0d9b08_79);
xor \U$175 ( \407 , \405 , \406 );
buf \U$176 ( \408 , \407 );
buf \U$177 ( \409 , \408 );
nand \U$178 ( \410 , \404 , \409 );
buf \U$179 ( \411 , \410 );
buf \U$180 ( \412 , \411 );
nand \U$181 ( \413 , \400 , \412 );
buf \U$182 ( \414 , \413 );
buf \U$183 ( \415 , RIc0d7a38_9);
buf \U$184 ( \416 , RIc0d9fb8_89);
xor \U$185 ( \417 , \415 , \416 );
buf \U$186 ( \418 , \417 );
buf \U$187 ( \419 , \418 );
not \U$188 ( \420 , \419 );
buf \U$189 ( \421 , RIc0da030_90);
buf \U$190 ( \422 , RIc0da0a8_91);
xor \U$191 ( \423 , \421 , \422 );
buf \U$192 ( \424 , \423 );
buf \U$193 ( \425 , \424 );
not \U$194 ( \426 , \425 );
buf \U$195 ( \427 , \426 );
buf \U$196 ( \428 , \427 );
xor \U$197 ( \429 , RIc0da030_90, RIc0d9fb8_89);
buf \U$198 ( \430 , \429 );
nand \U$199 ( \431 , \428 , \430 );
buf \U$200 ( \432 , \431 );
buf \U$203 ( \433 , \432 );
buf \U$204 ( \434 , \433 );
not \U$205 ( \435 , \434 );
buf \U$206 ( \436 , \435 );
buf \U$209 ( \437 , \436 );
buf \U$210 ( \438 , \437 );
not \U$211 ( \439 , \438 );
or \U$212 ( \440 , \420 , \439 );
buf \U$215 ( \441 , \424 );
buf \U$218 ( \442 , \441 );
buf \U$219 ( \443 , \442 );
buf \U$220 ( \444 , RIc0d79c0_8);
buf \U$221 ( \445 , RIc0d9fb8_89);
xor \U$222 ( \446 , \444 , \445 );
buf \U$223 ( \447 , \446 );
buf \U$224 ( \448 , \447 );
nand \U$225 ( \449 , \443 , \448 );
buf \U$226 ( \450 , \449 );
buf \U$227 ( \451 , \450 );
nand \U$228 ( \452 , \440 , \451 );
buf \U$229 ( \453 , \452 );
xor \U$230 ( \454 , \414 , \453 );
buf \U$231 ( \455 , RIc0d7858_5);
buf \U$232 ( \456 , RIc0da198_93);
xor \U$233 ( \457 , \455 , \456 );
buf \U$234 ( \458 , \457 );
buf \U$235 ( \459 , \458 );
not \U$236 ( \460 , \459 );
buf \U$237 ( \461 , RIc0da210_94);
buf \U$238 ( \462 , RIc0da288_95);
xor \U$239 ( \463 , \461 , \462 );
buf \U$240 ( \464 , \463 );
buf \U$241 ( \465 , \464 );
not \U$242 ( \466 , \465 );
buf \U$243 ( \467 , \466 );
buf \U$244 ( \468 , \467 );
xor \U$245 ( \469 , RIc0da210_94, RIc0da198_93);
buf \U$246 ( \470 , \469 );
nand \U$247 ( \471 , \468 , \470 );
buf \U$248 ( \472 , \471 );
buf \U$251 ( \473 , \472 );
buf \U$252 ( \474 , \473 );
not \U$253 ( \475 , \474 );
buf \U$254 ( \476 , \475 );
buf \U$255 ( \477 , \476 );
not \U$256 ( \478 , \477 );
or \U$257 ( \479 , \460 , \478 );
buf \U$260 ( \480 , \464 );
buf \U$263 ( \481 , \480 );
buf \U$264 ( \482 , \481 );
buf \U$265 ( \483 , RIc0da198_93);
buf \U$266 ( \484 , RIc0d77e0_4);
and \U$267 ( \485 , \483 , \484 );
not \U$268 ( \486 , \483 );
buf \U$269 ( \487 , RIc0d77e0_4);
not \U$270 ( \488 , \487 );
buf \U$271 ( \489 , \488 );
buf \U$272 ( \490 , \489 );
and \U$273 ( \491 , \486 , \490 );
nor \U$274 ( \492 , \485 , \491 );
buf \U$275 ( \493 , \492 );
buf \U$276 ( \494 , \493 );
nand \U$277 ( \495 , \482 , \494 );
buf \U$278 ( \496 , \495 );
buf \U$279 ( \497 , \496 );
nand \U$280 ( \498 , \479 , \497 );
buf \U$281 ( \499 , \498 );
xor \U$282 ( \500 , \454 , \499 );
buf \U$283 ( \501 , \500 );
xor \U$284 ( \502 , \366 , \501 );
buf \U$285 ( \503 , RIc0d7948_7);
buf \U$286 ( \504 , RIc0da0a8_91);
xor \U$287 ( \505 , \503 , \504 );
buf \U$288 ( \506 , \505 );
buf \U$289 ( \507 , \506 );
not \U$290 ( \508 , \507 );
buf \U$291 ( \509 , RIc0da120_92);
buf \U$292 ( \510 , RIc0da198_93);
xor \U$293 ( \511 , \509 , \510 );
buf \U$294 ( \512 , \511 );
buf \U$295 ( \513 , \512 );
not \U$296 ( \514 , \513 );
buf \U$297 ( \515 , \514 );
buf \U$298 ( \516 , \515 );
xor \U$299 ( \517 , RIc0da120_92, RIc0da0a8_91);
buf \U$300 ( \518 , \517 );
nand \U$301 ( \519 , \516 , \518 );
buf \U$302 ( \520 , \519 );
buf \U$305 ( \521 , \520 );
buf \U$306 ( \522 , \521 );
not \U$307 ( \523 , \522 );
buf \U$308 ( \524 , \523 );
buf \U$309 ( \525 , \524 );
not \U$310 ( \526 , \525 );
or \U$311 ( \527 , \508 , \526 );
buf \U$312 ( \528 , \512 );
not \U$313 ( \529 , \528 );
buf \U$314 ( \530 , \529 );
buf \U$315 ( \531 , \530 );
not \U$316 ( \532 , \531 );
buf \U$317 ( \533 , \532 );
buf \U$318 ( \534 , \533 );
buf \U$319 ( \535 , RIc0d78d0_6);
buf \U$320 ( \536 , RIc0da0a8_91);
xor \U$321 ( \537 , \535 , \536 );
buf \U$322 ( \538 , \537 );
buf \U$323 ( \539 , \538 );
nand \U$324 ( \540 , \534 , \539 );
buf \U$325 ( \541 , \540 );
buf \U$326 ( \542 , \541 );
nand \U$327 ( \543 , \527 , \542 );
buf \U$328 ( \544 , \543 );
buf \U$329 ( \545 , \544 );
buf \U$330 ( \546 , RIc0d7d08_15);
buf \U$331 ( \547 , RIc0d9ce8_83);
xnor \U$332 ( \548 , \546 , \547 );
buf \U$333 ( \549 , \548 );
buf \U$334 ( \550 , \549 );
not \U$335 ( \551 , \550 );
buf \U$336 ( \552 , \551 );
buf \U$337 ( \553 , \552 );
not \U$338 ( \554 , \553 );
buf \U$339 ( \555 , RIc0d9d60_84);
buf \U$340 ( \556 , RIc0d9dd8_85);
xor \U$341 ( \557 , \555 , \556 );
buf \U$342 ( \558 , \557 );
buf \U$343 ( \559 , \558 );
not \U$344 ( \560 , \559 );
buf \U$345 ( \561 , \560 );
buf \U$346 ( \562 , \561 );
buf \U$347 ( \563 , RIc0d9ce8_83);
buf \U$348 ( \564 , RIc0d9d60_84);
xor \U$349 ( \565 , \563 , \564 );
buf \U$350 ( \566 , \565 );
buf \U$351 ( \567 , \566 );
nand \U$352 ( \568 , \562 , \567 );
buf \U$353 ( \569 , \568 );
buf \U$354 ( \570 , \569 );
not \U$355 ( \571 , \570 );
buf \U$356 ( \572 , \571 );
buf \U$359 ( \573 , \572 );
buf \U$362 ( \574 , \573 );
buf \U$363 ( \575 , \574 );
not \U$364 ( \576 , \575 );
or \U$365 ( \577 , \554 , \576 );
buf \U$366 ( \578 , RIc0d7c90_14);
buf \U$367 ( \579 , RIc0d9ce8_83);
xnor \U$368 ( \580 , \578 , \579 );
buf \U$369 ( \581 , \580 );
buf \U$370 ( \582 , \581 );
not \U$371 ( \583 , \582 );
buf \U$374 ( \584 , \558 );
buf \U$375 ( \585 , \584 );
nand \U$376 ( \586 , \583 , \585 );
buf \U$377 ( \587 , \586 );
buf \U$378 ( \588 , \587 );
nand \U$379 ( \589 , \577 , \588 );
buf \U$380 ( \590 , \589 );
buf \U$381 ( \591 , \590 );
xor \U$382 ( \592 , \545 , \591 );
buf \U$383 ( \593 , RIc0d9f40_88);
buf \U$384 ( \594 , RIc0d9fb8_89);
and \U$385 ( \595 , \593 , \594 );
not \U$386 ( \596 , \593 );
buf \U$387 ( \597 , RIc0d9fb8_89);
not \U$388 ( \598 , \597 );
buf \U$389 ( \599 , \598 );
buf \U$390 ( \600 , \599 );
and \U$391 ( \601 , \596 , \600 );
nor \U$392 ( \602 , \595 , \601 );
buf \U$393 ( \603 , \602 );
buf \U$394 ( \604 , \603 );
not \U$395 ( \605 , \604 );
xor \U$396 ( \606 , RIc0d9f40_88, RIc0d9ec8_87);
buf \U$397 ( \607 , \606 );
nand \U$398 ( \608 , \605 , \607 );
buf \U$399 ( \609 , \608 );
buf \U$400 ( \610 , \609 );
not \U$401 ( \611 , \610 );
buf \U$402 ( \612 , \611 );
buf \U$403 ( \613 , \612 );
not \U$404 ( \614 , \613 );
buf \U$405 ( \615 , \614 );
buf \U$406 ( \616 , \615 );
not \U$407 ( \617 , \616 );
buf \U$408 ( \618 , \617 );
buf \U$409 ( \619 , \618 );
buf \U$410 ( \620 , RIc0d7b28_11);
buf \U$411 ( \621 , RIc0d9ec8_87);
xor \U$412 ( \622 , \620 , \621 );
buf \U$413 ( \623 , \622 );
buf \U$414 ( \624 , \623 );
and \U$415 ( \625 , \619 , \624 );
buf \U$416 ( \626 , \625 );
buf \U$417 ( \627 , \626 );
buf \U$418 ( \628 , RIc0d9f40_88);
buf \U$419 ( \629 , RIc0d9fb8_89);
xor \U$420 ( \630 , \628 , \629 );
buf \U$421 ( \631 , \630 );
buf \U$422 ( \632 , \631 );
not \U$423 ( \633 , \632 );
buf \U$424 ( \634 , \633 );
buf \U$425 ( \635 , \634 );
buf \U$426 ( \636 , RIc0d7ab0_10);
buf \U$427 ( \637 , RIc0d9ec8_87);
xnor \U$428 ( \638 , \636 , \637 );
buf \U$429 ( \639 , \638 );
buf \U$430 ( \640 , \639 );
nor \U$431 ( \641 , \635 , \640 );
buf \U$432 ( \642 , \641 );
buf \U$433 ( \643 , \642 );
nor \U$434 ( \644 , \627 , \643 );
buf \U$435 ( \645 , \644 );
buf \U$436 ( \646 , \645 );
xor \U$437 ( \647 , \592 , \646 );
buf \U$438 ( \648 , \647 );
buf \U$439 ( \649 , \648 );
and \U$440 ( \650 , \502 , \649 );
and \U$441 ( \651 , \366 , \501 );
or \U$442 ( \652 , \650 , \651 );
buf \U$443 ( \653 , \652 );
buf \U$444 ( \654 , \653 );
buf \U$445 ( \655 , RIc0d9478_65);
buf \U$446 ( \656 , RIc0d8578_33);
and \U$447 ( \657 , \655 , \656 );
buf \U$448 ( \658 , \657 );
buf \U$449 ( \659 , \658 );
buf \U$450 ( \660 , RIc0d8410_30);
buf \U$451 ( \661 , RIc0d9568_67);
xor \U$452 ( \662 , \660 , \661 );
buf \U$453 ( \663 , \662 );
buf \U$454 ( \664 , \663 );
not \U$455 ( \665 , \664 );
xor \U$456 ( \666 , RIc0d95e0_68, RIc0d9568_67);
buf \U$457 ( \667 , \666 );
buf \U$458 ( \668 , RIc0d95e0_68);
buf \U$459 ( \669 , RIc0d9658_69);
xnor \U$460 ( \670 , \668 , \669 );
buf \U$461 ( \671 , \670 );
buf \U$462 ( \672 , \671 );
nand \U$463 ( \673 , \667 , \672 );
buf \U$464 ( \674 , \673 );
buf \U$467 ( \675 , \674 );
buf \U$468 ( \676 , \675 );
not \U$469 ( \677 , \676 );
buf \U$470 ( \678 , \677 );
buf \U$471 ( \679 , \678 );
not \U$472 ( \680 , \679 );
or \U$473 ( \681 , \665 , \680 );
buf \U$474 ( \682 , RIc0d95e0_68);
buf \U$475 ( \683 , RIc0d9658_69);
xor \U$476 ( \684 , \682 , \683 );
buf \U$477 ( \685 , \684 );
buf \U$480 ( \686 , \685 );
buf \U$481 ( \687 , \686 );
buf \U$482 ( \688 , RIc0d9568_67);
buf \U$483 ( \689 , RIc0d8398_29);
xor \U$484 ( \690 , \688 , \689 );
buf \U$485 ( \691 , \690 );
buf \U$486 ( \692 , \691 );
nand \U$487 ( \693 , \687 , \692 );
buf \U$488 ( \694 , \693 );
buf \U$489 ( \695 , \694 );
nand \U$490 ( \696 , \681 , \695 );
buf \U$491 ( \697 , \696 );
buf \U$492 ( \698 , \697 );
xor \U$493 ( \699 , \659 , \698 );
buf \U$494 ( \700 , \538 );
not \U$495 ( \701 , \700 );
buf \U$496 ( \702 , \521 );
not \U$497 ( \703 , \702 );
buf \U$498 ( \704 , \703 );
buf \U$499 ( \705 , \704 );
not \U$500 ( \706 , \705 );
or \U$501 ( \707 , \701 , \706 );
buf \U$502 ( \708 , \512 );
not \U$503 ( \709 , \708 );
buf \U$504 ( \710 , \709 );
buf \U$507 ( \711 , \710 );
buf \U$508 ( \712 , \711 );
not \U$509 ( \713 , \712 );
buf \U$510 ( \714 , \713 );
buf \U$511 ( \715 , \714 );
buf \U$512 ( \716 , RIc0d7858_5);
buf \U$513 ( \717 , RIc0da0a8_91);
xor \U$514 ( \718 , \716 , \717 );
buf \U$515 ( \719 , \718 );
buf \U$516 ( \720 , \719 );
nand \U$517 ( \721 , \715 , \720 );
buf \U$518 ( \722 , \721 );
buf \U$519 ( \723 , \722 );
nand \U$520 ( \724 , \707 , \723 );
buf \U$521 ( \725 , \724 );
buf \U$522 ( \726 , \725 );
xor \U$523 ( \727 , \699 , \726 );
buf \U$524 ( \728 , \727 );
buf \U$525 ( \729 , \728 );
buf \U$526 ( \730 , RIc0da3f0_98);
buf \U$527 ( \731 , RIc0da468_99);
xor \U$528 ( \732 , \730 , \731 );
buf \U$529 ( \733 , \732 );
buf \U$532 ( \734 , \733 );
buf \U$533 ( \735 , \734 );
not \U$534 ( \736 , \735 );
buf \U$535 ( \737 , \736 );
buf \U$536 ( \738 , \737 );
not \U$537 ( \739 , \738 );
buf \U$538 ( \740 , RIc0da3f0_98);
buf \U$539 ( \741 , RIc0da468_99);
xnor \U$540 ( \742 , \740 , \741 );
buf \U$541 ( \743 , \742 );
buf \U$542 ( \744 , \743 );
xor \U$543 ( \745 , RIc0da3f0_98, RIc0da378_97);
buf \U$544 ( \746 , \745 );
nand \U$545 ( \747 , \744 , \746 );
buf \U$546 ( \748 , \747 );
buf \U$549 ( \749 , \748 );
buf \U$550 ( \750 , \749 );
not \U$551 ( \751 , \750 );
or \U$552 ( \752 , \739 , \751 );
buf \U$553 ( \753 , RIc0da378_97);
nand \U$554 ( \754 , \752 , \753 );
buf \U$555 ( \755 , \754 );
buf \U$556 ( \756 , \755 );
buf \U$557 ( \757 , RIc0d98b0_74);
buf \U$558 ( \758 , RIc0d9928_75);
and \U$559 ( \759 , \757 , \758 );
not \U$560 ( \760 , \757 );
buf \U$561 ( \761 , RIc0d9928_75);
not \U$562 ( \762 , \761 );
buf \U$563 ( \763 , \762 );
buf \U$564 ( \764 , \763 );
and \U$565 ( \765 , \760 , \764 );
or \U$566 ( \766 , \759 , \765 );
buf \U$567 ( \767 , \766 );
buf \U$568 ( \768 , \767 );
xor \U$569 ( \769 , RIc0d98b0_74, RIc0d9838_73);
buf \U$570 ( \770 , \769 );
nand \U$571 ( \771 , \768 , \770 );
buf \U$572 ( \772 , \771 );
buf \U$575 ( \773 , \772 );
buf \U$576 ( \774 , \773 );
not \U$577 ( \775 , \774 );
buf \U$578 ( \776 , \775 );
buf \U$579 ( \777 , \776 );
not \U$580 ( \778 , \777 );
buf \U$581 ( \779 , \778 );
buf \U$582 ( \780 , \779 );
buf \U$583 ( \781 , RIc0d8140_24);
buf \U$584 ( \782 , RIc0d9838_73);
xnor \U$585 ( \783 , \781 , \782 );
buf \U$586 ( \784 , \783 );
buf \U$587 ( \785 , \784 );
or \U$588 ( \786 , \780 , \785 );
buf \U$589 ( \787 , RIc0d98b0_74);
buf \U$590 ( \788 , RIc0d9928_75);
xor \U$591 ( \789 , \787 , \788 );
buf \U$592 ( \790 , \789 );
buf \U$595 ( \791 , \790 );
buf \U$598 ( \792 , \791 );
buf \U$599 ( \793 , \792 );
not \U$600 ( \794 , \793 );
buf \U$601 ( \795 , \794 );
buf \U$602 ( \796 , \795 );
buf \U$603 ( \797 , RIc0d80c8_23);
buf \U$604 ( \798 , RIc0d9838_73);
xnor \U$605 ( \799 , \797 , \798 );
buf \U$606 ( \800 , \799 );
buf \U$607 ( \801 , \800 );
or \U$608 ( \802 , \796 , \801 );
nand \U$609 ( \803 , \786 , \802 );
buf \U$610 ( \804 , \803 );
buf \U$611 ( \805 , \804 );
xor \U$612 ( \806 , \756 , \805 );
buf \U$613 ( \807 , \615 );
not \U$614 ( \808 , \807 );
buf \U$615 ( \809 , \808 );
buf \U$616 ( \810 , \809 );
not \U$617 ( \811 , \810 );
buf \U$618 ( \812 , \811 );
buf \U$619 ( \813 , \812 );
buf \U$620 ( \814 , \639 );
or \U$621 ( \815 , \813 , \814 );
buf \U$624 ( \816 , \631 );
buf \U$625 ( \817 , \816 );
not \U$626 ( \818 , \817 );
buf \U$627 ( \819 , \818 );
buf \U$628 ( \820 , \819 );
buf \U$629 ( \821 , RIc0d7a38_9);
buf \U$630 ( \822 , RIc0d9ec8_87);
xor \U$631 ( \823 , \821 , \822 );
buf \U$632 ( \824 , \823 );
buf \U$633 ( \825 , \824 );
not \U$634 ( \826 , \825 );
buf \U$635 ( \827 , \826 );
buf \U$636 ( \828 , \827 );
or \U$637 ( \829 , \820 , \828 );
nand \U$638 ( \830 , \815 , \829 );
buf \U$639 ( \831 , \830 );
buf \U$640 ( \832 , \831 );
xor \U$641 ( \833 , \806 , \832 );
buf \U$642 ( \834 , \833 );
buf \U$643 ( \835 , \834 );
xor \U$644 ( \836 , \729 , \835 );
buf \U$645 ( \837 , \447 );
not \U$646 ( \838 , \837 );
buf \U$647 ( \839 , \433 );
not \U$648 ( \840 , \839 );
buf \U$649 ( \841 , \840 );
buf \U$652 ( \842 , \841 );
buf \U$653 ( \843 , \842 );
not \U$654 ( \844 , \843 );
or \U$655 ( \845 , \838 , \844 );
buf \U$658 ( \846 , \441 );
buf \U$659 ( \847 , \846 );
buf \U$660 ( \848 , RIc0d7948_7);
buf \U$661 ( \849 , RIc0d9fb8_89);
xor \U$662 ( \850 , \848 , \849 );
buf \U$663 ( \851 , \850 );
buf \U$664 ( \852 , \851 );
nand \U$665 ( \853 , \847 , \852 );
buf \U$666 ( \854 , \853 );
buf \U$667 ( \855 , \854 );
nand \U$668 ( \856 , \845 , \855 );
buf \U$669 ( \857 , \856 );
buf \U$670 ( \858 , \857 );
buf \U$671 ( \859 , \289 );
not \U$672 ( \860 , \859 );
buf \U$675 ( \861 , \275 );
buf \U$676 ( \862 , \861 );
not \U$677 ( \863 , \862 );
buf \U$678 ( \864 , \863 );
buf \U$679 ( \865 , \864 );
not \U$680 ( \866 , \865 );
or \U$681 ( \867 , \860 , \866 );
buf \U$682 ( \868 , RIc0d9658_69);
buf \U$683 ( \869 , RIc0d82a8_27);
xnor \U$684 ( \870 , \868 , \869 );
buf \U$685 ( \871 , \870 );
buf \U$686 ( \872 , \871 );
not \U$687 ( \873 , \872 );
buf \U$690 ( \874 , \283 );
buf \U$691 ( \875 , \874 );
nand \U$692 ( \876 , \873 , \875 );
buf \U$693 ( \877 , \876 );
buf \U$694 ( \878 , \877 );
nand \U$695 ( \879 , \867 , \878 );
buf \U$696 ( \880 , \879 );
buf \U$697 ( \881 , \880 );
xor \U$698 ( \882 , \858 , \881 );
buf \U$699 ( \883 , \882 );
buf \U$700 ( \884 , \883 );
buf \U$701 ( \885 , \493 );
not \U$702 ( \886 , \885 );
buf \U$703 ( \887 , \473 );
not \U$704 ( \888 , \887 );
buf \U$705 ( \889 , \888 );
buf \U$706 ( \890 , \889 );
not \U$707 ( \891 , \890 );
or \U$708 ( \892 , \886 , \891 );
buf \U$709 ( \893 , \481 );
buf \U$710 ( \894 , RIc0d7768_3);
buf \U$711 ( \895 , RIc0da198_93);
xor \U$712 ( \896 , \894 , \895 );
buf \U$713 ( \897 , \896 );
buf \U$714 ( \898 , \897 );
nand \U$715 ( \899 , \893 , \898 );
buf \U$716 ( \900 , \899 );
buf \U$717 ( \901 , \900 );
nand \U$718 ( \902 , \892 , \901 );
buf \U$719 ( \903 , \902 );
buf \U$720 ( \904 , \903 );
xor \U$721 ( \905 , \884 , \904 );
buf \U$722 ( \906 , \905 );
buf \U$723 ( \907 , \906 );
xor \U$724 ( \908 , \836 , \907 );
buf \U$725 ( \909 , \908 );
buf \U$726 ( \910 , \909 );
xor \U$727 ( \911 , \654 , \910 );
buf \U$728 ( \912 , RIc0d9e50_86);
buf \U$729 ( \913 , RIc0d9ec8_87);
xor \U$730 ( \914 , \912 , \913 );
buf \U$731 ( \915 , \914 );
buf \U$732 ( \916 , \915 );
not \U$733 ( \917 , \916 );
buf \U$734 ( \918 , \917 );
buf \U$735 ( \919 , \918 );
not \U$736 ( \920 , \919 );
buf \U$737 ( \921 , \920 );
not \U$738 ( \922 , \921 );
buf \U$739 ( \923 , RIc0d7b28_11);
buf \U$740 ( \924 , RIc0d9dd8_85);
xor \U$741 ( \925 , \923 , \924 );
buf \U$742 ( \926 , \925 );
not \U$743 ( \927 , \926 );
or \U$744 ( \928 , \922 , \927 );
buf \U$745 ( \929 , RIc0d9e50_86);
not \U$746 ( \930 , \929 );
buf \U$747 ( \931 , RIc0d9dd8_85);
nand \U$748 ( \932 , \930 , \931 );
buf \U$749 ( \933 , \932 );
not \U$750 ( \934 , \933 );
buf \U$751 ( \935 , RIc0d9dd8_85);
not \U$752 ( \936 , \935 );
buf \U$753 ( \937 , RIc0d9e50_86);
nand \U$754 ( \938 , \936 , \937 );
buf \U$755 ( \939 , \938 );
not \U$756 ( \940 , \939 );
or \U$757 ( \941 , \934 , \940 );
buf \U$758 ( \942 , RIc0d9e50_86);
buf \U$759 ( \943 , RIc0d9ec8_87);
xnor \U$760 ( \944 , \942 , \943 );
buf \U$761 ( \945 , \944 );
nand \U$762 ( \946 , \941 , \945 );
buf \U$763 ( \947 , \946 );
buf \U$765 ( \948 , \947 );
buf \U$766 ( \949 , \948 );
not \U$767 ( \950 , \949 );
buf \U$768 ( \951 , \950 );
buf \U$769 ( \952 , \951 );
not \U$770 ( \953 , \952 );
buf \U$771 ( \954 , \953 );
buf \U$772 ( \955 , RIc0d7ba0_12);
buf \U$773 ( \956 , RIc0d9dd8_85);
xnor \U$774 ( \957 , \955 , \956 );
buf \U$775 ( \958 , \957 );
or \U$776 ( \959 , \954 , \958 );
nand \U$777 ( \960 , \928 , \959 );
buf \U$778 ( \961 , \960 );
buf \U$779 ( \962 , \356 );
not \U$780 ( \963 , \962 );
buf \U$781 ( \964 , \330 );
not \U$782 ( \965 , \964 );
or \U$783 ( \966 , \963 , \965 );
buf \U$784 ( \967 , \344 );
buf \U$785 ( \968 , RIc0da288_95);
buf \U$786 ( \969 , RIc0d7678_1);
and \U$787 ( \970 , \968 , \969 );
not \U$788 ( \971 , \968 );
buf \U$789 ( \972 , RIc0d7678_1);
not \U$790 ( \973 , \972 );
buf \U$791 ( \974 , \973 );
buf \U$792 ( \975 , \974 );
and \U$793 ( \976 , \971 , \975 );
nor \U$794 ( \977 , \970 , \976 );
buf \U$795 ( \978 , \977 );
buf \U$796 ( \979 , \978 );
nand \U$797 ( \980 , \967 , \979 );
buf \U$798 ( \981 , \980 );
buf \U$799 ( \982 , \981 );
nand \U$800 ( \983 , \966 , \982 );
buf \U$801 ( \984 , \983 );
buf \U$802 ( \985 , \984 );
xor \U$803 ( \986 , \961 , \985 );
buf \U$804 ( \987 , \574 );
not \U$805 ( \988 , \987 );
buf \U$806 ( \989 , \988 );
buf \U$807 ( \990 , \989 );
buf \U$808 ( \991 , \581 );
or \U$809 ( \992 , \990 , \991 );
buf \U$812 ( \993 , \558 );
buf \U$813 ( \994 , \993 );
not \U$814 ( \995 , \994 );
buf \U$815 ( \996 , \995 );
buf \U$816 ( \997 , \996 );
buf \U$817 ( \998 , RIc0d9ce8_83);
buf \U$818 ( \999 , RIc0d7c18_13);
not \U$819 ( \1000 , \999 );
buf \U$820 ( \1001 , \1000 );
buf \U$821 ( \1002 , \1001 );
and \U$822 ( \1003 , \998 , \1002 );
not \U$823 ( \1004 , \998 );
buf \U$824 ( \1005 , RIc0d7c18_13);
and \U$825 ( \1006 , \1004 , \1005 );
nor \U$826 ( \1007 , \1003 , \1006 );
buf \U$827 ( \1008 , \1007 );
buf \U$828 ( \1009 , \1008 );
or \U$829 ( \1010 , \997 , \1009 );
nand \U$830 ( \1011 , \992 , \1010 );
buf \U$831 ( \1012 , \1011 );
buf \U$832 ( \1013 , \1012 );
xor \U$833 ( \1014 , \986 , \1013 );
buf \U$834 ( \1015 , \1014 );
buf \U$835 ( \1016 , \1015 );
buf \U$836 ( \1017 , \408 );
not \U$837 ( \1018 , \1017 );
buf \U$838 ( \1019 , \393 );
not \U$839 ( \1020 , \1019 );
buf \U$840 ( \1021 , \1020 );
buf \U$841 ( \1022 , \1021 );
not \U$842 ( \1023 , \1022 );
or \U$843 ( \1024 , \1018 , \1023 );
buf \U$844 ( \1025 , \401 );
buf \U$845 ( \1026 , \1025 );
buf \U$846 ( \1027 , \1026 );
buf \U$847 ( \1028 , RIc0d7df8_17);
buf \U$848 ( \1029 , RIc0d9b08_79);
xor \U$849 ( \1030 , \1028 , \1029 );
buf \U$850 ( \1031 , \1030 );
buf \U$851 ( \1032 , \1031 );
nand \U$852 ( \1033 , \1027 , \1032 );
buf \U$853 ( \1034 , \1033 );
buf \U$854 ( \1035 , \1034 );
nand \U$855 ( \1036 , \1024 , \1035 );
buf \U$856 ( \1037 , \1036 );
buf \U$857 ( \1038 , RIc0d7d80_16);
buf \U$858 ( \1039 , RIc0d9bf8_81);
xor \U$859 ( \1040 , \1038 , \1039 );
buf \U$860 ( \1041 , \1040 );
buf \U$861 ( \1042 , \1041 );
not \U$862 ( \1043 , \1042 );
buf \U$863 ( \1044 , RIc0d9c70_82);
buf \U$864 ( \1045 , RIc0d9ce8_83);
and \U$865 ( \1046 , \1044 , \1045 );
not \U$866 ( \1047 , \1044 );
buf \U$867 ( \1048 , RIc0d9ce8_83);
not \U$868 ( \1049 , \1048 );
buf \U$869 ( \1050 , \1049 );
buf \U$870 ( \1051 , \1050 );
and \U$871 ( \1052 , \1047 , \1051 );
or \U$872 ( \1053 , \1046 , \1052 );
buf \U$873 ( \1054 , \1053 );
buf \U$874 ( \1055 , \1054 );
xor \U$875 ( \1056 , RIc0d9c70_82, RIc0d9bf8_81);
buf \U$876 ( \1057 , \1056 );
nand \U$877 ( \1058 , \1055 , \1057 );
buf \U$878 ( \1059 , \1058 );
buf \U$881 ( \1060 , \1059 );
buf \U$882 ( \1061 , \1060 );
not \U$883 ( \1062 , \1061 );
buf \U$884 ( \1063 , \1062 );
buf \U$887 ( \1064 , \1063 );
buf \U$888 ( \1065 , \1064 );
not \U$889 ( \1066 , \1065 );
or \U$890 ( \1067 , \1043 , \1066 );
buf \U$891 ( \1068 , RIc0d7d08_15);
buf \U$892 ( \1069 , RIc0d9bf8_81);
xnor \U$893 ( \1070 , \1068 , \1069 );
buf \U$894 ( \1071 , \1070 );
buf \U$895 ( \1072 , \1071 );
not \U$896 ( \1073 , \1072 );
buf \U$897 ( \1074 , RIc0d9c70_82);
buf \U$898 ( \1075 , RIc0d9ce8_83);
xor \U$899 ( \1076 , \1074 , \1075 );
buf \U$900 ( \1077 , \1076 );
buf \U$903 ( \1078 , \1077 );
buf \U$904 ( \1079 , \1078 );
nand \U$905 ( \1080 , \1073 , \1079 );
buf \U$906 ( \1081 , \1080 );
buf \U$907 ( \1082 , \1081 );
nand \U$908 ( \1083 , \1067 , \1082 );
buf \U$909 ( \1084 , \1083 );
xor \U$910 ( \1085 , \1037 , \1084 );
buf \U$911 ( \1086 , RIc0d8050_22);
buf \U$912 ( \1087 , RIc0d9928_75);
xor \U$913 ( \1088 , \1086 , \1087 );
buf \U$914 ( \1089 , \1088 );
buf \U$915 ( \1090 , \1089 );
not \U$916 ( \1091 , \1090 );
buf \U$917 ( \1092 , RIc0d99a0_76);
not \U$918 ( \1093 , \1092 );
buf \U$919 ( \1094 , RIc0d9928_75);
nand \U$920 ( \1095 , \1093 , \1094 );
buf \U$921 ( \1096 , \1095 );
buf \U$922 ( \1097 , \1096 );
buf \U$923 ( \1098 , RIc0d9928_75);
not \U$924 ( \1099 , \1098 );
buf \U$925 ( \1100 , RIc0d99a0_76);
nand \U$926 ( \1101 , \1099 , \1100 );
buf \U$927 ( \1102 , \1101 );
buf \U$928 ( \1103 , \1102 );
nand \U$929 ( \1104 , \1097 , \1103 );
buf \U$930 ( \1105 , \1104 );
buf \U$931 ( \1106 , \1105 );
buf \U$932 ( \1107 , RIc0d99a0_76);
buf \U$933 ( \1108 , RIc0d9a18_77);
and \U$934 ( \1109 , \1107 , \1108 );
not \U$935 ( \1110 , \1107 );
buf \U$936 ( \1111 , RIc0d9a18_77);
not \U$937 ( \1112 , \1111 );
buf \U$938 ( \1113 , \1112 );
buf \U$939 ( \1114 , \1113 );
and \U$940 ( \1115 , \1110 , \1114 );
nor \U$941 ( \1116 , \1109 , \1115 );
buf \U$942 ( \1117 , \1116 );
buf \U$943 ( \1118 , \1117 );
not \U$944 ( \1119 , \1118 );
buf \U$945 ( \1120 , \1119 );
buf \U$946 ( \1121 , \1120 );
nand \U$947 ( \1122 , \1106 , \1121 );
buf \U$948 ( \1123 , \1122 );
buf \U$951 ( \1124 , \1123 );
buf \U$954 ( \1125 , \1124 );
buf \U$957 ( \1126 , \1125 );
buf \U$958 ( \1127 , \1126 );
not \U$959 ( \1128 , \1127 );
buf \U$960 ( \1129 , \1128 );
buf \U$961 ( \1130 , \1129 );
not \U$962 ( \1131 , \1130 );
or \U$963 ( \1132 , \1091 , \1131 );
buf \U$964 ( \1133 , RIc0d7fd8_21);
buf \U$965 ( \1134 , RIc0d9928_75);
xnor \U$966 ( \1135 , \1133 , \1134 );
buf \U$967 ( \1136 , \1135 );
buf \U$968 ( \1137 , \1136 );
not \U$969 ( \1138 , \1137 );
buf \U$970 ( \1139 , RIc0d99a0_76);
buf \U$971 ( \1140 , RIc0d9a18_77);
xor \U$972 ( \1141 , \1139 , \1140 );
buf \U$973 ( \1142 , \1141 );
buf \U$976 ( \1143 , \1142 );
buf \U$977 ( \1144 , \1143 );
nand \U$978 ( \1145 , \1138 , \1144 );
buf \U$979 ( \1146 , \1145 );
buf \U$980 ( \1147 , \1146 );
nand \U$981 ( \1148 , \1132 , \1147 );
buf \U$982 ( \1149 , \1148 );
xnor \U$983 ( \1150 , \1085 , \1149 );
buf \U$984 ( \1151 , \1150 );
not \U$985 ( \1152 , \1151 );
buf \U$986 ( \1153 , \1152 );
buf \U$987 ( \1154 , \1153 );
and \U$988 ( \1155 , \1016 , \1154 );
not \U$989 ( \1156 , \1016 );
buf \U$990 ( \1157 , \1150 );
and \U$991 ( \1158 , \1156 , \1157 );
nor \U$992 ( \1159 , \1155 , \1158 );
buf \U$993 ( \1160 , \1159 );
buf \U$994 ( \1161 , \1160 );
buf \U$995 ( \1162 , RIc0d7f60_20);
buf \U$996 ( \1163 , RIc0d9a18_77);
xor \U$997 ( \1164 , \1162 , \1163 );
buf \U$998 ( \1165 , \1164 );
buf \U$999 ( \1166 , \1165 );
not \U$1000 ( \1167 , \1166 );
buf \U$1001 ( \1168 , RIc0d9a90_78);
buf \U$1002 ( \1169 , RIc0d9b08_79);
xor \U$1003 ( \1170 , \1168 , \1169 );
buf \U$1004 ( \1171 , \1170 );
buf \U$1005 ( \1172 , \1171 );
not \U$1006 ( \1173 , \1172 );
buf \U$1007 ( \1174 , \1173 );
buf \U$1008 ( \1175 , \1174 );
xor \U$1009 ( \1176 , RIc0d9a90_78, RIc0d9a18_77);
buf \U$1010 ( \1177 , \1176 );
nand \U$1011 ( \1178 , \1175 , \1177 );
buf \U$1012 ( \1179 , \1178 );
buf \U$1013 ( \1180 , \1179 );
not \U$1014 ( \1181 , \1180 );
buf \U$1015 ( \1182 , \1181 );
buf \U$1018 ( \1183 , \1182 );
buf \U$1019 ( \1184 , \1183 );
not \U$1020 ( \1185 , \1184 );
or \U$1021 ( \1186 , \1167 , \1185 );
buf \U$1022 ( \1187 , RIc0d9a18_77);
buf \U$1023 ( \1188 , RIc0d7ee8_19);
xnor \U$1024 ( \1189 , \1187 , \1188 );
buf \U$1025 ( \1190 , \1189 );
buf \U$1026 ( \1191 , \1190 );
not \U$1027 ( \1192 , \1191 );
buf \U$1030 ( \1193 , \1174 );
buf \U$1031 ( \1194 , \1193 );
not \U$1032 ( \1195 , \1194 );
buf \U$1033 ( \1196 , \1195 );
buf \U$1034 ( \1197 , \1196 );
nand \U$1035 ( \1198 , \1192 , \1197 );
buf \U$1036 ( \1199 , \1198 );
buf \U$1037 ( \1200 , \1199 );
nand \U$1038 ( \1201 , \1186 , \1200 );
buf \U$1039 ( \1202 , \1201 );
buf \U$1040 ( \1203 , RIc0d9478_65);
buf \U$1041 ( \1204 , RIc0d8500_32);
xor \U$1042 ( \1205 , \1203 , \1204 );
buf \U$1043 ( \1206 , \1205 );
buf \U$1044 ( \1207 , \1206 );
not \U$1045 ( \1208 , \1207 );
buf \U$1046 ( \1209 , RIc0d94f0_66);
buf \U$1047 ( \1210 , RIc0d9568_67);
xor \U$1048 ( \1211 , \1209 , \1210 );
buf \U$1049 ( \1212 , \1211 );
buf \U$1050 ( \1213 , \1212 );
not \U$1051 ( \1214 , \1213 );
buf \U$1052 ( \1215 , \1214 );
buf \U$1053 ( \1216 , \1215 );
xor \U$1054 ( \1217 , RIc0d9478_65, RIc0d94f0_66);
buf \U$1055 ( \1218 , \1217 );
nand \U$1056 ( \1219 , \1216 , \1218 );
buf \U$1057 ( \1220 , \1219 );
buf \U$1060 ( \1221 , \1220 );
buf \U$1061 ( \1222 , \1221 );
not \U$1062 ( \1223 , \1222 );
buf \U$1063 ( \1224 , \1223 );
buf \U$1066 ( \1225 , \1224 );
buf \U$1067 ( \1226 , \1225 );
not \U$1068 ( \1227 , \1226 );
or \U$1069 ( \1228 , \1208 , \1227 );
buf \U$1072 ( \1229 , \1212 );
buf \U$1073 ( \1230 , \1229 );
not \U$1074 ( \1231 , \1230 );
buf \U$1075 ( \1232 , \1231 );
buf \U$1076 ( \1233 , \1232 );
not \U$1077 ( \1234 , \1233 );
buf \U$1078 ( \1235 , \1234 );
buf \U$1079 ( \1236 , \1235 );
buf \U$1080 ( \1237 , RIc0d9478_65);
buf \U$1081 ( \1238 , RIc0d8488_31);
xor \U$1082 ( \1239 , \1237 , \1238 );
buf \U$1083 ( \1240 , \1239 );
buf \U$1084 ( \1241 , \1240 );
nand \U$1085 ( \1242 , \1236 , \1241 );
buf \U$1086 ( \1243 , \1242 );
buf \U$1087 ( \1244 , \1243 );
nand \U$1088 ( \1245 , \1228 , \1244 );
buf \U$1089 ( \1246 , \1245 );
xor \U$1090 ( \1247 , \1202 , \1246 );
buf \U$1091 ( \1248 , RIc0d8230_26);
buf \U$1092 ( \1249 , RIc0d9748_71);
xor \U$1093 ( \1250 , \1248 , \1249 );
buf \U$1094 ( \1251 , \1250 );
buf \U$1095 ( \1252 , \1251 );
not \U$1096 ( \1253 , \1252 );
xnor \U$1097 ( \1254 , RIc0d97c0_72, RIc0d9838_73);
buf \U$1098 ( \1255 , \1254 );
xor \U$1099 ( \1256 , RIc0d9748_71, RIc0d97c0_72);
buf \U$1100 ( \1257 , \1256 );
nand \U$1101 ( \1258 , \1255 , \1257 );
buf \U$1102 ( \1259 , \1258 );
buf \U$1105 ( \1260 , \1259 );
buf \U$1106 ( \1261 , \1260 );
not \U$1107 ( \1262 , \1261 );
buf \U$1108 ( \1263 , \1262 );
buf \U$1109 ( \1264 , \1263 );
not \U$1110 ( \1265 , \1264 );
or \U$1111 ( \1266 , \1253 , \1265 );
buf \U$1112 ( \1267 , RIc0d81b8_25);
buf \U$1113 ( \1268 , RIc0d9748_71);
xnor \U$1114 ( \1269 , \1267 , \1268 );
buf \U$1115 ( \1270 , \1269 );
buf \U$1116 ( \1271 , \1270 );
not \U$1117 ( \1272 , \1271 );
buf \U$1118 ( \1273 , RIc0d97c0_72);
buf \U$1119 ( \1274 , RIc0d9838_73);
xor \U$1120 ( \1275 , \1273 , \1274 );
buf \U$1121 ( \1276 , \1275 );
buf \U$1122 ( \1277 , \1276 );
not \U$1123 ( \1278 , \1277 );
buf \U$1124 ( \1279 , \1278 );
buf \U$1125 ( \1280 , \1279 );
not \U$1126 ( \1281 , \1280 );
buf \U$1127 ( \1282 , \1281 );
buf \U$1128 ( \1283 , \1282 );
nand \U$1129 ( \1284 , \1272 , \1283 );
buf \U$1130 ( \1285 , \1284 );
buf \U$1131 ( \1286 , \1285 );
nand \U$1132 ( \1287 , \1266 , \1286 );
buf \U$1133 ( \1288 , \1287 );
xnor \U$1134 ( \1289 , \1247 , \1288 );
buf \U$1135 ( \1290 , \1289 );
not \U$1136 ( \1291 , \1290 );
buf \U$1137 ( \1292 , \1291 );
buf \U$1138 ( \1293 , \1292 );
and \U$1139 ( \1294 , \1161 , \1293 );
not \U$1140 ( \1295 , \1161 );
buf \U$1141 ( \1296 , \1289 );
and \U$1142 ( \1297 , \1295 , \1296 );
nor \U$1143 ( \1298 , \1294 , \1297 );
buf \U$1144 ( \1299 , \1298 );
buf \U$1145 ( \1300 , \1299 );
and \U$1146 ( \1301 , \911 , \1300 );
and \U$1147 ( \1302 , \654 , \910 );
or \U$1148 ( \1303 , \1301 , \1302 );
buf \U$1149 ( \1304 , \1303 );
buf \U$1150 ( \1305 , \1304 );
xor \U$1151 ( \1306 , \659 , \698 );
and \U$1152 ( \1307 , \1306 , \726 );
and \U$1153 ( \1308 , \659 , \698 );
or \U$1154 ( \1309 , \1307 , \1308 );
buf \U$1155 ( \1310 , \1309 );
buf \U$1156 ( \1311 , \1310 );
buf \U$1157 ( \1312 , \857 );
buf \U$1158 ( \1313 , \880 );
or \U$1159 ( \1314 , \1312 , \1313 );
buf \U$1160 ( \1315 , \903 );
nand \U$1161 ( \1316 , \1314 , \1315 );
buf \U$1162 ( \1317 , \1316 );
buf \U$1163 ( \1318 , \1317 );
buf \U$1164 ( \1319 , \857 );
buf \U$1165 ( \1320 , \880 );
nand \U$1166 ( \1321 , \1319 , \1320 );
buf \U$1167 ( \1322 , \1321 );
buf \U$1168 ( \1323 , \1322 );
nand \U$1169 ( \1324 , \1318 , \1323 );
buf \U$1170 ( \1325 , \1324 );
buf \U$1171 ( \1326 , \1325 );
xor \U$1172 ( \1327 , \1311 , \1326 );
xor \U$1173 ( \1328 , \756 , \805 );
and \U$1174 ( \1329 , \1328 , \832 );
and \U$1175 ( \1330 , \756 , \805 );
or \U$1176 ( \1331 , \1329 , \1330 );
buf \U$1177 ( \1332 , \1331 );
buf \U$1178 ( \1333 , \1332 );
xor \U$1179 ( \1334 , \1327 , \1333 );
buf \U$1180 ( \1335 , \1334 );
buf \U$1181 ( \1336 , \1335 );
xor \U$1182 ( \1337 , \729 , \835 );
and \U$1183 ( \1338 , \1337 , \907 );
and \U$1184 ( \1339 , \729 , \835 );
or \U$1185 ( \1340 , \1338 , \1339 );
buf \U$1186 ( \1341 , \1340 );
buf \U$1187 ( \1342 , \1341 );
xor \U$1188 ( \1343 , \1336 , \1342 );
and \U$1189 ( \1344 , \1203 , \1204 );
buf \U$1190 ( \1345 , \1344 );
buf \U$1191 ( \1346 , \1345 );
buf \U$1192 ( \1347 , \1031 );
not \U$1193 ( \1348 , \1347 );
buf \U$1194 ( \1349 , \393 );
not \U$1195 ( \1350 , \1349 );
buf \U$1196 ( \1351 , \1350 );
buf \U$1197 ( \1352 , \1351 );
not \U$1198 ( \1353 , \1352 );
or \U$1199 ( \1354 , \1348 , \1353 );
buf \U$1200 ( \1355 , \1026 );
xor \U$1201 ( \1356 , RIc0d9b08_79, RIc0d7d80_16);
buf \U$1202 ( \1357 , \1356 );
nand \U$1203 ( \1358 , \1355 , \1357 );
buf \U$1204 ( \1359 , \1358 );
buf \U$1205 ( \1360 , \1359 );
nand \U$1206 ( \1361 , \1354 , \1360 );
buf \U$1207 ( \1362 , \1361 );
buf \U$1208 ( \1363 , \1362 );
xor \U$1209 ( \1364 , \1346 , \1363 );
buf \U$1210 ( \1365 , \1124 );
buf \U$1211 ( \1366 , \1136 );
or \U$1212 ( \1367 , \1365 , \1366 );
buf \U$1213 ( \1368 , \1143 );
not \U$1214 ( \1369 , \1368 );
buf \U$1215 ( \1370 , \1369 );
buf \U$1216 ( \1371 , \1370 );
buf \U$1217 ( \1372 , RIc0d7f60_20);
buf \U$1218 ( \1373 , RIc0d9928_75);
xnor \U$1219 ( \1374 , \1372 , \1373 );
buf \U$1220 ( \1375 , \1374 );
buf \U$1221 ( \1376 , \1375 );
or \U$1222 ( \1377 , \1371 , \1376 );
nand \U$1223 ( \1378 , \1367 , \1377 );
buf \U$1224 ( \1379 , \1378 );
buf \U$1225 ( \1380 , \1379 );
xor \U$1226 ( \1381 , \1364 , \1380 );
buf \U$1227 ( \1382 , \1381 );
buf \U$1228 ( \1383 , \1382 );
buf \U$1229 ( \1384 , \926 );
not \U$1230 ( \1385 , \1384 );
buf \U$1231 ( \1386 , \948 );
not \U$1232 ( \1387 , \1386 );
buf \U$1233 ( \1388 , \1387 );
buf \U$1236 ( \1389 , \1388 );
buf \U$1237 ( \1390 , \1389 );
not \U$1238 ( \1391 , \1390 );
or \U$1239 ( \1392 , \1385 , \1391 );
buf \U$1240 ( \1393 , RIc0d9dd8_85);
buf \U$1241 ( \1394 , RIc0d7ab0_10);
xnor \U$1242 ( \1395 , \1393 , \1394 );
buf \U$1243 ( \1396 , \1395 );
buf \U$1244 ( \1397 , \1396 );
not \U$1245 ( \1398 , \1397 );
buf \U$1246 ( \1399 , \918 );
not \U$1247 ( \1400 , \1399 );
buf \U$1248 ( \1401 , \1400 );
buf \U$1249 ( \1402 , \1401 );
nand \U$1250 ( \1403 , \1398 , \1402 );
buf \U$1251 ( \1404 , \1403 );
buf \U$1252 ( \1405 , \1404 );
nand \U$1253 ( \1406 , \1392 , \1405 );
buf \U$1254 ( \1407 , \1406 );
buf \U$1255 ( \1408 , \1407 );
xor \U$1256 ( \1409 , RIc0d9568_67, RIc0d8320_28);
and \U$1257 ( \1410 , \686 , \1409 );
not \U$1258 ( \1411 , \691 );
buf \U$1259 ( \1412 , \675 );
not \U$1260 ( \1413 , \1412 );
buf \U$1261 ( \1414 , \1413 );
buf \U$1262 ( \1415 , \1414 );
not \U$1263 ( \1416 , \1415 );
buf \U$1264 ( \1417 , \1416 );
nor \U$1265 ( \1418 , \1411 , \1417 );
nor \U$1266 ( \1419 , \1410 , \1418 );
buf \U$1267 ( \1420 , \1419 );
not \U$1268 ( \1421 , \1420 );
buf \U$1269 ( \1422 , \1421 );
buf \U$1270 ( \1423 , \1422 );
and \U$1271 ( \1424 , \1408 , \1423 );
not \U$1272 ( \1425 , \1408 );
buf \U$1273 ( \1426 , \1419 );
and \U$1274 ( \1427 , \1425 , \1426 );
nor \U$1275 ( \1428 , \1424 , \1427 );
buf \U$1276 ( \1429 , \1428 );
buf \U$1277 ( \1430 , \1429 );
buf \U$1280 ( \1431 , \1182 );
buf \U$1283 ( \1432 , \1431 );
buf \U$1284 ( \1433 , \1432 );
not \U$1285 ( \1434 , \1433 );
buf \U$1286 ( \1435 , \1434 );
buf \U$1287 ( \1436 , \1435 );
buf \U$1288 ( \1437 , \1190 );
or \U$1289 ( \1438 , \1436 , \1437 );
buf \U$1290 ( \1439 , \1193 );
xnor \U$1291 ( \1440 , RIc0d9a18_77, RIc0d7e70_18);
buf \U$1292 ( \1441 , \1440 );
or \U$1293 ( \1442 , \1439 , \1441 );
nand \U$1294 ( \1443 , \1438 , \1442 );
buf \U$1295 ( \1444 , \1443 );
buf \U$1296 ( \1445 , \1444 );
xor \U$1297 ( \1446 , \1430 , \1445 );
buf \U$1298 ( \1447 , \1446 );
buf \U$1299 ( \1448 , \1447 );
xor \U$1300 ( \1449 , \1383 , \1448 );
buf \U$1301 ( \1450 , \279 );
not \U$1302 ( \1451 , \1450 );
buf \U$1303 ( \1452 , \1451 );
not \U$1304 ( \1453 , \1452 );
not \U$1305 ( \1454 , \871 );
and \U$1306 ( \1455 , \1453 , \1454 );
buf \U$1307 ( \1456 , RIc0d8230_26);
buf \U$1308 ( \1457 , RIc0d9658_69);
xor \U$1309 ( \1458 , \1456 , \1457 );
buf \U$1310 ( \1459 , \1458 );
and \U$1311 ( \1460 , \284 , \1459 );
nor \U$1312 ( \1461 , \1455 , \1460 );
buf \U$1313 ( \1462 , \1461 );
not \U$1314 ( \1463 , \1462 );
buf \U$1315 ( \1464 , \1463 );
buf \U$1316 ( \1465 , \1464 );
not \U$1317 ( \1466 , \1465 );
buf \U$1318 ( \1467 , \851 );
not \U$1319 ( \1468 , \1467 );
buf \U$1320 ( \1469 , \842 );
not \U$1321 ( \1470 , \1469 );
or \U$1322 ( \1471 , \1468 , \1470 );
buf \U$1323 ( \1472 , \846 );
buf \U$1324 ( \1473 , RIc0d78d0_6);
buf \U$1325 ( \1474 , RIc0d9fb8_89);
xor \U$1326 ( \1475 , \1473 , \1474 );
buf \U$1327 ( \1476 , \1475 );
buf \U$1328 ( \1477 , \1476 );
nand \U$1329 ( \1478 , \1472 , \1477 );
buf \U$1330 ( \1479 , \1478 );
buf \U$1331 ( \1480 , \1479 );
nand \U$1332 ( \1481 , \1471 , \1480 );
buf \U$1333 ( \1482 , \1481 );
buf \U$1334 ( \1483 , \1482 );
not \U$1335 ( \1484 , \1483 );
buf \U$1336 ( \1485 , \1484 );
buf \U$1337 ( \1486 , \1485 );
buf \U$1338 ( \1487 , \897 );
not \U$1339 ( \1488 , \1487 );
buf \U$1340 ( \1489 , \476 );
not \U$1341 ( \1490 , \1489 );
or \U$1342 ( \1491 , \1488 , \1490 );
buf \U$1343 ( \1492 , \481 );
buf \U$1344 ( \1493 , RIc0da198_93);
buf \U$1345 ( \1494 , RIc0d76f0_2);
and \U$1346 ( \1495 , \1493 , \1494 );
not \U$1347 ( \1496 , \1493 );
buf \U$1348 ( \1497 , \352 );
and \U$1349 ( \1498 , \1496 , \1497 );
nor \U$1350 ( \1499 , \1495 , \1498 );
buf \U$1351 ( \1500 , \1499 );
buf \U$1352 ( \1501 , \1500 );
nand \U$1353 ( \1502 , \1492 , \1501 );
buf \U$1354 ( \1503 , \1502 );
buf \U$1355 ( \1504 , \1503 );
nand \U$1356 ( \1505 , \1491 , \1504 );
buf \U$1357 ( \1506 , \1505 );
buf \U$1358 ( \1507 , \1506 );
xor \U$1359 ( \1508 , \1486 , \1507 );
buf \U$1360 ( \1509 , \1508 );
buf \U$1361 ( \1510 , \1509 );
not \U$1362 ( \1511 , \1510 );
or \U$1363 ( \1512 , \1466 , \1511 );
buf \U$1364 ( \1513 , \1509 );
buf \U$1365 ( \1514 , \1464 );
or \U$1366 ( \1515 , \1513 , \1514 );
nand \U$1367 ( \1516 , \1512 , \1515 );
buf \U$1368 ( \1517 , \1516 );
buf \U$1369 ( \1518 , \1517 );
xor \U$1370 ( \1519 , \1449 , \1518 );
buf \U$1371 ( \1520 , \1519 );
buf \U$1372 ( \1521 , \1520 );
xor \U$1373 ( \1522 , \1343 , \1521 );
buf \U$1374 ( \1523 , \1522 );
buf \U$1375 ( \1524 , \1523 );
xor \U$1376 ( \1525 , \1305 , \1524 );
xor \U$1377 ( \1526 , \250 , \296 );
and \U$1378 ( \1527 , \1526 , \363 );
and \U$1379 ( \1528 , \250 , \296 );
or \U$1380 ( \1529 , \1527 , \1528 );
buf \U$1381 ( \1530 , \1529 );
buf \U$1382 ( \1531 , \1530 );
buf \U$1383 ( \1532 , \414 );
not \U$1384 ( \1533 , \1532 );
buf \U$1385 ( \1534 , \453 );
not \U$1386 ( \1535 , \1534 );
or \U$1387 ( \1536 , \1533 , \1535 );
buf \U$1388 ( \1537 , \453 );
buf \U$1389 ( \1538 , \414 );
or \U$1390 ( \1539 , \1537 , \1538 );
buf \U$1391 ( \1540 , \499 );
nand \U$1392 ( \1541 , \1539 , \1540 );
buf \U$1393 ( \1542 , \1541 );
buf \U$1394 ( \1543 , \1542 );
nand \U$1395 ( \1544 , \1536 , \1543 );
buf \U$1396 ( \1545 , \1544 );
buf \U$1397 ( \1546 , \1545 );
xor \U$1398 ( \1547 , \1531 , \1546 );
buf \U$1399 ( \1548 , RIc0d80c8_23);
buf \U$1400 ( \1549 , RIc0d9928_75);
xor \U$1401 ( \1550 , \1548 , \1549 );
buf \U$1402 ( \1551 , \1550 );
buf \U$1403 ( \1552 , \1551 );
not \U$1404 ( \1553 , \1552 );
buf \U$1405 ( \1554 , \1124 );
not \U$1406 ( \1555 , \1554 );
buf \U$1407 ( \1556 , \1555 );
buf \U$1408 ( \1557 , \1556 );
not \U$1409 ( \1558 , \1557 );
or \U$1410 ( \1559 , \1553 , \1558 );
buf \U$1411 ( \1560 , \1142 );
not \U$1412 ( \1561 , \1560 );
buf \U$1413 ( \1562 , \1561 );
buf \U$1414 ( \1563 , \1562 );
not \U$1415 ( \1564 , \1563 );
buf \U$1416 ( \1565 , \1564 );
buf \U$1417 ( \1566 , \1565 );
buf \U$1418 ( \1567 , \1089 );
nand \U$1419 ( \1568 , \1566 , \1567 );
buf \U$1420 ( \1569 , \1568 );
buf \U$1421 ( \1570 , \1569 );
nand \U$1422 ( \1571 , \1559 , \1570 );
buf \U$1423 ( \1572 , \1571 );
buf \U$1424 ( \1573 , \1572 );
buf \U$1425 ( \1574 , RIc0d7fd8_21);
buf \U$1426 ( \1575 , RIc0d9a18_77);
xor \U$1427 ( \1576 , \1574 , \1575 );
buf \U$1428 ( \1577 , \1576 );
buf \U$1429 ( \1578 , \1577 );
not \U$1430 ( \1579 , \1578 );
buf \U$1431 ( \1580 , \1183 );
not \U$1432 ( \1581 , \1580 );
or \U$1433 ( \1582 , \1579 , \1581 );
buf \U$1434 ( \1583 , \1171 );
not \U$1435 ( \1584 , \1583 );
buf \U$1436 ( \1585 , \1584 );
buf \U$1437 ( \1586 , \1585 );
not \U$1438 ( \1587 , \1586 );
buf \U$1439 ( \1588 , \1587 );
buf \U$1440 ( \1589 , \1588 );
buf \U$1441 ( \1590 , \1165 );
nand \U$1442 ( \1591 , \1589 , \1590 );
buf \U$1443 ( \1592 , \1591 );
buf \U$1444 ( \1593 , \1592 );
nand \U$1445 ( \1594 , \1582 , \1593 );
buf \U$1446 ( \1595 , \1594 );
buf \U$1447 ( \1596 , \1595 );
xor \U$1448 ( \1597 , \1573 , \1596 );
buf \U$1449 ( \1598 , \1063 );
not \U$1450 ( \1599 , \1598 );
buf \U$1451 ( \1600 , \1599 );
buf \U$1452 ( \1601 , \1600 );
buf \U$1453 ( \1602 , RIc0d7df8_17);
buf \U$1454 ( \1603 , RIc0d9bf8_81);
xnor \U$1455 ( \1604 , \1602 , \1603 );
buf \U$1456 ( \1605 , \1604 );
buf \U$1457 ( \1606 , \1605 );
or \U$1458 ( \1607 , \1601 , \1606 );
buf \U$1459 ( \1608 , \1078 );
not \U$1460 ( \1609 , \1608 );
buf \U$1461 ( \1610 , \1609 );
buf \U$1462 ( \1611 , \1610 );
buf \U$1463 ( \1612 , \1041 );
not \U$1464 ( \1613 , \1612 );
buf \U$1465 ( \1614 , \1613 );
buf \U$1466 ( \1615 , \1614 );
or \U$1467 ( \1616 , \1611 , \1615 );
nand \U$1468 ( \1617 , \1607 , \1616 );
buf \U$1469 ( \1618 , \1617 );
buf \U$1470 ( \1619 , \1618 );
and \U$1471 ( \1620 , \1597 , \1619 );
and \U$1472 ( \1621 , \1573 , \1596 );
or \U$1473 ( \1622 , \1620 , \1621 );
buf \U$1474 ( \1623 , \1622 );
buf \U$1475 ( \1624 , \1623 );
and \U$1476 ( \1625 , \1547 , \1624 );
and \U$1477 ( \1626 , \1531 , \1546 );
or \U$1478 ( \1627 , \1625 , \1626 );
buf \U$1479 ( \1628 , \1627 );
buf \U$1480 ( \1629 , \1628 );
buf \U$1481 ( \1630 , \1292 );
not \U$1482 ( \1631 , \1630 );
buf \U$1483 ( \1632 , \1153 );
not \U$1484 ( \1633 , \1632 );
or \U$1485 ( \1634 , \1631 , \1633 );
buf \U$1486 ( \1635 , \1289 );
not \U$1487 ( \1636 , \1635 );
buf \U$1488 ( \1637 , \1150 );
not \U$1489 ( \1638 , \1637 );
or \U$1490 ( \1639 , \1636 , \1638 );
buf \U$1491 ( \1640 , \1015 );
nand \U$1492 ( \1641 , \1639 , \1640 );
buf \U$1493 ( \1642 , \1641 );
buf \U$1494 ( \1643 , \1642 );
nand \U$1495 ( \1644 , \1634 , \1643 );
buf \U$1496 ( \1645 , \1644 );
buf \U$1497 ( \1646 , \1645 );
xor \U$1498 ( \1647 , \1629 , \1646 );
buf \U$1499 ( \1648 , \1037 );
not \U$1500 ( \1649 , \1648 );
buf \U$1501 ( \1650 , \1084 );
not \U$1502 ( \1651 , \1650 );
or \U$1503 ( \1652 , \1649 , \1651 );
buf \U$1504 ( \1653 , \1084 );
buf \U$1505 ( \1654 , \1037 );
or \U$1506 ( \1655 , \1653 , \1654 );
buf \U$1507 ( \1656 , \1149 );
nand \U$1508 ( \1657 , \1655 , \1656 );
buf \U$1509 ( \1658 , \1657 );
buf \U$1510 ( \1659 , \1658 );
nand \U$1511 ( \1660 , \1652 , \1659 );
buf \U$1512 ( \1661 , \1660 );
buf \U$1513 ( \1662 , \1661 );
xor \U$1514 ( \1663 , \961 , \985 );
and \U$1515 ( \1664 , \1663 , \1013 );
and \U$1516 ( \1665 , \961 , \985 );
or \U$1517 ( \1666 , \1664 , \1665 );
buf \U$1518 ( \1667 , \1666 );
buf \U$1519 ( \1668 , \1667 );
xor \U$1520 ( \1669 , \1662 , \1668 );
buf \U$1521 ( \1670 , \800 );
not \U$1522 ( \1671 , \1670 );
buf \U$1523 ( \1672 , \1671 );
buf \U$1524 ( \1673 , \1672 );
not \U$1525 ( \1674 , \1673 );
buf \U$1526 ( \1675 , \773 );
not \U$1527 ( \1676 , \1675 );
buf \U$1528 ( \1677 , \1676 );
buf \U$1529 ( \1678 , \1677 );
not \U$1530 ( \1679 , \1678 );
or \U$1531 ( \1680 , \1674 , \1679 );
buf \U$1532 ( \1681 , \792 );
buf \U$1533 ( \1682 , RIc0d8050_22);
buf \U$1534 ( \1683 , RIc0d9838_73);
xor \U$1535 ( \1684 , \1682 , \1683 );
buf \U$1536 ( \1685 , \1684 );
buf \U$1537 ( \1686 , \1685 );
nand \U$1538 ( \1687 , \1681 , \1686 );
buf \U$1539 ( \1688 , \1687 );
buf \U$1540 ( \1689 , \1688 );
nand \U$1541 ( \1690 , \1680 , \1689 );
buf \U$1542 ( \1691 , \1690 );
buf \U$1543 ( \1692 , \1240 );
not \U$1544 ( \1693 , \1692 );
buf \U$1545 ( \1694 , \1225 );
not \U$1546 ( \1695 , \1694 );
or \U$1547 ( \1696 , \1693 , \1695 );
buf \U$1548 ( \1697 , RIc0d8410_30);
buf \U$1549 ( \1698 , RIc0d9478_65);
xnor \U$1550 ( \1699 , \1697 , \1698 );
buf \U$1551 ( \1700 , \1699 );
buf \U$1552 ( \1701 , \1700 );
not \U$1553 ( \1702 , \1701 );
buf \U$1554 ( \1703 , \1232 );
not \U$1555 ( \1704 , \1703 );
buf \U$1556 ( \1705 , \1704 );
buf \U$1557 ( \1706 , \1705 );
nand \U$1558 ( \1707 , \1702 , \1706 );
buf \U$1559 ( \1708 , \1707 );
buf \U$1560 ( \1709 , \1708 );
nand \U$1561 ( \1710 , \1696 , \1709 );
buf \U$1562 ( \1711 , \1710 );
xor \U$1563 ( \1712 , \1691 , \1711 );
buf \U$1564 ( \1713 , \978 );
not \U$1565 ( \1714 , \1713 );
buf \U$1566 ( \1715 , \330 );
not \U$1567 ( \1716 , \1715 );
or \U$1568 ( \1717 , \1714 , \1716 );
buf \U$1569 ( \1718 , \344 );
buf \U$1570 ( \1719 , RIc0da288_95);
nand \U$1571 ( \1720 , \1718 , \1719 );
buf \U$1572 ( \1721 , \1720 );
buf \U$1573 ( \1722 , \1721 );
nand \U$1574 ( \1723 , \1717 , \1722 );
buf \U$1575 ( \1724 , \1723 );
xor \U$1576 ( \1725 , \1712 , \1724 );
buf \U$1577 ( \1726 , \1725 );
xor \U$1578 ( \1727 , \1669 , \1726 );
buf \U$1579 ( \1728 , \1727 );
buf \U$1580 ( \1729 , \1728 );
xor \U$1581 ( \1730 , \1647 , \1729 );
buf \U$1582 ( \1731 , \1730 );
buf \U$1583 ( \1732 , \1731 );
xor \U$1584 ( \1733 , \1525 , \1732 );
buf \U$1585 ( \1734 , \1733 );
buf \U$1586 ( \1735 , \1734 );
buf \U$1589 ( \1736 , \572 );
buf \U$1590 ( \1737 , \1736 );
not \U$1591 ( \1738 , \1737 );
buf \U$1592 ( \1739 , \1738 );
buf \U$1593 ( \1740 , \1739 );
buf \U$1594 ( \1741 , RIc0d9ce8_83);
buf \U$1595 ( \1742 , RIc0d7d80_16);
not \U$1596 ( \1743 , \1742 );
buf \U$1597 ( \1744 , \1743 );
buf \U$1598 ( \1745 , \1744 );
and \U$1599 ( \1746 , \1741 , \1745 );
not \U$1600 ( \1747 , \1741 );
buf \U$1601 ( \1748 , RIc0d7d80_16);
and \U$1602 ( \1749 , \1747 , \1748 );
nor \U$1603 ( \1750 , \1746 , \1749 );
buf \U$1604 ( \1751 , \1750 );
buf \U$1605 ( \1752 , \1751 );
or \U$1606 ( \1753 , \1740 , \1752 );
buf \U$1607 ( \1754 , \584 );
not \U$1608 ( \1755 , \1754 );
buf \U$1609 ( \1756 , \1755 );
buf \U$1610 ( \1757 , \1756 );
buf \U$1611 ( \1758 , \549 );
or \U$1612 ( \1759 , \1757 , \1758 );
nand \U$1613 ( \1760 , \1753 , \1759 );
buf \U$1614 ( \1761 , \1760 );
buf \U$1615 ( \1762 , \1761 );
buf \U$1616 ( \1763 , \615 );
not \U$1617 ( \1764 , \1763 );
buf \U$1618 ( \1765 , \1764 );
buf \U$1619 ( \1766 , \1765 );
not \U$1620 ( \1767 , \1766 );
buf \U$1621 ( \1768 , RIc0d7c18_13);
buf \U$1622 ( \1769 , RIc0d9ec8_87);
xnor \U$1623 ( \1770 , \1768 , \1769 );
buf \U$1624 ( \1771 , \1770 );
buf \U$1625 ( \1772 , \1771 );
nor \U$1626 ( \1773 , \1767 , \1772 );
buf \U$1627 ( \1774 , \1773 );
buf \U$1628 ( \1775 , \1774 );
buf \U$1629 ( \1776 , \816 );
buf \U$1630 ( \1777 , RIc0d7ba0_12);
buf \U$1631 ( \1778 , RIc0d9ec8_87);
xor \U$1632 ( \1779 , \1777 , \1778 );
buf \U$1633 ( \1780 , \1779 );
buf \U$1634 ( \1781 , \1780 );
and \U$1635 ( \1782 , \1776 , \1781 );
buf \U$1636 ( \1783 , \1782 );
buf \U$1637 ( \1784 , \1783 );
nor \U$1638 ( \1785 , \1775 , \1784 );
buf \U$1639 ( \1786 , \1785 );
buf \U$1640 ( \1787 , \1786 );
not \U$1641 ( \1788 , \1787 );
buf \U$1642 ( \1789 , \1788 );
buf \U$1643 ( \1790 , \1789 );
xor \U$1644 ( \1791 , \1762 , \1790 );
buf \U$1645 ( \1792 , RIc0d9478_65);
buf \U$1646 ( \1793 , RIc0d8668_35);
xor \U$1647 ( \1794 , \1792 , \1793 );
buf \U$1648 ( \1795 , \1794 );
buf \U$1649 ( \1796 , \1795 );
not \U$1650 ( \1797 , \1796 );
buf \U$1651 ( \1798 , \1224 );
not \U$1652 ( \1799 , \1798 );
or \U$1653 ( \1800 , \1797 , \1799 );
buf \U$1654 ( \1801 , RIc0d9478_65);
buf \U$1655 ( \1802 , RIc0d85f0_34);
xnor \U$1656 ( \1803 , \1801 , \1802 );
buf \U$1657 ( \1804 , \1803 );
buf \U$1658 ( \1805 , \1804 );
not \U$1659 ( \1806 , \1805 );
buf \U$1660 ( \1807 , \1229 );
nand \U$1661 ( \1808 , \1806 , \1807 );
buf \U$1662 ( \1809 , \1808 );
buf \U$1663 ( \1810 , \1809 );
nand \U$1664 ( \1811 , \1800 , \1810 );
buf \U$1665 ( \1812 , \1811 );
buf \U$1666 ( \1813 , \1812 );
buf \U$1667 ( \1814 , RIc0d8578_33);
buf \U$1668 ( \1815 , RIc0d9568_67);
xor \U$1669 ( \1816 , \1814 , \1815 );
buf \U$1670 ( \1817 , \1816 );
buf \U$1671 ( \1818 , \1817 );
not \U$1672 ( \1819 , \1818 );
buf \U$1673 ( \1820 , \674 );
not \U$1674 ( \1821 , \1820 );
buf \U$1675 ( \1822 , \1821 );
buf \U$1678 ( \1823 , \1822 );
buf \U$1679 ( \1824 , \1823 );
not \U$1680 ( \1825 , \1824 );
or \U$1681 ( \1826 , \1819 , \1825 );
buf \U$1682 ( \1827 , RIc0d9568_67);
buf \U$1683 ( \1828 , RIc0d8500_32);
xnor \U$1684 ( \1829 , \1827 , \1828 );
buf \U$1685 ( \1830 , \1829 );
buf \U$1686 ( \1831 , \1830 );
not \U$1687 ( \1832 , \1831 );
buf \U$1688 ( \1833 , \686 );
nand \U$1689 ( \1834 , \1832 , \1833 );
buf \U$1690 ( \1835 , \1834 );
buf \U$1691 ( \1836 , \1835 );
nand \U$1692 ( \1837 , \1826 , \1836 );
buf \U$1693 ( \1838 , \1837 );
buf \U$1694 ( \1839 , \1838 );
xor \U$1695 ( \1840 , \1813 , \1839 );
buf \U$1696 ( \1841 , RIc0d82a8_27);
buf \U$1697 ( \1842 , RIc0d9838_73);
xor \U$1698 ( \1843 , \1841 , \1842 );
buf \U$1699 ( \1844 , \1843 );
buf \U$1700 ( \1845 , \1844 );
not \U$1701 ( \1846 , \1845 );
buf \U$1702 ( \1847 , \776 );
not \U$1703 ( \1848 , \1847 );
or \U$1704 ( \1849 , \1846 , \1848 );
buf \U$1705 ( \1850 , RIc0d8230_26);
buf \U$1706 ( \1851 , RIc0d9838_73);
xnor \U$1707 ( \1852 , \1850 , \1851 );
buf \U$1708 ( \1853 , \1852 );
buf \U$1709 ( \1854 , \1853 );
not \U$1710 ( \1855 , \1854 );
buf \U$1713 ( \1856 , \790 );
buf \U$1714 ( \1857 , \1856 );
nand \U$1715 ( \1858 , \1855 , \1857 );
buf \U$1716 ( \1859 , \1858 );
buf \U$1717 ( \1860 , \1859 );
nand \U$1718 ( \1861 , \1849 , \1860 );
buf \U$1719 ( \1862 , \1861 );
buf \U$1720 ( \1863 , \1862 );
and \U$1721 ( \1864 , \1840 , \1863 );
and \U$1722 ( \1865 , \1813 , \1839 );
or \U$1723 ( \1866 , \1864 , \1865 );
buf \U$1724 ( \1867 , \1866 );
buf \U$1725 ( \1868 , \1867 );
and \U$1726 ( \1869 , \1791 , \1868 );
and \U$1727 ( \1870 , \1762 , \1790 );
or \U$1728 ( \1871 , \1869 , \1870 );
buf \U$1729 ( \1872 , \1871 );
buf \U$1730 ( \1873 , \1872 );
not \U$1731 ( \1874 , \1282 );
buf \U$1732 ( \1875 , RIc0d8320_28);
buf \U$1733 ( \1876 , RIc0d9748_71);
xor \U$1734 ( \1877 , \1875 , \1876 );
buf \U$1735 ( \1878 , \1877 );
not \U$1736 ( \1879 , \1878 );
or \U$1737 ( \1880 , \1874 , \1879 );
buf \U$1738 ( \1881 , RIc0d9748_71);
buf \U$1739 ( \1882 , RIc0d8398_29);
xnor \U$1740 ( \1883 , \1881 , \1882 );
buf \U$1741 ( \1884 , \1883 );
not \U$1742 ( \1885 , \1884 );
buf \U$1743 ( \1886 , \1260 );
not \U$1744 ( \1887 , \1886 );
buf \U$1745 ( \1888 , \1887 );
nand \U$1746 ( \1889 , \1885 , \1888 );
nand \U$1747 ( \1890 , \1880 , \1889 );
buf \U$1748 ( \1891 , \1890 );
not \U$1749 ( \1892 , \1891 );
buf \U$1750 ( \1893 , RIc0d7948_7);
buf \U$1751 ( \1894 , RIc0da198_93);
xor \U$1752 ( \1895 , \1893 , \1894 );
buf \U$1753 ( \1896 , \1895 );
buf \U$1754 ( \1897 , \1896 );
not \U$1755 ( \1898 , \1897 );
buf \U$1756 ( \1899 , \473 );
not \U$1757 ( \1900 , \1899 );
buf \U$1758 ( \1901 , \1900 );
buf \U$1759 ( \1902 , \1901 );
not \U$1760 ( \1903 , \1902 );
or \U$1761 ( \1904 , \1898 , \1903 );
buf \U$1762 ( \1905 , \481 );
xor \U$1763 ( \1906 , RIc0da198_93, RIc0d78d0_6);
buf \U$1764 ( \1907 , \1906 );
nand \U$1765 ( \1908 , \1905 , \1907 );
buf \U$1766 ( \1909 , \1908 );
buf \U$1767 ( \1910 , \1909 );
nand \U$1768 ( \1911 , \1904 , \1910 );
buf \U$1769 ( \1912 , \1911 );
buf \U$1770 ( \1913 , \1912 );
not \U$1771 ( \1914 , \1913 );
or \U$1772 ( \1915 , \1892 , \1914 );
buf \U$1773 ( \1916 , \1890 );
buf \U$1774 ( \1917 , \1912 );
or \U$1775 ( \1918 , \1916 , \1917 );
buf \U$1776 ( \1919 , RIc0d7a38_9);
buf \U$1777 ( \1920 , RIc0da0a8_91);
xor \U$1778 ( \1921 , \1919 , \1920 );
buf \U$1779 ( \1922 , \1921 );
buf \U$1780 ( \1923 , \1922 );
not \U$1781 ( \1924 , \1923 );
buf \U$1782 ( \1925 , \521 );
not \U$1783 ( \1926 , \1925 );
buf \U$1784 ( \1927 , \1926 );
buf \U$1785 ( \1928 , \1927 );
not \U$1786 ( \1929 , \1928 );
or \U$1787 ( \1930 , \1924 , \1929 );
buf \U$1788 ( \1931 , \710 );
not \U$1789 ( \1932 , \1931 );
buf \U$1790 ( \1933 , \1932 );
buf \U$1791 ( \1934 , \1933 );
buf \U$1792 ( \1935 , RIc0d79c0_8);
buf \U$1793 ( \1936 , RIc0da0a8_91);
xor \U$1794 ( \1937 , \1935 , \1936 );
buf \U$1795 ( \1938 , \1937 );
buf \U$1796 ( \1939 , \1938 );
nand \U$1797 ( \1940 , \1934 , \1939 );
buf \U$1798 ( \1941 , \1940 );
buf \U$1799 ( \1942 , \1941 );
nand \U$1800 ( \1943 , \1930 , \1942 );
buf \U$1801 ( \1944 , \1943 );
buf \U$1802 ( \1945 , \1944 );
nand \U$1803 ( \1946 , \1918 , \1945 );
buf \U$1804 ( \1947 , \1946 );
buf \U$1805 ( \1948 , \1947 );
nand \U$1806 ( \1949 , \1915 , \1948 );
buf \U$1807 ( \1950 , \1949 );
buf \U$1808 ( \1951 , \1950 );
not \U$1809 ( \1952 , \1600 );
buf \U$1810 ( \1953 , RIc0d7ee8_19);
buf \U$1811 ( \1954 , RIc0d9bf8_81);
xnor \U$1812 ( \1955 , \1953 , \1954 );
buf \U$1813 ( \1956 , \1955 );
not \U$1814 ( \1957 , \1956 );
and \U$1815 ( \1958 , \1952 , \1957 );
buf \U$1816 ( \1959 , RIc0d7e70_18);
buf \U$1817 ( \1960 , RIc0d9bf8_81);
xor \U$1818 ( \1961 , \1959 , \1960 );
buf \U$1819 ( \1962 , \1961 );
and \U$1820 ( \1963 , \1078 , \1962 );
nor \U$1821 ( \1964 , \1958 , \1963 );
buf \U$1822 ( \1965 , \1964 );
not \U$1823 ( \1966 , \1965 );
buf \U$1824 ( \1967 , \874 );
not \U$1825 ( \1968 , \1967 );
buf \U$1826 ( \1969 , \1968 );
not \U$1827 ( \1970 , \1969 );
xnor \U$1828 ( \1971 , RIc0d9658_69, RIc0d8410_30);
not \U$1829 ( \1972 , \1971 );
and \U$1830 ( \1973 , \1970 , \1972 );
not \U$1831 ( \1974 , \864 );
buf \U$1832 ( \1975 , RIc0d9658_69);
buf \U$1833 ( \1976 , RIc0d8488_31);
xnor \U$1834 ( \1977 , \1975 , \1976 );
buf \U$1835 ( \1978 , \1977 );
nor \U$1836 ( \1979 , \1974 , \1978 );
nor \U$1837 ( \1980 , \1973 , \1979 );
buf \U$1838 ( \1981 , \1980 );
not \U$1839 ( \1982 , \1981 );
or \U$1840 ( \1983 , \1966 , \1982 );
buf \U$1841 ( \1984 , RIc0da288_95);
buf \U$1842 ( \1985 , RIc0d7858_5);
and \U$1843 ( \1986 , \1984 , \1985 );
not \U$1844 ( \1987 , \1984 );
buf \U$1845 ( \1988 , RIc0d7858_5);
not \U$1846 ( \1989 , \1988 );
buf \U$1847 ( \1990 , \1989 );
buf \U$1848 ( \1991 , \1990 );
and \U$1849 ( \1992 , \1987 , \1991 );
nor \U$1850 ( \1993 , \1986 , \1992 );
buf \U$1851 ( \1994 , \1993 );
buf \U$1852 ( \1995 , \1994 );
not \U$1853 ( \1996 , \1995 );
buf \U$1854 ( \1997 , \336 );
not \U$1855 ( \1998 , \1997 );
or \U$1856 ( \1999 , \1996 , \1998 );
buf \U$1857 ( \2000 , \344 );
buf \U$1858 ( \2001 , RIc0da288_95);
buf \U$1859 ( \2002 , RIc0d77e0_4);
and \U$1860 ( \2003 , \2001 , \2002 );
not \U$1861 ( \2004 , \2001 );
buf \U$1862 ( \2005 , \489 );
and \U$1863 ( \2006 , \2004 , \2005 );
nor \U$1864 ( \2007 , \2003 , \2006 );
buf \U$1865 ( \2008 , \2007 );
buf \U$1866 ( \2009 , \2008 );
nand \U$1867 ( \2010 , \2000 , \2009 );
buf \U$1868 ( \2011 , \2010 );
buf \U$1869 ( \2012 , \2011 );
nand \U$1870 ( \2013 , \1999 , \2012 );
buf \U$1871 ( \2014 , \2013 );
buf \U$1872 ( \2015 , \2014 );
nand \U$1873 ( \2016 , \1983 , \2015 );
buf \U$1874 ( \2017 , \2016 );
buf \U$1875 ( \2018 , \2017 );
buf \U$1876 ( \2019 , \1980 );
buf \U$1877 ( \2020 , \1964 );
or \U$1878 ( \2021 , \2019 , \2020 );
buf \U$1879 ( \2022 , \2021 );
buf \U$1880 ( \2023 , \2022 );
nand \U$1881 ( \2024 , \2018 , \2023 );
buf \U$1882 ( \2025 , \2024 );
buf \U$1883 ( \2026 , \2025 );
xor \U$1884 ( \2027 , \1951 , \2026 );
buf \U$1885 ( \2028 , RIc0d7b28_11);
buf \U$1886 ( \2029 , RIc0d9fb8_89);
xor \U$1887 ( \2030 , \2028 , \2029 );
buf \U$1888 ( \2031 , \2030 );
buf \U$1889 ( \2032 , \2031 );
not \U$1890 ( \2033 , \2032 );
buf \U$1893 ( \2034 , \432 );
buf \U$1894 ( \2035 , \2034 );
not \U$1895 ( \2036 , \2035 );
buf \U$1896 ( \2037 , \2036 );
buf \U$1899 ( \2038 , \2037 );
buf \U$1900 ( \2039 , \2038 );
not \U$1901 ( \2040 , \2039 );
or \U$1902 ( \2041 , \2033 , \2040 );
buf \U$1903 ( \2042 , \846 );
buf \U$1904 ( \2043 , RIc0d7ab0_10);
buf \U$1905 ( \2044 , RIc0d9fb8_89);
xor \U$1906 ( \2045 , \2043 , \2044 );
buf \U$1907 ( \2046 , \2045 );
buf \U$1908 ( \2047 , \2046 );
nand \U$1909 ( \2048 , \2042 , \2047 );
buf \U$1910 ( \2049 , \2048 );
buf \U$1911 ( \2050 , \2049 );
nand \U$1912 ( \2051 , \2041 , \2050 );
buf \U$1913 ( \2052 , \2051 );
buf \U$1914 ( \2053 , \2052 );
buf \U$1915 ( \2054 , RIc0da378_97);
buf \U$1916 ( \2055 , RIc0d7768_3);
and \U$1917 ( \2056 , \2054 , \2055 );
not \U$1918 ( \2057 , \2054 );
buf \U$1919 ( \2058 , \304 );
and \U$1920 ( \2059 , \2057 , \2058 );
nor \U$1921 ( \2060 , \2056 , \2059 );
buf \U$1922 ( \2061 , \2060 );
buf \U$1923 ( \2062 , \2061 );
not \U$1924 ( \2063 , \2062 );
buf \U$1925 ( \2064 , \749 );
not \U$1926 ( \2065 , \2064 );
buf \U$1927 ( \2066 , \2065 );
buf \U$1928 ( \2067 , \2066 );
not \U$1929 ( \2068 , \2067 );
or \U$1930 ( \2069 , \2063 , \2068 );
buf \U$1933 ( \2070 , \733 );
buf \U$1934 ( \2071 , \2070 );
buf \U$1935 ( \2072 , RIc0da378_97);
buf \U$1936 ( \2073 , RIc0d76f0_2);
and \U$1937 ( \2074 , \2072 , \2073 );
not \U$1938 ( \2075 , \2072 );
buf \U$1939 ( \2076 , \352 );
and \U$1940 ( \2077 , \2075 , \2076 );
nor \U$1941 ( \2078 , \2074 , \2077 );
buf \U$1942 ( \2079 , \2078 );
buf \U$1943 ( \2080 , \2079 );
nand \U$1944 ( \2081 , \2071 , \2080 );
buf \U$1945 ( \2082 , \2081 );
buf \U$1946 ( \2083 , \2082 );
nand \U$1947 ( \2084 , \2069 , \2083 );
buf \U$1948 ( \2085 , \2084 );
buf \U$1949 ( \2086 , \2085 );
xor \U$1950 ( \2087 , \2053 , \2086 );
buf \U$1953 ( \2088 , \572 );
buf \U$1954 ( \2089 , \2088 );
not \U$1955 ( \2090 , \2089 );
buf \U$1956 ( \2091 , \2090 );
buf \U$1957 ( \2092 , \2091 );
buf \U$1958 ( \2093 , RIc0d7df8_17);
buf \U$1959 ( \2094 , RIc0d9ce8_83);
xnor \U$1960 ( \2095 , \2093 , \2094 );
buf \U$1961 ( \2096 , \2095 );
buf \U$1962 ( \2097 , \2096 );
or \U$1963 ( \2098 , \2092 , \2097 );
buf \U$1964 ( \2099 , \996 );
buf \U$1965 ( \2100 , \1751 );
or \U$1966 ( \2101 , \2099 , \2100 );
nand \U$1967 ( \2102 , \2098 , \2101 );
buf \U$1968 ( \2103 , \2102 );
buf \U$1969 ( \2104 , \2103 );
and \U$1970 ( \2105 , \2087 , \2104 );
and \U$1971 ( \2106 , \2053 , \2086 );
or \U$1972 ( \2107 , \2105 , \2106 );
buf \U$1973 ( \2108 , \2107 );
buf \U$1974 ( \2109 , \2108 );
and \U$1975 ( \2110 , \2027 , \2109 );
and \U$1976 ( \2111 , \1951 , \2026 );
or \U$1977 ( \2112 , \2110 , \2111 );
buf \U$1978 ( \2113 , \2112 );
buf \U$1979 ( \2114 , \2113 );
xor \U$1980 ( \2115 , \1873 , \2114 );
buf \U$1981 ( \2116 , RIc0d8140_24);
buf \U$1982 ( \2117 , RIc0d9928_75);
xor \U$1983 ( \2118 , \2116 , \2117 );
buf \U$1984 ( \2119 , \2118 );
buf \U$1985 ( \2120 , \2119 );
not \U$1986 ( \2121 , \2120 );
buf \U$1987 ( \2122 , \1124 );
not \U$1988 ( \2123 , \2122 );
buf \U$1989 ( \2124 , \2123 );
buf \U$1990 ( \2125 , \2124 );
not \U$1991 ( \2126 , \2125 );
or \U$1992 ( \2127 , \2121 , \2126 );
buf \U$1993 ( \2128 , \1565 );
buf \U$1994 ( \2129 , \1551 );
nand \U$1995 ( \2130 , \2128 , \2129 );
buf \U$1996 ( \2131 , \2130 );
buf \U$1997 ( \2132 , \2131 );
nand \U$1998 ( \2133 , \2127 , \2132 );
buf \U$1999 ( \2134 , \2133 );
buf \U$2000 ( \2135 , \2134 );
not \U$2001 ( \2136 , \2135 );
buf \U$2002 ( \2137 , RIc0d8050_22);
buf \U$2003 ( \2138 , RIc0d9a18_77);
xor \U$2004 ( \2139 , \2137 , \2138 );
buf \U$2005 ( \2140 , \2139 );
buf \U$2006 ( \2141 , \2140 );
not \U$2007 ( \2142 , \2141 );
buf \U$2008 ( \2143 , \1431 );
not \U$2009 ( \2144 , \2143 );
or \U$2010 ( \2145 , \2142 , \2144 );
buf \U$2011 ( \2146 , \1588 );
buf \U$2012 ( \2147 , \1577 );
nand \U$2013 ( \2148 , \2146 , \2147 );
buf \U$2014 ( \2149 , \2148 );
buf \U$2015 ( \2150 , \2149 );
nand \U$2016 ( \2151 , \2145 , \2150 );
buf \U$2017 ( \2152 , \2151 );
buf \U$2018 ( \2153 , \2152 );
not \U$2019 ( \2154 , \2153 );
or \U$2020 ( \2155 , \2136 , \2154 );
buf \U$2021 ( \2156 , \2152 );
buf \U$2022 ( \2157 , \2134 );
or \U$2023 ( \2158 , \2156 , \2157 );
buf \U$2024 ( \2159 , \1962 );
not \U$2025 ( \2160 , \2159 );
buf \U$2026 ( \2161 , \1064 );
not \U$2027 ( \2162 , \2161 );
or \U$2028 ( \2163 , \2160 , \2162 );
buf \U$2029 ( \2164 , \1605 );
not \U$2030 ( \2165 , \2164 );
buf \U$2031 ( \2166 , \1078 );
nand \U$2032 ( \2167 , \2165 , \2166 );
buf \U$2033 ( \2168 , \2167 );
buf \U$2034 ( \2169 , \2168 );
nand \U$2035 ( \2170 , \2163 , \2169 );
buf \U$2036 ( \2171 , \2170 );
buf \U$2037 ( \2172 , \2171 );
nand \U$2038 ( \2173 , \2158 , \2172 );
buf \U$2039 ( \2174 , \2173 );
buf \U$2040 ( \2175 , \2174 );
nand \U$2041 ( \2176 , \2155 , \2175 );
buf \U$2042 ( \2177 , \2176 );
buf \U$2043 ( \2178 , \2177 );
buf \U$2044 ( \2179 , \1906 );
not \U$2045 ( \2180 , \2179 );
buf \U$2046 ( \2181 , \476 );
not \U$2047 ( \2182 , \2181 );
or \U$2048 ( \2183 , \2180 , \2182 );
buf \U$2049 ( \2184 , \481 );
buf \U$2050 ( \2185 , \458 );
nand \U$2051 ( \2186 , \2184 , \2185 );
buf \U$2052 ( \2187 , \2186 );
buf \U$2053 ( \2188 , \2187 );
nand \U$2054 ( \2189 , \2183 , \2188 );
buf \U$2055 ( \2190 , \2189 );
buf \U$2056 ( \2191 , \2190 );
buf \U$2057 ( \2192 , RIc0da4e0_100);
buf \U$2058 ( \2193 , RIc0da558_101);
xor \U$2059 ( \2194 , \2192 , \2193 );
buf \U$2060 ( \2195 , \2194 );
buf \U$2061 ( \2196 , \2195 );
not \U$2062 ( \2197 , \2196 );
buf \U$2063 ( \2198 , \2197 );
buf \U$2066 ( \2199 , \2198 );
buf \U$2067 ( \2200 , \2199 );
not \U$2068 ( \2201 , \2200 );
buf \U$2069 ( \2202 , \2198 );
xor \U$2070 ( \2203 , RIc0da4e0_100, RIc0da468_99);
buf \U$2071 ( \2204 , \2203 );
nand \U$2072 ( \2205 , \2202 , \2204 );
buf \U$2073 ( \2206 , \2205 );
buf \U$2076 ( \2207 , \2206 );
buf \U$2077 ( \2208 , \2207 );
not \U$2078 ( \2209 , \2208 );
or \U$2079 ( \2210 , \2201 , \2209 );
buf \U$2080 ( \2211 , RIc0da468_99);
nand \U$2081 ( \2212 , \2210 , \2211 );
buf \U$2082 ( \2213 , \2212 );
buf \U$2083 ( \2214 , \2213 );
nor \U$2084 ( \2215 , \2191 , \2214 );
buf \U$2085 ( \2216 , \2215 );
buf \U$2086 ( \2217 , \2216 );
buf \U$2087 ( \2218 , RIc0d7f60_20);
buf \U$2088 ( \2219 , RIc0d9b08_79);
xnor \U$2089 ( \2220 , \2218 , \2219 );
buf \U$2090 ( \2221 , \2220 );
buf \U$2091 ( \2222 , \2221 );
not \U$2092 ( \2223 , \2222 );
buf \U$2093 ( \2224 , \2223 );
buf \U$2094 ( \2225 , \2224 );
not \U$2095 ( \2226 , \2225 );
buf \U$2096 ( \2227 , \1351 );
not \U$2097 ( \2228 , \2227 );
or \U$2098 ( \2229 , \2226 , \2228 );
buf \U$2099 ( \2230 , \1026 );
buf \U$2100 ( \2231 , \370 );
nand \U$2101 ( \2232 , \2230 , \2231 );
buf \U$2102 ( \2233 , \2232 );
buf \U$2103 ( \2234 , \2233 );
nand \U$2104 ( \2235 , \2229 , \2234 );
buf \U$2105 ( \2236 , \2235 );
buf \U$2106 ( \2237 , \2236 );
not \U$2107 ( \2238 , \2237 );
buf \U$2108 ( \2239 , \2238 );
buf \U$2109 ( \2240 , \2239 );
or \U$2110 ( \2241 , \2217 , \2240 );
buf \U$2111 ( \2242 , \2190 );
buf \U$2112 ( \2243 , \2213 );
nand \U$2113 ( \2244 , \2242 , \2243 );
buf \U$2114 ( \2245 , \2244 );
buf \U$2115 ( \2246 , \2245 );
nand \U$2116 ( \2247 , \2241 , \2246 );
buf \U$2117 ( \2248 , \2247 );
buf \U$2118 ( \2249 , \2248 );
xor \U$2119 ( \2250 , \2178 , \2249 );
buf \U$2120 ( \2251 , \1221 );
buf \U$2121 ( \2252 , \1804 );
or \U$2122 ( \2253 , \2251 , \2252 );
buf \U$2123 ( \2254 , \1232 );
xor \U$2124 ( \2255 , \655 , \656 );
buf \U$2125 ( \2256 , \2255 );
buf \U$2126 ( \2257 , \2256 );
not \U$2127 ( \2258 , \2257 );
buf \U$2128 ( \2259 , \2258 );
buf \U$2129 ( \2260 , \2259 );
or \U$2130 ( \2261 , \2254 , \2260 );
nand \U$2131 ( \2262 , \2253 , \2261 );
buf \U$2132 ( \2263 , \2262 );
buf \U$2133 ( \2264 , \2263 );
buf \U$2134 ( \2265 , \1878 );
not \U$2135 ( \2266 , \2265 );
buf \U$2136 ( \2267 , \1260 );
not \U$2137 ( \2268 , \2267 );
buf \U$2138 ( \2269 , \2268 );
buf \U$2139 ( \2270 , \2269 );
not \U$2140 ( \2271 , \2270 );
or \U$2141 ( \2272 , \2266 , \2271 );
buf \U$2142 ( \2273 , \1282 );
buf \U$2143 ( \2274 , RIc0d82a8_27);
buf \U$2144 ( \2275 , RIc0d9748_71);
xor \U$2145 ( \2276 , \2274 , \2275 );
buf \U$2146 ( \2277 , \2276 );
buf \U$2147 ( \2278 , \2277 );
nand \U$2148 ( \2279 , \2273 , \2278 );
buf \U$2149 ( \2280 , \2279 );
buf \U$2150 ( \2281 , \2280 );
nand \U$2151 ( \2282 , \2272 , \2281 );
buf \U$2152 ( \2283 , \2282 );
buf \U$2153 ( \2284 , \2283 );
xor \U$2154 ( \2285 , \2264 , \2284 );
buf \U$2155 ( \2286 , \2008 );
not \U$2156 ( \2287 , \2286 );
buf \U$2157 ( \2288 , \336 );
not \U$2158 ( \2289 , \2288 );
or \U$2159 ( \2290 , \2287 , \2289 );
buf \U$2160 ( \2291 , \344 );
buf \U$2161 ( \2292 , \308 );
nand \U$2162 ( \2293 , \2291 , \2292 );
buf \U$2163 ( \2294 , \2293 );
buf \U$2164 ( \2295 , \2294 );
nand \U$2165 ( \2296 , \2290 , \2295 );
buf \U$2166 ( \2297 , \2296 );
buf \U$2167 ( \2298 , \2297 );
and \U$2168 ( \2299 , \2285 , \2298 );
and \U$2169 ( \2300 , \2264 , \2284 );
or \U$2170 ( \2301 , \2299 , \2300 );
buf \U$2171 ( \2302 , \2301 );
buf \U$2172 ( \2303 , \2302 );
xor \U$2173 ( \2304 , \2250 , \2303 );
buf \U$2174 ( \2305 , \2304 );
buf \U$2175 ( \2306 , \2305 );
and \U$2176 ( \2307 , \2115 , \2306 );
and \U$2177 ( \2308 , \1873 , \2114 );
or \U$2178 ( \2309 , \2307 , \2308 );
buf \U$2179 ( \2310 , \2309 );
buf \U$2180 ( \2311 , \2310 );
buf \U$2181 ( \2312 , \954 );
not \U$2182 ( \2313 , \2312 );
xnor \U$2183 ( \2314 , RIc0d9dd8_85, RIc0d7d08_15);
buf \U$2184 ( \2315 , \2314 );
not \U$2185 ( \2316 , \2315 );
and \U$2186 ( \2317 , \2313 , \2316 );
buf \U$2187 ( \2318 , \1401 );
buf \U$2188 ( \2319 , RIc0d7c90_14);
buf \U$2189 ( \2320 , RIc0d9dd8_85);
xor \U$2190 ( \2321 , \2319 , \2320 );
buf \U$2191 ( \2322 , \2321 );
buf \U$2192 ( \2323 , \2322 );
and \U$2193 ( \2324 , \2318 , \2323 );
buf \U$2194 ( \2325 , \2324 );
buf \U$2195 ( \2326 , \2325 );
nor \U$2196 ( \2327 , \2317 , \2326 );
buf \U$2197 ( \2328 , \2327 );
buf \U$2198 ( \2329 , \2328 );
not \U$2199 ( \2330 , \2329 );
buf \U$2200 ( \2331 , \2330 );
buf \U$2201 ( \2332 , \2331 );
not \U$2202 ( \2333 , \2332 );
buf \U$2203 ( \2334 , RIc0d80c8_23);
buf \U$2204 ( \2335 , RIc0d9a18_77);
xor \U$2205 ( \2336 , \2334 , \2335 );
buf \U$2206 ( \2337 , \2336 );
buf \U$2207 ( \2338 , \2337 );
not \U$2208 ( \2339 , \2338 );
buf \U$2209 ( \2340 , \1183 );
not \U$2210 ( \2341 , \2340 );
or \U$2211 ( \2342 , \2339 , \2341 );
buf \U$2212 ( \2343 , \1196 );
buf \U$2213 ( \2344 , \2140 );
nand \U$2214 ( \2345 , \2343 , \2344 );
buf \U$2215 ( \2346 , \2345 );
buf \U$2216 ( \2347 , \2346 );
nand \U$2217 ( \2348 , \2342 , \2347 );
buf \U$2218 ( \2349 , \2348 );
buf \U$2219 ( \2350 , \2349 );
not \U$2220 ( \2351 , \2350 );
or \U$2221 ( \2352 , \2333 , \2351 );
buf \U$2222 ( \2353 , \2331 );
buf \U$2223 ( \2354 , \2349 );
or \U$2224 ( \2355 , \2353 , \2354 );
buf \U$2225 ( \2356 , \1123 );
not \U$2226 ( \2357 , \2356 );
buf \U$2227 ( \2358 , \2357 );
buf \U$2230 ( \2359 , \2358 );
buf \U$2231 ( \2360 , \2359 );
not \U$2232 ( \2361 , \2360 );
buf \U$2233 ( \2362 , \2361 );
buf \U$2234 ( \2363 , \2362 );
buf \U$2235 ( \2364 , RIc0d81b8_25);
buf \U$2236 ( \2365 , RIc0d9928_75);
xnor \U$2237 ( \2366 , \2364 , \2365 );
buf \U$2238 ( \2367 , \2366 );
buf \U$2239 ( \2368 , \2367 );
or \U$2240 ( \2369 , \2363 , \2368 );
buf \U$2241 ( \2370 , \1143 );
not \U$2242 ( \2371 , \2370 );
buf \U$2243 ( \2372 , \2371 );
buf \U$2244 ( \2373 , \2372 );
buf \U$2245 ( \2374 , \2119 );
not \U$2246 ( \2375 , \2374 );
buf \U$2247 ( \2376 , \2375 );
buf \U$2248 ( \2377 , \2376 );
or \U$2249 ( \2378 , \2373 , \2377 );
nand \U$2250 ( \2379 , \2369 , \2378 );
buf \U$2251 ( \2380 , \2379 );
buf \U$2252 ( \2381 , \2380 );
nand \U$2253 ( \2382 , \2355 , \2381 );
buf \U$2254 ( \2383 , \2382 );
buf \U$2255 ( \2384 , \2383 );
nand \U$2256 ( \2385 , \2352 , \2384 );
buf \U$2257 ( \2386 , \2385 );
buf \U$2258 ( \2387 , \2386 );
not \U$2259 ( \2388 , \2387 );
buf \U$2260 ( \2389 , \2322 );
not \U$2261 ( \2390 , \2389 );
buf \U$2262 ( \2391 , \946 );
not \U$2263 ( \2392 , \2391 );
buf \U$2264 ( \2393 , \2392 );
buf \U$2265 ( \2394 , \2393 );
not \U$2266 ( \2395 , \2394 );
buf \U$2267 ( \2396 , \2395 );
buf \U$2268 ( \2397 , \2396 );
not \U$2269 ( \2398 , \2397 );
buf \U$2270 ( \2399 , \2398 );
buf \U$2271 ( \2400 , \2399 );
not \U$2272 ( \2401 , \2400 );
or \U$2273 ( \2402 , \2390 , \2401 );
buf \U$2274 ( \2403 , RIc0d9dd8_85);
buf \U$2275 ( \2404 , RIc0d7c18_13);
xnor \U$2276 ( \2405 , \2403 , \2404 );
buf \U$2277 ( \2406 , \2405 );
buf \U$2278 ( \2407 , \2406 );
not \U$2279 ( \2408 , \2407 );
buf \U$2280 ( \2409 , \1401 );
nand \U$2281 ( \2410 , \2408 , \2409 );
buf \U$2282 ( \2411 , \2410 );
buf \U$2283 ( \2412 , \2411 );
nand \U$2284 ( \2413 , \2402 , \2412 );
buf \U$2285 ( \2414 , \2413 );
buf \U$2286 ( \2415 , \2414 );
not \U$2287 ( \2416 , \2415 );
buf \U$2288 ( \2417 , \2416 );
buf \U$2289 ( \2418 , \2079 );
not \U$2290 ( \2419 , \2418 );
buf \U$2291 ( \2420 , \2066 );
not \U$2292 ( \2421 , \2420 );
or \U$2293 ( \2422 , \2419 , \2421 );
buf \U$2294 ( \2423 , \2070 );
buf \U$2295 ( \2424 , RIc0da378_97);
buf \U$2296 ( \2425 , RIc0d7678_1);
and \U$2297 ( \2426 , \2424 , \2425 );
not \U$2298 ( \2427 , \2424 );
buf \U$2299 ( \2428 , \974 );
and \U$2300 ( \2429 , \2427 , \2428 );
nor \U$2301 ( \2430 , \2426 , \2429 );
buf \U$2302 ( \2431 , \2430 );
buf \U$2303 ( \2432 , \2431 );
nand \U$2304 ( \2433 , \2423 , \2432 );
buf \U$2305 ( \2434 , \2433 );
buf \U$2306 ( \2435 , \2434 );
nand \U$2307 ( \2436 , \2422 , \2435 );
buf \U$2308 ( \2437 , \2436 );
xor \U$2309 ( \2438 , \2417 , \2437 );
not \U$2310 ( \2439 , \773 );
not \U$2311 ( \2440 , \1853 );
and \U$2312 ( \2441 , \2439 , \2440 );
buf \U$2313 ( \2442 , RIc0d81b8_25);
buf \U$2314 ( \2443 , RIc0d9838_73);
xor \U$2315 ( \2444 , \2442 , \2443 );
buf \U$2316 ( \2445 , \2444 );
and \U$2317 ( \2446 , \1856 , \2445 );
nor \U$2318 ( \2447 , \2441 , \2446 );
xnor \U$2319 ( \2448 , \2438 , \2447 );
buf \U$2320 ( \2449 , \2448 );
nand \U$2321 ( \2450 , \2388 , \2449 );
buf \U$2322 ( \2451 , \2450 );
buf \U$2323 ( \2452 , \2451 );
buf \U$2324 ( \2453 , RIc0d9478_65);
buf \U$2325 ( \2454 , RIc0d86e0_36);
and \U$2326 ( \2455 , \2453 , \2454 );
buf \U$2327 ( \2456 , \2455 );
buf \U$2328 ( \2457 , \2456 );
buf \U$2329 ( \2458 , RIc0da468_99);
buf \U$2330 ( \2459 , RIc0d7678_1);
and \U$2331 ( \2460 , \2458 , \2459 );
not \U$2332 ( \2461 , \2458 );
buf \U$2333 ( \2462 , \974 );
and \U$2334 ( \2463 , \2461 , \2462 );
nor \U$2335 ( \2464 , \2460 , \2463 );
buf \U$2336 ( \2465 , \2464 );
buf \U$2337 ( \2466 , \2465 );
not \U$2338 ( \2467 , \2466 );
buf \U$2339 ( \2468 , \2207 );
not \U$2340 ( \2469 , \2468 );
buf \U$2341 ( \2470 , \2469 );
buf \U$2342 ( \2471 , \2470 );
not \U$2343 ( \2472 , \2471 );
or \U$2344 ( \2473 , \2467 , \2472 );
buf \U$2345 ( \2474 , \2199 );
not \U$2346 ( \2475 , \2474 );
buf \U$2347 ( \2476 , \2475 );
buf \U$2348 ( \2477 , \2476 );
buf \U$2349 ( \2478 , RIc0da468_99);
nand \U$2350 ( \2479 , \2477 , \2478 );
buf \U$2351 ( \2480 , \2479 );
buf \U$2352 ( \2481 , \2480 );
nand \U$2353 ( \2482 , \2473 , \2481 );
buf \U$2354 ( \2483 , \2482 );
buf \U$2355 ( \2484 , \2483 );
xor \U$2356 ( \2485 , \2457 , \2484 );
buf \U$2357 ( \2486 , \393 );
buf \U$2358 ( \2487 , RIc0d9b08_79);
buf \U$2359 ( \2488 , RIc0d7fd8_21);
xnor \U$2360 ( \2489 , \2487 , \2488 );
buf \U$2361 ( \2490 , \2489 );
buf \U$2362 ( \2491 , \2490 );
or \U$2363 ( \2492 , \2486 , \2491 );
not \U$2364 ( \2493 , \1026 );
buf \U$2365 ( \2494 , \2493 );
buf \U$2366 ( \2495 , \2221 );
or \U$2367 ( \2496 , \2494 , \2495 );
nand \U$2368 ( \2497 , \2492 , \2496 );
buf \U$2369 ( \2498 , \2497 );
buf \U$2370 ( \2499 , \2498 );
and \U$2371 ( \2500 , \2485 , \2499 );
and \U$2372 ( \2501 , \2457 , \2484 );
or \U$2373 ( \2502 , \2500 , \2501 );
buf \U$2374 ( \2503 , \2502 );
buf \U$2375 ( \2504 , \2503 );
and \U$2376 ( \2505 , \2452 , \2504 );
buf \U$2377 ( \2506 , \2386 );
not \U$2378 ( \2507 , \2506 );
buf \U$2379 ( \2508 , \2448 );
nor \U$2380 ( \2509 , \2507 , \2508 );
buf \U$2381 ( \2510 , \2509 );
buf \U$2382 ( \2511 , \2510 );
nor \U$2383 ( \2512 , \2505 , \2511 );
buf \U$2384 ( \2513 , \2512 );
buf \U$2385 ( \2514 , \2513 );
not \U$2386 ( \2515 , \2514 );
buf \U$2387 ( \2516 , \2515 );
buf \U$2388 ( \2517 , \2516 );
not \U$2389 ( \2518 , \2517 );
and \U$2390 ( \2519 , \1792 , \1793 );
buf \U$2391 ( \2520 , \2519 );
buf \U$2392 ( \2521 , \2520 );
not \U$2393 ( \2522 , \686 );
xor \U$2394 ( \2523 , RIc0d9568_67, RIc0d8488_31);
not \U$2395 ( \2524 , \2523 );
or \U$2396 ( \2525 , \2522 , \2524 );
not \U$2397 ( \2526 , \1830 );
nand \U$2398 ( \2527 , \2526 , \678 );
nand \U$2399 ( \2528 , \2525 , \2527 );
buf \U$2400 ( \2529 , \2528 );
xor \U$2401 ( \2530 , \2521 , \2529 );
buf \U$2402 ( \2531 , \1938 );
not \U$2403 ( \2532 , \2531 );
buf \U$2404 ( \2533 , \521 );
not \U$2405 ( \2534 , \2533 );
buf \U$2406 ( \2535 , \2534 );
buf \U$2407 ( \2536 , \2535 );
not \U$2408 ( \2537 , \2536 );
or \U$2409 ( \2538 , \2532 , \2537 );
buf \U$2410 ( \2539 , \1933 );
buf \U$2411 ( \2540 , \506 );
nand \U$2412 ( \2541 , \2539 , \2540 );
buf \U$2413 ( \2542 , \2541 );
buf \U$2414 ( \2543 , \2542 );
nand \U$2415 ( \2544 , \2538 , \2543 );
buf \U$2416 ( \2545 , \2544 );
buf \U$2417 ( \2546 , \2545 );
and \U$2418 ( \2547 , \2530 , \2546 );
and \U$2419 ( \2548 , \2521 , \2529 );
or \U$2420 ( \2549 , \2547 , \2548 );
buf \U$2421 ( \2550 , \2549 );
buf \U$2422 ( \2551 , \2550 );
not \U$2423 ( \2552 , \2551 );
buf \U$2424 ( \2553 , \2447 );
not \U$2425 ( \2554 , \2553 );
buf \U$2426 ( \2555 , \2417 );
not \U$2427 ( \2556 , \2555 );
or \U$2428 ( \2557 , \2554 , \2556 );
buf \U$2429 ( \2558 , \2437 );
nand \U$2430 ( \2559 , \2557 , \2558 );
buf \U$2431 ( \2560 , \2559 );
buf \U$2432 ( \2561 , \2560 );
buf \U$2433 ( \2562 , \2447 );
not \U$2434 ( \2563 , \2562 );
buf \U$2435 ( \2564 , \2414 );
nand \U$2436 ( \2565 , \2563 , \2564 );
buf \U$2437 ( \2566 , \2565 );
buf \U$2438 ( \2567 , \2566 );
nand \U$2439 ( \2568 , \2561 , \2567 );
buf \U$2440 ( \2569 , \2568 );
buf \U$2441 ( \2570 , \2569 );
not \U$2442 ( \2571 , \2570 );
buf \U$2443 ( \2572 , \2571 );
buf \U$2444 ( \2573 , \2572 );
not \U$2445 ( \2574 , \2573 );
or \U$2446 ( \2575 , \2552 , \2574 );
buf \U$2447 ( \2576 , \2550 );
not \U$2448 ( \2577 , \2576 );
buf \U$2449 ( \2578 , \2569 );
nand \U$2450 ( \2579 , \2577 , \2578 );
buf \U$2451 ( \2580 , \2579 );
buf \U$2452 ( \2581 , \2580 );
nand \U$2453 ( \2582 , \2575 , \2581 );
buf \U$2454 ( \2583 , \2582 );
buf \U$2455 ( \2584 , \2583 );
buf \U$2456 ( \2585 , \861 );
not \U$2457 ( \2586 , \2585 );
buf \U$2458 ( \2587 , \1971 );
not \U$2459 ( \2588 , \2587 );
and \U$2460 ( \2589 , \2586 , \2588 );
buf \U$2461 ( \2590 , \283 );
not \U$2462 ( \2591 , \2590 );
buf \U$2463 ( \2592 , \2591 );
buf \U$2464 ( \2593 , \2592 );
buf \U$2465 ( \2594 , \251 );
nor \U$2466 ( \2595 , \2593 , \2594 );
buf \U$2467 ( \2596 , \2595 );
buf \U$2468 ( \2597 , \2596 );
nor \U$2469 ( \2598 , \2589 , \2597 );
buf \U$2470 ( \2599 , \2598 );
buf \U$2471 ( \2600 , \2599 );
not \U$2472 ( \2601 , \2600 );
buf \U$2473 ( \2602 , \2601 );
buf \U$2474 ( \2603 , \2602 );
not \U$2475 ( \2604 , \2603 );
buf \U$2476 ( \2605 , \1780 );
not \U$2477 ( \2606 , \2605 );
buf \U$2480 ( \2607 , \612 );
buf \U$2481 ( \2608 , \2607 );
not \U$2482 ( \2609 , \2608 );
or \U$2483 ( \2610 , \2606 , \2609 );
buf \U$2484 ( \2611 , \816 );
buf \U$2485 ( \2612 , \623 );
nand \U$2486 ( \2613 , \2611 , \2612 );
buf \U$2487 ( \2614 , \2613 );
buf \U$2488 ( \2615 , \2614 );
nand \U$2489 ( \2616 , \2610 , \2615 );
buf \U$2490 ( \2617 , \2616 );
buf \U$2491 ( \2618 , \2617 );
not \U$2492 ( \2619 , \2618 );
or \U$2493 ( \2620 , \2604 , \2619 );
buf \U$2494 ( \2621 , \2617 );
buf \U$2495 ( \2622 , \2602 );
or \U$2496 ( \2623 , \2621 , \2622 );
buf \U$2497 ( \2624 , \418 );
not \U$2498 ( \2625 , \2624 );
buf \U$2499 ( \2626 , \846 );
not \U$2500 ( \2627 , \2626 );
or \U$2501 ( \2628 , \2625 , \2627 );
buf \U$2502 ( \2629 , \2038 );
buf \U$2503 ( \2630 , \2046 );
nand \U$2504 ( \2631 , \2629 , \2630 );
buf \U$2505 ( \2632 , \2631 );
buf \U$2506 ( \2633 , \2632 );
nand \U$2507 ( \2634 , \2628 , \2633 );
buf \U$2508 ( \2635 , \2634 );
buf \U$2509 ( \2636 , \2635 );
nand \U$2510 ( \2637 , \2623 , \2636 );
buf \U$2511 ( \2638 , \2637 );
buf \U$2512 ( \2639 , \2638 );
nand \U$2513 ( \2640 , \2620 , \2639 );
buf \U$2514 ( \2641 , \2640 );
buf \U$2515 ( \2642 , \2641 );
xnor \U$2516 ( \2643 , \2584 , \2642 );
buf \U$2517 ( \2644 , \2643 );
buf \U$2518 ( \2645 , \2644 );
not \U$2519 ( \2646 , \2645 );
buf \U$2520 ( \2647 , \2646 );
buf \U$2521 ( \2648 , \2647 );
not \U$2522 ( \2649 , \2648 );
or \U$2523 ( \2650 , \2518 , \2649 );
buf \U$2524 ( \2651 , \2644 );
not \U$2525 ( \2652 , \2651 );
buf \U$2526 ( \2653 , \2513 );
not \U$2527 ( \2654 , \2653 );
or \U$2528 ( \2655 , \2652 , \2654 );
xor \U$2529 ( \2656 , \2521 , \2529 );
xor \U$2530 ( \2657 , \2656 , \2546 );
buf \U$2531 ( \2658 , \2657 );
buf \U$2532 ( \2659 , \2658 );
xor \U$2533 ( \2660 , \2617 , \2599 );
xnor \U$2534 ( \2661 , \2660 , \2635 );
buf \U$2535 ( \2662 , \2661 );
xor \U$2536 ( \2663 , \2659 , \2662 );
xor \U$2537 ( \2664 , \2264 , \2284 );
xor \U$2538 ( \2665 , \2664 , \2298 );
buf \U$2539 ( \2666 , \2665 );
buf \U$2540 ( \2667 , \2666 );
and \U$2541 ( \2668 , \2663 , \2667 );
and \U$2542 ( \2669 , \2659 , \2662 );
or \U$2543 ( \2670 , \2668 , \2669 );
buf \U$2544 ( \2671 , \2670 );
buf \U$2545 ( \2672 , \2671 );
nand \U$2546 ( \2673 , \2655 , \2672 );
buf \U$2547 ( \2674 , \2673 );
buf \U$2548 ( \2675 , \2674 );
nand \U$2549 ( \2676 , \2650 , \2675 );
buf \U$2550 ( \2677 , \2676 );
buf \U$2551 ( \2678 , \2677 );
xor \U$2552 ( \2679 , \2311 , \2678 );
xor \U$2553 ( \2680 , \545 , \591 );
and \U$2554 ( \2681 , \2680 , \646 );
and \U$2555 ( \2682 , \545 , \591 );
or \U$2556 ( \2683 , \2681 , \2682 );
buf \U$2557 ( \2684 , \2683 );
buf \U$2558 ( \2685 , \2684 );
buf \U$2559 ( \2686 , \2641 );
buf \U$2560 ( \2687 , \2550 );
or \U$2561 ( \2688 , \2686 , \2687 );
buf \U$2562 ( \2689 , \2569 );
nand \U$2563 ( \2690 , \2688 , \2689 );
buf \U$2564 ( \2691 , \2690 );
buf \U$2565 ( \2692 , \2691 );
buf \U$2566 ( \2693 , \2550 );
buf \U$2567 ( \2694 , \2641 );
nand \U$2568 ( \2695 , \2693 , \2694 );
buf \U$2569 ( \2696 , \2695 );
buf \U$2570 ( \2697 , \2696 );
nand \U$2571 ( \2698 , \2692 , \2697 );
buf \U$2572 ( \2699 , \2698 );
buf \U$2573 ( \2700 , \2699 );
xor \U$2574 ( \2701 , \2685 , \2700 );
xor \U$2575 ( \2702 , \2178 , \2249 );
and \U$2576 ( \2703 , \2702 , \2303 );
and \U$2577 ( \2704 , \2178 , \2249 );
or \U$2578 ( \2705 , \2703 , \2704 );
buf \U$2579 ( \2706 , \2705 );
buf \U$2580 ( \2707 , \2706 );
xor \U$2581 ( \2708 , \2701 , \2707 );
buf \U$2582 ( \2709 , \2708 );
buf \U$2583 ( \2710 , \2709 );
and \U$2584 ( \2711 , \2679 , \2710 );
and \U$2585 ( \2712 , \2311 , \2678 );
or \U$2586 ( \2713 , \2711 , \2712 );
buf \U$2587 ( \2714 , \2713 );
buf \U$2588 ( \2715 , \2714 );
xor \U$2589 ( \2716 , \2685 , \2700 );
and \U$2590 ( \2717 , \2716 , \2707 );
and \U$2591 ( \2718 , \2685 , \2700 );
or \U$2592 ( \2719 , \2717 , \2718 );
buf \U$2593 ( \2720 , \2719 );
buf \U$2594 ( \2721 , \2720 );
buf \U$2595 ( \2722 , \719 );
not \U$2596 ( \2723 , \2722 );
buf \U$2597 ( \2724 , \521 );
not \U$2598 ( \2725 , \2724 );
buf \U$2599 ( \2726 , \2725 );
buf \U$2600 ( \2727 , \2726 );
not \U$2601 ( \2728 , \2727 );
or \U$2602 ( \2729 , \2723 , \2728 );
buf \U$2603 ( \2730 , RIc0da0a8_91);
buf \U$2604 ( \2731 , RIc0d77e0_4);
xnor \U$2605 ( \2732 , \2730 , \2731 );
buf \U$2606 ( \2733 , \2732 );
buf \U$2607 ( \2734 , \2733 );
not \U$2608 ( \2735 , \2734 );
buf \U$2609 ( \2736 , \1933 );
nand \U$2610 ( \2737 , \2735 , \2736 );
buf \U$2611 ( \2738 , \2737 );
buf \U$2612 ( \2739 , \2738 );
nand \U$2613 ( \2740 , \2729 , \2739 );
buf \U$2614 ( \2741 , \2740 );
buf \U$2615 ( \2742 , \2741 );
buf \U$2616 ( \2743 , \1008 );
not \U$2617 ( \2744 , \2743 );
buf \U$2618 ( \2745 , \2744 );
buf \U$2619 ( \2746 , \2745 );
not \U$2620 ( \2747 , \2746 );
buf \U$2621 ( \2748 , \574 );
not \U$2622 ( \2749 , \2748 );
or \U$2623 ( \2750 , \2747 , \2749 );
buf \U$2624 ( \2751 , \993 );
buf \U$2625 ( \2752 , RIc0d7ba0_12);
buf \U$2626 ( \2753 , RIc0d9ce8_83);
xor \U$2627 ( \2754 , \2752 , \2753 );
buf \U$2628 ( \2755 , \2754 );
buf \U$2629 ( \2756 , \2755 );
nand \U$2630 ( \2757 , \2751 , \2756 );
buf \U$2631 ( \2758 , \2757 );
buf \U$2632 ( \2759 , \2758 );
nand \U$2633 ( \2760 , \2750 , \2759 );
buf \U$2634 ( \2761 , \2760 );
buf \U$2635 ( \2762 , \2761 );
xor \U$2636 ( \2763 , \2742 , \2762 );
buf \U$2637 ( \2764 , \1060 );
not \U$2638 ( \2765 , \2764 );
buf \U$2639 ( \2766 , \2765 );
buf \U$2640 ( \2767 , \2766 );
not \U$2641 ( \2768 , \2767 );
buf \U$2642 ( \2769 , \2768 );
buf \U$2643 ( \2770 , \2769 );
buf \U$2644 ( \2771 , \1071 );
or \U$2645 ( \2772 , \2770 , \2771 );
buf \U$2646 ( \2773 , \1078 );
not \U$2647 ( \2774 , \2773 );
buf \U$2648 ( \2775 , \2774 );
buf \U$2649 ( \2776 , \2775 );
buf \U$2650 ( \2777 , RIc0d7c90_14);
buf \U$2651 ( \2778 , RIc0d9bf8_81);
xnor \U$2652 ( \2779 , \2777 , \2778 );
buf \U$2653 ( \2780 , \2779 );
buf \U$2654 ( \2781 , \2780 );
or \U$2655 ( \2782 , \2776 , \2781 );
nand \U$2656 ( \2783 , \2772 , \2782 );
buf \U$2657 ( \2784 , \2783 );
buf \U$2658 ( \2785 , \2784 );
xor \U$2659 ( \2786 , \2763 , \2785 );
buf \U$2660 ( \2787 , \2786 );
buf \U$2661 ( \2788 , \2787 );
buf \U$2662 ( \2789 , \824 );
not \U$2663 ( \2790 , \2789 );
buf \U$2664 ( \2791 , \618 );
not \U$2665 ( \2792 , \2791 );
or \U$2666 ( \2793 , \2790 , \2792 );
buf \U$2667 ( \2794 , RIc0d79c0_8);
buf \U$2668 ( \2795 , RIc0d9ec8_87);
xnor \U$2669 ( \2796 , \2794 , \2795 );
buf \U$2670 ( \2797 , \2796 );
buf \U$2671 ( \2798 , \2797 );
not \U$2672 ( \2799 , \2798 );
buf \U$2673 ( \2800 , \816 );
nand \U$2674 ( \2801 , \2799 , \2800 );
buf \U$2675 ( \2802 , \2801 );
buf \U$2676 ( \2803 , \2802 );
nand \U$2677 ( \2804 , \2793 , \2803 );
buf \U$2678 ( \2805 , \2804 );
buf \U$2679 ( \2806 , \2805 );
not \U$2680 ( \2807 , \2806 );
buf \U$2681 ( \2808 , \2807 );
buf \U$2682 ( \2809 , \2808 );
buf \U$2683 ( \2810 , \1260 );
not \U$2684 ( \2811 , \2810 );
buf \U$2685 ( \2812 , \2811 );
buf \U$2686 ( \2813 , \2812 );
not \U$2687 ( \2814 , \2813 );
buf \U$2688 ( \2815 , \2814 );
buf \U$2689 ( \2816 , \2815 );
buf \U$2690 ( \2817 , \1270 );
or \U$2691 ( \2818 , \2816 , \2817 );
buf \U$2692 ( \2819 , \1279 );
buf \U$2693 ( \2820 , RIc0d8140_24);
buf \U$2694 ( \2821 , RIc0d9748_71);
xnor \U$2695 ( \2822 , \2820 , \2821 );
buf \U$2696 ( \2823 , \2822 );
buf \U$2697 ( \2824 , \2823 );
or \U$2698 ( \2825 , \2819 , \2824 );
nand \U$2699 ( \2826 , \2818 , \2825 );
buf \U$2700 ( \2827 , \2826 );
buf \U$2701 ( \2828 , \2827 );
xor \U$2702 ( \2829 , \2809 , \2828 );
buf \U$2703 ( \2830 , \1246 );
not \U$2704 ( \2831 , \2830 );
buf \U$2705 ( \2832 , \1202 );
not \U$2706 ( \2833 , \2832 );
or \U$2707 ( \2834 , \2831 , \2833 );
buf \U$2708 ( \2835 , \1202 );
buf \U$2709 ( \2836 , \1246 );
or \U$2710 ( \2837 , \2835 , \2836 );
buf \U$2711 ( \2838 , \1288 );
nand \U$2712 ( \2839 , \2837 , \2838 );
buf \U$2713 ( \2840 , \2839 );
buf \U$2714 ( \2841 , \2840 );
nand \U$2715 ( \2842 , \2834 , \2841 );
buf \U$2716 ( \2843 , \2842 );
buf \U$2717 ( \2844 , \2843 );
xor \U$2718 ( \2845 , \2829 , \2844 );
buf \U$2719 ( \2846 , \2845 );
buf \U$2720 ( \2847 , \2846 );
xor \U$2721 ( \2848 , \2788 , \2847 );
buf \U$2722 ( \2849 , \645 );
not \U$2723 ( \2850 , \2849 );
buf \U$2724 ( \2851 , \2850 );
buf \U$2725 ( \2852 , \2851 );
buf \U$2726 ( \2853 , \2256 );
not \U$2727 ( \2854 , \2853 );
buf \U$2728 ( \2855 , \1224 );
not \U$2729 ( \2856 , \2855 );
or \U$2730 ( \2857 , \2854 , \2856 );
buf \U$2731 ( \2858 , \1229 );
buf \U$2732 ( \2859 , \1206 );
nand \U$2733 ( \2860 , \2858 , \2859 );
buf \U$2734 ( \2861 , \2860 );
buf \U$2735 ( \2862 , \2861 );
nand \U$2736 ( \2863 , \2857 , \2862 );
buf \U$2737 ( \2864 , \2863 );
buf \U$2738 ( \2865 , \2864 );
not \U$2739 ( \2866 , \2865 );
buf \U$2740 ( \2867 , \2445 );
not \U$2741 ( \2868 , \2867 );
buf \U$2742 ( \2869 , \773 );
not \U$2743 ( \2870 , \2869 );
buf \U$2744 ( \2871 , \2870 );
buf \U$2745 ( \2872 , \2871 );
not \U$2746 ( \2873 , \2872 );
or \U$2747 ( \2874 , \2868 , \2873 );
buf \U$2748 ( \2875 , \784 );
not \U$2749 ( \2876 , \2875 );
buf \U$2750 ( \2877 , \791 );
not \U$2751 ( \2878 , \2877 );
buf \U$2752 ( \2879 , \2878 );
buf \U$2753 ( \2880 , \2879 );
not \U$2754 ( \2881 , \2880 );
buf \U$2755 ( \2882 , \2881 );
buf \U$2756 ( \2883 , \2882 );
nand \U$2757 ( \2884 , \2876 , \2883 );
buf \U$2758 ( \2885 , \2884 );
buf \U$2759 ( \2886 , \2885 );
nand \U$2760 ( \2887 , \2874 , \2886 );
buf \U$2761 ( \2888 , \2887 );
buf \U$2762 ( \2889 , \2888 );
not \U$2763 ( \2890 , \2889 );
or \U$2764 ( \2891 , \2866 , \2890 );
buf \U$2765 ( \2892 , \2864 );
buf \U$2766 ( \2893 , \2888 );
or \U$2767 ( \2894 , \2892 , \2893 );
buf \U$2768 ( \2895 , \2523 );
not \U$2769 ( \2896 , \2895 );
buf \U$2770 ( \2897 , \675 );
not \U$2771 ( \2898 , \2897 );
buf \U$2772 ( \2899 , \2898 );
buf \U$2775 ( \2900 , \2899 );
buf \U$2776 ( \2901 , \2900 );
not \U$2777 ( \2902 , \2901 );
or \U$2778 ( \2903 , \2896 , \2902 );
buf \U$2779 ( \2904 , \686 );
buf \U$2780 ( \2905 , \663 );
nand \U$2781 ( \2906 , \2904 , \2905 );
buf \U$2782 ( \2907 , \2906 );
buf \U$2783 ( \2908 , \2907 );
nand \U$2784 ( \2909 , \2903 , \2908 );
buf \U$2785 ( \2910 , \2909 );
buf \U$2786 ( \2911 , \2910 );
nand \U$2787 ( \2912 , \2894 , \2911 );
buf \U$2788 ( \2913 , \2912 );
buf \U$2789 ( \2914 , \2913 );
nand \U$2790 ( \2915 , \2891 , \2914 );
buf \U$2791 ( \2916 , \2915 );
buf \U$2792 ( \2917 , \2916 );
xor \U$2793 ( \2918 , \2852 , \2917 );
buf \U$2794 ( \2919 , \2277 );
not \U$2795 ( \2920 , \2919 );
buf \U$2796 ( \2921 , \1260 );
not \U$2797 ( \2922 , \2921 );
buf \U$2798 ( \2923 , \2922 );
buf \U$2799 ( \2924 , \2923 );
not \U$2800 ( \2925 , \2924 );
or \U$2801 ( \2926 , \2920 , \2925 );
buf \U$2804 ( \2927 , \1276 );
buf \U$2805 ( \2928 , \2927 );
buf \U$2806 ( \2929 , \1251 );
nand \U$2807 ( \2930 , \2928 , \2929 );
buf \U$2808 ( \2931 , \2930 );
buf \U$2809 ( \2932 , \2931 );
nand \U$2810 ( \2933 , \2926 , \2932 );
buf \U$2811 ( \2934 , \2933 );
buf \U$2812 ( \2935 , \2934 );
buf \U$2813 ( \2936 , \2431 );
not \U$2814 ( \2937 , \2936 );
buf \U$2817 ( \2938 , \748 );
buf \U$2818 ( \2939 , \2938 );
not \U$2819 ( \2940 , \2939 );
buf \U$2820 ( \2941 , \2940 );
buf \U$2821 ( \2942 , \2941 );
not \U$2822 ( \2943 , \2942 );
or \U$2823 ( \2944 , \2937 , \2943 );
buf \U$2824 ( \2945 , \734 );
buf \U$2825 ( \2946 , RIc0da378_97);
nand \U$2826 ( \2947 , \2945 , \2946 );
buf \U$2827 ( \2948 , \2947 );
buf \U$2828 ( \2949 , \2948 );
nand \U$2829 ( \2950 , \2944 , \2949 );
buf \U$2830 ( \2951 , \2950 );
buf \U$2831 ( \2952 , \2951 );
xor \U$2832 ( \2953 , \2935 , \2952 );
buf \U$2833 ( \2954 , \1389 );
not \U$2834 ( \2955 , \2954 );
buf \U$2835 ( \2956 , \2955 );
buf \U$2836 ( \2957 , \2956 );
buf \U$2837 ( \2958 , \2406 );
or \U$2838 ( \2959 , \2957 , \2958 );
buf \U$2841 ( \2960 , \915 );
buf \U$2842 ( \2961 , \2960 );
not \U$2843 ( \2962 , \2961 );
buf \U$2844 ( \2963 , \2962 );
buf \U$2845 ( \2964 , \2963 );
buf \U$2846 ( \2965 , \958 );
or \U$2847 ( \2966 , \2964 , \2965 );
nand \U$2848 ( \2967 , \2959 , \2966 );
buf \U$2849 ( \2968 , \2967 );
buf \U$2850 ( \2969 , \2968 );
and \U$2851 ( \2970 , \2953 , \2969 );
and \U$2852 ( \2971 , \2935 , \2952 );
or \U$2853 ( \2972 , \2970 , \2971 );
buf \U$2854 ( \2973 , \2972 );
buf \U$2855 ( \2974 , \2973 );
and \U$2856 ( \2975 , \2918 , \2974 );
and \U$2857 ( \2976 , \2852 , \2917 );
or \U$2858 ( \2977 , \2975 , \2976 );
buf \U$2859 ( \2978 , \2977 );
buf \U$2860 ( \2979 , \2978 );
xor \U$2861 ( \2980 , \2848 , \2979 );
buf \U$2862 ( \2981 , \2980 );
buf \U$2863 ( \2982 , \2981 );
xor \U$2864 ( \2983 , \2721 , \2982 );
xor \U$2865 ( \2984 , \2852 , \2917 );
xor \U$2866 ( \2985 , \2984 , \2974 );
buf \U$2867 ( \2986 , \2985 );
buf \U$2868 ( \2987 , \2986 );
xor \U$2869 ( \2988 , \1573 , \1596 );
xor \U$2870 ( \2989 , \2988 , \1619 );
buf \U$2871 ( \2990 , \2989 );
buf \U$2872 ( \2991 , \2990 );
not \U$2873 ( \2992 , \2991 );
xor \U$2874 ( \2993 , \2888 , \2864 );
xnor \U$2875 ( \2994 , \2993 , \2910 );
buf \U$2876 ( \2995 , \2994 );
not \U$2877 ( \2996 , \2995 );
buf \U$2878 ( \2997 , \2996 );
buf \U$2879 ( \2998 , \2997 );
not \U$2880 ( \2999 , \2998 );
or \U$2881 ( \3000 , \2992 , \2999 );
buf \U$2882 ( \3001 , \2997 );
buf \U$2883 ( \3002 , \2990 );
or \U$2884 ( \3003 , \3001 , \3002 );
xor \U$2885 ( \3004 , \2935 , \2952 );
xor \U$2886 ( \3005 , \3004 , \2969 );
buf \U$2887 ( \3006 , \3005 );
buf \U$2888 ( \3007 , \3006 );
nand \U$2889 ( \3008 , \3003 , \3007 );
buf \U$2890 ( \3009 , \3008 );
buf \U$2891 ( \3010 , \3009 );
nand \U$2892 ( \3011 , \3000 , \3010 );
buf \U$2893 ( \3012 , \3011 );
buf \U$2894 ( \3013 , \3012 );
xor \U$2895 ( \3014 , \2987 , \3013 );
xor \U$2896 ( \3015 , \1531 , \1546 );
xor \U$2897 ( \3016 , \3015 , \1624 );
buf \U$2898 ( \3017 , \3016 );
buf \U$2899 ( \3018 , \3017 );
and \U$2900 ( \3019 , \3014 , \3018 );
and \U$2901 ( \3020 , \2987 , \3013 );
or \U$2902 ( \3021 , \3019 , \3020 );
buf \U$2903 ( \3022 , \3021 );
buf \U$2904 ( \3023 , \3022 );
xor \U$2905 ( \3024 , \2983 , \3023 );
buf \U$2906 ( \3025 , \3024 );
buf \U$2907 ( \3026 , \3025 );
xor \U$2908 ( \3027 , \2715 , \3026 );
xor \U$2909 ( \3028 , \2987 , \3013 );
xor \U$2910 ( \3029 , \3028 , \3018 );
buf \U$2911 ( \3030 , \3029 );
buf \U$2912 ( \3031 , \3030 );
xor \U$2913 ( \3032 , \366 , \501 );
xor \U$2914 ( \3033 , \3032 , \649 );
buf \U$2915 ( \3034 , \3033 );
buf \U$2916 ( \3035 , \3034 );
not \U$2917 ( \3036 , \3035 );
buf \U$2918 ( \3037 , \2994 );
not \U$2919 ( \3038 , \3037 );
buf \U$2920 ( \3039 , \3006 );
not \U$2921 ( \3040 , \3039 );
or \U$2922 ( \3041 , \3038 , \3040 );
buf \U$2923 ( \3042 , \2994 );
buf \U$2924 ( \3043 , \3006 );
or \U$2925 ( \3044 , \3042 , \3043 );
nand \U$2926 ( \3045 , \3041 , \3044 );
buf \U$2927 ( \3046 , \3045 );
buf \U$2928 ( \3047 , \3046 );
buf \U$2929 ( \3048 , \2990 );
and \U$2930 ( \3049 , \3047 , \3048 );
not \U$2931 ( \3050 , \3047 );
buf \U$2932 ( \3051 , \2990 );
not \U$2933 ( \3052 , \3051 );
buf \U$2934 ( \3053 , \3052 );
buf \U$2935 ( \3054 , \3053 );
and \U$2936 ( \3055 , \3050 , \3054 );
nor \U$2937 ( \3056 , \3049 , \3055 );
buf \U$2938 ( \3057 , \3056 );
buf \U$2939 ( \3058 , \3057 );
not \U$2940 ( \3059 , \3058 );
or \U$2941 ( \3060 , \3036 , \3059 );
buf \U$2942 ( \3061 , \3034 );
buf \U$2943 ( \3062 , \3057 );
or \U$2944 ( \3063 , \3061 , \3062 );
xor \U$2945 ( \3064 , \2152 , \2134 );
xor \U$2946 ( \3065 , \3064 , \2171 );
buf \U$2947 ( \3066 , \3065 );
buf \U$2948 ( \3067 , \2216 );
not \U$2949 ( \3068 , \3067 );
buf \U$2950 ( \3069 , \2245 );
nand \U$2951 ( \3070 , \3068 , \3069 );
buf \U$2952 ( \3071 , \3070 );
buf \U$2953 ( \3072 , \3071 );
buf \U$2954 ( \3073 , \2236 );
and \U$2955 ( \3074 , \3072 , \3073 );
not \U$2956 ( \3075 , \3072 );
buf \U$2957 ( \3076 , \2239 );
and \U$2958 ( \3077 , \3075 , \3076 );
or \U$2959 ( \3078 , \3074 , \3077 );
buf \U$2960 ( \3079 , \3078 );
buf \U$2961 ( \3080 , \3079 );
xor \U$2962 ( \3081 , \3066 , \3080 );
xor \U$2963 ( \3082 , \1762 , \1790 );
xor \U$2964 ( \3083 , \3082 , \1868 );
buf \U$2965 ( \3084 , \3083 );
buf \U$2966 ( \3085 , \3084 );
and \U$2967 ( \3086 , \3081 , \3085 );
and \U$2968 ( \3087 , \3066 , \3080 );
or \U$2969 ( \3088 , \3086 , \3087 );
buf \U$2970 ( \3089 , \3088 );
buf \U$2971 ( \3090 , \3089 );
nand \U$2972 ( \3091 , \3063 , \3090 );
buf \U$2973 ( \3092 , \3091 );
buf \U$2974 ( \3093 , \3092 );
nand \U$2975 ( \3094 , \3060 , \3093 );
buf \U$2976 ( \3095 , \3094 );
buf \U$2977 ( \3096 , \3095 );
xor \U$2978 ( \3097 , \3031 , \3096 );
xor \U$2979 ( \3098 , \654 , \910 );
xor \U$2980 ( \3099 , \3098 , \1300 );
buf \U$2981 ( \3100 , \3099 );
buf \U$2982 ( \3101 , \3100 );
and \U$2983 ( \3102 , \3097 , \3101 );
and \U$2984 ( \3103 , \3031 , \3096 );
or \U$2985 ( \3104 , \3102 , \3103 );
buf \U$2986 ( \3105 , \3104 );
buf \U$2987 ( \3106 , \3105 );
xor \U$2988 ( \3107 , \3027 , \3106 );
buf \U$2989 ( \3108 , \3107 );
buf \U$2990 ( \3109 , \3108 );
xor \U$2991 ( \3110 , \1735 , \3109 );
xor \U$2992 ( \3111 , \1951 , \2026 );
xor \U$2993 ( \3112 , \3111 , \2109 );
buf \U$2994 ( \3113 , \3112 );
buf \U$2995 ( \3114 , \3113 );
xor \U$2996 ( \3115 , \1964 , \1980 );
xor \U$2997 ( \3116 , \3115 , \2014 );
buf \U$2998 ( \3117 , \3116 );
not \U$2999 ( \3118 , \3117 );
xor \U$3000 ( \3119 , \1813 , \1839 );
xor \U$3001 ( \3120 , \3119 , \1863 );
buf \U$3002 ( \3121 , \3120 );
buf \U$3003 ( \3122 , \3121 );
not \U$3004 ( \3123 , \3122 );
or \U$3005 ( \3124 , \3118 , \3123 );
buf \U$3006 ( \3125 , \3121 );
buf \U$3007 ( \3126 , \3116 );
or \U$3008 ( \3127 , \3125 , \3126 );
xor \U$3009 ( \3128 , \2053 , \2086 );
xor \U$3010 ( \3129 , \3128 , \2104 );
buf \U$3011 ( \3130 , \3129 );
buf \U$3012 ( \3131 , \3130 );
nand \U$3013 ( \3132 , \3127 , \3131 );
buf \U$3014 ( \3133 , \3132 );
buf \U$3015 ( \3134 , \3133 );
nand \U$3016 ( \3135 , \3124 , \3134 );
buf \U$3017 ( \3136 , \3135 );
buf \U$3018 ( \3137 , \3136 );
or \U$3019 ( \3138 , \3114 , \3137 );
buf \U$3020 ( \3139 , RIc0d8500_32);
buf \U$3021 ( \3140 , RIc0d9658_69);
xor \U$3022 ( \3141 , \3139 , \3140 );
buf \U$3023 ( \3142 , \3141 );
buf \U$3024 ( \3143 , \3142 );
not \U$3025 ( \3144 , \3143 );
buf \U$3026 ( \3145 , \279 );
not \U$3027 ( \3146 , \3145 );
or \U$3028 ( \3147 , \3144 , \3146 );
buf \U$3029 ( \3148 , \1978 );
not \U$3030 ( \3149 , \3148 );
buf \U$3031 ( \3150 , \284 );
nand \U$3032 ( \3151 , \3149 , \3150 );
buf \U$3033 ( \3152 , \3151 );
buf \U$3034 ( \3153 , \3152 );
nand \U$3035 ( \3154 , \3147 , \3153 );
buf \U$3036 ( \3155 , \3154 );
buf \U$3037 ( \3156 , \3155 );
not \U$3038 ( \3157 , \3156 );
buf \U$3039 ( \3158 , \3157 );
buf \U$3040 ( \3159 , \3158 );
not \U$3041 ( \3160 , \3159 );
buf \U$3042 ( \3161 , RIc0d8320_28);
buf \U$3043 ( \3162 , RIc0d9838_73);
xor \U$3044 ( \3163 , \3161 , \3162 );
buf \U$3045 ( \3164 , \3163 );
buf \U$3046 ( \3165 , \3164 );
not \U$3047 ( \3166 , \3165 );
buf \U$3048 ( \3167 , \776 );
not \U$3049 ( \3168 , \3167 );
or \U$3050 ( \3169 , \3166 , \3168 );
buf \U$3051 ( \3170 , \792 );
buf \U$3052 ( \3171 , \1844 );
nand \U$3053 ( \3172 , \3170 , \3171 );
buf \U$3054 ( \3173 , \3172 );
buf \U$3055 ( \3174 , \3173 );
nand \U$3056 ( \3175 , \3169 , \3174 );
buf \U$3057 ( \3176 , \3175 );
buf \U$3058 ( \3177 , \3176 );
not \U$3059 ( \3178 , \3177 );
buf \U$3060 ( \3179 , \3178 );
buf \U$3061 ( \3180 , \3179 );
not \U$3062 ( \3181 , \3180 );
or \U$3063 ( \3182 , \3160 , \3181 );
buf \U$3064 ( \3183 , \812 );
buf \U$3065 ( \3184 , RIc0d9ec8_87);
buf \U$3066 ( \3185 , RIc0d7c90_14);
xnor \U$3067 ( \3186 , \3184 , \3185 );
buf \U$3068 ( \3187 , \3186 );
buf \U$3069 ( \3188 , \3187 );
or \U$3070 ( \3189 , \3183 , \3188 );
buf \U$3071 ( \3190 , \819 );
buf \U$3072 ( \3191 , \1771 );
or \U$3073 ( \3192 , \3190 , \3191 );
nand \U$3074 ( \3193 , \3189 , \3192 );
buf \U$3075 ( \3194 , \3193 );
buf \U$3076 ( \3195 , \3194 );
nand \U$3077 ( \3196 , \3182 , \3195 );
buf \U$3078 ( \3197 , \3196 );
buf \U$3079 ( \3198 , \3197 );
buf \U$3080 ( \3199 , \3176 );
buf \U$3081 ( \3200 , \3155 );
nand \U$3082 ( \3201 , \3199 , \3200 );
buf \U$3083 ( \3202 , \3201 );
buf \U$3084 ( \3203 , \3202 );
nand \U$3085 ( \3204 , \3198 , \3203 );
buf \U$3086 ( \3205 , \3204 );
buf \U$3087 ( \3206 , \3205 );
xor \U$3088 ( \3207 , \1890 , \1944 );
xor \U$3089 ( \3208 , \3207 , \1912 );
buf \U$3090 ( \3209 , \3208 );
xor \U$3091 ( \3210 , \3206 , \3209 );
buf \U$3092 ( \3211 , \2349 );
not \U$3093 ( \3212 , \3211 );
buf \U$3094 ( \3213 , \2328 );
not \U$3095 ( \3214 , \3213 );
or \U$3096 ( \3215 , \3212 , \3214 );
buf \U$3097 ( \3216 , \2328 );
buf \U$3098 ( \3217 , \2349 );
or \U$3099 ( \3218 , \3216 , \3217 );
nand \U$3100 ( \3219 , \3215 , \3218 );
buf \U$3101 ( \3220 , \3219 );
xor \U$3102 ( \3221 , \2380 , \3220 );
buf \U$3103 ( \3222 , \3221 );
and \U$3104 ( \3223 , \3210 , \3222 );
and \U$3105 ( \3224 , \3206 , \3209 );
or \U$3106 ( \3225 , \3223 , \3224 );
buf \U$3107 ( \3226 , \3225 );
buf \U$3108 ( \3227 , \3226 );
nand \U$3109 ( \3228 , \3138 , \3227 );
buf \U$3110 ( \3229 , \3228 );
buf \U$3111 ( \3230 , \3229 );
buf \U$3112 ( \3231 , \3113 );
buf \U$3113 ( \3232 , \3136 );
nand \U$3114 ( \3233 , \3231 , \3232 );
buf \U$3115 ( \3234 , \3233 );
buf \U$3116 ( \3235 , \3234 );
nand \U$3117 ( \3236 , \3230 , \3235 );
buf \U$3118 ( \3237 , \3236 );
buf \U$3119 ( \3238 , \3237 );
buf \U$3120 ( \3239 , \1786 );
buf \U$3121 ( \3240 , RIc0d9478_65);
buf \U$3122 ( \3241 , RIc0d8758_37);
and \U$3123 ( \3242 , \3240 , \3241 );
buf \U$3124 ( \3243 , \3242 );
buf \U$3125 ( \3244 , \3243 );
buf \U$3126 ( \3245 , RIc0d85f0_34);
buf \U$3127 ( \3246 , RIc0d9568_67);
xor \U$3128 ( \3247 , \3245 , \3246 );
buf \U$3129 ( \3248 , \3247 );
buf \U$3130 ( \3249 , \3248 );
not \U$3131 ( \3250 , \3249 );
buf \U$3132 ( \3251 , \2900 );
not \U$3133 ( \3252 , \3251 );
or \U$3134 ( \3253 , \3250 , \3252 );
buf \U$3135 ( \3254 , \686 );
buf \U$3136 ( \3255 , \1817 );
nand \U$3137 ( \3256 , \3254 , \3255 );
buf \U$3138 ( \3257 , \3256 );
buf \U$3139 ( \3258 , \3257 );
nand \U$3140 ( \3259 , \3253 , \3258 );
buf \U$3141 ( \3260 , \3259 );
buf \U$3142 ( \3261 , \3260 );
xor \U$3143 ( \3262 , \3244 , \3261 );
buf \U$3144 ( \3263 , \521 );
buf \U$3145 ( \3264 , RIc0da0a8_91);
buf \U$3146 ( \3265 , RIc0d7ab0_10);
xnor \U$3147 ( \3266 , \3264 , \3265 );
buf \U$3148 ( \3267 , \3266 );
buf \U$3149 ( \3268 , \3267 );
or \U$3150 ( \3269 , \3263 , \3268 );
buf \U$3151 ( \3270 , \711 );
buf \U$3152 ( \3271 , \1922 );
not \U$3153 ( \3272 , \3271 );
buf \U$3154 ( \3273 , \3272 );
buf \U$3155 ( \3274 , \3273 );
or \U$3156 ( \3275 , \3270 , \3274 );
nand \U$3157 ( \3276 , \3269 , \3275 );
buf \U$3158 ( \3277 , \3276 );
buf \U$3159 ( \3278 , \3277 );
and \U$3160 ( \3279 , \3262 , \3278 );
and \U$3161 ( \3280 , \3244 , \3261 );
or \U$3162 ( \3281 , \3279 , \3280 );
buf \U$3163 ( \3282 , \3281 );
buf \U$3164 ( \3283 , \3282 );
xor \U$3165 ( \3284 , \3239 , \3283 );
buf \U$3166 ( \3285 , RIc0d9dd8_85);
buf \U$3167 ( \3286 , RIc0d7d80_16);
xnor \U$3168 ( \3287 , \3285 , \3286 );
buf \U$3169 ( \3288 , \3287 );
buf \U$3170 ( \3289 , \3288 );
buf \U$3171 ( \3290 , \948 );
not \U$3172 ( \3291 , \3290 );
buf \U$3173 ( \3292 , \3291 );
buf \U$3174 ( \3293 , \3292 );
not \U$3175 ( \3294 , \3293 );
buf \U$3176 ( \3295 , \3294 );
buf \U$3177 ( \3296 , \3295 );
or \U$3178 ( \3297 , \3289 , \3296 );
buf \U$3179 ( \3298 , \2963 );
buf \U$3180 ( \3299 , \2314 );
or \U$3181 ( \3300 , \3298 , \3299 );
nand \U$3182 ( \3301 , \3297 , \3300 );
buf \U$3183 ( \3302 , \3301 );
buf \U$3184 ( \3303 , \3302 );
not \U$3185 ( \3304 , \3303 );
buf \U$3186 ( \3305 , RIc0da378_97);
buf \U$3187 ( \3306 , RIc0d77e0_4);
and \U$3188 ( \3307 , \3305 , \3306 );
not \U$3189 ( \3308 , \3305 );
buf \U$3190 ( \3309 , \489 );
and \U$3191 ( \3310 , \3308 , \3309 );
nor \U$3192 ( \3311 , \3307 , \3310 );
buf \U$3193 ( \3312 , \3311 );
buf \U$3194 ( \3313 , \3312 );
not \U$3195 ( \3314 , \3313 );
buf \U$3196 ( \3315 , \2066 );
not \U$3197 ( \3316 , \3315 );
or \U$3198 ( \3317 , \3314 , \3316 );
buf \U$3199 ( \3318 , \734 );
buf \U$3200 ( \3319 , \2061 );
nand \U$3201 ( \3320 , \3318 , \3319 );
buf \U$3202 ( \3321 , \3320 );
buf \U$3203 ( \3322 , \3321 );
nand \U$3204 ( \3323 , \3317 , \3322 );
buf \U$3205 ( \3324 , \3323 );
buf \U$3206 ( \3325 , \3324 );
not \U$3207 ( \3326 , \3325 );
or \U$3208 ( \3327 , \3304 , \3326 );
buf \U$3209 ( \3328 , \3324 );
buf \U$3210 ( \3329 , \3302 );
or \U$3211 ( \3330 , \3328 , \3329 );
buf \U$3212 ( \3331 , RIc0d7e70_18);
buf \U$3213 ( \3332 , RIc0d9ce8_83);
xor \U$3214 ( \3333 , \3331 , \3332 );
buf \U$3215 ( \3334 , \3333 );
buf \U$3216 ( \3335 , \3334 );
not \U$3217 ( \3336 , \3335 );
buf \U$3218 ( \3337 , \1736 );
not \U$3219 ( \3338 , \3337 );
or \U$3220 ( \3339 , \3336 , \3338 );
buf \U$3221 ( \3340 , \2096 );
not \U$3222 ( \3341 , \3340 );
buf \U$3223 ( \3342 , \993 );
nand \U$3224 ( \3343 , \3341 , \3342 );
buf \U$3225 ( \3344 , \3343 );
buf \U$3226 ( \3345 , \3344 );
nand \U$3227 ( \3346 , \3339 , \3345 );
buf \U$3228 ( \3347 , \3346 );
buf \U$3229 ( \3348 , \3347 );
nand \U$3230 ( \3349 , \3330 , \3348 );
buf \U$3231 ( \3350 , \3349 );
buf \U$3232 ( \3351 , \3350 );
nand \U$3233 ( \3352 , \3327 , \3351 );
buf \U$3234 ( \3353 , \3352 );
buf \U$3235 ( \3354 , \3353 );
and \U$3236 ( \3355 , \3284 , \3354 );
and \U$3237 ( \3356 , \3239 , \3283 );
or \U$3238 ( \3357 , \3355 , \3356 );
buf \U$3239 ( \3358 , \3357 );
buf \U$3240 ( \3359 , \3358 );
buf \U$3241 ( \3360 , RIc0d8050_22);
buf \U$3242 ( \3361 , RIc0d9b08_79);
xor \U$3243 ( \3362 , \3360 , \3361 );
buf \U$3244 ( \3363 , \3362 );
buf \U$3245 ( \3364 , \3363 );
not \U$3246 ( \3365 , \3364 );
buf \U$3247 ( \3366 , \397 );
not \U$3248 ( \3367 , \3366 );
or \U$3249 ( \3368 , \3365 , \3367 );
buf \U$3250 ( \3369 , \2490 );
not \U$3251 ( \3370 , \3369 );
buf \U$3252 ( \3371 , \1026 );
nand \U$3253 ( \3372 , \3370 , \3371 );
buf \U$3254 ( \3373 , \3372 );
buf \U$3255 ( \3374 , \3373 );
nand \U$3256 ( \3375 , \3368 , \3374 );
buf \U$3257 ( \3376 , \3375 );
buf \U$3258 ( \3377 , \3376 );
not \U$3259 ( \3378 , \3377 );
buf \U$3260 ( \3379 , \3378 );
buf \U$3261 ( \3380 , \3379 );
not \U$3262 ( \3381 , \3380 );
buf \U$3263 ( \3382 , \2034 );
not \U$3264 ( \3383 , \3382 );
buf \U$3265 ( \3384 , \3383 );
buf \U$3266 ( \3385 , \3384 );
not \U$3267 ( \3386 , \3385 );
buf \U$3268 ( \3387 , \3386 );
buf \U$3269 ( \3388 , \3387 );
not \U$3270 ( \3389 , \3388 );
buf \U$3271 ( \3390 , RIc0d9fb8_89);
buf \U$3272 ( \3391 , RIc0d7ba0_12);
xnor \U$3273 ( \3392 , \3390 , \3391 );
buf \U$3274 ( \3393 , \3392 );
buf \U$3275 ( \3394 , \3393 );
not \U$3276 ( \3395 , \3394 );
and \U$3277 ( \3396 , \3389 , \3395 );
buf \U$3278 ( \3397 , \442 );
buf \U$3279 ( \3398 , \2031 );
and \U$3280 ( \3399 , \3397 , \3398 );
buf \U$3281 ( \3400 , \3399 );
buf \U$3282 ( \3401 , \3400 );
nor \U$3283 ( \3402 , \3396 , \3401 );
buf \U$3284 ( \3403 , \3402 );
buf \U$3285 ( \3404 , \3403 );
not \U$3286 ( \3405 , \3404 );
or \U$3287 ( \3406 , \3381 , \3405 );
buf \U$3288 ( \3407 , RIc0d79c0_8);
buf \U$3289 ( \3408 , RIc0da198_93);
xor \U$3290 ( \3409 , \3407 , \3408 );
buf \U$3291 ( \3410 , \3409 );
buf \U$3292 ( \3411 , \3410 );
not \U$3293 ( \3412 , \3411 );
buf \U$3294 ( \3413 , \473 );
not \U$3295 ( \3414 , \3413 );
buf \U$3296 ( \3415 , \3414 );
buf \U$3297 ( \3416 , \3415 );
not \U$3298 ( \3417 , \3416 );
or \U$3299 ( \3418 , \3412 , \3417 );
buf \U$3300 ( \3419 , \481 );
buf \U$3301 ( \3420 , \1896 );
nand \U$3302 ( \3421 , \3419 , \3420 );
buf \U$3303 ( \3422 , \3421 );
buf \U$3304 ( \3423 , \3422 );
nand \U$3305 ( \3424 , \3418 , \3423 );
buf \U$3306 ( \3425 , \3424 );
buf \U$3307 ( \3426 , \3425 );
nand \U$3308 ( \3427 , \3406 , \3426 );
buf \U$3309 ( \3428 , \3427 );
buf \U$3310 ( \3429 , \3428 );
buf \U$3311 ( \3430 , \3403 );
not \U$3312 ( \3431 , \3430 );
buf \U$3313 ( \3432 , \3376 );
nand \U$3314 ( \3433 , \3431 , \3432 );
buf \U$3315 ( \3434 , \3433 );
buf \U$3316 ( \3435 , \3434 );
nand \U$3317 ( \3436 , \3429 , \3435 );
buf \U$3318 ( \3437 , \3436 );
buf \U$3319 ( \3438 , \3437 );
buf \U$3320 ( \3439 , RIc0d8230_26);
buf \U$3321 ( \3440 , RIc0d9928_75);
xnor \U$3322 ( \3441 , \3439 , \3440 );
buf \U$3323 ( \3442 , \3441 );
buf \U$3324 ( \3443 , \3442 );
not \U$3325 ( \3444 , \3443 );
buf \U$3326 ( \3445 , \3444 );
buf \U$3327 ( \3446 , \3445 );
not \U$3328 ( \3447 , \3446 );
buf \U$3329 ( \3448 , \1129 );
not \U$3330 ( \3449 , \3448 );
or \U$3331 ( \3450 , \3447 , \3449 );
buf \U$3332 ( \3451 , \2367 );
not \U$3333 ( \3452 , \3451 );
buf \U$3334 ( \3453 , \1565 );
nand \U$3335 ( \3454 , \3452 , \3453 );
buf \U$3336 ( \3455 , \3454 );
buf \U$3337 ( \3456 , \3455 );
nand \U$3338 ( \3457 , \3450 , \3456 );
buf \U$3339 ( \3458 , \3457 );
buf \U$3340 ( \3459 , \3458 );
not \U$3341 ( \3460 , \3459 );
buf \U$3342 ( \3461 , RIc0d8140_24);
buf \U$3343 ( \3462 , RIc0d9a18_77);
xor \U$3344 ( \3463 , \3461 , \3462 );
buf \U$3345 ( \3464 , \3463 );
buf \U$3346 ( \3465 , \3464 );
not \U$3347 ( \3466 , \3465 );
buf \U$3348 ( \3467 , \1183 );
not \U$3349 ( \3468 , \3467 );
or \U$3350 ( \3469 , \3466 , \3468 );
buf \U$3351 ( \3470 , \1196 );
buf \U$3352 ( \3471 , \2337 );
nand \U$3353 ( \3472 , \3470 , \3471 );
buf \U$3354 ( \3473 , \3472 );
buf \U$3355 ( \3474 , \3473 );
nand \U$3356 ( \3475 , \3469 , \3474 );
buf \U$3357 ( \3476 , \3475 );
buf \U$3358 ( \3477 , \3476 );
not \U$3359 ( \3478 , \3477 );
or \U$3360 ( \3479 , \3460 , \3478 );
buf \U$3361 ( \3480 , \3476 );
buf \U$3362 ( \3481 , \3458 );
or \U$3363 ( \3482 , \3480 , \3481 );
buf \U$3364 ( \3483 , RIc0da468_99);
buf \U$3365 ( \3484 , RIc0d76f0_2);
and \U$3366 ( \3485 , \3483 , \3484 );
not \U$3367 ( \3486 , \3483 );
buf \U$3368 ( \3487 , \352 );
and \U$3369 ( \3488 , \3486 , \3487 );
nor \U$3370 ( \3489 , \3485 , \3488 );
buf \U$3371 ( \3490 , \3489 );
buf \U$3372 ( \3491 , \3490 );
not \U$3373 ( \3492 , \3491 );
buf \U$3374 ( \3493 , \2470 );
not \U$3375 ( \3494 , \3493 );
or \U$3376 ( \3495 , \3492 , \3494 );
buf \U$3377 ( \3496 , \2476 );
buf \U$3378 ( \3497 , \2465 );
nand \U$3379 ( \3498 , \3496 , \3497 );
buf \U$3380 ( \3499 , \3498 );
buf \U$3381 ( \3500 , \3499 );
nand \U$3382 ( \3501 , \3495 , \3500 );
buf \U$3383 ( \3502 , \3501 );
buf \U$3384 ( \3503 , \3502 );
nand \U$3385 ( \3504 , \3482 , \3503 );
buf \U$3386 ( \3505 , \3504 );
buf \U$3387 ( \3506 , \3505 );
nand \U$3388 ( \3507 , \3479 , \3506 );
buf \U$3389 ( \3508 , \3507 );
buf \U$3390 ( \3509 , \3508 );
xor \U$3391 ( \3510 , \3438 , \3509 );
buf \U$3392 ( \3511 , RIc0da5d0_102);
buf \U$3393 ( \3512 , RIc0da648_103);
xor \U$3394 ( \3513 , \3511 , \3512 );
buf \U$3395 ( \3514 , \3513 );
buf \U$3398 ( \3515 , \3514 );
buf \U$3399 ( \3516 , \3515 );
not \U$3400 ( \3517 , \3516 );
buf \U$3401 ( \3518 , \3517 );
buf \U$3402 ( \3519 , \3518 );
not \U$3403 ( \3520 , \3519 );
xor \U$3404 ( \3521 , RIc0da558_101, RIc0da5d0_102);
buf \U$3405 ( \3522 , \3521 );
buf \U$3406 ( \3523 , \3514 );
not \U$3407 ( \3524 , \3523 );
buf \U$3408 ( \3525 , \3524 );
buf \U$3409 ( \3526 , \3525 );
and \U$3410 ( \3527 , \3522 , \3526 );
buf \U$3411 ( \3528 , \3527 );
buf \U$3412 ( \3529 , \3528 );
not \U$3413 ( \3530 , \3529 );
buf \U$3414 ( \3531 , \3530 );
buf \U$3415 ( \3532 , \3531 );
not \U$3416 ( \3533 , \3532 );
buf \U$3417 ( \3534 , \3533 );
buf \U$3420 ( \3535 , \3534 );
buf \U$3421 ( \3536 , \3535 );
not \U$3422 ( \3537 , \3536 );
buf \U$3423 ( \3538 , \3537 );
buf \U$3424 ( \3539 , \3538 );
not \U$3425 ( \3540 , \3539 );
or \U$3426 ( \3541 , \3520 , \3540 );
buf \U$3427 ( \3542 , RIc0da558_101);
nand \U$3428 ( \3543 , \3541 , \3542 );
buf \U$3429 ( \3544 , \3543 );
buf \U$3430 ( \3545 , \3544 );
buf \U$3431 ( \3546 , RIc0d78d0_6);
buf \U$3432 ( \3547 , RIc0da288_95);
xor \U$3433 ( \3548 , \3546 , \3547 );
buf \U$3434 ( \3549 , \3548 );
buf \U$3435 ( \3550 , \3549 );
not \U$3436 ( \3551 , \3550 );
buf \U$3437 ( \3552 , \330 );
not \U$3438 ( \3553 , \3552 );
or \U$3439 ( \3554 , \3551 , \3553 );
buf \U$3440 ( \3555 , \344 );
buf \U$3441 ( \3556 , \1994 );
nand \U$3442 ( \3557 , \3555 , \3556 );
buf \U$3443 ( \3558 , \3557 );
buf \U$3444 ( \3559 , \3558 );
nand \U$3445 ( \3560 , \3554 , \3559 );
buf \U$3446 ( \3561 , \3560 );
buf \U$3447 ( \3562 , \3561 );
xor \U$3448 ( \3563 , \3545 , \3562 );
buf \U$3449 ( \3564 , \1064 );
not \U$3450 ( \3565 , \3564 );
buf \U$3451 ( \3566 , \3565 );
buf \U$3452 ( \3567 , \3566 );
buf \U$3453 ( \3568 , RIc0d9bf8_81);
buf \U$3454 ( \3569 , RIc0d7f60_20);
xnor \U$3455 ( \3570 , \3568 , \3569 );
buf \U$3456 ( \3571 , \3570 );
buf \U$3457 ( \3572 , \3571 );
or \U$3458 ( \3573 , \3567 , \3572 );
buf \U$3459 ( \3574 , \2775 );
buf \U$3460 ( \3575 , \1956 );
or \U$3461 ( \3576 , \3574 , \3575 );
nand \U$3462 ( \3577 , \3573 , \3576 );
buf \U$3463 ( \3578 , \3577 );
buf \U$3464 ( \3579 , \3578 );
and \U$3465 ( \3580 , \3563 , \3579 );
and \U$3466 ( \3581 , \3545 , \3562 );
or \U$3467 ( \3582 , \3580 , \3581 );
buf \U$3468 ( \3583 , \3582 );
buf \U$3469 ( \3584 , \3583 );
and \U$3470 ( \3585 , \3510 , \3584 );
and \U$3471 ( \3586 , \3438 , \3509 );
or \U$3472 ( \3587 , \3585 , \3586 );
buf \U$3473 ( \3588 , \3587 );
buf \U$3474 ( \3589 , \3588 );
xor \U$3475 ( \3590 , \3359 , \3589 );
xor \U$3476 ( \3591 , \2386 , \2503 );
xnor \U$3477 ( \3592 , \3591 , \2448 );
buf \U$3478 ( \3593 , \3592 );
and \U$3479 ( \3594 , \3590 , \3593 );
and \U$3480 ( \3595 , \3359 , \3589 );
or \U$3481 ( \3596 , \3594 , \3595 );
buf \U$3482 ( \3597 , \3596 );
buf \U$3483 ( \3598 , \3597 );
xor \U$3484 ( \3599 , \3238 , \3598 );
xor \U$3485 ( \3600 , \1873 , \2114 );
xor \U$3486 ( \3601 , \3600 , \2306 );
buf \U$3487 ( \3602 , \3601 );
buf \U$3488 ( \3603 , \3602 );
and \U$3489 ( \3604 , \3599 , \3603 );
and \U$3490 ( \3605 , \3238 , \3598 );
or \U$3491 ( \3606 , \3604 , \3605 );
buf \U$3492 ( \3607 , \3606 );
buf \U$3493 ( \3608 , \3607 );
xor \U$3494 ( \3609 , \2311 , \2678 );
xor \U$3495 ( \3610 , \3609 , \2710 );
buf \U$3496 ( \3611 , \3610 );
buf \U$3497 ( \3612 , \3611 );
xor \U$3498 ( \3613 , \3608 , \3612 );
xor \U$3499 ( \3614 , \2659 , \2662 );
xor \U$3500 ( \3615 , \3614 , \2667 );
buf \U$3501 ( \3616 , \3615 );
buf \U$3502 ( \3617 , \3616 );
buf \U$3503 ( \3618 , RIc0d7d08_15);
buf \U$3504 ( \3619 , RIc0d9ec8_87);
xor \U$3505 ( \3620 , \3618 , \3619 );
buf \U$3506 ( \3621 , \3620 );
buf \U$3507 ( \3622 , \3621 );
not \U$3508 ( \3623 , \3622 );
buf \U$3509 ( \3624 , \809 );
not \U$3510 ( \3625 , \3624 );
or \U$3511 ( \3626 , \3623 , \3625 );
buf \U$3512 ( \3627 , \3187 );
not \U$3513 ( \3628 , \3627 );
buf \U$3514 ( \3629 , \634 );
not \U$3515 ( \3630 , \3629 );
buf \U$3516 ( \3631 , \3630 );
buf \U$3517 ( \3632 , \3631 );
nand \U$3518 ( \3633 , \3628 , \3632 );
buf \U$3519 ( \3634 , \3633 );
buf \U$3520 ( \3635 , \3634 );
nand \U$3521 ( \3636 , \3626 , \3635 );
buf \U$3522 ( \3637 , \3636 );
buf \U$3523 ( \3638 , \3637 );
not \U$3524 ( \3639 , \3638 );
xor \U$3525 ( \3640 , \2453 , \2454 );
buf \U$3526 ( \3641 , \3640 );
buf \U$3527 ( \3642 , \3641 );
not \U$3528 ( \3643 , \3642 );
buf \U$3529 ( \3644 , \1225 );
not \U$3530 ( \3645 , \3644 );
or \U$3531 ( \3646 , \3643 , \3645 );
buf \U$3532 ( \3647 , \1705 );
buf \U$3533 ( \3648 , \1795 );
nand \U$3534 ( \3649 , \3647 , \3648 );
buf \U$3535 ( \3650 , \3649 );
buf \U$3536 ( \3651 , \3650 );
nand \U$3537 ( \3652 , \3646 , \3651 );
buf \U$3538 ( \3653 , \3652 );
buf \U$3539 ( \3654 , \3653 );
not \U$3540 ( \3655 , \3654 );
or \U$3541 ( \3656 , \3639 , \3655 );
buf \U$3542 ( \3657 , \3637 );
buf \U$3543 ( \3658 , \3653 );
or \U$3544 ( \3659 , \3657 , \3658 );
buf \U$3545 ( \3660 , RIc0d8410_30);
buf \U$3546 ( \3661 , RIc0d9748_71);
xor \U$3547 ( \3662 , \3660 , \3661 );
buf \U$3548 ( \3663 , \3662 );
buf \U$3549 ( \3664 , \3663 );
not \U$3550 ( \3665 , \3664 );
buf \U$3551 ( \3666 , \2269 );
not \U$3552 ( \3667 , \3666 );
or \U$3553 ( \3668 , \3665 , \3667 );
buf \U$3554 ( \3669 , \1884 );
not \U$3555 ( \3670 , \3669 );
buf \U$3556 ( \3671 , \1282 );
nand \U$3557 ( \3672 , \3670 , \3671 );
buf \U$3558 ( \3673 , \3672 );
buf \U$3559 ( \3674 , \3673 );
nand \U$3560 ( \3675 , \3668 , \3674 );
buf \U$3561 ( \3676 , \3675 );
buf \U$3562 ( \3677 , \3676 );
nand \U$3563 ( \3678 , \3659 , \3677 );
buf \U$3564 ( \3679 , \3678 );
buf \U$3565 ( \3680 , \3679 );
nand \U$3566 ( \3681 , \3656 , \3680 );
buf \U$3567 ( \3682 , \3681 );
buf \U$3568 ( \3683 , \3682 );
xor \U$3569 ( \3684 , \2457 , \2484 );
xor \U$3570 ( \3685 , \3684 , \2499 );
buf \U$3571 ( \3686 , \3685 );
buf \U$3572 ( \3687 , \3686 );
xor \U$3573 ( \3688 , \3683 , \3687 );
buf \U$3574 ( \3689 , RIc0d7fd8_21);
buf \U$3575 ( \3690 , RIc0d9bf8_81);
xor \U$3576 ( \3691 , \3689 , \3690 );
buf \U$3577 ( \3692 , \3691 );
buf \U$3578 ( \3693 , \3692 );
not \U$3579 ( \3694 , \3693 );
buf \U$3580 ( \3695 , \2766 );
not \U$3581 ( \3696 , \3695 );
or \U$3582 ( \3697 , \3694 , \3696 );
buf \U$3583 ( \3698 , \3571 );
not \U$3584 ( \3699 , \3698 );
buf \U$3585 ( \3700 , \1078 );
nand \U$3586 ( \3701 , \3699 , \3700 );
buf \U$3587 ( \3702 , \3701 );
buf \U$3588 ( \3703 , \3702 );
nand \U$3589 ( \3704 , \3697 , \3703 );
buf \U$3590 ( \3705 , \3704 );
buf \U$3591 ( \3706 , \3705 );
not \U$3592 ( \3707 , \3706 );
buf \U$3593 ( \3708 , RIc0d7948_7);
buf \U$3594 ( \3709 , RIc0da288_95);
xor \U$3595 ( \3710 , \3708 , \3709 );
buf \U$3596 ( \3711 , \3710 );
buf \U$3597 ( \3712 , \3711 );
not \U$3598 ( \3713 , \3712 );
buf \U$3601 ( \3714 , \329 );
buf \U$3602 ( \3715 , \3714 );
not \U$3603 ( \3716 , \3715 );
or \U$3604 ( \3717 , \3713 , \3716 );
buf \U$3605 ( \3718 , \344 );
buf \U$3606 ( \3719 , \3549 );
nand \U$3607 ( \3720 , \3718 , \3719 );
buf \U$3608 ( \3721 , \3720 );
buf \U$3609 ( \3722 , \3721 );
nand \U$3610 ( \3723 , \3717 , \3722 );
buf \U$3611 ( \3724 , \3723 );
buf \U$3612 ( \3725 , \3724 );
not \U$3613 ( \3726 , \3725 );
or \U$3614 ( \3727 , \3707 , \3726 );
buf \U$3615 ( \3728 , \3724 );
buf \U$3616 ( \3729 , \3705 );
or \U$3617 ( \3730 , \3728 , \3729 );
buf \U$3618 ( \3731 , RIc0d81b8_25);
buf \U$3619 ( \3732 , RIc0d9a18_77);
xor \U$3620 ( \3733 , \3731 , \3732 );
buf \U$3621 ( \3734 , \3733 );
buf \U$3622 ( \3735 , \3734 );
not \U$3623 ( \3736 , \3735 );
buf \U$3624 ( \3737 , \1183 );
not \U$3625 ( \3738 , \3737 );
or \U$3626 ( \3739 , \3736 , \3738 );
buf \U$3627 ( \3740 , \1585 );
not \U$3628 ( \3741 , \3740 );
buf \U$3629 ( \3742 , \3741 );
buf \U$3630 ( \3743 , \3742 );
buf \U$3631 ( \3744 , \3464 );
nand \U$3632 ( \3745 , \3743 , \3744 );
buf \U$3633 ( \3746 , \3745 );
buf \U$3634 ( \3747 , \3746 );
nand \U$3635 ( \3748 , \3739 , \3747 );
buf \U$3636 ( \3749 , \3748 );
buf \U$3637 ( \3750 , \3749 );
nand \U$3638 ( \3751 , \3730 , \3750 );
buf \U$3639 ( \3752 , \3751 );
buf \U$3640 ( \3753 , \3752 );
nand \U$3641 ( \3754 , \3727 , \3753 );
buf \U$3642 ( \3755 , \3754 );
buf \U$3643 ( \3756 , \3755 );
buf \U$3644 ( \3757 , RIc0d7b28_11);
buf \U$3645 ( \3758 , RIc0da0a8_91);
xor \U$3646 ( \3759 , \3757 , \3758 );
buf \U$3647 ( \3760 , \3759 );
buf \U$3648 ( \3761 , \3760 );
not \U$3649 ( \3762 , \3761 );
buf \U$3650 ( \3763 , \2726 );
not \U$3651 ( \3764 , \3763 );
or \U$3652 ( \3765 , \3762 , \3764 );
buf \U$3653 ( \3766 , \3267 );
not \U$3654 ( \3767 , \3766 );
buf \U$3655 ( \3768 , \1933 );
nand \U$3656 ( \3769 , \3767 , \3768 );
buf \U$3657 ( \3770 , \3769 );
buf \U$3658 ( \3771 , \3770 );
nand \U$3659 ( \3772 , \3765 , \3771 );
buf \U$3660 ( \3773 , \3772 );
xor \U$3661 ( \3774 , \3240 , \3241 );
buf \U$3662 ( \3775 , \3774 );
buf \U$3663 ( \3776 , \3775 );
not \U$3664 ( \3777 , \3776 );
buf \U$3665 ( \3778 , \1221 );
not \U$3666 ( \3779 , \3778 );
buf \U$3667 ( \3780 , \3779 );
buf \U$3670 ( \3781 , \3780 );
buf \U$3671 ( \3782 , \3781 );
not \U$3672 ( \3783 , \3782 );
or \U$3673 ( \3784 , \3777 , \3783 );
buf \U$3674 ( \3785 , \1229 );
buf \U$3675 ( \3786 , \3641 );
nand \U$3676 ( \3787 , \3785 , \3786 );
buf \U$3677 ( \3788 , \3787 );
buf \U$3678 ( \3789 , \3788 );
nand \U$3679 ( \3790 , \3784 , \3789 );
buf \U$3680 ( \3791 , \3790 );
xor \U$3681 ( \3792 , \3773 , \3791 );
buf \U$3682 ( \3793 , RIc0d8668_35);
buf \U$3683 ( \3794 , RIc0d9568_67);
xor \U$3684 ( \3795 , \3793 , \3794 );
buf \U$3685 ( \3796 , \3795 );
buf \U$3686 ( \3797 , \3796 );
not \U$3687 ( \3798 , \3797 );
buf \U$3688 ( \3799 , \1823 );
not \U$3689 ( \3800 , \3799 );
or \U$3690 ( \3801 , \3798 , \3800 );
buf \U$3691 ( \3802 , \686 );
buf \U$3692 ( \3803 , \3248 );
nand \U$3693 ( \3804 , \3802 , \3803 );
buf \U$3694 ( \3805 , \3804 );
buf \U$3695 ( \3806 , \3805 );
nand \U$3696 ( \3807 , \3801 , \3806 );
buf \U$3697 ( \3808 , \3807 );
and \U$3698 ( \3809 , \3792 , \3808 );
and \U$3699 ( \3810 , \3773 , \3791 );
or \U$3700 ( \3811 , \3809 , \3810 );
buf \U$3701 ( \3812 , \3811 );
xor \U$3702 ( \3813 , \3756 , \3812 );
buf \U$3703 ( \3814 , \2124 );
not \U$3704 ( \3815 , \3814 );
buf \U$3705 ( \3816 , \3815 );
buf \U$3706 ( \3817 , \3816 );
buf \U$3707 ( \3818 , RIc0d9928_75);
buf \U$3708 ( \3819 , RIc0d82a8_27);
xnor \U$3709 ( \3820 , \3818 , \3819 );
buf \U$3710 ( \3821 , \3820 );
buf \U$3711 ( \3822 , \3821 );
or \U$3712 ( \3823 , \3817 , \3822 );
buf \U$3713 ( \3824 , \1370 );
buf \U$3714 ( \3825 , \3442 );
or \U$3715 ( \3826 , \3824 , \3825 );
nand \U$3716 ( \3827 , \3823 , \3826 );
buf \U$3717 ( \3828 , \3827 );
buf \U$3718 ( \3829 , \3828 );
buf \U$3719 ( \3830 , RIc0da468_99);
buf \U$3720 ( \3831 , \304 );
and \U$3721 ( \3832 , \3830 , \3831 );
not \U$3722 ( \3833 , \3830 );
buf \U$3723 ( \3834 , RIc0d7768_3);
and \U$3724 ( \3835 , \3833 , \3834 );
nor \U$3725 ( \3836 , \3832 , \3835 );
buf \U$3726 ( \3837 , \3836 );
buf \U$3727 ( \3838 , \3837 );
not \U$3728 ( \3839 , \3838 );
buf \U$3729 ( \3840 , \3839 );
buf \U$3730 ( \3841 , \3840 );
not \U$3731 ( \3842 , \3841 );
buf \U$3732 ( \3843 , \2470 );
not \U$3733 ( \3844 , \3843 );
or \U$3734 ( \3845 , \3842 , \3844 );
buf \U$3735 ( \3846 , \2476 );
buf \U$3736 ( \3847 , \3490 );
nand \U$3737 ( \3848 , \3846 , \3847 );
buf \U$3738 ( \3849 , \3848 );
buf \U$3739 ( \3850 , \3849 );
nand \U$3740 ( \3851 , \3845 , \3850 );
buf \U$3741 ( \3852 , \3851 );
buf \U$3742 ( \3853 , \3852 );
or \U$3743 ( \3854 , \3829 , \3853 );
buf \U$3744 ( \3855 , \3312 );
not \U$3745 ( \3856 , \3855 );
buf \U$3746 ( \3857 , \2070 );
not \U$3747 ( \3858 , \3857 );
or \U$3748 ( \3859 , \3856 , \3858 );
buf \U$3749 ( \3860 , RIc0d7858_5);
buf \U$3750 ( \3861 , RIc0da378_97);
xnor \U$3751 ( \3862 , \3860 , \3861 );
buf \U$3752 ( \3863 , \3862 );
buf \U$3753 ( \3864 , \3863 );
not \U$3754 ( \3865 , \3864 );
buf \U$3755 ( \3866 , \2066 );
nand \U$3756 ( \3867 , \3865 , \3866 );
buf \U$3757 ( \3868 , \3867 );
buf \U$3758 ( \3869 , \3868 );
nand \U$3759 ( \3870 , \3859 , \3869 );
buf \U$3760 ( \3871 , \3870 );
buf \U$3761 ( \3872 , \3871 );
nand \U$3762 ( \3873 , \3854 , \3872 );
buf \U$3763 ( \3874 , \3873 );
buf \U$3764 ( \3875 , \3874 );
buf \U$3765 ( \3876 , \3828 );
buf \U$3766 ( \3877 , \3852 );
nand \U$3767 ( \3878 , \3876 , \3877 );
buf \U$3768 ( \3879 , \3878 );
buf \U$3769 ( \3880 , \3879 );
nand \U$3770 ( \3881 , \3875 , \3880 );
buf \U$3771 ( \3882 , \3881 );
buf \U$3772 ( \3883 , \3882 );
and \U$3773 ( \3884 , \3813 , \3883 );
and \U$3774 ( \3885 , \3756 , \3812 );
or \U$3775 ( \3886 , \3884 , \3885 );
buf \U$3776 ( \3887 , \3886 );
buf \U$3777 ( \3888 , \3887 );
and \U$3778 ( \3889 , \3688 , \3888 );
and \U$3779 ( \3890 , \3683 , \3687 );
or \U$3780 ( \3891 , \3889 , \3890 );
buf \U$3781 ( \3892 , \3891 );
buf \U$3782 ( \3893 , \3892 );
xor \U$3783 ( \3894 , \3617 , \3893 );
xor \U$3784 ( \3895 , \3066 , \3080 );
xor \U$3785 ( \3896 , \3895 , \3085 );
buf \U$3786 ( \3897 , \3896 );
buf \U$3787 ( \3898 , \3897 );
and \U$3788 ( \3899 , \3894 , \3898 );
and \U$3789 ( \3900 , \3617 , \3893 );
or \U$3790 ( \3901 , \3899 , \3900 );
buf \U$3791 ( \3902 , \3901 );
buf \U$3792 ( \3903 , \3902 );
buf \U$3793 ( \3904 , \2644 );
not \U$3794 ( \3905 , \3904 );
buf \U$3795 ( \3906 , \2671 );
not \U$3796 ( \3907 , \3906 );
or \U$3797 ( \3908 , \3905 , \3907 );
buf \U$3798 ( \3909 , \2644 );
buf \U$3799 ( \3910 , \2671 );
or \U$3800 ( \3911 , \3909 , \3910 );
nand \U$3801 ( \3912 , \3908 , \3911 );
buf \U$3802 ( \3913 , \3912 );
buf \U$3803 ( \3914 , \3913 );
buf \U$3804 ( \3915 , \2516 );
and \U$3805 ( \3916 , \3914 , \3915 );
not \U$3806 ( \3917 , \3914 );
buf \U$3807 ( \3918 , \2513 );
and \U$3808 ( \3919 , \3917 , \3918 );
nor \U$3809 ( \3920 , \3916 , \3919 );
buf \U$3810 ( \3921 , \3920 );
buf \U$3811 ( \3922 , \3921 );
xor \U$3812 ( \3923 , \3903 , \3922 );
buf \U$3813 ( \3924 , \3057 );
buf \U$3814 ( \3925 , \3034 );
xor \U$3815 ( \3926 , \3924 , \3925 );
buf \U$3816 ( \3927 , \3926 );
buf \U$3817 ( \3928 , \3927 );
buf \U$3818 ( \3929 , \3089 );
xor \U$3819 ( \3930 , \3928 , \3929 );
buf \U$3820 ( \3931 , \3930 );
buf \U$3821 ( \3932 , \3931 );
and \U$3822 ( \3933 , \3923 , \3932 );
and \U$3823 ( \3934 , \3903 , \3922 );
or \U$3824 ( \3935 , \3933 , \3934 );
buf \U$3825 ( \3936 , \3935 );
buf \U$3826 ( \3937 , \3936 );
and \U$3827 ( \3938 , \3613 , \3937 );
and \U$3828 ( \3939 , \3608 , \3612 );
or \U$3829 ( \3940 , \3938 , \3939 );
buf \U$3830 ( \3941 , \3940 );
buf \U$3831 ( \3942 , \3941 );
xor \U$3832 ( \3943 , \3110 , \3942 );
buf \U$3833 ( \3944 , \3943 );
buf \U$3834 ( \3945 , \3944 );
xor \U$3835 ( \3946 , \3031 , \3096 );
xor \U$3836 ( \3947 , \3946 , \3101 );
buf \U$3837 ( \3948 , \3947 );
buf \U$3838 ( \3949 , \3948 );
buf \U$3839 ( \3950 , RIc0d9fb8_89);
buf \U$3840 ( \3951 , RIc0d7c18_13);
and \U$3841 ( \3952 , \3950 , \3951 );
not \U$3842 ( \3953 , \3950 );
buf \U$3843 ( \3954 , \1001 );
and \U$3844 ( \3955 , \3953 , \3954 );
nor \U$3845 ( \3956 , \3952 , \3955 );
buf \U$3846 ( \3957 , \3956 );
buf \U$3847 ( \3958 , \3957 );
not \U$3848 ( \3959 , \3958 );
buf \U$3849 ( \3960 , \842 );
not \U$3850 ( \3961 , \3960 );
or \U$3851 ( \3962 , \3959 , \3961 );
buf \U$3852 ( \3963 , \3393 );
not \U$3853 ( \3964 , \3963 );
buf \U$3854 ( \3965 , \846 );
nand \U$3855 ( \3966 , \3964 , \3965 );
buf \U$3856 ( \3967 , \3966 );
buf \U$3857 ( \3968 , \3967 );
nand \U$3858 ( \3969 , \3962 , \3968 );
buf \U$3859 ( \3970 , \3969 );
buf \U$3860 ( \3971 , \3970 );
not \U$3861 ( \3972 , \3971 );
buf \U$3862 ( \3973 , \3972 );
buf \U$3863 ( \3974 , \3973 );
not \U$3864 ( \3975 , \3974 );
buf \U$3865 ( \3976 , RIc0d80c8_23);
buf \U$3866 ( \3977 , RIc0d9b08_79);
xor \U$3867 ( \3978 , \3976 , \3977 );
buf \U$3868 ( \3979 , \3978 );
buf \U$3869 ( \3980 , \3979 );
not \U$3870 ( \3981 , \3980 );
buf \U$3871 ( \3982 , \397 );
not \U$3872 ( \3983 , \3982 );
or \U$3873 ( \3984 , \3981 , \3983 );
buf \U$3874 ( \3985 , \401 );
buf \U$3875 ( \3986 , \3985 );
buf \U$3876 ( \3987 , \3363 );
nand \U$3877 ( \3988 , \3986 , \3987 );
buf \U$3878 ( \3989 , \3988 );
buf \U$3879 ( \3990 , \3989 );
nand \U$3880 ( \3991 , \3984 , \3990 );
buf \U$3881 ( \3992 , \3991 );
buf \U$3882 ( \3993 , \3992 );
not \U$3883 ( \3994 , \3993 );
buf \U$3884 ( \3995 , \3994 );
buf \U$3885 ( \3996 , \3995 );
not \U$3886 ( \3997 , \3996 );
or \U$3887 ( \3998 , \3975 , \3997 );
buf \U$3888 ( \3999 , RIc0d7a38_9);
buf \U$3889 ( \4000 , RIc0da198_93);
xor \U$3890 ( \4001 , \3999 , \4000 );
buf \U$3891 ( \4002 , \4001 );
buf \U$3892 ( \4003 , \4002 );
not \U$3893 ( \4004 , \4003 );
buf \U$3894 ( \4005 , \3415 );
not \U$3895 ( \4006 , \4005 );
or \U$3896 ( \4007 , \4004 , \4006 );
buf \U$3899 ( \4008 , \480 );
buf \U$3900 ( \4009 , \4008 );
buf \U$3901 ( \4010 , \3410 );
nand \U$3902 ( \4011 , \4009 , \4010 );
buf \U$3903 ( \4012 , \4011 );
buf \U$3904 ( \4013 , \4012 );
nand \U$3905 ( \4014 , \4007 , \4013 );
buf \U$3906 ( \4015 , \4014 );
buf \U$3907 ( \4016 , \4015 );
nand \U$3908 ( \4017 , \3998 , \4016 );
buf \U$3909 ( \4018 , \4017 );
buf \U$3910 ( \4019 , \4018 );
buf \U$3911 ( \4020 , \3992 );
buf \U$3912 ( \4021 , \3970 );
nand \U$3913 ( \4022 , \4020 , \4021 );
buf \U$3914 ( \4023 , \4022 );
buf \U$3915 ( \4024 , \4023 );
nand \U$3916 ( \4025 , \4019 , \4024 );
buf \U$3917 ( \4026 , \4025 );
buf \U$3918 ( \4027 , RIc0d9478_65);
buf \U$3919 ( \4028 , RIc0d87d0_38);
and \U$3920 ( \4029 , \4027 , \4028 );
buf \U$3921 ( \4030 , \4029 );
buf \U$3922 ( \4031 , \4030 );
buf \U$3923 ( \4032 , RIc0da558_101);
buf \U$3924 ( \4033 , RIc0d7678_1);
and \U$3925 ( \4034 , \4032 , \4033 );
not \U$3926 ( \4035 , \4032 );
buf \U$3927 ( \4036 , \974 );
and \U$3928 ( \4037 , \4035 , \4036 );
nor \U$3929 ( \4038 , \4034 , \4037 );
buf \U$3930 ( \4039 , \4038 );
buf \U$3931 ( \4040 , \4039 );
not \U$3932 ( \4041 , \4040 );
buf \U$3935 ( \4042 , \3528 );
buf \U$3938 ( \4043 , \4042 );
buf \U$3939 ( \4044 , \4043 );
not \U$3940 ( \4045 , \4044 );
or \U$3941 ( \4046 , \4041 , \4045 );
buf \U$3942 ( \4047 , \3518 );
not \U$3943 ( \4048 , \4047 );
buf \U$3944 ( \4049 , \4048 );
buf \U$3945 ( \4050 , \4049 );
buf \U$3946 ( \4051 , RIc0da558_101);
nand \U$3947 ( \4052 , \4050 , \4051 );
buf \U$3948 ( \4053 , \4052 );
buf \U$3949 ( \4054 , \4053 );
nand \U$3950 ( \4055 , \4046 , \4054 );
buf \U$3951 ( \4056 , \4055 );
buf \U$3952 ( \4057 , \4056 );
xor \U$3953 ( \4058 , \4031 , \4057 );
buf \U$3954 ( \4059 , \1739 );
buf \U$3955 ( \4060 , RIc0d9ce8_83);
buf \U$3956 ( \4061 , RIc0d7ee8_19);
xnor \U$3957 ( \4062 , \4060 , \4061 );
buf \U$3958 ( \4063 , \4062 );
buf \U$3959 ( \4064 , \4063 );
or \U$3960 ( \4065 , \4059 , \4064 );
buf \U$3961 ( \4066 , \996 );
buf \U$3962 ( \4067 , \3334 );
not \U$3963 ( \4068 , \4067 );
buf \U$3964 ( \4069 , \4068 );
buf \U$3965 ( \4070 , \4069 );
or \U$3966 ( \4071 , \4066 , \4070 );
nand \U$3967 ( \4072 , \4065 , \4071 );
buf \U$3968 ( \4073 , \4072 );
buf \U$3969 ( \4074 , \4073 );
and \U$3970 ( \4075 , \4058 , \4074 );
and \U$3971 ( \4076 , \4031 , \4057 );
or \U$3972 ( \4077 , \4075 , \4076 );
buf \U$3973 ( \4078 , \4077 );
xor \U$3974 ( \4079 , \4026 , \4078 );
buf \U$3975 ( \4080 , RIc0d7df8_17);
buf \U$3976 ( \4081 , RIc0d9dd8_85);
xor \U$3977 ( \4082 , \4080 , \4081 );
buf \U$3978 ( \4083 , \4082 );
buf \U$3979 ( \4084 , \4083 );
not \U$3980 ( \4085 , \4084 );
buf \U$3981 ( \4086 , \1389 );
not \U$3982 ( \4087 , \4086 );
or \U$3983 ( \4088 , \4085 , \4087 );
buf \U$3984 ( \4089 , \3288 );
not \U$3985 ( \4090 , \4089 );
buf \U$3986 ( \4091 , \2960 );
nand \U$3987 ( \4092 , \4090 , \4091 );
buf \U$3988 ( \4093 , \4092 );
buf \U$3989 ( \4094 , \4093 );
nand \U$3990 ( \4095 , \4088 , \4094 );
buf \U$3991 ( \4096 , \4095 );
not \U$3992 ( \4097 , \4096 );
buf \U$3993 ( \4098 , RIc0d8488_31);
buf \U$3994 ( \4099 , RIc0d9748_71);
xor \U$3995 ( \4100 , \4098 , \4099 );
buf \U$3996 ( \4101 , \4100 );
buf \U$3997 ( \4102 , \4101 );
not \U$3998 ( \4103 , \4102 );
buf \U$3999 ( \4104 , \2269 );
not \U$4000 ( \4105 , \4104 );
or \U$4001 ( \4106 , \4103 , \4105 );
buf \U$4002 ( \4107 , \2927 );
buf \U$4003 ( \4108 , \3663 );
nand \U$4004 ( \4109 , \4107 , \4108 );
buf \U$4005 ( \4110 , \4109 );
buf \U$4006 ( \4111 , \4110 );
nand \U$4007 ( \4112 , \4106 , \4111 );
buf \U$4008 ( \4113 , \4112 );
buf \U$4009 ( \4114 , \4113 );
not \U$4010 ( \4115 , \4114 );
buf \U$4011 ( \4116 , \4115 );
nand \U$4012 ( \4117 , \4097 , \4116 );
not \U$4013 ( \4118 , \4117 );
buf \U$4014 ( \4119 , \773 );
buf \U$4015 ( \4120 , RIc0d8398_29);
buf \U$4016 ( \4121 , RIc0d9838_73);
xnor \U$4017 ( \4122 , \4120 , \4121 );
buf \U$4018 ( \4123 , \4122 );
buf \U$4019 ( \4124 , \4123 );
or \U$4020 ( \4125 , \4119 , \4124 );
buf \U$4021 ( \4126 , \2879 );
buf \U$4022 ( \4127 , \3164 );
not \U$4023 ( \4128 , \4127 );
buf \U$4024 ( \4129 , \4128 );
buf \U$4025 ( \4130 , \4129 );
or \U$4026 ( \4131 , \4126 , \4130 );
nand \U$4027 ( \4132 , \4125 , \4131 );
buf \U$4028 ( \4133 , \4132 );
not \U$4029 ( \4134 , \4133 );
or \U$4030 ( \4135 , \4118 , \4134 );
buf \U$4031 ( \4136 , \4096 );
buf \U$4032 ( \4137 , \4113 );
nand \U$4033 ( \4138 , \4136 , \4137 );
buf \U$4034 ( \4139 , \4138 );
nand \U$4035 ( \4140 , \4135 , \4139 );
and \U$4036 ( \4141 , \4079 , \4140 );
and \U$4037 ( \4142 , \4026 , \4078 );
or \U$4038 ( \4143 , \4141 , \4142 );
buf \U$4039 ( \4144 , \4143 );
xor \U$4040 ( \4145 , \3239 , \3283 );
xor \U$4041 ( \4146 , \4145 , \3354 );
buf \U$4042 ( \4147 , \4146 );
buf \U$4043 ( \4148 , \4147 );
xor \U$4044 ( \4149 , \4144 , \4148 );
xor \U$4045 ( \4150 , \3438 , \3509 );
xor \U$4046 ( \4151 , \4150 , \3584 );
buf \U$4047 ( \4152 , \4151 );
buf \U$4048 ( \4153 , \4152 );
and \U$4049 ( \4154 , \4149 , \4153 );
and \U$4050 ( \4155 , \4144 , \4148 );
or \U$4051 ( \4156 , \4154 , \4155 );
buf \U$4052 ( \4157 , \4156 );
buf \U$4053 ( \4158 , \4157 );
xor \U$4054 ( \4159 , \3359 , \3589 );
xor \U$4055 ( \4160 , \4159 , \3593 );
buf \U$4056 ( \4161 , \4160 );
buf \U$4057 ( \4162 , \4161 );
xor \U$4058 ( \4163 , \4158 , \4162 );
xor \U$4059 ( \4164 , \3226 , \3113 );
xor \U$4060 ( \4165 , \4164 , \3136 );
buf \U$4061 ( \4166 , \4165 );
and \U$4062 ( \4167 , \4163 , \4166 );
and \U$4063 ( \4168 , \4158 , \4162 );
or \U$4064 ( \4169 , \4167 , \4168 );
buf \U$4065 ( \4170 , \4169 );
buf \U$4066 ( \4171 , \4170 );
not \U$4067 ( \4172 , \4171 );
xor \U$4068 ( \4173 , \3238 , \3598 );
xor \U$4069 ( \4174 , \4173 , \3603 );
buf \U$4070 ( \4175 , \4174 );
buf \U$4071 ( \4176 , \4175 );
not \U$4072 ( \4177 , \4176 );
or \U$4073 ( \4178 , \4172 , \4177 );
buf \U$4074 ( \4179 , \4175 );
buf \U$4075 ( \4180 , \4170 );
or \U$4076 ( \4181 , \4179 , \4180 );
xor \U$4077 ( \4182 , \3244 , \3261 );
xor \U$4078 ( \4183 , \4182 , \3278 );
buf \U$4079 ( \4184 , \4183 );
buf \U$4080 ( \4185 , \4184 );
not \U$4081 ( \4186 , \4185 );
xor \U$4082 ( \4187 , \3403 , \3425 );
xor \U$4083 ( \4188 , \4187 , \3379 );
buf \U$4084 ( \4189 , \4188 );
not \U$4085 ( \4190 , \4189 );
or \U$4086 ( \4191 , \4186 , \4190 );
buf \U$4087 ( \4192 , \4184 );
buf \U$4088 ( \4193 , \4188 );
or \U$4089 ( \4194 , \4192 , \4193 );
buf \U$4090 ( \4195 , \3179 );
buf \U$4091 ( \4196 , \3158 );
and \U$4092 ( \4197 , \4195 , \4196 );
not \U$4093 ( \4198 , \4195 );
buf \U$4094 ( \4199 , \3155 );
and \U$4095 ( \4200 , \4198 , \4199 );
nor \U$4096 ( \4201 , \4197 , \4200 );
buf \U$4097 ( \4202 , \4201 );
buf \U$4098 ( \4203 , \4202 );
buf \U$4099 ( \4204 , \3194 );
xor \U$4100 ( \4205 , \4203 , \4204 );
buf \U$4101 ( \4206 , \4205 );
buf \U$4102 ( \4207 , \4206 );
nand \U$4103 ( \4208 , \4194 , \4207 );
buf \U$4104 ( \4209 , \4208 );
buf \U$4105 ( \4210 , \4209 );
nand \U$4106 ( \4211 , \4191 , \4210 );
buf \U$4107 ( \4212 , \4211 );
buf \U$4108 ( \4213 , \4212 );
xor \U$4109 ( \4214 , \3458 , \3502 );
buf \U$4110 ( \4215 , \4214 );
buf \U$4111 ( \4216 , \3476 );
not \U$4112 ( \4217 , \4216 );
buf \U$4113 ( \4218 , \4217 );
buf \U$4114 ( \4219 , \4218 );
and \U$4115 ( \4220 , \4215 , \4219 );
not \U$4116 ( \4221 , \4215 );
buf \U$4117 ( \4222 , \3476 );
and \U$4118 ( \4223 , \4221 , \4222 );
nor \U$4119 ( \4224 , \4220 , \4223 );
buf \U$4120 ( \4225 , \4224 );
buf \U$4121 ( \4226 , \4225 );
not \U$4122 ( \4227 , \4226 );
buf \U$4123 ( \4228 , \4227 );
buf \U$4124 ( \4229 , \4228 );
not \U$4125 ( \4230 , \4229 );
xor \U$4126 ( \4231 , \3324 , \3347 );
xnor \U$4127 ( \4232 , \4231 , \3302 );
buf \U$4128 ( \4233 , \4232 );
not \U$4129 ( \4234 , \4233 );
buf \U$4130 ( \4235 , \4234 );
buf \U$4131 ( \4236 , \4235 );
not \U$4132 ( \4237 , \4236 );
or \U$4133 ( \4238 , \4230 , \4237 );
buf \U$4134 ( \4239 , \4232 );
buf \U$4135 ( \4240 , \4225 );
nand \U$4136 ( \4241 , \4239 , \4240 );
buf \U$4137 ( \4242 , \4241 );
buf \U$4138 ( \4243 , \4242 );
xor \U$4139 ( \4244 , \3545 , \3562 );
xor \U$4140 ( \4245 , \4244 , \3579 );
buf \U$4141 ( \4246 , \4245 );
buf \U$4142 ( \4247 , \4246 );
nand \U$4143 ( \4248 , \4243 , \4247 );
buf \U$4144 ( \4249 , \4248 );
buf \U$4145 ( \4250 , \4249 );
nand \U$4146 ( \4251 , \4238 , \4250 );
buf \U$4147 ( \4252 , \4251 );
buf \U$4148 ( \4253 , \4252 );
xor \U$4149 ( \4254 , \4213 , \4253 );
xor \U$4150 ( \4255 , \3121 , \3130 );
xor \U$4151 ( \4256 , \4255 , \3116 );
buf \U$4152 ( \4257 , \4256 );
and \U$4153 ( \4258 , \4254 , \4257 );
and \U$4154 ( \4259 , \4213 , \4253 );
or \U$4155 ( \4260 , \4258 , \4259 );
buf \U$4156 ( \4261 , \4260 );
buf \U$4157 ( \4262 , \4261 );
xor \U$4158 ( \4263 , \3206 , \3209 );
xor \U$4159 ( \4264 , \4263 , \3222 );
buf \U$4160 ( \4265 , \4264 );
buf \U$4161 ( \4266 , \4265 );
xor \U$4162 ( \4267 , \3683 , \3687 );
xor \U$4163 ( \4268 , \4267 , \3888 );
buf \U$4164 ( \4269 , \4268 );
buf \U$4165 ( \4270 , \4269 );
xor \U$4166 ( \4271 , \4266 , \4270 );
buf \U$4167 ( \4272 , \3637 );
not \U$4168 ( \4273 , \4272 );
buf \U$4169 ( \4274 , \4273 );
buf \U$4170 ( \4275 , \4274 );
not \U$4171 ( \4276 , \4275 );
xor \U$4172 ( \4277 , \3653 , \3676 );
buf \U$4173 ( \4278 , \4277 );
not \U$4174 ( \4279 , \4278 );
or \U$4175 ( \4280 , \4276 , \4279 );
buf \U$4176 ( \4281 , \4277 );
buf \U$4177 ( \4282 , \4274 );
or \U$4178 ( \4283 , \4281 , \4282 );
nand \U$4179 ( \4284 , \4280 , \4283 );
buf \U$4180 ( \4285 , \4284 );
buf \U$4181 ( \4286 , \4285 );
buf \U$4182 ( \4287 , \4274 );
buf \U$4183 ( \4288 , \1452 );
buf \U$4184 ( \4289 , RIc0d8578_33);
buf \U$4185 ( \4290 , RIc0d9658_69);
xnor \U$4186 ( \4291 , \4289 , \4290 );
buf \U$4187 ( \4292 , \4291 );
buf \U$4188 ( \4293 , \4292 );
or \U$4189 ( \4294 , \4288 , \4293 );
buf \U$4190 ( \4295 , \284 );
not \U$4191 ( \4296 , \4295 );
buf \U$4192 ( \4297 , \4296 );
buf \U$4193 ( \4298 , \4297 );
buf \U$4194 ( \4299 , \3142 );
not \U$4195 ( \4300 , \4299 );
buf \U$4196 ( \4301 , \4300 );
buf \U$4197 ( \4302 , \4301 );
or \U$4198 ( \4303 , \4298 , \4302 );
nand \U$4199 ( \4304 , \4294 , \4303 );
buf \U$4200 ( \4305 , \4304 );
buf \U$4201 ( \4306 , \4305 );
xor \U$4202 ( \4307 , \4287 , \4306 );
buf \U$4203 ( \4308 , RIc0d8500_32);
buf \U$4204 ( \4309 , RIc0d9748_71);
xor \U$4205 ( \4310 , \4308 , \4309 );
buf \U$4206 ( \4311 , \4310 );
buf \U$4207 ( \4312 , \4311 );
not \U$4208 ( \4313 , \4312 );
buf \U$4209 ( \4314 , \2269 );
not \U$4210 ( \4315 , \4314 );
or \U$4211 ( \4316 , \4313 , \4315 );
buf \U$4212 ( \4317 , \2927 );
buf \U$4213 ( \4318 , \4101 );
nand \U$4214 ( \4319 , \4317 , \4318 );
buf \U$4215 ( \4320 , \4319 );
buf \U$4216 ( \4321 , \4320 );
nand \U$4217 ( \4322 , \4316 , \4321 );
buf \U$4218 ( \4323 , \4322 );
buf \U$4219 ( \4324 , \4323 );
not \U$4220 ( \4325 , \4324 );
xor \U$4221 ( \4326 , RIc0da378_97, RIc0d78d0_6);
buf \U$4222 ( \4327 , \4326 );
not \U$4223 ( \4328 , \4327 );
buf \U$4224 ( \4329 , \2941 );
not \U$4225 ( \4330 , \4329 );
or \U$4226 ( \4331 , \4328 , \4330 );
buf \U$4227 ( \4332 , \3863 );
not \U$4228 ( \4333 , \4332 );
buf \U$4229 ( \4334 , \734 );
nand \U$4230 ( \4335 , \4333 , \4334 );
buf \U$4231 ( \4336 , \4335 );
buf \U$4232 ( \4337 , \4336 );
nand \U$4233 ( \4338 , \4331 , \4337 );
buf \U$4234 ( \4339 , \4338 );
buf \U$4235 ( \4340 , \4339 );
not \U$4236 ( \4341 , \4340 );
or \U$4237 ( \4342 , \4325 , \4341 );
buf \U$4238 ( \4343 , \4339 );
buf \U$4239 ( \4344 , \4323 );
or \U$4240 ( \4345 , \4343 , \4344 );
buf \U$4241 ( \4346 , RIc0d7f60_20);
buf \U$4242 ( \4347 , RIc0d9ce8_83);
xnor \U$4243 ( \4348 , \4346 , \4347 );
buf \U$4244 ( \4349 , \4348 );
buf \U$4245 ( \4350 , \4349 );
not \U$4246 ( \4351 , \4350 );
buf \U$4247 ( \4352 , \4351 );
buf \U$4248 ( \4353 , \4352 );
not \U$4249 ( \4354 , \4353 );
buf \U$4250 ( \4355 , \1736 );
not \U$4251 ( \4356 , \4355 );
or \U$4252 ( \4357 , \4354 , \4356 );
buf \U$4253 ( \4358 , \4063 );
not \U$4254 ( \4359 , \4358 );
buf \U$4255 ( \4360 , \993 );
nand \U$4256 ( \4361 , \4359 , \4360 );
buf \U$4257 ( \4362 , \4361 );
buf \U$4258 ( \4363 , \4362 );
nand \U$4259 ( \4364 , \4357 , \4363 );
buf \U$4260 ( \4365 , \4364 );
buf \U$4261 ( \4366 , \4365 );
nand \U$4262 ( \4367 , \4345 , \4366 );
buf \U$4263 ( \4368 , \4367 );
buf \U$4264 ( \4369 , \4368 );
nand \U$4265 ( \4370 , \4342 , \4369 );
buf \U$4266 ( \4371 , \4370 );
buf \U$4267 ( \4372 , \4371 );
and \U$4268 ( \4373 , \4307 , \4372 );
and \U$4269 ( \4374 , \4287 , \4306 );
or \U$4270 ( \4375 , \4373 , \4374 );
buf \U$4271 ( \4376 , \4375 );
buf \U$4272 ( \4377 , \4376 );
xor \U$4273 ( \4378 , \4286 , \4377 );
buf \U$4274 ( \4379 , RIc0d9478_65);
buf \U$4275 ( \4380 , RIc0d8848_39);
and \U$4276 ( \4381 , \4379 , \4380 );
buf \U$4277 ( \4382 , \4381 );
buf \U$4278 ( \4383 , \4382 );
buf \U$4279 ( \4384 , RIc0d86e0_36);
buf \U$4280 ( \4385 , RIc0d9568_67);
xor \U$4281 ( \4386 , \4384 , \4385 );
buf \U$4282 ( \4387 , \4386 );
buf \U$4283 ( \4388 , \4387 );
not \U$4284 ( \4389 , \4388 );
buf \U$4285 ( \4390 , \678 );
not \U$4286 ( \4391 , \4390 );
or \U$4287 ( \4392 , \4389 , \4391 );
buf \U$4288 ( \4393 , \686 );
buf \U$4289 ( \4394 , \3796 );
nand \U$4290 ( \4395 , \4393 , \4394 );
buf \U$4291 ( \4396 , \4395 );
buf \U$4292 ( \4397 , \4396 );
nand \U$4293 ( \4398 , \4392 , \4397 );
buf \U$4294 ( \4399 , \4398 );
buf \U$4295 ( \4400 , \4399 );
xor \U$4296 ( \4401 , \4383 , \4400 );
buf \U$4297 ( \4402 , \521 );
buf \U$4298 ( \4403 , RIc0d7ba0_12);
buf \U$4299 ( \4404 , RIc0da0a8_91);
xnor \U$4300 ( \4405 , \4403 , \4404 );
buf \U$4301 ( \4406 , \4405 );
buf \U$4302 ( \4407 , \4406 );
or \U$4303 ( \4408 , \4402 , \4407 );
buf \U$4304 ( \4409 , \711 );
buf \U$4305 ( \4410 , \3760 );
not \U$4306 ( \4411 , \4410 );
buf \U$4307 ( \4412 , \4411 );
buf \U$4308 ( \4413 , \4412 );
or \U$4309 ( \4414 , \4409 , \4413 );
nand \U$4310 ( \4415 , \4408 , \4414 );
buf \U$4311 ( \4416 , \4415 );
buf \U$4312 ( \4417 , \4416 );
and \U$4313 ( \4418 , \4401 , \4417 );
and \U$4314 ( \4419 , \4383 , \4400 );
or \U$4315 ( \4420 , \4418 , \4419 );
buf \U$4316 ( \4421 , \4420 );
buf \U$4317 ( \4422 , \4421 );
buf \U$4318 ( \4423 , \3775 );
not \U$4319 ( \4424 , \4423 );
buf \U$4320 ( \4425 , \1232 );
not \U$4321 ( \4426 , \4425 );
buf \U$4322 ( \4427 , \4426 );
buf \U$4323 ( \4428 , \4427 );
not \U$4324 ( \4429 , \4428 );
or \U$4325 ( \4430 , \4424 , \4429 );
buf \U$4326 ( \4431 , \1225 );
xor \U$4327 ( \4432 , \4027 , \4028 );
buf \U$4328 ( \4433 , \4432 );
buf \U$4329 ( \4434 , \4433 );
nand \U$4330 ( \4435 , \4431 , \4434 );
buf \U$4331 ( \4436 , \4435 );
buf \U$4332 ( \4437 , \4436 );
nand \U$4333 ( \4438 , \4430 , \4437 );
buf \U$4334 ( \4439 , \4438 );
buf \U$4335 ( \4440 , \4439 );
not \U$4336 ( \4441 , \4440 );
buf \U$4337 ( \4442 , RIc0da288_95);
buf \U$4338 ( \4443 , RIc0d79c0_8);
and \U$4339 ( \4444 , \4442 , \4443 );
not \U$4340 ( \4445 , \4442 );
buf \U$4341 ( \4446 , RIc0d79c0_8);
not \U$4342 ( \4447 , \4446 );
buf \U$4343 ( \4448 , \4447 );
buf \U$4344 ( \4449 , \4448 );
and \U$4345 ( \4450 , \4445 , \4449 );
nor \U$4346 ( \4451 , \4444 , \4450 );
buf \U$4347 ( \4452 , \4451 );
buf \U$4348 ( \4453 , \4452 );
not \U$4349 ( \4454 , \4453 );
buf \U$4350 ( \4455 , \336 );
not \U$4351 ( \4456 , \4455 );
or \U$4352 ( \4457 , \4454 , \4456 );
buf \U$4353 ( \4458 , \343 );
buf \U$4354 ( \4459 , \3711 );
nand \U$4355 ( \4460 , \4458 , \4459 );
buf \U$4356 ( \4461 , \4460 );
buf \U$4357 ( \4462 , \4461 );
nand \U$4358 ( \4463 , \4457 , \4462 );
buf \U$4359 ( \4464 , \4463 );
buf \U$4360 ( \4465 , \4464 );
not \U$4361 ( \4466 , \4465 );
or \U$4362 ( \4467 , \4441 , \4466 );
buf \U$4363 ( \4468 , \4464 );
buf \U$4364 ( \4469 , \4439 );
or \U$4365 ( \4470 , \4468 , \4469 );
buf \U$4366 ( \4471 , RIc0da6c0_104);
buf \U$4367 ( \4472 , RIc0da738_105);
xnor \U$4368 ( \4473 , \4471 , \4472 );
buf \U$4369 ( \4474 , \4473 );
buf \U$4372 ( \4475 , \4474 );
buf \U$4373 ( \4476 , \4475 );
not \U$4374 ( \4477 , \4476 );
buf \U$4375 ( \4478 , \4474 );
xor \U$4376 ( \4479 , RIc0da6c0_104, RIc0da648_103);
buf \U$4377 ( \4480 , \4479 );
nand \U$4378 ( \4481 , \4478 , \4480 );
buf \U$4379 ( \4482 , \4481 );
buf \U$4382 ( \4483 , \4482 );
buf \U$4383 ( \4484 , \4483 );
not \U$4384 ( \4485 , \4484 );
or \U$4385 ( \4486 , \4477 , \4485 );
buf \U$4386 ( \4487 , RIc0da648_103);
nand \U$4387 ( \4488 , \4486 , \4487 );
buf \U$4388 ( \4489 , \4488 );
buf \U$4389 ( \4490 , \4489 );
nand \U$4390 ( \4491 , \4470 , \4490 );
buf \U$4391 ( \4492 , \4491 );
buf \U$4392 ( \4493 , \4492 );
nand \U$4393 ( \4494 , \4467 , \4493 );
buf \U$4394 ( \4495 , \4494 );
buf \U$4395 ( \4496 , \4495 );
xor \U$4396 ( \4497 , \4422 , \4496 );
buf \U$4397 ( \4498 , RIc0d8140_24);
buf \U$4398 ( \4499 , RIc0d9b08_79);
xnor \U$4399 ( \4500 , \4498 , \4499 );
buf \U$4400 ( \4501 , \4500 );
buf \U$4401 ( \4502 , \4501 );
not \U$4402 ( \4503 , \4502 );
buf \U$4403 ( \4504 , \4503 );
buf \U$4404 ( \4505 , \4504 );
not \U$4405 ( \4506 , \4505 );
buf \U$4406 ( \4507 , \393 );
not \U$4407 ( \4508 , \4507 );
buf \U$4408 ( \4509 , \4508 );
buf \U$4409 ( \4510 , \4509 );
not \U$4410 ( \4511 , \4510 );
or \U$4411 ( \4512 , \4506 , \4511 );
buf \U$4412 ( \4513 , \1026 );
buf \U$4413 ( \4514 , \3979 );
nand \U$4414 ( \4515 , \4513 , \4514 );
buf \U$4415 ( \4516 , \4515 );
buf \U$4416 ( \4517 , \4516 );
nand \U$4417 ( \4518 , \4512 , \4517 );
buf \U$4418 ( \4519 , \4518 );
buf \U$4419 ( \4520 , \4519 );
buf \U$4420 ( \4521 , RIc0d7d80_16);
buf \U$4421 ( \4522 , RIc0d9ec8_87);
xor \U$4422 ( \4523 , \4521 , \4522 );
buf \U$4423 ( \4524 , \4523 );
buf \U$4424 ( \4525 , \4524 );
not \U$4425 ( \4526 , \4525 );
buf \U$4428 ( \4527 , \612 );
buf \U$4429 ( \4528 , \4527 );
not \U$4430 ( \4529 , \4528 );
or \U$4431 ( \4530 , \4526 , \4529 );
buf \U$4432 ( \4531 , \3631 );
buf \U$4433 ( \4532 , \3621 );
nand \U$4434 ( \4533 , \4531 , \4532 );
buf \U$4435 ( \4534 , \4533 );
buf \U$4436 ( \4535 , \4534 );
nand \U$4437 ( \4536 , \4530 , \4535 );
buf \U$4438 ( \4537 , \4536 );
buf \U$4439 ( \4538 , \4537 );
or \U$4440 ( \4539 , \4520 , \4538 );
buf \U$4441 ( \4540 , RIc0da198_93);
buf \U$4442 ( \4541 , RIc0d7ab0_10);
and \U$4443 ( \4542 , \4540 , \4541 );
not \U$4444 ( \4543 , \4540 );
buf \U$4445 ( \4544 , RIc0d7ab0_10);
not \U$4446 ( \4545 , \4544 );
buf \U$4447 ( \4546 , \4545 );
buf \U$4448 ( \4547 , \4546 );
and \U$4449 ( \4548 , \4543 , \4547 );
nor \U$4450 ( \4549 , \4542 , \4548 );
buf \U$4451 ( \4550 , \4549 );
buf \U$4452 ( \4551 , \4550 );
not \U$4453 ( \4552 , \4551 );
buf \U$4454 ( \4553 , \3415 );
not \U$4455 ( \4554 , \4553 );
or \U$4456 ( \4555 , \4552 , \4554 );
buf \U$4457 ( \4556 , \481 );
buf \U$4458 ( \4557 , \4002 );
nand \U$4459 ( \4558 , \4556 , \4557 );
buf \U$4460 ( \4559 , \4558 );
buf \U$4461 ( \4560 , \4559 );
nand \U$4462 ( \4561 , \4555 , \4560 );
buf \U$4463 ( \4562 , \4561 );
buf \U$4464 ( \4563 , \4562 );
nand \U$4465 ( \4564 , \4539 , \4563 );
buf \U$4466 ( \4565 , \4564 );
buf \U$4467 ( \4566 , \4565 );
buf \U$4468 ( \4567 , \4519 );
buf \U$4469 ( \4568 , \4537 );
nand \U$4470 ( \4569 , \4567 , \4568 );
buf \U$4471 ( \4570 , \4569 );
buf \U$4472 ( \4571 , \4570 );
nand \U$4473 ( \4572 , \4566 , \4571 );
buf \U$4474 ( \4573 , \4572 );
buf \U$4475 ( \4574 , \4573 );
and \U$4476 ( \4575 , \4497 , \4574 );
and \U$4477 ( \4576 , \4422 , \4496 );
or \U$4478 ( \4577 , \4575 , \4576 );
buf \U$4479 ( \4578 , \4577 );
buf \U$4480 ( \4579 , \4578 );
and \U$4481 ( \4580 , \4378 , \4579 );
and \U$4482 ( \4581 , \4286 , \4377 );
or \U$4483 ( \4582 , \4580 , \4581 );
buf \U$4484 ( \4583 , \4582 );
buf \U$4485 ( \4584 , \4583 );
and \U$4486 ( \4585 , \4271 , \4584 );
and \U$4487 ( \4586 , \4266 , \4270 );
or \U$4488 ( \4587 , \4585 , \4586 );
buf \U$4489 ( \4588 , \4587 );
buf \U$4490 ( \4589 , \4588 );
xor \U$4491 ( \4590 , \4262 , \4589 );
xor \U$4492 ( \4591 , \3617 , \3893 );
xor \U$4493 ( \4592 , \4591 , \3898 );
buf \U$4494 ( \4593 , \4592 );
buf \U$4495 ( \4594 , \4593 );
and \U$4496 ( \4595 , \4590 , \4594 );
and \U$4497 ( \4596 , \4262 , \4589 );
or \U$4498 ( \4597 , \4595 , \4596 );
buf \U$4499 ( \4598 , \4597 );
buf \U$4500 ( \4599 , \4598 );
nand \U$4501 ( \4600 , \4181 , \4599 );
buf \U$4502 ( \4601 , \4600 );
buf \U$4503 ( \4602 , \4601 );
nand \U$4504 ( \4603 , \4178 , \4602 );
buf \U$4505 ( \4604 , \4603 );
buf \U$4506 ( \4605 , \4604 );
xor \U$4507 ( \4606 , \3949 , \4605 );
xor \U$4508 ( \4607 , \3608 , \3612 );
xor \U$4509 ( \4608 , \4607 , \3937 );
buf \U$4510 ( \4609 , \4608 );
buf \U$4511 ( \4610 , \4609 );
and \U$4512 ( \4611 , \4606 , \4610 );
and \U$4513 ( \4612 , \3949 , \4605 );
or \U$4514 ( \4613 , \4611 , \4612 );
buf \U$4515 ( \4614 , \4613 );
buf \U$4516 ( \4615 , \4614 );
or \U$4517 ( \4616 , \3945 , \4615 );
buf \U$4518 ( \4617 , \4616 );
buf \U$4519 ( \4618 , \4617 );
xor \U$4520 ( \4619 , \2809 , \2828 );
and \U$4521 ( \4620 , \4619 , \2844 );
and \U$4522 ( \4621 , \2809 , \2828 );
or \U$4523 ( \4622 , \4620 , \4621 );
buf \U$4524 ( \4623 , \4622 );
buf \U$4525 ( \4624 , \4623 );
buf \U$4526 ( \4625 , \1419 );
not \U$4527 ( \4626 , \4625 );
buf \U$4528 ( \4627 , \1407 );
not \U$4529 ( \4628 , \4627 );
buf \U$4530 ( \4629 , \4628 );
buf \U$4531 ( \4630 , \4629 );
not \U$4532 ( \4631 , \4630 );
or \U$4533 ( \4632 , \4626 , \4631 );
buf \U$4534 ( \4633 , \1444 );
nand \U$4535 ( \4634 , \4632 , \4633 );
buf \U$4536 ( \4635 , \4634 );
buf \U$4537 ( \4636 , \4635 );
buf \U$4538 ( \4637 , \1407 );
buf \U$4539 ( \4638 , \1422 );
nand \U$4540 ( \4639 , \4637 , \4638 );
buf \U$4541 ( \4640 , \4639 );
buf \U$4542 ( \4641 , \4640 );
nand \U$4543 ( \4642 , \4636 , \4641 );
buf \U$4544 ( \4643 , \4642 );
buf \U$4545 ( \4644 , \4643 );
buf \U$4546 ( \4645 , \1711 );
not \U$4547 ( \4646 , \4645 );
buf \U$4548 ( \4647 , \1691 );
not \U$4549 ( \4648 , \4647 );
or \U$4550 ( \4649 , \4646 , \4648 );
buf \U$4551 ( \4650 , \1691 );
buf \U$4552 ( \4651 , \1711 );
or \U$4553 ( \4652 , \4650 , \4651 );
buf \U$4554 ( \4653 , \1724 );
nand \U$4555 ( \4654 , \4652 , \4653 );
buf \U$4556 ( \4655 , \4654 );
buf \U$4557 ( \4656 , \4655 );
nand \U$4558 ( \4657 , \4649 , \4656 );
buf \U$4559 ( \4658 , \4657 );
buf \U$4560 ( \4659 , \4658 );
xor \U$4561 ( \4660 , \4644 , \4659 );
xor \U$4562 ( \4661 , \2742 , \2762 );
and \U$4563 ( \4662 , \4661 , \2785 );
and \U$4564 ( \4663 , \2742 , \2762 );
or \U$4565 ( \4664 , \4662 , \4663 );
buf \U$4566 ( \4665 , \4664 );
buf \U$4567 ( \4666 , \4665 );
xor \U$4568 ( \4667 , \4660 , \4666 );
buf \U$4569 ( \4668 , \4667 );
buf \U$4570 ( \4669 , \4668 );
xor \U$4571 ( \4670 , \4624 , \4669 );
xor \U$4572 ( \4671 , \1346 , \1363 );
and \U$4573 ( \4672 , \4671 , \1380 );
and \U$4574 ( \4673 , \1346 , \1363 );
or \U$4575 ( \4674 , \4672 , \4673 );
buf \U$4576 ( \4675 , \4674 );
buf \U$4577 ( \4676 , \4675 );
not \U$4578 ( \4677 , \1482 );
not \U$4579 ( \4678 , \1464 );
or \U$4580 ( \4679 , \4677 , \4678 );
not \U$4581 ( \4680 , \1461 );
not \U$4582 ( \4681 , \1485 );
or \U$4583 ( \4682 , \4680 , \4681 );
nand \U$4584 ( \4683 , \4682 , \1506 );
nand \U$4585 ( \4684 , \4679 , \4683 );
buf \U$4586 ( \4685 , \4684 );
xor \U$4587 ( \4686 , \4676 , \4685 );
buf \U$4588 ( \4687 , \1459 );
not \U$4589 ( \4688 , \4687 );
buf \U$4590 ( \4689 , \861 );
not \U$4591 ( \4690 , \4689 );
buf \U$4592 ( \4691 , \4690 );
buf \U$4595 ( \4692 , \4691 );
buf \U$4596 ( \4693 , \4692 );
not \U$4597 ( \4694 , \4693 );
or \U$4598 ( \4695 , \4688 , \4694 );
buf \U$4599 ( \4696 , \284 );
buf \U$4600 ( \4697 , RIc0d81b8_25);
buf \U$4601 ( \4698 , RIc0d9658_69);
xor \U$4602 ( \4699 , \4697 , \4698 );
buf \U$4603 ( \4700 , \4699 );
buf \U$4604 ( \4701 , \4700 );
nand \U$4605 ( \4702 , \4696 , \4701 );
buf \U$4606 ( \4703 , \4702 );
buf \U$4607 ( \4704 , \4703 );
nand \U$4608 ( \4705 , \4695 , \4704 );
buf \U$4609 ( \4706 , \4705 );
buf \U$4610 ( \4707 , \4706 );
buf \U$4611 ( \4708 , \1476 );
not \U$4612 ( \4709 , \4708 );
buf \U$4613 ( \4710 , \437 );
not \U$4614 ( \4711 , \4710 );
or \U$4615 ( \4712 , \4709 , \4711 );
buf \U$4616 ( \4713 , RIc0d7858_5);
buf \U$4617 ( \4714 , RIc0d9fb8_89);
xnor \U$4618 ( \4715 , \4713 , \4714 );
buf \U$4619 ( \4716 , \4715 );
buf \U$4620 ( \4717 , \4716 );
not \U$4621 ( \4718 , \4717 );
buf \U$4622 ( \4719 , \442 );
nand \U$4623 ( \4720 , \4718 , \4719 );
buf \U$4624 ( \4721 , \4720 );
buf \U$4625 ( \4722 , \4721 );
nand \U$4626 ( \4723 , \4712 , \4722 );
buf \U$4627 ( \4724 , \4723 );
buf \U$4628 ( \4725 , \4724 );
xor \U$4629 ( \4726 , \4707 , \4725 );
buf \U$4630 ( \4727 , \812 );
buf \U$4631 ( \4728 , \2797 );
or \U$4632 ( \4729 , \4727 , \4728 );
buf \U$4633 ( \4730 , \819 );
buf \U$4634 ( \4731 , RIc0d7948_7);
buf \U$4635 ( \4732 , RIc0d9ec8_87);
xor \U$4636 ( \4733 , \4731 , \4732 );
buf \U$4637 ( \4734 , \4733 );
buf \U$4638 ( \4735 , \4734 );
not \U$4639 ( \4736 , \4735 );
buf \U$4640 ( \4737 , \4736 );
buf \U$4641 ( \4738 , \4737 );
or \U$4642 ( \4739 , \4730 , \4738 );
nand \U$4643 ( \4740 , \4729 , \4739 );
buf \U$4644 ( \4741 , \4740 );
buf \U$4645 ( \4742 , \4741 );
xor \U$4646 ( \4743 , \4726 , \4742 );
buf \U$4647 ( \4744 , \4743 );
buf \U$4648 ( \4745 , \4744 );
xor \U$4649 ( \4746 , \4686 , \4745 );
buf \U$4650 ( \4747 , \4746 );
buf \U$4651 ( \4748 , \4747 );
xor \U$4652 ( \4749 , \4670 , \4748 );
buf \U$4653 ( \4750 , \4749 );
buf \U$4654 ( \4751 , \4750 );
xor \U$4655 ( \4752 , \1336 , \1342 );
and \U$4656 ( \4753 , \4752 , \1521 );
and \U$4657 ( \4754 , \1336 , \1342 );
or \U$4658 ( \4755 , \4753 , \4754 );
buf \U$4659 ( \4756 , \4755 );
buf \U$4660 ( \4757 , \4756 );
xor \U$4661 ( \4758 , \4751 , \4757 );
xor \U$4662 ( \4759 , \1662 , \1668 );
and \U$4663 ( \4760 , \4759 , \1726 );
and \U$4664 ( \4761 , \1662 , \1668 );
or \U$4665 ( \4762 , \4760 , \4761 );
buf \U$4666 ( \4763 , \4762 );
buf \U$4667 ( \4764 , \4763 );
xor \U$4668 ( \4765 , \1383 , \1448 );
and \U$4669 ( \4766 , \4765 , \1518 );
and \U$4670 ( \4767 , \1383 , \1448 );
or \U$4671 ( \4768 , \4766 , \4767 );
buf \U$4672 ( \4769 , \4768 );
buf \U$4673 ( \4770 , \4769 );
xor \U$4674 ( \4771 , \4764 , \4770 );
buf \U$4675 ( \4772 , \1356 );
not \U$4676 ( \4773 , \4772 );
buf \U$4677 ( \4774 , \397 );
not \U$4678 ( \4775 , \4774 );
or \U$4679 ( \4776 , \4773 , \4775 );
buf \U$4680 ( \4777 , \403 );
buf \U$4681 ( \4778 , RIc0d7d08_15);
buf \U$4682 ( \4779 , RIc0d9b08_79);
xor \U$4683 ( \4780 , \4778 , \4779 );
buf \U$4684 ( \4781 , \4780 );
buf \U$4685 ( \4782 , \4781 );
nand \U$4686 ( \4783 , \4777 , \4782 );
buf \U$4687 ( \4784 , \4783 );
buf \U$4688 ( \4785 , \4784 );
nand \U$4689 ( \4786 , \4776 , \4785 );
buf \U$4690 ( \4787 , \4786 );
buf \U$4691 ( \4788 , \1500 );
not \U$4692 ( \4789 , \4788 );
buf \U$4693 ( \4790 , \476 );
not \U$4694 ( \4791 , \4790 );
or \U$4695 ( \4792 , \4789 , \4791 );
buf \U$4696 ( \4793 , \4008 );
buf \U$4697 ( \4794 , RIc0d7678_1);
buf \U$4698 ( \4795 , RIc0da198_93);
xor \U$4699 ( \4796 , \4794 , \4795 );
buf \U$4700 ( \4797 , \4796 );
buf \U$4701 ( \4798 , \4797 );
nand \U$4702 ( \4799 , \4793 , \4798 );
buf \U$4703 ( \4800 , \4799 );
buf \U$4704 ( \4801 , \4800 );
nand \U$4705 ( \4802 , \4792 , \4801 );
buf \U$4706 ( \4803 , \4802 );
xor \U$4707 ( \4804 , \4787 , \4803 );
buf \U$4708 ( \4805 , \4804 );
buf \U$4709 ( \4806 , \2780 );
not \U$4710 ( \4807 , \4806 );
buf \U$4711 ( \4808 , \4807 );
buf \U$4712 ( \4809 , \4808 );
not \U$4713 ( \4810 , \4809 );
buf \U$4714 ( \4811 , \1064 );
not \U$4715 ( \4812 , \4811 );
or \U$4716 ( \4813 , \4810 , \4812 );
buf \U$4717 ( \4814 , \1078 );
buf \U$4718 ( \4815 , RIc0d7c18_13);
buf \U$4719 ( \4816 , RIc0d9bf8_81);
xor \U$4720 ( \4817 , \4815 , \4816 );
buf \U$4721 ( \4818 , \4817 );
buf \U$4722 ( \4819 , \4818 );
nand \U$4723 ( \4820 , \4814 , \4819 );
buf \U$4724 ( \4821 , \4820 );
buf \U$4725 ( \4822 , \4821 );
nand \U$4726 ( \4823 , \4813 , \4822 );
buf \U$4727 ( \4824 , \4823 );
buf \U$4728 ( \4825 , \4824 );
xnor \U$4729 ( \4826 , \4805 , \4825 );
buf \U$4730 ( \4827 , \4826 );
buf \U$4731 ( \4828 , \4827 );
not \U$4732 ( \4829 , \4828 );
buf \U$4733 ( \4830 , \2755 );
not \U$4734 ( \4831 , \4830 );
buf \U$4735 ( \4832 , \574 );
not \U$4736 ( \4833 , \4832 );
or \U$4737 ( \4834 , \4831 , \4833 );
buf \U$4738 ( \4835 , RIc0d7b28_11);
buf \U$4739 ( \4836 , RIc0d9ce8_83);
xnor \U$4740 ( \4837 , \4835 , \4836 );
buf \U$4741 ( \4838 , \4837 );
buf \U$4742 ( \4839 , \4838 );
not \U$4743 ( \4840 , \4839 );
buf \U$4744 ( \4841 , \993 );
nand \U$4745 ( \4842 , \4840 , \4841 );
buf \U$4746 ( \4843 , \4842 );
buf \U$4747 ( \4844 , \4843 );
nand \U$4748 ( \4845 , \4834 , \4844 );
buf \U$4749 ( \4846 , \4845 );
buf \U$4750 ( \4847 , \344 );
not \U$4751 ( \4848 , \4847 );
buf \U$4752 ( \4849 , \4848 );
buf \U$4753 ( \4850 , \4849 );
not \U$4754 ( \4851 , \4850 );
buf \U$4755 ( \4852 , \333 );
not \U$4756 ( \4853 , \4852 );
or \U$4757 ( \4854 , \4851 , \4853 );
buf \U$4758 ( \4855 , RIc0da288_95);
nand \U$4759 ( \4856 , \4854 , \4855 );
buf \U$4760 ( \4857 , \4856 );
buf \U$4761 ( \4858 , \4857 );
not \U$4762 ( \4859 , \4858 );
buf \U$4763 ( \4860 , \4859 );
and \U$4764 ( \4861 , \4846 , \4860 );
not \U$4765 ( \4862 , \4846 );
and \U$4766 ( \4863 , \4862 , \4857 );
or \U$4767 ( \4864 , \4861 , \4863 );
buf \U$4768 ( \4865 , \4864 );
buf \U$4769 ( \4866 , \2269 );
not \U$4770 ( \4867 , \4866 );
buf \U$4771 ( \4868 , \4867 );
buf \U$4772 ( \4869 , \4868 );
not \U$4773 ( \4870 , \4869 );
buf \U$4774 ( \4871 , \2823 );
not \U$4775 ( \4872 , \4871 );
and \U$4776 ( \4873 , \4870 , \4872 );
buf \U$4777 ( \4874 , \2927 );
buf \U$4778 ( \4875 , RIc0d80c8_23);
buf \U$4779 ( \4876 , RIc0d9748_71);
xor \U$4780 ( \4877 , \4875 , \4876 );
buf \U$4781 ( \4878 , \4877 );
buf \U$4782 ( \4879 , \4878 );
and \U$4783 ( \4880 , \4874 , \4879 );
buf \U$4784 ( \4881 , \4880 );
buf \U$4785 ( \4882 , \4881 );
nor \U$4786 ( \4883 , \4873 , \4882 );
buf \U$4787 ( \4884 , \4883 );
buf \U$4788 ( \4885 , \4884 );
xnor \U$4789 ( \4886 , \4865 , \4885 );
buf \U$4790 ( \4887 , \4886 );
buf \U$4791 ( \4888 , \4887 );
not \U$4792 ( \4889 , \4888 );
or \U$4793 ( \4890 , \4829 , \4889 );
buf \U$4794 ( \4891 , \4887 );
buf \U$4795 ( \4892 , \4827 );
or \U$4796 ( \4893 , \4891 , \4892 );
nand \U$4797 ( \4894 , \4890 , \4893 );
buf \U$4798 ( \4895 , \4894 );
buf \U$4799 ( \4896 , \4895 );
and \U$4800 ( \4897 , \1237 , \1238 );
buf \U$4801 ( \4898 , \4897 );
buf \U$4802 ( \4899 , \4898 );
buf \U$4803 ( \4900 , \1409 );
not \U$4804 ( \4901 , \4900 );
buf \U$4805 ( \4902 , \1822 );
not \U$4806 ( \4903 , \4902 );
buf \U$4807 ( \4904 , \4903 );
buf \U$4808 ( \4905 , \4904 );
not \U$4809 ( \4906 , \4905 );
buf \U$4810 ( \4907 , \4906 );
buf \U$4811 ( \4908 , \4907 );
not \U$4812 ( \4909 , \4908 );
or \U$4813 ( \4910 , \4901 , \4909 );
buf \U$4814 ( \4911 , \686 );
buf \U$4815 ( \4912 , RIc0d82a8_27);
buf \U$4816 ( \4913 , RIc0d9568_67);
xor \U$4817 ( \4914 , \4912 , \4913 );
buf \U$4818 ( \4915 , \4914 );
buf \U$4819 ( \4916 , \4915 );
nand \U$4820 ( \4917 , \4911 , \4916 );
buf \U$4821 ( \4918 , \4917 );
buf \U$4822 ( \4919 , \4918 );
nand \U$4823 ( \4920 , \4910 , \4919 );
buf \U$4824 ( \4921 , \4920 );
buf \U$4825 ( \4922 , \4921 );
xor \U$4826 ( \4923 , \4899 , \4922 );
buf \U$4827 ( \4924 , \521 );
buf \U$4828 ( \4925 , \2733 );
or \U$4829 ( \4926 , \4924 , \4925 );
buf \U$4830 ( \4927 , \711 );
buf \U$4831 ( \4928 , RIc0d7768_3);
buf \U$4832 ( \4929 , RIc0da0a8_91);
xnor \U$4833 ( \4930 , \4928 , \4929 );
buf \U$4834 ( \4931 , \4930 );
buf \U$4835 ( \4932 , \4931 );
or \U$4836 ( \4933 , \4927 , \4932 );
nand \U$4837 ( \4934 , \4926 , \4933 );
buf \U$4838 ( \4935 , \4934 );
buf \U$4839 ( \4936 , \4935 );
xor \U$4840 ( \4937 , \4923 , \4936 );
buf \U$4841 ( \4938 , \4937 );
buf \U$4842 ( \4939 , \4938 );
and \U$4843 ( \4940 , \4896 , \4939 );
not \U$4844 ( \4941 , \4896 );
buf \U$4845 ( \4942 , \4938 );
not \U$4846 ( \4943 , \4942 );
buf \U$4847 ( \4944 , \4943 );
buf \U$4848 ( \4945 , \4944 );
and \U$4849 ( \4946 , \4941 , \4945 );
nor \U$4850 ( \4947 , \4940 , \4946 );
buf \U$4851 ( \4948 , \4947 );
buf \U$4852 ( \4949 , \4948 );
xor \U$4853 ( \4950 , \4771 , \4949 );
buf \U$4854 ( \4951 , \4950 );
buf \U$4855 ( \4952 , \4951 );
xor \U$4856 ( \4953 , \4758 , \4952 );
buf \U$4857 ( \4954 , \4953 );
buf \U$4858 ( \4955 , \4954 );
xor \U$4859 ( \4956 , \2715 , \3026 );
and \U$4860 ( \4957 , \4956 , \3106 );
and \U$4861 ( \4958 , \2715 , \3026 );
or \U$4862 ( \4959 , \4957 , \4958 );
buf \U$4863 ( \4960 , \4959 );
buf \U$4864 ( \4961 , \4960 );
xor \U$4865 ( \4962 , \4955 , \4961 );
xor \U$4866 ( \4963 , \2721 , \2982 );
and \U$4867 ( \4964 , \4963 , \3023 );
and \U$4868 ( \4965 , \2721 , \2982 );
or \U$4869 ( \4966 , \4964 , \4965 );
buf \U$4870 ( \4967 , \4966 );
buf \U$4871 ( \4968 , \4967 );
xor \U$4872 ( \4969 , \2788 , \2847 );
and \U$4873 ( \4970 , \4969 , \2979 );
and \U$4874 ( \4971 , \2788 , \2847 );
or \U$4875 ( \4972 , \4970 , \4971 );
buf \U$4876 ( \4973 , \4972 );
buf \U$4877 ( \4974 , \4973 );
buf \U$4878 ( \4975 , RIc0d9478_65);
buf \U$4879 ( \4976 , RIc0d8398_29);
xor \U$4880 ( \4977 , \4975 , \4976 );
buf \U$4881 ( \4978 , \4977 );
buf \U$4882 ( \4979 , \4978 );
not \U$4883 ( \4980 , \4979 );
buf \U$4884 ( \4981 , \1235 );
not \U$4885 ( \4982 , \4981 );
or \U$4886 ( \4983 , \4980 , \4982 );
buf \U$4887 ( \4984 , \1700 );
not \U$4888 ( \4985 , \4984 );
buf \U$4889 ( \4986 , \1224 );
nand \U$4890 ( \4987 , \4985 , \4986 );
buf \U$4891 ( \4988 , \4987 );
buf \U$4892 ( \4989 , \4988 );
nand \U$4893 ( \4990 , \4983 , \4989 );
buf \U$4894 ( \4991 , \4990 );
buf \U$4895 ( \4992 , \4991 );
buf \U$4896 ( \4993 , \3816 );
not \U$4897 ( \4994 , \4993 );
buf \U$4898 ( \4995 , \1375 );
not \U$4899 ( \4996 , \4995 );
and \U$4900 ( \4997 , \4994 , \4996 );
buf \U$4901 ( \4998 , \1143 );
xor \U$4902 ( \4999 , RIc0d9928_75, RIc0d7ee8_19);
buf \U$4903 ( \5000 , \4999 );
and \U$4904 ( \5001 , \4998 , \5000 );
buf \U$4905 ( \5002 , \5001 );
buf \U$4906 ( \5003 , \5002 );
nor \U$4907 ( \5004 , \4997 , \5003 );
buf \U$4908 ( \5005 , \5004 );
buf \U$4909 ( \5006 , \5005 );
not \U$4910 ( \5007 , \5006 );
buf \U$4911 ( \5008 , \5007 );
buf \U$4912 ( \5009 , \5008 );
and \U$4913 ( \5010 , \4992 , \5009 );
not \U$4914 ( \5011 , \4992 );
buf \U$4915 ( \5012 , \5005 );
and \U$4916 ( \5013 , \5011 , \5012 );
nor \U$4917 ( \5014 , \5010 , \5013 );
buf \U$4918 ( \5015 , \5014 );
buf \U$4919 ( \5016 , \5015 );
buf \U$4920 ( \5017 , \1431 );
not \U$4921 ( \5018 , \5017 );
buf \U$4922 ( \5019 , \5018 );
not \U$4923 ( \5020 , \5019 );
not \U$4924 ( \5021 , \1440 );
and \U$4925 ( \5022 , \5020 , \5021 );
buf \U$4926 ( \5023 , RIc0d7df8_17);
buf \U$4927 ( \5024 , RIc0d9a18_77);
xor \U$4928 ( \5025 , \5023 , \5024 );
buf \U$4929 ( \5026 , \5025 );
and \U$4930 ( \5027 , \3742 , \5026 );
nor \U$4931 ( \5028 , \5022 , \5027 );
buf \U$4932 ( \5029 , \5028 );
not \U$4933 ( \5030 , \5029 );
buf \U$4934 ( \5031 , \5030 );
buf \U$4935 ( \5032 , \5031 );
and \U$4936 ( \5033 , \5016 , \5032 );
not \U$4937 ( \5034 , \5016 );
buf \U$4938 ( \5035 , \5028 );
and \U$4939 ( \5036 , \5034 , \5035 );
nor \U$4940 ( \5037 , \5033 , \5036 );
buf \U$4941 ( \5038 , \5037 );
buf \U$4942 ( \5039 , \5038 );
buf \U$4943 ( \5040 , \1685 );
not \U$4944 ( \5041 , \5040 );
buf \U$4945 ( \5042 , \1677 );
not \U$4946 ( \5043 , \5042 );
or \U$4947 ( \5044 , \5041 , \5043 );
buf \U$4948 ( \5045 , \2882 );
buf \U$4949 ( \5046 , RIc0d7fd8_21);
buf \U$4950 ( \5047 , RIc0d9838_73);
xor \U$4951 ( \5048 , \5046 , \5047 );
buf \U$4952 ( \5049 , \5048 );
buf \U$4953 ( \5050 , \5049 );
nand \U$4954 ( \5051 , \5045 , \5050 );
buf \U$4955 ( \5052 , \5051 );
buf \U$4956 ( \5053 , \5052 );
nand \U$4957 ( \5054 , \5044 , \5053 );
buf \U$4958 ( \5055 , \5054 );
buf \U$4959 ( \5056 , \5055 );
not \U$4960 ( \5057 , \954 );
not \U$4961 ( \5058 , \1396 );
and \U$4962 ( \5059 , \5057 , \5058 );
buf \U$4963 ( \5060 , RIc0d7a38_9);
buf \U$4964 ( \5061 , RIc0d9dd8_85);
xor \U$4965 ( \5062 , \5060 , \5061 );
buf \U$4966 ( \5063 , \5062 );
and \U$4967 ( \5064 , \921 , \5063 );
nor \U$4968 ( \5065 , \5059 , \5064 );
buf \U$4969 ( \5066 , \5065 );
not \U$4970 ( \5067 , \5066 );
buf \U$4971 ( \5068 , \5067 );
buf \U$4972 ( \5069 , \5068 );
and \U$4973 ( \5070 , \5056 , \5069 );
not \U$4974 ( \5071 , \5056 );
buf \U$4975 ( \5072 , \5065 );
and \U$4976 ( \5073 , \5071 , \5072 );
nor \U$4977 ( \5074 , \5070 , \5073 );
buf \U$4978 ( \5075 , \5074 );
buf \U$4979 ( \5076 , \5075 );
buf \U$4980 ( \5077 , \2805 );
and \U$4981 ( \5078 , \5076 , \5077 );
not \U$4982 ( \5079 , \5076 );
buf \U$4983 ( \5080 , \2808 );
and \U$4984 ( \5081 , \5079 , \5080 );
nor \U$4985 ( \5082 , \5078 , \5081 );
buf \U$4986 ( \5083 , \5082 );
buf \U$4987 ( \5084 , \5083 );
xor \U$4988 ( \5085 , \5039 , \5084 );
xor \U$4989 ( \5086 , \1311 , \1326 );
and \U$4990 ( \5087 , \5086 , \1333 );
and \U$4991 ( \5088 , \1311 , \1326 );
or \U$4992 ( \5089 , \5087 , \5088 );
buf \U$4993 ( \5090 , \5089 );
buf \U$4994 ( \5091 , \5090 );
xor \U$4995 ( \5092 , \5085 , \5091 );
buf \U$4996 ( \5093 , \5092 );
buf \U$4997 ( \5094 , \5093 );
xor \U$4998 ( \5095 , \4974 , \5094 );
xor \U$4999 ( \5096 , \1629 , \1646 );
and \U$5000 ( \5097 , \5096 , \1729 );
and \U$5001 ( \5098 , \1629 , \1646 );
or \U$5002 ( \5099 , \5097 , \5098 );
buf \U$5003 ( \5100 , \5099 );
buf \U$5004 ( \5101 , \5100 );
xor \U$5005 ( \5102 , \5095 , \5101 );
buf \U$5006 ( \5103 , \5102 );
buf \U$5007 ( \5104 , \5103 );
xor \U$5008 ( \5105 , \4968 , \5104 );
xor \U$5009 ( \5106 , \1305 , \1524 );
and \U$5010 ( \5107 , \5106 , \1732 );
and \U$5011 ( \5108 , \1305 , \1524 );
or \U$5012 ( \5109 , \5107 , \5108 );
buf \U$5013 ( \5110 , \5109 );
buf \U$5014 ( \5111 , \5110 );
xor \U$5015 ( \5112 , \5105 , \5111 );
buf \U$5016 ( \5113 , \5112 );
buf \U$5017 ( \5114 , \5113 );
xor \U$5018 ( \5115 , \4962 , \5114 );
buf \U$5019 ( \5116 , \5115 );
buf \U$5020 ( \5117 , \5116 );
not \U$5021 ( \5118 , \5117 );
buf \U$5022 ( \5119 , \5118 );
buf \U$5023 ( \5120 , \5119 );
xor \U$5024 ( \5121 , \1735 , \3109 );
and \U$5025 ( \5122 , \5121 , \3942 );
and \U$5026 ( \5123 , \1735 , \3109 );
or \U$5027 ( \5124 , \5122 , \5123 );
buf \U$5028 ( \5125 , \5124 );
buf \U$5029 ( \5126 , \5125 );
not \U$5030 ( \5127 , \5126 );
buf \U$5031 ( \5128 , \5127 );
buf \U$5032 ( \5129 , \5128 );
nand \U$5033 ( \5130 , \5120 , \5129 );
buf \U$5034 ( \5131 , \5130 );
buf \U$5035 ( \5132 , \5131 );
nand \U$5036 ( \5133 , \4618 , \5132 );
buf \U$5037 ( \5134 , \5133 );
buf \U$5038 ( \5135 , \5134 );
not \U$5039 ( \5136 , \5135 );
buf \U$5040 ( \5137 , \4734 );
not \U$5041 ( \5138 , \5137 );
buf \U$5042 ( \5139 , \4527 );
not \U$5043 ( \5140 , \5139 );
or \U$5044 ( \5141 , \5138 , \5140 );
buf \U$5045 ( \5142 , \816 );
buf \U$5046 ( \5143 , RIc0d78d0_6);
buf \U$5047 ( \5144 , RIc0d9ec8_87);
xor \U$5048 ( \5145 , \5143 , \5144 );
buf \U$5049 ( \5146 , \5145 );
buf \U$5050 ( \5147 , \5146 );
nand \U$5051 ( \5148 , \5142 , \5147 );
buf \U$5052 ( \5149 , \5148 );
buf \U$5053 ( \5150 , \5149 );
nand \U$5054 ( \5151 , \5141 , \5150 );
buf \U$5055 ( \5152 , \5151 );
buf \U$5056 ( \5153 , \5152 );
not \U$5057 ( \5154 , \5153 );
buf \U$5058 ( \5155 , \5154 );
buf \U$5059 ( \5156 , \5155 );
xor \U$5060 ( \5157 , \4899 , \4922 );
and \U$5061 ( \5158 , \5157 , \4936 );
and \U$5062 ( \5159 , \4899 , \4922 );
or \U$5063 ( \5160 , \5158 , \5159 );
buf \U$5064 ( \5161 , \5160 );
buf \U$5065 ( \5162 , \5161 );
xor \U$5066 ( \5163 , \5156 , \5162 );
xor \U$5067 ( \5164 , \4707 , \4725 );
and \U$5068 ( \5165 , \5164 , \4742 );
and \U$5069 ( \5166 , \4707 , \4725 );
or \U$5070 ( \5167 , \5165 , \5166 );
buf \U$5071 ( \5168 , \5167 );
buf \U$5072 ( \5169 , \5168 );
xor \U$5073 ( \5170 , \5163 , \5169 );
buf \U$5074 ( \5171 , \5170 );
buf \U$5075 ( \5172 , \5171 );
xor \U$5076 ( \5173 , \4644 , \4659 );
and \U$5077 ( \5174 , \5173 , \4666 );
and \U$5078 ( \5175 , \4644 , \4659 );
or \U$5079 ( \5176 , \5174 , \5175 );
buf \U$5080 ( \5177 , \5176 );
buf \U$5081 ( \5178 , \5177 );
xor \U$5082 ( \5179 , \5172 , \5178 );
buf \U$5083 ( \5180 , \4824 );
not \U$5084 ( \5181 , \5180 );
buf \U$5085 ( \5182 , \4787 );
not \U$5086 ( \5183 , \5182 );
or \U$5087 ( \5184 , \5181 , \5183 );
buf \U$5088 ( \5185 , \4787 );
buf \U$5089 ( \5186 , \4824 );
or \U$5090 ( \5187 , \5185 , \5186 );
buf \U$5091 ( \5188 , \4803 );
nand \U$5092 ( \5189 , \5187 , \5188 );
buf \U$5093 ( \5190 , \5189 );
buf \U$5094 ( \5191 , \5190 );
nand \U$5095 ( \5192 , \5184 , \5191 );
buf \U$5096 ( \5193 , \5192 );
buf \U$5097 ( \5194 , \5008 );
not \U$5098 ( \5195 , \5194 );
buf \U$5099 ( \5196 , \5031 );
not \U$5100 ( \5197 , \5196 );
or \U$5101 ( \5198 , \5195 , \5197 );
buf \U$5102 ( \5199 , \5005 );
not \U$5103 ( \5200 , \5199 );
buf \U$5104 ( \5201 , \5028 );
not \U$5105 ( \5202 , \5201 );
or \U$5106 ( \5203 , \5200 , \5202 );
buf \U$5107 ( \5204 , \4991 );
nand \U$5108 ( \5205 , \5203 , \5204 );
buf \U$5109 ( \5206 , \5205 );
buf \U$5110 ( \5207 , \5206 );
nand \U$5111 ( \5208 , \5198 , \5207 );
buf \U$5112 ( \5209 , \5208 );
xor \U$5113 ( \5210 , \5193 , \5209 );
buf \U$5114 ( \5211 , \4884 );
not \U$5115 ( \5212 , \5211 );
buf \U$5116 ( \5213 , \4860 );
not \U$5117 ( \5214 , \5213 );
or \U$5118 ( \5215 , \5212 , \5214 );
buf \U$5119 ( \5216 , \4846 );
nand \U$5120 ( \5217 , \5215 , \5216 );
buf \U$5121 ( \5218 , \5217 );
buf \U$5122 ( \5219 , \5218 );
buf \U$5123 ( \5220 , \4884 );
not \U$5124 ( \5221 , \5220 );
buf \U$5125 ( \5222 , \4857 );
nand \U$5126 ( \5223 , \5221 , \5222 );
buf \U$5127 ( \5224 , \5223 );
buf \U$5128 ( \5225 , \5224 );
nand \U$5129 ( \5226 , \5219 , \5225 );
buf \U$5130 ( \5227 , \5226 );
xor \U$5131 ( \5228 , \5210 , \5227 );
buf \U$5132 ( \5229 , \5228 );
xor \U$5133 ( \5230 , \5179 , \5229 );
buf \U$5134 ( \5231 , \5230 );
buf \U$5135 ( \5232 , \5231 );
xor \U$5136 ( \5233 , \4764 , \4770 );
and \U$5137 ( \5234 , \5233 , \4949 );
and \U$5138 ( \5235 , \4764 , \4770 );
or \U$5139 ( \5236 , \5234 , \5235 );
buf \U$5140 ( \5237 , \5236 );
buf \U$5141 ( \5238 , \5237 );
xor \U$5142 ( \5239 , \5232 , \5238 );
xor \U$5143 ( \5240 , \4676 , \4685 );
and \U$5144 ( \5241 , \5240 , \4745 );
and \U$5145 ( \5242 , \4676 , \4685 );
or \U$5146 ( \5243 , \5241 , \5242 );
buf \U$5147 ( \5244 , \5243 );
buf \U$5148 ( \5245 , \5244 );
buf \U$5149 ( \5246 , \4944 );
not \U$5150 ( \5247 , \5246 );
buf \U$5151 ( \5248 , \4827 );
not \U$5152 ( \5249 , \5248 );
or \U$5153 ( \5250 , \5247 , \5249 );
buf \U$5154 ( \5251 , \4887 );
nand \U$5155 ( \5252 , \5250 , \5251 );
buf \U$5156 ( \5253 , \5252 );
buf \U$5157 ( \5254 , \5253 );
buf \U$5158 ( \5255 , \4827 );
not \U$5159 ( \5256 , \5255 );
buf \U$5160 ( \5257 , \4938 );
nand \U$5161 ( \5258 , \5256 , \5257 );
buf \U$5162 ( \5259 , \5258 );
buf \U$5163 ( \5260 , \5259 );
nand \U$5164 ( \5261 , \5254 , \5260 );
buf \U$5165 ( \5262 , \5261 );
buf \U$5166 ( \5263 , \5262 );
xor \U$5167 ( \5264 , \5245 , \5263 );
buf \U$5168 ( \5265 , \4915 );
not \U$5169 ( \5266 , \5265 );
buf \U$5170 ( \5267 , \4907 );
not \U$5171 ( \5268 , \5267 );
or \U$5172 ( \5269 , \5266 , \5268 );
buf \U$5173 ( \5270 , \686 );
buf \U$5174 ( \5271 , RIc0d8230_26);
buf \U$5175 ( \5272 , RIc0d9568_67);
xor \U$5176 ( \5273 , \5271 , \5272 );
buf \U$5177 ( \5274 , \5273 );
buf \U$5178 ( \5275 , \5274 );
nand \U$5179 ( \5276 , \5270 , \5275 );
buf \U$5180 ( \5277 , \5276 );
buf \U$5181 ( \5278 , \5277 );
nand \U$5182 ( \5279 , \5269 , \5278 );
buf \U$5183 ( \5280 , \5279 );
buf \U$5184 ( \5281 , \5280 );
buf \U$5185 ( \5282 , \4878 );
not \U$5186 ( \5283 , \5282 );
buf \U$5187 ( \5284 , \1263 );
not \U$5188 ( \5285 , \5284 );
or \U$5189 ( \5286 , \5283 , \5285 );
buf \U$5190 ( \5287 , \2927 );
buf \U$5191 ( \5288 , RIc0d8050_22);
buf \U$5192 ( \5289 , RIc0d9748_71);
xor \U$5193 ( \5290 , \5288 , \5289 );
buf \U$5194 ( \5291 , \5290 );
buf \U$5195 ( \5292 , \5291 );
nand \U$5196 ( \5293 , \5287 , \5292 );
buf \U$5197 ( \5294 , \5293 );
buf \U$5198 ( \5295 , \5294 );
nand \U$5199 ( \5296 , \5286 , \5295 );
buf \U$5200 ( \5297 , \5296 );
buf \U$5201 ( \5298 , \5297 );
xor \U$5202 ( \5299 , \5281 , \5298 );
buf \U$5203 ( \5300 , \5063 );
not \U$5204 ( \5301 , \5300 );
buf \U$5205 ( \5302 , \2396 );
not \U$5206 ( \5303 , \5302 );
buf \U$5207 ( \5304 , \5303 );
buf \U$5210 ( \5305 , \5304 );
buf \U$5211 ( \5306 , \5305 );
not \U$5212 ( \5307 , \5306 );
or \U$5213 ( \5308 , \5301 , \5307 );
buf \U$5214 ( \5309 , \2960 );
buf \U$5215 ( \5310 , RIc0d79c0_8);
buf \U$5216 ( \5311 , RIc0d9dd8_85);
xor \U$5217 ( \5312 , \5310 , \5311 );
buf \U$5218 ( \5313 , \5312 );
buf \U$5219 ( \5314 , \5313 );
nand \U$5220 ( \5315 , \5309 , \5314 );
buf \U$5221 ( \5316 , \5315 );
buf \U$5222 ( \5317 , \5316 );
nand \U$5223 ( \5318 , \5308 , \5317 );
buf \U$5224 ( \5319 , \5318 );
buf \U$5225 ( \5320 , \5319 );
xor \U$5226 ( \5321 , \5299 , \5320 );
buf \U$5227 ( \5322 , \5321 );
buf \U$5228 ( \5323 , \5322 );
buf \U$5229 ( \5324 , \4999 );
not \U$5230 ( \5325 , \5324 );
buf \U$5231 ( \5326 , \2124 );
not \U$5232 ( \5327 , \5326 );
or \U$5233 ( \5328 , \5325 , \5327 );
buf \U$5234 ( \5329 , \1565 );
buf \U$5235 ( \5330 , RIc0d7e70_18);
buf \U$5236 ( \5331 , RIc0d9928_75);
xor \U$5237 ( \5332 , \5330 , \5331 );
buf \U$5238 ( \5333 , \5332 );
buf \U$5239 ( \5334 , \5333 );
nand \U$5240 ( \5335 , \5329 , \5334 );
buf \U$5241 ( \5336 , \5335 );
buf \U$5242 ( \5337 , \5336 );
nand \U$5243 ( \5338 , \5328 , \5337 );
buf \U$5244 ( \5339 , \5338 );
buf \U$5245 ( \5340 , \5339 );
buf \U$5246 ( \5341 , \5026 );
not \U$5247 ( \5342 , \5341 );
buf \U$5248 ( \5343 , \1432 );
not \U$5249 ( \5344 , \5343 );
or \U$5250 ( \5345 , \5342 , \5344 );
buf \U$5251 ( \5346 , RIc0d7d80_16);
buf \U$5252 ( \5347 , RIc0d9a18_77);
xnor \U$5253 ( \5348 , \5346 , \5347 );
buf \U$5254 ( \5349 , \5348 );
buf \U$5255 ( \5350 , \5349 );
not \U$5256 ( \5351 , \5350 );
buf \U$5257 ( \5352 , \1196 );
nand \U$5258 ( \5353 , \5351 , \5352 );
buf \U$5259 ( \5354 , \5353 );
buf \U$5260 ( \5355 , \5354 );
nand \U$5261 ( \5356 , \5345 , \5355 );
buf \U$5262 ( \5357 , \5356 );
buf \U$5263 ( \5358 , \5357 );
xor \U$5264 ( \5359 , \5340 , \5358 );
buf \U$5265 ( \5360 , \842 );
not \U$5266 ( \5361 , \5360 );
buf \U$5267 ( \5362 , \5361 );
buf \U$5268 ( \5363 , \5362 );
buf \U$5269 ( \5364 , \4716 );
or \U$5270 ( \5365 , \5363 , \5364 );
buf \U$5271 ( \5366 , \846 );
not \U$5272 ( \5367 , \5366 );
buf \U$5273 ( \5368 , \5367 );
buf \U$5274 ( \5369 , \5368 );
buf \U$5275 ( \5370 , RIc0d9fb8_89);
buf \U$5276 ( \5371 , \489 );
and \U$5277 ( \5372 , \5370 , \5371 );
not \U$5278 ( \5373 , \5370 );
buf \U$5279 ( \5374 , RIc0d77e0_4);
and \U$5280 ( \5375 , \5373 , \5374 );
nor \U$5281 ( \5376 , \5372 , \5375 );
buf \U$5282 ( \5377 , \5376 );
buf \U$5283 ( \5378 , \5377 );
or \U$5284 ( \5379 , \5369 , \5378 );
nand \U$5285 ( \5380 , \5365 , \5379 );
buf \U$5286 ( \5381 , \5380 );
buf \U$5287 ( \5382 , \5381 );
xor \U$5288 ( \5383 , \5359 , \5382 );
buf \U$5289 ( \5384 , \5383 );
buf \U$5290 ( \5385 , \5384 );
xor \U$5291 ( \5386 , \5323 , \5385 );
buf \U$5292 ( \5387 , \5049 );
not \U$5293 ( \5388 , \5387 );
buf \U$5294 ( \5389 , \2871 );
not \U$5295 ( \5390 , \5389 );
or \U$5296 ( \5391 , \5388 , \5390 );
buf \U$5297 ( \5392 , \1856 );
buf \U$5298 ( \5393 , RIc0d7f60_20);
buf \U$5299 ( \5394 , RIc0d9838_73);
xor \U$5300 ( \5395 , \5393 , \5394 );
buf \U$5301 ( \5396 , \5395 );
buf \U$5302 ( \5397 , \5396 );
nand \U$5303 ( \5398 , \5392 , \5397 );
buf \U$5304 ( \5399 , \5398 );
buf \U$5305 ( \5400 , \5399 );
nand \U$5306 ( \5401 , \5391 , \5400 );
buf \U$5307 ( \5402 , \5401 );
buf \U$5308 ( \5403 , \4978 );
not \U$5309 ( \5404 , \5403 );
buf \U$5310 ( \5405 , \3781 );
not \U$5311 ( \5406 , \5405 );
or \U$5312 ( \5407 , \5404 , \5406 );
buf \U$5313 ( \5408 , \1229 );
buf \U$5314 ( \5409 , RIc0d9478_65);
buf \U$5315 ( \5410 , RIc0d8320_28);
xor \U$5316 ( \5411 , \5409 , \5410 );
buf \U$5317 ( \5412 , \5411 );
buf \U$5318 ( \5413 , \5412 );
nand \U$5319 ( \5414 , \5408 , \5413 );
buf \U$5320 ( \5415 , \5414 );
buf \U$5321 ( \5416 , \5415 );
nand \U$5322 ( \5417 , \5407 , \5416 );
buf \U$5323 ( \5418 , \5417 );
xor \U$5324 ( \5419 , \5402 , \5418 );
buf \U$5325 ( \5420 , \4931 );
not \U$5326 ( \5421 , \5420 );
buf \U$5327 ( \5422 , \5421 );
buf \U$5328 ( \5423 , \5422 );
not \U$5329 ( \5424 , \5423 );
buf \U$5330 ( \5425 , \524 );
not \U$5331 ( \5426 , \5425 );
or \U$5332 ( \5427 , \5424 , \5426 );
buf \U$5333 ( \5428 , \1933 );
buf \U$5334 ( \5429 , RIc0d76f0_2);
buf \U$5335 ( \5430 , RIc0da0a8_91);
xor \U$5336 ( \5431 , \5429 , \5430 );
buf \U$5337 ( \5432 , \5431 );
buf \U$5338 ( \5433 , \5432 );
nand \U$5339 ( \5434 , \5428 , \5433 );
buf \U$5340 ( \5435 , \5434 );
buf \U$5341 ( \5436 , \5435 );
nand \U$5342 ( \5437 , \5427 , \5436 );
buf \U$5343 ( \5438 , \5437 );
xor \U$5344 ( \5439 , \5419 , \5438 );
buf \U$5345 ( \5440 , \5439 );
xor \U$5346 ( \5441 , \5386 , \5440 );
buf \U$5347 ( \5442 , \5441 );
buf \U$5348 ( \5443 , \5442 );
xor \U$5349 ( \5444 , \5264 , \5443 );
buf \U$5350 ( \5445 , \5444 );
buf \U$5351 ( \5446 , \5445 );
xor \U$5352 ( \5447 , \5239 , \5446 );
buf \U$5353 ( \5448 , \5447 );
buf \U$5354 ( \5449 , \5448 );
xor \U$5355 ( \5450 , \4974 , \5094 );
and \U$5356 ( \5451 , \5450 , \5101 );
and \U$5357 ( \5452 , \4974 , \5094 );
or \U$5358 ( \5453 , \5451 , \5452 );
buf \U$5359 ( \5454 , \5453 );
buf \U$5360 ( \5455 , \5454 );
buf \U$5361 ( \5456 , \5065 );
not \U$5362 ( \5457 , \5456 );
buf \U$5363 ( \5458 , \2808 );
not \U$5364 ( \5459 , \5458 );
or \U$5365 ( \5460 , \5457 , \5459 );
buf \U$5366 ( \5461 , \5055 );
nand \U$5367 ( \5462 , \5460 , \5461 );
buf \U$5368 ( \5463 , \5462 );
buf \U$5369 ( \5464 , \5463 );
buf \U$5370 ( \5465 , \2805 );
buf \U$5371 ( \5466 , \5068 );
nand \U$5372 ( \5467 , \5465 , \5466 );
buf \U$5373 ( \5468 , \5467 );
buf \U$5374 ( \5469 , \5468 );
nand \U$5375 ( \5470 , \5464 , \5469 );
buf \U$5376 ( \5471 , \5470 );
buf \U$5377 ( \5472 , \5471 );
buf \U$5378 ( \5473 , RIc0d8410_30);
buf \U$5379 ( \5474 , RIc0d9478_65);
nand \U$5380 ( \5475 , \5473 , \5474 );
buf \U$5381 ( \5476 , \5475 );
buf \U$5382 ( \5477 , \4700 );
not \U$5383 ( \5478 , \5477 );
buf \U$5384 ( \5479 , \4692 );
not \U$5385 ( \5480 , \5479 );
or \U$5386 ( \5481 , \5478 , \5480 );
buf \U$5387 ( \5482 , \284 );
buf \U$5388 ( \5483 , RIc0d8140_24);
buf \U$5389 ( \5484 , RIc0d9658_69);
xor \U$5390 ( \5485 , \5483 , \5484 );
buf \U$5391 ( \5486 , \5485 );
buf \U$5392 ( \5487 , \5486 );
nand \U$5393 ( \5488 , \5482 , \5487 );
buf \U$5394 ( \5489 , \5488 );
buf \U$5395 ( \5490 , \5489 );
nand \U$5396 ( \5491 , \5481 , \5490 );
buf \U$5397 ( \5492 , \5491 );
xor \U$5398 ( \5493 , \5476 , \5492 );
buf \U$5399 ( \5494 , \4797 );
not \U$5400 ( \5495 , \5494 );
buf \U$5401 ( \5496 , \889 );
not \U$5402 ( \5497 , \5496 );
or \U$5403 ( \5498 , \5495 , \5497 );
buf \U$5404 ( \5499 , \481 );
buf \U$5405 ( \5500 , RIc0da198_93);
nand \U$5406 ( \5501 , \5499 , \5500 );
buf \U$5407 ( \5502 , \5501 );
buf \U$5408 ( \5503 , \5502 );
nand \U$5409 ( \5504 , \5498 , \5503 );
buf \U$5410 ( \5505 , \5504 );
xnor \U$5411 ( \5506 , \5493 , \5505 );
buf \U$5412 ( \5507 , \5506 );
xor \U$5413 ( \5508 , \5472 , \5507 );
buf \U$5414 ( \5509 , \989 );
buf \U$5415 ( \5510 , \4838 );
or \U$5416 ( \5511 , \5509 , \5510 );
buf \U$5417 ( \5512 , \996 );
buf \U$5418 ( \5513 , RIc0d7ab0_10);
buf \U$5419 ( \5514 , RIc0d9ce8_83);
xnor \U$5420 ( \5515 , \5513 , \5514 );
buf \U$5421 ( \5516 , \5515 );
buf \U$5422 ( \5517 , \5516 );
or \U$5423 ( \5518 , \5512 , \5517 );
nand \U$5424 ( \5519 , \5511 , \5518 );
buf \U$5425 ( \5520 , \5519 );
buf \U$5426 ( \5521 , \5520 );
not \U$5427 ( \5522 , \5521 );
buf \U$5428 ( \5523 , \5522 );
buf \U$5429 ( \5524 , \5523 );
not \U$5430 ( \5525 , \5524 );
buf \U$5431 ( \5526 , \4818 );
not \U$5432 ( \5527 , \5526 );
buf \U$5433 ( \5528 , \1064 );
not \U$5434 ( \5529 , \5528 );
or \U$5435 ( \5530 , \5527 , \5529 );
buf \U$5436 ( \5531 , RIc0d7ba0_12);
buf \U$5437 ( \5532 , RIc0d9bf8_81);
xnor \U$5438 ( \5533 , \5531 , \5532 );
buf \U$5439 ( \5534 , \5533 );
buf \U$5440 ( \5535 , \5534 );
not \U$5441 ( \5536 , \5535 );
buf \U$5442 ( \5537 , \1078 );
nand \U$5443 ( \5538 , \5536 , \5537 );
buf \U$5444 ( \5539 , \5538 );
buf \U$5445 ( \5540 , \5539 );
nand \U$5446 ( \5541 , \5530 , \5540 );
buf \U$5447 ( \5542 , \5541 );
buf \U$5448 ( \5543 , \4781 );
not \U$5449 ( \5544 , \5543 );
buf \U$5450 ( \5545 , \4509 );
not \U$5451 ( \5546 , \5545 );
or \U$5452 ( \5547 , \5544 , \5546 );
buf \U$5453 ( \5548 , \1026 );
buf \U$5454 ( \5549 , RIc0d7c90_14);
buf \U$5455 ( \5550 , RIc0d9b08_79);
xor \U$5456 ( \5551 , \5549 , \5550 );
buf \U$5457 ( \5552 , \5551 );
buf \U$5458 ( \5553 , \5552 );
nand \U$5459 ( \5554 , \5548 , \5553 );
buf \U$5460 ( \5555 , \5554 );
buf \U$5461 ( \5556 , \5555 );
nand \U$5462 ( \5557 , \5547 , \5556 );
buf \U$5463 ( \5558 , \5557 );
xor \U$5464 ( \5559 , \5542 , \5558 );
buf \U$5465 ( \5560 , \5559 );
not \U$5466 ( \5561 , \5560 );
or \U$5467 ( \5562 , \5525 , \5561 );
buf \U$5468 ( \5563 , \5559 );
buf \U$5469 ( \5564 , \5523 );
or \U$5470 ( \5565 , \5563 , \5564 );
nand \U$5471 ( \5566 , \5562 , \5565 );
buf \U$5472 ( \5567 , \5566 );
buf \U$5473 ( \5568 , \5567 );
xor \U$5474 ( \5569 , \5508 , \5568 );
buf \U$5475 ( \5570 , \5569 );
buf \U$5476 ( \5571 , \5570 );
xor \U$5477 ( \5572 , \5039 , \5084 );
and \U$5478 ( \5573 , \5572 , \5091 );
and \U$5479 ( \5574 , \5039 , \5084 );
or \U$5480 ( \5575 , \5573 , \5574 );
buf \U$5481 ( \5576 , \5575 );
buf \U$5482 ( \5577 , \5576 );
xor \U$5483 ( \5578 , \5571 , \5577 );
xor \U$5484 ( \5579 , \4624 , \4669 );
and \U$5485 ( \5580 , \5579 , \4748 );
and \U$5486 ( \5581 , \4624 , \4669 );
or \U$5487 ( \5582 , \5580 , \5581 );
buf \U$5488 ( \5583 , \5582 );
buf \U$5489 ( \5584 , \5583 );
xor \U$5490 ( \5585 , \5578 , \5584 );
buf \U$5491 ( \5586 , \5585 );
buf \U$5492 ( \5587 , \5586 );
xor \U$5493 ( \5588 , \5455 , \5587 );
xor \U$5494 ( \5589 , \4751 , \4757 );
and \U$5495 ( \5590 , \5589 , \4952 );
and \U$5496 ( \5591 , \4751 , \4757 );
or \U$5497 ( \5592 , \5590 , \5591 );
buf \U$5498 ( \5593 , \5592 );
buf \U$5499 ( \5594 , \5593 );
xor \U$5500 ( \5595 , \5588 , \5594 );
buf \U$5501 ( \5596 , \5595 );
buf \U$5502 ( \5597 , \5596 );
xor \U$5503 ( \5598 , \5449 , \5597 );
xor \U$5504 ( \5599 , \4968 , \5104 );
and \U$5505 ( \5600 , \5599 , \5111 );
and \U$5506 ( \5601 , \4968 , \5104 );
or \U$5507 ( \5602 , \5600 , \5601 );
buf \U$5508 ( \5603 , \5602 );
buf \U$5509 ( \5604 , \5603 );
xor \U$5510 ( \5605 , \5598 , \5604 );
buf \U$5511 ( \5606 , \5605 );
buf \U$5512 ( \5607 , \5606 );
xor \U$5513 ( \5608 , \4955 , \4961 );
and \U$5514 ( \5609 , \5608 , \5114 );
and \U$5515 ( \5610 , \4955 , \4961 );
or \U$5516 ( \5611 , \5609 , \5610 );
buf \U$5517 ( \5612 , \5611 );
buf \U$5518 ( \5613 , \5612 );
or \U$5519 ( \5614 , \5607 , \5613 );
buf \U$5520 ( \5615 , \5614 );
buf \U$5521 ( \5616 , \5615 );
nand \U$5522 ( \5617 , \5136 , \5616 );
buf \U$5523 ( \5618 , \5617 );
buf \U$5524 ( \5619 , \5618 );
buf \U$5525 ( \5620 , \5155 );
not \U$5526 ( \5621 , \5620 );
buf \U$5527 ( \5622 , \5146 );
not \U$5528 ( \5623 , \5622 );
buf \U$5529 ( \5624 , \618 );
not \U$5530 ( \5625 , \5624 );
or \U$5531 ( \5626 , \5623 , \5625 );
xnor \U$5532 ( \5627 , RIc0d9ec8_87, RIc0d7858_5);
buf \U$5533 ( \5628 , \5627 );
not \U$5534 ( \5629 , \5628 );
buf \U$5535 ( \5630 , \816 );
nand \U$5536 ( \5631 , \5629 , \5630 );
buf \U$5537 ( \5632 , \5631 );
buf \U$5538 ( \5633 , \5632 );
nand \U$5539 ( \5634 , \5626 , \5633 );
buf \U$5540 ( \5635 , \5634 );
buf \U$5541 ( \5636 , \5635 );
not \U$5542 ( \5637 , \5636 );
and \U$5543 ( \5638 , \5621 , \5637 );
buf \U$5544 ( \5639 , \5635 );
buf \U$5545 ( \5640 , \5155 );
and \U$5546 ( \5641 , \5639 , \5640 );
nor \U$5547 ( \5642 , \5638 , \5641 );
buf \U$5548 ( \5643 , \5642 );
buf \U$5549 ( \5644 , \5643 );
not \U$5550 ( \5645 , \5644 );
buf \U$5551 ( \5646 , \5418 );
not \U$5552 ( \5647 , \5646 );
buf \U$5553 ( \5648 , \5402 );
not \U$5554 ( \5649 , \5648 );
or \U$5555 ( \5650 , \5647 , \5649 );
buf \U$5556 ( \5651 , \5402 );
buf \U$5557 ( \5652 , \5418 );
or \U$5558 ( \5653 , \5651 , \5652 );
buf \U$5559 ( \5654 , \5438 );
nand \U$5560 ( \5655 , \5653 , \5654 );
buf \U$5561 ( \5656 , \5655 );
buf \U$5562 ( \5657 , \5656 );
nand \U$5563 ( \5658 , \5650 , \5657 );
buf \U$5564 ( \5659 , \5658 );
buf \U$5565 ( \5660 , \5659 );
not \U$5566 ( \5661 , \5660 );
or \U$5567 ( \5662 , \5645 , \5661 );
buf \U$5568 ( \5663 , \5659 );
buf \U$5569 ( \5664 , \5643 );
or \U$5570 ( \5665 , \5663 , \5664 );
nand \U$5571 ( \5666 , \5662 , \5665 );
buf \U$5572 ( \5667 , \5666 );
buf \U$5573 ( \5668 , \5667 );
xor \U$5574 ( \5669 , \5156 , \5162 );
and \U$5575 ( \5670 , \5669 , \5169 );
and \U$5576 ( \5671 , \5156 , \5162 );
or \U$5577 ( \5672 , \5670 , \5671 );
buf \U$5578 ( \5673 , \5672 );
buf \U$5579 ( \5674 , \5673 );
xor \U$5580 ( \5675 , \5668 , \5674 );
buf \U$5581 ( \5676 , \5209 );
not \U$5582 ( \5677 , \5676 );
buf \U$5583 ( \5678 , \5227 );
not \U$5584 ( \5679 , \5678 );
or \U$5585 ( \5680 , \5677 , \5679 );
buf \U$5586 ( \5681 , \5227 );
buf \U$5587 ( \5682 , \5209 );
or \U$5588 ( \5683 , \5681 , \5682 );
buf \U$5589 ( \5684 , \5193 );
nand \U$5590 ( \5685 , \5683 , \5684 );
buf \U$5591 ( \5686 , \5685 );
buf \U$5592 ( \5687 , \5686 );
nand \U$5593 ( \5688 , \5680 , \5687 );
buf \U$5594 ( \5689 , \5688 );
buf \U$5595 ( \5690 , \5689 );
xor \U$5596 ( \5691 , \5675 , \5690 );
buf \U$5597 ( \5692 , \5691 );
buf \U$5598 ( \5693 , \5692 );
xor \U$5599 ( \5694 , \5245 , \5263 );
and \U$5600 ( \5695 , \5694 , \5443 );
and \U$5601 ( \5696 , \5245 , \5263 );
or \U$5602 ( \5697 , \5695 , \5696 );
buf \U$5603 ( \5698 , \5697 );
buf \U$5604 ( \5699 , \5698 );
xor \U$5605 ( \5700 , \5693 , \5699 );
buf \U$5606 ( \5701 , \5476 );
not \U$5607 ( \5702 , \5701 );
buf \U$5608 ( \5703 , \5702 );
buf \U$5609 ( \5704 , \5703 );
not \U$5610 ( \5705 , \5704 );
buf \U$5611 ( \5706 , \5492 );
not \U$5612 ( \5707 , \5706 );
or \U$5613 ( \5708 , \5705 , \5707 );
buf \U$5614 ( \5709 , \5492 );
buf \U$5615 ( \5710 , \5703 );
or \U$5616 ( \5711 , \5709 , \5710 );
buf \U$5617 ( \5712 , \5505 );
nand \U$5618 ( \5713 , \5711 , \5712 );
buf \U$5619 ( \5714 , \5713 );
buf \U$5620 ( \5715 , \5714 );
nand \U$5621 ( \5716 , \5708 , \5715 );
buf \U$5622 ( \5717 , \5716 );
buf \U$5623 ( \5718 , \5717 );
xor \U$5624 ( \5719 , \5340 , \5358 );
and \U$5625 ( \5720 , \5719 , \5382 );
and \U$5626 ( \5721 , \5340 , \5358 );
or \U$5627 ( \5722 , \5720 , \5721 );
buf \U$5628 ( \5723 , \5722 );
buf \U$5629 ( \5724 , \5723 );
xor \U$5630 ( \5725 , \5718 , \5724 );
buf \U$5631 ( \5726 , \5558 );
not \U$5632 ( \5727 , \5726 );
buf \U$5633 ( \5728 , \5542 );
not \U$5634 ( \5729 , \5728 );
or \U$5635 ( \5730 , \5727 , \5729 );
buf \U$5636 ( \5731 , \5542 );
buf \U$5637 ( \5732 , \5558 );
or \U$5638 ( \5733 , \5731 , \5732 );
buf \U$5639 ( \5734 , \5520 );
nand \U$5640 ( \5735 , \5733 , \5734 );
buf \U$5641 ( \5736 , \5735 );
buf \U$5642 ( \5737 , \5736 );
nand \U$5643 ( \5738 , \5730 , \5737 );
buf \U$5644 ( \5739 , \5738 );
buf \U$5645 ( \5740 , \5739 );
xor \U$5646 ( \5741 , \5725 , \5740 );
buf \U$5647 ( \5742 , \5741 );
buf \U$5648 ( \5743 , \5742 );
xor \U$5649 ( \5744 , \5472 , \5507 );
and \U$5650 ( \5745 , \5744 , \5568 );
and \U$5651 ( \5746 , \5472 , \5507 );
or \U$5652 ( \5747 , \5745 , \5746 );
buf \U$5653 ( \5748 , \5747 );
buf \U$5654 ( \5749 , \5748 );
xor \U$5655 ( \5750 , \5743 , \5749 );
xor \U$5656 ( \5751 , \5323 , \5385 );
and \U$5657 ( \5752 , \5751 , \5440 );
and \U$5658 ( \5753 , \5323 , \5385 );
or \U$5659 ( \5754 , \5752 , \5753 );
buf \U$5660 ( \5755 , \5754 );
buf \U$5661 ( \5756 , \5755 );
xor \U$5662 ( \5757 , \5750 , \5756 );
buf \U$5663 ( \5758 , \5757 );
buf \U$5664 ( \5759 , \5758 );
xor \U$5665 ( \5760 , \5700 , \5759 );
buf \U$5666 ( \5761 , \5760 );
buf \U$5667 ( \5762 , \5761 );
xor \U$5668 ( \5763 , \5455 , \5587 );
and \U$5669 ( \5764 , \5763 , \5594 );
and \U$5670 ( \5765 , \5455 , \5587 );
or \U$5671 ( \5766 , \5764 , \5765 );
buf \U$5672 ( \5767 , \5766 );
buf \U$5673 ( \5768 , \5767 );
xor \U$5674 ( \5769 , \5762 , \5768 );
xor \U$5675 ( \5770 , \5571 , \5577 );
and \U$5676 ( \5771 , \5770 , \5584 );
and \U$5677 ( \5772 , \5571 , \5577 );
or \U$5678 ( \5773 , \5771 , \5772 );
buf \U$5679 ( \5774 , \5773 );
buf \U$5680 ( \5775 , \5774 );
xor \U$5681 ( \5776 , \5281 , \5298 );
and \U$5682 ( \5777 , \5776 , \5320 );
and \U$5683 ( \5778 , \5281 , \5298 );
or \U$5684 ( \5779 , \5777 , \5778 );
buf \U$5685 ( \5780 , \5779 );
buf \U$5686 ( \5781 , \5780 );
and \U$5687 ( \5782 , \4975 , \4976 );
buf \U$5688 ( \5783 , \5782 );
buf \U$5689 ( \5784 , \5783 );
buf \U$5690 ( \5785 , \5274 );
not \U$5691 ( \5786 , \5785 );
buf \U$5692 ( \5787 , \678 );
not \U$5693 ( \5788 , \5787 );
or \U$5694 ( \5789 , \5786 , \5788 );
buf \U$5695 ( \5790 , \686 );
buf \U$5696 ( \5791 , RIc0d81b8_25);
buf \U$5697 ( \5792 , RIc0d9568_67);
xor \U$5698 ( \5793 , \5791 , \5792 );
buf \U$5699 ( \5794 , \5793 );
buf \U$5700 ( \5795 , \5794 );
nand \U$5701 ( \5796 , \5790 , \5795 );
buf \U$5702 ( \5797 , \5796 );
buf \U$5703 ( \5798 , \5797 );
nand \U$5704 ( \5799 , \5789 , \5798 );
buf \U$5705 ( \5800 , \5799 );
buf \U$5706 ( \5801 , \5800 );
xor \U$5707 ( \5802 , \5784 , \5801 );
buf \U$5708 ( \5803 , \5432 );
not \U$5709 ( \5804 , \5803 );
buf \U$5710 ( \5805 , \2726 );
not \U$5711 ( \5806 , \5805 );
or \U$5712 ( \5807 , \5804 , \5806 );
buf \U$5713 ( \5808 , \1933 );
buf \U$5714 ( \5809 , RIc0d7678_1);
buf \U$5715 ( \5810 , RIc0da0a8_91);
xor \U$5716 ( \5811 , \5809 , \5810 );
buf \U$5717 ( \5812 , \5811 );
buf \U$5718 ( \5813 , \5812 );
nand \U$5719 ( \5814 , \5808 , \5813 );
buf \U$5720 ( \5815 , \5814 );
buf \U$5721 ( \5816 , \5815 );
nand \U$5722 ( \5817 , \5807 , \5816 );
buf \U$5723 ( \5818 , \5817 );
buf \U$5724 ( \5819 , \5818 );
xor \U$5725 ( \5820 , \5802 , \5819 );
buf \U$5726 ( \5821 , \5820 );
buf \U$5727 ( \5822 , \5821 );
xor \U$5728 ( \5823 , \5781 , \5822 );
buf \U$5729 ( \5824 , \2769 );
buf \U$5730 ( \5825 , \5534 );
or \U$5731 ( \5826 , \5824 , \5825 );
buf \U$5732 ( \5827 , \2775 );
buf \U$5733 ( \5828 , RIc0d7b28_11);
buf \U$5734 ( \5829 , RIc0d9bf8_81);
xor \U$5735 ( \5830 , \5828 , \5829 );
buf \U$5736 ( \5831 , \5830 );
buf \U$5737 ( \5832 , \5831 );
not \U$5738 ( \5833 , \5832 );
buf \U$5739 ( \5834 , \5833 );
buf \U$5740 ( \5835 , \5834 );
or \U$5741 ( \5836 , \5827 , \5835 );
nand \U$5742 ( \5837 , \5826 , \5836 );
buf \U$5743 ( \5838 , \5837 );
buf \U$5744 ( \5839 , \5377 );
not \U$5745 ( \5840 , \5839 );
buf \U$5746 ( \5841 , \5840 );
buf \U$5747 ( \5842 , \5841 );
not \U$5748 ( \5843 , \5842 );
buf \U$5749 ( \5844 , \842 );
not \U$5750 ( \5845 , \5844 );
or \U$5751 ( \5846 , \5843 , \5845 );
buf \U$5752 ( \5847 , \846 );
buf \U$5753 ( \5848 , RIc0d9fb8_89);
buf \U$5754 ( \5849 , RIc0d7768_3);
and \U$5755 ( \5850 , \5848 , \5849 );
not \U$5756 ( \5851 , \5848 );
buf \U$5757 ( \5852 , \304 );
and \U$5758 ( \5853 , \5851 , \5852 );
nor \U$5759 ( \5854 , \5850 , \5853 );
buf \U$5760 ( \5855 , \5854 );
buf \U$5761 ( \5856 , \5855 );
nand \U$5762 ( \5857 , \5847 , \5856 );
buf \U$5763 ( \5858 , \5857 );
buf \U$5764 ( \5859 , \5858 );
nand \U$5765 ( \5860 , \5846 , \5859 );
buf \U$5766 ( \5861 , \5860 );
xor \U$5767 ( \5862 , \5838 , \5861 );
buf \U$5768 ( \5863 , \5552 );
not \U$5769 ( \5864 , \5863 );
buf \U$5770 ( \5865 , \1021 );
not \U$5771 ( \5866 , \5865 );
or \U$5772 ( \5867 , \5864 , \5866 );
buf \U$5773 ( \5868 , \3985 );
buf \U$5774 ( \5869 , RIc0d7c18_13);
buf \U$5775 ( \5870 , RIc0d9b08_79);
xor \U$5776 ( \5871 , \5869 , \5870 );
buf \U$5777 ( \5872 , \5871 );
buf \U$5778 ( \5873 , \5872 );
nand \U$5779 ( \5874 , \5868 , \5873 );
buf \U$5780 ( \5875 , \5874 );
buf \U$5781 ( \5876 , \5875 );
nand \U$5782 ( \5877 , \5867 , \5876 );
buf \U$5783 ( \5878 , \5877 );
xor \U$5784 ( \5879 , \5862 , \5878 );
buf \U$5785 ( \5880 , \5879 );
xor \U$5786 ( \5881 , \5823 , \5880 );
buf \U$5787 ( \5882 , \5881 );
buf \U$5788 ( \5883 , \5882 );
buf \U$5789 ( \5884 , \4008 );
not \U$5790 ( \5885 , \5884 );
buf \U$5791 ( \5886 , \5885 );
buf \U$5792 ( \5887 , \5886 );
not \U$5793 ( \5888 , \5887 );
buf \U$5794 ( \5889 , \473 );
not \U$5795 ( \5890 , \5889 );
or \U$5796 ( \5891 , \5888 , \5890 );
buf \U$5797 ( \5892 , RIc0da198_93);
nand \U$5798 ( \5893 , \5891 , \5892 );
buf \U$5799 ( \5894 , \5893 );
buf \U$5800 ( \5895 , \5412 );
not \U$5801 ( \5896 , \5895 );
buf \U$5802 ( \5897 , \3781 );
not \U$5803 ( \5898 , \5897 );
or \U$5804 ( \5899 , \5896 , \5898 );
buf \U$5805 ( \5900 , \1229 );
buf \U$5806 ( \5901 , RIc0d9478_65);
buf \U$5807 ( \5902 , RIc0d82a8_27);
xor \U$5808 ( \5903 , \5901 , \5902 );
buf \U$5809 ( \5904 , \5903 );
buf \U$5810 ( \5905 , \5904 );
nand \U$5811 ( \5906 , \5900 , \5905 );
buf \U$5812 ( \5907 , \5906 );
buf \U$5813 ( \5908 , \5907 );
nand \U$5814 ( \5909 , \5899 , \5908 );
buf \U$5815 ( \5910 , \5909 );
buf \U$5816 ( \5911 , \5910 );
not \U$5817 ( \5912 , \5911 );
buf \U$5818 ( \5913 , \5912 );
and \U$5819 ( \5914 , \5894 , \5913 );
not \U$5820 ( \5915 , \5894 );
and \U$5821 ( \5916 , \5915 , \5910 );
or \U$5822 ( \5917 , \5914 , \5916 );
buf \U$5823 ( \5918 , \5917 );
buf \U$5824 ( \5919 , \5291 );
not \U$5825 ( \5920 , \5919 );
buf \U$5826 ( \5921 , \2269 );
not \U$5827 ( \5922 , \5921 );
or \U$5828 ( \5923 , \5920 , \5922 );
buf \U$5829 ( \5924 , \2927 );
buf \U$5830 ( \5925 , RIc0d7fd8_21);
buf \U$5831 ( \5926 , RIc0d9748_71);
xor \U$5832 ( \5927 , \5925 , \5926 );
buf \U$5833 ( \5928 , \5927 );
buf \U$5834 ( \5929 , \5928 );
nand \U$5835 ( \5930 , \5924 , \5929 );
buf \U$5836 ( \5931 , \5930 );
buf \U$5837 ( \5932 , \5931 );
nand \U$5838 ( \5933 , \5923 , \5932 );
buf \U$5839 ( \5934 , \5933 );
buf \U$5840 ( \5935 , \5934 );
and \U$5841 ( \5936 , \5918 , \5935 );
not \U$5842 ( \5937 , \5918 );
buf \U$5843 ( \5938 , \5934 );
not \U$5844 ( \5939 , \5938 );
buf \U$5845 ( \5940 , \5939 );
buf \U$5846 ( \5941 , \5940 );
and \U$5847 ( \5942 , \5937 , \5941 );
nor \U$5848 ( \5943 , \5936 , \5942 );
buf \U$5849 ( \5944 , \5943 );
buf \U$5850 ( \5945 , \5944 );
buf \U$5851 ( \5946 , \5333 );
not \U$5852 ( \5947 , \5946 );
buf \U$5853 ( \5948 , \2359 );
not \U$5854 ( \5949 , \5948 );
or \U$5855 ( \5950 , \5947 , \5949 );
buf \U$5856 ( \5951 , \1143 );
buf \U$5857 ( \5952 , RIc0d7df8_17);
buf \U$5858 ( \5953 , RIc0d9928_75);
xor \U$5859 ( \5954 , \5952 , \5953 );
buf \U$5860 ( \5955 , \5954 );
buf \U$5861 ( \5956 , \5955 );
nand \U$5862 ( \5957 , \5951 , \5956 );
buf \U$5863 ( \5958 , \5957 );
buf \U$5864 ( \5959 , \5958 );
nand \U$5865 ( \5960 , \5950 , \5959 );
buf \U$5866 ( \5961 , \5960 );
buf \U$5867 ( \5962 , \5961 );
buf \U$5868 ( \5963 , \5516 );
not \U$5869 ( \5964 , \5963 );
buf \U$5870 ( \5965 , \5964 );
buf \U$5871 ( \5966 , \5965 );
not \U$5872 ( \5967 , \5966 );
buf \U$5873 ( \5968 , \2088 );
not \U$5874 ( \5969 , \5968 );
or \U$5875 ( \5970 , \5967 , \5969 );
buf \U$5876 ( \5971 , \1050 );
buf \U$5877 ( \5972 , RIc0d7a38_9);
and \U$5878 ( \5973 , \5971 , \5972 );
buf \U$5879 ( \5974 , RIc0d7a38_9);
not \U$5880 ( \5975 , \5974 );
buf \U$5881 ( \5976 , \5975 );
buf \U$5882 ( \5977 , \5976 );
buf \U$5883 ( \5978 , RIc0d9ce8_83);
and \U$5884 ( \5979 , \5977 , \5978 );
nor \U$5885 ( \5980 , \5973 , \5979 );
buf \U$5886 ( \5981 , \5980 );
buf \U$5887 ( \5982 , \5981 );
not \U$5888 ( \5983 , \5982 );
buf \U$5889 ( \5984 , \993 );
nand \U$5890 ( \5985 , \5983 , \5984 );
buf \U$5891 ( \5986 , \5985 );
buf \U$5892 ( \5987 , \5986 );
nand \U$5893 ( \5988 , \5970 , \5987 );
buf \U$5894 ( \5989 , \5988 );
buf \U$5895 ( \5990 , \5989 );
xor \U$5896 ( \5991 , \5962 , \5990 );
buf \U$5897 ( \5992 , \1435 );
buf \U$5898 ( \5993 , \5349 );
or \U$5899 ( \5994 , \5992 , \5993 );
buf \U$5900 ( \5995 , \1193 );
buf \U$5901 ( \5996 , RIc0d7d08_15);
buf \U$5902 ( \5997 , RIc0d9a18_77);
xnor \U$5903 ( \5998 , \5996 , \5997 );
buf \U$5904 ( \5999 , \5998 );
buf \U$5905 ( \6000 , \5999 );
or \U$5906 ( \6001 , \5995 , \6000 );
nand \U$5907 ( \6002 , \5994 , \6001 );
buf \U$5908 ( \6003 , \6002 );
buf \U$5909 ( \6004 , \6003 );
xor \U$5910 ( \6005 , \5991 , \6004 );
buf \U$5911 ( \6006 , \6005 );
buf \U$5912 ( \6007 , \6006 );
xor \U$5913 ( \6008 , \5945 , \6007 );
buf \U$5914 ( \6009 , \5396 );
not \U$5915 ( \6010 , \6009 );
buf \U$5916 ( \6011 , \1677 );
not \U$5917 ( \6012 , \6011 );
or \U$5918 ( \6013 , \6010 , \6012 );
buf \U$5919 ( \6014 , \2882 );
buf \U$5920 ( \6015 , RIc0d7ee8_19);
buf \U$5921 ( \6016 , RIc0d9838_73);
xor \U$5922 ( \6017 , \6015 , \6016 );
buf \U$5923 ( \6018 , \6017 );
buf \U$5924 ( \6019 , \6018 );
nand \U$5925 ( \6020 , \6014 , \6019 );
buf \U$5926 ( \6021 , \6020 );
buf \U$5927 ( \6022 , \6021 );
nand \U$5928 ( \6023 , \6013 , \6022 );
buf \U$5929 ( \6024 , \6023 );
buf \U$5930 ( \6025 , \5313 );
not \U$5931 ( \6026 , \6025 );
buf \U$5932 ( \6027 , \3295 );
not \U$5933 ( \6028 , \6027 );
buf \U$5934 ( \6029 , \6028 );
buf \U$5935 ( \6030 , \6029 );
not \U$5936 ( \6031 , \6030 );
or \U$5937 ( \6032 , \6026 , \6031 );
buf \U$5938 ( \6033 , \921 );
buf \U$5939 ( \6034 , RIc0d7948_7);
buf \U$5940 ( \6035 , RIc0d9dd8_85);
xor \U$5941 ( \6036 , \6034 , \6035 );
buf \U$5942 ( \6037 , \6036 );
buf \U$5943 ( \6038 , \6037 );
nand \U$5944 ( \6039 , \6033 , \6038 );
buf \U$5945 ( \6040 , \6039 );
buf \U$5946 ( \6041 , \6040 );
nand \U$5947 ( \6042 , \6032 , \6041 );
buf \U$5948 ( \6043 , \6042 );
buf \U$5949 ( \6044 , \6043 );
buf \U$5950 ( \6045 , \5486 );
not \U$5951 ( \6046 , \6045 );
buf \U$5952 ( \6047 , \864 );
not \U$5953 ( \6048 , \6047 );
or \U$5954 ( \6049 , \6046 , \6048 );
buf \U$5955 ( \6050 , RIc0d80c8_23);
buf \U$5956 ( \6051 , RIc0d9658_69);
xnor \U$5957 ( \6052 , \6050 , \6051 );
buf \U$5958 ( \6053 , \6052 );
buf \U$5959 ( \6054 , \6053 );
not \U$5960 ( \6055 , \6054 );
buf \U$5961 ( \6056 , \284 );
nand \U$5962 ( \6057 , \6055 , \6056 );
buf \U$5963 ( \6058 , \6057 );
buf \U$5964 ( \6059 , \6058 );
nand \U$5965 ( \6060 , \6049 , \6059 );
buf \U$5966 ( \6061 , \6060 );
buf \U$5967 ( \6062 , \6061 );
xor \U$5968 ( \6063 , \6044 , \6062 );
buf \U$5969 ( \6064 , \6063 );
xor \U$5970 ( \6065 , \6024 , \6064 );
buf \U$5971 ( \6066 , \6065 );
xor \U$5972 ( \6067 , \6008 , \6066 );
buf \U$5973 ( \6068 , \6067 );
buf \U$5974 ( \6069 , \6068 );
xor \U$5975 ( \6070 , \5883 , \6069 );
xor \U$5976 ( \6071 , \5172 , \5178 );
and \U$5977 ( \6072 , \6071 , \5229 );
and \U$5978 ( \6073 , \5172 , \5178 );
or \U$5979 ( \6074 , \6072 , \6073 );
buf \U$5980 ( \6075 , \6074 );
buf \U$5981 ( \6076 , \6075 );
xor \U$5982 ( \6077 , \6070 , \6076 );
buf \U$5983 ( \6078 , \6077 );
buf \U$5984 ( \6079 , \6078 );
xor \U$5985 ( \6080 , \5775 , \6079 );
xor \U$5986 ( \6081 , \5232 , \5238 );
and \U$5987 ( \6082 , \6081 , \5446 );
and \U$5988 ( \6083 , \5232 , \5238 );
or \U$5989 ( \6084 , \6082 , \6083 );
buf \U$5990 ( \6085 , \6084 );
buf \U$5991 ( \6086 , \6085 );
xor \U$5992 ( \6087 , \6080 , \6086 );
buf \U$5993 ( \6088 , \6087 );
buf \U$5994 ( \6089 , \6088 );
xor \U$5995 ( \6090 , \5769 , \6089 );
buf \U$5996 ( \6091 , \6090 );
buf \U$5997 ( \6092 , \6091 );
xor \U$5998 ( \6093 , \5449 , \5597 );
and \U$5999 ( \6094 , \6093 , \5604 );
and \U$6000 ( \6095 , \5449 , \5597 );
or \U$6001 ( \6096 , \6094 , \6095 );
buf \U$6002 ( \6097 , \6096 );
buf \U$6003 ( \6098 , \6097 );
nor \U$6004 ( \6099 , \6092 , \6098 );
buf \U$6005 ( \6100 , \6099 );
buf \U$6006 ( \6101 , \6100 );
nor \U$6007 ( \6102 , \5619 , \6101 );
buf \U$6008 ( \6103 , \6102 );
buf \U$6009 ( \6104 , \6103 );
buf \U$6010 ( \6105 , \5155 );
not \U$6011 ( \6106 , \6105 );
buf \U$6012 ( \6107 , \5635 );
not \U$6013 ( \6108 , \6107 );
buf \U$6014 ( \6109 , \6108 );
buf \U$6015 ( \6110 , \6109 );
not \U$6016 ( \6111 , \6110 );
or \U$6017 ( \6112 , \6106 , \6111 );
buf \U$6018 ( \6113 , \5659 );
nand \U$6019 ( \6114 , \6112 , \6113 );
buf \U$6020 ( \6115 , \6114 );
buf \U$6021 ( \6116 , \6115 );
buf \U$6022 ( \6117 , \5152 );
buf \U$6023 ( \6118 , \5635 );
nand \U$6024 ( \6119 , \6117 , \6118 );
buf \U$6025 ( \6120 , \6119 );
buf \U$6026 ( \6121 , \6120 );
nand \U$6027 ( \6122 , \6116 , \6121 );
buf \U$6028 ( \6123 , \6122 );
buf \U$6029 ( \6124 , \6123 );
buf \U$6030 ( \6125 , \5999 );
not \U$6031 ( \6126 , \6125 );
buf \U$6032 ( \6127 , \6126 );
buf \U$6033 ( \6128 , \6127 );
not \U$6034 ( \6129 , \6128 );
buf \U$6035 ( \6130 , \1432 );
not \U$6036 ( \6131 , \6130 );
or \U$6037 ( \6132 , \6129 , \6131 );
buf \U$6038 ( \6133 , RIc0d7c90_14);
buf \U$6039 ( \6134 , RIc0d9a18_77);
xnor \U$6040 ( \6135 , \6133 , \6134 );
buf \U$6041 ( \6136 , \6135 );
buf \U$6042 ( \6137 , \6136 );
not \U$6043 ( \6138 , \6137 );
buf \U$6044 ( \6139 , \1193 );
not \U$6045 ( \6140 , \6139 );
buf \U$6046 ( \6141 , \6140 );
buf \U$6047 ( \6142 , \6141 );
nand \U$6048 ( \6143 , \6138 , \6142 );
buf \U$6049 ( \6144 , \6143 );
buf \U$6050 ( \6145 , \6144 );
nand \U$6051 ( \6146 , \6132 , \6145 );
buf \U$6052 ( \6147 , \6146 );
buf \U$6053 ( \6148 , \6037 );
not \U$6054 ( \6149 , \6148 );
buf \U$6055 ( \6150 , \5305 );
not \U$6056 ( \6151 , \6150 );
or \U$6057 ( \6152 , \6149 , \6151 );
buf \U$6058 ( \6153 , \2960 );
buf \U$6059 ( \6154 , RIc0d78d0_6);
buf \U$6060 ( \6155 , RIc0d9dd8_85);
xor \U$6061 ( \6156 , \6154 , \6155 );
buf \U$6062 ( \6157 , \6156 );
buf \U$6063 ( \6158 , \6157 );
nand \U$6064 ( \6159 , \6153 , \6158 );
buf \U$6065 ( \6160 , \6159 );
buf \U$6066 ( \6161 , \6160 );
nand \U$6067 ( \6162 , \6152 , \6161 );
buf \U$6068 ( \6163 , \6162 );
xor \U$6069 ( \6164 , \6147 , \6163 );
buf \U$6070 ( \6165 , \5812 );
not \U$6071 ( \6166 , \6165 );
buf \U$6072 ( \6167 , \2535 );
not \U$6073 ( \6168 , \6167 );
or \U$6074 ( \6169 , \6166 , \6168 );
buf \U$6075 ( \6170 , \533 );
buf \U$6076 ( \6171 , RIc0da0a8_91);
nand \U$6077 ( \6172 , \6170 , \6171 );
buf \U$6078 ( \6173 , \6172 );
buf \U$6079 ( \6174 , \6173 );
nand \U$6080 ( \6175 , \6169 , \6174 );
buf \U$6081 ( \6176 , \6175 );
not \U$6082 ( \6177 , \6176 );
xor \U$6083 ( \6178 , \6164 , \6177 );
buf \U$6084 ( \6179 , \6178 );
xor \U$6085 ( \6180 , \6124 , \6179 );
xor \U$6086 ( \6181 , \5718 , \5724 );
and \U$6087 ( \6182 , \6181 , \5740 );
and \U$6088 ( \6183 , \5718 , \5724 );
or \U$6089 ( \6184 , \6182 , \6183 );
buf \U$6090 ( \6185 , \6184 );
buf \U$6091 ( \6186 , \6185 );
xor \U$6092 ( \6187 , \6180 , \6186 );
buf \U$6093 ( \6188 , \6187 );
buf \U$6094 ( \6189 , \6188 );
xor \U$6095 ( \6190 , \5743 , \5749 );
and \U$6096 ( \6191 , \6190 , \5756 );
and \U$6097 ( \6192 , \5743 , \5749 );
or \U$6098 ( \6193 , \6191 , \6192 );
buf \U$6099 ( \6194 , \6193 );
buf \U$6100 ( \6195 , \6194 );
xor \U$6101 ( \6196 , \6189 , \6195 );
xor \U$6102 ( \6197 , \5781 , \5822 );
and \U$6103 ( \6198 , \6197 , \5880 );
and \U$6104 ( \6199 , \5781 , \5822 );
or \U$6105 ( \6200 , \6198 , \6199 );
buf \U$6106 ( \6201 , \6200 );
buf \U$6107 ( \6202 , \6201 );
xor \U$6108 ( \6203 , \5784 , \5801 );
and \U$6109 ( \6204 , \6203 , \5819 );
and \U$6110 ( \6205 , \5784 , \5801 );
or \U$6111 ( \6206 , \6204 , \6205 );
buf \U$6112 ( \6207 , \6206 );
buf \U$6113 ( \6208 , \6207 );
buf \U$6114 ( \6209 , \5913 );
not \U$6115 ( \6210 , \6209 );
buf \U$6116 ( \6211 , \5940 );
not \U$6117 ( \6212 , \6211 );
or \U$6118 ( \6213 , \6210 , \6212 );
buf \U$6119 ( \6214 , \5894 );
nand \U$6120 ( \6215 , \6213 , \6214 );
buf \U$6121 ( \6216 , \6215 );
buf \U$6122 ( \6217 , \6216 );
buf \U$6123 ( \6218 , \5934 );
buf \U$6124 ( \6219 , \5910 );
nand \U$6125 ( \6220 , \6218 , \6219 );
buf \U$6126 ( \6221 , \6220 );
buf \U$6127 ( \6222 , \6221 );
nand \U$6128 ( \6223 , \6217 , \6222 );
buf \U$6129 ( \6224 , \6223 );
buf \U$6130 ( \6225 , \6224 );
xor \U$6131 ( \6226 , \6208 , \6225 );
buf \U$6132 ( \6227 , \5878 );
not \U$6133 ( \6228 , \6227 );
buf \U$6134 ( \6229 , \5861 );
not \U$6135 ( \6230 , \6229 );
or \U$6136 ( \6231 , \6228 , \6230 );
buf \U$6137 ( \6232 , \5861 );
buf \U$6138 ( \6233 , \5878 );
or \U$6139 ( \6234 , \6232 , \6233 );
buf \U$6140 ( \6235 , \5838 );
nand \U$6141 ( \6236 , \6234 , \6235 );
buf \U$6142 ( \6237 , \6236 );
buf \U$6143 ( \6238 , \6237 );
nand \U$6144 ( \6239 , \6231 , \6238 );
buf \U$6145 ( \6240 , \6239 );
buf \U$6146 ( \6241 , \6240 );
xor \U$6147 ( \6242 , \6226 , \6241 );
buf \U$6148 ( \6243 , \6242 );
buf \U$6149 ( \6244 , \6243 );
xor \U$6150 ( \6245 , \6202 , \6244 );
buf \U$6151 ( \6246 , \6043 );
not \U$6152 ( \6247 , \6246 );
buf \U$6153 ( \6248 , \6061 );
not \U$6154 ( \6249 , \6248 );
or \U$6155 ( \6250 , \6247 , \6249 );
buf \U$6156 ( \6251 , \6061 );
buf \U$6157 ( \6252 , \6043 );
or \U$6158 ( \6253 , \6251 , \6252 );
buf \U$6159 ( \6254 , \6024 );
nand \U$6160 ( \6255 , \6253 , \6254 );
buf \U$6161 ( \6256 , \6255 );
buf \U$6162 ( \6257 , \6256 );
nand \U$6163 ( \6258 , \6250 , \6257 );
buf \U$6164 ( \6259 , \6258 );
buf \U$6165 ( \6260 , \6259 );
xor \U$6166 ( \6261 , \5962 , \5990 );
and \U$6167 ( \6262 , \6261 , \6004 );
and \U$6168 ( \6263 , \5962 , \5990 );
or \U$6169 ( \6264 , \6262 , \6263 );
buf \U$6170 ( \6265 , \6264 );
buf \U$6171 ( \6266 , \6265 );
xor \U$6172 ( \6267 , \6260 , \6266 );
buf \U$6173 ( \6268 , \2607 );
not \U$6174 ( \6269 , \6268 );
buf \U$6175 ( \6270 , \6269 );
buf \U$6176 ( \6271 , \6270 );
buf \U$6177 ( \6272 , \5627 );
or \U$6178 ( \6273 , \6271 , \6272 );
buf \U$6179 ( \6274 , \819 );
buf \U$6180 ( \6275 , RIc0d77e0_4);
buf \U$6181 ( \6276 , RIc0d9ec8_87);
xnor \U$6182 ( \6277 , \6275 , \6276 );
buf \U$6183 ( \6278 , \6277 );
buf \U$6184 ( \6279 , \6278 );
or \U$6185 ( \6280 , \6274 , \6279 );
nand \U$6186 ( \6281 , \6273 , \6280 );
buf \U$6187 ( \6282 , \6281 );
buf \U$6188 ( \6283 , \6018 );
not \U$6189 ( \6284 , \6283 );
buf \U$6190 ( \6285 , \1677 );
not \U$6191 ( \6286 , \6285 );
or \U$6192 ( \6287 , \6284 , \6286 );
buf \U$6193 ( \6288 , \792 );
buf \U$6194 ( \6289 , RIc0d7e70_18);
buf \U$6195 ( \6290 , RIc0d9838_73);
xor \U$6196 ( \6291 , \6289 , \6290 );
buf \U$6197 ( \6292 , \6291 );
buf \U$6198 ( \6293 , \6292 );
nand \U$6199 ( \6294 , \6288 , \6293 );
buf \U$6200 ( \6295 , \6294 );
buf \U$6201 ( \6296 , \6295 );
nand \U$6202 ( \6297 , \6287 , \6296 );
buf \U$6203 ( \6298 , \6297 );
buf \U$6204 ( \6299 , \5872 );
not \U$6205 ( \6300 , \6299 );
buf \U$6206 ( \6301 , \1021 );
not \U$6207 ( \6302 , \6301 );
or \U$6208 ( \6303 , \6300 , \6302 );
buf \U$6209 ( \6304 , \3985 );
buf \U$6210 ( \6305 , RIc0d7ba0_12);
buf \U$6211 ( \6306 , RIc0d9b08_79);
xor \U$6212 ( \6307 , \6305 , \6306 );
buf \U$6213 ( \6308 , \6307 );
buf \U$6214 ( \6309 , \6308 );
nand \U$6215 ( \6310 , \6304 , \6309 );
buf \U$6216 ( \6311 , \6310 );
buf \U$6217 ( \6312 , \6311 );
nand \U$6218 ( \6313 , \6303 , \6312 );
buf \U$6219 ( \6314 , \6313 );
xor \U$6220 ( \6315 , \6298 , \6314 );
xor \U$6221 ( \6316 , \6282 , \6315 );
buf \U$6222 ( \6317 , \6316 );
xor \U$6223 ( \6318 , \6267 , \6317 );
buf \U$6224 ( \6319 , \6318 );
buf \U$6225 ( \6320 , \6319 );
xor \U$6226 ( \6321 , \6245 , \6320 );
buf \U$6227 ( \6322 , \6321 );
buf \U$6228 ( \6323 , \6322 );
xor \U$6229 ( \6324 , \6196 , \6323 );
buf \U$6230 ( \6325 , \6324 );
buf \U$6231 ( \6326 , \6325 );
not \U$6232 ( \6327 , \6326 );
xor \U$6233 ( \6328 , \5945 , \6007 );
and \U$6234 ( \6329 , \6328 , \6066 );
and \U$6235 ( \6330 , \5945 , \6007 );
or \U$6236 ( \6331 , \6329 , \6330 );
buf \U$6237 ( \6332 , \6331 );
buf \U$6238 ( \6333 , \6332 );
and \U$6239 ( \6334 , \5409 , \5410 );
buf \U$6240 ( \6335 , \6334 );
buf \U$6241 ( \6336 , \6335 );
buf \U$6242 ( \6337 , \5955 );
not \U$6243 ( \6338 , \6337 );
buf \U$6244 ( \6339 , \1556 );
not \U$6245 ( \6340 , \6339 );
or \U$6246 ( \6341 , \6338 , \6340 );
xnor \U$6247 ( \6342 , RIc0d9928_75, RIc0d7d80_16);
buf \U$6248 ( \6343 , \6342 );
not \U$6249 ( \6344 , \6343 );
buf \U$6250 ( \6345 , \1143 );
nand \U$6251 ( \6346 , \6344 , \6345 );
buf \U$6252 ( \6347 , \6346 );
buf \U$6253 ( \6348 , \6347 );
nand \U$6254 ( \6349 , \6341 , \6348 );
buf \U$6255 ( \6350 , \6349 );
buf \U$6256 ( \6351 , \6350 );
xor \U$6257 ( \6352 , \6336 , \6351 );
buf \U$6258 ( \6353 , \861 );
buf \U$6259 ( \6354 , \6053 );
or \U$6260 ( \6355 , \6353 , \6354 );
buf \U$6261 ( \6356 , \1969 );
buf \U$6262 ( \6357 , RIc0d8050_22);
buf \U$6263 ( \6358 , RIc0d9658_69);
xor \U$6264 ( \6359 , \6357 , \6358 );
buf \U$6265 ( \6360 , \6359 );
buf \U$6266 ( \6361 , \6360 );
not \U$6267 ( \6362 , \6361 );
buf \U$6268 ( \6363 , \6362 );
buf \U$6269 ( \6364 , \6363 );
or \U$6270 ( \6365 , \6356 , \6364 );
nand \U$6271 ( \6366 , \6355 , \6365 );
buf \U$6272 ( \6367 , \6366 );
buf \U$6273 ( \6368 , \6367 );
xor \U$6274 ( \6369 , \6352 , \6368 );
buf \U$6275 ( \6370 , \6369 );
buf \U$6276 ( \6371 , \6370 );
buf \U$6277 ( \6372 , \5928 );
not \U$6278 ( \6373 , \6372 );
buf \U$6279 ( \6374 , \1263 );
not \U$6280 ( \6375 , \6374 );
or \U$6281 ( \6376 , \6373 , \6375 );
buf \U$6282 ( \6377 , \1282 );
buf \U$6283 ( \6378 , RIc0d7f60_20);
buf \U$6284 ( \6379 , RIc0d9748_71);
xor \U$6285 ( \6380 , \6378 , \6379 );
buf \U$6286 ( \6381 , \6380 );
buf \U$6287 ( \6382 , \6381 );
nand \U$6288 ( \6383 , \6377 , \6382 );
buf \U$6289 ( \6384 , \6383 );
buf \U$6290 ( \6385 , \6384 );
nand \U$6291 ( \6386 , \6376 , \6385 );
buf \U$6292 ( \6387 , \6386 );
buf \U$6293 ( \6388 , \6387 );
buf \U$6294 ( \6389 , \5855 );
not \U$6295 ( \6390 , \6389 );
buf \U$6296 ( \6391 , \3384 );
not \U$6297 ( \6392 , \6391 );
or \U$6298 ( \6393 , \6390 , \6392 );
and \U$6299 ( \6394 , RIc0d9fb8_89, \352 );
not \U$6300 ( \6395 , RIc0d9fb8_89);
and \U$6301 ( \6396 , \6395 , RIc0d76f0_2);
nor \U$6302 ( \6397 , \6394 , \6396 );
buf \U$6303 ( \6398 , \6397 );
not \U$6304 ( \6399 , \6398 );
buf \U$6305 ( \6400 , \442 );
nand \U$6306 ( \6401 , \6399 , \6400 );
buf \U$6307 ( \6402 , \6401 );
buf \U$6308 ( \6403 , \6402 );
nand \U$6309 ( \6404 , \6393 , \6403 );
buf \U$6310 ( \6405 , \6404 );
buf \U$6311 ( \6406 , \6405 );
xor \U$6312 ( \6407 , \6388 , \6406 );
buf \U$6313 ( \6408 , \1739 );
buf \U$6314 ( \6409 , \5981 );
or \U$6315 ( \6410 , \6408 , \6409 );
buf \U$6316 ( \6411 , \996 );
buf \U$6317 ( \6412 , \1050 );
buf \U$6318 ( \6413 , RIc0d79c0_8);
and \U$6319 ( \6414 , \6412 , \6413 );
buf \U$6320 ( \6415 , \4448 );
buf \U$6321 ( \6416 , RIc0d9ce8_83);
and \U$6322 ( \6417 , \6415 , \6416 );
nor \U$6323 ( \6418 , \6414 , \6417 );
buf \U$6324 ( \6419 , \6418 );
buf \U$6325 ( \6420 , \6419 );
or \U$6326 ( \6421 , \6411 , \6420 );
nand \U$6327 ( \6422 , \6410 , \6421 );
buf \U$6328 ( \6423 , \6422 );
buf \U$6329 ( \6424 , \6423 );
xor \U$6330 ( \6425 , \6407 , \6424 );
buf \U$6331 ( \6426 , \6425 );
buf \U$6332 ( \6427 , \6426 );
xor \U$6333 ( \6428 , \6371 , \6427 );
buf \U$6334 ( \6429 , \1417 );
buf \U$6335 ( \6430 , \5794 );
not \U$6336 ( \6431 , \6430 );
buf \U$6337 ( \6432 , \6431 );
buf \U$6338 ( \6433 , \6432 );
or \U$6339 ( \6434 , \6429 , \6433 );
buf \U$6340 ( \6435 , \686 );
not \U$6341 ( \6436 , \6435 );
buf \U$6342 ( \6437 , \6436 );
buf \U$6343 ( \6438 , \6437 );
buf \U$6344 ( \6439 , RIc0d8140_24);
buf \U$6345 ( \6440 , RIc0d9568_67);
xor \U$6346 ( \6441 , \6439 , \6440 );
buf \U$6347 ( \6442 , \6441 );
buf \U$6348 ( \6443 , \6442 );
not \U$6349 ( \6444 , \6443 );
buf \U$6350 ( \6445 , \6444 );
buf \U$6351 ( \6446 , \6445 );
or \U$6352 ( \6447 , \6438 , \6446 );
nand \U$6353 ( \6448 , \6434 , \6447 );
buf \U$6354 ( \6449 , \6448 );
buf \U$6355 ( \6450 , \5831 );
not \U$6356 ( \6451 , \6450 );
buf \U$6357 ( \6452 , \1064 );
not \U$6358 ( \6453 , \6452 );
or \U$6359 ( \6454 , \6451 , \6453 );
buf \U$6360 ( \6455 , \1078 );
buf \U$6361 ( \6456 , RIc0d7ab0_10);
buf \U$6362 ( \6457 , RIc0d9bf8_81);
xor \U$6363 ( \6458 , \6456 , \6457 );
buf \U$6364 ( \6459 , \6458 );
buf \U$6365 ( \6460 , \6459 );
nand \U$6366 ( \6461 , \6455 , \6460 );
buf \U$6367 ( \6462 , \6461 );
buf \U$6368 ( \6463 , \6462 );
nand \U$6369 ( \6464 , \6454 , \6463 );
buf \U$6370 ( \6465 , \6464 );
buf \U$6371 ( \6466 , \5904 );
not \U$6372 ( \6467 , \6466 );
buf \U$6373 ( \6468 , \1225 );
not \U$6374 ( \6469 , \6468 );
or \U$6375 ( \6470 , \6467 , \6469 );
buf \U$6376 ( \6471 , \1229 );
buf \U$6377 ( \6472 , RIc0d9478_65);
buf \U$6378 ( \6473 , RIc0d8230_26);
xor \U$6379 ( \6474 , \6472 , \6473 );
buf \U$6380 ( \6475 , \6474 );
buf \U$6381 ( \6476 , \6475 );
nand \U$6382 ( \6477 , \6471 , \6476 );
buf \U$6383 ( \6478 , \6477 );
buf \U$6384 ( \6479 , \6478 );
nand \U$6385 ( \6480 , \6470 , \6479 );
buf \U$6386 ( \6481 , \6480 );
xor \U$6387 ( \6482 , \6465 , \6481 );
xor \U$6388 ( \6483 , \6449 , \6482 );
buf \U$6389 ( \6484 , \6483 );
xor \U$6390 ( \6485 , \6428 , \6484 );
buf \U$6391 ( \6486 , \6485 );
buf \U$6392 ( \6487 , \6486 );
xor \U$6393 ( \6488 , \6333 , \6487 );
xor \U$6394 ( \6489 , \5668 , \5674 );
and \U$6395 ( \6490 , \6489 , \5690 );
and \U$6396 ( \6491 , \5668 , \5674 );
or \U$6397 ( \6492 , \6490 , \6491 );
buf \U$6398 ( \6493 , \6492 );
buf \U$6399 ( \6494 , \6493 );
xor \U$6400 ( \6495 , \6488 , \6494 );
buf \U$6401 ( \6496 , \6495 );
buf \U$6402 ( \6497 , \6496 );
xor \U$6403 ( \6498 , \5883 , \6069 );
and \U$6404 ( \6499 , \6498 , \6076 );
and \U$6405 ( \6500 , \5883 , \6069 );
or \U$6406 ( \6501 , \6499 , \6500 );
buf \U$6407 ( \6502 , \6501 );
buf \U$6408 ( \6503 , \6502 );
xor \U$6409 ( \6504 , \6497 , \6503 );
xor \U$6410 ( \6505 , \5693 , \5699 );
and \U$6411 ( \6506 , \6505 , \5759 );
and \U$6412 ( \6507 , \5693 , \5699 );
or \U$6413 ( \6508 , \6506 , \6507 );
buf \U$6414 ( \6509 , \6508 );
buf \U$6415 ( \6510 , \6509 );
xor \U$6416 ( \6511 , \6504 , \6510 );
buf \U$6417 ( \6512 , \6511 );
buf \U$6418 ( \6513 , \6512 );
not \U$6419 ( \6514 , \6513 );
or \U$6420 ( \6515 , \6327 , \6514 );
buf \U$6421 ( \6516 , \6512 );
buf \U$6422 ( \6517 , \6325 );
or \U$6423 ( \6518 , \6516 , \6517 );
xor \U$6424 ( \6519 , \5775 , \6079 );
and \U$6425 ( \6520 , \6519 , \6086 );
and \U$6426 ( \6521 , \5775 , \6079 );
or \U$6427 ( \6522 , \6520 , \6521 );
buf \U$6428 ( \6523 , \6522 );
buf \U$6429 ( \6524 , \6523 );
nand \U$6430 ( \6525 , \6518 , \6524 );
buf \U$6431 ( \6526 , \6525 );
buf \U$6432 ( \6527 , \6526 );
nand \U$6433 ( \6528 , \6515 , \6527 );
buf \U$6434 ( \6529 , \6528 );
xor \U$6435 ( \6530 , \6124 , \6179 );
and \U$6436 ( \6531 , \6530 , \6186 );
and \U$6437 ( \6532 , \6124 , \6179 );
or \U$6438 ( \6533 , \6531 , \6532 );
buf \U$6439 ( \6534 , \6533 );
buf \U$6440 ( \6535 , \6534 );
xor \U$6441 ( \6536 , \6202 , \6244 );
and \U$6442 ( \6537 , \6536 , \6320 );
and \U$6443 ( \6538 , \6202 , \6244 );
or \U$6444 ( \6539 , \6537 , \6538 );
buf \U$6445 ( \6540 , \6539 );
buf \U$6446 ( \6541 , \6540 );
xor \U$6447 ( \6542 , \6535 , \6541 );
buf \U$6448 ( \6543 , \6176 );
xor \U$6449 ( \6544 , \6336 , \6351 );
and \U$6450 ( \6545 , \6544 , \6368 );
and \U$6451 ( \6546 , \6336 , \6351 );
or \U$6452 ( \6547 , \6545 , \6546 );
buf \U$6453 ( \6548 , \6547 );
buf \U$6454 ( \6549 , \6548 );
xor \U$6455 ( \6550 , \6543 , \6549 );
buf \U$6456 ( \6551 , \6314 );
not \U$6457 ( \6552 , \6551 );
buf \U$6458 ( \6553 , \6298 );
not \U$6459 ( \6554 , \6553 );
or \U$6460 ( \6555 , \6552 , \6554 );
buf \U$6461 ( \6556 , \6298 );
buf \U$6462 ( \6557 , \6314 );
or \U$6463 ( \6558 , \6556 , \6557 );
buf \U$6464 ( \6559 , \6282 );
nand \U$6465 ( \6560 , \6558 , \6559 );
buf \U$6466 ( \6561 , \6560 );
buf \U$6467 ( \6562 , \6561 );
nand \U$6468 ( \6563 , \6555 , \6562 );
buf \U$6469 ( \6564 , \6563 );
buf \U$6470 ( \6565 , \6564 );
xor \U$6471 ( \6566 , \6550 , \6565 );
buf \U$6472 ( \6567 , \6566 );
buf \U$6473 ( \6568 , \6567 );
xor \U$6474 ( \6569 , \6371 , \6427 );
and \U$6475 ( \6570 , \6569 , \6484 );
and \U$6476 ( \6571 , \6371 , \6427 );
or \U$6477 ( \6572 , \6570 , \6571 );
buf \U$6478 ( \6573 , \6572 );
buf \U$6479 ( \6574 , \6573 );
xor \U$6480 ( \6575 , \6568 , \6574 );
buf \U$6481 ( \6576 , \6481 );
not \U$6482 ( \6577 , \6576 );
buf \U$6483 ( \6578 , \6465 );
not \U$6484 ( \6579 , \6578 );
or \U$6485 ( \6580 , \6577 , \6579 );
buf \U$6486 ( \6581 , \6465 );
buf \U$6487 ( \6582 , \6481 );
or \U$6488 ( \6583 , \6581 , \6582 );
buf \U$6489 ( \6584 , \6449 );
nand \U$6490 ( \6585 , \6583 , \6584 );
buf \U$6491 ( \6586 , \6585 );
buf \U$6492 ( \6587 , \6586 );
nand \U$6493 ( \6588 , \6580 , \6587 );
buf \U$6494 ( \6589 , \6588 );
buf \U$6495 ( \6590 , \6589 );
xor \U$6496 ( \6591 , \6388 , \6406 );
and \U$6497 ( \6592 , \6591 , \6424 );
and \U$6498 ( \6593 , \6388 , \6406 );
or \U$6499 ( \6594 , \6592 , \6593 );
buf \U$6500 ( \6595 , \6594 );
buf \U$6501 ( \6596 , \6595 );
xor \U$6502 ( \6597 , \6590 , \6596 );
buf \U$6503 ( \6598 , \6459 );
not \U$6504 ( \6599 , \6598 );
buf \U$6505 ( \6600 , \1064 );
not \U$6506 ( \6601 , \6600 );
or \U$6507 ( \6602 , \6599 , \6601 );
buf \U$6508 ( \6603 , \1078 );
buf \U$6509 ( \6604 , RIc0d7a38_9);
buf \U$6510 ( \6605 , RIc0d9bf8_81);
xor \U$6511 ( \6606 , \6604 , \6605 );
buf \U$6512 ( \6607 , \6606 );
buf \U$6513 ( \6608 , \6607 );
nand \U$6514 ( \6609 , \6603 , \6608 );
buf \U$6515 ( \6610 , \6609 );
buf \U$6516 ( \6611 , \6610 );
nand \U$6517 ( \6612 , \6602 , \6611 );
buf \U$6518 ( \6613 , \6612 );
buf \U$6519 ( \6614 , \6613 );
not \U$6520 ( \6615 , \6614 );
buf \U$6521 ( \6616 , \6475 );
not \U$6522 ( \6617 , \6616 );
buf \U$6523 ( \6618 , \3781 );
not \U$6524 ( \6619 , \6618 );
or \U$6525 ( \6620 , \6617 , \6619 );
buf \U$6526 ( \6621 , \4427 );
buf \U$6527 ( \6622 , RIc0d9478_65);
buf \U$6528 ( \6623 , RIc0d81b8_25);
xor \U$6529 ( \6624 , \6622 , \6623 );
buf \U$6530 ( \6625 , \6624 );
buf \U$6531 ( \6626 , \6625 );
nand \U$6532 ( \6627 , \6621 , \6626 );
buf \U$6533 ( \6628 , \6627 );
buf \U$6534 ( \6629 , \6628 );
nand \U$6535 ( \6630 , \6620 , \6629 );
buf \U$6536 ( \6631 , \6630 );
buf \U$6537 ( \6632 , \6631 );
not \U$6538 ( \6633 , \6632 );
buf \U$6539 ( \6634 , \6633 );
buf \U$6540 ( \6635 , \6634 );
not \U$6541 ( \6636 , \6635 );
or \U$6542 ( \6637 , \6615 , \6636 );
buf \U$6543 ( \6638 , \6634 );
buf \U$6544 ( \6639 , \6613 );
or \U$6545 ( \6640 , \6638 , \6639 );
nand \U$6546 ( \6641 , \6637 , \6640 );
buf \U$6547 ( \6642 , \6641 );
buf \U$6548 ( \6643 , \6642 );
buf \U$6549 ( \6644 , \1435 );
buf \U$6550 ( \6645 , \6136 );
or \U$6551 ( \6646 , \6644 , \6645 );
buf \U$6552 ( \6647 , \1585 );
buf \U$6553 ( \6648 , RIc0d7c18_13);
buf \U$6554 ( \6649 , RIc0d9a18_77);
xnor \U$6555 ( \6650 , \6648 , \6649 );
buf \U$6556 ( \6651 , \6650 );
buf \U$6557 ( \6652 , \6651 );
or \U$6558 ( \6653 , \6647 , \6652 );
nand \U$6559 ( \6654 , \6646 , \6653 );
buf \U$6560 ( \6655 , \6654 );
buf \U$6561 ( \6656 , \6655 );
xor \U$6562 ( \6657 , \6643 , \6656 );
buf \U$6563 ( \6658 , \6657 );
buf \U$6564 ( \6659 , \6658 );
xor \U$6565 ( \6660 , \6597 , \6659 );
buf \U$6566 ( \6661 , \6660 );
buf \U$6567 ( \6662 , \6661 );
xor \U$6568 ( \6663 , \6575 , \6662 );
buf \U$6569 ( \6664 , \6663 );
buf \U$6570 ( \6665 , \6664 );
xor \U$6571 ( \6666 , \6542 , \6665 );
buf \U$6572 ( \6667 , \6666 );
buf \U$6573 ( \6668 , \6667 );
xor \U$6574 ( \6669 , \6497 , \6503 );
and \U$6575 ( \6670 , \6669 , \6510 );
and \U$6576 ( \6671 , \6497 , \6503 );
or \U$6577 ( \6672 , \6670 , \6671 );
buf \U$6578 ( \6673 , \6672 );
buf \U$6579 ( \6674 , \6673 );
xor \U$6580 ( \6675 , \6668 , \6674 );
xor \U$6581 ( \6676 , \6260 , \6266 );
and \U$6582 ( \6677 , \6676 , \6317 );
and \U$6583 ( \6678 , \6260 , \6266 );
or \U$6584 ( \6679 , \6677 , \6678 );
buf \U$6585 ( \6680 , \6679 );
buf \U$6586 ( \6681 , \6680 );
buf \U$6587 ( \6682 , \6381 );
not \U$6588 ( \6683 , \6682 );
buf \U$6589 ( \6684 , \1263 );
not \U$6590 ( \6685 , \6684 );
or \U$6591 ( \6686 , \6683 , \6685 );
buf \U$6592 ( \6687 , \2927 );
buf \U$6593 ( \6688 , RIc0d7ee8_19);
buf \U$6594 ( \6689 , RIc0d9748_71);
xor \U$6595 ( \6690 , \6688 , \6689 );
buf \U$6596 ( \6691 , \6690 );
buf \U$6597 ( \6692 , \6691 );
nand \U$6598 ( \6693 , \6687 , \6692 );
buf \U$6599 ( \6694 , \6693 );
buf \U$6600 ( \6695 , \6694 );
nand \U$6601 ( \6696 , \6686 , \6695 );
buf \U$6602 ( \6697 , \6696 );
buf \U$6603 ( \6698 , \6697 );
buf \U$6604 ( \6699 , \3816 );
buf \U$6605 ( \6700 , \6342 );
or \U$6606 ( \6701 , \6699 , \6700 );
buf \U$6607 ( \6702 , \1562 );
buf \U$6608 ( \6703 , RIc0d7d08_15);
buf \U$6609 ( \6704 , RIc0d9928_75);
xnor \U$6610 ( \6705 , \6703 , \6704 );
buf \U$6611 ( \6706 , \6705 );
buf \U$6612 ( \6707 , \6706 );
or \U$6613 ( \6708 , \6702 , \6707 );
nand \U$6614 ( \6709 , \6701 , \6708 );
buf \U$6615 ( \6710 , \6709 );
buf \U$6616 ( \6711 , \6710 );
xor \U$6617 ( \6712 , \6698 , \6711 );
buf \U$6618 ( \6713 , \1739 );
buf \U$6619 ( \6714 , \6419 );
or \U$6620 ( \6715 , \6713 , \6714 );
buf \U$6621 ( \6716 , \996 );
buf \U$6622 ( \6717 , RIc0d7948_7);
buf \U$6623 ( \6718 , RIc0d9ce8_83);
xnor \U$6624 ( \6719 , \6717 , \6718 );
buf \U$6625 ( \6720 , \6719 );
buf \U$6626 ( \6721 , \6720 );
or \U$6627 ( \6722 , \6716 , \6721 );
nand \U$6628 ( \6723 , \6715 , \6722 );
buf \U$6629 ( \6724 , \6723 );
buf \U$6630 ( \6725 , \6724 );
xor \U$6631 ( \6726 , \6712 , \6725 );
buf \U$6632 ( \6727 , \6726 );
buf \U$6633 ( \6728 , \6727 );
xor \U$6634 ( \6729 , \6147 , \6163 );
not \U$6635 ( \6730 , \6176 );
and \U$6636 ( \6731 , \6729 , \6730 );
and \U$6637 ( \6732 , \6147 , \6163 );
or \U$6638 ( \6733 , \6731 , \6732 );
buf \U$6639 ( \6734 , \6733 );
xor \U$6640 ( \6735 , \6728 , \6734 );
xor \U$6641 ( \6736 , \6208 , \6225 );
and \U$6642 ( \6737 , \6736 , \6241 );
and \U$6643 ( \6738 , \6208 , \6225 );
or \U$6644 ( \6739 , \6737 , \6738 );
buf \U$6645 ( \6740 , \6739 );
buf \U$6646 ( \6741 , \6740 );
xor \U$6647 ( \6742 , \6735 , \6741 );
buf \U$6648 ( \6743 , \6742 );
buf \U$6649 ( \6744 , \6743 );
xor \U$6650 ( \6745 , \6681 , \6744 );
and \U$6651 ( \6746 , \5901 , \5902 );
buf \U$6652 ( \6747 , \6746 );
buf \U$6653 ( \6748 , \6747 );
buf \U$6654 ( \6749 , \6442 );
not \U$6655 ( \6750 , \6749 );
buf \U$6656 ( \6751 , \1823 );
not \U$6657 ( \6752 , \6751 );
or \U$6658 ( \6753 , \6750 , \6752 );
buf \U$6659 ( \6754 , \686 );
buf \U$6660 ( \6755 , RIc0d80c8_23);
buf \U$6661 ( \6756 , RIc0d9568_67);
xor \U$6662 ( \6757 , \6755 , \6756 );
buf \U$6663 ( \6758 , \6757 );
buf \U$6664 ( \6759 , \6758 );
nand \U$6665 ( \6760 , \6754 , \6759 );
buf \U$6666 ( \6761 , \6760 );
buf \U$6667 ( \6762 , \6761 );
nand \U$6668 ( \6763 , \6753 , \6762 );
buf \U$6669 ( \6764 , \6763 );
buf \U$6670 ( \6765 , \6764 );
xor \U$6671 ( \6766 , \6748 , \6765 );
buf \U$6672 ( \6767 , \711 );
not \U$6673 ( \6768 , \6767 );
buf \U$6674 ( \6769 , \521 );
not \U$6675 ( \6770 , \6769 );
or \U$6676 ( \6771 , \6768 , \6770 );
buf \U$6677 ( \6772 , RIc0da0a8_91);
nand \U$6678 ( \6773 , \6771 , \6772 );
buf \U$6679 ( \6774 , \6773 );
buf \U$6680 ( \6775 , \6774 );
xnor \U$6681 ( \6776 , \6766 , \6775 );
buf \U$6682 ( \6777 , \6776 );
buf \U$6683 ( \6778 , \6308 );
not \U$6684 ( \6779 , \6778 );
buf \U$6685 ( \6780 , \397 );
not \U$6686 ( \6781 , \6780 );
or \U$6687 ( \6782 , \6779 , \6781 );
buf \U$6688 ( \6783 , RIc0d9b08_79);
buf \U$6689 ( \6784 , RIc0d7b28_11);
xnor \U$6690 ( \6785 , \6783 , \6784 );
buf \U$6691 ( \6786 , \6785 );
buf \U$6692 ( \6787 , \6786 );
not \U$6693 ( \6788 , \6787 );
buf \U$6694 ( \6789 , \403 );
nand \U$6695 ( \6790 , \6788 , \6789 );
buf \U$6696 ( \6791 , \6790 );
buf \U$6697 ( \6792 , \6791 );
nand \U$6698 ( \6793 , \6782 , \6792 );
buf \U$6699 ( \6794 , \6793 );
buf \U$6700 ( \6795 , \6794 );
buf \U$6701 ( \6796 , \6278 );
not \U$6702 ( \6797 , \6796 );
buf \U$6703 ( \6798 , \6797 );
buf \U$6704 ( \6799 , \6798 );
not \U$6705 ( \6800 , \6799 );
buf \U$6706 ( \6801 , \2607 );
not \U$6707 ( \6802 , \6801 );
or \U$6708 ( \6803 , \6800 , \6802 );
buf \U$6709 ( \6804 , \816 );
buf \U$6710 ( \6805 , RIc0d9ec8_87);
buf \U$6711 ( \6806 , RIc0d7768_3);
and \U$6712 ( \6807 , \6805 , \6806 );
not \U$6713 ( \6808 , \6805 );
buf \U$6714 ( \6809 , \304 );
and \U$6715 ( \6810 , \6808 , \6809 );
nor \U$6716 ( \6811 , \6807 , \6810 );
buf \U$6717 ( \6812 , \6811 );
buf \U$6718 ( \6813 , \6812 );
nand \U$6719 ( \6814 , \6804 , \6813 );
buf \U$6720 ( \6815 , \6814 );
buf \U$6721 ( \6816 , \6815 );
nand \U$6722 ( \6817 , \6803 , \6816 );
buf \U$6723 ( \6818 , \6817 );
buf \U$6724 ( \6819 , \6818 );
xor \U$6725 ( \6820 , \6795 , \6819 );
buf \U$6726 ( \6821 , \437 );
not \U$6727 ( \6822 , \6821 );
buf \U$6728 ( \6823 , \6822 );
buf \U$6729 ( \6824 , \6823 );
buf \U$6730 ( \6825 , \6397 );
or \U$6731 ( \6826 , \6824 , \6825 );
buf \U$6732 ( \6827 , \442 );
not \U$6733 ( \6828 , \6827 );
buf \U$6734 ( \6829 , \6828 );
buf \U$6735 ( \6830 , \6829 );
buf \U$6736 ( \6831 , \599 );
buf \U$6737 ( \6832 , RIc0d7678_1);
and \U$6738 ( \6833 , \6831 , \6832 );
buf \U$6739 ( \6834 , \974 );
buf \U$6740 ( \6835 , RIc0d9fb8_89);
and \U$6741 ( \6836 , \6834 , \6835 );
nor \U$6742 ( \6837 , \6833 , \6836 );
buf \U$6743 ( \6838 , \6837 );
buf \U$6744 ( \6839 , \6838 );
or \U$6745 ( \6840 , \6830 , \6839 );
nand \U$6746 ( \6841 , \6826 , \6840 );
buf \U$6747 ( \6842 , \6841 );
buf \U$6748 ( \6843 , \6842 );
xor \U$6749 ( \6844 , \6820 , \6843 );
buf \U$6750 ( \6845 , \6844 );
xnor \U$6751 ( \6846 , \6777 , \6845 );
buf \U$6752 ( \6847 , \6846 );
buf \U$6753 ( \6848 , \6360 );
not \U$6754 ( \6849 , \6848 );
buf \U$6755 ( \6850 , \279 );
not \U$6756 ( \6851 , \6850 );
or \U$6757 ( \6852 , \6849 , \6851 );
buf \U$6758 ( \6853 , RIc0d9658_69);
buf \U$6759 ( \6854 , RIc0d7fd8_21);
xnor \U$6760 ( \6855 , \6853 , \6854 );
buf \U$6761 ( \6856 , \6855 );
buf \U$6762 ( \6857 , \6856 );
not \U$6763 ( \6858 , \6857 );
buf \U$6764 ( \6859 , \874 );
nand \U$6765 ( \6860 , \6858 , \6859 );
buf \U$6766 ( \6861 , \6860 );
buf \U$6767 ( \6862 , \6861 );
nand \U$6768 ( \6863 , \6852 , \6862 );
buf \U$6769 ( \6864 , \6863 );
buf \U$6770 ( \6865 , \6157 );
not \U$6771 ( \6866 , \6865 );
buf \U$6772 ( \6867 , \6029 );
not \U$6773 ( \6868 , \6867 );
or \U$6774 ( \6869 , \6866 , \6868 );
buf \U$6775 ( \6870 , \2960 );
buf \U$6776 ( \6871 , RIc0d7858_5);
buf \U$6777 ( \6872 , RIc0d9dd8_85);
xor \U$6778 ( \6873 , \6871 , \6872 );
buf \U$6779 ( \6874 , \6873 );
buf \U$6780 ( \6875 , \6874 );
nand \U$6781 ( \6876 , \6870 , \6875 );
buf \U$6782 ( \6877 , \6876 );
buf \U$6783 ( \6878 , \6877 );
nand \U$6784 ( \6879 , \6869 , \6878 );
buf \U$6785 ( \6880 , \6879 );
xor \U$6786 ( \6881 , \6864 , \6880 );
buf \U$6787 ( \6882 , RIc0d7df8_17);
buf \U$6788 ( \6883 , RIc0d9838_73);
xor \U$6789 ( \6884 , \6882 , \6883 );
buf \U$6790 ( \6885 , \6884 );
buf \U$6791 ( \6886 , \6885 );
not \U$6792 ( \6887 , \6886 );
buf \U$6793 ( \6888 , \2882 );
not \U$6794 ( \6889 , \6888 );
or \U$6795 ( \6890 , \6887 , \6889 );
buf \U$6796 ( \6891 , \1677 );
buf \U$6797 ( \6892 , \6292 );
nand \U$6798 ( \6893 , \6891 , \6892 );
buf \U$6799 ( \6894 , \6893 );
buf \U$6800 ( \6895 , \6894 );
nand \U$6801 ( \6896 , \6890 , \6895 );
buf \U$6802 ( \6897 , \6896 );
xnor \U$6803 ( \6898 , \6881 , \6897 );
buf \U$6804 ( \6899 , \6898 );
not \U$6805 ( \6900 , \6899 );
buf \U$6806 ( \6901 , \6900 );
buf \U$6807 ( \6902 , \6901 );
and \U$6808 ( \6903 , \6847 , \6902 );
not \U$6809 ( \6904 , \6847 );
buf \U$6810 ( \6905 , \6898 );
and \U$6811 ( \6906 , \6904 , \6905 );
nor \U$6812 ( \6907 , \6903 , \6906 );
buf \U$6813 ( \6908 , \6907 );
buf \U$6814 ( \6909 , \6908 );
xor \U$6815 ( \6910 , \6745 , \6909 );
buf \U$6816 ( \6911 , \6910 );
buf \U$6817 ( \6912 , \6911 );
xor \U$6818 ( \6913 , \6333 , \6487 );
and \U$6819 ( \6914 , \6913 , \6494 );
and \U$6820 ( \6915 , \6333 , \6487 );
or \U$6821 ( \6916 , \6914 , \6915 );
buf \U$6822 ( \6917 , \6916 );
buf \U$6823 ( \6918 , \6917 );
xor \U$6824 ( \6919 , \6912 , \6918 );
xor \U$6825 ( \6920 , \6189 , \6195 );
and \U$6826 ( \6921 , \6920 , \6323 );
and \U$6827 ( \6922 , \6189 , \6195 );
or \U$6828 ( \6923 , \6921 , \6922 );
buf \U$6829 ( \6924 , \6923 );
buf \U$6830 ( \6925 , \6924 );
xor \U$6831 ( \6926 , \6919 , \6925 );
buf \U$6832 ( \6927 , \6926 );
buf \U$6833 ( \6928 , \6927 );
xor \U$6834 ( \6929 , \6675 , \6928 );
buf \U$6835 ( \6930 , \6929 );
or \U$6836 ( \6931 , \6529 , \6930 );
buf \U$6837 ( \6932 , \6931 );
xor \U$6838 ( \6933 , \5762 , \5768 );
and \U$6839 ( \6934 , \6933 , \6089 );
and \U$6840 ( \6935 , \5762 , \5768 );
or \U$6841 ( \6936 , \6934 , \6935 );
buf \U$6842 ( \6937 , \6936 );
buf \U$6843 ( \6938 , \6937 );
not \U$6844 ( \6939 , \6938 );
buf \U$6845 ( \6940 , \6512 );
not \U$6846 ( \6941 , \6940 );
buf \U$6847 ( \6942 , \6941 );
xor \U$6848 ( \6943 , \6325 , \6942 );
xor \U$6849 ( \6944 , \6943 , \6523 );
buf \U$6850 ( \6945 , \6944 );
nand \U$6851 ( \6946 , \6939 , \6945 );
buf \U$6852 ( \6947 , \6946 );
buf \U$6853 ( \6948 , \6947 );
and \U$6854 ( \6949 , \6932 , \6948 );
buf \U$6855 ( \6950 , \6949 );
buf \U$6856 ( \6951 , \6950 );
xor \U$6857 ( \6952 , \6568 , \6574 );
and \U$6858 ( \6953 , \6952 , \6662 );
and \U$6859 ( \6954 , \6568 , \6574 );
or \U$6860 ( \6955 , \6953 , \6954 );
buf \U$6861 ( \6956 , \6955 );
buf \U$6862 ( \6957 , \6956 );
xor \U$6863 ( \6958 , \6728 , \6734 );
and \U$6864 ( \6959 , \6958 , \6741 );
and \U$6865 ( \6960 , \6728 , \6734 );
or \U$6866 ( \6961 , \6959 , \6960 );
buf \U$6867 ( \6962 , \6961 );
buf \U$6868 ( \6963 , \6962 );
xor \U$6869 ( \6964 , \6957 , \6963 );
buf \U$6870 ( \6965 , \393 );
buf \U$6871 ( \6966 , \6786 );
or \U$6872 ( \6967 , \6965 , \6966 );
buf \U$6873 ( \6968 , \2493 );
buf \U$6874 ( \6969 , RIc0d7ab0_10);
buf \U$6875 ( \6970 , RIc0d9b08_79);
xnor \U$6876 ( \6971 , \6969 , \6970 );
buf \U$6877 ( \6972 , \6971 );
buf \U$6878 ( \6973 , \6972 );
or \U$6879 ( \6974 , \6968 , \6973 );
nand \U$6880 ( \6975 , \6967 , \6974 );
buf \U$6881 ( \6976 , \6975 );
buf \U$6882 ( \6977 , \6976 );
buf \U$6883 ( \6978 , \6812 );
not \U$6884 ( \6979 , \6978 );
buf \U$6885 ( \6980 , \809 );
not \U$6886 ( \6981 , \6980 );
or \U$6887 ( \6982 , \6979 , \6981 );
buf \U$6888 ( \6983 , RIc0d76f0_2);
buf \U$6889 ( \6984 , RIc0d9ec8_87);
xnor \U$6890 ( \6985 , \6983 , \6984 );
buf \U$6891 ( \6986 , \6985 );
buf \U$6892 ( \6987 , \6986 );
not \U$6893 ( \6988 , \6987 );
buf \U$6894 ( \6989 , \3631 );
nand \U$6895 ( \6990 , \6988 , \6989 );
buf \U$6896 ( \6991 , \6990 );
buf \U$6897 ( \6992 , \6991 );
nand \U$6898 ( \6993 , \6982 , \6992 );
buf \U$6899 ( \6994 , \6993 );
buf \U$6900 ( \6995 , \6994 );
not \U$6901 ( \6996 , \6995 );
buf \U$6902 ( \6997 , \6996 );
buf \U$6903 ( \6998 , \6997 );
xor \U$6904 ( \6999 , \6977 , \6998 );
xor \U$6905 ( \7000 , \6795 , \6819 );
and \U$6906 ( \7001 , \7000 , \6843 );
and \U$6907 ( \7002 , \6795 , \6819 );
or \U$6908 ( \7003 , \7001 , \7002 );
buf \U$6909 ( \7004 , \7003 );
buf \U$6910 ( \7005 , \7004 );
xor \U$6911 ( \7006 , \6999 , \7005 );
buf \U$6912 ( \7007 , \7006 );
buf \U$6913 ( \7008 , \7007 );
buf \U$6914 ( \7009 , \6777 );
not \U$6915 ( \7010 , \7009 );
buf \U$6916 ( \7011 , \7010 );
buf \U$6917 ( \7012 , \7011 );
not \U$6918 ( \7013 , \7012 );
buf \U$6919 ( \7014 , \6901 );
not \U$6920 ( \7015 , \7014 );
or \U$6921 ( \7016 , \7013 , \7015 );
buf \U$6922 ( \7017 , \6777 );
not \U$6923 ( \7018 , \7017 );
buf \U$6924 ( \7019 , \6898 );
not \U$6925 ( \7020 , \7019 );
or \U$6926 ( \7021 , \7018 , \7020 );
buf \U$6927 ( \7022 , \6845 );
nand \U$6928 ( \7023 , \7021 , \7022 );
buf \U$6929 ( \7024 , \7023 );
buf \U$6930 ( \7025 , \7024 );
nand \U$6931 ( \7026 , \7016 , \7025 );
buf \U$6932 ( \7027 , \7026 );
buf \U$6933 ( \7028 , \7027 );
xor \U$6934 ( \7029 , \7008 , \7028 );
xor \U$6935 ( \7030 , \6698 , \6711 );
and \U$6936 ( \7031 , \7030 , \6725 );
and \U$6937 ( \7032 , \6698 , \6711 );
or \U$6938 ( \7033 , \7031 , \7032 );
buf \U$6939 ( \7034 , \7033 );
not \U$6940 ( \7035 , \6613 );
nand \U$6941 ( \7036 , \7035 , \6634 );
not \U$6942 ( \7037 , \7036 );
not \U$6943 ( \7038 , \6655 );
or \U$6944 ( \7039 , \7037 , \7038 );
buf \U$6945 ( \7040 , \6613 );
buf \U$6946 ( \7041 , \6631 );
nand \U$6947 ( \7042 , \7040 , \7041 );
buf \U$6948 ( \7043 , \7042 );
nand \U$6949 ( \7044 , \7039 , \7043 );
xor \U$6950 ( \7045 , \7034 , \7044 );
buf \U$6951 ( \7046 , \6880 );
not \U$6952 ( \7047 , \7046 );
buf \U$6953 ( \7048 , \6864 );
not \U$6954 ( \7049 , \7048 );
or \U$6955 ( \7050 , \7047 , \7049 );
buf \U$6956 ( \7051 , \6880 );
buf \U$6957 ( \7052 , \6864 );
or \U$6958 ( \7053 , \7051 , \7052 );
buf \U$6959 ( \7054 , \6897 );
nand \U$6960 ( \7055 , \7053 , \7054 );
buf \U$6961 ( \7056 , \7055 );
buf \U$6962 ( \7057 , \7056 );
nand \U$6963 ( \7058 , \7050 , \7057 );
buf \U$6964 ( \7059 , \7058 );
xor \U$6965 ( \7060 , \7045 , \7059 );
buf \U$6966 ( \7061 , \7060 );
xor \U$6967 ( \7062 , \7029 , \7061 );
buf \U$6968 ( \7063 , \7062 );
buf \U$6969 ( \7064 , \7063 );
xor \U$6970 ( \7065 , \6964 , \7064 );
buf \U$6971 ( \7066 , \7065 );
buf \U$6972 ( \7067 , \7066 );
xor \U$6973 ( \7068 , \6912 , \6918 );
and \U$6974 ( \7069 , \7068 , \6925 );
and \U$6975 ( \7070 , \6912 , \6918 );
or \U$6976 ( \7071 , \7069 , \7070 );
buf \U$6977 ( \7072 , \7071 );
buf \U$6978 ( \7073 , \7072 );
xor \U$6979 ( \7074 , \7067 , \7073 );
xor \U$6980 ( \7075 , \6681 , \6744 );
and \U$6981 ( \7076 , \7075 , \6909 );
and \U$6982 ( \7077 , \6681 , \6744 );
or \U$6983 ( \7078 , \7076 , \7077 );
buf \U$6984 ( \7079 , \7078 );
buf \U$6985 ( \7080 , \7079 );
xor \U$6986 ( \7081 , \6590 , \6596 );
and \U$6987 ( \7082 , \7081 , \6659 );
and \U$6988 ( \7083 , \6590 , \6596 );
or \U$6989 ( \7084 , \7082 , \7083 );
buf \U$6990 ( \7085 , \7084 );
buf \U$6991 ( \7086 , \7085 );
buf \U$6992 ( \7087 , \6747 );
not \U$6993 ( \7088 , \7087 );
buf \U$6994 ( \7089 , \6764 );
not \U$6995 ( \7090 , \7089 );
or \U$6996 ( \7091 , \7088 , \7090 );
buf \U$6997 ( \7092 , \6764 );
buf \U$6998 ( \7093 , \6747 );
or \U$6999 ( \7094 , \7092 , \7093 );
buf \U$7000 ( \7095 , \6774 );
nand \U$7001 ( \7096 , \7094 , \7095 );
buf \U$7002 ( \7097 , \7096 );
buf \U$7003 ( \7098 , \7097 );
nand \U$7004 ( \7099 , \7091 , \7098 );
buf \U$7005 ( \7100 , \7099 );
buf \U$7006 ( \7101 , \7100 );
buf \U$7007 ( \7102 , \6691 );
not \U$7008 ( \7103 , \7102 );
buf \U$7009 ( \7104 , \2269 );
not \U$7010 ( \7105 , \7104 );
or \U$7011 ( \7106 , \7103 , \7105 );
buf \U$7012 ( \7107 , \2927 );
buf \U$7013 ( \7108 , RIc0d7e70_18);
buf \U$7014 ( \7109 , RIc0d9748_71);
xor \U$7015 ( \7110 , \7108 , \7109 );
buf \U$7016 ( \7111 , \7110 );
buf \U$7017 ( \7112 , \7111 );
nand \U$7018 ( \7113 , \7107 , \7112 );
buf \U$7019 ( \7114 , \7113 );
buf \U$7020 ( \7115 , \7114 );
nand \U$7021 ( \7116 , \7106 , \7115 );
buf \U$7022 ( \7117 , \7116 );
buf \U$7023 ( \7118 , \7117 );
buf \U$7024 ( \7119 , \6651 );
not \U$7025 ( \7120 , \7119 );
buf \U$7026 ( \7121 , \7120 );
buf \U$7027 ( \7122 , \7121 );
not \U$7028 ( \7123 , \7122 );
buf \U$7029 ( \7124 , \1432 );
not \U$7030 ( \7125 , \7124 );
or \U$7031 ( \7126 , \7123 , \7125 );
buf \U$7032 ( \7127 , \6141 );
buf \U$7033 ( \7128 , RIc0d7ba0_12);
buf \U$7034 ( \7129 , RIc0d9a18_77);
xor \U$7035 ( \7130 , \7128 , \7129 );
buf \U$7036 ( \7131 , \7130 );
buf \U$7037 ( \7132 , \7131 );
nand \U$7038 ( \7133 , \7127 , \7132 );
buf \U$7039 ( \7134 , \7133 );
buf \U$7040 ( \7135 , \7134 );
nand \U$7041 ( \7136 , \7126 , \7135 );
buf \U$7042 ( \7137 , \7136 );
buf \U$7043 ( \7138 , \7137 );
xor \U$7044 ( \7139 , \7118 , \7138 );
buf \U$7045 ( \7140 , \6823 );
buf \U$7046 ( \7141 , \6838 );
or \U$7047 ( \7142 , \7140 , \7141 );
buf \U$7048 ( \7143 , \6829 );
buf \U$7049 ( \7144 , \599 );
or \U$7050 ( \7145 , \7143 , \7144 );
nand \U$7051 ( \7146 , \7142 , \7145 );
buf \U$7052 ( \7147 , \7146 );
buf \U$7053 ( \7148 , \7147 );
xor \U$7054 ( \7149 , \7139 , \7148 );
buf \U$7055 ( \7150 , \7149 );
buf \U$7056 ( \7151 , \7150 );
xor \U$7057 ( \7152 , \7101 , \7151 );
and \U$7058 ( \7153 , \6472 , \6473 );
buf \U$7059 ( \7154 , \7153 );
buf \U$7060 ( \7155 , \7154 );
buf \U$7061 ( \7156 , \6885 );
not \U$7062 ( \7157 , \7156 );
buf \U$7063 ( \7158 , \1677 );
not \U$7064 ( \7159 , \7158 );
or \U$7065 ( \7160 , \7157 , \7159 );
buf \U$7066 ( \7161 , \2882 );
buf \U$7067 ( \7162 , RIc0d7d80_16);
buf \U$7068 ( \7163 , RIc0d9838_73);
xor \U$7069 ( \7164 , \7162 , \7163 );
buf \U$7070 ( \7165 , \7164 );
buf \U$7071 ( \7166 , \7165 );
nand \U$7072 ( \7167 , \7161 , \7166 );
buf \U$7073 ( \7168 , \7167 );
buf \U$7074 ( \7169 , \7168 );
nand \U$7075 ( \7170 , \7160 , \7169 );
buf \U$7076 ( \7171 , \7170 );
buf \U$7077 ( \7172 , \7171 );
xor \U$7078 ( \7173 , \7155 , \7172 );
buf \U$7079 ( \7174 , \3816 );
buf \U$7080 ( \7175 , \6706 );
or \U$7081 ( \7176 , \7174 , \7175 );
buf \U$7082 ( \7177 , \2372 );
buf \U$7083 ( \7178 , RIc0d7c90_14);
buf \U$7084 ( \7179 , RIc0d9928_75);
xnor \U$7085 ( \7180 , \7178 , \7179 );
buf \U$7086 ( \7181 , \7180 );
buf \U$7087 ( \7182 , \7181 );
or \U$7088 ( \7183 , \7177 , \7182 );
nand \U$7089 ( \7184 , \7176 , \7183 );
buf \U$7090 ( \7185 , \7184 );
buf \U$7091 ( \7186 , \7185 );
xor \U$7092 ( \7187 , \7173 , \7186 );
buf \U$7093 ( \7188 , \7187 );
buf \U$7094 ( \7189 , \7188 );
xor \U$7095 ( \7190 , \7152 , \7189 );
buf \U$7096 ( \7191 , \7190 );
buf \U$7097 ( \7192 , \7191 );
xor \U$7098 ( \7193 , \7086 , \7192 );
buf \U$7099 ( \7194 , \6874 );
not \U$7100 ( \7195 , \7194 );
buf \U$7101 ( \7196 , \951 );
not \U$7102 ( \7197 , \7196 );
or \U$7103 ( \7198 , \7195 , \7197 );
buf \U$7104 ( \7199 , \2960 );
buf \U$7105 ( \7200 , RIc0d77e0_4);
buf \U$7106 ( \7201 , RIc0d9dd8_85);
xor \U$7107 ( \7202 , \7200 , \7201 );
buf \U$7108 ( \7203 , \7202 );
buf \U$7109 ( \7204 , \7203 );
nand \U$7110 ( \7205 , \7199 , \7204 );
buf \U$7111 ( \7206 , \7205 );
buf \U$7112 ( \7207 , \7206 );
nand \U$7113 ( \7208 , \7198 , \7207 );
buf \U$7114 ( \7209 , \7208 );
buf \U$7115 ( \7210 , \7209 );
buf \U$7116 ( \7211 , \6625 );
not \U$7117 ( \7212 , \7211 );
buf \U$7118 ( \7213 , \1225 );
not \U$7119 ( \7214 , \7213 );
or \U$7120 ( \7215 , \7212 , \7214 );
buf \U$7121 ( \7216 , RIc0d8140_24);
buf \U$7122 ( \7217 , RIc0d9478_65);
xnor \U$7123 ( \7218 , \7216 , \7217 );
buf \U$7124 ( \7219 , \7218 );
buf \U$7125 ( \7220 , \7219 );
not \U$7126 ( \7221 , \7220 );
buf \U$7127 ( \7222 , \4427 );
nand \U$7128 ( \7223 , \7221 , \7222 );
buf \U$7129 ( \7224 , \7223 );
buf \U$7130 ( \7225 , \7224 );
nand \U$7131 ( \7226 , \7215 , \7225 );
buf \U$7132 ( \7227 , \7226 );
buf \U$7133 ( \7228 , \7227 );
xor \U$7134 ( \7229 , \7210 , \7228 );
buf \U$7135 ( \7230 , \6720 );
not \U$7136 ( \7231 , \7230 );
buf \U$7137 ( \7232 , \7231 );
buf \U$7138 ( \7233 , \7232 );
not \U$7139 ( \7234 , \7233 );
buf \U$7140 ( \7235 , \574 );
not \U$7141 ( \7236 , \7235 );
or \U$7142 ( \7237 , \7234 , \7236 );
buf \U$7143 ( \7238 , \993 );
buf \U$7144 ( \7239 , RIc0d78d0_6);
buf \U$7145 ( \7240 , RIc0d9ce8_83);
xor \U$7146 ( \7241 , \7239 , \7240 );
buf \U$7147 ( \7242 , \7241 );
buf \U$7148 ( \7243 , \7242 );
nand \U$7149 ( \7244 , \7238 , \7243 );
buf \U$7150 ( \7245 , \7244 );
buf \U$7151 ( \7246 , \7245 );
nand \U$7152 ( \7247 , \7237 , \7246 );
buf \U$7153 ( \7248 , \7247 );
buf \U$7154 ( \7249 , \7248 );
xor \U$7155 ( \7250 , \7229 , \7249 );
buf \U$7156 ( \7251 , \7250 );
buf \U$7157 ( \7252 , \7251 );
buf \U$7158 ( \7253 , \6758 );
not \U$7159 ( \7254 , \7253 );
buf \U$7160 ( \7255 , \678 );
not \U$7161 ( \7256 , \7255 );
or \U$7162 ( \7257 , \7254 , \7256 );
buf \U$7163 ( \7258 , \686 );
buf \U$7164 ( \7259 , RIc0d8050_22);
buf \U$7165 ( \7260 , RIc0d9568_67);
xor \U$7166 ( \7261 , \7259 , \7260 );
buf \U$7167 ( \7262 , \7261 );
buf \U$7168 ( \7263 , \7262 );
nand \U$7169 ( \7264 , \7258 , \7263 );
buf \U$7170 ( \7265 , \7264 );
buf \U$7171 ( \7266 , \7265 );
nand \U$7172 ( \7267 , \7257 , \7266 );
buf \U$7173 ( \7268 , \7267 );
buf \U$7174 ( \7269 , \7268 );
buf \U$7175 ( \7270 , \6607 );
not \U$7176 ( \7271 , \7270 );
buf \U$7177 ( \7272 , \2766 );
not \U$7178 ( \7273 , \7272 );
or \U$7179 ( \7274 , \7271 , \7273 );
buf \U$7180 ( \7275 , \1078 );
buf \U$7181 ( \7276 , RIc0d79c0_8);
buf \U$7182 ( \7277 , RIc0d9bf8_81);
xor \U$7183 ( \7278 , \7276 , \7277 );
buf \U$7184 ( \7279 , \7278 );
buf \U$7185 ( \7280 , \7279 );
nand \U$7186 ( \7281 , \7275 , \7280 );
buf \U$7187 ( \7282 , \7281 );
buf \U$7188 ( \7283 , \7282 );
nand \U$7189 ( \7284 , \7274 , \7283 );
buf \U$7190 ( \7285 , \7284 );
buf \U$7191 ( \7286 , \7285 );
xor \U$7192 ( \7287 , \7269 , \7286 );
buf \U$7193 ( \7288 , \1452 );
buf \U$7194 ( \7289 , \6856 );
or \U$7195 ( \7290 , \7288 , \7289 );
buf \U$7196 ( \7291 , \4297 );
buf \U$7197 ( \7292 , RIc0d7f60_20);
buf \U$7198 ( \7293 , RIc0d9658_69);
xnor \U$7199 ( \7294 , \7292 , \7293 );
buf \U$7200 ( \7295 , \7294 );
buf \U$7201 ( \7296 , \7295 );
or \U$7202 ( \7297 , \7291 , \7296 );
nand \U$7203 ( \7298 , \7290 , \7297 );
buf \U$7204 ( \7299 , \7298 );
buf \U$7205 ( \7300 , \7299 );
xor \U$7206 ( \7301 , \7287 , \7300 );
buf \U$7207 ( \7302 , \7301 );
buf \U$7208 ( \7303 , \7302 );
xor \U$7209 ( \7304 , \7252 , \7303 );
xor \U$7210 ( \7305 , \6543 , \6549 );
and \U$7211 ( \7306 , \7305 , \6565 );
and \U$7212 ( \7307 , \6543 , \6549 );
or \U$7213 ( \7308 , \7306 , \7307 );
buf \U$7214 ( \7309 , \7308 );
buf \U$7215 ( \7310 , \7309 );
xor \U$7216 ( \7311 , \7304 , \7310 );
buf \U$7217 ( \7312 , \7311 );
buf \U$7218 ( \7313 , \7312 );
xor \U$7219 ( \7314 , \7193 , \7313 );
buf \U$7220 ( \7315 , \7314 );
buf \U$7221 ( \7316 , \7315 );
xor \U$7222 ( \7317 , \7080 , \7316 );
xor \U$7223 ( \7318 , \6535 , \6541 );
and \U$7224 ( \7319 , \7318 , \6665 );
and \U$7225 ( \7320 , \6535 , \6541 );
or \U$7226 ( \7321 , \7319 , \7320 );
buf \U$7227 ( \7322 , \7321 );
buf \U$7228 ( \7323 , \7322 );
xor \U$7229 ( \7324 , \7317 , \7323 );
buf \U$7230 ( \7325 , \7324 );
buf \U$7231 ( \7326 , \7325 );
xor \U$7232 ( \7327 , \7074 , \7326 );
buf \U$7233 ( \7328 , \7327 );
buf \U$7234 ( \7329 , \7328 );
xor \U$7235 ( \7330 , \6668 , \6674 );
and \U$7236 ( \7331 , \7330 , \6928 );
and \U$7237 ( \7332 , \6668 , \6674 );
or \U$7238 ( \7333 , \7331 , \7332 );
buf \U$7239 ( \7334 , \7333 );
buf \U$7240 ( \7335 , \7334 );
or \U$7241 ( \7336 , \7329 , \7335 );
buf \U$7242 ( \7337 , \7336 );
buf \U$7243 ( \7338 , \7337 );
xor \U$7244 ( \7339 , \6957 , \6963 );
and \U$7245 ( \7340 , \7339 , \7064 );
and \U$7246 ( \7341 , \6957 , \6963 );
or \U$7247 ( \7342 , \7340 , \7341 );
buf \U$7248 ( \7343 , \7342 );
buf \U$7249 ( \7344 , \7343 );
xor \U$7250 ( \7345 , \7080 , \7316 );
and \U$7251 ( \7346 , \7345 , \7323 );
and \U$7252 ( \7347 , \7080 , \7316 );
or \U$7253 ( \7348 , \7346 , \7347 );
buf \U$7254 ( \7349 , \7348 );
buf \U$7255 ( \7350 , \7349 );
xor \U$7256 ( \7351 , \7344 , \7350 );
xor \U$7257 ( \7352 , \7086 , \7192 );
and \U$7258 ( \7353 , \7352 , \7313 );
and \U$7259 ( \7354 , \7086 , \7192 );
or \U$7260 ( \7355 , \7353 , \7354 );
buf \U$7261 ( \7356 , \7355 );
buf \U$7262 ( \7357 , \7356 );
xor \U$7263 ( \7358 , \7101 , \7151 );
and \U$7264 ( \7359 , \7358 , \7189 );
and \U$7265 ( \7360 , \7101 , \7151 );
or \U$7266 ( \7361 , \7359 , \7360 );
buf \U$7267 ( \7362 , \7361 );
buf \U$7268 ( \7363 , \7362 );
xor \U$7269 ( \7364 , \7210 , \7228 );
and \U$7270 ( \7365 , \7364 , \7249 );
and \U$7271 ( \7366 , \7210 , \7228 );
or \U$7272 ( \7367 , \7365 , \7366 );
buf \U$7273 ( \7368 , \7367 );
buf \U$7274 ( \7369 , \7368 );
and \U$7275 ( \7370 , \6622 , \6623 );
buf \U$7276 ( \7371 , \7370 );
buf \U$7277 ( \7372 , \7371 );
buf \U$7278 ( \7373 , \7262 );
not \U$7279 ( \7374 , \7373 );
buf \U$7280 ( \7375 , \2900 );
not \U$7281 ( \7376 , \7375 );
or \U$7282 ( \7377 , \7374 , \7376 );
buf \U$7283 ( \7378 , RIc0d9568_67);
buf \U$7284 ( \7379 , RIc0d7fd8_21);
xnor \U$7285 ( \7380 , \7378 , \7379 );
buf \U$7286 ( \7381 , \7380 );
buf \U$7287 ( \7382 , \7381 );
not \U$7288 ( \7383 , \7382 );
buf \U$7289 ( \7384 , \686 );
nand \U$7290 ( \7385 , \7383 , \7384 );
buf \U$7291 ( \7386 , \7385 );
buf \U$7292 ( \7387 , \7386 );
nand \U$7293 ( \7388 , \7377 , \7387 );
buf \U$7294 ( \7389 , \7388 );
buf \U$7295 ( \7390 , \7389 );
xor \U$7296 ( \7391 , \7372 , \7390 );
buf \U$7297 ( \7392 , \7131 );
not \U$7298 ( \7393 , \7392 );
buf \U$7299 ( \7394 , \1432 );
not \U$7300 ( \7395 , \7394 );
or \U$7301 ( \7396 , \7393 , \7395 );
buf \U$7302 ( \7397 , \6141 );
buf \U$7303 ( \7398 , RIc0d7b28_11);
buf \U$7304 ( \7399 , RIc0d9a18_77);
xor \U$7305 ( \7400 , \7398 , \7399 );
buf \U$7306 ( \7401 , \7400 );
buf \U$7307 ( \7402 , \7401 );
nand \U$7308 ( \7403 , \7397 , \7402 );
buf \U$7309 ( \7404 , \7403 );
buf \U$7310 ( \7405 , \7404 );
nand \U$7311 ( \7406 , \7396 , \7405 );
buf \U$7312 ( \7407 , \7406 );
buf \U$7313 ( \7408 , \7407 );
xor \U$7314 ( \7409 , \7391 , \7408 );
buf \U$7315 ( \7410 , \7409 );
buf \U$7316 ( \7411 , \7410 );
xor \U$7317 ( \7412 , \7369 , \7411 );
buf \U$7318 ( \7413 , \7111 );
not \U$7319 ( \7414 , \7413 );
buf \U$7320 ( \7415 , \2269 );
not \U$7321 ( \7416 , \7415 );
or \U$7322 ( \7417 , \7414 , \7416 );
buf \U$7323 ( \7418 , \2927 );
buf \U$7324 ( \7419 , RIc0d7df8_17);
buf \U$7325 ( \7420 , RIc0d9748_71);
xor \U$7326 ( \7421 , \7419 , \7420 );
buf \U$7327 ( \7422 , \7421 );
buf \U$7328 ( \7423 , \7422 );
nand \U$7329 ( \7424 , \7418 , \7423 );
buf \U$7330 ( \7425 , \7424 );
buf \U$7331 ( \7426 , \7425 );
nand \U$7332 ( \7427 , \7417 , \7426 );
buf \U$7333 ( \7428 , \7427 );
buf \U$7334 ( \7429 , \7428 );
buf \U$7335 ( \7430 , \4692 );
not \U$7336 ( \7431 , \7430 );
buf \U$7337 ( \7432 , \7431 );
buf \U$7338 ( \7433 , \7432 );
buf \U$7339 ( \7434 , \7295 );
or \U$7340 ( \7435 , \7433 , \7434 );
buf \U$7341 ( \7436 , \4297 );
buf \U$7342 ( \7437 , RIc0d7ee8_19);
buf \U$7343 ( \7438 , RIc0d9658_69);
xnor \U$7344 ( \7439 , \7437 , \7438 );
buf \U$7345 ( \7440 , \7439 );
buf \U$7346 ( \7441 , \7440 );
or \U$7347 ( \7442 , \7436 , \7441 );
nand \U$7348 ( \7443 , \7435 , \7442 );
buf \U$7349 ( \7444 , \7443 );
buf \U$7350 ( \7445 , \7444 );
xor \U$7351 ( \7446 , \7429 , \7445 );
buf \U$7352 ( \7447 , \3781 );
not \U$7353 ( \7448 , \7447 );
buf \U$7354 ( \7449 , \7448 );
buf \U$7355 ( \7450 , \7449 );
buf \U$7356 ( \7451 , \7219 );
or \U$7357 ( \7452 , \7450 , \7451 );
buf \U$7358 ( \7453 , \1232 );
buf \U$7359 ( \7454 , RIc0d9478_65);
not \U$7360 ( \7455 , \7454 );
buf \U$7361 ( \7456 , \7455 );
buf \U$7362 ( \7457 , \7456 );
buf \U$7363 ( \7458 , RIc0d80c8_23);
and \U$7364 ( \7459 , \7457 , \7458 );
buf \U$7365 ( \7460 , RIc0d80c8_23);
not \U$7366 ( \7461 , \7460 );
buf \U$7367 ( \7462 , \7461 );
buf \U$7368 ( \7463 , \7462 );
buf \U$7369 ( \7464 , RIc0d9478_65);
and \U$7370 ( \7465 , \7463 , \7464 );
nor \U$7371 ( \7466 , \7459 , \7465 );
buf \U$7372 ( \7467 , \7466 );
buf \U$7373 ( \7468 , \7467 );
or \U$7374 ( \7469 , \7453 , \7468 );
nand \U$7375 ( \7470 , \7452 , \7469 );
buf \U$7376 ( \7471 , \7470 );
buf \U$7377 ( \7472 , \7471 );
xor \U$7378 ( \7473 , \7446 , \7472 );
buf \U$7379 ( \7474 , \7473 );
buf \U$7380 ( \7475 , \7474 );
xor \U$7381 ( \7476 , \7412 , \7475 );
buf \U$7382 ( \7477 , \7476 );
buf \U$7383 ( \7478 , \7477 );
xor \U$7384 ( \7479 , \7363 , \7478 );
buf \U$7385 ( \7480 , \5368 );
not \U$7386 ( \7481 , \7480 );
buf \U$7387 ( \7482 , \3387 );
not \U$7388 ( \7483 , \7482 );
or \U$7389 ( \7484 , \7481 , \7483 );
buf \U$7390 ( \7485 , RIc0d9fb8_89);
nand \U$7391 ( \7486 , \7484 , \7485 );
buf \U$7392 ( \7487 , \7486 );
buf \U$7393 ( \7488 , \7487 );
buf \U$7394 ( \7489 , \7279 );
not \U$7395 ( \7490 , \7489 );
buf \U$7396 ( \7491 , \2766 );
not \U$7397 ( \7492 , \7491 );
or \U$7398 ( \7493 , \7490 , \7492 );
buf \U$7399 ( \7494 , \1078 );
buf \U$7400 ( \7495 , RIc0d7948_7);
buf \U$7401 ( \7496 , RIc0d9bf8_81);
xor \U$7402 ( \7497 , \7495 , \7496 );
buf \U$7403 ( \7498 , \7497 );
buf \U$7404 ( \7499 , \7498 );
nand \U$7405 ( \7500 , \7494 , \7499 );
buf \U$7406 ( \7501 , \7500 );
buf \U$7407 ( \7502 , \7501 );
nand \U$7408 ( \7503 , \7493 , \7502 );
buf \U$7409 ( \7504 , \7503 );
buf \U$7410 ( \7505 , \7504 );
xor \U$7411 ( \7506 , \7488 , \7505 );
buf \U$7412 ( \7507 , \6994 );
xor \U$7413 ( \7508 , \7506 , \7507 );
buf \U$7414 ( \7509 , \7508 );
buf \U$7415 ( \7510 , \7509 );
buf \U$7416 ( \7511 , \6972 );
not \U$7417 ( \7512 , \7511 );
buf \U$7418 ( \7513 , \7512 );
buf \U$7419 ( \7514 , \7513 );
not \U$7420 ( \7515 , \7514 );
buf \U$7421 ( \7516 , \1351 );
not \U$7422 ( \7517 , \7516 );
or \U$7423 ( \7518 , \7515 , \7517 );
buf \U$7424 ( \7519 , RIc0d7a38_9);
buf \U$7425 ( \7520 , RIc0d9b08_79);
xnor \U$7426 ( \7521 , \7519 , \7520 );
buf \U$7427 ( \7522 , \7521 );
buf \U$7428 ( \7523 , \7522 );
not \U$7429 ( \7524 , \7523 );
buf \U$7430 ( \7525 , \403 );
nand \U$7431 ( \7526 , \7524 , \7525 );
buf \U$7432 ( \7527 , \7526 );
buf \U$7433 ( \7528 , \7527 );
nand \U$7434 ( \7529 , \7518 , \7528 );
buf \U$7435 ( \7530 , \7529 );
buf \U$7436 ( \7531 , \7530 );
buf \U$7437 ( \7532 , \7165 );
not \U$7438 ( \7533 , \7532 );
buf \U$7439 ( \7534 , \2871 );
not \U$7440 ( \7535 , \7534 );
or \U$7441 ( \7536 , \7533 , \7535 );
buf \U$7442 ( \7537 , \2882 );
buf \U$7443 ( \7538 , RIc0d7d08_15);
buf \U$7444 ( \7539 , RIc0d9838_73);
xor \U$7445 ( \7540 , \7538 , \7539 );
buf \U$7446 ( \7541 , \7540 );
buf \U$7447 ( \7542 , \7541 );
nand \U$7448 ( \7543 , \7537 , \7542 );
buf \U$7449 ( \7544 , \7543 );
buf \U$7450 ( \7545 , \7544 );
nand \U$7451 ( \7546 , \7536 , \7545 );
buf \U$7452 ( \7547 , \7546 );
buf \U$7453 ( \7548 , \7547 );
xor \U$7454 ( \7549 , \7531 , \7548 );
buf \U$7455 ( \7550 , \812 );
buf \U$7456 ( \7551 , \6986 );
or \U$7457 ( \7552 , \7550 , \7551 );
buf \U$7458 ( \7553 , \819 );
buf \U$7459 ( \7554 , RIc0d9ec8_87);
not \U$7460 ( \7555 , \7554 );
buf \U$7461 ( \7556 , \7555 );
buf \U$7462 ( \7557 , \7556 );
buf \U$7463 ( \7558 , RIc0d7678_1);
and \U$7464 ( \7559 , \7557 , \7558 );
buf \U$7465 ( \7560 , \974 );
buf \U$7466 ( \7561 , RIc0d9ec8_87);
and \U$7467 ( \7562 , \7560 , \7561 );
nor \U$7468 ( \7563 , \7559 , \7562 );
buf \U$7469 ( \7564 , \7563 );
buf \U$7470 ( \7565 , \7564 );
or \U$7471 ( \7566 , \7553 , \7565 );
nand \U$7472 ( \7567 , \7552 , \7566 );
buf \U$7473 ( \7568 , \7567 );
buf \U$7474 ( \7569 , \7568 );
xor \U$7475 ( \7570 , \7549 , \7569 );
buf \U$7476 ( \7571 , \7570 );
buf \U$7477 ( \7572 , \7571 );
xor \U$7478 ( \7573 , \7510 , \7572 );
buf \U$7479 ( \7574 , \7181 );
not \U$7480 ( \7575 , \7574 );
buf \U$7481 ( \7576 , \7575 );
buf \U$7482 ( \7577 , \7576 );
not \U$7483 ( \7578 , \7577 );
buf \U$7484 ( \7579 , \1129 );
not \U$7485 ( \7580 , \7579 );
or \U$7486 ( \7581 , \7578 , \7580 );
buf \U$7487 ( \7582 , \1143 );
buf \U$7488 ( \7583 , RIc0d9928_75);
buf \U$7489 ( \7584 , RIc0d7c18_13);
and \U$7490 ( \7585 , \7583 , \7584 );
not \U$7491 ( \7586 , \7583 );
buf \U$7492 ( \7587 , \1001 );
and \U$7493 ( \7588 , \7586 , \7587 );
nor \U$7494 ( \7589 , \7585 , \7588 );
buf \U$7495 ( \7590 , \7589 );
buf \U$7496 ( \7591 , \7590 );
nand \U$7497 ( \7592 , \7582 , \7591 );
buf \U$7498 ( \7593 , \7592 );
buf \U$7499 ( \7594 , \7593 );
nand \U$7500 ( \7595 , \7581 , \7594 );
buf \U$7501 ( \7596 , \7595 );
buf \U$7502 ( \7597 , \7242 );
not \U$7503 ( \7598 , \7597 );
buf \U$7504 ( \7599 , \574 );
not \U$7505 ( \7600 , \7599 );
or \U$7506 ( \7601 , \7598 , \7600 );
buf \U$7507 ( \7602 , \584 );
buf \U$7508 ( \7603 , RIc0d7858_5);
buf \U$7509 ( \7604 , RIc0d9ce8_83);
xor \U$7510 ( \7605 , \7603 , \7604 );
buf \U$7511 ( \7606 , \7605 );
buf \U$7512 ( \7607 , \7606 );
nand \U$7513 ( \7608 , \7602 , \7607 );
buf \U$7514 ( \7609 , \7608 );
buf \U$7515 ( \7610 , \7609 );
nand \U$7516 ( \7611 , \7601 , \7610 );
buf \U$7517 ( \7612 , \7611 );
buf \U$7518 ( \7613 , \7203 );
not \U$7519 ( \7614 , \7613 );
buf \U$7520 ( \7615 , \1389 );
not \U$7521 ( \7616 , \7615 );
or \U$7522 ( \7617 , \7614 , \7616 );
buf \U$7523 ( \7618 , \921 );
buf \U$7524 ( \7619 , RIc0d7768_3);
buf \U$7525 ( \7620 , RIc0d9dd8_85);
xor \U$7526 ( \7621 , \7619 , \7620 );
buf \U$7527 ( \7622 , \7621 );
buf \U$7528 ( \7623 , \7622 );
nand \U$7529 ( \7624 , \7618 , \7623 );
buf \U$7530 ( \7625 , \7624 );
buf \U$7531 ( \7626 , \7625 );
nand \U$7532 ( \7627 , \7617 , \7626 );
buf \U$7533 ( \7628 , \7627 );
xor \U$7534 ( \7629 , \7612 , \7628 );
xor \U$7535 ( \7630 , \7596 , \7629 );
buf \U$7536 ( \7631 , \7630 );
xor \U$7537 ( \7632 , \7573 , \7631 );
buf \U$7538 ( \7633 , \7632 );
buf \U$7539 ( \7634 , \7633 );
xor \U$7540 ( \7635 , \7479 , \7634 );
buf \U$7541 ( \7636 , \7635 );
buf \U$7542 ( \7637 , \7636 );
xor \U$7543 ( \7638 , \7357 , \7637 );
xor \U$7544 ( \7639 , \7252 , \7303 );
and \U$7545 ( \7640 , \7639 , \7310 );
and \U$7546 ( \7641 , \7252 , \7303 );
or \U$7547 ( \7642 , \7640 , \7641 );
buf \U$7548 ( \7643 , \7642 );
buf \U$7549 ( \7644 , \7643 );
xor \U$7550 ( \7645 , \7008 , \7028 );
and \U$7551 ( \7646 , \7645 , \7061 );
and \U$7552 ( \7647 , \7008 , \7028 );
or \U$7553 ( \7648 , \7646 , \7647 );
buf \U$7554 ( \7649 , \7648 );
buf \U$7555 ( \7650 , \7649 );
xor \U$7556 ( \7651 , \7644 , \7650 );
xor \U$7557 ( \7652 , \6977 , \6998 );
and \U$7558 ( \7653 , \7652 , \7005 );
and \U$7559 ( \7654 , \6977 , \6998 );
or \U$7560 ( \7655 , \7653 , \7654 );
buf \U$7561 ( \7656 , \7655 );
buf \U$7562 ( \7657 , \7656 );
buf \U$7563 ( \7658 , \7059 );
not \U$7564 ( \7659 , \7658 );
buf \U$7565 ( \7660 , \7044 );
not \U$7566 ( \7661 , \7660 );
or \U$7567 ( \7662 , \7659 , \7661 );
buf \U$7568 ( \7663 , \7059 );
buf \U$7569 ( \7664 , \7044 );
or \U$7570 ( \7665 , \7663 , \7664 );
buf \U$7571 ( \7666 , \7034 );
nand \U$7572 ( \7667 , \7665 , \7666 );
buf \U$7573 ( \7668 , \7667 );
buf \U$7574 ( \7669 , \7668 );
nand \U$7575 ( \7670 , \7662 , \7669 );
buf \U$7576 ( \7671 , \7670 );
buf \U$7577 ( \7672 , \7671 );
xor \U$7578 ( \7673 , \7657 , \7672 );
xor \U$7579 ( \7674 , \7269 , \7286 );
and \U$7580 ( \7675 , \7674 , \7300 );
and \U$7581 ( \7676 , \7269 , \7286 );
or \U$7582 ( \7677 , \7675 , \7676 );
buf \U$7583 ( \7678 , \7677 );
buf \U$7584 ( \7679 , \7678 );
xor \U$7585 ( \7680 , \7118 , \7138 );
and \U$7586 ( \7681 , \7680 , \7148 );
and \U$7587 ( \7682 , \7118 , \7138 );
or \U$7588 ( \7683 , \7681 , \7682 );
buf \U$7589 ( \7684 , \7683 );
buf \U$7590 ( \7685 , \7684 );
xor \U$7591 ( \7686 , \7679 , \7685 );
xor \U$7592 ( \7687 , \7155 , \7172 );
and \U$7593 ( \7688 , \7687 , \7186 );
and \U$7594 ( \7689 , \7155 , \7172 );
or \U$7595 ( \7690 , \7688 , \7689 );
buf \U$7596 ( \7691 , \7690 );
buf \U$7597 ( \7692 , \7691 );
xor \U$7598 ( \7693 , \7686 , \7692 );
buf \U$7599 ( \7694 , \7693 );
buf \U$7600 ( \7695 , \7694 );
xor \U$7601 ( \7696 , \7673 , \7695 );
buf \U$7602 ( \7697 , \7696 );
buf \U$7603 ( \7698 , \7697 );
xor \U$7604 ( \7699 , \7651 , \7698 );
buf \U$7605 ( \7700 , \7699 );
buf \U$7606 ( \7701 , \7700 );
xor \U$7607 ( \7702 , \7638 , \7701 );
buf \U$7608 ( \7703 , \7702 );
buf \U$7609 ( \7704 , \7703 );
xor \U$7610 ( \7705 , \7351 , \7704 );
buf \U$7611 ( \7706 , \7705 );
buf \U$7612 ( \7707 , \7706 );
xor \U$7613 ( \7708 , \7067 , \7073 );
and \U$7614 ( \7709 , \7708 , \7326 );
and \U$7615 ( \7710 , \7067 , \7073 );
or \U$7616 ( \7711 , \7709 , \7710 );
buf \U$7617 ( \7712 , \7711 );
buf \U$7618 ( \7713 , \7712 );
or \U$7619 ( \7714 , \7707 , \7713 );
buf \U$7620 ( \7715 , \7714 );
buf \U$7621 ( \7716 , \7715 );
and \U$7622 ( \7717 , \6951 , \7338 , \7716 );
buf \U$7623 ( \7718 , \7717 );
buf \U$7624 ( \7719 , \7718 );
and \U$7625 ( \7720 , \6104 , \7719 );
buf \U$7626 ( \7721 , \7720 );
buf \U$7627 ( \7722 , \7721 );
buf \U$7628 ( \7723 , RIc0d80c8_23);
buf \U$7629 ( \7724 , RIc0d9478_65);
and \U$7630 ( \7725 , \7723 , \7724 );
buf \U$7631 ( \7726 , \7725 );
buf \U$7632 ( \7727 , \7726 );
buf \U$7633 ( \7728 , RIc0d7f60_20);
buf \U$7634 ( \7729 , RIc0d9568_67);
xor \U$7635 ( \7730 , \7728 , \7729 );
buf \U$7636 ( \7731 , \7730 );
buf \U$7637 ( \7732 , \7731 );
not \U$7638 ( \7733 , \7732 );
buf \U$7639 ( \7734 , \2900 );
not \U$7640 ( \7735 , \7734 );
or \U$7641 ( \7736 , \7733 , \7735 );
buf \U$7642 ( \7737 , RIc0d9568_67);
buf \U$7643 ( \7738 , RIc0d7ee8_19);
xnor \U$7644 ( \7739 , \7737 , \7738 );
buf \U$7645 ( \7740 , \7739 );
buf \U$7646 ( \7741 , \7740 );
not \U$7647 ( \7742 , \7741 );
buf \U$7648 ( \7743 , \686 );
nand \U$7649 ( \7744 , \7742 , \7743 );
buf \U$7650 ( \7745 , \7744 );
buf \U$7651 ( \7746 , \7745 );
nand \U$7652 ( \7747 , \7736 , \7746 );
buf \U$7653 ( \7748 , \7747 );
buf \U$7654 ( \7749 , \7748 );
xor \U$7655 ( \7750 , \7727 , \7749 );
buf \U$7656 ( \7751 , \1183 );
not \U$7657 ( \7752 , \7751 );
buf \U$7658 ( \7753 , \7752 );
buf \U$7659 ( \7754 , \7753 );
buf \U$7660 ( \7755 , RIc0d9a18_77);
buf \U$7661 ( \7756 , RIc0d7ab0_10);
xnor \U$7662 ( \7757 , \7755 , \7756 );
buf \U$7663 ( \7758 , \7757 );
buf \U$7664 ( \7759 , \7758 );
or \U$7665 ( \7760 , \7754 , \7759 );
buf \U$7666 ( \7761 , \1585 );
buf \U$7667 ( \7762 , RIc0d7a38_9);
buf \U$7668 ( \7763 , RIc0d9a18_77);
xnor \U$7669 ( \7764 , \7762 , \7763 );
buf \U$7670 ( \7765 , \7764 );
buf \U$7671 ( \7766 , \7765 );
or \U$7672 ( \7767 , \7761 , \7766 );
nand \U$7673 ( \7768 , \7760 , \7767 );
buf \U$7674 ( \7769 , \7768 );
buf \U$7675 ( \7770 , \7769 );
xor \U$7676 ( \7771 , \7750 , \7770 );
buf \U$7677 ( \7772 , \7771 );
buf \U$7678 ( \7773 , \7772 );
buf \U$7679 ( \7774 , \2815 );
buf \U$7680 ( \7775 , RIc0d7d80_16);
buf \U$7681 ( \7776 , RIc0d9748_71);
xnor \U$7682 ( \7777 , \7775 , \7776 );
buf \U$7683 ( \7778 , \7777 );
buf \U$7684 ( \7779 , \7778 );
or \U$7685 ( \7780 , \7774 , \7779 );
buf \U$7686 ( \7781 , \2927 );
not \U$7687 ( \7782 , \7781 );
buf \U$7688 ( \7783 , \7782 );
buf \U$7689 ( \7784 , \7783 );
xnor \U$7690 ( \7785 , RIc0d9748_71, RIc0d7d08_15);
buf \U$7691 ( \7786 , \7785 );
or \U$7692 ( \7787 , \7784 , \7786 );
nand \U$7693 ( \7788 , \7780 , \7787 );
buf \U$7694 ( \7789 , \7788 );
buf \U$7695 ( \7790 , \7789 );
buf \U$7696 ( \7791 , RIc0d8050_22);
buf \U$7697 ( \7792 , RIc0d9478_65);
xnor \U$7698 ( \7793 , \7791 , \7792 );
buf \U$7699 ( \7794 , \7793 );
buf \U$7700 ( \7795 , \7794 );
not \U$7701 ( \7796 , \7795 );
buf \U$7702 ( \7797 , \7796 );
buf \U$7703 ( \7798 , \7797 );
not \U$7704 ( \7799 , \7798 );
buf \U$7705 ( \7800 , \1225 );
not \U$7706 ( \7801 , \7800 );
or \U$7707 ( \7802 , \7799 , \7801 );
buf \U$7708 ( \7803 , \1229 );
buf \U$7709 ( \7804 , RIc0d9478_65);
buf \U$7710 ( \7805 , RIc0d7fd8_21);
xor \U$7711 ( \7806 , \7804 , \7805 );
buf \U$7712 ( \7807 , \7806 );
buf \U$7713 ( \7808 , \7807 );
nand \U$7714 ( \7809 , \7803 , \7808 );
buf \U$7715 ( \7810 , \7809 );
buf \U$7716 ( \7811 , \7810 );
nand \U$7717 ( \7812 , \7802 , \7811 );
buf \U$7718 ( \7813 , \7812 );
buf \U$7719 ( \7814 , \7813 );
xor \U$7720 ( \7815 , \7790 , \7814 );
buf \U$7721 ( \7816 , \1452 );
buf \U$7722 ( \7817 , RIc0d9658_69);
buf \U$7723 ( \7818 , RIc0d7e70_18);
not \U$7724 ( \7819 , \7818 );
buf \U$7725 ( \7820 , \7819 );
buf \U$7726 ( \7821 , \7820 );
and \U$7727 ( \7822 , \7817 , \7821 );
not \U$7728 ( \7823 , \7817 );
buf \U$7729 ( \7824 , RIc0d7e70_18);
and \U$7730 ( \7825 , \7823 , \7824 );
nor \U$7731 ( \7826 , \7822 , \7825 );
buf \U$7732 ( \7827 , \7826 );
buf \U$7733 ( \7828 , \7827 );
or \U$7734 ( \7829 , \7816 , \7828 );
buf \U$7735 ( \7830 , \1969 );
buf \U$7736 ( \7831 , RIc0d9658_69);
buf \U$7737 ( \7832 , RIc0d7df8_17);
not \U$7738 ( \7833 , \7832 );
buf \U$7739 ( \7834 , \7833 );
buf \U$7740 ( \7835 , \7834 );
and \U$7741 ( \7836 , \7831 , \7835 );
not \U$7742 ( \7837 , \7831 );
buf \U$7743 ( \7838 , RIc0d7df8_17);
and \U$7744 ( \7839 , \7837 , \7838 );
nor \U$7745 ( \7840 , \7836 , \7839 );
buf \U$7746 ( \7841 , \7840 );
buf \U$7747 ( \7842 , \7841 );
or \U$7748 ( \7843 , \7830 , \7842 );
nand \U$7749 ( \7844 , \7829 , \7843 );
buf \U$7750 ( \7845 , \7844 );
buf \U$7751 ( \7846 , \7845 );
xor \U$7752 ( \7847 , \7815 , \7846 );
buf \U$7753 ( \7848 , \7847 );
buf \U$7754 ( \7849 , \7848 );
xor \U$7755 ( \7850 , \7773 , \7849 );
buf \U$7756 ( \7851 , \3816 );
buf \U$7757 ( \7852 , RIc0d7ba0_12);
buf \U$7758 ( \7853 , RIc0d9928_75);
xnor \U$7759 ( \7854 , \7852 , \7853 );
buf \U$7760 ( \7855 , \7854 );
buf \U$7761 ( \7856 , \7855 );
or \U$7762 ( \7857 , \7851 , \7856 );
buf \U$7763 ( \7858 , \2372 );
buf \U$7764 ( \7859 , RIc0d7b28_11);
buf \U$7765 ( \7860 , RIc0d9928_75);
xnor \U$7766 ( \7861 , \7859 , \7860 );
buf \U$7767 ( \7862 , \7861 );
buf \U$7768 ( \7863 , \7862 );
or \U$7769 ( \7864 , \7858 , \7863 );
nand \U$7770 ( \7865 , \7857 , \7864 );
buf \U$7771 ( \7866 , \7865 );
buf \U$7772 ( \7867 , \7866 );
not \U$7773 ( \7868 , \7867 );
buf \U$7774 ( \7869 , RIc0d76f0_2);
buf \U$7775 ( \7870 , RIc0d9dd8_85);
xor \U$7776 ( \7871 , \7869 , \7870 );
buf \U$7777 ( \7872 , \7871 );
buf \U$7778 ( \7873 , \7872 );
not \U$7779 ( \7874 , \7873 );
buf \U$7780 ( \7875 , \1389 );
not \U$7781 ( \7876 , \7875 );
or \U$7782 ( \7877 , \7874 , \7876 );
buf \U$7783 ( \7878 , \921 );
buf \U$7784 ( \7879 , RIc0d7678_1);
buf \U$7785 ( \7880 , RIc0d9dd8_85);
xor \U$7786 ( \7881 , \7879 , \7880 );
buf \U$7787 ( \7882 , \7881 );
buf \U$7788 ( \7883 , \7882 );
nand \U$7789 ( \7884 , \7878 , \7883 );
buf \U$7790 ( \7885 , \7884 );
buf \U$7791 ( \7886 , \7885 );
nand \U$7792 ( \7887 , \7877 , \7886 );
buf \U$7793 ( \7888 , \7887 );
buf \U$7794 ( \7889 , RIc0d77e0_4);
buf \U$7795 ( \7890 , RIc0d9ce8_83);
xor \U$7796 ( \7891 , \7889 , \7890 );
buf \U$7797 ( \7892 , \7891 );
buf \U$7798 ( \7893 , \7892 );
not \U$7799 ( \7894 , \7893 );
buf \U$7800 ( \7895 , \574 );
not \U$7801 ( \7896 , \7895 );
or \U$7802 ( \7897 , \7894 , \7896 );
buf \U$7803 ( \7898 , RIc0d7768_3);
buf \U$7804 ( \7899 , RIc0d9ce8_83);
xnor \U$7805 ( \7900 , \7898 , \7899 );
buf \U$7806 ( \7901 , \7900 );
buf \U$7807 ( \7902 , \7901 );
not \U$7808 ( \7903 , \7902 );
buf \U$7809 ( \7904 , \584 );
nand \U$7810 ( \7905 , \7903 , \7904 );
buf \U$7811 ( \7906 , \7905 );
buf \U$7812 ( \7907 , \7906 );
nand \U$7813 ( \7908 , \7897 , \7907 );
buf \U$7814 ( \7909 , \7908 );
xnor \U$7815 ( \7910 , \7888 , \7909 );
buf \U$7816 ( \7911 , \7910 );
not \U$7817 ( \7912 , \7911 );
or \U$7818 ( \7913 , \7868 , \7912 );
buf \U$7819 ( \7914 , \7910 );
buf \U$7820 ( \7915 , \7866 );
or \U$7821 ( \7916 , \7914 , \7915 );
nand \U$7822 ( \7917 , \7913 , \7916 );
buf \U$7823 ( \7918 , \7917 );
buf \U$7824 ( \7919 , \7918 );
xor \U$7825 ( \7920 , \7850 , \7919 );
buf \U$7826 ( \7921 , \7920 );
buf \U$7827 ( \7922 , \7921 );
buf \U$7828 ( \7923 , \819 );
not \U$7829 ( \7924 , \7923 );
buf \U$7830 ( \7925 , \812 );
not \U$7831 ( \7926 , \7925 );
or \U$7832 ( \7927 , \7924 , \7926 );
buf \U$7833 ( \7928 , RIc0d9ec8_87);
nand \U$7834 ( \7929 , \7927 , \7928 );
buf \U$7835 ( \7930 , \7929 );
buf \U$7836 ( \7931 , RIc0d7c90_14);
buf \U$7837 ( \7932 , RIc0d9838_73);
xor \U$7838 ( \7933 , \7931 , \7932 );
buf \U$7839 ( \7934 , \7933 );
buf \U$7840 ( \7935 , \7934 );
not \U$7841 ( \7936 , \7935 );
buf \U$7842 ( \7937 , \1677 );
not \U$7843 ( \7938 , \7937 );
or \U$7844 ( \7939 , \7936 , \7938 );
buf \U$7845 ( \7940 , RIc0d7c18_13);
buf \U$7846 ( \7941 , RIc0d9838_73);
xnor \U$7847 ( \7942 , \7940 , \7941 );
buf \U$7848 ( \7943 , \7942 );
buf \U$7849 ( \7944 , \7943 );
not \U$7850 ( \7945 , \7944 );
buf \U$7851 ( \7946 , \1856 );
nand \U$7852 ( \7947 , \7945 , \7946 );
buf \U$7853 ( \7948 , \7947 );
buf \U$7854 ( \7949 , \7948 );
nand \U$7855 ( \7950 , \7939 , \7949 );
buf \U$7856 ( \7951 , \7950 );
buf \U$7857 ( \7952 , RIc0d79c0_8);
buf \U$7858 ( \7953 , RIc0d9b08_79);
xnor \U$7859 ( \7954 , \7952 , \7953 );
buf \U$7860 ( \7955 , \7954 );
buf \U$7861 ( \7956 , \7955 );
not \U$7862 ( \7957 , \7956 );
buf \U$7863 ( \7958 , \7957 );
buf \U$7864 ( \7959 , \7958 );
not \U$7865 ( \7960 , \7959 );
buf \U$7866 ( \7961 , \1351 );
not \U$7867 ( \7962 , \7961 );
or \U$7868 ( \7963 , \7960 , \7962 );
buf \U$7869 ( \7964 , RIc0d7948_7);
buf \U$7870 ( \7965 , RIc0d9b08_79);
xnor \U$7871 ( \7966 , \7964 , \7965 );
buf \U$7872 ( \7967 , \7966 );
buf \U$7873 ( \7968 , \7967 );
not \U$7874 ( \7969 , \7968 );
buf \U$7875 ( \7970 , \3985 );
nand \U$7876 ( \7971 , \7969 , \7970 );
buf \U$7877 ( \7972 , \7971 );
buf \U$7878 ( \7973 , \7972 );
nand \U$7879 ( \7974 , \7963 , \7973 );
buf \U$7880 ( \7975 , \7974 );
xor \U$7881 ( \7976 , \7951 , \7975 );
xor \U$7882 ( \7977 , \7930 , \7976 );
buf \U$7883 ( \7978 , \7977 );
buf \U$7884 ( \7979 , \6270 );
buf \U$7885 ( \7980 , \7564 );
or \U$7886 ( \7981 , \7979 , \7980 );
buf \U$7887 ( \7982 , \819 );
buf \U$7888 ( \7983 , \7556 );
or \U$7889 ( \7984 , \7982 , \7983 );
nand \U$7890 ( \7985 , \7981 , \7984 );
buf \U$7891 ( \7986 , \7985 );
buf \U$7892 ( \7987 , \7986 );
buf \U$7893 ( \7988 , \2769 );
buf \U$7894 ( \7989 , RIc0d78d0_6);
buf \U$7895 ( \7990 , RIc0d9bf8_81);
xnor \U$7896 ( \7991 , \7989 , \7990 );
buf \U$7897 ( \7992 , \7991 );
buf \U$7898 ( \7993 , \7992 );
or \U$7899 ( \7994 , \7988 , \7993 );
buf \U$7900 ( \7995 , \1610 );
buf \U$7901 ( \7996 , RIc0d9bf8_81);
not \U$7902 ( \7997 , \7996 );
buf \U$7903 ( \7998 , \7997 );
buf \U$7904 ( \7999 , \7998 );
buf \U$7905 ( \8000 , RIc0d7858_5);
and \U$7906 ( \8001 , \7999 , \8000 );
buf \U$7907 ( \8002 , \1990 );
buf \U$7908 ( \8003 , RIc0d9bf8_81);
and \U$7909 ( \8004 , \8002 , \8003 );
nor \U$7910 ( \8005 , \8001 , \8004 );
buf \U$7911 ( \8006 , \8005 );
buf \U$7912 ( \8007 , \8006 );
or \U$7913 ( \8008 , \7995 , \8007 );
nand \U$7914 ( \8009 , \7994 , \8008 );
buf \U$7915 ( \8010 , \8009 );
buf \U$7916 ( \8011 , \8010 );
xor \U$7917 ( \8012 , \7987 , \8011 );
buf \U$7918 ( \8013 , \7622 );
not \U$7919 ( \8014 , \8013 );
buf \U$7920 ( \8015 , \1389 );
not \U$7921 ( \8016 , \8015 );
or \U$7922 ( \8017 , \8014 , \8016 );
buf \U$7923 ( \8018 , \2960 );
buf \U$7924 ( \8019 , \7872 );
nand \U$7925 ( \8020 , \8018 , \8019 );
buf \U$7926 ( \8021 , \8020 );
buf \U$7927 ( \8022 , \8021 );
nand \U$7928 ( \8023 , \8017 , \8022 );
buf \U$7929 ( \8024 , \8023 );
buf \U$7930 ( \8025 , \8024 );
not \U$7931 ( \8026 , \8025 );
buf \U$7932 ( \8027 , \7498 );
not \U$7933 ( \8028 , \8027 );
buf \U$7934 ( \8029 , \1064 );
not \U$7935 ( \8030 , \8029 );
or \U$7936 ( \8031 , \8028 , \8030 );
buf \U$7937 ( \8032 , \7992 );
not \U$7938 ( \8033 , \8032 );
buf \U$7939 ( \8034 , \1078 );
nand \U$7940 ( \8035 , \8033 , \8034 );
buf \U$7941 ( \8036 , \8035 );
buf \U$7942 ( \8037 , \8036 );
nand \U$7943 ( \8038 , \8031 , \8037 );
buf \U$7944 ( \8039 , \8038 );
buf \U$7945 ( \8040 , \8039 );
not \U$7946 ( \8041 , \8040 );
or \U$7947 ( \8042 , \8026 , \8041 );
buf \U$7948 ( \8043 , \8039 );
buf \U$7949 ( \8044 , \8024 );
or \U$7950 ( \8045 , \8043 , \8044 );
buf \U$7951 ( \8046 , \7606 );
not \U$7952 ( \8047 , \8046 );
buf \U$7953 ( \8048 , \2088 );
not \U$7954 ( \8049 , \8048 );
or \U$7955 ( \8050 , \8047 , \8049 );
buf \U$7956 ( \8051 , \993 );
buf \U$7957 ( \8052 , \7892 );
nand \U$7958 ( \8053 , \8051 , \8052 );
buf \U$7959 ( \8054 , \8053 );
buf \U$7960 ( \8055 , \8054 );
nand \U$7961 ( \8056 , \8050 , \8055 );
buf \U$7962 ( \8057 , \8056 );
buf \U$7963 ( \8058 , \8057 );
nand \U$7964 ( \8059 , \8045 , \8058 );
buf \U$7965 ( \8060 , \8059 );
buf \U$7966 ( \8061 , \8060 );
nand \U$7967 ( \8062 , \8042 , \8061 );
buf \U$7968 ( \8063 , \8062 );
buf \U$7969 ( \8064 , \8063 );
xor \U$7970 ( \8065 , \8012 , \8064 );
buf \U$7971 ( \8066 , \8065 );
buf \U$7972 ( \8067 , \8066 );
xor \U$7973 ( \8068 , \7978 , \8067 );
buf \U$7974 ( \8069 , \7986 );
not \U$7975 ( \8070 , \8069 );
buf \U$7976 ( \8071 , \8070 );
buf \U$7977 ( \8072 , \8071 );
buf \U$7978 ( \8073 , \7628 );
buf \U$7979 ( \8074 , \7596 );
or \U$7980 ( \8075 , \8073 , \8074 );
buf \U$7981 ( \8076 , \7612 );
nand \U$7982 ( \8077 , \8075 , \8076 );
buf \U$7983 ( \8078 , \8077 );
buf \U$7984 ( \8079 , \8078 );
buf \U$7985 ( \8080 , \7628 );
buf \U$7986 ( \8081 , \7596 );
nand \U$7987 ( \8082 , \8080 , \8081 );
buf \U$7988 ( \8083 , \8082 );
buf \U$7989 ( \8084 , \8083 );
nand \U$7990 ( \8085 , \8079 , \8084 );
buf \U$7991 ( \8086 , \8085 );
buf \U$7992 ( \8087 , \8086 );
xor \U$7993 ( \8088 , \8072 , \8087 );
xor \U$7994 ( \8089 , \7531 , \7548 );
and \U$7995 ( \8090 , \8089 , \7569 );
and \U$7996 ( \8091 , \7531 , \7548 );
or \U$7997 ( \8092 , \8090 , \8091 );
buf \U$7998 ( \8093 , \8092 );
buf \U$7999 ( \8094 , \8093 );
and \U$8000 ( \8095 , \8088 , \8094 );
and \U$8001 ( \8096 , \8072 , \8087 );
or \U$8002 ( \8097 , \8095 , \8096 );
buf \U$8003 ( \8098 , \8097 );
buf \U$8004 ( \8099 , \8098 );
xor \U$8005 ( \8100 , \8068 , \8099 );
buf \U$8006 ( \8101 , \8100 );
buf \U$8007 ( \8102 , \8101 );
xor \U$8008 ( \8103 , \7922 , \8102 );
xor \U$8009 ( \8104 , \7488 , \7505 );
and \U$8010 ( \8105 , \8104 , \7507 );
and \U$8011 ( \8106 , \7488 , \7505 );
or \U$8012 ( \8107 , \8105 , \8106 );
buf \U$8013 ( \8108 , \8107 );
buf \U$8014 ( \8109 , \8108 );
xor \U$8015 ( \8110 , \7679 , \7685 );
and \U$8016 ( \8111 , \8110 , \7692 );
and \U$8017 ( \8112 , \7679 , \7685 );
or \U$8018 ( \8113 , \8111 , \8112 );
buf \U$8019 ( \8114 , \8113 );
buf \U$8020 ( \8115 , \8114 );
xor \U$8021 ( \8116 , \8109 , \8115 );
xor \U$8022 ( \8117 , \8072 , \8087 );
xor \U$8023 ( \8118 , \8117 , \8094 );
buf \U$8024 ( \8119 , \8118 );
buf \U$8025 ( \8120 , \8119 );
and \U$8026 ( \8121 , \8116 , \8120 );
and \U$8027 ( \8122 , \8109 , \8115 );
or \U$8028 ( \8123 , \8121 , \8122 );
buf \U$8029 ( \8124 , \8123 );
buf \U$8030 ( \8125 , \8124 );
xor \U$8031 ( \8126 , \8103 , \8125 );
buf \U$8032 ( \8127 , \8126 );
buf \U$8033 ( \8128 , \8127 );
xor \U$8034 ( \8129 , \7369 , \7411 );
and \U$8035 ( \8130 , \8129 , \7475 );
and \U$8036 ( \8131 , \7369 , \7411 );
or \U$8037 ( \8132 , \8130 , \8131 );
buf \U$8038 ( \8133 , \8132 );
buf \U$8039 ( \8134 , \8133 );
xor \U$8040 ( \8135 , \7510 , \7572 );
and \U$8041 ( \8136 , \8135 , \7631 );
and \U$8042 ( \8137 , \7510 , \7572 );
or \U$8043 ( \8138 , \8136 , \8137 );
buf \U$8044 ( \8139 , \8138 );
buf \U$8045 ( \8140 , \8139 );
xor \U$8046 ( \8141 , \8134 , \8140 );
xor \U$8047 ( \8142 , \7372 , \7390 );
and \U$8048 ( \8143 , \8142 , \7408 );
and \U$8049 ( \8144 , \7372 , \7390 );
or \U$8050 ( \8145 , \8143 , \8144 );
buf \U$8051 ( \8146 , \8145 );
buf \U$8052 ( \8147 , \8146 );
xor \U$8053 ( \8148 , \7429 , \7445 );
and \U$8054 ( \8149 , \8148 , \7472 );
and \U$8055 ( \8150 , \7429 , \7445 );
or \U$8056 ( \8151 , \8149 , \8150 );
buf \U$8057 ( \8152 , \8151 );
buf \U$8058 ( \8153 , \8152 );
xor \U$8059 ( \8154 , \8147 , \8153 );
buf \U$8060 ( \8155 , RIc0d8140_24);
buf \U$8061 ( \8156 , RIc0d9478_65);
and \U$8062 ( \8157 , \8155 , \8156 );
buf \U$8063 ( \8158 , \8157 );
buf \U$8064 ( \8159 , \8158 );
buf \U$8065 ( \8160 , \7401 );
not \U$8066 ( \8161 , \8160 );
buf \U$8067 ( \8162 , \1183 );
not \U$8068 ( \8163 , \8162 );
or \U$8069 ( \8164 , \8161 , \8163 );
buf \U$8070 ( \8165 , \7758 );
not \U$8071 ( \8166 , \8165 );
buf \U$8072 ( \8167 , \1588 );
nand \U$8073 ( \8168 , \8166 , \8167 );
buf \U$8074 ( \8169 , \8168 );
buf \U$8075 ( \8170 , \8169 );
nand \U$8076 ( \8171 , \8164 , \8170 );
buf \U$8077 ( \8172 , \8171 );
buf \U$8078 ( \8173 , \8172 );
xor \U$8079 ( \8174 , \8159 , \8173 );
buf \U$8080 ( \8175 , \393 );
buf \U$8081 ( \8176 , \7522 );
or \U$8082 ( \8177 , \8175 , \8176 );
not \U$8083 ( \8178 , \403 );
buf \U$8084 ( \8179 , \8178 );
buf \U$8085 ( \8180 , \7955 );
or \U$8086 ( \8181 , \8179 , \8180 );
nand \U$8087 ( \8182 , \8177 , \8181 );
buf \U$8088 ( \8183 , \8182 );
buf \U$8089 ( \8184 , \8183 );
xor \U$8090 ( \8185 , \8174 , \8184 );
buf \U$8091 ( \8186 , \8185 );
buf \U$8092 ( \8187 , \8186 );
xor \U$8093 ( \8188 , \8154 , \8187 );
buf \U$8094 ( \8189 , \8188 );
buf \U$8095 ( \8190 , \8189 );
and \U$8096 ( \8191 , \8141 , \8190 );
and \U$8097 ( \8192 , \8134 , \8140 );
or \U$8098 ( \8193 , \8191 , \8192 );
buf \U$8099 ( \8194 , \8193 );
buf \U$8100 ( \8195 , \8194 );
xor \U$8101 ( \8196 , \8147 , \8153 );
and \U$8102 ( \8197 , \8196 , \8187 );
and \U$8103 ( \8198 , \8147 , \8153 );
or \U$8104 ( \8199 , \8197 , \8198 );
buf \U$8105 ( \8200 , \8199 );
buf \U$8106 ( \8201 , \8200 );
buf \U$8107 ( \8202 , \7731 );
not \U$8108 ( \8203 , \8202 );
buf \U$8109 ( \8204 , \686 );
not \U$8110 ( \8205 , \8204 );
or \U$8111 ( \8206 , \8203 , \8205 );
buf \U$8112 ( \8207 , \1823 );
not \U$8113 ( \8208 , \8207 );
buf \U$8114 ( \8209 , \8208 );
buf \U$8115 ( \8210 , \8209 );
buf \U$8116 ( \8211 , \7381 );
or \U$8117 ( \8212 , \8210 , \8211 );
nand \U$8118 ( \8213 , \8206 , \8212 );
buf \U$8119 ( \8214 , \8213 );
buf \U$8120 ( \8215 , \8214 );
buf \U$8121 ( \8216 , \7541 );
not \U$8122 ( \8217 , \8216 );
buf \U$8123 ( \8218 , \2871 );
not \U$8124 ( \8219 , \8218 );
or \U$8125 ( \8220 , \8217 , \8219 );
buf \U$8126 ( \8221 , \2882 );
buf \U$8127 ( \8222 , \7934 );
nand \U$8128 ( \8223 , \8221 , \8222 );
buf \U$8129 ( \8224 , \8223 );
buf \U$8130 ( \8225 , \8224 );
nand \U$8131 ( \8226 , \8220 , \8225 );
buf \U$8132 ( \8227 , \8226 );
buf \U$8133 ( \8228 , \8227 );
xor \U$8134 ( \8229 , \8215 , \8228 );
buf \U$8135 ( \8230 , \1452 );
buf \U$8136 ( \8231 , \7440 );
or \U$8137 ( \8232 , \8230 , \8231 );
buf \U$8138 ( \8233 , \1969 );
buf \U$8139 ( \8234 , \7827 );
or \U$8140 ( \8235 , \8233 , \8234 );
nand \U$8141 ( \8236 , \8232 , \8235 );
buf \U$8142 ( \8237 , \8236 );
buf \U$8143 ( \8238 , \8237 );
xor \U$8144 ( \8239 , \8229 , \8238 );
buf \U$8145 ( \8240 , \8239 );
buf \U$8146 ( \8241 , \8240 );
buf \U$8147 ( \8242 , \7422 );
not \U$8148 ( \8243 , \8242 );
buf \U$8149 ( \8244 , \1263 );
not \U$8150 ( \8245 , \8244 );
or \U$8151 ( \8246 , \8243 , \8245 );
buf \U$8152 ( \8247 , \7778 );
not \U$8153 ( \8248 , \8247 );
buf \U$8154 ( \8249 , \2927 );
nand \U$8155 ( \8250 , \8248 , \8249 );
buf \U$8156 ( \8251 , \8250 );
buf \U$8157 ( \8252 , \8251 );
nand \U$8158 ( \8253 , \8246 , \8252 );
buf \U$8159 ( \8254 , \8253 );
buf \U$8160 ( \8255 , \8254 );
buf \U$8161 ( \8256 , \7590 );
not \U$8162 ( \8257 , \8256 );
buf \U$8163 ( \8258 , \1129 );
not \U$8164 ( \8259 , \8258 );
or \U$8165 ( \8260 , \8257 , \8259 );
buf \U$8166 ( \8261 , \7855 );
not \U$8167 ( \8262 , \8261 );
buf \U$8168 ( \8263 , \1143 );
nand \U$8169 ( \8264 , \8262 , \8263 );
buf \U$8170 ( \8265 , \8264 );
buf \U$8171 ( \8266 , \8265 );
nand \U$8172 ( \8267 , \8260 , \8266 );
buf \U$8173 ( \8268 , \8267 );
buf \U$8174 ( \8269 , \8268 );
xor \U$8175 ( \8270 , \8255 , \8269 );
buf \U$8176 ( \8271 , \1224 );
not \U$8177 ( \8272 , \8271 );
buf \U$8178 ( \8273 , \8272 );
buf \U$8179 ( \8274 , \8273 );
buf \U$8180 ( \8275 , \7467 );
or \U$8181 ( \8276 , \8274 , \8275 );
buf \U$8182 ( \8277 , \1232 );
buf \U$8183 ( \8278 , \7794 );
or \U$8184 ( \8279 , \8277 , \8278 );
nand \U$8185 ( \8280 , \8276 , \8279 );
buf \U$8186 ( \8281 , \8280 );
buf \U$8187 ( \8282 , \8281 );
xor \U$8188 ( \8283 , \8270 , \8282 );
buf \U$8189 ( \8284 , \8283 );
buf \U$8190 ( \8285 , \8284 );
or \U$8191 ( \8286 , \8241 , \8285 );
xor \U$8192 ( \8287 , \8039 , \8024 );
xor \U$8193 ( \8288 , \8287 , \8057 );
buf \U$8194 ( \8289 , \8288 );
nand \U$8195 ( \8290 , \8286 , \8289 );
buf \U$8196 ( \8291 , \8290 );
buf \U$8197 ( \8292 , \8291 );
buf \U$8198 ( \8293 , \8240 );
buf \U$8199 ( \8294 , \8284 );
nand \U$8200 ( \8295 , \8293 , \8294 );
buf \U$8201 ( \8296 , \8295 );
buf \U$8202 ( \8297 , \8296 );
nand \U$8203 ( \8298 , \8292 , \8297 );
buf \U$8204 ( \8299 , \8298 );
buf \U$8205 ( \8300 , \8299 );
xor \U$8206 ( \8301 , \8201 , \8300 );
xor \U$8207 ( \8302 , \8159 , \8173 );
and \U$8208 ( \8303 , \8302 , \8184 );
and \U$8209 ( \8304 , \8159 , \8173 );
or \U$8210 ( \8305 , \8303 , \8304 );
buf \U$8211 ( \8306 , \8305 );
buf \U$8212 ( \8307 , \8306 );
xor \U$8213 ( \8308 , \8255 , \8269 );
and \U$8214 ( \8309 , \8308 , \8282 );
and \U$8215 ( \8310 , \8255 , \8269 );
or \U$8216 ( \8311 , \8309 , \8310 );
buf \U$8217 ( \8312 , \8311 );
buf \U$8218 ( \8313 , \8312 );
xor \U$8219 ( \8314 , \8307 , \8313 );
xor \U$8220 ( \8315 , \8215 , \8228 );
and \U$8221 ( \8316 , \8315 , \8238 );
and \U$8222 ( \8317 , \8215 , \8228 );
or \U$8223 ( \8318 , \8316 , \8317 );
buf \U$8224 ( \8319 , \8318 );
buf \U$8225 ( \8320 , \8319 );
xor \U$8226 ( \8321 , \8314 , \8320 );
buf \U$8227 ( \8322 , \8321 );
buf \U$8228 ( \8323 , \8322 );
xor \U$8229 ( \8324 , \8301 , \8323 );
buf \U$8230 ( \8325 , \8324 );
buf \U$8231 ( \8326 , \8325 );
xor \U$8232 ( \8327 , \8195 , \8326 );
buf \U$8233 ( \8328 , \8288 );
not \U$8234 ( \8329 , \8328 );
buf \U$8235 ( \8330 , \8240 );
buf \U$8236 ( \8331 , \8284 );
not \U$8237 ( \8332 , \8331 );
xor \U$8238 ( \8333 , \8330 , \8332 );
buf \U$8239 ( \8334 , \8333 );
buf \U$8240 ( \8335 , \8334 );
not \U$8241 ( \8336 , \8335 );
or \U$8242 ( \8337 , \8329 , \8336 );
buf \U$8243 ( \8338 , \8334 );
buf \U$8244 ( \8339 , \8288 );
or \U$8245 ( \8340 , \8338 , \8339 );
nand \U$8246 ( \8341 , \8337 , \8340 );
buf \U$8247 ( \8342 , \8341 );
buf \U$8248 ( \8343 , \8342 );
xor \U$8249 ( \8344 , \7657 , \7672 );
and \U$8250 ( \8345 , \8344 , \7695 );
and \U$8251 ( \8346 , \7657 , \7672 );
or \U$8252 ( \8347 , \8345 , \8346 );
buf \U$8253 ( \8348 , \8347 );
buf \U$8254 ( \8349 , \8348 );
xor \U$8255 ( \8350 , \8343 , \8349 );
xor \U$8256 ( \8351 , \8109 , \8115 );
xor \U$8257 ( \8352 , \8351 , \8120 );
buf \U$8258 ( \8353 , \8352 );
buf \U$8259 ( \8354 , \8353 );
and \U$8260 ( \8355 , \8350 , \8354 );
and \U$8261 ( \8356 , \8343 , \8349 );
or \U$8262 ( \8357 , \8355 , \8356 );
buf \U$8263 ( \8358 , \8357 );
buf \U$8264 ( \8359 , \8358 );
xor \U$8265 ( \8360 , \8327 , \8359 );
buf \U$8266 ( \8361 , \8360 );
buf \U$8267 ( \8362 , \8361 );
xor \U$8268 ( \8363 , \8128 , \8362 );
xor \U$8269 ( \8364 , \7363 , \7478 );
and \U$8270 ( \8365 , \8364 , \7634 );
and \U$8271 ( \8366 , \7363 , \7478 );
or \U$8272 ( \8367 , \8365 , \8366 );
buf \U$8273 ( \8368 , \8367 );
buf \U$8274 ( \8369 , \8368 );
xor \U$8275 ( \8370 , \8134 , \8140 );
xor \U$8276 ( \8371 , \8370 , \8190 );
buf \U$8277 ( \8372 , \8371 );
buf \U$8278 ( \8373 , \8372 );
xor \U$8279 ( \8374 , \8369 , \8373 );
xor \U$8280 ( \8375 , \7644 , \7650 );
and \U$8281 ( \8376 , \8375 , \7698 );
and \U$8282 ( \8377 , \7644 , \7650 );
or \U$8283 ( \8378 , \8376 , \8377 );
buf \U$8284 ( \8379 , \8378 );
buf \U$8285 ( \8380 , \8379 );
and \U$8286 ( \8381 , \8374 , \8380 );
and \U$8287 ( \8382 , \8369 , \8373 );
or \U$8288 ( \8383 , \8381 , \8382 );
buf \U$8289 ( \8384 , \8383 );
buf \U$8290 ( \8385 , \8384 );
xor \U$8291 ( \8386 , \8363 , \8385 );
buf \U$8292 ( \8387 , \8386 );
buf \U$8293 ( \8388 , \8387 );
xor \U$8294 ( \8389 , \8343 , \8349 );
xor \U$8295 ( \8390 , \8389 , \8354 );
buf \U$8296 ( \8391 , \8390 );
buf \U$8297 ( \8392 , \8391 );
xor \U$8298 ( \8393 , \7357 , \7637 );
and \U$8299 ( \8394 , \8393 , \7701 );
and \U$8300 ( \8395 , \7357 , \7637 );
or \U$8301 ( \8396 , \8394 , \8395 );
buf \U$8302 ( \8397 , \8396 );
buf \U$8303 ( \8398 , \8397 );
xor \U$8304 ( \8399 , \8392 , \8398 );
xor \U$8305 ( \8400 , \8369 , \8373 );
xor \U$8306 ( \8401 , \8400 , \8380 );
buf \U$8307 ( \8402 , \8401 );
buf \U$8308 ( \8403 , \8402 );
and \U$8309 ( \8404 , \8399 , \8403 );
and \U$8310 ( \8405 , \8392 , \8398 );
or \U$8311 ( \8406 , \8404 , \8405 );
buf \U$8312 ( \8407 , \8406 );
buf \U$8313 ( \8408 , \8407 );
or \U$8314 ( \8409 , \8388 , \8408 );
buf \U$8315 ( \8410 , \8409 );
buf \U$8316 ( \8411 , \8410 );
not \U$8317 ( \8412 , \8411 );
buf \U$8318 ( \8413 , \7975 );
not \U$8319 ( \8414 , \8413 );
buf \U$8320 ( \8415 , \7951 );
not \U$8321 ( \8416 , \8415 );
or \U$8322 ( \8417 , \8414 , \8416 );
buf \U$8323 ( \8418 , \7951 );
buf \U$8324 ( \8419 , \7975 );
or \U$8325 ( \8420 , \8418 , \8419 );
buf \U$8326 ( \8421 , \7930 );
nand \U$8327 ( \8422 , \8420 , \8421 );
buf \U$8328 ( \8423 , \8422 );
buf \U$8329 ( \8424 , \8423 );
nand \U$8330 ( \8425 , \8417 , \8424 );
buf \U$8331 ( \8426 , \8425 );
buf \U$8332 ( \8427 , \8426 );
buf \U$8333 ( \8428 , \7785 );
not \U$8334 ( \8429 , \8428 );
buf \U$8335 ( \8430 , \8429 );
buf \U$8336 ( \8431 , \8430 );
not \U$8337 ( \8432 , \8431 );
buf \U$8338 ( \8433 , \2923 );
not \U$8339 ( \8434 , \8433 );
or \U$8340 ( \8435 , \8432 , \8434 );
buf \U$8341 ( \8436 , RIc0d7c90_14);
buf \U$8342 ( \8437 , RIc0d9748_71);
xnor \U$8343 ( \8438 , \8436 , \8437 );
buf \U$8344 ( \8439 , \8438 );
buf \U$8345 ( \8440 , \8439 );
not \U$8346 ( \8441 , \8440 );
buf \U$8347 ( \8442 , \1282 );
nand \U$8348 ( \8443 , \8441 , \8442 );
buf \U$8349 ( \8444 , \8443 );
buf \U$8350 ( \8445 , \8444 );
nand \U$8351 ( \8446 , \8435 , \8445 );
buf \U$8352 ( \8447 , \8446 );
buf \U$8353 ( \8448 , \8447 );
buf \U$8354 ( \8449 , \7807 );
not \U$8355 ( \8450 , \8449 );
buf \U$8356 ( \8451 , \3781 );
not \U$8357 ( \8452 , \8451 );
or \U$8358 ( \8453 , \8450 , \8452 );
buf \U$8359 ( \8454 , RIc0d7f60_20);
buf \U$8360 ( \8455 , RIc0d9478_65);
xnor \U$8361 ( \8456 , \8454 , \8455 );
buf \U$8362 ( \8457 , \8456 );
buf \U$8363 ( \8458 , \8457 );
not \U$8364 ( \8459 , \8458 );
buf \U$8365 ( \8460 , \1229 );
nand \U$8366 ( \8461 , \8459 , \8460 );
buf \U$8367 ( \8462 , \8461 );
buf \U$8368 ( \8463 , \8462 );
nand \U$8369 ( \8464 , \8453 , \8463 );
buf \U$8370 ( \8465 , \8464 );
buf \U$8371 ( \8466 , \8465 );
xor \U$8372 ( \8467 , \8448 , \8466 );
buf \U$8373 ( \8468 , \1739 );
buf \U$8374 ( \8469 , \7901 );
or \U$8375 ( \8470 , \8468 , \8469 );
buf \U$8376 ( \8471 , \996 );
buf \U$8377 ( \8472 , RIc0d76f0_2);
buf \U$8378 ( \8473 , RIc0d9ce8_83);
xnor \U$8379 ( \8474 , \8472 , \8473 );
buf \U$8380 ( \8475 , \8474 );
buf \U$8381 ( \8476 , \8475 );
or \U$8382 ( \8477 , \8471 , \8476 );
nand \U$8383 ( \8478 , \8470 , \8477 );
buf \U$8384 ( \8479 , \8478 );
buf \U$8385 ( \8480 , \8479 );
xor \U$8386 ( \8481 , \8467 , \8480 );
buf \U$8387 ( \8482 , \8481 );
buf \U$8388 ( \8483 , \8482 );
xor \U$8389 ( \8484 , \8427 , \8483 );
buf \U$8390 ( \8485 , \4904 );
buf \U$8391 ( \8486 , \7740 );
or \U$8392 ( \8487 , \8485 , \8486 );
buf \U$8393 ( \8488 , \6437 );
buf \U$8394 ( \8489 , RIc0d7e70_18);
buf \U$8395 ( \8490 , RIc0d9568_67);
xnor \U$8396 ( \8491 , \8489 , \8490 );
buf \U$8397 ( \8492 , \8491 );
buf \U$8398 ( \8493 , \8492 );
or \U$8399 ( \8494 , \8488 , \8493 );
nand \U$8400 ( \8495 , \8487 , \8494 );
buf \U$8401 ( \8496 , \8495 );
buf \U$8402 ( \8497 , \8496 );
buf \U$8403 ( \8498 , \779 );
buf \U$8404 ( \8499 , \7943 );
or \U$8405 ( \8500 , \8498 , \8499 );
buf \U$8406 ( \8501 , \795 );
buf \U$8407 ( \8502 , RIc0d7ba0_12);
buf \U$8408 ( \8503 , RIc0d9838_73);
xor \U$8409 ( \8504 , \8502 , \8503 );
buf \U$8410 ( \8505 , \8504 );
buf \U$8411 ( \8506 , \8505 );
not \U$8412 ( \8507 , \8506 );
buf \U$8413 ( \8508 , \8507 );
buf \U$8414 ( \8509 , \8508 );
or \U$8415 ( \8510 , \8501 , \8509 );
nand \U$8416 ( \8511 , \8500 , \8510 );
buf \U$8417 ( \8512 , \8511 );
buf \U$8418 ( \8513 , \8512 );
xor \U$8419 ( \8514 , \8497 , \8513 );
buf \U$8420 ( \8515 , \1452 );
buf \U$8421 ( \8516 , \7841 );
or \U$8422 ( \8517 , \8515 , \8516 );
buf \U$8423 ( \8518 , \1969 );
buf \U$8424 ( \8519 , RIc0d9658_69);
buf \U$8425 ( \8520 , \1744 );
and \U$8426 ( \8521 , \8519 , \8520 );
not \U$8427 ( \8522 , \8519 );
buf \U$8428 ( \8523 , RIc0d7d80_16);
and \U$8429 ( \8524 , \8522 , \8523 );
nor \U$8430 ( \8525 , \8521 , \8524 );
buf \U$8431 ( \8526 , \8525 );
buf \U$8432 ( \8527 , \8526 );
or \U$8433 ( \8528 , \8518 , \8527 );
nand \U$8434 ( \8529 , \8517 , \8528 );
buf \U$8435 ( \8530 , \8529 );
buf \U$8436 ( \8531 , \8530 );
xor \U$8437 ( \8532 , \8514 , \8531 );
buf \U$8438 ( \8533 , \8532 );
buf \U$8439 ( \8534 , \8533 );
xor \U$8440 ( \8535 , \8484 , \8534 );
buf \U$8441 ( \8536 , \8535 );
buf \U$8442 ( \8537 , \8536 );
xor \U$8443 ( \8538 , \7978 , \8067 );
and \U$8444 ( \8539 , \8538 , \8099 );
and \U$8445 ( \8540 , \7978 , \8067 );
or \U$8446 ( \8541 , \8539 , \8540 );
buf \U$8447 ( \8542 , \8541 );
buf \U$8448 ( \8543 , \8542 );
xor \U$8449 ( \8544 , \8537 , \8543 );
buf \U$8450 ( \8545 , \7862 );
not \U$8451 ( \8546 , \8545 );
buf \U$8452 ( \8547 , \8546 );
buf \U$8453 ( \8548 , \8547 );
not \U$8454 ( \8549 , \8548 );
buf \U$8455 ( \8550 , \1129 );
not \U$8456 ( \8551 , \8550 );
or \U$8457 ( \8552 , \8549 , \8551 );
buf \U$8458 ( \8553 , RIc0d7ab0_10);
buf \U$8459 ( \8554 , RIc0d9928_75);
xnor \U$8460 ( \8555 , \8553 , \8554 );
buf \U$8461 ( \8556 , \8555 );
buf \U$8462 ( \8557 , \8556 );
not \U$8463 ( \8558 , \8557 );
buf \U$8464 ( \8559 , \1143 );
nand \U$8465 ( \8560 , \8558 , \8559 );
buf \U$8466 ( \8561 , \8560 );
buf \U$8467 ( \8562 , \8561 );
nand \U$8468 ( \8563 , \8552 , \8562 );
buf \U$8469 ( \8564 , \8563 );
buf \U$8470 ( \8565 , \8564 );
buf \U$8471 ( \8566 , \7765 );
not \U$8472 ( \8567 , \8566 );
buf \U$8473 ( \8568 , \8567 );
buf \U$8474 ( \8569 , \8568 );
not \U$8475 ( \8570 , \8569 );
buf \U$8476 ( \8571 , \1183 );
not \U$8477 ( \8572 , \8571 );
or \U$8478 ( \8573 , \8570 , \8572 );
buf \U$8479 ( \8574 , RIc0d79c0_8);
buf \U$8480 ( \8575 , RIc0d9a18_77);
xnor \U$8481 ( \8576 , \8574 , \8575 );
buf \U$8482 ( \8577 , \8576 );
buf \U$8483 ( \8578 , \8577 );
not \U$8484 ( \8579 , \8578 );
buf \U$8485 ( \8580 , \3742 );
nand \U$8486 ( \8581 , \8579 , \8580 );
buf \U$8487 ( \8582 , \8581 );
buf \U$8488 ( \8583 , \8582 );
nand \U$8489 ( \8584 , \8573 , \8583 );
buf \U$8490 ( \8585 , \8584 );
buf \U$8491 ( \8586 , \8585 );
xor \U$8492 ( \8587 , \8565 , \8586 );
buf \U$8493 ( \8588 , \2769 );
buf \U$8494 ( \8589 , \8006 );
or \U$8495 ( \8590 , \8588 , \8589 );
buf \U$8496 ( \8591 , \1610 );
buf \U$8497 ( \8592 , RIc0d77e0_4);
buf \U$8498 ( \8593 , RIc0d9bf8_81);
xor \U$8499 ( \8594 , \8592 , \8593 );
buf \U$8500 ( \8595 , \8594 );
buf \U$8501 ( \8596 , \8595 );
not \U$8502 ( \8597 , \8596 );
buf \U$8503 ( \8598 , \8597 );
buf \U$8504 ( \8599 , \8598 );
or \U$8505 ( \8600 , \8591 , \8599 );
nand \U$8506 ( \8601 , \8590 , \8600 );
buf \U$8507 ( \8602 , \8601 );
buf \U$8508 ( \8603 , \8602 );
xor \U$8509 ( \8604 , \8587 , \8603 );
buf \U$8510 ( \8605 , \8604 );
buf \U$8511 ( \8606 , \8605 );
buf \U$8512 ( \8607 , RIc0d8050_22);
buf \U$8513 ( \8608 , RIc0d9478_65);
and \U$8514 ( \8609 , \8607 , \8608 );
buf \U$8515 ( \8610 , \8609 );
buf \U$8516 ( \8611 , \8610 );
buf \U$8517 ( \8612 , \7882 );
not \U$8518 ( \8613 , \8612 );
buf \U$8519 ( \8614 , \6029 );
not \U$8520 ( \8615 , \8614 );
or \U$8521 ( \8616 , \8613 , \8615 );
buf \U$8522 ( \8617 , \2960 );
buf \U$8523 ( \8618 , RIc0d9dd8_85);
nand \U$8524 ( \8619 , \8617 , \8618 );
buf \U$8525 ( \8620 , \8619 );
buf \U$8526 ( \8621 , \8620 );
nand \U$8527 ( \8622 , \8616 , \8621 );
buf \U$8528 ( \8623 , \8622 );
buf \U$8529 ( \8624 , \8623 );
not \U$8530 ( \8625 , \8624 );
buf \U$8531 ( \8626 , \8625 );
buf \U$8532 ( \8627 , \8626 );
xor \U$8533 ( \8628 , \8611 , \8627 );
buf \U$8534 ( \8629 , \393 );
buf \U$8535 ( \8630 , \7967 );
or \U$8536 ( \8631 , \8629 , \8630 );
buf \U$8537 ( \8632 , \8178 );
buf \U$8538 ( \8633 , RIc0d78d0_6);
buf \U$8539 ( \8634 , RIc0d9b08_79);
xor \U$8540 ( \8635 , \8633 , \8634 );
buf \U$8541 ( \8636 , \8635 );
buf \U$8542 ( \8637 , \8636 );
not \U$8543 ( \8638 , \8637 );
buf \U$8544 ( \8639 , \8638 );
buf \U$8545 ( \8640 , \8639 );
or \U$8546 ( \8641 , \8632 , \8640 );
nand \U$8547 ( \8642 , \8631 , \8641 );
buf \U$8548 ( \8643 , \8642 );
buf \U$8549 ( \8644 , \8643 );
xor \U$8550 ( \8645 , \8628 , \8644 );
buf \U$8551 ( \8646 , \8645 );
buf \U$8552 ( \8647 , \8646 );
xor \U$8553 ( \8648 , \8606 , \8647 );
xor \U$8554 ( \8649 , \8307 , \8313 );
and \U$8555 ( \8650 , \8649 , \8320 );
and \U$8556 ( \8651 , \8307 , \8313 );
or \U$8557 ( \8652 , \8650 , \8651 );
buf \U$8558 ( \8653 , \8652 );
buf \U$8559 ( \8654 , \8653 );
xor \U$8560 ( \8655 , \8648 , \8654 );
buf \U$8561 ( \8656 , \8655 );
buf \U$8562 ( \8657 , \8656 );
xor \U$8563 ( \8658 , \8544 , \8657 );
buf \U$8564 ( \8659 , \8658 );
buf \U$8565 ( \8660 , \8659 );
xor \U$8566 ( \8661 , \7987 , \8011 );
and \U$8567 ( \8662 , \8661 , \8064 );
and \U$8568 ( \8663 , \7987 , \8011 );
or \U$8569 ( \8664 , \8662 , \8663 );
buf \U$8570 ( \8665 , \8664 );
buf \U$8571 ( \8666 , \8665 );
xor \U$8572 ( \8667 , \7727 , \7749 );
and \U$8573 ( \8668 , \8667 , \7770 );
and \U$8574 ( \8669 , \7727 , \7749 );
or \U$8575 ( \8670 , \8668 , \8669 );
buf \U$8576 ( \8671 , \8670 );
buf \U$8577 ( \8672 , \8671 );
buf \U$8578 ( \8673 , \7888 );
not \U$8579 ( \8674 , \8673 );
buf \U$8580 ( \8675 , \7866 );
not \U$8581 ( \8676 , \8675 );
or \U$8582 ( \8677 , \8674 , \8676 );
buf \U$8583 ( \8678 , \7866 );
buf \U$8584 ( \8679 , \7888 );
or \U$8585 ( \8680 , \8678 , \8679 );
buf \U$8586 ( \8681 , \7909 );
nand \U$8587 ( \8682 , \8680 , \8681 );
buf \U$8588 ( \8683 , \8682 );
buf \U$8589 ( \8684 , \8683 );
nand \U$8590 ( \8685 , \8677 , \8684 );
buf \U$8591 ( \8686 , \8685 );
buf \U$8592 ( \8687 , \8686 );
xor \U$8593 ( \8688 , \8672 , \8687 );
xor \U$8594 ( \8689 , \7790 , \7814 );
and \U$8595 ( \8690 , \8689 , \7846 );
and \U$8596 ( \8691 , \7790 , \7814 );
or \U$8597 ( \8692 , \8690 , \8691 );
buf \U$8598 ( \8693 , \8692 );
buf \U$8599 ( \8694 , \8693 );
xor \U$8600 ( \8695 , \8688 , \8694 );
buf \U$8601 ( \8696 , \8695 );
buf \U$8602 ( \8697 , \8696 );
xor \U$8603 ( \8698 , \8666 , \8697 );
xor \U$8604 ( \8699 , \7773 , \7849 );
and \U$8605 ( \8700 , \8699 , \7919 );
and \U$8606 ( \8701 , \7773 , \7849 );
or \U$8607 ( \8702 , \8700 , \8701 );
buf \U$8608 ( \8703 , \8702 );
buf \U$8609 ( \8704 , \8703 );
xor \U$8610 ( \8705 , \8698 , \8704 );
buf \U$8611 ( \8706 , \8705 );
buf \U$8612 ( \8707 , \8706 );
xor \U$8613 ( \8708 , \8201 , \8300 );
and \U$8614 ( \8709 , \8708 , \8323 );
and \U$8615 ( \8710 , \8201 , \8300 );
or \U$8616 ( \8711 , \8709 , \8710 );
buf \U$8617 ( \8712 , \8711 );
buf \U$8618 ( \8713 , \8712 );
xor \U$8619 ( \8714 , \8707 , \8713 );
xor \U$8620 ( \8715 , \7922 , \8102 );
and \U$8621 ( \8716 , \8715 , \8125 );
and \U$8622 ( \8717 , \7922 , \8102 );
or \U$8623 ( \8718 , \8716 , \8717 );
buf \U$8624 ( \8719 , \8718 );
buf \U$8625 ( \8720 , \8719 );
xor \U$8626 ( \8721 , \8714 , \8720 );
buf \U$8627 ( \8722 , \8721 );
buf \U$8628 ( \8723 , \8722 );
xor \U$8629 ( \8724 , \8660 , \8723 );
xor \U$8630 ( \8725 , \8195 , \8326 );
and \U$8631 ( \8726 , \8725 , \8359 );
and \U$8632 ( \8727 , \8195 , \8326 );
or \U$8633 ( \8728 , \8726 , \8727 );
buf \U$8634 ( \8729 , \8728 );
buf \U$8635 ( \8730 , \8729 );
xor \U$8636 ( \8731 , \8724 , \8730 );
buf \U$8637 ( \8732 , \8731 );
buf \U$8638 ( \8733 , \8732 );
xor \U$8639 ( \8734 , \8128 , \8362 );
and \U$8640 ( \8735 , \8734 , \8385 );
and \U$8641 ( \8736 , \8128 , \8362 );
or \U$8642 ( \8737 , \8735 , \8736 );
buf \U$8643 ( \8738 , \8737 );
buf \U$8644 ( \8739 , \8738 );
nor \U$8645 ( \8740 , \8733 , \8739 );
buf \U$8646 ( \8741 , \8740 );
buf \U$8647 ( \8742 , \8741 );
nor \U$8648 ( \8743 , \8412 , \8742 );
buf \U$8649 ( \8744 , \8743 );
buf \U$8650 ( \8745 , \8744 );
xor \U$8651 ( \8746 , \8392 , \8398 );
xor \U$8652 ( \8747 , \8746 , \8403 );
buf \U$8653 ( \8748 , \8747 );
buf \U$8654 ( \8749 , \8748 );
xor \U$8655 ( \8750 , \7344 , \7350 );
and \U$8656 ( \8751 , \8750 , \7704 );
and \U$8657 ( \8752 , \7344 , \7350 );
or \U$8658 ( \8753 , \8751 , \8752 );
buf \U$8659 ( \8754 , \8753 );
buf \U$8660 ( \8755 , \8754 );
or \U$8661 ( \8756 , \8749 , \8755 );
buf \U$8662 ( \8757 , \8756 );
buf \U$8663 ( \8758 , \8757 );
xor \U$8664 ( \8759 , \8660 , \8723 );
and \U$8665 ( \8760 , \8759 , \8730 );
and \U$8666 ( \8761 , \8660 , \8723 );
or \U$8667 ( \8762 , \8760 , \8761 );
buf \U$8668 ( \8763 , \8762 );
buf \U$8669 ( \8764 , \8763 );
xor \U$8670 ( \8765 , \8707 , \8713 );
and \U$8671 ( \8766 , \8765 , \8720 );
and \U$8672 ( \8767 , \8707 , \8713 );
or \U$8673 ( \8768 , \8766 , \8767 );
buf \U$8674 ( \8769 , \8768 );
buf \U$8675 ( \8770 , \8769 );
xor \U$8676 ( \8771 , \8448 , \8466 );
and \U$8677 ( \8772 , \8771 , \8480 );
and \U$8678 ( \8773 , \8448 , \8466 );
or \U$8679 ( \8774 , \8772 , \8773 );
buf \U$8680 ( \8775 , \8774 );
buf \U$8681 ( \8776 , \8505 );
not \U$8682 ( \8777 , \8776 );
buf \U$8683 ( \8778 , \2871 );
not \U$8684 ( \8779 , \8778 );
or \U$8685 ( \8780 , \8777 , \8779 );
buf \U$8686 ( \8781 , \792 );
buf \U$8687 ( \8782 , RIc0d7b28_11);
buf \U$8688 ( \8783 , RIc0d9838_73);
xor \U$8689 ( \8784 , \8782 , \8783 );
buf \U$8690 ( \8785 , \8784 );
buf \U$8691 ( \8786 , \8785 );
nand \U$8692 ( \8787 , \8781 , \8786 );
buf \U$8693 ( \8788 , \8787 );
buf \U$8694 ( \8789 , \8788 );
nand \U$8695 ( \8790 , \8780 , \8789 );
buf \U$8696 ( \8791 , \8790 );
buf \U$8697 ( \8792 , \8636 );
not \U$8698 ( \8793 , \8792 );
buf \U$8699 ( \8794 , \1351 );
not \U$8700 ( \8795 , \8794 );
or \U$8701 ( \8796 , \8793 , \8795 );
buf \U$8702 ( \8797 , \1026 );
buf \U$8703 ( \8798 , RIc0d7858_5);
buf \U$8704 ( \8799 , RIc0d9b08_79);
xor \U$8705 ( \8800 , \8798 , \8799 );
buf \U$8706 ( \8801 , \8800 );
buf \U$8707 ( \8802 , \8801 );
nand \U$8708 ( \8803 , \8797 , \8802 );
buf \U$8709 ( \8804 , \8803 );
buf \U$8710 ( \8805 , \8804 );
nand \U$8711 ( \8806 , \8796 , \8805 );
buf \U$8712 ( \8807 , \8806 );
xor \U$8713 ( \8808 , \8791 , \8807 );
buf \U$8714 ( \8809 , \8595 );
not \U$8715 ( \8810 , \8809 );
buf \U$8716 ( \8811 , \1064 );
not \U$8717 ( \8812 , \8811 );
or \U$8718 ( \8813 , \8810 , \8812 );
buf \U$8719 ( \8814 , \1078 );
buf \U$8720 ( \8815 , RIc0d7768_3);
buf \U$8721 ( \8816 , RIc0d9bf8_81);
xor \U$8722 ( \8817 , \8815 , \8816 );
buf \U$8723 ( \8818 , \8817 );
buf \U$8724 ( \8819 , \8818 );
nand \U$8725 ( \8820 , \8814 , \8819 );
buf \U$8726 ( \8821 , \8820 );
buf \U$8727 ( \8822 , \8821 );
nand \U$8728 ( \8823 , \8813 , \8822 );
buf \U$8729 ( \8824 , \8823 );
xor \U$8730 ( \8825 , \8808 , \8824 );
xor \U$8731 ( \8826 , \8775 , \8825 );
buf \U$8732 ( \8827 , RIc0d7a38_9);
buf \U$8733 ( \8828 , RIc0d9928_75);
xor \U$8734 ( \8829 , \8827 , \8828 );
buf \U$8735 ( \8830 , \8829 );
buf \U$8736 ( \8831 , \8830 );
not \U$8737 ( \8832 , \8831 );
buf \U$8738 ( \8833 , \1143 );
not \U$8739 ( \8834 , \8833 );
or \U$8740 ( \8835 , \8832 , \8834 );
buf \U$8741 ( \8836 , \3816 );
buf \U$8742 ( \8837 , \8556 );
or \U$8743 ( \8838 , \8836 , \8837 );
nand \U$8744 ( \8839 , \8835 , \8838 );
buf \U$8745 ( \8840 , \8839 );
buf \U$8746 ( \8841 , RIc0d7678_1);
buf \U$8747 ( \8842 , RIc0d9ce8_83);
xor \U$8748 ( \8843 , \8841 , \8842 );
buf \U$8749 ( \8844 , \8843 );
buf \U$8750 ( \8845 , \8844 );
not \U$8751 ( \8846 , \8845 );
buf \U$8752 ( \8847 , \993 );
not \U$8753 ( \8848 , \8847 );
or \U$8754 ( \8849 , \8846 , \8848 );
buf \U$8755 ( \8850 , \8475 );
not \U$8756 ( \8851 , \8850 );
buf \U$8757 ( \8852 , \574 );
nand \U$8758 ( \8853 , \8851 , \8852 );
buf \U$8759 ( \8854 , \8853 );
buf \U$8760 ( \8855 , \8854 );
nand \U$8761 ( \8856 , \8849 , \8855 );
buf \U$8762 ( \8857 , \8856 );
xor \U$8763 ( \8858 , \8840 , \8857 );
buf \U$8764 ( \8859 , \2963 );
not \U$8765 ( \8860 , \8859 );
buf \U$8766 ( \8861 , \5305 );
not \U$8767 ( \8862 , \8861 );
buf \U$8768 ( \8863 , \8862 );
buf \U$8769 ( \8864 , \8863 );
not \U$8770 ( \8865 , \8864 );
or \U$8771 ( \8866 , \8860 , \8865 );
buf \U$8772 ( \8867 , RIc0d9dd8_85);
nand \U$8773 ( \8868 , \8866 , \8867 );
buf \U$8774 ( \8869 , \8868 );
xor \U$8775 ( \8870 , \8858 , \8869 );
xor \U$8776 ( \8871 , \8826 , \8870 );
and \U$8777 ( \8872 , \7804 , \7805 );
buf \U$8778 ( \8873 , \8872 );
buf \U$8779 ( \8874 , \8873 );
buf \U$8780 ( \8875 , \8492 );
not \U$8781 ( \8876 , \8875 );
buf \U$8782 ( \8877 , \8876 );
buf \U$8783 ( \8878 , \8877 );
not \U$8784 ( \8879 , \8878 );
buf \U$8785 ( \8880 , \4907 );
not \U$8786 ( \8881 , \8880 );
or \U$8787 ( \8882 , \8879 , \8881 );
buf \U$8788 ( \8883 , \686 );
buf \U$8789 ( \8884 , RIc0d7df8_17);
buf \U$8790 ( \8885 , RIc0d9568_67);
xor \U$8791 ( \8886 , \8884 , \8885 );
buf \U$8792 ( \8887 , \8886 );
buf \U$8793 ( \8888 , \8887 );
nand \U$8794 ( \8889 , \8883 , \8888 );
buf \U$8795 ( \8890 , \8889 );
buf \U$8796 ( \8891 , \8890 );
nand \U$8797 ( \8892 , \8882 , \8891 );
buf \U$8798 ( \8893 , \8892 );
buf \U$8799 ( \8894 , \8893 );
xor \U$8800 ( \8895 , \8874 , \8894 );
buf \U$8801 ( \8896 , \7753 );
buf \U$8802 ( \8897 , \8577 );
or \U$8803 ( \8898 , \8896 , \8897 );
buf \U$8804 ( \8899 , \1193 );
buf \U$8805 ( \8900 , RIc0d7948_7);
buf \U$8806 ( \8901 , RIc0d9a18_77);
xnor \U$8807 ( \8902 , \8900 , \8901 );
buf \U$8808 ( \8903 , \8902 );
buf \U$8809 ( \8904 , \8903 );
or \U$8810 ( \8905 , \8899 , \8904 );
nand \U$8811 ( \8906 , \8898 , \8905 );
buf \U$8812 ( \8907 , \8906 );
buf \U$8813 ( \8908 , \8907 );
xor \U$8814 ( \8909 , \8895 , \8908 );
buf \U$8815 ( \8910 , \8909 );
buf \U$8816 ( \8911 , \8910 );
xor \U$8817 ( \8912 , \8611 , \8627 );
and \U$8818 ( \8913 , \8912 , \8644 );
and \U$8819 ( \8914 , \8611 , \8627 );
or \U$8820 ( \8915 , \8913 , \8914 );
buf \U$8821 ( \8916 , \8915 );
buf \U$8822 ( \8917 , \8916 );
xor \U$8823 ( \8918 , \8911 , \8917 );
buf \U$8824 ( \8919 , \8273 );
buf \U$8825 ( \8920 , \8457 );
or \U$8826 ( \8921 , \8919 , \8920 );
buf \U$8827 ( \8922 , \1232 );
buf \U$8828 ( \8923 , RIc0d7ee8_19);
buf \U$8829 ( \8924 , RIc0d9478_65);
xnor \U$8830 ( \8925 , \8923 , \8924 );
buf \U$8831 ( \8926 , \8925 );
buf \U$8832 ( \8927 , \8926 );
or \U$8833 ( \8928 , \8922 , \8927 );
nand \U$8834 ( \8929 , \8921 , \8928 );
buf \U$8835 ( \8930 , \8929 );
buf \U$8836 ( \8931 , \8930 );
buf \U$8837 ( \8932 , \4868 );
buf \U$8838 ( \8933 , \8439 );
or \U$8839 ( \8934 , \8932 , \8933 );
buf \U$8840 ( \8935 , \1279 );
buf \U$8841 ( \8936 , RIc0d7c18_13);
buf \U$8842 ( \8937 , RIc0d9748_71);
xnor \U$8843 ( \8938 , \8936 , \8937 );
buf \U$8844 ( \8939 , \8938 );
buf \U$8845 ( \8940 , \8939 );
or \U$8846 ( \8941 , \8935 , \8940 );
nand \U$8847 ( \8942 , \8934 , \8941 );
buf \U$8848 ( \8943 , \8942 );
buf \U$8849 ( \8944 , \8943 );
xor \U$8850 ( \8945 , \8931 , \8944 );
buf \U$8851 ( \8946 , \1452 );
buf \U$8852 ( \8947 , \8526 );
or \U$8853 ( \8948 , \8946 , \8947 );
buf \U$8854 ( \8949 , \1969 );
buf \U$8855 ( \8950 , RIc0d7d08_15);
buf \U$8856 ( \8951 , RIc0d9658_69);
xnor \U$8857 ( \8952 , \8950 , \8951 );
buf \U$8858 ( \8953 , \8952 );
buf \U$8859 ( \8954 , \8953 );
or \U$8860 ( \8955 , \8949 , \8954 );
nand \U$8861 ( \8956 , \8948 , \8955 );
buf \U$8862 ( \8957 , \8956 );
buf \U$8863 ( \8958 , \8957 );
xor \U$8864 ( \8959 , \8945 , \8958 );
buf \U$8865 ( \8960 , \8959 );
buf \U$8866 ( \8961 , \8960 );
xor \U$8867 ( \8962 , \8918 , \8961 );
buf \U$8868 ( \8963 , \8962 );
xor \U$8869 ( \8964 , \8606 , \8647 );
and \U$8870 ( \8965 , \8964 , \8654 );
and \U$8871 ( \8966 , \8606 , \8647 );
or \U$8872 ( \8967 , \8965 , \8966 );
buf \U$8873 ( \8968 , \8967 );
xor \U$8874 ( \8969 , \8963 , \8968 );
xor \U$8875 ( \8970 , \8871 , \8969 );
buf \U$8876 ( \8971 , \8970 );
xor \U$8877 ( \8972 , \8770 , \8971 );
xor \U$8878 ( \8973 , \8672 , \8687 );
and \U$8879 ( \8974 , \8973 , \8694 );
and \U$8880 ( \8975 , \8672 , \8687 );
or \U$8881 ( \8976 , \8974 , \8975 );
buf \U$8882 ( \8977 , \8976 );
buf \U$8883 ( \8978 , \8977 );
buf \U$8884 ( \8979 , \8623 );
xor \U$8885 ( \8980 , \8565 , \8586 );
and \U$8886 ( \8981 , \8980 , \8603 );
and \U$8887 ( \8982 , \8565 , \8586 );
or \U$8888 ( \8983 , \8981 , \8982 );
buf \U$8889 ( \8984 , \8983 );
buf \U$8890 ( \8985 , \8984 );
xor \U$8891 ( \8986 , \8979 , \8985 );
xor \U$8892 ( \8987 , \8497 , \8513 );
and \U$8893 ( \8988 , \8987 , \8531 );
and \U$8894 ( \8989 , \8497 , \8513 );
or \U$8895 ( \8990 , \8988 , \8989 );
buf \U$8896 ( \8991 , \8990 );
buf \U$8897 ( \8992 , \8991 );
xor \U$8898 ( \8993 , \8986 , \8992 );
buf \U$8899 ( \8994 , \8993 );
buf \U$8900 ( \8995 , \8994 );
xor \U$8901 ( \8996 , \8978 , \8995 );
xor \U$8902 ( \8997 , \8427 , \8483 );
and \U$8903 ( \8998 , \8997 , \8534 );
and \U$8904 ( \8999 , \8427 , \8483 );
or \U$8905 ( \9000 , \8998 , \8999 );
buf \U$8906 ( \9001 , \9000 );
buf \U$8907 ( \9002 , \9001 );
xor \U$8908 ( \9003 , \8996 , \9002 );
buf \U$8909 ( \9004 , \9003 );
buf \U$8910 ( \9005 , \9004 );
xor \U$8911 ( \9006 , \8666 , \8697 );
and \U$8912 ( \9007 , \9006 , \8704 );
and \U$8913 ( \9008 , \8666 , \8697 );
or \U$8914 ( \9009 , \9007 , \9008 );
buf \U$8915 ( \9010 , \9009 );
buf \U$8916 ( \9011 , \9010 );
xor \U$8917 ( \9012 , \9005 , \9011 );
xor \U$8918 ( \9013 , \8537 , \8543 );
and \U$8919 ( \9014 , \9013 , \8657 );
and \U$8920 ( \9015 , \8537 , \8543 );
or \U$8921 ( \9016 , \9014 , \9015 );
buf \U$8922 ( \9017 , \9016 );
buf \U$8923 ( \9018 , \9017 );
xor \U$8924 ( \9019 , \9012 , \9018 );
buf \U$8925 ( \9020 , \9019 );
buf \U$8926 ( \9021 , \9020 );
xor \U$8927 ( \9022 , \8972 , \9021 );
buf \U$8928 ( \9023 , \9022 );
buf \U$8929 ( \9024 , \9023 );
or \U$8930 ( \9025 , \8764 , \9024 );
buf \U$8931 ( \9026 , \9025 );
buf \U$8932 ( \9027 , \9026 );
and \U$8933 ( \9028 , \8745 , \8758 , \9027 );
buf \U$8934 ( \9029 , \9028 );
buf \U$8935 ( \9030 , \9029 );
and \U$8936 ( \9031 , \7722 , \9030 );
buf \U$8937 ( \9032 , \9031 );
buf \U$8938 ( \9033 , \9032 );
xor \U$8939 ( \9034 , \9005 , \9011 );
and \U$8940 ( \9035 , \9034 , \9018 );
and \U$8941 ( \9036 , \9005 , \9011 );
or \U$8942 ( \9037 , \9035 , \9036 );
buf \U$8943 ( \9038 , \9037 );
buf \U$8944 ( \9039 , \9038 );
xor \U$8945 ( \9040 , \8775 , \8825 );
xor \U$8946 ( \9041 , \9040 , \8870 );
and \U$8947 ( \9042 , \8963 , \9041 );
xor \U$8948 ( \9043 , \8775 , \8825 );
xor \U$8949 ( \9044 , \9043 , \8870 );
and \U$8950 ( \9045 , \8968 , \9044 );
and \U$8951 ( \9046 , \8963 , \8968 );
or \U$8952 ( \9047 , \9042 , \9045 , \9046 );
buf \U$8953 ( \9048 , \9047 );
xor \U$8954 ( \9049 , \9039 , \9048 );
buf \U$8955 ( \9050 , RIc0d7f60_20);
buf \U$8956 ( \9051 , RIc0d9478_65);
and \U$8957 ( \9052 , \9050 , \9051 );
buf \U$8958 ( \9053 , \9052 );
buf \U$8959 ( \9054 , \9053 );
buf \U$8960 ( \9055 , \8939 );
not \U$8961 ( \9056 , \9055 );
buf \U$8962 ( \9057 , \9056 );
buf \U$8963 ( \9058 , \9057 );
not \U$8964 ( \9059 , \9058 );
buf \U$8965 ( \9060 , \1263 );
not \U$8966 ( \9061 , \9060 );
or \U$8967 ( \9062 , \9059 , \9061 );
buf \U$8968 ( \9063 , \1282 );
buf \U$8969 ( \9064 , RIc0d7ba0_12);
buf \U$8970 ( \9065 , RIc0d9748_71);
xor \U$8971 ( \9066 , \9064 , \9065 );
buf \U$8972 ( \9067 , \9066 );
buf \U$8973 ( \9068 , \9067 );
nand \U$8974 ( \9069 , \9063 , \9068 );
buf \U$8975 ( \9070 , \9069 );
buf \U$8976 ( \9071 , \9070 );
nand \U$8977 ( \9072 , \9062 , \9071 );
buf \U$8978 ( \9073 , \9072 );
buf \U$8979 ( \9074 , \9073 );
not \U$8980 ( \9075 , \9074 );
buf \U$8981 ( \9076 , \9075 );
buf \U$8982 ( \9077 , \9076 );
xor \U$8983 ( \9078 , \9054 , \9077 );
xor \U$8984 ( \9079 , \8874 , \8894 );
and \U$8985 ( \9080 , \9079 , \8908 );
and \U$8986 ( \9081 , \8874 , \8894 );
or \U$8987 ( \9082 , \9080 , \9081 );
buf \U$8988 ( \9083 , \9082 );
buf \U$8989 ( \9084 , \9083 );
xor \U$8990 ( \9085 , \9078 , \9084 );
buf \U$8991 ( \9086 , \9085 );
xor \U$8992 ( \9087 , \8979 , \8985 );
and \U$8993 ( \9088 , \9087 , \8992 );
and \U$8994 ( \9089 , \8979 , \8985 );
or \U$8995 ( \9090 , \9088 , \9089 );
buf \U$8996 ( \9091 , \9090 );
xor \U$8997 ( \9092 , \9086 , \9091 );
xor \U$8998 ( \9093 , \8775 , \8825 );
and \U$8999 ( \9094 , \9093 , \8870 );
and \U$9000 ( \9095 , \8775 , \8825 );
or \U$9001 ( \9096 , \9094 , \9095 );
xor \U$9002 ( \9097 , \9092 , \9096 );
xor \U$9003 ( \9098 , \8978 , \8995 );
and \U$9004 ( \9099 , \9098 , \9002 );
and \U$9005 ( \9100 , \8978 , \8995 );
or \U$9006 ( \9101 , \9099 , \9100 );
buf \U$9007 ( \9102 , \9101 );
xor \U$9008 ( \9103 , \8791 , \8807 );
and \U$9009 ( \9104 , \9103 , \8824 );
and \U$9010 ( \9105 , \8791 , \8807 );
or \U$9011 ( \9106 , \9104 , \9105 );
buf \U$9012 ( \9107 , \9106 );
xor \U$9013 ( \9108 , \8840 , \8857 );
and \U$9014 ( \9109 , \9108 , \8869 );
and \U$9015 ( \9110 , \8840 , \8857 );
or \U$9016 ( \9111 , \9109 , \9110 );
buf \U$9017 ( \9112 , \9111 );
xor \U$9018 ( \9113 , \9107 , \9112 );
xor \U$9019 ( \9114 , \8931 , \8944 );
and \U$9020 ( \9115 , \9114 , \8958 );
and \U$9021 ( \9116 , \8931 , \8944 );
or \U$9022 ( \9117 , \9115 , \9116 );
buf \U$9023 ( \9118 , \9117 );
buf \U$9024 ( \9119 , \9118 );
xor \U$9025 ( \9120 , \9113 , \9119 );
buf \U$9026 ( \9121 , \9120 );
buf \U$9027 ( \9122 , \9121 );
xor \U$9028 ( \9123 , \8911 , \8917 );
and \U$9029 ( \9124 , \9123 , \8961 );
and \U$9030 ( \9125 , \8911 , \8917 );
or \U$9031 ( \9126 , \9124 , \9125 );
buf \U$9032 ( \9127 , \9126 );
buf \U$9033 ( \9128 , \9127 );
xor \U$9034 ( \9129 , \9122 , \9128 );
buf \U$9035 ( \9130 , \8926 );
not \U$9036 ( \9131 , \9130 );
buf \U$9037 ( \9132 , \9131 );
buf \U$9038 ( \9133 , \9132 );
not \U$9039 ( \9134 , \9133 );
buf \U$9040 ( \9135 , \1225 );
not \U$9041 ( \9136 , \9135 );
or \U$9042 ( \9137 , \9134 , \9136 );
buf \U$9043 ( \9138 , \1705 );
buf \U$9044 ( \9139 , RIc0d9478_65);
buf \U$9045 ( \9140 , RIc0d7e70_18);
xor \U$9046 ( \9141 , \9139 , \9140 );
buf \U$9047 ( \9142 , \9141 );
buf \U$9048 ( \9143 , \9142 );
nand \U$9049 ( \9144 , \9138 , \9143 );
buf \U$9050 ( \9145 , \9144 );
buf \U$9051 ( \9146 , \9145 );
nand \U$9052 ( \9147 , \9137 , \9146 );
buf \U$9053 ( \9148 , \9147 );
buf \U$9054 ( \9149 , \8887 );
not \U$9055 ( \9150 , \9149 );
buf \U$9056 ( \9151 , \1823 );
not \U$9057 ( \9152 , \9151 );
or \U$9058 ( \9153 , \9150 , \9152 );
buf \U$9059 ( \9154 , \686 );
buf \U$9060 ( \9155 , RIc0d7d80_16);
buf \U$9061 ( \9156 , RIc0d9568_67);
xor \U$9062 ( \9157 , \9155 , \9156 );
buf \U$9063 ( \9158 , \9157 );
buf \U$9064 ( \9159 , \9158 );
nand \U$9065 ( \9160 , \9154 , \9159 );
buf \U$9066 ( \9161 , \9160 );
buf \U$9067 ( \9162 , \9161 );
nand \U$9068 ( \9163 , \9153 , \9162 );
buf \U$9069 ( \9164 , \9163 );
xor \U$9070 ( \9165 , \9148 , \9164 );
buf \U$9071 ( \9166 , RIc0d7c90_14);
buf \U$9072 ( \9167 , RIc0d9658_69);
xor \U$9073 ( \9168 , \9166 , \9167 );
buf \U$9074 ( \9169 , \9168 );
buf \U$9075 ( \9170 , \9169 );
not \U$9076 ( \9171 , \9170 );
buf \U$9077 ( \9172 , \874 );
not \U$9078 ( \9173 , \9172 );
or \U$9079 ( \9174 , \9171 , \9173 );
buf \U$9080 ( \9175 , \8953 );
not \U$9081 ( \9176 , \9175 );
buf \U$9082 ( \9177 , \4692 );
nand \U$9083 ( \9178 , \9176 , \9177 );
buf \U$9084 ( \9179 , \9178 );
buf \U$9085 ( \9180 , \9179 );
nand \U$9086 ( \9181 , \9174 , \9180 );
buf \U$9087 ( \9182 , \9181 );
xnor \U$9088 ( \9183 , \9165 , \9182 );
buf \U$9089 ( \9184 , \9183 );
not \U$9090 ( \9185 , \9184 );
buf \U$9091 ( \9186 , \9185 );
buf \U$9092 ( \9187 , \9186 );
not \U$9093 ( \9188 , \9187 );
buf \U$9094 ( \9189 , \8903 );
not \U$9095 ( \9190 , \9189 );
buf \U$9096 ( \9191 , \9190 );
buf \U$9097 ( \9192 , \9191 );
not \U$9098 ( \9193 , \9192 );
buf \U$9099 ( \9194 , \1432 );
not \U$9100 ( \9195 , \9194 );
or \U$9101 ( \9196 , \9193 , \9195 );
buf \U$9102 ( \9197 , \1588 );
buf \U$9103 ( \9198 , RIc0d78d0_6);
buf \U$9104 ( \9199 , RIc0d9a18_77);
xor \U$9105 ( \9200 , \9198 , \9199 );
buf \U$9106 ( \9201 , \9200 );
buf \U$9107 ( \9202 , \9201 );
nand \U$9108 ( \9203 , \9197 , \9202 );
buf \U$9109 ( \9204 , \9203 );
buf \U$9110 ( \9205 , \9204 );
nand \U$9111 ( \9206 , \9196 , \9205 );
buf \U$9112 ( \9207 , \9206 );
buf \U$9113 ( \9208 , \8818 );
not \U$9114 ( \9209 , \9208 );
buf \U$9115 ( \9210 , \2766 );
not \U$9116 ( \9211 , \9210 );
or \U$9117 ( \9212 , \9209 , \9211 );
buf \U$9118 ( \9213 , RIc0d76f0_2);
buf \U$9119 ( \9214 , RIc0d9bf8_81);
xnor \U$9120 ( \9215 , \9213 , \9214 );
buf \U$9121 ( \9216 , \9215 );
buf \U$9122 ( \9217 , \9216 );
not \U$9123 ( \9218 , \9217 );
buf \U$9124 ( \9219 , \1078 );
nand \U$9125 ( \9220 , \9218 , \9219 );
buf \U$9126 ( \9221 , \9220 );
buf \U$9127 ( \9222 , \9221 );
nand \U$9128 ( \9223 , \9212 , \9222 );
buf \U$9129 ( \9224 , \9223 );
xor \U$9130 ( \9225 , \9207 , \9224 );
buf \U$9131 ( \9226 , \8801 );
not \U$9132 ( \9227 , \9226 );
buf \U$9133 ( \9228 , \1351 );
not \U$9134 ( \9229 , \9228 );
or \U$9135 ( \9230 , \9227 , \9229 );
buf \U$9136 ( \9231 , RIc0d77e0_4);
buf \U$9137 ( \9232 , RIc0d9b08_79);
xnor \U$9138 ( \9233 , \9231 , \9232 );
buf \U$9139 ( \9234 , \9233 );
buf \U$9140 ( \9235 , \9234 );
not \U$9141 ( \9236 , \9235 );
buf \U$9142 ( \9237 , \403 );
nand \U$9143 ( \9238 , \9236 , \9237 );
buf \U$9144 ( \9239 , \9238 );
buf \U$9145 ( \9240 , \9239 );
nand \U$9146 ( \9241 , \9230 , \9240 );
buf \U$9147 ( \9242 , \9241 );
xnor \U$9148 ( \9243 , \9225 , \9242 );
buf \U$9149 ( \9244 , \9243 );
not \U$9150 ( \9245 , \9244 );
buf \U$9151 ( \9246 , \9245 );
buf \U$9152 ( \9247 , \9246 );
buf \U$9153 ( \9248 , \8830 );
not \U$9154 ( \9249 , \9248 );
buf \U$9155 ( \9250 , \1556 );
not \U$9156 ( \9251 , \9250 );
or \U$9157 ( \9252 , \9249 , \9251 );
buf \U$9158 ( \9253 , \1565 );
buf \U$9159 ( \9254 , RIc0d79c0_8);
buf \U$9160 ( \9255 , RIc0d9928_75);
xor \U$9161 ( \9256 , \9254 , \9255 );
buf \U$9162 ( \9257 , \9256 );
buf \U$9163 ( \9258 , \9257 );
nand \U$9164 ( \9259 , \9253 , \9258 );
buf \U$9165 ( \9260 , \9259 );
buf \U$9166 ( \9261 , \9260 );
nand \U$9167 ( \9262 , \9252 , \9261 );
buf \U$9168 ( \9263 , \9262 );
buf \U$9169 ( \9264 , \9263 );
buf \U$9170 ( \9265 , \8785 );
not \U$9171 ( \9266 , \9265 );
buf \U$9172 ( \9267 , \776 );
not \U$9173 ( \9268 , \9267 );
or \U$9174 ( \9269 , \9266 , \9268 );
buf \U$9175 ( \9270 , RIc0d7ab0_10);
buf \U$9176 ( \9271 , RIc0d9838_73);
xnor \U$9177 ( \9272 , \9270 , \9271 );
buf \U$9178 ( \9273 , \9272 );
buf \U$9179 ( \9274 , \9273 );
not \U$9180 ( \9275 , \9274 );
buf \U$9181 ( \9276 , \2882 );
nand \U$9182 ( \9277 , \9275 , \9276 );
buf \U$9183 ( \9278 , \9277 );
buf \U$9184 ( \9279 , \9278 );
nand \U$9185 ( \9280 , \9269 , \9279 );
buf \U$9186 ( \9281 , \9280 );
buf \U$9187 ( \9282 , \9281 );
xor \U$9188 ( \9283 , \9264 , \9282 );
buf \U$9189 ( \9284 , \1739 );
buf \U$9190 ( \9285 , \8844 );
not \U$9191 ( \9286 , \9285 );
buf \U$9192 ( \9287 , \9286 );
buf \U$9193 ( \9288 , \9287 );
or \U$9194 ( \9289 , \9284 , \9288 );
buf \U$9195 ( \9290 , \996 );
buf \U$9196 ( \9291 , \1050 );
or \U$9197 ( \9292 , \9290 , \9291 );
nand \U$9198 ( \9293 , \9289 , \9292 );
buf \U$9199 ( \9294 , \9293 );
buf \U$9200 ( \9295 , \9294 );
xor \U$9201 ( \9296 , \9283 , \9295 );
buf \U$9202 ( \9297 , \9296 );
buf \U$9203 ( \9298 , \9297 );
xnor \U$9204 ( \9299 , \9247 , \9298 );
buf \U$9205 ( \9300 , \9299 );
buf \U$9206 ( \9301 , \9300 );
not \U$9207 ( \9302 , \9301 );
or \U$9208 ( \9303 , \9188 , \9302 );
buf \U$9209 ( \9304 , \9300 );
buf \U$9210 ( \9305 , \9186 );
or \U$9211 ( \9306 , \9304 , \9305 );
nand \U$9212 ( \9307 , \9303 , \9306 );
buf \U$9213 ( \9308 , \9307 );
buf \U$9214 ( \9309 , \9308 );
xor \U$9215 ( \9310 , \9129 , \9309 );
buf \U$9216 ( \9311 , \9310 );
xor \U$9217 ( \9312 , \9102 , \9311 );
xor \U$9218 ( \9313 , \9097 , \9312 );
buf \U$9219 ( \9314 , \9313 );
and \U$9220 ( \9315 , \9049 , \9314 );
and \U$9221 ( \9316 , \9039 , \9048 );
or \U$9222 ( \9317 , \9315 , \9316 );
buf \U$9223 ( \9318 , \9317 );
buf \U$9224 ( \9319 , \9318 );
xor \U$9225 ( \9320 , \9086 , \9091 );
and \U$9226 ( \9321 , \9320 , \9096 );
and \U$9227 ( \9322 , \9086 , \9091 );
or \U$9228 ( \9323 , \9321 , \9322 );
buf \U$9229 ( \9324 , \403 );
not \U$9230 ( \9325 , \9324 );
buf \U$9231 ( \9326 , RIc0d7768_3);
buf \U$9232 ( \9327 , RIc0d9b08_79);
xor \U$9233 ( \9328 , \9326 , \9327 );
buf \U$9234 ( \9329 , \9328 );
buf \U$9235 ( \9330 , \9329 );
not \U$9236 ( \9331 , \9330 );
or \U$9237 ( \9332 , \9325 , \9331 );
buf \U$9238 ( \9333 , \393 );
buf \U$9239 ( \9334 , \9234 );
or \U$9240 ( \9335 , \9333 , \9334 );
nand \U$9241 ( \9336 , \9332 , \9335 );
buf \U$9242 ( \9337 , \9336 );
xor \U$9243 ( \9338 , \9073 , \9337 );
buf \U$9244 ( \9339 , \2769 );
buf \U$9245 ( \9340 , \9216 );
or \U$9246 ( \9341 , \9339 , \9340 );
buf \U$9247 ( \9342 , \1610 );
buf \U$9248 ( \9343 , RIc0d7678_1);
buf \U$9249 ( \9344 , RIc0d9bf8_81);
xnor \U$9250 ( \9345 , \9343 , \9344 );
buf \U$9251 ( \9346 , \9345 );
buf \U$9252 ( \9347 , \9346 );
or \U$9253 ( \9348 , \9342 , \9347 );
nand \U$9254 ( \9349 , \9341 , \9348 );
buf \U$9255 ( \9350 , \9349 );
xor \U$9256 ( \9351 , \9338 , \9350 );
xor \U$9257 ( \9352 , \9054 , \9077 );
and \U$9258 ( \9353 , \9352 , \9084 );
and \U$9259 ( \9354 , \9054 , \9077 );
or \U$9260 ( \9355 , \9353 , \9354 );
buf \U$9261 ( \9356 , \9355 );
xor \U$9262 ( \9357 , \9107 , \9112 );
and \U$9263 ( \9358 , \9357 , \9119 );
and \U$9264 ( \9359 , \9107 , \9112 );
or \U$9265 ( \9360 , \9358 , \9359 );
buf \U$9266 ( \9361 , \9360 );
xor \U$9267 ( \9362 , \9356 , \9361 );
xor \U$9268 ( \9363 , \9351 , \9362 );
xor \U$9269 ( \9364 , \9323 , \9363 );
buf \U$9270 ( \9365 , \9186 );
not \U$9271 ( \9366 , \9365 );
buf \U$9272 ( \9367 , \9246 );
not \U$9273 ( \9368 , \9367 );
or \U$9274 ( \9369 , \9366 , \9368 );
buf \U$9275 ( \9370 , \9243 );
buf \U$9276 ( \9371 , \9183 );
nand \U$9277 ( \9372 , \9370 , \9371 );
buf \U$9278 ( \9373 , \9372 );
buf \U$9279 ( \9374 , \9373 );
buf \U$9280 ( \9375 , \9297 );
nand \U$9281 ( \9376 , \9374 , \9375 );
buf \U$9282 ( \9377 , \9376 );
buf \U$9283 ( \9378 , \9377 );
nand \U$9284 ( \9379 , \9369 , \9378 );
buf \U$9285 ( \9380 , \9379 );
buf \U$9286 ( \9381 , \9380 );
buf \U$9287 ( \9382 , \9148 );
buf \U$9288 ( \9383 , \9164 );
or \U$9289 ( \9384 , \9382 , \9383 );
buf \U$9290 ( \9385 , \9182 );
nand \U$9291 ( \9386 , \9384 , \9385 );
buf \U$9292 ( \9387 , \9386 );
buf \U$9293 ( \9388 , \9387 );
buf \U$9294 ( \9389 , \9148 );
buf \U$9295 ( \9390 , \9164 );
nand \U$9296 ( \9391 , \9389 , \9390 );
buf \U$9297 ( \9392 , \9391 );
buf \U$9298 ( \9393 , \9392 );
nand \U$9299 ( \9394 , \9388 , \9393 );
buf \U$9300 ( \9395 , \9394 );
buf \U$9301 ( \9396 , \9395 );
xor \U$9302 ( \9397 , \9264 , \9282 );
and \U$9303 ( \9398 , \9397 , \9295 );
and \U$9304 ( \9399 , \9264 , \9282 );
or \U$9305 ( \9400 , \9398 , \9399 );
buf \U$9306 ( \9401 , \9400 );
buf \U$9307 ( \9402 , \9401 );
xor \U$9308 ( \9403 , \9396 , \9402 );
buf \U$9309 ( \9404 , \9224 );
not \U$9310 ( \9405 , \9404 );
buf \U$9311 ( \9406 , \9207 );
not \U$9312 ( \9407 , \9406 );
or \U$9313 ( \9408 , \9405 , \9407 );
buf \U$9314 ( \9409 , \9207 );
buf \U$9315 ( \9410 , \9224 );
or \U$9316 ( \9411 , \9409 , \9410 );
buf \U$9317 ( \9412 , \9242 );
nand \U$9318 ( \9413 , \9411 , \9412 );
buf \U$9319 ( \9414 , \9413 );
buf \U$9320 ( \9415 , \9414 );
nand \U$9321 ( \9416 , \9408 , \9415 );
buf \U$9322 ( \9417 , \9416 );
buf \U$9323 ( \9418 , \9417 );
xor \U$9324 ( \9419 , \9403 , \9418 );
buf \U$9325 ( \9420 , \9419 );
buf \U$9326 ( \9421 , \9420 );
xor \U$9327 ( \9422 , \9381 , \9421 );
buf \U$9328 ( \9423 , RIc0d7ee8_19);
buf \U$9329 ( \9424 , RIc0d9478_65);
and \U$9330 ( \9425 , \9423 , \9424 );
buf \U$9331 ( \9426 , \9425 );
buf \U$9332 ( \9427 , \9158 );
not \U$9333 ( \9428 , \9427 );
buf \U$9334 ( \9429 , \2900 );
not \U$9335 ( \9430 , \9429 );
or \U$9336 ( \9431 , \9428 , \9430 );
buf \U$9337 ( \9432 , \686 );
buf \U$9338 ( \9433 , RIc0d7d08_15);
buf \U$9339 ( \9434 , RIc0d9568_67);
xor \U$9340 ( \9435 , \9433 , \9434 );
buf \U$9341 ( \9436 , \9435 );
buf \U$9342 ( \9437 , \9436 );
nand \U$9343 ( \9438 , \9432 , \9437 );
buf \U$9344 ( \9439 , \9438 );
buf \U$9345 ( \9440 , \9439 );
nand \U$9346 ( \9441 , \9431 , \9440 );
buf \U$9347 ( \9442 , \9441 );
xor \U$9348 ( \9443 , \9426 , \9442 );
buf \U$9349 ( \9444 , \9201 );
not \U$9350 ( \9445 , \9444 );
buf \U$9351 ( \9446 , \1432 );
not \U$9352 ( \9447 , \9446 );
or \U$9353 ( \9448 , \9445 , \9447 );
buf \U$9354 ( \9449 , \3742 );
buf \U$9355 ( \9450 , RIc0d7858_5);
buf \U$9356 ( \9451 , RIc0d9a18_77);
xor \U$9357 ( \9452 , \9450 , \9451 );
buf \U$9358 ( \9453 , \9452 );
buf \U$9359 ( \9454 , \9453 );
nand \U$9360 ( \9455 , \9449 , \9454 );
buf \U$9361 ( \9456 , \9455 );
buf \U$9362 ( \9457 , \9456 );
nand \U$9363 ( \9458 , \9448 , \9457 );
buf \U$9364 ( \9459 , \9458 );
xor \U$9365 ( \9460 , \9443 , \9459 );
buf \U$9366 ( \9461 , \9257 );
not \U$9367 ( \9462 , \9461 );
buf \U$9368 ( \9463 , \2124 );
not \U$9369 ( \9464 , \9463 );
or \U$9370 ( \9465 , \9462 , \9464 );
buf \U$9371 ( \9466 , \1565 );
buf \U$9372 ( \9467 , RIc0d7948_7);
buf \U$9373 ( \9468 , RIc0d9928_75);
xor \U$9374 ( \9469 , \9467 , \9468 );
buf \U$9375 ( \9470 , \9469 );
buf \U$9376 ( \9471 , \9470 );
nand \U$9377 ( \9472 , \9466 , \9471 );
buf \U$9378 ( \9473 , \9472 );
buf \U$9379 ( \9474 , \9473 );
nand \U$9380 ( \9475 , \9465 , \9474 );
buf \U$9381 ( \9476 , \9475 );
buf \U$9382 ( \9477 , \9476 );
buf \U$9383 ( \9478 , \996 );
not \U$9384 ( \9479 , \9478 );
buf \U$9385 ( \9480 , \2091 );
not \U$9386 ( \9481 , \9480 );
or \U$9387 ( \9482 , \9479 , \9481 );
buf \U$9388 ( \9483 , RIc0d9ce8_83);
nand \U$9389 ( \9484 , \9482 , \9483 );
buf \U$9390 ( \9485 , \9484 );
buf \U$9391 ( \9486 , \9485 );
xor \U$9392 ( \9487 , \9477 , \9486 );
buf \U$9393 ( \9488 , \779 );
buf \U$9394 ( \9489 , \9273 );
or \U$9395 ( \9490 , \9488 , \9489 );
buf \U$9396 ( \9491 , \1856 );
not \U$9397 ( \9492 , \9491 );
buf \U$9398 ( \9493 , \9492 );
buf \U$9399 ( \9494 , \9493 );
buf \U$9400 ( \9495 , RIc0d7a38_9);
buf \U$9401 ( \9496 , RIc0d9838_73);
xor \U$9402 ( \9497 , \9495 , \9496 );
buf \U$9403 ( \9498 , \9497 );
buf \U$9404 ( \9499 , \9498 );
not \U$9405 ( \9500 , \9499 );
buf \U$9406 ( \9501 , \9500 );
buf \U$9407 ( \9502 , \9501 );
or \U$9408 ( \9503 , \9494 , \9502 );
nand \U$9409 ( \9504 , \9490 , \9503 );
buf \U$9410 ( \9505 , \9504 );
buf \U$9411 ( \9506 , \9505 );
xor \U$9412 ( \9507 , \9487 , \9506 );
buf \U$9413 ( \9508 , \9507 );
buf \U$9414 ( \9509 , \9142 );
not \U$9415 ( \9510 , \9509 );
buf \U$9416 ( \9511 , \1225 );
not \U$9417 ( \9512 , \9511 );
or \U$9418 ( \9513 , \9510 , \9512 );
buf \U$9419 ( \9514 , \1705 );
buf \U$9420 ( \9515 , RIc0d9478_65);
buf \U$9421 ( \9516 , RIc0d7df8_17);
xor \U$9422 ( \9517 , \9515 , \9516 );
buf \U$9423 ( \9518 , \9517 );
buf \U$9424 ( \9519 , \9518 );
nand \U$9425 ( \9520 , \9514 , \9519 );
buf \U$9426 ( \9521 , \9520 );
buf \U$9427 ( \9522 , \9521 );
nand \U$9428 ( \9523 , \9513 , \9522 );
buf \U$9429 ( \9524 , \9523 );
buf \U$9430 ( \9525 , \9067 );
not \U$9431 ( \9526 , \9525 );
buf \U$9432 ( \9527 , \1263 );
not \U$9433 ( \9528 , \9527 );
or \U$9434 ( \9529 , \9526 , \9528 );
buf \U$9435 ( \9530 , RIc0d9748_71);
buf \U$9436 ( \9531 , RIc0d7b28_11);
xnor \U$9437 ( \9532 , \9530 , \9531 );
buf \U$9438 ( \9533 , \9532 );
buf \U$9439 ( \9534 , \9533 );
not \U$9440 ( \9535 , \9534 );
buf \U$9441 ( \9536 , \1282 );
nand \U$9442 ( \9537 , \9535 , \9536 );
buf \U$9443 ( \9538 , \9537 );
buf \U$9444 ( \9539 , \9538 );
nand \U$9445 ( \9540 , \9529 , \9539 );
buf \U$9446 ( \9541 , \9540 );
xor \U$9447 ( \9542 , \9524 , \9541 );
buf \U$9448 ( \9543 , \9542 );
buf \U$9449 ( \9544 , \9169 );
not \U$9450 ( \9545 , \9544 );
buf \U$9451 ( \9546 , \279 );
not \U$9452 ( \9547 , \9546 );
or \U$9453 ( \9548 , \9545 , \9547 );
buf \U$9454 ( \9549 , \874 );
buf \U$9455 ( \9550 , RIc0d7c18_13);
buf \U$9456 ( \9551 , RIc0d9658_69);
xor \U$9457 ( \9552 , \9550 , \9551 );
buf \U$9458 ( \9553 , \9552 );
buf \U$9459 ( \9554 , \9553 );
nand \U$9460 ( \9555 , \9549 , \9554 );
buf \U$9461 ( \9556 , \9555 );
buf \U$9462 ( \9557 , \9556 );
nand \U$9463 ( \9558 , \9548 , \9557 );
buf \U$9464 ( \9559 , \9558 );
buf \U$9465 ( \9560 , \9559 );
xor \U$9466 ( \9561 , \9543 , \9560 );
buf \U$9467 ( \9562 , \9561 );
xor \U$9468 ( \9563 , \9508 , \9562 );
xor \U$9469 ( \9564 , \9460 , \9563 );
buf \U$9470 ( \9565 , \9564 );
xor \U$9471 ( \9566 , \9422 , \9565 );
buf \U$9472 ( \9567 , \9566 );
xor \U$9473 ( \9568 , \9364 , \9567 );
xor \U$9474 ( \9569 , \9122 , \9128 );
and \U$9475 ( \9570 , \9569 , \9309 );
and \U$9476 ( \9571 , \9122 , \9128 );
or \U$9477 ( \9572 , \9570 , \9571 );
buf \U$9478 ( \9573 , \9572 );
xor \U$9479 ( \9574 , \9086 , \9091 );
xor \U$9480 ( \9575 , \9574 , \9096 );
and \U$9481 ( \9576 , \9102 , \9575 );
xor \U$9482 ( \9577 , \9086 , \9091 );
xor \U$9483 ( \9578 , \9577 , \9096 );
and \U$9484 ( \9579 , \9311 , \9578 );
and \U$9485 ( \9580 , \9102 , \9311 );
or \U$9486 ( \9581 , \9576 , \9579 , \9580 );
xor \U$9487 ( \9582 , \9573 , \9581 );
xor \U$9488 ( \9583 , \9568 , \9582 );
buf \U$9489 ( \9584 , \9583 );
nor \U$9490 ( \9585 , \9319 , \9584 );
buf \U$9491 ( \9586 , \9585 );
buf \U$9492 ( \9587 , \9586 );
xor \U$9493 ( \9588 , \9039 , \9048 );
xor \U$9494 ( \9589 , \9588 , \9314 );
buf \U$9495 ( \9590 , \9589 );
buf \U$9496 ( \9591 , \9590 );
xor \U$9497 ( \9592 , \8770 , \8971 );
and \U$9498 ( \9593 , \9592 , \9021 );
and \U$9499 ( \9594 , \8770 , \8971 );
or \U$9500 ( \9595 , \9593 , \9594 );
buf \U$9501 ( \9596 , \9595 );
buf \U$9502 ( \9597 , \9596 );
nor \U$9503 ( \9598 , \9591 , \9597 );
buf \U$9504 ( \9599 , \9598 );
buf \U$9505 ( \9600 , \9599 );
nor \U$9506 ( \9601 , \9587 , \9600 );
buf \U$9507 ( \9602 , \9601 );
buf \U$9508 ( \9603 , \9602 );
xor \U$9509 ( \9604 , \9073 , \9337 );
xor \U$9510 ( \9605 , \9604 , \9350 );
and \U$9511 ( \9606 , \9356 , \9605 );
xor \U$9512 ( \9607 , \9073 , \9337 );
xor \U$9513 ( \9608 , \9607 , \9350 );
and \U$9514 ( \9609 , \9361 , \9608 );
and \U$9515 ( \9610 , \9356 , \9361 );
or \U$9516 ( \9611 , \9606 , \9609 , \9610 );
xor \U$9517 ( \9612 , \9073 , \9337 );
and \U$9518 ( \9613 , \9612 , \9350 );
and \U$9519 ( \9614 , \9073 , \9337 );
or \U$9520 ( \9615 , \9613 , \9614 );
buf \U$9521 ( \9616 , \9615 );
and \U$9522 ( \9617 , \9139 , \9140 );
buf \U$9523 ( \9618 , \9617 );
buf \U$9524 ( \9619 , \9618 );
buf \U$9525 ( \9620 , \9498 );
not \U$9526 ( \9621 , \9620 );
buf \U$9527 ( \9622 , \776 );
not \U$9528 ( \9623 , \9622 );
or \U$9529 ( \9624 , \9621 , \9623 );
buf \U$9530 ( \9625 , RIc0d9838_73);
buf \U$9531 ( \9626 , RIc0d79c0_8);
xnor \U$9532 ( \9627 , \9625 , \9626 );
buf \U$9533 ( \9628 , \9627 );
buf \U$9534 ( \9629 , \9628 );
not \U$9535 ( \9630 , \9629 );
buf \U$9536 ( \9631 , \792 );
nand \U$9537 ( \9632 , \9630 , \9631 );
buf \U$9538 ( \9633 , \9632 );
buf \U$9539 ( \9634 , \9633 );
nand \U$9540 ( \9635 , \9624 , \9634 );
buf \U$9541 ( \9636 , \9635 );
buf \U$9542 ( \9637 , \9636 );
xor \U$9543 ( \9638 , \9619 , \9637 );
buf \U$9544 ( \9639 , \1124 );
buf \U$9545 ( \9640 , \9470 );
not \U$9546 ( \9641 , \9640 );
buf \U$9547 ( \9642 , \9641 );
buf \U$9548 ( \9643 , \9642 );
or \U$9549 ( \9644 , \9639 , \9643 );
buf \U$9550 ( \9645 , \1370 );
buf \U$9551 ( \9646 , RIc0d78d0_6);
buf \U$9552 ( \9647 , RIc0d9928_75);
xnor \U$9553 ( \9648 , \9646 , \9647 );
buf \U$9554 ( \9649 , \9648 );
buf \U$9555 ( \9650 , \9649 );
or \U$9556 ( \9651 , \9645 , \9650 );
nand \U$9557 ( \9652 , \9644 , \9651 );
buf \U$9558 ( \9653 , \9652 );
buf \U$9559 ( \9654 , \9653 );
xor \U$9560 ( \9655 , \9638 , \9654 );
buf \U$9561 ( \9656 , \9655 );
buf \U$9562 ( \9657 , \9656 );
xor \U$9563 ( \9658 , \9616 , \9657 );
xor \U$9564 ( \9659 , \9396 , \9402 );
and \U$9565 ( \9660 , \9659 , \9418 );
and \U$9566 ( \9661 , \9396 , \9402 );
or \U$9567 ( \9662 , \9660 , \9661 );
buf \U$9568 ( \9663 , \9662 );
buf \U$9569 ( \9664 , \9663 );
xor \U$9570 ( \9665 , \9658 , \9664 );
buf \U$9571 ( \9666 , \9665 );
xor \U$9572 ( \9667 , \9611 , \9666 );
xor \U$9573 ( \9668 , \9381 , \9421 );
and \U$9574 ( \9669 , \9668 , \9565 );
and \U$9575 ( \9670 , \9381 , \9421 );
or \U$9576 ( \9671 , \9669 , \9670 );
buf \U$9577 ( \9672 , \9671 );
xor \U$9578 ( \9673 , \9667 , \9672 );
buf \U$9579 ( \9674 , \1263 );
not \U$9580 ( \9675 , \9674 );
buf \U$9581 ( \9676 , \9675 );
buf \U$9582 ( \9677 , \9676 );
buf \U$9583 ( \9678 , \9533 );
or \U$9584 ( \9679 , \9677 , \9678 );
buf \U$9585 ( \9680 , \1279 );
buf \U$9586 ( \9681 , RIc0d7ab0_10);
buf \U$9587 ( \9682 , RIc0d9748_71);
xor \U$9588 ( \9683 , \9681 , \9682 );
buf \U$9589 ( \9684 , \9683 );
buf \U$9590 ( \9685 , \9684 );
not \U$9591 ( \9686 , \9685 );
buf \U$9592 ( \9687 , \9686 );
buf \U$9593 ( \9688 , \9687 );
or \U$9594 ( \9689 , \9680 , \9688 );
nand \U$9595 ( \9690 , \9679 , \9689 );
buf \U$9596 ( \9691 , \9690 );
buf \U$9597 ( \9692 , \9691 );
not \U$9598 ( \9693 , \9692 );
buf \U$9599 ( \9694 , \9693 );
buf \U$9600 ( \9695 , \9694 );
buf \U$9601 ( \9696 , \9524 );
buf \U$9602 ( \9697 , \9541 );
or \U$9603 ( \9698 , \9696 , \9697 );
buf \U$9604 ( \9699 , \9559 );
nand \U$9605 ( \9700 , \9698 , \9699 );
buf \U$9606 ( \9701 , \9700 );
buf \U$9607 ( \9702 , \9701 );
buf \U$9608 ( \9703 , \9524 );
buf \U$9609 ( \9704 , \9541 );
nand \U$9610 ( \9705 , \9703 , \9704 );
buf \U$9611 ( \9706 , \9705 );
buf \U$9612 ( \9707 , \9706 );
nand \U$9613 ( \9708 , \9702 , \9707 );
buf \U$9614 ( \9709 , \9708 );
buf \U$9615 ( \9710 , \9709 );
xor \U$9616 ( \9711 , \9695 , \9710 );
xor \U$9617 ( \9712 , \9477 , \9486 );
and \U$9618 ( \9713 , \9712 , \9506 );
and \U$9619 ( \9714 , \9477 , \9486 );
or \U$9620 ( \9715 , \9713 , \9714 );
buf \U$9621 ( \9716 , \9715 );
buf \U$9622 ( \9717 , \9716 );
xor \U$9623 ( \9718 , \9711 , \9717 );
buf \U$9624 ( \9719 , \9718 );
buf \U$9625 ( \9720 , \9719 );
xor \U$9626 ( \9721 , \9426 , \9442 );
xor \U$9627 ( \9722 , \9721 , \9459 );
and \U$9628 ( \9723 , \9508 , \9722 );
xor \U$9629 ( \9724 , \9426 , \9442 );
xor \U$9630 ( \9725 , \9724 , \9459 );
and \U$9631 ( \9726 , \9562 , \9725 );
and \U$9632 ( \9727 , \9508 , \9562 );
or \U$9633 ( \9728 , \9723 , \9726 , \9727 );
buf \U$9634 ( \9729 , \9728 );
xor \U$9635 ( \9730 , \9720 , \9729 );
xor \U$9636 ( \9731 , \9426 , \9442 );
and \U$9637 ( \9732 , \9731 , \9459 );
and \U$9638 ( \9733 , \9426 , \9442 );
or \U$9639 ( \9734 , \9732 , \9733 );
buf \U$9640 ( \9735 , \9734 );
buf \U$9641 ( \9736 , \9329 );
not \U$9642 ( \9737 , \9736 );
buf \U$9643 ( \9738 , \4509 );
not \U$9644 ( \9739 , \9738 );
or \U$9645 ( \9740 , \9737 , \9739 );
buf \U$9646 ( \9741 , \1026 );
buf \U$9647 ( \9742 , RIc0d76f0_2);
buf \U$9648 ( \9743 , RIc0d9b08_79);
xor \U$9649 ( \9744 , \9742 , \9743 );
buf \U$9650 ( \9745 , \9744 );
buf \U$9651 ( \9746 , \9745 );
nand \U$9652 ( \9747 , \9741 , \9746 );
buf \U$9653 ( \9748 , \9747 );
buf \U$9654 ( \9749 , \9748 );
nand \U$9655 ( \9750 , \9740 , \9749 );
buf \U$9656 ( \9751 , \9750 );
buf \U$9657 ( \9752 , \9751 );
buf \U$9658 ( \9753 , \9453 );
not \U$9659 ( \9754 , \9753 );
buf \U$9660 ( \9755 , \1183 );
not \U$9661 ( \9756 , \9755 );
or \U$9662 ( \9757 , \9754 , \9756 );
xnor \U$9663 ( \9758 , RIc0d9a18_77, RIc0d77e0_4);
buf \U$9664 ( \9759 , \9758 );
not \U$9665 ( \9760 , \9759 );
buf \U$9666 ( \9761 , \1588 );
nand \U$9667 ( \9762 , \9760 , \9761 );
buf \U$9668 ( \9763 , \9762 );
buf \U$9669 ( \9764 , \9763 );
nand \U$9670 ( \9765 , \9757 , \9764 );
buf \U$9671 ( \9766 , \9765 );
buf \U$9672 ( \9767 , \9766 );
xor \U$9673 ( \9768 , \9752 , \9767 );
buf \U$9674 ( \9769 , \3566 );
buf \U$9675 ( \9770 , \9346 );
or \U$9676 ( \9771 , \9769 , \9770 );
buf \U$9677 ( \9772 , \2775 );
buf \U$9678 ( \9773 , \7998 );
or \U$9679 ( \9774 , \9772 , \9773 );
nand \U$9680 ( \9775 , \9771 , \9774 );
buf \U$9681 ( \9776 , \9775 );
buf \U$9682 ( \9777 , \9776 );
xor \U$9683 ( \9778 , \9768 , \9777 );
buf \U$9684 ( \9779 , \9778 );
buf \U$9685 ( \9780 , \9779 );
xor \U$9686 ( \9781 , \9735 , \9780 );
buf \U$9687 ( \9782 , \9553 );
not \U$9688 ( \9783 , \9782 );
buf \U$9689 ( \9784 , \279 );
not \U$9690 ( \9785 , \9784 );
or \U$9691 ( \9786 , \9783 , \9785 );
buf \U$9692 ( \9787 , \874 );
buf \U$9693 ( \9788 , RIc0d7ba0_12);
buf \U$9694 ( \9789 , RIc0d9658_69);
xor \U$9695 ( \9790 , \9788 , \9789 );
buf \U$9696 ( \9791 , \9790 );
buf \U$9697 ( \9792 , \9791 );
nand \U$9698 ( \9793 , \9787 , \9792 );
buf \U$9699 ( \9794 , \9793 );
buf \U$9700 ( \9795 , \9794 );
nand \U$9701 ( \9796 , \9786 , \9795 );
buf \U$9702 ( \9797 , \9796 );
buf \U$9703 ( \9798 , \9518 );
not \U$9704 ( \9799 , \9798 );
buf \U$9705 ( \9800 , \1224 );
not \U$9706 ( \9801 , \9800 );
or \U$9707 ( \9802 , \9799 , \9801 );
buf \U$9708 ( \9803 , \1229 );
buf \U$9709 ( \9804 , RIc0d9478_65);
buf \U$9710 ( \9805 , RIc0d7d80_16);
xor \U$9711 ( \9806 , \9804 , \9805 );
buf \U$9712 ( \9807 , \9806 );
buf \U$9713 ( \9808 , \9807 );
nand \U$9714 ( \9809 , \9803 , \9808 );
buf \U$9715 ( \9810 , \9809 );
buf \U$9716 ( \9811 , \9810 );
nand \U$9717 ( \9812 , \9802 , \9811 );
buf \U$9718 ( \9813 , \9812 );
xor \U$9719 ( \9814 , \9797 , \9813 );
buf \U$9720 ( \9815 , \9436 );
not \U$9721 ( \9816 , \9815 );
buf \U$9722 ( \9817 , \2900 );
not \U$9723 ( \9818 , \9817 );
or \U$9724 ( \9819 , \9816 , \9818 );
buf \U$9725 ( \9820 , \686 );
buf \U$9726 ( \9821 , RIc0d7c90_14);
buf \U$9727 ( \9822 , RIc0d9568_67);
xor \U$9728 ( \9823 , \9821 , \9822 );
buf \U$9729 ( \9824 , \9823 );
buf \U$9730 ( \9825 , \9824 );
nand \U$9731 ( \9826 , \9820 , \9825 );
buf \U$9732 ( \9827 , \9826 );
buf \U$9733 ( \9828 , \9827 );
nand \U$9734 ( \9829 , \9819 , \9828 );
buf \U$9735 ( \9830 , \9829 );
xor \U$9736 ( \9831 , \9814 , \9830 );
buf \U$9737 ( \9832 , \9831 );
xor \U$9738 ( \9833 , \9781 , \9832 );
buf \U$9739 ( \9834 , \9833 );
buf \U$9740 ( \9835 , \9834 );
xor \U$9741 ( \9836 , \9730 , \9835 );
buf \U$9742 ( \9837 , \9836 );
xor \U$9743 ( \9838 , \9323 , \9363 );
and \U$9744 ( \9839 , \9838 , \9567 );
and \U$9745 ( \9840 , \9323 , \9363 );
or \U$9746 ( \9841 , \9839 , \9840 );
xor \U$9747 ( \9842 , \9837 , \9841 );
xor \U$9748 ( \9843 , \9673 , \9842 );
buf \U$9749 ( \9844 , \9843 );
xor \U$9750 ( \9845 , \9323 , \9363 );
xor \U$9751 ( \9846 , \9845 , \9567 );
and \U$9752 ( \9847 , \9573 , \9846 );
xor \U$9753 ( \9848 , \9323 , \9363 );
xor \U$9754 ( \9849 , \9848 , \9567 );
and \U$9755 ( \9850 , \9581 , \9849 );
and \U$9756 ( \9851 , \9573 , \9581 );
or \U$9757 ( \9852 , \9847 , \9850 , \9851 );
buf \U$9758 ( \9853 , \9852 );
or \U$9759 ( \9854 , \9844 , \9853 );
buf \U$9760 ( \9855 , \9854 );
buf \U$9761 ( \9856 , \9855 );
and \U$9762 ( \9857 , \9603 , \9856 );
buf \U$9763 ( \9858 , \9857 );
buf \U$9764 ( \9859 , \9858 );
xor \U$9765 ( \9860 , \9611 , \9666 );
xor \U$9766 ( \9861 , \9860 , \9672 );
and \U$9767 ( \9862 , \9837 , \9861 );
xor \U$9768 ( \9863 , \9611 , \9666 );
xor \U$9769 ( \9864 , \9863 , \9672 );
and \U$9770 ( \9865 , \9841 , \9864 );
and \U$9771 ( \9866 , \9837 , \9841 );
or \U$9772 ( \9867 , \9862 , \9865 , \9866 );
buf \U$9773 ( \9868 , \9867 );
xor \U$9774 ( \9869 , \9695 , \9710 );
and \U$9775 ( \9870 , \9869 , \9717 );
and \U$9776 ( \9871 , \9695 , \9710 );
or \U$9777 ( \9872 , \9870 , \9871 );
buf \U$9778 ( \9873 , \9872 );
buf \U$9779 ( \9874 , \9873 );
xor \U$9780 ( \9875 , \9735 , \9780 );
and \U$9781 ( \9876 , \9875 , \9832 );
and \U$9782 ( \9877 , \9735 , \9780 );
or \U$9783 ( \9878 , \9876 , \9877 );
buf \U$9784 ( \9879 , \9878 );
buf \U$9785 ( \9880 , \9879 );
xor \U$9786 ( \9881 , \9874 , \9880 );
buf \U$9787 ( \9882 , \9649 );
not \U$9788 ( \9883 , \9882 );
buf \U$9789 ( \9884 , \9883 );
buf \U$9790 ( \9885 , \9884 );
not \U$9791 ( \9886 , \9885 );
buf \U$9792 ( \9887 , \2359 );
not \U$9793 ( \9888 , \9887 );
or \U$9794 ( \9889 , \9886 , \9888 );
buf \U$9795 ( \9890 , \1143 );
buf \U$9796 ( \9891 , RIc0d7858_5);
buf \U$9797 ( \9892 , RIc0d9928_75);
xor \U$9798 ( \9893 , \9891 , \9892 );
buf \U$9799 ( \9894 , \9893 );
buf \U$9800 ( \9895 , \9894 );
nand \U$9801 ( \9896 , \9890 , \9895 );
buf \U$9802 ( \9897 , \9896 );
buf \U$9803 ( \9898 , \9897 );
nand \U$9804 ( \9899 , \9889 , \9898 );
buf \U$9805 ( \9900 , \9899 );
buf \U$9806 ( \9901 , \9900 );
buf \U$9807 ( \9902 , \9745 );
not \U$9808 ( \9903 , \9902 );
buf \U$9809 ( \9904 , \1351 );
not \U$9810 ( \9905 , \9904 );
or \U$9811 ( \9906 , \9903 , \9905 );
buf \U$9812 ( \9907 , \403 );
buf \U$9813 ( \9908 , RIc0d7678_1);
buf \U$9814 ( \9909 , RIc0d9b08_79);
xor \U$9815 ( \9910 , \9908 , \9909 );
buf \U$9816 ( \9911 , \9910 );
buf \U$9817 ( \9912 , \9911 );
nand \U$9818 ( \9913 , \9907 , \9912 );
buf \U$9819 ( \9914 , \9913 );
buf \U$9820 ( \9915 , \9914 );
nand \U$9821 ( \9916 , \9906 , \9915 );
buf \U$9822 ( \9917 , \9916 );
buf \U$9823 ( \9918 , \9917 );
xor \U$9824 ( \9919 , \9901 , \9918 );
buf \U$9825 ( \9920 , \2871 );
not \U$9826 ( \9921 , \9920 );
buf \U$9827 ( \9922 , \9921 );
buf \U$9828 ( \9923 , \9922 );
buf \U$9829 ( \9924 , \9628 );
or \U$9830 ( \9925 , \9923 , \9924 );
buf \U$9831 ( \9926 , \2879 );
buf \U$9832 ( \9927 , RIc0d7948_7);
buf \U$9833 ( \9928 , RIc0d9838_73);
xnor \U$9834 ( \9929 , \9927 , \9928 );
buf \U$9835 ( \9930 , \9929 );
buf \U$9836 ( \9931 , \9930 );
or \U$9837 ( \9932 , \9926 , \9931 );
nand \U$9838 ( \9933 , \9925 , \9932 );
buf \U$9839 ( \9934 , \9933 );
buf \U$9840 ( \9935 , \9934 );
xor \U$9841 ( \9936 , \9919 , \9935 );
buf \U$9842 ( \9937 , \9936 );
xor \U$9843 ( \9938 , \9752 , \9767 );
and \U$9844 ( \9939 , \9938 , \9777 );
and \U$9845 ( \9940 , \9752 , \9767 );
or \U$9846 ( \9941 , \9939 , \9940 );
buf \U$9847 ( \9942 , \9941 );
xor \U$9848 ( \9943 , \9937 , \9942 );
buf \U$9849 ( \9944 , \9830 );
not \U$9850 ( \9945 , \9944 );
buf \U$9851 ( \9946 , \9813 );
not \U$9852 ( \9947 , \9946 );
or \U$9853 ( \9948 , \9945 , \9947 );
buf \U$9854 ( \9949 , \9813 );
buf \U$9855 ( \9950 , \9830 );
or \U$9856 ( \9951 , \9949 , \9950 );
buf \U$9857 ( \9952 , \9797 );
nand \U$9858 ( \9953 , \9951 , \9952 );
buf \U$9859 ( \9954 , \9953 );
buf \U$9860 ( \9955 , \9954 );
nand \U$9861 ( \9956 , \9948 , \9955 );
buf \U$9862 ( \9957 , \9956 );
xor \U$9863 ( \9958 , \9943 , \9957 );
buf \U$9864 ( \9959 , \9958 );
xor \U$9865 ( \9960 , \9881 , \9959 );
buf \U$9866 ( \9961 , \9960 );
buf \U$9867 ( \9962 , \9961 );
xor \U$9868 ( \9963 , \9611 , \9666 );
and \U$9869 ( \9964 , \9963 , \9672 );
and \U$9870 ( \9965 , \9611 , \9666 );
or \U$9871 ( \9966 , \9964 , \9965 );
buf \U$9872 ( \9967 , \9966 );
xor \U$9873 ( \9968 , \9962 , \9967 );
xor \U$9874 ( \9969 , \9616 , \9657 );
and \U$9875 ( \9970 , \9969 , \9664 );
and \U$9876 ( \9971 , \9616 , \9657 );
or \U$9877 ( \9972 , \9970 , \9971 );
buf \U$9878 ( \9973 , \9972 );
buf \U$9879 ( \9974 , \9973 );
buf \U$9880 ( \9975 , \9807 );
not \U$9881 ( \9976 , \9975 );
buf \U$9882 ( \9977 , \3781 );
not \U$9883 ( \9978 , \9977 );
or \U$9884 ( \9979 , \9976 , \9978 );
buf \U$9885 ( \9980 , \1229 );
buf \U$9886 ( \9981 , RIc0d9478_65);
buf \U$9887 ( \9982 , RIc0d7d08_15);
xor \U$9888 ( \9983 , \9981 , \9982 );
buf \U$9889 ( \9984 , \9983 );
buf \U$9890 ( \9985 , \9984 );
nand \U$9891 ( \9986 , \9980 , \9985 );
buf \U$9892 ( \9987 , \9986 );
buf \U$9893 ( \9988 , \9987 );
nand \U$9894 ( \9989 , \9979 , \9988 );
buf \U$9895 ( \9990 , \9989 );
buf \U$9896 ( \9991 , \9684 );
not \U$9897 ( \9992 , \9991 );
buf \U$9898 ( \9993 , \1263 );
not \U$9899 ( \9994 , \9993 );
or \U$9900 ( \9995 , \9992 , \9994 );
buf \U$9901 ( \9996 , \2927 );
buf \U$9902 ( \9997 , RIc0d7a38_9);
buf \U$9903 ( \9998 , RIc0d9748_71);
xor \U$9904 ( \9999 , \9997 , \9998 );
buf \U$9905 ( \10000 , \9999 );
buf \U$9906 ( \10001 , \10000 );
nand \U$9907 ( \10002 , \9996 , \10001 );
buf \U$9908 ( \10003 , \10002 );
buf \U$9909 ( \10004 , \10003 );
nand \U$9910 ( \10005 , \9995 , \10004 );
buf \U$9911 ( \10006 , \10005 );
xor \U$9912 ( \10007 , \9990 , \10006 );
buf \U$9913 ( \10008 , \9791 );
not \U$9914 ( \10009 , \10008 );
buf \U$9915 ( \10010 , \4692 );
not \U$9916 ( \10011 , \10010 );
or \U$9917 ( \10012 , \10009 , \10011 );
buf \U$9918 ( \10013 , RIc0d7b28_11);
buf \U$9919 ( \10014 , RIc0d9658_69);
xnor \U$9920 ( \10015 , \10013 , \10014 );
buf \U$9921 ( \10016 , \10015 );
buf \U$9922 ( \10017 , \10016 );
not \U$9923 ( \10018 , \10017 );
buf \U$9924 ( \10019 , \284 );
nand \U$9925 ( \10020 , \10018 , \10019 );
buf \U$9926 ( \10021 , \10020 );
buf \U$9927 ( \10022 , \10021 );
nand \U$9928 ( \10023 , \10012 , \10022 );
buf \U$9929 ( \10024 , \10023 );
xor \U$9930 ( \10025 , \10007 , \10024 );
buf \U$9931 ( \10026 , \10025 );
and \U$9932 ( \10027 , \9515 , \9516 );
buf \U$9933 ( \10028 , \10027 );
buf \U$9934 ( \10029 , \10028 );
buf \U$9935 ( \10030 , \9824 );
not \U$9936 ( \10031 , \10030 );
buf \U$9937 ( \10032 , \1417 );
not \U$9938 ( \10033 , \10032 );
buf \U$9939 ( \10034 , \10033 );
buf \U$9940 ( \10035 , \10034 );
not \U$9941 ( \10036 , \10035 );
or \U$9942 ( \10037 , \10031 , \10036 );
buf \U$9943 ( \10038 , \686 );
buf \U$9944 ( \10039 , RIc0d7c18_13);
buf \U$9945 ( \10040 , RIc0d9568_67);
xor \U$9946 ( \10041 , \10039 , \10040 );
buf \U$9947 ( \10042 , \10041 );
buf \U$9948 ( \10043 , \10042 );
nand \U$9949 ( \10044 , \10038 , \10043 );
buf \U$9950 ( \10045 , \10044 );
buf \U$9951 ( \10046 , \10045 );
nand \U$9952 ( \10047 , \10037 , \10046 );
buf \U$9953 ( \10048 , \10047 );
buf \U$9954 ( \10049 , \10048 );
xor \U$9955 ( \10050 , \10029 , \10049 );
buf \U$9956 ( \10051 , \1435 );
buf \U$9957 ( \10052 , \9758 );
or \U$9958 ( \10053 , \10051 , \10052 );
buf \U$9959 ( \10054 , \1193 );
buf \U$9960 ( \10055 , RIc0d7768_3);
buf \U$9961 ( \10056 , RIc0d9a18_77);
xnor \U$9962 ( \10057 , \10055 , \10056 );
buf \U$9963 ( \10058 , \10057 );
buf \U$9964 ( \10059 , \10058 );
or \U$9965 ( \10060 , \10054 , \10059 );
nand \U$9966 ( \10061 , \10053 , \10060 );
buf \U$9967 ( \10062 , \10061 );
buf \U$9968 ( \10063 , \10062 );
xor \U$9969 ( \10064 , \10050 , \10063 );
buf \U$9970 ( \10065 , \10064 );
buf \U$9971 ( \10066 , \10065 );
xor \U$9972 ( \10067 , \10026 , \10066 );
buf \U$9973 ( \10068 , \1610 );
not \U$9974 ( \10069 , \10068 );
buf \U$9975 ( \10070 , \3566 );
not \U$9976 ( \10071 , \10070 );
or \U$9977 ( \10072 , \10069 , \10071 );
buf \U$9978 ( \10073 , RIc0d9bf8_81);
nand \U$9979 ( \10074 , \10072 , \10073 );
buf \U$9980 ( \10075 , \10074 );
buf \U$9981 ( \10076 , \10075 );
buf \U$9982 ( \10077 , \9691 );
xor \U$9983 ( \10078 , \10076 , \10077 );
xor \U$9984 ( \10079 , \9619 , \9637 );
and \U$9985 ( \10080 , \10079 , \9654 );
and \U$9986 ( \10081 , \9619 , \9637 );
or \U$9987 ( \10082 , \10080 , \10081 );
buf \U$9988 ( \10083 , \10082 );
buf \U$9989 ( \10084 , \10083 );
xor \U$9990 ( \10085 , \10078 , \10084 );
buf \U$9991 ( \10086 , \10085 );
buf \U$9992 ( \10087 , \10086 );
xor \U$9993 ( \10088 , \10067 , \10087 );
buf \U$9994 ( \10089 , \10088 );
buf \U$9995 ( \10090 , \10089 );
xor \U$9996 ( \10091 , \9974 , \10090 );
xor \U$9997 ( \10092 , \9720 , \9729 );
and \U$9998 ( \10093 , \10092 , \9835 );
and \U$9999 ( \10094 , \9720 , \9729 );
or \U$10000 ( \10095 , \10093 , \10094 );
buf \U$10001 ( \10096 , \10095 );
buf \U$10002 ( \10097 , \10096 );
xor \U$10003 ( \10098 , \10091 , \10097 );
buf \U$10004 ( \10099 , \10098 );
buf \U$10005 ( \10100 , \10099 );
xor \U$10006 ( \10101 , \9968 , \10100 );
buf \U$10007 ( \10102 , \10101 );
buf \U$10008 ( \10103 , \10102 );
or \U$10009 ( \10104 , \9868 , \10103 );
buf \U$10010 ( \10105 , \10104 );
buf \U$10011 ( \10106 , \10105 );
and \U$10012 ( \10107 , \9859 , \10106 );
buf \U$10013 ( \10108 , \10107 );
buf \U$10014 ( \10109 , \10108 );
and \U$10015 ( \10110 , \9033 , \10109 );
buf \U$10016 ( \10111 , \10110 );
buf \U$10017 ( \10112 , \10111 );
xor \U$10018 ( \10113 , \10076 , \10077 );
and \U$10019 ( \10114 , \10113 , \10084 );
and \U$10020 ( \10115 , \10076 , \10077 );
or \U$10021 ( \10116 , \10114 , \10115 );
buf \U$10022 ( \10117 , \10116 );
buf \U$10023 ( \10118 , \10117 );
buf \U$10024 ( \10119 , \9942 );
buf \U$10025 ( \10120 , \9957 );
or \U$10026 ( \10121 , \10119 , \10120 );
buf \U$10027 ( \10122 , \9937 );
nand \U$10028 ( \10123 , \10121 , \10122 );
buf \U$10029 ( \10124 , \10123 );
buf \U$10030 ( \10125 , \10124 );
buf \U$10031 ( \10126 , \9942 );
buf \U$10032 ( \10127 , \9957 );
nand \U$10033 ( \10128 , \10126 , \10127 );
buf \U$10034 ( \10129 , \10128 );
buf \U$10035 ( \10130 , \10129 );
nand \U$10036 ( \10131 , \10125 , \10130 );
buf \U$10037 ( \10132 , \10131 );
buf \U$10038 ( \10133 , \10132 );
xor \U$10039 ( \10134 , \10118 , \10133 );
buf \U$10040 ( \10135 , \9990 );
buf \U$10041 ( \10136 , \10006 );
or \U$10042 ( \10137 , \10135 , \10136 );
buf \U$10043 ( \10138 , \10024 );
nand \U$10044 ( \10139 , \10137 , \10138 );
buf \U$10045 ( \10140 , \10139 );
buf \U$10046 ( \10141 , \10140 );
buf \U$10047 ( \10142 , \9990 );
buf \U$10048 ( \10143 , \10006 );
nand \U$10049 ( \10144 , \10142 , \10143 );
buf \U$10050 ( \10145 , \10144 );
buf \U$10051 ( \10146 , \10145 );
nand \U$10052 ( \10147 , \10141 , \10146 );
buf \U$10053 ( \10148 , \10147 );
buf \U$10054 ( \10149 , \10148 );
xor \U$10055 ( \10150 , \10029 , \10049 );
and \U$10056 ( \10151 , \10150 , \10063 );
and \U$10057 ( \10152 , \10029 , \10049 );
or \U$10058 ( \10153 , \10151 , \10152 );
buf \U$10059 ( \10154 , \10153 );
buf \U$10060 ( \10155 , \10154 );
xor \U$10061 ( \10156 , \10149 , \10155 );
xor \U$10062 ( \10157 , \9901 , \9918 );
and \U$10063 ( \10158 , \10157 , \9935 );
and \U$10064 ( \10159 , \9901 , \9918 );
or \U$10065 ( \10160 , \10158 , \10159 );
buf \U$10066 ( \10161 , \10160 );
buf \U$10067 ( \10162 , \10161 );
xor \U$10068 ( \10163 , \10156 , \10162 );
buf \U$10069 ( \10164 , \10163 );
buf \U$10070 ( \10165 , \10164 );
xor \U$10071 ( \10166 , \10134 , \10165 );
buf \U$10072 ( \10167 , \10166 );
buf \U$10073 ( \10168 , \10167 );
xor \U$10074 ( \10169 , \10026 , \10066 );
and \U$10075 ( \10170 , \10169 , \10087 );
and \U$10076 ( \10171 , \10026 , \10066 );
or \U$10077 ( \10172 , \10170 , \10171 );
buf \U$10078 ( \10173 , \10172 );
buf \U$10079 ( \10174 , \10173 );
and \U$10080 ( \10175 , \9804 , \9805 );
buf \U$10081 ( \10176 , \10175 );
buf \U$10082 ( \10177 , \10176 );
buf \U$10083 ( \10178 , \10000 );
not \U$10084 ( \10179 , \10178 );
buf \U$10085 ( \10180 , \1263 );
not \U$10086 ( \10181 , \10180 );
or \U$10087 ( \10182 , \10179 , \10181 );
buf \U$10088 ( \10183 , \2927 );
buf \U$10089 ( \10184 , RIc0d79c0_8);
buf \U$10090 ( \10185 , RIc0d9748_71);
xor \U$10091 ( \10186 , \10184 , \10185 );
buf \U$10092 ( \10187 , \10186 );
buf \U$10093 ( \10188 , \10187 );
nand \U$10094 ( \10189 , \10183 , \10188 );
buf \U$10095 ( \10190 , \10189 );
buf \U$10096 ( \10191 , \10190 );
nand \U$10097 ( \10192 , \10182 , \10191 );
buf \U$10098 ( \10193 , \10192 );
buf \U$10099 ( \10194 , \10193 );
not \U$10100 ( \10195 , \10194 );
buf \U$10101 ( \10196 , \10195 );
buf \U$10102 ( \10197 , \10196 );
xor \U$10103 ( \10198 , \10177 , \10197 );
buf \U$10104 ( \10199 , \9930 );
not \U$10105 ( \10200 , \10199 );
buf \U$10106 ( \10201 , \10200 );
buf \U$10107 ( \10202 , \10201 );
not \U$10108 ( \10203 , \10202 );
buf \U$10109 ( \10204 , \1677 );
not \U$10110 ( \10205 , \10204 );
or \U$10111 ( \10206 , \10203 , \10205 );
buf \U$10112 ( \10207 , \2882 );
buf \U$10113 ( \10208 , RIc0d78d0_6);
buf \U$10114 ( \10209 , RIc0d9838_73);
xor \U$10115 ( \10210 , \10208 , \10209 );
buf \U$10116 ( \10211 , \10210 );
buf \U$10117 ( \10212 , \10211 );
nand \U$10118 ( \10213 , \10207 , \10212 );
buf \U$10119 ( \10214 , \10213 );
buf \U$10120 ( \10215 , \10214 );
nand \U$10121 ( \10216 , \10206 , \10215 );
buf \U$10122 ( \10217 , \10216 );
buf \U$10123 ( \10218 , \10217 );
xor \U$10124 ( \10219 , \10198 , \10218 );
buf \U$10125 ( \10220 , \10219 );
buf \U$10126 ( \10221 , \10220 );
buf \U$10127 ( \10222 , \10042 );
not \U$10128 ( \10223 , \10222 );
buf \U$10129 ( \10224 , \4907 );
not \U$10130 ( \10225 , \10224 );
or \U$10131 ( \10226 , \10223 , \10225 );
buf \U$10132 ( \10227 , \686 );
buf \U$10133 ( \10228 , RIc0d7ba0_12);
buf \U$10134 ( \10229 , RIc0d9568_67);
xor \U$10135 ( \10230 , \10228 , \10229 );
buf \U$10136 ( \10231 , \10230 );
buf \U$10137 ( \10232 , \10231 );
nand \U$10138 ( \10233 , \10227 , \10232 );
buf \U$10139 ( \10234 , \10233 );
buf \U$10140 ( \10235 , \10234 );
nand \U$10141 ( \10236 , \10226 , \10235 );
buf \U$10142 ( \10237 , \10236 );
buf \U$10143 ( \10238 , \10237 );
buf \U$10144 ( \10239 , \9894 );
not \U$10145 ( \10240 , \10239 );
buf \U$10146 ( \10241 , \1129 );
not \U$10147 ( \10242 , \10241 );
or \U$10148 ( \10243 , \10240 , \10242 );
buf \U$10149 ( \10244 , RIc0d9928_75);
buf \U$10150 ( \10245 , RIc0d77e0_4);
xnor \U$10151 ( \10246 , \10244 , \10245 );
buf \U$10152 ( \10247 , \10246 );
buf \U$10153 ( \10248 , \10247 );
not \U$10154 ( \10249 , \10248 );
buf \U$10155 ( \10250 , \1143 );
nand \U$10156 ( \10251 , \10249 , \10250 );
buf \U$10157 ( \10252 , \10251 );
buf \U$10158 ( \10253 , \10252 );
nand \U$10159 ( \10254 , \10243 , \10253 );
buf \U$10160 ( \10255 , \10254 );
buf \U$10161 ( \10256 , \10255 );
xor \U$10162 ( \10257 , \10238 , \10256 );
buf \U$10163 ( \10258 , \7753 );
buf \U$10164 ( \10259 , \10058 );
or \U$10165 ( \10260 , \10258 , \10259 );
buf \U$10166 ( \10261 , \1193 );
buf \U$10167 ( \10262 , RIc0d76f0_2);
buf \U$10168 ( \10263 , RIc0d9a18_77);
xnor \U$10169 ( \10264 , \10262 , \10263 );
buf \U$10170 ( \10265 , \10264 );
buf \U$10171 ( \10266 , \10265 );
or \U$10172 ( \10267 , \10261 , \10266 );
nand \U$10173 ( \10268 , \10260 , \10267 );
buf \U$10174 ( \10269 , \10268 );
buf \U$10175 ( \10270 , \10269 );
xor \U$10176 ( \10271 , \10257 , \10270 );
buf \U$10177 ( \10272 , \10271 );
buf \U$10178 ( \10273 , \10272 );
xor \U$10179 ( \10274 , \10221 , \10273 );
buf \U$10180 ( \10275 , \9911 );
not \U$10181 ( \10276 , \10275 );
buf \U$10182 ( \10277 , \1021 );
not \U$10183 ( \10278 , \10277 );
or \U$10184 ( \10279 , \10276 , \10278 );
buf \U$10185 ( \10280 , \403 );
buf \U$10186 ( \10281 , RIc0d9b08_79);
nand \U$10187 ( \10282 , \10280 , \10281 );
buf \U$10188 ( \10283 , \10282 );
buf \U$10189 ( \10284 , \10283 );
nand \U$10190 ( \10285 , \10279 , \10284 );
buf \U$10191 ( \10286 , \10285 );
buf \U$10192 ( \10287 , \9984 );
not \U$10193 ( \10288 , \10287 );
buf \U$10194 ( \10289 , \1225 );
not \U$10195 ( \10290 , \10289 );
or \U$10196 ( \10291 , \10288 , \10290 );
buf \U$10197 ( \10292 , RIc0d7c90_14);
buf \U$10198 ( \10293 , RIc0d9478_65);
xnor \U$10199 ( \10294 , \10292 , \10293 );
buf \U$10200 ( \10295 , \10294 );
buf \U$10201 ( \10296 , \10295 );
not \U$10202 ( \10297 , \10296 );
buf \U$10203 ( \10298 , \1229 );
nand \U$10204 ( \10299 , \10297 , \10298 );
buf \U$10205 ( \10300 , \10299 );
buf \U$10206 ( \10301 , \10300 );
nand \U$10207 ( \10302 , \10291 , \10301 );
buf \U$10208 ( \10303 , \10302 );
xor \U$10209 ( \10304 , \10286 , \10303 );
buf \U$10210 ( \10305 , \1452 );
buf \U$10211 ( \10306 , \10016 );
or \U$10212 ( \10307 , \10305 , \10306 );
buf \U$10213 ( \10308 , \4297 );
buf \U$10214 ( \10309 , RIc0d7ab0_10);
buf \U$10215 ( \10310 , RIc0d9658_69);
xnor \U$10216 ( \10311 , \10309 , \10310 );
buf \U$10217 ( \10312 , \10311 );
buf \U$10218 ( \10313 , \10312 );
or \U$10219 ( \10314 , \10308 , \10313 );
nand \U$10220 ( \10315 , \10307 , \10314 );
buf \U$10221 ( \10316 , \10315 );
xor \U$10222 ( \10317 , \10304 , \10316 );
buf \U$10223 ( \10318 , \10317 );
xor \U$10224 ( \10319 , \10274 , \10318 );
buf \U$10225 ( \10320 , \10319 );
buf \U$10226 ( \10321 , \10320 );
xor \U$10227 ( \10322 , \10174 , \10321 );
xor \U$10228 ( \10323 , \9874 , \9880 );
and \U$10229 ( \10324 , \10323 , \9959 );
and \U$10230 ( \10325 , \9874 , \9880 );
or \U$10231 ( \10326 , \10324 , \10325 );
buf \U$10232 ( \10327 , \10326 );
buf \U$10233 ( \10328 , \10327 );
xor \U$10234 ( \10329 , \10322 , \10328 );
buf \U$10235 ( \10330 , \10329 );
buf \U$10236 ( \10331 , \10330 );
xor \U$10237 ( \10332 , \10168 , \10331 );
xor \U$10238 ( \10333 , \9974 , \10090 );
and \U$10239 ( \10334 , \10333 , \10097 );
and \U$10240 ( \10335 , \9974 , \10090 );
or \U$10241 ( \10336 , \10334 , \10335 );
buf \U$10242 ( \10337 , \10336 );
buf \U$10243 ( \10338 , \10337 );
xor \U$10244 ( \10339 , \10332 , \10338 );
buf \U$10245 ( \10340 , \10339 );
buf \U$10246 ( \10341 , \10340 );
xor \U$10247 ( \10342 , \9962 , \9967 );
and \U$10248 ( \10343 , \10342 , \10100 );
and \U$10249 ( \10344 , \9962 , \9967 );
or \U$10250 ( \10345 , \10343 , \10344 );
buf \U$10251 ( \10346 , \10345 );
buf \U$10252 ( \10347 , \10346 );
nor \U$10253 ( \10348 , \10341 , \10347 );
buf \U$10254 ( \10349 , \10348 );
buf \U$10255 ( \10350 , \10349 );
xor \U$10256 ( \10351 , \10177 , \10197 );
and \U$10257 ( \10352 , \10351 , \10218 );
and \U$10258 ( \10353 , \10177 , \10197 );
or \U$10259 ( \10354 , \10352 , \10353 );
buf \U$10260 ( \10355 , \10354 );
buf \U$10261 ( \10356 , \10355 );
xor \U$10262 ( \10357 , \10149 , \10155 );
and \U$10263 ( \10358 , \10357 , \10162 );
and \U$10264 ( \10359 , \10149 , \10155 );
or \U$10265 ( \10360 , \10358 , \10359 );
buf \U$10266 ( \10361 , \10360 );
buf \U$10267 ( \10362 , \10361 );
xor \U$10268 ( \10363 , \10356 , \10362 );
buf \U$10269 ( \10364 , \10193 );
buf \U$10270 ( \10365 , \10303 );
not \U$10271 ( \10366 , \10365 );
buf \U$10272 ( \10367 , \10286 );
not \U$10273 ( \10368 , \10367 );
or \U$10274 ( \10369 , \10366 , \10368 );
buf \U$10275 ( \10370 , \10286 );
buf \U$10276 ( \10371 , \10303 );
or \U$10277 ( \10372 , \10370 , \10371 );
buf \U$10278 ( \10373 , \10316 );
nand \U$10279 ( \10374 , \10372 , \10373 );
buf \U$10280 ( \10375 , \10374 );
buf \U$10281 ( \10376 , \10375 );
nand \U$10282 ( \10377 , \10369 , \10376 );
buf \U$10283 ( \10378 , \10377 );
buf \U$10284 ( \10379 , \10378 );
xor \U$10285 ( \10380 , \10364 , \10379 );
xor \U$10286 ( \10381 , \10238 , \10256 );
and \U$10287 ( \10382 , \10381 , \10270 );
and \U$10288 ( \10383 , \10238 , \10256 );
or \U$10289 ( \10384 , \10382 , \10383 );
buf \U$10290 ( \10385 , \10384 );
buf \U$10291 ( \10386 , \10385 );
xor \U$10292 ( \10387 , \10380 , \10386 );
buf \U$10293 ( \10388 , \10387 );
buf \U$10294 ( \10389 , \10388 );
xor \U$10295 ( \10390 , \10363 , \10389 );
buf \U$10296 ( \10391 , \10390 );
buf \U$10297 ( \10392 , \10391 );
and \U$10298 ( \10393 , \9981 , \9982 );
buf \U$10299 ( \10394 , \10393 );
buf \U$10300 ( \10395 , \10394 );
buf \U$10301 ( \10396 , \10231 );
not \U$10302 ( \10397 , \10396 );
buf \U$10303 ( \10398 , \2900 );
not \U$10304 ( \10399 , \10398 );
or \U$10305 ( \10400 , \10397 , \10399 );
buf \U$10306 ( \10401 , \686 );
buf \U$10307 ( \10402 , RIc0d7b28_11);
buf \U$10308 ( \10403 , RIc0d9568_67);
xor \U$10309 ( \10404 , \10402 , \10403 );
buf \U$10310 ( \10405 , \10404 );
buf \U$10311 ( \10406 , \10405 );
nand \U$10312 ( \10407 , \10401 , \10406 );
buf \U$10313 ( \10408 , \10407 );
buf \U$10314 ( \10409 , \10408 );
nand \U$10315 ( \10410 , \10400 , \10409 );
buf \U$10316 ( \10411 , \10410 );
buf \U$10317 ( \10412 , \10411 );
xor \U$10318 ( \10413 , \10395 , \10412 );
buf \U$10319 ( \10414 , \6141 );
not \U$10320 ( \10415 , \10414 );
buf \U$10321 ( \10416 , RIc0d7678_1);
buf \U$10322 ( \10417 , RIc0d9a18_77);
xor \U$10323 ( \10418 , \10416 , \10417 );
buf \U$10324 ( \10419 , \10418 );
buf \U$10325 ( \10420 , \10419 );
not \U$10326 ( \10421 , \10420 );
or \U$10327 ( \10422 , \10415 , \10421 );
buf \U$10328 ( \10423 , \1435 );
buf \U$10329 ( \10424 , \10265 );
or \U$10330 ( \10425 , \10423 , \10424 );
nand \U$10331 ( \10426 , \10422 , \10425 );
buf \U$10332 ( \10427 , \10426 );
buf \U$10333 ( \10428 , \10427 );
xor \U$10334 ( \10429 , \10413 , \10428 );
buf \U$10335 ( \10430 , \10429 );
buf \U$10336 ( \10431 , \10430 );
buf \U$10337 ( \10432 , \8178 );
not \U$10338 ( \10433 , \10432 );
buf \U$10339 ( \10434 , \393 );
not \U$10340 ( \10435 , \10434 );
or \U$10341 ( \10436 , \10433 , \10435 );
buf \U$10342 ( \10437 , RIc0d9b08_79);
nand \U$10343 ( \10438 , \10436 , \10437 );
buf \U$10344 ( \10439 , \10438 );
buf \U$10345 ( \10440 , \10439 );
buf \U$10346 ( \10441 , \1556 );
not \U$10347 ( \10442 , \10441 );
buf \U$10348 ( \10443 , \10442 );
buf \U$10349 ( \10444 , \10443 );
buf \U$10350 ( \10445 , \10247 );
or \U$10351 ( \10446 , \10444 , \10445 );
buf \U$10352 ( \10447 , \2372 );
buf \U$10353 ( \10448 , RIc0d7768_3);
buf \U$10354 ( \10449 , RIc0d9928_75);
xor \U$10355 ( \10450 , \10448 , \10449 );
buf \U$10356 ( \10451 , \10450 );
buf \U$10357 ( \10452 , \10451 );
not \U$10358 ( \10453 , \10452 );
buf \U$10359 ( \10454 , \10453 );
buf \U$10360 ( \10455 , \10454 );
or \U$10361 ( \10456 , \10447 , \10455 );
nand \U$10362 ( \10457 , \10446 , \10456 );
buf \U$10363 ( \10458 , \10457 );
buf \U$10364 ( \10459 , \10458 );
xor \U$10365 ( \10460 , \10440 , \10459 );
buf \U$10366 ( \10461 , \7449 );
buf \U$10367 ( \10462 , \10295 );
or \U$10368 ( \10463 , \10461 , \10462 );
buf \U$10369 ( \10464 , \1232 );
buf \U$10370 ( \10465 , RIc0d7c18_13);
buf \U$10371 ( \10466 , RIc0d9478_65);
xnor \U$10372 ( \10467 , \10465 , \10466 );
buf \U$10373 ( \10468 , \10467 );
buf \U$10374 ( \10469 , \10468 );
or \U$10375 ( \10470 , \10464 , \10469 );
nand \U$10376 ( \10471 , \10463 , \10470 );
buf \U$10377 ( \10472 , \10471 );
buf \U$10378 ( \10473 , \10472 );
xor \U$10379 ( \10474 , \10460 , \10473 );
buf \U$10380 ( \10475 , \10474 );
buf \U$10381 ( \10476 , \10475 );
xor \U$10382 ( \10477 , \10431 , \10476 );
buf \U$10383 ( \10478 , \10211 );
not \U$10384 ( \10479 , \10478 );
buf \U$10385 ( \10480 , \2871 );
not \U$10386 ( \10481 , \10480 );
or \U$10387 ( \10482 , \10479 , \10481 );
buf \U$10388 ( \10483 , RIc0d7858_5);
buf \U$10389 ( \10484 , RIc0d9838_73);
xnor \U$10390 ( \10485 , \10483 , \10484 );
buf \U$10391 ( \10486 , \10485 );
buf \U$10392 ( \10487 , \10486 );
not \U$10393 ( \10488 , \10487 );
buf \U$10394 ( \10489 , \792 );
nand \U$10395 ( \10490 , \10488 , \10489 );
buf \U$10396 ( \10491 , \10490 );
buf \U$10397 ( \10492 , \10491 );
nand \U$10398 ( \10493 , \10482 , \10492 );
buf \U$10399 ( \10494 , \10493 );
buf \U$10400 ( \10495 , \10494 );
not \U$10401 ( \10496 , \10495 );
buf \U$10402 ( \10497 , \10187 );
not \U$10403 ( \10498 , \10497 );
buf \U$10404 ( \10499 , \1888 );
not \U$10405 ( \10500 , \10499 );
or \U$10406 ( \10501 , \10498 , \10500 );
buf \U$10407 ( \10502 , \2927 );
buf \U$10408 ( \10503 , RIc0d7948_7);
buf \U$10409 ( \10504 , RIc0d9748_71);
xor \U$10410 ( \10505 , \10503 , \10504 );
buf \U$10411 ( \10506 , \10505 );
buf \U$10412 ( \10507 , \10506 );
nand \U$10413 ( \10508 , \10502 , \10507 );
buf \U$10414 ( \10509 , \10508 );
buf \U$10415 ( \10510 , \10509 );
nand \U$10416 ( \10511 , \10501 , \10510 );
buf \U$10417 ( \10512 , \10511 );
buf \U$10418 ( \10513 , \10512 );
not \U$10419 ( \10514 , \10513 );
buf \U$10420 ( \10515 , \10514 );
buf \U$10421 ( \10516 , \10515 );
not \U$10422 ( \10517 , \10516 );
or \U$10423 ( \10518 , \10496 , \10517 );
buf \U$10424 ( \10519 , \10515 );
buf \U$10425 ( \10520 , \10494 );
or \U$10426 ( \10521 , \10519 , \10520 );
nand \U$10427 ( \10522 , \10518 , \10521 );
buf \U$10428 ( \10523 , \10522 );
buf \U$10429 ( \10524 , \10523 );
buf \U$10430 ( \10525 , \1452 );
buf \U$10431 ( \10526 , \10312 );
or \U$10432 ( \10527 , \10525 , \10526 );
buf \U$10433 ( \10528 , \4297 );
buf \U$10434 ( \10529 , RIc0d7a38_9);
buf \U$10435 ( \10530 , RIc0d9658_69);
xnor \U$10436 ( \10531 , \10529 , \10530 );
buf \U$10437 ( \10532 , \10531 );
buf \U$10438 ( \10533 , \10532 );
or \U$10439 ( \10534 , \10528 , \10533 );
nand \U$10440 ( \10535 , \10527 , \10534 );
buf \U$10441 ( \10536 , \10535 );
buf \U$10442 ( \10537 , \10536 );
xor \U$10443 ( \10538 , \10524 , \10537 );
buf \U$10444 ( \10539 , \10538 );
buf \U$10445 ( \10540 , \10539 );
xor \U$10446 ( \10541 , \10477 , \10540 );
buf \U$10447 ( \10542 , \10541 );
buf \U$10448 ( \10543 , \10542 );
xor \U$10449 ( \10544 , \10221 , \10273 );
and \U$10450 ( \10545 , \10544 , \10318 );
and \U$10451 ( \10546 , \10221 , \10273 );
or \U$10452 ( \10547 , \10545 , \10546 );
buf \U$10453 ( \10548 , \10547 );
buf \U$10454 ( \10549 , \10548 );
xor \U$10455 ( \10550 , \10543 , \10549 );
xor \U$10456 ( \10551 , \10118 , \10133 );
and \U$10457 ( \10552 , \10551 , \10165 );
and \U$10458 ( \10553 , \10118 , \10133 );
or \U$10459 ( \10554 , \10552 , \10553 );
buf \U$10460 ( \10555 , \10554 );
buf \U$10461 ( \10556 , \10555 );
xor \U$10462 ( \10557 , \10550 , \10556 );
buf \U$10463 ( \10558 , \10557 );
buf \U$10464 ( \10559 , \10558 );
xor \U$10465 ( \10560 , \10392 , \10559 );
xor \U$10466 ( \10561 , \10174 , \10321 );
and \U$10467 ( \10562 , \10561 , \10328 );
and \U$10468 ( \10563 , \10174 , \10321 );
or \U$10469 ( \10564 , \10562 , \10563 );
buf \U$10470 ( \10565 , \10564 );
buf \U$10471 ( \10566 , \10565 );
xor \U$10472 ( \10567 , \10560 , \10566 );
buf \U$10473 ( \10568 , \10567 );
buf \U$10474 ( \10569 , \10568 );
xor \U$10475 ( \10570 , \10168 , \10331 );
and \U$10476 ( \10571 , \10570 , \10338 );
and \U$10477 ( \10572 , \10168 , \10331 );
or \U$10478 ( \10573 , \10571 , \10572 );
buf \U$10479 ( \10574 , \10573 );
buf \U$10480 ( \10575 , \10574 );
nor \U$10481 ( \10576 , \10569 , \10575 );
buf \U$10482 ( \10577 , \10576 );
buf \U$10483 ( \10578 , \10577 );
nor \U$10484 ( \10579 , \10350 , \10578 );
buf \U$10485 ( \10580 , \10579 );
buf \U$10486 ( \10581 , \10580 );
buf \U$10487 ( \10582 , \10515 );
not \U$10488 ( \10583 , \10582 );
buf \U$10489 ( \10584 , \10494 );
not \U$10490 ( \10585 , \10584 );
buf \U$10491 ( \10586 , \10585 );
buf \U$10492 ( \10587 , \10586 );
not \U$10493 ( \10588 , \10587 );
or \U$10494 ( \10589 , \10583 , \10588 );
buf \U$10495 ( \10590 , \10536 );
nand \U$10496 ( \10591 , \10589 , \10590 );
buf \U$10497 ( \10592 , \10591 );
buf \U$10498 ( \10593 , \10592 );
buf \U$10499 ( \10594 , \10512 );
buf \U$10500 ( \10595 , \10494 );
nand \U$10501 ( \10596 , \10594 , \10595 );
buf \U$10502 ( \10597 , \10596 );
buf \U$10503 ( \10598 , \10597 );
nand \U$10504 ( \10599 , \10593 , \10598 );
buf \U$10505 ( \10600 , \10599 );
buf \U$10506 ( \10601 , \10600 );
not \U$10507 ( \10602 , \10601 );
buf \U$10508 ( \10603 , \1452 );
buf \U$10509 ( \10604 , \10532 );
or \U$10510 ( \10605 , \10603 , \10604 );
buf \U$10511 ( \10606 , \1969 );
buf \U$10512 ( \10607 , RIc0d79c0_8);
buf \U$10513 ( \10608 , RIc0d9658_69);
xor \U$10514 ( \10609 , \10607 , \10608 );
buf \U$10515 ( \10610 , \10609 );
buf \U$10516 ( \10611 , \10610 );
not \U$10517 ( \10612 , \10611 );
buf \U$10518 ( \10613 , \10612 );
buf \U$10519 ( \10614 , \10613 );
or \U$10520 ( \10615 , \10606 , \10614 );
nand \U$10521 ( \10616 , \10605 , \10615 );
buf \U$10522 ( \10617 , \10616 );
buf \U$10523 ( \10618 , \10617 );
not \U$10524 ( \10619 , \10618 );
buf \U$10525 ( \10620 , \10419 );
not \U$10526 ( \10621 , \10620 );
buf \U$10527 ( \10622 , \1432 );
not \U$10528 ( \10623 , \10622 );
or \U$10529 ( \10624 , \10621 , \10623 );
buf \U$10530 ( \10625 , \1196 );
buf \U$10531 ( \10626 , RIc0d9a18_77);
nand \U$10532 ( \10627 , \10625 , \10626 );
buf \U$10533 ( \10628 , \10627 );
buf \U$10534 ( \10629 , \10628 );
nand \U$10535 ( \10630 , \10624 , \10629 );
buf \U$10536 ( \10631 , \10630 );
buf \U$10537 ( \10632 , \10631 );
not \U$10538 ( \10633 , \10632 );
and \U$10539 ( \10634 , \10619 , \10633 );
buf \U$10540 ( \10635 , \10631 );
buf \U$10541 ( \10636 , \10617 );
and \U$10542 ( \10637 , \10635 , \10636 );
nor \U$10543 ( \10638 , \10634 , \10637 );
buf \U$10544 ( \10639 , \10638 );
buf \U$10545 ( \10640 , \10639 );
not \U$10546 ( \10641 , \10640 );
and \U$10547 ( \10642 , \10602 , \10641 );
buf \U$10548 ( \10643 , \10600 );
buf \U$10549 ( \10644 , \10639 );
and \U$10550 ( \10645 , \10643 , \10644 );
nor \U$10551 ( \10646 , \10642 , \10645 );
buf \U$10552 ( \10647 , \10646 );
buf \U$10553 ( \10648 , \10647 );
not \U$10554 ( \10649 , \10648 );
buf \U$10555 ( \10650 , \10649 );
buf \U$10556 ( \10651 , \10650 );
not \U$10557 ( \10652 , \10651 );
xor \U$10558 ( \10653 , \10364 , \10379 );
and \U$10559 ( \10654 , \10653 , \10386 );
and \U$10560 ( \10655 , \10364 , \10379 );
or \U$10561 ( \10656 , \10654 , \10655 );
buf \U$10562 ( \10657 , \10656 );
buf \U$10563 ( \10658 , \10657 );
buf \U$10564 ( \10659 , RIc0d7c90_14);
buf \U$10565 ( \10660 , RIc0d9478_65);
nand \U$10566 ( \10661 , \10659 , \10660 );
buf \U$10567 ( \10662 , \10661 );
buf \U$10568 ( \10663 , \10662 );
not \U$10569 ( \10664 , \10663 );
buf \U$10570 ( \10665 , \10451 );
not \U$10571 ( \10666 , \10665 );
buf \U$10572 ( \10667 , \1129 );
not \U$10573 ( \10668 , \10667 );
or \U$10574 ( \10669 , \10666 , \10668 );
buf \U$10575 ( \10670 , RIc0d9928_75);
buf \U$10576 ( \10671 , RIc0d76f0_2);
xnor \U$10577 ( \10672 , \10670 , \10671 );
buf \U$10578 ( \10673 , \10672 );
buf \U$10579 ( \10674 , \10673 );
not \U$10580 ( \10675 , \10674 );
buf \U$10581 ( \10676 , \1143 );
nand \U$10582 ( \10677 , \10675 , \10676 );
buf \U$10583 ( \10678 , \10677 );
buf \U$10584 ( \10679 , \10678 );
nand \U$10585 ( \10680 , \10669 , \10679 );
buf \U$10586 ( \10681 , \10680 );
buf \U$10587 ( \10682 , \10506 );
not \U$10588 ( \10683 , \10682 );
buf \U$10589 ( \10684 , \2269 );
not \U$10590 ( \10685 , \10684 );
or \U$10591 ( \10686 , \10683 , \10685 );
buf \U$10592 ( \10687 , \1282 );
buf \U$10593 ( \10688 , RIc0d78d0_6);
buf \U$10594 ( \10689 , RIc0d9748_71);
xor \U$10595 ( \10690 , \10688 , \10689 );
buf \U$10596 ( \10691 , \10690 );
buf \U$10597 ( \10692 , \10691 );
nand \U$10598 ( \10693 , \10687 , \10692 );
buf \U$10599 ( \10694 , \10693 );
buf \U$10600 ( \10695 , \10694 );
nand \U$10601 ( \10696 , \10686 , \10695 );
buf \U$10602 ( \10697 , \10696 );
xor \U$10603 ( \10698 , \10681 , \10697 );
buf \U$10604 ( \10699 , \10698 );
not \U$10605 ( \10700 , \10699 );
or \U$10606 ( \10701 , \10664 , \10700 );
buf \U$10607 ( \10702 , \10698 );
buf \U$10608 ( \10703 , \10662 );
or \U$10609 ( \10704 , \10702 , \10703 );
nand \U$10610 ( \10705 , \10701 , \10704 );
buf \U$10611 ( \10706 , \10705 );
buf \U$10612 ( \10707 , \10706 );
xnor \U$10613 ( \10708 , \10658 , \10707 );
buf \U$10614 ( \10709 , \10708 );
buf \U$10615 ( \10710 , \10709 );
not \U$10616 ( \10711 , \10710 );
or \U$10617 ( \10712 , \10652 , \10711 );
buf \U$10618 ( \10713 , \10709 );
buf \U$10619 ( \10714 , \10650 );
or \U$10620 ( \10715 , \10713 , \10714 );
nand \U$10621 ( \10716 , \10712 , \10715 );
buf \U$10622 ( \10717 , \10716 );
buf \U$10623 ( \10718 , \10717 );
xor \U$10624 ( \10719 , \10431 , \10476 );
and \U$10625 ( \10720 , \10719 , \10540 );
and \U$10626 ( \10721 , \10431 , \10476 );
or \U$10627 ( \10722 , \10720 , \10721 );
buf \U$10628 ( \10723 , \10722 );
buf \U$10629 ( \10724 , \10723 );
xor \U$10630 ( \10725 , \10395 , \10412 );
and \U$10631 ( \10726 , \10725 , \10428 );
and \U$10632 ( \10727 , \10395 , \10412 );
or \U$10633 ( \10728 , \10726 , \10727 );
buf \U$10634 ( \10729 , \10728 );
buf \U$10635 ( \10730 , \10729 );
xor \U$10636 ( \10731 , \10440 , \10459 );
and \U$10637 ( \10732 , \10731 , \10473 );
and \U$10638 ( \10733 , \10440 , \10459 );
or \U$10639 ( \10734 , \10732 , \10733 );
buf \U$10640 ( \10735 , \10734 );
buf \U$10641 ( \10736 , \10735 );
xor \U$10642 ( \10737 , \10730 , \10736 );
buf \U$10643 ( \10738 , \10405 );
not \U$10644 ( \10739 , \10738 );
buf \U$10645 ( \10740 , \1414 );
not \U$10646 ( \10741 , \10740 );
or \U$10647 ( \10742 , \10739 , \10741 );
buf \U$10648 ( \10743 , \686 );
buf \U$10649 ( \10744 , RIc0d7ab0_10);
buf \U$10650 ( \10745 , RIc0d9568_67);
xor \U$10651 ( \10746 , \10744 , \10745 );
buf \U$10652 ( \10747 , \10746 );
buf \U$10653 ( \10748 , \10747 );
nand \U$10654 ( \10749 , \10743 , \10748 );
buf \U$10655 ( \10750 , \10749 );
buf \U$10656 ( \10751 , \10750 );
nand \U$10657 ( \10752 , \10742 , \10751 );
buf \U$10658 ( \10753 , \10752 );
buf \U$10659 ( \10754 , \10753 );
buf \U$10660 ( \10755 , \10468 );
not \U$10661 ( \10756 , \10755 );
buf \U$10662 ( \10757 , \10756 );
buf \U$10663 ( \10758 , \10757 );
not \U$10664 ( \10759 , \10758 );
buf \U$10665 ( \10760 , \3781 );
not \U$10666 ( \10761 , \10760 );
or \U$10667 ( \10762 , \10759 , \10761 );
buf \U$10668 ( \10763 , \1229 );
buf \U$10669 ( \10764 , RIc0d9478_65);
buf \U$10670 ( \10765 , RIc0d7ba0_12);
xor \U$10671 ( \10766 , \10764 , \10765 );
buf \U$10672 ( \10767 , \10766 );
buf \U$10673 ( \10768 , \10767 );
nand \U$10674 ( \10769 , \10763 , \10768 );
buf \U$10675 ( \10770 , \10769 );
buf \U$10676 ( \10771 , \10770 );
nand \U$10677 ( \10772 , \10762 , \10771 );
buf \U$10678 ( \10773 , \10772 );
buf \U$10679 ( \10774 , \10773 );
xor \U$10680 ( \10775 , \10754 , \10774 );
buf \U$10681 ( \10776 , \773 );
buf \U$10682 ( \10777 , \10486 );
or \U$10683 ( \10778 , \10776 , \10777 );
buf \U$10684 ( \10779 , \9493 );
buf \U$10685 ( \10780 , RIc0d77e0_4);
buf \U$10686 ( \10781 , RIc0d9838_73);
xor \U$10687 ( \10782 , \10780 , \10781 );
buf \U$10688 ( \10783 , \10782 );
buf \U$10689 ( \10784 , \10783 );
not \U$10690 ( \10785 , \10784 );
buf \U$10691 ( \10786 , \10785 );
buf \U$10692 ( \10787 , \10786 );
or \U$10693 ( \10788 , \10779 , \10787 );
nand \U$10694 ( \10789 , \10778 , \10788 );
buf \U$10695 ( \10790 , \10789 );
buf \U$10696 ( \10791 , \10790 );
xor \U$10697 ( \10792 , \10775 , \10791 );
buf \U$10698 ( \10793 , \10792 );
buf \U$10699 ( \10794 , \10793 );
xor \U$10700 ( \10795 , \10737 , \10794 );
buf \U$10701 ( \10796 , \10795 );
buf \U$10702 ( \10797 , \10796 );
xor \U$10703 ( \10798 , \10724 , \10797 );
xor \U$10704 ( \10799 , \10356 , \10362 );
and \U$10705 ( \10800 , \10799 , \10389 );
and \U$10706 ( \10801 , \10356 , \10362 );
or \U$10707 ( \10802 , \10800 , \10801 );
buf \U$10708 ( \10803 , \10802 );
buf \U$10709 ( \10804 , \10803 );
xor \U$10710 ( \10805 , \10798 , \10804 );
buf \U$10711 ( \10806 , \10805 );
buf \U$10712 ( \10807 , \10806 );
xor \U$10713 ( \10808 , \10718 , \10807 );
xor \U$10714 ( \10809 , \10543 , \10549 );
and \U$10715 ( \10810 , \10809 , \10556 );
and \U$10716 ( \10811 , \10543 , \10549 );
or \U$10717 ( \10812 , \10810 , \10811 );
buf \U$10718 ( \10813 , \10812 );
buf \U$10719 ( \10814 , \10813 );
xor \U$10720 ( \10815 , \10808 , \10814 );
buf \U$10721 ( \10816 , \10815 );
buf \U$10722 ( \10817 , \10816 );
xor \U$10723 ( \10818 , \10392 , \10559 );
and \U$10724 ( \10819 , \10818 , \10566 );
and \U$10725 ( \10820 , \10392 , \10559 );
or \U$10726 ( \10821 , \10819 , \10820 );
buf \U$10727 ( \10822 , \10821 );
buf \U$10728 ( \10823 , \10822 );
or \U$10729 ( \10824 , \10817 , \10823 );
buf \U$10730 ( \10825 , \10824 );
buf \U$10731 ( \10826 , \10825 );
nand \U$10732 ( \10827 , \10581 , \10826 );
buf \U$10733 ( \10828 , \10827 );
buf \U$10734 ( \10829 , \10828 );
xor \U$10735 ( \10830 , \10718 , \10807 );
and \U$10736 ( \10831 , \10830 , \10814 );
and \U$10737 ( \10832 , \10718 , \10807 );
or \U$10738 ( \10833 , \10831 , \10832 );
buf \U$10739 ( \10834 , \10833 );
buf \U$10740 ( \10835 , \10834 );
buf \U$10741 ( \10836 , \10631 );
not \U$10742 ( \10837 , \10836 );
buf \U$10743 ( \10838 , \10837 );
buf \U$10744 ( \10839 , \10838 );
not \U$10745 ( \10840 , \10839 );
buf \U$10746 ( \10841 , \10767 );
not \U$10747 ( \10842 , \10841 );
buf \U$10748 ( \10843 , \1225 );
not \U$10749 ( \10844 , \10843 );
or \U$10750 ( \10845 , \10842 , \10844 );
buf \U$10751 ( \10846 , RIc0d7b28_11);
buf \U$10752 ( \10847 , RIc0d9478_65);
xnor \U$10753 ( \10848 , \10846 , \10847 );
buf \U$10754 ( \10849 , \10848 );
buf \U$10755 ( \10850 , \10849 );
not \U$10756 ( \10851 , \10850 );
buf \U$10757 ( \10852 , \1229 );
nand \U$10758 ( \10853 , \10851 , \10852 );
buf \U$10759 ( \10854 , \10853 );
buf \U$10760 ( \10855 , \10854 );
nand \U$10761 ( \10856 , \10845 , \10855 );
buf \U$10762 ( \10857 , \10856 );
buf \U$10763 ( \10858 , \10691 );
not \U$10764 ( \10859 , \10858 );
buf \U$10765 ( \10860 , \2812 );
not \U$10766 ( \10861 , \10860 );
or \U$10767 ( \10862 , \10859 , \10861 );
buf \U$10768 ( \10863 , RIc0d7858_5);
buf \U$10769 ( \10864 , RIc0d9748_71);
xnor \U$10770 ( \10865 , \10863 , \10864 );
buf \U$10771 ( \10866 , \10865 );
buf \U$10772 ( \10867 , \10866 );
not \U$10773 ( \10868 , \10867 );
buf \U$10774 ( \10869 , \1282 );
nand \U$10775 ( \10870 , \10868 , \10869 );
buf \U$10776 ( \10871 , \10870 );
buf \U$10777 ( \10872 , \10871 );
nand \U$10778 ( \10873 , \10862 , \10872 );
buf \U$10779 ( \10874 , \10873 );
xor \U$10780 ( \10875 , \10857 , \10874 );
buf \U$10781 ( \10876 , \10875 );
not \U$10782 ( \10877 , \10876 );
or \U$10783 ( \10878 , \10840 , \10877 );
buf \U$10784 ( \10879 , \10875 );
buf \U$10785 ( \10880 , \10838 );
or \U$10786 ( \10881 , \10879 , \10880 );
nand \U$10787 ( \10882 , \10878 , \10881 );
buf \U$10788 ( \10883 , \10882 );
buf \U$10789 ( \10884 , \10883 );
buf \U$10790 ( \10885 , \1126 );
buf \U$10791 ( \10886 , \10673 );
or \U$10792 ( \10887 , \10885 , \10886 );
buf \U$10793 ( \10888 , \1370 );
buf \U$10794 ( \10889 , RIc0d7678_1);
buf \U$10795 ( \10890 , RIc0d9928_75);
xnor \U$10796 ( \10891 , \10889 , \10890 );
buf \U$10797 ( \10892 , \10891 );
buf \U$10798 ( \10893 , \10892 );
or \U$10799 ( \10894 , \10888 , \10893 );
nand \U$10800 ( \10895 , \10887 , \10894 );
buf \U$10801 ( \10896 , \10895 );
buf \U$10802 ( \10897 , \10610 );
not \U$10803 ( \10898 , \10897 );
buf \U$10804 ( \10899 , \279 );
not \U$10805 ( \10900 , \10899 );
or \U$10806 ( \10901 , \10898 , \10900 );
buf \U$10807 ( \10902 , RIc0d7948_7);
buf \U$10808 ( \10903 , RIc0d9658_69);
xnor \U$10809 ( \10904 , \10902 , \10903 );
buf \U$10810 ( \10905 , \10904 );
buf \U$10811 ( \10906 , \10905 );
not \U$10812 ( \10907 , \10906 );
buf \U$10813 ( \10908 , \284 );
nand \U$10814 ( \10909 , \10907 , \10908 );
buf \U$10815 ( \10910 , \10909 );
buf \U$10816 ( \10911 , \10910 );
nand \U$10817 ( \10912 , \10901 , \10911 );
buf \U$10818 ( \10913 , \10912 );
buf \U$10819 ( \10914 , \10783 );
not \U$10820 ( \10915 , \10914 );
buf \U$10821 ( \10916 , \1677 );
not \U$10822 ( \10917 , \10916 );
or \U$10823 ( \10918 , \10915 , \10917 );
buf \U$10824 ( \10919 , \1856 );
buf \U$10825 ( \10920 , RIc0d7768_3);
buf \U$10826 ( \10921 , RIc0d9838_73);
xor \U$10827 ( \10922 , \10920 , \10921 );
buf \U$10828 ( \10923 , \10922 );
buf \U$10829 ( \10924 , \10923 );
nand \U$10830 ( \10925 , \10919 , \10924 );
buf \U$10831 ( \10926 , \10925 );
buf \U$10832 ( \10927 , \10926 );
nand \U$10833 ( \10928 , \10918 , \10927 );
buf \U$10834 ( \10929 , \10928 );
xor \U$10835 ( \10930 , \10913 , \10929 );
xor \U$10836 ( \10931 , \10896 , \10930 );
buf \U$10837 ( \10932 , \10931 );
xor \U$10838 ( \10933 , \10884 , \10932 );
buf \U$10839 ( \10934 , \10617 );
not \U$10840 ( \10935 , \10934 );
buf \U$10841 ( \10936 , \10838 );
not \U$10842 ( \10937 , \10936 );
or \U$10843 ( \10938 , \10935 , \10937 );
buf \U$10844 ( \10939 , \10838 );
buf \U$10845 ( \10940 , \10617 );
or \U$10846 ( \10941 , \10939 , \10940 );
buf \U$10847 ( \10942 , \10600 );
nand \U$10848 ( \10943 , \10941 , \10942 );
buf \U$10849 ( \10944 , \10943 );
buf \U$10850 ( \10945 , \10944 );
nand \U$10851 ( \10946 , \10938 , \10945 );
buf \U$10852 ( \10947 , \10946 );
buf \U$10853 ( \10948 , \10947 );
xor \U$10854 ( \10949 , \10933 , \10948 );
buf \U$10855 ( \10950 , \10949 );
buf \U$10856 ( \10951 , \10950 );
xor \U$10857 ( \10952 , \10730 , \10736 );
and \U$10858 ( \10953 , \10952 , \10794 );
and \U$10859 ( \10954 , \10730 , \10736 );
or \U$10860 ( \10955 , \10953 , \10954 );
buf \U$10861 ( \10956 , \10955 );
buf \U$10862 ( \10957 , \10956 );
buf \U$10863 ( \10958 , \10681 );
buf \U$10864 ( \10959 , \10662 );
not \U$10865 ( \10960 , \10959 );
buf \U$10866 ( \10961 , \10960 );
buf \U$10867 ( \10962 , \10961 );
or \U$10868 ( \10963 , \10958 , \10962 );
buf \U$10869 ( \10964 , \10697 );
nand \U$10870 ( \10965 , \10963 , \10964 );
buf \U$10871 ( \10966 , \10965 );
buf \U$10872 ( \10967 , \10966 );
buf \U$10873 ( \10968 , \10681 );
buf \U$10874 ( \10969 , \10961 );
nand \U$10875 ( \10970 , \10968 , \10969 );
buf \U$10876 ( \10971 , \10970 );
buf \U$10877 ( \10972 , \10971 );
nand \U$10878 ( \10973 , \10967 , \10972 );
buf \U$10879 ( \10974 , \10973 );
buf \U$10880 ( \10975 , \10974 );
buf \U$10881 ( \10976 , RIc0d7c18_13);
buf \U$10882 ( \10977 , RIc0d9478_65);
and \U$10883 ( \10978 , \10976 , \10977 );
buf \U$10884 ( \10979 , \10978 );
buf \U$10885 ( \10980 , \10979 );
buf \U$10886 ( \10981 , \10747 );
not \U$10887 ( \10982 , \10981 );
buf \U$10888 ( \10983 , \10034 );
not \U$10889 ( \10984 , \10983 );
or \U$10890 ( \10985 , \10982 , \10984 );
buf \U$10891 ( \10986 , \686 );
buf \U$10892 ( \10987 , RIc0d7a38_9);
buf \U$10893 ( \10988 , RIc0d9568_67);
xor \U$10894 ( \10989 , \10987 , \10988 );
buf \U$10895 ( \10990 , \10989 );
buf \U$10896 ( \10991 , \10990 );
nand \U$10897 ( \10992 , \10986 , \10991 );
buf \U$10898 ( \10993 , \10992 );
buf \U$10899 ( \10994 , \10993 );
nand \U$10900 ( \10995 , \10985 , \10994 );
buf \U$10901 ( \10996 , \10995 );
buf \U$10902 ( \10997 , \10996 );
xor \U$10903 ( \10998 , \10980 , \10997 );
buf \U$10904 ( \10999 , \1193 );
not \U$10905 ( \11000 , \10999 );
buf \U$10906 ( \11001 , \1435 );
not \U$10907 ( \11002 , \11001 );
or \U$10908 ( \11003 , \11000 , \11002 );
buf \U$10909 ( \11004 , RIc0d9a18_77);
nand \U$10910 ( \11005 , \11003 , \11004 );
buf \U$10911 ( \11006 , \11005 );
buf \U$10912 ( \11007 , \11006 );
xor \U$10913 ( \11008 , \10998 , \11007 );
buf \U$10914 ( \11009 , \11008 );
buf \U$10915 ( \11010 , \11009 );
xor \U$10916 ( \11011 , \10975 , \11010 );
xor \U$10917 ( \11012 , \10754 , \10774 );
and \U$10918 ( \11013 , \11012 , \10791 );
and \U$10919 ( \11014 , \10754 , \10774 );
or \U$10920 ( \11015 , \11013 , \11014 );
buf \U$10921 ( \11016 , \11015 );
buf \U$10922 ( \11017 , \11016 );
xor \U$10923 ( \11018 , \11011 , \11017 );
buf \U$10924 ( \11019 , \11018 );
buf \U$10925 ( \11020 , \11019 );
xor \U$10926 ( \11021 , \10957 , \11020 );
buf \U$10927 ( \11022 , \10706 );
not \U$10928 ( \11023 , \11022 );
buf \U$10929 ( \11024 , \10650 );
not \U$10930 ( \11025 , \11024 );
or \U$10931 ( \11026 , \11023 , \11025 );
buf \U$10932 ( \11027 , \10706 );
not \U$10933 ( \11028 , \11027 );
buf \U$10934 ( \11029 , \10647 );
nand \U$10935 ( \11030 , \11028 , \11029 );
buf \U$10936 ( \11031 , \11030 );
buf \U$10937 ( \11032 , \11031 );
buf \U$10938 ( \11033 , \10657 );
nand \U$10939 ( \11034 , \11032 , \11033 );
buf \U$10940 ( \11035 , \11034 );
buf \U$10941 ( \11036 , \11035 );
nand \U$10942 ( \11037 , \11026 , \11036 );
buf \U$10943 ( \11038 , \11037 );
buf \U$10944 ( \11039 , \11038 );
xor \U$10945 ( \11040 , \11021 , \11039 );
buf \U$10946 ( \11041 , \11040 );
buf \U$10947 ( \11042 , \11041 );
xor \U$10948 ( \11043 , \10951 , \11042 );
xor \U$10949 ( \11044 , \10724 , \10797 );
and \U$10950 ( \11045 , \11044 , \10804 );
and \U$10951 ( \11046 , \10724 , \10797 );
or \U$10952 ( \11047 , \11045 , \11046 );
buf \U$10953 ( \11048 , \11047 );
buf \U$10954 ( \11049 , \11048 );
xor \U$10955 ( \11050 , \11043 , \11049 );
buf \U$10956 ( \11051 , \11050 );
buf \U$10957 ( \11052 , \11051 );
nor \U$10958 ( \11053 , \10835 , \11052 );
buf \U$10959 ( \11054 , \11053 );
buf \U$10960 ( \11055 , \11054 );
nor \U$10961 ( \11056 , \10829 , \11055 );
buf \U$10962 ( \11057 , \11056 );
buf \U$10963 ( \11058 , \11057 );
buf \U$10964 ( \11059 , \2362 );
buf \U$10965 ( \11060 , \10892 );
or \U$10966 ( \11061 , \11059 , \11060 );
buf \U$10967 ( \11062 , \1370 );
buf \U$10968 ( \11063 , \763 );
or \U$10969 ( \11064 , \11062 , \11063 );
nand \U$10970 ( \11065 , \11061 , \11064 );
buf \U$10971 ( \11066 , \11065 );
buf \U$10972 ( \11067 , \11066 );
buf \U$10973 ( \11068 , \9922 );
buf \U$10974 ( \11069 , RIc0d76f0_2);
buf \U$10975 ( \11070 , RIc0d9838_73);
xnor \U$10976 ( \11071 , \11069 , \11070 );
buf \U$10977 ( \11072 , \11071 );
buf \U$10978 ( \11073 , \11072 );
or \U$10979 ( \11074 , \11068 , \11073 );
buf \U$10980 ( \11075 , \2879 );
buf \U$10981 ( \11076 , RIc0d9838_73);
buf \U$10982 ( \11077 , \974 );
and \U$10983 ( \11078 , \11076 , \11077 );
not \U$10984 ( \11079 , \11076 );
buf \U$10985 ( \11080 , RIc0d7678_1);
and \U$10986 ( \11081 , \11079 , \11080 );
nor \U$10987 ( \11082 , \11078 , \11081 );
buf \U$10988 ( \11083 , \11082 );
buf \U$10989 ( \11084 , \11083 );
or \U$10990 ( \11085 , \11075 , \11084 );
nand \U$10991 ( \11086 , \11074 , \11085 );
buf \U$10992 ( \11087 , \11086 );
buf \U$10993 ( \11088 , \11087 );
xor \U$10994 ( \11089 , \11067 , \11088 );
and \U$10995 ( \11090 , \10764 , \10765 );
buf \U$10996 ( \11091 , \11090 );
buf \U$10997 ( \11092 , \11091 );
buf \U$10998 ( \11093 , \10990 );
not \U$10999 ( \11094 , \11093 );
buf \U$11000 ( \11095 , \2900 );
not \U$11001 ( \11096 , \11095 );
or \U$11002 ( \11097 , \11094 , \11096 );
buf \U$11003 ( \11098 , RIc0d9568_67);
buf \U$11004 ( \11099 , RIc0d79c0_8);
xnor \U$11005 ( \11100 , \11098 , \11099 );
buf \U$11006 ( \11101 , \11100 );
buf \U$11007 ( \11102 , \11101 );
not \U$11008 ( \11103 , \11102 );
buf \U$11009 ( \11104 , \686 );
nand \U$11010 ( \11105 , \11103 , \11104 );
buf \U$11011 ( \11106 , \11105 );
buf \U$11012 ( \11107 , \11106 );
nand \U$11013 ( \11108 , \11097 , \11107 );
buf \U$11014 ( \11109 , \11108 );
buf \U$11015 ( \11110 , \11109 );
xor \U$11016 ( \11111 , \11092 , \11110 );
buf \U$11017 ( \11112 , \10923 );
not \U$11018 ( \11113 , \11112 );
buf \U$11019 ( \11114 , \776 );
not \U$11020 ( \11115 , \11114 );
or \U$11021 ( \11116 , \11113 , \11115 );
buf \U$11022 ( \11117 , \11072 );
not \U$11023 ( \11118 , \11117 );
buf \U$11024 ( \11119 , \1856 );
nand \U$11025 ( \11120 , \11118 , \11119 );
buf \U$11026 ( \11121 , \11120 );
buf \U$11027 ( \11122 , \11121 );
nand \U$11028 ( \11123 , \11116 , \11122 );
buf \U$11029 ( \11124 , \11123 );
buf \U$11030 ( \11125 , \11124 );
and \U$11031 ( \11126 , \11111 , \11125 );
and \U$11032 ( \11127 , \11092 , \11110 );
or \U$11033 ( \11128 , \11126 , \11127 );
buf \U$11034 ( \11129 , \11128 );
buf \U$11035 ( \11130 , \11129 );
xor \U$11036 ( \11131 , \11089 , \11130 );
buf \U$11037 ( \11132 , \11131 );
buf \U$11038 ( \11133 , \11132 );
buf \U$11039 ( \11134 , \11066 );
not \U$11040 ( \11135 , \11134 );
buf \U$11041 ( \11136 , \11135 );
buf \U$11042 ( \11137 , \11136 );
buf \U$11043 ( \11138 , \10929 );
not \U$11044 ( \11139 , \11138 );
buf \U$11045 ( \11140 , \10913 );
not \U$11046 ( \11141 , \11140 );
or \U$11047 ( \11142 , \11139 , \11141 );
buf \U$11048 ( \11143 , \10913 );
buf \U$11049 ( \11144 , \10929 );
or \U$11050 ( \11145 , \11143 , \11144 );
buf \U$11051 ( \11146 , \10896 );
nand \U$11052 ( \11147 , \11145 , \11146 );
buf \U$11053 ( \11148 , \11147 );
buf \U$11054 ( \11149 , \11148 );
nand \U$11055 ( \11150 , \11142 , \11149 );
buf \U$11056 ( \11151 , \11150 );
buf \U$11057 ( \11152 , \11151 );
xor \U$11058 ( \11153 , \11137 , \11152 );
xor \U$11059 ( \11154 , \10980 , \10997 );
and \U$11060 ( \11155 , \11154 , \11007 );
and \U$11061 ( \11156 , \10980 , \10997 );
or \U$11062 ( \11157 , \11155 , \11156 );
buf \U$11063 ( \11158 , \11157 );
buf \U$11064 ( \11159 , \11158 );
and \U$11065 ( \11160 , \11153 , \11159 );
and \U$11066 ( \11161 , \11137 , \11152 );
or \U$11067 ( \11162 , \11160 , \11161 );
buf \U$11068 ( \11163 , \11162 );
buf \U$11069 ( \11164 , \11163 );
xor \U$11070 ( \11165 , \11133 , \11164 );
buf \U$11071 ( \11166 , \10631 );
buf \U$11072 ( \11167 , \10874 );
or \U$11073 ( \11168 , \11166 , \11167 );
buf \U$11074 ( \11169 , \10857 );
nand \U$11075 ( \11170 , \11168 , \11169 );
buf \U$11076 ( \11171 , \11170 );
buf \U$11077 ( \11172 , \11171 );
buf \U$11078 ( \11173 , \10631 );
buf \U$11079 ( \11174 , \10874 );
nand \U$11080 ( \11175 , \11173 , \11174 );
buf \U$11081 ( \11176 , \11175 );
buf \U$11082 ( \11177 , \11176 );
nand \U$11083 ( \11178 , \11172 , \11177 );
buf \U$11084 ( \11179 , \11178 );
buf \U$11085 ( \11180 , \11179 );
xor \U$11086 ( \11181 , \11092 , \11110 );
xor \U$11087 ( \11182 , \11181 , \11125 );
buf \U$11088 ( \11183 , \11182 );
buf \U$11089 ( \11184 , \11183 );
xor \U$11090 ( \11185 , \11180 , \11184 );
buf \U$11091 ( \11186 , \7449 );
buf \U$11092 ( \11187 , \10849 );
or \U$11093 ( \11188 , \11186 , \11187 );
buf \U$11094 ( \11189 , \1232 );
buf \U$11095 ( \11190 , RIc0d7ab0_10);
buf \U$11096 ( \11191 , RIc0d9478_65);
xnor \U$11097 ( \11192 , \11190 , \11191 );
buf \U$11098 ( \11193 , \11192 );
buf \U$11099 ( \11194 , \11193 );
or \U$11100 ( \11195 , \11189 , \11194 );
nand \U$11101 ( \11196 , \11188 , \11195 );
buf \U$11102 ( \11197 , \11196 );
buf \U$11103 ( \11198 , \11197 );
buf \U$11104 ( \11199 , \1260 );
buf \U$11105 ( \11200 , \10866 );
or \U$11106 ( \11201 , \11199 , \11200 );
buf \U$11107 ( \11202 , \1279 );
buf \U$11108 ( \11203 , \263 );
buf \U$11109 ( \11204 , RIc0d77e0_4);
and \U$11110 ( \11205 , \11203 , \11204 );
buf \U$11111 ( \11206 , \489 );
buf \U$11112 ( \11207 , RIc0d9748_71);
and \U$11113 ( \11208 , \11206 , \11207 );
nor \U$11114 ( \11209 , \11205 , \11208 );
buf \U$11115 ( \11210 , \11209 );
buf \U$11116 ( \11211 , \11210 );
or \U$11117 ( \11212 , \11202 , \11211 );
nand \U$11118 ( \11213 , \11201 , \11212 );
buf \U$11119 ( \11214 , \11213 );
buf \U$11120 ( \11215 , \11214 );
xor \U$11121 ( \11216 , \11198 , \11215 );
buf \U$11122 ( \11217 , \1452 );
buf \U$11123 ( \11218 , \10905 );
or \U$11124 ( \11219 , \11217 , \11218 );
buf \U$11125 ( \11220 , \1969 );
buf \U$11126 ( \11221 , RIc0d9658_69);
buf \U$11127 ( \11222 , RIc0d78d0_6);
not \U$11128 ( \11223 , \11222 );
buf \U$11129 ( \11224 , \11223 );
buf \U$11130 ( \11225 , \11224 );
and \U$11131 ( \11226 , \11221 , \11225 );
not \U$11132 ( \11227 , \11221 );
buf \U$11133 ( \11228 , RIc0d78d0_6);
and \U$11134 ( \11229 , \11227 , \11228 );
nor \U$11135 ( \11230 , \11226 , \11229 );
buf \U$11136 ( \11231 , \11230 );
buf \U$11137 ( \11232 , \11231 );
or \U$11138 ( \11233 , \11220 , \11232 );
nand \U$11139 ( \11234 , \11219 , \11233 );
buf \U$11140 ( \11235 , \11234 );
buf \U$11141 ( \11236 , \11235 );
xor \U$11142 ( \11237 , \11216 , \11236 );
buf \U$11143 ( \11238 , \11237 );
buf \U$11144 ( \11239 , \11238 );
and \U$11145 ( \11240 , \11185 , \11239 );
and \U$11146 ( \11241 , \11180 , \11184 );
or \U$11147 ( \11242 , \11240 , \11241 );
buf \U$11148 ( \11243 , \11242 );
buf \U$11149 ( \11244 , \11243 );
and \U$11150 ( \11245 , \11165 , \11244 );
and \U$11151 ( \11246 , \11133 , \11164 );
or \U$11152 ( \11247 , \11245 , \11246 );
buf \U$11153 ( \11248 , \11247 );
buf \U$11154 ( \11249 , \11248 );
buf \U$11155 ( \11250 , \7449 );
buf \U$11156 ( \11251 , \11193 );
or \U$11157 ( \11252 , \11250 , \11251 );
buf \U$11158 ( \11253 , \1232 );
buf \U$11159 ( \11254 , \7456 );
buf \U$11160 ( \11255 , RIc0d7a38_9);
and \U$11161 ( \11256 , \11254 , \11255 );
buf \U$11162 ( \11257 , \5976 );
buf \U$11163 ( \11258 , RIc0d9478_65);
and \U$11164 ( \11259 , \11257 , \11258 );
nor \U$11165 ( \11260 , \11256 , \11259 );
buf \U$11166 ( \11261 , \11260 );
buf \U$11167 ( \11262 , \11261 );
or \U$11168 ( \11263 , \11253 , \11262 );
nand \U$11169 ( \11264 , \11252 , \11263 );
buf \U$11170 ( \11265 , \11264 );
buf \U$11171 ( \11266 , \11265 );
buf \U$11172 ( \11267 , \2372 );
not \U$11173 ( \11268 , \11267 );
buf \U$11174 ( \11269 , \3816 );
not \U$11175 ( \11270 , \11269 );
or \U$11176 ( \11271 , \11268 , \11270 );
buf \U$11177 ( \11272 , RIc0d9928_75);
nand \U$11178 ( \11273 , \11271 , \11272 );
buf \U$11179 ( \11274 , \11273 );
buf \U$11180 ( \11275 , \11274 );
xor \U$11181 ( \11276 , \11266 , \11275 );
buf \U$11182 ( \11277 , RIc0d7768_3);
buf \U$11183 ( \11278 , RIc0d9748_71);
xor \U$11184 ( \11279 , \11277 , \11278 );
buf \U$11185 ( \11280 , \11279 );
buf \U$11186 ( \11281 , \11280 );
not \U$11187 ( \11282 , \11281 );
buf \U$11188 ( \11283 , \1282 );
not \U$11189 ( \11284 , \11283 );
or \U$11190 ( \11285 , \11282 , \11284 );
buf \U$11191 ( \11286 , \4868 );
buf \U$11192 ( \11287 , \11210 );
or \U$11193 ( \11288 , \11286 , \11287 );
nand \U$11194 ( \11289 , \11285 , \11288 );
buf \U$11195 ( \11290 , \11289 );
buf \U$11196 ( \11291 , \11290 );
and \U$11197 ( \11292 , \11276 , \11291 );
and \U$11198 ( \11293 , \11266 , \11275 );
or \U$11199 ( \11294 , \11292 , \11293 );
buf \U$11200 ( \11295 , \11294 );
buf \U$11201 ( \11296 , \11295 );
buf \U$11202 ( \11297 , RIc0d7b28_11);
buf \U$11203 ( \11298 , RIc0d9478_65);
and \U$11204 ( \11299 , \11297 , \11298 );
buf \U$11205 ( \11300 , \11299 );
buf \U$11206 ( \11301 , \1417 );
buf \U$11207 ( \11302 , \11101 );
or \U$11208 ( \11303 , \11301 , \11302 );
buf \U$11209 ( \11304 , \6437 );
buf \U$11210 ( \11305 , RIc0d9568_67);
not \U$11211 ( \11306 , \11305 );
buf \U$11212 ( \11307 , \11306 );
buf \U$11213 ( \11308 , \11307 );
buf \U$11214 ( \11309 , RIc0d7948_7);
and \U$11215 ( \11310 , \11308 , \11309 );
buf \U$11216 ( \11311 , RIc0d7948_7);
not \U$11217 ( \11312 , \11311 );
buf \U$11218 ( \11313 , \11312 );
buf \U$11219 ( \11314 , \11313 );
buf \U$11220 ( \11315 , RIc0d9568_67);
and \U$11221 ( \11316 , \11314 , \11315 );
nor \U$11222 ( \11317 , \11310 , \11316 );
buf \U$11223 ( \11318 , \11317 );
buf \U$11224 ( \11319 , \11318 );
or \U$11225 ( \11320 , \11304 , \11319 );
nand \U$11226 ( \11321 , \11303 , \11320 );
buf \U$11227 ( \11322 , \11321 );
xor \U$11228 ( \11323 , \11300 , \11322 );
buf \U$11229 ( \11324 , \1452 );
buf \U$11230 ( \11325 , \11231 );
or \U$11231 ( \11326 , \11324 , \11325 );
buf \U$11232 ( \11327 , \1969 );
buf \U$11233 ( \11328 , RIc0d9658_69);
buf \U$11234 ( \11329 , \1990 );
and \U$11235 ( \11330 , \11328 , \11329 );
not \U$11236 ( \11331 , \11328 );
buf \U$11237 ( \11332 , RIc0d7858_5);
and \U$11238 ( \11333 , \11331 , \11332 );
nor \U$11239 ( \11334 , \11330 , \11333 );
buf \U$11240 ( \11335 , \11334 );
buf \U$11241 ( \11336 , \11335 );
or \U$11242 ( \11337 , \11327 , \11336 );
nand \U$11243 ( \11338 , \11326 , \11337 );
buf \U$11244 ( \11339 , \11338 );
and \U$11245 ( \11340 , \11323 , \11339 );
and \U$11246 ( \11341 , \11300 , \11322 );
or \U$11247 ( \11342 , \11340 , \11341 );
buf \U$11248 ( \11343 , \11342 );
xor \U$11249 ( \11344 , \11296 , \11343 );
buf \U$11250 ( \11345 , \773 );
buf \U$11251 ( \11346 , \11083 );
or \U$11252 ( \11347 , \11345 , \11346 );
buf \U$11253 ( \11348 , \9493 );
buf \U$11254 ( \11349 , RIc0d9838_73);
not \U$11255 ( \11350 , \11349 );
buf \U$11256 ( \11351 , \11350 );
buf \U$11257 ( \11352 , \11351 );
or \U$11258 ( \11353 , \11348 , \11352 );
nand \U$11259 ( \11354 , \11347 , \11353 );
buf \U$11260 ( \11355 , \11354 );
buf \U$11261 ( \11356 , \11355 );
buf \U$11262 ( \11357 , RIc0d7ab0_10);
buf \U$11263 ( \11358 , RIc0d9478_65);
and \U$11264 ( \11359 , \11357 , \11358 );
buf \U$11265 ( \11360 , \11359 );
buf \U$11266 ( \11361 , \11360 );
xor \U$11267 ( \11362 , \11356 , \11361 );
buf \U$11268 ( \11363 , \1452 );
buf \U$11269 ( \11364 , \11335 );
or \U$11270 ( \11365 , \11363 , \11364 );
buf \U$11271 ( \11366 , \1969 );
buf \U$11272 ( \11367 , RIc0d9658_69);
buf \U$11273 ( \11368 , \489 );
and \U$11274 ( \11369 , \11367 , \11368 );
not \U$11275 ( \11370 , \11367 );
buf \U$11276 ( \11371 , RIc0d77e0_4);
and \U$11277 ( \11372 , \11370 , \11371 );
nor \U$11278 ( \11373 , \11369 , \11372 );
buf \U$11279 ( \11374 , \11373 );
buf \U$11280 ( \11375 , \11374 );
or \U$11281 ( \11376 , \11366 , \11375 );
nand \U$11282 ( \11377 , \11365 , \11376 );
buf \U$11283 ( \11378 , \11377 );
buf \U$11284 ( \11379 , \11378 );
xor \U$11285 ( \11380 , \11362 , \11379 );
buf \U$11286 ( \11381 , \11380 );
buf \U$11287 ( \11382 , \11381 );
xor \U$11288 ( \11383 , \11344 , \11382 );
buf \U$11289 ( \11384 , \11383 );
buf \U$11290 ( \11385 , \11384 );
xor \U$11291 ( \11386 , \11249 , \11385 );
xor \U$11292 ( \11387 , \11067 , \11088 );
and \U$11293 ( \11388 , \11387 , \11130 );
and \U$11294 ( \11389 , \11067 , \11088 );
or \U$11295 ( \11390 , \11388 , \11389 );
buf \U$11296 ( \11391 , \11390 );
buf \U$11297 ( \11392 , \11391 );
buf \U$11298 ( \11393 , \7449 );
buf \U$11299 ( \11394 , \11261 );
or \U$11300 ( \11395 , \11393 , \11394 );
buf \U$11301 ( \11396 , \1232 );
buf \U$11302 ( \11397 , \7456 );
buf \U$11303 ( \11398 , RIc0d79c0_8);
and \U$11304 ( \11399 , \11397 , \11398 );
buf \U$11305 ( \11400 , \4448 );
buf \U$11306 ( \11401 , RIc0d9478_65);
and \U$11307 ( \11402 , \11400 , \11401 );
nor \U$11308 ( \11403 , \11399 , \11402 );
buf \U$11309 ( \11404 , \11403 );
buf \U$11310 ( \11405 , \11404 );
or \U$11311 ( \11406 , \11396 , \11405 );
nand \U$11312 ( \11407 , \11395 , \11406 );
buf \U$11313 ( \11408 , \11407 );
buf \U$11314 ( \11409 , \11408 );
buf \U$11315 ( \11410 , \1417 );
buf \U$11316 ( \11411 , \11318 );
or \U$11317 ( \11412 , \11410 , \11411 );
buf \U$11318 ( \11413 , \6437 );
buf \U$11319 ( \11414 , \11307 );
buf \U$11320 ( \11415 , RIc0d78d0_6);
and \U$11321 ( \11416 , \11414 , \11415 );
buf \U$11322 ( \11417 , \11224 );
buf \U$11323 ( \11418 , RIc0d9568_67);
and \U$11324 ( \11419 , \11417 , \11418 );
nor \U$11325 ( \11420 , \11416 , \11419 );
buf \U$11326 ( \11421 , \11420 );
buf \U$11327 ( \11422 , \11421 );
or \U$11328 ( \11423 , \11413 , \11422 );
nand \U$11329 ( \11424 , \11412 , \11423 );
buf \U$11330 ( \11425 , \11424 );
buf \U$11331 ( \11426 , \11425 );
xor \U$11332 ( \11427 , \11409 , \11426 );
buf \U$11333 ( \11428 , \1279 );
not \U$11334 ( \11429 , \11428 );
buf \U$11335 ( \11430 , \263 );
buf \U$11336 ( \11431 , RIc0d76f0_2);
and \U$11337 ( \11432 , \11430 , \11431 );
buf \U$11338 ( \11433 , \352 );
buf \U$11339 ( \11434 , RIc0d9748_71);
and \U$11340 ( \11435 , \11433 , \11434 );
nor \U$11341 ( \11436 , \11432 , \11435 );
buf \U$11342 ( \11437 , \11436 );
buf \U$11343 ( \11438 , \11437 );
not \U$11344 ( \11439 , \11438 );
and \U$11345 ( \11440 , \11429 , \11439 );
buf \U$11346 ( \11441 , \2269 );
buf \U$11347 ( \11442 , \11280 );
and \U$11348 ( \11443 , \11441 , \11442 );
nor \U$11349 ( \11444 , \11440 , \11443 );
buf \U$11350 ( \11445 , \11444 );
buf \U$11351 ( \11446 , \11445 );
xor \U$11352 ( \11447 , \11427 , \11446 );
buf \U$11353 ( \11448 , \11447 );
buf \U$11354 ( \11449 , \11448 );
xor \U$11355 ( \11450 , \11392 , \11449 );
xor \U$11356 ( \11451 , \11198 , \11215 );
and \U$11357 ( \11452 , \11451 , \11236 );
and \U$11358 ( \11453 , \11198 , \11215 );
or \U$11359 ( \11454 , \11452 , \11453 );
buf \U$11360 ( \11455 , \11454 );
xor \U$11361 ( \11456 , \11300 , \11322 );
xor \U$11362 ( \11457 , \11456 , \11339 );
and \U$11363 ( \11458 , \11455 , \11457 );
xor \U$11364 ( \11459 , \11266 , \11275 );
xor \U$11365 ( \11460 , \11459 , \11291 );
buf \U$11366 ( \11461 , \11460 );
xor \U$11367 ( \11462 , \11300 , \11322 );
xor \U$11368 ( \11463 , \11462 , \11339 );
and \U$11369 ( \11464 , \11461 , \11463 );
and \U$11370 ( \11465 , \11455 , \11461 );
or \U$11371 ( \11466 , \11458 , \11464 , \11465 );
buf \U$11372 ( \11467 , \11466 );
xor \U$11373 ( \11468 , \11450 , \11467 );
buf \U$11374 ( \11469 , \11468 );
buf \U$11375 ( \11470 , \11469 );
xor \U$11376 ( \11471 , \11386 , \11470 );
buf \U$11377 ( \11472 , \11471 );
buf \U$11378 ( \11473 , \11472 );
xor \U$11379 ( \11474 , \11300 , \11322 );
xor \U$11380 ( \11475 , \11474 , \11339 );
xor \U$11381 ( \11476 , \11455 , \11461 );
xor \U$11382 ( \11477 , \11475 , \11476 );
buf \U$11383 ( \11478 , \11477 );
xor \U$11384 ( \11479 , \11133 , \11164 );
xor \U$11385 ( \11480 , \11479 , \11244 );
buf \U$11386 ( \11481 , \11480 );
buf \U$11387 ( \11482 , \11481 );
xor \U$11388 ( \11483 , \11478 , \11482 );
xor \U$11389 ( \11484 , \10975 , \11010 );
and \U$11390 ( \11485 , \11484 , \11017 );
and \U$11391 ( \11486 , \10975 , \11010 );
or \U$11392 ( \11487 , \11485 , \11486 );
buf \U$11393 ( \11488 , \11487 );
buf \U$11394 ( \11489 , \11488 );
xor \U$11395 ( \11490 , \11137 , \11152 );
xor \U$11396 ( \11491 , \11490 , \11159 );
buf \U$11397 ( \11492 , \11491 );
buf \U$11398 ( \11493 , \11492 );
xor \U$11399 ( \11494 , \11489 , \11493 );
xor \U$11400 ( \11495 , \11180 , \11184 );
xor \U$11401 ( \11496 , \11495 , \11239 );
buf \U$11402 ( \11497 , \11496 );
buf \U$11403 ( \11498 , \11497 );
and \U$11404 ( \11499 , \11494 , \11498 );
and \U$11405 ( \11500 , \11489 , \11493 );
or \U$11406 ( \11501 , \11499 , \11500 );
buf \U$11407 ( \11502 , \11501 );
buf \U$11408 ( \11503 , \11502 );
and \U$11409 ( \11504 , \11483 , \11503 );
and \U$11410 ( \11505 , \11478 , \11482 );
or \U$11411 ( \11506 , \11504 , \11505 );
buf \U$11412 ( \11507 , \11506 );
buf \U$11413 ( \11508 , \11507 );
nor \U$11414 ( \11509 , \11473 , \11508 );
buf \U$11415 ( \11510 , \11509 );
buf \U$11416 ( \11511 , \11510 );
not \U$11417 ( \11512 , \11511 );
xor \U$11418 ( \11513 , \10884 , \10932 );
and \U$11419 ( \11514 , \11513 , \10948 );
and \U$11420 ( \11515 , \10884 , \10932 );
or \U$11421 ( \11516 , \11514 , \11515 );
buf \U$11422 ( \11517 , \11516 );
buf \U$11423 ( \11518 , \11517 );
xor \U$11424 ( \11519 , \10957 , \11020 );
and \U$11425 ( \11520 , \11519 , \11039 );
and \U$11426 ( \11521 , \10957 , \11020 );
or \U$11427 ( \11522 , \11520 , \11521 );
buf \U$11428 ( \11523 , \11522 );
buf \U$11429 ( \11524 , \11523 );
xor \U$11430 ( \11525 , \11518 , \11524 );
xor \U$11431 ( \11526 , \11489 , \11493 );
xor \U$11432 ( \11527 , \11526 , \11498 );
buf \U$11433 ( \11528 , \11527 );
buf \U$11434 ( \11529 , \11528 );
xor \U$11435 ( \11530 , \11525 , \11529 );
buf \U$11436 ( \11531 , \11530 );
buf \U$11437 ( \11532 , \11531 );
xor \U$11438 ( \11533 , \10951 , \11042 );
and \U$11439 ( \11534 , \11533 , \11049 );
and \U$11440 ( \11535 , \10951 , \11042 );
or \U$11441 ( \11536 , \11534 , \11535 );
buf \U$11442 ( \11537 , \11536 );
buf \U$11443 ( \11538 , \11537 );
nor \U$11444 ( \11539 , \11532 , \11538 );
buf \U$11445 ( \11540 , \11539 );
buf \U$11446 ( \11541 , \11540 );
xor \U$11447 ( \11542 , \11478 , \11482 );
xor \U$11448 ( \11543 , \11542 , \11503 );
buf \U$11449 ( \11544 , \11543 );
buf \U$11450 ( \11545 , \11544 );
xor \U$11451 ( \11546 , \11518 , \11524 );
and \U$11452 ( \11547 , \11546 , \11529 );
and \U$11453 ( \11548 , \11518 , \11524 );
or \U$11454 ( \11549 , \11547 , \11548 );
buf \U$11455 ( \11550 , \11549 );
buf \U$11456 ( \11551 , \11550 );
nor \U$11457 ( \11552 , \11545 , \11551 );
buf \U$11458 ( \11553 , \11552 );
buf \U$11459 ( \11554 , \11553 );
nor \U$11460 ( \11555 , \11541 , \11554 );
buf \U$11461 ( \11556 , \11555 );
buf \U$11462 ( \11557 , \11556 );
nand \U$11463 ( \11558 , \11512 , \11557 );
buf \U$11464 ( \11559 , \11558 );
buf \U$11465 ( \11560 , \11559 );
xor \U$11466 ( \11561 , \11249 , \11385 );
and \U$11467 ( \11562 , \11561 , \11470 );
and \U$11468 ( \11563 , \11249 , \11385 );
or \U$11469 ( \11564 , \11562 , \11563 );
buf \U$11470 ( \11565 , \11564 );
buf \U$11471 ( \11566 , \11565 );
xor \U$11472 ( \11567 , \11392 , \11449 );
and \U$11473 ( \11568 , \11567 , \11467 );
and \U$11474 ( \11569 , \11392 , \11449 );
or \U$11475 ( \11570 , \11568 , \11569 );
buf \U$11476 ( \11571 , \11570 );
buf \U$11477 ( \11572 , \11571 );
xor \U$11478 ( \11573 , \11296 , \11343 );
and \U$11479 ( \11574 , \11573 , \11382 );
and \U$11480 ( \11575 , \11296 , \11343 );
or \U$11481 ( \11576 , \11574 , \11575 );
buf \U$11482 ( \11577 , \11576 );
buf \U$11483 ( \11578 , \11577 );
xor \U$11484 ( \11579 , \11572 , \11578 );
buf \U$11485 ( \11580 , \1417 );
buf \U$11486 ( \11581 , \11421 );
or \U$11487 ( \11582 , \11580 , \11581 );
buf \U$11488 ( \11583 , \6437 );
buf \U$11489 ( \11584 , \11307 );
buf \U$11490 ( \11585 , RIc0d7858_5);
and \U$11491 ( \11586 , \11584 , \11585 );
buf \U$11492 ( \11587 , \1990 );
buf \U$11493 ( \11588 , RIc0d9568_67);
and \U$11494 ( \11589 , \11587 , \11588 );
nor \U$11495 ( \11590 , \11586 , \11589 );
buf \U$11496 ( \11591 , \11590 );
buf \U$11497 ( \11592 , \11591 );
or \U$11498 ( \11593 , \11583 , \11592 );
nand \U$11499 ( \11594 , \11582 , \11593 );
buf \U$11500 ( \11595 , \11594 );
buf \U$11501 ( \11596 , \5976 );
buf \U$11502 ( \11597 , \7456 );
nor \U$11503 ( \11598 , \11596 , \11597 );
buf \U$11504 ( \11599 , \11598 );
xor \U$11505 ( \11600 , \11595 , \11599 );
buf \U$11506 ( \11601 , \7449 );
buf \U$11507 ( \11602 , \11404 );
or \U$11508 ( \11603 , \11601 , \11602 );
buf \U$11509 ( \11604 , \1232 );
buf \U$11510 ( \11605 , \7456 );
buf \U$11511 ( \11606 , RIc0d7948_7);
and \U$11512 ( \11607 , \11605 , \11606 );
buf \U$11513 ( \11608 , \11313 );
buf \U$11514 ( \11609 , RIc0d9478_65);
and \U$11515 ( \11610 , \11608 , \11609 );
nor \U$11516 ( \11611 , \11607 , \11610 );
buf \U$11517 ( \11612 , \11611 );
buf \U$11518 ( \11613 , \11612 );
or \U$11519 ( \11614 , \11604 , \11613 );
nand \U$11520 ( \11615 , \11603 , \11614 );
buf \U$11521 ( \11616 , \11615 );
xor \U$11522 ( \11617 , \11600 , \11616 );
xor \U$11523 ( \11618 , \11409 , \11426 );
and \U$11524 ( \11619 , \11618 , \11446 );
and \U$11525 ( \11620 , \11409 , \11426 );
or \U$11526 ( \11621 , \11619 , \11620 );
buf \U$11527 ( \11622 , \11621 );
xor \U$11528 ( \11623 , \11356 , \11361 );
and \U$11529 ( \11624 , \11623 , \11379 );
and \U$11530 ( \11625 , \11356 , \11361 );
or \U$11531 ( \11626 , \11624 , \11625 );
buf \U$11532 ( \11627 , \11626 );
buf \U$11533 ( \11628 , \11627 );
buf \U$11534 ( \11629 , \11445 );
not \U$11535 ( \11630 , \11629 );
buf \U$11536 ( \11631 , \11630 );
buf \U$11537 ( \11632 , \11631 );
xor \U$11538 ( \11633 , \11628 , \11632 );
buf \U$11539 ( \11634 , \4868 );
buf \U$11540 ( \11635 , \11437 );
or \U$11541 ( \11636 , \11634 , \11635 );
buf \U$11542 ( \11637 , \1279 );
buf \U$11543 ( \11638 , \263 );
buf \U$11544 ( \11639 , RIc0d7678_1);
and \U$11545 ( \11640 , \11638 , \11639 );
buf \U$11546 ( \11641 , \974 );
buf \U$11547 ( \11642 , RIc0d9748_71);
and \U$11548 ( \11643 , \11641 , \11642 );
nor \U$11549 ( \11644 , \11640 , \11643 );
buf \U$11550 ( \11645 , \11644 );
buf \U$11551 ( \11646 , \11645 );
or \U$11552 ( \11647 , \11637 , \11646 );
nand \U$11553 ( \11648 , \11636 , \11647 );
buf \U$11554 ( \11649 , \11648 );
buf \U$11555 ( \11650 , \11649 );
buf \U$11556 ( \11651 , \2871 );
buf \U$11557 ( \11652 , \2882 );
or \U$11558 ( \11653 , \11651 , \11652 );
buf \U$11559 ( \11654 , RIc0d9838_73);
nand \U$11560 ( \11655 , \11653 , \11654 );
buf \U$11561 ( \11656 , \11655 );
buf \U$11562 ( \11657 , \11656 );
xor \U$11563 ( \11658 , \11650 , \11657 );
buf \U$11564 ( \11659 , \1452 );
buf \U$11565 ( \11660 , \11374 );
or \U$11566 ( \11661 , \11659 , \11660 );
buf \U$11567 ( \11662 , \1969 );
buf \U$11568 ( \11663 , RIc0d9658_69);
buf \U$11569 ( \11664 , \304 );
and \U$11570 ( \11665 , \11663 , \11664 );
not \U$11571 ( \11666 , \11663 );
buf \U$11572 ( \11667 , RIc0d7768_3);
and \U$11573 ( \11668 , \11666 , \11667 );
nor \U$11574 ( \11669 , \11665 , \11668 );
buf \U$11575 ( \11670 , \11669 );
buf \U$11576 ( \11671 , \11670 );
or \U$11577 ( \11672 , \11662 , \11671 );
nand \U$11578 ( \11673 , \11661 , \11672 );
buf \U$11579 ( \11674 , \11673 );
buf \U$11580 ( \11675 , \11674 );
xor \U$11581 ( \11676 , \11658 , \11675 );
buf \U$11582 ( \11677 , \11676 );
buf \U$11583 ( \11678 , \11677 );
xor \U$11584 ( \11679 , \11633 , \11678 );
buf \U$11585 ( \11680 , \11679 );
xor \U$11586 ( \11681 , \11622 , \11680 );
xor \U$11587 ( \11682 , \11617 , \11681 );
buf \U$11588 ( \11683 , \11682 );
xor \U$11589 ( \11684 , \11579 , \11683 );
buf \U$11590 ( \11685 , \11684 );
buf \U$11591 ( \11686 , \11685 );
nor \U$11592 ( \11687 , \11566 , \11686 );
buf \U$11593 ( \11688 , \11687 );
buf \U$11594 ( \11689 , \11688 );
nor \U$11595 ( \11690 , \11560 , \11689 );
buf \U$11596 ( \11691 , \11690 );
buf \U$11597 ( \11692 , \11691 );
nand \U$11598 ( \11693 , \11058 , \11692 );
buf \U$11599 ( \11694 , \11693 );
buf \U$11600 ( \11695 , \11694 );
not \U$11601 ( \11696 , \11695 );
buf \U$11602 ( \11697 , \11696 );
buf \U$11603 ( \11698 , \11697 );
and \U$11604 ( \11699 , \10112 , \11698 );
buf \U$11605 ( \11700 , \11699 );
buf \U$11606 ( \11701 , \11700 );
buf \U$11607 ( \11702 , \1417 );
buf \U$11608 ( \11703 , \11307 );
buf \U$11609 ( \11704 , RIc0d76f0_2);
and \U$11610 ( \11705 , \11703 , \11704 );
buf \U$11611 ( \11706 , \352 );
buf \U$11612 ( \11707 , RIc0d9568_67);
and \U$11613 ( \11708 , \11706 , \11707 );
nor \U$11614 ( \11709 , \11705 , \11708 );
buf \U$11615 ( \11710 , \11709 );
buf \U$11616 ( \11711 , \11710 );
or \U$11617 ( \11712 , \11702 , \11711 );
buf \U$11618 ( \11713 , \6437 );
buf \U$11619 ( \11714 , \11307 );
buf \U$11620 ( \11715 , RIc0d7678_1);
and \U$11621 ( \11716 , \11714 , \11715 );
buf \U$11622 ( \11717 , \974 );
buf \U$11623 ( \11718 , RIc0d9568_67);
and \U$11624 ( \11719 , \11717 , \11718 );
nor \U$11625 ( \11720 , \11716 , \11719 );
buf \U$11626 ( \11721 , \11720 );
buf \U$11627 ( \11722 , \11721 );
or \U$11628 ( \11723 , \11713 , \11722 );
nand \U$11629 ( \11724 , \11712 , \11723 );
buf \U$11630 ( \11725 , \11724 );
buf \U$11631 ( \11726 , \11725 );
buf \U$11632 ( \11727 , \7456 );
buf \U$11633 ( \11728 , \1990 );
nor \U$11634 ( \11729 , \11727 , \11728 );
buf \U$11635 ( \11730 , \11729 );
buf \U$11636 ( \11731 , \11730 );
xor \U$11637 ( \11732 , \11726 , \11731 );
buf \U$11638 ( \11733 , \7449 );
buf \U$11639 ( \11734 , \7456 );
buf \U$11640 ( \11735 , RIc0d77e0_4);
and \U$11641 ( \11736 , \11734 , \11735 );
buf \U$11642 ( \11737 , \489 );
buf \U$11643 ( \11738 , RIc0d9478_65);
and \U$11644 ( \11739 , \11737 , \11738 );
nor \U$11645 ( \11740 , \11736 , \11739 );
buf \U$11646 ( \11741 , \11740 );
buf \U$11647 ( \11742 , \11741 );
or \U$11648 ( \11743 , \11733 , \11742 );
buf \U$11649 ( \11744 , \1232 );
buf \U$11650 ( \11745 , \7456 );
buf \U$11651 ( \11746 , RIc0d7768_3);
and \U$11652 ( \11747 , \11745 , \11746 );
buf \U$11653 ( \11748 , \304 );
buf \U$11654 ( \11749 , RIc0d9478_65);
and \U$11655 ( \11750 , \11748 , \11749 );
nor \U$11656 ( \11751 , \11747 , \11750 );
buf \U$11657 ( \11752 , \11751 );
buf \U$11658 ( \11753 , \11752 );
or \U$11659 ( \11754 , \11744 , \11753 );
nand \U$11660 ( \11755 , \11743 , \11754 );
buf \U$11661 ( \11756 , \11755 );
buf \U$11662 ( \11757 , \11756 );
xor \U$11663 ( \11758 , \11732 , \11757 );
buf \U$11664 ( \11759 , \11758 );
buf \U$11665 ( \11760 , \1452 );
not \U$11666 ( \11761 , \11760 );
buf \U$11667 ( \11762 , RIc0d9658_69);
buf \U$11668 ( \11763 , \974 );
and \U$11669 ( \11764 , \11762 , \11763 );
not \U$11670 ( \11765 , \11762 );
buf \U$11671 ( \11766 , RIc0d7678_1);
and \U$11672 ( \11767 , \11765 , \11766 );
nor \U$11673 ( \11768 , \11764 , \11767 );
buf \U$11674 ( \11769 , \11768 );
buf \U$11675 ( \11770 , \11769 );
not \U$11676 ( \11771 , \11770 );
and \U$11677 ( \11772 , \11761 , \11771 );
buf \U$11678 ( \11773 , \874 );
buf \U$11679 ( \11774 , RIc0d9658_69);
and \U$11680 ( \11775 , \11773 , \11774 );
nor \U$11681 ( \11776 , \11772 , \11775 );
buf \U$11682 ( \11777 , \11776 );
buf \U$11683 ( \11778 , \11777 );
not \U$11684 ( \11779 , \11778 );
buf \U$11685 ( \11780 , \11779 );
buf \U$11686 ( \11781 , \279 );
buf \U$11687 ( \11782 , \874 );
or \U$11688 ( \11783 , \11781 , \11782 );
buf \U$11689 ( \11784 , RIc0d9658_69);
nand \U$11690 ( \11785 , \11783 , \11784 );
buf \U$11691 ( \11786 , \11785 );
xor \U$11692 ( \11787 , \11780 , \11786 );
buf \U$11693 ( \11788 , \1417 );
buf \U$11694 ( \11789 , \11307 );
buf \U$11695 ( \11790 , RIc0d7768_3);
and \U$11696 ( \11791 , \11789 , \11790 );
buf \U$11697 ( \11792 , \304 );
buf \U$11698 ( \11793 , RIc0d9568_67);
and \U$11699 ( \11794 , \11792 , \11793 );
nor \U$11700 ( \11795 , \11791 , \11794 );
buf \U$11701 ( \11796 , \11795 );
buf \U$11702 ( \11797 , \11796 );
or \U$11703 ( \11798 , \11788 , \11797 );
buf \U$11704 ( \11799 , \6437 );
buf \U$11705 ( \11800 , \11710 );
or \U$11706 ( \11801 , \11799 , \11800 );
nand \U$11707 ( \11802 , \11798 , \11801 );
buf \U$11708 ( \11803 , \11802 );
buf \U$11709 ( \11804 , \11803 );
buf \U$11710 ( \11805 , \11224 );
buf \U$11711 ( \11806 , \7456 );
nor \U$11712 ( \11807 , \11805 , \11806 );
buf \U$11713 ( \11808 , \11807 );
buf \U$11714 ( \11809 , \11808 );
xor \U$11715 ( \11810 , \11804 , \11809 );
buf \U$11716 ( \11811 , \7449 );
buf \U$11717 ( \11812 , \7456 );
buf \U$11718 ( \11813 , RIc0d7858_5);
and \U$11719 ( \11814 , \11812 , \11813 );
buf \U$11720 ( \11815 , \1990 );
buf \U$11721 ( \11816 , RIc0d9478_65);
and \U$11722 ( \11817 , \11815 , \11816 );
nor \U$11723 ( \11818 , \11814 , \11817 );
buf \U$11724 ( \11819 , \11818 );
buf \U$11725 ( \11820 , \11819 );
or \U$11726 ( \11821 , \11811 , \11820 );
buf \U$11727 ( \11822 , \1232 );
buf \U$11728 ( \11823 , \11741 );
or \U$11729 ( \11824 , \11822 , \11823 );
nand \U$11730 ( \11825 , \11821 , \11824 );
buf \U$11731 ( \11826 , \11825 );
buf \U$11732 ( \11827 , \11826 );
and \U$11733 ( \11828 , \11810 , \11827 );
and \U$11734 ( \11829 , \11804 , \11809 );
or \U$11735 ( \11830 , \11828 , \11829 );
buf \U$11736 ( \11831 , \11830 );
xor \U$11737 ( \11832 , \11787 , \11831 );
and \U$11738 ( \11833 , \11759 , \11832 );
buf \U$11739 ( \11834 , \1417 );
buf \U$11740 ( \11835 , \11307 );
buf \U$11741 ( \11836 , RIc0d77e0_4);
and \U$11742 ( \11837 , \11835 , \11836 );
buf \U$11743 ( \11838 , \489 );
buf \U$11744 ( \11839 , RIc0d9568_67);
and \U$11745 ( \11840 , \11838 , \11839 );
nor \U$11746 ( \11841 , \11837 , \11840 );
buf \U$11747 ( \11842 , \11841 );
buf \U$11748 ( \11843 , \11842 );
or \U$11749 ( \11844 , \11834 , \11843 );
buf \U$11750 ( \11845 , \6437 );
buf \U$11751 ( \11846 , \11796 );
or \U$11752 ( \11847 , \11845 , \11846 );
nand \U$11753 ( \11848 , \11844 , \11847 );
buf \U$11754 ( \11849 , \11848 );
buf \U$11755 ( \11850 , \11849 );
buf \U$11756 ( \11851 , \11313 );
buf \U$11757 ( \11852 , \7456 );
nor \U$11758 ( \11853 , \11851 , \11852 );
buf \U$11759 ( \11854 , \11853 );
buf \U$11760 ( \11855 , \11854 );
xor \U$11761 ( \11856 , \11850 , \11855 );
buf \U$11762 ( \11857 , \7449 );
buf \U$11763 ( \11858 , \7456 );
buf \U$11764 ( \11859 , RIc0d78d0_6);
and \U$11765 ( \11860 , \11858 , \11859 );
buf \U$11766 ( \11861 , \11224 );
buf \U$11767 ( \11862 , RIc0d9478_65);
and \U$11768 ( \11863 , \11861 , \11862 );
nor \U$11769 ( \11864 , \11860 , \11863 );
buf \U$11770 ( \11865 , \11864 );
buf \U$11771 ( \11866 , \11865 );
or \U$11772 ( \11867 , \11857 , \11866 );
buf \U$11773 ( \11868 , \1232 );
buf \U$11774 ( \11869 , \11819 );
or \U$11775 ( \11870 , \11868 , \11869 );
nand \U$11776 ( \11871 , \11867 , \11870 );
buf \U$11777 ( \11872 , \11871 );
buf \U$11778 ( \11873 , \11872 );
and \U$11779 ( \11874 , \11856 , \11873 );
and \U$11780 ( \11875 , \11850 , \11855 );
or \U$11781 ( \11876 , \11874 , \11875 );
buf \U$11782 ( \11877 , \11876 );
xor \U$11783 ( \11878 , \11877 , \11777 );
xor \U$11784 ( \11879 , \11804 , \11809 );
xor \U$11785 ( \11880 , \11879 , \11827 );
buf \U$11786 ( \11881 , \11880 );
and \U$11787 ( \11882 , \11878 , \11881 );
and \U$11788 ( \11883 , \11877 , \11777 );
or \U$11789 ( \11884 , \11882 , \11883 );
xor \U$11790 ( \11885 , \11780 , \11786 );
xor \U$11791 ( \11886 , \11885 , \11831 );
and \U$11792 ( \11887 , \11884 , \11886 );
and \U$11793 ( \11888 , \11759 , \11884 );
or \U$11794 ( \11889 , \11833 , \11887 , \11888 );
buf \U$11795 ( \11890 , \11889 );
buf \U$11796 ( \11891 , \7449 );
buf \U$11797 ( \11892 , \11752 );
or \U$11798 ( \11893 , \11891 , \11892 );
buf \U$11799 ( \11894 , \1232 );
buf \U$11800 ( \11895 , \7456 );
buf \U$11801 ( \11896 , RIc0d76f0_2);
and \U$11802 ( \11897 , \11895 , \11896 );
buf \U$11803 ( \11898 , \352 );
buf \U$11804 ( \11899 , RIc0d9478_65);
and \U$11805 ( \11900 , \11898 , \11899 );
nor \U$11806 ( \11901 , \11897 , \11900 );
buf \U$11807 ( \11902 , \11901 );
buf \U$11808 ( \11903 , \11902 );
or \U$11809 ( \11904 , \11894 , \11903 );
nand \U$11810 ( \11905 , \11893 , \11904 );
buf \U$11811 ( \11906 , \11905 );
buf \U$11812 ( \11907 , RIc0d77e0_4);
buf \U$11813 ( \11908 , RIc0d9478_65);
nand \U$11814 ( \11909 , \11907 , \11908 );
buf \U$11815 ( \11910 , \11909 );
xor \U$11816 ( \11911 , \11906 , \11910 );
buf \U$11817 ( \11912 , \1417 );
buf \U$11818 ( \11913 , \11721 );
or \U$11819 ( \11914 , \11912 , \11913 );
buf \U$11820 ( \11915 , \6437 );
buf \U$11821 ( \11916 , \11307 );
or \U$11822 ( \11917 , \11915 , \11916 );
nand \U$11823 ( \11918 , \11914 , \11917 );
buf \U$11824 ( \11919 , \11918 );
xor \U$11825 ( \11920 , \11911 , \11919 );
xor \U$11826 ( \11921 , \11726 , \11731 );
and \U$11827 ( \11922 , \11921 , \11757 );
and \U$11828 ( \11923 , \11726 , \11731 );
or \U$11829 ( \11924 , \11922 , \11923 );
buf \U$11830 ( \11925 , \11924 );
xor \U$11831 ( \11926 , \11780 , \11786 );
and \U$11832 ( \11927 , \11926 , \11831 );
and \U$11833 ( \11928 , \11780 , \11786 );
or \U$11834 ( \11929 , \11927 , \11928 );
xor \U$11835 ( \11930 , \11925 , \11929 );
xor \U$11836 ( \11931 , \11920 , \11930 );
buf \U$11837 ( \11932 , \11931 );
nor \U$11838 ( \11933 , \11890 , \11932 );
buf \U$11839 ( \11934 , \11933 );
buf \U$11840 ( \11935 , \11934 );
xor \U$11841 ( \11936 , \11906 , \11910 );
xor \U$11842 ( \11937 , \11936 , \11919 );
and \U$11843 ( \11938 , \11925 , \11937 );
xor \U$11844 ( \11939 , \11906 , \11910 );
xor \U$11845 ( \11940 , \11939 , \11919 );
and \U$11846 ( \11941 , \11929 , \11940 );
and \U$11847 ( \11942 , \11925 , \11929 );
or \U$11848 ( \11943 , \11938 , \11941 , \11942 );
buf \U$11849 ( \11944 , \11943 );
xor \U$11850 ( \11945 , \11906 , \11910 );
and \U$11851 ( \11946 , \11945 , \11919 );
and \U$11852 ( \11947 , \11906 , \11910 );
or \U$11853 ( \11948 , \11946 , \11947 );
buf \U$11854 ( \11949 , \11948 );
buf \U$11855 ( \11950 , \11910 );
not \U$11856 ( \11951 , \11950 );
buf \U$11857 ( \11952 , \11951 );
buf \U$11858 ( \11953 , \11952 );
xor \U$11859 ( \11954 , \11949 , \11953 );
buf \U$11860 ( \11955 , \10034 );
buf \U$11861 ( \11956 , \686 );
or \U$11862 ( \11957 , \11955 , \11956 );
buf \U$11863 ( \11958 , RIc0d9568_67);
nand \U$11864 ( \11959 , \11957 , \11958 );
buf \U$11865 ( \11960 , \11959 );
buf \U$11866 ( \11961 , \11960 );
buf \U$11867 ( \11962 , \7456 );
buf \U$11868 ( \11963 , \304 );
nor \U$11869 ( \11964 , \11962 , \11963 );
buf \U$11870 ( \11965 , \11964 );
buf \U$11871 ( \11966 , \11965 );
xor \U$11872 ( \11967 , \11961 , \11966 );
buf \U$11873 ( \11968 , \7449 );
buf \U$11874 ( \11969 , \11902 );
or \U$11875 ( \11970 , \11968 , \11969 );
buf \U$11876 ( \11971 , \1232 );
buf \U$11877 ( \11972 , \7456 );
buf \U$11878 ( \11973 , RIc0d7678_1);
and \U$11879 ( \11974 , \11972 , \11973 );
buf \U$11880 ( \11975 , \974 );
buf \U$11881 ( \11976 , RIc0d9478_65);
and \U$11882 ( \11977 , \11975 , \11976 );
nor \U$11883 ( \11978 , \11974 , \11977 );
buf \U$11884 ( \11979 , \11978 );
buf \U$11885 ( \11980 , \11979 );
or \U$11886 ( \11981 , \11971 , \11980 );
nand \U$11887 ( \11982 , \11970 , \11981 );
buf \U$11888 ( \11983 , \11982 );
buf \U$11889 ( \11984 , \11983 );
xor \U$11890 ( \11985 , \11967 , \11984 );
buf \U$11891 ( \11986 , \11985 );
buf \U$11892 ( \11987 , \11986 );
xor \U$11893 ( \11988 , \11954 , \11987 );
buf \U$11894 ( \11989 , \11988 );
buf \U$11895 ( \11990 , \11989 );
nor \U$11896 ( \11991 , \11944 , \11990 );
buf \U$11897 ( \11992 , \11991 );
buf \U$11898 ( \11993 , \11992 );
nor \U$11899 ( \11994 , \11935 , \11993 );
buf \U$11900 ( \11995 , \11994 );
buf \U$11901 ( \11996 , \11995 );
not \U$11902 ( \11997 , \11996 );
buf \U$11903 ( \11998 , \1417 );
buf \U$11904 ( \11999 , \11591 );
or \U$11905 ( \12000 , \11998 , \11999 );
buf \U$11906 ( \12001 , \6437 );
buf \U$11907 ( \12002 , \11842 );
or \U$11908 ( \12003 , \12001 , \12002 );
nand \U$11909 ( \12004 , \12000 , \12003 );
buf \U$11910 ( \12005 , \12004 );
buf \U$11911 ( \12006 , \12005 );
buf \U$11912 ( \12007 , \7449 );
buf \U$11913 ( \12008 , \11612 );
or \U$11914 ( \12009 , \12007 , \12008 );
buf \U$11915 ( \12010 , \1232 );
buf \U$11916 ( \12011 , \11865 );
or \U$11917 ( \12012 , \12010 , \12011 );
nand \U$11918 ( \12013 , \12009 , \12012 );
buf \U$11919 ( \12014 , \12013 );
buf \U$11920 ( \12015 , \12014 );
xor \U$11921 ( \12016 , \12006 , \12015 );
buf \U$11922 ( \12017 , \1452 );
buf \U$11923 ( \12018 , \11670 );
or \U$11924 ( \12019 , \12017 , \12018 );
buf \U$11925 ( \12020 , \1969 );
buf \U$11926 ( \12021 , RIc0d9658_69);
buf \U$11927 ( \12022 , \352 );
and \U$11928 ( \12023 , \12021 , \12022 );
not \U$11929 ( \12024 , \12021 );
buf \U$11930 ( \12025 , RIc0d76f0_2);
and \U$11931 ( \12026 , \12024 , \12025 );
nor \U$11932 ( \12027 , \12023 , \12026 );
buf \U$11933 ( \12028 , \12027 );
buf \U$11934 ( \12029 , \12028 );
or \U$11935 ( \12030 , \12020 , \12029 );
nand \U$11936 ( \12031 , \12019 , \12030 );
buf \U$11937 ( \12032 , \12031 );
buf \U$11938 ( \12033 , \12032 );
xor \U$11939 ( \12034 , \12016 , \12033 );
buf \U$11940 ( \12035 , \12034 );
xor \U$11941 ( \12036 , \11595 , \11599 );
and \U$11942 ( \12037 , \12036 , \11616 );
and \U$11943 ( \12038 , \11595 , \11599 );
or \U$11944 ( \12039 , \12037 , \12038 );
xor \U$11945 ( \12040 , \12035 , \12039 );
buf \U$11946 ( \12041 , \4868 );
buf \U$11947 ( \12042 , \11645 );
or \U$11948 ( \12043 , \12041 , \12042 );
buf \U$11949 ( \12044 , \1279 );
buf \U$11950 ( \12045 , \263 );
or \U$11951 ( \12046 , \12044 , \12045 );
nand \U$11952 ( \12047 , \12043 , \12046 );
buf \U$11953 ( \12048 , \12047 );
buf \U$11954 ( \12049 , \12048 );
not \U$11955 ( \12050 , \12049 );
buf \U$11956 ( \12051 , \12050 );
buf \U$11957 ( \12052 , \12051 );
buf \U$11958 ( \12053 , \4448 );
buf \U$11959 ( \12054 , \7456 );
nor \U$11960 ( \12055 , \12053 , \12054 );
buf \U$11961 ( \12056 , \12055 );
buf \U$11962 ( \12057 , \12056 );
xor \U$11963 ( \12058 , \12052 , \12057 );
xor \U$11964 ( \12059 , \11650 , \11657 );
and \U$11965 ( \12060 , \12059 , \11675 );
and \U$11966 ( \12061 , \11650 , \11657 );
or \U$11967 ( \12062 , \12060 , \12061 );
buf \U$11968 ( \12063 , \12062 );
buf \U$11969 ( \12064 , \12063 );
xor \U$11970 ( \12065 , \12058 , \12064 );
buf \U$11971 ( \12066 , \12065 );
xor \U$11972 ( \12067 , \12040 , \12066 );
xor \U$11973 ( \12068 , \11628 , \11632 );
and \U$11974 ( \12069 , \12068 , \11678 );
and \U$11975 ( \12070 , \11628 , \11632 );
or \U$11976 ( \12071 , \12069 , \12070 );
buf \U$11977 ( \12072 , \12071 );
xor \U$11978 ( \12073 , \11595 , \11599 );
xor \U$11979 ( \12074 , \12073 , \11616 );
and \U$11980 ( \12075 , \11622 , \12074 );
xor \U$11981 ( \12076 , \11595 , \11599 );
xor \U$11982 ( \12077 , \12076 , \11616 );
and \U$11983 ( \12078 , \11680 , \12077 );
and \U$11984 ( \12079 , \11622 , \11680 );
or \U$11985 ( \12080 , \12075 , \12078 , \12079 );
xor \U$11986 ( \12081 , \12072 , \12080 );
xor \U$11987 ( \12082 , \12067 , \12081 );
buf \U$11988 ( \12083 , \12082 );
xor \U$11989 ( \12084 , \11572 , \11578 );
and \U$11990 ( \12085 , \12084 , \11683 );
and \U$11991 ( \12086 , \11572 , \11578 );
or \U$11992 ( \12087 , \12085 , \12086 );
buf \U$11993 ( \12088 , \12087 );
buf \U$11994 ( \12089 , \12088 );
or \U$11995 ( \12090 , \12083 , \12089 );
buf \U$11996 ( \12091 , \12090 );
buf \U$11997 ( \12092 , \12091 );
not \U$11998 ( \12093 , \12092 );
xor \U$11999 ( \12094 , \11850 , \11855 );
xor \U$12000 ( \12095 , \12094 , \11873 );
buf \U$12001 ( \12096 , \12095 );
xor \U$12002 ( \12097 , \12006 , \12015 );
and \U$12003 ( \12098 , \12097 , \12033 );
and \U$12004 ( \12099 , \12006 , \12015 );
or \U$12005 ( \12100 , \12098 , \12099 );
buf \U$12006 ( \12101 , \12100 );
xor \U$12007 ( \12102 , \12096 , \12101 );
buf \U$12008 ( \12103 , \12048 );
buf \U$12009 ( \12104 , \1279 );
not \U$12010 ( \12105 , \12104 );
buf \U$12011 ( \12106 , \4868 );
not \U$12012 ( \12107 , \12106 );
or \U$12013 ( \12108 , \12105 , \12107 );
buf \U$12014 ( \12109 , RIc0d9748_71);
nand \U$12015 ( \12110 , \12108 , \12109 );
buf \U$12016 ( \12111 , \12110 );
buf \U$12017 ( \12112 , \12111 );
xor \U$12018 ( \12113 , \12103 , \12112 );
buf \U$12019 ( \12114 , \1452 );
buf \U$12020 ( \12115 , \12028 );
or \U$12021 ( \12116 , \12114 , \12115 );
buf \U$12022 ( \12117 , \1969 );
buf \U$12023 ( \12118 , \11769 );
or \U$12024 ( \12119 , \12117 , \12118 );
nand \U$12025 ( \12120 , \12116 , \12119 );
buf \U$12026 ( \12121 , \12120 );
buf \U$12027 ( \12122 , \12121 );
xor \U$12028 ( \12123 , \12113 , \12122 );
buf \U$12029 ( \12124 , \12123 );
xor \U$12030 ( \12125 , \12102 , \12124 );
xor \U$12031 ( \12126 , \12052 , \12057 );
and \U$12032 ( \12127 , \12126 , \12064 );
and \U$12033 ( \12128 , \12052 , \12057 );
or \U$12034 ( \12129 , \12127 , \12128 );
buf \U$12035 ( \12130 , \12129 );
xor \U$12036 ( \12131 , \12035 , \12039 );
and \U$12037 ( \12132 , \12131 , \12066 );
and \U$12038 ( \12133 , \12035 , \12039 );
or \U$12039 ( \12134 , \12132 , \12133 );
xor \U$12040 ( \12135 , \12130 , \12134 );
xor \U$12041 ( \12136 , \12125 , \12135 );
buf \U$12042 ( \12137 , \12136 );
xor \U$12043 ( \12138 , \12035 , \12039 );
xor \U$12044 ( \12139 , \12138 , \12066 );
and \U$12045 ( \12140 , \12072 , \12139 );
xor \U$12046 ( \12141 , \12035 , \12039 );
xor \U$12047 ( \12142 , \12141 , \12066 );
and \U$12048 ( \12143 , \12080 , \12142 );
and \U$12049 ( \12144 , \12072 , \12080 );
or \U$12050 ( \12145 , \12140 , \12143 , \12144 );
buf \U$12051 ( \12146 , \12145 );
nor \U$12052 ( \12147 , \12137 , \12146 );
buf \U$12053 ( \12148 , \12147 );
buf \U$12054 ( \12149 , \12148 );
nor \U$12055 ( \12150 , \12093 , \12149 );
buf \U$12056 ( \12151 , \12150 );
buf \U$12057 ( \12152 , \12151 );
xor \U$12058 ( \12153 , \11877 , \11777 );
xor \U$12059 ( \12154 , \12153 , \11881 );
xor \U$12060 ( \12155 , \12103 , \12112 );
and \U$12061 ( \12156 , \12155 , \12122 );
and \U$12062 ( \12157 , \12103 , \12112 );
or \U$12063 ( \12158 , \12156 , \12157 );
buf \U$12064 ( \12159 , \12158 );
xor \U$12065 ( \12160 , \12096 , \12101 );
and \U$12066 ( \12161 , \12160 , \12124 );
and \U$12067 ( \12162 , \12096 , \12101 );
or \U$12068 ( \12163 , \12161 , \12162 );
xor \U$12069 ( \12164 , \12159 , \12163 );
xor \U$12070 ( \12165 , \12154 , \12164 );
buf \U$12071 ( \12166 , \12165 );
xor \U$12072 ( \12167 , \12096 , \12101 );
xor \U$12073 ( \12168 , \12167 , \12124 );
and \U$12074 ( \12169 , \12130 , \12168 );
xor \U$12075 ( \12170 , \12096 , \12101 );
xor \U$12076 ( \12171 , \12170 , \12124 );
and \U$12077 ( \12172 , \12134 , \12171 );
and \U$12078 ( \12173 , \12130 , \12134 );
or \U$12079 ( \12174 , \12169 , \12172 , \12173 );
buf \U$12080 ( \12175 , \12174 );
or \U$12081 ( \12176 , \12166 , \12175 );
buf \U$12082 ( \12177 , \12176 );
buf \U$12083 ( \12178 , \12177 );
nand \U$12084 ( \12179 , \12152 , \12178 );
buf \U$12085 ( \12180 , \12179 );
buf \U$12086 ( \12181 , \12180 );
xor \U$12087 ( \12182 , \11877 , \11777 );
xor \U$12088 ( \12183 , \12182 , \11881 );
and \U$12089 ( \12184 , \12159 , \12183 );
xor \U$12090 ( \12185 , \11877 , \11777 );
xor \U$12091 ( \12186 , \12185 , \11881 );
and \U$12092 ( \12187 , \12163 , \12186 );
and \U$12093 ( \12188 , \12159 , \12163 );
or \U$12094 ( \12189 , \12184 , \12187 , \12188 );
buf \U$12095 ( \12190 , \12189 );
xor \U$12096 ( \12191 , \11780 , \11786 );
xor \U$12097 ( \12192 , \12191 , \11831 );
xor \U$12098 ( \12193 , \11759 , \11884 );
xor \U$12099 ( \12194 , \12192 , \12193 );
buf \U$12100 ( \12195 , \12194 );
nor \U$12101 ( \12196 , \12190 , \12195 );
buf \U$12102 ( \12197 , \12196 );
buf \U$12103 ( \12198 , \12197 );
nor \U$12104 ( \12199 , \12181 , \12198 );
buf \U$12105 ( \12200 , \12199 );
not \U$12106 ( \12201 , \12200 );
buf \U$12107 ( \12202 , \12201 );
xor \U$12108 ( \12203 , \11949 , \11953 );
and \U$12109 ( \12204 , \12203 , \11987 );
and \U$12110 ( \12205 , \11949 , \11953 );
or \U$12111 ( \12206 , \12204 , \12205 );
buf \U$12112 ( \12207 , \12206 );
buf \U$12113 ( \12208 , \12207 );
buf \U$12114 ( \12209 , \7449 );
buf \U$12115 ( \12210 , \11979 );
or \U$12116 ( \12211 , \12209 , \12210 );
buf \U$12117 ( \12212 , \1235 );
buf \U$12118 ( \12213 , RIc0d9478_65);
nand \U$12119 ( \12214 , \12212 , \12213 );
buf \U$12120 ( \12215 , \12214 );
buf \U$12121 ( \12216 , \12215 );
nand \U$12122 ( \12217 , \12211 , \12216 );
buf \U$12123 ( \12218 , \12217 );
buf \U$12124 ( \12219 , \12218 );
buf \U$12125 ( \12220 , RIc0d76f0_2);
buf \U$12126 ( \12221 , RIc0d9478_65);
nand \U$12127 ( \12222 , \12220 , \12221 );
buf \U$12128 ( \12223 , \12222 );
buf \U$12129 ( \12224 , \12223 );
xor \U$12130 ( \12225 , \12219 , \12224 );
xor \U$12131 ( \12226 , \11961 , \11966 );
and \U$12132 ( \12227 , \12226 , \11984 );
and \U$12133 ( \12228 , \11961 , \11966 );
or \U$12134 ( \12229 , \12227 , \12228 );
buf \U$12135 ( \12230 , \12229 );
buf \U$12136 ( \12231 , \12230 );
xor \U$12137 ( \12232 , \12225 , \12231 );
buf \U$12138 ( \12233 , \12232 );
buf \U$12139 ( \12234 , \12233 );
nor \U$12140 ( \12235 , \12208 , \12234 );
buf \U$12141 ( \12236 , \12235 );
buf \U$12142 ( \12237 , \12236 );
nor \U$12143 ( \12238 , \11997 , \12202 , \12237 );
buf \U$12144 ( \12239 , \12238 );
buf \U$12145 ( \12240 , \12239 );
and \U$12146 ( \12241 , \11701 , \12240 );
buf \U$12147 ( \12242 , \12241 );
buf \U$12148 ( \12243 , \12242 );
not \U$12149 ( \12244 , \12243 );
xor \U$12150 ( \12245 , RIc0d9ce8_83, RIc0d8b90_46);
buf \U$12151 ( \12246 , \12245 );
not \U$12152 ( \12247 , \12246 );
buf \U$12153 ( \12248 , \561 );
buf \U$12154 ( \12249 , \566 );
nand \U$12155 ( \12250 , \12248 , \12249 );
buf \U$12156 ( \12251 , \12250 );
buf \U$12157 ( \12252 , \12251 );
not \U$12158 ( \12253 , \12252 );
buf \U$12159 ( \12254 , \12253 );
buf \U$12160 ( \12255 , \12254 );
not \U$12161 ( \12256 , \12255 );
or \U$12162 ( \12257 , \12247 , \12256 );
buf \U$12163 ( \12258 , \993 );
xor \U$12164 ( \12259 , RIc0d9ce8_83, RIc0d8b18_45);
buf \U$12165 ( \12260 , \12259 );
nand \U$12166 ( \12261 , \12258 , \12260 );
buf \U$12167 ( \12262 , \12261 );
buf \U$12168 ( \12263 , \12262 );
nand \U$12169 ( \12264 , \12257 , \12263 );
buf \U$12170 ( \12265 , \12264 );
buf \U$12171 ( \12266 , RIc0d7c90_14);
buf \U$12172 ( \12267 , RIc0dabe8_115);
xor \U$12173 ( \12268 , \12266 , \12267 );
buf \U$12174 ( \12269 , \12268 );
buf \U$12175 ( \12270 , \12269 );
not \U$12176 ( \12271 , \12270 );
buf \U$12177 ( \12272 , RIc0dac60_116);
buf \U$12178 ( \12273 , RIc0dacd8_117);
xor \U$12179 ( \12274 , \12272 , \12273 );
buf \U$12180 ( \12275 , \12274 );
buf \U$12181 ( \12276 , \12275 );
not \U$12182 ( \12277 , \12276 );
buf \U$12183 ( \12278 , \12277 );
buf \U$12184 ( \12279 , \12278 );
buf \U$12185 ( \12280 , RIc0dac60_116);
not \U$12186 ( \12281 , \12280 );
buf \U$12187 ( \12282 , RIc0dabe8_115);
nand \U$12188 ( \12283 , \12281 , \12282 );
buf \U$12189 ( \12284 , \12283 );
buf \U$12190 ( \12285 , \12284 );
buf \U$12191 ( \12286 , RIc0dabe8_115);
not \U$12192 ( \12287 , \12286 );
buf \U$12193 ( \12288 , RIc0dac60_116);
nand \U$12194 ( \12289 , \12287 , \12288 );
buf \U$12195 ( \12290 , \12289 );
buf \U$12196 ( \12291 , \12290 );
nand \U$12197 ( \12292 , \12285 , \12291 );
buf \U$12198 ( \12293 , \12292 );
buf \U$12199 ( \12294 , \12293 );
nand \U$12200 ( \12295 , \12279 , \12294 );
buf \U$12201 ( \12296 , \12295 );
buf \U$12202 ( \12297 , \12296 );
not \U$12203 ( \12298 , \12297 );
buf \U$12204 ( \12299 , \12298 );
buf \U$12205 ( \12300 , \12299 );
not \U$12206 ( \12301 , \12300 );
or \U$12207 ( \12302 , \12271 , \12301 );
buf \U$12210 ( \12303 , \12275 );
buf \U$12211 ( \12304 , \12303 );
buf \U$12212 ( \12305 , RIc0d7c18_13);
buf \U$12213 ( \12306 , RIc0dabe8_115);
xor \U$12214 ( \12307 , \12305 , \12306 );
buf \U$12215 ( \12308 , \12307 );
buf \U$12216 ( \12309 , \12308 );
nand \U$12217 ( \12310 , \12304 , \12309 );
buf \U$12218 ( \12311 , \12310 );
buf \U$12219 ( \12312 , \12311 );
nand \U$12220 ( \12313 , \12302 , \12312 );
buf \U$12221 ( \12314 , \12313 );
xor \U$12222 ( \12315 , \12265 , \12314 );
buf \U$12223 ( \12316 , RIc0da828_107);
buf \U$12224 ( \12317 , RIc0d8050_22);
xor \U$12225 ( \12318 , \12316 , \12317 );
buf \U$12226 ( \12319 , \12318 );
buf \U$12227 ( \12320 , \12319 );
not \U$12228 ( \12321 , \12320 );
buf \U$12229 ( \12322 , RIc0da8a0_108);
buf \U$12230 ( \12323 , RIc0da918_109);
xnor \U$12231 ( \12324 , \12322 , \12323 );
buf \U$12232 ( \12325 , \12324 );
buf \U$12233 ( \12326 , \12325 );
xor \U$12234 ( \12327 , RIc0da8a0_108, RIc0da828_107);
buf \U$12235 ( \12328 , \12327 );
nand \U$12236 ( \12329 , \12326 , \12328 );
buf \U$12237 ( \12330 , \12329 );
buf \U$12240 ( \12331 , \12330 );
buf \U$12241 ( \12332 , \12331 );
not \U$12242 ( \12333 , \12332 );
buf \U$12243 ( \12334 , \12333 );
buf \U$12244 ( \12335 , \12334 );
not \U$12245 ( \12336 , \12335 );
or \U$12246 ( \12337 , \12321 , \12336 );
buf \U$12247 ( \12338 , RIc0da8a0_108);
buf \U$12248 ( \12339 , RIc0da918_109);
xor \U$12249 ( \12340 , \12338 , \12339 );
buf \U$12250 ( \12341 , \12340 );
buf \U$12253 ( \12342 , \12341 );
buf \U$12254 ( \12343 , \12342 );
xor \U$12255 ( \12344 , RIc0da828_107, RIc0d7fd8_21);
buf \U$12256 ( \12345 , \12344 );
nand \U$12257 ( \12346 , \12343 , \12345 );
buf \U$12258 ( \12347 , \12346 );
buf \U$12259 ( \12348 , \12347 );
nand \U$12260 ( \12349 , \12337 , \12348 );
buf \U$12261 ( \12350 , \12349 );
xor \U$12262 ( \12351 , \12315 , \12350 );
xor \U$12263 ( \12352 , RIc0d9b08_79, RIc0d8d70_50);
buf \U$12264 ( \12353 , \12352 );
not \U$12265 ( \12354 , \12353 );
not \U$12266 ( \12355 , RIc0d9b80_80);
nand \U$12267 ( \12356 , \12355 , RIc0d9b08_79);
not \U$12268 ( \12357 , \12356 );
not \U$12269 ( \12358 , \383 );
or \U$12270 ( \12359 , \12357 , \12358 );
nand \U$12271 ( \12360 , \12359 , \390 );
not \U$12272 ( \12361 , \12360 );
buf \U$12273 ( \12362 , \12361 );
not \U$12274 ( \12363 , \12362 );
or \U$12275 ( \12364 , \12354 , \12363 );
buf \U$12276 ( \12365 , \3985 );
xor \U$12277 ( \12366 , RIc0d9b08_79, RIc0d8cf8_49);
buf \U$12278 ( \12367 , \12366 );
nand \U$12279 ( \12368 , \12365 , \12367 );
buf \U$12280 ( \12369 , \12368 );
buf \U$12281 ( \12370 , \12369 );
nand \U$12282 ( \12371 , \12364 , \12370 );
buf \U$12283 ( \12372 , \12371 );
buf \U$12284 ( \12373 , \12372 );
not \U$12285 ( \12374 , \12373 );
buf \U$12286 ( \12375 , RIc0d7d80_16);
buf \U$12287 ( \12376 , RIc0daaf8_113);
xor \U$12288 ( \12377 , \12375 , \12376 );
buf \U$12289 ( \12378 , \12377 );
buf \U$12290 ( \12379 , \12378 );
not \U$12291 ( \12380 , \12379 );
buf \U$12292 ( \12381 , RIc0dab70_114);
buf \U$12293 ( \12382 , RIc0dabe8_115);
and \U$12294 ( \12383 , \12381 , \12382 );
not \U$12295 ( \12384 , \12381 );
buf \U$12296 ( \12385 , RIc0dabe8_115);
not \U$12297 ( \12386 , \12385 );
buf \U$12298 ( \12387 , \12386 );
buf \U$12299 ( \12388 , \12387 );
and \U$12300 ( \12389 , \12384 , \12388 );
nor \U$12301 ( \12390 , \12383 , \12389 );
buf \U$12302 ( \12391 , \12390 );
buf \U$12303 ( \12392 , \12391 );
not \U$12304 ( \12393 , \12392 );
buf \U$12305 ( \12394 , \12393 );
buf \U$12306 ( \12395 , \12394 );
xor \U$12307 ( \12396 , RIc0dab70_114, RIc0daaf8_113);
buf \U$12308 ( \12397 , \12396 );
nand \U$12309 ( \12398 , \12395 , \12397 );
buf \U$12310 ( \12399 , \12398 );
buf \U$12311 ( \12400 , \12399 );
not \U$12312 ( \12401 , \12400 );
buf \U$12313 ( \12402 , \12401 );
buf \U$12314 ( \12403 , \12402 );
not \U$12315 ( \12404 , \12403 );
or \U$12316 ( \12405 , \12380 , \12404 );
buf \U$12317 ( \12406 , RIc0dabe8_115);
buf \U$12318 ( \12407 , RIc0dab70_114);
xor \U$12319 ( \12408 , \12406 , \12407 );
buf \U$12320 ( \12409 , \12408 );
buf \U$12323 ( \12410 , \12409 );
buf \U$12324 ( \12411 , \12410 );
buf \U$12325 ( \12412 , RIc0d7d08_15);
buf \U$12326 ( \12413 , RIc0daaf8_113);
xor \U$12327 ( \12414 , \12412 , \12413 );
buf \U$12328 ( \12415 , \12414 );
buf \U$12329 ( \12416 , \12415 );
nand \U$12330 ( \12417 , \12411 , \12416 );
buf \U$12331 ( \12418 , \12417 );
buf \U$12332 ( \12419 , \12418 );
nand \U$12333 ( \12420 , \12405 , \12419 );
buf \U$12334 ( \12421 , \12420 );
not \U$12335 ( \12422 , \12421 );
buf \U$12336 ( \12423 , \12422 );
not \U$12337 ( \12424 , \12423 );
or \U$12338 ( \12425 , \12374 , \12424 );
buf \U$12339 ( \12426 , \12372 );
not \U$12340 ( \12427 , \12426 );
buf \U$12341 ( \12428 , \12427 );
buf \U$12342 ( \12429 , \12428 );
buf \U$12343 ( \12430 , \12421 );
nand \U$12344 ( \12431 , \12429 , \12430 );
buf \U$12345 ( \12432 , \12431 );
buf \U$12346 ( \12433 , \12432 );
nand \U$12347 ( \12434 , \12425 , \12433 );
buf \U$12348 ( \12435 , \12434 );
buf \U$12349 ( \12436 , \12435 );
xor \U$12350 ( \12437 , RIc0d9838_73, RIc0d9040_56);
buf \U$12351 ( \12438 , \12437 );
not \U$12352 ( \12439 , \12438 );
buf \U$12353 ( \12440 , \773 );
not \U$12354 ( \12441 , \12440 );
buf \U$12355 ( \12442 , \12441 );
buf \U$12356 ( \12443 , \12442 );
not \U$12357 ( \12444 , \12443 );
or \U$12358 ( \12445 , \12439 , \12444 );
buf \U$12359 ( \12446 , \1856 );
xor \U$12360 ( \12447 , RIc0d9838_73, RIc0d8fc8_55);
buf \U$12361 ( \12448 , \12447 );
nand \U$12362 ( \12449 , \12446 , \12448 );
buf \U$12363 ( \12450 , \12449 );
buf \U$12364 ( \12451 , \12450 );
nand \U$12365 ( \12452 , \12445 , \12451 );
buf \U$12366 ( \12453 , \12452 );
buf \U$12367 ( \12454 , \12453 );
xnor \U$12368 ( \12455 , \12436 , \12454 );
buf \U$12369 ( \12456 , \12455 );
xor \U$12370 ( \12457 , \12351 , \12456 );
buf \U$12371 ( \12458 , RIc0d9220_60);
buf \U$12372 ( \12459 , RIc0d9658_69);
xor \U$12373 ( \12460 , \12458 , \12459 );
buf \U$12374 ( \12461 , \12460 );
buf \U$12375 ( \12462 , \12461 );
not \U$12376 ( \12463 , \12462 );
buf \U$12377 ( \12464 , \4691 );
not \U$12378 ( \12465 , \12464 );
or \U$12379 ( \12466 , \12463 , \12465 );
buf \U$12380 ( \12467 , \284 );
buf \U$12381 ( \12468 , RIc0d91a8_59);
buf \U$12382 ( \12469 , RIc0d9658_69);
xor \U$12383 ( \12470 , \12468 , \12469 );
buf \U$12384 ( \12471 , \12470 );
buf \U$12385 ( \12472 , \12471 );
nand \U$12386 ( \12473 , \12467 , \12472 );
buf \U$12387 ( \12474 , \12473 );
buf \U$12388 ( \12475 , \12474 );
nand \U$12389 ( \12476 , \12466 , \12475 );
buf \U$12390 ( \12477 , \12476 );
buf \U$12391 ( \12478 , \12477 );
not \U$12392 ( \12479 , \12478 );
buf \U$12393 ( \12480 , RIc0d8aa0_44);
buf \U$12394 ( \12481 , RIc0d9dd8_85);
xor \U$12395 ( \12482 , \12480 , \12481 );
buf \U$12396 ( \12483 , \12482 );
buf \U$12397 ( \12484 , \12483 );
not \U$12398 ( \12485 , \12484 );
buf \U$12399 ( \12486 , \5304 );
not \U$12400 ( \12487 , \12486 );
or \U$12401 ( \12488 , \12485 , \12487 );
buf \U$12402 ( \12489 , \2960 );
buf \U$12403 ( \12490 , RIc0d8a28_43);
buf \U$12404 ( \12491 , RIc0d9dd8_85);
xor \U$12405 ( \12492 , \12490 , \12491 );
buf \U$12406 ( \12493 , \12492 );
buf \U$12407 ( \12494 , \12493 );
nand \U$12408 ( \12495 , \12489 , \12494 );
buf \U$12409 ( \12496 , \12495 );
buf \U$12410 ( \12497 , \12496 );
nand \U$12411 ( \12498 , \12488 , \12497 );
buf \U$12412 ( \12499 , \12498 );
buf \U$12413 ( \12500 , \12499 );
not \U$12414 ( \12501 , \12500 );
buf \U$12415 ( \12502 , \12501 );
buf \U$12416 ( \12503 , \12502 );
not \U$12417 ( \12504 , \12503 );
or \U$12418 ( \12505 , \12479 , \12504 );
buf \U$12419 ( \12506 , \12499 );
buf \U$12420 ( \12507 , \12477 );
not \U$12421 ( \12508 , \12507 );
buf \U$12422 ( \12509 , \12508 );
buf \U$12423 ( \12510 , \12509 );
nand \U$12424 ( \12511 , \12506 , \12510 );
buf \U$12425 ( \12512 , \12511 );
buf \U$12426 ( \12513 , \12512 );
nand \U$12427 ( \12514 , \12505 , \12513 );
buf \U$12428 ( \12515 , \12514 );
buf \U$12429 ( \12516 , \12515 );
xor \U$12430 ( \12517 , RIc0daa08_111, RIc0daa80_112);
buf \U$12431 ( \12518 , \12517 );
buf \U$12432 ( \12519 , RIc0daa80_112);
buf \U$12433 ( \12520 , RIc0daaf8_113);
xor \U$12434 ( \12521 , \12519 , \12520 );
buf \U$12435 ( \12522 , \12521 );
buf \U$12436 ( \12523 , \12522 );
not \U$12437 ( \12524 , \12523 );
buf \U$12438 ( \12525 , \12524 );
buf \U$12439 ( \12526 , \12525 );
and \U$12440 ( \12527 , \12518 , \12526 );
buf \U$12441 ( \12528 , \12527 );
buf \U$12444 ( \12529 , \12528 );
buf \U$12445 ( \12530 , \12529 );
not \U$12446 ( \12531 , \12530 );
buf \U$12447 ( \12532 , \12531 );
buf \U$12448 ( \12533 , \12532 );
xor \U$12449 ( \12534 , RIc0daa08_111, RIc0d7e70_18);
buf \U$12450 ( \12535 , \12534 );
not \U$12451 ( \12536 , \12535 );
buf \U$12452 ( \12537 , \12536 );
buf \U$12453 ( \12538 , \12537 );
or \U$12454 ( \12539 , \12533 , \12538 );
buf \U$12457 ( \12540 , \12525 );
buf \U$12460 ( \12541 , \12540 );
buf \U$12461 ( \12542 , \12541 );
buf \U$12462 ( \12543 , RIc0daa08_111);
buf \U$12463 ( \12544 , RIc0d7df8_17);
xor \U$12464 ( \12545 , \12543 , \12544 );
buf \U$12465 ( \12546 , \12545 );
buf \U$12466 ( \12547 , \12546 );
not \U$12467 ( \12548 , \12547 );
buf \U$12468 ( \12549 , \12548 );
buf \U$12469 ( \12550 , \12549 );
or \U$12470 ( \12551 , \12542 , \12550 );
nand \U$12471 ( \12552 , \12539 , \12551 );
buf \U$12472 ( \12553 , \12552 );
buf \U$12473 ( \12554 , \12553 );
not \U$12474 ( \12555 , \12554 );
buf \U$12475 ( \12556 , \12555 );
buf \U$12476 ( \12557 , \12556 );
and \U$12477 ( \12558 , \12516 , \12557 );
not \U$12478 ( \12559 , \12516 );
buf \U$12479 ( \12560 , \12553 );
and \U$12480 ( \12561 , \12559 , \12560 );
nor \U$12481 ( \12562 , \12558 , \12561 );
buf \U$12482 ( \12563 , \12562 );
buf \U$12483 ( \12564 , \12563 );
not \U$12484 ( \12565 , \12564 );
buf \U$12485 ( \12566 , \12565 );
xnor \U$12486 ( \12567 , \12457 , \12566 );
buf \U$12487 ( \12568 , \12567 );
buf \U$12488 ( \12569 , RIc0d8410_30);
buf \U$12489 ( \12570 , RIc0da468_99);
xor \U$12490 ( \12571 , \12569 , \12570 );
buf \U$12491 ( \12572 , \12571 );
buf \U$12492 ( \12573 , \12572 );
not \U$12493 ( \12574 , \12573 );
buf \U$12494 ( \12575 , \2195 );
not \U$12495 ( \12576 , \12575 );
buf \U$12496 ( \12577 , \12576 );
and \U$12497 ( \12578 , \12577 , \2203 );
buf \U$12498 ( \12579 , \12578 );
not \U$12499 ( \12580 , \12579 );
or \U$12500 ( \12581 , \12574 , \12580 );
buf \U$12501 ( \12582 , \12577 );
not \U$12502 ( \12583 , \12582 );
buf \U$12503 ( \12584 , \12583 );
buf \U$12504 ( \12585 , \12584 );
buf \U$12505 ( \12586 , RIc0d8398_29);
buf \U$12506 ( \12587 , RIc0da468_99);
xor \U$12507 ( \12588 , \12586 , \12587 );
buf \U$12508 ( \12589 , \12588 );
buf \U$12509 ( \12590 , \12589 );
nand \U$12510 ( \12591 , \12585 , \12590 );
buf \U$12511 ( \12592 , \12591 );
buf \U$12512 ( \12593 , \12592 );
nand \U$12513 ( \12594 , \12581 , \12593 );
buf \U$12514 ( \12595 , \12594 );
buf \U$12515 ( \12596 , \12595 );
buf \U$12516 ( \12597 , RIc0d86e0_36);
buf \U$12517 ( \12598 , RIc0da198_93);
xor \U$12518 ( \12599 , \12597 , \12598 );
buf \U$12519 ( \12600 , \12599 );
buf \U$12520 ( \12601 , \12600 );
not \U$12521 ( \12602 , \12601 );
buf \U$12522 ( \12603 , \889 );
not \U$12523 ( \12604 , \12603 );
or \U$12524 ( \12605 , \12602 , \12604 );
buf \U$12525 ( \12606 , \481 );
buf \U$12526 ( \12607 , RIc0d8668_35);
buf \U$12527 ( \12608 , RIc0da198_93);
xor \U$12528 ( \12609 , \12607 , \12608 );
buf \U$12529 ( \12610 , \12609 );
buf \U$12530 ( \12611 , \12610 );
nand \U$12531 ( \12612 , \12606 , \12611 );
buf \U$12532 ( \12613 , \12612 );
buf \U$12533 ( \12614 , \12613 );
nand \U$12534 ( \12615 , \12605 , \12614 );
buf \U$12535 ( \12616 , \12615 );
buf \U$12536 ( \12617 , \12616 );
xor \U$12537 ( \12618 , \12596 , \12617 );
buf \U$12538 ( \12619 , RIc0d89b0_42);
buf \U$12539 ( \12620 , RIc0d9ec8_87);
xor \U$12540 ( \12621 , \12619 , \12620 );
buf \U$12541 ( \12622 , \12621 );
buf \U$12542 ( \12623 , \12622 );
not \U$12543 ( \12624 , \12623 );
buf \U$12544 ( \12625 , \4527 );
not \U$12545 ( \12626 , \12625 );
or \U$12546 ( \12627 , \12624 , \12626 );
buf \U$12547 ( \12628 , \816 );
xor \U$12548 ( \12629 , RIc0d9ec8_87, RIc0d8938_41);
buf \U$12549 ( \12630 , \12629 );
nand \U$12550 ( \12631 , \12628 , \12630 );
buf \U$12551 ( \12632 , \12631 );
buf \U$12552 ( \12633 , \12632 );
nand \U$12553 ( \12634 , \12627 , \12633 );
buf \U$12554 ( \12635 , \12634 );
buf \U$12555 ( \12636 , \12635 );
xor \U$12556 ( \12637 , \12618 , \12636 );
buf \U$12557 ( \12638 , \12637 );
buf \U$12558 ( \12639 , RIc0d76f0_2);
buf \U$12559 ( \12640 , RIc0db188_127);
xor \U$12560 ( \12641 , \12639 , \12640 );
buf \U$12561 ( \12642 , \12641 );
buf \U$12562 ( \12643 , \12642 );
not \U$12563 ( \12644 , \12643 );
buf \U$12564 ( \12645 , RIc0db200_128);
not \U$12565 ( \12646 , \12645 );
buf \U$12566 ( \12647 , \12646 );
buf \U$12567 ( \12648 , \12647 );
buf \U$12568 ( \12649 , RIc0db188_127);
nand \U$12569 ( \12650 , \12648 , \12649 );
buf \U$12570 ( \12651 , \12650 );
buf \U$12571 ( \12652 , \12651 );
not \U$12572 ( \12653 , \12652 );
buf \U$12573 ( \12654 , \12653 );
buf \U$12574 ( \12655 , \12654 );
not \U$12575 ( \12656 , \12655 );
or \U$12576 ( \12657 , \12644 , \12656 );
buf \U$12577 ( \12658 , RIc0d7678_1);
buf \U$12578 ( \12659 , RIc0db188_127);
xor \U$12579 ( \12660 , \12658 , \12659 );
buf \U$12580 ( \12661 , \12660 );
buf \U$12581 ( \12662 , \12661 );
buf \U$12582 ( \12663 , RIc0db200_128);
nand \U$12583 ( \12664 , \12662 , \12663 );
buf \U$12584 ( \12665 , \12664 );
buf \U$12585 ( \12666 , \12665 );
nand \U$12586 ( \12667 , \12657 , \12666 );
buf \U$12587 ( \12668 , \12667 );
buf \U$12588 ( \12669 , \12668 );
buf \U$12589 ( \12670 , RIc0d9130_58);
buf \U$12590 ( \12671 , RIc0d9748_71);
xor \U$12591 ( \12672 , \12670 , \12671 );
buf \U$12592 ( \12673 , \12672 );
buf \U$12593 ( \12674 , \12673 );
not \U$12594 ( \12675 , \12674 );
and \U$12595 ( \12676 , \1254 , \1256 );
buf \U$12596 ( \12677 , \12676 );
not \U$12597 ( \12678 , \12677 );
or \U$12598 ( \12679 , \12675 , \12678 );
buf \U$12599 ( \12680 , RIc0d97c0_72);
buf \U$12600 ( \12681 , RIc0d9838_73);
xor \U$12601 ( \12682 , \12680 , \12681 );
buf \U$12602 ( \12683 , \12682 );
buf \U$12603 ( \12684 , \12683 );
buf \U$12604 ( \12685 , RIc0d90b8_57);
buf \U$12605 ( \12686 , RIc0d9748_71);
xor \U$12606 ( \12687 , \12685 , \12686 );
buf \U$12607 ( \12688 , \12687 );
buf \U$12608 ( \12689 , \12688 );
nand \U$12609 ( \12690 , \12684 , \12689 );
buf \U$12610 ( \12691 , \12690 );
buf \U$12611 ( \12692 , \12691 );
nand \U$12612 ( \12693 , \12679 , \12692 );
buf \U$12613 ( \12694 , \12693 );
buf \U$12614 ( \12695 , \12694 );
xor \U$12615 ( \12696 , \12669 , \12695 );
buf \U$12616 ( \12697 , RIc0d85f0_34);
buf \U$12617 ( \12698 , RIc0da288_95);
xor \U$12618 ( \12699 , \12697 , \12698 );
buf \U$12619 ( \12700 , \12699 );
buf \U$12620 ( \12701 , \12700 );
not \U$12621 ( \12702 , \12701 );
buf \U$12622 ( \12703 , \330 );
not \U$12623 ( \12704 , \12703 );
or \U$12624 ( \12705 , \12702 , \12704 );
buf \U$12625 ( \12706 , \344 );
buf \U$12626 ( \12707 , RIc0da288_95);
buf \U$12627 ( \12708 , RIc0d8578_33);
xor \U$12628 ( \12709 , \12707 , \12708 );
buf \U$12629 ( \12710 , \12709 );
buf \U$12630 ( \12711 , \12710 );
nand \U$12631 ( \12712 , \12706 , \12711 );
buf \U$12632 ( \12713 , \12712 );
buf \U$12633 ( \12714 , \12713 );
nand \U$12634 ( \12715 , \12705 , \12714 );
buf \U$12635 ( \12716 , \12715 );
buf \U$12636 ( \12717 , \12716 );
xnor \U$12637 ( \12718 , \12696 , \12717 );
buf \U$12638 ( \12719 , \12718 );
xnor \U$12639 ( \12720 , \12638 , \12719 );
buf \U$12640 ( \12721 , \12720 );
buf \U$12641 ( \12722 , RIc0d8140_24);
buf \U$12642 ( \12723 , RIc0da738_105);
xor \U$12643 ( \12724 , \12722 , \12723 );
buf \U$12644 ( \12725 , \12724 );
buf \U$12645 ( \12726 , \12725 );
not \U$12646 ( \12727 , \12726 );
buf \U$12647 ( \12728 , RIc0da738_105);
buf \U$12648 ( \12729 , RIc0da7b0_106);
xor \U$12649 ( \12730 , \12728 , \12729 );
buf \U$12650 ( \12731 , \12730 );
not \U$12651 ( \12732 , \12731 );
xor \U$12652 ( \12733 , RIc0da828_107, RIc0da7b0_106);
nor \U$12653 ( \12734 , \12732 , \12733 );
buf \U$12654 ( \12735 , \12734 );
buf \U$12656 ( \12736 , \12735 );
buf \U$12657 ( \12737 , \12736 );
not \U$12658 ( \12738 , \12737 );
or \U$12659 ( \12739 , \12727 , \12738 );
buf \U$12660 ( \12740 , RIc0da7b0_106);
buf \U$12661 ( \12741 , RIc0da828_107);
xor \U$12662 ( \12742 , \12740 , \12741 );
buf \U$12663 ( \12743 , \12742 );
buf \U$12666 ( \12744 , \12743 );
buf \U$12667 ( \12745 , \12744 );
buf \U$12668 ( \12746 , RIc0da738_105);
buf \U$12669 ( \12747 , RIc0d80c8_23);
xor \U$12670 ( \12748 , \12746 , \12747 );
buf \U$12671 ( \12749 , \12748 );
buf \U$12672 ( \12750 , \12749 );
nand \U$12673 ( \12751 , \12745 , \12750 );
buf \U$12674 ( \12752 , \12751 );
buf \U$12675 ( \12753 , \12752 );
nand \U$12676 ( \12754 , \12739 , \12753 );
buf \U$12677 ( \12755 , \12754 );
buf \U$12678 ( \12756 , \12755 );
not \U$12679 ( \12757 , \12756 );
buf \U$12680 ( \12758 , RIc0d9a18_77);
buf \U$12681 ( \12759 , RIc0d8e60_52);
xor \U$12682 ( \12760 , \12758 , \12759 );
buf \U$12683 ( \12761 , \12760 );
buf \U$12684 ( \12762 , \12761 );
not \U$12685 ( \12763 , \12762 );
buf \U$12686 ( \12764 , \1431 );
not \U$12687 ( \12765 , \12764 );
or \U$12688 ( \12766 , \12763 , \12765 );
buf \U$12689 ( \12767 , \1196 );
xor \U$12690 ( \12768 , RIc0d9a18_77, RIc0d8de8_51);
buf \U$12691 ( \12769 , \12768 );
nand \U$12692 ( \12770 , \12767 , \12769 );
buf \U$12693 ( \12771 , \12770 );
buf \U$12694 ( \12772 , \12771 );
nand \U$12695 ( \12773 , \12766 , \12772 );
buf \U$12696 ( \12774 , \12773 );
buf \U$12697 ( \12775 , \12774 );
not \U$12698 ( \12776 , \12775 );
buf \U$12699 ( \12777 , \12776 );
buf \U$12700 ( \12778 , \12777 );
not \U$12701 ( \12779 , \12778 );
or \U$12702 ( \12780 , \12757 , \12779 );
buf \U$12703 ( \12781 , \12755 );
buf \U$12704 ( \12782 , \12777 );
or \U$12705 ( \12783 , \12781 , \12782 );
nand \U$12706 ( \12784 , \12780 , \12783 );
buf \U$12707 ( \12785 , \12784 );
buf \U$12708 ( \12786 , \12785 );
buf \U$12709 ( \12787 , RIc0d9478_65);
buf \U$12710 ( \12788 , RIc0d9400_64);
xor \U$12711 ( \12789 , \12787 , \12788 );
buf \U$12712 ( \12790 , \12789 );
buf \U$12713 ( \12791 , \12790 );
not \U$12714 ( \12792 , \12791 );
buf \U$12715 ( \12793 , \1221 );
not \U$12716 ( \12794 , \12793 );
buf \U$12717 ( \12795 , \12794 );
buf \U$12718 ( \12796 , \12795 );
not \U$12719 ( \12797 , \12796 );
or \U$12720 ( \12798 , \12792 , \12797 );
buf \U$12721 ( \12799 , \1229 );
buf \U$12722 ( \12800 , RIc0d9478_65);
buf \U$12723 ( \12801 , RIc0d9388_63);
xor \U$12724 ( \12802 , \12800 , \12801 );
buf \U$12725 ( \12803 , \12802 );
buf \U$12726 ( \12804 , \12803 );
nand \U$12727 ( \12805 , \12799 , \12804 );
buf \U$12728 ( \12806 , \12805 );
buf \U$12729 ( \12807 , \12806 );
nand \U$12730 ( \12808 , \12798 , \12807 );
buf \U$12731 ( \12809 , \12808 );
buf \U$12732 ( \12810 , \12809 );
and \U$12733 ( \12811 , \12786 , \12810 );
not \U$12734 ( \12812 , \12786 );
buf \U$12735 ( \12813 , \12809 );
not \U$12736 ( \12814 , \12813 );
buf \U$12737 ( \12815 , \12814 );
buf \U$12738 ( \12816 , \12815 );
and \U$12739 ( \12817 , \12812 , \12816 );
nor \U$12740 ( \12818 , \12811 , \12817 );
buf \U$12741 ( \12819 , \12818 );
buf \U$12742 ( \12820 , \12819 );
xor \U$12743 ( \12821 , \12721 , \12820 );
buf \U$12744 ( \12822 , \12821 );
buf \U$12745 ( \12823 , \12822 );
xor \U$12746 ( \12824 , \12568 , \12823 );
buf \U$12747 ( \12825 , RIc0d8320_28);
buf \U$12748 ( \12826 , RIc0da558_101);
xor \U$12749 ( \12827 , \12825 , \12826 );
buf \U$12750 ( \12828 , \12827 );
buf \U$12751 ( \12829 , \12828 );
not \U$12752 ( \12830 , \12829 );
buf \U$12753 ( \12831 , \3531 );
not \U$12754 ( \12832 , \12831 );
buf \U$12755 ( \12833 , \12832 );
buf \U$12756 ( \12834 , \12833 );
not \U$12757 ( \12835 , \12834 );
or \U$12758 ( \12836 , \12830 , \12835 );
buf \U$12759 ( \12837 , \3518 );
not \U$12760 ( \12838 , \12837 );
buf \U$12761 ( \12839 , \12838 );
buf \U$12762 ( \12840 , \12839 );
buf \U$12763 ( \12841 , RIc0d82a8_27);
buf \U$12764 ( \12842 , RIc0da558_101);
xor \U$12765 ( \12843 , \12841 , \12842 );
buf \U$12766 ( \12844 , \12843 );
buf \U$12767 ( \12845 , \12844 );
nand \U$12768 ( \12846 , \12840 , \12845 );
buf \U$12769 ( \12847 , \12846 );
buf \U$12770 ( \12848 , \12847 );
nand \U$12771 ( \12849 , \12836 , \12848 );
buf \U$12772 ( \12850 , \12849 );
not \U$12773 ( \12851 , \12850 );
buf \U$12774 ( \12852 , RIc0d78d0_6);
buf \U$12775 ( \12853 , RIc0dafa8_123);
xor \U$12776 ( \12854 , \12852 , \12853 );
buf \U$12777 ( \12855 , \12854 );
buf \U$12778 ( \12856 , \12855 );
not \U$12779 ( \12857 , \12856 );
buf \U$12780 ( \12858 , RIc0dafa8_123);
buf \U$12781 ( \12859 , RIc0db020_124);
xor \U$12782 ( \12860 , \12858 , \12859 );
buf \U$12783 ( \12861 , \12860 );
buf \U$12784 ( \12862 , \12861 );
not \U$12785 ( \12863 , \12862 );
buf \U$12786 ( \12864 , RIc0db020_124);
buf \U$12787 ( \12865 , RIc0db098_125);
xor \U$12788 ( \12866 , \12864 , \12865 );
buf \U$12789 ( \12867 , \12866 );
buf \U$12790 ( \12868 , \12867 );
nor \U$12791 ( \12869 , \12863 , \12868 );
buf \U$12792 ( \12870 , \12869 );
buf \U$12793 ( \12871 , \12870 );
not \U$12794 ( \12872 , \12871 );
or \U$12795 ( \12873 , \12857 , \12872 );
buf \U$12796 ( \12874 , RIc0db020_124);
buf \U$12797 ( \12875 , RIc0db098_125);
xor \U$12798 ( \12876 , \12874 , \12875 );
buf \U$12799 ( \12877 , \12876 );
buf \U$12800 ( \12878 , \12877 );
buf \U$12801 ( \12879 , RIc0d7858_5);
buf \U$12802 ( \12880 , RIc0dafa8_123);
xor \U$12803 ( \12881 , \12879 , \12880 );
buf \U$12804 ( \12882 , \12881 );
buf \U$12805 ( \12883 , \12882 );
nand \U$12806 ( \12884 , \12878 , \12883 );
buf \U$12807 ( \12885 , \12884 );
buf \U$12808 ( \12886 , \12885 );
nand \U$12809 ( \12887 , \12873 , \12886 );
buf \U$12810 ( \12888 , \12887 );
buf \U$12811 ( \12889 , \12888 );
not \U$12812 ( \12890 , \12889 );
buf \U$12813 ( \12891 , \12890 );
not \U$12814 ( \12892 , \12891 );
or \U$12815 ( \12893 , \12851 , \12892 );
buf \U$12816 ( \12894 , \12850 );
not \U$12817 ( \12895 , \12894 );
buf \U$12818 ( \12896 , \12895 );
buf \U$12819 ( \12897 , \12896 );
buf \U$12820 ( \12898 , \12888 );
nand \U$12821 ( \12899 , \12897 , \12898 );
buf \U$12822 ( \12900 , \12899 );
nand \U$12823 ( \12901 , \12893 , \12900 );
xor \U$12824 ( \12902 , RIc0dacd8_117, RIc0d7ba0_12);
buf \U$12825 ( \12903 , \12902 );
not \U$12826 ( \12904 , \12903 );
buf \U$12827 ( \12905 , RIc0dad50_118);
buf \U$12828 ( \12906 , RIc0dadc8_119);
and \U$12829 ( \12907 , \12905 , \12906 );
not \U$12830 ( \12908 , \12905 );
buf \U$12831 ( \12909 , RIc0dadc8_119);
not \U$12832 ( \12910 , \12909 );
buf \U$12833 ( \12911 , \12910 );
buf \U$12834 ( \12912 , \12911 );
and \U$12835 ( \12913 , \12908 , \12912 );
or \U$12836 ( \12914 , \12907 , \12913 );
buf \U$12837 ( \12915 , \12914 );
buf \U$12838 ( \12916 , \12915 );
xor \U$12839 ( \12917 , RIc0dad50_118, RIc0dacd8_117);
buf \U$12840 ( \12918 , \12917 );
nand \U$12841 ( \12919 , \12916 , \12918 );
buf \U$12842 ( \12920 , \12919 );
buf \U$12843 ( \12921 , \12920 );
not \U$12844 ( \12922 , \12921 );
buf \U$12845 ( \12923 , \12922 );
buf \U$12846 ( \12924 , \12923 );
not \U$12847 ( \12925 , \12924 );
buf \U$12848 ( \12926 , \12925 );
buf \U$12849 ( \12927 , \12926 );
not \U$12850 ( \12928 , \12927 );
buf \U$12851 ( \12929 , \12928 );
buf \U$12852 ( \12930 , \12929 );
not \U$12853 ( \12931 , \12930 );
or \U$12854 ( \12932 , \12904 , \12931 );
buf \U$12855 ( \12933 , RIc0dad50_118);
buf \U$12856 ( \12934 , RIc0dadc8_119);
xor \U$12857 ( \12935 , \12933 , \12934 );
buf \U$12858 ( \12936 , \12935 );
buf \U$12861 ( \12937 , \12936 );
buf \U$12862 ( \12938 , \12937 );
buf \U$12863 ( \12939 , RIc0d7b28_11);
buf \U$12864 ( \12940 , RIc0dacd8_117);
xor \U$12865 ( \12941 , \12939 , \12940 );
buf \U$12866 ( \12942 , \12941 );
buf \U$12867 ( \12943 , \12942 );
nand \U$12868 ( \12944 , \12938 , \12943 );
buf \U$12869 ( \12945 , \12944 );
buf \U$12870 ( \12946 , \12945 );
nand \U$12871 ( \12947 , \12932 , \12946 );
buf \U$12872 ( \12948 , \12947 );
xnor \U$12873 ( \12949 , \12901 , \12948 );
buf \U$12874 ( \12950 , RIc0d79c0_8);
buf \U$12875 ( \12951 , RIc0daeb8_121);
xor \U$12876 ( \12952 , \12950 , \12951 );
buf \U$12877 ( \12953 , \12952 );
buf \U$12878 ( \12954 , \12953 );
not \U$12879 ( \12955 , \12954 );
buf \U$12880 ( \12956 , RIc0daf30_122);
buf \U$12881 ( \12957 , RIc0dafa8_123);
xor \U$12882 ( \12958 , \12956 , \12957 );
buf \U$12883 ( \12959 , \12958 );
buf \U$12884 ( \12960 , \12959 );
not \U$12885 ( \12961 , \12960 );
buf \U$12886 ( \12962 , \12961 );
buf \U$12887 ( \12963 , \12962 );
xor \U$12888 ( \12964 , RIc0daf30_122, RIc0daeb8_121);
buf \U$12889 ( \12965 , \12964 );
nand \U$12890 ( \12966 , \12963 , \12965 );
buf \U$12891 ( \12967 , \12966 );
buf \U$12894 ( \12968 , \12967 );
buf \U$12895 ( \12969 , \12968 );
not \U$12896 ( \12970 , \12969 );
buf \U$12897 ( \12971 , \12970 );
buf \U$12898 ( \12972 , \12971 );
not \U$12899 ( \12973 , \12972 );
or \U$12900 ( \12974 , \12955 , \12973 );
buf \U$12903 ( \12975 , \12959 );
buf \U$12904 ( \12976 , \12975 );
buf \U$12905 ( \12977 , RIc0d7948_7);
buf \U$12906 ( \12978 , RIc0daeb8_121);
xor \U$12907 ( \12979 , \12977 , \12978 );
buf \U$12908 ( \12980 , \12979 );
buf \U$12909 ( \12981 , \12980 );
nand \U$12910 ( \12982 , \12976 , \12981 );
buf \U$12911 ( \12983 , \12982 );
buf \U$12912 ( \12984 , \12983 );
nand \U$12913 ( \12985 , \12974 , \12984 );
buf \U$12914 ( \12986 , \12985 );
buf \U$12915 ( \12987 , \12986 );
not \U$12916 ( \12988 , \12987 );
buf \U$12917 ( \12989 , RIc0d7ab0_10);
buf \U$12918 ( \12990 , RIc0dadc8_119);
xor \U$12919 ( \12991 , \12989 , \12990 );
buf \U$12920 ( \12992 , \12991 );
buf \U$12921 ( \12993 , \12992 );
not \U$12922 ( \12994 , \12993 );
xor \U$12923 ( \12995 , RIc0dae40_120, RIc0dadc8_119);
not \U$12924 ( \12996 , \12995 );
buf \U$12925 ( \12997 , RIc0dae40_120);
buf \U$12926 ( \12998 , RIc0daeb8_121);
xor \U$12927 ( \12999 , \12997 , \12998 );
buf \U$12928 ( \13000 , \12999 );
nor \U$12929 ( \13001 , \12996 , \13000 );
buf \U$12930 ( \13002 , \13001 );
not \U$12931 ( \13003 , \13002 );
or \U$12932 ( \13004 , \12994 , \13003 );
buf \U$12935 ( \13005 , \13000 );
buf \U$12936 ( \13006 , \13005 );
buf \U$12937 ( \13007 , RIc0d7a38_9);
buf \U$12938 ( \13008 , RIc0dadc8_119);
xor \U$12939 ( \13009 , \13007 , \13008 );
buf \U$12940 ( \13010 , \13009 );
buf \U$12941 ( \13011 , \13010 );
nand \U$12942 ( \13012 , \13006 , \13011 );
buf \U$12943 ( \13013 , \13012 );
buf \U$12944 ( \13014 , \13013 );
nand \U$12945 ( \13015 , \13004 , \13014 );
buf \U$12946 ( \13016 , \13015 );
buf \U$12947 ( \13017 , \13016 );
not \U$12948 ( \13018 , \13017 );
buf \U$12949 ( \13019 , \13018 );
buf \U$12950 ( \13020 , \13019 );
not \U$12951 ( \13021 , \13020 );
or \U$12952 ( \13022 , \12988 , \13021 );
buf \U$12953 ( \13023 , \12986 );
not \U$12954 ( \13024 , \13023 );
buf \U$12955 ( \13025 , \13024 );
buf \U$12956 ( \13026 , \13025 );
buf \U$12957 ( \13027 , \13016 );
nand \U$12958 ( \13028 , \13026 , \13027 );
buf \U$12959 ( \13029 , \13028 );
buf \U$12960 ( \13030 , \13029 );
nand \U$12961 ( \13031 , \13022 , \13030 );
buf \U$12962 ( \13032 , \13031 );
buf \U$12963 ( \13033 , \13032 );
buf \U$12964 ( \13034 , RIc0da648_103);
buf \U$12965 ( \13035 , RIc0d8230_26);
xor \U$12966 ( \13036 , \13034 , \13035 );
buf \U$12967 ( \13037 , \13036 );
buf \U$12968 ( \13038 , \13037 );
not \U$12969 ( \13039 , \13038 );
buf \U$12970 ( \13040 , \4483 );
not \U$12971 ( \13041 , \13040 );
buf \U$12972 ( \13042 , \13041 );
buf \U$12973 ( \13043 , \13042 );
not \U$12974 ( \13044 , \13043 );
or \U$12975 ( \13045 , \13039 , \13044 );
buf \U$12976 ( \13046 , \4475 );
not \U$12977 ( \13047 , \13046 );
buf \U$12978 ( \13048 , \13047 );
buf \U$12979 ( \13049 , \13048 );
buf \U$12980 ( \13050 , RIc0d81b8_25);
buf \U$12981 ( \13051 , RIc0da648_103);
xor \U$12982 ( \13052 , \13050 , \13051 );
buf \U$12983 ( \13053 , \13052 );
buf \U$12984 ( \13054 , \13053 );
nand \U$12985 ( \13055 , \13049 , \13054 );
buf \U$12986 ( \13056 , \13055 );
buf \U$12987 ( \13057 , \13056 );
nand \U$12988 ( \13058 , \13045 , \13057 );
buf \U$12989 ( \13059 , \13058 );
buf \U$12990 ( \13060 , \13059 );
xnor \U$12991 ( \13061 , \13033 , \13060 );
buf \U$12992 ( \13062 , \13061 );
buf \U$12993 ( \13063 , \13062 );
not \U$12994 ( \13064 , \13063 );
buf \U$12995 ( \13065 , \13064 );
xor \U$12996 ( \13066 , \12949 , \13065 );
buf \U$12997 ( \13067 , RIc0d9bf8_81);
buf \U$12998 ( \13068 , RIc0d8c80_48);
xor \U$12999 ( \13069 , \13067 , \13068 );
buf \U$13000 ( \13070 , \13069 );
buf \U$13001 ( \13071 , \13070 );
not \U$13002 ( \13072 , \13071 );
buf \U$13003 ( \13073 , \1060 );
not \U$13004 ( \13074 , \13073 );
buf \U$13005 ( \13075 , \13074 );
buf \U$13006 ( \13076 , \13075 );
not \U$13007 ( \13077 , \13076 );
or \U$13008 ( \13078 , \13072 , \13077 );
buf \U$13009 ( \13079 , \1078 );
xor \U$13010 ( \13080 , RIc0d9bf8_81, RIc0d8c08_47);
buf \U$13011 ( \13081 , \13080 );
nand \U$13012 ( \13082 , \13079 , \13081 );
buf \U$13013 ( \13083 , \13082 );
buf \U$13014 ( \13084 , \13083 );
nand \U$13015 ( \13085 , \13078 , \13084 );
buf \U$13016 ( \13086 , \13085 );
xor \U$13017 ( \13087 , RIc0da378_97, RIc0d8500_32);
buf \U$13018 ( \13088 , \13087 );
not \U$13019 ( \13089 , \13088 );
buf \U$13020 ( \13090 , \2938 );
not \U$13021 ( \13091 , \13090 );
buf \U$13022 ( \13092 , \13091 );
buf \U$13023 ( \13093 , \13092 );
not \U$13024 ( \13094 , \13093 );
or \U$13025 ( \13095 , \13089 , \13094 );
buf \U$13026 ( \13096 , \734 );
buf \U$13027 ( \13097 , RIc0d8488_31);
buf \U$13028 ( \13098 , RIc0da378_97);
xor \U$13029 ( \13099 , \13097 , \13098 );
buf \U$13030 ( \13100 , \13099 );
buf \U$13031 ( \13101 , \13100 );
nand \U$13032 ( \13102 , \13096 , \13101 );
buf \U$13033 ( \13103 , \13102 );
buf \U$13034 ( \13104 , \13103 );
nand \U$13035 ( \13105 , \13095 , \13104 );
buf \U$13036 ( \13106 , \13105 );
buf \U$13037 ( \13107 , \13106 );
not \U$13038 ( \13108 , \13107 );
buf \U$13039 ( \13109 , \13108 );
xor \U$13040 ( \13110 , \13086 , \13109 );
buf \U$13041 ( \13111 , RIc0da0a8_91);
buf \U$13042 ( \13112 , RIc0d87d0_38);
xor \U$13043 ( \13113 , \13111 , \13112 );
buf \U$13044 ( \13114 , \13113 );
buf \U$13045 ( \13115 , \13114 );
not \U$13046 ( \13116 , \13115 );
buf \U$13047 ( \13117 , \524 );
not \U$13048 ( \13118 , \13117 );
or \U$13049 ( \13119 , \13116 , \13118 );
buf \U$13050 ( \13120 , \533 );
buf \U$13051 ( \13121 , RIc0d8758_37);
buf \U$13052 ( \13122 , RIc0da0a8_91);
xor \U$13053 ( \13123 , \13121 , \13122 );
buf \U$13054 ( \13124 , \13123 );
buf \U$13055 ( \13125 , \13124 );
nand \U$13056 ( \13126 , \13120 , \13125 );
buf \U$13057 ( \13127 , \13126 );
buf \U$13058 ( \13128 , \13127 );
nand \U$13059 ( \13129 , \13119 , \13128 );
buf \U$13060 ( \13130 , \13129 );
xnor \U$13061 ( \13131 , \13110 , \13130 );
not \U$13062 ( \13132 , \13131 );
xor \U$13063 ( \13133 , \13066 , \13132 );
buf \U$13064 ( \13134 , \13133 );
xor \U$13065 ( \13135 , \12824 , \13134 );
buf \U$13066 ( \13136 , \13135 );
buf \U$13067 ( \13137 , \13136 );
xor \U$13068 ( \13138 , RIc0dacd8_117, RIc0d7c18_13);
buf \U$13069 ( \13139 , \13138 );
not \U$13070 ( \13140 , \13139 );
buf \U$13071 ( \13141 , \12923 );
not \U$13072 ( \13142 , \13141 );
buf \U$13073 ( \13143 , \13142 );
buf \U$13074 ( \13144 , \13143 );
not \U$13075 ( \13145 , \13144 );
buf \U$13076 ( \13146 , \13145 );
buf \U$13077 ( \13147 , \13146 );
not \U$13078 ( \13148 , \13147 );
or \U$13079 ( \13149 , \13140 , \13148 );
buf \U$13080 ( \13150 , \12937 );
buf \U$13081 ( \13151 , \12902 );
nand \U$13082 ( \13152 , \13150 , \13151 );
buf \U$13083 ( \13153 , \13152 );
buf \U$13084 ( \13154 , \13153 );
nand \U$13085 ( \13155 , \13149 , \13154 );
buf \U$13086 ( \13156 , \13155 );
xor \U$13087 ( \13157 , RIc0dadc8_119, RIc0d7b28_11);
buf \U$13088 ( \13158 , \13157 );
not \U$13089 ( \13159 , \13158 );
buf \U$13090 ( \13160 , RIc0dae40_120);
buf \U$13091 ( \13161 , RIc0daeb8_121);
and \U$13092 ( \13162 , \13160 , \13161 );
not \U$13093 ( \13163 , \13160 );
buf \U$13094 ( \13164 , RIc0daeb8_121);
not \U$13095 ( \13165 , \13164 );
buf \U$13096 ( \13166 , \13165 );
buf \U$13097 ( \13167 , \13166 );
and \U$13098 ( \13168 , \13163 , \13167 );
nor \U$13099 ( \13169 , \13162 , \13168 );
buf \U$13100 ( \13170 , \13169 );
buf \U$13101 ( \13171 , \13170 );
not \U$13102 ( \13172 , \13171 );
buf \U$13103 ( \13173 , \13172 );
buf \U$13104 ( \13174 , \13173 );
buf \U$13105 ( \13175 , \12995 );
nand \U$13106 ( \13176 , \13174 , \13175 );
buf \U$13107 ( \13177 , \13176 );
buf \U$13110 ( \13178 , \13177 );
buf \U$13111 ( \13179 , \13178 );
not \U$13112 ( \13180 , \13179 );
buf \U$13113 ( \13181 , \13180 );
buf \U$13114 ( \13182 , \13181 );
not \U$13115 ( \13183 , \13182 );
or \U$13116 ( \13184 , \13159 , \13183 );
buf \U$13117 ( \13185 , \13005 );
buf \U$13118 ( \13186 , \12992 );
nand \U$13119 ( \13187 , \13185 , \13186 );
buf \U$13120 ( \13188 , \13187 );
buf \U$13121 ( \13189 , \13188 );
nand \U$13122 ( \13190 , \13184 , \13189 );
buf \U$13123 ( \13191 , \13190 );
xor \U$13124 ( \13192 , \13156 , \13191 );
buf \U$13125 ( \13193 , \13192 );
buf \U$13126 ( \13194 , RIc0d8c08_47);
buf \U$13127 ( \13195 , RIc0d9ce8_83);
xor \U$13128 ( \13196 , \13194 , \13195 );
buf \U$13129 ( \13197 , \13196 );
buf \U$13130 ( \13198 , \13197 );
not \U$13131 ( \13199 , \13198 );
buf \U$13132 ( \13200 , \1736 );
not \U$13133 ( \13201 , \13200 );
or \U$13134 ( \13202 , \13199 , \13201 );
buf \U$13135 ( \13203 , \584 );
buf \U$13136 ( \13204 , \12245 );
nand \U$13137 ( \13205 , \13203 , \13204 );
buf \U$13138 ( \13206 , \13205 );
buf \U$13139 ( \13207 , \13206 );
nand \U$13140 ( \13208 , \13202 , \13207 );
buf \U$13141 ( \13209 , \13208 );
buf \U$13142 ( \13210 , \13209 );
xor \U$13143 ( \13211 , \13193 , \13210 );
buf \U$13144 ( \13212 , \13211 );
buf \U$13145 ( \13213 , \13212 );
buf \U$13146 ( \13214 , \4904 );
buf \U$13147 ( \13215 , RIc0d9388_63);
buf \U$13148 ( \13216 , RIc0d9568_67);
xor \U$13149 ( \13217 , \13215 , \13216 );
buf \U$13150 ( \13218 , \13217 );
buf \U$13151 ( \13219 , \13218 );
not \U$13152 ( \13220 , \13219 );
buf \U$13153 ( \13221 , \13220 );
buf \U$13154 ( \13222 , \13221 );
or \U$13155 ( \13223 , \13214 , \13222 );
buf \U$13156 ( \13224 , \685 );
not \U$13157 ( \13225 , \13224 );
buf \U$13158 ( \13226 , \13225 );
buf \U$13159 ( \13227 , \13226 );
buf \U$13160 ( \13228 , RIc0d9310_62);
buf \U$13161 ( \13229 , RIc0d9568_67);
xor \U$13162 ( \13230 , \13228 , \13229 );
buf \U$13163 ( \13231 , \13230 );
buf \U$13164 ( \13232 , \13231 );
not \U$13165 ( \13233 , \13232 );
buf \U$13166 ( \13234 , \13233 );
buf \U$13167 ( \13235 , \13234 );
or \U$13168 ( \13236 , \13227 , \13235 );
nand \U$13169 ( \13237 , \13223 , \13236 );
buf \U$13170 ( \13238 , \13237 );
buf \U$13171 ( \13239 , \13238 );
buf \U$13172 ( \13240 , RIc0d8578_33);
buf \U$13173 ( \13241 , RIc0da378_97);
xor \U$13174 ( \13242 , \13240 , \13241 );
buf \U$13175 ( \13243 , \13242 );
buf \U$13176 ( \13244 , \13243 );
not \U$13177 ( \13245 , \13244 );
buf \U$13178 ( \13246 , \2941 );
not \U$13179 ( \13247 , \13246 );
or \U$13180 ( \13248 , \13245 , \13247 );
buf \U$13181 ( \13249 , \734 );
buf \U$13182 ( \13250 , \13087 );
nand \U$13183 ( \13251 , \13249 , \13250 );
buf \U$13184 ( \13252 , \13251 );
buf \U$13185 ( \13253 , \13252 );
nand \U$13186 ( \13254 , \13248 , \13253 );
buf \U$13187 ( \13255 , \13254 );
buf \U$13188 ( \13256 , \13255 );
xor \U$13189 ( \13257 , \13239 , \13256 );
buf \U$13190 ( \13258 , \12331 );
buf \U$13191 ( \13259 , RIc0d80c8_23);
buf \U$13192 ( \13260 , RIc0da828_107);
xor \U$13193 ( \13261 , \13259 , \13260 );
buf \U$13194 ( \13262 , \13261 );
buf \U$13195 ( \13263 , \13262 );
not \U$13196 ( \13264 , \13263 );
buf \U$13197 ( \13265 , \13264 );
buf \U$13198 ( \13266 , \13265 );
or \U$13199 ( \13267 , \13258 , \13266 );
buf \U$13200 ( \13268 , \12342 );
not \U$13201 ( \13269 , \13268 );
buf \U$13202 ( \13270 , \13269 );
buf \U$13203 ( \13271 , \13270 );
buf \U$13204 ( \13272 , \12319 );
not \U$13205 ( \13273 , \13272 );
buf \U$13206 ( \13274 , \13273 );
buf \U$13207 ( \13275 , \13274 );
or \U$13208 ( \13276 , \13271 , \13275 );
nand \U$13209 ( \13277 , \13267 , \13276 );
buf \U$13210 ( \13278 , \13277 );
buf \U$13211 ( \13279 , \13278 );
xor \U$13212 ( \13280 , \13257 , \13279 );
buf \U$13213 ( \13281 , \13280 );
buf \U$13214 ( \13282 , \13281 );
xor \U$13215 ( \13283 , \13213 , \13282 );
buf \U$13216 ( \13284 , RIc0d8848_39);
buf \U$13217 ( \13285 , RIc0da0a8_91);
xor \U$13218 ( \13286 , \13284 , \13285 );
buf \U$13219 ( \13287 , \13286 );
buf \U$13220 ( \13288 , \13287 );
not \U$13221 ( \13289 , \13288 );
buf \U$13222 ( \13290 , \704 );
not \U$13223 ( \13291 , \13290 );
or \U$13224 ( \13292 , \13289 , \13291 );
buf \U$13227 ( \13293 , \533 );
buf \U$13228 ( \13294 , \13293 );
buf \U$13229 ( \13295 , \13114 );
nand \U$13230 ( \13296 , \13294 , \13295 );
buf \U$13231 ( \13297 , \13296 );
buf \U$13232 ( \13298 , \13297 );
nand \U$13233 ( \13299 , \13292 , \13298 );
buf \U$13234 ( \13300 , \13299 );
buf \U$13235 ( \13301 , \13300 );
buf \U$13236 ( \13302 , RIc0d7a38_9);
buf \U$13237 ( \13303 , RIc0daeb8_121);
xor \U$13238 ( \13304 , \13302 , \13303 );
buf \U$13239 ( \13305 , \13304 );
buf \U$13240 ( \13306 , \13305 );
not \U$13241 ( \13307 , \13306 );
buf \U$13242 ( \13308 , \12968 );
not \U$13243 ( \13309 , \13308 );
buf \U$13244 ( \13310 , \13309 );
buf \U$13245 ( \13311 , \13310 );
not \U$13246 ( \13312 , \13311 );
or \U$13247 ( \13313 , \13307 , \13312 );
buf \U$13250 ( \13314 , \12975 );
buf \U$13251 ( \13315 , \13314 );
buf \U$13252 ( \13316 , \12953 );
nand \U$13253 ( \13317 , \13315 , \13316 );
buf \U$13254 ( \13318 , \13317 );
buf \U$13255 ( \13319 , \13318 );
nand \U$13256 ( \13320 , \13313 , \13319 );
buf \U$13257 ( \13321 , \13320 );
buf \U$13258 ( \13322 , \13321 );
xor \U$13259 ( \13323 , \13301 , \13322 );
buf \U$13260 ( \13324 , RIc0d9310_62);
buf \U$13261 ( \13325 , RIc0d9658_69);
xor \U$13262 ( \13326 , \13324 , \13325 );
buf \U$13263 ( \13327 , \13326 );
buf \U$13264 ( \13328 , \13327 );
not \U$13265 ( \13329 , \13328 );
buf \U$13266 ( \13330 , \861 );
not \U$13267 ( \13331 , \13330 );
buf \U$13268 ( \13332 , \13331 );
buf \U$13269 ( \13333 , \13332 );
not \U$13270 ( \13334 , \13333 );
or \U$13271 ( \13335 , \13329 , \13334 );
buf \U$13272 ( \13336 , \874 );
xor \U$13273 ( \13337 , RIc0d9658_69, RIc0d9298_61);
buf \U$13274 ( \13338 , \13337 );
nand \U$13275 ( \13339 , \13336 , \13338 );
buf \U$13276 ( \13340 , \13339 );
buf \U$13277 ( \13341 , \13340 );
nand \U$13278 ( \13342 , \13335 , \13341 );
buf \U$13279 ( \13343 , \13342 );
buf \U$13280 ( \13344 , \13343 );
not \U$13281 ( \13345 , \13344 );
buf \U$13282 ( \13346 , RIc0d9400_64);
buf \U$13283 ( \13347 , RIc0d95e0_68);
nand \U$13284 ( \13348 , \13346 , \13347 );
buf \U$13285 ( \13349 , \13348 );
buf \U$13286 ( \13350 , RIc0d9400_64);
buf \U$13287 ( \13351 , RIc0d95e0_68);
or \U$13288 ( \13352 , \13350 , \13351 );
buf \U$13289 ( \13353 , RIc0d9658_69);
nand \U$13290 ( \13354 , \13352 , \13353 );
buf \U$13291 ( \13355 , \13354 );
nand \U$13292 ( \13356 , \13349 , RIc0d9568_67, \13355 );
buf \U$13293 ( \13357 , \13356 );
nor \U$13294 ( \13358 , \13345 , \13357 );
buf \U$13295 ( \13359 , \13358 );
buf \U$13296 ( \13360 , \13359 );
xor \U$13297 ( \13361 , \13323 , \13360 );
buf \U$13298 ( \13362 , \13361 );
buf \U$13299 ( \13363 , \13362 );
and \U$13300 ( \13364 , \13283 , \13363 );
and \U$13301 ( \13365 , \13213 , \13282 );
or \U$13302 ( \13366 , \13364 , \13365 );
buf \U$13303 ( \13367 , \13366 );
buf \U$13304 ( \13368 , \13367 );
xor \U$13305 ( \13369 , \13301 , \13322 );
and \U$13306 ( \13370 , \13369 , \13360 );
and \U$13307 ( \13371 , \13301 , \13322 );
or \U$13308 ( \13372 , \13370 , \13371 );
buf \U$13309 ( \13373 , \13372 );
buf \U$13310 ( \13374 , \13373 );
buf \U$13311 ( \13375 , RIc0d8f50_54);
buf \U$13312 ( \13376 , RIc0d9928_75);
xor \U$13313 ( \13377 , \13375 , \13376 );
buf \U$13314 ( \13378 , \13377 );
buf \U$13315 ( \13379 , \13378 );
not \U$13316 ( \13380 , \13379 );
buf \U$13317 ( \13381 , \1124 );
not \U$13318 ( \13382 , \13381 );
buf \U$13319 ( \13383 , \13382 );
buf \U$13320 ( \13384 , \13383 );
not \U$13321 ( \13385 , \13384 );
or \U$13322 ( \13386 , \13380 , \13385 );
buf \U$13323 ( \13387 , \1562 );
not \U$13324 ( \13388 , \13387 );
buf \U$13325 ( \13389 , \13388 );
buf \U$13326 ( \13390 , \13389 );
buf \U$13327 ( \13391 , RIc0d8ed8_53);
buf \U$13328 ( \13392 , RIc0d9928_75);
xor \U$13329 ( \13393 , \13391 , \13392 );
buf \U$13330 ( \13394 , \13393 );
buf \U$13331 ( \13395 , \13394 );
nand \U$13332 ( \13396 , \13390 , \13395 );
buf \U$13333 ( \13397 , \13396 );
buf \U$13334 ( \13398 , \13397 );
nand \U$13335 ( \13399 , \13386 , \13398 );
buf \U$13336 ( \13400 , \13399 );
buf \U$13337 ( \13401 , \13400 );
xor \U$13338 ( \13402 , RIc0da918_109, RIc0d7f60_20);
buf \U$13339 ( \13403 , \13402 );
not \U$13340 ( \13404 , \13403 );
buf \U$13341 ( \13405 , RIc0da990_110);
buf \U$13342 ( \13406 , RIc0daa08_111);
xor \U$13343 ( \13407 , \13405 , \13406 );
buf \U$13344 ( \13408 , \13407 );
buf \U$13345 ( \13409 , \13408 );
not \U$13346 ( \13410 , \13409 );
buf \U$13347 ( \13411 , \13410 );
buf \U$13348 ( \13412 , \13411 );
xor \U$13349 ( \13413 , RIc0da990_110, RIc0da918_109);
buf \U$13350 ( \13414 , \13413 );
nand \U$13351 ( \13415 , \13412 , \13414 );
buf \U$13352 ( \13416 , \13415 );
buf \U$13353 ( \13417 , \13416 );
not \U$13354 ( \13418 , \13417 );
buf \U$13355 ( \13419 , \13418 );
buf \U$13356 ( \13420 , \13419 );
not \U$13357 ( \13421 , \13420 );
or \U$13358 ( \13422 , \13404 , \13421 );
buf \U$13361 ( \13423 , \13411 );
buf \U$13362 ( \13424 , \13423 );
not \U$13363 ( \13425 , \13424 );
buf \U$13364 ( \13426 , \13425 );
buf \U$13365 ( \13427 , \13426 );
buf \U$13366 ( \13428 , RIc0d7ee8_19);
buf \U$13367 ( \13429 , RIc0da918_109);
xor \U$13368 ( \13430 , \13428 , \13429 );
buf \U$13369 ( \13431 , \13430 );
buf \U$13370 ( \13432 , \13431 );
nand \U$13371 ( \13433 , \13427 , \13432 );
buf \U$13372 ( \13434 , \13433 );
buf \U$13373 ( \13435 , \13434 );
nand \U$13374 ( \13436 , \13422 , \13435 );
buf \U$13375 ( \13437 , \13436 );
buf \U$13376 ( \13438 , \13437 );
xor \U$13377 ( \13439 , \13401 , \13438 );
buf \U$13378 ( \13440 , RIc0d77e0_4);
buf \U$13379 ( \13441 , RIc0db098_125);
xor \U$13380 ( \13442 , \13440 , \13441 );
buf \U$13381 ( \13443 , \13442 );
buf \U$13382 ( \13444 , \13443 );
not \U$13383 ( \13445 , \13444 );
buf \U$13384 ( \13446 , RIc0db110_126);
buf \U$13385 ( \13447 , RIc0db188_127);
xor \U$13386 ( \13448 , \13446 , \13447 );
buf \U$13387 ( \13449 , \13448 );
buf \U$13388 ( \13450 , \13449 );
not \U$13389 ( \13451 , \13450 );
buf \U$13390 ( \13452 , \13451 );
buf \U$13391 ( \13453 , \13452 );
xor \U$13392 ( \13454 , RIc0db110_126, RIc0db098_125);
buf \U$13393 ( \13455 , \13454 );
nand \U$13394 ( \13456 , \13453 , \13455 );
buf \U$13395 ( \13457 , \13456 );
buf \U$13396 ( \13458 , \13457 );
not \U$13397 ( \13459 , \13458 );
buf \U$13398 ( \13460 , \13459 );
buf \U$13401 ( \13461 , \13460 );
buf \U$13402 ( \13462 , \13461 );
not \U$13403 ( \13463 , \13462 );
or \U$13404 ( \13464 , \13445 , \13463 );
buf \U$13407 ( \13465 , \13449 );
buf \U$13408 ( \13466 , \13465 );
buf \U$13409 ( \13467 , RIc0d7768_3);
buf \U$13410 ( \13468 , RIc0db098_125);
xor \U$13411 ( \13469 , \13467 , \13468 );
buf \U$13412 ( \13470 , \13469 );
buf \U$13413 ( \13471 , \13470 );
nand \U$13414 ( \13472 , \13466 , \13471 );
buf \U$13415 ( \13473 , \13472 );
buf \U$13416 ( \13474 , \13473 );
nand \U$13417 ( \13475 , \13464 , \13474 );
buf \U$13418 ( \13476 , \13475 );
buf \U$13419 ( \13477 , \13476 );
xor \U$13420 ( \13478 , \13439 , \13477 );
buf \U$13421 ( \13479 , \13478 );
buf \U$13422 ( \13480 , \13479 );
xor \U$13423 ( \13481 , \13374 , \13480 );
buf \U$13424 ( \13482 , \6823 );
buf \U$13425 ( \13483 , RIc0d88c0_40);
buf \U$13426 ( \13484 , RIc0d9fb8_89);
xor \U$13427 ( \13485 , \13483 , \13484 );
buf \U$13428 ( \13486 , \13485 );
buf \U$13429 ( \13487 , \13486 );
not \U$13430 ( \13488 , \13487 );
buf \U$13431 ( \13489 , \13488 );
buf \U$13432 ( \13490 , \13489 );
or \U$13433 ( \13491 , \13482 , \13490 );
buf \U$13434 ( \13492 , \441 );
not \U$13435 ( \13493 , \13492 );
buf \U$13436 ( \13494 , \13493 );
buf \U$13437 ( \13495 , \13494 );
buf \U$13438 ( \13496 , RIc0d8848_39);
buf \U$13439 ( \13497 , RIc0d9fb8_89);
xor \U$13440 ( \13498 , \13496 , \13497 );
buf \U$13441 ( \13499 , \13498 );
buf \U$13442 ( \13500 , \13499 );
not \U$13443 ( \13501 , \13500 );
buf \U$13444 ( \13502 , \13501 );
buf \U$13445 ( \13503 , \13502 );
or \U$13446 ( \13504 , \13495 , \13503 );
nand \U$13447 ( \13505 , \13491 , \13504 );
buf \U$13448 ( \13506 , \13505 );
buf \U$13449 ( \13507 , \13506 );
buf \U$13450 ( \13508 , RIc0d9400_64);
buf \U$13451 ( \13509 , RIc0d94f0_66);
or \U$13452 ( \13510 , \13508 , \13509 );
buf \U$13453 ( \13511 , RIc0d9568_67);
nand \U$13454 ( \13512 , \13510 , \13511 );
buf \U$13455 ( \13513 , \13512 );
buf \U$13456 ( \13514 , \13513 );
buf \U$13457 ( \13515 , RIc0d9400_64);
buf \U$13458 ( \13516 , RIc0d94f0_66);
nand \U$13459 ( \13517 , \13515 , \13516 );
buf \U$13460 ( \13518 , \13517 );
buf \U$13461 ( \13519 , \13518 );
buf \U$13462 ( \13520 , RIc0d9478_65);
and \U$13463 ( \13521 , \13514 , \13519 , \13520 );
buf \U$13464 ( \13522 , \13521 );
buf \U$13465 ( \13523 , \13522 );
buf \U$13466 ( \13524 , \13231 );
not \U$13467 ( \13525 , \13524 );
buf \U$13468 ( \13526 , \678 );
not \U$13469 ( \13527 , \13526 );
or \U$13470 ( \13528 , \13525 , \13527 );
buf \U$13471 ( \13529 , \686 );
buf \U$13472 ( \13530 , RIc0d9298_61);
buf \U$13473 ( \13531 , RIc0d9568_67);
xor \U$13474 ( \13532 , \13530 , \13531 );
buf \U$13475 ( \13533 , \13532 );
buf \U$13476 ( \13534 , \13533 );
nand \U$13477 ( \13535 , \13529 , \13534 );
buf \U$13478 ( \13536 , \13535 );
buf \U$13479 ( \13537 , \13536 );
nand \U$13480 ( \13538 , \13528 , \13537 );
buf \U$13481 ( \13539 , \13538 );
buf \U$13482 ( \13540 , \13539 );
xor \U$13483 ( \13541 , \13523 , \13540 );
buf \U$13484 ( \13542 , \13541 );
buf \U$13485 ( \13543 , \13542 );
xor \U$13486 ( \13544 , \13507 , \13543 );
buf \U$13487 ( \13545 , \1229 );
buf \U$13488 ( \13546 , RIc0d9400_64);
and \U$13489 ( \13547 , \13545 , \13546 );
buf \U$13490 ( \13548 , \13547 );
buf \U$13491 ( \13549 , \13548 );
buf \U$13492 ( \13550 , \13337 );
not \U$13493 ( \13551 , \13550 );
buf \U$13494 ( \13552 , \4691 );
not \U$13495 ( \13553 , \13552 );
or \U$13496 ( \13554 , \13551 , \13553 );
buf \U$13497 ( \13555 , \284 );
buf \U$13498 ( \13556 , \12461 );
nand \U$13499 ( \13557 , \13555 , \13556 );
buf \U$13500 ( \13558 , \13557 );
buf \U$13501 ( \13559 , \13558 );
nand \U$13502 ( \13560 , \13554 , \13559 );
buf \U$13503 ( \13561 , \13560 );
buf \U$13504 ( \13562 , \13561 );
xor \U$13505 ( \13563 , \13549 , \13562 );
xor \U$13506 ( \13564 , RIc0da198_93, RIc0d8758_37);
buf \U$13507 ( \13565 , \13564 );
not \U$13508 ( \13566 , \13565 );
buf \U$13509 ( \13567 , \473 );
not \U$13510 ( \13568 , \13567 );
buf \U$13511 ( \13569 , \13568 );
buf \U$13512 ( \13570 , \13569 );
not \U$13513 ( \13571 , \13570 );
or \U$13514 ( \13572 , \13566 , \13571 );
buf \U$13515 ( \13573 , \4008 );
buf \U$13516 ( \13574 , \12600 );
nand \U$13517 ( \13575 , \13573 , \13574 );
buf \U$13518 ( \13576 , \13575 );
buf \U$13519 ( \13577 , \13576 );
nand \U$13520 ( \13578 , \13572 , \13577 );
buf \U$13521 ( \13579 , \13578 );
buf \U$13522 ( \13580 , \13579 );
and \U$13523 ( \13581 , \13563 , \13580 );
and \U$13524 ( \13582 , \13549 , \13562 );
or \U$13525 ( \13583 , \13581 , \13582 );
buf \U$13526 ( \13584 , \13583 );
buf \U$13527 ( \13585 , \13584 );
xor \U$13528 ( \13586 , \13544 , \13585 );
buf \U$13529 ( \13587 , \13586 );
buf \U$13530 ( \13588 , \13587 );
xor \U$13531 ( \13589 , \13481 , \13588 );
buf \U$13532 ( \13590 , \13589 );
buf \U$13533 ( \13591 , \13590 );
xor \U$13534 ( \13592 , \13368 , \13591 );
buf \U$13535 ( \13593 , \12396 );
buf \U$13536 ( \13594 , RIc0d7ee8_19);
buf \U$13537 ( \13595 , RIc0daaf8_113);
xor \U$13538 ( \13596 , \13594 , \13595 );
buf \U$13539 ( \13597 , \13596 );
buf \U$13540 ( \13598 , \13597 );
nand \U$13541 ( \13599 , \13593 , \13598 );
buf \U$13542 ( \13600 , \13599 );
buf \U$13543 ( \13601 , \13600 );
buf \U$13544 ( \13602 , \12409 );
or \U$13545 ( \13603 , \13601 , \13602 );
buf \U$13546 ( \13604 , \12409 );
xor \U$13547 ( \13605 , RIc0daaf8_113, RIc0d7e70_18);
buf \U$13548 ( \13606 , \13605 );
nand \U$13549 ( \13607 , \13604 , \13606 );
buf \U$13550 ( \13608 , \13607 );
buf \U$13551 ( \13609 , \13608 );
nand \U$13552 ( \13610 , \13603 , \13609 );
buf \U$13553 ( \13611 , \13610 );
buf \U$13554 ( \13612 , \13611 );
xor \U$13555 ( \13613 , RIc0d9fb8_89, RIc0d89b0_42);
buf \U$13556 ( \13614 , \13613 );
not \U$13557 ( \13615 , \13614 );
buf \U$13558 ( \13616 , \427 );
not \U$13559 ( \13617 , \13616 );
buf \U$13560 ( \13618 , \13617 );
buf \U$13561 ( \13619 , \13618 );
not \U$13562 ( \13620 , \13619 );
or \U$13563 ( \13621 , \13615 , \13620 );
buf \U$13564 ( \13622 , \429 );
buf \U$13565 ( \13623 , RIc0d8a28_43);
buf \U$13566 ( \13624 , RIc0d9fb8_89);
xor \U$13567 ( \13625 , \13623 , \13624 );
buf \U$13568 ( \13626 , \13625 );
buf \U$13569 ( \13627 , \13626 );
nand \U$13570 ( \13628 , \13622 , \13627 );
buf \U$13571 ( \13629 , \13628 );
buf \U$13572 ( \13630 , \13629 );
buf \U$13573 ( \13631 , \441 );
or \U$13574 ( \13632 , \13630 , \13631 );
nand \U$13575 ( \13633 , \13621 , \13632 );
buf \U$13576 ( \13634 , \13633 );
buf \U$13577 ( \13635 , \13634 );
xor \U$13578 ( \13636 , \13612 , \13635 );
xor \U$13579 ( \13637 , RIc0d9ce8_83, RIc0d8cf8_49);
buf \U$13580 ( \13638 , \13637 );
not \U$13581 ( \13639 , \13638 );
buf \U$13582 ( \13640 , \12254 );
not \U$13583 ( \13641 , \13640 );
or \U$13584 ( \13642 , \13639 , \13641 );
buf \U$13585 ( \13643 , \993 );
xor \U$13586 ( \13644 , RIc0d9ce8_83, RIc0d8c80_48);
buf \U$13587 ( \13645 , \13644 );
nand \U$13588 ( \13646 , \13643 , \13645 );
buf \U$13589 ( \13647 , \13646 );
buf \U$13590 ( \13648 , \13647 );
nand \U$13591 ( \13649 , \13642 , \13648 );
buf \U$13592 ( \13650 , \13649 );
buf \U$13593 ( \13651 , \13650 );
and \U$13594 ( \13652 , \13636 , \13651 );
and \U$13595 ( \13653 , \13612 , \13635 );
or \U$13596 ( \13654 , \13652 , \13653 );
buf \U$13597 ( \13655 , \13654 );
buf \U$13598 ( \13656 , \13655 );
buf \U$13599 ( \13657 , \1176 );
buf \U$13600 ( \13658 , RIc0d8fc8_55);
buf \U$13601 ( \13659 , RIc0d9a18_77);
xor \U$13602 ( \13660 , \13658 , \13659 );
buf \U$13603 ( \13661 , \13660 );
buf \U$13604 ( \13662 , \13661 );
nand \U$13605 ( \13663 , \13657 , \13662 );
buf \U$13606 ( \13664 , \13663 );
buf \U$13607 ( \13665 , \13664 );
buf \U$13608 ( \13666 , \1588 );
or \U$13609 ( \13667 , \13665 , \13666 );
buf \U$13610 ( \13668 , \3742 );
xor \U$13611 ( \13669 , RIc0d9a18_77, RIc0d8f50_54);
buf \U$13612 ( \13670 , \13669 );
nand \U$13613 ( \13671 , \13668 , \13670 );
buf \U$13614 ( \13672 , \13671 );
buf \U$13615 ( \13673 , \13672 );
nand \U$13616 ( \13674 , \13667 , \13673 );
buf \U$13617 ( \13675 , \13674 );
buf \U$13618 ( \13676 , \13675 );
xor \U$13619 ( \13677 , RIc0dacd8_117, RIc0d7d08_15);
buf \U$13620 ( \13678 , \13677 );
not \U$13621 ( \13679 , \13678 );
not \U$13622 ( \13680 , \12936 );
nand \U$13623 ( \13681 , \13680 , \12917 );
buf \U$13624 ( \13682 , \13681 );
not \U$13625 ( \13683 , \13682 );
buf \U$13626 ( \13684 , \13683 );
buf \U$13627 ( \13685 , \13684 );
not \U$13628 ( \13686 , \13685 );
or \U$13629 ( \13687 , \13679 , \13686 );
buf \U$13630 ( \13688 , \12937 );
xor \U$13631 ( \13689 , RIc0dacd8_117, RIc0d7c90_14);
buf \U$13632 ( \13690 , \13689 );
nand \U$13633 ( \13691 , \13688 , \13690 );
buf \U$13634 ( \13692 , \13691 );
buf \U$13635 ( \13693 , \13692 );
nand \U$13636 ( \13694 , \13687 , \13693 );
buf \U$13637 ( \13695 , \13694 );
buf \U$13638 ( \13696 , \13695 );
xor \U$13639 ( \13697 , \13676 , \13696 );
buf \U$13640 ( \13698 , RIc0da648_103);
buf \U$13641 ( \13699 , RIc0d8398_29);
xor \U$13642 ( \13700 , \13698 , \13699 );
buf \U$13643 ( \13701 , \13700 );
buf \U$13644 ( \13702 , \13701 );
not \U$13645 ( \13703 , \13702 );
buf \U$13646 ( \13704 , \4483 );
not \U$13647 ( \13705 , \13704 );
buf \U$13648 ( \13706 , \13705 );
buf \U$13649 ( \13707 , \13706 );
not \U$13650 ( \13708 , \13707 );
or \U$13651 ( \13709 , \13703 , \13708 );
buf \U$13652 ( \13710 , \4475 );
not \U$13653 ( \13711 , \13710 );
buf \U$13654 ( \13712 , \13711 );
buf \U$13655 ( \13713 , \13712 );
buf \U$13656 ( \13714 , RIc0d8320_28);
buf \U$13657 ( \13715 , RIc0da648_103);
xor \U$13658 ( \13716 , \13714 , \13715 );
buf \U$13659 ( \13717 , \13716 );
buf \U$13660 ( \13718 , \13717 );
nand \U$13661 ( \13719 , \13713 , \13718 );
buf \U$13662 ( \13720 , \13719 );
buf \U$13663 ( \13721 , \13720 );
nand \U$13664 ( \13722 , \13709 , \13721 );
buf \U$13665 ( \13723 , \13722 );
buf \U$13666 ( \13724 , \13723 );
and \U$13667 ( \13725 , \13697 , \13724 );
and \U$13668 ( \13726 , \13676 , \13696 );
or \U$13669 ( \13727 , \13725 , \13726 );
buf \U$13670 ( \13728 , \13727 );
buf \U$13671 ( \13729 , \13728 );
xor \U$13672 ( \13730 , \13656 , \13729 );
buf \U$13673 ( \13731 , RIc0d8c08_47);
buf \U$13674 ( \13732 , RIc0d9dd8_85);
xor \U$13675 ( \13733 , \13731 , \13732 );
buf \U$13676 ( \13734 , \13733 );
buf \U$13677 ( \13735 , \13734 );
not \U$13678 ( \13736 , \13735 );
buf \U$13681 ( \13737 , \2393 );
buf \U$13682 ( \13738 , \13737 );
not \U$13683 ( \13739 , \13738 );
or \U$13684 ( \13740 , \13736 , \13739 );
buf \U$13685 ( \13741 , \2960 );
buf \U$13686 ( \13742 , RIc0d8b90_46);
buf \U$13687 ( \13743 , RIc0d9dd8_85);
xor \U$13688 ( \13744 , \13742 , \13743 );
buf \U$13689 ( \13745 , \13744 );
buf \U$13690 ( \13746 , \13745 );
nand \U$13691 ( \13747 , \13741 , \13746 );
buf \U$13692 ( \13748 , \13747 );
buf \U$13693 ( \13749 , \13748 );
nand \U$13694 ( \13750 , \13740 , \13749 );
buf \U$13695 ( \13751 , \13750 );
buf \U$13696 ( \13752 , \13751 );
xor \U$13697 ( \13753 , RIc0d9bf8_81, RIc0d8de8_51);
buf \U$13698 ( \13754 , \13753 );
not \U$13699 ( \13755 , \13754 );
buf \U$13700 ( \13756 , \2766 );
not \U$13701 ( \13757 , \13756 );
or \U$13702 ( \13758 , \13755 , \13757 );
buf \U$13703 ( \13759 , \1078 );
buf \U$13704 ( \13760 , RIc0d8d70_50);
buf \U$13705 ( \13761 , RIc0d9bf8_81);
xor \U$13706 ( \13762 , \13760 , \13761 );
buf \U$13707 ( \13763 , \13762 );
buf \U$13708 ( \13764 , \13763 );
nand \U$13709 ( \13765 , \13759 , \13764 );
buf \U$13710 ( \13766 , \13765 );
buf \U$13711 ( \13767 , \13766 );
nand \U$13712 ( \13768 , \13758 , \13767 );
buf \U$13713 ( \13769 , \13768 );
buf \U$13714 ( \13770 , \13769 );
xor \U$13715 ( \13771 , \13752 , \13770 );
buf \U$13716 ( \13772 , RIc0d7b28_11);
buf \U$13717 ( \13773 , RIc0daeb8_121);
xor \U$13718 ( \13774 , \13772 , \13773 );
buf \U$13719 ( \13775 , \13774 );
buf \U$13720 ( \13776 , \13775 );
not \U$13721 ( \13777 , \13776 );
buf \U$13722 ( \13778 , \13310 );
not \U$13723 ( \13779 , \13778 );
or \U$13724 ( \13780 , \13777 , \13779 );
buf \U$13725 ( \13781 , \13314 );
buf \U$13726 ( \13782 , RIc0daeb8_121);
buf \U$13727 ( \13783 , RIc0d7ab0_10);
xor \U$13728 ( \13784 , \13782 , \13783 );
buf \U$13729 ( \13785 , \13784 );
buf \U$13730 ( \13786 , \13785 );
nand \U$13731 ( \13787 , \13781 , \13786 );
buf \U$13732 ( \13788 , \13787 );
buf \U$13733 ( \13789 , \13788 );
nand \U$13734 ( \13790 , \13780 , \13789 );
buf \U$13735 ( \13791 , \13790 );
buf \U$13736 ( \13792 , \13791 );
and \U$13737 ( \13793 , \13771 , \13792 );
and \U$13738 ( \13794 , \13752 , \13770 );
or \U$13739 ( \13795 , \13793 , \13794 );
buf \U$13740 ( \13796 , \13795 );
buf \U$13741 ( \13797 , \13796 );
and \U$13742 ( \13798 , \13730 , \13797 );
and \U$13743 ( \13799 , \13656 , \13729 );
or \U$13744 ( \13800 , \13798 , \13799 );
buf \U$13745 ( \13801 , \13800 );
buf \U$13746 ( \13802 , \13801 );
buf \U$13747 ( \13803 , \13343 );
not \U$13748 ( \13804 , \13803 );
buf \U$13749 ( \13805 , \13356 );
not \U$13750 ( \13806 , \13805 );
and \U$13751 ( \13807 , \13804 , \13806 );
buf \U$13752 ( \13808 , \13343 );
buf \U$13753 ( \13809 , \13356 );
and \U$13754 ( \13810 , \13808 , \13809 );
nor \U$13755 ( \13811 , \13807 , \13810 );
buf \U$13756 ( \13812 , \13811 );
buf \U$13757 ( \13813 , \13812 );
not \U$13758 ( \13814 , \13813 );
buf \U$13759 ( \13815 , \13814 );
buf \U$13760 ( \13816 , \13815 );
not \U$13761 ( \13817 , \13816 );
buf \U$13762 ( \13818 , \685 );
buf \U$13763 ( \13819 , RIc0d9400_64);
and \U$13764 ( \13820 , \13818 , \13819 );
buf \U$13765 ( \13821 , \13820 );
buf \U$13766 ( \13822 , \13821 );
not \U$13767 ( \13823 , \13822 );
buf \U$13768 ( \13824 , RIc0d9298_61);
buf \U$13769 ( \13825 , RIc0d9748_71);
xor \U$13770 ( \13826 , \13824 , \13825 );
buf \U$13771 ( \13827 , \13826 );
buf \U$13772 ( \13828 , \13827 );
not \U$13773 ( \13829 , \13828 );
buf \U$13774 ( \13830 , \12676 );
not \U$13775 ( \13831 , \13830 );
or \U$13776 ( \13832 , \13829 , \13831 );
buf \U$13777 ( \13833 , \12683 );
buf \U$13778 ( \13834 , RIc0d9220_60);
buf \U$13779 ( \13835 , RIc0d9748_71);
xor \U$13780 ( \13836 , \13834 , \13835 );
buf \U$13781 ( \13837 , \13836 );
buf \U$13782 ( \13838 , \13837 );
nand \U$13783 ( \13839 , \13833 , \13838 );
buf \U$13784 ( \13840 , \13839 );
buf \U$13785 ( \13841 , \13840 );
nand \U$13786 ( \13842 , \13832 , \13841 );
buf \U$13787 ( \13843 , \13842 );
buf \U$13788 ( \13844 , \13843 );
not \U$13789 ( \13845 , \13844 );
or \U$13790 ( \13846 , \13823 , \13845 );
buf \U$13791 ( \13847 , \13821 );
buf \U$13792 ( \13848 , \13843 );
or \U$13793 ( \13849 , \13847 , \13848 );
buf \U$13794 ( \13850 , RIc0d8758_37);
buf \U$13795 ( \13851 , RIc0da288_95);
xor \U$13796 ( \13852 , \13850 , \13851 );
buf \U$13797 ( \13853 , \13852 );
buf \U$13798 ( \13854 , \13853 );
not \U$13799 ( \13855 , \13854 );
buf \U$13800 ( \13856 , \326 );
buf \U$13801 ( \13857 , \320 );
buf \U$13802 ( \13858 , \314 );
and \U$13803 ( \13859 , \13856 , \13857 , \13858 );
buf \U$13804 ( \13860 , \13859 );
buf \U$13805 ( \13861 , \13860 );
not \U$13806 ( \13862 , \13861 );
or \U$13807 ( \13863 , \13855 , \13862 );
buf \U$13808 ( \13864 , RIc0d86e0_36);
buf \U$13809 ( \13865 , RIc0da288_95);
xnor \U$13810 ( \13866 , \13864 , \13865 );
buf \U$13811 ( \13867 , \13866 );
buf \U$13812 ( \13868 , \13867 );
not \U$13813 ( \13869 , \13868 );
buf \U$13814 ( \13870 , RIc0da300_96);
buf \U$13815 ( \13871 , RIc0da378_97);
xor \U$13816 ( \13872 , \13870 , \13871 );
buf \U$13817 ( \13873 , \13872 );
buf \U$13818 ( \13874 , \13873 );
nand \U$13819 ( \13875 , \13869 , \13874 );
buf \U$13820 ( \13876 , \13875 );
buf \U$13821 ( \13877 , \13876 );
nand \U$13822 ( \13878 , \13863 , \13877 );
buf \U$13823 ( \13879 , \13878 );
buf \U$13824 ( \13880 , \13879 );
nand \U$13825 ( \13881 , \13849 , \13880 );
buf \U$13826 ( \13882 , \13881 );
buf \U$13827 ( \13883 , \13882 );
nand \U$13828 ( \13884 , \13846 , \13883 );
buf \U$13829 ( \13885 , \13884 );
buf \U$13830 ( \13886 , \13885 );
not \U$13831 ( \13887 , \13886 );
or \U$13832 ( \13888 , \13817 , \13887 );
buf \U$13833 ( \13889 , \13885 );
buf \U$13834 ( \13890 , \13815 );
or \U$13835 ( \13891 , \13889 , \13890 );
buf \U$13836 ( \13892 , RIc0d88c0_40);
buf \U$13837 ( \13893 , RIc0da0a8_91);
xor \U$13838 ( \13894 , \13892 , \13893 );
buf \U$13839 ( \13895 , \13894 );
buf \U$13840 ( \13896 , \13895 );
not \U$13841 ( \13897 , \13896 );
buf \U$13842 ( \13898 , \533 );
not \U$13843 ( \13899 , \13898 );
or \U$13844 ( \13900 , \13897 , \13899 );
buf \U$13845 ( \13901 , \530 );
buf \U$13846 ( \13902 , RIc0d8938_41);
buf \U$13847 ( \13903 , RIc0da0a8_91);
xor \U$13848 ( \13904 , \13902 , \13903 );
buf \U$13849 ( \13905 , \13904 );
buf \U$13850 ( \13906 , \13905 );
buf \U$13851 ( \13907 , \517 );
nand \U$13852 ( \13908 , \13901 , \13906 , \13907 );
buf \U$13853 ( \13909 , \13908 );
buf \U$13854 ( \13910 , \13909 );
nand \U$13855 ( \13911 , \13900 , \13910 );
buf \U$13856 ( \13912 , \13911 );
buf \U$13857 ( \13913 , \13912 );
not \U$13858 ( \13914 , \13913 );
buf \U$13859 ( \13915 , \13914 );
buf \U$13860 ( \13916 , \13915 );
not \U$13861 ( \13917 , \13916 );
xor \U$13862 ( \13918 , RIc0da738_105, RIc0d82a8_27);
buf \U$13863 ( \13919 , \13918 );
not \U$13864 ( \13920 , \13919 );
buf \U$13865 ( \13921 , \12736 );
not \U$13866 ( \13922 , \13921 );
or \U$13867 ( \13923 , \13920 , \13922 );
buf \U$13868 ( \13924 , \12744 );
buf \U$13869 ( \13925 , RIc0d8230_26);
buf \U$13870 ( \13926 , RIc0da738_105);
xor \U$13871 ( \13927 , \13925 , \13926 );
buf \U$13872 ( \13928 , \13927 );
buf \U$13873 ( \13929 , \13928 );
nand \U$13874 ( \13930 , \13924 , \13929 );
buf \U$13875 ( \13931 , \13930 );
buf \U$13876 ( \13932 , \13931 );
nand \U$13877 ( \13933 , \13923 , \13932 );
buf \U$13878 ( \13934 , \13933 );
buf \U$13879 ( \13935 , \13934 );
not \U$13880 ( \13936 , \13935 );
buf \U$13881 ( \13937 , \13936 );
buf \U$13882 ( \13938 , \13937 );
not \U$13883 ( \13939 , \13938 );
or \U$13884 ( \13940 , \13917 , \13939 );
buf \U$13885 ( \13941 , RIc0dadc8_119);
buf \U$13886 ( \13942 , RIc0d7c18_13);
xor \U$13887 ( \13943 , \13941 , \13942 );
buf \U$13888 ( \13944 , \13943 );
buf \U$13889 ( \13945 , \13944 );
not \U$13890 ( \13946 , \13945 );
buf \U$13891 ( \13947 , \13178 );
not \U$13892 ( \13948 , \13947 );
buf \U$13893 ( \13949 , \13948 );
buf \U$13894 ( \13950 , \13949 );
not \U$13895 ( \13951 , \13950 );
or \U$13896 ( \13952 , \13946 , \13951 );
buf \U$13899 ( \13953 , \13005 );
buf \U$13900 ( \13954 , \13953 );
xor \U$13901 ( \13955 , RIc0dadc8_119, RIc0d7ba0_12);
buf \U$13902 ( \13956 , \13955 );
nand \U$13903 ( \13957 , \13954 , \13956 );
buf \U$13904 ( \13958 , \13957 );
buf \U$13905 ( \13959 , \13958 );
nand \U$13906 ( \13960 , \13952 , \13959 );
buf \U$13907 ( \13961 , \13960 );
buf \U$13908 ( \13962 , \13961 );
nand \U$13909 ( \13963 , \13940 , \13962 );
buf \U$13910 ( \13964 , \13963 );
buf \U$13911 ( \13965 , \13964 );
buf \U$13912 ( \13966 , \13937 );
not \U$13913 ( \13967 , \13966 );
buf \U$13914 ( \13968 , \13912 );
nand \U$13915 ( \13969 , \13967 , \13968 );
buf \U$13916 ( \13970 , \13969 );
buf \U$13917 ( \13971 , \13970 );
nand \U$13918 ( \13972 , \13965 , \13971 );
buf \U$13919 ( \13973 , \13972 );
buf \U$13920 ( \13974 , \13973 );
nand \U$13921 ( \13975 , \13891 , \13974 );
buf \U$13922 ( \13976 , \13975 );
buf \U$13923 ( \13977 , \13976 );
nand \U$13924 ( \13978 , \13888 , \13977 );
buf \U$13925 ( \13979 , \13978 );
buf \U$13926 ( \13980 , \13979 );
xor \U$13927 ( \13981 , \13802 , \13980 );
buf \U$13928 ( \13982 , RIc0d90b8_57);
buf \U$13929 ( \13983 , RIc0d9928_75);
xor \U$13930 ( \13984 , \13982 , \13983 );
buf \U$13931 ( \13985 , \13984 );
buf \U$13932 ( \13986 , \13985 );
not \U$13933 ( \13987 , \13986 );
buf \U$13934 ( \13988 , \1120 );
buf \U$13935 ( \13989 , \1105 );
and \U$13936 ( \13990 , \13988 , \13989 );
buf \U$13937 ( \13991 , \13990 );
buf \U$13938 ( \13992 , \13991 );
not \U$13939 ( \13993 , \13992 );
or \U$13940 ( \13994 , \13987 , \13993 );
buf \U$13941 ( \13995 , RIc0d99a0_76);
buf \U$13942 ( \13996 , RIc0d9a18_77);
xor \U$13943 ( \13997 , \13995 , \13996 );
buf \U$13944 ( \13998 , \13997 );
buf \U$13945 ( \13999 , \13998 );
buf \U$13946 ( \14000 , RIc0d9040_56);
buf \U$13947 ( \14001 , RIc0d9928_75);
xor \U$13948 ( \14002 , \14000 , \14001 );
buf \U$13949 ( \14003 , \14002 );
buf \U$13950 ( \14004 , \14003 );
nand \U$13951 ( \14005 , \13999 , \14004 );
buf \U$13952 ( \14006 , \14005 );
buf \U$13953 ( \14007 , \14006 );
nand \U$13954 ( \14008 , \13994 , \14007 );
buf \U$13955 ( \14009 , \14008 );
buf \U$13956 ( \14010 , \14009 );
not \U$13957 ( \14011 , \14010 );
buf \U$13958 ( \14012 , \14011 );
buf \U$13959 ( \14013 , \14012 );
not \U$13960 ( \14014 , \14013 );
xor \U$13961 ( \14015 , RIc0d9ec8_87, RIc0d8b18_45);
buf \U$13962 ( \14016 , \14015 );
not \U$13963 ( \14017 , \14016 );
buf \U$13964 ( \14018 , \4527 );
not \U$13965 ( \14019 , \14018 );
or \U$13966 ( \14020 , \14017 , \14019 );
buf \U$13967 ( \14021 , \3631 );
xor \U$13968 ( \14022 , RIc0d9ec8_87, RIc0d8aa0_44);
buf \U$13969 ( \14023 , \14022 );
nand \U$13970 ( \14024 , \14021 , \14023 );
buf \U$13971 ( \14025 , \14024 );
buf \U$13972 ( \14026 , \14025 );
nand \U$13973 ( \14027 , \14020 , \14026 );
buf \U$13974 ( \14028 , \14027 );
buf \U$13975 ( \14029 , \14028 );
not \U$13976 ( \14030 , \14029 );
buf \U$13977 ( \14031 , \14030 );
buf \U$13978 ( \14032 , \14031 );
not \U$13979 ( \14033 , \14032 );
or \U$13980 ( \14034 , \14014 , \14033 );
buf \U$13981 ( \14035 , RIc0d8488_31);
buf \U$13982 ( \14036 , RIc0da558_101);
xor \U$13983 ( \14037 , \14035 , \14036 );
buf \U$13984 ( \14038 , \14037 );
buf \U$13985 ( \14039 , \14038 );
not \U$13986 ( \14040 , \14039 );
buf \U$13987 ( \14041 , \12833 );
not \U$13988 ( \14042 , \14041 );
or \U$13989 ( \14043 , \14040 , \14042 );
buf \U$13990 ( \14044 , \12839 );
buf \U$13991 ( \14045 , RIc0d8410_30);
buf \U$13992 ( \14046 , RIc0da558_101);
xor \U$13993 ( \14047 , \14045 , \14046 );
buf \U$13994 ( \14048 , \14047 );
buf \U$13995 ( \14049 , \14048 );
nand \U$13996 ( \14050 , \14044 , \14049 );
buf \U$13997 ( \14051 , \14050 );
buf \U$13998 ( \14052 , \14051 );
nand \U$13999 ( \14053 , \14043 , \14052 );
buf \U$14000 ( \14054 , \14053 );
buf \U$14001 ( \14055 , \14054 );
nand \U$14002 ( \14056 , \14034 , \14055 );
buf \U$14003 ( \14057 , \14056 );
buf \U$14004 ( \14058 , \14057 );
buf \U$14005 ( \14059 , \14028 );
buf \U$14006 ( \14060 , \14009 );
nand \U$14007 ( \14061 , \14059 , \14060 );
buf \U$14008 ( \14062 , \14061 );
buf \U$14009 ( \14063 , \14062 );
nand \U$14010 ( \14064 , \14058 , \14063 );
buf \U$14011 ( \14065 , \14064 );
buf \U$14012 ( \14066 , \14065 );
buf \U$14013 ( \14067 , RIc0d91a8_59);
buf \U$14014 ( \14068 , RIc0d9838_73);
xor \U$14015 ( \14069 , \14067 , \14068 );
buf \U$14016 ( \14070 , \14069 );
buf \U$14017 ( \14071 , \14070 );
not \U$14018 ( \14072 , \14071 );
buf \U$14019 ( \14073 , \773 );
not \U$14020 ( \14074 , \14073 );
buf \U$14021 ( \14075 , \14074 );
buf \U$14022 ( \14076 , \14075 );
not \U$14023 ( \14077 , \14076 );
or \U$14024 ( \14078 , \14072 , \14077 );
buf \U$14025 ( \14079 , \1856 );
buf \U$14026 ( \14080 , RIc0d9130_58);
buf \U$14027 ( \14081 , RIc0d9838_73);
xor \U$14028 ( \14082 , \14080 , \14081 );
buf \U$14029 ( \14083 , \14082 );
buf \U$14030 ( \14084 , \14083 );
nand \U$14031 ( \14085 , \14079 , \14084 );
buf \U$14032 ( \14086 , \14085 );
buf \U$14033 ( \14087 , \14086 );
nand \U$14034 ( \14088 , \14078 , \14087 );
buf \U$14035 ( \14089 , \14088 );
not \U$14036 ( \14090 , \14089 );
buf \U$14037 ( \14091 , RIc0d7fd8_21);
buf \U$14038 ( \14092 , RIc0daa08_111);
xor \U$14039 ( \14093 , \14091 , \14092 );
buf \U$14040 ( \14094 , \14093 );
buf \U$14041 ( \14095 , \14094 );
not \U$14042 ( \14096 , \14095 );
buf \U$14043 ( \14097 , \12525 );
buf \U$14044 ( \14098 , \12517 );
and \U$14045 ( \14099 , \14097 , \14098 );
buf \U$14046 ( \14100 , \14099 );
buf \U$14047 ( \14101 , \14100 );
not \U$14048 ( \14102 , \14101 );
or \U$14049 ( \14103 , \14096 , \14102 );
buf \U$14050 ( \14104 , \12540 );
not \U$14051 ( \14105 , \14104 );
buf \U$14052 ( \14106 , \14105 );
buf \U$14053 ( \14107 , \14106 );
buf \U$14054 ( \14108 , RIc0d7f60_20);
buf \U$14055 ( \14109 , RIc0daa08_111);
xor \U$14056 ( \14110 , \14108 , \14109 );
buf \U$14057 ( \14111 , \14110 );
buf \U$14058 ( \14112 , \14111 );
nand \U$14059 ( \14113 , \14107 , \14112 );
buf \U$14060 ( \14114 , \14113 );
buf \U$14061 ( \14115 , \14114 );
nand \U$14062 ( \14116 , \14103 , \14115 );
buf \U$14063 ( \14117 , \14116 );
not \U$14064 ( \14118 , \14117 );
or \U$14065 ( \14119 , \14090 , \14118 );
buf \U$14066 ( \14120 , \14117 );
not \U$14067 ( \14121 , \14120 );
buf \U$14068 ( \14122 , \14121 );
not \U$14069 ( \14123 , \14122 );
buf \U$14070 ( \14124 , \14089 );
not \U$14071 ( \14125 , \14124 );
buf \U$14072 ( \14126 , \14125 );
not \U$14073 ( \14127 , \14126 );
or \U$14074 ( \14128 , \14123 , \14127 );
buf \U$14075 ( \14129 , RIc0d8578_33);
buf \U$14076 ( \14130 , RIc0da468_99);
xor \U$14077 ( \14131 , \14129 , \14130 );
buf \U$14078 ( \14132 , \14131 );
buf \U$14079 ( \14133 , \14132 );
not \U$14080 ( \14134 , \14133 );
buf \U$14081 ( \14135 , \12578 );
not \U$14082 ( \14136 , \14135 );
or \U$14083 ( \14137 , \14134 , \14136 );
buf \U$14084 ( \14138 , \2198 );
not \U$14085 ( \14139 , \14138 );
buf \U$14086 ( \14140 , \14139 );
buf \U$14087 ( \14141 , \14140 );
buf \U$14088 ( \14142 , RIc0d8500_32);
buf \U$14089 ( \14143 , RIc0da468_99);
xor \U$14090 ( \14144 , \14142 , \14143 );
buf \U$14091 ( \14145 , \14144 );
buf \U$14092 ( \14146 , \14145 );
nand \U$14093 ( \14147 , \14141 , \14146 );
buf \U$14094 ( \14148 , \14147 );
buf \U$14095 ( \14149 , \14148 );
nand \U$14096 ( \14150 , \14137 , \14149 );
buf \U$14097 ( \14151 , \14150 );
nand \U$14098 ( \14152 , \14128 , \14151 );
nand \U$14099 ( \14153 , \14119 , \14152 );
buf \U$14100 ( \14154 , \14153 );
xor \U$14101 ( \14155 , \14066 , \14154 );
buf \U$14102 ( \14156 , RIc0d9388_63);
buf \U$14103 ( \14157 , RIc0d9658_69);
xor \U$14104 ( \14158 , \14156 , \14157 );
buf \U$14105 ( \14159 , \14158 );
buf \U$14106 ( \14160 , \14159 );
not \U$14107 ( \14161 , \14160 );
buf \U$14108 ( \14162 , \13332 );
not \U$14109 ( \14163 , \14162 );
or \U$14110 ( \14164 , \14161 , \14163 );
buf \U$14111 ( \14165 , \284 );
buf \U$14112 ( \14166 , \13327 );
nand \U$14113 ( \14167 , \14165 , \14166 );
buf \U$14114 ( \14168 , \14167 );
buf \U$14115 ( \14169 , \14168 );
nand \U$14116 ( \14170 , \14164 , \14169 );
buf \U$14117 ( \14171 , \14170 );
buf \U$14118 ( \14172 , \14171 );
xor \U$14119 ( \14173 , RIc0dabe8_115, RIc0d7df8_17);
buf \U$14120 ( \14174 , \14173 );
not \U$14121 ( \14175 , \14174 );
buf \U$14122 ( \14176 , RIc0dac60_116);
buf \U$14123 ( \14177 , RIc0dacd8_117);
xnor \U$14124 ( \14178 , \14176 , \14177 );
buf \U$14125 ( \14179 , \14178 );
buf \U$14126 ( \14180 , \14179 );
buf \U$14127 ( \14181 , \12293 );
nand \U$14128 ( \14182 , \14180 , \14181 );
buf \U$14129 ( \14183 , \14182 );
buf \U$14130 ( \14184 , \14183 );
not \U$14131 ( \14185 , \14184 );
buf \U$14132 ( \14186 , \14185 );
buf \U$14133 ( \14187 , \14186 );
not \U$14134 ( \14188 , \14187 );
or \U$14135 ( \14189 , \14175 , \14188 );
buf \U$14136 ( \14190 , \12303 );
xor \U$14137 ( \14191 , RIc0dabe8_115, RIc0d7d80_16);
buf \U$14138 ( \14192 , \14191 );
nand \U$14139 ( \14193 , \14190 , \14192 );
buf \U$14140 ( \14194 , \14193 );
buf \U$14141 ( \14195 , \14194 );
nand \U$14142 ( \14196 , \14189 , \14195 );
buf \U$14143 ( \14197 , \14196 );
buf \U$14144 ( \14198 , \14197 );
xor \U$14145 ( \14199 , \14172 , \14198 );
xor \U$14146 ( \14200 , RIc0da918_109, RIc0d80c8_23);
buf \U$14147 ( \14201 , \14200 );
not \U$14148 ( \14202 , \14201 );
buf \U$14149 ( \14203 , \13411 );
buf \U$14150 ( \14204 , \13413 );
nand \U$14151 ( \14205 , \14203 , \14204 );
buf \U$14152 ( \14206 , \14205 );
buf \U$14155 ( \14207 , \14206 );
buf \U$14156 ( \14208 , \14207 );
not \U$14157 ( \14209 , \14208 );
buf \U$14158 ( \14210 , \14209 );
buf \U$14159 ( \14211 , \14210 );
not \U$14160 ( \14212 , \14211 );
or \U$14161 ( \14213 , \14202 , \14212 );
buf \U$14162 ( \14214 , \13411 );
not \U$14163 ( \14215 , \14214 );
buf \U$14164 ( \14216 , \14215 );
buf \U$14165 ( \14217 , \14216 );
buf \U$14166 ( \14218 , RIc0da918_109);
buf \U$14167 ( \14219 , RIc0d8050_22);
xor \U$14168 ( \14220 , \14218 , \14219 );
buf \U$14169 ( \14221 , \14220 );
buf \U$14170 ( \14222 , \14221 );
nand \U$14171 ( \14223 , \14217 , \14222 );
buf \U$14172 ( \14224 , \14223 );
buf \U$14173 ( \14225 , \14224 );
nand \U$14174 ( \14226 , \14213 , \14225 );
buf \U$14175 ( \14227 , \14226 );
buf \U$14176 ( \14228 , \14227 );
and \U$14177 ( \14229 , \14199 , \14228 );
and \U$14178 ( \14230 , \14172 , \14198 );
or \U$14179 ( \14231 , \14229 , \14230 );
buf \U$14180 ( \14232 , \14231 );
buf \U$14181 ( \14233 , \14232 );
and \U$14182 ( \14234 , \14155 , \14233 );
and \U$14183 ( \14235 , \14066 , \14154 );
or \U$14184 ( \14236 , \14234 , \14235 );
buf \U$14185 ( \14237 , \14236 );
buf \U$14186 ( \14238 , \14237 );
and \U$14187 ( \14239 , \13981 , \14238 );
and \U$14188 ( \14240 , \13802 , \13980 );
or \U$14189 ( \14241 , \14239 , \14240 );
buf \U$14190 ( \14242 , \14241 );
buf \U$14191 ( \14243 , \14242 );
xor \U$14192 ( \14244 , \13592 , \14243 );
buf \U$14193 ( \14245 , \14244 );
buf \U$14194 ( \14246 , \14245 );
xor \U$14195 ( \14247 , \13137 , \14246 );
buf \U$14196 ( \14248 , RIc0d8398_29);
buf \U$14197 ( \14249 , RIc0da558_101);
xor \U$14198 ( \14250 , \14248 , \14249 );
buf \U$14199 ( \14251 , \14250 );
buf \U$14200 ( \14252 , \14251 );
not \U$14201 ( \14253 , \14252 );
buf \U$14202 ( \14254 , \4042 );
not \U$14203 ( \14255 , \14254 );
or \U$14204 ( \14256 , \14253 , \14255 );
buf \U$14205 ( \14257 , \12839 );
buf \U$14206 ( \14258 , \12828 );
nand \U$14207 ( \14259 , \14257 , \14258 );
buf \U$14208 ( \14260 , \14259 );
buf \U$14209 ( \14261 , \14260 );
nand \U$14210 ( \14262 , \14256 , \14261 );
buf \U$14211 ( \14263 , \14262 );
buf \U$14212 ( \14264 , RIc0d7948_7);
buf \U$14213 ( \14265 , RIc0dafa8_123);
xor \U$14214 ( \14266 , \14264 , \14265 );
buf \U$14215 ( \14267 , \14266 );
buf \U$14216 ( \14268 , \14267 );
not \U$14217 ( \14269 , \14268 );
buf \U$14218 ( \14270 , \12870 );
not \U$14219 ( \14271 , \14270 );
or \U$14220 ( \14272 , \14269 , \14271 );
buf \U$14221 ( \14273 , \12877 );
not \U$14222 ( \14274 , \14273 );
buf \U$14223 ( \14275 , \14274 );
buf \U$14224 ( \14276 , \14275 );
not \U$14225 ( \14277 , \14276 );
buf \U$14226 ( \14278 , \14277 );
buf \U$14227 ( \14279 , \14278 );
buf \U$14228 ( \14280 , \12855 );
nand \U$14229 ( \14281 , \14279 , \14280 );
buf \U$14230 ( \14282 , \14281 );
buf \U$14231 ( \14283 , \14282 );
nand \U$14232 ( \14284 , \14272 , \14283 );
buf \U$14233 ( \14285 , \14284 );
xor \U$14234 ( \14286 , \14263 , \14285 );
buf \U$14235 ( \14287 , RIc0d9928_75);
buf \U$14236 ( \14288 , RIc0d8fc8_55);
xor \U$14237 ( \14289 , \14287 , \14288 );
buf \U$14238 ( \14290 , \14289 );
buf \U$14239 ( \14291 , \14290 );
not \U$14240 ( \14292 , \14291 );
buf \U$14241 ( \14293 , \2358 );
not \U$14242 ( \14294 , \14293 );
or \U$14243 ( \14295 , \14292 , \14294 );
buf \U$14244 ( \14296 , \1143 );
buf \U$14245 ( \14297 , \13378 );
nand \U$14246 ( \14298 , \14296 , \14297 );
buf \U$14247 ( \14299 , \14298 );
buf \U$14248 ( \14300 , \14299 );
nand \U$14249 ( \14301 , \14295 , \14300 );
buf \U$14250 ( \14302 , \14301 );
buf \U$14251 ( \14303 , \14302 );
not \U$14252 ( \14304 , \14303 );
buf \U$14253 ( \14305 , \14304 );
and \U$14254 ( \14306 , \14286 , \14305 );
not \U$14255 ( \14307 , \14286 );
and \U$14256 ( \14308 , \14307 , \14302 );
nor \U$14257 ( \14309 , \14306 , \14308 );
buf \U$14258 ( \14310 , \14309 );
not \U$14259 ( \14311 , \14310 );
buf \U$14260 ( \14312 , RIc0d8a28_43);
buf \U$14261 ( \14313 , RIc0d9ec8_87);
xor \U$14262 ( \14314 , \14312 , \14313 );
buf \U$14263 ( \14315 , \14314 );
buf \U$14264 ( \14316 , \14315 );
not \U$14265 ( \14317 , \14316 );
buf \U$14266 ( \14318 , \631 );
not \U$14267 ( \14319 , \14318 );
buf \U$14268 ( \14320 , \606 );
nand \U$14269 ( \14321 , \14319 , \14320 );
buf \U$14270 ( \14322 , \14321 );
buf \U$14271 ( \14323 , \14322 );
not \U$14272 ( \14324 , \14323 );
buf \U$14273 ( \14325 , \14324 );
buf \U$14274 ( \14326 , \14325 );
not \U$14275 ( \14327 , \14326 );
or \U$14276 ( \14328 , \14317 , \14327 );
buf \U$14277 ( \14329 , \634 );
not \U$14278 ( \14330 , \14329 );
buf \U$14279 ( \14331 , \14330 );
buf \U$14280 ( \14332 , \14331 );
buf \U$14281 ( \14333 , \12622 );
nand \U$14282 ( \14334 , \14332 , \14333 );
buf \U$14283 ( \14335 , \14334 );
buf \U$14284 ( \14336 , \14335 );
nand \U$14285 ( \14337 , \14328 , \14336 );
buf \U$14286 ( \14338 , \14337 );
buf \U$14287 ( \14339 , \14338 );
buf \U$14288 ( \14340 , RIc0daa08_111);
buf \U$14289 ( \14341 , RIc0d7ee8_19);
xor \U$14290 ( \14342 , \14340 , \14341 );
buf \U$14291 ( \14343 , \14342 );
buf \U$14292 ( \14344 , \14343 );
not \U$14293 ( \14345 , \14344 );
buf \U$14296 ( \14346 , \12528 );
buf \U$14297 ( \14347 , \14346 );
not \U$14298 ( \14348 , \14347 );
or \U$14299 ( \14349 , \14345 , \14348 );
buf \U$14300 ( \14350 , \12525 );
not \U$14301 ( \14351 , \14350 );
buf \U$14302 ( \14352 , \14351 );
buf \U$14305 ( \14353 , \14352 );
buf \U$14306 ( \14354 , \14353 );
buf \U$14307 ( \14355 , \12534 );
nand \U$14308 ( \14356 , \14354 , \14355 );
buf \U$14309 ( \14357 , \14356 );
buf \U$14310 ( \14358 , \14357 );
nand \U$14311 ( \14359 , \14349 , \14358 );
buf \U$14312 ( \14360 , \14359 );
buf \U$14313 ( \14361 , \14360 );
xor \U$14314 ( \14362 , \14339 , \14361 );
buf \U$14315 ( \14363 , RIc0d9a18_77);
buf \U$14316 ( \14364 , RIc0d8ed8_53);
xor \U$14317 ( \14365 , \14363 , \14364 );
buf \U$14318 ( \14366 , \14365 );
buf \U$14319 ( \14367 , \14366 );
not \U$14320 ( \14368 , \14367 );
buf \U$14321 ( \14369 , \1431 );
not \U$14322 ( \14370 , \14369 );
or \U$14323 ( \14371 , \14368 , \14370 );
buf \U$14324 ( \14372 , \1193 );
not \U$14325 ( \14373 , \14372 );
buf \U$14326 ( \14374 , \14373 );
buf \U$14327 ( \14375 , \14374 );
buf \U$14328 ( \14376 , \12761 );
nand \U$14329 ( \14377 , \14375 , \14376 );
buf \U$14330 ( \14378 , \14377 );
buf \U$14331 ( \14379 , \14378 );
nand \U$14332 ( \14380 , \14371 , \14379 );
buf \U$14333 ( \14381 , \14380 );
buf \U$14334 ( \14382 , \14381 );
xor \U$14335 ( \14383 , \14362 , \14382 );
buf \U$14336 ( \14384 , \14383 );
buf \U$14337 ( \14385 , \14384 );
not \U$14338 ( \14386 , \14385 );
or \U$14339 ( \14387 , \14311 , \14386 );
buf \U$14340 ( \14388 , \14384 );
buf \U$14341 ( \14389 , \14309 );
or \U$14342 ( \14390 , \14388 , \14389 );
nand \U$14343 ( \14391 , \14387 , \14390 );
buf \U$14344 ( \14392 , \14391 );
buf \U$14345 ( \14393 , \14392 );
xor \U$14346 ( \14394 , RIc0daaf8_113, RIc0d7df8_17);
buf \U$14347 ( \14395 , \14394 );
not \U$14348 ( \14396 , \14395 );
buf \U$14349 ( \14397 , \12402 );
not \U$14350 ( \14398 , \14397 );
or \U$14351 ( \14399 , \14396 , \14398 );
buf \U$14352 ( \14400 , \12409 );
not \U$14353 ( \14401 , \14400 );
buf \U$14354 ( \14402 , \14401 );
buf \U$14355 ( \14403 , \14402 );
not \U$14356 ( \14404 , \14403 );
buf \U$14357 ( \14405 , \14404 );
buf \U$14358 ( \14406 , \14405 );
buf \U$14359 ( \14407 , \12378 );
nand \U$14360 ( \14408 , \14406 , \14407 );
buf \U$14361 ( \14409 , \14408 );
buf \U$14362 ( \14410 , \14409 );
nand \U$14363 ( \14411 , \14399 , \14410 );
buf \U$14364 ( \14412 , \14411 );
buf \U$14365 ( \14413 , \14412 );
xor \U$14366 ( \14414 , RIc0da468_99, RIc0d8488_31);
buf \U$14367 ( \14415 , \14414 );
not \U$14368 ( \14416 , \14415 );
buf \U$14369 ( \14417 , \2207 );
not \U$14370 ( \14418 , \14417 );
buf \U$14371 ( \14419 , \14418 );
buf \U$14372 ( \14420 , \14419 );
not \U$14373 ( \14421 , \14420 );
or \U$14374 ( \14422 , \14416 , \14421 );
buf \U$14375 ( \14423 , \12584 );
buf \U$14376 ( \14424 , \12572 );
nand \U$14377 ( \14425 , \14423 , \14424 );
buf \U$14378 ( \14426 , \14425 );
buf \U$14379 ( \14427 , \14426 );
nand \U$14380 ( \14428 , \14422 , \14427 );
buf \U$14381 ( \14429 , \14428 );
buf \U$14382 ( \14430 , \14429 );
xor \U$14383 ( \14431 , \14413 , \14430 );
buf \U$14384 ( \14432 , \14431 );
xor \U$14385 ( \14433 , RIc0d9bf8_81, RIc0d8cf8_49);
buf \U$14386 ( \14434 , \14433 );
not \U$14387 ( \14435 , \14434 );
buf \U$14388 ( \14436 , \1063 );
not \U$14389 ( \14437 , \14436 );
or \U$14390 ( \14438 , \14435 , \14437 );
buf \U$14391 ( \14439 , \1078 );
buf \U$14392 ( \14440 , \13070 );
nand \U$14393 ( \14441 , \14439 , \14440 );
buf \U$14394 ( \14442 , \14441 );
buf \U$14395 ( \14443 , \14442 );
nand \U$14396 ( \14444 , \14438 , \14443 );
buf \U$14397 ( \14445 , \14444 );
xnor \U$14398 ( \14446 , \14432 , \14445 );
buf \U$14399 ( \14447 , \14446 );
not \U$14400 ( \14448 , \14447 );
buf \U$14401 ( \14449 , \14448 );
buf \U$14402 ( \14450 , \14449 );
and \U$14403 ( \14451 , \14393 , \14450 );
not \U$14404 ( \14452 , \14393 );
buf \U$14405 ( \14453 , \14446 );
and \U$14406 ( \14454 , \14452 , \14453 );
nor \U$14407 ( \14455 , \14451 , \14454 );
buf \U$14408 ( \14456 , \14455 );
buf \U$14409 ( \14457 , \14456 );
xor \U$14410 ( \14458 , \13213 , \13282 );
xor \U$14411 ( \14459 , \14458 , \13363 );
buf \U$14412 ( \14460 , \14459 );
buf \U$14413 ( \14461 , \14460 );
xor \U$14414 ( \14462 , \14457 , \14461 );
xor \U$14415 ( \14463 , RIc0db098_125, RIc0d7948_7);
buf \U$14416 ( \14464 , \14463 );
not \U$14417 ( \14465 , \14464 );
buf \U$14418 ( \14466 , \13460 );
not \U$14419 ( \14467 , \14466 );
buf \U$14420 ( \14468 , \14467 );
buf \U$14421 ( \14469 , \14468 );
not \U$14422 ( \14470 , \14469 );
buf \U$14423 ( \14471 , \14470 );
buf \U$14424 ( \14472 , \14471 );
not \U$14425 ( \14473 , \14472 );
or \U$14426 ( \14474 , \14465 , \14473 );
buf \U$14427 ( \14475 , \13465 );
buf \U$14428 ( \14476 , RIc0db098_125);
buf \U$14429 ( \14477 , RIc0d78d0_6);
xor \U$14430 ( \14478 , \14476 , \14477 );
buf \U$14431 ( \14479 , \14478 );
buf \U$14432 ( \14480 , \14479 );
nand \U$14433 ( \14481 , \14475 , \14480 );
buf \U$14434 ( \14482 , \14481 );
buf \U$14435 ( \14483 , \14482 );
nand \U$14436 ( \14484 , \14474 , \14483 );
buf \U$14437 ( \14485 , \14484 );
buf \U$14438 ( \14486 , \14485 );
buf \U$14439 ( \14487 , RIc0d9400_64);
buf \U$14440 ( \14488 , RIc0d96d0_70);
or \U$14441 ( \14489 , \14487 , \14488 );
buf \U$14442 ( \14490 , RIc0d9748_71);
nand \U$14443 ( \14491 , \14489 , \14490 );
buf \U$14444 ( \14492 , \14491 );
buf \U$14445 ( \14493 , \14492 );
buf \U$14446 ( \14494 , RIc0d9400_64);
buf \U$14447 ( \14495 , RIc0d96d0_70);
nand \U$14448 ( \14496 , \14494 , \14495 );
buf \U$14449 ( \14497 , \14496 );
buf \U$14450 ( \14498 , \14497 );
buf \U$14451 ( \14499 , RIc0d9658_69);
and \U$14452 ( \14500 , \14493 , \14498 , \14499 );
buf \U$14453 ( \14501 , \14500 );
buf \U$14454 ( \14502 , \14501 );
buf \U$14455 ( \14503 , RIc0d9310_62);
buf \U$14456 ( \14504 , RIc0d9748_71);
xor \U$14457 ( \14505 , \14503 , \14504 );
buf \U$14458 ( \14506 , \14505 );
buf \U$14459 ( \14507 , \14506 );
not \U$14460 ( \14508 , \14507 );
buf \U$14461 ( \14509 , \2923 );
not \U$14462 ( \14510 , \14509 );
or \U$14463 ( \14511 , \14508 , \14510 );
buf \U$14464 ( \14512 , \2927 );
buf \U$14465 ( \14513 , \13827 );
nand \U$14466 ( \14514 , \14512 , \14513 );
buf \U$14467 ( \14515 , \14514 );
buf \U$14468 ( \14516 , \14515 );
nand \U$14469 ( \14517 , \14511 , \14516 );
buf \U$14470 ( \14518 , \14517 );
buf \U$14471 ( \14519 , \14518 );
and \U$14472 ( \14520 , \14502 , \14519 );
buf \U$14473 ( \14521 , \14520 );
buf \U$14474 ( \14522 , \14521 );
xor \U$14475 ( \14523 , \14486 , \14522 );
buf \U$14476 ( \14524 , RIc0d8e60_52);
buf \U$14477 ( \14525 , RIc0d9bf8_81);
xor \U$14478 ( \14526 , \14524 , \14525 );
buf \U$14479 ( \14527 , \14526 );
buf \U$14480 ( \14528 , \14527 );
not \U$14481 ( \14529 , \14528 );
buf \U$14482 ( \14530 , \1060 );
not \U$14483 ( \14531 , \14530 );
buf \U$14484 ( \14532 , \14531 );
buf \U$14485 ( \14533 , \14532 );
not \U$14486 ( \14534 , \14533 );
or \U$14487 ( \14535 , \14529 , \14534 );
buf \U$14488 ( \14536 , \1078 );
buf \U$14489 ( \14537 , \13753 );
nand \U$14490 ( \14538 , \14536 , \14537 );
buf \U$14491 ( \14539 , \14538 );
buf \U$14492 ( \14540 , \14539 );
nand \U$14493 ( \14541 , \14535 , \14540 );
buf \U$14494 ( \14542 , \14541 );
buf \U$14495 ( \14543 , \14542 );
xor \U$14496 ( \14544 , RIc0d9dd8_85, RIc0d8c80_48);
buf \U$14497 ( \14545 , \14544 );
not \U$14498 ( \14546 , \14545 );
buf \U$14499 ( \14547 , \5304 );
not \U$14500 ( \14548 , \14547 );
or \U$14501 ( \14549 , \14546 , \14548 );
buf \U$14502 ( \14550 , \1401 );
buf \U$14503 ( \14551 , \13734 );
nand \U$14504 ( \14552 , \14550 , \14551 );
buf \U$14505 ( \14553 , \14552 );
buf \U$14506 ( \14554 , \14553 );
nand \U$14507 ( \14555 , \14549 , \14554 );
buf \U$14508 ( \14556 , \14555 );
buf \U$14509 ( \14557 , \14556 );
nor \U$14510 ( \14558 , \14543 , \14557 );
buf \U$14511 ( \14559 , \14558 );
buf \U$14512 ( \14560 , \14559 );
buf \U$14513 ( \14561 , RIc0d7c90_14);
buf \U$14514 ( \14562 , RIc0dadc8_119);
xor \U$14515 ( \14563 , \14561 , \14562 );
buf \U$14516 ( \14564 , \14563 );
buf \U$14517 ( \14565 , \14564 );
not \U$14518 ( \14566 , \14565 );
buf \U$14519 ( \14567 , \13178 );
not \U$14520 ( \14568 , \14567 );
buf \U$14521 ( \14569 , \14568 );
buf \U$14522 ( \14570 , \14569 );
not \U$14523 ( \14571 , \14570 );
or \U$14524 ( \14572 , \14566 , \14571 );
buf \U$14525 ( \14573 , \13953 );
buf \U$14526 ( \14574 , \13944 );
nand \U$14527 ( \14575 , \14573 , \14574 );
buf \U$14528 ( \14576 , \14575 );
buf \U$14529 ( \14577 , \14576 );
nand \U$14530 ( \14578 , \14572 , \14577 );
buf \U$14531 ( \14579 , \14578 );
buf \U$14532 ( \14580 , \14579 );
not \U$14533 ( \14581 , \14580 );
buf \U$14534 ( \14582 , \14581 );
buf \U$14535 ( \14583 , \14582 );
or \U$14536 ( \14584 , \14560 , \14583 );
buf \U$14537 ( \14585 , \14542 );
buf \U$14538 ( \14586 , \14556 );
nand \U$14539 ( \14587 , \14585 , \14586 );
buf \U$14540 ( \14588 , \14587 );
buf \U$14541 ( \14589 , \14588 );
nand \U$14542 ( \14590 , \14584 , \14589 );
buf \U$14543 ( \14591 , \14590 );
buf \U$14544 ( \14592 , \14591 );
and \U$14545 ( \14593 , \14523 , \14592 );
and \U$14546 ( \14594 , \14486 , \14522 );
or \U$14547 ( \14595 , \14593 , \14594 );
buf \U$14548 ( \14596 , \14595 );
buf \U$14549 ( \14597 , \14596 );
buf \U$14550 ( \14598 , RIc0d9220_60);
buf \U$14551 ( \14599 , RIc0d9838_73);
xor \U$14552 ( \14600 , \14598 , \14599 );
buf \U$14553 ( \14601 , \14600 );
buf \U$14554 ( \14602 , \14601 );
not \U$14555 ( \14603 , \14602 );
buf \U$14556 ( \14604 , \769 );
not \U$14557 ( \14605 , \14604 );
buf \U$14558 ( \14606 , \790 );
nor \U$14559 ( \14607 , \14605 , \14606 );
buf \U$14560 ( \14608 , \14607 );
buf \U$14561 ( \14609 , \14608 );
not \U$14562 ( \14610 , \14609 );
or \U$14563 ( \14611 , \14603 , \14610 );
buf \U$14564 ( \14612 , \791 );
buf \U$14565 ( \14613 , \14070 );
nand \U$14566 ( \14614 , \14612 , \14613 );
buf \U$14567 ( \14615 , \14614 );
buf \U$14568 ( \14616 , \14615 );
nand \U$14569 ( \14617 , \14611 , \14616 );
buf \U$14570 ( \14618 , \14617 );
buf \U$14571 ( \14619 , \14618 );
not \U$14572 ( \14620 , \14619 );
xor \U$14573 ( \14621 , RIc0d9ec8_87, RIc0d8b90_46);
buf \U$14574 ( \14622 , \14621 );
not \U$14575 ( \14623 , \14622 );
buf \U$14576 ( \14624 , \14325 );
not \U$14577 ( \14625 , \14624 );
or \U$14578 ( \14626 , \14623 , \14625 );
buf \U$14579 ( \14627 , \816 );
buf \U$14580 ( \14628 , \14015 );
nand \U$14581 ( \14629 , \14627 , \14628 );
buf \U$14582 ( \14630 , \14629 );
buf \U$14583 ( \14631 , \14630 );
nand \U$14584 ( \14632 , \14626 , \14631 );
buf \U$14585 ( \14633 , \14632 );
buf \U$14586 ( \14634 , \14633 );
not \U$14587 ( \14635 , \14634 );
or \U$14588 ( \14636 , \14620 , \14635 );
buf \U$14589 ( \14637 , \14633 );
buf \U$14590 ( \14638 , \14618 );
or \U$14591 ( \14639 , \14637 , \14638 );
xor \U$14592 ( \14640 , RIc0da468_99, RIc0d85f0_34);
buf \U$14593 ( \14641 , \14640 );
not \U$14594 ( \14642 , \14641 );
buf \U$14595 ( \14643 , \12578 );
not \U$14596 ( \14644 , \14643 );
or \U$14597 ( \14645 , \14642 , \14644 );
buf \U$14598 ( \14646 , \2199 );
not \U$14599 ( \14647 , \14646 );
buf \U$14600 ( \14648 , \14647 );
buf \U$14601 ( \14649 , \14648 );
buf \U$14602 ( \14650 , \14132 );
nand \U$14603 ( \14651 , \14649 , \14650 );
buf \U$14604 ( \14652 , \14651 );
buf \U$14605 ( \14653 , \14652 );
nand \U$14606 ( \14654 , \14645 , \14653 );
buf \U$14607 ( \14655 , \14654 );
buf \U$14608 ( \14656 , \14655 );
nand \U$14609 ( \14657 , \14639 , \14656 );
buf \U$14610 ( \14658 , \14657 );
buf \U$14611 ( \14659 , \14658 );
nand \U$14612 ( \14660 , \14636 , \14659 );
buf \U$14613 ( \14661 , \14660 );
buf \U$14614 ( \14662 , \14661 );
not \U$14615 ( \14663 , \14662 );
xor \U$14616 ( \14664 , RIc0da918_109, RIc0d8140_24);
buf \U$14617 ( \14665 , \14664 );
not \U$14618 ( \14666 , \14665 );
buf \U$14619 ( \14667 , \13419 );
not \U$14620 ( \14668 , \14667 );
or \U$14621 ( \14669 , \14666 , \14668 );
buf \U$14622 ( \14670 , \14216 );
buf \U$14623 ( \14671 , \14200 );
nand \U$14624 ( \14672 , \14670 , \14671 );
buf \U$14625 ( \14673 , \14672 );
buf \U$14626 ( \14674 , \14673 );
nand \U$14627 ( \14675 , \14669 , \14674 );
buf \U$14628 ( \14676 , \14675 );
buf \U$14629 ( \14677 , \14676 );
xor \U$14630 ( \14678 , RIc0dabe8_115, RIc0d7e70_18);
buf \U$14631 ( \14679 , \14678 );
not \U$14632 ( \14680 , \14679 );
buf \U$14635 ( \14681 , \14183 );
buf \U$14636 ( \14682 , \14681 );
not \U$14637 ( \14683 , \14682 );
buf \U$14638 ( \14684 , \14683 );
buf \U$14639 ( \14685 , \14684 );
not \U$14640 ( \14686 , \14685 );
or \U$14641 ( \14687 , \14680 , \14686 );
buf \U$14642 ( \14688 , \12278 );
not \U$14643 ( \14689 , \14688 );
buf \U$14644 ( \14690 , \14689 );
buf \U$14645 ( \14691 , \14690 );
buf \U$14646 ( \14692 , \14173 );
nand \U$14647 ( \14693 , \14691 , \14692 );
buf \U$14648 ( \14694 , \14693 );
buf \U$14649 ( \14695 , \14694 );
nand \U$14650 ( \14696 , \14687 , \14695 );
buf \U$14651 ( \14697 , \14696 );
buf \U$14652 ( \14698 , \14697 );
xor \U$14653 ( \14699 , \14677 , \14698 );
buf \U$14654 ( \14700 , \13853 );
not \U$14655 ( \14701 , \14700 );
buf \U$14656 ( \14702 , \343 );
not \U$14657 ( \14703 , \14702 );
buf \U$14658 ( \14704 , \14703 );
buf \U$14659 ( \14705 , \14704 );
not \U$14660 ( \14706 , \14705 );
buf \U$14661 ( \14707 , \14706 );
buf \U$14662 ( \14708 , \14707 );
not \U$14663 ( \14709 , \14708 );
or \U$14664 ( \14710 , \14701 , \14709 );
buf \U$14665 ( \14711 , \3714 );
not \U$14666 ( \14712 , \14711 );
buf \U$14667 ( \14713 , \14712 );
buf \U$14668 ( \14714 , \14713 );
xnor \U$14669 ( \14715 , RIc0da288_95, RIc0d87d0_38);
buf \U$14670 ( \14716 , \14715 );
or \U$14671 ( \14717 , \14714 , \14716 );
nand \U$14672 ( \14718 , \14710 , \14717 );
buf \U$14673 ( \14719 , \14718 );
buf \U$14674 ( \14720 , \14719 );
and \U$14675 ( \14721 , \14699 , \14720 );
and \U$14676 ( \14722 , \14677 , \14698 );
or \U$14677 ( \14723 , \14721 , \14722 );
buf \U$14678 ( \14724 , \14723 );
buf \U$14679 ( \14725 , \14724 );
not \U$14680 ( \14726 , \14725 );
or \U$14681 ( \14727 , \14663 , \14726 );
buf \U$14682 ( \14728 , \14724 );
buf \U$14683 ( \14729 , \14661 );
or \U$14684 ( \14730 , \14728 , \14729 );
buf \U$14685 ( \14731 , RIc0d9130_58);
buf \U$14686 ( \14732 , RIc0d9928_75);
xor \U$14687 ( \14733 , \14731 , \14732 );
buf \U$14688 ( \14734 , \14733 );
buf \U$14689 ( \14735 , \14734 );
not \U$14690 ( \14736 , \14735 );
buf \U$14691 ( \14737 , \13991 );
not \U$14692 ( \14738 , \14737 );
or \U$14693 ( \14739 , \14736 , \14738 );
buf \U$14694 ( \14740 , \13998 );
buf \U$14695 ( \14741 , \13985 );
nand \U$14696 ( \14742 , \14740 , \14741 );
buf \U$14697 ( \14743 , \14742 );
buf \U$14698 ( \14744 , \14743 );
nand \U$14699 ( \14745 , \14739 , \14744 );
buf \U$14700 ( \14746 , \14745 );
buf \U$14701 ( \14747 , \14746 );
not \U$14702 ( \14748 , \14747 );
buf \U$14703 ( \14749 , RIc0d9400_64);
buf \U$14704 ( \14750 , RIc0d9658_69);
xor \U$14705 ( \14751 , \14749 , \14750 );
buf \U$14706 ( \14752 , \14751 );
buf \U$14707 ( \14753 , \14752 );
not \U$14708 ( \14754 , \14753 );
buf \U$14709 ( \14755 , \278 );
not \U$14710 ( \14756 , \14755 );
or \U$14711 ( \14757 , \14754 , \14756 );
buf \U$14712 ( \14758 , \283 );
buf \U$14713 ( \14759 , \14159 );
nand \U$14714 ( \14760 , \14758 , \14759 );
buf \U$14715 ( \14761 , \14760 );
buf \U$14716 ( \14762 , \14761 );
nand \U$14717 ( \14763 , \14757 , \14762 );
buf \U$14718 ( \14764 , \14763 );
buf \U$14719 ( \14765 , \14764 );
not \U$14720 ( \14766 , \14765 );
or \U$14721 ( \14767 , \14748 , \14766 );
or \U$14722 ( \14768 , \14764 , \14746 );
buf \U$14723 ( \14769 , RIc0d8500_32);
buf \U$14724 ( \14770 , RIc0da558_101);
xor \U$14725 ( \14771 , \14769 , \14770 );
buf \U$14726 ( \14772 , \14771 );
buf \U$14727 ( \14773 , \14772 );
not \U$14728 ( \14774 , \14773 );
buf \U$14729 ( \14775 , \4042 );
not \U$14730 ( \14776 , \14775 );
or \U$14731 ( \14777 , \14774 , \14776 );
buf \U$14732 ( \14778 , \4049 );
buf \U$14733 ( \14779 , \14038 );
nand \U$14734 ( \14780 , \14778 , \14779 );
buf \U$14735 ( \14781 , \14780 );
buf \U$14736 ( \14782 , \14781 );
nand \U$14737 ( \14783 , \14777 , \14782 );
buf \U$14738 ( \14784 , \14783 );
nand \U$14739 ( \14785 , \14768 , \14784 );
buf \U$14740 ( \14786 , \14785 );
nand \U$14741 ( \14787 , \14767 , \14786 );
buf \U$14742 ( \14788 , \14787 );
buf \U$14743 ( \14789 , \14788 );
nand \U$14744 ( \14790 , \14730 , \14789 );
buf \U$14745 ( \14791 , \14790 );
buf \U$14746 ( \14792 , \14791 );
nand \U$14747 ( \14793 , \14727 , \14792 );
buf \U$14748 ( \14794 , \14793 );
buf \U$14749 ( \14795 , \14794 );
xor \U$14750 ( \14796 , \14597 , \14795 );
xor \U$14751 ( \14797 , RIc0da738_105, RIc0d8320_28);
buf \U$14752 ( \14798 , \14797 );
not \U$14753 ( \14799 , \14798 );
buf \U$14754 ( \14800 , \12731 );
not \U$14755 ( \14801 , \14800 );
buf \U$14756 ( \14802 , \12743 );
nor \U$14757 ( \14803 , \14801 , \14802 );
buf \U$14758 ( \14804 , \14803 );
buf \U$14759 ( \14805 , \14804 );
not \U$14760 ( \14806 , \14805 );
or \U$14761 ( \14807 , \14799 , \14806 );
buf \U$14762 ( \14808 , \12744 );
buf \U$14763 ( \14809 , \13918 );
nand \U$14764 ( \14810 , \14808 , \14809 );
buf \U$14765 ( \14811 , \14810 );
buf \U$14766 ( \14812 , \14811 );
nand \U$14767 ( \14813 , \14807 , \14812 );
buf \U$14768 ( \14814 , \14813 );
not \U$14769 ( \14815 , \14814 );
buf \U$14770 ( \14816 , RIc0d9040_56);
buf \U$14771 ( \14817 , RIc0d9a18_77);
xor \U$14772 ( \14818 , \14816 , \14817 );
buf \U$14773 ( \14819 , \14818 );
buf \U$14774 ( \14820 , \14819 );
not \U$14775 ( \14821 , \14820 );
buf \U$14776 ( \14822 , \1174 );
buf \U$14777 ( \14823 , \1176 );
and \U$14778 ( \14824 , \14822 , \14823 );
buf \U$14779 ( \14825 , \14824 );
buf \U$14780 ( \14826 , \14825 );
not \U$14781 ( \14827 , \14826 );
or \U$14782 ( \14828 , \14821 , \14827 );
buf \U$14783 ( \14829 , \3742 );
buf \U$14784 ( \14830 , \13661 );
nand \U$14785 ( \14831 , \14829 , \14830 );
buf \U$14786 ( \14832 , \14831 );
buf \U$14787 ( \14833 , \14832 );
nand \U$14788 ( \14834 , \14828 , \14833 );
buf \U$14789 ( \14835 , \14834 );
not \U$14790 ( \14836 , \14835 );
or \U$14791 ( \14837 , \14815 , \14836 );
buf \U$14792 ( \14838 , \14835 );
not \U$14793 ( \14839 , \14838 );
buf \U$14794 ( \14840 , \14839 );
not \U$14795 ( \14841 , \14840 );
buf \U$14796 ( \14842 , \14814 );
not \U$14797 ( \14843 , \14842 );
buf \U$14798 ( \14844 , \14843 );
not \U$14799 ( \14845 , \14844 );
or \U$14800 ( \14846 , \14841 , \14845 );
xor \U$14801 ( \14847 , RIc0da0a8_91, RIc0d89b0_42);
buf \U$14802 ( \14848 , \14847 );
not \U$14803 ( \14849 , \14848 );
buf \U$14804 ( \14850 , \1927 );
not \U$14805 ( \14851 , \14850 );
or \U$14806 ( \14852 , \14849 , \14851 );
buf \U$14807 ( \14853 , \533 );
buf \U$14808 ( \14854 , \13905 );
nand \U$14809 ( \14855 , \14853 , \14854 );
buf \U$14810 ( \14856 , \14855 );
buf \U$14811 ( \14857 , \14856 );
nand \U$14812 ( \14858 , \14852 , \14857 );
buf \U$14813 ( \14859 , \14858 );
nand \U$14814 ( \14860 , \14846 , \14859 );
nand \U$14815 ( \14861 , \14837 , \14860 );
buf \U$14816 ( \14862 , \14861 );
buf \U$14817 ( \14863 , RIc0d8050_22);
buf \U$14818 ( \14864 , RIc0daa08_111);
xor \U$14819 ( \14865 , \14863 , \14864 );
buf \U$14820 ( \14866 , \14865 );
buf \U$14821 ( \14867 , \14866 );
not \U$14822 ( \14868 , \14867 );
buf \U$14823 ( \14869 , \14100 );
not \U$14824 ( \14870 , \14869 );
or \U$14825 ( \14871 , \14868 , \14870 );
buf \U$14826 ( \14872 , \14353 );
buf \U$14827 ( \14873 , \14094 );
nand \U$14828 ( \14874 , \14872 , \14873 );
buf \U$14829 ( \14875 , \14874 );
buf \U$14830 ( \14876 , \14875 );
nand \U$14831 ( \14877 , \14871 , \14876 );
buf \U$14832 ( \14878 , \14877 );
buf \U$14833 ( \14879 , \14878 );
not \U$14834 ( \14880 , \14879 );
xor \U$14835 ( \14881 , RIc0daaf8_113, RIc0d7f60_20);
buf \U$14836 ( \14882 , \14881 );
not \U$14837 ( \14883 , \14882 );
buf \U$14838 ( \14884 , \12394 );
buf \U$14839 ( \14885 , \12396 );
nand \U$14840 ( \14886 , \14884 , \14885 );
buf \U$14841 ( \14887 , \14886 );
buf \U$14844 ( \14888 , \14887 );
buf \U$14845 ( \14889 , \14888 );
not \U$14846 ( \14890 , \14889 );
buf \U$14847 ( \14891 , \14890 );
buf \U$14848 ( \14892 , \14891 );
not \U$14849 ( \14893 , \14892 );
or \U$14850 ( \14894 , \14883 , \14893 );
buf \U$14851 ( \14895 , \12410 );
buf \U$14852 ( \14896 , \13597 );
nand \U$14853 ( \14897 , \14895 , \14896 );
buf \U$14854 ( \14898 , \14897 );
buf \U$14855 ( \14899 , \14898 );
nand \U$14856 ( \14900 , \14894 , \14899 );
buf \U$14857 ( \14901 , \14900 );
buf \U$14858 ( \14902 , \14901 );
not \U$14859 ( \14903 , \14902 );
or \U$14860 ( \14904 , \14880 , \14903 );
buf \U$14861 ( \14905 , \14901 );
buf \U$14862 ( \14906 , \14878 );
or \U$14863 ( \14907 , \14905 , \14906 );
buf \U$14864 ( \14908 , RIc0d8d70_50);
buf \U$14865 ( \14909 , RIc0d9ce8_83);
xor \U$14866 ( \14910 , \14908 , \14909 );
buf \U$14867 ( \14911 , \14910 );
buf \U$14868 ( \14912 , \14911 );
not \U$14869 ( \14913 , \14912 );
buf \U$14870 ( \14914 , \12254 );
not \U$14871 ( \14915 , \14914 );
or \U$14872 ( \14916 , \14913 , \14915 );
buf \U$14873 ( \14917 , \584 );
buf \U$14874 ( \14918 , \13637 );
nand \U$14875 ( \14919 , \14917 , \14918 );
buf \U$14876 ( \14920 , \14919 );
buf \U$14877 ( \14921 , \14920 );
nand \U$14878 ( \14922 , \14916 , \14921 );
buf \U$14879 ( \14923 , \14922 );
buf \U$14880 ( \14924 , \14923 );
nand \U$14881 ( \14925 , \14907 , \14924 );
buf \U$14882 ( \14926 , \14925 );
buf \U$14883 ( \14927 , \14926 );
nand \U$14884 ( \14928 , \14904 , \14927 );
buf \U$14885 ( \14929 , \14928 );
buf \U$14886 ( \14930 , \14929 );
xor \U$14887 ( \14931 , \14862 , \14930 );
buf \U$14888 ( \14932 , RIc0d9b08_79);
buf \U$14889 ( \14933 , RIc0d8f50_54);
xor \U$14890 ( \14934 , \14932 , \14933 );
buf \U$14891 ( \14935 , \14934 );
buf \U$14892 ( \14936 , \14935 );
not \U$14893 ( \14937 , \14936 );
buf \U$14894 ( \14938 , \393 );
not \U$14895 ( \14939 , \14938 );
buf \U$14896 ( \14940 , \14939 );
buf \U$14897 ( \14941 , \14940 );
not \U$14898 ( \14942 , \14941 );
or \U$14899 ( \14943 , \14937 , \14942 );
buf \U$14900 ( \14944 , \402 );
buf \U$14901 ( \14945 , RIc0d8ed8_53);
buf \U$14902 ( \14946 , RIc0d9b08_79);
xor \U$14903 ( \14947 , \14945 , \14946 );
buf \U$14904 ( \14948 , \14947 );
buf \U$14905 ( \14949 , \14948 );
nand \U$14906 ( \14950 , \14944 , \14949 );
buf \U$14907 ( \14951 , \14950 );
buf \U$14908 ( \14952 , \14951 );
nand \U$14909 ( \14953 , \14943 , \14952 );
buf \U$14910 ( \14954 , \14953 );
buf \U$14911 ( \14955 , \14954 );
buf \U$14912 ( \14956 , RIc0d8aa0_44);
buf \U$14913 ( \14957 , RIc0d9fb8_89);
xor \U$14914 ( \14958 , \14956 , \14957 );
buf \U$14915 ( \14959 , \14958 );
buf \U$14916 ( \14960 , \14959 );
not \U$14917 ( \14961 , \14960 );
buf \U$14918 ( \14962 , \842 );
not \U$14919 ( \14963 , \14962 );
or \U$14920 ( \14964 , \14961 , \14963 );
buf \U$14921 ( \14965 , \846 );
buf \U$14922 ( \14966 , \13626 );
nand \U$14923 ( \14967 , \14965 , \14966 );
buf \U$14924 ( \14968 , \14967 );
buf \U$14925 ( \14969 , \14968 );
nand \U$14926 ( \14970 , \14964 , \14969 );
buf \U$14927 ( \14971 , \14970 );
buf \U$14928 ( \14972 , \14971 );
or \U$14929 ( \14973 , \14955 , \14972 );
xor \U$14930 ( \14974 , RIc0dafa8_123, RIc0d7ab0_10);
buf \U$14931 ( \14975 , \14974 );
not \U$14932 ( \14976 , \14975 );
buf \U$14933 ( \14977 , \12861 );
not \U$14934 ( \14978 , \14977 );
buf \U$14935 ( \14979 , \12867 );
nor \U$14936 ( \14980 , \14978 , \14979 );
buf \U$14937 ( \14981 , \14980 );
buf \U$14940 ( \14982 , \14981 );
buf \U$14941 ( \14983 , \14982 );
not \U$14942 ( \14984 , \14983 );
or \U$14943 ( \14985 , \14976 , \14984 );
buf \U$14944 ( \14986 , \14278 );
buf \U$14945 ( \14987 , RIc0d7a38_9);
buf \U$14946 ( \14988 , RIc0dafa8_123);
xor \U$14947 ( \14989 , \14987 , \14988 );
buf \U$14948 ( \14990 , \14989 );
buf \U$14949 ( \14991 , \14990 );
nand \U$14950 ( \14992 , \14986 , \14991 );
buf \U$14951 ( \14993 , \14992 );
buf \U$14952 ( \14994 , \14993 );
nand \U$14953 ( \14995 , \14985 , \14994 );
buf \U$14954 ( \14996 , \14995 );
buf \U$14955 ( \14997 , \14996 );
nand \U$14956 ( \14998 , \14973 , \14997 );
buf \U$14957 ( \14999 , \14998 );
buf \U$14958 ( \15000 , \14999 );
buf \U$14959 ( \15001 , \14971 );
buf \U$14960 ( \15002 , \14954 );
nand \U$14961 ( \15003 , \15001 , \15002 );
buf \U$14962 ( \15004 , \15003 );
buf \U$14963 ( \15005 , \15004 );
nand \U$14964 ( \15006 , \15000 , \15005 );
buf \U$14965 ( \15007 , \15006 );
buf \U$14966 ( \15008 , \15007 );
and \U$14967 ( \15009 , \14931 , \15008 );
and \U$14968 ( \15010 , \14862 , \14930 );
or \U$14969 ( \15011 , \15009 , \15010 );
buf \U$14970 ( \15012 , \15011 );
buf \U$14971 ( \15013 , \15012 );
and \U$14972 ( \15014 , \14796 , \15013 );
and \U$14973 ( \15015 , \14597 , \14795 );
or \U$14974 ( \15016 , \15014 , \15015 );
buf \U$14975 ( \15017 , \15016 );
buf \U$14976 ( \15018 , \15017 );
and \U$14977 ( \15019 , \14462 , \15018 );
and \U$14978 ( \15020 , \14457 , \14461 );
or \U$14979 ( \15021 , \15019 , \15020 );
buf \U$14980 ( \15022 , \15021 );
buf \U$14981 ( \15023 , \15022 );
and \U$14982 ( \15024 , \14247 , \15023 );
and \U$14983 ( \15025 , \13137 , \14246 );
or \U$14984 ( \15026 , \15024 , \15025 );
buf \U$14985 ( \15027 , \15026 );
buf \U$14986 ( \15028 , \15027 );
not \U$14987 ( \15029 , \15028 );
buf \U$14988 ( \15030 , \15029 );
buf \U$14989 ( \15031 , \15030 );
not \U$14990 ( \15032 , \12850 );
not \U$14991 ( \15033 , \12888 );
or \U$14992 ( \15034 , \15032 , \15033 );
not \U$14993 ( \15035 , \12891 );
not \U$14994 ( \15036 , \12896 );
or \U$14995 ( \15037 , \15035 , \15036 );
nand \U$14996 ( \15038 , \15037 , \12948 );
nand \U$14997 ( \15039 , \15034 , \15038 );
buf \U$14998 ( \15040 , \15039 );
not \U$14999 ( \15041 , \12499 );
not \U$15000 ( \15042 , \12477 );
or \U$15001 ( \15043 , \15041 , \15042 );
not \U$15002 ( \15044 , \12509 );
not \U$15003 ( \15045 , \12502 );
or \U$15004 ( \15046 , \15044 , \15045 );
nand \U$15005 ( \15047 , \15046 , \12553 );
nand \U$15006 ( \15048 , \15043 , \15047 );
buf \U$15007 ( \15049 , \15048 );
xor \U$15008 ( \15050 , \15040 , \15049 );
xor \U$15009 ( \15051 , \12596 , \12617 );
and \U$15010 ( \15052 , \15051 , \12636 );
and \U$15011 ( \15053 , \12596 , \12617 );
or \U$15012 ( \15054 , \15052 , \15053 );
buf \U$15013 ( \15055 , \15054 );
buf \U$15014 ( \15056 , \15055 );
xor \U$15015 ( \15057 , \15050 , \15056 );
buf \U$15016 ( \15058 , \15057 );
buf \U$15017 ( \15059 , \12428 );
not \U$15018 ( \15060 , \15059 );
buf \U$15019 ( \15061 , \12422 );
not \U$15020 ( \15062 , \15061 );
or \U$15021 ( \15063 , \15060 , \15062 );
buf \U$15022 ( \15064 , \12453 );
nand \U$15023 ( \15065 , \15063 , \15064 );
buf \U$15024 ( \15066 , \15065 );
buf \U$15025 ( \15067 , \15066 );
buf \U$15026 ( \15068 , \12428 );
not \U$15027 ( \15069 , \15068 );
buf \U$15028 ( \15070 , \12421 );
nand \U$15029 ( \15071 , \15069 , \15070 );
buf \U$15030 ( \15072 , \15071 );
buf \U$15031 ( \15073 , \15072 );
nand \U$15032 ( \15074 , \15067 , \15073 );
buf \U$15033 ( \15075 , \15074 );
buf \U$15034 ( \15076 , \15075 );
not \U$15035 ( \15077 , \15076 );
buf \U$15036 ( \15078 , \15077 );
buf \U$15037 ( \15079 , \12716 );
not \U$15038 ( \15080 , \15079 );
buf \U$15039 ( \15081 , \12694 );
buf \U$15040 ( \15082 , \12668 );
or \U$15041 ( \15083 , \15081 , \15082 );
buf \U$15042 ( \15084 , \15083 );
buf \U$15043 ( \15085 , \15084 );
not \U$15044 ( \15086 , \15085 );
or \U$15045 ( \15087 , \15080 , \15086 );
buf \U$15046 ( \15088 , \12694 );
buf \U$15047 ( \15089 , \12668 );
nand \U$15048 ( \15090 , \15088 , \15089 );
buf \U$15049 ( \15091 , \15090 );
buf \U$15050 ( \15092 , \15091 );
nand \U$15051 ( \15093 , \15087 , \15092 );
buf \U$15052 ( \15094 , \15093 );
xor \U$15053 ( \15095 , \15078 , \15094 );
and \U$15054 ( \15096 , \12787 , \12788 );
buf \U$15055 ( \15097 , \15096 );
buf \U$15056 ( \15098 , \15097 );
buf \U$15057 ( \15099 , \13124 );
not \U$15058 ( \15100 , \15099 );
buf \U$15059 ( \15101 , \524 );
not \U$15060 ( \15102 , \15101 );
or \U$15061 ( \15103 , \15100 , \15102 );
buf \U$15062 ( \15104 , \714 );
xor \U$15063 ( \15105 , RIc0da0a8_91, RIc0d86e0_36);
buf \U$15064 ( \15106 , \15105 );
nand \U$15065 ( \15107 , \15104 , \15106 );
buf \U$15066 ( \15108 , \15107 );
buf \U$15067 ( \15109 , \15108 );
nand \U$15068 ( \15110 , \15103 , \15109 );
buf \U$15069 ( \15111 , \15110 );
buf \U$15070 ( \15112 , \15111 );
xor \U$15071 ( \15113 , \15098 , \15112 );
buf \U$15072 ( \15114 , \13533 );
not \U$15073 ( \15115 , \15114 );
buf \U$15074 ( \15116 , \2900 );
not \U$15075 ( \15117 , \15116 );
or \U$15076 ( \15118 , \15115 , \15117 );
buf \U$15077 ( \15119 , \686 );
buf \U$15078 ( \15120 , RIc0d9220_60);
buf \U$15079 ( \15121 , RIc0d9568_67);
xor \U$15080 ( \15122 , \15120 , \15121 );
buf \U$15081 ( \15123 , \15122 );
buf \U$15082 ( \15124 , \15123 );
nand \U$15083 ( \15125 , \15119 , \15124 );
buf \U$15084 ( \15126 , \15125 );
buf \U$15085 ( \15127 , \15126 );
nand \U$15086 ( \15128 , \15118 , \15127 );
buf \U$15087 ( \15129 , \15128 );
buf \U$15088 ( \15130 , \15129 );
xor \U$15089 ( \15131 , \15113 , \15130 );
buf \U$15090 ( \15132 , \15131 );
xor \U$15091 ( \15133 , \15095 , \15132 );
and \U$15092 ( \15134 , \15058 , \15133 );
not \U$15093 ( \15135 , \15058 );
buf \U$15094 ( \15136 , \15133 );
not \U$15095 ( \15137 , \15136 );
buf \U$15096 ( \15138 , \15137 );
and \U$15097 ( \15139 , \15135 , \15138 );
or \U$15098 ( \15140 , \15134 , \15139 );
buf \U$15099 ( \15141 , \15140 );
xor \U$15100 ( \15142 , \12265 , \12314 );
and \U$15101 ( \15143 , \15142 , \12350 );
and \U$15102 ( \15144 , \12265 , \12314 );
or \U$15103 ( \15145 , \15143 , \15144 );
or \U$15104 ( \15146 , \13400 , \13437 );
nand \U$15105 ( \15147 , \15146 , \13476 );
buf \U$15106 ( \15148 , \15147 );
buf \U$15107 ( \15149 , \13437 );
buf \U$15108 ( \15150 , \13400 );
nand \U$15109 ( \15151 , \15149 , \15150 );
buf \U$15110 ( \15152 , \15151 );
buf \U$15111 ( \15153 , \15152 );
nand \U$15112 ( \15154 , \15148 , \15153 );
buf \U$15113 ( \15155 , \15154 );
xor \U$15114 ( \15156 , \15145 , \15155 );
buf \U$15115 ( \15157 , \15156 );
buf \U$15116 ( \15158 , \12777 );
not \U$15117 ( \15159 , \15158 );
buf \U$15118 ( \15160 , \12815 );
not \U$15119 ( \15161 , \15160 );
or \U$15120 ( \15162 , \15159 , \15161 );
buf \U$15121 ( \15163 , \12755 );
nand \U$15122 ( \15164 , \15162 , \15163 );
buf \U$15123 ( \15165 , \15164 );
buf \U$15124 ( \15166 , \15165 );
buf \U$15125 ( \15167 , \12774 );
buf \U$15126 ( \15168 , \12809 );
nand \U$15127 ( \15169 , \15167 , \15168 );
buf \U$15128 ( \15170 , \15169 );
buf \U$15129 ( \15171 , \15170 );
nand \U$15130 ( \15172 , \15166 , \15171 );
buf \U$15131 ( \15173 , \15172 );
buf \U$15134 ( \15174 , \15173 );
buf \U$15135 ( \15175 , \15174 );
not \U$15136 ( \15176 , \15175 );
buf \U$15137 ( \15177 , \15176 );
buf \U$15138 ( \15178 , \15177 );
and \U$15139 ( \15179 , \15157 , \15178 );
not \U$15140 ( \15180 , \15157 );
buf \U$15141 ( \15181 , \15174 );
and \U$15142 ( \15182 , \15180 , \15181 );
nor \U$15143 ( \15183 , \15179 , \15182 );
buf \U$15144 ( \15184 , \15183 );
buf \U$15145 ( \15185 , \15184 );
not \U$15146 ( \15186 , \15185 );
buf \U$15147 ( \15187 , \15186 );
buf \U$15148 ( \15188 , \15187 );
and \U$15149 ( \15189 , \15141 , \15188 );
not \U$15150 ( \15190 , \15141 );
buf \U$15151 ( \15191 , \15184 );
and \U$15152 ( \15192 , \15190 , \15191 );
nor \U$15153 ( \15193 , \15189 , \15192 );
buf \U$15154 ( \15194 , \15193 );
buf \U$15155 ( \15195 , \15194 );
buf \U$15156 ( \15196 , \13065 );
not \U$15157 ( \15197 , \15196 );
buf \U$15158 ( \15198 , \12949 );
not \U$15159 ( \15199 , \15198 );
buf \U$15160 ( \15200 , \15199 );
buf \U$15161 ( \15201 , \15200 );
not \U$15162 ( \15202 , \15201 );
or \U$15163 ( \15203 , \15197 , \15202 );
buf \U$15164 ( \15204 , \13062 );
not \U$15165 ( \15205 , \15204 );
buf \U$15166 ( \15206 , \12949 );
not \U$15167 ( \15207 , \15206 );
or \U$15168 ( \15208 , \15205 , \15207 );
buf \U$15169 ( \15209 , \13131 );
nand \U$15170 ( \15210 , \15208 , \15209 );
buf \U$15171 ( \15211 , \15210 );
buf \U$15172 ( \15212 , \15211 );
nand \U$15173 ( \15213 , \15203 , \15212 );
buf \U$15174 ( \15214 , \15213 );
buf \U$15175 ( \15215 , \15214 );
not \U$15176 ( \15216 , \15215 );
buf \U$15177 ( \15217 , \12638 );
not \U$15178 ( \15218 , \15217 );
buf \U$15179 ( \15219 , \12719 );
not \U$15180 ( \15220 , \15219 );
buf \U$15181 ( \15221 , \15220 );
buf \U$15182 ( \15222 , \15221 );
not \U$15183 ( \15223 , \15222 );
or \U$15184 ( \15224 , \15218 , \15223 );
buf \U$15185 ( \15225 , \12638 );
not \U$15186 ( \15226 , \15225 );
buf \U$15187 ( \15227 , \15226 );
buf \U$15188 ( \15228 , \15227 );
not \U$15189 ( \15229 , \15228 );
buf \U$15190 ( \15230 , \12719 );
not \U$15191 ( \15231 , \15230 );
or \U$15192 ( \15232 , \15229 , \15231 );
buf \U$15193 ( \15233 , \12819 );
nand \U$15194 ( \15234 , \15232 , \15233 );
buf \U$15195 ( \15235 , \15234 );
buf \U$15196 ( \15236 , \15235 );
nand \U$15197 ( \15237 , \15224 , \15236 );
buf \U$15198 ( \15238 , \15237 );
buf \U$15199 ( \15239 , \15238 );
not \U$15200 ( \15240 , \15239 );
buf \U$15201 ( \15241 , \15240 );
buf \U$15202 ( \15242 , \15241 );
not \U$15203 ( \15243 , \15242 );
or \U$15204 ( \15244 , \15216 , \15243 );
buf \U$15205 ( \15245 , \15214 );
buf \U$15206 ( \15246 , \15241 );
or \U$15207 ( \15247 , \15245 , \15246 );
nand \U$15208 ( \15248 , \15244 , \15247 );
buf \U$15209 ( \15249 , \15248 );
buf \U$15210 ( \15250 , \15249 );
buf \U$15211 ( \15251 , \12456 );
not \U$15212 ( \15252 , \15251 );
buf \U$15213 ( \15253 , \12563 );
not \U$15214 ( \15254 , \15253 );
or \U$15215 ( \15255 , \15252 , \15254 );
buf \U$15216 ( \15256 , \12351 );
nand \U$15217 ( \15257 , \15255 , \15256 );
buf \U$15218 ( \15258 , \15257 );
buf \U$15219 ( \15259 , \15258 );
buf \U$15220 ( \15260 , \12456 );
not \U$15221 ( \15261 , \15260 );
buf \U$15222 ( \15262 , \12566 );
nand \U$15223 ( \15263 , \15261 , \15262 );
buf \U$15224 ( \15264 , \15263 );
buf \U$15225 ( \15265 , \15264 );
nand \U$15226 ( \15266 , \15259 , \15265 );
buf \U$15227 ( \15267 , \15266 );
buf \U$15228 ( \15268 , \15267 );
and \U$15229 ( \15269 , \15250 , \15268 );
not \U$15230 ( \15270 , \15250 );
buf \U$15231 ( \15271 , \15267 );
not \U$15232 ( \15272 , \15271 );
buf \U$15233 ( \15273 , \15272 );
buf \U$15234 ( \15274 , \15273 );
and \U$15235 ( \15275 , \15270 , \15274 );
nor \U$15236 ( \15276 , \15269 , \15275 );
buf \U$15237 ( \15277 , \15276 );
buf \U$15238 ( \15278 , \15277 );
not \U$15239 ( \15279 , \15278 );
buf \U$15240 ( \15280 , \15279 );
buf \U$15241 ( \15281 , \15280 );
and \U$15242 ( \15282 , \15195 , \15281 );
not \U$15243 ( \15283 , \15195 );
buf \U$15244 ( \15284 , \15277 );
and \U$15245 ( \15285 , \15283 , \15284 );
nor \U$15246 ( \15286 , \15282 , \15285 );
buf \U$15247 ( \15287 , \15286 );
buf \U$15248 ( \15288 , \15287 );
xor \U$15249 ( \15289 , \12568 , \12823 );
and \U$15250 ( \15290 , \15289 , \13134 );
and \U$15251 ( \15291 , \12568 , \12823 );
or \U$15252 ( \15292 , \15290 , \15291 );
buf \U$15253 ( \15293 , \15292 );
buf \U$15254 ( \15294 , \15293 );
not \U$15255 ( \15295 , \15294 );
buf \U$15256 ( \15296 , \15295 );
buf \U$15257 ( \15297 , \15296 );
and \U$15258 ( \15298 , \15288 , \15297 );
not \U$15259 ( \15299 , \15288 );
buf \U$15260 ( \15300 , \15293 );
and \U$15261 ( \15301 , \15299 , \15300 );
nor \U$15262 ( \15302 , \15298 , \15301 );
buf \U$15263 ( \15303 , \15302 );
not \U$15264 ( \15304 , \15303 );
buf \U$15265 ( \15305 , \15304 );
and \U$15266 ( \15306 , \15031 , \15305 );
not \U$15267 ( \15307 , \15031 );
buf \U$15268 ( \15308 , \15303 );
and \U$15269 ( \15309 , \15307 , \15308 );
nor \U$15270 ( \15310 , \15306 , \15309 );
buf \U$15271 ( \15311 , \15310 );
buf \U$15272 ( \15312 , \15311 );
xor \U$15273 ( \15313 , \13368 , \13591 );
and \U$15274 ( \15314 , \15313 , \14243 );
and \U$15275 ( \15315 , \13368 , \13591 );
or \U$15276 ( \15316 , \15314 , \15315 );
buf \U$15277 ( \15317 , \15316 );
buf \U$15278 ( \15318 , \15317 );
not \U$15279 ( \15319 , \15318 );
buf \U$15280 ( \15320 , \13100 );
not \U$15281 ( \15321 , \15320 );
buf \U$15282 ( \15322 , \733 );
not \U$15283 ( \15323 , \15322 );
buf \U$15284 ( \15324 , \745 );
nand \U$15285 ( \15325 , \15323 , \15324 );
buf \U$15286 ( \15326 , \15325 );
buf \U$15287 ( \15327 , \15326 );
not \U$15288 ( \15328 , \15327 );
buf \U$15289 ( \15329 , \15328 );
buf \U$15290 ( \15330 , \15329 );
not \U$15291 ( \15331 , \15330 );
or \U$15292 ( \15332 , \15321 , \15331 );
buf \U$15293 ( \15333 , \734 );
buf \U$15294 ( \15334 , RIc0d8410_30);
buf \U$15295 ( \15335 , RIc0da378_97);
xor \U$15296 ( \15336 , \15334 , \15335 );
buf \U$15297 ( \15337 , \15336 );
buf \U$15298 ( \15338 , \15337 );
nand \U$15299 ( \15339 , \15333 , \15338 );
buf \U$15300 ( \15340 , \15339 );
buf \U$15301 ( \15341 , \15340 );
nand \U$15302 ( \15342 , \15332 , \15341 );
buf \U$15303 ( \15343 , \15342 );
buf \U$15304 ( \15344 , \13010 );
not \U$15305 ( \15345 , \15344 );
buf \U$15306 ( \15346 , \13001 );
not \U$15307 ( \15347 , \15346 );
or \U$15308 ( \15348 , \15345 , \15347 );
buf \U$15309 ( \15349 , \13005 );
buf \U$15310 ( \15350 , RIc0d79c0_8);
buf \U$15311 ( \15351 , RIc0dadc8_119);
xor \U$15312 ( \15352 , \15350 , \15351 );
buf \U$15313 ( \15353 , \15352 );
buf \U$15314 ( \15354 , \15353 );
nand \U$15315 ( \15355 , \15349 , \15354 );
buf \U$15316 ( \15356 , \15355 );
buf \U$15317 ( \15357 , \15356 );
nand \U$15318 ( \15358 , \15348 , \15357 );
buf \U$15319 ( \15359 , \15358 );
buf \U$15320 ( \15360 , \15359 );
not \U$15321 ( \15361 , \15360 );
buf \U$15322 ( \15362 , \15361 );
and \U$15323 ( \15363 , \15343 , \15362 );
not \U$15324 ( \15364 , \15343 );
and \U$15325 ( \15365 , \15364 , \15359 );
or \U$15326 ( \15366 , \15363 , \15365 );
buf \U$15327 ( \15367 , \15366 );
buf \U$15328 ( \15368 , \13080 );
not \U$15329 ( \15369 , \15368 );
buf \U$15330 ( \15370 , \14532 );
not \U$15331 ( \15371 , \15370 );
or \U$15332 ( \15372 , \15369 , \15371 );
buf \U$15333 ( \15373 , \1078 );
xor \U$15334 ( \15374 , RIc0d9bf8_81, RIc0d8b90_46);
buf \U$15335 ( \15375 , \15374 );
nand \U$15336 ( \15376 , \15373 , \15375 );
buf \U$15337 ( \15377 , \15376 );
buf \U$15338 ( \15378 , \15377 );
nand \U$15339 ( \15379 , \15372 , \15378 );
buf \U$15340 ( \15380 , \15379 );
buf \U$15341 ( \15381 , \15380 );
not \U$15342 ( \15382 , \15381 );
buf \U$15343 ( \15383 , \15382 );
buf \U$15344 ( \15384 , \15383 );
and \U$15345 ( \15385 , \15367 , \15384 );
not \U$15346 ( \15386 , \15367 );
buf \U$15347 ( \15387 , \15380 );
and \U$15348 ( \15388 , \15386 , \15387 );
nor \U$15349 ( \15389 , \15385 , \15388 );
buf \U$15350 ( \15390 , \15389 );
buf \U$15351 ( \15391 , \15390 );
not \U$15352 ( \15392 , \15391 );
buf \U$15353 ( \15393 , \13053 );
not \U$15354 ( \15394 , \15393 );
buf \U$15355 ( \15395 , \4482 );
not \U$15356 ( \15396 , \15395 );
buf \U$15357 ( \15397 , \15396 );
buf \U$15358 ( \15398 , \15397 );
not \U$15359 ( \15399 , \15398 );
or \U$15360 ( \15400 , \15394 , \15399 );
buf \U$15361 ( \15401 , \4475 );
not \U$15362 ( \15402 , \15401 );
buf \U$15363 ( \15403 , \15402 );
buf \U$15364 ( \15404 , \15403 );
buf \U$15365 ( \15405 , RIc0d8140_24);
buf \U$15366 ( \15406 , RIc0da648_103);
xor \U$15367 ( \15407 , \15405 , \15406 );
buf \U$15368 ( \15408 , \15407 );
buf \U$15369 ( \15409 , \15408 );
nand \U$15370 ( \15410 , \15404 , \15409 );
buf \U$15371 ( \15411 , \15410 );
buf \U$15372 ( \15412 , \15411 );
nand \U$15373 ( \15413 , \15400 , \15412 );
buf \U$15374 ( \15414 , \15413 );
buf \U$15375 ( \15415 , \15414 );
buf \U$15376 ( \15416 , \12980 );
not \U$15377 ( \15417 , \15416 );
buf \U$15378 ( \15418 , \12968 );
not \U$15379 ( \15419 , \15418 );
buf \U$15380 ( \15420 , \15419 );
buf \U$15381 ( \15421 , \15420 );
not \U$15382 ( \15422 , \15421 );
or \U$15383 ( \15423 , \15417 , \15422 );
buf \U$15384 ( \15424 , \13314 );
xor \U$15385 ( \15425 , RIc0daeb8_121, RIc0d78d0_6);
buf \U$15386 ( \15426 , \15425 );
nand \U$15387 ( \15427 , \15424 , \15426 );
buf \U$15388 ( \15428 , \15427 );
buf \U$15389 ( \15429 , \15428 );
nand \U$15390 ( \15430 , \15423 , \15429 );
buf \U$15391 ( \15431 , \15430 );
buf \U$15392 ( \15432 , \15431 );
xor \U$15393 ( \15433 , \15415 , \15432 );
buf \U$15394 ( \15434 , \12768 );
not \U$15395 ( \15435 , \15434 );
buf \U$15396 ( \15436 , \1183 );
not \U$15397 ( \15437 , \15436 );
or \U$15398 ( \15438 , \15435 , \15437 );
buf \U$15399 ( \15439 , \14374 );
xor \U$15400 ( \15440 , RIc0d9a18_77, RIc0d8d70_50);
buf \U$15401 ( \15441 , \15440 );
nand \U$15402 ( \15442 , \15439 , \15441 );
buf \U$15403 ( \15443 , \15442 );
buf \U$15404 ( \15444 , \15443 );
nand \U$15405 ( \15445 , \15438 , \15444 );
buf \U$15406 ( \15446 , \15445 );
buf \U$15407 ( \15447 , \15446 );
xor \U$15408 ( \15448 , \15433 , \15447 );
buf \U$15409 ( \15449 , \15448 );
buf \U$15410 ( \15450 , \15449 );
not \U$15411 ( \15451 , \15450 );
or \U$15412 ( \15452 , \15392 , \15451 );
buf \U$15413 ( \15453 , \15390 );
buf \U$15414 ( \15454 , \15449 );
or \U$15415 ( \15455 , \15453 , \15454 );
nand \U$15416 ( \15456 , \15452 , \15455 );
buf \U$15417 ( \15457 , \15456 );
buf \U$15418 ( \15458 , \15457 );
buf \U$15419 ( \15459 , \12688 );
not \U$15420 ( \15460 , \15459 );
buf \U$15421 ( \15461 , \12676 );
not \U$15422 ( \15462 , \15461 );
or \U$15423 ( \15463 , \15460 , \15462 );
buf \U$15424 ( \15464 , \2927 );
buf \U$15425 ( \15465 , RIc0d9040_56);
buf \U$15426 ( \15466 , RIc0d9748_71);
xor \U$15427 ( \15467 , \15465 , \15466 );
buf \U$15428 ( \15468 , \15467 );
buf \U$15429 ( \15469 , \15468 );
nand \U$15430 ( \15470 , \15464 , \15469 );
buf \U$15431 ( \15471 , \15470 );
buf \U$15432 ( \15472 , \15471 );
nand \U$15433 ( \15473 , \15463 , \15472 );
buf \U$15434 ( \15474 , \15473 );
buf \U$15435 ( \15475 , \15474 );
buf \U$15436 ( \15476 , \12710 );
not \U$15437 ( \15477 , \15476 );
buf \U$15438 ( \15478 , \330 );
not \U$15439 ( \15479 , \15478 );
or \U$15440 ( \15480 , \15477 , \15479 );
buf \U$15441 ( \15481 , \344 );
buf \U$15442 ( \15482 , RIc0da288_95);
buf \U$15443 ( \15483 , RIc0d8500_32);
xor \U$15444 ( \15484 , \15482 , \15483 );
buf \U$15445 ( \15485 , \15484 );
buf \U$15446 ( \15486 , \15485 );
nand \U$15447 ( \15487 , \15481 , \15486 );
buf \U$15448 ( \15488 , \15487 );
buf \U$15449 ( \15489 , \15488 );
nand \U$15450 ( \15490 , \15480 , \15489 );
buf \U$15451 ( \15491 , \15490 );
buf \U$15452 ( \15492 , \15491 );
xor \U$15453 ( \15493 , \15475 , \15492 );
buf \U$15454 ( \15494 , \1739 );
buf \U$15455 ( \15495 , \12259 );
not \U$15456 ( \15496 , \15495 );
buf \U$15457 ( \15497 , \15496 );
buf \U$15458 ( \15498 , \15497 );
or \U$15459 ( \15499 , \15494 , \15498 );
buf \U$15460 ( \15500 , \996 );
buf \U$15461 ( \15501 , RIc0d8aa0_44);
buf \U$15462 ( \15502 , RIc0d9ce8_83);
xor \U$15463 ( \15503 , \15501 , \15502 );
buf \U$15464 ( \15504 , \15503 );
buf \U$15465 ( \15505 , \15504 );
not \U$15466 ( \15506 , \15505 );
buf \U$15467 ( \15507 , \15506 );
buf \U$15468 ( \15508 , \15507 );
or \U$15469 ( \15509 , \15500 , \15508 );
nand \U$15470 ( \15510 , \15499 , \15509 );
buf \U$15471 ( \15511 , \15510 );
buf \U$15472 ( \15512 , \15511 );
xor \U$15473 ( \15513 , \15493 , \15512 );
buf \U$15474 ( \15514 , \15513 );
buf \U$15475 ( \15515 , \15514 );
not \U$15476 ( \15516 , \15515 );
buf \U$15477 ( \15517 , \15516 );
buf \U$15478 ( \15518 , \15517 );
and \U$15479 ( \15519 , \15458 , \15518 );
not \U$15480 ( \15520 , \15458 );
buf \U$15481 ( \15521 , \15514 );
and \U$15482 ( \15522 , \15520 , \15521 );
nor \U$15483 ( \15523 , \15519 , \15522 );
buf \U$15484 ( \15524 , \15523 );
buf \U$15485 ( \15525 , \15524 );
not \U$15486 ( \15526 , \15525 );
buf \U$15487 ( \15527 , \12942 );
not \U$15488 ( \15528 , \15527 );
buf \U$15489 ( \15529 , \13684 );
not \U$15490 ( \15530 , \15529 );
or \U$15491 ( \15531 , \15528 , \15530 );
buf \U$15492 ( \15532 , \12937 );
buf \U$15493 ( \15533 , RIc0d7ab0_10);
buf \U$15494 ( \15534 , RIc0dacd8_117);
xor \U$15495 ( \15535 , \15533 , \15534 );
buf \U$15496 ( \15536 , \15535 );
buf \U$15497 ( \15537 , \15536 );
nand \U$15498 ( \15538 , \15532 , \15537 );
buf \U$15499 ( \15539 , \15538 );
buf \U$15500 ( \15540 , \15539 );
nand \U$15501 ( \15541 , \15531 , \15540 );
buf \U$15502 ( \15542 , \15541 );
buf \U$15503 ( \15543 , \15542 );
not \U$15504 ( \15544 , \15543 );
buf \U$15505 ( \15545 , \12844 );
not \U$15506 ( \15546 , \15545 );
buf \U$15507 ( \15547 , \4042 );
not \U$15508 ( \15548 , \15547 );
or \U$15509 ( \15549 , \15546 , \15548 );
buf \U$15512 ( \15550 , \3515 );
buf \U$15513 ( \15551 , \15550 );
buf \U$15514 ( \15552 , RIc0d8230_26);
buf \U$15515 ( \15553 , RIc0da558_101);
xor \U$15516 ( \15554 , \15552 , \15553 );
buf \U$15517 ( \15555 , \15554 );
buf \U$15518 ( \15556 , \15555 );
nand \U$15519 ( \15557 , \15551 , \15556 );
buf \U$15520 ( \15558 , \15557 );
buf \U$15521 ( \15559 , \15558 );
nand \U$15522 ( \15560 , \15549 , \15559 );
buf \U$15523 ( \15561 , \15560 );
buf \U$15524 ( \15562 , \15561 );
not \U$15525 ( \15563 , \15562 );
buf \U$15526 ( \15564 , \15563 );
buf \U$15527 ( \15565 , \15564 );
not \U$15528 ( \15566 , \15565 );
or \U$15529 ( \15567 , \15544 , \15566 );
buf \U$15530 ( \15568 , \15542 );
buf \U$15531 ( \15569 , \15564 );
or \U$15532 ( \15570 , \15568 , \15569 );
nand \U$15533 ( \15571 , \15567 , \15570 );
buf \U$15534 ( \15572 , \15571 );
buf \U$15535 ( \15573 , \15572 );
buf \U$15536 ( \15574 , \13499 );
not \U$15537 ( \15575 , \15574 );
buf \U$15538 ( \15576 , \841 );
not \U$15539 ( \15577 , \15576 );
or \U$15540 ( \15578 , \15575 , \15577 );
buf \U$15541 ( \15579 , \442 );
buf \U$15542 ( \15580 , RIc0d87d0_38);
buf \U$15543 ( \15581 , RIc0d9fb8_89);
xor \U$15544 ( \15582 , \15580 , \15581 );
buf \U$15545 ( \15583 , \15582 );
buf \U$15546 ( \15584 , \15583 );
nand \U$15547 ( \15585 , \15579 , \15584 );
buf \U$15548 ( \15586 , \15585 );
buf \U$15549 ( \15587 , \15586 );
nand \U$15550 ( \15588 , \15578 , \15587 );
buf \U$15551 ( \15589 , \15588 );
buf \U$15552 ( \15590 , \15589 );
not \U$15553 ( \15591 , \15590 );
buf \U$15554 ( \15592 , \15591 );
buf \U$15555 ( \15593 , \15592 );
and \U$15556 ( \15594 , \15573 , \15593 );
not \U$15557 ( \15595 , \15573 );
buf \U$15558 ( \15596 , \15589 );
and \U$15559 ( \15597 , \15595 , \15596 );
nor \U$15560 ( \15598 , \15594 , \15597 );
buf \U$15561 ( \15599 , \15598 );
buf \U$15562 ( \15600 , \15599 );
not \U$15563 ( \15601 , \15600 );
buf \U$15564 ( \15602 , \12661 );
not \U$15565 ( \15603 , \15602 );
buf \U$15566 ( \15604 , RIc0db188_127);
not \U$15567 ( \15605 , \15604 );
buf \U$15568 ( \15606 , RIc0db200_128);
nor \U$15569 ( \15607 , \15605 , \15606 );
buf \U$15570 ( \15608 , \15607 );
buf \U$15571 ( \15609 , \15608 );
buf \U$15572 ( \15610 , \15609 );
not \U$15573 ( \15611 , \15610 );
or \U$15574 ( \15612 , \15603 , \15611 );
buf \U$15575 ( \15613 , RIc0db188_127);
buf \U$15576 ( \15614 , RIc0db200_128);
nand \U$15577 ( \15615 , \15613 , \15614 );
buf \U$15578 ( \15616 , \15615 );
buf \U$15579 ( \15617 , \15616 );
nand \U$15580 ( \15618 , \15612 , \15617 );
buf \U$15581 ( \15619 , \15618 );
buf \U$15582 ( \15620 , \15619 );
buf \U$15583 ( \15621 , \12803 );
not \U$15584 ( \15622 , \15621 );
buf \U$15585 ( \15623 , \3780 );
not \U$15586 ( \15624 , \15623 );
or \U$15587 ( \15625 , \15622 , \15624 );
buf \U$15588 ( \15626 , \1229 );
buf \U$15589 ( \15627 , RIc0d9478_65);
buf \U$15590 ( \15628 , RIc0d9310_62);
xor \U$15591 ( \15629 , \15627 , \15628 );
buf \U$15592 ( \15630 , \15629 );
buf \U$15593 ( \15631 , \15630 );
nand \U$15594 ( \15632 , \15626 , \15631 );
buf \U$15595 ( \15633 , \15632 );
buf \U$15596 ( \15634 , \15633 );
nand \U$15597 ( \15635 , \15625 , \15634 );
buf \U$15598 ( \15636 , \15635 );
buf \U$15599 ( \15637 , \15636 );
xor \U$15600 ( \15638 , \15620 , \15637 );
buf \U$15601 ( \15639 , \12749 );
not \U$15602 ( \15640 , \15639 );
not \U$15603 ( \15641 , \12731 );
xor \U$15604 ( \15642 , RIc0da828_107, RIc0da7b0_106);
nor \U$15605 ( \15643 , \15641 , \15642 );
buf \U$15606 ( \15644 , \15643 );
buf \U$15607 ( \15645 , \15644 );
not \U$15608 ( \15646 , \15645 );
or \U$15609 ( \15647 , \15640 , \15646 );
buf \U$15610 ( \15648 , \12743 );
not \U$15611 ( \15649 , \15648 );
buf \U$15612 ( \15650 , \15649 );
buf \U$15613 ( \15651 , \15650 );
not \U$15614 ( \15652 , \15651 );
buf \U$15615 ( \15653 , \15652 );
buf \U$15616 ( \15654 , \15653 );
buf \U$15617 ( \15655 , RIc0d8050_22);
buf \U$15618 ( \15656 , RIc0da738_105);
xor \U$15619 ( \15657 , \15655 , \15656 );
buf \U$15620 ( \15658 , \15657 );
buf \U$15621 ( \15659 , \15658 );
nand \U$15622 ( \15660 , \15654 , \15659 );
buf \U$15623 ( \15661 , \15660 );
buf \U$15624 ( \15662 , \15661 );
nand \U$15625 ( \15663 , \15647 , \15662 );
buf \U$15626 ( \15664 , \15663 );
buf \U$15627 ( \15665 , \15664 );
xor \U$15628 ( \15666 , \15638 , \15665 );
buf \U$15629 ( \15667 , \15666 );
buf \U$15630 ( \15668 , \15667 );
not \U$15631 ( \15669 , \15668 );
or \U$15632 ( \15670 , \15601 , \15669 );
buf \U$15633 ( \15671 , \15667 );
buf \U$15634 ( \15672 , \15599 );
or \U$15635 ( \15673 , \15671 , \15672 );
nand \U$15636 ( \15674 , \15670 , \15673 );
buf \U$15637 ( \15675 , \15674 );
buf \U$15638 ( \15676 , \15675 );
buf \U$15639 ( \15677 , \12415 );
not \U$15640 ( \15678 , \15677 );
buf \U$15641 ( \15679 , \12402 );
not \U$15642 ( \15680 , \15679 );
or \U$15643 ( \15681 , \15678 , \15680 );
buf \U$15644 ( \15682 , \14405 );
buf \U$15645 ( \15683 , RIc0d7c90_14);
buf \U$15646 ( \15684 , RIc0daaf8_113);
xor \U$15647 ( \15685 , \15683 , \15684 );
buf \U$15648 ( \15686 , \15685 );
buf \U$15649 ( \15687 , \15686 );
nand \U$15650 ( \15688 , \15682 , \15687 );
buf \U$15651 ( \15689 , \15688 );
buf \U$15652 ( \15690 , \15689 );
nand \U$15653 ( \15691 , \15681 , \15690 );
buf \U$15654 ( \15692 , \15691 );
buf \U$15655 ( \15693 , \12610 );
not \U$15656 ( \15694 , \15693 );
buf \U$15657 ( \15695 , \3415 );
not \U$15658 ( \15696 , \15695 );
or \U$15659 ( \15697 , \15694 , \15696 );
buf \U$15660 ( \15698 , \481 );
buf \U$15661 ( \15699 , RIc0d85f0_34);
buf \U$15662 ( \15700 , RIc0da198_93);
xor \U$15663 ( \15701 , \15699 , \15700 );
buf \U$15664 ( \15702 , \15701 );
buf \U$15665 ( \15703 , \15702 );
nand \U$15666 ( \15704 , \15698 , \15703 );
buf \U$15667 ( \15705 , \15704 );
buf \U$15668 ( \15706 , \15705 );
nand \U$15669 ( \15707 , \15697 , \15706 );
buf \U$15670 ( \15708 , \15707 );
xor \U$15671 ( \15709 , \15692 , \15708 );
buf \U$15672 ( \15710 , \12447 );
not \U$15673 ( \15711 , \15710 );
buf \U$15674 ( \15712 , \14075 );
not \U$15675 ( \15713 , \15712 );
or \U$15676 ( \15714 , \15711 , \15713 );
buf \U$15677 ( \15715 , \791 );
xor \U$15678 ( \15716 , RIc0d9838_73, RIc0d8f50_54);
buf \U$15679 ( \15717 , \15716 );
nand \U$15680 ( \15718 , \15715 , \15717 );
buf \U$15681 ( \15719 , \15718 );
buf \U$15682 ( \15720 , \15719 );
nand \U$15683 ( \15721 , \15714 , \15720 );
buf \U$15684 ( \15722 , \15721 );
xnor \U$15685 ( \15723 , \15709 , \15722 );
buf \U$15686 ( \15724 , \15723 );
not \U$15687 ( \15725 , \15724 );
buf \U$15688 ( \15726 , \15725 );
buf \U$15689 ( \15727 , \15726 );
and \U$15690 ( \15728 , \15676 , \15727 );
not \U$15691 ( \15729 , \15676 );
buf \U$15692 ( \15730 , \15723 );
and \U$15693 ( \15731 , \15729 , \15730 );
nor \U$15694 ( \15732 , \15728 , \15731 );
buf \U$15695 ( \15733 , \15732 );
buf \U$15696 ( \15734 , \15733 );
not \U$15697 ( \15735 , \15734 );
or \U$15698 ( \15736 , \15526 , \15735 );
buf \U$15699 ( \15737 , \15733 );
buf \U$15700 ( \15738 , \15524 );
or \U$15701 ( \15739 , \15737 , \15738 );
nand \U$15702 ( \15740 , \15736 , \15739 );
buf \U$15703 ( \15741 , \15740 );
buf \U$15704 ( \15742 , \15741 );
buf \U$15705 ( \15743 , \12471 );
not \U$15706 ( \15744 , \15743 );
buf \U$15707 ( \15745 , \13332 );
not \U$15708 ( \15746 , \15745 );
or \U$15709 ( \15747 , \15744 , \15746 );
buf \U$15710 ( \15748 , \874 );
buf \U$15711 ( \15749 , RIc0d9130_58);
buf \U$15712 ( \15750 , RIc0d9658_69);
xor \U$15713 ( \15751 , \15749 , \15750 );
buf \U$15714 ( \15752 , \15751 );
buf \U$15715 ( \15753 , \15752 );
nand \U$15716 ( \15754 , \15748 , \15753 );
buf \U$15717 ( \15755 , \15754 );
buf \U$15718 ( \15756 , \15755 );
nand \U$15719 ( \15757 , \15747 , \15756 );
buf \U$15720 ( \15758 , \15757 );
buf \U$15721 ( \15759 , \15758 );
not \U$15722 ( \15760 , \15759 );
buf \U$15723 ( \15761 , \15760 );
buf \U$15724 ( \15762 , \15761 );
not \U$15725 ( \15763 , \15762 );
buf \U$15726 ( \15764 , \13394 );
not \U$15727 ( \15765 , \15764 );
buf \U$15728 ( \15766 , \2358 );
not \U$15729 ( \15767 , \15766 );
or \U$15730 ( \15768 , \15765 , \15767 );
buf \U$15731 ( \15769 , \1143 );
buf \U$15732 ( \15770 , RIc0d8e60_52);
buf \U$15733 ( \15771 , RIc0d9928_75);
xor \U$15734 ( \15772 , \15770 , \15771 );
buf \U$15735 ( \15773 , \15772 );
buf \U$15736 ( \15774 , \15773 );
nand \U$15737 ( \15775 , \15769 , \15774 );
buf \U$15738 ( \15776 , \15775 );
buf \U$15739 ( \15777 , \15776 );
nand \U$15740 ( \15778 , \15768 , \15777 );
buf \U$15741 ( \15779 , \15778 );
buf \U$15742 ( \15780 , \15779 );
not \U$15743 ( \15781 , \15780 );
buf \U$15744 ( \15782 , \15781 );
buf \U$15745 ( \15783 , \15782 );
not \U$15746 ( \15784 , \15783 );
buf \U$15747 ( \15785 , \13470 );
not \U$15748 ( \15786 , \15785 );
buf \U$15749 ( \15787 , \13457 );
not \U$15750 ( \15788 , \15787 );
buf \U$15751 ( \15789 , \15788 );
buf \U$15752 ( \15790 , \15789 );
not \U$15753 ( \15791 , \15790 );
or \U$15754 ( \15792 , \15786 , \15791 );
buf \U$15757 ( \15793 , \13449 );
buf \U$15758 ( \15794 , \15793 );
buf \U$15759 ( \15795 , RIc0d76f0_2);
buf \U$15760 ( \15796 , RIc0db098_125);
xor \U$15761 ( \15797 , \15795 , \15796 );
buf \U$15762 ( \15798 , \15797 );
buf \U$15763 ( \15799 , \15798 );
nand \U$15764 ( \15800 , \15794 , \15799 );
buf \U$15765 ( \15801 , \15800 );
buf \U$15766 ( \15802 , \15801 );
nand \U$15767 ( \15803 , \15792 , \15802 );
buf \U$15768 ( \15804 , \15803 );
buf \U$15769 ( \15805 , \15804 );
not \U$15770 ( \15806 , \15805 );
or \U$15771 ( \15807 , \15784 , \15806 );
buf \U$15772 ( \15808 , \15804 );
buf \U$15773 ( \15809 , \15782 );
or \U$15774 ( \15810 , \15808 , \15809 );
nand \U$15775 ( \15811 , \15807 , \15810 );
buf \U$15776 ( \15812 , \15811 );
buf \U$15777 ( \15813 , \15812 );
not \U$15778 ( \15814 , \15813 );
or \U$15779 ( \15815 , \15763 , \15814 );
buf \U$15780 ( \15816 , \15812 );
buf \U$15781 ( \15817 , \15761 );
or \U$15782 ( \15818 , \15816 , \15817 );
nand \U$15783 ( \15819 , \15815 , \15818 );
buf \U$15784 ( \15820 , \15819 );
buf \U$15785 ( \15821 , \15820 );
buf \U$15786 ( \15822 , \12493 );
not \U$15787 ( \15823 , \15822 );
buf \U$15788 ( \15824 , \2399 );
not \U$15789 ( \15825 , \15824 );
or \U$15790 ( \15826 , \15823 , \15825 );
buf \U$15791 ( \15827 , \2960 );
buf \U$15792 ( \15828 , RIc0d89b0_42);
buf \U$15793 ( \15829 , RIc0d9dd8_85);
xor \U$15794 ( \15830 , \15828 , \15829 );
buf \U$15795 ( \15831 , \15830 );
buf \U$15796 ( \15832 , \15831 );
nand \U$15797 ( \15833 , \15827 , \15832 );
buf \U$15798 ( \15834 , \15833 );
buf \U$15799 ( \15835 , \15834 );
nand \U$15800 ( \15836 , \15826 , \15835 );
buf \U$15801 ( \15837 , \15836 );
buf \U$15802 ( \15838 , \15837 );
buf \U$15803 ( \15839 , \12366 );
not \U$15804 ( \15840 , \15839 );
buf \U$15805 ( \15841 , \396 );
not \U$15806 ( \15842 , \15841 );
or \U$15807 ( \15843 , \15840 , \15842 );
buf \U$15808 ( \15844 , \403 );
buf \U$15809 ( \15845 , RIc0d8c80_48);
buf \U$15810 ( \15846 , RIc0d9b08_79);
xor \U$15811 ( \15847 , \15845 , \15846 );
buf \U$15812 ( \15848 , \15847 );
buf \U$15813 ( \15849 , \15848 );
nand \U$15814 ( \15850 , \15844 , \15849 );
buf \U$15815 ( \15851 , \15850 );
buf \U$15816 ( \15852 , \15851 );
nand \U$15817 ( \15853 , \15843 , \15852 );
buf \U$15818 ( \15854 , \15853 );
buf \U$15819 ( \15855 , \15854 );
xor \U$15820 ( \15856 , \15838 , \15855 );
buf \U$15821 ( \15857 , \12546 );
not \U$15822 ( \15858 , \15857 );
buf \U$15823 ( \15859 , \12529 );
not \U$15824 ( \15860 , \15859 );
or \U$15825 ( \15861 , \15858 , \15860 );
buf \U$15826 ( \15862 , \12541 );
not \U$15827 ( \15863 , \15862 );
buf \U$15828 ( \15864 , \15863 );
buf \U$15829 ( \15865 , \15864 );
buf \U$15830 ( \15866 , RIc0d7d80_16);
buf \U$15831 ( \15867 , RIc0daa08_111);
xor \U$15832 ( \15868 , \15866 , \15867 );
buf \U$15833 ( \15869 , \15868 );
buf \U$15834 ( \15870 , \15869 );
nand \U$15835 ( \15871 , \15865 , \15870 );
buf \U$15836 ( \15872 , \15871 );
buf \U$15837 ( \15873 , \15872 );
nand \U$15838 ( \15874 , \15861 , \15873 );
buf \U$15839 ( \15875 , \15874 );
buf \U$15840 ( \15876 , \15875 );
xor \U$15841 ( \15877 , \15856 , \15876 );
buf \U$15842 ( \15878 , \15877 );
buf \U$15843 ( \15879 , \15878 );
xor \U$15844 ( \15880 , \15821 , \15879 );
buf \U$15845 ( \15881 , \12344 );
not \U$15846 ( \15882 , \15881 );
buf \U$15847 ( \15883 , \12334 );
not \U$15848 ( \15884 , \15883 );
or \U$15849 ( \15885 , \15882 , \15884 );
buf \U$15850 ( \15886 , \12342 );
buf \U$15851 ( \15887 , RIc0d7f60_20);
buf \U$15852 ( \15888 , RIc0da828_107);
xor \U$15853 ( \15889 , \15887 , \15888 );
buf \U$15854 ( \15890 , \15889 );
buf \U$15855 ( \15891 , \15890 );
nand \U$15856 ( \15892 , \15886 , \15891 );
buf \U$15857 ( \15893 , \15892 );
buf \U$15858 ( \15894 , \15893 );
nand \U$15859 ( \15895 , \15885 , \15894 );
buf \U$15860 ( \15896 , \15895 );
buf \U$15861 ( \15897 , \15896 );
not \U$15862 ( \15898 , \15897 );
buf \U$15863 ( \15899 , \15898 );
buf \U$15864 ( \15900 , \15899 );
not \U$15865 ( \15901 , \15900 );
buf \U$15866 ( \15902 , \13431 );
not \U$15867 ( \15903 , \15902 );
buf \U$15868 ( \15904 , \14210 );
not \U$15869 ( \15905 , \15904 );
or \U$15870 ( \15906 , \15903 , \15905 );
buf \U$15871 ( \15907 , \13423 );
not \U$15872 ( \15908 , \15907 );
buf \U$15873 ( \15909 , \15908 );
buf \U$15874 ( \15910 , \15909 );
buf \U$15875 ( \15911 , RIc0da918_109);
buf \U$15876 ( \15912 , RIc0d7e70_18);
xor \U$15877 ( \15913 , \15911 , \15912 );
buf \U$15878 ( \15914 , \15913 );
buf \U$15879 ( \15915 , \15914 );
nand \U$15880 ( \15916 , \15910 , \15915 );
buf \U$15881 ( \15917 , \15916 );
buf \U$15882 ( \15918 , \15917 );
nand \U$15883 ( \15919 , \15906 , \15918 );
buf \U$15884 ( \15920 , \15919 );
buf \U$15885 ( \15921 , \15920 );
not \U$15886 ( \15922 , \15921 );
or \U$15887 ( \15923 , \15901 , \15922 );
buf \U$15888 ( \15924 , \15920 );
buf \U$15889 ( \15925 , \15899 );
or \U$15890 ( \15926 , \15924 , \15925 );
nand \U$15891 ( \15927 , \15923 , \15926 );
buf \U$15892 ( \15928 , \15927 );
buf \U$15893 ( \15929 , \15928 );
buf \U$15894 ( \15930 , RIc0d7ba0_12);
buf \U$15895 ( \15931 , RIc0dabe8_115);
xor \U$15896 ( \15932 , \15930 , \15931 );
buf \U$15897 ( \15933 , \15932 );
and \U$15898 ( \15934 , \12303 , \15933 );
not \U$15899 ( \15935 , \12308 );
nor \U$15900 ( \15936 , \15935 , \14681 );
nor \U$15901 ( \15937 , \15934 , \15936 );
buf \U$15902 ( \15938 , \15937 );
not \U$15903 ( \15939 , \15938 );
buf \U$15904 ( \15940 , \15939 );
buf \U$15905 ( \15941 , \15940 );
and \U$15906 ( \15942 , \15929 , \15941 );
not \U$15907 ( \15943 , \15929 );
buf \U$15908 ( \15944 , \15937 );
and \U$15909 ( \15945 , \15943 , \15944 );
nor \U$15910 ( \15946 , \15942 , \15945 );
buf \U$15911 ( \15947 , \15946 );
buf \U$15912 ( \15948 , \15947 );
xnor \U$15913 ( \15949 , \15880 , \15948 );
buf \U$15914 ( \15950 , \15949 );
buf \U$15915 ( \15951 , \15950 );
and \U$15916 ( \15952 , \15742 , \15951 );
not \U$15917 ( \15953 , \15742 );
buf \U$15918 ( \15954 , \15950 );
not \U$15919 ( \15955 , \15954 );
buf \U$15920 ( \15956 , \15955 );
buf \U$15921 ( \15957 , \15956 );
and \U$15922 ( \15958 , \15953 , \15957 );
nor \U$15923 ( \15959 , \15952 , \15958 );
buf \U$15924 ( \15960 , \15959 );
buf \U$15925 ( \15961 , \15960 );
not \U$15926 ( \15962 , \15961 );
and \U$15927 ( \15963 , \15319 , \15962 );
buf \U$15928 ( \15964 , \15317 );
buf \U$15929 ( \15965 , \15960 );
and \U$15930 ( \15966 , \15964 , \15965 );
nor \U$15931 ( \15967 , \15963 , \15966 );
buf \U$15932 ( \15968 , \15967 );
buf \U$15933 ( \15969 , \15968 );
xor \U$15934 ( \15970 , RIc0d9b08_79, RIc0d8e60_52);
buf \U$15935 ( \15971 , \15970 );
not \U$15936 ( \15972 , \15971 );
buf \U$15937 ( \15973 , \12361 );
not \U$15938 ( \15974 , \15973 );
or \U$15939 ( \15975 , \15972 , \15974 );
buf \U$15940 ( \15976 , \3985 );
xor \U$15941 ( \15977 , RIc0d9b08_79, RIc0d8de8_51);
buf \U$15942 ( \15978 , \15977 );
nand \U$15943 ( \15979 , \15976 , \15978 );
buf \U$15944 ( \15980 , \15979 );
buf \U$15945 ( \15981 , \15980 );
nand \U$15946 ( \15982 , \15975 , \15981 );
buf \U$15947 ( \15983 , \15982 );
buf \U$15948 ( \15984 , \15983 );
not \U$15949 ( \15985 , \15984 );
xor \U$15950 ( \15986 , RIc0da198_93, RIc0d87d0_38);
buf \U$15951 ( \15987 , \15986 );
not \U$15952 ( \15988 , \15987 );
buf \U$15953 ( \15989 , \467 );
buf \U$15954 ( \15990 , \469 );
nand \U$15955 ( \15991 , \15989 , \15990 );
buf \U$15956 ( \15992 , \15991 );
buf \U$15957 ( \15993 , \15992 );
not \U$15958 ( \15994 , \15993 );
buf \U$15959 ( \15995 , \15994 );
buf \U$15960 ( \15996 , \15995 );
not \U$15961 ( \15997 , \15996 );
or \U$15962 ( \15998 , \15988 , \15997 );
buf \U$15963 ( \15999 , \4008 );
buf \U$15964 ( \16000 , \13564 );
nand \U$15965 ( \16001 , \15999 , \16000 );
buf \U$15966 ( \16002 , \16001 );
buf \U$15967 ( \16003 , \16002 );
nand \U$15968 ( \16004 , \15998 , \16003 );
buf \U$15969 ( \16005 , \16004 );
buf \U$15970 ( \16006 , \16005 );
not \U$15971 ( \16007 , \16006 );
or \U$15972 ( \16008 , \15985 , \16007 );
buf \U$15973 ( \16009 , \16005 );
buf \U$15974 ( \16010 , \15983 );
or \U$15975 ( \16011 , \16009 , \16010 );
buf \U$15976 ( \16012 , \13928 );
not \U$15977 ( \16013 , \16012 );
buf \U$15978 ( \16014 , \15643 );
buf \U$15979 ( \16015 , \16014 );
not \U$15980 ( \16016 , \16015 );
or \U$15981 ( \16017 , \16013 , \16016 );
buf \U$15982 ( \16018 , \12744 );
buf \U$15983 ( \16019 , RIc0d81b8_25);
buf \U$15984 ( \16020 , RIc0da738_105);
xor \U$15985 ( \16021 , \16019 , \16020 );
buf \U$15986 ( \16022 , \16021 );
buf \U$15987 ( \16023 , \16022 );
nand \U$15988 ( \16024 , \16018 , \16023 );
buf \U$15989 ( \16025 , \16024 );
buf \U$15990 ( \16026 , \16025 );
nand \U$15991 ( \16027 , \16017 , \16026 );
buf \U$15992 ( \16028 , \16027 );
buf \U$15993 ( \16029 , \16028 );
nand \U$15994 ( \16030 , \16011 , \16029 );
buf \U$15995 ( \16031 , \16030 );
buf \U$15996 ( \16032 , \16031 );
nand \U$15997 ( \16033 , \16008 , \16032 );
buf \U$15998 ( \16034 , \16033 );
buf \U$15999 ( \16035 , RIc0d77e0_4);
buf \U$16000 ( \16036 , RIc0db188_127);
xor \U$16001 ( \16037 , \16035 , \16036 );
buf \U$16002 ( \16038 , \16037 );
buf \U$16003 ( \16039 , \16038 );
not \U$16004 ( \16040 , \16039 );
buf \U$16005 ( \16041 , \12654 );
not \U$16006 ( \16042 , \16041 );
or \U$16007 ( \16043 , \16040 , \16042 );
buf \U$16008 ( \16044 , RIc0d7768_3);
buf \U$16009 ( \16045 , RIc0db188_127);
xor \U$16010 ( \16046 , \16044 , \16045 );
buf \U$16011 ( \16047 , \16046 );
buf \U$16012 ( \16048 , \16047 );
buf \U$16013 ( \16049 , RIc0db200_128);
nand \U$16014 ( \16050 , \16048 , \16049 );
buf \U$16015 ( \16051 , \16050 );
buf \U$16016 ( \16052 , \16051 );
nand \U$16017 ( \16053 , \16043 , \16052 );
buf \U$16018 ( \16054 , \16053 );
buf \U$16019 ( \16055 , \16054 );
buf \U$16020 ( \16056 , RIc0d8140_24);
buf \U$16021 ( \16057 , RIc0da828_107);
xor \U$16022 ( \16058 , \16056 , \16057 );
buf \U$16023 ( \16059 , \16058 );
buf \U$16024 ( \16060 , \16059 );
not \U$16025 ( \16061 , \16060 );
buf \U$16026 ( \16062 , \12341 );
not \U$16027 ( \16063 , \16062 );
buf \U$16028 ( \16064 , \16063 );
and \U$16029 ( \16065 , \16064 , \12327 );
buf \U$16030 ( \16066 , \16065 );
not \U$16031 ( \16067 , \16066 );
or \U$16032 ( \16068 , \16061 , \16067 );
buf \U$16033 ( \16069 , \16064 );
not \U$16034 ( \16070 , \16069 );
buf \U$16035 ( \16071 , \16070 );
buf \U$16036 ( \16072 , \16071 );
buf \U$16037 ( \16073 , \13262 );
nand \U$16038 ( \16074 , \16072 , \16073 );
buf \U$16039 ( \16075 , \16074 );
buf \U$16040 ( \16076 , \16075 );
nand \U$16041 ( \16077 , \16068 , \16076 );
buf \U$16042 ( \16078 , \16077 );
buf \U$16043 ( \16079 , \16078 );
xor \U$16044 ( \16080 , \16055 , \16079 );
xor \U$16045 ( \16081 , RIc0da378_97, RIc0d85f0_34);
buf \U$16046 ( \16082 , \16081 );
not \U$16047 ( \16083 , \16082 );
buf \U$16048 ( \16084 , \748 );
not \U$16049 ( \16085 , \16084 );
buf \U$16050 ( \16086 , \16085 );
buf \U$16051 ( \16087 , \16086 );
not \U$16052 ( \16088 , \16087 );
or \U$16053 ( \16089 , \16083 , \16088 );
buf \U$16054 ( \16090 , \734 );
buf \U$16055 ( \16091 , \13243 );
nand \U$16056 ( \16092 , \16090 , \16091 );
buf \U$16057 ( \16093 , \16092 );
buf \U$16058 ( \16094 , \16093 );
nand \U$16059 ( \16095 , \16089 , \16094 );
buf \U$16060 ( \16096 , \16095 );
buf \U$16061 ( \16097 , \16096 );
and \U$16062 ( \16098 , \16080 , \16097 );
and \U$16063 ( \16099 , \16055 , \16079 );
or \U$16064 ( \16100 , \16098 , \16099 );
buf \U$16065 ( \16101 , \16100 );
xor \U$16066 ( \16102 , \16034 , \16101 );
buf \U$16067 ( \16103 , RIc0d9400_64);
buf \U$16068 ( \16104 , RIc0d9568_67);
xor \U$16069 ( \16105 , \16103 , \16104 );
buf \U$16070 ( \16106 , \16105 );
buf \U$16071 ( \16107 , \16106 );
not \U$16072 ( \16108 , \16107 );
buf \U$16073 ( \16109 , \1823 );
not \U$16074 ( \16110 , \16109 );
or \U$16075 ( \16111 , \16108 , \16110 );
buf \U$16076 ( \16112 , \686 );
buf \U$16077 ( \16113 , \13218 );
nand \U$16078 ( \16114 , \16112 , \16113 );
buf \U$16079 ( \16115 , \16114 );
buf \U$16080 ( \16116 , \16115 );
nand \U$16081 ( \16117 , \16111 , \16116 );
buf \U$16082 ( \16118 , \16117 );
buf \U$16083 ( \16119 , \16118 );
not \U$16084 ( \16120 , \16119 );
buf \U$16085 ( \16121 , \16120 );
buf \U$16086 ( \16122 , \16121 );
not \U$16087 ( \16123 , \16122 );
buf \U$16088 ( \16124 , \14083 );
not \U$16089 ( \16125 , \16124 );
buf \U$16090 ( \16126 , \12442 );
not \U$16091 ( \16127 , \16126 );
or \U$16092 ( \16128 , \16125 , \16127 );
buf \U$16093 ( \16129 , \1856 );
buf \U$16094 ( \16130 , RIc0d90b8_57);
buf \U$16095 ( \16131 , RIc0d9838_73);
xor \U$16096 ( \16132 , \16130 , \16131 );
buf \U$16097 ( \16133 , \16132 );
buf \U$16098 ( \16134 , \16133 );
nand \U$16099 ( \16135 , \16129 , \16134 );
buf \U$16100 ( \16136 , \16135 );
buf \U$16101 ( \16137 , \16136 );
nand \U$16102 ( \16138 , \16128 , \16137 );
buf \U$16103 ( \16139 , \16138 );
buf \U$16104 ( \16140 , \16139 );
not \U$16105 ( \16141 , \16140 );
buf \U$16106 ( \16142 , \16141 );
buf \U$16107 ( \16143 , \16142 );
not \U$16108 ( \16144 , \16143 );
or \U$16109 ( \16145 , \16123 , \16144 );
buf \U$16110 ( \16146 , \14479 );
not \U$16111 ( \16147 , \16146 );
buf \U$16112 ( \16148 , \13461 );
not \U$16113 ( \16149 , \16148 );
or \U$16114 ( \16150 , \16147 , \16149 );
buf \U$16115 ( \16151 , \13465 );
buf \U$16116 ( \16152 , RIc0d7858_5);
buf \U$16117 ( \16153 , RIc0db098_125);
xor \U$16118 ( \16154 , \16152 , \16153 );
buf \U$16119 ( \16155 , \16154 );
buf \U$16120 ( \16156 , \16155 );
nand \U$16121 ( \16157 , \16151 , \16156 );
buf \U$16122 ( \16158 , \16157 );
buf \U$16123 ( \16159 , \16158 );
nand \U$16124 ( \16160 , \16150 , \16159 );
buf \U$16125 ( \16161 , \16160 );
buf \U$16126 ( \16162 , \16161 );
nand \U$16127 ( \16163 , \16145 , \16162 );
buf \U$16128 ( \16164 , \16163 );
buf \U$16129 ( \16165 , \16164 );
buf \U$16130 ( \16166 , \16139 );
buf \U$16131 ( \16167 , \16118 );
nand \U$16132 ( \16168 , \16166 , \16167 );
buf \U$16133 ( \16169 , \16168 );
buf \U$16134 ( \16170 , \16169 );
nand \U$16135 ( \16171 , \16165 , \16170 );
buf \U$16136 ( \16172 , \16171 );
xnor \U$16137 ( \16173 , \16102 , \16172 );
buf \U$16138 ( \16174 , \16173 );
not \U$16139 ( \16175 , \16174 );
buf \U$16140 ( \16176 , \16175 );
buf \U$16141 ( \16177 , \16176 );
not \U$16142 ( \16178 , \16177 );
xor \U$16143 ( \16179 , \16055 , \16079 );
xor \U$16144 ( \16180 , \16179 , \16097 );
buf \U$16145 ( \16181 , \16180 );
buf \U$16146 ( \16182 , \16181 );
xor \U$16147 ( \16183 , \16005 , \16028 );
buf \U$16148 ( \16184 , \16183 );
buf \U$16149 ( \16185 , \15983 );
xor \U$16150 ( \16186 , \16184 , \16185 );
buf \U$16151 ( \16187 , \16186 );
buf \U$16152 ( \16188 , \16187 );
xor \U$16153 ( \16189 , \16182 , \16188 );
buf \U$16154 ( \16190 , \13745 );
not \U$16155 ( \16191 , \16190 );
buf \U$16156 ( \16192 , \951 );
not \U$16157 ( \16193 , \16192 );
or \U$16158 ( \16194 , \16191 , \16193 );
buf \U$16159 ( \16195 , \2960 );
buf \U$16160 ( \16196 , RIc0d8b18_45);
buf \U$16161 ( \16197 , RIc0d9dd8_85);
xor \U$16162 ( \16198 , \16196 , \16197 );
buf \U$16163 ( \16199 , \16198 );
buf \U$16164 ( \16200 , \16199 );
nand \U$16165 ( \16201 , \16195 , \16200 );
buf \U$16166 ( \16202 , \16201 );
buf \U$16167 ( \16203 , \16202 );
nand \U$16168 ( \16204 , \16194 , \16203 );
buf \U$16169 ( \16205 , \16204 );
buf \U$16170 ( \16206 , \16205 );
buf \U$16171 ( \16207 , \14191 );
not \U$16172 ( \16208 , \16207 );
buf \U$16173 ( \16209 , \14186 );
not \U$16174 ( \16210 , \16209 );
or \U$16175 ( \16211 , \16208 , \16210 );
buf \U$16176 ( \16212 , \12303 );
buf \U$16177 ( \16213 , RIc0dabe8_115);
buf \U$16178 ( \16214 , RIc0d7d08_15);
xor \U$16179 ( \16215 , \16213 , \16214 );
buf \U$16180 ( \16216 , \16215 );
buf \U$16181 ( \16217 , \16216 );
nand \U$16182 ( \16218 , \16212 , \16217 );
buf \U$16183 ( \16219 , \16218 );
buf \U$16184 ( \16220 , \16219 );
nand \U$16185 ( \16221 , \16211 , \16220 );
buf \U$16186 ( \16222 , \16221 );
buf \U$16187 ( \16223 , \16222 );
xor \U$16188 ( \16224 , \16206 , \16223 );
buf \U$16189 ( \16225 , \14221 );
not \U$16190 ( \16226 , \16225 );
buf \U$16191 ( \16227 , \14210 );
not \U$16192 ( \16228 , \16227 );
or \U$16193 ( \16229 , \16226 , \16228 );
buf \U$16194 ( \16230 , \13423 );
not \U$16195 ( \16231 , \16230 );
buf \U$16196 ( \16232 , \16231 );
buf \U$16197 ( \16233 , \16232 );
buf \U$16198 ( \16234 , RIc0da918_109);
buf \U$16199 ( \16235 , RIc0d7fd8_21);
and \U$16200 ( \16236 , \16234 , \16235 );
not \U$16201 ( \16237 , \16234 );
buf \U$16202 ( \16238 , RIc0d7fd8_21);
not \U$16203 ( \16239 , \16238 );
buf \U$16204 ( \16240 , \16239 );
buf \U$16205 ( \16241 , \16240 );
and \U$16206 ( \16242 , \16237 , \16241 );
nor \U$16207 ( \16243 , \16236 , \16242 );
buf \U$16208 ( \16244 , \16243 );
buf \U$16209 ( \16245 , \16244 );
nand \U$16210 ( \16246 , \16233 , \16245 );
buf \U$16211 ( \16247 , \16246 );
buf \U$16212 ( \16248 , \16247 );
nand \U$16213 ( \16249 , \16229 , \16248 );
buf \U$16214 ( \16250 , \16249 );
buf \U$16215 ( \16251 , \16250 );
xor \U$16216 ( \16252 , \16224 , \16251 );
buf \U$16217 ( \16253 , \16252 );
buf \U$16218 ( \16254 , \16253 );
and \U$16219 ( \16255 , \16189 , \16254 );
and \U$16220 ( \16256 , \16182 , \16188 );
or \U$16221 ( \16257 , \16255 , \16256 );
buf \U$16222 ( \16258 , \16257 );
buf \U$16223 ( \16259 , \16258 );
not \U$16224 ( \16260 , \16259 );
or \U$16225 ( \16261 , \16178 , \16260 );
buf \U$16226 ( \16262 , \16176 );
buf \U$16227 ( \16263 , \16258 );
or \U$16228 ( \16264 , \16262 , \16263 );
xor \U$16229 ( \16265 , RIc0db188_127, RIc0d7858_5);
buf \U$16230 ( \16266 , \16265 );
not \U$16231 ( \16267 , \16266 );
buf \U$16232 ( \16268 , \12654 );
not \U$16233 ( \16269 , \16268 );
or \U$16234 ( \16270 , \16267 , \16269 );
buf \U$16235 ( \16271 , \16038 );
buf \U$16236 ( \16272 , RIc0db200_128);
nand \U$16237 ( \16273 , \16271 , \16272 );
buf \U$16238 ( \16274 , \16273 );
buf \U$16239 ( \16275 , \16274 );
nand \U$16240 ( \16276 , \16270 , \16275 );
buf \U$16241 ( \16277 , \16276 );
buf \U$16242 ( \16278 , \16277 );
buf \U$16243 ( \16279 , RIc0d81b8_25);
buf \U$16244 ( \16280 , RIc0da828_107);
xor \U$16245 ( \16281 , \16279 , \16280 );
buf \U$16246 ( \16282 , \16281 );
buf \U$16247 ( \16283 , \16282 );
not \U$16248 ( \16284 , \16283 );
buf \U$16249 ( \16285 , \16065 );
not \U$16250 ( \16286 , \16285 );
or \U$16251 ( \16287 , \16284 , \16286 );
buf \U$16252 ( \16288 , \12342 );
buf \U$16253 ( \16289 , \16059 );
nand \U$16254 ( \16290 , \16288 , \16289 );
buf \U$16255 ( \16291 , \16290 );
buf \U$16256 ( \16292 , \16291 );
nand \U$16257 ( \16293 , \16287 , \16292 );
buf \U$16258 ( \16294 , \16293 );
buf \U$16259 ( \16295 , \16294 );
xor \U$16260 ( \16296 , \16278 , \16295 );
xor \U$16261 ( \16297 , RIc0da198_93, RIc0d8848_39);
buf \U$16262 ( \16298 , \16297 );
not \U$16263 ( \16299 , \16298 );
buf \U$16264 ( \16300 , \1901 );
not \U$16265 ( \16301 , \16300 );
or \U$16266 ( \16302 , \16299 , \16301 );
buf \U$16267 ( \16303 , \481 );
buf \U$16268 ( \16304 , \15986 );
nand \U$16269 ( \16305 , \16303 , \16304 );
buf \U$16270 ( \16306 , \16305 );
buf \U$16271 ( \16307 , \16306 );
nand \U$16272 ( \16308 , \16302 , \16307 );
buf \U$16273 ( \16309 , \16308 );
buf \U$16274 ( \16310 , \16309 );
and \U$16275 ( \16311 , \16296 , \16310 );
and \U$16276 ( \16312 , \16278 , \16295 );
or \U$16277 ( \16313 , \16311 , \16312 );
buf \U$16278 ( \16314 , \16313 );
buf \U$16279 ( \16315 , \16314 );
buf \U$16280 ( \16316 , \14990 );
not \U$16281 ( \16317 , \16316 );
buf \U$16282 ( \16318 , \12870 );
not \U$16283 ( \16319 , \16318 );
or \U$16284 ( \16320 , \16317 , \16319 );
buf \U$16285 ( \16321 , RIc0d79c0_8);
buf \U$16286 ( \16322 , RIc0dafa8_123);
xnor \U$16287 ( \16323 , \16321 , \16322 );
buf \U$16288 ( \16324 , \16323 );
buf \U$16289 ( \16325 , \16324 );
not \U$16290 ( \16326 , \16325 );
buf \U$16291 ( \16327 , \12877 );
nand \U$16292 ( \16328 , \16326 , \16327 );
buf \U$16293 ( \16329 , \16328 );
buf \U$16294 ( \16330 , \16329 );
nand \U$16295 ( \16331 , \16320 , \16330 );
buf \U$16296 ( \16332 , \16331 );
buf \U$16297 ( \16333 , \16332 );
buf \U$16298 ( \16334 , \14948 );
not \U$16299 ( \16335 , \16334 );
buf \U$16300 ( \16336 , \1021 );
not \U$16301 ( \16337 , \16336 );
or \U$16302 ( \16338 , \16335 , \16337 );
buf \U$16303 ( \16339 , \3985 );
buf \U$16304 ( \16340 , \15970 );
nand \U$16305 ( \16341 , \16339 , \16340 );
buf \U$16306 ( \16342 , \16341 );
buf \U$16307 ( \16343 , \16342 );
nand \U$16308 ( \16344 , \16338 , \16343 );
buf \U$16309 ( \16345 , \16344 );
buf \U$16310 ( \16346 , \16345 );
or \U$16311 ( \16347 , \16333 , \16346 );
buf \U$16312 ( \16348 , \16347 );
not \U$16313 ( \16349 , \16348 );
buf \U$16314 ( \16350 , RIc0d8668_35);
buf \U$16315 ( \16351 , RIc0da378_97);
xor \U$16316 ( \16352 , \16350 , \16351 );
buf \U$16317 ( \16353 , \16352 );
buf \U$16318 ( \16354 , \16353 );
not \U$16319 ( \16355 , \16354 );
buf \U$16320 ( \16356 , \2938 );
not \U$16321 ( \16357 , \16356 );
buf \U$16322 ( \16358 , \16357 );
buf \U$16323 ( \16359 , \16358 );
not \U$16324 ( \16360 , \16359 );
or \U$16325 ( \16361 , \16355 , \16360 );
buf \U$16326 ( \16362 , \734 );
buf \U$16327 ( \16363 , \16081 );
nand \U$16328 ( \16364 , \16362 , \16363 );
buf \U$16329 ( \16365 , \16364 );
buf \U$16330 ( \16366 , \16365 );
nand \U$16331 ( \16367 , \16361 , \16366 );
buf \U$16332 ( \16368 , \16367 );
not \U$16333 ( \16369 , \16368 );
or \U$16334 ( \16370 , \16349 , \16369 );
buf \U$16335 ( \16371 , \16332 );
buf \U$16336 ( \16372 , \16345 );
nand \U$16337 ( \16373 , \16371 , \16372 );
buf \U$16338 ( \16374 , \16373 );
nand \U$16339 ( \16375 , \16370 , \16374 );
buf \U$16340 ( \16376 , \16375 );
xor \U$16341 ( \16377 , \16315 , \16376 );
buf \U$16342 ( \16378 , \13785 );
not \U$16343 ( \16379 , \16378 );
buf \U$16344 ( \16380 , \12968 );
not \U$16345 ( \16381 , \16380 );
buf \U$16346 ( \16382 , \16381 );
buf \U$16347 ( \16383 , \16382 );
not \U$16348 ( \16384 , \16383 );
or \U$16349 ( \16385 , \16379 , \16384 );
buf \U$16352 ( \16386 , \12975 );
buf \U$16353 ( \16387 , \16386 );
buf \U$16354 ( \16388 , \13305 );
nand \U$16355 ( \16389 , \16387 , \16388 );
buf \U$16356 ( \16390 , \16389 );
buf \U$16357 ( \16391 , \16390 );
nand \U$16358 ( \16392 , \16385 , \16391 );
buf \U$16359 ( \16393 , \16392 );
buf \U$16360 ( \16394 , \13895 );
not \U$16361 ( \16395 , \16394 );
buf \U$16362 ( \16396 , \710 );
buf \U$16363 ( \16397 , \517 );
nand \U$16364 ( \16398 , \16396 , \16397 );
buf \U$16365 ( \16399 , \16398 );
buf \U$16366 ( \16400 , \16399 );
not \U$16367 ( \16401 , \16400 );
buf \U$16368 ( \16402 , \16401 );
buf \U$16369 ( \16403 , \16402 );
not \U$16370 ( \16404 , \16403 );
or \U$16371 ( \16405 , \16395 , \16404 );
buf \U$16372 ( \16406 , \533 );
buf \U$16373 ( \16407 , \13287 );
nand \U$16374 ( \16408 , \16406 , \16407 );
buf \U$16375 ( \16409 , \16408 );
buf \U$16376 ( \16410 , \16409 );
nand \U$16377 ( \16411 , \16405 , \16410 );
buf \U$16378 ( \16412 , \16411 );
buf \U$16379 ( \16413 , \16412 );
not \U$16380 ( \16414 , \16413 );
buf \U$16381 ( \16415 , \13644 );
not \U$16382 ( \16416 , \16415 );
buf \U$16383 ( \16417 , \12254 );
not \U$16384 ( \16418 , \16417 );
or \U$16385 ( \16419 , \16416 , \16418 );
buf \U$16386 ( \16420 , \584 );
buf \U$16387 ( \16421 , \13197 );
nand \U$16388 ( \16422 , \16420 , \16421 );
buf \U$16389 ( \16423 , \16422 );
buf \U$16390 ( \16424 , \16423 );
nand \U$16391 ( \16425 , \16419 , \16424 );
buf \U$16392 ( \16426 , \16425 );
buf \U$16393 ( \16427 , \16426 );
not \U$16394 ( \16428 , \16427 );
buf \U$16395 ( \16429 , \16428 );
buf \U$16396 ( \16430 , \16429 );
not \U$16397 ( \16431 , \16430 );
or \U$16398 ( \16432 , \16414 , \16431 );
buf \U$16399 ( \16433 , \16426 );
buf \U$16400 ( \16434 , \16412 );
not \U$16401 ( \16435 , \16434 );
buf \U$16402 ( \16436 , \16435 );
buf \U$16403 ( \16437 , \16436 );
nand \U$16404 ( \16438 , \16433 , \16437 );
buf \U$16405 ( \16439 , \16438 );
buf \U$16406 ( \16440 , \16439 );
nand \U$16407 ( \16441 , \16432 , \16440 );
buf \U$16408 ( \16442 , \16441 );
xor \U$16409 ( \16443 , \16393 , \16442 );
buf \U$16410 ( \16444 , \16443 );
and \U$16411 ( \16445 , \16377 , \16444 );
and \U$16412 ( \16446 , \16315 , \16376 );
or \U$16413 ( \16447 , \16445 , \16446 );
buf \U$16414 ( \16448 , \16447 );
buf \U$16415 ( \16449 , \16448 );
nand \U$16416 ( \16450 , \16264 , \16449 );
buf \U$16417 ( \16451 , \16450 );
buf \U$16418 ( \16452 , \16451 );
nand \U$16419 ( \16453 , \16261 , \16452 );
buf \U$16420 ( \16454 , \16453 );
buf \U$16421 ( \16455 , \16454 );
buf \U$16422 ( \16456 , \16101 );
not \U$16423 ( \16457 , \16456 );
buf \U$16424 ( \16458 , \16172 );
not \U$16425 ( \16459 , \16458 );
or \U$16426 ( \16460 , \16457 , \16459 );
buf \U$16427 ( \16461 , \16172 );
buf \U$16428 ( \16462 , \16101 );
or \U$16429 ( \16463 , \16461 , \16462 );
buf \U$16430 ( \16464 , \16034 );
nand \U$16431 ( \16465 , \16463 , \16464 );
buf \U$16432 ( \16466 , \16465 );
buf \U$16433 ( \16467 , \16466 );
nand \U$16434 ( \16468 , \16460 , \16467 );
buf \U$16435 ( \16469 , \16468 );
buf \U$16436 ( \16470 , \16469 );
not \U$16437 ( \16471 , \16470 );
buf \U$16438 ( \16472 , \13613 );
not \U$16439 ( \16473 , \16472 );
buf \U$16440 ( \16474 , \2037 );
not \U$16441 ( \16475 , \16474 );
or \U$16442 ( \16476 , \16473 , \16475 );
buf \U$16445 ( \16477 , \441 );
buf \U$16446 ( \16478 , \16477 );
buf \U$16447 ( \16479 , RIc0d8938_41);
buf \U$16448 ( \16480 , RIc0d9fb8_89);
xor \U$16449 ( \16481 , \16479 , \16480 );
buf \U$16450 ( \16482 , \16481 );
buf \U$16451 ( \16483 , \16482 );
nand \U$16452 ( \16484 , \16478 , \16483 );
buf \U$16453 ( \16485 , \16484 );
buf \U$16454 ( \16486 , \16485 );
nand \U$16455 ( \16487 , \16476 , \16486 );
buf \U$16456 ( \16488 , \16487 );
buf \U$16457 ( \16489 , \16488 );
buf \U$16458 ( \16490 , \14003 );
not \U$16459 ( \16491 , \16490 );
buf \U$16460 ( \16492 , \1124 );
not \U$16461 ( \16493 , \16492 );
buf \U$16462 ( \16494 , \16493 );
buf \U$16463 ( \16495 , \16494 );
not \U$16464 ( \16496 , \16495 );
or \U$16465 ( \16497 , \16491 , \16496 );
buf \U$16466 ( \16498 , \1562 );
not \U$16467 ( \16499 , \16498 );
buf \U$16468 ( \16500 , \16499 );
buf \U$16469 ( \16501 , \16500 );
buf \U$16470 ( \16502 , \14290 );
nand \U$16471 ( \16503 , \16501 , \16502 );
buf \U$16472 ( \16504 , \16503 );
buf \U$16473 ( \16505 , \16504 );
nand \U$16474 ( \16506 , \16497 , \16505 );
buf \U$16475 ( \16507 , \16506 );
buf \U$16476 ( \16508 , \16507 );
nor \U$16477 ( \16509 , \16489 , \16508 );
buf \U$16478 ( \16510 , \16509 );
buf \U$16479 ( \16511 , \16510 );
not \U$16480 ( \16512 , \14713 );
not \U$16481 ( \16513 , \13867 );
and \U$16482 ( \16514 , \16512 , \16513 );
buf \U$16483 ( \16515 , \14707 );
xor \U$16484 ( \16516 , RIc0da288_95, RIc0d8668_35);
buf \U$16485 ( \16517 , \16516 );
and \U$16486 ( \16518 , \16515 , \16517 );
buf \U$16487 ( \16519 , \16518 );
nor \U$16488 ( \16520 , \16514 , \16519 );
buf \U$16489 ( \16521 , \16520 );
or \U$16490 ( \16522 , \16511 , \16521 );
buf \U$16491 ( \16523 , \16488 );
buf \U$16492 ( \16524 , \16507 );
nand \U$16493 ( \16525 , \16523 , \16524 );
buf \U$16494 ( \16526 , \16525 );
buf \U$16495 ( \16527 , \16526 );
nand \U$16496 ( \16528 , \16522 , \16527 );
buf \U$16497 ( \16529 , \16528 );
buf \U$16498 ( \16530 , \16529 );
not \U$16499 ( \16531 , \16530 );
buf \U$16500 ( \16532 , \13955 );
not \U$16501 ( \16533 , \16532 );
buf \U$16502 ( \16534 , \14569 );
not \U$16503 ( \16535 , \16534 );
or \U$16504 ( \16536 , \16533 , \16535 );
buf \U$16505 ( \16537 , \13005 );
buf \U$16506 ( \16538 , \13157 );
nand \U$16507 ( \16539 , \16537 , \16538 );
buf \U$16508 ( \16540 , \16539 );
buf \U$16509 ( \16541 , \16540 );
nand \U$16510 ( \16542 , \16536 , \16541 );
buf \U$16511 ( \16543 , \16542 );
buf \U$16512 ( \16544 , \16543 );
not \U$16513 ( \16545 , \16544 );
buf \U$16514 ( \16546 , \16545 );
buf \U$16515 ( \16547 , \16546 );
not \U$16516 ( \16548 , \16547 );
buf \U$16517 ( \16549 , \13689 );
not \U$16518 ( \16550 , \16549 );
buf \U$16519 ( \16551 , \13684 );
not \U$16520 ( \16552 , \16551 );
or \U$16521 ( \16553 , \16550 , \16552 );
buf \U$16522 ( \16554 , \12936 );
not \U$16523 ( \16555 , \16554 );
buf \U$16524 ( \16556 , \16555 );
buf \U$16525 ( \16557 , \16556 );
not \U$16526 ( \16558 , \16557 );
buf \U$16527 ( \16559 , \16558 );
buf \U$16528 ( \16560 , \16559 );
buf \U$16529 ( \16561 , \13138 );
nand \U$16530 ( \16562 , \16560 , \16561 );
buf \U$16531 ( \16563 , \16562 );
buf \U$16532 ( \16564 , \16563 );
nand \U$16533 ( \16565 , \16553 , \16564 );
buf \U$16534 ( \16566 , \16565 );
buf \U$16535 ( \16567 , \16566 );
not \U$16536 ( \16568 , \16567 );
buf \U$16537 ( \16569 , \16568 );
buf \U$16538 ( \16570 , \16569 );
not \U$16539 ( \16571 , \16570 );
or \U$16540 ( \16572 , \16548 , \16571 );
buf \U$16541 ( \16573 , \13717 );
not \U$16542 ( \16574 , \16573 );
buf \U$16545 ( \16575 , \4482 );
buf \U$16546 ( \16576 , \16575 );
not \U$16547 ( \16577 , \16576 );
buf \U$16548 ( \16578 , \16577 );
buf \U$16549 ( \16579 , \16578 );
not \U$16550 ( \16580 , \16579 );
or \U$16551 ( \16581 , \16574 , \16580 );
buf \U$16552 ( \16582 , \4475 );
not \U$16553 ( \16583 , \16582 );
buf \U$16554 ( \16584 , \16583 );
buf \U$16555 ( \16585 , \16584 );
buf \U$16556 ( \16586 , RIc0da648_103);
buf \U$16557 ( \16587 , RIc0d82a8_27);
xor \U$16558 ( \16588 , \16586 , \16587 );
buf \U$16559 ( \16589 , \16588 );
buf \U$16560 ( \16590 , \16589 );
nand \U$16561 ( \16591 , \16585 , \16590 );
buf \U$16562 ( \16592 , \16591 );
buf \U$16563 ( \16593 , \16592 );
nand \U$16564 ( \16594 , \16581 , \16593 );
buf \U$16565 ( \16595 , \16594 );
buf \U$16566 ( \16596 , \16595 );
nand \U$16567 ( \16597 , \16572 , \16596 );
buf \U$16568 ( \16598 , \16597 );
buf \U$16569 ( \16599 , \16598 );
buf \U$16570 ( \16600 , \16566 );
buf \U$16571 ( \16601 , \16543 );
nand \U$16572 ( \16602 , \16600 , \16601 );
buf \U$16573 ( \16603 , \16602 );
buf \U$16574 ( \16604 , \16603 );
nand \U$16575 ( \16605 , \16599 , \16604 );
buf \U$16576 ( \16606 , \16605 );
buf \U$16577 ( \16607 , \16606 );
not \U$16578 ( \16608 , \16607 );
or \U$16579 ( \16609 , \16531 , \16608 );
buf \U$16580 ( \16610 , \16606 );
buf \U$16581 ( \16611 , \16529 );
or \U$16582 ( \16612 , \16610 , \16611 );
buf \U$16583 ( \16613 , \16436 );
not \U$16584 ( \16614 , \16613 );
buf \U$16585 ( \16615 , \16429 );
not \U$16586 ( \16616 , \16615 );
or \U$16587 ( \16617 , \16614 , \16616 );
buf \U$16588 ( \16618 , \16393 );
nand \U$16589 ( \16619 , \16617 , \16618 );
buf \U$16590 ( \16620 , \16619 );
buf \U$16591 ( \16621 , \16620 );
buf \U$16592 ( \16622 , \16426 );
buf \U$16593 ( \16623 , \16412 );
nand \U$16594 ( \16624 , \16622 , \16623 );
buf \U$16595 ( \16625 , \16624 );
buf \U$16596 ( \16626 , \16625 );
nand \U$16597 ( \16627 , \16621 , \16626 );
buf \U$16598 ( \16628 , \16627 );
buf \U$16599 ( \16629 , \16628 );
nand \U$16600 ( \16630 , \16612 , \16629 );
buf \U$16601 ( \16631 , \16630 );
buf \U$16602 ( \16632 , \16631 );
nand \U$16603 ( \16633 , \16609 , \16632 );
buf \U$16604 ( \16634 , \16633 );
buf \U$16605 ( \16635 , \16634 );
not \U$16606 ( \16636 , \16635 );
buf \U$16607 ( \16637 , \16636 );
buf \U$16608 ( \16638 , \16637 );
not \U$16609 ( \16639 , \16638 );
or \U$16610 ( \16640 , \16471 , \16639 );
buf \U$16611 ( \16641 , \16634 );
buf \U$16612 ( \16642 , \16469 );
not \U$16613 ( \16643 , \16642 );
buf \U$16614 ( \16644 , \16643 );
buf \U$16615 ( \16645 , \16644 );
nand \U$16616 ( \16646 , \16641 , \16645 );
buf \U$16617 ( \16647 , \16646 );
buf \U$16618 ( \16648 , \16647 );
nand \U$16619 ( \16649 , \16640 , \16648 );
buf \U$16620 ( \16650 , \16649 );
buf \U$16621 ( \16651 , \16650 );
buf \U$16622 ( \16652 , \13605 );
not \U$16623 ( \16653 , \16652 );
buf \U$16624 ( \16654 , \14888 );
not \U$16625 ( \16655 , \16654 );
buf \U$16626 ( \16656 , \16655 );
buf \U$16627 ( \16657 , \16656 );
not \U$16628 ( \16658 , \16657 );
or \U$16629 ( \16659 , \16653 , \16658 );
buf \U$16630 ( \16660 , \14402 );
not \U$16631 ( \16661 , \16660 );
buf \U$16632 ( \16662 , \16661 );
buf \U$16633 ( \16663 , \16662 );
buf \U$16634 ( \16664 , \14394 );
nand \U$16635 ( \16665 , \16663 , \16664 );
buf \U$16636 ( \16666 , \16665 );
buf \U$16637 ( \16667 , \16666 );
nand \U$16638 ( \16668 , \16659 , \16667 );
buf \U$16639 ( \16669 , \16668 );
buf \U$16640 ( \16670 , \16669 );
buf \U$16641 ( \16671 , \14048 );
not \U$16642 ( \16672 , \16671 );
buf \U$16643 ( \16673 , \4043 );
not \U$16644 ( \16674 , \16673 );
or \U$16645 ( \16675 , \16672 , \16674 );
buf \U$16648 ( \16676 , \15550 );
buf \U$16649 ( \16677 , \16676 );
buf \U$16650 ( \16678 , \14251 );
nand \U$16651 ( \16679 , \16677 , \16678 );
buf \U$16652 ( \16680 , \16679 );
buf \U$16653 ( \16681 , \16680 );
nand \U$16654 ( \16682 , \16675 , \16681 );
buf \U$16655 ( \16683 , \16682 );
buf \U$16656 ( \16684 , \16683 );
xor \U$16657 ( \16685 , \16670 , \16684 );
buf \U$16658 ( \16686 , \14982 );
not \U$16659 ( \16687 , \16686 );
buf \U$16660 ( \16688 , \16687 );
buf \U$16661 ( \16689 , \16688 );
buf \U$16662 ( \16690 , \16324 );
or \U$16663 ( \16691 , \16689 , \16690 );
buf \U$16666 ( \16692 , \12877 );
buf \U$16667 ( \16693 , \16692 );
not \U$16668 ( \16694 , \16693 );
buf \U$16669 ( \16695 , \16694 );
buf \U$16670 ( \16696 , \16695 );
buf \U$16671 ( \16697 , \14267 );
not \U$16672 ( \16698 , \16697 );
buf \U$16673 ( \16699 , \16698 );
buf \U$16674 ( \16700 , \16699 );
or \U$16675 ( \16701 , \16696 , \16700 );
nand \U$16676 ( \16702 , \16691 , \16701 );
buf \U$16677 ( \16703 , \16702 );
buf \U$16678 ( \16704 , \16703 );
and \U$16679 ( \16705 , \16685 , \16704 );
and \U$16680 ( \16706 , \16670 , \16684 );
or \U$16681 ( \16707 , \16705 , \16706 );
buf \U$16682 ( \16708 , \16707 );
not \U$16683 ( \16709 , \16708 );
and \U$16684 ( \16710 , \1078 , \14433 );
not \U$16685 ( \16711 , \13763 );
nor \U$16686 ( \16712 , \16711 , \1600 );
nor \U$16687 ( \16713 , \16710 , \16712 );
not \U$16688 ( \16714 , \16713 );
buf \U$16689 ( \16715 , \16714 );
not \U$16690 ( \16716 , \16715 );
buf \U$16691 ( \16717 , \13669 );
not \U$16692 ( \16718 , \16717 );
buf \U$16693 ( \16719 , \1431 );
not \U$16694 ( \16720 , \16719 );
or \U$16695 ( \16721 , \16718 , \16720 );
buf \U$16696 ( \16722 , \14374 );
buf \U$16697 ( \16723 , \14366 );
nand \U$16698 ( \16724 , \16722 , \16723 );
buf \U$16699 ( \16725 , \16724 );
buf \U$16700 ( \16726 , \16725 );
nand \U$16701 ( \16727 , \16721 , \16726 );
buf \U$16702 ( \16728 , \16727 );
buf \U$16703 ( \16729 , \16728 );
not \U$16704 ( \16730 , \16729 );
or \U$16705 ( \16731 , \16716 , \16730 );
buf \U$16706 ( \16732 , \16713 );
not \U$16707 ( \16733 , \16732 );
buf \U$16708 ( \16734 , \16728 );
not \U$16709 ( \16735 , \16734 );
buf \U$16710 ( \16736 , \16735 );
buf \U$16711 ( \16737 , \16736 );
not \U$16712 ( \16738 , \16737 );
or \U$16713 ( \16739 , \16733 , \16738 );
buf \U$16714 ( \16740 , \14145 );
not \U$16715 ( \16741 , \16740 );
buf \U$16716 ( \16742 , \2207 );
not \U$16717 ( \16743 , \16742 );
buf \U$16718 ( \16744 , \16743 );
buf \U$16719 ( \16745 , \16744 );
not \U$16720 ( \16746 , \16745 );
or \U$16721 ( \16747 , \16741 , \16746 );
buf \U$16722 ( \16748 , \2199 );
not \U$16723 ( \16749 , \16748 );
buf \U$16724 ( \16750 , \16749 );
buf \U$16725 ( \16751 , \16750 );
buf \U$16726 ( \16752 , \14414 );
nand \U$16727 ( \16753 , \16751 , \16752 );
buf \U$16728 ( \16754 , \16753 );
buf \U$16729 ( \16755 , \16754 );
nand \U$16730 ( \16756 , \16747 , \16755 );
buf \U$16731 ( \16757 , \16756 );
buf \U$16732 ( \16758 , \16757 );
nand \U$16733 ( \16759 , \16739 , \16758 );
buf \U$16734 ( \16760 , \16759 );
buf \U$16735 ( \16761 , \16760 );
nand \U$16736 ( \16762 , \16731 , \16761 );
buf \U$16737 ( \16763 , \16762 );
not \U$16738 ( \16764 , \16763 );
xor \U$16739 ( \16765 , \16206 , \16223 );
and \U$16740 ( \16766 , \16765 , \16251 );
and \U$16741 ( \16767 , \16206 , \16223 );
or \U$16742 ( \16768 , \16766 , \16767 );
buf \U$16743 ( \16769 , \16768 );
buf \U$16744 ( \16770 , \16769 );
not \U$16745 ( \16771 , \16770 );
buf \U$16746 ( \16772 , \16771 );
nand \U$16747 ( \16773 , \16764 , \16772 );
not \U$16748 ( \16774 , \16773 );
or \U$16749 ( \16775 , \16709 , \16774 );
buf \U$16750 ( \16776 , \16769 );
buf \U$16751 ( \16777 , \16763 );
nand \U$16752 ( \16778 , \16776 , \16777 );
buf \U$16753 ( \16779 , \16778 );
nand \U$16754 ( \16780 , \16775 , \16779 );
buf \U$16755 ( \16781 , \16780 );
xor \U$16756 ( \16782 , \16651 , \16781 );
buf \U$16757 ( \16783 , \16782 );
buf \U$16758 ( \16784 , \16783 );
xor \U$16759 ( \16785 , \16455 , \16784 );
buf \U$16760 ( \16786 , \16628 );
not \U$16761 ( \16787 , \16786 );
buf \U$16762 ( \16788 , \16787 );
xor \U$16763 ( \16789 , \16606 , \16788 );
xnor \U$16764 ( \16790 , \16789 , \16529 );
buf \U$16765 ( \16791 , \16790 );
buf \U$16766 ( \16792 , \16142 );
buf \U$16767 ( \16793 , \16121 );
and \U$16768 ( \16794 , \16792 , \16793 );
not \U$16769 ( \16795 , \16792 );
buf \U$16770 ( \16796 , \16118 );
and \U$16771 ( \16797 , \16795 , \16796 );
nor \U$16772 ( \16798 , \16794 , \16797 );
buf \U$16773 ( \16799 , \16798 );
xor \U$16774 ( \16800 , \16161 , \16799 );
buf \U$16775 ( \16801 , \16800 );
buf \U$16776 ( \16802 , \16520 );
not \U$16777 ( \16803 , \16802 );
buf \U$16778 ( \16804 , \16488 );
not \U$16779 ( \16805 , \16804 );
buf \U$16780 ( \16806 , \16507 );
not \U$16781 ( \16807 , \16806 );
buf \U$16782 ( \16808 , \16807 );
buf \U$16783 ( \16809 , \16808 );
not \U$16784 ( \16810 , \16809 );
or \U$16785 ( \16811 , \16805 , \16810 );
buf \U$16786 ( \16812 , \16488 );
buf \U$16787 ( \16813 , \16808 );
or \U$16788 ( \16814 , \16812 , \16813 );
nand \U$16789 ( \16815 , \16811 , \16814 );
buf \U$16790 ( \16816 , \16815 );
buf \U$16791 ( \16817 , \16816 );
not \U$16792 ( \16818 , \16817 );
or \U$16793 ( \16819 , \16803 , \16818 );
buf \U$16794 ( \16820 , \16816 );
buf \U$16795 ( \16821 , \16520 );
or \U$16796 ( \16822 , \16820 , \16821 );
nand \U$16797 ( \16823 , \16819 , \16822 );
buf \U$16798 ( \16824 , \16823 );
buf \U$16799 ( \16825 , \16824 );
xor \U$16800 ( \16826 , \16801 , \16825 );
xor \U$16801 ( \16827 , \16670 , \16684 );
xor \U$16802 ( \16828 , \16827 , \16704 );
buf \U$16803 ( \16829 , \16828 );
buf \U$16804 ( \16830 , \16829 );
and \U$16805 ( \16831 , \16826 , \16830 );
and \U$16806 ( \16832 , \16801 , \16825 );
or \U$16807 ( \16833 , \16831 , \16832 );
buf \U$16808 ( \16834 , \16833 );
buf \U$16809 ( \16835 , \16834 );
xor \U$16810 ( \16836 , \16791 , \16835 );
xor \U$16811 ( \16837 , \16763 , \16772 );
xnor \U$16812 ( \16838 , \16837 , \16708 );
buf \U$16813 ( \16839 , \16838 );
and \U$16814 ( \16840 , \16836 , \16839 );
and \U$16815 ( \16841 , \16791 , \16835 );
or \U$16816 ( \16842 , \16840 , \16841 );
buf \U$16817 ( \16843 , \16842 );
buf \U$16818 ( \16844 , \16843 );
and \U$16819 ( \16845 , \16785 , \16844 );
and \U$16820 ( \16846 , \16455 , \16784 );
or \U$16821 ( \16847 , \16845 , \16846 );
buf \U$16822 ( \16848 , \16847 );
buf \U$16823 ( \16849 , \16848 );
and \U$16824 ( \16850 , \15969 , \16849 );
not \U$16825 ( \16851 , \15969 );
buf \U$16826 ( \16852 , \16848 );
not \U$16827 ( \16853 , \16852 );
buf \U$16828 ( \16854 , \16853 );
buf \U$16829 ( \16855 , \16854 );
and \U$16830 ( \16856 , \16851 , \16855 );
nor \U$16831 ( \16857 , \16850 , \16856 );
buf \U$16832 ( \16858 , \16857 );
buf \U$16833 ( \16859 , \16858 );
not \U$16834 ( \16860 , \16859 );
buf \U$16835 ( \16861 , \16860 );
buf \U$16836 ( \16862 , \16861 );
and \U$16837 ( \16863 , \15312 , \16862 );
not \U$16838 ( \16864 , \15312 );
buf \U$16839 ( \16865 , \16858 );
and \U$16840 ( \16866 , \16864 , \16865 );
nor \U$16841 ( \16867 , \16863 , \16866 );
buf \U$16842 ( \16868 , \16867 );
buf \U$16843 ( \16869 , \16868 );
xor \U$16844 ( \16870 , RIc0da0a8_91, RIc0d8a28_43);
buf \U$16845 ( \16871 , \16870 );
not \U$16846 ( \16872 , \16871 );
buf \U$16847 ( \16873 , \16402 );
not \U$16848 ( \16874 , \16873 );
or \U$16849 ( \16875 , \16872 , \16874 );
buf \U$16850 ( \16876 , \530 );
not \U$16851 ( \16877 , \16876 );
buf \U$16852 ( \16878 , \14847 );
nand \U$16853 ( \16879 , \16877 , \16878 );
buf \U$16854 ( \16880 , \16879 );
buf \U$16855 ( \16881 , \16880 );
nand \U$16856 ( \16882 , \16875 , \16881 );
buf \U$16857 ( \16883 , \16882 );
buf \U$16858 ( \16884 , \16883 );
not \U$16859 ( \16885 , \16884 );
xor \U$16860 ( \16886 , RIc0da738_105, RIc0d8398_29);
buf \U$16861 ( \16887 , \16886 );
not \U$16862 ( \16888 , \16887 );
buf \U$16863 ( \16889 , \14804 );
not \U$16864 ( \16890 , \16889 );
or \U$16865 ( \16891 , \16888 , \16890 );
buf \U$16866 ( \16892 , \12744 );
buf \U$16867 ( \16893 , \14797 );
nand \U$16868 ( \16894 , \16892 , \16893 );
buf \U$16869 ( \16895 , \16894 );
buf \U$16870 ( \16896 , \16895 );
nand \U$16871 ( \16897 , \16891 , \16896 );
buf \U$16872 ( \16898 , \16897 );
buf \U$16873 ( \16899 , \16898 );
not \U$16874 ( \16900 , \16899 );
or \U$16875 ( \16901 , \16885 , \16900 );
buf \U$16876 ( \16902 , \16898 );
buf \U$16877 ( \16903 , \16883 );
or \U$16878 ( \16904 , \16902 , \16903 );
buf \U$16879 ( \16905 , RIc0d7a38_9);
buf \U$16880 ( \16906 , RIc0db098_125);
xor \U$16881 ( \16907 , \16905 , \16906 );
buf \U$16882 ( \16908 , \16907 );
buf \U$16883 ( \16909 , \16908 );
not \U$16884 ( \16910 , \16909 );
buf \U$16885 ( \16911 , \13452 );
buf \U$16886 ( \16912 , \13454 );
and \U$16887 ( \16913 , \16911 , \16912 );
buf \U$16888 ( \16914 , \16913 );
buf \U$16889 ( \16915 , \16914 );
not \U$16890 ( \16916 , \16915 );
or \U$16891 ( \16917 , \16910 , \16916 );
buf \U$16892 ( \16918 , \15793 );
buf \U$16893 ( \16919 , RIc0d79c0_8);
buf \U$16894 ( \16920 , RIc0db098_125);
xor \U$16895 ( \16921 , \16919 , \16920 );
buf \U$16896 ( \16922 , \16921 );
buf \U$16897 ( \16923 , \16922 );
nand \U$16898 ( \16924 , \16918 , \16923 );
buf \U$16899 ( \16925 , \16924 );
buf \U$16900 ( \16926 , \16925 );
nand \U$16901 ( \16927 , \16917 , \16926 );
buf \U$16902 ( \16928 , \16927 );
buf \U$16903 ( \16929 , \16928 );
nand \U$16904 ( \16930 , \16904 , \16929 );
buf \U$16905 ( \16931 , \16930 );
buf \U$16906 ( \16932 , \16931 );
nand \U$16907 ( \16933 , \16901 , \16932 );
buf \U$16908 ( \16934 , \16933 );
buf \U$16909 ( \16935 , \16934 );
buf \U$16910 ( \16936 , RIc0d8b18_45);
buf \U$16911 ( \16937 , RIc0d9fb8_89);
xor \U$16912 ( \16938 , \16936 , \16937 );
buf \U$16913 ( \16939 , \16938 );
buf \U$16914 ( \16940 , \16939 );
not \U$16915 ( \16941 , \16940 );
and \U$16916 ( \16942 , \427 , \429 );
buf \U$16917 ( \16943 , \16942 );
not \U$16918 ( \16944 , \16943 );
or \U$16919 ( \16945 , \16941 , \16944 );
buf \U$16920 ( \16946 , \13618 );
buf \U$16921 ( \16947 , \14959 );
nand \U$16922 ( \16948 , \16946 , \16947 );
buf \U$16923 ( \16949 , \16948 );
buf \U$16924 ( \16950 , \16949 );
nand \U$16925 ( \16951 , \16945 , \16950 );
buf \U$16926 ( \16952 , \16951 );
not \U$16927 ( \16953 , \16952 );
buf \U$16928 ( \16954 , RIc0d91a8_59);
not \U$16929 ( \16955 , \16954 );
buf \U$16930 ( \16956 , \16955 );
and \U$16931 ( \16957 , RIc0d9928_75, \16956 );
not \U$16932 ( \16958 , RIc0d9928_75);
and \U$16933 ( \16959 , \16958 , RIc0d91a8_59);
or \U$16934 ( \16960 , \16957 , \16959 );
buf \U$16935 ( \16961 , \16960 );
not \U$16936 ( \16962 , \16961 );
buf \U$16937 ( \16963 , \13991 );
not \U$16938 ( \16964 , \16963 );
or \U$16939 ( \16965 , \16962 , \16964 );
buf \U$16940 ( \16966 , \13998 );
buf \U$16941 ( \16967 , \14734 );
nand \U$16942 ( \16968 , \16966 , \16967 );
buf \U$16943 ( \16969 , \16968 );
buf \U$16944 ( \16970 , \16969 );
nand \U$16945 ( \16971 , \16965 , \16970 );
buf \U$16946 ( \16972 , \16971 );
not \U$16947 ( \16973 , \16972 );
or \U$16948 ( \16974 , \16953 , \16973 );
buf \U$16949 ( \16975 , \16972 );
not \U$16950 ( \16976 , \16975 );
buf \U$16951 ( \16977 , \16976 );
not \U$16952 ( \16978 , \16977 );
buf \U$16953 ( \16979 , \16952 );
not \U$16954 ( \16980 , \16979 );
buf \U$16955 ( \16981 , \16980 );
not \U$16956 ( \16982 , \16981 );
or \U$16957 ( \16983 , \16978 , \16982 );
xor \U$16958 ( \16984 , RIc0daaf8_113, RIc0d7fd8_21);
buf \U$16959 ( \16985 , \16984 );
not \U$16960 ( \16986 , \16985 );
buf \U$16961 ( \16987 , \14888 );
not \U$16962 ( \16988 , \16987 );
buf \U$16963 ( \16989 , \16988 );
buf \U$16964 ( \16990 , \16989 );
not \U$16965 ( \16991 , \16990 );
or \U$16966 ( \16992 , \16986 , \16991 );
buf \U$16967 ( \16993 , \14402 );
not \U$16968 ( \16994 , \16993 );
buf \U$16969 ( \16995 , \16994 );
buf \U$16970 ( \16996 , \16995 );
buf \U$16971 ( \16997 , \14881 );
nand \U$16972 ( \16998 , \16996 , \16997 );
buf \U$16973 ( \16999 , \16998 );
buf \U$16974 ( \17000 , \16999 );
nand \U$16975 ( \17001 , \16992 , \17000 );
buf \U$16976 ( \17002 , \17001 );
nand \U$16977 ( \17003 , \16983 , \17002 );
nand \U$16978 ( \17004 , \16974 , \17003 );
buf \U$16979 ( \17005 , \17004 );
xor \U$16980 ( \17006 , \16935 , \17005 );
buf \U$16981 ( \17007 , RIc0d9e50_86);
buf \U$16982 ( \17008 , RIc0d9ec8_87);
xor \U$16983 ( \17009 , \17007 , \17008 );
buf \U$16984 ( \17010 , \17009 );
not \U$16985 ( \17011 , \17010 );
not \U$16986 ( \17012 , \14544 );
or \U$16987 ( \17013 , \17011 , \17012 );
buf \U$16988 ( \17014 , RIc0d8cf8_49);
buf \U$16989 ( \17015 , RIc0d9dd8_85);
xnor \U$16990 ( \17016 , \17014 , \17015 );
buf \U$16991 ( \17017 , \17016 );
or \U$16992 ( \17018 , \2396 , \17017 );
nand \U$16993 ( \17019 , \17013 , \17018 );
buf \U$16994 ( \17020 , \17019 );
xor \U$16995 ( \17021 , RIc0da468_99, RIc0d8668_35);
buf \U$16996 ( \17022 , \17021 );
not \U$16997 ( \17023 , \17022 );
buf \U$16998 ( \17024 , \14419 );
not \U$16999 ( \17025 , \17024 );
or \U$17000 ( \17026 , \17023 , \17025 );
buf \U$17001 ( \17027 , \12584 );
buf \U$17002 ( \17028 , \14640 );
nand \U$17003 ( \17029 , \17027 , \17028 );
buf \U$17004 ( \17030 , \17029 );
buf \U$17005 ( \17031 , \17030 );
nand \U$17006 ( \17032 , \17026 , \17031 );
buf \U$17007 ( \17033 , \17032 );
buf \U$17008 ( \17034 , \17033 );
xor \U$17009 ( \17035 , \17020 , \17034 );
buf \U$17010 ( \17036 , RIc0d7ee8_19);
buf \U$17011 ( \17037 , RIc0dabe8_115);
xor \U$17012 ( \17038 , \17036 , \17037 );
buf \U$17013 ( \17039 , \17038 );
buf \U$17014 ( \17040 , \17039 );
not \U$17015 ( \17041 , \17040 );
buf \U$17016 ( \17042 , \14186 );
not \U$17017 ( \17043 , \17042 );
or \U$17018 ( \17044 , \17041 , \17043 );
buf \U$17019 ( \17045 , \12303 );
buf \U$17020 ( \17046 , \14678 );
nand \U$17021 ( \17047 , \17045 , \17046 );
buf \U$17022 ( \17048 , \17047 );
buf \U$17023 ( \17049 , \17048 );
nand \U$17024 ( \17050 , \17044 , \17049 );
buf \U$17025 ( \17051 , \17050 );
buf \U$17026 ( \17052 , \17051 );
and \U$17027 ( \17053 , \17035 , \17052 );
and \U$17028 ( \17054 , \17020 , \17034 );
or \U$17029 ( \17055 , \17053 , \17054 );
buf \U$17030 ( \17056 , \17055 );
buf \U$17031 ( \17057 , \17056 );
and \U$17032 ( \17058 , \17006 , \17057 );
and \U$17033 ( \17059 , \16935 , \17005 );
or \U$17034 ( \17060 , \17058 , \17059 );
buf \U$17035 ( \17061 , \17060 );
not \U$17036 ( \17062 , \17061 );
buf \U$17037 ( \17063 , RIc0d8c08_47);
buf \U$17038 ( \17064 , RIc0d9ec8_87);
xor \U$17039 ( \17065 , \17063 , \17064 );
buf \U$17040 ( \17066 , \17065 );
buf \U$17041 ( \17067 , \17066 );
not \U$17042 ( \17068 , \17067 );
buf \U$17043 ( \17069 , \4527 );
not \U$17044 ( \17070 , \17069 );
or \U$17045 ( \17071 , \17068 , \17070 );
buf \U$17046 ( \17072 , \14331 );
buf \U$17047 ( \17073 , \14621 );
nand \U$17048 ( \17074 , \17072 , \17073 );
buf \U$17049 ( \17075 , \17074 );
buf \U$17050 ( \17076 , \17075 );
nand \U$17051 ( \17077 , \17071 , \17076 );
buf \U$17052 ( \17078 , \17077 );
buf \U$17053 ( \17079 , \17078 );
not \U$17054 ( \17080 , \17079 );
buf \U$17055 ( \17081 , RIc0d7c18_13);
buf \U$17056 ( \17082 , RIc0daeb8_121);
xor \U$17057 ( \17083 , \17081 , \17082 );
buf \U$17058 ( \17084 , \17083 );
buf \U$17059 ( \17085 , \17084 );
not \U$17060 ( \17086 , \17085 );
buf \U$17061 ( \17087 , \12968 );
not \U$17062 ( \17088 , \17087 );
buf \U$17063 ( \17089 , \17088 );
buf \U$17064 ( \17090 , \17089 );
not \U$17065 ( \17091 , \17090 );
or \U$17066 ( \17092 , \17086 , \17091 );
buf \U$17067 ( \17093 , \13314 );
buf \U$17068 ( \17094 , RIc0d7ba0_12);
buf \U$17069 ( \17095 , RIc0daeb8_121);
xor \U$17070 ( \17096 , \17094 , \17095 );
buf \U$17071 ( \17097 , \17096 );
buf \U$17072 ( \17098 , \17097 );
nand \U$17073 ( \17099 , \17093 , \17098 );
buf \U$17074 ( \17100 , \17099 );
buf \U$17075 ( \17101 , \17100 );
nand \U$17076 ( \17102 , \17092 , \17101 );
buf \U$17077 ( \17103 , \17102 );
buf \U$17078 ( \17104 , \17103 );
not \U$17079 ( \17105 , \17104 );
or \U$17080 ( \17106 , \17080 , \17105 );
buf \U$17081 ( \17107 , \17103 );
buf \U$17082 ( \17108 , \17078 );
or \U$17083 ( \17109 , \17107 , \17108 );
buf \U$17084 ( \17110 , RIc0d7b28_11);
buf \U$17085 ( \17111 , RIc0dafa8_123);
xor \U$17086 ( \17112 , \17110 , \17111 );
buf \U$17087 ( \17113 , \17112 );
buf \U$17088 ( \17114 , \17113 );
not \U$17089 ( \17115 , \17114 );
buf \U$17090 ( \17116 , \14982 );
not \U$17091 ( \17117 , \17116 );
or \U$17092 ( \17118 , \17115 , \17117 );
buf \U$17093 ( \17119 , \16692 );
buf \U$17094 ( \17120 , \14974 );
nand \U$17095 ( \17121 , \17119 , \17120 );
buf \U$17096 ( \17122 , \17121 );
buf \U$17097 ( \17123 , \17122 );
nand \U$17098 ( \17124 , \17118 , \17123 );
buf \U$17099 ( \17125 , \17124 );
buf \U$17100 ( \17126 , \17125 );
nand \U$17101 ( \17127 , \17109 , \17126 );
buf \U$17102 ( \17128 , \17127 );
buf \U$17103 ( \17129 , \17128 );
nand \U$17104 ( \17130 , \17106 , \17129 );
buf \U$17105 ( \17131 , \17130 );
buf \U$17106 ( \17132 , \17131 );
buf \U$17107 ( \17133 , RIc0d8ed8_53);
buf \U$17108 ( \17134 , RIc0d9bf8_81);
xor \U$17109 ( \17135 , \17133 , \17134 );
buf \U$17110 ( \17136 , \17135 );
buf \U$17111 ( \17137 , \17136 );
not \U$17112 ( \17138 , \17137 );
buf \U$17113 ( \17139 , \1060 );
not \U$17114 ( \17140 , \17139 );
buf \U$17115 ( \17141 , \17140 );
buf \U$17116 ( \17142 , \17141 );
not \U$17117 ( \17143 , \17142 );
or \U$17118 ( \17144 , \17138 , \17143 );
buf \U$17119 ( \17145 , \1078 );
buf \U$17120 ( \17146 , \14527 );
nand \U$17121 ( \17147 , \17145 , \17146 );
buf \U$17122 ( \17148 , \17147 );
buf \U$17123 ( \17149 , \17148 );
nand \U$17124 ( \17150 , \17144 , \17149 );
buf \U$17125 ( \17151 , \17150 );
buf \U$17126 ( \17152 , \17151 );
not \U$17127 ( \17153 , \17152 );
buf \U$17128 ( \17154 , RIc0d7d08_15);
buf \U$17129 ( \17155 , RIc0dadc8_119);
xor \U$17130 ( \17156 , \17154 , \17155 );
buf \U$17131 ( \17157 , \17156 );
buf \U$17132 ( \17158 , \17157 );
not \U$17133 ( \17159 , \17158 );
buf \U$17134 ( \17160 , \13001 );
not \U$17135 ( \17161 , \17160 );
or \U$17136 ( \17162 , \17159 , \17161 );
buf \U$17137 ( \17163 , \13005 );
buf \U$17138 ( \17164 , \14564 );
nand \U$17139 ( \17165 , \17163 , \17164 );
buf \U$17140 ( \17166 , \17165 );
buf \U$17141 ( \17167 , \17166 );
nand \U$17142 ( \17168 , \17162 , \17167 );
buf \U$17143 ( \17169 , \17168 );
buf \U$17144 ( \17170 , \17169 );
not \U$17145 ( \17171 , \17170 );
or \U$17146 ( \17172 , \17153 , \17171 );
buf \U$17147 ( \17173 , \17151 );
buf \U$17148 ( \17174 , \17169 );
or \U$17149 ( \17175 , \17173 , \17174 );
buf \U$17150 ( \17176 , RIc0d8de8_51);
buf \U$17151 ( \17177 , RIc0d9ce8_83);
xor \U$17152 ( \17178 , \17176 , \17177 );
buf \U$17153 ( \17179 , \17178 );
buf \U$17154 ( \17180 , \17179 );
not \U$17155 ( \17181 , \17180 );
buf \U$17156 ( \17182 , \2088 );
not \U$17157 ( \17183 , \17182 );
or \U$17158 ( \17184 , \17181 , \17183 );
buf \U$17159 ( \17185 , \993 );
buf \U$17160 ( \17186 , \14911 );
nand \U$17161 ( \17187 , \17185 , \17186 );
buf \U$17162 ( \17188 , \17187 );
buf \U$17163 ( \17189 , \17188 );
nand \U$17164 ( \17190 , \17184 , \17189 );
buf \U$17165 ( \17191 , \17190 );
buf \U$17166 ( \17192 , \17191 );
nand \U$17167 ( \17193 , \17175 , \17192 );
buf \U$17168 ( \17194 , \17193 );
buf \U$17169 ( \17195 , \17194 );
nand \U$17170 ( \17196 , \17172 , \17195 );
buf \U$17171 ( \17197 , \17196 );
buf \U$17172 ( \17198 , \17197 );
or \U$17173 ( \17199 , \17132 , \17198 );
buf \U$17174 ( \17200 , RIc0d7948_7);
buf \U$17175 ( \17201 , RIc0db188_127);
xor \U$17176 ( \17202 , \17200 , \17201 );
buf \U$17177 ( \17203 , \17202 );
buf \U$17178 ( \17204 , \17203 );
not \U$17179 ( \17205 , \17204 );
buf \U$17180 ( \17206 , \12654 );
not \U$17181 ( \17207 , \17206 );
or \U$17182 ( \17208 , \17205 , \17207 );
buf \U$17183 ( \17209 , RIc0d78d0_6);
buf \U$17184 ( \17210 , RIc0db188_127);
xor \U$17185 ( \17211 , \17209 , \17210 );
buf \U$17186 ( \17212 , \17211 );
buf \U$17187 ( \17213 , \17212 );
buf \U$17188 ( \17214 , RIc0db200_128);
nand \U$17189 ( \17215 , \17213 , \17214 );
buf \U$17190 ( \17216 , \17215 );
buf \U$17191 ( \17217 , \17216 );
nand \U$17192 ( \17218 , \17208 , \17217 );
buf \U$17193 ( \17219 , \17218 );
buf \U$17194 ( \17220 , \17219 );
buf \U$17195 ( \17221 , RIc0d80c8_23);
buf \U$17196 ( \17222 , RIc0daa08_111);
xor \U$17197 ( \17223 , \17221 , \17222 );
buf \U$17198 ( \17224 , \17223 );
buf \U$17199 ( \17225 , \17224 );
not \U$17200 ( \17226 , \17225 );
buf \U$17201 ( \17227 , \14100 );
not \U$17202 ( \17228 , \17227 );
or \U$17203 ( \17229 , \17226 , \17228 );
buf \U$17204 ( \17230 , \14353 );
buf \U$17205 ( \17231 , \14866 );
nand \U$17206 ( \17232 , \17230 , \17231 );
buf \U$17207 ( \17233 , \17232 );
buf \U$17208 ( \17234 , \17233 );
nand \U$17209 ( \17235 , \17229 , \17234 );
buf \U$17210 ( \17236 , \17235 );
buf \U$17211 ( \17237 , \17236 );
xor \U$17212 ( \17238 , \17220 , \17237 );
buf \U$17213 ( \17239 , RIc0d8578_33);
buf \U$17214 ( \17240 , RIc0da558_101);
xor \U$17215 ( \17241 , \17239 , \17240 );
buf \U$17216 ( \17242 , \17241 );
buf \U$17217 ( \17243 , \17242 );
not \U$17218 ( \17244 , \17243 );
buf \U$17219 ( \17245 , \4042 );
not \U$17220 ( \17246 , \17245 );
or \U$17221 ( \17247 , \17244 , \17246 );
buf \U$17222 ( \17248 , \4049 );
buf \U$17223 ( \17249 , \14772 );
nand \U$17224 ( \17250 , \17248 , \17249 );
buf \U$17225 ( \17251 , \17250 );
buf \U$17226 ( \17252 , \17251 );
nand \U$17227 ( \17253 , \17247 , \17252 );
buf \U$17228 ( \17254 , \17253 );
buf \U$17229 ( \17255 , \17254 );
and \U$17230 ( \17256 , \17238 , \17255 );
and \U$17231 ( \17257 , \17220 , \17237 );
or \U$17232 ( \17258 , \17256 , \17257 );
buf \U$17233 ( \17259 , \17258 );
buf \U$17234 ( \17260 , \17259 );
nand \U$17235 ( \17261 , \17199 , \17260 );
buf \U$17236 ( \17262 , \17261 );
buf \U$17237 ( \17263 , \17262 );
buf \U$17238 ( \17264 , \17131 );
buf \U$17239 ( \17265 , \17197 );
nand \U$17240 ( \17266 , \17264 , \17265 );
buf \U$17241 ( \17267 , \17266 );
buf \U$17242 ( \17268 , \17267 );
nand \U$17243 ( \17269 , \17263 , \17268 );
buf \U$17244 ( \17270 , \17269 );
not \U$17245 ( \17271 , \17270 );
or \U$17246 ( \17272 , \17062 , \17271 );
buf \U$17247 ( \17273 , \17061 );
not \U$17248 ( \17274 , \17273 );
buf \U$17249 ( \17275 , \17274 );
not \U$17250 ( \17276 , \17275 );
buf \U$17251 ( \17277 , \17270 );
not \U$17252 ( \17278 , \17277 );
buf \U$17253 ( \17279 , \17278 );
not \U$17254 ( \17280 , \17279 );
or \U$17255 ( \17281 , \17276 , \17280 );
xor \U$17256 ( \17282 , \14862 , \14930 );
xor \U$17257 ( \17283 , \17282 , \15008 );
buf \U$17258 ( \17284 , \17283 );
nand \U$17259 ( \17285 , \17281 , \17284 );
nand \U$17260 ( \17286 , \17272 , \17285 );
buf \U$17261 ( \17287 , \17286 );
xor \U$17262 ( \17288 , \14597 , \14795 );
xor \U$17263 ( \17289 , \17288 , \15013 );
buf \U$17264 ( \17290 , \17289 );
buf \U$17265 ( \17291 , \17290 );
xor \U$17266 ( \17292 , \17287 , \17291 );
buf \U$17267 ( \17293 , \14788 );
buf \U$17268 ( \17294 , \14661 );
xor \U$17269 ( \17295 , \17293 , \17294 );
buf \U$17270 ( \17296 , \14724 );
xnor \U$17271 ( \17297 , \17295 , \17296 );
buf \U$17272 ( \17298 , \17297 );
buf \U$17273 ( \17299 , \17298 );
not \U$17274 ( \17300 , \17299 );
buf \U$17275 ( \17301 , \17300 );
buf \U$17276 ( \17302 , \17301 );
not \U$17277 ( \17303 , \17302 );
xor \U$17278 ( \17304 , RIc0da198_93, RIc0d88c0_40);
buf \U$17279 ( \17305 , \17304 );
not \U$17280 ( \17306 , \17305 );
buf \U$17281 ( \17307 , \15995 );
not \U$17282 ( \17308 , \17307 );
or \U$17283 ( \17309 , \17306 , \17308 );
buf \U$17284 ( \17310 , \481 );
buf \U$17285 ( \17311 , \16297 );
nand \U$17286 ( \17312 , \17310 , \17311 );
buf \U$17287 ( \17313 , \17312 );
buf \U$17288 ( \17314 , \17313 );
nand \U$17289 ( \17315 , \17309 , \17314 );
buf \U$17290 ( \17316 , \17315 );
buf \U$17291 ( \17317 , \17316 );
buf \U$17292 ( \17318 , RIc0d8230_26);
buf \U$17293 ( \17319 , RIc0da828_107);
xor \U$17294 ( \17320 , \17318 , \17319 );
buf \U$17295 ( \17321 , \17320 );
buf \U$17296 ( \17322 , \17321 );
not \U$17297 ( \17323 , \17322 );
buf \U$17298 ( \17324 , \16065 );
not \U$17299 ( \17325 , \17324 );
or \U$17300 ( \17326 , \17323 , \17325 );
buf \U$17301 ( \17327 , \12342 );
buf \U$17302 ( \17328 , \16282 );
nand \U$17303 ( \17329 , \17327 , \17328 );
buf \U$17304 ( \17330 , \17329 );
buf \U$17305 ( \17331 , \17330 );
nand \U$17306 ( \17332 , \17326 , \17331 );
buf \U$17307 ( \17333 , \17332 );
buf \U$17308 ( \17334 , \17333 );
or \U$17309 ( \17335 , \17317 , \17334 );
buf \U$17310 ( \17336 , \17097 );
not \U$17311 ( \17337 , \17336 );
buf \U$17312 ( \17338 , \15420 );
not \U$17313 ( \17339 , \17338 );
or \U$17314 ( \17340 , \17337 , \17339 );
buf \U$17315 ( \17341 , \16386 );
buf \U$17316 ( \17342 , \13775 );
nand \U$17317 ( \17343 , \17341 , \17342 );
buf \U$17318 ( \17344 , \17343 );
buf \U$17319 ( \17345 , \17344 );
nand \U$17320 ( \17346 , \17340 , \17345 );
buf \U$17321 ( \17347 , \17346 );
buf \U$17322 ( \17348 , \17347 );
nand \U$17323 ( \17349 , \17335 , \17348 );
buf \U$17324 ( \17350 , \17349 );
buf \U$17325 ( \17351 , \17350 );
buf \U$17326 ( \17352 , \17316 );
buf \U$17327 ( \17353 , \17333 );
nand \U$17328 ( \17354 , \17352 , \17353 );
buf \U$17329 ( \17355 , \17354 );
buf \U$17330 ( \17356 , \17355 );
nand \U$17331 ( \17357 , \17351 , \17356 );
buf \U$17332 ( \17358 , \17357 );
buf \U$17333 ( \17359 , \17358 );
buf \U$17334 ( \17360 , RIc0d86e0_36);
buf \U$17335 ( \17361 , RIc0da378_97);
xor \U$17336 ( \17362 , \17360 , \17361 );
buf \U$17337 ( \17363 , \17362 );
buf \U$17338 ( \17364 , \17363 );
not \U$17339 ( \17365 , \17364 );
buf \U$17340 ( \17366 , \15329 );
not \U$17341 ( \17367 , \17366 );
or \U$17342 ( \17368 , \17365 , \17367 );
buf \U$17343 ( \17369 , \734 );
buf \U$17344 ( \17370 , \16353 );
nand \U$17345 ( \17371 , \17369 , \17370 );
buf \U$17346 ( \17372 , \17371 );
buf \U$17347 ( \17373 , \17372 );
nand \U$17348 ( \17374 , \17368 , \17373 );
buf \U$17349 ( \17375 , \17374 );
buf \U$17350 ( \17376 , \17375 );
not \U$17351 ( \17377 , \17376 );
xor \U$17352 ( \17378 , RIc0dacd8_117, RIc0d7d80_16);
buf \U$17353 ( \17379 , \17378 );
not \U$17354 ( \17380 , \17379 );
buf \U$17355 ( \17381 , \13684 );
not \U$17356 ( \17382 , \17381 );
or \U$17357 ( \17383 , \17380 , \17382 );
buf \U$17358 ( \17384 , \12937 );
buf \U$17359 ( \17385 , \13677 );
nand \U$17360 ( \17386 , \17384 , \17385 );
buf \U$17361 ( \17387 , \17386 );
buf \U$17362 ( \17388 , \17387 );
nand \U$17363 ( \17389 , \17383 , \17388 );
buf \U$17364 ( \17390 , \17389 );
buf \U$17365 ( \17391 , \17390 );
not \U$17366 ( \17392 , \17391 );
or \U$17367 ( \17393 , \17377 , \17392 );
buf \U$17368 ( \17394 , \17390 );
buf \U$17369 ( \17395 , \17375 );
or \U$17370 ( \17396 , \17394 , \17395 );
buf \U$17371 ( \17397 , RIc0d8410_30);
buf \U$17372 ( \17398 , RIc0da648_103);
xor \U$17373 ( \17399 , \17397 , \17398 );
buf \U$17374 ( \17400 , \17399 );
buf \U$17375 ( \17401 , \17400 );
not \U$17376 ( \17402 , \17401 );
buf \U$17377 ( \17403 , \16575 );
not \U$17378 ( \17404 , \17403 );
buf \U$17379 ( \17405 , \17404 );
buf \U$17380 ( \17406 , \17405 );
not \U$17381 ( \17407 , \17406 );
or \U$17382 ( \17408 , \17402 , \17407 );
buf \U$17383 ( \17409 , \13048 );
buf \U$17384 ( \17410 , \13701 );
nand \U$17385 ( \17411 , \17409 , \17410 );
buf \U$17386 ( \17412 , \17411 );
buf \U$17387 ( \17413 , \17412 );
nand \U$17388 ( \17414 , \17408 , \17413 );
buf \U$17389 ( \17415 , \17414 );
buf \U$17390 ( \17416 , \17415 );
nand \U$17391 ( \17417 , \17396 , \17416 );
buf \U$17392 ( \17418 , \17417 );
buf \U$17393 ( \17419 , \17418 );
nand \U$17394 ( \17420 , \17393 , \17419 );
buf \U$17395 ( \17421 , \17420 );
buf \U$17396 ( \17422 , \17421 );
xor \U$17397 ( \17423 , \17359 , \17422 );
xor \U$17398 ( \17424 , \14172 , \14198 );
xor \U$17399 ( \17425 , \17424 , \14228 );
buf \U$17400 ( \17426 , \17425 );
buf \U$17401 ( \17427 , \17426 );
xor \U$17402 ( \17428 , \17423 , \17427 );
buf \U$17403 ( \17429 , \17428 );
buf \U$17404 ( \17430 , \17429 );
not \U$17405 ( \17431 , \17430 );
or \U$17406 ( \17432 , \17303 , \17431 );
buf \U$17407 ( \17433 , \17429 );
not \U$17408 ( \17434 , \17433 );
buf \U$17409 ( \17435 , \17298 );
nand \U$17410 ( \17436 , \17434 , \17435 );
buf \U$17411 ( \17437 , \17436 );
buf \U$17412 ( \17438 , \17437 );
buf \U$17413 ( \17439 , \14954 );
buf \U$17414 ( \17440 , \14971 );
xor \U$17415 ( \17441 , \17439 , \17440 );
buf \U$17416 ( \17442 , \14996 );
xnor \U$17417 ( \17443 , \17441 , \17442 );
buf \U$17418 ( \17444 , \17443 );
buf \U$17419 ( \17445 , \17444 );
not \U$17420 ( \17446 , \17445 );
buf \U$17421 ( \17447 , \17446 );
buf \U$17422 ( \17448 , \17447 );
not \U$17423 ( \17449 , \17448 );
buf \U$17424 ( \17450 , \14844 );
buf \U$17425 ( \17451 , \14835 );
and \U$17426 ( \17452 , \17450 , \17451 );
not \U$17427 ( \17453 , \17450 );
buf \U$17428 ( \17454 , \14840 );
and \U$17429 ( \17455 , \17453 , \17454 );
or \U$17430 ( \17456 , \17452 , \17455 );
buf \U$17431 ( \17457 , \17456 );
buf \U$17432 ( \17458 , \17457 );
not \U$17433 ( \17459 , \17458 );
buf \U$17434 ( \17460 , \14859 );
not \U$17435 ( \17461 , \17460 );
buf \U$17436 ( \17462 , \17461 );
buf \U$17437 ( \17463 , \17462 );
not \U$17438 ( \17464 , \17463 );
and \U$17439 ( \17465 , \17459 , \17464 );
buf \U$17440 ( \17466 , \17457 );
buf \U$17441 ( \17467 , \17462 );
and \U$17442 ( \17468 , \17466 , \17467 );
nor \U$17443 ( \17469 , \17465 , \17468 );
buf \U$17444 ( \17470 , \17469 );
buf \U$17445 ( \17471 , \17470 );
not \U$17446 ( \17472 , \17471 );
buf \U$17447 ( \17473 , \17472 );
buf \U$17448 ( \17474 , \17473 );
not \U$17449 ( \17475 , \17474 );
or \U$17450 ( \17476 , \17449 , \17475 );
buf \U$17451 ( \17477 , \17444 );
not \U$17452 ( \17478 , \17477 );
buf \U$17453 ( \17479 , \17470 );
not \U$17454 ( \17480 , \17479 );
or \U$17455 ( \17481 , \17478 , \17480 );
buf \U$17456 ( \17482 , \17390 );
not \U$17457 ( \17483 , \17482 );
buf \U$17458 ( \17484 , \17375 );
not \U$17459 ( \17485 , \17484 );
buf \U$17460 ( \17486 , \17485 );
buf \U$17461 ( \17487 , \17486 );
not \U$17462 ( \17488 , \17487 );
or \U$17463 ( \17489 , \17483 , \17488 );
buf \U$17464 ( \17490 , \17486 );
buf \U$17465 ( \17491 , \17390 );
or \U$17466 ( \17492 , \17490 , \17491 );
nand \U$17467 ( \17493 , \17489 , \17492 );
buf \U$17468 ( \17494 , \17493 );
buf \U$17469 ( \17495 , \17494 );
buf \U$17470 ( \17496 , \17415 );
xor \U$17471 ( \17497 , \17495 , \17496 );
buf \U$17472 ( \17498 , \17497 );
buf \U$17473 ( \17499 , \17498 );
nand \U$17474 ( \17500 , \17481 , \17499 );
buf \U$17475 ( \17501 , \17500 );
buf \U$17476 ( \17502 , \17501 );
nand \U$17477 ( \17503 , \17476 , \17502 );
buf \U$17478 ( \17504 , \17503 );
buf \U$17479 ( \17505 , \17504 );
nand \U$17480 ( \17506 , \17438 , \17505 );
buf \U$17481 ( \17507 , \17506 );
buf \U$17482 ( \17508 , \17507 );
nand \U$17483 ( \17509 , \17432 , \17508 );
buf \U$17484 ( \17510 , \17509 );
buf \U$17485 ( \17511 , \17510 );
and \U$17486 ( \17512 , \17292 , \17511 );
and \U$17487 ( \17513 , \17287 , \17291 );
or \U$17488 ( \17514 , \17512 , \17513 );
buf \U$17489 ( \17515 , \17514 );
buf \U$17490 ( \17516 , \17515 );
buf \U$17491 ( \17517 , \14764 );
buf \U$17492 ( \17518 , \14746 );
xor \U$17493 ( \17519 , \17517 , \17518 );
buf \U$17494 ( \17520 , \14784 );
not \U$17495 ( \17521 , \17520 );
xor \U$17496 ( \17522 , \17519 , \17521 );
buf \U$17497 ( \17523 , \17522 );
buf \U$17498 ( \17524 , \17523 );
not \U$17499 ( \17525 , \17524 );
buf \U$17500 ( \17526 , \17525 );
not \U$17501 ( \17527 , \17526 );
buf \U$17502 ( \17528 , \14618 );
buf \U$17503 ( \17529 , \14633 );
xor \U$17504 ( \17530 , \17528 , \17529 );
buf \U$17505 ( \17531 , \14655 );
xnor \U$17506 ( \17532 , \17530 , \17531 );
buf \U$17507 ( \17533 , \17532 );
buf \U$17508 ( \17534 , \17533 );
not \U$17509 ( \17535 , \17534 );
buf \U$17510 ( \17536 , \17535 );
not \U$17511 ( \17537 , \17536 );
or \U$17512 ( \17538 , \17527 , \17537 );
not \U$17513 ( \17539 , \17533 );
not \U$17514 ( \17540 , \17523 );
or \U$17515 ( \17541 , \17539 , \17540 );
buf \U$17516 ( \17542 , \17347 );
buf \U$17517 ( \17543 , \17333 );
xor \U$17518 ( \17544 , \17542 , \17543 );
buf \U$17519 ( \17545 , \17544 );
buf \U$17520 ( \17546 , \17545 );
buf \U$17521 ( \17547 , \17316 );
xor \U$17522 ( \17548 , \17546 , \17547 );
buf \U$17523 ( \17549 , \17548 );
nand \U$17524 ( \17550 , \17541 , \17549 );
nand \U$17525 ( \17551 , \17538 , \17550 );
buf \U$17526 ( \17552 , \17551 );
xor \U$17527 ( \17553 , \13612 , \13635 );
xor \U$17528 ( \17554 , \17553 , \13651 );
buf \U$17529 ( \17555 , \17554 );
buf \U$17530 ( \17556 , \17555 );
xor \U$17531 ( \17557 , \13676 , \13696 );
xor \U$17532 ( \17558 , \17557 , \13724 );
buf \U$17533 ( \17559 , \17558 );
buf \U$17534 ( \17560 , \17559 );
xor \U$17535 ( \17561 , \17556 , \17560 );
buf \U$17536 ( \17562 , \16332 );
buf \U$17537 ( \17563 , \16345 );
xor \U$17538 ( \17564 , \17562 , \17563 );
buf \U$17539 ( \17565 , \16368 );
xor \U$17540 ( \17566 , \17564 , \17565 );
buf \U$17541 ( \17567 , \17566 );
buf \U$17542 ( \17568 , \17567 );
xor \U$17543 ( \17569 , \17561 , \17568 );
buf \U$17544 ( \17570 , \17569 );
buf \U$17545 ( \17571 , \17570 );
xor \U$17546 ( \17572 , \17552 , \17571 );
xor \U$17547 ( \17573 , RIc0d9b08_79, RIc0d8fc8_55);
buf \U$17548 ( \17574 , \17573 );
not \U$17549 ( \17575 , \17574 );
buf \U$17550 ( \17576 , \1351 );
not \U$17551 ( \17577 , \17576 );
or \U$17552 ( \17578 , \17575 , \17577 );
buf \U$17553 ( \17579 , \1026 );
buf \U$17554 ( \17580 , \14935 );
nand \U$17555 ( \17581 , \17579 , \17580 );
buf \U$17556 ( \17582 , \17581 );
buf \U$17557 ( \17583 , \17582 );
nand \U$17558 ( \17584 , \17578 , \17583 );
buf \U$17559 ( \17585 , \17584 );
buf \U$17560 ( \17586 , \17585 );
buf \U$17561 ( \17587 , RIc0da828_107);
buf \U$17562 ( \17588 , RIc0d82a8_27);
xor \U$17563 ( \17589 , \17587 , \17588 );
buf \U$17564 ( \17590 , \17589 );
buf \U$17565 ( \17591 , \17590 );
not \U$17566 ( \17592 , \17591 );
buf \U$17567 ( \17593 , \12331 );
not \U$17568 ( \17594 , \17593 );
buf \U$17569 ( \17595 , \17594 );
buf \U$17570 ( \17596 , \17595 );
not \U$17571 ( \17597 , \17596 );
or \U$17572 ( \17598 , \17592 , \17597 );
buf \U$17573 ( \17599 , \12342 );
buf \U$17574 ( \17600 , \17321 );
nand \U$17575 ( \17601 , \17599 , \17600 );
buf \U$17576 ( \17602 , \17601 );
buf \U$17577 ( \17603 , \17602 );
nand \U$17578 ( \17604 , \17598 , \17603 );
buf \U$17579 ( \17605 , \17604 );
buf \U$17580 ( \17606 , \17605 );
nor \U$17581 ( \17607 , \17586 , \17606 );
buf \U$17582 ( \17608 , \17607 );
buf \U$17583 ( \17609 , \17608 );
buf \U$17584 ( \17610 , RIc0d8938_41);
buf \U$17585 ( \17611 , RIc0da198_93);
xor \U$17586 ( \17612 , \17610 , \17611 );
buf \U$17587 ( \17613 , \17612 );
buf \U$17588 ( \17614 , \17613 );
not \U$17589 ( \17615 , \17614 );
buf \U$17590 ( \17616 , \3415 );
not \U$17591 ( \17617 , \17616 );
or \U$17592 ( \17618 , \17615 , \17617 );
buf \U$17593 ( \17619 , \481 );
buf \U$17594 ( \17620 , \17304 );
nand \U$17595 ( \17621 , \17619 , \17620 );
buf \U$17596 ( \17622 , \17621 );
buf \U$17597 ( \17623 , \17622 );
nand \U$17598 ( \17624 , \17618 , \17623 );
buf \U$17599 ( \17625 , \17624 );
buf \U$17600 ( \17626 , \17625 );
not \U$17601 ( \17627 , \17626 );
buf \U$17602 ( \17628 , \17627 );
buf \U$17603 ( \17629 , \17628 );
or \U$17604 ( \17630 , \17609 , \17629 );
buf \U$17605 ( \17631 , \17585 );
buf \U$17606 ( \17632 , \17605 );
nand \U$17607 ( \17633 , \17631 , \17632 );
buf \U$17608 ( \17634 , \17633 );
buf \U$17609 ( \17635 , \17634 );
nand \U$17610 ( \17636 , \17630 , \17635 );
buf \U$17611 ( \17637 , \17636 );
buf \U$17612 ( \17638 , \17637 );
xor \U$17613 ( \17639 , \14677 , \14698 );
xor \U$17614 ( \17640 , \17639 , \14720 );
buf \U$17615 ( \17641 , \17640 );
buf \U$17616 ( \17642 , \17641 );
xor \U$17617 ( \17643 , \17638 , \17642 );
xor \U$17618 ( \17644 , \14923 , \14878 );
xor \U$17619 ( \17645 , \17644 , \14901 );
buf \U$17620 ( \17646 , \17645 );
and \U$17621 ( \17647 , \17643 , \17646 );
and \U$17622 ( \17648 , \17638 , \17642 );
or \U$17623 ( \17649 , \17647 , \17648 );
buf \U$17624 ( \17650 , \17649 );
buf \U$17625 ( \17651 , \17650 );
and \U$17626 ( \17652 , \17572 , \17651 );
and \U$17627 ( \17653 , \17552 , \17571 );
or \U$17628 ( \17654 , \17652 , \17653 );
buf \U$17629 ( \17655 , \17654 );
buf \U$17630 ( \17656 , \17655 );
not \U$17631 ( \17657 , \17656 );
xor \U$17632 ( \17658 , \13656 , \13729 );
xor \U$17633 ( \17659 , \17658 , \13797 );
buf \U$17634 ( \17660 , \17659 );
buf \U$17635 ( \17661 , \17660 );
xor \U$17636 ( \17662 , \16315 , \16376 );
xor \U$17637 ( \17663 , \17662 , \16444 );
buf \U$17638 ( \17664 , \17663 );
buf \U$17639 ( \17665 , \17664 );
xor \U$17640 ( \17666 , \17661 , \17665 );
xor \U$17641 ( \17667 , \14066 , \14154 );
xor \U$17642 ( \17668 , \17667 , \14233 );
buf \U$17643 ( \17669 , \17668 );
buf \U$17644 ( \17670 , \17669 );
xor \U$17645 ( \17671 , \17666 , \17670 );
buf \U$17646 ( \17672 , \17671 );
buf \U$17647 ( \17673 , \17672 );
not \U$17648 ( \17674 , \17673 );
or \U$17649 ( \17675 , \17657 , \17674 );
buf \U$17650 ( \17676 , \17655 );
buf \U$17651 ( \17677 , \17672 );
or \U$17652 ( \17678 , \17676 , \17677 );
xor \U$17653 ( \17679 , \13812 , \13885 );
xor \U$17654 ( \17680 , \17679 , \13973 );
buf \U$17655 ( \17681 , \13912 );
not \U$17656 ( \17682 , \17681 );
buf \U$17657 ( \17683 , \13937 );
not \U$17658 ( \17684 , \17683 );
or \U$17659 ( \17685 , \17682 , \17684 );
buf \U$17660 ( \17686 , \13934 );
buf \U$17661 ( \17687 , \13915 );
nand \U$17662 ( \17688 , \17686 , \17687 );
buf \U$17663 ( \17689 , \17688 );
buf \U$17664 ( \17690 , \17689 );
nand \U$17665 ( \17691 , \17685 , \17690 );
buf \U$17666 ( \17692 , \17691 );
buf \U$17667 ( \17693 , \17692 );
buf \U$17668 ( \17694 , \13961 );
not \U$17669 ( \17695 , \17694 );
buf \U$17670 ( \17696 , \17695 );
buf \U$17671 ( \17697 , \17696 );
and \U$17672 ( \17698 , \17693 , \17697 );
not \U$17673 ( \17699 , \17693 );
buf \U$17674 ( \17700 , \13961 );
and \U$17675 ( \17701 , \17699 , \17700 );
nor \U$17676 ( \17702 , \17698 , \17701 );
buf \U$17677 ( \17703 , \17702 );
buf \U$17678 ( \17704 , \17703 );
not \U$17679 ( \17705 , \17704 );
buf \U$17680 ( \17706 , \17705 );
buf \U$17681 ( \17707 , \17706 );
not \U$17682 ( \17708 , \17707 );
buf \U$17683 ( \17709 , \14151 );
not \U$17684 ( \17710 , \17709 );
buf \U$17685 ( \17711 , \14122 );
not \U$17686 ( \17712 , \17711 );
or \U$17687 ( \17713 , \17710 , \17712 );
buf \U$17688 ( \17714 , \14151 );
buf \U$17689 ( \17715 , \14122 );
or \U$17690 ( \17716 , \17714 , \17715 );
nand \U$17691 ( \17717 , \17713 , \17716 );
buf \U$17692 ( \17718 , \17717 );
buf \U$17693 ( \17719 , \17718 );
buf \U$17694 ( \17720 , \14126 );
and \U$17695 ( \17721 , \17719 , \17720 );
not \U$17696 ( \17722 , \17719 );
buf \U$17697 ( \17723 , \14089 );
and \U$17698 ( \17724 , \17722 , \17723 );
nor \U$17699 ( \17725 , \17721 , \17724 );
buf \U$17700 ( \17726 , \17725 );
buf \U$17701 ( \17727 , \17726 );
not \U$17702 ( \17728 , \17727 );
buf \U$17703 ( \17729 , \17728 );
buf \U$17704 ( \17730 , \17729 );
not \U$17705 ( \17731 , \17730 );
or \U$17706 ( \17732 , \17708 , \17731 );
buf \U$17707 ( \17733 , \17726 );
not \U$17708 ( \17734 , \17733 );
buf \U$17709 ( \17735 , \17703 );
not \U$17710 ( \17736 , \17735 );
or \U$17711 ( \17737 , \17734 , \17736 );
xor \U$17712 ( \17738 , \13752 , \13770 );
xor \U$17713 ( \17739 , \17738 , \13792 );
buf \U$17714 ( \17740 , \17739 );
buf \U$17715 ( \17741 , \17740 );
nand \U$17716 ( \17742 , \17737 , \17741 );
buf \U$17717 ( \17743 , \17742 );
buf \U$17718 ( \17744 , \17743 );
nand \U$17719 ( \17745 , \17732 , \17744 );
buf \U$17720 ( \17746 , \17745 );
xor \U$17721 ( \17747 , \17680 , \17746 );
buf \U$17722 ( \17748 , \14054 );
not \U$17723 ( \17749 , \17748 );
buf \U$17724 ( \17750 , \14012 );
not \U$17725 ( \17751 , \17750 );
or \U$17726 ( \17752 , \17749 , \17751 );
buf \U$17727 ( \17753 , \14054 );
buf \U$17728 ( \17754 , \14012 );
or \U$17729 ( \17755 , \17753 , \17754 );
nand \U$17730 ( \17756 , \17752 , \17755 );
buf \U$17731 ( \17757 , \17756 );
buf \U$17732 ( \17758 , \17757 );
not \U$17733 ( \17759 , \17758 );
buf \U$17734 ( \17760 , \14028 );
not \U$17735 ( \17761 , \17760 );
buf \U$17736 ( \17762 , \17761 );
buf \U$17737 ( \17763 , \17762 );
not \U$17738 ( \17764 , \17763 );
and \U$17739 ( \17765 , \17759 , \17764 );
buf \U$17740 ( \17766 , \17757 );
buf \U$17741 ( \17767 , \17762 );
and \U$17742 ( \17768 , \17766 , \17767 );
nor \U$17743 ( \17769 , \17765 , \17768 );
buf \U$17744 ( \17770 , \17769 );
buf \U$17745 ( \17771 , \17770 );
not \U$17746 ( \17772 , \17771 );
buf \U$17747 ( \17773 , \17772 );
not \U$17748 ( \17774 , \17773 );
buf \U$17749 ( \17775 , \13821 );
buf \U$17750 ( \17776 , \13843 );
xor \U$17751 ( \17777 , \17775 , \17776 );
buf \U$17752 ( \17778 , \13879 );
xnor \U$17753 ( \17779 , \17777 , \17778 );
buf \U$17754 ( \17780 , \17779 );
buf \U$17755 ( \17781 , \17780 );
not \U$17756 ( \17782 , \17781 );
buf \U$17757 ( \17783 , \17782 );
not \U$17758 ( \17784 , \17783 );
or \U$17759 ( \17785 , \17774 , \17784 );
not \U$17760 ( \17786 , \17780 );
not \U$17761 ( \17787 , \17770 );
or \U$17762 ( \17788 , \17786 , \17787 );
xor \U$17763 ( \17789 , \16278 , \16295 );
xor \U$17764 ( \17790 , \17789 , \16310 );
buf \U$17765 ( \17791 , \17790 );
nand \U$17766 ( \17792 , \17788 , \17791 );
nand \U$17767 ( \17793 , \17785 , \17792 );
xnor \U$17768 ( \17794 , \17747 , \17793 );
buf \U$17769 ( \17795 , \17794 );
nand \U$17770 ( \17796 , \17678 , \17795 );
buf \U$17771 ( \17797 , \17796 );
buf \U$17772 ( \17798 , \17797 );
nand \U$17773 ( \17799 , \17675 , \17798 );
buf \U$17774 ( \17800 , \17799 );
buf \U$17775 ( \17801 , \17800 );
xor \U$17776 ( \17802 , \17516 , \17801 );
buf \U$17777 ( \17803 , \17793 );
not \U$17778 ( \17804 , \17803 );
buf \U$17779 ( \17805 , \17746 );
not \U$17780 ( \17806 , \17805 );
or \U$17781 ( \17807 , \17804 , \17806 );
buf \U$17782 ( \17808 , \17746 );
buf \U$17783 ( \17809 , \17793 );
or \U$17784 ( \17810 , \17808 , \17809 );
buf \U$17785 ( \17811 , \17680 );
not \U$17786 ( \17812 , \17811 );
buf \U$17787 ( \17813 , \17812 );
buf \U$17788 ( \17814 , \17813 );
nand \U$17789 ( \17815 , \17810 , \17814 );
buf \U$17790 ( \17816 , \17815 );
buf \U$17791 ( \17817 , \17816 );
nand \U$17792 ( \17818 , \17807 , \17817 );
buf \U$17793 ( \17819 , \17818 );
buf \U$17794 ( \17820 , \17819 );
xor \U$17795 ( \17821 , \13802 , \13980 );
xor \U$17796 ( \17822 , \17821 , \14238 );
buf \U$17797 ( \17823 , \17822 );
buf \U$17798 ( \17824 , \17823 );
xor \U$17799 ( \17825 , \17820 , \17824 );
xor \U$17800 ( \17826 , \17661 , \17665 );
and \U$17801 ( \17827 , \17826 , \17670 );
and \U$17802 ( \17828 , \17661 , \17665 );
or \U$17803 ( \17829 , \17827 , \17828 );
buf \U$17804 ( \17830 , \17829 );
buf \U$17805 ( \17831 , \17830 );
xor \U$17806 ( \17832 , \17825 , \17831 );
buf \U$17807 ( \17833 , \17832 );
buf \U$17808 ( \17834 , \17833 );
and \U$17809 ( \17835 , \17802 , \17834 );
and \U$17810 ( \17836 , \17516 , \17801 );
or \U$17811 ( \17837 , \17835 , \17836 );
buf \U$17812 ( \17838 , \17837 );
buf \U$17813 ( \17839 , \17838 );
xor \U$17814 ( \17840 , \17820 , \17824 );
and \U$17815 ( \17841 , \17840 , \17831 );
and \U$17816 ( \17842 , \17820 , \17824 );
or \U$17817 ( \17843 , \17841 , \17842 );
buf \U$17818 ( \17844 , \17843 );
buf \U$17819 ( \17845 , \17844 );
xor \U$17820 ( \17846 , \16182 , \16188 );
xor \U$17821 ( \17847 , \17846 , \16254 );
buf \U$17822 ( \17848 , \17847 );
buf \U$17823 ( \17849 , \17848 );
not \U$17824 ( \17850 , \17849 );
xor \U$17825 ( \17851 , \17359 , \17422 );
and \U$17826 ( \17852 , \17851 , \17427 );
and \U$17827 ( \17853 , \17359 , \17422 );
or \U$17828 ( \17854 , \17852 , \17853 );
buf \U$17829 ( \17855 , \17854 );
buf \U$17830 ( \17856 , \17855 );
not \U$17831 ( \17857 , \17856 );
or \U$17832 ( \17858 , \17850 , \17857 );
buf \U$17833 ( \17859 , \17855 );
buf \U$17834 ( \17860 , \17848 );
or \U$17835 ( \17861 , \17859 , \17860 );
xor \U$17836 ( \17862 , \17556 , \17560 );
and \U$17837 ( \17863 , \17862 , \17568 );
and \U$17838 ( \17864 , \17556 , \17560 );
or \U$17839 ( \17865 , \17863 , \17864 );
buf \U$17840 ( \17866 , \17865 );
buf \U$17841 ( \17867 , \17866 );
nand \U$17842 ( \17868 , \17861 , \17867 );
buf \U$17843 ( \17869 , \17868 );
buf \U$17844 ( \17870 , \17869 );
nand \U$17845 ( \17871 , \17858 , \17870 );
buf \U$17846 ( \17872 , \17871 );
buf \U$17847 ( \17873 , \17872 );
not \U$17848 ( \17874 , \17873 );
buf \U$17849 ( \17875 , \16173 );
buf \U$17850 ( \17876 , \16448 );
or \U$17851 ( \17877 , \17875 , \17876 );
buf \U$17852 ( \17878 , \16173 );
buf \U$17853 ( \17879 , \16448 );
nand \U$17854 ( \17880 , \17878 , \17879 );
buf \U$17855 ( \17881 , \17880 );
buf \U$17856 ( \17882 , \17881 );
nand \U$17857 ( \17883 , \17877 , \17882 );
buf \U$17858 ( \17884 , \17883 );
buf \U$17859 ( \17885 , \17884 );
buf \U$17860 ( \17886 , \16258 );
not \U$17861 ( \17887 , \17886 );
buf \U$17862 ( \17888 , \17887 );
buf \U$17863 ( \17889 , \17888 );
and \U$17864 ( \17890 , \17885 , \17889 );
not \U$17865 ( \17891 , \17885 );
buf \U$17866 ( \17892 , \16258 );
and \U$17867 ( \17893 , \17891 , \17892 );
nor \U$17868 ( \17894 , \17890 , \17893 );
buf \U$17869 ( \17895 , \17894 );
buf \U$17870 ( \17896 , \17895 );
not \U$17871 ( \17897 , \17896 );
buf \U$17872 ( \17898 , \17897 );
buf \U$17873 ( \17899 , \17898 );
not \U$17874 ( \17900 , \17899 );
or \U$17875 ( \17901 , \17874 , \17900 );
buf \U$17876 ( \17902 , \17898 );
buf \U$17877 ( \17903 , \17872 );
or \U$17878 ( \17904 , \17902 , \17903 );
xor \U$17879 ( \17905 , \16791 , \16835 );
xor \U$17880 ( \17906 , \17905 , \16839 );
buf \U$17881 ( \17907 , \17906 );
buf \U$17882 ( \17908 , \17907 );
nand \U$17883 ( \17909 , \17904 , \17908 );
buf \U$17884 ( \17910 , \17909 );
buf \U$17885 ( \17911 , \17910 );
nand \U$17886 ( \17912 , \17901 , \17911 );
buf \U$17887 ( \17913 , \17912 );
buf \U$17888 ( \17914 , \17913 );
xor \U$17889 ( \17915 , \17845 , \17914 );
xor \U$17890 ( \17916 , \16455 , \16784 );
xor \U$17891 ( \17917 , \17916 , \16844 );
buf \U$17892 ( \17918 , \17917 );
buf \U$17893 ( \17919 , \17918 );
xor \U$17894 ( \17920 , \17915 , \17919 );
buf \U$17895 ( \17921 , \17920 );
buf \U$17896 ( \17922 , \17921 );
xor \U$17897 ( \17923 , \17839 , \17922 );
buf \U$17898 ( \17924 , \17895 );
not \U$17899 ( \17925 , \17924 );
buf \U$17900 ( \17926 , \17872 );
not \U$17901 ( \17927 , \17926 );
and \U$17902 ( \17928 , \17925 , \17927 );
buf \U$17903 ( \17929 , \17872 );
buf \U$17904 ( \17930 , \17895 );
and \U$17905 ( \17931 , \17929 , \17930 );
nor \U$17906 ( \17932 , \17928 , \17931 );
buf \U$17907 ( \17933 , \17932 );
buf \U$17908 ( \17934 , \17933 );
buf \U$17909 ( \17935 , \17907 );
not \U$17910 ( \17936 , \17935 );
buf \U$17911 ( \17937 , \17936 );
buf \U$17912 ( \17938 , \17937 );
and \U$17913 ( \17939 , \17934 , \17938 );
not \U$17914 ( \17940 , \17934 );
buf \U$17915 ( \17941 , \17907 );
and \U$17916 ( \17942 , \17940 , \17941 );
nor \U$17917 ( \17943 , \17939 , \17942 );
buf \U$17918 ( \17944 , \17943 );
buf \U$17919 ( \17945 , \17944 );
buf \U$17920 ( \17946 , \17791 );
buf \U$17921 ( \17947 , \17783 );
and \U$17922 ( \17948 , \17946 , \17947 );
not \U$17923 ( \17949 , \17946 );
buf \U$17924 ( \17950 , \17780 );
and \U$17925 ( \17951 , \17949 , \17950 );
nor \U$17926 ( \17952 , \17948 , \17951 );
buf \U$17927 ( \17953 , \17952 );
buf \U$17928 ( \17954 , \17953 );
buf \U$17929 ( \17955 , \17773 );
and \U$17930 ( \17956 , \17954 , \17955 );
not \U$17931 ( \17957 , \17954 );
buf \U$17932 ( \17958 , \17770 );
and \U$17933 ( \17959 , \17957 , \17958 );
nor \U$17934 ( \17960 , \17956 , \17959 );
buf \U$17935 ( \17961 , \17960 );
buf \U$17936 ( \17962 , \17961 );
buf \U$17937 ( \17963 , \17706 );
not \U$17938 ( \17964 , \17963 );
buf \U$17939 ( \17965 , \17740 );
buf \U$17940 ( \17966 , \17726 );
and \U$17941 ( \17967 , \17965 , \17966 );
not \U$17942 ( \17968 , \17965 );
buf \U$17943 ( \17969 , \17729 );
and \U$17944 ( \17970 , \17968 , \17969 );
nor \U$17945 ( \17971 , \17967 , \17970 );
buf \U$17946 ( \17972 , \17971 );
buf \U$17947 ( \17973 , \17972 );
not \U$17948 ( \17974 , \17973 );
or \U$17949 ( \17975 , \17964 , \17974 );
buf \U$17950 ( \17976 , \17972 );
not \U$17951 ( \17977 , \17976 );
buf \U$17952 ( \17978 , \17703 );
nand \U$17953 ( \17979 , \17977 , \17978 );
buf \U$17954 ( \17980 , \17979 );
buf \U$17955 ( \17981 , \17980 );
nand \U$17956 ( \17982 , \17975 , \17981 );
buf \U$17957 ( \17983 , \17982 );
buf \U$17958 ( \17984 , \17983 );
xor \U$17959 ( \17985 , \17962 , \17984 );
xor \U$17960 ( \17986 , \14502 , \14519 );
buf \U$17961 ( \17987 , \17986 );
buf \U$17962 ( \17988 , \17987 );
not \U$17963 ( \17989 , \17988 );
buf \U$17964 ( \17990 , \16922 );
not \U$17965 ( \17991 , \17990 );
buf \U$17968 ( \17992 , \13457 );
buf \U$17969 ( \17993 , \17992 );
not \U$17970 ( \17994 , \17993 );
buf \U$17971 ( \17995 , \17994 );
buf \U$17972 ( \17996 , \17995 );
not \U$17973 ( \17997 , \17996 );
or \U$17974 ( \17998 , \17991 , \17997 );
buf \U$17975 ( \17999 , \15793 );
buf \U$17976 ( \18000 , \14463 );
nand \U$17977 ( \18001 , \17999 , \18000 );
buf \U$17978 ( \18002 , \18001 );
buf \U$17979 ( \18003 , \18002 );
nand \U$17980 ( \18004 , \17998 , \18003 );
buf \U$17981 ( \18005 , \18004 );
buf \U$17982 ( \18006 , \18005 );
not \U$17983 ( \18007 , \18006 );
not \U$17984 ( \18008 , \15609 );
buf \U$17985 ( \18009 , \18008 );
not \U$17986 ( \18010 , \18009 );
buf \U$17987 ( \18011 , \17212 );
not \U$17988 ( \18012 , \18011 );
buf \U$17989 ( \18013 , \18012 );
buf \U$17990 ( \18014 , \18013 );
not \U$17991 ( \18015 , \18014 );
and \U$17992 ( \18016 , \18010 , \18015 );
buf \U$17993 ( \18017 , \16265 );
buf \U$17994 ( \18018 , RIc0db200_128);
and \U$17995 ( \18019 , \18017 , \18018 );
nor \U$17996 ( \18020 , \18016 , \18019 );
buf \U$17997 ( \18021 , \18020 );
buf \U$17998 ( \18022 , \18021 );
not \U$17999 ( \18023 , \18022 );
and \U$18000 ( \18024 , \18007 , \18023 );
buf \U$18001 ( \18025 , \18005 );
buf \U$18002 ( \18026 , \18021 );
and \U$18003 ( \18027 , \18025 , \18026 );
nor \U$18004 ( \18028 , \18024 , \18027 );
buf \U$18005 ( \18029 , \18028 );
buf \U$18006 ( \18030 , \18029 );
not \U$18007 ( \18031 , \18030 );
or \U$18008 ( \18032 , \17989 , \18031 );
buf \U$18009 ( \18033 , \17987 );
buf \U$18010 ( \18034 , \18029 );
or \U$18011 ( \18035 , \18033 , \18034 );
nand \U$18012 ( \18036 , \18032 , \18035 );
buf \U$18013 ( \18037 , \18036 );
buf \U$18014 ( \18038 , \18037 );
and \U$18015 ( \18039 , \14542 , \14582 );
not \U$18016 ( \18040 , \14542 );
and \U$18017 ( \18041 , \18040 , \14579 );
or \U$18018 ( \18042 , \18039 , \18041 );
buf \U$18019 ( \18043 , \18042 );
buf \U$18020 ( \18044 , \14556 );
xor \U$18021 ( \18045 , \18043 , \18044 );
buf \U$18022 ( \18046 , \18045 );
buf \U$18023 ( \18047 , \18046 );
xor \U$18024 ( \18048 , \18038 , \18047 );
buf \U$18025 ( \18049 , RIc0d9310_62);
buf \U$18026 ( \18050 , RIc0d9838_73);
xor \U$18027 ( \18051 , \18049 , \18050 );
buf \U$18028 ( \18052 , \18051 );
buf \U$18029 ( \18053 , \18052 );
not \U$18030 ( \18054 , \18053 );
buf \U$18031 ( \18055 , \773 );
not \U$18032 ( \18056 , \18055 );
buf \U$18033 ( \18057 , \18056 );
buf \U$18034 ( \18058 , \18057 );
not \U$18035 ( \18059 , \18058 );
or \U$18036 ( \18060 , \18054 , \18059 );
buf \U$18037 ( \18061 , \791 );
buf \U$18038 ( \18062 , RIc0d9298_61);
buf \U$18039 ( \18063 , RIc0d9838_73);
xor \U$18040 ( \18064 , \18062 , \18063 );
buf \U$18041 ( \18065 , \18064 );
buf \U$18042 ( \18066 , \18065 );
nand \U$18043 ( \18067 , \18061 , \18066 );
buf \U$18044 ( \18068 , \18067 );
buf \U$18045 ( \18069 , \18068 );
nand \U$18046 ( \18070 , \18060 , \18069 );
buf \U$18047 ( \18071 , \18070 );
buf \U$18048 ( \18072 , \18071 );
buf \U$18049 ( \18073 , RIc0d9400_64);
buf \U$18050 ( \18074 , RIc0d97c0_72);
or \U$18051 ( \18075 , \18073 , \18074 );
buf \U$18052 ( \18076 , RIc0d9838_73);
nand \U$18053 ( \18077 , \18075 , \18076 );
buf \U$18054 ( \18078 , \18077 );
buf \U$18055 ( \18079 , \18078 );
buf \U$18056 ( \18080 , RIc0d9400_64);
buf \U$18057 ( \18081 , RIc0d97c0_72);
nand \U$18058 ( \18082 , \18080 , \18081 );
buf \U$18059 ( \18083 , \18082 );
buf \U$18060 ( \18084 , \18083 );
buf \U$18061 ( \18085 , RIc0d9748_71);
and \U$18062 ( \18086 , \18079 , \18084 , \18085 );
buf \U$18063 ( \18087 , \18086 );
buf \U$18064 ( \18088 , \18087 );
and \U$18065 ( \18089 , \18072 , \18088 );
buf \U$18066 ( \18090 , \18089 );
buf \U$18067 ( \18091 , \18090 );
buf \U$18068 ( \18092 , RIc0d9130_58);
buf \U$18069 ( \18093 , RIc0d9a18_77);
xor \U$18070 ( \18094 , \18092 , \18093 );
buf \U$18071 ( \18095 , \18094 );
buf \U$18072 ( \18096 , \18095 );
not \U$18073 ( \18097 , \18096 );
buf \U$18074 ( \18098 , \14825 );
not \U$18075 ( \18099 , \18098 );
or \U$18076 ( \18100 , \18097 , \18099 );
buf \U$18077 ( \18101 , \1588 );
buf \U$18078 ( \18102 , RIc0d90b8_57);
buf \U$18079 ( \18103 , RIc0d9a18_77);
xor \U$18080 ( \18104 , \18102 , \18103 );
buf \U$18081 ( \18105 , \18104 );
buf \U$18082 ( \18106 , \18105 );
nand \U$18083 ( \18107 , \18101 , \18106 );
buf \U$18084 ( \18108 , \18107 );
buf \U$18085 ( \18109 , \18108 );
nand \U$18086 ( \18110 , \18100 , \18109 );
buf \U$18087 ( \18111 , \18110 );
buf \U$18088 ( \18112 , \18111 );
not \U$18089 ( \18113 , \18112 );
buf \U$18090 ( \18114 , RIc0d9220_60);
buf \U$18091 ( \18115 , RIc0d9928_75);
xor \U$18092 ( \18116 , \18114 , \18115 );
buf \U$18093 ( \18117 , \18116 );
not \U$18094 ( \18118 , \18117 );
buf \U$18095 ( \18119 , \2358 );
not \U$18096 ( \18120 , \18119 );
buf \U$18097 ( \18121 , \18120 );
nor \U$18098 ( \18122 , \18118 , \18121 );
buf \U$18099 ( \18123 , \18122 );
buf \U$18100 ( \18124 , \13998 );
buf \U$18101 ( \18125 , \16960 );
and \U$18102 ( \18126 , \18124 , \18125 );
buf \U$18103 ( \18127 , \18126 );
buf \U$18104 ( \18128 , \18127 );
nor \U$18105 ( \18129 , \18123 , \18128 );
buf \U$18106 ( \18130 , \18129 );
buf \U$18107 ( \18131 , \18130 );
not \U$18108 ( \18132 , \18131 );
buf \U$18109 ( \18133 , \18132 );
buf \U$18110 ( \18134 , \18133 );
not \U$18111 ( \18135 , \18134 );
or \U$18112 ( \18136 , \18113 , \18135 );
buf \U$18113 ( \18137 , \18111 );
not \U$18114 ( \18138 , \18137 );
buf \U$18115 ( \18139 , \18138 );
buf \U$18116 ( \18140 , \18139 );
not \U$18117 ( \18141 , \18140 );
buf \U$18118 ( \18142 , \18130 );
not \U$18119 ( \18143 , \18142 );
or \U$18120 ( \18144 , \18141 , \18143 );
xor \U$18121 ( \18145 , RIc0d9fb8_89, RIc0d8b90_46);
buf \U$18122 ( \18146 , \18145 );
not \U$18123 ( \18147 , \18146 );
buf \U$18124 ( \18148 , \2034 );
not \U$18125 ( \18149 , \18148 );
buf \U$18126 ( \18150 , \18149 );
buf \U$18127 ( \18151 , \18150 );
not \U$18128 ( \18152 , \18151 );
or \U$18129 ( \18153 , \18147 , \18152 );
buf \U$18130 ( \18154 , \846 );
buf \U$18131 ( \18155 , \16939 );
nand \U$18132 ( \18156 , \18154 , \18155 );
buf \U$18133 ( \18157 , \18156 );
buf \U$18134 ( \18158 , \18157 );
nand \U$18135 ( \18159 , \18153 , \18158 );
buf \U$18136 ( \18160 , \18159 );
buf \U$18137 ( \18161 , \18160 );
nand \U$18138 ( \18162 , \18144 , \18161 );
buf \U$18139 ( \18163 , \18162 );
buf \U$18140 ( \18164 , \18163 );
nand \U$18141 ( \18165 , \18136 , \18164 );
buf \U$18142 ( \18166 , \18165 );
buf \U$18143 ( \18167 , \18166 );
xor \U$18144 ( \18168 , \18091 , \18167 );
buf \U$18145 ( \18169 , RIc0d9400_64);
buf \U$18146 ( \18170 , RIc0d9748_71);
xor \U$18147 ( \18171 , \18169 , \18170 );
buf \U$18148 ( \18172 , \18171 );
buf \U$18149 ( \18173 , \18172 );
not \U$18150 ( \18174 , \18173 );
buf \U$18151 ( \18175 , \1888 );
not \U$18152 ( \18176 , \18175 );
or \U$18153 ( \18177 , \18174 , \18176 );
buf \U$18154 ( \18178 , \2927 );
buf \U$18155 ( \18179 , RIc0d9388_63);
buf \U$18156 ( \18180 , RIc0d9748_71);
xor \U$18157 ( \18181 , \18179 , \18180 );
buf \U$18158 ( \18182 , \18181 );
buf \U$18159 ( \18183 , \18182 );
nand \U$18160 ( \18184 , \18178 , \18183 );
buf \U$18161 ( \18185 , \18184 );
buf \U$18162 ( \18186 , \18185 );
nand \U$18163 ( \18187 , \18177 , \18186 );
buf \U$18164 ( \18188 , \18187 );
buf \U$18165 ( \18189 , \18188 );
buf \U$18166 ( \18190 , RIc0d87d0_38);
buf \U$18167 ( \18191 , RIc0da378_97);
xor \U$18168 ( \18192 , \18190 , \18191 );
buf \U$18169 ( \18193 , \18192 );
buf \U$18170 ( \18194 , \18193 );
not \U$18171 ( \18195 , \18194 );
buf \U$18172 ( \18196 , \15329 );
not \U$18173 ( \18197 , \18196 );
or \U$18174 ( \18198 , \18195 , \18197 );
buf \U$18175 ( \18199 , \2070 );
buf \U$18176 ( \18200 , RIc0d8758_37);
buf \U$18177 ( \18201 , RIc0da378_97);
xor \U$18178 ( \18202 , \18200 , \18201 );
buf \U$18179 ( \18203 , \18202 );
buf \U$18180 ( \18204 , \18203 );
nand \U$18181 ( \18205 , \18199 , \18204 );
buf \U$18182 ( \18206 , \18205 );
buf \U$18183 ( \18207 , \18206 );
nand \U$18184 ( \18208 , \18198 , \18207 );
buf \U$18185 ( \18209 , \18208 );
buf \U$18186 ( \18210 , \18209 );
or \U$18187 ( \18211 , \18189 , \18210 );
buf \U$18188 ( \18212 , RIc0d8500_32);
buf \U$18189 ( \18213 , RIc0da648_103);
xor \U$18190 ( \18214 , \18212 , \18213 );
buf \U$18191 ( \18215 , \18214 );
buf \U$18192 ( \18216 , \18215 );
not \U$18193 ( \18217 , \18216 );
buf \U$18194 ( \18218 , \4483 );
not \U$18195 ( \18219 , \18218 );
buf \U$18196 ( \18220 , \18219 );
buf \U$18197 ( \18221 , \18220 );
not \U$18198 ( \18222 , \18221 );
or \U$18199 ( \18223 , \18217 , \18222 );
buf \U$18200 ( \18224 , \13048 );
xor \U$18201 ( \18225 , RIc0da648_103, RIc0d8488_31);
buf \U$18202 ( \18226 , \18225 );
nand \U$18203 ( \18227 , \18224 , \18226 );
buf \U$18204 ( \18228 , \18227 );
buf \U$18205 ( \18229 , \18228 );
nand \U$18206 ( \18230 , \18223 , \18229 );
buf \U$18207 ( \18231 , \18230 );
buf \U$18208 ( \18232 , \18231 );
nand \U$18209 ( \18233 , \18211 , \18232 );
buf \U$18210 ( \18234 , \18233 );
buf \U$18211 ( \18235 , \18234 );
buf \U$18212 ( \18236 , \18209 );
buf \U$18213 ( \18237 , \18188 );
nand \U$18214 ( \18238 , \18236 , \18237 );
buf \U$18215 ( \18239 , \18238 );
buf \U$18216 ( \18240 , \18239 );
nand \U$18217 ( \18241 , \18235 , \18240 );
buf \U$18218 ( \18242 , \18241 );
buf \U$18219 ( \18243 , \18242 );
and \U$18220 ( \18244 , \18168 , \18243 );
and \U$18221 ( \18245 , \18091 , \18167 );
or \U$18222 ( \18246 , \18244 , \18245 );
buf \U$18223 ( \18247 , \18246 );
buf \U$18224 ( \18248 , \18247 );
and \U$18225 ( \18249 , \18048 , \18248 );
and \U$18226 ( \18250 , \18038 , \18047 );
or \U$18227 ( \18251 , \18249 , \18250 );
buf \U$18228 ( \18252 , \18251 );
buf \U$18229 ( \18253 , \18252 );
and \U$18230 ( \18254 , \17985 , \18253 );
and \U$18231 ( \18255 , \17962 , \17984 );
or \U$18232 ( \18256 , \18254 , \18255 );
buf \U$18233 ( \18257 , \18256 );
buf \U$18234 ( \18258 , \18257 );
xor \U$18235 ( \18259 , \17866 , \17855 );
xor \U$18236 ( \18260 , \18259 , \17848 );
buf \U$18237 ( \18261 , \18260 );
xor \U$18238 ( \18262 , \18258 , \18261 );
xor \U$18239 ( \18263 , \16801 , \16825 );
xor \U$18240 ( \18264 , \18263 , \16830 );
buf \U$18241 ( \18265 , \18264 );
buf \U$18242 ( \18266 , \18265 );
buf \U$18243 ( \18267 , \13837 );
not \U$18244 ( \18268 , \18267 );
buf \U$18245 ( \18269 , \2812 );
not \U$18246 ( \18270 , \18269 );
or \U$18247 ( \18271 , \18268 , \18270 );
buf \U$18248 ( \18272 , \1276 );
not \U$18249 ( \18273 , \18272 );
buf \U$18250 ( \18274 , \18273 );
buf \U$18251 ( \18275 , \18274 );
not \U$18252 ( \18276 , \18275 );
buf \U$18253 ( \18277 , \18276 );
buf \U$18254 ( \18278 , \18277 );
buf \U$18255 ( \18279 , RIc0d91a8_59);
buf \U$18256 ( \18280 , RIc0d9748_71);
xor \U$18257 ( \18281 , \18279 , \18280 );
buf \U$18258 ( \18282 , \18281 );
buf \U$18259 ( \18283 , \18282 );
nand \U$18260 ( \18284 , \18278 , \18283 );
buf \U$18261 ( \18285 , \18284 );
buf \U$18262 ( \18286 , \18285 );
nand \U$18263 ( \18287 , \18271 , \18286 );
buf \U$18264 ( \18288 , \18287 );
buf \U$18265 ( \18289 , \18288 );
buf \U$18266 ( \18290 , \14022 );
not \U$18267 ( \18291 , \18290 );
buf \U$18268 ( \18292 , \1765 );
not \U$18269 ( \18293 , \18292 );
or \U$18270 ( \18294 , \18291 , \18293 );
buf \U$18271 ( \18295 , \816 );
buf \U$18272 ( \18296 , \14315 );
nand \U$18273 ( \18297 , \18295 , \18296 );
buf \U$18274 ( \18298 , \18297 );
buf \U$18275 ( \18299 , \18298 );
nand \U$18276 ( \18300 , \18294 , \18299 );
buf \U$18277 ( \18301 , \18300 );
buf \U$18278 ( \18302 , \18301 );
xor \U$18279 ( \18303 , \18289 , \18302 );
buf \U$18280 ( \18304 , \14111 );
not \U$18281 ( \18305 , \18304 );
buf \U$18284 ( \18306 , \14346 );
buf \U$18285 ( \18307 , \18306 );
not \U$18286 ( \18308 , \18307 );
or \U$18287 ( \18309 , \18305 , \18308 );
buf \U$18288 ( \18310 , \12540 );
not \U$18289 ( \18311 , \18310 );
buf \U$18290 ( \18312 , \18311 );
buf \U$18291 ( \18313 , \18312 );
buf \U$18292 ( \18314 , \14343 );
nand \U$18293 ( \18315 , \18313 , \18314 );
buf \U$18294 ( \18316 , \18315 );
buf \U$18295 ( \18317 , \18316 );
nand \U$18296 ( \18318 , \18309 , \18317 );
buf \U$18297 ( \18319 , \18318 );
buf \U$18298 ( \18320 , \18319 );
xnor \U$18299 ( \18321 , \18303 , \18320 );
buf \U$18300 ( \18322 , \18321 );
buf \U$18301 ( \18323 , \18322 );
not \U$18302 ( \18324 , \18323 );
xor \U$18303 ( \18325 , \16736 , \16757 );
and \U$18304 ( \18326 , \18325 , \16713 );
not \U$18305 ( \18327 , \18325 );
and \U$18306 ( \18328 , \18327 , \16714 );
nor \U$18307 ( \18329 , \18326 , \18328 );
buf \U$18308 ( \18330 , \18329 );
not \U$18309 ( \18331 , \18330 );
or \U$18310 ( \18332 , \18324 , \18331 );
buf \U$18311 ( \18333 , \18329 );
not \U$18312 ( \18334 , \18333 );
buf \U$18313 ( \18335 , \18322 );
not \U$18314 ( \18336 , \18335 );
buf \U$18315 ( \18337 , \18336 );
buf \U$18316 ( \18338 , \18337 );
nand \U$18317 ( \18339 , \18334 , \18338 );
buf \U$18318 ( \18340 , \18339 );
buf \U$18319 ( \18341 , \18340 );
nand \U$18320 ( \18342 , \18332 , \18341 );
buf \U$18321 ( \18343 , \18342 );
buf \U$18322 ( \18344 , \18343 );
buf \U$18323 ( \18345 , \16543 );
not \U$18324 ( \18346 , \18345 );
buf \U$18325 ( \18347 , \16569 );
not \U$18326 ( \18348 , \18347 );
or \U$18327 ( \18349 , \18346 , \18348 );
buf \U$18328 ( \18350 , \16566 );
buf \U$18329 ( \18351 , \16546 );
nand \U$18330 ( \18352 , \18350 , \18351 );
buf \U$18331 ( \18353 , \18352 );
buf \U$18332 ( \18354 , \18353 );
nand \U$18333 ( \18355 , \18349 , \18354 );
buf \U$18334 ( \18356 , \18355 );
buf \U$18335 ( \18357 , \18356 );
buf \U$18336 ( \18358 , \16595 );
xnor \U$18337 ( \18359 , \18357 , \18358 );
buf \U$18338 ( \18360 , \18359 );
buf \U$18339 ( \18361 , \18360 );
not \U$18340 ( \18362 , \18361 );
buf \U$18341 ( \18363 , \18362 );
buf \U$18342 ( \18364 , \18363 );
and \U$18343 ( \18365 , \18344 , \18364 );
not \U$18344 ( \18366 , \18344 );
buf \U$18345 ( \18367 , \18360 );
and \U$18346 ( \18368 , \18366 , \18367 );
nor \U$18347 ( \18369 , \18365 , \18368 );
buf \U$18348 ( \18370 , \18369 );
buf \U$18349 ( \18371 , \18370 );
xor \U$18350 ( \18372 , \18266 , \18371 );
buf \U$18351 ( \18373 , \18105 );
not \U$18352 ( \18374 , \18373 );
buf \U$18353 ( \18375 , \1183 );
not \U$18354 ( \18376 , \18375 );
or \U$18355 ( \18377 , \18374 , \18376 );
buf \U$18356 ( \18378 , \14374 );
buf \U$18357 ( \18379 , \14819 );
nand \U$18358 ( \18380 , \18378 , \18379 );
buf \U$18359 ( \18381 , \18380 );
buf \U$18360 ( \18382 , \18381 );
nand \U$18361 ( \18383 , \18377 , \18382 );
buf \U$18362 ( \18384 , \18383 );
not \U$18363 ( \18385 , \18384 );
buf \U$18364 ( \18386 , \18182 );
not \U$18365 ( \18387 , \18386 );
buf \U$18366 ( \18388 , \1888 );
not \U$18367 ( \18389 , \18388 );
or \U$18368 ( \18390 , \18387 , \18389 );
buf \U$18369 ( \18391 , \2927 );
buf \U$18370 ( \18392 , \14506 );
nand \U$18371 ( \18393 , \18391 , \18392 );
buf \U$18372 ( \18394 , \18393 );
buf \U$18373 ( \18395 , \18394 );
nand \U$18374 ( \18396 , \18390 , \18395 );
buf \U$18375 ( \18397 , \18396 );
not \U$18376 ( \18398 , \18397 );
or \U$18377 ( \18399 , \18385 , \18398 );
buf \U$18378 ( \18400 , \18397 );
not \U$18379 ( \18401 , \18400 );
buf \U$18380 ( \18402 , \18401 );
not \U$18381 ( \18403 , \18402 );
buf \U$18382 ( \18404 , \18384 );
not \U$18383 ( \18405 , \18404 );
buf \U$18384 ( \18406 , \18405 );
not \U$18385 ( \18407 , \18406 );
or \U$18386 ( \18408 , \18403 , \18407 );
buf \U$18387 ( \18409 , \18225 );
not \U$18388 ( \18410 , \18409 );
buf \U$18389 ( \18411 , \15397 );
not \U$18390 ( \18412 , \18411 );
or \U$18391 ( \18413 , \18410 , \18412 );
buf \U$18392 ( \18414 , \4475 );
not \U$18393 ( \18415 , \18414 );
buf \U$18394 ( \18416 , \18415 );
buf \U$18395 ( \18417 , \18416 );
buf \U$18396 ( \18418 , \17400 );
nand \U$18397 ( \18419 , \18417 , \18418 );
buf \U$18398 ( \18420 , \18419 );
buf \U$18399 ( \18421 , \18420 );
nand \U$18400 ( \18422 , \18413 , \18421 );
buf \U$18401 ( \18423 , \18422 );
nand \U$18402 ( \18424 , \18408 , \18423 );
nand \U$18403 ( \18425 , \18399 , \18424 );
buf \U$18404 ( \18426 , \18425 );
not \U$18405 ( \18427 , \18426 );
buf \U$18406 ( \18428 , RIc0d81b8_25);
buf \U$18407 ( \18429 , RIc0da918_109);
xor \U$18408 ( \18430 , \18428 , \18429 );
buf \U$18409 ( \18431 , \18430 );
buf \U$18410 ( \18432 , \18431 );
not \U$18411 ( \18433 , \18432 );
buf \U$18412 ( \18434 , \13419 );
not \U$18413 ( \18435 , \18434 );
or \U$18414 ( \18436 , \18433 , \18435 );
buf \U$18415 ( \18437 , \13426 );
buf \U$18416 ( \18438 , \14664 );
nand \U$18417 ( \18439 , \18437 , \18438 );
buf \U$18418 ( \18440 , \18439 );
buf \U$18419 ( \18441 , \18440 );
nand \U$18420 ( \18442 , \18436 , \18441 );
buf \U$18421 ( \18443 , \18442 );
buf \U$18422 ( \18444 , RIc0d7df8_17);
buf \U$18423 ( \18445 , RIc0dacd8_117);
xor \U$18424 ( \18446 , \18444 , \18445 );
buf \U$18425 ( \18447 , \18446 );
buf \U$18426 ( \18448 , \18447 );
not \U$18427 ( \18449 , \18448 );
buf \U$18428 ( \18450 , \13684 );
not \U$18429 ( \18451 , \18450 );
or \U$18430 ( \18452 , \18449 , \18451 );
buf \U$18431 ( \18453 , \12936 );
buf \U$18432 ( \18454 , \17378 );
nand \U$18433 ( \18455 , \18453 , \18454 );
buf \U$18434 ( \18456 , \18455 );
buf \U$18435 ( \18457 , \18456 );
nand \U$18436 ( \18458 , \18452 , \18457 );
buf \U$18437 ( \18459 , \18458 );
xor \U$18438 ( \18460 , \18443 , \18459 );
buf \U$18439 ( \18461 , \14713 );
buf \U$18440 ( \18462 , RIc0d8848_39);
buf \U$18441 ( \18463 , RIc0da288_95);
xor \U$18442 ( \18464 , \18462 , \18463 );
buf \U$18443 ( \18465 , \18464 );
buf \U$18444 ( \18466 , \18465 );
not \U$18445 ( \18467 , \18466 );
buf \U$18446 ( \18468 , \18467 );
buf \U$18447 ( \18469 , \18468 );
or \U$18448 ( \18470 , \18461 , \18469 );
buf \U$18449 ( \18471 , \14704 );
buf \U$18450 ( \18472 , \14715 );
or \U$18451 ( \18473 , \18471 , \18472 );
nand \U$18452 ( \18474 , \18470 , \18473 );
buf \U$18453 ( \18475 , \18474 );
and \U$18454 ( \18476 , \18460 , \18475 );
and \U$18455 ( \18477 , \18443 , \18459 );
or \U$18456 ( \18478 , \18476 , \18477 );
buf \U$18457 ( \18479 , \18478 );
not \U$18458 ( \18480 , \18479 );
or \U$18459 ( \18481 , \18427 , \18480 );
buf \U$18460 ( \18482 , \18478 );
buf \U$18461 ( \18483 , \18425 );
or \U$18462 ( \18484 , \18482 , \18483 );
buf \U$18463 ( \18485 , \874 );
buf \U$18464 ( \18486 , RIc0d9400_64);
and \U$18465 ( \18487 , \18485 , \18486 );
buf \U$18466 ( \18488 , \18487 );
buf \U$18467 ( \18489 , \18488 );
buf \U$18468 ( \18490 , \18065 );
not \U$18469 ( \18491 , \18490 );
buf \U$18470 ( \18492 , \12442 );
not \U$18471 ( \18493 , \18492 );
or \U$18472 ( \18494 , \18491 , \18493 );
buf \U$18473 ( \18495 , \791 );
buf \U$18474 ( \18496 , \14601 );
nand \U$18475 ( \18497 , \18495 , \18496 );
buf \U$18476 ( \18498 , \18497 );
buf \U$18477 ( \18499 , \18498 );
nand \U$18478 ( \18500 , \18494 , \18499 );
buf \U$18479 ( \18501 , \18500 );
buf \U$18480 ( \18502 , \18501 );
xor \U$18481 ( \18503 , \18489 , \18502 );
buf \U$18482 ( \18504 , \18203 );
not \U$18483 ( \18505 , \18504 );
buf \U$18484 ( \18506 , \16086 );
not \U$18485 ( \18507 , \18506 );
or \U$18486 ( \18508 , \18505 , \18507 );
buf \U$18487 ( \18509 , \2070 );
buf \U$18488 ( \18510 , \17363 );
nand \U$18489 ( \18511 , \18509 , \18510 );
buf \U$18490 ( \18512 , \18511 );
buf \U$18491 ( \18513 , \18512 );
nand \U$18492 ( \18514 , \18508 , \18513 );
buf \U$18493 ( \18515 , \18514 );
buf \U$18494 ( \18516 , \18515 );
and \U$18495 ( \18517 , \18503 , \18516 );
and \U$18496 ( \18518 , \18489 , \18502 );
or \U$18497 ( \18519 , \18517 , \18518 );
buf \U$18498 ( \18520 , \18519 );
buf \U$18499 ( \18521 , \18520 );
nand \U$18500 ( \18522 , \18484 , \18521 );
buf \U$18501 ( \18523 , \18522 );
buf \U$18502 ( \18524 , \18523 );
nand \U$18503 ( \18525 , \18481 , \18524 );
buf \U$18504 ( \18526 , \18525 );
buf \U$18505 ( \18527 , \18526 );
buf \U$18506 ( \18528 , \18005 );
not \U$18507 ( \18529 , \18528 );
buf \U$18508 ( \18530 , \18529 );
buf \U$18509 ( \18531 , \18530 );
buf \U$18510 ( \18532 , \18021 );
nand \U$18511 ( \18533 , \18531 , \18532 );
buf \U$18512 ( \18534 , \18533 );
buf \U$18513 ( \18535 , \18534 );
not \U$18514 ( \18536 , \18535 );
buf \U$18515 ( \18537 , \17987 );
not \U$18516 ( \18538 , \18537 );
or \U$18517 ( \18539 , \18536 , \18538 );
buf \U$18518 ( \18540 , \18021 );
buf \U$18519 ( \18541 , \18530 );
or \U$18520 ( \18542 , \18540 , \18541 );
buf \U$18521 ( \18543 , \18542 );
buf \U$18522 ( \18544 , \18543 );
nand \U$18523 ( \18545 , \18539 , \18544 );
buf \U$18524 ( \18546 , \18545 );
buf \U$18525 ( \18547 , \18546 );
or \U$18526 ( \18548 , \18527 , \18547 );
xor \U$18527 ( \18549 , \14486 , \14522 );
xor \U$18528 ( \18550 , \18549 , \14592 );
buf \U$18529 ( \18551 , \18550 );
buf \U$18530 ( \18552 , \18551 );
nand \U$18531 ( \18553 , \18548 , \18552 );
buf \U$18532 ( \18554 , \18553 );
buf \U$18533 ( \18555 , \18554 );
buf \U$18534 ( \18556 , \18526 );
buf \U$18535 ( \18557 , \18546 );
nand \U$18536 ( \18558 , \18556 , \18557 );
buf \U$18537 ( \18559 , \18558 );
buf \U$18538 ( \18560 , \18559 );
nand \U$18539 ( \18561 , \18555 , \18560 );
buf \U$18540 ( \18562 , \18561 );
buf \U$18541 ( \18563 , \18562 );
xor \U$18542 ( \18564 , \18372 , \18563 );
buf \U$18543 ( \18565 , \18564 );
buf \U$18544 ( \18566 , \18565 );
and \U$18545 ( \18567 , \18262 , \18566 );
and \U$18546 ( \18568 , \18258 , \18261 );
or \U$18547 ( \18569 , \18567 , \18568 );
buf \U$18548 ( \18570 , \18569 );
buf \U$18549 ( \18571 , \18570 );
xor \U$18550 ( \18572 , \17945 , \18571 );
buf \U$18551 ( \18573 , \15977 );
not \U$18552 ( \18574 , \18573 );
buf \U$18553 ( \18575 , \12361 );
not \U$18554 ( \18576 , \18575 );
or \U$18555 ( \18577 , \18574 , \18576 );
buf \U$18556 ( \18578 , \1025 );
buf \U$18557 ( \18579 , \12352 );
nand \U$18558 ( \18580 , \18578 , \18579 );
buf \U$18559 ( \18581 , \18580 );
buf \U$18560 ( \18582 , \18581 );
nand \U$18561 ( \18583 , \18577 , \18582 );
buf \U$18562 ( \18584 , \18583 );
buf \U$18563 ( \18585 , \18584 );
not \U$18564 ( \18586 , \18585 );
buf \U$18565 ( \18587 , \16047 );
not \U$18566 ( \18588 , \18587 );
buf \U$18567 ( \18589 , \12654 );
not \U$18568 ( \18590 , \18589 );
or \U$18569 ( \18591 , \18588 , \18590 );
buf \U$18570 ( \18592 , \12642 );
buf \U$18571 ( \18593 , RIc0db200_128);
nand \U$18572 ( \18594 , \18592 , \18593 );
buf \U$18573 ( \18595 , \18594 );
buf \U$18574 ( \18596 , \18595 );
nand \U$18575 ( \18597 , \18591 , \18596 );
buf \U$18576 ( \18598 , \18597 );
buf \U$18577 ( \18599 , \18598 );
not \U$18578 ( \18600 , \18599 );
buf \U$18579 ( \18601 , \18600 );
buf \U$18580 ( \18602 , \18601 );
not \U$18581 ( \18603 , \18602 );
buf \U$18582 ( \18604 , \15650 );
not \U$18583 ( \18605 , \18604 );
buf \U$18584 ( \18606 , \12731 );
buf \U$18585 ( \18607 , \16022 );
and \U$18586 ( \18608 , \18606 , \18607 );
buf \U$18587 ( \18609 , \18608 );
buf \U$18588 ( \18610 , \18609 );
not \U$18589 ( \18611 , \18610 );
or \U$18590 ( \18612 , \18605 , \18611 );
buf \U$18591 ( \18613 , \12743 );
buf \U$18592 ( \18614 , \12725 );
nand \U$18593 ( \18615 , \18613 , \18614 );
buf \U$18594 ( \18616 , \18615 );
buf \U$18595 ( \18617 , \18616 );
nand \U$18596 ( \18618 , \18612 , \18617 );
buf \U$18597 ( \18619 , \18618 );
buf \U$18598 ( \18620 , \18619 );
not \U$18599 ( \18621 , \18620 );
and \U$18600 ( \18622 , \18603 , \18621 );
buf \U$18601 ( \18623 , \18601 );
buf \U$18602 ( \18624 , \18619 );
and \U$18603 ( \18625 , \18623 , \18624 );
nor \U$18604 ( \18626 , \18622 , \18625 );
buf \U$18605 ( \18627 , \18626 );
buf \U$18606 ( \18628 , \18627 );
not \U$18607 ( \18629 , \18628 );
or \U$18608 ( \18630 , \18586 , \18629 );
buf \U$18609 ( \18631 , \18627 );
buf \U$18610 ( \18632 , \18584 );
or \U$18611 ( \18633 , \18631 , \18632 );
nand \U$18612 ( \18634 , \18630 , \18633 );
buf \U$18613 ( \18635 , \18634 );
buf \U$18614 ( \18636 , \18635 );
buf \U$18615 ( \18637 , \16482 );
not \U$18616 ( \18638 , \18637 );
buf \U$18617 ( \18639 , \841 );
not \U$18618 ( \18640 , \18639 );
or \U$18619 ( \18641 , \18638 , \18640 );
buf \U$18620 ( \18642 , \441 );
buf \U$18621 ( \18643 , \13486 );
nand \U$18622 ( \18644 , \18642 , \18643 );
buf \U$18623 ( \18645 , \18644 );
buf \U$18624 ( \18646 , \18645 );
nand \U$18625 ( \18647 , \18641 , \18646 );
buf \U$18626 ( \18648 , \18647 );
buf \U$18627 ( \18649 , \18648 );
not \U$18628 ( \18650 , \16516 );
not \U$18629 ( \18651 , \3714 );
or \U$18630 ( \18652 , \18650 , \18651 );
buf \U$18631 ( \18653 , \344 );
buf \U$18632 ( \18654 , \12700 );
nand \U$18633 ( \18655 , \18653 , \18654 );
buf \U$18634 ( \18656 , \18655 );
nand \U$18635 ( \18657 , \18652 , \18656 );
buf \U$18636 ( \18658 , \18657 );
xor \U$18637 ( \18659 , \18649 , \18658 );
buf \U$18638 ( \18660 , \16589 );
not \U$18639 ( \18661 , \18660 );
buf \U$18640 ( \18662 , \17405 );
not \U$18641 ( \18663 , \18662 );
or \U$18642 ( \18664 , \18661 , \18663 );
buf \U$18643 ( \18665 , \18416 );
buf \U$18644 ( \18666 , \13037 );
nand \U$18645 ( \18667 , \18665 , \18666 );
buf \U$18646 ( \18668 , \18667 );
buf \U$18647 ( \18669 , \18668 );
nand \U$18648 ( \18670 , \18664 , \18669 );
buf \U$18649 ( \18671 , \18670 );
buf \U$18650 ( \18672 , \18671 );
xor \U$18651 ( \18673 , \18659 , \18672 );
buf \U$18652 ( \18674 , \18673 );
buf \U$18653 ( \18675 , \18674 );
xor \U$18654 ( \18676 , \18636 , \18675 );
buf \U$18655 ( \18677 , \769 );
buf \U$18656 ( \18678 , \16133 );
nand \U$18657 ( \18679 , \18677 , \18678 );
buf \U$18658 ( \18680 , \18679 );
buf \U$18659 ( \18681 , \18680 );
buf \U$18660 ( \18682 , \1856 );
or \U$18661 ( \18683 , \18681 , \18682 );
buf \U$18662 ( \18684 , \791 );
buf \U$18663 ( \18685 , \12437 );
nand \U$18664 ( \18686 , \18684 , \18685 );
buf \U$18665 ( \18687 , \18686 );
buf \U$18666 ( \18688 , \18687 );
nand \U$18667 ( \18689 , \18683 , \18688 );
buf \U$18668 ( \18690 , \18689 );
buf \U$18669 ( \18691 , \18690 );
buf \U$18670 ( \18692 , \13443 );
not \U$18671 ( \18693 , \18692 );
buf \U$18672 ( \18694 , \15793 );
not \U$18673 ( \18695 , \18694 );
or \U$18674 ( \18696 , \18693 , \18695 );
buf \U$18675 ( \18697 , \13465 );
not \U$18676 ( \18698 , \18697 );
buf \U$18677 ( \18699 , \18698 );
buf \U$18678 ( \18700 , \18699 );
buf \U$18679 ( \18701 , \16155 );
buf \U$18680 ( \18702 , \13454 );
buf \U$18681 ( \18703 , \18702 );
nand \U$18682 ( \18704 , \18700 , \18701 , \18703 );
buf \U$18683 ( \18705 , \18704 );
buf \U$18684 ( \18706 , \18705 );
nand \U$18685 ( \18707 , \18696 , \18706 );
buf \U$18686 ( \18708 , \18707 );
buf \U$18687 ( \18709 , \18708 );
xor \U$18688 ( \18710 , \18691 , \18709 );
buf \U$18689 ( \18711 , \16216 );
not \U$18690 ( \18712 , \18711 );
buf \U$18691 ( \18713 , \14186 );
not \U$18692 ( \18714 , \18713 );
or \U$18693 ( \18715 , \18712 , \18714 );
buf \U$18694 ( \18716 , \12303 );
buf \U$18695 ( \18717 , \12269 );
nand \U$18696 ( \18718 , \18716 , \18717 );
buf \U$18697 ( \18719 , \18718 );
buf \U$18698 ( \18720 , \18719 );
nand \U$18699 ( \18721 , \18715 , \18720 );
buf \U$18700 ( \18722 , \18721 );
buf \U$18701 ( \18723 , \18722 );
xor \U$18702 ( \18724 , \18710 , \18723 );
buf \U$18703 ( \18725 , \18724 );
buf \U$18704 ( \18726 , \18725 );
xor \U$18705 ( \18727 , \18676 , \18726 );
buf \U$18706 ( \18728 , \18727 );
buf \U$18707 ( \18729 , \18728 );
buf \U$18708 ( \18730 , \18363 );
not \U$18709 ( \18731 , \18730 );
buf \U$18710 ( \18732 , \18337 );
not \U$18711 ( \18733 , \18732 );
or \U$18712 ( \18734 , \18731 , \18733 );
buf \U$18713 ( \18735 , \18360 );
not \U$18714 ( \18736 , \18735 );
buf \U$18715 ( \18737 , \18322 );
not \U$18716 ( \18738 , \18737 );
or \U$18717 ( \18739 , \18736 , \18738 );
buf \U$18718 ( \18740 , \18329 );
nand \U$18719 ( \18741 , \18739 , \18740 );
buf \U$18720 ( \18742 , \18741 );
buf \U$18721 ( \18743 , \18742 );
nand \U$18722 ( \18744 , \18734 , \18743 );
buf \U$18723 ( \18745 , \18744 );
buf \U$18724 ( \18746 , \18745 );
xor \U$18725 ( \18747 , \18729 , \18746 );
buf \U$18726 ( \18748 , \18301 );
buf \U$18727 ( \18749 , \18288 );
or \U$18728 ( \18750 , \18748 , \18749 );
buf \U$18729 ( \18751 , \18319 );
nand \U$18730 ( \18752 , \18750 , \18751 );
buf \U$18731 ( \18753 , \18752 );
buf \U$18732 ( \18754 , \18753 );
buf \U$18733 ( \18755 , \18301 );
buf \U$18734 ( \18756 , \18288 );
nand \U$18735 ( \18757 , \18755 , \18756 );
buf \U$18736 ( \18758 , \18757 );
buf \U$18737 ( \18759 , \18758 );
nand \U$18738 ( \18760 , \18754 , \18759 );
buf \U$18739 ( \18761 , \18760 );
buf \U$18740 ( \18762 , \18761 );
buf \U$18741 ( \18763 , \16199 );
not \U$18742 ( \18764 , \18763 );
buf \U$18743 ( \18765 , \948 );
not \U$18744 ( \18766 , \18765 );
buf \U$18745 ( \18767 , \18766 );
buf \U$18746 ( \18768 , \18767 );
not \U$18747 ( \18769 , \18768 );
or \U$18748 ( \18770 , \18764 , \18769 );
buf \U$18749 ( \18771 , \17010 );
buf \U$18750 ( \18772 , \12483 );
nand \U$18751 ( \18773 , \18771 , \18772 );
buf \U$18752 ( \18774 , \18773 );
buf \U$18753 ( \18775 , \18774 );
nand \U$18754 ( \18776 , \18770 , \18775 );
buf \U$18755 ( \18777 , \18776 );
buf \U$18756 ( \18778 , \18777 );
buf \U$18757 ( \18779 , \16244 );
not \U$18758 ( \18780 , \18779 );
buf \U$18759 ( \18781 , \14210 );
not \U$18760 ( \18782 , \18781 );
or \U$18761 ( \18783 , \18780 , \18782 );
buf \U$18762 ( \18784 , \15909 );
buf \U$18763 ( \18785 , \13402 );
nand \U$18764 ( \18786 , \18784 , \18785 );
buf \U$18765 ( \18787 , \18786 );
buf \U$18766 ( \18788 , \18787 );
nand \U$18767 ( \18789 , \18783 , \18788 );
buf \U$18768 ( \18790 , \18789 );
buf \U$18769 ( \18791 , \18790 );
xor \U$18770 ( \18792 , \18778 , \18791 );
not \U$18771 ( \18793 , \1282 );
not \U$18772 ( \18794 , \12673 );
or \U$18773 ( \18795 , \18793 , \18794 );
buf \U$18774 ( \18796 , \18282 );
not \U$18775 ( \18797 , \18796 );
buf \U$18776 ( \18798 , \18797 );
or \U$18777 ( \18799 , \2815 , \18798 );
nand \U$18778 ( \18800 , \18795 , \18799 );
buf \U$18779 ( \18801 , \18800 );
xnor \U$18780 ( \18802 , \18792 , \18801 );
buf \U$18781 ( \18803 , \18802 );
not \U$18782 ( \18804 , \18803 );
buf \U$18783 ( \18805 , \18804 );
xor \U$18784 ( \18806 , \18762 , \18805 );
xor \U$18785 ( \18807 , \13549 , \13562 );
xor \U$18786 ( \18808 , \18807 , \13580 );
buf \U$18787 ( \18809 , \18808 );
buf \U$18788 ( \18810 , \18809 );
xor \U$18789 ( \18811 , \18806 , \18810 );
buf \U$18790 ( \18812 , \18811 );
buf \U$18791 ( \18813 , \18812 );
xor \U$18792 ( \18814 , \18747 , \18813 );
buf \U$18793 ( \18815 , \18814 );
buf \U$18794 ( \18816 , \18815 );
xor \U$18795 ( \18817 , \14457 , \14461 );
xor \U$18796 ( \18818 , \18817 , \15018 );
buf \U$18797 ( \18819 , \18818 );
buf \U$18798 ( \18820 , \18819 );
xor \U$18799 ( \18821 , \18816 , \18820 );
xor \U$18800 ( \18822 , \18266 , \18371 );
and \U$18801 ( \18823 , \18822 , \18563 );
and \U$18802 ( \18824 , \18266 , \18371 );
or \U$18803 ( \18825 , \18823 , \18824 );
buf \U$18804 ( \18826 , \18825 );
buf \U$18805 ( \18827 , \18826 );
xor \U$18806 ( \18828 , \18821 , \18827 );
buf \U$18807 ( \18829 , \18828 );
buf \U$18808 ( \18830 , \18829 );
and \U$18809 ( \18831 , \18572 , \18830 );
and \U$18810 ( \18832 , \17945 , \18571 );
or \U$18811 ( \18833 , \18831 , \18832 );
buf \U$18812 ( \18834 , \18833 );
buf \U$18813 ( \18835 , \18834 );
and \U$18814 ( \18836 , \17923 , \18835 );
and \U$18815 ( \18837 , \17839 , \17922 );
or \U$18816 ( \18838 , \18836 , \18837 );
buf \U$18817 ( \18839 , \18838 );
buf \U$18818 ( \18840 , \18839 );
xor \U$18819 ( \18841 , \16869 , \18840 );
xor \U$18820 ( \18842 , \17845 , \17914 );
and \U$18821 ( \18843 , \18842 , \17919 );
and \U$18822 ( \18844 , \17845 , \17914 );
or \U$18823 ( \18845 , \18843 , \18844 );
buf \U$18824 ( \18846 , \18845 );
buf \U$18825 ( \18847 , \18846 );
buf \U$18826 ( \18848 , \18598 );
not \U$18827 ( \18849 , \18848 );
buf \U$18828 ( \18850 , \18619 );
not \U$18829 ( \18851 , \18850 );
or \U$18830 ( \18852 , \18849 , \18851 );
buf \U$18831 ( \18853 , \18619 );
not \U$18832 ( \18854 , \18853 );
buf \U$18833 ( \18855 , \18601 );
nand \U$18834 ( \18856 , \18854 , \18855 );
buf \U$18835 ( \18857 , \18856 );
buf \U$18836 ( \18858 , \18857 );
buf \U$18837 ( \18859 , \18584 );
nand \U$18838 ( \18860 , \18858 , \18859 );
buf \U$18839 ( \18861 , \18860 );
buf \U$18840 ( \18862 , \18861 );
nand \U$18841 ( \18863 , \18852 , \18862 );
buf \U$18842 ( \18864 , \18863 );
buf \U$18843 ( \18865 , \18864 );
buf \U$18844 ( \18866 , \18690 );
not \U$18845 ( \18867 , \18866 );
buf \U$18846 ( \18868 , \18867 );
buf \U$18847 ( \18869 , \18868 );
buf \U$18848 ( \18870 , \18708 );
not \U$18849 ( \18871 , \18870 );
buf \U$18850 ( \18872 , \18871 );
buf \U$18851 ( \18873 , \18872 );
nand \U$18852 ( \18874 , \18869 , \18873 );
buf \U$18853 ( \18875 , \18874 );
buf \U$18854 ( \18876 , \18875 );
not \U$18855 ( \18877 , \18876 );
buf \U$18856 ( \18878 , \18722 );
not \U$18857 ( \18879 , \18878 );
or \U$18858 ( \18880 , \18877 , \18879 );
buf \U$18859 ( \18881 , \18690 );
buf \U$18860 ( \18882 , \18708 );
nand \U$18861 ( \18883 , \18881 , \18882 );
buf \U$18862 ( \18884 , \18883 );
buf \U$18863 ( \18885 , \18884 );
nand \U$18864 ( \18886 , \18880 , \18885 );
buf \U$18865 ( \18887 , \18886 );
buf \U$18866 ( \18888 , \18887 );
xor \U$18867 ( \18889 , \18865 , \18888 );
xor \U$18868 ( \18890 , \13239 , \13256 );
and \U$18869 ( \18891 , \18890 , \13279 );
and \U$18870 ( \18892 , \13239 , \13256 );
or \U$18871 ( \18893 , \18891 , \18892 );
buf \U$18872 ( \18894 , \18893 );
buf \U$18873 ( \18895 , \18894 );
xor \U$18874 ( \18896 , \18889 , \18895 );
buf \U$18875 ( \18897 , \18896 );
buf \U$18876 ( \18898 , \18897 );
not \U$18877 ( \18899 , \18761 );
nand \U$18878 ( \18900 , \18899 , \18803 );
not \U$18879 ( \18901 , \18900 );
not \U$18880 ( \18902 , \18809 );
or \U$18881 ( \18903 , \18901 , \18902 );
buf \U$18882 ( \18904 , \18804 );
buf \U$18883 ( \18905 , \18761 );
nand \U$18884 ( \18906 , \18904 , \18905 );
buf \U$18885 ( \18907 , \18906 );
nand \U$18886 ( \18908 , \18903 , \18907 );
buf \U$18887 ( \18909 , \18908 );
or \U$18888 ( \18910 , \18898 , \18909 );
buf \U$18889 ( \18911 , \14309 );
not \U$18890 ( \18912 , \18911 );
buf \U$18891 ( \18913 , \18912 );
buf \U$18892 ( \18914 , \18913 );
not \U$18893 ( \18915 , \18914 );
buf \U$18894 ( \18916 , \14449 );
not \U$18895 ( \18917 , \18916 );
or \U$18896 ( \18918 , \18915 , \18917 );
buf \U$18897 ( \18919 , \14309 );
not \U$18898 ( \18920 , \18919 );
buf \U$18899 ( \18921 , \14446 );
not \U$18900 ( \18922 , \18921 );
or \U$18901 ( \18923 , \18920 , \18922 );
buf \U$18902 ( \18924 , \14384 );
nand \U$18903 ( \18925 , \18923 , \18924 );
buf \U$18904 ( \18926 , \18925 );
buf \U$18905 ( \18927 , \18926 );
nand \U$18906 ( \18928 , \18918 , \18927 );
buf \U$18907 ( \18929 , \18928 );
buf \U$18908 ( \18930 , \18929 );
nand \U$18909 ( \18931 , \18910 , \18930 );
buf \U$18910 ( \18932 , \18931 );
buf \U$18911 ( \18933 , \18932 );
buf \U$18912 ( \18934 , \18897 );
buf \U$18913 ( \18935 , \18908 );
nand \U$18914 ( \18936 , \18934 , \18935 );
buf \U$18915 ( \18937 , \18936 );
buf \U$18916 ( \18938 , \18937 );
nand \U$18917 ( \18939 , \18933 , \18938 );
buf \U$18918 ( \18940 , \18939 );
buf \U$18919 ( \18941 , \18940 );
xor \U$18920 ( \18942 , \18865 , \18888 );
and \U$18921 ( \18943 , \18942 , \18895 );
and \U$18922 ( \18944 , \18865 , \18888 );
or \U$18923 ( \18945 , \18943 , \18944 );
buf \U$18924 ( \18946 , \18945 );
buf \U$18925 ( \18947 , \18946 );
buf \U$18926 ( \18948 , \13156 );
not \U$18927 ( \18949 , \18948 );
buf \U$18928 ( \18950 , \13191 );
not \U$18929 ( \18951 , \18950 );
or \U$18930 ( \18952 , \18949 , \18951 );
buf \U$18931 ( \18953 , \13191 );
buf \U$18932 ( \18954 , \13156 );
or \U$18933 ( \18955 , \18953 , \18954 );
buf \U$18934 ( \18956 , \13209 );
nand \U$18935 ( \18957 , \18955 , \18956 );
buf \U$18936 ( \18958 , \18957 );
buf \U$18937 ( \18959 , \18958 );
nand \U$18938 ( \18960 , \18952 , \18959 );
buf \U$18939 ( \18961 , \18960 );
buf \U$18940 ( \18962 , \18961 );
xor \U$18941 ( \18963 , \18649 , \18658 );
and \U$18942 ( \18964 , \18963 , \18672 );
and \U$18943 ( \18965 , \18649 , \18658 );
or \U$18944 ( \18966 , \18964 , \18965 );
buf \U$18945 ( \18967 , \18966 );
buf \U$18946 ( \18968 , \18967 );
or \U$18947 ( \18969 , \18962 , \18968 );
buf \U$18948 ( \18970 , \18777 );
not \U$18949 ( \18971 , \18970 );
buf \U$18950 ( \18972 , \18800 );
not \U$18951 ( \18973 , \18972 );
or \U$18952 ( \18974 , \18971 , \18973 );
buf \U$18953 ( \18975 , \18800 );
buf \U$18954 ( \18976 , \18777 );
or \U$18955 ( \18977 , \18975 , \18976 );
buf \U$18956 ( \18978 , \18790 );
nand \U$18957 ( \18979 , \18977 , \18978 );
buf \U$18958 ( \18980 , \18979 );
buf \U$18959 ( \18981 , \18980 );
nand \U$18960 ( \18982 , \18974 , \18981 );
buf \U$18961 ( \18983 , \18982 );
buf \U$18962 ( \18984 , \18983 );
nand \U$18963 ( \18985 , \18969 , \18984 );
buf \U$18964 ( \18986 , \18985 );
buf \U$18965 ( \18987 , \18986 );
buf \U$18966 ( \18988 , \18961 );
buf \U$18967 ( \18989 , \18967 );
nand \U$18968 ( \18990 , \18988 , \18989 );
buf \U$18969 ( \18991 , \18990 );
buf \U$18970 ( \18992 , \18991 );
nand \U$18971 ( \18993 , \18987 , \18992 );
buf \U$18972 ( \18994 , \18993 );
buf \U$18973 ( \18995 , \18994 );
xor \U$18974 ( \18996 , \18947 , \18995 );
and \U$18975 ( \18997 , \13523 , \13540 );
buf \U$18976 ( \18998 , \18997 );
buf \U$18977 ( \18999 , \18998 );
buf \U$18978 ( \19000 , \12986 );
not \U$18979 ( \19001 , \19000 );
buf \U$18980 ( \19002 , \13016 );
not \U$18981 ( \19003 , \19002 );
or \U$18982 ( \19004 , \19001 , \19003 );
buf \U$18983 ( \19005 , \13059 );
buf \U$18984 ( \19006 , \13025 );
buf \U$18985 ( \19007 , \13019 );
nand \U$18986 ( \19008 , \19006 , \19007 );
buf \U$18987 ( \19009 , \19008 );
buf \U$18988 ( \19010 , \19009 );
nand \U$18989 ( \19011 , \19005 , \19010 );
buf \U$18990 ( \19012 , \19011 );
buf \U$18991 ( \19013 , \19012 );
nand \U$18992 ( \19014 , \19004 , \19013 );
buf \U$18993 ( \19015 , \19014 );
buf \U$18994 ( \19016 , \19015 );
xor \U$18995 ( \19017 , \18999 , \19016 );
buf \U$18996 ( \19018 , \13106 );
buf \U$18997 ( \19019 , \13086 );
nor \U$18998 ( \19020 , \19018 , \19019 );
buf \U$18999 ( \19021 , \19020 );
buf \U$19000 ( \19022 , \19021 );
buf \U$19001 ( \19023 , \13130 );
not \U$19002 ( \19024 , \19023 );
buf \U$19003 ( \19025 , \19024 );
buf \U$19004 ( \19026 , \19025 );
or \U$19005 ( \19027 , \19022 , \19026 );
buf \U$19006 ( \19028 , \13106 );
buf \U$19007 ( \19029 , \13086 );
nand \U$19008 ( \19030 , \19028 , \19029 );
buf \U$19009 ( \19031 , \19030 );
buf \U$19010 ( \19032 , \19031 );
nand \U$19011 ( \19033 , \19027 , \19032 );
buf \U$19012 ( \19034 , \19033 );
buf \U$19013 ( \19035 , \19034 );
xor \U$19014 ( \19036 , \19017 , \19035 );
buf \U$19015 ( \19037 , \19036 );
buf \U$19016 ( \19038 , \19037 );
xor \U$19017 ( \19039 , \18996 , \19038 );
buf \U$19018 ( \19040 , \19039 );
buf \U$19019 ( \19041 , \19040 );
xor \U$19020 ( \19042 , \18941 , \19041 );
buf \U$19021 ( \19043 , \12882 );
not \U$19022 ( \19044 , \19043 );
buf \U$19023 ( \19045 , \14982 );
not \U$19024 ( \19046 , \19045 );
or \U$19025 ( \19047 , \19044 , \19046 );
buf \U$19026 ( \19048 , \16692 );
xor \U$19027 ( \19049 , RIc0dafa8_123, RIc0d77e0_4);
buf \U$19028 ( \19050 , \19049 );
nand \U$19029 ( \19051 , \19048 , \19050 );
buf \U$19030 ( \19052 , \19051 );
buf \U$19031 ( \19053 , \19052 );
nand \U$19032 ( \19054 , \19047 , \19053 );
buf \U$19033 ( \19055 , \19054 );
buf \U$19034 ( \19056 , \12589 );
not \U$19035 ( \19057 , \19056 );
buf \U$19036 ( \19058 , \12578 );
not \U$19037 ( \19059 , \19058 );
or \U$19038 ( \19060 , \19057 , \19059 );
buf \U$19039 ( \19061 , \14140 );
xor \U$19040 ( \19062 , RIc0da468_99, RIc0d8320_28);
buf \U$19041 ( \19063 , \19062 );
nand \U$19042 ( \19064 , \19061 , \19063 );
buf \U$19043 ( \19065 , \19064 );
buf \U$19044 ( \19066 , \19065 );
nand \U$19045 ( \19067 , \19060 , \19066 );
buf \U$19046 ( \19068 , \19067 );
xor \U$19047 ( \19069 , \19055 , \19068 );
buf \U$19048 ( \19070 , \12629 );
not \U$19049 ( \19071 , \19070 );
buf \U$19050 ( \19072 , \14325 );
not \U$19051 ( \19073 , \19072 );
or \U$19052 ( \19074 , \19071 , \19073 );
buf \U$19053 ( \19075 , \14331 );
xor \U$19054 ( \19076 , RIc0d9ec8_87, RIc0d88c0_40);
buf \U$19055 ( \19077 , \19076 );
nand \U$19056 ( \19078 , \19075 , \19077 );
buf \U$19057 ( \19079 , \19078 );
buf \U$19058 ( \19080 , \19079 );
nand \U$19059 ( \19081 , \19074 , \19080 );
buf \U$19060 ( \19082 , \19081 );
xor \U$19061 ( \19083 , \19069 , \19082 );
buf \U$19062 ( \19084 , \19083 );
xor \U$19063 ( \19085 , \13507 , \13543 );
and \U$19064 ( \19086 , \19085 , \13585 );
and \U$19065 ( \19087 , \13507 , \13543 );
or \U$19066 ( \19088 , \19086 , \19087 );
buf \U$19067 ( \19089 , \19088 );
buf \U$19068 ( \19090 , \19089 );
xor \U$19069 ( \19091 , \19084 , \19090 );
buf \U$19070 ( \19092 , \14412 );
not \U$19071 ( \19093 , \19092 );
buf \U$19072 ( \19094 , \14445 );
not \U$19073 ( \19095 , \19094 );
or \U$19074 ( \19096 , \19093 , \19095 );
buf \U$19075 ( \19097 , \14445 );
buf \U$19076 ( \19098 , \14412 );
or \U$19077 ( \19099 , \19097 , \19098 );
buf \U$19078 ( \19100 , \14429 );
nand \U$19079 ( \19101 , \19099 , \19100 );
buf \U$19080 ( \19102 , \19101 );
buf \U$19081 ( \19103 , \19102 );
nand \U$19082 ( \19104 , \19096 , \19103 );
buf \U$19083 ( \19105 , \19104 );
buf \U$19084 ( \19106 , \19105 );
xor \U$19085 ( \19107 , \14339 , \14361 );
and \U$19086 ( \19108 , \19107 , \14382 );
and \U$19087 ( \19109 , \14339 , \14361 );
or \U$19088 ( \19110 , \19108 , \19109 );
buf \U$19089 ( \19111 , \19110 );
buf \U$19090 ( \19112 , \19111 );
nor \U$19091 ( \19113 , \19106 , \19112 );
buf \U$19092 ( \19114 , \19113 );
buf \U$19093 ( \19115 , \19114 );
buf \U$19094 ( \19116 , \14263 );
not \U$19095 ( \19117 , \19116 );
buf \U$19096 ( \19118 , \19117 );
buf \U$19097 ( \19119 , \19118 );
not \U$19098 ( \19120 , \19119 );
buf \U$19099 ( \19121 , \14305 );
not \U$19100 ( \19122 , \19121 );
or \U$19101 ( \19123 , \19120 , \19122 );
buf \U$19102 ( \19124 , \14285 );
nand \U$19103 ( \19125 , \19123 , \19124 );
buf \U$19104 ( \19126 , \19125 );
buf \U$19105 ( \19127 , \19126 );
buf \U$19106 ( \19128 , \14302 );
buf \U$19107 ( \19129 , \14263 );
nand \U$19108 ( \19130 , \19128 , \19129 );
buf \U$19109 ( \19131 , \19130 );
buf \U$19110 ( \19132 , \19131 );
nand \U$19111 ( \19133 , \19127 , \19132 );
buf \U$19112 ( \19134 , \19133 );
buf \U$19113 ( \19135 , \19134 );
not \U$19114 ( \19136 , \19135 );
buf \U$19115 ( \19137 , \19136 );
buf \U$19116 ( \19138 , \19137 );
or \U$19117 ( \19139 , \19115 , \19138 );
buf \U$19118 ( \19140 , \19105 );
buf \U$19119 ( \19141 , \19111 );
nand \U$19120 ( \19142 , \19140 , \19141 );
buf \U$19121 ( \19143 , \19142 );
buf \U$19122 ( \19144 , \19143 );
nand \U$19123 ( \19145 , \19139 , \19144 );
buf \U$19124 ( \19146 , \19145 );
buf \U$19125 ( \19147 , \19146 );
xor \U$19126 ( \19148 , \19091 , \19147 );
buf \U$19127 ( \19149 , \19148 );
buf \U$19128 ( \19150 , \19149 );
xor \U$19129 ( \19151 , \19042 , \19150 );
buf \U$19130 ( \19152 , \19151 );
buf \U$19131 ( \19153 , \19152 );
not \U$19132 ( \19154 , \19153 );
buf \U$19133 ( \19155 , \16644 );
not \U$19134 ( \19156 , \19155 );
buf \U$19135 ( \19157 , \16637 );
not \U$19136 ( \19158 , \19157 );
or \U$19137 ( \19159 , \19156 , \19158 );
buf \U$19138 ( \19160 , \16780 );
nand \U$19139 ( \19161 , \19159 , \19160 );
buf \U$19140 ( \19162 , \19161 );
buf \U$19141 ( \19163 , \19162 );
buf \U$19142 ( \19164 , \16634 );
buf \U$19143 ( \19165 , \16469 );
nand \U$19144 ( \19166 , \19164 , \19165 );
buf \U$19145 ( \19167 , \19166 );
buf \U$19146 ( \19168 , \19167 );
nand \U$19147 ( \19169 , \19163 , \19168 );
buf \U$19148 ( \19170 , \19169 );
buf \U$19149 ( \19171 , \19170 );
not \U$19150 ( \19172 , \19171 );
buf \U$19151 ( \19173 , \19172 );
buf \U$19152 ( \19174 , \19173 );
xor \U$19153 ( \19175 , \13374 , \13480 );
and \U$19154 ( \19176 , \19175 , \13588 );
and \U$19155 ( \19177 , \13374 , \13480 );
or \U$19156 ( \19178 , \19176 , \19177 );
buf \U$19157 ( \19179 , \19178 );
buf \U$19158 ( \19180 , \19179 );
not \U$19159 ( \19181 , \19180 );
buf \U$19160 ( \19182 , \19181 );
buf \U$19161 ( \19183 , \19182 );
and \U$19162 ( \19184 , \19174 , \19183 );
not \U$19163 ( \19185 , \19174 );
buf \U$19164 ( \19186 , \19179 );
and \U$19165 ( \19187 , \19185 , \19186 );
nor \U$19166 ( \19188 , \19184 , \19187 );
buf \U$19167 ( \19189 , \19188 );
buf \U$19168 ( \19190 , \19189 );
xor \U$19169 ( \19191 , \18636 , \18675 );
and \U$19170 ( \19192 , \19191 , \18726 );
and \U$19171 ( \19193 , \18636 , \18675 );
or \U$19172 ( \19194 , \19192 , \19193 );
buf \U$19173 ( \19195 , \19194 );
buf \U$19174 ( \19196 , \19195 );
buf \U$19175 ( \19197 , \18983 );
not \U$19176 ( \19198 , \19197 );
buf \U$19177 ( \19199 , \18961 );
not \U$19178 ( \19200 , \19199 );
buf \U$19179 ( \19201 , \19200 );
buf \U$19180 ( \19202 , \19201 );
not \U$19181 ( \19203 , \19202 );
or \U$19182 ( \19204 , \19198 , \19203 );
buf \U$19183 ( \19205 , \19201 );
buf \U$19184 ( \19206 , \18983 );
or \U$19185 ( \19207 , \19205 , \19206 );
nand \U$19186 ( \19208 , \19204 , \19207 );
buf \U$19187 ( \19209 , \19208 );
buf \U$19188 ( \19210 , \19209 );
buf \U$19189 ( \19211 , \18967 );
and \U$19190 ( \19212 , \19210 , \19211 );
not \U$19191 ( \19213 , \19210 );
buf \U$19192 ( \19214 , \18967 );
not \U$19193 ( \19215 , \19214 );
buf \U$19194 ( \19216 , \19215 );
buf \U$19195 ( \19217 , \19216 );
and \U$19196 ( \19218 , \19213 , \19217 );
nor \U$19197 ( \19219 , \19212 , \19218 );
buf \U$19198 ( \19220 , \19219 );
buf \U$19199 ( \19221 , \19220 );
xor \U$19200 ( \19222 , \19196 , \19221 );
xor \U$19201 ( \19223 , \19111 , \19105 );
buf \U$19202 ( \19224 , \19223 );
buf \U$19203 ( \19225 , \19134 );
and \U$19204 ( \19226 , \19224 , \19225 );
not \U$19205 ( \19227 , \19224 );
buf \U$19206 ( \19228 , \19137 );
and \U$19207 ( \19229 , \19227 , \19228 );
nor \U$19208 ( \19230 , \19226 , \19229 );
buf \U$19209 ( \19231 , \19230 );
buf \U$19210 ( \19232 , \19231 );
and \U$19211 ( \19233 , \19222 , \19232 );
and \U$19212 ( \19234 , \19196 , \19221 );
or \U$19213 ( \19235 , \19233 , \19234 );
buf \U$19214 ( \19236 , \19235 );
buf \U$19215 ( \19237 , \19236 );
not \U$19216 ( \19238 , \19237 );
buf \U$19217 ( \19239 , \19238 );
buf \U$19218 ( \19240 , \19239 );
and \U$19219 ( \19241 , \19190 , \19240 );
not \U$19220 ( \19242 , \19190 );
buf \U$19221 ( \19243 , \19236 );
and \U$19222 ( \19244 , \19242 , \19243 );
nor \U$19223 ( \19245 , \19241 , \19244 );
buf \U$19224 ( \19246 , \19245 );
buf \U$19225 ( \19247 , \19246 );
not \U$19226 ( \19248 , \19247 );
or \U$19227 ( \19249 , \19154 , \19248 );
buf \U$19228 ( \19250 , \19246 );
buf \U$19229 ( \19251 , \19152 );
or \U$19230 ( \19252 , \19250 , \19251 );
nand \U$19231 ( \19253 , \19249 , \19252 );
buf \U$19232 ( \19254 , \19253 );
buf \U$19233 ( \19255 , \19254 );
xor \U$19234 ( \19256 , \19196 , \19221 );
xor \U$19235 ( \19257 , \19256 , \19232 );
buf \U$19236 ( \19258 , \19257 );
buf \U$19237 ( \19259 , \19258 );
xor \U$19238 ( \19260 , \18729 , \18746 );
and \U$19239 ( \19261 , \19260 , \18813 );
and \U$19240 ( \19262 , \18729 , \18746 );
or \U$19241 ( \19263 , \19261 , \19262 );
buf \U$19242 ( \19264 , \19263 );
buf \U$19243 ( \19265 , \19264 );
xor \U$19244 ( \19266 , \19259 , \19265 );
xor \U$19245 ( \19267 , \18908 , \18929 );
xor \U$19246 ( \19268 , \19267 , \18897 );
buf \U$19247 ( \19269 , \19268 );
and \U$19248 ( \19270 , \19266 , \19269 );
and \U$19249 ( \19271 , \19259 , \19265 );
or \U$19250 ( \19272 , \19270 , \19271 );
buf \U$19251 ( \19273 , \19272 );
buf \U$19252 ( \19274 , \19273 );
xor \U$19253 ( \19275 , \19255 , \19274 );
buf \U$19254 ( \19276 , \19275 );
buf \U$19255 ( \19277 , \19276 );
xor \U$19256 ( \19278 , \18847 , \19277 );
xor \U$19257 ( \19279 , \19259 , \19265 );
xor \U$19258 ( \19280 , \19279 , \19269 );
buf \U$19259 ( \19281 , \19280 );
buf \U$19260 ( \19282 , \19281 );
xor \U$19261 ( \19283 , \18816 , \18820 );
and \U$19262 ( \19284 , \19283 , \18827 );
and \U$19263 ( \19285 , \18816 , \18820 );
or \U$19264 ( \19286 , \19284 , \19285 );
buf \U$19265 ( \19287 , \19286 );
buf \U$19266 ( \19288 , \19287 );
xor \U$19267 ( \19289 , \19282 , \19288 );
xor \U$19268 ( \19290 , \13137 , \14246 );
xor \U$19269 ( \19291 , \19290 , \15023 );
buf \U$19270 ( \19292 , \19291 );
buf \U$19271 ( \19293 , \19292 );
and \U$19272 ( \19294 , \19289 , \19293 );
and \U$19273 ( \19295 , \19282 , \19288 );
or \U$19274 ( \19296 , \19294 , \19295 );
buf \U$19275 ( \19297 , \19296 );
buf \U$19276 ( \19298 , \19297 );
xor \U$19277 ( \19299 , \19278 , \19298 );
buf \U$19278 ( \19300 , \19299 );
buf \U$19279 ( \19301 , \19300 );
xor \U$19280 ( \19302 , \18841 , \19301 );
buf \U$19281 ( \19303 , \19302 );
buf \U$19282 ( \19304 , \19303 );
xor \U$19283 ( \19305 , \19282 , \19288 );
xor \U$19284 ( \19306 , \19305 , \19293 );
buf \U$19285 ( \19307 , \19306 );
buf \U$19286 ( \19308 , \19307 );
not \U$19287 ( \19309 , \19308 );
buf \U$19288 ( \19310 , RIc0d8230_26);
buf \U$19289 ( \19311 , RIc0da918_109);
xor \U$19290 ( \19312 , \19310 , \19311 );
buf \U$19291 ( \19313 , \19312 );
buf \U$19292 ( \19314 , \19313 );
not \U$19293 ( \19315 , \19314 );
buf \U$19294 ( \19316 , \13419 );
not \U$19295 ( \19317 , \19316 );
or \U$19296 ( \19318 , \19315 , \19317 );
buf \U$19297 ( \19319 , \14216 );
buf \U$19298 ( \19320 , \18431 );
nand \U$19299 ( \19321 , \19319 , \19320 );
buf \U$19300 ( \19322 , \19321 );
buf \U$19301 ( \19323 , \19322 );
nand \U$19302 ( \19324 , \19318 , \19323 );
buf \U$19303 ( \19325 , \19324 );
buf \U$19304 ( \19326 , \19325 );
not \U$19305 ( \19327 , \19326 );
buf \U$19306 ( \19328 , RIc0d7e70_18);
buf \U$19307 ( \19329 , RIc0dacd8_117);
xor \U$19308 ( \19330 , \19328 , \19329 );
buf \U$19309 ( \19331 , \19330 );
buf \U$19310 ( \19332 , \19331 );
not \U$19311 ( \19333 , \19332 );
buf \U$19312 ( \19334 , \13684 );
not \U$19313 ( \19335 , \19334 );
or \U$19314 ( \19336 , \19333 , \19335 );
buf \U$19315 ( \19337 , \12937 );
buf \U$19316 ( \19338 , \18447 );
nand \U$19317 ( \19339 , \19337 , \19338 );
buf \U$19318 ( \19340 , \19339 );
buf \U$19319 ( \19341 , \19340 );
nand \U$19320 ( \19342 , \19336 , \19341 );
buf \U$19321 ( \19343 , \19342 );
buf \U$19322 ( \19344 , \19343 );
not \U$19323 ( \19345 , \19344 );
or \U$19324 ( \19346 , \19327 , \19345 );
buf \U$19325 ( \19347 , \19343 );
buf \U$19326 ( \19348 , \19325 );
or \U$19327 ( \19349 , \19347 , \19348 );
buf \U$19328 ( \19350 , RIc0d7ba0_12);
buf \U$19329 ( \19351 , RIc0dafa8_123);
xor \U$19330 ( \19352 , \19350 , \19351 );
buf \U$19331 ( \19353 , \19352 );
buf \U$19332 ( \19354 , \19353 );
not \U$19333 ( \19355 , \19354 );
buf \U$19334 ( \19356 , \14982 );
not \U$19335 ( \19357 , \19356 );
or \U$19336 ( \19358 , \19355 , \19357 );
buf \U$19337 ( \19359 , \16692 );
buf \U$19338 ( \19360 , \17113 );
nand \U$19339 ( \19361 , \19359 , \19360 );
buf \U$19340 ( \19362 , \19361 );
buf \U$19341 ( \19363 , \19362 );
nand \U$19342 ( \19364 , \19358 , \19363 );
buf \U$19343 ( \19365 , \19364 );
buf \U$19344 ( \19366 , \19365 );
nand \U$19345 ( \19367 , \19349 , \19366 );
buf \U$19346 ( \19368 , \19367 );
buf \U$19347 ( \19369 , \19368 );
nand \U$19348 ( \19370 , \19346 , \19369 );
buf \U$19349 ( \19371 , \19370 );
buf \U$19350 ( \19372 , \19371 );
not \U$19351 ( \19373 , \19372 );
buf \U$19352 ( \19374 , RIc0d8e60_52);
buf \U$19353 ( \19375 , RIc0d9ce8_83);
xor \U$19354 ( \19376 , \19374 , \19375 );
buf \U$19355 ( \19377 , \19376 );
buf \U$19356 ( \19378 , \19377 );
not \U$19357 ( \19379 , \19378 );
buf \U$19358 ( \19380 , \12254 );
not \U$19359 ( \19381 , \19380 );
or \U$19360 ( \19382 , \19379 , \19381 );
buf \U$19361 ( \19383 , \993 );
buf \U$19362 ( \19384 , \17179 );
nand \U$19363 ( \19385 , \19383 , \19384 );
buf \U$19364 ( \19386 , \19385 );
buf \U$19365 ( \19387 , \19386 );
nand \U$19366 ( \19388 , \19382 , \19387 );
buf \U$19367 ( \19389 , \19388 );
buf \U$19368 ( \19390 , \19389 );
xor \U$19369 ( \19391 , RIc0d9b08_79, RIc0d9040_56);
buf \U$19370 ( \19392 , \19391 );
not \U$19371 ( \19393 , \19392 );
buf \U$19372 ( \19394 , \14940 );
not \U$19373 ( \19395 , \19394 );
or \U$19374 ( \19396 , \19393 , \19395 );
buf \U$19375 ( \19397 , \1025 );
buf \U$19376 ( \19398 , \17573 );
nand \U$19377 ( \19399 , \19397 , \19398 );
buf \U$19378 ( \19400 , \19399 );
buf \U$19379 ( \19401 , \19400 );
nand \U$19380 ( \19402 , \19396 , \19401 );
buf \U$19381 ( \19403 , \19402 );
buf \U$19382 ( \19404 , \19403 );
xor \U$19383 ( \19405 , \19390 , \19404 );
buf \U$19384 ( \19406 , RIc0d8320_28);
buf \U$19385 ( \19407 , RIc0da828_107);
xor \U$19386 ( \19408 , \19406 , \19407 );
buf \U$19387 ( \19409 , \19408 );
buf \U$19388 ( \19410 , \19409 );
not \U$19389 ( \19411 , \19410 );
buf \U$19390 ( \19412 , \12331 );
not \U$19391 ( \19413 , \19412 );
buf \U$19392 ( \19414 , \19413 );
buf \U$19393 ( \19415 , \19414 );
not \U$19394 ( \19416 , \19415 );
or \U$19395 ( \19417 , \19411 , \19416 );
buf \U$19396 ( \19418 , \12342 );
buf \U$19397 ( \19419 , \17590 );
nand \U$19398 ( \19420 , \19418 , \19419 );
buf \U$19399 ( \19421 , \19420 );
buf \U$19400 ( \19422 , \19421 );
nand \U$19401 ( \19423 , \19417 , \19422 );
buf \U$19402 ( \19424 , \19423 );
buf \U$19403 ( \19425 , \19424 );
and \U$19404 ( \19426 , \19405 , \19425 );
and \U$19405 ( \19427 , \19390 , \19404 );
or \U$19406 ( \19428 , \19426 , \19427 );
buf \U$19407 ( \19429 , \19428 );
buf \U$19408 ( \19430 , \19429 );
not \U$19409 ( \19431 , \19430 );
or \U$19410 ( \19432 , \19373 , \19431 );
buf \U$19411 ( \19433 , \19429 );
buf \U$19412 ( \19434 , \19371 );
or \U$19413 ( \19435 , \19433 , \19434 );
buf \U$19414 ( \19436 , RIc0d8c80_48);
buf \U$19415 ( \19437 , RIc0d9ec8_87);
xor \U$19416 ( \19438 , \19436 , \19437 );
buf \U$19417 ( \19439 , \19438 );
buf \U$19418 ( \19440 , \19439 );
not \U$19419 ( \19441 , \19440 );
buf \U$19420 ( \19442 , \14325 );
not \U$19421 ( \19443 , \19442 );
or \U$19422 ( \19444 , \19441 , \19443 );
buf \U$19423 ( \19445 , \816 );
buf \U$19424 ( \19446 , \17066 );
nand \U$19425 ( \19447 , \19445 , \19446 );
buf \U$19426 ( \19448 , \19447 );
buf \U$19427 ( \19449 , \19448 );
nand \U$19428 ( \19450 , \19444 , \19449 );
buf \U$19429 ( \19451 , \19450 );
buf \U$19430 ( \19452 , \19451 );
not \U$19431 ( \19453 , \19452 );
buf \U$19432 ( \19454 , \19453 );
buf \U$19433 ( \19455 , \19454 );
not \U$19434 ( \19456 , \19455 );
buf \U$19435 ( \19457 , RIc0d89b0_42);
buf \U$19436 ( \19458 , RIc0da198_93);
xor \U$19437 ( \19459 , \19457 , \19458 );
buf \U$19438 ( \19460 , \19459 );
buf \U$19439 ( \19461 , \19460 );
not \U$19440 ( \19462 , \19461 );
buf \U$19441 ( \19463 , \15995 );
not \U$19442 ( \19464 , \19463 );
or \U$19443 ( \19465 , \19462 , \19464 );
buf \U$19444 ( \19466 , \481 );
buf \U$19445 ( \19467 , \17613 );
nand \U$19446 ( \19468 , \19466 , \19467 );
buf \U$19447 ( \19469 , \19468 );
buf \U$19448 ( \19470 , \19469 );
nand \U$19449 ( \19471 , \19465 , \19470 );
buf \U$19450 ( \19472 , \19471 );
buf \U$19451 ( \19473 , \19472 );
not \U$19452 ( \19474 , \19473 );
buf \U$19453 ( \19475 , \19474 );
buf \U$19454 ( \19476 , \19475 );
not \U$19455 ( \19477 , \19476 );
or \U$19456 ( \19478 , \19456 , \19477 );
buf \U$19457 ( \19479 , RIc0d7c90_14);
buf \U$19458 ( \19480 , RIc0daeb8_121);
xor \U$19459 ( \19481 , \19479 , \19480 );
buf \U$19460 ( \19482 , \19481 );
buf \U$19461 ( \19483 , \19482 );
not \U$19462 ( \19484 , \19483 );
buf \U$19463 ( \19485 , \12968 );
not \U$19464 ( \19486 , \19485 );
buf \U$19465 ( \19487 , \19486 );
buf \U$19466 ( \19488 , \19487 );
not \U$19467 ( \19489 , \19488 );
or \U$19468 ( \19490 , \19484 , \19489 );
buf \U$19469 ( \19491 , \16386 );
buf \U$19470 ( \19492 , \17084 );
nand \U$19471 ( \19493 , \19491 , \19492 );
buf \U$19472 ( \19494 , \19493 );
buf \U$19473 ( \19495 , \19494 );
nand \U$19474 ( \19496 , \19490 , \19495 );
buf \U$19475 ( \19497 , \19496 );
buf \U$19476 ( \19498 , \19497 );
nand \U$19477 ( \19499 , \19478 , \19498 );
buf \U$19478 ( \19500 , \19499 );
buf \U$19479 ( \19501 , \19500 );
buf \U$19480 ( \19502 , \19472 );
buf \U$19481 ( \19503 , \19451 );
nand \U$19482 ( \19504 , \19502 , \19503 );
buf \U$19483 ( \19505 , \19504 );
buf \U$19484 ( \19506 , \19505 );
nand \U$19485 ( \19507 , \19501 , \19506 );
buf \U$19486 ( \19508 , \19507 );
buf \U$19487 ( \19509 , \19508 );
nand \U$19488 ( \19510 , \19435 , \19509 );
buf \U$19489 ( \19511 , \19510 );
buf \U$19490 ( \19512 , \19511 );
nand \U$19491 ( \19513 , \19432 , \19512 );
buf \U$19492 ( \19514 , \19513 );
buf \U$19493 ( \19515 , \19514 );
not \U$19494 ( \19516 , \19515 );
buf \U$19495 ( \19517 , \19516 );
buf \U$19496 ( \19518 , \19517 );
not \U$19497 ( \19519 , \19518 );
buf \U$19498 ( \19520 , RIc0d7ab0_10);
buf \U$19499 ( \19521 , RIc0db098_125);
xor \U$19500 ( \19522 , \19520 , \19521 );
buf \U$19501 ( \19523 , \19522 );
buf \U$19502 ( \19524 , \19523 );
not \U$19503 ( \19525 , \19524 );
buf \U$19504 ( \19526 , \16914 );
not \U$19505 ( \19527 , \19526 );
or \U$19506 ( \19528 , \19525 , \19527 );
buf \U$19507 ( \19529 , \15793 );
buf \U$19508 ( \19530 , \16908 );
nand \U$19509 ( \19531 , \19529 , \19530 );
buf \U$19510 ( \19532 , \19531 );
buf \U$19511 ( \19533 , \19532 );
nand \U$19512 ( \19534 , \19528 , \19533 );
buf \U$19513 ( \19535 , \19534 );
buf \U$19514 ( \19536 , \19535 );
buf \U$19515 ( \19537 , RIc0d8f50_54);
buf \U$19516 ( \19538 , RIc0d9bf8_81);
xor \U$19517 ( \19539 , \19537 , \19538 );
buf \U$19518 ( \19540 , \19539 );
buf \U$19519 ( \19541 , \19540 );
not \U$19520 ( \19542 , \19541 );
not \U$19521 ( \19543 , \1056 );
nor \U$19522 ( \19544 , \19543 , \1077 );
buf \U$19523 ( \19545 , \19544 );
not \U$19524 ( \19546 , \19545 );
or \U$19525 ( \19547 , \19542 , \19546 );
buf \U$19526 ( \19548 , \1078 );
buf \U$19527 ( \19549 , \17136 );
nand \U$19528 ( \19550 , \19548 , \19549 );
buf \U$19529 ( \19551 , \19550 );
buf \U$19530 ( \19552 , \19551 );
nand \U$19531 ( \19553 , \19547 , \19552 );
buf \U$19532 ( \19554 , \19553 );
buf \U$19533 ( \19555 , \19554 );
xor \U$19534 ( \19556 , \19536 , \19555 );
buf \U$19535 ( \19557 , RIc0d7d80_16);
buf \U$19536 ( \19558 , RIc0dadc8_119);
xor \U$19537 ( \19559 , \19557 , \19558 );
buf \U$19538 ( \19560 , \19559 );
buf \U$19539 ( \19561 , \19560 );
not \U$19540 ( \19562 , \19561 );
buf \U$19541 ( \19563 , \13181 );
not \U$19542 ( \19564 , \19563 );
or \U$19543 ( \19565 , \19562 , \19564 );
buf \U$19544 ( \19566 , \13005 );
buf \U$19545 ( \19567 , \17157 );
nand \U$19546 ( \19568 , \19566 , \19567 );
buf \U$19547 ( \19569 , \19568 );
buf \U$19548 ( \19570 , \19569 );
nand \U$19549 ( \19571 , \19565 , \19570 );
buf \U$19550 ( \19572 , \19571 );
buf \U$19551 ( \19573 , \19572 );
and \U$19552 ( \19574 , \19556 , \19573 );
and \U$19553 ( \19575 , \19536 , \19555 );
or \U$19554 ( \19576 , \19574 , \19575 );
buf \U$19555 ( \19577 , \19576 );
buf \U$19556 ( \19578 , RIc0d7f60_20);
buf \U$19557 ( \19579 , RIc0dabe8_115);
xor \U$19558 ( \19580 , \19578 , \19579 );
buf \U$19559 ( \19581 , \19580 );
buf \U$19560 ( \19582 , \19581 );
not \U$19561 ( \19583 , \19582 );
buf \U$19562 ( \19584 , \12299 );
not \U$19563 ( \19585 , \19584 );
or \U$19564 ( \19586 , \19583 , \19585 );
buf \U$19565 ( \19587 , \12303 );
buf \U$19566 ( \19588 , \17039 );
nand \U$19567 ( \19589 , \19587 , \19588 );
buf \U$19568 ( \19590 , \19589 );
buf \U$19569 ( \19591 , \19590 );
nand \U$19570 ( \19592 , \19586 , \19591 );
buf \U$19571 ( \19593 , \19592 );
buf \U$19572 ( \19594 , \19593 );
not \U$19573 ( \19595 , \19594 );
buf \U$19574 ( \19596 , RIc0d8aa0_44);
buf \U$19575 ( \19597 , RIc0da0a8_91);
xor \U$19576 ( \19598 , \19596 , \19597 );
buf \U$19577 ( \19599 , \19598 );
buf \U$19578 ( \19600 , \19599 );
not \U$19579 ( \19601 , \19600 );
buf \U$19580 ( \19602 , \16402 );
not \U$19581 ( \19603 , \19602 );
or \U$19582 ( \19604 , \19601 , \19603 );
buf \U$19583 ( \19605 , \533 );
buf \U$19584 ( \19606 , \16870 );
nand \U$19585 ( \19607 , \19605 , \19606 );
buf \U$19586 ( \19608 , \19607 );
buf \U$19587 ( \19609 , \19608 );
nand \U$19588 ( \19610 , \19604 , \19609 );
buf \U$19589 ( \19611 , \19610 );
buf \U$19590 ( \19612 , \19611 );
not \U$19591 ( \19613 , \19612 );
or \U$19592 ( \19614 , \19595 , \19613 );
buf \U$19593 ( \19615 , \19593 );
not \U$19594 ( \19616 , \19615 );
buf \U$19595 ( \19617 , \19616 );
buf \U$19596 ( \19618 , \19617 );
not \U$19597 ( \19619 , \19618 );
buf \U$19598 ( \19620 , \19611 );
not \U$19599 ( \19621 , \19620 );
buf \U$19600 ( \19622 , \19621 );
buf \U$19601 ( \19623 , \19622 );
not \U$19602 ( \19624 , \19623 );
or \U$19603 ( \19625 , \19619 , \19624 );
buf \U$19604 ( \19626 , RIc0d8410_30);
buf \U$19605 ( \19627 , RIc0da738_105);
xor \U$19606 ( \19628 , \19626 , \19627 );
buf \U$19607 ( \19629 , \19628 );
buf \U$19608 ( \19630 , \19629 );
not \U$19609 ( \19631 , \19630 );
buf \U$19610 ( \19632 , \12736 );
not \U$19611 ( \19633 , \19632 );
or \U$19612 ( \19634 , \19631 , \19633 );
buf \U$19613 ( \19635 , \12744 );
buf \U$19614 ( \19636 , \16886 );
nand \U$19615 ( \19637 , \19635 , \19636 );
buf \U$19616 ( \19638 , \19637 );
buf \U$19617 ( \19639 , \19638 );
nand \U$19618 ( \19640 , \19634 , \19639 );
buf \U$19619 ( \19641 , \19640 );
buf \U$19620 ( \19642 , \19641 );
nand \U$19621 ( \19643 , \19625 , \19642 );
buf \U$19622 ( \19644 , \19643 );
buf \U$19623 ( \19645 , \19644 );
nand \U$19624 ( \19646 , \19614 , \19645 );
buf \U$19625 ( \19647 , \19646 );
xor \U$19626 ( \19648 , \19577 , \19647 );
buf \U$19627 ( \19649 , RIc0d8d70_50);
buf \U$19628 ( \19650 , RIc0d9dd8_85);
xor \U$19629 ( \19651 , \19649 , \19650 );
buf \U$19630 ( \19652 , \19651 );
buf \U$19631 ( \19653 , \19652 );
not \U$19632 ( \19654 , \19653 );
buf \U$19633 ( \19655 , \5304 );
not \U$19634 ( \19656 , \19655 );
or \U$19635 ( \19657 , \19654 , \19656 );
buf \U$19636 ( \19658 , \17017 );
not \U$19637 ( \19659 , \19658 );
buf \U$19638 ( \19660 , \921 );
nand \U$19639 ( \19661 , \19659 , \19660 );
buf \U$19640 ( \19662 , \19661 );
buf \U$19641 ( \19663 , \19662 );
nand \U$19642 ( \19664 , \19657 , \19663 );
buf \U$19643 ( \19665 , \19664 );
buf \U$19644 ( \19666 , \19665 );
not \U$19645 ( \19667 , \19666 );
buf \U$19646 ( \19668 , \19667 );
buf \U$19647 ( \19669 , \19668 );
not \U$19648 ( \19670 , \19669 );
xor \U$19649 ( \19671 , RIc0daaf8_113, RIc0d8050_22);
buf \U$19650 ( \19672 , \19671 );
not \U$19651 ( \19673 , \19672 );
buf \U$19652 ( \19674 , \14891 );
not \U$19653 ( \19675 , \19674 );
or \U$19654 ( \19676 , \19673 , \19675 );
buf \U$19655 ( \19677 , \12410 );
buf \U$19656 ( \19678 , \16984 );
nand \U$19657 ( \19679 , \19677 , \19678 );
buf \U$19658 ( \19680 , \19679 );
buf \U$19659 ( \19681 , \19680 );
nand \U$19660 ( \19682 , \19676 , \19681 );
buf \U$19661 ( \19683 , \19682 );
buf \U$19662 ( \19684 , \19683 );
not \U$19663 ( \19685 , \19684 );
buf \U$19664 ( \19686 , \19685 );
buf \U$19665 ( \19687 , \19686 );
not \U$19666 ( \19688 , \19687 );
or \U$19667 ( \19689 , \19670 , \19688 );
xor \U$19668 ( \19690 , RIc0da468_99, RIc0d86e0_36);
buf \U$19669 ( \19691 , \19690 );
not \U$19670 ( \19692 , \19691 );
buf \U$19671 ( \19693 , \2207 );
not \U$19672 ( \19694 , \19693 );
buf \U$19673 ( \19695 , \19694 );
buf \U$19674 ( \19696 , \19695 );
not \U$19675 ( \19697 , \19696 );
or \U$19676 ( \19698 , \19692 , \19697 );
buf \U$19677 ( \19699 , \16750 );
buf \U$19678 ( \19700 , \17021 );
nand \U$19679 ( \19701 , \19699 , \19700 );
buf \U$19680 ( \19702 , \19701 );
buf \U$19681 ( \19703 , \19702 );
nand \U$19682 ( \19704 , \19698 , \19703 );
buf \U$19683 ( \19705 , \19704 );
buf \U$19684 ( \19706 , \19705 );
nand \U$19685 ( \19707 , \19689 , \19706 );
buf \U$19686 ( \19708 , \19707 );
buf \U$19687 ( \19709 , \19708 );
buf \U$19688 ( \19710 , \19683 );
buf \U$19689 ( \19711 , \19665 );
nand \U$19690 ( \19712 , \19710 , \19711 );
buf \U$19691 ( \19713 , \19712 );
buf \U$19692 ( \19714 , \19713 );
nand \U$19693 ( \19715 , \19709 , \19714 );
buf \U$19694 ( \19716 , \19715 );
and \U$19695 ( \19717 , \19648 , \19716 );
and \U$19696 ( \19718 , \19577 , \19647 );
or \U$19697 ( \19719 , \19717 , \19718 );
buf \U$19698 ( \19720 , \19719 );
not \U$19699 ( \19721 , \19720 );
buf \U$19700 ( \19722 , \19721 );
buf \U$19701 ( \19723 , \19722 );
not \U$19702 ( \19724 , \19723 );
or \U$19703 ( \19725 , \19519 , \19724 );
xor \U$19704 ( \19726 , \17259 , \17131 );
xor \U$19705 ( \19727 , \19726 , \17197 );
buf \U$19706 ( \19728 , \19727 );
nand \U$19707 ( \19729 , \19725 , \19728 );
buf \U$19708 ( \19730 , \19729 );
buf \U$19709 ( \19731 , \19730 );
buf \U$19710 ( \19732 , \19719 );
buf \U$19711 ( \19733 , \19514 );
nand \U$19712 ( \19734 , \19732 , \19733 );
buf \U$19713 ( \19735 , \19734 );
buf \U$19714 ( \19736 , \19735 );
nand \U$19715 ( \19737 , \19731 , \19736 );
buf \U$19716 ( \19738 , \19737 );
buf \U$19717 ( \19739 , \19738 );
buf \U$19718 ( \19740 , \17061 );
not \U$19719 ( \19741 , \19740 );
buf \U$19720 ( \19742 , \17279 );
not \U$19721 ( \19743 , \19742 );
or \U$19722 ( \19744 , \19741 , \19743 );
buf \U$19723 ( \19745 , \17275 );
buf \U$19724 ( \19746 , \17270 );
nand \U$19725 ( \19747 , \19745 , \19746 );
buf \U$19726 ( \19748 , \19747 );
buf \U$19727 ( \19749 , \19748 );
nand \U$19728 ( \19750 , \19744 , \19749 );
buf \U$19729 ( \19751 , \19750 );
buf \U$19730 ( \19752 , \19751 );
buf \U$19731 ( \19753 , \17284 );
xor \U$19732 ( \19754 , \19752 , \19753 );
buf \U$19733 ( \19755 , \19754 );
buf \U$19734 ( \19756 , \19755 );
xor \U$19735 ( \19757 , \19739 , \19756 );
xor \U$19736 ( \19758 , \16935 , \17005 );
xor \U$19737 ( \19759 , \19758 , \17057 );
buf \U$19738 ( \19760 , \19759 );
buf \U$19739 ( \19761 , \19760 );
buf \U$19740 ( \19762 , \18520 );
buf \U$19741 ( \19763 , \18478 );
xor \U$19742 ( \19764 , \19762 , \19763 );
buf \U$19743 ( \19765 , \18425 );
xor \U$19744 ( \19766 , \19764 , \19765 );
buf \U$19745 ( \19767 , \19766 );
buf \U$19746 ( \19768 , \19767 );
xor \U$19747 ( \19769 , \19761 , \19768 );
xor \U$19748 ( \19770 , \18443 , \18459 );
xor \U$19749 ( \19771 , \19770 , \18475 );
buf \U$19750 ( \19772 , \19771 );
buf \U$19751 ( \19773 , \16972 );
not \U$19752 ( \19774 , \19773 );
buf \U$19753 ( \19775 , \16981 );
not \U$19754 ( \19776 , \19775 );
or \U$19755 ( \19777 , \19774 , \19776 );
buf \U$19756 ( \19778 , \16952 );
buf \U$19757 ( \19779 , \16977 );
nand \U$19758 ( \19780 , \19778 , \19779 );
buf \U$19759 ( \19781 , \19780 );
buf \U$19760 ( \19782 , \19781 );
nand \U$19761 ( \19783 , \19777 , \19782 );
buf \U$19762 ( \19784 , \19783 );
buf \U$19763 ( \19785 , \19784 );
buf \U$19764 ( \19786 , \17002 );
xnor \U$19765 ( \19787 , \19785 , \19786 );
buf \U$19766 ( \19788 , \19787 );
buf \U$19767 ( \19789 , \19788 );
not \U$19768 ( \19790 , \19789 );
buf \U$19769 ( \19791 , \19790 );
buf \U$19770 ( \19792 , \19791 );
or \U$19771 ( \19793 , \19772 , \19792 );
xor \U$19772 ( \19794 , \18489 , \18502 );
xor \U$19773 ( \19795 , \19794 , \18516 );
buf \U$19774 ( \19796 , \19795 );
buf \U$19775 ( \19797 , \19796 );
nand \U$19776 ( \19798 , \19793 , \19797 );
buf \U$19777 ( \19799 , \19798 );
buf \U$19778 ( \19800 , \19799 );
buf \U$19779 ( \19801 , \19771 );
buf \U$19780 ( \19802 , \19791 );
nand \U$19781 ( \19803 , \19801 , \19802 );
buf \U$19782 ( \19804 , \19803 );
buf \U$19783 ( \19805 , \19804 );
nand \U$19784 ( \19806 , \19800 , \19805 );
buf \U$19785 ( \19807 , \19806 );
buf \U$19786 ( \19808 , \19807 );
and \U$19787 ( \19809 , \19769 , \19808 );
and \U$19788 ( \19810 , \19761 , \19768 );
or \U$19789 ( \19811 , \19809 , \19810 );
buf \U$19790 ( \19812 , \19811 );
buf \U$19791 ( \19813 , \19812 );
and \U$19792 ( \19814 , \19757 , \19813 );
and \U$19793 ( \19815 , \19739 , \19756 );
or \U$19794 ( \19816 , \19814 , \19815 );
buf \U$19795 ( \19817 , \19816 );
buf \U$19796 ( \19818 , \19817 );
buf \U$19797 ( \19819 , \18546 );
buf \U$19798 ( \19820 , \18526 );
xor \U$19799 ( \19821 , \19819 , \19820 );
buf \U$19800 ( \19822 , \18551 );
xnor \U$19801 ( \19823 , \19821 , \19822 );
buf \U$19802 ( \19824 , \19823 );
buf \U$19803 ( \19825 , \19824 );
not \U$19804 ( \19826 , \19825 );
buf \U$19805 ( \19827 , \17429 );
not \U$19806 ( \19828 , \19827 );
buf \U$19807 ( \19829 , \17298 );
not \U$19808 ( \19830 , \19829 );
or \U$19809 ( \19831 , \19828 , \19830 );
buf \U$19810 ( \19832 , \17298 );
buf \U$19811 ( \19833 , \17429 );
or \U$19812 ( \19834 , \19832 , \19833 );
nand \U$19813 ( \19835 , \19831 , \19834 );
buf \U$19814 ( \19836 , \19835 );
buf \U$19815 ( \19837 , \19836 );
buf \U$19816 ( \19838 , \17504 );
not \U$19817 ( \19839 , \19838 );
buf \U$19818 ( \19840 , \19839 );
buf \U$19819 ( \19841 , \19840 );
and \U$19820 ( \19842 , \19837 , \19841 );
not \U$19821 ( \19843 , \19837 );
buf \U$19822 ( \19844 , \17504 );
and \U$19823 ( \19845 , \19843 , \19844 );
nor \U$19824 ( \19846 , \19842 , \19845 );
buf \U$19825 ( \19847 , \19846 );
buf \U$19826 ( \19848 , \19847 );
not \U$19827 ( \19849 , \19848 );
or \U$19828 ( \19850 , \19826 , \19849 );
xor \U$19829 ( \19851 , \17552 , \17571 );
xor \U$19830 ( \19852 , \19851 , \17651 );
buf \U$19831 ( \19853 , \19852 );
buf \U$19832 ( \19854 , \19853 );
nand \U$19833 ( \19855 , \19850 , \19854 );
buf \U$19834 ( \19856 , \19855 );
buf \U$19835 ( \19857 , \19856 );
buf \U$19836 ( \19858 , \19847 );
not \U$19837 ( \19859 , \19858 );
buf \U$19838 ( \19860 , \19824 );
not \U$19839 ( \19861 , \19860 );
buf \U$19840 ( \19862 , \19861 );
buf \U$19841 ( \19863 , \19862 );
nand \U$19842 ( \19864 , \19859 , \19863 );
buf \U$19843 ( \19865 , \19864 );
buf \U$19844 ( \19866 , \19865 );
nand \U$19845 ( \19867 , \19857 , \19866 );
buf \U$19846 ( \19868 , \19867 );
buf \U$19847 ( \19869 , \19868 );
or \U$19848 ( \19870 , \19818 , \19869 );
xor \U$19849 ( \19871 , \17287 , \17291 );
xor \U$19850 ( \19872 , \19871 , \17511 );
buf \U$19851 ( \19873 , \19872 );
buf \U$19852 ( \19874 , \19873 );
nand \U$19853 ( \19875 , \19870 , \19874 );
buf \U$19854 ( \19876 , \19875 );
buf \U$19855 ( \19877 , \19876 );
buf \U$19856 ( \19878 , \19817 );
buf \U$19857 ( \19879 , \19868 );
nand \U$19858 ( \19880 , \19878 , \19879 );
buf \U$19859 ( \19881 , \19880 );
buf \U$19860 ( \19882 , \19881 );
nand \U$19861 ( \19883 , \19877 , \19882 );
buf \U$19862 ( \19884 , \19883 );
buf \U$19863 ( \19885 , \19884 );
not \U$19864 ( \19886 , \19885 );
buf \U$19865 ( \19887 , \19886 );
buf \U$19866 ( \19888 , \19887 );
not \U$19867 ( \19889 , \19888 );
xor \U$19868 ( \19890 , \17516 , \17801 );
xor \U$19869 ( \19891 , \19890 , \17834 );
buf \U$19870 ( \19892 , \19891 );
buf \U$19871 ( \19893 , \19892 );
not \U$19872 ( \19894 , \19893 );
buf \U$19873 ( \19895 , \19894 );
buf \U$19874 ( \19896 , \19895 );
not \U$19875 ( \19897 , \19896 );
or \U$19876 ( \19898 , \19889 , \19897 );
xor \U$19877 ( \19899 , \17962 , \17984 );
xor \U$19878 ( \19900 , \19899 , \18253 );
buf \U$19879 ( \19901 , \19900 );
buf \U$19880 ( \19902 , \19901 );
buf \U$19881 ( \19903 , \17549 );
not \U$19882 ( \19904 , \19903 );
buf \U$19883 ( \19905 , \17523 );
not \U$19884 ( \19906 , \19905 );
or \U$19885 ( \19907 , \19904 , \19906 );
buf \U$19886 ( \19908 , \17549 );
not \U$19887 ( \19909 , \19908 );
buf \U$19888 ( \19910 , \17526 );
nand \U$19889 ( \19911 , \19909 , \19910 );
buf \U$19890 ( \19912 , \19911 );
buf \U$19891 ( \19913 , \19912 );
nand \U$19892 ( \19914 , \19907 , \19913 );
buf \U$19893 ( \19915 , \19914 );
buf \U$19894 ( \19916 , \19915 );
buf \U$19895 ( \19917 , \17533 );
and \U$19896 ( \19918 , \19916 , \19917 );
not \U$19897 ( \19919 , \19916 );
buf \U$19898 ( \19920 , \17536 );
and \U$19899 ( \19921 , \19919 , \19920 );
nor \U$19900 ( \19922 , \19918 , \19921 );
buf \U$19901 ( \19923 , \19922 );
buf \U$19902 ( \19924 , \19923 );
not \U$19903 ( \19925 , \19924 );
buf \U$19904 ( \19926 , \19925 );
not \U$19905 ( \19927 , \19926 );
xor \U$19906 ( \19928 , \17220 , \17237 );
xor \U$19907 ( \19929 , \19928 , \17255 );
buf \U$19908 ( \19930 , \19929 );
buf \U$19909 ( \19931 , \19930 );
buf \U$19910 ( \19932 , RIc0d85f0_34);
buf \U$19911 ( \19933 , RIc0da558_101);
xor \U$19912 ( \19934 , \19932 , \19933 );
buf \U$19913 ( \19935 , \19934 );
buf \U$19914 ( \19936 , \19935 );
not \U$19915 ( \19937 , \19936 );
buf \U$19916 ( \19938 , \4042 );
not \U$19917 ( \19939 , \19938 );
or \U$19918 ( \19940 , \19937 , \19939 );
buf \U$19919 ( \19941 , \4049 );
buf \U$19920 ( \19942 , \17242 );
nand \U$19921 ( \19943 , \19941 , \19942 );
buf \U$19922 ( \19944 , \19943 );
buf \U$19923 ( \19945 , \19944 );
nand \U$19924 ( \19946 , \19940 , \19945 );
buf \U$19925 ( \19947 , \19946 );
buf \U$19926 ( \19948 , \19947 );
buf \U$19927 ( \19949 , \14713 );
buf \U$19928 ( \19950 , RIc0d88c0_40);
buf \U$19929 ( \19951 , RIc0da288_95);
xnor \U$19930 ( \19952 , \19950 , \19951 );
buf \U$19931 ( \19953 , \19952 );
buf \U$19932 ( \19954 , \19953 );
or \U$19933 ( \19955 , \19949 , \19954 );
buf \U$19934 ( \19956 , \344 );
buf \U$19935 ( \19957 , \18465 );
nand \U$19936 ( \19958 , \19956 , \19957 );
buf \U$19937 ( \19959 , \19958 );
buf \U$19938 ( \19960 , \19959 );
nand \U$19939 ( \19961 , \19955 , \19960 );
buf \U$19940 ( \19962 , \19961 );
buf \U$19941 ( \19963 , \19962 );
xor \U$19942 ( \19964 , \19948 , \19963 );
buf \U$19943 ( \19965 , RIc0daa08_111);
buf \U$19944 ( \19966 , RIc0d8140_24);
xor \U$19945 ( \19967 , \19965 , \19966 );
buf \U$19946 ( \19968 , \19967 );
buf \U$19947 ( \19969 , \19968 );
not \U$19948 ( \19970 , \19969 );
buf \U$19949 ( \19971 , \14346 );
not \U$19950 ( \19972 , \19971 );
or \U$19951 ( \19973 , \19970 , \19972 );
buf \U$19952 ( \19974 , \14353 );
buf \U$19953 ( \19975 , \17224 );
nand \U$19954 ( \19976 , \19974 , \19975 );
buf \U$19955 ( \19977 , \19976 );
buf \U$19956 ( \19978 , \19977 );
nand \U$19957 ( \19979 , \19973 , \19978 );
buf \U$19958 ( \19980 , \19979 );
buf \U$19959 ( \19981 , \19980 );
and \U$19960 ( \19982 , \19964 , \19981 );
and \U$19961 ( \19983 , \19948 , \19963 );
or \U$19962 ( \19984 , \19982 , \19983 );
buf \U$19963 ( \19985 , \19984 );
buf \U$19964 ( \19986 , \19985 );
xor \U$19965 ( \19987 , \19931 , \19986 );
xnor \U$19966 ( \19988 , \18423 , \18402 );
buf \U$19967 ( \19989 , \19988 );
buf \U$19968 ( \19990 , \18384 );
and \U$19969 ( \19991 , \19989 , \19990 );
not \U$19970 ( \19992 , \19989 );
buf \U$19971 ( \19993 , \18406 );
and \U$19972 ( \19994 , \19992 , \19993 );
nor \U$19973 ( \19995 , \19991 , \19994 );
buf \U$19974 ( \19996 , \19995 );
buf \U$19975 ( \19997 , \19996 );
and \U$19976 ( \19998 , \19987 , \19997 );
and \U$19977 ( \19999 , \19931 , \19986 );
or \U$19978 ( \20000 , \19998 , \19999 );
buf \U$19979 ( \20001 , \20000 );
not \U$19980 ( \20002 , \20001 );
or \U$19981 ( \20003 , \19927 , \20002 );
buf \U$19982 ( \20004 , \20001 );
not \U$19983 ( \20005 , \20004 );
buf \U$19984 ( \20006 , \20005 );
not \U$19985 ( \20007 , \20006 );
not \U$19986 ( \20008 , \19923 );
or \U$19987 ( \20009 , \20007 , \20008 );
xor \U$19988 ( \20010 , \17020 , \17034 );
xor \U$19989 ( \20011 , \20010 , \17052 );
buf \U$19990 ( \20012 , \20011 );
buf \U$19991 ( \20013 , \20012 );
not \U$19992 ( \20014 , \20013 );
xor \U$19993 ( \20015 , \17605 , \17628 );
xnor \U$19994 ( \20016 , \20015 , \17585 );
buf \U$19995 ( \20017 , \20016 );
not \U$19996 ( \20018 , \20017 );
or \U$19997 ( \20019 , \20014 , \20018 );
buf \U$19998 ( \20020 , \20016 );
buf \U$19999 ( \20021 , \20012 );
or \U$20000 ( \20022 , \20020 , \20021 );
buf \U$20001 ( \20023 , \17125 );
buf \U$20002 ( \20024 , \17103 );
and \U$20003 ( \20025 , \20023 , \20024 );
not \U$20004 ( \20026 , \20023 );
buf \U$20005 ( \20027 , \17103 );
not \U$20006 ( \20028 , \20027 );
buf \U$20007 ( \20029 , \20028 );
buf \U$20008 ( \20030 , \20029 );
and \U$20009 ( \20031 , \20026 , \20030 );
nor \U$20010 ( \20032 , \20025 , \20031 );
buf \U$20011 ( \20033 , \20032 );
buf \U$20012 ( \20034 , \20033 );
buf \U$20013 ( \20035 , \17078 );
not \U$20014 ( \20036 , \20035 );
buf \U$20015 ( \20037 , \20036 );
buf \U$20016 ( \20038 , \20037 );
and \U$20017 ( \20039 , \20034 , \20038 );
not \U$20018 ( \20040 , \20034 );
buf \U$20019 ( \20041 , \17078 );
and \U$20020 ( \20042 , \20040 , \20041 );
nor \U$20021 ( \20043 , \20039 , \20042 );
buf \U$20022 ( \20044 , \20043 );
buf \U$20023 ( \20045 , \20044 );
not \U$20024 ( \20046 , \20045 );
buf \U$20025 ( \20047 , \20046 );
buf \U$20026 ( \20048 , \20047 );
nand \U$20027 ( \20049 , \20022 , \20048 );
buf \U$20028 ( \20050 , \20049 );
buf \U$20029 ( \20051 , \20050 );
nand \U$20030 ( \20052 , \20019 , \20051 );
buf \U$20031 ( \20053 , \20052 );
nand \U$20032 ( \20054 , \20009 , \20053 );
nand \U$20033 ( \20055 , \20003 , \20054 );
buf \U$20034 ( \20056 , \20055 );
xor \U$20035 ( \20057 , \19902 , \20056 );
xor \U$20036 ( \20058 , \17638 , \17642 );
xor \U$20037 ( \20059 , \20058 , \17646 );
buf \U$20038 ( \20060 , \20059 );
buf \U$20039 ( \20061 , \20060 );
buf \U$20040 ( \20062 , \17470 );
not \U$20041 ( \20063 , \20062 );
buf \U$20042 ( \20064 , \17498 );
not \U$20043 ( \20065 , \20064 );
or \U$20044 ( \20066 , \20063 , \20065 );
buf \U$20045 ( \20067 , \17470 );
buf \U$20046 ( \20068 , \17498 );
or \U$20047 ( \20069 , \20067 , \20068 );
nand \U$20048 ( \20070 , \20066 , \20069 );
buf \U$20049 ( \20071 , \20070 );
buf \U$20050 ( \20072 , \20071 );
buf \U$20051 ( \20073 , \17447 );
and \U$20052 ( \20074 , \20072 , \20073 );
not \U$20053 ( \20075 , \20072 );
buf \U$20054 ( \20076 , \17444 );
and \U$20055 ( \20077 , \20075 , \20076 );
nor \U$20056 ( \20078 , \20074 , \20077 );
buf \U$20057 ( \20079 , \20078 );
buf \U$20058 ( \20080 , \20079 );
xor \U$20059 ( \20081 , \20061 , \20080 );
xor \U$20060 ( \20082 , \17191 , \17169 );
xor \U$20061 ( \20083 , \20082 , \17151 );
buf \U$20062 ( \20084 , \20083 );
xor \U$20063 ( \20085 , \16898 , \16883 );
xor \U$20064 ( \20086 , \20085 , \16928 );
buf \U$20065 ( \20087 , \20086 );
xor \U$20066 ( \20088 , \20084 , \20087 );
buf \U$20067 ( \20089 , RIc0d7d08_15);
buf \U$20068 ( \20090 , RIc0daeb8_121);
xor \U$20069 ( \20091 , \20089 , \20090 );
buf \U$20070 ( \20092 , \20091 );
buf \U$20071 ( \20093 , \20092 );
not \U$20072 ( \20094 , \20093 );
buf \U$20073 ( \20095 , \12962 );
buf \U$20074 ( \20096 , \12964 );
and \U$20075 ( \20097 , \20095 , \20096 );
buf \U$20076 ( \20098 , \20097 );
buf \U$20077 ( \20099 , \20098 );
not \U$20078 ( \20100 , \20099 );
or \U$20079 ( \20101 , \20094 , \20100 );
buf \U$20080 ( \20102 , \12975 );
buf \U$20081 ( \20103 , \19482 );
nand \U$20082 ( \20104 , \20102 , \20103 );
buf \U$20083 ( \20105 , \20104 );
buf \U$20084 ( \20106 , \20105 );
nand \U$20085 ( \20107 , \20101 , \20106 );
buf \U$20086 ( \20108 , \20107 );
buf \U$20087 ( \20109 , \20108 );
buf \U$20088 ( \20110 , RIc0d8de8_51);
buf \U$20089 ( \20111 , RIc0d9dd8_85);
xor \U$20090 ( \20112 , \20110 , \20111 );
buf \U$20091 ( \20113 , \20112 );
buf \U$20092 ( \20114 , \20113 );
not \U$20093 ( \20115 , \20114 );
buf \U$20094 ( \20116 , \2393 );
not \U$20095 ( \20117 , \20116 );
or \U$20096 ( \20118 , \20115 , \20117 );
buf \U$20097 ( \20119 , \17010 );
buf \U$20098 ( \20120 , \19652 );
nand \U$20099 ( \20121 , \20119 , \20120 );
buf \U$20100 ( \20122 , \20121 );
buf \U$20101 ( \20123 , \20122 );
nand \U$20102 ( \20124 , \20118 , \20123 );
buf \U$20103 ( \20125 , \20124 );
buf \U$20104 ( \20126 , \20125 );
or \U$20105 ( \20127 , \20109 , \20126 );
buf \U$20106 ( \20128 , RIc0d8ed8_53);
buf \U$20107 ( \20129 , RIc0d9ce8_83);
xor \U$20108 ( \20130 , \20128 , \20129 );
buf \U$20109 ( \20131 , \20130 );
buf \U$20110 ( \20132 , \20131 );
not \U$20111 ( \20133 , \20132 );
buf \U$20112 ( \20134 , \12254 );
not \U$20113 ( \20135 , \20134 );
or \U$20114 ( \20136 , \20133 , \20135 );
buf \U$20115 ( \20137 , \584 );
buf \U$20116 ( \20138 , \19377 );
nand \U$20117 ( \20139 , \20137 , \20138 );
buf \U$20118 ( \20140 , \20139 );
buf \U$20119 ( \20141 , \20140 );
nand \U$20120 ( \20142 , \20136 , \20141 );
buf \U$20121 ( \20143 , \20142 );
buf \U$20122 ( \20144 , \20143 );
nand \U$20123 ( \20145 , \20127 , \20144 );
buf \U$20124 ( \20146 , \20145 );
buf \U$20125 ( \20147 , \20146 );
buf \U$20126 ( \20148 , \20108 );
buf \U$20127 ( \20149 , \20125 );
nand \U$20128 ( \20150 , \20148 , \20149 );
buf \U$20129 ( \20151 , \20150 );
buf \U$20130 ( \20152 , \20151 );
nand \U$20131 ( \20153 , \20147 , \20152 );
buf \U$20132 ( \20154 , \20153 );
buf \U$20133 ( \20155 , \20154 );
buf \U$20134 ( \20156 , RIc0d8fc8_55);
buf \U$20135 ( \20157 , RIc0d9bf8_81);
xor \U$20136 ( \20158 , \20156 , \20157 );
buf \U$20137 ( \20159 , \20158 );
buf \U$20138 ( \20160 , \20159 );
not \U$20139 ( \20161 , \20160 );
buf \U$20140 ( \20162 , \19544 );
not \U$20141 ( \20163 , \20162 );
or \U$20142 ( \20164 , \20161 , \20163 );
buf \U$20143 ( \20165 , \1077 );
buf \U$20144 ( \20166 , \19540 );
nand \U$20145 ( \20167 , \20165 , \20166 );
buf \U$20146 ( \20168 , \20167 );
buf \U$20147 ( \20169 , \20168 );
nand \U$20148 ( \20170 , \20164 , \20169 );
buf \U$20149 ( \20171 , \20170 );
buf \U$20150 ( \20172 , \20171 );
not \U$20151 ( \20173 , \20172 );
buf \U$20152 ( \20174 , \20173 );
buf \U$20153 ( \20175 , \20174 );
not \U$20154 ( \20176 , \20175 );
buf \U$20155 ( \20177 , \13860 );
not \U$20156 ( \20178 , \20177 );
buf \U$20157 ( \20179 , \20178 );
buf \U$20158 ( \20180 , \20179 );
buf \U$20159 ( \20181 , RIc0d8938_41);
buf \U$20160 ( \20182 , RIc0da288_95);
xor \U$20161 ( \20183 , \20181 , \20182 );
buf \U$20162 ( \20184 , \20183 );
buf \U$20163 ( \20185 , \20184 );
not \U$20164 ( \20186 , \20185 );
buf \U$20165 ( \20187 , \20186 );
buf \U$20166 ( \20188 , \20187 );
or \U$20167 ( \20189 , \20180 , \20188 );
buf \U$20168 ( \20190 , \13873 );
not \U$20169 ( \20191 , \20190 );
buf \U$20170 ( \20192 , \20191 );
buf \U$20171 ( \20193 , \20192 );
buf \U$20172 ( \20194 , \19953 );
or \U$20173 ( \20195 , \20193 , \20194 );
nand \U$20174 ( \20196 , \20189 , \20195 );
buf \U$20175 ( \20197 , \20196 );
not \U$20176 ( \20198 , \20197 );
buf \U$20177 ( \20199 , \20198 );
not \U$20178 ( \20200 , \20199 );
or \U$20179 ( \20201 , \20176 , \20200 );
buf \U$20180 ( \20202 , RIc0d82a8_27);
buf \U$20181 ( \20203 , RIc0da918_109);
xor \U$20182 ( \20204 , \20202 , \20203 );
buf \U$20183 ( \20205 , \20204 );
buf \U$20184 ( \20206 , \20205 );
not \U$20185 ( \20207 , \20206 );
buf \U$20186 ( \20208 , \13419 );
not \U$20187 ( \20209 , \20208 );
or \U$20188 ( \20210 , \20207 , \20209 );
buf \U$20191 ( \20211 , \13408 );
buf \U$20192 ( \20212 , \20211 );
buf \U$20193 ( \20213 , \19313 );
nand \U$20194 ( \20214 , \20212 , \20213 );
buf \U$20195 ( \20215 , \20214 );
buf \U$20196 ( \20216 , \20215 );
nand \U$20197 ( \20217 , \20210 , \20216 );
buf \U$20198 ( \20218 , \20217 );
buf \U$20199 ( \20219 , \20218 );
nand \U$20200 ( \20220 , \20201 , \20219 );
buf \U$20201 ( \20221 , \20220 );
buf \U$20202 ( \20222 , \20221 );
buf \U$20203 ( \20223 , \20197 );
buf \U$20204 ( \20224 , \20171 );
nand \U$20205 ( \20225 , \20223 , \20224 );
buf \U$20206 ( \20226 , \20225 );
buf \U$20207 ( \20227 , \20226 );
nand \U$20208 ( \20228 , \20222 , \20227 );
buf \U$20209 ( \20229 , \20228 );
buf \U$20210 ( \20230 , \20229 );
xor \U$20211 ( \20231 , \20155 , \20230 );
buf \U$20212 ( \20232 , RIc0d8578_33);
buf \U$20213 ( \20233 , RIc0da648_103);
xor \U$20214 ( \20234 , \20232 , \20233 );
buf \U$20215 ( \20235 , \20234 );
buf \U$20216 ( \20236 , \20235 );
not \U$20217 ( \20237 , \20236 );
buf \U$20218 ( \20238 , \15397 );
not \U$20219 ( \20239 , \20238 );
or \U$20220 ( \20240 , \20237 , \20239 );
buf \U$20221 ( \20241 , \4475 );
not \U$20222 ( \20242 , \20241 );
buf \U$20223 ( \20243 , \20242 );
buf \U$20224 ( \20244 , \20243 );
buf \U$20225 ( \20245 , \18215 );
nand \U$20226 ( \20246 , \20244 , \20245 );
buf \U$20227 ( \20247 , \20246 );
buf \U$20228 ( \20248 , \20247 );
nand \U$20229 ( \20249 , \20240 , \20248 );
buf \U$20230 ( \20250 , \20249 );
buf \U$20231 ( \20251 , \20250 );
buf \U$20232 ( \20252 , RIc0d81b8_25);
buf \U$20233 ( \20253 , RIc0daa08_111);
xor \U$20234 ( \20254 , \20252 , \20253 );
buf \U$20235 ( \20255 , \20254 );
buf \U$20236 ( \20256 , \20255 );
not \U$20237 ( \20257 , \20256 );
buf \U$20238 ( \20258 , \12529 );
not \U$20239 ( \20259 , \20258 );
or \U$20240 ( \20260 , \20257 , \20259 );
buf \U$20241 ( \20261 , \14106 );
buf \U$20242 ( \20262 , \19968 );
nand \U$20243 ( \20263 , \20261 , \20262 );
buf \U$20244 ( \20264 , \20263 );
buf \U$20245 ( \20265 , \20264 );
nand \U$20246 ( \20266 , \20260 , \20265 );
buf \U$20247 ( \20267 , \20266 );
buf \U$20248 ( \20268 , \20267 );
xor \U$20249 ( \20269 , \20251 , \20268 );
buf \U$20250 ( \20270 , RIc0da378_97);
buf \U$20251 ( \20271 , RIc0d8848_39);
xor \U$20252 ( \20272 , \20270 , \20271 );
buf \U$20253 ( \20273 , \20272 );
buf \U$20254 ( \20274 , \20273 );
not \U$20255 ( \20275 , \20274 );
buf \U$20256 ( \20276 , \2066 );
not \U$20257 ( \20277 , \20276 );
or \U$20258 ( \20278 , \20275 , \20277 );
buf \U$20259 ( \20279 , \734 );
buf \U$20260 ( \20280 , \18193 );
nand \U$20261 ( \20281 , \20279 , \20280 );
buf \U$20262 ( \20282 , \20281 );
buf \U$20263 ( \20283 , \20282 );
nand \U$20264 ( \20284 , \20278 , \20283 );
buf \U$20265 ( \20285 , \20284 );
buf \U$20266 ( \20286 , \20285 );
and \U$20267 ( \20287 , \20269 , \20286 );
and \U$20268 ( \20288 , \20251 , \20268 );
or \U$20269 ( \20289 , \20287 , \20288 );
buf \U$20270 ( \20290 , \20289 );
buf \U$20271 ( \20291 , \20290 );
and \U$20272 ( \20292 , \20231 , \20291 );
and \U$20273 ( \20293 , \20155 , \20230 );
or \U$20274 ( \20294 , \20292 , \20293 );
buf \U$20275 ( \20295 , \20294 );
buf \U$20276 ( \20296 , \20295 );
and \U$20277 ( \20297 , \20088 , \20296 );
and \U$20278 ( \20298 , \20084 , \20087 );
or \U$20279 ( \20299 , \20297 , \20298 );
buf \U$20280 ( \20300 , \20299 );
buf \U$20281 ( \20301 , \20300 );
and \U$20282 ( \20302 , \20081 , \20301 );
and \U$20283 ( \20303 , \20061 , \20080 );
or \U$20284 ( \20304 , \20302 , \20303 );
buf \U$20285 ( \20305 , \20304 );
buf \U$20286 ( \20306 , \20305 );
and \U$20287 ( \20307 , \20057 , \20306 );
and \U$20288 ( \20308 , \19902 , \20056 );
or \U$20289 ( \20309 , \20307 , \20308 );
buf \U$20290 ( \20310 , \20309 );
buf \U$20291 ( \20311 , \20310 );
not \U$20292 ( \20312 , \20311 );
xor \U$20293 ( \20313 , \18258 , \18261 );
xor \U$20294 ( \20314 , \20313 , \18566 );
buf \U$20295 ( \20315 , \20314 );
buf \U$20296 ( \20316 , \20315 );
not \U$20297 ( \20317 , \20316 );
or \U$20298 ( \20318 , \20312 , \20317 );
buf \U$20299 ( \20319 , \20315 );
buf \U$20300 ( \20320 , \20310 );
or \U$20301 ( \20321 , \20319 , \20320 );
xor \U$20302 ( \20322 , \17794 , \17655 );
xor \U$20303 ( \20323 , \20322 , \17672 );
buf \U$20304 ( \20324 , \20323 );
nand \U$20305 ( \20325 , \20321 , \20324 );
buf \U$20306 ( \20326 , \20325 );
buf \U$20307 ( \20327 , \20326 );
nand \U$20308 ( \20328 , \20318 , \20327 );
buf \U$20309 ( \20329 , \20328 );
buf \U$20310 ( \20330 , \20329 );
nand \U$20311 ( \20331 , \19898 , \20330 );
buf \U$20312 ( \20332 , \20331 );
buf \U$20313 ( \20333 , \20332 );
buf \U$20314 ( \20334 , \19895 );
buf \U$20315 ( \20335 , \19887 );
or \U$20316 ( \20336 , \20334 , \20335 );
buf \U$20317 ( \20337 , \20336 );
buf \U$20318 ( \20338 , \20337 );
nand \U$20319 ( \20339 , \20333 , \20338 );
buf \U$20320 ( \20340 , \20339 );
buf \U$20321 ( \20341 , \20340 );
not \U$20322 ( \20342 , \20341 );
or \U$20323 ( \20343 , \19309 , \20342 );
xor \U$20324 ( \20344 , \17839 , \17922 );
xor \U$20325 ( \20345 , \20344 , \18835 );
buf \U$20326 ( \20346 , \20345 );
buf \U$20327 ( \20347 , \20346 );
buf \U$20328 ( \20348 , \19307 );
not \U$20329 ( \20349 , \20348 );
buf \U$20330 ( \20350 , \20340 );
not \U$20331 ( \20351 , \20350 );
buf \U$20332 ( \20352 , \20351 );
buf \U$20333 ( \20353 , \20352 );
nand \U$20334 ( \20354 , \20349 , \20353 );
buf \U$20335 ( \20355 , \20354 );
buf \U$20336 ( \20356 , \20355 );
nand \U$20337 ( \20357 , \20347 , \20356 );
buf \U$20338 ( \20358 , \20357 );
buf \U$20339 ( \20359 , \20358 );
nand \U$20340 ( \20360 , \20343 , \20359 );
buf \U$20341 ( \20361 , \20360 );
buf \U$20342 ( \20362 , \20361 );
nand \U$20343 ( \20363 , \19304 , \20362 );
buf \U$20344 ( \20364 , \20363 );
buf \U$20345 ( \20365 , \20364 );
buf \U$20346 ( \20366 , \15524 );
not \U$20347 ( \20367 , \20366 );
buf \U$20348 ( \20368 , \20367 );
buf \U$20349 ( \20369 , \20368 );
not \U$20350 ( \20370 , \20369 );
buf \U$20351 ( \20371 , \15956 );
not \U$20352 ( \20372 , \20371 );
or \U$20353 ( \20373 , \20370 , \20372 );
buf \U$20354 ( \20374 , \15524 );
not \U$20355 ( \20375 , \20374 );
buf \U$20356 ( \20376 , \15950 );
not \U$20357 ( \20377 , \20376 );
or \U$20358 ( \20378 , \20375 , \20377 );
buf \U$20359 ( \20379 , \15733 );
nand \U$20360 ( \20380 , \20378 , \20379 );
buf \U$20361 ( \20381 , \20380 );
buf \U$20362 ( \20382 , \20381 );
nand \U$20363 ( \20383 , \20373 , \20382 );
buf \U$20364 ( \20384 , \20383 );
buf \U$20365 ( \20385 , \20384 );
not \U$20366 ( \20386 , \20385 );
buf \U$20367 ( \20387 , \15599 );
not \U$20368 ( \20388 , \20387 );
buf \U$20369 ( \20389 , \15723 );
not \U$20370 ( \20390 , \20389 );
or \U$20371 ( \20391 , \20388 , \20390 );
buf \U$20372 ( \20392 , \15667 );
nand \U$20373 ( \20393 , \20391 , \20392 );
buf \U$20374 ( \20394 , \20393 );
buf \U$20375 ( \20395 , \20394 );
buf \U$20376 ( \20396 , \15599 );
not \U$20377 ( \20397 , \20396 );
buf \U$20378 ( \20398 , \15726 );
nand \U$20379 ( \20399 , \20397 , \20398 );
buf \U$20380 ( \20400 , \20399 );
buf \U$20381 ( \20401 , \20400 );
nand \U$20382 ( \20402 , \20395 , \20401 );
buf \U$20383 ( \20403 , \20402 );
buf \U$20384 ( \20404 , \20403 );
not \U$20385 ( \20405 , \20404 );
buf \U$20386 ( \20406 , \15820 );
not \U$20387 ( \20407 , \20406 );
buf \U$20388 ( \20408 , \15878 );
not \U$20389 ( \20409 , \20408 );
or \U$20390 ( \20410 , \20407 , \20409 );
buf \U$20391 ( \20411 , \15878 );
buf \U$20392 ( \20412 , \15820 );
or \U$20393 ( \20413 , \20411 , \20412 );
buf \U$20394 ( \20414 , \15947 );
nand \U$20395 ( \20415 , \20413 , \20414 );
buf \U$20396 ( \20416 , \20415 );
buf \U$20397 ( \20417 , \20416 );
nand \U$20398 ( \20418 , \20410 , \20417 );
buf \U$20399 ( \20419 , \20418 );
buf \U$20400 ( \20420 , \20419 );
not \U$20401 ( \20421 , \20420 );
buf \U$20402 ( \20422 , \20421 );
buf \U$20403 ( \20423 , \20422 );
not \U$20404 ( \20424 , \20423 );
or \U$20405 ( \20425 , \20405 , \20424 );
buf \U$20406 ( \20426 , \20403 );
buf \U$20407 ( \20427 , \20422 );
or \U$20408 ( \20428 , \20426 , \20427 );
buf \U$20409 ( \20429 , \20428 );
buf \U$20410 ( \20430 , \20429 );
nand \U$20411 ( \20431 , \20425 , \20430 );
buf \U$20412 ( \20432 , \20431 );
buf \U$20413 ( \20433 , \20432 );
not \U$20414 ( \20434 , \15094 );
nand \U$20415 ( \20435 , \20434 , \15078 );
not \U$20416 ( \20436 , \20435 );
not \U$20417 ( \20437 , \15132 );
or \U$20418 ( \20438 , \20436 , \20437 );
buf \U$20419 ( \20439 , \15094 );
buf \U$20420 ( \20440 , \15075 );
nand \U$20421 ( \20441 , \20439 , \20440 );
buf \U$20422 ( \20442 , \20441 );
nand \U$20423 ( \20443 , \20438 , \20442 );
buf \U$20424 ( \20444 , \20443 );
not \U$20425 ( \20445 , \20444 );
buf \U$20426 ( \20446 , \20445 );
buf \U$20427 ( \20447 , \20446 );
and \U$20428 ( \20448 , \20433 , \20447 );
not \U$20429 ( \20449 , \20433 );
buf \U$20430 ( \20450 , \20443 );
and \U$20431 ( \20451 , \20449 , \20450 );
nor \U$20432 ( \20452 , \20448 , \20451 );
buf \U$20433 ( \20453 , \20452 );
buf \U$20434 ( \20454 , \20453 );
not \U$20435 ( \20455 , \20454 );
or \U$20436 ( \20456 , \20386 , \20455 );
buf \U$20437 ( \20457 , \20453 );
buf \U$20438 ( \20458 , \20384 );
or \U$20439 ( \20459 , \20457 , \20458 );
nand \U$20440 ( \20460 , \20456 , \20459 );
buf \U$20441 ( \20461 , \20460 );
buf \U$20442 ( \20462 , \20461 );
not \U$20443 ( \20463 , \15514 );
buf \U$20444 ( \20464 , \15449 );
not \U$20445 ( \20465 , \20464 );
buf \U$20446 ( \20466 , \15390 );
nand \U$20447 ( \20467 , \20465 , \20466 );
buf \U$20448 ( \20468 , \20467 );
not \U$20449 ( \20469 , \20468 );
or \U$20450 ( \20470 , \20463 , \20469 );
buf \U$20451 ( \20471 , \15390 );
not \U$20452 ( \20472 , \20471 );
buf \U$20453 ( \20473 , \15449 );
nand \U$20454 ( \20474 , \20472 , \20473 );
buf \U$20455 ( \20475 , \20474 );
nand \U$20456 ( \20476 , \20470 , \20475 );
not \U$20457 ( \20477 , \15561 );
not \U$20458 ( \20478 , \15589 );
or \U$20459 ( \20479 , \20477 , \20478 );
not \U$20460 ( \20480 , \15592 );
not \U$20461 ( \20481 , \15564 );
or \U$20462 ( \20482 , \20480 , \20481 );
nand \U$20463 ( \20483 , \20482 , \15542 );
nand \U$20464 ( \20484 , \20479 , \20483 );
buf \U$20465 ( \20485 , \20484 );
not \U$20466 ( \20486 , \20485 );
buf \U$20467 ( \20487 , \20486 );
buf \U$20468 ( \20488 , \20487 );
buf \U$20469 ( \20489 , \19082 );
not \U$20470 ( \20490 , \20489 );
buf \U$20471 ( \20491 , \19068 );
not \U$20472 ( \20492 , \20491 );
or \U$20473 ( \20493 , \20490 , \20492 );
buf \U$20474 ( \20494 , \19068 );
buf \U$20475 ( \20495 , \19082 );
or \U$20476 ( \20496 , \20494 , \20495 );
buf \U$20477 ( \20497 , \19055 );
nand \U$20478 ( \20498 , \20496 , \20497 );
buf \U$20479 ( \20499 , \20498 );
buf \U$20480 ( \20500 , \20499 );
nand \U$20481 ( \20501 , \20493 , \20500 );
buf \U$20482 ( \20502 , \20501 );
buf \U$20483 ( \20503 , \20502 );
not \U$20484 ( \20504 , \20503 );
buf \U$20485 ( \20505 , \20504 );
buf \U$20486 ( \20506 , \20505 );
and \U$20487 ( \20507 , \20488 , \20506 );
not \U$20488 ( \20508 , \20488 );
buf \U$20489 ( \20509 , \20502 );
and \U$20490 ( \20510 , \20508 , \20509 );
nor \U$20491 ( \20511 , \20507 , \20510 );
buf \U$20492 ( \20512 , \20511 );
buf \U$20493 ( \20513 , \20512 );
xor \U$20494 ( \20514 , \15098 , \15112 );
and \U$20495 ( \20515 , \20514 , \15130 );
and \U$20496 ( \20516 , \15098 , \15112 );
or \U$20497 ( \20517 , \20515 , \20516 );
buf \U$20498 ( \20518 , \20517 );
buf \U$20499 ( \20519 , \20518 );
not \U$20500 ( \20520 , \20519 );
buf \U$20501 ( \20521 , \20520 );
buf \U$20502 ( \20522 , \20521 );
and \U$20503 ( \20523 , \20513 , \20522 );
not \U$20504 ( \20524 , \20513 );
buf \U$20505 ( \20525 , \20518 );
and \U$20506 ( \20526 , \20524 , \20525 );
nor \U$20507 ( \20527 , \20523 , \20526 );
buf \U$20508 ( \20528 , \20527 );
and \U$20509 ( \20529 , \20476 , \20528 );
not \U$20510 ( \20530 , \20476 );
buf \U$20511 ( \20531 , \20528 );
not \U$20512 ( \20532 , \20531 );
buf \U$20513 ( \20533 , \20532 );
and \U$20514 ( \20534 , \20530 , \20533 );
or \U$20515 ( \20535 , \20529 , \20534 );
buf \U$20516 ( \20536 , \20535 );
buf \U$20517 ( \20537 , \15380 );
buf \U$20518 ( \20538 , \15343 );
nor \U$20519 ( \20539 , \20537 , \20538 );
buf \U$20520 ( \20540 , \20539 );
buf \U$20521 ( \20541 , \20540 );
buf \U$20522 ( \20542 , \15362 );
or \U$20523 ( \20543 , \20541 , \20542 );
buf \U$20524 ( \20544 , \15380 );
buf \U$20525 ( \20545 , \15343 );
nand \U$20526 ( \20546 , \20544 , \20545 );
buf \U$20527 ( \20547 , \20546 );
buf \U$20528 ( \20548 , \20547 );
nand \U$20529 ( \20549 , \20543 , \20548 );
buf \U$20530 ( \20550 , \20549 );
xor \U$20531 ( \20551 , \15415 , \15432 );
and \U$20532 ( \20552 , \20551 , \15447 );
and \U$20533 ( \20553 , \15415 , \15432 );
or \U$20534 ( \20554 , \20552 , \20553 );
buf \U$20535 ( \20555 , \20554 );
xor \U$20536 ( \20556 , \20550 , \20555 );
xor \U$20537 ( \20557 , \15620 , \15637 );
and \U$20538 ( \20558 , \20557 , \15665 );
and \U$20539 ( \20559 , \15620 , \15637 );
or \U$20540 ( \20560 , \20558 , \20559 );
buf \U$20541 ( \20561 , \20560 );
xnor \U$20542 ( \20562 , \20556 , \20561 );
buf \U$20543 ( \20563 , \20562 );
and \U$20544 ( \20564 , \20536 , \20563 );
not \U$20545 ( \20565 , \20536 );
buf \U$20546 ( \20566 , \20562 );
not \U$20547 ( \20567 , \20566 );
buf \U$20548 ( \20568 , \20567 );
buf \U$20549 ( \20569 , \20568 );
and \U$20550 ( \20570 , \20565 , \20569 );
nor \U$20551 ( \20571 , \20564 , \20570 );
buf \U$20552 ( \20572 , \20571 );
buf \U$20553 ( \20573 , \20572 );
and \U$20554 ( \20574 , \20462 , \20573 );
not \U$20555 ( \20575 , \20462 );
buf \U$20556 ( \20576 , \20572 );
not \U$20557 ( \20577 , \20576 );
buf \U$20558 ( \20578 , \20577 );
buf \U$20559 ( \20579 , \20578 );
and \U$20560 ( \20580 , \20575 , \20579 );
nor \U$20561 ( \20581 , \20574 , \20580 );
buf \U$20562 ( \20582 , \20581 );
buf \U$20563 ( \20583 , \20582 );
buf \U$20564 ( \20584 , \15317 );
not \U$20565 ( \20585 , \20584 );
buf \U$20566 ( \20586 , \15960 );
nand \U$20567 ( \20587 , \20585 , \20586 );
buf \U$20568 ( \20588 , \20587 );
buf \U$20569 ( \20589 , \20588 );
not \U$20570 ( \20590 , \20589 );
buf \U$20571 ( \20591 , \16848 );
not \U$20572 ( \20592 , \20591 );
or \U$20573 ( \20593 , \20590 , \20592 );
buf \U$20574 ( \20594 , \15960 );
not \U$20575 ( \20595 , \20594 );
buf \U$20576 ( \20596 , \15317 );
nand \U$20577 ( \20597 , \20595 , \20596 );
buf \U$20578 ( \20598 , \20597 );
buf \U$20579 ( \20599 , \20598 );
nand \U$20580 ( \20600 , \20593 , \20599 );
buf \U$20581 ( \20601 , \20600 );
buf \U$20582 ( \20602 , \20601 );
not \U$20583 ( \20603 , \20602 );
buf \U$20584 ( \20604 , \20603 );
buf \U$20585 ( \20605 , \20604 );
xor \U$20586 ( \20606 , \20583 , \20605 );
buf \U$20587 ( \20607 , \15702 );
not \U$20588 ( \20608 , \20607 );
buf \U$20589 ( \20609 , \15995 );
not \U$20590 ( \20610 , \20609 );
or \U$20591 ( \20611 , \20608 , \20610 );
buf \U$20592 ( \20612 , \481 );
buf \U$20593 ( \20613 , RIc0d8578_33);
buf \U$20594 ( \20614 , RIc0da198_93);
xor \U$20595 ( \20615 , \20613 , \20614 );
buf \U$20596 ( \20616 , \20615 );
buf \U$20597 ( \20617 , \20616 );
nand \U$20598 ( \20618 , \20612 , \20617 );
buf \U$20599 ( \20619 , \20618 );
buf \U$20600 ( \20620 , \20619 );
nand \U$20601 ( \20621 , \20611 , \20620 );
buf \U$20602 ( \20622 , \20621 );
buf \U$20603 ( \20623 , \15583 );
not \U$20604 ( \20624 , \20623 );
buf \U$20605 ( \20625 , \16942 );
not \U$20606 ( \20626 , \20625 );
or \U$20607 ( \20627 , \20624 , \20626 );
buf \U$20608 ( \20628 , \442 );
buf \U$20609 ( \20629 , RIc0d8758_37);
buf \U$20610 ( \20630 , RIc0d9fb8_89);
xor \U$20611 ( \20631 , \20629 , \20630 );
buf \U$20612 ( \20632 , \20631 );
buf \U$20613 ( \20633 , \20632 );
nand \U$20614 ( \20634 , \20628 , \20633 );
buf \U$20615 ( \20635 , \20634 );
buf \U$20616 ( \20636 , \20635 );
nand \U$20617 ( \20637 , \20627 , \20636 );
buf \U$20618 ( \20638 , \20637 );
xnor \U$20619 ( \20639 , \20622 , \20638 );
buf \U$20620 ( \20640 , \15374 );
not \U$20621 ( \20641 , \20640 );
buf \U$20622 ( \20642 , \14532 );
not \U$20623 ( \20643 , \20642 );
or \U$20624 ( \20644 , \20641 , \20643 );
buf \U$20625 ( \20645 , \1078 );
buf \U$20626 ( \20646 , RIc0d8b18_45);
buf \U$20627 ( \20647 , RIc0d9bf8_81);
xor \U$20628 ( \20648 , \20646 , \20647 );
buf \U$20629 ( \20649 , \20648 );
buf \U$20630 ( \20650 , \20649 );
nand \U$20631 ( \20651 , \20645 , \20650 );
buf \U$20632 ( \20652 , \20651 );
buf \U$20633 ( \20653 , \20652 );
nand \U$20634 ( \20654 , \20644 , \20653 );
buf \U$20635 ( \20655 , \20654 );
buf \U$20636 ( \20656 , \20655 );
not \U$20637 ( \20657 , \20656 );
buf \U$20638 ( \20658 , \20657 );
and \U$20639 ( \20659 , \20639 , \20658 );
not \U$20640 ( \20660 , \20639 );
and \U$20641 ( \20661 , \20660 , \20655 );
nor \U$20642 ( \20662 , \20659 , \20661 );
buf \U$20643 ( \20663 , \20662 );
buf \U$20644 ( \20664 , \15752 );
not \U$20645 ( \20665 , \20664 );
buf \U$20646 ( \20666 , \13332 );
not \U$20647 ( \20667 , \20666 );
or \U$20648 ( \20668 , \20665 , \20667 );
buf \U$20649 ( \20669 , \874 );
buf \U$20650 ( \20670 , RIc0d90b8_57);
buf \U$20651 ( \20671 , RIc0d9658_69);
xor \U$20652 ( \20672 , \20670 , \20671 );
buf \U$20653 ( \20673 , \20672 );
buf \U$20654 ( \20674 , \20673 );
nand \U$20655 ( \20675 , \20669 , \20674 );
buf \U$20656 ( \20676 , \20675 );
buf \U$20657 ( \20677 , \20676 );
nand \U$20658 ( \20678 , \20668 , \20677 );
buf \U$20659 ( \20679 , \20678 );
buf \U$20660 ( \20680 , \20679 );
buf \U$20661 ( \20681 , \15773 );
not \U$20662 ( \20682 , \20681 );
buf \U$20663 ( \20683 , \2358 );
not \U$20664 ( \20684 , \20683 );
or \U$20665 ( \20685 , \20682 , \20684 );
buf \U$20666 ( \20686 , \1143 );
buf \U$20667 ( \20687 , RIc0d8de8_51);
buf \U$20668 ( \20688 , RIc0d9928_75);
xor \U$20669 ( \20689 , \20687 , \20688 );
buf \U$20670 ( \20690 , \20689 );
buf \U$20671 ( \20691 , \20690 );
nand \U$20672 ( \20692 , \20686 , \20691 );
buf \U$20673 ( \20693 , \20692 );
buf \U$20674 ( \20694 , \20693 );
nand \U$20675 ( \20695 , \20685 , \20694 );
buf \U$20676 ( \20696 , \20695 );
buf \U$20677 ( \20697 , \20696 );
xor \U$20678 ( \20698 , \20680 , \20697 );
buf \U$20679 ( \20699 , \15485 );
not \U$20680 ( \20700 , \20699 );
buf \U$20681 ( \20701 , \330 );
not \U$20682 ( \20702 , \20701 );
or \U$20683 ( \20703 , \20700 , \20702 );
buf \U$20684 ( \20704 , \343 );
buf \U$20685 ( \20705 , RIc0da288_95);
buf \U$20686 ( \20706 , RIc0d8488_31);
xor \U$20687 ( \20707 , \20705 , \20706 );
buf \U$20688 ( \20708 , \20707 );
buf \U$20689 ( \20709 , \20708 );
nand \U$20690 ( \20710 , \20704 , \20709 );
buf \U$20691 ( \20711 , \20710 );
buf \U$20692 ( \20712 , \20711 );
nand \U$20693 ( \20713 , \20703 , \20712 );
buf \U$20694 ( \20714 , \20713 );
buf \U$20695 ( \20715 , \20714 );
xor \U$20696 ( \20716 , \20698 , \20715 );
buf \U$20697 ( \20717 , \20716 );
buf \U$20698 ( \20718 , \20717 );
xor \U$20699 ( \20719 , \20663 , \20718 );
buf \U$20700 ( \20720 , \15630 );
not \U$20701 ( \20721 , \20720 );
buf \U$20702 ( \20722 , \12795 );
not \U$20703 ( \20723 , \20722 );
or \U$20704 ( \20724 , \20721 , \20723 );
buf \U$20705 ( \20725 , \1229 );
buf \U$20706 ( \20726 , RIc0d9298_61);
buf \U$20707 ( \20727 , RIc0d9478_65);
xor \U$20708 ( \20728 , \20726 , \20727 );
buf \U$20709 ( \20729 , \20728 );
buf \U$20710 ( \20730 , \20729 );
nand \U$20711 ( \20731 , \20725 , \20730 );
buf \U$20712 ( \20732 , \20731 );
buf \U$20713 ( \20733 , \20732 );
nand \U$20714 ( \20734 , \20724 , \20733 );
buf \U$20715 ( \20735 , \20734 );
buf \U$20716 ( \20736 , \20735 );
buf \U$20717 ( \20737 , \15890 );
not \U$20718 ( \20738 , \20737 );
buf \U$20719 ( \20739 , \12331 );
not \U$20720 ( \20740 , \20739 );
buf \U$20721 ( \20741 , \20740 );
buf \U$20722 ( \20742 , \20741 );
not \U$20723 ( \20743 , \20742 );
or \U$20724 ( \20744 , \20738 , \20743 );
buf \U$20725 ( \20745 , \12342 );
xor \U$20726 ( \20746 , RIc0da828_107, RIc0d7ee8_19);
buf \U$20727 ( \20747 , \20746 );
nand \U$20728 ( \20748 , \20745 , \20747 );
buf \U$20729 ( \20749 , \20748 );
buf \U$20730 ( \20750 , \20749 );
nand \U$20731 ( \20751 , \20744 , \20750 );
buf \U$20732 ( \20752 , \20751 );
buf \U$20733 ( \20753 , \20752 );
xor \U$20734 ( \20754 , \20736 , \20753 );
buf \U$20735 ( \20755 , \15914 );
not \U$20736 ( \20756 , \20755 );
buf \U$20737 ( \20757 , \14207 );
not \U$20738 ( \20758 , \20757 );
buf \U$20739 ( \20759 , \20758 );
buf \U$20740 ( \20760 , \20759 );
not \U$20741 ( \20761 , \20760 );
or \U$20742 ( \20762 , \20756 , \20761 );
buf \U$20743 ( \20763 , \20211 );
xor \U$20744 ( \20764 , RIc0da918_109, RIc0d7df8_17);
buf \U$20745 ( \20765 , \20764 );
nand \U$20746 ( \20766 , \20763 , \20765 );
buf \U$20747 ( \20767 , \20766 );
buf \U$20748 ( \20768 , \20767 );
nand \U$20749 ( \20769 , \20762 , \20768 );
buf \U$20750 ( \20770 , \20769 );
buf \U$20751 ( \20771 , \20770 );
xor \U$20752 ( \20772 , \20754 , \20771 );
buf \U$20753 ( \20773 , \20772 );
buf \U$20754 ( \20774 , \20773 );
xor \U$20755 ( \20775 , \20719 , \20774 );
buf \U$20756 ( \20776 , \20775 );
buf \U$20757 ( \20777 , \20776 );
not \U$20758 ( \20778 , \20777 );
buf \U$20759 ( \20779 , \15425 );
not \U$20760 ( \20780 , \20779 );
buf \U$20761 ( \20781 , \20098 );
not \U$20762 ( \20782 , \20781 );
or \U$20763 ( \20783 , \20780 , \20782 );
buf \U$20764 ( \20784 , \12975 );
xor \U$20765 ( \20785 , RIc0daeb8_121, RIc0d7858_5);
buf \U$20766 ( \20786 , \20785 );
nand \U$20767 ( \20787 , \20784 , \20786 );
buf \U$20768 ( \20788 , \20787 );
buf \U$20769 ( \20789 , \20788 );
nand \U$20770 ( \20790 , \20783 , \20789 );
buf \U$20771 ( \20791 , \20790 );
buf \U$20772 ( \20792 , \15555 );
not \U$20773 ( \20793 , \20792 );
buf \U$20774 ( \20794 , \3521 );
not \U$20775 ( \20795 , \20794 );
buf \U$20776 ( \20796 , \3515 );
nor \U$20777 ( \20797 , \20795 , \20796 );
buf \U$20778 ( \20798 , \20797 );
buf \U$20779 ( \20799 , \20798 );
not \U$20780 ( \20800 , \20799 );
or \U$20781 ( \20801 , \20793 , \20800 );
buf \U$20782 ( \20802 , \15550 );
buf \U$20783 ( \20803 , RIc0d81b8_25);
buf \U$20784 ( \20804 , RIc0da558_101);
xor \U$20785 ( \20805 , \20803 , \20804 );
buf \U$20786 ( \20806 , \20805 );
buf \U$20787 ( \20807 , \20806 );
nand \U$20788 ( \20808 , \20802 , \20807 );
buf \U$20789 ( \20809 , \20808 );
buf \U$20790 ( \20810 , \20809 );
nand \U$20791 ( \20811 , \20801 , \20810 );
buf \U$20792 ( \20812 , \20811 );
xor \U$20793 ( \20813 , \20791 , \20812 );
buf \U$20794 ( \20814 , \15105 );
not \U$20795 ( \20815 , \20814 );
buf \U$20796 ( \20816 , \16402 );
not \U$20797 ( \20817 , \20816 );
or \U$20798 ( \20818 , \20815 , \20817 );
buf \U$20799 ( \20819 , \1933 );
buf \U$20800 ( \20820 , RIc0d8668_35);
buf \U$20801 ( \20821 , RIc0da0a8_91);
xor \U$20802 ( \20822 , \20820 , \20821 );
buf \U$20803 ( \20823 , \20822 );
buf \U$20804 ( \20824 , \20823 );
nand \U$20805 ( \20825 , \20819 , \20824 );
buf \U$20806 ( \20826 , \20825 );
buf \U$20807 ( \20827 , \20826 );
nand \U$20808 ( \20828 , \20818 , \20827 );
buf \U$20809 ( \20829 , \20828 );
xnor \U$20810 ( \20830 , \20813 , \20829 );
buf \U$20811 ( \20831 , \20830 );
not \U$20812 ( \20832 , \20831 );
buf \U$20813 ( \20833 , \15504 );
not \U$20814 ( \20834 , \20833 );
buf \U$20815 ( \20835 , \573 );
not \U$20816 ( \20836 , \20835 );
or \U$20817 ( \20837 , \20834 , \20836 );
buf \U$20818 ( \20838 , \993 );
buf \U$20819 ( \20839 , RIc0d8a28_43);
buf \U$20820 ( \20840 , RIc0d9ce8_83);
xor \U$20821 ( \20841 , \20839 , \20840 );
buf \U$20822 ( \20842 , \20841 );
buf \U$20823 ( \20843 , \20842 );
nand \U$20824 ( \20844 , \20838 , \20843 );
buf \U$20825 ( \20845 , \20844 );
buf \U$20826 ( \20846 , \20845 );
nand \U$20827 ( \20847 , \20837 , \20846 );
buf \U$20828 ( \20848 , \20847 );
buf \U$20829 ( \20849 , \20848 );
buf \U$20830 ( \20850 , \15869 );
not \U$20831 ( \20851 , \20850 );
buf \U$20832 ( \20852 , \14100 );
not \U$20833 ( \20853 , \20852 );
or \U$20834 ( \20854 , \20851 , \20853 );
buf \U$20835 ( \20855 , \14353 );
buf \U$20836 ( \20856 , RIc0d7d08_15);
buf \U$20837 ( \20857 , RIc0daa08_111);
xor \U$20838 ( \20858 , \20856 , \20857 );
buf \U$20839 ( \20859 , \20858 );
buf \U$20840 ( \20860 , \20859 );
nand \U$20841 ( \20861 , \20855 , \20860 );
buf \U$20842 ( \20862 , \20861 );
buf \U$20843 ( \20863 , \20862 );
nand \U$20844 ( \20864 , \20854 , \20863 );
buf \U$20845 ( \20865 , \20864 );
buf \U$20846 ( \20866 , \20865 );
xor \U$20847 ( \20867 , \20849 , \20866 );
buf \U$20848 ( \20868 , \15686 );
not \U$20849 ( \20869 , \20868 );
buf \U$20850 ( \20870 , \12402 );
not \U$20851 ( \20871 , \20870 );
or \U$20852 ( \20872 , \20869 , \20871 );
buf \U$20853 ( \20873 , \16995 );
buf \U$20854 ( \20874 , RIc0d7c18_13);
buf \U$20855 ( \20875 , RIc0daaf8_113);
xor \U$20856 ( \20876 , \20874 , \20875 );
buf \U$20857 ( \20877 , \20876 );
buf \U$20858 ( \20878 , \20877 );
nand \U$20859 ( \20879 , \20873 , \20878 );
buf \U$20860 ( \20880 , \20879 );
buf \U$20861 ( \20881 , \20880 );
nand \U$20862 ( \20882 , \20872 , \20881 );
buf \U$20863 ( \20883 , \20882 );
buf \U$20864 ( \20884 , \20883 );
xor \U$20865 ( \20885 , \20867 , \20884 );
buf \U$20866 ( \20886 , \20885 );
buf \U$20867 ( \20887 , \20886 );
not \U$20868 ( \20888 , \20887 );
or \U$20869 ( \20889 , \20832 , \20888 );
buf \U$20870 ( \20890 , \20830 );
buf \U$20871 ( \20891 , \20886 );
or \U$20872 ( \20892 , \20890 , \20891 );
nand \U$20873 ( \20893 , \20889 , \20892 );
buf \U$20874 ( \20894 , \20893 );
buf \U$20875 ( \20895 , \20894 );
buf \U$20876 ( \20896 , \15408 );
not \U$20877 ( \20897 , \20896 );
buf \U$20878 ( \20898 , \15397 );
not \U$20879 ( \20899 , \20898 );
or \U$20880 ( \20900 , \20897 , \20899 );
buf \U$20881 ( \20901 , \18416 );
buf \U$20882 ( \20902 , RIc0d80c8_23);
buf \U$20883 ( \20903 , RIc0da648_103);
xor \U$20884 ( \20904 , \20902 , \20903 );
buf \U$20885 ( \20905 , \20904 );
buf \U$20886 ( \20906 , \20905 );
nand \U$20887 ( \20907 , \20901 , \20906 );
buf \U$20888 ( \20908 , \20907 );
buf \U$20889 ( \20909 , \20908 );
nand \U$20890 ( \20910 , \20900 , \20909 );
buf \U$20891 ( \20911 , \20910 );
buf \U$20892 ( \20912 , \20911 );
not \U$20893 ( \20913 , \20912 );
buf \U$20894 ( \20914 , \15658 );
not \U$20895 ( \20915 , \20914 );
buf \U$20896 ( \20916 , \12736 );
not \U$20897 ( \20917 , \20916 );
or \U$20898 ( \20918 , \20915 , \20917 );
buf \U$20899 ( \20919 , \12744 );
buf \U$20900 ( \20920 , RIc0d7fd8_21);
buf \U$20901 ( \20921 , RIc0da738_105);
xor \U$20902 ( \20922 , \20920 , \20921 );
buf \U$20903 ( \20923 , \20922 );
buf \U$20904 ( \20924 , \20923 );
nand \U$20905 ( \20925 , \20919 , \20924 );
buf \U$20906 ( \20926 , \20925 );
buf \U$20907 ( \20927 , \20926 );
nand \U$20908 ( \20928 , \20918 , \20927 );
buf \U$20909 ( \20929 , \20928 );
buf \U$20910 ( \20930 , \20929 );
not \U$20911 ( \20931 , \20930 );
buf \U$20912 ( \20932 , \20931 );
buf \U$20913 ( \20933 , \20932 );
not \U$20914 ( \20934 , \20933 );
or \U$20915 ( \20935 , \20913 , \20934 );
buf \U$20916 ( \20936 , \20932 );
buf \U$20917 ( \20937 , \20911 );
or \U$20918 ( \20938 , \20936 , \20937 );
nand \U$20919 ( \20939 , \20935 , \20938 );
buf \U$20920 ( \20940 , \20939 );
buf \U$20921 ( \20941 , \20940 );
buf \U$20922 ( \20942 , \4527 );
buf \U$20923 ( \20943 , \19076 );
and \U$20924 ( \20944 , \20942 , \20943 );
buf \U$20925 ( \20945 , RIc0d8848_39);
buf \U$20926 ( \20946 , RIc0d9ec8_87);
xor \U$20927 ( \20947 , \20945 , \20946 );
buf \U$20928 ( \20948 , \20947 );
buf \U$20929 ( \20949 , \20948 );
not \U$20930 ( \20950 , \20949 );
buf \U$20931 ( \20951 , \634 );
nor \U$20932 ( \20952 , \20950 , \20951 );
buf \U$20933 ( \20953 , \20952 );
buf \U$20934 ( \20954 , \20953 );
nor \U$20935 ( \20955 , \20944 , \20954 );
buf \U$20936 ( \20956 , \20955 );
buf \U$20937 ( \20957 , \20956 );
and \U$20938 ( \20958 , \20941 , \20957 );
not \U$20939 ( \20959 , \20941 );
buf \U$20940 ( \20960 , \20956 );
not \U$20941 ( \20961 , \20960 );
buf \U$20942 ( \20962 , \20961 );
buf \U$20943 ( \20963 , \20962 );
and \U$20944 ( \20964 , \20959 , \20963 );
nor \U$20945 ( \20965 , \20958 , \20964 );
buf \U$20946 ( \20966 , \20965 );
buf \U$20947 ( \20967 , \20966 );
and \U$20948 ( \20968 , \20895 , \20967 );
not \U$20949 ( \20969 , \20895 );
buf \U$20950 ( \20970 , \20966 );
not \U$20951 ( \20971 , \20970 );
buf \U$20952 ( \20972 , \20971 );
buf \U$20953 ( \20973 , \20972 );
and \U$20954 ( \20974 , \20969 , \20973 );
nor \U$20955 ( \20975 , \20968 , \20974 );
buf \U$20956 ( \20976 , \20975 );
buf \U$20957 ( \20977 , \20976 );
not \U$20958 ( \20978 , \20977 );
or \U$20959 ( \20979 , \20778 , \20978 );
buf \U$20960 ( \20980 , \20976 );
buf \U$20961 ( \20981 , \20776 );
or \U$20962 ( \20982 , \20980 , \20981 );
nand \U$20963 ( \20983 , \20979 , \20982 );
buf \U$20964 ( \20984 , \20983 );
buf \U$20965 ( \20985 , \20984 );
and \U$20966 ( \20986 , \12800 , \12801 );
buf \U$20967 ( \20987 , \20986 );
buf \U$20968 ( \20988 , \20987 );
buf \U$20969 ( \20989 , \15468 );
not \U$20970 ( \20990 , \20989 );
buf \U$20971 ( \20991 , \12676 );
not \U$20972 ( \20992 , \20991 );
or \U$20973 ( \20993 , \20990 , \20992 );
buf \U$20974 ( \20994 , \12683 );
buf \U$20975 ( \20995 , RIc0d8fc8_55);
buf \U$20976 ( \20996 , RIc0d9748_71);
xor \U$20977 ( \20997 , \20995 , \20996 );
buf \U$20978 ( \20998 , \20997 );
buf \U$20979 ( \20999 , \20998 );
nand \U$20980 ( \21000 , \20994 , \20999 );
buf \U$20981 ( \21001 , \21000 );
buf \U$20982 ( \21002 , \21001 );
nand \U$20983 ( \21003 , \20993 , \21002 );
buf \U$20984 ( \21004 , \21003 );
buf \U$20985 ( \21005 , \21004 );
xor \U$20986 ( \21006 , \20988 , \21005 );
buf \U$20987 ( \21007 , \15353 );
not \U$20988 ( \21008 , \21007 );
buf \U$20989 ( \21009 , \13181 );
not \U$20990 ( \21010 , \21009 );
or \U$20991 ( \21011 , \21008 , \21010 );
buf \U$20992 ( \21012 , \13005 );
buf \U$20993 ( \21013 , RIc0d7948_7);
buf \U$20994 ( \21014 , RIc0dadc8_119);
xor \U$20995 ( \21015 , \21013 , \21014 );
buf \U$20996 ( \21016 , \21015 );
buf \U$20997 ( \21017 , \21016 );
nand \U$20998 ( \21018 , \21012 , \21017 );
buf \U$20999 ( \21019 , \21018 );
buf \U$21000 ( \21020 , \21019 );
nand \U$21001 ( \21021 , \21011 , \21020 );
buf \U$21002 ( \21022 , \21021 );
buf \U$21003 ( \21023 , \21022 );
xnor \U$21004 ( \21024 , \21006 , \21023 );
buf \U$21005 ( \21025 , \21024 );
buf \U$21006 ( \21026 , \21025 );
not \U$21007 ( \21027 , \21026 );
buf \U$21008 ( \21028 , \15123 );
not \U$21009 ( \21029 , \21028 );
buf \U$21010 ( \21030 , \2899 );
not \U$21011 ( \21031 , \21030 );
or \U$21012 ( \21032 , \21029 , \21031 );
buf \U$21013 ( \21033 , \686 );
buf \U$21014 ( \21034 , RIc0d91a8_59);
buf \U$21015 ( \21035 , RIc0d9568_67);
xor \U$21016 ( \21036 , \21034 , \21035 );
buf \U$21017 ( \21037 , \21036 );
buf \U$21018 ( \21038 , \21037 );
nand \U$21019 ( \21039 , \21033 , \21038 );
buf \U$21020 ( \21040 , \21039 );
buf \U$21021 ( \21041 , \21040 );
nand \U$21022 ( \21042 , \21032 , \21041 );
buf \U$21023 ( \21043 , \21042 );
buf \U$21024 ( \21044 , \21043 );
not \U$21025 ( \21045 , \21044 );
buf \U$21026 ( \21046 , \15848 );
not \U$21027 ( \21047 , \21046 );
buf \U$21028 ( \21048 , \12361 );
not \U$21029 ( \21049 , \21048 );
or \U$21030 ( \21050 , \21047 , \21049 );
buf \U$21031 ( \21051 , \402 );
buf \U$21032 ( \21052 , RIc0d8c08_47);
buf \U$21033 ( \21053 , RIc0d9b08_79);
xor \U$21034 ( \21054 , \21052 , \21053 );
buf \U$21035 ( \21055 , \21054 );
buf \U$21036 ( \21056 , \21055 );
nand \U$21037 ( \21057 , \21051 , \21056 );
buf \U$21038 ( \21058 , \21057 );
buf \U$21039 ( \21059 , \21058 );
nand \U$21040 ( \21060 , \21050 , \21059 );
buf \U$21041 ( \21061 , \21060 );
buf \U$21042 ( \21062 , \21061 );
not \U$21043 ( \21063 , \21062 );
buf \U$21044 ( \21064 , \21063 );
buf \U$21045 ( \21065 , \21064 );
not \U$21046 ( \21066 , \21065 );
or \U$21047 ( \21067 , \21045 , \21066 );
buf \U$21048 ( \21068 , \21043 );
not \U$21049 ( \21069 , \21068 );
buf \U$21050 ( \21070 , \21069 );
buf \U$21051 ( \21071 , \21070 );
buf \U$21052 ( \21072 , \21061 );
nand \U$21053 ( \21073 , \21071 , \21072 );
buf \U$21054 ( \21074 , \21073 );
buf \U$21055 ( \21075 , \21074 );
nand \U$21056 ( \21076 , \21067 , \21075 );
buf \U$21057 ( \21077 , \21076 );
buf \U$21058 ( \21078 , \21077 );
buf \U$21059 ( \21079 , \15337 );
not \U$21060 ( \21080 , \21079 );
buf \U$21061 ( \21081 , \2941 );
not \U$21062 ( \21082 , \21081 );
or \U$21063 ( \21083 , \21080 , \21082 );
buf \U$21064 ( \21084 , \2070 );
buf \U$21065 ( \21085 , RIc0da378_97);
buf \U$21066 ( \21086 , RIc0d8398_29);
xor \U$21067 ( \21087 , \21085 , \21086 );
buf \U$21068 ( \21088 , \21087 );
buf \U$21069 ( \21089 , \21088 );
nand \U$21070 ( \21090 , \21084 , \21089 );
buf \U$21071 ( \21091 , \21090 );
buf \U$21072 ( \21092 , \21091 );
nand \U$21073 ( \21093 , \21083 , \21092 );
buf \U$21074 ( \21094 , \21093 );
buf \U$21075 ( \21095 , \21094 );
not \U$21076 ( \21096 , \21095 );
buf \U$21077 ( \21097 , \21096 );
buf \U$21078 ( \21098 , \21097 );
and \U$21079 ( \21099 , \21078 , \21098 );
not \U$21080 ( \21100 , \21078 );
buf \U$21081 ( \21101 , \21094 );
and \U$21082 ( \21102 , \21100 , \21101 );
nor \U$21083 ( \21103 , \21099 , \21102 );
buf \U$21084 ( \21104 , \21103 );
buf \U$21085 ( \21105 , \21104 );
not \U$21086 ( \21106 , \21105 );
buf \U$21087 ( \21107 , \21106 );
buf \U$21088 ( \21108 , \21107 );
not \U$21089 ( \21109 , \21108 );
or \U$21090 ( \21110 , \21027 , \21109 );
buf \U$21091 ( \21111 , \21104 );
buf \U$21092 ( \21112 , \21025 );
not \U$21093 ( \21113 , \21112 );
buf \U$21094 ( \21114 , \21113 );
buf \U$21095 ( \21115 , \21114 );
nand \U$21096 ( \21116 , \21111 , \21115 );
buf \U$21097 ( \21117 , \21116 );
buf \U$21098 ( \21118 , \21117 );
nand \U$21099 ( \21119 , \21110 , \21118 );
buf \U$21100 ( \21120 , \21119 );
buf \U$21101 ( \21121 , \21120 );
buf \U$21102 ( \21122 , \15798 );
not \U$21103 ( \21123 , \21122 );
buf \U$21104 ( \21124 , \16914 );
not \U$21105 ( \21125 , \21124 );
or \U$21106 ( \21126 , \21123 , \21125 );
buf \U$21107 ( \21127 , \15793 );
buf \U$21108 ( \21128 , RIc0d7678_1);
buf \U$21109 ( \21129 , RIc0db098_125);
xor \U$21110 ( \21130 , \21128 , \21129 );
buf \U$21111 ( \21131 , \21130 );
buf \U$21112 ( \21132 , \21131 );
nand \U$21113 ( \21133 , \21127 , \21132 );
buf \U$21114 ( \21134 , \21133 );
buf \U$21115 ( \21135 , \21134 );
nand \U$21116 ( \21136 , \21126 , \21135 );
buf \U$21117 ( \21137 , \21136 );
buf \U$21118 ( \21138 , \15933 );
not \U$21119 ( \21139 , \21138 );
buf \U$21120 ( \21140 , \14684 );
not \U$21121 ( \21141 , \21140 );
or \U$21122 ( \21142 , \21139 , \21141 );
buf \U$21123 ( \21143 , \12303 );
buf \U$21124 ( \21144 , RIc0d7b28_11);
buf \U$21125 ( \21145 , RIc0dabe8_115);
xor \U$21126 ( \21146 , \21144 , \21145 );
buf \U$21127 ( \21147 , \21146 );
buf \U$21128 ( \21148 , \21147 );
nand \U$21129 ( \21149 , \21143 , \21148 );
buf \U$21130 ( \21150 , \21149 );
buf \U$21131 ( \21151 , \21150 );
nand \U$21132 ( \21152 , \21142 , \21151 );
buf \U$21133 ( \21153 , \21152 );
xor \U$21134 ( \21154 , \21137 , \21153 );
buf \U$21135 ( \21155 , \21154 );
buf \U$21136 ( \21156 , \15536 );
not \U$21137 ( \21157 , \21156 );
buf \U$21138 ( \21158 , \13143 );
nor \U$21139 ( \21159 , \21157 , \21158 );
buf \U$21140 ( \21160 , \21159 );
buf \U$21141 ( \21161 , \21160 );
buf \U$21142 ( \21162 , \16559 );
xor \U$21143 ( \21163 , RIc0dacd8_117, RIc0d7a38_9);
buf \U$21144 ( \21164 , \21163 );
and \U$21145 ( \21165 , \21162 , \21164 );
buf \U$21146 ( \21166 , \21165 );
buf \U$21147 ( \21167 , \21166 );
nor \U$21148 ( \21168 , \21161 , \21167 );
buf \U$21149 ( \21169 , \21168 );
buf \U$21150 ( \21170 , \21169 );
not \U$21151 ( \21171 , \21170 );
buf \U$21152 ( \21172 , \21171 );
buf \U$21153 ( \21173 , \21172 );
and \U$21154 ( \21174 , \21155 , \21173 );
not \U$21155 ( \21175 , \21155 );
buf \U$21156 ( \21176 , \21169 );
and \U$21157 ( \21177 , \21175 , \21176 );
nor \U$21158 ( \21178 , \21174 , \21177 );
buf \U$21159 ( \21179 , \21178 );
buf \U$21160 ( \21180 , \21179 );
not \U$21161 ( \21181 , \21180 );
buf \U$21162 ( \21182 , \21181 );
buf \U$21163 ( \21183 , \21182 );
and \U$21164 ( \21184 , \21121 , \21183 );
not \U$21165 ( \21185 , \21121 );
buf \U$21166 ( \21186 , \21179 );
and \U$21167 ( \21187 , \21185 , \21186 );
nor \U$21168 ( \21188 , \21184 , \21187 );
buf \U$21169 ( \21189 , \21188 );
buf \U$21170 ( \21190 , \21189 );
not \U$21171 ( \21191 , \21190 );
buf \U$21172 ( \21192 , \21191 );
buf \U$21173 ( \21193 , \21192 );
and \U$21174 ( \21194 , \20985 , \21193 );
not \U$21175 ( \21195 , \20985 );
buf \U$21176 ( \21196 , \21189 );
and \U$21177 ( \21197 , \21195 , \21196 );
nor \U$21178 ( \21198 , \21194 , \21197 );
buf \U$21179 ( \21199 , \21198 );
buf \U$21180 ( \21200 , \19179 );
not \U$21181 ( \21201 , \21200 );
buf \U$21182 ( \21202 , \19170 );
not \U$21183 ( \21203 , \21202 );
or \U$21184 ( \21204 , \21201 , \21203 );
buf \U$21185 ( \21205 , \19182 );
not \U$21186 ( \21206 , \21205 );
buf \U$21187 ( \21207 , \19173 );
not \U$21188 ( \21208 , \21207 );
or \U$21189 ( \21209 , \21206 , \21208 );
buf \U$21190 ( \21210 , \19236 );
nand \U$21191 ( \21211 , \21209 , \21210 );
buf \U$21192 ( \21212 , \21211 );
buf \U$21193 ( \21213 , \21212 );
nand \U$21194 ( \21214 , \21204 , \21213 );
buf \U$21195 ( \21215 , \21214 );
xor \U$21196 ( \21216 , \21199 , \21215 );
xor \U$21197 ( \21217 , \18941 , \19041 );
and \U$21198 ( \21218 , \21217 , \19150 );
and \U$21199 ( \21219 , \18941 , \19041 );
or \U$21200 ( \21220 , \21218 , \21219 );
buf \U$21201 ( \21221 , \21220 );
xnor \U$21202 ( \21222 , \21216 , \21221 );
buf \U$21203 ( \21223 , \21222 );
xor \U$21204 ( \21224 , \20606 , \21223 );
buf \U$21205 ( \21225 , \21224 );
buf \U$21206 ( \21226 , \21225 );
xor \U$21207 ( \21227 , \18847 , \19277 );
and \U$21208 ( \21228 , \21227 , \19298 );
and \U$21209 ( \21229 , \18847 , \19277 );
or \U$21210 ( \21230 , \21228 , \21229 );
buf \U$21211 ( \21231 , \21230 );
buf \U$21212 ( \21232 , \21231 );
not \U$21213 ( \21233 , \21232 );
buf \U$21214 ( \21234 , \21233 );
buf \U$21215 ( \21235 , \21234 );
xor \U$21216 ( \21236 , \21226 , \21235 );
buf \U$21217 ( \21237 , \19246 );
not \U$21218 ( \21238 , \21237 );
buf \U$21219 ( \21239 , \21238 );
and \U$21220 ( \21240 , \19152 , \21239 );
buf \U$21221 ( \21241 , \19152 );
not \U$21222 ( \21242 , \21241 );
buf \U$21223 ( \21243 , \21242 );
buf \U$21224 ( \21244 , \21243 );
buf \U$21225 ( \21245 , \19246 );
nand \U$21226 ( \21246 , \21244 , \21245 );
buf \U$21227 ( \21247 , \21246 );
and \U$21228 ( \21248 , \21247 , \19273 );
nor \U$21229 ( \21249 , \21240 , \21248 );
buf \U$21230 ( \21250 , \21249 );
buf \U$21231 ( \21251 , \15293 );
not \U$21232 ( \21252 , \21251 );
buf \U$21233 ( \21253 , \15277 );
not \U$21234 ( \21254 , \21253 );
or \U$21235 ( \21255 , \21252 , \21254 );
buf \U$21236 ( \21256 , \15293 );
buf \U$21237 ( \21257 , \15277 );
or \U$21238 ( \21258 , \21256 , \21257 );
buf \U$21239 ( \21259 , \15194 );
nand \U$21240 ( \21260 , \21258 , \21259 );
buf \U$21241 ( \21261 , \21260 );
buf \U$21242 ( \21262 , \21261 );
nand \U$21243 ( \21263 , \21255 , \21262 );
buf \U$21244 ( \21264 , \21263 );
xor \U$21245 ( \21265 , \19084 , \19090 );
and \U$21246 ( \21266 , \21265 , \19147 );
and \U$21247 ( \21267 , \19084 , \19090 );
or \U$21248 ( \21268 , \21266 , \21267 );
buf \U$21249 ( \21269 , \21268 );
xor \U$21250 ( \21270 , \18947 , \18995 );
and \U$21251 ( \21271 , \21270 , \19038 );
and \U$21252 ( \21272 , \18947 , \18995 );
or \U$21253 ( \21273 , \21271 , \21272 );
buf \U$21254 ( \21274 , \21273 );
xor \U$21255 ( \21275 , \21269 , \21274 );
buf \U$21256 ( \21276 , RIc0db188_127);
not \U$21257 ( \21277 , \21276 );
buf \U$21258 ( \21278 , \21277 );
buf \U$21259 ( \21279 , \21278 );
buf \U$21260 ( \21280 , \15831 );
not \U$21261 ( \21281 , \21280 );
buf \U$21262 ( \21282 , \951 );
not \U$21263 ( \21283 , \21282 );
or \U$21264 ( \21284 , \21281 , \21283 );
buf \U$21265 ( \21285 , \2960 );
buf \U$21266 ( \21286 , RIc0d8938_41);
buf \U$21267 ( \21287 , RIc0d9dd8_85);
xor \U$21268 ( \21288 , \21286 , \21287 );
buf \U$21269 ( \21289 , \21288 );
buf \U$21270 ( \21290 , \21289 );
nand \U$21271 ( \21291 , \21285 , \21290 );
buf \U$21272 ( \21292 , \21291 );
buf \U$21273 ( \21293 , \21292 );
nand \U$21274 ( \21294 , \21284 , \21293 );
buf \U$21275 ( \21295 , \21294 );
buf \U$21276 ( \21296 , \21295 );
xor \U$21277 ( \21297 , \21279 , \21296 );
buf \U$21278 ( \21298 , \19049 );
not \U$21279 ( \21299 , \21298 );
buf \U$21280 ( \21300 , \14982 );
not \U$21281 ( \21301 , \21300 );
or \U$21282 ( \21302 , \21299 , \21301 );
buf \U$21283 ( \21303 , \16692 );
xor \U$21284 ( \21304 , RIc0dafa8_123, RIc0d7768_3);
buf \U$21285 ( \21305 , \21304 );
nand \U$21286 ( \21306 , \21303 , \21305 );
buf \U$21287 ( \21307 , \21306 );
buf \U$21288 ( \21308 , \21307 );
nand \U$21289 ( \21309 , \21302 , \21308 );
buf \U$21290 ( \21310 , \21309 );
buf \U$21291 ( \21311 , \21310 );
not \U$21292 ( \21312 , \21311 );
buf \U$21293 ( \21313 , \21312 );
buf \U$21294 ( \21314 , \21313 );
xor \U$21295 ( \21315 , \21297 , \21314 );
buf \U$21296 ( \21316 , \21315 );
buf \U$21297 ( \21317 , \21316 );
xor \U$21298 ( \21318 , \18999 , \19016 );
and \U$21299 ( \21319 , \21318 , \19035 );
and \U$21300 ( \21320 , \18999 , \19016 );
or \U$21301 ( \21321 , \21319 , \21320 );
buf \U$21302 ( \21322 , \21321 );
buf \U$21303 ( \21323 , \21322 );
xor \U$21304 ( \21324 , \21317 , \21323 );
xor \U$21305 ( \21325 , \15040 , \15049 );
and \U$21306 ( \21326 , \21325 , \15056 );
and \U$21307 ( \21327 , \15040 , \15049 );
or \U$21308 ( \21328 , \21326 , \21327 );
buf \U$21309 ( \21329 , \21328 );
buf \U$21310 ( \21330 , \21329 );
xor \U$21311 ( \21331 , \21324 , \21330 );
buf \U$21312 ( \21332 , \21331 );
xnor \U$21313 ( \21333 , \21275 , \21332 );
and \U$21314 ( \21334 , \21264 , \21333 );
not \U$21315 ( \21335 , \21264 );
not \U$21316 ( \21336 , \21333 );
and \U$21317 ( \21337 , \21335 , \21336 );
nor \U$21318 ( \21338 , \21334 , \21337 );
buf \U$21319 ( \21339 , \15267 );
not \U$21320 ( \21340 , \21339 );
buf \U$21321 ( \21341 , \15238 );
not \U$21322 ( \21342 , \21341 );
or \U$21323 ( \21343 , \21340 , \21342 );
buf \U$21324 ( \21344 , \15241 );
not \U$21325 ( \21345 , \21344 );
buf \U$21326 ( \21346 , \15273 );
not \U$21327 ( \21347 , \21346 );
or \U$21328 ( \21348 , \21345 , \21347 );
buf \U$21329 ( \21349 , \15214 );
nand \U$21330 ( \21350 , \21348 , \21349 );
buf \U$21331 ( \21351 , \21350 );
buf \U$21332 ( \21352 , \21351 );
nand \U$21333 ( \21353 , \21343 , \21352 );
buf \U$21334 ( \21354 , \21353 );
buf \U$21335 ( \21355 , \21354 );
not \U$21336 ( \21356 , \21355 );
not \U$21337 ( \21357 , \15138 );
not \U$21338 ( \21358 , \15187 );
or \U$21339 ( \21359 , \21357 , \21358 );
not \U$21340 ( \21360 , \15133 );
not \U$21341 ( \21361 , \15184 );
or \U$21342 ( \21362 , \21360 , \21361 );
nand \U$21343 ( \21363 , \21362 , \15058 );
nand \U$21344 ( \21364 , \21359 , \21363 );
buf \U$21345 ( \21365 , \21364 );
not \U$21346 ( \21366 , \21365 );
buf \U$21347 ( \21367 , \21366 );
buf \U$21348 ( \21368 , \21367 );
not \U$21349 ( \21369 , \21368 );
or \U$21350 ( \21370 , \21356 , \21369 );
buf \U$21351 ( \21371 , \21367 );
buf \U$21352 ( \21372 , \21354 );
or \U$21353 ( \21373 , \21371 , \21372 );
nand \U$21354 ( \21374 , \21370 , \21373 );
buf \U$21355 ( \21375 , \21374 );
buf \U$21356 ( \21376 , \21375 );
buf \U$21357 ( \21377 , \15145 );
not \U$21358 ( \21378 , \21377 );
buf \U$21359 ( \21379 , \15173 );
not \U$21360 ( \21380 , \21379 );
or \U$21361 ( \21381 , \21378 , \21380 );
buf \U$21362 ( \21382 , \15173 );
buf \U$21363 ( \21383 , \15145 );
or \U$21364 ( \21384 , \21382 , \21383 );
buf \U$21365 ( \21385 , \15155 );
nand \U$21366 ( \21386 , \21384 , \21385 );
buf \U$21367 ( \21387 , \21386 );
buf \U$21368 ( \21388 , \21387 );
nand \U$21369 ( \21389 , \21381 , \21388 );
buf \U$21370 ( \21390 , \21389 );
buf \U$21371 ( \21391 , \21390 );
buf \U$21372 ( \21392 , \15761 );
not \U$21373 ( \21393 , \21392 );
buf \U$21374 ( \21394 , \15782 );
not \U$21375 ( \21395 , \21394 );
or \U$21376 ( \21396 , \21393 , \21395 );
buf \U$21377 ( \21397 , \15804 );
nand \U$21378 ( \21398 , \21396 , \21397 );
buf \U$21379 ( \21399 , \21398 );
buf \U$21380 ( \21400 , \21399 );
buf \U$21381 ( \21401 , \15779 );
buf \U$21382 ( \21402 , \15758 );
nand \U$21383 ( \21403 , \21401 , \21402 );
buf \U$21384 ( \21404 , \21403 );
buf \U$21385 ( \21405 , \21404 );
nand \U$21386 ( \21406 , \21400 , \21405 );
buf \U$21387 ( \21407 , \21406 );
buf \U$21388 ( \21408 , \21407 );
buf \U$21389 ( \21409 , \15722 );
not \U$21390 ( \21410 , \21409 );
buf \U$21391 ( \21411 , \15692 );
not \U$21392 ( \21412 , \21411 );
or \U$21393 ( \21413 , \21410 , \21412 );
buf \U$21394 ( \21414 , \15692 );
buf \U$21395 ( \21415 , \15722 );
or \U$21396 ( \21416 , \21414 , \21415 );
buf \U$21397 ( \21417 , \15708 );
nand \U$21398 ( \21418 , \21416 , \21417 );
buf \U$21399 ( \21419 , \21418 );
buf \U$21400 ( \21420 , \21419 );
nand \U$21401 ( \21421 , \21413 , \21420 );
buf \U$21402 ( \21422 , \21421 );
buf \U$21403 ( \21423 , \21422 );
xor \U$21404 ( \21424 , \21408 , \21423 );
buf \U$21405 ( \21425 , \15440 );
not \U$21406 ( \21426 , \21425 );
buf \U$21407 ( \21427 , \1182 );
not \U$21408 ( \21428 , \21427 );
or \U$21409 ( \21429 , \21426 , \21428 );
buf \U$21410 ( \21430 , \1588 );
buf \U$21411 ( \21431 , RIc0d8cf8_49);
buf \U$21412 ( \21432 , RIc0d9a18_77);
xor \U$21413 ( \21433 , \21431 , \21432 );
buf \U$21414 ( \21434 , \21433 );
buf \U$21415 ( \21435 , \21434 );
nand \U$21416 ( \21436 , \21430 , \21435 );
buf \U$21417 ( \21437 , \21436 );
buf \U$21418 ( \21438 , \21437 );
nand \U$21419 ( \21439 , \21429 , \21438 );
buf \U$21420 ( \21440 , \21439 );
buf \U$21421 ( \21441 , \21440 );
buf \U$21422 ( \21442 , \15716 );
not \U$21423 ( \21443 , \21442 );
buf \U$21424 ( \21444 , \12442 );
not \U$21425 ( \21445 , \21444 );
or \U$21426 ( \21446 , \21443 , \21445 );
buf \U$21427 ( \21447 , \791 );
xor \U$21428 ( \21448 , RIc0d9838_73, RIc0d8ed8_53);
buf \U$21429 ( \21449 , \21448 );
nand \U$21430 ( \21450 , \21447 , \21449 );
buf \U$21431 ( \21451 , \21450 );
buf \U$21432 ( \21452 , \21451 );
nand \U$21433 ( \21453 , \21446 , \21452 );
buf \U$21434 ( \21454 , \21453 );
buf \U$21435 ( \21455 , \21454 );
xor \U$21436 ( \21456 , \21441 , \21455 );
buf \U$21437 ( \21457 , \19062 );
not \U$21438 ( \21458 , \21457 );
buf \U$21439 ( \21459 , \2207 );
not \U$21440 ( \21460 , \21459 );
buf \U$21441 ( \21461 , \21460 );
buf \U$21442 ( \21462 , \21461 );
not \U$21443 ( \21463 , \21462 );
or \U$21444 ( \21464 , \21458 , \21463 );
buf \U$21445 ( \21465 , \16750 );
buf \U$21446 ( \21466 , RIc0da468_99);
buf \U$21447 ( \21467 , RIc0d82a8_27);
xor \U$21448 ( \21468 , \21466 , \21467 );
buf \U$21449 ( \21469 , \21468 );
buf \U$21450 ( \21470 , \21469 );
nand \U$21451 ( \21471 , \21465 , \21470 );
buf \U$21452 ( \21472 , \21471 );
buf \U$21453 ( \21473 , \21472 );
nand \U$21454 ( \21474 , \21464 , \21473 );
buf \U$21455 ( \21475 , \21474 );
buf \U$21456 ( \21476 , \21475 );
xor \U$21457 ( \21477 , \21456 , \21476 );
buf \U$21458 ( \21478 , \21477 );
buf \U$21459 ( \21479 , \21478 );
xor \U$21460 ( \21480 , \21424 , \21479 );
buf \U$21461 ( \21481 , \21480 );
buf \U$21462 ( \21482 , \21481 );
xor \U$21463 ( \21483 , \21391 , \21482 );
not \U$21464 ( \21484 , \15896 );
not \U$21465 ( \21485 , \15940 );
or \U$21466 ( \21486 , \21484 , \21485 );
not \U$21467 ( \21487 , \15937 );
not \U$21468 ( \21488 , \15899 );
or \U$21469 ( \21489 , \21487 , \21488 );
nand \U$21470 ( \21490 , \21489 , \15920 );
nand \U$21471 ( \21491 , \21486 , \21490 );
buf \U$21472 ( \21492 , \21491 );
xor \U$21473 ( \21493 , \15475 , \15492 );
and \U$21474 ( \21494 , \21493 , \15512 );
and \U$21475 ( \21495 , \15475 , \15492 );
or \U$21476 ( \21496 , \21494 , \21495 );
buf \U$21477 ( \21497 , \21496 );
buf \U$21478 ( \21498 , \21497 );
xor \U$21479 ( \21499 , \21492 , \21498 );
xor \U$21480 ( \21500 , \15838 , \15855 );
and \U$21481 ( \21501 , \21500 , \15876 );
and \U$21482 ( \21502 , \15838 , \15855 );
or \U$21483 ( \21503 , \21501 , \21502 );
buf \U$21484 ( \21504 , \21503 );
buf \U$21485 ( \21505 , \21504 );
xor \U$21486 ( \21506 , \21499 , \21505 );
buf \U$21487 ( \21507 , \21506 );
buf \U$21488 ( \21508 , \21507 );
xnor \U$21489 ( \21509 , \21483 , \21508 );
buf \U$21490 ( \21510 , \21509 );
buf \U$21494 ( \21511 , \21510 );
and \U$21495 ( \21512 , \21376 , \21511 );
not \U$21496 ( \21513 , \21376 );
buf \U$21497 ( \21514 , \21510 );
not \U$21498 ( \21515 , \21514 );
buf \U$21499 ( \21516 , \21515 );
buf \U$21500 ( \21517 , \21516 );
and \U$21501 ( \21518 , \21513 , \21517 );
nor \U$21502 ( \21519 , \21512 , \21518 );
buf \U$21503 ( \21520 , \21519 );
buf \U$21504 ( \21521 , \21520 );
not \U$21505 ( \21522 , \21521 );
buf \U$21506 ( \21523 , \21522 );
buf \U$21509 ( \21524 , \21523 );
xor \U$21510 ( \21525 , \21338 , \21524 );
buf \U$21511 ( \21526 , \21525 );
xor \U$21512 ( \21527 , \21250 , \21526 );
buf \U$21513 ( \21528 , \15027 );
not \U$21514 ( \21529 , \21528 );
buf \U$21515 ( \21530 , \16858 );
nand \U$21516 ( \21531 , \21529 , \21530 );
buf \U$21517 ( \21532 , \21531 );
buf \U$21518 ( \21533 , \21532 );
not \U$21519 ( \21534 , \15304 );
buf \U$21520 ( \21535 , \21534 );
and \U$21521 ( \21536 , \21533 , \21535 );
buf \U$21522 ( \21537 , \16858 );
buf \U$21523 ( \21538 , \15030 );
nor \U$21524 ( \21539 , \21537 , \21538 );
buf \U$21525 ( \21540 , \21539 );
buf \U$21526 ( \21541 , \21540 );
nor \U$21527 ( \21542 , \21536 , \21541 );
buf \U$21528 ( \21543 , \21542 );
buf \U$21529 ( \21544 , \21543 );
xor \U$21530 ( \21545 , \21527 , \21544 );
buf \U$21531 ( \21546 , \21545 );
buf \U$21532 ( \21547 , \21546 );
xor \U$21533 ( \21548 , \21236 , \21547 );
buf \U$21534 ( \21549 , \21548 );
buf \U$21535 ( \21550 , \21549 );
not \U$21536 ( \21551 , \21550 );
buf \U$21537 ( \21552 , \21551 );
buf \U$21538 ( \21553 , \21552 );
xor \U$21539 ( \21554 , \16869 , \18840 );
and \U$21540 ( \21555 , \21554 , \19301 );
and \U$21541 ( \21556 , \16869 , \18840 );
or \U$21542 ( \21557 , \21555 , \21556 );
buf \U$21543 ( \21558 , \21557 );
buf \U$21544 ( \21559 , \21558 );
nand \U$21545 ( \21560 , \21553 , \21559 );
buf \U$21546 ( \21561 , \21560 );
buf \U$21547 ( \21562 , \21561 );
and \U$21548 ( \21563 , \20365 , \21562 );
buf \U$21549 ( \21564 , \21558 );
not \U$21550 ( \21565 , \21564 );
buf \U$21551 ( \21566 , \21549 );
nand \U$21552 ( \21567 , \21565 , \21566 );
buf \U$21553 ( \21568 , \21567 );
buf \U$21554 ( \21569 , \21568 );
not \U$21555 ( \21570 , \21569 );
buf \U$21556 ( \21571 , \21570 );
buf \U$21557 ( \21572 , \21571 );
nor \U$21558 ( \21573 , \21563 , \21572 );
buf \U$21559 ( \21574 , \21573 );
buf \U$21560 ( \21575 , \21574 );
not \U$21561 ( \21576 , \21575 );
buf \U$21562 ( \21577 , \20877 );
not \U$21563 ( \21578 , \21577 );
buf \U$21564 ( \21579 , \12402 );
not \U$21565 ( \21580 , \21579 );
or \U$21566 ( \21581 , \21578 , \21580 );
buf \U$21567 ( \21582 , \14405 );
buf \U$21568 ( \21583 , RIc0d7ba0_12);
buf \U$21569 ( \21584 , RIc0daaf8_113);
xor \U$21570 ( \21585 , \21583 , \21584 );
buf \U$21571 ( \21586 , \21585 );
buf \U$21572 ( \21587 , \21586 );
nand \U$21573 ( \21588 , \21582 , \21587 );
buf \U$21574 ( \21589 , \21588 );
buf \U$21575 ( \21590 , \21589 );
nand \U$21576 ( \21591 , \21581 , \21590 );
buf \U$21577 ( \21592 , \21591 );
buf \U$21578 ( \21593 , \21592 );
buf \U$21579 ( \21594 , \20649 );
not \U$21580 ( \21595 , \21594 );
buf \U$21581 ( \21596 , \13075 );
not \U$21582 ( \21597 , \21596 );
or \U$21583 ( \21598 , \21595 , \21597 );
buf \U$21584 ( \21599 , \1078 );
xor \U$21585 ( \21600 , RIc0d9bf8_81, RIc0d8aa0_44);
buf \U$21586 ( \21601 , \21600 );
nand \U$21587 ( \21602 , \21599 , \21601 );
buf \U$21588 ( \21603 , \21602 );
buf \U$21589 ( \21604 , \21603 );
nand \U$21590 ( \21605 , \21598 , \21604 );
buf \U$21591 ( \21606 , \21605 );
buf \U$21592 ( \21607 , \21606 );
xor \U$21593 ( \21608 , \21593 , \21607 );
buf \U$21594 ( \21609 , \21304 );
not \U$21595 ( \21610 , \21609 );
buf \U$21596 ( \21611 , \14982 );
not \U$21597 ( \21612 , \21611 );
or \U$21598 ( \21613 , \21610 , \21612 );
buf \U$21599 ( \21614 , \16692 );
buf \U$21600 ( \21615 , RIc0d76f0_2);
buf \U$21601 ( \21616 , RIc0dafa8_123);
xor \U$21602 ( \21617 , \21615 , \21616 );
buf \U$21603 ( \21618 , \21617 );
buf \U$21604 ( \21619 , \21618 );
nand \U$21605 ( \21620 , \21614 , \21619 );
buf \U$21606 ( \21621 , \21620 );
buf \U$21607 ( \21622 , \21621 );
nand \U$21608 ( \21623 , \21613 , \21622 );
buf \U$21609 ( \21624 , \21623 );
buf \U$21610 ( \21625 , \21624 );
xor \U$21611 ( \21626 , \21608 , \21625 );
buf \U$21612 ( \21627 , \21626 );
buf \U$21613 ( \21628 , \21627 );
and \U$21614 ( \21629 , \15627 , \15628 );
buf \U$21615 ( \21630 , \21629 );
buf \U$21616 ( \21631 , \21630 );
buf \U$21617 ( \21632 , \20616 );
not \U$21618 ( \21633 , \21632 );
buf \U$21619 ( \21634 , \15995 );
not \U$21620 ( \21635 , \21634 );
or \U$21621 ( \21636 , \21633 , \21635 );
buf \U$21622 ( \21637 , \481 );
buf \U$21623 ( \21638 , RIc0d8500_32);
buf \U$21624 ( \21639 , RIc0da198_93);
xor \U$21625 ( \21640 , \21638 , \21639 );
buf \U$21626 ( \21641 , \21640 );
buf \U$21627 ( \21642 , \21641 );
nand \U$21628 ( \21643 , \21637 , \21642 );
buf \U$21629 ( \21644 , \21643 );
buf \U$21630 ( \21645 , \21644 );
nand \U$21631 ( \21646 , \21636 , \21645 );
buf \U$21632 ( \21647 , \21646 );
buf \U$21633 ( \21648 , \21647 );
xor \U$21634 ( \21649 , \21631 , \21648 );
buf \U$21635 ( \21650 , \20673 );
not \U$21636 ( \21651 , \21650 );
buf \U$21637 ( \21652 , \4691 );
not \U$21638 ( \21653 , \21652 );
or \U$21639 ( \21654 , \21651 , \21653 );
buf \U$21640 ( \21655 , \2592 );
not \U$21641 ( \21656 , \21655 );
buf \U$21642 ( \21657 , \21656 );
buf \U$21643 ( \21658 , \21657 );
xor \U$21644 ( \21659 , RIc0d9658_69, RIc0d9040_56);
buf \U$21645 ( \21660 , \21659 );
nand \U$21646 ( \21661 , \21658 , \21660 );
buf \U$21647 ( \21662 , \21661 );
buf \U$21648 ( \21663 , \21662 );
nand \U$21649 ( \21664 , \21654 , \21663 );
buf \U$21650 ( \21665 , \21664 );
buf \U$21651 ( \21666 , \21665 );
xnor \U$21652 ( \21667 , \21649 , \21666 );
buf \U$21653 ( \21668 , \21667 );
buf \U$21654 ( \21669 , \21668 );
not \U$21655 ( \21670 , \21669 );
buf \U$21656 ( \21671 , \21670 );
buf \U$21657 ( \21672 , \21671 );
or \U$21658 ( \21673 , \21628 , \21672 );
buf \U$21659 ( \21674 , \21147 );
not \U$21660 ( \21675 , \21674 );
buf \U$21661 ( \21676 , \14186 );
not \U$21662 ( \21677 , \21676 );
or \U$21663 ( \21678 , \21675 , \21677 );
buf \U$21664 ( \21679 , \14690 );
buf \U$21665 ( \21680 , RIc0d7ab0_10);
buf \U$21666 ( \21681 , RIc0dabe8_115);
xor \U$21667 ( \21682 , \21680 , \21681 );
buf \U$21668 ( \21683 , \21682 );
buf \U$21669 ( \21684 , \21683 );
nand \U$21670 ( \21685 , \21679 , \21684 );
buf \U$21671 ( \21686 , \21685 );
buf \U$21672 ( \21687 , \21686 );
nand \U$21673 ( \21688 , \21678 , \21687 );
buf \U$21674 ( \21689 , \21688 );
buf \U$21675 ( \21690 , \21055 );
not \U$21676 ( \21691 , \21690 );
buf \U$21677 ( \21692 , \12361 );
not \U$21678 ( \21693 , \21692 );
or \U$21679 ( \21694 , \21691 , \21693 );
buf \U$21680 ( \21695 , \402 );
buf \U$21681 ( \21696 , RIc0d8b90_46);
buf \U$21682 ( \21697 , RIc0d9b08_79);
xor \U$21683 ( \21698 , \21696 , \21697 );
buf \U$21684 ( \21699 , \21698 );
buf \U$21685 ( \21700 , \21699 );
nand \U$21686 ( \21701 , \21695 , \21700 );
buf \U$21687 ( \21702 , \21701 );
buf \U$21688 ( \21703 , \21702 );
nand \U$21689 ( \21704 , \21694 , \21703 );
buf \U$21690 ( \21705 , \21704 );
buf \U$21691 ( \21706 , \21705 );
not \U$21692 ( \21707 , \21706 );
buf \U$21693 ( \21708 , \21707 );
xor \U$21694 ( \21709 , \21689 , \21708 );
buf \U$21695 ( \21710 , \20948 );
not \U$21696 ( \21711 , \21710 );
buf \U$21697 ( \21712 , \14325 );
not \U$21698 ( \21713 , \21712 );
or \U$21699 ( \21714 , \21711 , \21713 );
buf \U$21700 ( \21715 , \816 );
buf \U$21701 ( \21716 , RIc0d87d0_38);
buf \U$21702 ( \21717 , RIc0d9ec8_87);
xor \U$21703 ( \21718 , \21716 , \21717 );
buf \U$21704 ( \21719 , \21718 );
buf \U$21705 ( \21720 , \21719 );
nand \U$21706 ( \21721 , \21715 , \21720 );
buf \U$21707 ( \21722 , \21721 );
buf \U$21708 ( \21723 , \21722 );
nand \U$21709 ( \21724 , \21714 , \21723 );
buf \U$21710 ( \21725 , \21724 );
buf \U$21711 ( \21726 , \21725 );
not \U$21712 ( \21727 , \21726 );
buf \U$21713 ( \21728 , \21727 );
and \U$21714 ( \21729 , \21709 , \21728 );
not \U$21715 ( \21730 , \21709 );
and \U$21716 ( \21731 , \21730 , \21725 );
nor \U$21717 ( \21732 , \21729 , \21731 );
buf \U$21718 ( \21733 , \21732 );
nand \U$21719 ( \21734 , \21673 , \21733 );
buf \U$21720 ( \21735 , \21734 );
buf \U$21721 ( \21736 , \21735 );
buf \U$21722 ( \21737 , \21627 );
buf \U$21723 ( \21738 , \21671 );
nand \U$21724 ( \21739 , \21737 , \21738 );
buf \U$21725 ( \21740 , \21739 );
buf \U$21726 ( \21741 , \21740 );
nand \U$21727 ( \21742 , \21736 , \21741 );
buf \U$21728 ( \21743 , \21742 );
buf \U$21729 ( \21744 , \21743 );
buf \U$21730 ( \21745 , \20690 );
not \U$21731 ( \21746 , \21745 );
buf \U$21732 ( \21747 , \13991 );
not \U$21733 ( \21748 , \21747 );
or \U$21734 ( \21749 , \21746 , \21748 );
buf \U$21735 ( \21750 , \13998 );
buf \U$21736 ( \21751 , RIc0d8d70_50);
buf \U$21737 ( \21752 , RIc0d9928_75);
xor \U$21738 ( \21753 , \21751 , \21752 );
buf \U$21739 ( \21754 , \21753 );
buf \U$21740 ( \21755 , \21754 );
nand \U$21741 ( \21756 , \21750 , \21755 );
buf \U$21742 ( \21757 , \21756 );
buf \U$21743 ( \21758 , \21757 );
nand \U$21744 ( \21759 , \21749 , \21758 );
buf \U$21745 ( \21760 , \21759 );
buf \U$21746 ( \21761 , \21760 );
buf \U$21747 ( \21762 , \20905 );
not \U$21748 ( \21763 , \21762 );
buf \U$21749 ( \21764 , \15397 );
not \U$21750 ( \21765 , \21764 );
or \U$21751 ( \21766 , \21763 , \21765 );
buf \U$21752 ( \21767 , \18416 );
buf \U$21753 ( \21768 , RIc0d8050_22);
buf \U$21754 ( \21769 , RIc0da648_103);
xor \U$21755 ( \21770 , \21768 , \21769 );
buf \U$21756 ( \21771 , \21770 );
buf \U$21757 ( \21772 , \21771 );
nand \U$21758 ( \21773 , \21767 , \21772 );
buf \U$21759 ( \21774 , \21773 );
buf \U$21760 ( \21775 , \21774 );
nand \U$21761 ( \21776 , \21766 , \21775 );
buf \U$21762 ( \21777 , \21776 );
buf \U$21763 ( \21778 , \21777 );
xor \U$21764 ( \21779 , \21761 , \21778 );
buf \U$21765 ( \21780 , \20806 );
not \U$21766 ( \21781 , \21780 );
buf \U$21767 ( \21782 , \3534 );
not \U$21768 ( \21783 , \21782 );
or \U$21769 ( \21784 , \21781 , \21783 );
buf \U$21770 ( \21785 , \16676 );
buf \U$21771 ( \21786 , RIc0da558_101);
buf \U$21772 ( \21787 , RIc0d8140_24);
xor \U$21773 ( \21788 , \21786 , \21787 );
buf \U$21774 ( \21789 , \21788 );
buf \U$21775 ( \21790 , \21789 );
nand \U$21776 ( \21791 , \21785 , \21790 );
buf \U$21777 ( \21792 , \21791 );
buf \U$21778 ( \21793 , \21792 );
nand \U$21779 ( \21794 , \21784 , \21793 );
buf \U$21780 ( \21795 , \21794 );
buf \U$21781 ( \21796 , \21795 );
and \U$21782 ( \21797 , \21779 , \21796 );
and \U$21783 ( \21798 , \21761 , \21778 );
or \U$21784 ( \21799 , \21797 , \21798 );
buf \U$21785 ( \21800 , \21799 );
buf \U$21786 ( \21801 , \21800 );
buf \U$21787 ( \21802 , \20729 );
not \U$21788 ( \21803 , \21802 );
buf \U$21789 ( \21804 , \3780 );
not \U$21790 ( \21805 , \21804 );
or \U$21791 ( \21806 , \21803 , \21805 );
buf \U$21792 ( \21807 , \1229 );
buf \U$21793 ( \21808 , RIc0d9478_65);
buf \U$21794 ( \21809 , RIc0d9220_60);
xor \U$21795 ( \21810 , \21808 , \21809 );
buf \U$21796 ( \21811 , \21810 );
buf \U$21797 ( \21812 , \21811 );
nand \U$21798 ( \21813 , \21807 , \21812 );
buf \U$21799 ( \21814 , \21813 );
buf \U$21800 ( \21815 , \21814 );
nand \U$21801 ( \21816 , \21806 , \21815 );
buf \U$21802 ( \21817 , \21816 );
buf \U$21803 ( \21818 , \21817 );
buf \U$21804 ( \21819 , \21448 );
not \U$21805 ( \21820 , \21819 );
buf \U$21806 ( \21821 , \14075 );
not \U$21807 ( \21822 , \21821 );
or \U$21808 ( \21823 , \21820 , \21822 );
buf \U$21809 ( \21824 , \792 );
buf \U$21810 ( \21825 , RIc0d8e60_52);
buf \U$21811 ( \21826 , RIc0d9838_73);
xor \U$21812 ( \21827 , \21825 , \21826 );
buf \U$21813 ( \21828 , \21827 );
buf \U$21814 ( \21829 , \21828 );
nand \U$21815 ( \21830 , \21824 , \21829 );
buf \U$21816 ( \21831 , \21830 );
buf \U$21817 ( \21832 , \21831 );
nand \U$21818 ( \21833 , \21823 , \21832 );
buf \U$21819 ( \21834 , \21833 );
buf \U$21820 ( \21835 , \21834 );
xor \U$21821 ( \21836 , \21818 , \21835 );
buf \U$21822 ( \21837 , \21131 );
not \U$21823 ( \21838 , \21837 );
buf \U$21824 ( \21839 , \14471 );
not \U$21825 ( \21840 , \21839 );
or \U$21826 ( \21841 , \21838 , \21840 );
buf \U$21827 ( \21842 , \15793 );
buf \U$21828 ( \21843 , RIc0db098_125);
nand \U$21829 ( \21844 , \21842 , \21843 );
buf \U$21830 ( \21845 , \21844 );
buf \U$21831 ( \21846 , \21845 );
nand \U$21832 ( \21847 , \21841 , \21846 );
buf \U$21833 ( \21848 , \21847 );
buf \U$21834 ( \21849 , \21848 );
and \U$21835 ( \21850 , \21836 , \21849 );
and \U$21836 ( \21851 , \21818 , \21835 );
or \U$21837 ( \21852 , \21850 , \21851 );
buf \U$21838 ( \21853 , \21852 );
buf \U$21839 ( \21854 , \21853 );
xor \U$21840 ( \21855 , \21801 , \21854 );
buf \U$21841 ( \21856 , \21037 );
not \U$21842 ( \21857 , \21856 );
buf \U$21843 ( \21858 , \1823 );
not \U$21844 ( \21859 , \21858 );
or \U$21845 ( \21860 , \21857 , \21859 );
buf \U$21846 ( \21861 , \686 );
buf \U$21847 ( \21862 , RIc0d9130_58);
buf \U$21848 ( \21863 , RIc0d9568_67);
xor \U$21849 ( \21864 , \21862 , \21863 );
buf \U$21850 ( \21865 , \21864 );
buf \U$21851 ( \21866 , \21865 );
nand \U$21852 ( \21867 , \21861 , \21866 );
buf \U$21853 ( \21868 , \21867 );
buf \U$21854 ( \21869 , \21868 );
nand \U$21855 ( \21870 , \21860 , \21869 );
buf \U$21856 ( \21871 , \21870 );
buf \U$21857 ( \21872 , \21871 );
buf \U$21858 ( \21873 , \20923 );
not \U$21859 ( \21874 , \21873 );
buf \U$21860 ( \21875 , \15644 );
not \U$21861 ( \21876 , \21875 );
or \U$21862 ( \21877 , \21874 , \21876 );
buf \U$21863 ( \21878 , \15650 );
not \U$21864 ( \21879 , \21878 );
buf \U$21865 ( \21880 , \21879 );
buf \U$21866 ( \21881 , \21880 );
buf \U$21867 ( \21882 , RIc0da738_105);
buf \U$21868 ( \21883 , RIc0d7f60_20);
xor \U$21869 ( \21884 , \21882 , \21883 );
buf \U$21870 ( \21885 , \21884 );
buf \U$21871 ( \21886 , \21885 );
nand \U$21872 ( \21887 , \21881 , \21886 );
buf \U$21873 ( \21888 , \21887 );
buf \U$21874 ( \21889 , \21888 );
nand \U$21875 ( \21890 , \21877 , \21889 );
buf \U$21876 ( \21891 , \21890 );
buf \U$21877 ( \21892 , \21891 );
xor \U$21878 ( \21893 , \21872 , \21892 );
buf \U$21879 ( \21894 , \20746 );
not \U$21880 ( \21895 , \21894 );
buf \U$21881 ( \21896 , \12331 );
not \U$21882 ( \21897 , \21896 );
buf \U$21883 ( \21898 , \21897 );
buf \U$21884 ( \21899 , \21898 );
not \U$21885 ( \21900 , \21899 );
or \U$21886 ( \21901 , \21895 , \21900 );
buf \U$21887 ( \21902 , \16071 );
xor \U$21888 ( \21903 , RIc0da828_107, RIc0d7e70_18);
buf \U$21889 ( \21904 , \21903 );
nand \U$21890 ( \21905 , \21902 , \21904 );
buf \U$21891 ( \21906 , \21905 );
buf \U$21892 ( \21907 , \21906 );
nand \U$21893 ( \21908 , \21901 , \21907 );
buf \U$21894 ( \21909 , \21908 );
buf \U$21895 ( \21910 , \21909 );
and \U$21896 ( \21911 , \21893 , \21910 );
and \U$21897 ( \21912 , \21872 , \21892 );
or \U$21898 ( \21913 , \21911 , \21912 );
buf \U$21899 ( \21914 , \21913 );
buf \U$21900 ( \21915 , \21914 );
xor \U$21901 ( \21916 , \21855 , \21915 );
buf \U$21902 ( \21917 , \21916 );
buf \U$21903 ( \21918 , \21917 );
xor \U$21904 ( \21919 , \21744 , \21918 );
buf \U$21905 ( \21920 , \21434 );
not \U$21906 ( \21921 , \21920 );
buf \U$21907 ( \21922 , \14825 );
not \U$21908 ( \21923 , \21922 );
or \U$21909 ( \21924 , \21921 , \21923 );
buf \U$21910 ( \21925 , \3742 );
buf \U$21911 ( \21926 , RIc0d8c80_48);
buf \U$21912 ( \21927 , RIc0d9a18_77);
xor \U$21913 ( \21928 , \21926 , \21927 );
buf \U$21914 ( \21929 , \21928 );
buf \U$21915 ( \21930 , \21929 );
nand \U$21916 ( \21931 , \21925 , \21930 );
buf \U$21917 ( \21932 , \21931 );
buf \U$21918 ( \21933 , \21932 );
nand \U$21919 ( \21934 , \21924 , \21933 );
buf \U$21920 ( \21935 , \21934 );
buf \U$21921 ( \21936 , \21935 );
buf \U$21922 ( \21937 , \20859 );
not \U$21923 ( \21938 , \21937 );
buf \U$21924 ( \21939 , \14346 );
not \U$21925 ( \21940 , \21939 );
or \U$21926 ( \21941 , \21938 , \21940 );
buf \U$21927 ( \21942 , \18312 );
buf \U$21928 ( \21943 , RIc0d7c90_14);
buf \U$21929 ( \21944 , RIc0daa08_111);
xor \U$21930 ( \21945 , \21943 , \21944 );
buf \U$21931 ( \21946 , \21945 );
buf \U$21932 ( \21947 , \21946 );
nand \U$21933 ( \21948 , \21942 , \21947 );
buf \U$21934 ( \21949 , \21948 );
buf \U$21935 ( \21950 , \21949 );
nand \U$21936 ( \21951 , \21941 , \21950 );
buf \U$21937 ( \21952 , \21951 );
buf \U$21938 ( \21953 , \21952 );
xor \U$21939 ( \21954 , \21936 , \21953 );
buf \U$21940 ( \21955 , \20764 );
not \U$21941 ( \21956 , \21955 );
buf \U$21942 ( \21957 , \14207 );
not \U$21943 ( \21958 , \21957 );
buf \U$21944 ( \21959 , \21958 );
buf \U$21945 ( \21960 , \21959 );
not \U$21946 ( \21961 , \21960 );
or \U$21947 ( \21962 , \21956 , \21961 );
buf \U$21948 ( \21963 , \20211 );
buf \U$21949 ( \21964 , RIc0d7d80_16);
buf \U$21950 ( \21965 , RIc0da918_109);
xor \U$21951 ( \21966 , \21964 , \21965 );
buf \U$21952 ( \21967 , \21966 );
buf \U$21953 ( \21968 , \21967 );
nand \U$21954 ( \21969 , \21963 , \21968 );
buf \U$21955 ( \21970 , \21969 );
buf \U$21956 ( \21971 , \21970 );
nand \U$21957 ( \21972 , \21962 , \21971 );
buf \U$21958 ( \21973 , \21972 );
buf \U$21959 ( \21974 , \21973 );
xor \U$21960 ( \21975 , \21954 , \21974 );
buf \U$21961 ( \21976 , \21975 );
buf \U$21962 ( \21977 , \21976 );
xor \U$21963 ( \21978 , \21872 , \21892 );
xor \U$21964 ( \21979 , \21978 , \21910 );
buf \U$21965 ( \21980 , \21979 );
buf \U$21966 ( \21981 , \21980 );
xor \U$21967 ( \21982 , \21977 , \21981 );
buf \U$21968 ( \21983 , \20708 );
not \U$21969 ( \21984 , \21983 );
buf \U$21970 ( \21985 , \330 );
not \U$21971 ( \21986 , \21985 );
or \U$21972 ( \21987 , \21984 , \21986 );
buf \U$21973 ( \21988 , \14707 );
buf \U$21974 ( \21989 , RIc0d8410_30);
buf \U$21975 ( \21990 , RIc0da288_95);
xor \U$21976 ( \21991 , \21989 , \21990 );
buf \U$21977 ( \21992 , \21991 );
buf \U$21978 ( \21993 , \21992 );
nand \U$21979 ( \21994 , \21988 , \21993 );
buf \U$21980 ( \21995 , \21994 );
buf \U$21981 ( \21996 , \21995 );
nand \U$21982 ( \21997 , \21987 , \21996 );
buf \U$21983 ( \21998 , \21997 );
buf \U$21984 ( \21999 , \21469 );
not \U$21985 ( \22000 , \21999 );
buf \U$21986 ( \22001 , \2470 );
not \U$21987 ( \22002 , \22001 );
or \U$21988 ( \22003 , \22000 , \22002 );
buf \U$21989 ( \22004 , \2199 );
not \U$21990 ( \22005 , \22004 );
buf \U$21991 ( \22006 , \22005 );
buf \U$21992 ( \22007 , \22006 );
buf \U$21993 ( \22008 , RIc0da468_99);
buf \U$21994 ( \22009 , RIc0d8230_26);
xor \U$21995 ( \22010 , \22008 , \22009 );
buf \U$21996 ( \22011 , \22010 );
buf \U$21997 ( \22012 , \22011 );
nand \U$21998 ( \22013 , \22007 , \22012 );
buf \U$21999 ( \22014 , \22013 );
buf \U$22000 ( \22015 , \22014 );
nand \U$22001 ( \22016 , \22003 , \22015 );
buf \U$22002 ( \22017 , \22016 );
xor \U$22003 ( \22018 , \21998 , \22017 );
buf \U$22004 ( \22019 , \20785 );
not \U$22005 ( \22020 , \22019 );
buf \U$22006 ( \22021 , \19487 );
not \U$22007 ( \22022 , \22021 );
or \U$22008 ( \22023 , \22020 , \22022 );
buf \U$22009 ( \22024 , \13314 );
xor \U$22010 ( \22025 , RIc0daeb8_121, RIc0d77e0_4);
buf \U$22011 ( \22026 , \22025 );
nand \U$22012 ( \22027 , \22024 , \22026 );
buf \U$22013 ( \22028 , \22027 );
buf \U$22014 ( \22029 , \22028 );
nand \U$22015 ( \22030 , \22023 , \22029 );
buf \U$22016 ( \22031 , \22030 );
xor \U$22017 ( \22032 , \22018 , \22031 );
buf \U$22018 ( \22033 , \22032 );
and \U$22019 ( \22034 , \21982 , \22033 );
and \U$22020 ( \22035 , \21977 , \21981 );
or \U$22021 ( \22036 , \22034 , \22035 );
buf \U$22022 ( \22037 , \22036 );
buf \U$22023 ( \22038 , \22037 );
xor \U$22024 ( \22039 , \21919 , \22038 );
buf \U$22025 ( \22040 , \22039 );
buf \U$22026 ( \22041 , \22040 );
buf \U$22027 ( \22042 , \20561 );
not \U$22028 ( \22043 , \22042 );
buf \U$22029 ( \22044 , \20550 );
not \U$22030 ( \22045 , \22044 );
or \U$22031 ( \22046 , \22043 , \22045 );
buf \U$22032 ( \22047 , \20561 );
buf \U$22033 ( \22048 , \20550 );
or \U$22034 ( \22049 , \22047 , \22048 );
buf \U$22035 ( \22050 , \20555 );
nand \U$22036 ( \22051 , \22049 , \22050 );
buf \U$22037 ( \22052 , \22051 );
buf \U$22038 ( \22053 , \22052 );
nand \U$22039 ( \22054 , \22046 , \22053 );
buf \U$22040 ( \22055 , \22054 );
buf \U$22041 ( \22056 , \22055 );
buf \U$22042 ( \22057 , \20679 );
not \U$22043 ( \22058 , \22057 );
buf \U$22044 ( \22059 , \20714 );
not \U$22045 ( \22060 , \22059 );
or \U$22046 ( \22061 , \22058 , \22060 );
buf \U$22047 ( \22062 , \20714 );
buf \U$22048 ( \22063 , \20679 );
or \U$22049 ( \22064 , \22062 , \22063 );
buf \U$22050 ( \22065 , \20696 );
nand \U$22051 ( \22066 , \22064 , \22065 );
buf \U$22052 ( \22067 , \22066 );
buf \U$22053 ( \22068 , \22067 );
nand \U$22054 ( \22069 , \22061 , \22068 );
buf \U$22055 ( \22070 , \22069 );
buf \U$22056 ( \22071 , \22070 );
buf \U$22057 ( \22072 , \20638 );
not \U$22058 ( \22073 , \22072 );
buf \U$22059 ( \22074 , \20655 );
not \U$22060 ( \22075 , \22074 );
or \U$22061 ( \22076 , \22073 , \22075 );
buf \U$22062 ( \22077 , \20655 );
buf \U$22063 ( \22078 , \20638 );
or \U$22064 ( \22079 , \22077 , \22078 );
buf \U$22065 ( \22080 , \20622 );
nand \U$22066 ( \22081 , \22079 , \22080 );
buf \U$22067 ( \22082 , \22081 );
buf \U$22068 ( \22083 , \22082 );
nand \U$22069 ( \22084 , \22076 , \22083 );
buf \U$22070 ( \22085 , \22084 );
buf \U$22071 ( \22086 , \22085 );
and \U$22072 ( \22087 , \22071 , \22086 );
not \U$22073 ( \22088 , \22071 );
buf \U$22074 ( \22089 , \22085 );
not \U$22075 ( \22090 , \22089 );
buf \U$22076 ( \22091 , \22090 );
buf \U$22077 ( \22092 , \22091 );
and \U$22078 ( \22093 , \22088 , \22092 );
nor \U$22079 ( \22094 , \22087 , \22093 );
buf \U$22080 ( \22095 , \22094 );
buf \U$22081 ( \22096 , \22095 );
xor \U$22082 ( \22097 , \20849 , \20866 );
and \U$22083 ( \22098 , \22097 , \20884 );
and \U$22084 ( \22099 , \20849 , \20866 );
or \U$22085 ( \22100 , \22098 , \22099 );
buf \U$22086 ( \22101 , \22100 );
buf \U$22087 ( \22102 , \22101 );
xor \U$22088 ( \22103 , \22096 , \22102 );
buf \U$22089 ( \22104 , \22103 );
buf \U$22090 ( \22105 , \22104 );
xor \U$22091 ( \22106 , \22056 , \22105 );
xor \U$22092 ( \22107 , \20663 , \20718 );
and \U$22093 ( \22108 , \22107 , \20774 );
and \U$22094 ( \22109 , \20663 , \20718 );
or \U$22095 ( \22110 , \22108 , \22109 );
buf \U$22096 ( \22111 , \22110 );
buf \U$22097 ( \22112 , \22111 );
and \U$22098 ( \22113 , \22106 , \22112 );
and \U$22099 ( \22114 , \22056 , \22105 );
or \U$22100 ( \22115 , \22113 , \22114 );
buf \U$22101 ( \22116 , \22115 );
buf \U$22102 ( \22117 , \22116 );
and \U$22103 ( \22118 , \22041 , \22117 );
not \U$22104 ( \22119 , \22041 );
buf \U$22105 ( \22120 , \22116 );
not \U$22106 ( \22121 , \22120 );
buf \U$22107 ( \22122 , \22121 );
buf \U$22108 ( \22123 , \22122 );
and \U$22109 ( \22124 , \22119 , \22123 );
nor \U$22110 ( \22125 , \22118 , \22124 );
buf \U$22111 ( \22126 , \22125 );
buf \U$22112 ( \22127 , \22126 );
buf \U$22113 ( \22128 , \20842 );
not \U$22114 ( \22129 , \22128 );
buf \U$22115 ( \22130 , \12254 );
not \U$22116 ( \22131 , \22130 );
or \U$22117 ( \22132 , \22129 , \22131 );
buf \U$22118 ( \22133 , \584 );
buf \U$22119 ( \22134 , RIc0d89b0_42);
buf \U$22120 ( \22135 , RIc0d9ce8_83);
xor \U$22121 ( \22136 , \22134 , \22135 );
buf \U$22122 ( \22137 , \22136 );
buf \U$22123 ( \22138 , \22137 );
nand \U$22124 ( \22139 , \22133 , \22138 );
buf \U$22125 ( \22140 , \22139 );
buf \U$22126 ( \22141 , \22140 );
nand \U$22127 ( \22142 , \22132 , \22141 );
buf \U$22128 ( \22143 , \22142 );
buf \U$22129 ( \22144 , \22143 );
buf \U$22130 ( \22145 , \20823 );
not \U$22131 ( \22146 , \22145 );
buf \U$22132 ( \22147 , \2535 );
not \U$22133 ( \22148 , \22147 );
or \U$22134 ( \22149 , \22146 , \22148 );
buf \U$22135 ( \22150 , \533 );
buf \U$22136 ( \22151 , RIc0d85f0_34);
buf \U$22137 ( \22152 , RIc0da0a8_91);
xor \U$22138 ( \22153 , \22151 , \22152 );
buf \U$22139 ( \22154 , \22153 );
buf \U$22140 ( \22155 , \22154 );
nand \U$22141 ( \22156 , \22150 , \22155 );
buf \U$22142 ( \22157 , \22156 );
buf \U$22143 ( \22158 , \22157 );
nand \U$22144 ( \22159 , \22149 , \22158 );
buf \U$22145 ( \22160 , \22159 );
buf \U$22146 ( \22161 , \22160 );
xor \U$22147 ( \22162 , \22144 , \22161 );
buf \U$22148 ( \22163 , \20632 );
not \U$22149 ( \22164 , \22163 );
buf \U$22150 ( \22165 , \842 );
not \U$22151 ( \22166 , \22165 );
or \U$22152 ( \22167 , \22164 , \22166 );
buf \U$22153 ( \22168 , \846 );
buf \U$22154 ( \22169 , RIc0d9fb8_89);
buf \U$22155 ( \22170 , RIc0d86e0_36);
xor \U$22156 ( \22171 , \22169 , \22170 );
buf \U$22157 ( \22172 , \22171 );
buf \U$22158 ( \22173 , \22172 );
nand \U$22159 ( \22174 , \22168 , \22173 );
buf \U$22160 ( \22175 , \22174 );
buf \U$22161 ( \22176 , \22175 );
nand \U$22162 ( \22177 , \22167 , \22176 );
buf \U$22163 ( \22178 , \22177 );
buf \U$22164 ( \22179 , \22178 );
xor \U$22165 ( \22180 , \22162 , \22179 );
buf \U$22166 ( \22181 , \22180 );
buf \U$22167 ( \22182 , \22181 );
not \U$22168 ( \22183 , \22182 );
buf \U$22169 ( \22184 , \22183 );
buf \U$22170 ( \22185 , \22184 );
not \U$22171 ( \22186 , \22185 );
buf \U$22172 ( \22187 , \20998 );
not \U$22173 ( \22188 , \22187 );
buf \U$22174 ( \22189 , \12676 );
not \U$22175 ( \22190 , \22189 );
or \U$22176 ( \22191 , \22188 , \22190 );
buf \U$22177 ( \22192 , \12683 );
buf \U$22178 ( \22193 , RIc0d8f50_54);
buf \U$22179 ( \22194 , RIc0d9748_71);
xor \U$22180 ( \22195 , \22193 , \22194 );
buf \U$22181 ( \22196 , \22195 );
buf \U$22182 ( \22197 , \22196 );
nand \U$22183 ( \22198 , \22192 , \22197 );
buf \U$22184 ( \22199 , \22198 );
buf \U$22185 ( \22200 , \22199 );
nand \U$22186 ( \22201 , \22191 , \22200 );
buf \U$22187 ( \22202 , \22201 );
buf \U$22188 ( \22203 , \21289 );
not \U$22189 ( \22204 , \22203 );
buf \U$22190 ( \22205 , \1388 );
not \U$22191 ( \22206 , \22205 );
or \U$22192 ( \22207 , \22204 , \22206 );
buf \U$22193 ( \22208 , \1401 );
buf \U$22194 ( \22209 , RIc0d88c0_40);
buf \U$22195 ( \22210 , RIc0d9dd8_85);
xor \U$22196 ( \22211 , \22209 , \22210 );
buf \U$22197 ( \22212 , \22211 );
buf \U$22198 ( \22213 , \22212 );
nand \U$22199 ( \22214 , \22208 , \22213 );
buf \U$22200 ( \22215 , \22214 );
buf \U$22201 ( \22216 , \22215 );
nand \U$22202 ( \22217 , \22207 , \22216 );
buf \U$22203 ( \22218 , \22217 );
xor \U$22204 ( \22219 , \22202 , \22218 );
buf \U$22205 ( \22220 , \21088 );
not \U$22206 ( \22221 , \22220 );
buf \U$22207 ( \22222 , \2941 );
not \U$22208 ( \22223 , \22222 );
or \U$22209 ( \22224 , \22221 , \22223 );
buf \U$22210 ( \22225 , \2070 );
buf \U$22211 ( \22226 , RIc0d8320_28);
buf \U$22212 ( \22227 , RIc0da378_97);
xor \U$22213 ( \22228 , \22226 , \22227 );
buf \U$22214 ( \22229 , \22228 );
buf \U$22215 ( \22230 , \22229 );
nand \U$22216 ( \22231 , \22225 , \22230 );
buf \U$22217 ( \22232 , \22231 );
buf \U$22218 ( \22233 , \22232 );
nand \U$22219 ( \22234 , \22224 , \22233 );
buf \U$22220 ( \22235 , \22234 );
xnor \U$22221 ( \22236 , \22219 , \22235 );
buf \U$22222 ( \22237 , \22236 );
not \U$22223 ( \22238 , \22237 );
buf \U$22224 ( \22239 , \22238 );
buf \U$22225 ( \22240 , \22239 );
not \U$22226 ( \22241 , \22240 );
or \U$22227 ( \22242 , \22186 , \22241 );
buf \U$22228 ( \22243 , \22236 );
buf \U$22229 ( \22244 , \22181 );
nand \U$22230 ( \22245 , \22243 , \22244 );
buf \U$22231 ( \22246 , \22245 );
buf \U$22232 ( \22247 , \22246 );
nand \U$22233 ( \22248 , \22242 , \22247 );
buf \U$22234 ( \22249 , \22248 );
buf \U$22235 ( \22250 , \22249 );
xor \U$22236 ( \22251 , \21279 , \21296 );
and \U$22237 ( \22252 , \22251 , \21314 );
and \U$22238 ( \22253 , \21279 , \21296 );
or \U$22239 ( \22254 , \22252 , \22253 );
buf \U$22240 ( \22255 , \22254 );
buf \U$22241 ( \22256 , \22255 );
not \U$22242 ( \22257 , \22256 );
buf \U$22243 ( \22258 , \22257 );
buf \U$22244 ( \22259 , \22258 );
and \U$22245 ( \22260 , \22250 , \22259 );
not \U$22246 ( \22261 , \22250 );
buf \U$22247 ( \22262 , \22255 );
and \U$22248 ( \22263 , \22261 , \22262 );
nor \U$22249 ( \22264 , \22260 , \22263 );
buf \U$22250 ( \22265 , \22264 );
buf \U$22251 ( \22266 , \22265 );
buf \U$22252 ( \22267 , \20735 );
not \U$22253 ( \22268 , \22267 );
buf \U$22254 ( \22269 , \20752 );
not \U$22255 ( \22270 , \22269 );
or \U$22256 ( \22271 , \22268 , \22270 );
buf \U$22257 ( \22272 , \20752 );
buf \U$22258 ( \22273 , \20735 );
or \U$22259 ( \22274 , \22272 , \22273 );
buf \U$22260 ( \22275 , \20770 );
nand \U$22261 ( \22276 , \22274 , \22275 );
buf \U$22262 ( \22277 , \22276 );
buf \U$22263 ( \22278 , \22277 );
nand \U$22264 ( \22279 , \22271 , \22278 );
buf \U$22265 ( \22280 , \22279 );
xor \U$22266 ( \22281 , \21761 , \21778 );
xor \U$22267 ( \22282 , \22281 , \21796 );
buf \U$22268 ( \22283 , \22282 );
xor \U$22269 ( \22284 , \22280 , \22283 );
xor \U$22270 ( \22285 , \21818 , \21835 );
xor \U$22271 ( \22286 , \22285 , \21849 );
buf \U$22272 ( \22287 , \22286 );
xnor \U$22273 ( \22288 , \22284 , \22287 );
buf \U$22274 ( \22289 , \22288 );
nand \U$22275 ( \22290 , \22266 , \22289 );
buf \U$22276 ( \22291 , \22290 );
not \U$22277 ( \22292 , \22291 );
xor \U$22278 ( \22293 , \21977 , \21981 );
xor \U$22279 ( \22294 , \22293 , \22033 );
buf \U$22280 ( \22295 , \22294 );
not \U$22281 ( \22296 , \22295 );
or \U$22282 ( \22297 , \22292 , \22296 );
buf \U$22283 ( \22298 , \22288 );
not \U$22284 ( \22299 , \22298 );
buf \U$22285 ( \22300 , \22265 );
not \U$22286 ( \22301 , \22300 );
buf \U$22287 ( \22302 , \22301 );
buf \U$22288 ( \22303 , \22302 );
nand \U$22289 ( \22304 , \22299 , \22303 );
buf \U$22290 ( \22305 , \22304 );
nand \U$22291 ( \22306 , \22297 , \22305 );
buf \U$22292 ( \22307 , \22306 );
not \U$22293 ( \22308 , \22307 );
buf \U$22294 ( \22309 , \22308 );
buf \U$22295 ( \22310 , \22309 );
not \U$22296 ( \22311 , \22310 );
buf \U$22297 ( \22312 , \22311 );
buf \U$22298 ( \22313 , \22312 );
and \U$22299 ( \22314 , \22127 , \22313 );
not \U$22300 ( \22315 , \22127 );
buf \U$22301 ( \22316 , \22309 );
and \U$22302 ( \22317 , \22315 , \22316 );
nor \U$22303 ( \22318 , \22314 , \22317 );
buf \U$22304 ( \22319 , \22318 );
buf \U$22305 ( \22320 , \22319 );
xor \U$22306 ( \22321 , \21317 , \21323 );
and \U$22307 ( \22322 , \22321 , \21330 );
and \U$22308 ( \22323 , \21317 , \21323 );
or \U$22309 ( \22324 , \22322 , \22323 );
buf \U$22310 ( \22325 , \22324 );
buf \U$22311 ( \22326 , \22325 );
buf \U$22312 ( \22327 , \21016 );
not \U$22313 ( \22328 , \22327 );
buf \U$22314 ( \22329 , \14569 );
not \U$22315 ( \22330 , \22329 );
or \U$22316 ( \22331 , \22328 , \22330 );
buf \U$22317 ( \22332 , RIc0d78d0_6);
buf \U$22318 ( \22333 , RIc0dadc8_119);
xnor \U$22319 ( \22334 , \22332 , \22333 );
buf \U$22320 ( \22335 , \22334 );
buf \U$22321 ( \22336 , \22335 );
not \U$22322 ( \22337 , \22336 );
buf \U$22323 ( \22338 , \13005 );
nand \U$22324 ( \22339 , \22337 , \22338 );
buf \U$22325 ( \22340 , \22339 );
buf \U$22326 ( \22341 , \22340 );
nand \U$22327 ( \22342 , \22331 , \22341 );
buf \U$22328 ( \22343 , \22342 );
buf \U$22329 ( \22344 , \22343 );
not \U$22330 ( \22345 , \22344 );
buf \U$22331 ( \22346 , \22345 );
buf \U$22332 ( \22347 , \22346 );
buf \U$22333 ( \22348 , \21163 );
not \U$22334 ( \22349 , \22348 );
buf \U$22337 ( \22350 , \12923 );
buf \U$22338 ( \22351 , \22350 );
not \U$22339 ( \22352 , \22351 );
or \U$22340 ( \22353 , \22349 , \22352 );
buf \U$22341 ( \22354 , \16556 );
not \U$22342 ( \22355 , \22354 );
buf \U$22343 ( \22356 , \22355 );
buf \U$22344 ( \22357 , \22356 );
xor \U$22345 ( \22358 , RIc0dacd8_117, RIc0d79c0_8);
buf \U$22346 ( \22359 , \22358 );
nand \U$22347 ( \22360 , \22357 , \22359 );
buf \U$22348 ( \22361 , \22360 );
buf \U$22349 ( \22362 , \22361 );
nand \U$22350 ( \22363 , \22353 , \22362 );
buf \U$22351 ( \22364 , \22363 );
buf \U$22352 ( \22365 , \22364 );
xor \U$22353 ( \22366 , \22347 , \22365 );
buf \U$22354 ( \22367 , \21310 );
xor \U$22355 ( \22368 , \22366 , \22367 );
buf \U$22356 ( \22369 , \22368 );
buf \U$22357 ( \22370 , \22369 );
buf \U$22358 ( \22371 , \20505 );
not \U$22359 ( \22372 , \22371 );
buf \U$22360 ( \22373 , \20487 );
not \U$22361 ( \22374 , \22373 );
or \U$22362 ( \22375 , \22372 , \22374 );
buf \U$22363 ( \22376 , \20518 );
nand \U$22364 ( \22377 , \22375 , \22376 );
buf \U$22365 ( \22378 , \22377 );
buf \U$22366 ( \22379 , \22378 );
buf \U$22367 ( \22380 , \20484 );
buf \U$22368 ( \22381 , \20502 );
nand \U$22369 ( \22382 , \22380 , \22381 );
buf \U$22370 ( \22383 , \22382 );
buf \U$22371 ( \22384 , \22383 );
nand \U$22372 ( \22385 , \22379 , \22384 );
buf \U$22373 ( \22386 , \22385 );
buf \U$22374 ( \22387 , \22386 );
xor \U$22375 ( \22388 , \22370 , \22387 );
buf \U$22376 ( \22389 , \21504 );
buf \U$22377 ( \22390 , \21497 );
or \U$22378 ( \22391 , \22389 , \22390 );
buf \U$22379 ( \22392 , \21491 );
nand \U$22380 ( \22393 , \22391 , \22392 );
buf \U$22381 ( \22394 , \22393 );
buf \U$22382 ( \22395 , \22394 );
buf \U$22383 ( \22396 , \21504 );
buf \U$22384 ( \22397 , \21497 );
nand \U$22385 ( \22398 , \22396 , \22397 );
buf \U$22386 ( \22399 , \22398 );
buf \U$22387 ( \22400 , \22399 );
nand \U$22388 ( \22401 , \22395 , \22400 );
buf \U$22389 ( \22402 , \22401 );
buf \U$22390 ( \22403 , \22402 );
xor \U$22391 ( \22404 , \22388 , \22403 );
buf \U$22392 ( \22405 , \22404 );
buf \U$22393 ( \22406 , \22405 );
xor \U$22394 ( \22407 , \22326 , \22406 );
not \U$22395 ( \22408 , \21507 );
not \U$22396 ( \22409 , \21481 );
buf \U$22397 ( \22410 , \21390 );
not \U$22398 ( \22411 , \22410 );
buf \U$22399 ( \22412 , \22411 );
nand \U$22400 ( \22413 , \22409 , \22412 );
not \U$22401 ( \22414 , \22413 );
or \U$22402 ( \22415 , \22408 , \22414 );
not \U$22403 ( \22416 , \22412 );
nand \U$22404 ( \22417 , \22416 , \21481 );
nand \U$22405 ( \22418 , \22415 , \22417 );
buf \U$22406 ( \22419 , \22418 );
xor \U$22407 ( \22420 , \22407 , \22419 );
buf \U$22408 ( \22421 , \22420 );
buf \U$22409 ( \22422 , \22421 );
buf \U$22410 ( \22423 , \21364 );
not \U$22411 ( \22424 , \22423 );
buf \U$22412 ( \22425 , \21516 );
not \U$22413 ( \22426 , \22425 );
or \U$22414 ( \22427 , \22424 , \22426 );
buf \U$22415 ( \22428 , \21367 );
not \U$22416 ( \22429 , \22428 );
buf \U$22417 ( \22430 , \21510 );
not \U$22418 ( \22431 , \22430 );
or \U$22419 ( \22432 , \22429 , \22431 );
buf \U$22420 ( \22433 , \21354 );
nand \U$22421 ( \22434 , \22432 , \22433 );
buf \U$22422 ( \22435 , \22434 );
buf \U$22423 ( \22436 , \22435 );
nand \U$22424 ( \22437 , \22427 , \22436 );
buf \U$22425 ( \22438 , \22437 );
buf \U$22426 ( \22439 , \22438 );
or \U$22427 ( \22440 , \22422 , \22439 );
not \U$22428 ( \22441 , \20419 );
not \U$22429 ( \22442 , \20443 );
or \U$22430 ( \22443 , \22441 , \22442 );
not \U$22431 ( \22444 , \20446 );
not \U$22432 ( \22445 , \20422 );
or \U$22433 ( \22446 , \22444 , \22445 );
nand \U$22434 ( \22447 , \22446 , \20403 );
nand \U$22435 ( \22448 , \22443 , \22447 );
buf \U$22436 ( \22449 , \22448 );
not \U$22437 ( \22450 , \20568 );
not \U$22438 ( \22451 , \20533 );
or \U$22439 ( \22452 , \22450 , \22451 );
not \U$22440 ( \22453 , \20528 );
not \U$22441 ( \22454 , \20562 );
or \U$22442 ( \22455 , \22453 , \22454 );
nand \U$22443 ( \22456 , \22455 , \20476 );
nand \U$22444 ( \22457 , \22452 , \22456 );
buf \U$22445 ( \22458 , \22457 );
xor \U$22446 ( \22459 , \22449 , \22458 );
xor \U$22447 ( \22460 , \22056 , \22105 );
xor \U$22448 ( \22461 , \22460 , \22112 );
buf \U$22449 ( \22462 , \22461 );
buf \U$22450 ( \22463 , \22462 );
xor \U$22451 ( \22464 , \22459 , \22463 );
buf \U$22452 ( \22465 , \22464 );
buf \U$22453 ( \22466 , \22465 );
nand \U$22454 ( \22467 , \22440 , \22466 );
buf \U$22455 ( \22468 , \22467 );
buf \U$22456 ( \22469 , \22468 );
buf \U$22457 ( \22470 , \22421 );
buf \U$22458 ( \22471 , \22438 );
nand \U$22459 ( \22472 , \22470 , \22471 );
buf \U$22460 ( \22473 , \22472 );
buf \U$22461 ( \22474 , \22473 );
nand \U$22462 ( \22475 , \22469 , \22474 );
buf \U$22463 ( \22476 , \22475 );
buf \U$22464 ( \22477 , \22476 );
xor \U$22465 ( \22478 , \22320 , \22477 );
buf \U$22466 ( \22479 , \22258 );
not \U$22467 ( \22480 , \22479 );
buf \U$22468 ( \22481 , \22184 );
not \U$22469 ( \22482 , \22481 );
or \U$22470 ( \22483 , \22480 , \22482 );
buf \U$22471 ( \22484 , \22239 );
nand \U$22472 ( \22485 , \22483 , \22484 );
buf \U$22473 ( \22486 , \22485 );
buf \U$22474 ( \22487 , \22486 );
buf \U$22475 ( \22488 , \22181 );
buf \U$22476 ( \22489 , \22255 );
nand \U$22477 ( \22490 , \22488 , \22489 );
buf \U$22478 ( \22491 , \22490 );
buf \U$22479 ( \22492 , \22491 );
nand \U$22480 ( \22493 , \22487 , \22492 );
buf \U$22481 ( \22494 , \22493 );
buf \U$22482 ( \22495 , \22494 );
buf \U$22483 ( \22496 , \21754 );
not \U$22484 ( \22497 , \22496 );
buf \U$22485 ( \22498 , \13383 );
not \U$22486 ( \22499 , \22498 );
or \U$22487 ( \22500 , \22497 , \22499 );
buf \U$22488 ( \22501 , \1143 );
buf \U$22489 ( \22502 , RIc0d8cf8_49);
not \U$22490 ( \22503 , \22502 );
buf \U$22491 ( \22504 , \22503 );
and \U$22492 ( \22505 , RIc0d9928_75, \22504 );
not \U$22493 ( \22506 , RIc0d9928_75);
and \U$22494 ( \22507 , \22506 , RIc0d8cf8_49);
or \U$22495 ( \22508 , \22505 , \22507 );
buf \U$22496 ( \22509 , \22508 );
nand \U$22497 ( \22510 , \22501 , \22509 );
buf \U$22498 ( \22511 , \22510 );
buf \U$22499 ( \22512 , \22511 );
nand \U$22500 ( \22513 , \22500 , \22512 );
buf \U$22501 ( \22514 , \22513 );
buf \U$22502 ( \22515 , \22514 );
not \U$22503 ( \22516 , \22515 );
buf \U$22504 ( \22517 , \21967 );
not \U$22505 ( \22518 , \22517 );
buf \U$22506 ( \22519 , \13419 );
not \U$22507 ( \22520 , \22519 );
or \U$22508 ( \22521 , \22518 , \22520 );
buf \U$22509 ( \22522 , \14216 );
buf \U$22510 ( \22523 , RIc0d7d08_15);
buf \U$22511 ( \22524 , RIc0da918_109);
xor \U$22512 ( \22525 , \22523 , \22524 );
buf \U$22513 ( \22526 , \22525 );
buf \U$22514 ( \22527 , \22526 );
nand \U$22515 ( \22528 , \22522 , \22527 );
buf \U$22516 ( \22529 , \22528 );
buf \U$22517 ( \22530 , \22529 );
nand \U$22518 ( \22531 , \22521 , \22530 );
buf \U$22519 ( \22532 , \22531 );
buf \U$22520 ( \22533 , \22532 );
buf \U$22521 ( \22534 , \22212 );
not \U$22522 ( \22535 , \22534 );
buf \U$22523 ( \22536 , \18767 );
not \U$22524 ( \22537 , \22536 );
or \U$22525 ( \22538 , \22535 , \22537 );
buf \U$22526 ( \22539 , \2960 );
buf \U$22527 ( \22540 , RIc0d8848_39);
buf \U$22528 ( \22541 , RIc0d9dd8_85);
xor \U$22529 ( \22542 , \22540 , \22541 );
buf \U$22530 ( \22543 , \22542 );
buf \U$22531 ( \22544 , \22543 );
nand \U$22532 ( \22545 , \22539 , \22544 );
buf \U$22533 ( \22546 , \22545 );
buf \U$22534 ( \22547 , \22546 );
nand \U$22535 ( \22548 , \22538 , \22547 );
buf \U$22536 ( \22549 , \22548 );
buf \U$22537 ( \22550 , \22549 );
xnor \U$22538 ( \22551 , \22533 , \22550 );
buf \U$22539 ( \22552 , \22551 );
buf \U$22540 ( \22553 , \22552 );
not \U$22541 ( \22554 , \22553 );
or \U$22542 ( \22555 , \22516 , \22554 );
buf \U$22543 ( \22556 , \22552 );
buf \U$22544 ( \22557 , \22514 );
or \U$22545 ( \22558 , \22556 , \22557 );
nand \U$22546 ( \22559 , \22555 , \22558 );
buf \U$22547 ( \22560 , \22559 );
buf \U$22548 ( \22561 , \22560 );
xor \U$22549 ( \22562 , RIc0d9bf8_81, RIc0d8a28_43);
buf \U$22550 ( \22563 , \22562 );
not \U$22551 ( \22564 , \22563 );
buf \U$22552 ( \22565 , \1077 );
not \U$22553 ( \22566 , \22565 );
or \U$22554 ( \22567 , \22564 , \22566 );
buf \U$22555 ( \22568 , \1056 );
buf \U$22556 ( \22569 , \21600 );
nand \U$22557 ( \22570 , \22568 , \22569 );
buf \U$22558 ( \22571 , \22570 );
buf \U$22559 ( \22572 , \22571 );
buf \U$22560 ( \22573 , \1078 );
or \U$22561 ( \22574 , \22572 , \22573 );
nand \U$22562 ( \22575 , \22567 , \22574 );
buf \U$22563 ( \22576 , \22575 );
buf \U$22564 ( \22577 , \22576 );
buf \U$22565 ( \22578 , \22358 );
not \U$22566 ( \22579 , \22578 );
buf \U$22567 ( \22580 , \13684 );
not \U$22568 ( \22581 , \22580 );
or \U$22569 ( \22582 , \22579 , \22581 );
buf \U$22570 ( \22583 , \12937 );
xor \U$22571 ( \22584 , RIc0dacd8_117, RIc0d7948_7);
buf \U$22572 ( \22585 , \22584 );
nand \U$22573 ( \22586 , \22583 , \22585 );
buf \U$22574 ( \22587 , \22586 );
buf \U$22575 ( \22588 , \22587 );
nand \U$22576 ( \22589 , \22582 , \22588 );
buf \U$22577 ( \22590 , \22589 );
buf \U$22578 ( \22591 , \22590 );
xor \U$22579 ( \22592 , \22577 , \22591 );
buf \U$22580 ( \22593 , \14186 );
not \U$22581 ( \22594 , \22593 );
buf \U$22582 ( \22595 , \22594 );
buf \U$22583 ( \22596 , \22595 );
buf \U$22584 ( \22597 , \21683 );
not \U$22585 ( \22598 , \22597 );
buf \U$22586 ( \22599 , \22598 );
buf \U$22587 ( \22600 , \22599 );
or \U$22588 ( \22601 , \22596 , \22600 );
buf \U$22589 ( \22602 , \12278 );
buf \U$22590 ( \22603 , RIc0d7a38_9);
buf \U$22591 ( \22604 , RIc0dabe8_115);
xnor \U$22592 ( \22605 , \22603 , \22604 );
buf \U$22593 ( \22606 , \22605 );
buf \U$22594 ( \22607 , \22606 );
or \U$22595 ( \22608 , \22602 , \22607 );
nand \U$22596 ( \22609 , \22601 , \22608 );
buf \U$22597 ( \22610 , \22609 );
buf \U$22598 ( \22611 , \22610 );
xor \U$22599 ( \22612 , \22592 , \22611 );
buf \U$22600 ( \22613 , \22612 );
buf \U$22601 ( \22614 , \22613 );
xor \U$22602 ( \22615 , \22561 , \22614 );
buf \U$22603 ( \22616 , \21641 );
not \U$22604 ( \22617 , \22616 );
buf \U$22605 ( \22618 , \13569 );
not \U$22606 ( \22619 , \22618 );
or \U$22607 ( \22620 , \22617 , \22619 );
buf \U$22608 ( \22621 , \4008 );
xor \U$22609 ( \22622 , RIc0da198_93, RIc0d8488_31);
buf \U$22610 ( \22623 , \22622 );
nand \U$22611 ( \22624 , \22621 , \22623 );
buf \U$22612 ( \22625 , \22624 );
buf \U$22613 ( \22626 , \22625 );
nand \U$22614 ( \22627 , \22620 , \22626 );
buf \U$22615 ( \22628 , \22627 );
buf \U$22616 ( \22629 , \21789 );
not \U$22617 ( \22630 , \22629 );
buf \U$22620 ( \22631 , \4042 );
buf \U$22621 ( \22632 , \22631 );
not \U$22622 ( \22633 , \22632 );
or \U$22623 ( \22634 , \22630 , \22633 );
buf \U$22624 ( \22635 , \16676 );
buf \U$22625 ( \22636 , RIc0da558_101);
buf \U$22626 ( \22637 , RIc0d80c8_23);
xor \U$22627 ( \22638 , \22636 , \22637 );
buf \U$22628 ( \22639 , \22638 );
buf \U$22629 ( \22640 , \22639 );
nand \U$22630 ( \22641 , \22635 , \22640 );
buf \U$22631 ( \22642 , \22641 );
buf \U$22632 ( \22643 , \22642 );
nand \U$22633 ( \22644 , \22634 , \22643 );
buf \U$22634 ( \22645 , \22644 );
xor \U$22635 ( \22646 , \22628 , \22645 );
buf \U$22636 ( \22647 , \21719 );
not \U$22637 ( \22648 , \22647 );
buf \U$22638 ( \22649 , \618 );
not \U$22639 ( \22650 , \22649 );
or \U$22640 ( \22651 , \22648 , \22650 );
buf \U$22641 ( \22652 , \816 );
buf \U$22642 ( \22653 , RIc0d8758_37);
buf \U$22643 ( \22654 , RIc0d9ec8_87);
xor \U$22644 ( \22655 , \22653 , \22654 );
buf \U$22645 ( \22656 , \22655 );
buf \U$22646 ( \22657 , \22656 );
nand \U$22647 ( \22658 , \22652 , \22657 );
buf \U$22648 ( \22659 , \22658 );
buf \U$22649 ( \22660 , \22659 );
nand \U$22650 ( \22661 , \22651 , \22660 );
buf \U$22651 ( \22662 , \22661 );
xor \U$22652 ( \22663 , \22646 , \22662 );
buf \U$22653 ( \22664 , \22663 );
xor \U$22654 ( \22665 , \22615 , \22664 );
buf \U$22655 ( \22666 , \22665 );
buf \U$22656 ( \22667 , \22666 );
xor \U$22657 ( \22668 , \22495 , \22667 );
buf \U$22658 ( \22669 , \21828 );
not \U$22659 ( \22670 , \22669 );
buf \U$22660 ( \22671 , \18057 );
not \U$22661 ( \22672 , \22671 );
or \U$22662 ( \22673 , \22670 , \22672 );
buf \U$22663 ( \22674 , \791 );
buf \U$22664 ( \22675 , RIc0d8de8_51);
buf \U$22665 ( \22676 , RIc0d9838_73);
xor \U$22666 ( \22677 , \22675 , \22676 );
buf \U$22667 ( \22678 , \22677 );
buf \U$22668 ( \22679 , \22678 );
nand \U$22669 ( \22680 , \22674 , \22679 );
buf \U$22670 ( \22681 , \22680 );
buf \U$22671 ( \22682 , \22681 );
nand \U$22672 ( \22683 , \22673 , \22682 );
buf \U$22673 ( \22684 , \22683 );
buf \U$22674 ( \22685 , \22684 );
buf \U$22675 ( \22686 , \21586 );
not \U$22676 ( \22687 , \22686 );
buf \U$22677 ( \22688 , \12402 );
not \U$22678 ( \22689 , \22688 );
or \U$22679 ( \22690 , \22687 , \22689 );
buf \U$22680 ( \22691 , \14405 );
buf \U$22681 ( \22692 , RIc0d7b28_11);
buf \U$22682 ( \22693 , RIc0daaf8_113);
xor \U$22683 ( \22694 , \22692 , \22693 );
buf \U$22684 ( \22695 , \22694 );
buf \U$22685 ( \22696 , \22695 );
nand \U$22686 ( \22697 , \22691 , \22696 );
buf \U$22687 ( \22698 , \22697 );
buf \U$22688 ( \22699 , \22698 );
nand \U$22689 ( \22700 , \22690 , \22699 );
buf \U$22690 ( \22701 , \22700 );
buf \U$22691 ( \22702 , \22701 );
not \U$22692 ( \22703 , \22702 );
buf \U$22693 ( \22704 , \22703 );
buf \U$22694 ( \22705 , \22704 );
xor \U$22695 ( \22706 , \22685 , \22705 );
buf \U$22696 ( \22707 , \22011 );
not \U$22697 ( \22708 , \22707 );
buf \U$22698 ( \22709 , \16744 );
not \U$22699 ( \22710 , \22709 );
or \U$22700 ( \22711 , \22708 , \22710 );
buf \U$22701 ( \22712 , \16750 );
buf \U$22702 ( \22713 , RIc0da468_99);
buf \U$22703 ( \22714 , RIc0d81b8_25);
xor \U$22704 ( \22715 , \22713 , \22714 );
buf \U$22705 ( \22716 , \22715 );
buf \U$22706 ( \22717 , \22716 );
nand \U$22707 ( \22718 , \22712 , \22717 );
buf \U$22708 ( \22719 , \22718 );
buf \U$22709 ( \22720 , \22719 );
nand \U$22710 ( \22721 , \22711 , \22720 );
buf \U$22711 ( \22722 , \22721 );
buf \U$22712 ( \22723 , \22722 );
xor \U$22713 ( \22724 , \22706 , \22723 );
buf \U$22714 ( \22725 , \22724 );
buf \U$22715 ( \22726 , \21946 );
not \U$22716 ( \22727 , \22726 );
buf \U$22717 ( \22728 , \14346 );
not \U$22718 ( \22729 , \22728 );
or \U$22719 ( \22730 , \22727 , \22729 );
buf \U$22720 ( \22731 , \14353 );
buf \U$22721 ( \22732 , RIc0daa08_111);
buf \U$22722 ( \22733 , RIc0d7c18_13);
xor \U$22723 ( \22734 , \22732 , \22733 );
buf \U$22724 ( \22735 , \22734 );
buf \U$22725 ( \22736 , \22735 );
nand \U$22726 ( \22737 , \22731 , \22736 );
buf \U$22727 ( \22738 , \22737 );
buf \U$22728 ( \22739 , \22738 );
nand \U$22729 ( \22740 , \22730 , \22739 );
buf \U$22730 ( \22741 , \22740 );
buf \U$22731 ( \22742 , \15793 );
not \U$22732 ( \22743 , \22742 );
buf \U$22733 ( \22744 , \22743 );
buf \U$22734 ( \22745 , \22744 );
not \U$22735 ( \22746 , \22745 );
buf \U$22736 ( \22747 , \14468 );
not \U$22737 ( \22748 , \22747 );
or \U$22738 ( \22749 , \22746 , \22748 );
buf \U$22739 ( \22750 , RIc0db098_125);
nand \U$22740 ( \22751 , \22749 , \22750 );
buf \U$22741 ( \22752 , \22751 );
xor \U$22742 ( \22753 , \22741 , \22752 );
buf \U$22743 ( \22754 , \1351 );
buf \U$22744 ( \22755 , \21699 );
and \U$22745 ( \22756 , \22754 , \22755 );
buf \U$22746 ( \22757 , \3985 );
buf \U$22747 ( \22758 , RIc0d8b18_45);
buf \U$22748 ( \22759 , RIc0d9b08_79);
xor \U$22749 ( \22760 , \22758 , \22759 );
buf \U$22750 ( \22761 , \22760 );
buf \U$22751 ( \22762 , \22761 );
and \U$22752 ( \22763 , \22757 , \22762 );
nor \U$22753 ( \22764 , \22756 , \22763 );
buf \U$22754 ( \22765 , \22764 );
buf \U$22755 ( \22766 , \22765 );
not \U$22756 ( \22767 , \22766 );
buf \U$22757 ( \22768 , \22767 );
and \U$22758 ( \22769 , \22753 , \22768 );
not \U$22759 ( \22770 , \22753 );
and \U$22760 ( \22771 , \22770 , \22765 );
nor \U$22761 ( \22772 , \22769 , \22771 );
xor \U$22762 ( \22773 , \22725 , \22772 );
buf \U$22763 ( \22774 , \22343 );
buf \U$22764 ( \22775 , \22172 );
not \U$22765 ( \22776 , \22775 );
buf \U$22766 ( \22777 , \437 );
not \U$22767 ( \22778 , \22777 );
or \U$22768 ( \22779 , \22776 , \22778 );
buf \U$22769 ( \22780 , \846 );
buf \U$22770 ( \22781 , RIc0d8668_35);
buf \U$22771 ( \22782 , RIc0d9fb8_89);
xor \U$22772 ( \22783 , \22781 , \22782 );
buf \U$22773 ( \22784 , \22783 );
buf \U$22774 ( \22785 , \22784 );
nand \U$22775 ( \22786 , \22780 , \22785 );
buf \U$22776 ( \22787 , \22786 );
buf \U$22777 ( \22788 , \22787 );
nand \U$22778 ( \22789 , \22779 , \22788 );
buf \U$22779 ( \22790 , \22789 );
buf \U$22780 ( \22791 , \22790 );
xor \U$22781 ( \22792 , \22774 , \22791 );
buf \U$22782 ( \22793 , \13178 );
buf \U$22783 ( \22794 , \22335 );
or \U$22784 ( \22795 , \22793 , \22794 );
buf \U$22785 ( \22796 , \13953 );
not \U$22786 ( \22797 , \22796 );
buf \U$22787 ( \22798 , \22797 );
buf \U$22788 ( \22799 , \22798 );
buf \U$22789 ( \22800 , RIc0dadc8_119);
buf \U$22790 ( \22801 , RIc0d7858_5);
xor \U$22791 ( \22802 , \22800 , \22801 );
buf \U$22792 ( \22803 , \22802 );
buf \U$22793 ( \22804 , \22803 );
not \U$22794 ( \22805 , \22804 );
buf \U$22795 ( \22806 , \22805 );
buf \U$22796 ( \22807 , \22806 );
or \U$22797 ( \22808 , \22799 , \22807 );
nand \U$22798 ( \22809 , \22795 , \22808 );
buf \U$22799 ( \22810 , \22809 );
buf \U$22800 ( \22811 , \22810 );
xor \U$22801 ( \22812 , \22792 , \22811 );
buf \U$22802 ( \22813 , \22812 );
xnor \U$22803 ( \22814 , \22773 , \22813 );
buf \U$22804 ( \22815 , \22814 );
xor \U$22805 ( \22816 , \22668 , \22815 );
buf \U$22806 ( \22817 , \22816 );
buf \U$22807 ( \22818 , \22817 );
xor \U$22808 ( \22819 , \22326 , \22406 );
and \U$22809 ( \22820 , \22819 , \22419 );
and \U$22810 ( \22821 , \22326 , \22406 );
or \U$22811 ( \22822 , \22820 , \22821 );
buf \U$22812 ( \22823 , \22822 );
buf \U$22813 ( \22824 , \22823 );
xor \U$22814 ( \22825 , \22818 , \22824 );
buf \U$22815 ( \22826 , \20976 );
not \U$22816 ( \22827 , \22826 );
buf \U$22817 ( \22828 , \21189 );
not \U$22818 ( \22829 , \22828 );
or \U$22819 ( \22830 , \22827 , \22829 );
buf \U$22820 ( \22831 , \20776 );
nand \U$22821 ( \22832 , \22830 , \22831 );
buf \U$22822 ( \22833 , \22832 );
buf \U$22823 ( \22834 , \22833 );
buf \U$22824 ( \22835 , \20976 );
not \U$22825 ( \22836 , \22835 );
buf \U$22826 ( \22837 , \21192 );
nand \U$22827 ( \22838 , \22836 , \22837 );
buf \U$22828 ( \22839 , \22838 );
buf \U$22829 ( \22840 , \22839 );
nand \U$22830 ( \22841 , \22834 , \22840 );
buf \U$22831 ( \22842 , \22841 );
buf \U$22832 ( \22843 , \22842 );
buf \U$22833 ( \22844 , \21070 );
not \U$22834 ( \22845 , \22844 );
buf \U$22835 ( \22846 , \21064 );
not \U$22836 ( \22847 , \22846 );
or \U$22837 ( \22848 , \22845 , \22847 );
buf \U$22838 ( \22849 , \21094 );
nand \U$22839 ( \22850 , \22848 , \22849 );
buf \U$22840 ( \22851 , \22850 );
buf \U$22841 ( \22852 , \22851 );
buf \U$22842 ( \22853 , \21061 );
buf \U$22843 ( \22854 , \21043 );
nand \U$22844 ( \22855 , \22853 , \22854 );
buf \U$22845 ( \22856 , \22855 );
buf \U$22846 ( \22857 , \22856 );
nand \U$22847 ( \22858 , \22852 , \22857 );
buf \U$22848 ( \22859 , \22858 );
buf \U$22849 ( \22860 , \22859 );
xor \U$22850 ( \22861 , \21441 , \21455 );
and \U$22851 ( \22862 , \22861 , \21476 );
and \U$22852 ( \22863 , \21441 , \21455 );
or \U$22853 ( \22864 , \22862 , \22863 );
buf \U$22854 ( \22865 , \22864 );
buf \U$22855 ( \22866 , \22865 );
xor \U$22856 ( \22867 , \22860 , \22866 );
buf \U$22857 ( \22868 , \20932 );
not \U$22858 ( \22869 , \22868 );
buf \U$22859 ( \22870 , \20956 );
not \U$22860 ( \22871 , \22870 );
or \U$22861 ( \22872 , \22869 , \22871 );
buf \U$22862 ( \22873 , \20911 );
nand \U$22863 ( \22874 , \22872 , \22873 );
buf \U$22864 ( \22875 , \22874 );
buf \U$22865 ( \22876 , \22875 );
buf \U$22866 ( \22877 , \20962 );
buf \U$22867 ( \22878 , \20929 );
nand \U$22868 ( \22879 , \22877 , \22878 );
buf \U$22869 ( \22880 , \22879 );
buf \U$22870 ( \22881 , \22880 );
nand \U$22871 ( \22882 , \22876 , \22881 );
buf \U$22872 ( \22883 , \22882 );
buf \U$22873 ( \22884 , \22883 );
xor \U$22874 ( \22885 , \22867 , \22884 );
buf \U$22875 ( \22886 , \22885 );
buf \U$22876 ( \22887 , \22886 );
not \U$22877 ( \22888 , \22887 );
buf \U$22878 ( \22889 , \21004 );
buf \U$22879 ( \22890 , \20987 );
or \U$22880 ( \22891 , \22889 , \22890 );
buf \U$22881 ( \22892 , \21022 );
nand \U$22882 ( \22893 , \22891 , \22892 );
buf \U$22883 ( \22894 , \22893 );
buf \U$22884 ( \22895 , \22894 );
buf \U$22885 ( \22896 , \21004 );
buf \U$22886 ( \22897 , \20987 );
nand \U$22887 ( \22898 , \22896 , \22897 );
buf \U$22888 ( \22899 , \22898 );
buf \U$22889 ( \22900 , \22899 );
nand \U$22890 ( \22901 , \22895 , \22900 );
buf \U$22891 ( \22902 , \22901 );
buf \U$22892 ( \22903 , \22902 );
buf \U$22893 ( \22904 , \20791 );
not \U$22894 ( \22905 , \22904 );
buf \U$22895 ( \22906 , \20812 );
not \U$22896 ( \22907 , \22906 );
or \U$22897 ( \22908 , \22905 , \22907 );
buf \U$22898 ( \22909 , \20812 );
buf \U$22899 ( \22910 , \20791 );
or \U$22900 ( \22911 , \22909 , \22910 );
buf \U$22901 ( \22912 , \20829 );
nand \U$22902 ( \22913 , \22911 , \22912 );
buf \U$22903 ( \22914 , \22913 );
buf \U$22904 ( \22915 , \22914 );
nand \U$22905 ( \22916 , \22908 , \22915 );
buf \U$22906 ( \22917 , \22916 );
buf \U$22907 ( \22918 , \22917 );
xor \U$22908 ( \22919 , \22903 , \22918 );
buf \U$22909 ( \22920 , \21153 );
buf \U$22910 ( \22921 , \21137 );
nor \U$22911 ( \22922 , \22920 , \22921 );
buf \U$22912 ( \22923 , \22922 );
buf \U$22913 ( \22924 , \22923 );
buf \U$22914 ( \22925 , \21169 );
or \U$22915 ( \22926 , \22924 , \22925 );
buf \U$22916 ( \22927 , \21153 );
buf \U$22917 ( \22928 , \21137 );
nand \U$22918 ( \22929 , \22927 , \22928 );
buf \U$22919 ( \22930 , \22929 );
buf \U$22920 ( \22931 , \22930 );
nand \U$22921 ( \22932 , \22926 , \22931 );
buf \U$22922 ( \22933 , \22932 );
buf \U$22923 ( \22934 , \22933 );
xor \U$22924 ( \22935 , \22919 , \22934 );
buf \U$22925 ( \22936 , \22935 );
buf \U$22926 ( \22937 , \21025 );
not \U$22927 ( \22938 , \22937 );
buf \U$22928 ( \22939 , \21104 );
not \U$22929 ( \22940 , \22939 );
or \U$22930 ( \22941 , \22938 , \22940 );
buf \U$22931 ( \22942 , \21179 );
nand \U$22932 ( \22943 , \22941 , \22942 );
buf \U$22933 ( \22944 , \22943 );
buf \U$22934 ( \22945 , \22944 );
buf \U$22935 ( \22946 , \21107 );
buf \U$22936 ( \22947 , \21114 );
nand \U$22937 ( \22948 , \22946 , \22947 );
buf \U$22938 ( \22949 , \22948 );
buf \U$22939 ( \22950 , \22949 );
nand \U$22940 ( \22951 , \22945 , \22950 );
buf \U$22941 ( \22952 , \22951 );
buf \U$22942 ( \22953 , \22952 );
not \U$22943 ( \22954 , \22953 );
buf \U$22944 ( \22955 , \22954 );
xor \U$22945 ( \22956 , \22936 , \22955 );
buf \U$22946 ( \22957 , \22956 );
not \U$22947 ( \22958 , \22957 );
or \U$22948 ( \22959 , \22888 , \22958 );
buf \U$22949 ( \22960 , \22956 );
buf \U$22950 ( \22961 , \22886 );
or \U$22951 ( \22962 , \22960 , \22961 );
nand \U$22952 ( \22963 , \22959 , \22962 );
buf \U$22953 ( \22964 , \22963 );
buf \U$22954 ( \22965 , \22964 );
xor \U$22955 ( \22966 , \22843 , \22965 );
xor \U$22956 ( \22967 , \21408 , \21423 );
and \U$22957 ( \22968 , \22967 , \21479 );
and \U$22958 ( \22969 , \21408 , \21423 );
or \U$22959 ( \22970 , \22968 , \22969 );
buf \U$22960 ( \22971 , \22970 );
buf \U$22961 ( \22972 , \22971 );
buf \U$22962 ( \22973 , \20830 );
not \U$22963 ( \22974 , \22973 );
buf \U$22964 ( \22975 , \20966 );
not \U$22965 ( \22976 , \22975 );
or \U$22966 ( \22977 , \22974 , \22976 );
buf \U$22967 ( \22978 , \20886 );
nand \U$22968 ( \22979 , \22977 , \22978 );
buf \U$22969 ( \22980 , \22979 );
buf \U$22970 ( \22981 , \22980 );
buf \U$22971 ( \22982 , \20830 );
not \U$22972 ( \22983 , \22982 );
buf \U$22973 ( \22984 , \20972 );
nand \U$22974 ( \22985 , \22983 , \22984 );
buf \U$22975 ( \22986 , \22985 );
buf \U$22976 ( \22987 , \22986 );
nand \U$22977 ( \22988 , \22981 , \22987 );
buf \U$22978 ( \22989 , \22988 );
buf \U$22979 ( \22990 , \22989 );
xor \U$22980 ( \22991 , \22972 , \22990 );
xor \U$22981 ( \22992 , \21668 , \21627 );
xnor \U$22982 ( \22993 , \22992 , \21732 );
buf \U$22983 ( \22994 , \22993 );
xor \U$22984 ( \22995 , \22991 , \22994 );
buf \U$22985 ( \22996 , \22995 );
buf \U$22986 ( \22997 , \22996 );
and \U$22987 ( \22998 , \22966 , \22997 );
and \U$22988 ( \22999 , \22843 , \22965 );
or \U$22989 ( \23000 , \22998 , \22999 );
buf \U$22990 ( \23001 , \23000 );
buf \U$22991 ( \23002 , \23001 );
xor \U$22992 ( \23003 , \22825 , \23002 );
buf \U$22993 ( \23004 , \23003 );
buf \U$22994 ( \23005 , \23004 );
xor \U$22995 ( \23006 , \22478 , \23005 );
buf \U$22996 ( \23007 , \23006 );
xor \U$22997 ( \23008 , \22370 , \22387 );
and \U$22998 ( \23009 , \23008 , \22403 );
and \U$22999 ( \23010 , \22370 , \22387 );
or \U$23000 ( \23011 , \23009 , \23010 );
buf \U$23001 ( \23012 , \23011 );
buf \U$23002 ( \23013 , \23012 );
xor \U$23003 ( \23014 , \22347 , \22365 );
and \U$23004 ( \23015 , \23014 , \22367 );
and \U$23005 ( \23016 , \22347 , \22365 );
or \U$23006 ( \23017 , \23015 , \23016 );
buf \U$23007 ( \23018 , \23017 );
buf \U$23008 ( \23019 , \23018 );
buf \U$23009 ( \23020 , \22085 );
not \U$23010 ( \23021 , \23020 );
buf \U$23011 ( \23022 , \22070 );
not \U$23012 ( \23023 , \23022 );
or \U$23013 ( \23024 , \23021 , \23023 );
buf \U$23014 ( \23025 , \22070 );
buf \U$23015 ( \23026 , \22085 );
or \U$23016 ( \23027 , \23025 , \23026 );
buf \U$23017 ( \23028 , \22101 );
nand \U$23018 ( \23029 , \23027 , \23028 );
buf \U$23019 ( \23030 , \23029 );
buf \U$23020 ( \23031 , \23030 );
nand \U$23021 ( \23032 , \23024 , \23031 );
buf \U$23022 ( \23033 , \23032 );
buf \U$23023 ( \23034 , \23033 );
xor \U$23024 ( \23035 , \23019 , \23034 );
xor \U$23025 ( \23036 , \22860 , \22866 );
and \U$23026 ( \23037 , \23036 , \22884 );
and \U$23027 ( \23038 , \22860 , \22866 );
or \U$23028 ( \23039 , \23037 , \23038 );
buf \U$23029 ( \23040 , \23039 );
buf \U$23030 ( \23041 , \23040 );
xor \U$23031 ( \23042 , \23035 , \23041 );
buf \U$23032 ( \23043 , \23042 );
buf \U$23033 ( \23044 , \23043 );
xor \U$23034 ( \23045 , \23013 , \23044 );
buf \U$23035 ( \23046 , \22936 );
buf \U$23036 ( \23047 , \22886 );
or \U$23037 ( \23048 , \23046 , \23047 );
buf \U$23038 ( \23049 , \22955 );
not \U$23039 ( \23050 , \23049 );
buf \U$23040 ( \23051 , \23050 );
buf \U$23041 ( \23052 , \23051 );
nand \U$23042 ( \23053 , \23048 , \23052 );
buf \U$23043 ( \23054 , \23053 );
buf \U$23044 ( \23055 , \23054 );
buf \U$23045 ( \23056 , \22936 );
buf \U$23046 ( \23057 , \22886 );
nand \U$23047 ( \23058 , \23056 , \23057 );
buf \U$23048 ( \23059 , \23058 );
buf \U$23049 ( \23060 , \23059 );
nand \U$23050 ( \23061 , \23055 , \23060 );
buf \U$23051 ( \23062 , \23061 );
buf \U$23052 ( \23063 , \23062 );
xor \U$23053 ( \23064 , \23045 , \23063 );
buf \U$23054 ( \23065 , \23064 );
buf \U$23055 ( \23066 , \23065 );
xor \U$23056 ( \23067 , \22449 , \22458 );
and \U$23057 ( \23068 , \23067 , \22463 );
and \U$23058 ( \23069 , \22449 , \22458 );
or \U$23059 ( \23070 , \23068 , \23069 );
buf \U$23060 ( \23071 , \23070 );
buf \U$23061 ( \23072 , \23071 );
xor \U$23062 ( \23073 , \23066 , \23072 );
not \U$23063 ( \23074 , \21705 );
not \U$23064 ( \23075 , \21725 );
or \U$23065 ( \23076 , \23074 , \23075 );
not \U$23066 ( \23077 , \21728 );
not \U$23067 ( \23078 , \21708 );
or \U$23068 ( \23079 , \23077 , \23078 );
nand \U$23069 ( \23080 , \23079 , \21689 );
nand \U$23070 ( \23081 , \23076 , \23080 );
buf \U$23071 ( \23082 , \23081 );
buf \U$23072 ( \23083 , \22218 );
buf \U$23073 ( \23084 , \22202 );
or \U$23074 ( \23085 , \23083 , \23084 );
buf \U$23075 ( \23086 , \23085 );
not \U$23076 ( \23087 , \23086 );
not \U$23077 ( \23088 , \22235 );
or \U$23078 ( \23089 , \23087 , \23088 );
buf \U$23079 ( \23090 , \22202 );
buf \U$23080 ( \23091 , \22218 );
nand \U$23081 ( \23092 , \23090 , \23091 );
buf \U$23082 ( \23093 , \23092 );
nand \U$23083 ( \23094 , \23089 , \23093 );
buf \U$23084 ( \23095 , \23094 );
xor \U$23085 ( \23096 , \23082 , \23095 );
xor \U$23086 ( \23097 , \21936 , \21953 );
and \U$23087 ( \23098 , \23097 , \21974 );
and \U$23088 ( \23099 , \21936 , \21953 );
or \U$23089 ( \23100 , \23098 , \23099 );
buf \U$23090 ( \23101 , \23100 );
buf \U$23091 ( \23102 , \23101 );
xor \U$23092 ( \23103 , \23096 , \23102 );
buf \U$23093 ( \23104 , \23103 );
buf \U$23094 ( \23105 , \23104 );
xor \U$23095 ( \23106 , \22903 , \22918 );
and \U$23096 ( \23107 , \23106 , \22934 );
and \U$23097 ( \23108 , \22903 , \22918 );
or \U$23098 ( \23109 , \23107 , \23108 );
buf \U$23099 ( \23110 , \23109 );
buf \U$23100 ( \23111 , \23110 );
and \U$23101 ( \23112 , \23105 , \23111 );
not \U$23102 ( \23113 , \23105 );
buf \U$23103 ( \23114 , \23110 );
not \U$23104 ( \23115 , \23114 );
buf \U$23105 ( \23116 , \23115 );
buf \U$23106 ( \23117 , \23116 );
and \U$23107 ( \23118 , \23113 , \23117 );
nor \U$23108 ( \23119 , \23112 , \23118 );
buf \U$23109 ( \23120 , \23119 );
buf \U$23110 ( \23121 , \23120 );
buf \U$23111 ( \23122 , \21665 );
buf \U$23112 ( \23123 , \21630 );
or \U$23113 ( \23124 , \23122 , \23123 );
buf \U$23114 ( \23125 , \21647 );
nand \U$23115 ( \23126 , \23124 , \23125 );
buf \U$23116 ( \23127 , \23126 );
buf \U$23117 ( \23128 , \23127 );
buf \U$23118 ( \23129 , \21665 );
buf \U$23119 ( \23130 , \21630 );
nand \U$23120 ( \23131 , \23129 , \23130 );
buf \U$23121 ( \23132 , \23131 );
buf \U$23122 ( \23133 , \23132 );
nand \U$23123 ( \23134 , \23128 , \23133 );
buf \U$23124 ( \23135 , \23134 );
buf \U$23125 ( \23136 , \23135 );
xor \U$23126 ( \23137 , \22144 , \22161 );
and \U$23127 ( \23138 , \23137 , \22179 );
and \U$23128 ( \23139 , \22144 , \22161 );
or \U$23129 ( \23140 , \23138 , \23139 );
buf \U$23130 ( \23141 , \23140 );
buf \U$23131 ( \23142 , \23141 );
xor \U$23132 ( \23143 , \23136 , \23142 );
xor \U$23133 ( \23144 , \21593 , \21607 );
and \U$23134 ( \23145 , \23144 , \21625 );
and \U$23135 ( \23146 , \21593 , \21607 );
or \U$23136 ( \23147 , \23145 , \23146 );
buf \U$23137 ( \23148 , \23147 );
buf \U$23138 ( \23149 , \23148 );
xor \U$23139 ( \23150 , \23143 , \23149 );
buf \U$23140 ( \23151 , \23150 );
buf \U$23141 ( \23152 , \23151 );
not \U$23142 ( \23153 , \23152 );
buf \U$23143 ( \23154 , \23153 );
buf \U$23144 ( \23155 , \23154 );
and \U$23145 ( \23156 , \23121 , \23155 );
not \U$23146 ( \23157 , \23121 );
buf \U$23147 ( \23158 , \23151 );
and \U$23148 ( \23159 , \23157 , \23158 );
nor \U$23149 ( \23160 , \23156 , \23159 );
buf \U$23150 ( \23161 , \23160 );
buf \U$23151 ( \23162 , \23161 );
not \U$23152 ( \23163 , \23162 );
buf \U$23153 ( \23164 , \23163 );
buf \U$23154 ( \23165 , \23164 );
not \U$23155 ( \23166 , \23165 );
buf \U$23156 ( \23167 , \22971 );
not \U$23157 ( \23168 , \23167 );
buf \U$23158 ( \23169 , \22989 );
not \U$23159 ( \23170 , \23169 );
or \U$23160 ( \23171 , \23168 , \23170 );
buf \U$23161 ( \23172 , \22989 );
buf \U$23162 ( \23173 , \22971 );
or \U$23163 ( \23174 , \23172 , \23173 );
buf \U$23164 ( \23175 , \22993 );
nand \U$23165 ( \23176 , \23174 , \23175 );
buf \U$23166 ( \23177 , \23176 );
buf \U$23167 ( \23178 , \23177 );
nand \U$23168 ( \23179 , \23171 , \23178 );
buf \U$23169 ( \23180 , \23179 );
buf \U$23170 ( \23181 , \23180 );
not \U$23171 ( \23182 , \23181 );
buf \U$23172 ( \23183 , \23182 );
buf \U$23173 ( \23184 , \23183 );
not \U$23174 ( \23185 , \23184 );
or \U$23175 ( \23186 , \23166 , \23185 );
buf \U$23176 ( \23187 , \23161 );
buf \U$23177 ( \23188 , \23180 );
nand \U$23178 ( \23189 , \23187 , \23188 );
buf \U$23179 ( \23190 , \23189 );
buf \U$23180 ( \23191 , \23190 );
nand \U$23181 ( \23192 , \23186 , \23191 );
buf \U$23182 ( \23193 , \23192 );
buf \U$23183 ( \23194 , \23193 );
buf \U$23184 ( \23195 , \22280 );
not \U$23185 ( \23196 , \23195 );
buf \U$23186 ( \23197 , \22287 );
not \U$23187 ( \23198 , \23197 );
or \U$23188 ( \23199 , \23196 , \23198 );
buf \U$23189 ( \23200 , \22280 );
buf \U$23190 ( \23201 , \22287 );
or \U$23191 ( \23202 , \23200 , \23201 );
buf \U$23192 ( \23203 , \22283 );
nand \U$23193 ( \23204 , \23202 , \23203 );
buf \U$23194 ( \23205 , \23204 );
buf \U$23195 ( \23206 , \23205 );
nand \U$23196 ( \23207 , \23199 , \23206 );
buf \U$23197 ( \23208 , \23207 );
buf \U$23198 ( \23209 , \23208 );
buf \U$23199 ( \23210 , \21865 );
not \U$23200 ( \23211 , \23210 );
buf \U$23201 ( \23212 , \1822 );
not \U$23202 ( \23213 , \23212 );
or \U$23203 ( \23214 , \23211 , \23213 );
buf \U$23204 ( \23215 , \685 );
buf \U$23205 ( \23216 , RIc0d90b8_57);
buf \U$23206 ( \23217 , RIc0d9568_67);
xor \U$23207 ( \23218 , \23216 , \23217 );
buf \U$23208 ( \23219 , \23218 );
buf \U$23209 ( \23220 , \23219 );
nand \U$23210 ( \23221 , \23215 , \23220 );
buf \U$23211 ( \23222 , \23221 );
buf \U$23212 ( \23223 , \23222 );
nand \U$23213 ( \23224 , \23214 , \23223 );
buf \U$23214 ( \23225 , \23224 );
buf \U$23215 ( \23226 , RIc0d9298_61);
buf \U$23216 ( \23227 , RIc0d9478_65);
nand \U$23217 ( \23228 , \23226 , \23227 );
buf \U$23218 ( \23229 , \23228 );
xor \U$23219 ( \23230 , \23225 , \23229 );
buf \U$23220 ( \23231 , \22154 );
not \U$23221 ( \23232 , \23231 );
buf \U$23222 ( \23233 , \16402 );
not \U$23223 ( \23234 , \23233 );
or \U$23224 ( \23235 , \23232 , \23234 );
buf \U$23225 ( \23236 , \533 );
buf \U$23226 ( \23237 , RIc0d8578_33);
buf \U$23227 ( \23238 , RIc0da0a8_91);
xor \U$23228 ( \23239 , \23237 , \23238 );
buf \U$23229 ( \23240 , \23239 );
buf \U$23230 ( \23241 , \23240 );
nand \U$23231 ( \23242 , \23236 , \23241 );
buf \U$23232 ( \23243 , \23242 );
buf \U$23233 ( \23244 , \23243 );
nand \U$23234 ( \23245 , \23235 , \23244 );
buf \U$23235 ( \23246 , \23245 );
xor \U$23236 ( \23247 , \23230 , \23246 );
buf \U$23237 ( \23248 , \23247 );
buf \U$23238 ( \23249 , \21811 );
not \U$23239 ( \23250 , \23249 );
buf \U$23240 ( \23251 , \1220 );
not \U$23241 ( \23252 , \23251 );
buf \U$23242 ( \23253 , \23252 );
buf \U$23243 ( \23254 , \23253 );
not \U$23244 ( \23255 , \23254 );
or \U$23245 ( \23256 , \23250 , \23255 );
buf \U$23246 ( \23257 , \1229 );
buf \U$23247 ( \23258 , RIc0d9478_65);
buf \U$23248 ( \23259 , RIc0d91a8_59);
xor \U$23249 ( \23260 , \23258 , \23259 );
buf \U$23250 ( \23261 , \23260 );
buf \U$23251 ( \23262 , \23261 );
nand \U$23252 ( \23263 , \23257 , \23262 );
buf \U$23253 ( \23264 , \23263 );
buf \U$23254 ( \23265 , \23264 );
nand \U$23255 ( \23266 , \23256 , \23265 );
buf \U$23256 ( \23267 , \23266 );
buf \U$23257 ( \23268 , \23267 );
buf \U$23258 ( \23269 , \21992 );
not \U$23259 ( \23270 , \23269 );
buf \U$23260 ( \23271 , \13860 );
not \U$23261 ( \23272 , \23271 );
or \U$23262 ( \23273 , \23270 , \23272 );
buf \U$23263 ( \23274 , \13873 );
buf \U$23264 ( \23275 , RIc0d8398_29);
buf \U$23265 ( \23276 , RIc0da288_95);
xor \U$23266 ( \23277 , \23275 , \23276 );
buf \U$23267 ( \23278 , \23277 );
buf \U$23268 ( \23279 , \23278 );
nand \U$23269 ( \23280 , \23274 , \23279 );
buf \U$23270 ( \23281 , \23280 );
buf \U$23271 ( \23282 , \23281 );
nand \U$23272 ( \23283 , \23273 , \23282 );
buf \U$23273 ( \23284 , \23283 );
buf \U$23274 ( \23285 , \23284 );
xor \U$23275 ( \23286 , \23268 , \23285 );
buf \U$23276 ( \23287 , \21885 );
not \U$23277 ( \23288 , \23287 );
buf \U$23278 ( \23289 , \12736 );
not \U$23279 ( \23290 , \23289 );
or \U$23280 ( \23291 , \23288 , \23290 );
buf \U$23281 ( \23292 , \21880 );
xor \U$23282 ( \23293 , RIc0da738_105, RIc0d7ee8_19);
buf \U$23283 ( \23294 , \23293 );
nand \U$23284 ( \23295 , \23292 , \23294 );
buf \U$23285 ( \23296 , \23295 );
buf \U$23286 ( \23297 , \23296 );
nand \U$23287 ( \23298 , \23291 , \23297 );
buf \U$23288 ( \23299 , \23298 );
buf \U$23289 ( \23300 , \23299 );
xor \U$23290 ( \23301 , \23286 , \23300 );
buf \U$23291 ( \23302 , \23301 );
buf \U$23292 ( \23303 , \23302 );
xor \U$23293 ( \23304 , \23248 , \23303 );
buf \U$23294 ( \23305 , \22017 );
not \U$23295 ( \23306 , \23305 );
buf \U$23296 ( \23307 , \21998 );
not \U$23297 ( \23308 , \23307 );
or \U$23298 ( \23309 , \23306 , \23308 );
buf \U$23299 ( \23310 , \21998 );
buf \U$23300 ( \23311 , \22017 );
or \U$23301 ( \23312 , \23310 , \23311 );
buf \U$23302 ( \23313 , \22031 );
nand \U$23303 ( \23314 , \23312 , \23313 );
buf \U$23304 ( \23315 , \23314 );
buf \U$23305 ( \23316 , \23315 );
nand \U$23306 ( \23317 , \23309 , \23316 );
buf \U$23307 ( \23318 , \23317 );
buf \U$23308 ( \23319 , \23318 );
xor \U$23309 ( \23320 , \23304 , \23319 );
buf \U$23310 ( \23321 , \23320 );
buf \U$23311 ( \23322 , \23321 );
not \U$23312 ( \23323 , \23322 );
buf \U$23313 ( \23324 , \23323 );
buf \U$23314 ( \23325 , \23324 );
xor \U$23315 ( \23326 , \23209 , \23325 );
buf \U$23316 ( \23327 , \22229 );
not \U$23317 ( \23328 , \23327 );
buf \U$23318 ( \23329 , \15329 );
not \U$23319 ( \23330 , \23329 );
or \U$23320 ( \23331 , \23328 , \23330 );
buf \U$23321 ( \23332 , \734 );
buf \U$23322 ( \23333 , RIc0d82a8_27);
buf \U$23323 ( \23334 , RIc0da378_97);
xor \U$23324 ( \23335 , \23333 , \23334 );
buf \U$23325 ( \23336 , \23335 );
buf \U$23326 ( \23337 , \23336 );
nand \U$23327 ( \23338 , \23332 , \23337 );
buf \U$23328 ( \23339 , \23338 );
buf \U$23329 ( \23340 , \23339 );
nand \U$23330 ( \23341 , \23331 , \23340 );
buf \U$23331 ( \23342 , \23341 );
buf \U$23332 ( \23343 , \23342 );
buf \U$23333 ( \23344 , \21618 );
not \U$23334 ( \23345 , \23344 );
buf \U$23335 ( \23346 , \12870 );
not \U$23336 ( \23347 , \23346 );
or \U$23337 ( \23348 , \23345 , \23347 );
buf \U$23338 ( \23349 , \12877 );
buf \U$23339 ( \23350 , RIc0d7678_1);
buf \U$23340 ( \23351 , RIc0dafa8_123);
xor \U$23341 ( \23352 , \23350 , \23351 );
buf \U$23342 ( \23353 , \23352 );
buf \U$23343 ( \23354 , \23353 );
nand \U$23344 ( \23355 , \23349 , \23354 );
buf \U$23345 ( \23356 , \23355 );
buf \U$23346 ( \23357 , \23356 );
nand \U$23347 ( \23358 , \23348 , \23357 );
buf \U$23348 ( \23359 , \23358 );
buf \U$23349 ( \23360 , \23359 );
xor \U$23350 ( \23361 , \23343 , \23360 );
buf \U$23351 ( \23362 , \23361 );
buf \U$23352 ( \23363 , \23362 );
buf \U$23353 ( \23364 , \22196 );
not \U$23354 ( \23365 , \23364 );
buf \U$23355 ( \23366 , \2923 );
not \U$23356 ( \23367 , \23366 );
or \U$23357 ( \23368 , \23365 , \23367 );
buf \U$23358 ( \23369 , \2927 );
buf \U$23359 ( \23370 , RIc0d8ed8_53);
not \U$23360 ( \23371 , \23370 );
buf \U$23361 ( \23372 , \23371 );
and \U$23362 ( \23373 , RIc0d9748_71, \23372 );
not \U$23363 ( \23374 , RIc0d9748_71);
and \U$23364 ( \23375 , \23374 , RIc0d8ed8_53);
or \U$23365 ( \23376 , \23373 , \23375 );
buf \U$23366 ( \23377 , \23376 );
nand \U$23367 ( \23378 , \23369 , \23377 );
buf \U$23368 ( \23379 , \23378 );
buf \U$23369 ( \23380 , \23379 );
nand \U$23370 ( \23381 , \23368 , \23380 );
buf \U$23371 ( \23382 , \23381 );
buf \U$23372 ( \23383 , \23382 );
xor \U$23373 ( \23384 , \23363 , \23383 );
buf \U$23374 ( \23385 , \23384 );
buf \U$23375 ( \23386 , \23385 );
buf \U$23376 ( \23387 , \21929 );
not \U$23377 ( \23388 , \23387 );
buf \U$23378 ( \23389 , \1431 );
not \U$23379 ( \23390 , \23389 );
or \U$23380 ( \23391 , \23388 , \23390 );
buf \U$23381 ( \23392 , \14374 );
buf \U$23382 ( \23393 , RIc0d9a18_77);
buf \U$23383 ( \23394 , RIc0d8c08_47);
xor \U$23384 ( \23395 , \23393 , \23394 );
buf \U$23385 ( \23396 , \23395 );
buf \U$23386 ( \23397 , \23396 );
nand \U$23387 ( \23398 , \23392 , \23397 );
buf \U$23388 ( \23399 , \23398 );
buf \U$23389 ( \23400 , \23399 );
nand \U$23390 ( \23401 , \23391 , \23400 );
buf \U$23391 ( \23402 , \23401 );
buf \U$23392 ( \23403 , \23402 );
not \U$23393 ( \23404 , \23403 );
buf \U$23394 ( \23405 , \23404 );
buf \U$23395 ( \23406 , \23405 );
not \U$23396 ( \23407 , \23406 );
buf \U$23397 ( \23408 , \22025 );
not \U$23398 ( \23409 , \23408 );
buf \U$23399 ( \23410 , \12971 );
not \U$23400 ( \23411 , \23410 );
or \U$23401 ( \23412 , \23409 , \23411 );
buf \U$23402 ( \23413 , \13314 );
xor \U$23403 ( \23414 , RIc0daeb8_121, RIc0d7768_3);
buf \U$23404 ( \23415 , \23414 );
nand \U$23405 ( \23416 , \23413 , \23415 );
buf \U$23406 ( \23417 , \23416 );
buf \U$23407 ( \23418 , \23417 );
nand \U$23408 ( \23419 , \23412 , \23418 );
buf \U$23409 ( \23420 , \23419 );
buf \U$23410 ( \23421 , \21771 );
not \U$23411 ( \23422 , \23421 );
buf \U$23412 ( \23423 , \15397 );
not \U$23413 ( \23424 , \23423 );
or \U$23414 ( \23425 , \23422 , \23424 );
buf \U$23415 ( \23426 , \13712 );
buf \U$23416 ( \23427 , RIc0d7fd8_21);
buf \U$23417 ( \23428 , RIc0da648_103);
xor \U$23418 ( \23429 , \23427 , \23428 );
buf \U$23419 ( \23430 , \23429 );
buf \U$23420 ( \23431 , \23430 );
nand \U$23421 ( \23432 , \23426 , \23431 );
buf \U$23422 ( \23433 , \23432 );
buf \U$23423 ( \23434 , \23433 );
nand \U$23424 ( \23435 , \23425 , \23434 );
buf \U$23425 ( \23436 , \23435 );
xor \U$23426 ( \23437 , \23420 , \23436 );
buf \U$23427 ( \23438 , \23437 );
not \U$23428 ( \23439 , \23438 );
or \U$23429 ( \23440 , \23407 , \23439 );
buf \U$23430 ( \23441 , \23437 );
buf \U$23431 ( \23442 , \23405 );
or \U$23432 ( \23443 , \23441 , \23442 );
nand \U$23433 ( \23444 , \23440 , \23443 );
buf \U$23434 ( \23445 , \23444 );
buf \U$23435 ( \23446 , \23445 );
xor \U$23436 ( \23447 , \23386 , \23446 );
buf \U$23437 ( \23448 , \22137 );
not \U$23438 ( \23449 , \23448 );
buf \U$23439 ( \23450 , \1736 );
not \U$23440 ( \23451 , \23450 );
or \U$23441 ( \23452 , \23449 , \23451 );
buf \U$23442 ( \23453 , \584 );
xor \U$23443 ( \23454 , RIc0d9ce8_83, RIc0d8938_41);
buf \U$23444 ( \23455 , \23454 );
nand \U$23445 ( \23456 , \23453 , \23455 );
buf \U$23446 ( \23457 , \23456 );
buf \U$23447 ( \23458 , \23457 );
nand \U$23448 ( \23459 , \23452 , \23458 );
buf \U$23449 ( \23460 , \23459 );
buf \U$23450 ( \23461 , \21903 );
not \U$23451 ( \23462 , \23461 );
buf \U$23452 ( \23463 , \21898 );
not \U$23453 ( \23464 , \23463 );
or \U$23454 ( \23465 , \23462 , \23464 );
buf \U$23455 ( \23466 , \12342 );
buf \U$23456 ( \23467 , RIc0da828_107);
buf \U$23457 ( \23468 , RIc0d7df8_17);
xor \U$23458 ( \23469 , \23467 , \23468 );
buf \U$23459 ( \23470 , \23469 );
buf \U$23460 ( \23471 , \23470 );
nand \U$23461 ( \23472 , \23466 , \23471 );
buf \U$23462 ( \23473 , \23472 );
buf \U$23463 ( \23474 , \23473 );
nand \U$23464 ( \23475 , \23465 , \23474 );
buf \U$23465 ( \23476 , \23475 );
xor \U$23466 ( \23477 , \23460 , \23476 );
buf \U$23467 ( \23478 , \21659 );
not \U$23468 ( \23479 , \23478 );
buf \U$23469 ( \23480 , \864 );
not \U$23470 ( \23481 , \23480 );
or \U$23471 ( \23482 , \23479 , \23481 );
buf \U$23472 ( \23483 , \284 );
buf \U$23473 ( \23484 , RIc0d8fc8_55);
buf \U$23474 ( \23485 , RIc0d9658_69);
xor \U$23475 ( \23486 , \23484 , \23485 );
buf \U$23476 ( \23487 , \23486 );
buf \U$23477 ( \23488 , \23487 );
nand \U$23478 ( \23489 , \23483 , \23488 );
buf \U$23479 ( \23490 , \23489 );
buf \U$23480 ( \23491 , \23490 );
nand \U$23481 ( \23492 , \23482 , \23491 );
buf \U$23482 ( \23493 , \23492 );
xor \U$23483 ( \23494 , \23477 , \23493 );
buf \U$23484 ( \23495 , \23494 );
xor \U$23485 ( \23496 , \23447 , \23495 );
buf \U$23486 ( \23497 , \23496 );
buf \U$23487 ( \23498 , \23497 );
xnor \U$23488 ( \23499 , \23326 , \23498 );
buf \U$23489 ( \23500 , \23499 );
buf \U$23490 ( \23501 , \23500 );
not \U$23491 ( \23502 , \23501 );
buf \U$23492 ( \23503 , \23502 );
buf \U$23493 ( \23504 , \23503 );
and \U$23494 ( \23505 , \23194 , \23504 );
not \U$23495 ( \23506 , \23194 );
buf \U$23496 ( \23507 , \23500 );
and \U$23497 ( \23508 , \23506 , \23507 );
nor \U$23498 ( \23509 , \23505 , \23508 );
buf \U$23499 ( \23510 , \23509 );
buf \U$23500 ( \23511 , \23510 );
xor \U$23501 ( \23512 , \23073 , \23511 );
buf \U$23502 ( \23513 , \23512 );
buf \U$23503 ( \23514 , \23513 );
not \U$23504 ( \23515 , \23514 );
buf \U$23505 ( \23516 , \22302 );
not \U$23506 ( \23517 , \23516 );
buf \U$23507 ( \23518 , \22295 );
not \U$23508 ( \23519 , \23518 );
buf \U$23509 ( \23520 , \22288 );
not \U$23510 ( \23521 , \23520 );
and \U$23511 ( \23522 , \23519 , \23521 );
buf \U$23512 ( \23523 , \22295 );
buf \U$23513 ( \23524 , \22288 );
and \U$23514 ( \23525 , \23523 , \23524 );
nor \U$23515 ( \23526 , \23522 , \23525 );
buf \U$23516 ( \23527 , \23526 );
buf \U$23517 ( \23528 , \23527 );
not \U$23518 ( \23529 , \23528 );
or \U$23519 ( \23530 , \23517 , \23529 );
buf \U$23520 ( \23531 , \23527 );
buf \U$23521 ( \23532 , \22302 );
or \U$23522 ( \23533 , \23531 , \23532 );
nand \U$23523 ( \23534 , \23530 , \23533 );
buf \U$23524 ( \23535 , \23534 );
buf \U$23525 ( \23536 , \23535 );
buf \U$23526 ( \23537 , \21269 );
not \U$23527 ( \23538 , \23537 );
buf \U$23528 ( \23539 , \21274 );
not \U$23529 ( \23540 , \23539 );
or \U$23530 ( \23541 , \23538 , \23540 );
buf \U$23531 ( \23542 , \21274 );
buf \U$23532 ( \23543 , \21269 );
or \U$23533 ( \23544 , \23542 , \23543 );
buf \U$23534 ( \23545 , \21332 );
nand \U$23535 ( \23546 , \23544 , \23545 );
buf \U$23536 ( \23547 , \23546 );
buf \U$23537 ( \23548 , \23547 );
nand \U$23538 ( \23549 , \23541 , \23548 );
buf \U$23539 ( \23550 , \23549 );
buf \U$23540 ( \23551 , \23550 );
xor \U$23541 ( \23552 , \23536 , \23551 );
buf \U$23542 ( \23553 , \20578 );
not \U$23543 ( \23554 , \23553 );
buf \U$23544 ( \23555 , \20453 );
not \U$23545 ( \23556 , \23555 );
buf \U$23546 ( \23557 , \23556 );
buf \U$23547 ( \23558 , \23557 );
not \U$23548 ( \23559 , \23558 );
or \U$23549 ( \23560 , \23554 , \23559 );
buf \U$23550 ( \23561 , \20572 );
not \U$23551 ( \23562 , \23561 );
buf \U$23552 ( \23563 , \20453 );
not \U$23553 ( \23564 , \23563 );
or \U$23554 ( \23565 , \23562 , \23564 );
buf \U$23555 ( \23566 , \20384 );
nand \U$23556 ( \23567 , \23565 , \23566 );
buf \U$23557 ( \23568 , \23567 );
buf \U$23558 ( \23569 , \23568 );
nand \U$23559 ( \23570 , \23560 , \23569 );
buf \U$23560 ( \23571 , \23570 );
buf \U$23561 ( \23572 , \23571 );
and \U$23562 ( \23573 , \23552 , \23572 );
and \U$23563 ( \23574 , \23536 , \23551 );
or \U$23564 ( \23575 , \23573 , \23574 );
buf \U$23565 ( \23576 , \23575 );
buf \U$23566 ( \23577 , \23576 );
not \U$23567 ( \23578 , \23577 );
buf \U$23568 ( \23579 , \23578 );
buf \U$23569 ( \23580 , \23579 );
not \U$23570 ( \23581 , \23580 );
and \U$23571 ( \23582 , \23515 , \23581 );
buf \U$23572 ( \23583 , \23513 );
buf \U$23573 ( \23584 , \23579 );
and \U$23574 ( \23585 , \23583 , \23584 );
nor \U$23575 ( \23586 , \23582 , \23585 );
buf \U$23576 ( \23587 , \23586 );
buf \U$23577 ( \23588 , \23587 );
not \U$23578 ( \23589 , \23588 );
xor \U$23579 ( \23590 , \22843 , \22965 );
xor \U$23580 ( \23591 , \23590 , \22997 );
buf \U$23581 ( \23592 , \23591 );
buf \U$23582 ( \23593 , \23592 );
buf \U$23583 ( \23594 , \21221 );
buf \U$23584 ( \23595 , \21199 );
or \U$23585 ( \23596 , \23594 , \23595 );
buf \U$23586 ( \23597 , \21215 );
nand \U$23587 ( \23598 , \23596 , \23597 );
buf \U$23588 ( \23599 , \23598 );
buf \U$23589 ( \23600 , \23599 );
buf \U$23590 ( \23601 , \21221 );
buf \U$23591 ( \23602 , \21199 );
nand \U$23592 ( \23603 , \23601 , \23602 );
buf \U$23593 ( \23604 , \23603 );
buf \U$23594 ( \23605 , \23604 );
nand \U$23595 ( \23606 , \23600 , \23605 );
buf \U$23596 ( \23607 , \23606 );
buf \U$23597 ( \23608 , \23607 );
xor \U$23598 ( \23609 , \23593 , \23608 );
buf \U$23599 ( \23610 , \21336 );
not \U$23600 ( \23611 , \23610 );
buf \U$23601 ( \23612 , \21523 );
not \U$23602 ( \23613 , \23612 );
or \U$23603 ( \23614 , \23611 , \23613 );
buf \U$23604 ( \23615 , \21333 );
not \U$23605 ( \23616 , \23615 );
buf \U$23606 ( \23617 , \21520 );
not \U$23607 ( \23618 , \23617 );
or \U$23608 ( \23619 , \23616 , \23618 );
buf \U$23609 ( \23620 , \21264 );
nand \U$23610 ( \23621 , \23619 , \23620 );
buf \U$23611 ( \23622 , \23621 );
buf \U$23612 ( \23623 , \23622 );
nand \U$23613 ( \23624 , \23614 , \23623 );
buf \U$23614 ( \23625 , \23624 );
buf \U$23615 ( \23626 , \23625 );
and \U$23616 ( \23627 , \23609 , \23626 );
and \U$23617 ( \23628 , \23593 , \23608 );
or \U$23618 ( \23629 , \23627 , \23628 );
buf \U$23619 ( \23630 , \23629 );
buf \U$23620 ( \23631 , \23630 );
not \U$23621 ( \23632 , \23631 );
and \U$23622 ( \23633 , \23589 , \23632 );
buf \U$23623 ( \23634 , \23587 );
buf \U$23624 ( \23635 , \23630 );
and \U$23625 ( \23636 , \23634 , \23635 );
nor \U$23626 ( \23637 , \23633 , \23636 );
buf \U$23627 ( \23638 , \23637 );
xor \U$23628 ( \23639 , \23007 , \23638 );
xor \U$23629 ( \23640 , \23536 , \23551 );
xor \U$23630 ( \23641 , \23640 , \23572 );
buf \U$23631 ( \23642 , \23641 );
buf \U$23632 ( \23643 , \23642 );
not \U$23633 ( \23644 , \23643 );
buf \U$23634 ( \23645 , \22421 );
buf \U$23635 ( \23646 , \22438 );
xor \U$23636 ( \23647 , \23645 , \23646 );
buf \U$23637 ( \23648 , \22465 );
xor \U$23638 ( \23649 , \23647 , \23648 );
buf \U$23639 ( \23650 , \23649 );
buf \U$23640 ( \23651 , \23650 );
not \U$23641 ( \23652 , \23651 );
or \U$23642 ( \23653 , \23644 , \23652 );
xor \U$23643 ( \23654 , \23593 , \23608 );
xor \U$23644 ( \23655 , \23654 , \23626 );
buf \U$23645 ( \23656 , \23655 );
buf \U$23646 ( \23657 , \23656 );
buf \U$23647 ( \23658 , \23650 );
not \U$23648 ( \23659 , \23658 );
buf \U$23649 ( \23660 , \23642 );
not \U$23650 ( \23661 , \23660 );
buf \U$23651 ( \23662 , \23661 );
buf \U$23652 ( \23663 , \23662 );
nand \U$23653 ( \23664 , \23659 , \23663 );
buf \U$23654 ( \23665 , \23664 );
buf \U$23655 ( \23666 , \23665 );
nand \U$23656 ( \23667 , \23657 , \23666 );
buf \U$23657 ( \23668 , \23667 );
buf \U$23658 ( \23669 , \23668 );
nand \U$23659 ( \23670 , \23653 , \23669 );
buf \U$23660 ( \23671 , \23670 );
xor \U$23661 ( \23672 , \23639 , \23671 );
buf \U$23662 ( \23673 , \23672 );
xor \U$23663 ( \23674 , \20583 , \20605 );
and \U$23664 ( \23675 , \23674 , \21223 );
and \U$23665 ( \23676 , \20583 , \20605 );
or \U$23666 ( \23677 , \23675 , \23676 );
buf \U$23667 ( \23678 , \23677 );
buf \U$23668 ( \23679 , \23678 );
xor \U$23669 ( \23680 , \21250 , \21526 );
and \U$23670 ( \23681 , \23680 , \21544 );
and \U$23671 ( \23682 , \21250 , \21526 );
or \U$23672 ( \23683 , \23681 , \23682 );
buf \U$23673 ( \23684 , \23683 );
buf \U$23674 ( \23685 , \23684 );
xor \U$23675 ( \23686 , \23679 , \23685 );
buf \U$23676 ( \23687 , \23650 );
buf \U$23677 ( \23688 , \23642 );
and \U$23678 ( \23689 , \23687 , \23688 );
not \U$23679 ( \23690 , \23687 );
buf \U$23680 ( \23691 , \23662 );
and \U$23681 ( \23692 , \23690 , \23691 );
nor \U$23682 ( \23693 , \23689 , \23692 );
buf \U$23683 ( \23694 , \23693 );
buf \U$23684 ( \23695 , \23694 );
buf \U$23685 ( \23696 , \23656 );
not \U$23686 ( \23697 , \23696 );
buf \U$23687 ( \23698 , \23697 );
buf \U$23688 ( \23699 , \23698 );
and \U$23689 ( \23700 , \23695 , \23699 );
not \U$23690 ( \23701 , \23695 );
buf \U$23691 ( \23702 , \23656 );
and \U$23692 ( \23703 , \23701 , \23702 );
nor \U$23693 ( \23704 , \23700 , \23703 );
buf \U$23694 ( \23705 , \23704 );
buf \U$23695 ( \23706 , \23705 );
and \U$23696 ( \23707 , \23686 , \23706 );
and \U$23697 ( \23708 , \23679 , \23685 );
or \U$23698 ( \23709 , \23707 , \23708 );
buf \U$23699 ( \23710 , \23709 );
buf \U$23700 ( \23711 , \23710 );
nand \U$23701 ( \23712 , \23673 , \23711 );
buf \U$23702 ( \23713 , \23712 );
buf \U$23703 ( \23714 , \23713 );
xor \U$23704 ( \23715 , \23679 , \23685 );
xor \U$23705 ( \23716 , \23715 , \23706 );
buf \U$23706 ( \23717 , \23716 );
buf \U$23707 ( \23718 , \23717 );
xor \U$23708 ( \23719 , \21226 , \21235 );
and \U$23709 ( \23720 , \23719 , \21547 );
and \U$23710 ( \23721 , \21226 , \21235 );
or \U$23711 ( \23722 , \23720 , \23721 );
buf \U$23712 ( \23723 , \23722 );
buf \U$23713 ( \23724 , \23723 );
nand \U$23714 ( \23725 , \23718 , \23724 );
buf \U$23715 ( \23726 , \23725 );
buf \U$23716 ( \23727 , \23726 );
and \U$23717 ( \23728 , \23714 , \23727 );
buf \U$23718 ( \23729 , \23728 );
buf \U$23719 ( \23730 , \23729 );
not \U$23720 ( \23731 , \23730 );
or \U$23721 ( \23732 , \21576 , \23731 );
not \U$23722 ( \23733 , \23713 );
buf \U$23723 ( \23734 , \23723 );
buf \U$23724 ( \23735 , \23717 );
nor \U$23725 ( \23736 , \23734 , \23735 );
buf \U$23726 ( \23737 , \23736 );
not \U$23727 ( \23738 , \23737 );
or \U$23728 ( \23739 , \23733 , \23738 );
buf \U$23729 ( \23740 , \23672 );
not \U$23730 ( \23741 , \23740 );
buf \U$23731 ( \23742 , \23741 );
buf \U$23732 ( \23743 , \23742 );
buf \U$23733 ( \23744 , \23710 );
not \U$23734 ( \23745 , \23744 );
buf \U$23735 ( \23746 , \23745 );
buf \U$23736 ( \23747 , \23746 );
nand \U$23737 ( \23748 , \23743 , \23747 );
buf \U$23738 ( \23749 , \23748 );
nand \U$23739 ( \23750 , \23739 , \23749 );
buf \U$23740 ( \23751 , \23750 );
not \U$23741 ( \23752 , \23751 );
buf \U$23742 ( \23753 , \23752 );
buf \U$23743 ( \23754 , \23753 );
nand \U$23744 ( \23755 , \23732 , \23754 );
buf \U$23745 ( \23756 , \23755 );
buf \U$23746 ( \23757 , \23756 );
xor \U$23747 ( \23758 , \22495 , \22667 );
and \U$23748 ( \23759 , \23758 , \22815 );
and \U$23749 ( \23760 , \22495 , \22667 );
or \U$23750 ( \23761 , \23759 , \23760 );
buf \U$23751 ( \23762 , \23761 );
buf \U$23752 ( \23763 , \23762 );
not \U$23753 ( \23764 , \23763 );
xor \U$23754 ( \23765 , \22774 , \22791 );
and \U$23755 ( \23766 , \23765 , \22811 );
and \U$23756 ( \23767 , \22774 , \22791 );
or \U$23757 ( \23768 , \23766 , \23767 );
buf \U$23758 ( \23769 , \23768 );
buf \U$23759 ( \23770 , \23769 );
xor \U$23760 ( \23771 , \23136 , \23142 );
and \U$23761 ( \23772 , \23771 , \23149 );
and \U$23762 ( \23773 , \23136 , \23142 );
or \U$23763 ( \23774 , \23772 , \23773 );
buf \U$23764 ( \23775 , \23774 );
buf \U$23765 ( \23776 , \23775 );
xor \U$23766 ( \23777 , \23770 , \23776 );
xor \U$23767 ( \23778 , \21801 , \21854 );
and \U$23768 ( \23779 , \23778 , \21915 );
and \U$23769 ( \23780 , \21801 , \21854 );
or \U$23770 ( \23781 , \23779 , \23780 );
buf \U$23771 ( \23782 , \23781 );
buf \U$23772 ( \23783 , \23782 );
xor \U$23773 ( \23784 , \23777 , \23783 );
buf \U$23774 ( \23785 , \23784 );
buf \U$23775 ( \23786 , \23324 );
not \U$23776 ( \23787 , \23786 );
buf \U$23777 ( \23788 , \23208 );
not \U$23778 ( \23789 , \23788 );
or \U$23779 ( \23790 , \23787 , \23789 );
buf \U$23780 ( \23791 , \23497 );
buf \U$23781 ( \23792 , \23208 );
not \U$23782 ( \23793 , \23792 );
buf \U$23783 ( \23794 , \23321 );
nand \U$23784 ( \23795 , \23793 , \23794 );
buf \U$23785 ( \23796 , \23795 );
buf \U$23786 ( \23797 , \23796 );
nand \U$23787 ( \23798 , \23791 , \23797 );
buf \U$23788 ( \23799 , \23798 );
buf \U$23789 ( \23800 , \23799 );
nand \U$23790 ( \23801 , \23790 , \23800 );
buf \U$23791 ( \23802 , \23801 );
xor \U$23792 ( \23803 , \23785 , \23802 );
buf \U$23793 ( \23804 , \23803 );
not \U$23794 ( \23805 , \23804 );
buf \U$23795 ( \23806 , \23805 );
buf \U$23796 ( \23807 , \23806 );
not \U$23797 ( \23808 , \23807 );
or \U$23798 ( \23809 , \23764 , \23808 );
buf \U$23799 ( \23810 , \23762 );
not \U$23800 ( \23811 , \23810 );
buf \U$23801 ( \23812 , \23803 );
nand \U$23802 ( \23813 , \23811 , \23812 );
buf \U$23803 ( \23814 , \23813 );
buf \U$23804 ( \23815 , \23814 );
nand \U$23805 ( \23816 , \23809 , \23815 );
buf \U$23806 ( \23817 , \23816 );
buf \U$23807 ( \23818 , \23817 );
xor \U$23808 ( \23819 , \22818 , \22824 );
and \U$23809 ( \23820 , \23819 , \23002 );
and \U$23810 ( \23821 , \22818 , \22824 );
or \U$23811 ( \23822 , \23820 , \23821 );
buf \U$23812 ( \23823 , \23822 );
buf \U$23814 ( \23824 , \23823 );
xor \U$23815 ( \23825 , \23818 , \23824 );
buf \U$23816 ( \23826 , \23454 );
not \U$23817 ( \23827 , \23826 );
buf \U$23818 ( \23828 , \573 );
not \U$23819 ( \23829 , \23828 );
or \U$23820 ( \23830 , \23827 , \23829 );
buf \U$23821 ( \23831 , \993 );
xor \U$23822 ( \23832 , RIc0d9ce8_83, RIc0d88c0_40);
buf \U$23823 ( \23833 , \23832 );
nand \U$23824 ( \23834 , \23831 , \23833 );
buf \U$23825 ( \23835 , \23834 );
buf \U$23826 ( \23836 , \23835 );
nand \U$23827 ( \23837 , \23830 , \23836 );
buf \U$23828 ( \23838 , \23837 );
buf \U$23829 ( \23839 , \23838 );
buf \U$23830 ( \23840 , \23396 );
not \U$23831 ( \23841 , \23840 );
buf \U$23832 ( \23842 , \1183 );
not \U$23833 ( \23843 , \23842 );
or \U$23834 ( \23844 , \23841 , \23843 );
buf \U$23835 ( \23845 , \14374 );
buf \U$23836 ( \23846 , RIc0d8b90_46);
buf \U$23837 ( \23847 , RIc0d9a18_77);
xor \U$23838 ( \23848 , \23846 , \23847 );
buf \U$23839 ( \23849 , \23848 );
buf \U$23840 ( \23850 , \23849 );
nand \U$23841 ( \23851 , \23845 , \23850 );
buf \U$23842 ( \23852 , \23851 );
buf \U$23843 ( \23853 , \23852 );
nand \U$23844 ( \23854 , \23844 , \23853 );
buf \U$23845 ( \23855 , \23854 );
buf \U$23846 ( \23856 , \23855 );
xor \U$23847 ( \23857 , \23839 , \23856 );
buf \U$23848 ( \23858 , \22526 );
not \U$23849 ( \23859 , \23858 );
buf \U$23850 ( \23860 , \14210 );
not \U$23851 ( \23861 , \23860 );
or \U$23852 ( \23862 , \23859 , \23861 );
buf \U$23853 ( \23863 , \20211 );
buf \U$23854 ( \23864 , RIc0d7c90_14);
buf \U$23855 ( \23865 , RIc0da918_109);
xor \U$23856 ( \23866 , \23864 , \23865 );
buf \U$23857 ( \23867 , \23866 );
buf \U$23858 ( \23868 , \23867 );
nand \U$23859 ( \23869 , \23863 , \23868 );
buf \U$23860 ( \23870 , \23869 );
buf \U$23861 ( \23871 , \23870 );
nand \U$23862 ( \23872 , \23862 , \23871 );
buf \U$23863 ( \23873 , \23872 );
buf \U$23864 ( \23874 , \23873 );
xor \U$23865 ( \23875 , \23857 , \23874 );
buf \U$23866 ( \23876 , \23875 );
buf \U$23867 ( \23877 , \23876 );
not \U$23868 ( \23878 , \23877 );
buf \U$23869 ( \23879 , \23878 );
buf \U$23870 ( \23880 , \23879 );
not \U$23871 ( \23881 , \23880 );
buf \U$23872 ( \23882 , \23240 );
not \U$23873 ( \23883 , \23882 );
buf \U$23874 ( \23884 , \16402 );
not \U$23875 ( \23885 , \23884 );
or \U$23876 ( \23886 , \23883 , \23885 );
buf \U$23877 ( \23887 , \1933 );
buf \U$23878 ( \23888 , RIc0d8500_32);
buf \U$23879 ( \23889 , RIc0da0a8_91);
xor \U$23880 ( \23890 , \23888 , \23889 );
buf \U$23881 ( \23891 , \23890 );
buf \U$23882 ( \23892 , \23891 );
nand \U$23883 ( \23893 , \23887 , \23892 );
buf \U$23884 ( \23894 , \23893 );
buf \U$23885 ( \23895 , \23894 );
nand \U$23886 ( \23896 , \23886 , \23895 );
buf \U$23887 ( \23897 , \23896 );
buf \U$23888 ( \23898 , \23336 );
not \U$23889 ( \23899 , \23898 );
buf \U$23890 ( \23900 , \16086 );
not \U$23891 ( \23901 , \23900 );
or \U$23892 ( \23902 , \23899 , \23901 );
buf \U$23893 ( \23903 , \734 );
buf \U$23894 ( \23904 , RIc0d8230_26);
buf \U$23895 ( \23905 , RIc0da378_97);
xor \U$23896 ( \23906 , \23904 , \23905 );
buf \U$23897 ( \23907 , \23906 );
buf \U$23898 ( \23908 , \23907 );
nand \U$23899 ( \23909 , \23903 , \23908 );
buf \U$23900 ( \23910 , \23909 );
buf \U$23901 ( \23911 , \23910 );
nand \U$23902 ( \23912 , \23902 , \23911 );
buf \U$23903 ( \23913 , \23912 );
xor \U$23904 ( \23914 , \23897 , \23913 );
buf \U$23905 ( \23915 , \23261 );
not \U$23906 ( \23916 , \23915 );
buf \U$23907 ( \23917 , \3781 );
not \U$23908 ( \23918 , \23917 );
or \U$23909 ( \23919 , \23916 , \23918 );
buf \U$23910 ( \23920 , \1229 );
buf \U$23911 ( \23921 , RIc0d9478_65);
buf \U$23912 ( \23922 , RIc0d9130_58);
xor \U$23913 ( \23923 , \23921 , \23922 );
buf \U$23914 ( \23924 , \23923 );
buf \U$23915 ( \23925 , \23924 );
nand \U$23916 ( \23926 , \23920 , \23925 );
buf \U$23917 ( \23927 , \23926 );
buf \U$23918 ( \23928 , \23927 );
nand \U$23919 ( \23929 , \23919 , \23928 );
buf \U$23920 ( \23930 , \23929 );
xnor \U$23921 ( \23931 , \23914 , \23930 );
buf \U$23922 ( \23932 , \23931 );
not \U$23923 ( \23933 , \23932 );
buf \U$23924 ( \23934 , \23933 );
buf \U$23925 ( \23935 , \23934 );
not \U$23926 ( \23936 , \23935 );
or \U$23927 ( \23937 , \23881 , \23936 );
buf \U$23928 ( \23938 , \23876 );
buf \U$23929 ( \23939 , \23931 );
nand \U$23930 ( \23940 , \23938 , \23939 );
buf \U$23931 ( \23941 , \23940 );
buf \U$23932 ( \23942 , \23941 );
nand \U$23933 ( \23943 , \23937 , \23942 );
buf \U$23934 ( \23944 , \23943 );
buf \U$23935 ( \23945 , \23944 );
buf \U$23936 ( \23946 , \2815 );
buf \U$23937 ( \23947 , \23376 );
not \U$23938 ( \23948 , \23947 );
buf \U$23939 ( \23949 , \23948 );
buf \U$23940 ( \23950 , \23949 );
or \U$23941 ( \23951 , \23946 , \23950 );
buf \U$23942 ( \23952 , \2927 );
buf \U$23943 ( \23953 , RIc0d9748_71);
buf \U$23944 ( \23954 , RIc0d8e60_52);
xor \U$23945 ( \23955 , \23953 , \23954 );
buf \U$23946 ( \23956 , \23955 );
buf \U$23947 ( \23957 , \23956 );
nand \U$23948 ( \23958 , \23952 , \23957 );
buf \U$23949 ( \23959 , \23958 );
buf \U$23950 ( \23960 , \23959 );
nand \U$23951 ( \23961 , \23951 , \23960 );
buf \U$23952 ( \23962 , \23961 );
buf \U$23953 ( \23963 , \22716 );
not \U$23954 ( \23964 , \23963 );
buf \U$23955 ( \23965 , \21461 );
not \U$23956 ( \23966 , \23965 );
or \U$23957 ( \23967 , \23964 , \23966 );
buf \U$23958 ( \23968 , RIc0d8140_24);
buf \U$23959 ( \23969 , RIc0da468_99);
xnor \U$23960 ( \23970 , \23968 , \23969 );
buf \U$23961 ( \23971 , \23970 );
buf \U$23962 ( \23972 , \23971 );
not \U$23963 ( \23973 , \23972 );
buf \U$23964 ( \23974 , \14140 );
nand \U$23965 ( \23975 , \23973 , \23974 );
buf \U$23966 ( \23976 , \23975 );
buf \U$23967 ( \23977 , \23976 );
nand \U$23968 ( \23978 , \23967 , \23977 );
buf \U$23969 ( \23979 , \23978 );
xor \U$23970 ( \23980 , \23962 , \23979 );
buf \U$23971 ( \23981 , \22803 );
not \U$23972 ( \23982 , \23981 );
buf \U$23973 ( \23983 , \13178 );
not \U$23974 ( \23984 , \23983 );
buf \U$23975 ( \23985 , \23984 );
buf \U$23976 ( \23986 , \23985 );
not \U$23977 ( \23987 , \23986 );
or \U$23978 ( \23988 , \23982 , \23987 );
buf \U$23979 ( \23989 , \13953 );
buf \U$23980 ( \23990 , RIc0dadc8_119);
buf \U$23981 ( \23991 , RIc0d77e0_4);
xor \U$23982 ( \23992 , \23990 , \23991 );
buf \U$23983 ( \23993 , \23992 );
buf \U$23984 ( \23994 , \23993 );
nand \U$23985 ( \23995 , \23989 , \23994 );
buf \U$23986 ( \23996 , \23995 );
buf \U$23987 ( \23997 , \23996 );
nand \U$23988 ( \23998 , \23988 , \23997 );
buf \U$23989 ( \23999 , \23998 );
xor \U$23990 ( \24000 , \23980 , \23999 );
buf \U$23991 ( \24001 , \24000 );
and \U$23992 ( \24002 , \23945 , \24001 );
not \U$23993 ( \24003 , \23945 );
buf \U$23994 ( \24004 , \24000 );
not \U$23995 ( \24005 , \24004 );
buf \U$23996 ( \24006 , \24005 );
buf \U$23997 ( \24007 , \24006 );
and \U$23998 ( \24008 , \24003 , \24007 );
nor \U$23999 ( \24009 , \24002 , \24008 );
buf \U$24000 ( \24010 , \24009 );
buf \U$24003 ( \24011 , \24010 );
buf \U$24004 ( \24012 , \24011 );
not \U$24005 ( \24013 , \24012 );
buf \U$24006 ( \24014 , \22725 );
not \U$24007 ( \24015 , \24014 );
buf \U$24008 ( \24016 , \24015 );
buf \U$24009 ( \24017 , \24016 );
not \U$24010 ( \24018 , \24017 );
buf \U$24011 ( \24019 , \22813 );
not \U$24012 ( \24020 , \24019 );
or \U$24013 ( \24021 , \24018 , \24020 );
buf \U$24014 ( \24022 , \24016 );
buf \U$24015 ( \24023 , \22813 );
or \U$24016 ( \24024 , \24022 , \24023 );
buf \U$24017 ( \24025 , \22772 );
nand \U$24018 ( \24026 , \24024 , \24025 );
buf \U$24019 ( \24027 , \24026 );
buf \U$24020 ( \24028 , \24027 );
nand \U$24021 ( \24029 , \24021 , \24028 );
buf \U$24022 ( \24030 , \24029 );
buf \U$24023 ( \24031 , \24030 );
buf \U$24024 ( \24032 , \22761 );
not \U$24025 ( \24033 , \24032 );
buf \U$24026 ( \24034 , \12361 );
not \U$24027 ( \24035 , \24034 );
or \U$24028 ( \24036 , \24033 , \24035 );
buf \U$24029 ( \24037 , \1025 );
buf \U$24030 ( \24038 , RIc0d8aa0_44);
buf \U$24031 ( \24039 , RIc0d9b08_79);
xor \U$24032 ( \24040 , \24038 , \24039 );
buf \U$24033 ( \24041 , \24040 );
buf \U$24034 ( \24042 , \24041 );
nand \U$24035 ( \24043 , \24037 , \24042 );
buf \U$24036 ( \24044 , \24043 );
buf \U$24037 ( \24045 , \24044 );
nand \U$24038 ( \24046 , \24036 , \24045 );
buf \U$24039 ( \24047 , \24046 );
buf \U$24040 ( \24048 , \24047 );
buf \U$24041 ( \24049 , \22656 );
not \U$24042 ( \24050 , \24049 );
buf \U$24043 ( \24051 , \2607 );
not \U$24044 ( \24052 , \24051 );
or \U$24045 ( \24053 , \24050 , \24052 );
buf \U$24046 ( \24054 , \816 );
buf \U$24047 ( \24055 , RIc0d86e0_36);
buf \U$24048 ( \24056 , RIc0d9ec8_87);
xor \U$24049 ( \24057 , \24055 , \24056 );
buf \U$24050 ( \24058 , \24057 );
buf \U$24051 ( \24059 , \24058 );
nand \U$24052 ( \24060 , \24054 , \24059 );
buf \U$24053 ( \24061 , \24060 );
buf \U$24054 ( \24062 , \24061 );
nand \U$24055 ( \24063 , \24053 , \24062 );
buf \U$24056 ( \24064 , \24063 );
buf \U$24057 ( \24065 , \24064 );
xor \U$24058 ( \24066 , \24048 , \24065 );
buf \U$24059 ( \24067 , \22606 );
not \U$24060 ( \24068 , \24067 );
buf \U$24061 ( \24069 , \24068 );
buf \U$24062 ( \24070 , \24069 );
not \U$24063 ( \24071 , \24070 );
buf \U$24064 ( \24072 , \14186 );
not \U$24065 ( \24073 , \24072 );
or \U$24066 ( \24074 , \24071 , \24073 );
buf \U$24067 ( \24075 , \12303 );
buf \U$24068 ( \24076 , RIc0d79c0_8);
buf \U$24069 ( \24077 , RIc0dabe8_115);
xor \U$24070 ( \24078 , \24076 , \24077 );
buf \U$24071 ( \24079 , \24078 );
buf \U$24072 ( \24080 , \24079 );
nand \U$24073 ( \24081 , \24075 , \24080 );
buf \U$24074 ( \24082 , \24081 );
buf \U$24075 ( \24083 , \24082 );
nand \U$24076 ( \24084 , \24074 , \24083 );
buf \U$24077 ( \24085 , \24084 );
buf \U$24078 ( \24086 , \24085 );
xor \U$24079 ( \24087 , \24066 , \24086 );
buf \U$24080 ( \24088 , \24087 );
buf \U$24081 ( \24089 , \24088 );
buf \U$24082 ( \24090 , \23487 );
not \U$24083 ( \24091 , \24090 );
buf \U$24084 ( \24092 , \13332 );
not \U$24085 ( \24093 , \24092 );
or \U$24086 ( \24094 , \24091 , \24093 );
buf \U$24087 ( \24095 , \284 );
buf \U$24088 ( \24096 , RIc0d8f50_54);
buf \U$24089 ( \24097 , RIc0d9658_69);
xor \U$24090 ( \24098 , \24096 , \24097 );
buf \U$24091 ( \24099 , \24098 );
buf \U$24092 ( \24100 , \24099 );
nand \U$24093 ( \24101 , \24095 , \24100 );
buf \U$24094 ( \24102 , \24101 );
buf \U$24095 ( \24103 , \24102 );
nand \U$24096 ( \24104 , \24094 , \24103 );
buf \U$24097 ( \24105 , \24104 );
buf \U$24098 ( \24106 , \24105 );
not \U$24099 ( \24107 , \24106 );
buf \U$24100 ( \24108 , \22562 );
not \U$24101 ( \24109 , \24108 );
buf \U$24102 ( \24110 , \2766 );
not \U$24103 ( \24111 , \24110 );
or \U$24104 ( \24112 , \24109 , \24111 );
buf \U$24105 ( \24113 , \1078 );
buf \U$24106 ( \24114 , RIc0d89b0_42);
buf \U$24107 ( \24115 , RIc0d9bf8_81);
xor \U$24108 ( \24116 , \24114 , \24115 );
buf \U$24109 ( \24117 , \24116 );
buf \U$24110 ( \24118 , \24117 );
nand \U$24111 ( \24119 , \24113 , \24118 );
buf \U$24112 ( \24120 , \24119 );
buf \U$24113 ( \24121 , \24120 );
nand \U$24114 ( \24122 , \24112 , \24121 );
buf \U$24115 ( \24123 , \24122 );
buf \U$24116 ( \24124 , \24123 );
not \U$24117 ( \24125 , \24124 );
buf \U$24118 ( \24126 , \24125 );
buf \U$24119 ( \24127 , \24126 );
not \U$24120 ( \24128 , \24127 );
or \U$24121 ( \24129 , \24107 , \24128 );
buf \U$24122 ( \24130 , \24105 );
not \U$24123 ( \24131 , \24130 );
buf \U$24124 ( \24132 , \24131 );
buf \U$24125 ( \24133 , \24132 );
buf \U$24126 ( \24134 , \24123 );
nand \U$24127 ( \24135 , \24133 , \24134 );
buf \U$24128 ( \24136 , \24135 );
buf \U$24129 ( \24137 , \24136 );
nand \U$24130 ( \24138 , \24129 , \24137 );
buf \U$24131 ( \24139 , \24138 );
buf \U$24132 ( \24140 , \24139 );
buf \U$24133 ( \24141 , \23278 );
not \U$24134 ( \24142 , \24141 );
buf \U$24135 ( \24143 , \3714 );
not \U$24136 ( \24144 , \24143 );
or \U$24137 ( \24145 , \24142 , \24144 );
buf \U$24138 ( \24146 , \344 );
buf \U$24139 ( \24147 , RIc0d8320_28);
buf \U$24140 ( \24148 , RIc0da288_95);
xor \U$24141 ( \24149 , \24147 , \24148 );
buf \U$24142 ( \24150 , \24149 );
buf \U$24143 ( \24151 , \24150 );
nand \U$24144 ( \24152 , \24146 , \24151 );
buf \U$24145 ( \24153 , \24152 );
buf \U$24146 ( \24154 , \24153 );
nand \U$24147 ( \24155 , \24145 , \24154 );
buf \U$24148 ( \24156 , \24155 );
buf \U$24149 ( \24157 , \24156 );
and \U$24150 ( \24158 , \24140 , \24157 );
not \U$24151 ( \24159 , \24140 );
buf \U$24152 ( \24160 , \24156 );
not \U$24153 ( \24161 , \24160 );
buf \U$24154 ( \24162 , \24161 );
buf \U$24155 ( \24163 , \24162 );
and \U$24156 ( \24164 , \24159 , \24163 );
nor \U$24157 ( \24165 , \24158 , \24164 );
buf \U$24158 ( \24166 , \24165 );
buf \U$24159 ( \24167 , \24166 );
xor \U$24160 ( \24168 , \24089 , \24167 );
buf \U$24161 ( \24169 , \22543 );
not \U$24162 ( \24170 , \24169 );
buf \U$24163 ( \24171 , \1389 );
not \U$24164 ( \24172 , \24171 );
or \U$24165 ( \24173 , \24170 , \24172 );
buf \U$24166 ( \24174 , \921 );
buf \U$24167 ( \24175 , RIc0d9dd8_85);
buf \U$24168 ( \24176 , RIc0d87d0_38);
xor \U$24169 ( \24177 , \24175 , \24176 );
buf \U$24170 ( \24178 , \24177 );
buf \U$24171 ( \24179 , \24178 );
nand \U$24172 ( \24180 , \24174 , \24179 );
buf \U$24173 ( \24181 , \24180 );
buf \U$24174 ( \24182 , \24181 );
nand \U$24175 ( \24183 , \24173 , \24182 );
buf \U$24176 ( \24184 , \24183 );
buf \U$24177 ( \24185 , \24184 );
buf \U$24178 ( \24186 , \22784 );
not \U$24179 ( \24187 , \24186 );
buf \U$24180 ( \24188 , \437 );
not \U$24181 ( \24189 , \24188 );
or \U$24182 ( \24190 , \24187 , \24189 );
buf \U$24183 ( \24191 , RIc0d9fb8_89);
buf \U$24184 ( \24192 , RIc0d85f0_34);
xnor \U$24185 ( \24193 , \24191 , \24192 );
buf \U$24186 ( \24194 , \24193 );
buf \U$24187 ( \24195 , \24194 );
not \U$24188 ( \24196 , \24195 );
buf \U$24189 ( \24197 , \16477 );
nand \U$24190 ( \24198 , \24196 , \24197 );
buf \U$24191 ( \24199 , \24198 );
buf \U$24192 ( \24200 , \24199 );
nand \U$24193 ( \24201 , \24190 , \24200 );
buf \U$24194 ( \24202 , \24201 );
buf \U$24195 ( \24203 , \24202 );
xor \U$24196 ( \24204 , \24185 , \24203 );
buf \U$24197 ( \24205 , \22695 );
not \U$24198 ( \24206 , \24205 );
buf \U$24199 ( \24207 , \16656 );
not \U$24200 ( \24208 , \24207 );
or \U$24201 ( \24209 , \24206 , \24208 );
buf \U$24202 ( \24210 , \16662 );
buf \U$24203 ( \24211 , RIc0d7ab0_10);
buf \U$24204 ( \24212 , RIc0daaf8_113);
xor \U$24205 ( \24213 , \24211 , \24212 );
buf \U$24206 ( \24214 , \24213 );
buf \U$24207 ( \24215 , \24214 );
nand \U$24208 ( \24216 , \24210 , \24215 );
buf \U$24209 ( \24217 , \24216 );
buf \U$24210 ( \24218 , \24217 );
nand \U$24211 ( \24219 , \24209 , \24218 );
buf \U$24212 ( \24220 , \24219 );
buf \U$24213 ( \24221 , \24220 );
xor \U$24214 ( \24222 , \24204 , \24221 );
buf \U$24215 ( \24223 , \24222 );
buf \U$24216 ( \24224 , \24223 );
xor \U$24217 ( \24225 , \24168 , \24224 );
buf \U$24218 ( \24226 , \24225 );
buf \U$24219 ( \24227 , \24226 );
xnor \U$24220 ( \24228 , \24031 , \24227 );
buf \U$24221 ( \24229 , \24228 );
buf \U$24222 ( \24230 , \24229 );
not \U$24223 ( \24231 , \24230 );
or \U$24224 ( \24232 , \24013 , \24231 );
buf \U$24225 ( \24233 , \24229 );
buf \U$24226 ( \24234 , \24011 );
or \U$24227 ( \24235 , \24233 , \24234 );
nand \U$24228 ( \24236 , \24232 , \24235 );
buf \U$24229 ( \24237 , \24236 );
buf \U$24230 ( \24238 , \24237 );
xor \U$24231 ( \24239 , \23013 , \23044 );
and \U$24232 ( \24240 , \24239 , \23063 );
and \U$24233 ( \24241 , \23013 , \23044 );
or \U$24234 ( \24242 , \24240 , \24241 );
buf \U$24235 ( \24243 , \24242 );
buf \U$24236 ( \24244 , \24243 );
xor \U$24237 ( \24245 , \24238 , \24244 );
xor \U$24238 ( \24246 , \23019 , \23034 );
and \U$24239 ( \24247 , \24246 , \23041 );
and \U$24240 ( \24248 , \23019 , \23034 );
or \U$24241 ( \24249 , \24247 , \24248 );
buf \U$24242 ( \24250 , \24249 );
buf \U$24243 ( \24251 , \24250 );
buf \U$24244 ( \24252 , \23110 );
not \U$24245 ( \24253 , \24252 );
buf \U$24246 ( \24254 , \23104 );
not \U$24247 ( \24255 , \24254 );
or \U$24248 ( \24256 , \24253 , \24255 );
buf \U$24249 ( \24257 , \23116 );
not \U$24250 ( \24258 , \24257 );
buf \U$24251 ( \24259 , \23104 );
not \U$24252 ( \24260 , \24259 );
buf \U$24253 ( \24261 , \24260 );
buf \U$24254 ( \24262 , \24261 );
not \U$24255 ( \24263 , \24262 );
or \U$24256 ( \24264 , \24258 , \24263 );
buf \U$24257 ( \24265 , \23151 );
nand \U$24258 ( \24266 , \24264 , \24265 );
buf \U$24259 ( \24267 , \24266 );
buf \U$24260 ( \24268 , \24267 );
nand \U$24261 ( \24269 , \24256 , \24268 );
buf \U$24262 ( \24270 , \24269 );
buf \U$24263 ( \24271 , \24270 );
xor \U$24264 ( \24272 , \24251 , \24271 );
xor \U$24265 ( \24273 , \21744 , \21918 );
and \U$24266 ( \24274 , \24273 , \22038 );
and \U$24267 ( \24275 , \21744 , \21918 );
or \U$24268 ( \24276 , \24274 , \24275 );
buf \U$24269 ( \24277 , \24276 );
buf \U$24270 ( \24278 , \24277 );
xor \U$24271 ( \24279 , \24272 , \24278 );
buf \U$24272 ( \24280 , \24279 );
buf \U$24273 ( \24281 , \24280 );
xor \U$24274 ( \24282 , \24245 , \24281 );
buf \U$24275 ( \24283 , \24282 );
buf \U$24276 ( \24284 , \24283 );
xor \U$24277 ( \24285 , \23825 , \24284 );
buf \U$24278 ( \24286 , \24285 );
buf \U$24279 ( \24287 , \24286 );
xor \U$24280 ( \24288 , \23066 , \23072 );
and \U$24281 ( \24289 , \24288 , \23511 );
and \U$24282 ( \24290 , \23066 , \23072 );
or \U$24283 ( \24291 , \24289 , \24290 );
buf \U$24284 ( \24292 , \24291 );
buf \U$24285 ( \24293 , \24292 );
buf \U$24286 ( \24294 , \23180 );
buf \U$24287 ( \24295 , \23164 );
nor \U$24288 ( \24296 , \24294 , \24295 );
buf \U$24289 ( \24297 , \24296 );
buf \U$24290 ( \24298 , \24297 );
buf \U$24291 ( \24299 , \23500 );
or \U$24292 ( \24300 , \24298 , \24299 );
buf \U$24293 ( \24301 , \23164 );
buf \U$24294 ( \24302 , \23180 );
nand \U$24295 ( \24303 , \24301 , \24302 );
buf \U$24296 ( \24304 , \24303 );
buf \U$24297 ( \24305 , \24304 );
nand \U$24298 ( \24306 , \24300 , \24305 );
buf \U$24299 ( \24307 , \24306 );
buf \U$24300 ( \24308 , \24307 );
buf \U$24301 ( \24309 , \22040 );
not \U$24302 ( \24310 , \24309 );
buf \U$24303 ( \24311 , \24310 );
buf \U$24304 ( \24312 , \24311 );
buf \U$24305 ( \24313 , \22309 );
nand \U$24306 ( \24314 , \24312 , \24313 );
buf \U$24307 ( \24315 , \24314 );
buf \U$24308 ( \24316 , \24315 );
buf \U$24309 ( \24317 , \22116 );
nand \U$24310 ( \24318 , \24316 , \24317 );
buf \U$24311 ( \24319 , \24318 );
buf \U$24312 ( \24320 , \24319 );
buf \U$24313 ( \24321 , \22040 );
buf \U$24314 ( \24322 , \22306 );
nand \U$24315 ( \24323 , \24321 , \24322 );
buf \U$24316 ( \24324 , \24323 );
buf \U$24317 ( \24325 , \24324 );
nand \U$24318 ( \24326 , \24320 , \24325 );
buf \U$24319 ( \24327 , \24326 );
buf \U$24320 ( \24328 , \24327 );
xor \U$24321 ( \24329 , \24308 , \24328 );
xor \U$24322 ( \24330 , \23082 , \23095 );
and \U$24323 ( \24331 , \24330 , \23102 );
and \U$24324 ( \24332 , \23082 , \23095 );
or \U$24325 ( \24333 , \24331 , \24332 );
buf \U$24326 ( \24334 , \24333 );
buf \U$24327 ( \24335 , \24334 );
not \U$24328 ( \24336 , \22514 );
not \U$24329 ( \24337 , \22549 );
or \U$24330 ( \24338 , \24336 , \24337 );
buf \U$24331 ( \24339 , \22514 );
buf \U$24332 ( \24340 , \22549 );
or \U$24333 ( \24341 , \24339 , \24340 );
buf \U$24334 ( \24342 , \22532 );
nand \U$24335 ( \24343 , \24341 , \24342 );
buf \U$24336 ( \24344 , \24343 );
nand \U$24337 ( \24345 , \24338 , \24344 );
buf \U$24338 ( \24346 , \24345 );
xor \U$24339 ( \24347 , \22577 , \22591 );
and \U$24340 ( \24348 , \24347 , \22611 );
and \U$24341 ( \24349 , \22577 , \22591 );
or \U$24342 ( \24350 , \24348 , \24349 );
buf \U$24343 ( \24351 , \24350 );
buf \U$24344 ( \24352 , \24351 );
xor \U$24345 ( \24353 , \24346 , \24352 );
and \U$24346 ( \24354 , \21808 , \21809 );
buf \U$24347 ( \24355 , \24354 );
buf \U$24348 ( \24356 , \24355 );
buf \U$24349 ( \24357 , \23430 );
not \U$24350 ( \24358 , \24357 );
buf \U$24351 ( \24359 , \18220 );
not \U$24352 ( \24360 , \24359 );
or \U$24353 ( \24361 , \24358 , \24360 );
buf \U$24354 ( \24362 , \13048 );
buf \U$24355 ( \24363 , RIc0d7f60_20);
buf \U$24356 ( \24364 , RIc0da648_103);
xor \U$24357 ( \24365 , \24363 , \24364 );
buf \U$24358 ( \24366 , \24365 );
buf \U$24359 ( \24367 , \24366 );
nand \U$24360 ( \24368 , \24362 , \24367 );
buf \U$24361 ( \24369 , \24368 );
buf \U$24362 ( \24370 , \24369 );
nand \U$24363 ( \24371 , \24361 , \24370 );
buf \U$24364 ( \24372 , \24371 );
buf \U$24365 ( \24373 , \24372 );
xor \U$24366 ( \24374 , \24356 , \24373 );
buf \U$24367 ( \24375 , \22735 );
not \U$24368 ( \24376 , \24375 );
buf \U$24369 ( \24377 , \12529 );
not \U$24370 ( \24378 , \24377 );
or \U$24371 ( \24379 , \24376 , \24378 );
buf \U$24372 ( \24380 , \14106 );
xor \U$24373 ( \24381 , RIc0daa08_111, RIc0d7ba0_12);
buf \U$24374 ( \24382 , \24381 );
nand \U$24375 ( \24383 , \24380 , \24382 );
buf \U$24376 ( \24384 , \24383 );
buf \U$24377 ( \24385 , \24384 );
nand \U$24378 ( \24386 , \24379 , \24385 );
buf \U$24379 ( \24387 , \24386 );
buf \U$24380 ( \24388 , \24387 );
xor \U$24381 ( \24389 , \24374 , \24388 );
buf \U$24382 ( \24390 , \24389 );
buf \U$24383 ( \24391 , \24390 );
xor \U$24384 ( \24392 , \24353 , \24391 );
buf \U$24385 ( \24393 , \24392 );
buf \U$24386 ( \24394 , \24393 );
xor \U$24387 ( \24395 , \24335 , \24394 );
buf \U$24388 ( \24396 , \22768 );
not \U$24389 ( \24397 , \24396 );
buf \U$24390 ( \24398 , \22741 );
not \U$24391 ( \24399 , \24398 );
or \U$24392 ( \24400 , \24397 , \24399 );
buf \U$24393 ( \24401 , \22765 );
not \U$24394 ( \24402 , \24401 );
buf \U$24395 ( \24403 , \22741 );
not \U$24396 ( \24404 , \24403 );
buf \U$24397 ( \24405 , \24404 );
buf \U$24398 ( \24406 , \24405 );
not \U$24399 ( \24407 , \24406 );
or \U$24400 ( \24408 , \24402 , \24407 );
buf \U$24401 ( \24409 , \22752 );
nand \U$24402 ( \24410 , \24408 , \24409 );
buf \U$24403 ( \24411 , \24410 );
buf \U$24404 ( \24412 , \24411 );
nand \U$24405 ( \24413 , \24400 , \24412 );
buf \U$24406 ( \24414 , \24413 );
buf \U$24407 ( \24415 , \24414 );
not \U$24408 ( \24416 , \24415 );
buf \U$24409 ( \24417 , \22684 );
not \U$24410 ( \24418 , \24417 );
buf \U$24411 ( \24419 , \24418 );
buf \U$24412 ( \24420 , \24419 );
not \U$24413 ( \24421 , \24420 );
buf \U$24414 ( \24422 , \22704 );
not \U$24415 ( \24423 , \24422 );
or \U$24416 ( \24424 , \24421 , \24423 );
buf \U$24417 ( \24425 , \22722 );
nand \U$24418 ( \24426 , \24424 , \24425 );
buf \U$24419 ( \24427 , \24426 );
buf \U$24420 ( \24428 , \24427 );
buf \U$24421 ( \24429 , \22701 );
buf \U$24422 ( \24430 , \22684 );
nand \U$24423 ( \24431 , \24429 , \24430 );
buf \U$24424 ( \24432 , \24431 );
buf \U$24425 ( \24433 , \24432 );
nand \U$24426 ( \24434 , \24428 , \24433 );
buf \U$24427 ( \24435 , \24434 );
buf \U$24428 ( \24436 , \24435 );
not \U$24429 ( \24437 , \24436 );
buf \U$24430 ( \24438 , \24437 );
buf \U$24431 ( \24439 , \24438 );
not \U$24432 ( \24440 , \24439 );
or \U$24433 ( \24441 , \24416 , \24440 );
buf \U$24434 ( \24442 , \24414 );
not \U$24435 ( \24443 , \24442 );
buf \U$24436 ( \24444 , \24435 );
nand \U$24437 ( \24445 , \24443 , \24444 );
buf \U$24438 ( \24446 , \24445 );
buf \U$24439 ( \24447 , \24446 );
nand \U$24440 ( \24448 , \24441 , \24447 );
buf \U$24441 ( \24449 , \24448 );
buf \U$24442 ( \24450 , \24449 );
buf \U$24443 ( \24451 , \22645 );
buf \U$24444 ( \24452 , \22662 );
or \U$24445 ( \24453 , \24451 , \24452 );
buf \U$24446 ( \24454 , \22628 );
nand \U$24447 ( \24455 , \24453 , \24454 );
buf \U$24448 ( \24456 , \24455 );
buf \U$24449 ( \24457 , \24456 );
buf \U$24450 ( \24458 , \22645 );
buf \U$24451 ( \24459 , \22662 );
nand \U$24452 ( \24460 , \24458 , \24459 );
buf \U$24453 ( \24461 , \24460 );
buf \U$24454 ( \24462 , \24461 );
nand \U$24455 ( \24463 , \24457 , \24462 );
buf \U$24456 ( \24464 , \24463 );
buf \U$24459 ( \24465 , \24464 );
buf \U$24460 ( \24466 , \24465 );
and \U$24461 ( \24467 , \24450 , \24466 );
not \U$24462 ( \24468 , \24450 );
buf \U$24463 ( \24469 , \24465 );
not \U$24464 ( \24470 , \24469 );
buf \U$24465 ( \24471 , \24470 );
buf \U$24466 ( \24472 , \24471 );
and \U$24467 ( \24473 , \24468 , \24472 );
nor \U$24468 ( \24474 , \24467 , \24473 );
buf \U$24469 ( \24475 , \24474 );
buf \U$24470 ( \24476 , \24475 );
xor \U$24471 ( \24477 , \24395 , \24476 );
buf \U$24472 ( \24478 , \24477 );
buf \U$24473 ( \24479 , \24478 );
buf \U$24474 ( \24480 , \23353 );
not \U$24475 ( \24481 , \24480 );
buf \U$24476 ( \24482 , \14982 );
not \U$24477 ( \24483 , \24482 );
or \U$24478 ( \24484 , \24481 , \24483 );
buf \U$24479 ( \24485 , \16692 );
buf \U$24480 ( \24486 , RIc0dafa8_123);
nand \U$24481 ( \24487 , \24485 , \24486 );
buf \U$24482 ( \24488 , \24487 );
buf \U$24483 ( \24489 , \24488 );
nand \U$24484 ( \24490 , \24484 , \24489 );
buf \U$24485 ( \24491 , \24490 );
buf \U$24486 ( \24492 , \24491 );
not \U$24487 ( \24493 , \24492 );
buf \U$24488 ( \24494 , \24493 );
buf \U$24489 ( \24495 , \24494 );
buf \U$24490 ( \24496 , \23229 );
not \U$24491 ( \24497 , \24496 );
buf \U$24492 ( \24498 , \23225 );
not \U$24493 ( \24499 , \24498 );
buf \U$24494 ( \24500 , \24499 );
buf \U$24495 ( \24501 , \24500 );
not \U$24496 ( \24502 , \24501 );
or \U$24497 ( \24503 , \24497 , \24502 );
buf \U$24498 ( \24504 , \23246 );
nand \U$24499 ( \24505 , \24503 , \24504 );
buf \U$24500 ( \24506 , \24505 );
buf \U$24501 ( \24507 , \24506 );
buf \U$24502 ( \24508 , \23229 );
not \U$24503 ( \24509 , \24508 );
buf \U$24504 ( \24510 , \23225 );
nand \U$24505 ( \24511 , \24509 , \24510 );
buf \U$24506 ( \24512 , \24511 );
buf \U$24507 ( \24513 , \24512 );
nand \U$24508 ( \24514 , \24507 , \24513 );
buf \U$24509 ( \24515 , \24514 );
buf \U$24510 ( \24516 , \24515 );
xor \U$24511 ( \24517 , \24495 , \24516 );
buf \U$24512 ( \24518 , \23436 );
buf \U$24513 ( \24519 , \23402 );
or \U$24514 ( \24520 , \24518 , \24519 );
buf \U$24515 ( \24521 , \23420 );
nand \U$24516 ( \24522 , \24520 , \24521 );
buf \U$24517 ( \24523 , \24522 );
buf \U$24518 ( \24524 , \24523 );
buf \U$24519 ( \24525 , \23436 );
buf \U$24520 ( \24526 , \23402 );
nand \U$24521 ( \24527 , \24525 , \24526 );
buf \U$24522 ( \24528 , \24527 );
buf \U$24523 ( \24529 , \24528 );
nand \U$24524 ( \24530 , \24524 , \24529 );
buf \U$24525 ( \24531 , \24530 );
buf \U$24526 ( \24532 , \24531 );
xor \U$24527 ( \24533 , \24517 , \24532 );
buf \U$24528 ( \24534 , \24533 );
buf \U$24529 ( \24535 , \24534 );
buf \U$24530 ( \24536 , \23382 );
not \U$24531 ( \24537 , \24536 );
buf \U$24532 ( \24538 , \23359 );
not \U$24533 ( \24539 , \24538 );
or \U$24534 ( \24540 , \24537 , \24539 );
buf \U$24535 ( \24541 , \23359 );
buf \U$24536 ( \24542 , \23382 );
or \U$24537 ( \24543 , \24541 , \24542 );
buf \U$24538 ( \24544 , \23342 );
nand \U$24539 ( \24545 , \24543 , \24544 );
buf \U$24540 ( \24546 , \24545 );
buf \U$24541 ( \24547 , \24546 );
nand \U$24542 ( \24548 , \24540 , \24547 );
buf \U$24543 ( \24549 , \24548 );
buf \U$24544 ( \24550 , \24549 );
xor \U$24545 ( \24551 , \23268 , \23285 );
and \U$24546 ( \24552 , \24551 , \23300 );
and \U$24547 ( \24553 , \23268 , \23285 );
or \U$24548 ( \24554 , \24552 , \24553 );
buf \U$24549 ( \24555 , \24554 );
buf \U$24550 ( \24556 , \24555 );
xor \U$24551 ( \24557 , \24550 , \24556 );
buf \U$24552 ( \24558 , \23493 );
not \U$24553 ( \24559 , \24558 );
buf \U$24554 ( \24560 , \23476 );
not \U$24555 ( \24561 , \24560 );
or \U$24556 ( \24562 , \24559 , \24561 );
buf \U$24557 ( \24563 , \23476 );
buf \U$24558 ( \24564 , \23493 );
or \U$24559 ( \24565 , \24563 , \24564 );
buf \U$24560 ( \24566 , \23460 );
nand \U$24561 ( \24567 , \24565 , \24566 );
buf \U$24562 ( \24568 , \24567 );
buf \U$24563 ( \24569 , \24568 );
nand \U$24564 ( \24570 , \24562 , \24569 );
buf \U$24565 ( \24571 , \24570 );
buf \U$24566 ( \24572 , \24571 );
xor \U$24567 ( \24573 , \24557 , \24572 );
buf \U$24568 ( \24574 , \24573 );
buf \U$24569 ( \24575 , \24574 );
xor \U$24570 ( \24576 , \24535 , \24575 );
xor \U$24571 ( \24577 , \23386 , \23446 );
and \U$24572 ( \24578 , \24577 , \23495 );
and \U$24573 ( \24579 , \23386 , \23446 );
or \U$24574 ( \24580 , \24578 , \24579 );
buf \U$24575 ( \24581 , \24580 );
buf \U$24576 ( \24582 , \24581 );
xor \U$24577 ( \24583 , \24576 , \24582 );
buf \U$24578 ( \24584 , \24583 );
buf \U$24579 ( \24585 , \24584 );
xor \U$24580 ( \24586 , \24479 , \24585 );
buf \U$24581 ( \24587 , \23247 );
not \U$24582 ( \24588 , \24587 );
buf \U$24583 ( \24589 , \23318 );
not \U$24584 ( \24590 , \24589 );
buf \U$24585 ( \24591 , \24590 );
buf \U$24586 ( \24592 , \24591 );
not \U$24587 ( \24593 , \24592 );
or \U$24588 ( \24594 , \24588 , \24593 );
buf \U$24589 ( \24595 , \23302 );
nand \U$24590 ( \24596 , \24594 , \24595 );
buf \U$24591 ( \24597 , \24596 );
buf \U$24592 ( \24598 , \24597 );
buf \U$24593 ( \24599 , \23247 );
not \U$24594 ( \24600 , \24599 );
buf \U$24595 ( \24601 , \23318 );
nand \U$24596 ( \24602 , \24600 , \24601 );
buf \U$24597 ( \24603 , \24602 );
buf \U$24598 ( \24604 , \24603 );
nand \U$24599 ( \24605 , \24598 , \24604 );
buf \U$24600 ( \24606 , \24605 );
buf \U$24601 ( \24607 , \24606 );
xor \U$24602 ( \24608 , \22561 , \22614 );
and \U$24603 ( \24609 , \24608 , \22664 );
and \U$24604 ( \24610 , \22561 , \22614 );
or \U$24605 ( \24611 , \24609 , \24610 );
buf \U$24606 ( \24612 , \24611 );
buf \U$24607 ( \24613 , \24612 );
xor \U$24608 ( \24614 , \24607 , \24613 );
buf \U$24609 ( \24615 , \22639 );
not \U$24610 ( \24616 , \24615 );
buf \U$24611 ( \24617 , \3534 );
not \U$24612 ( \24618 , \24617 );
or \U$24613 ( \24619 , \24616 , \24618 );
buf \U$24614 ( \24620 , \12839 );
buf \U$24615 ( \24621 , RIc0da558_101);
buf \U$24616 ( \24622 , RIc0d8050_22);
xor \U$24617 ( \24623 , \24621 , \24622 );
buf \U$24618 ( \24624 , \24623 );
buf \U$24619 ( \24625 , \24624 );
nand \U$24620 ( \24626 , \24620 , \24625 );
buf \U$24621 ( \24627 , \24626 );
buf \U$24622 ( \24628 , \24627 );
nand \U$24623 ( \24629 , \24619 , \24628 );
buf \U$24624 ( \24630 , \24629 );
buf \U$24625 ( \24631 , \22584 );
not \U$24626 ( \24632 , \24631 );
buf \U$24627 ( \24633 , \12923 );
not \U$24628 ( \24634 , \24633 );
or \U$24629 ( \24635 , \24632 , \24634 );
buf \U$24630 ( \24636 , \12936 );
buf \U$24631 ( \24637 , RIc0dacd8_117);
buf \U$24632 ( \24638 , RIc0d78d0_6);
xor \U$24633 ( \24639 , \24637 , \24638 );
buf \U$24634 ( \24640 , \24639 );
buf \U$24635 ( \24641 , \24640 );
nand \U$24636 ( \24642 , \24636 , \24641 );
buf \U$24637 ( \24643 , \24642 );
buf \U$24638 ( \24644 , \24643 );
nand \U$24639 ( \24645 , \24635 , \24644 );
buf \U$24640 ( \24646 , \24645 );
xor \U$24641 ( \24647 , \24630 , \24646 );
buf \U$24642 ( \24648 , \24647 );
buf \U$24643 ( \24649 , \22508 );
not \U$24644 ( \24650 , \24649 );
buf \U$24645 ( \24651 , \2124 );
not \U$24646 ( \24652 , \24651 );
or \U$24647 ( \24653 , \24650 , \24652 );
buf \U$24648 ( \24654 , \1143 );
xor \U$24649 ( \24655 , RIc0d9928_75, RIc0d8c80_48);
buf \U$24650 ( \24656 , \24655 );
nand \U$24651 ( \24657 , \24654 , \24656 );
buf \U$24652 ( \24658 , \24657 );
buf \U$24653 ( \24659 , \24658 );
nand \U$24654 ( \24660 , \24653 , \24659 );
buf \U$24655 ( \24661 , \24660 );
buf \U$24656 ( \24662 , \24661 );
xnor \U$24657 ( \24663 , \24648 , \24662 );
buf \U$24658 ( \24664 , \24663 );
buf \U$24659 ( \24665 , \24664 );
not \U$24660 ( \24666 , \24665 );
buf \U$24661 ( \24667 , \24666 );
buf \U$24662 ( \24668 , \23414 );
not \U$24663 ( \24669 , \24668 );
buf \U$24664 ( \24670 , \12968 );
not \U$24665 ( \24671 , \24670 );
buf \U$24666 ( \24672 , \24671 );
buf \U$24667 ( \24673 , \24672 );
not \U$24668 ( \24674 , \24673 );
or \U$24669 ( \24675 , \24669 , \24674 );
buf \U$24670 ( \24676 , \16386 );
buf \U$24671 ( \24677 , RIc0d76f0_2);
buf \U$24672 ( \24678 , RIc0daeb8_121);
xor \U$24673 ( \24679 , \24677 , \24678 );
buf \U$24674 ( \24680 , \24679 );
buf \U$24675 ( \24681 , \24680 );
nand \U$24676 ( \24682 , \24676 , \24681 );
buf \U$24677 ( \24683 , \24682 );
buf \U$24678 ( \24684 , \24683 );
nand \U$24679 ( \24685 , \24675 , \24684 );
buf \U$24680 ( \24686 , \24685 );
buf \U$24681 ( \24687 , \24686 );
not \U$24682 ( \24688 , \24687 );
buf \U$24683 ( \24689 , \24688 );
buf \U$24684 ( \24690 , \24689 );
not \U$24685 ( \24691 , \24690 );
buf \U$24686 ( \24692 , \22622 );
not \U$24687 ( \24693 , \24692 );
buf \U$24688 ( \24694 , \1901 );
not \U$24689 ( \24695 , \24694 );
or \U$24690 ( \24696 , \24693 , \24695 );
buf \U$24691 ( \24697 , \481 );
xor \U$24692 ( \24698 , RIc0da198_93, RIc0d8410_30);
buf \U$24693 ( \24699 , \24698 );
nand \U$24694 ( \24700 , \24697 , \24699 );
buf \U$24695 ( \24701 , \24700 );
buf \U$24696 ( \24702 , \24701 );
nand \U$24697 ( \24703 , \24696 , \24702 );
buf \U$24698 ( \24704 , \24703 );
buf \U$24699 ( \24705 , \24704 );
not \U$24700 ( \24706 , \24705 );
or \U$24701 ( \24707 , \24691 , \24706 );
buf \U$24702 ( \24708 , \24686 );
buf \U$24703 ( \24709 , \24704 );
not \U$24704 ( \24710 , \24709 );
buf \U$24705 ( \24711 , \24710 );
buf \U$24706 ( \24712 , \24711 );
nand \U$24707 ( \24713 , \24708 , \24712 );
buf \U$24708 ( \24714 , \24713 );
buf \U$24709 ( \24715 , \24714 );
nand \U$24710 ( \24716 , \24707 , \24715 );
buf \U$24711 ( \24717 , \24716 );
buf \U$24712 ( \24718 , \24717 );
buf \U$24713 ( \24719 , \22678 );
not \U$24714 ( \24720 , \24719 );
buf \U$24715 ( \24721 , \776 );
not \U$24716 ( \24722 , \24721 );
or \U$24717 ( \24723 , \24720 , \24722 );
buf \U$24718 ( \24724 , \791 );
xor \U$24719 ( \24725 , RIc0d9838_73, RIc0d8d70_50);
buf \U$24720 ( \24726 , \24725 );
nand \U$24721 ( \24727 , \24724 , \24726 );
buf \U$24722 ( \24728 , \24727 );
buf \U$24723 ( \24729 , \24728 );
nand \U$24724 ( \24730 , \24723 , \24729 );
buf \U$24725 ( \24731 , \24730 );
buf \U$24726 ( \24732 , \24731 );
not \U$24727 ( \24733 , \24732 );
buf \U$24728 ( \24734 , \24733 );
buf \U$24729 ( \24735 , \24734 );
and \U$24730 ( \24736 , \24718 , \24735 );
not \U$24731 ( \24737 , \24718 );
buf \U$24732 ( \24738 , \24731 );
and \U$24733 ( \24739 , \24737 , \24738 );
nor \U$24734 ( \24740 , \24736 , \24739 );
buf \U$24735 ( \24741 , \24740 );
buf \U$24736 ( \24742 , \24741 );
not \U$24737 ( \24743 , \24742 );
buf \U$24738 ( \24744 , \23293 );
not \U$24739 ( \24745 , \24744 );
buf \U$24740 ( \24746 , \16014 );
not \U$24741 ( \24747 , \24746 );
or \U$24742 ( \24748 , \24745 , \24747 );
buf \U$24743 ( \24749 , \12744 );
xor \U$24744 ( \24750 , RIc0da738_105, RIc0d7e70_18);
buf \U$24745 ( \24751 , \24750 );
nand \U$24746 ( \24752 , \24749 , \24751 );
buf \U$24747 ( \24753 , \24752 );
buf \U$24748 ( \24754 , \24753 );
nand \U$24749 ( \24755 , \24748 , \24754 );
buf \U$24750 ( \24756 , \24755 );
buf \U$24751 ( \24757 , \24756 );
not \U$24752 ( \24758 , \24757 );
buf \U$24753 ( \24759 , \23470 );
not \U$24754 ( \24760 , \24759 );
buf \U$24755 ( \24761 , \17595 );
not \U$24756 ( \24762 , \24761 );
or \U$24757 ( \24763 , \24760 , \24762 );
buf \U$24758 ( \24764 , \12342 );
buf \U$24759 ( \24765 , RIc0da828_107);
buf \U$24760 ( \24766 , RIc0d7d80_16);
xor \U$24761 ( \24767 , \24765 , \24766 );
buf \U$24762 ( \24768 , \24767 );
buf \U$24763 ( \24769 , \24768 );
nand \U$24764 ( \24770 , \24764 , \24769 );
buf \U$24765 ( \24771 , \24770 );
buf \U$24766 ( \24772 , \24771 );
nand \U$24767 ( \24773 , \24763 , \24772 );
buf \U$24768 ( \24774 , \24773 );
buf \U$24769 ( \24775 , \24774 );
not \U$24770 ( \24776 , \24775 );
buf \U$24771 ( \24777 , \24776 );
buf \U$24772 ( \24778 , \24777 );
not \U$24773 ( \24779 , \24778 );
or \U$24774 ( \24780 , \24758 , \24779 );
buf \U$24775 ( \24781 , \24756 );
not \U$24776 ( \24782 , \24781 );
buf \U$24777 ( \24783 , \24774 );
nand \U$24778 ( \24784 , \24782 , \24783 );
buf \U$24779 ( \24785 , \24784 );
buf \U$24780 ( \24786 , \24785 );
nand \U$24781 ( \24787 , \24780 , \24786 );
buf \U$24782 ( \24788 , \24787 );
buf \U$24783 ( \24789 , \24788 );
buf \U$24784 ( \24790 , \23219 );
not \U$24785 ( \24791 , \24790 );
buf \U$24786 ( \24792 , \1414 );
not \U$24787 ( \24793 , \24792 );
or \U$24788 ( \24794 , \24791 , \24793 );
buf \U$24789 ( \24795 , \686 );
xor \U$24790 ( \24796 , RIc0d9568_67, RIc0d9040_56);
buf \U$24791 ( \24797 , \24796 );
nand \U$24792 ( \24798 , \24795 , \24797 );
buf \U$24793 ( \24799 , \24798 );
buf \U$24794 ( \24800 , \24799 );
nand \U$24795 ( \24801 , \24794 , \24800 );
buf \U$24796 ( \24802 , \24801 );
buf \U$24797 ( \24803 , \24802 );
and \U$24798 ( \24804 , \24789 , \24803 );
not \U$24799 ( \24805 , \24789 );
buf \U$24800 ( \24806 , \24802 );
not \U$24801 ( \24807 , \24806 );
buf \U$24802 ( \24808 , \24807 );
buf \U$24803 ( \24809 , \24808 );
and \U$24804 ( \24810 , \24805 , \24809 );
nor \U$24805 ( \24811 , \24804 , \24810 );
buf \U$24806 ( \24812 , \24811 );
buf \U$24807 ( \24813 , \24812 );
not \U$24808 ( \24814 , \24813 );
or \U$24809 ( \24815 , \24743 , \24814 );
buf \U$24810 ( \24816 , \24812 );
buf \U$24811 ( \24817 , \24741 );
or \U$24812 ( \24818 , \24816 , \24817 );
nand \U$24813 ( \24819 , \24815 , \24818 );
buf \U$24814 ( \24820 , \24819 );
xor \U$24815 ( \24821 , \24667 , \24820 );
buf \U$24816 ( \24822 , \24821 );
xor \U$24817 ( \24823 , \24614 , \24822 );
buf \U$24818 ( \24824 , \24823 );
buf \U$24819 ( \24825 , \24824 );
xor \U$24820 ( \24826 , \24586 , \24825 );
buf \U$24821 ( \24827 , \24826 );
buf \U$24822 ( \24828 , \24827 );
xor \U$24823 ( \24829 , \24329 , \24828 );
buf \U$24824 ( \24830 , \24829 );
buf \U$24825 ( \24831 , \24830 );
xor \U$24826 ( \24832 , \24293 , \24831 );
xor \U$24827 ( \24833 , \22320 , \22477 );
and \U$24828 ( \24834 , \24833 , \23005 );
and \U$24829 ( \24835 , \22320 , \22477 );
or \U$24830 ( \24836 , \24834 , \24835 );
buf \U$24831 ( \24837 , \24836 );
buf \U$24832 ( \24838 , \24837 );
xor \U$24833 ( \24839 , \24832 , \24838 );
buf \U$24834 ( \24840 , \24839 );
buf \U$24835 ( \24841 , \24840 );
xor \U$24836 ( \24842 , \24287 , \24841 );
buf \U$24837 ( \24843 , \23579 );
not \U$24838 ( \24844 , \24843 );
buf \U$24839 ( \24845 , \24844 );
buf \U$24840 ( \24846 , \24845 );
not \U$24841 ( \24847 , \24846 );
buf \U$24842 ( \24848 , \23630 );
not \U$24843 ( \24849 , \24848 );
or \U$24844 ( \24850 , \24847 , \24849 );
buf \U$24845 ( \24851 , \23630 );
buf \U$24846 ( \24852 , \24845 );
or \U$24847 ( \24853 , \24851 , \24852 );
buf \U$24848 ( \24854 , \23513 );
nand \U$24849 ( \24855 , \24853 , \24854 );
buf \U$24850 ( \24856 , \24855 );
buf \U$24851 ( \24857 , \24856 );
nand \U$24852 ( \24858 , \24850 , \24857 );
buf \U$24853 ( \24859 , \24858 );
buf \U$24854 ( \24860 , \24859 );
xnor \U$24855 ( \24861 , \24842 , \24860 );
buf \U$24856 ( \24862 , \24861 );
buf \U$24857 ( \24863 , \24862 );
buf \U$24858 ( \24864 , \23007 );
not \U$24859 ( \24865 , \24864 );
buf \U$24860 ( \24866 , \24865 );
buf \U$24861 ( \24867 , \24866 );
not \U$24862 ( \24868 , \24867 );
buf \U$24863 ( \24869 , \23671 );
not \U$24864 ( \24870 , \24869 );
buf \U$24865 ( \24871 , \24870 );
buf \U$24866 ( \24872 , \24871 );
not \U$24867 ( \24873 , \24872 );
or \U$24868 ( \24874 , \24868 , \24873 );
buf \U$24869 ( \24875 , \23638 );
not \U$24870 ( \24876 , \24875 );
buf \U$24871 ( \24877 , \24876 );
buf \U$24872 ( \24878 , \24877 );
nand \U$24873 ( \24879 , \24874 , \24878 );
buf \U$24874 ( \24880 , \24879 );
buf \U$24875 ( \24881 , \24880 );
buf \U$24876 ( \24882 , \23671 );
buf \U$24877 ( \24883 , \23007 );
nand \U$24878 ( \24884 , \24882 , \24883 );
buf \U$24879 ( \24885 , \24884 );
buf \U$24880 ( \24886 , \24885 );
and \U$24881 ( \24887 , \24881 , \24886 );
buf \U$24882 ( \24888 , \24887 );
buf \U$24883 ( \24889 , \24888 );
nand \U$24884 ( \24890 , \24863 , \24889 );
buf \U$24885 ( \24891 , \24890 );
buf \U$24886 ( \24892 , \24891 );
buf \U$24887 ( \24893 , \24286 );
not \U$24888 ( \24894 , \24893 );
buf \U$24889 ( \24895 , \24894 );
buf \U$24890 ( \24896 , \24895 );
not \U$24891 ( \24897 , \24896 );
buf \U$24892 ( \24898 , \24840 );
not \U$24893 ( \24899 , \24898 );
buf \U$24894 ( \24900 , \24899 );
buf \U$24895 ( \24901 , \24900 );
not \U$24896 ( \24902 , \24901 );
or \U$24897 ( \24903 , \24897 , \24902 );
buf \U$24898 ( \24904 , \24859 );
nand \U$24899 ( \24905 , \24903 , \24904 );
buf \U$24900 ( \24906 , \24905 );
buf \U$24901 ( \24907 , \24906 );
buf \U$24902 ( \24908 , \24840 );
buf \U$24903 ( \24909 , \24286 );
nand \U$24904 ( \24910 , \24908 , \24909 );
buf \U$24905 ( \24911 , \24910 );
buf \U$24906 ( \24912 , \24911 );
nand \U$24907 ( \24913 , \24907 , \24912 );
buf \U$24908 ( \24914 , \24913 );
buf \U$24909 ( \24915 , \24914 );
not \U$24910 ( \24916 , \24915 );
xor \U$24911 ( \24917 , \24607 , \24613 );
and \U$24912 ( \24918 , \24917 , \24822 );
and \U$24913 ( \24919 , \24607 , \24613 );
or \U$24914 ( \24920 , \24918 , \24919 );
buf \U$24915 ( \24921 , \24920 );
buf \U$24918 ( \24922 , \24921 );
buf \U$24919 ( \24923 , \24922 );
not \U$24920 ( \24924 , \24923 );
not \U$24921 ( \24925 , \23934 );
not \U$24922 ( \24926 , \23876 );
or \U$24923 ( \24927 , \24925 , \24926 );
not \U$24924 ( \24928 , \23879 );
not \U$24925 ( \24929 , \23931 );
or \U$24926 ( \24930 , \24928 , \24929 );
nand \U$24927 ( \24931 , \24930 , \24000 );
nand \U$24928 ( \24932 , \24927 , \24931 );
buf \U$24929 ( \24933 , \24932 );
buf \U$24930 ( \24934 , \24646 );
not \U$24931 ( \24935 , \24934 );
buf \U$24932 ( \24936 , \24661 );
not \U$24933 ( \24937 , \24936 );
or \U$24934 ( \24938 , \24935 , \24937 );
buf \U$24935 ( \24939 , \24646 );
buf \U$24936 ( \24940 , \24661 );
or \U$24937 ( \24941 , \24939 , \24940 );
buf \U$24938 ( \24942 , \24630 );
nand \U$24939 ( \24943 , \24941 , \24942 );
buf \U$24940 ( \24944 , \24943 );
buf \U$24941 ( \24945 , \24944 );
nand \U$24942 ( \24946 , \24938 , \24945 );
buf \U$24943 ( \24947 , \24946 );
xor \U$24944 ( \24948 , \24048 , \24065 );
and \U$24945 ( \24949 , \24948 , \24086 );
and \U$24946 ( \24950 , \24048 , \24065 );
or \U$24947 ( \24951 , \24949 , \24950 );
buf \U$24948 ( \24952 , \24951 );
xor \U$24949 ( \24953 , \24947 , \24952 );
buf \U$24950 ( \24954 , \24953 );
buf \U$24951 ( \24955 , \23930 );
buf \U$24952 ( \24956 , \23897 );
or \U$24953 ( \24957 , \24955 , \24956 );
buf \U$24954 ( \24958 , \23913 );
nand \U$24955 ( \24959 , \24957 , \24958 );
buf \U$24956 ( \24960 , \24959 );
buf \U$24957 ( \24961 , \24960 );
buf \U$24958 ( \24962 , \23897 );
buf \U$24959 ( \24963 , \23930 );
nand \U$24960 ( \24964 , \24962 , \24963 );
buf \U$24961 ( \24965 , \24964 );
buf \U$24962 ( \24966 , \24965 );
nand \U$24963 ( \24967 , \24961 , \24966 );
buf \U$24964 ( \24968 , \24967 );
buf \U$24965 ( \24969 , \24968 );
xor \U$24966 ( \24970 , \24954 , \24969 );
buf \U$24967 ( \24971 , \24970 );
buf \U$24968 ( \24972 , \24971 );
xor \U$24969 ( \24973 , \24933 , \24972 );
buf \U$24970 ( \24974 , \23962 );
not \U$24971 ( \24975 , \24974 );
buf \U$24972 ( \24976 , \23999 );
not \U$24973 ( \24977 , \24976 );
or \U$24974 ( \24978 , \24975 , \24977 );
buf \U$24975 ( \24979 , \23999 );
buf \U$24976 ( \24980 , \23962 );
or \U$24977 ( \24981 , \24979 , \24980 );
buf \U$24978 ( \24982 , \23979 );
nand \U$24979 ( \24983 , \24981 , \24982 );
buf \U$24980 ( \24984 , \24983 );
buf \U$24981 ( \24985 , \24984 );
nand \U$24982 ( \24986 , \24978 , \24985 );
buf \U$24983 ( \24987 , \24986 );
xor \U$24984 ( \24988 , \23839 , \23856 );
and \U$24985 ( \24989 , \24988 , \23874 );
and \U$24986 ( \24990 , \23839 , \23856 );
or \U$24987 ( \24991 , \24989 , \24990 );
buf \U$24988 ( \24992 , \24991 );
xor \U$24989 ( \24993 , \24987 , \24992 );
xor \U$24990 ( \24994 , \24185 , \24203 );
and \U$24991 ( \24995 , \24994 , \24221 );
and \U$24992 ( \24996 , \24185 , \24203 );
or \U$24993 ( \24997 , \24995 , \24996 );
buf \U$24994 ( \24998 , \24997 );
xor \U$24995 ( \24999 , \24993 , \24998 );
buf \U$24996 ( \25000 , \24999 );
xor \U$24997 ( \25001 , \24973 , \25000 );
buf \U$24998 ( \25002 , \25001 );
buf \U$24999 ( \25003 , \25002 );
xor \U$25000 ( \25004 , \24346 , \24352 );
and \U$25001 ( \25005 , \25004 , \24391 );
and \U$25002 ( \25006 , \24346 , \24352 );
or \U$25003 ( \25007 , \25005 , \25006 );
buf \U$25004 ( \25008 , \25007 );
buf \U$25005 ( \25009 , \25008 );
buf \U$25006 ( \25010 , \24741 );
not \U$25007 ( \25011 , \25010 );
buf \U$25008 ( \25012 , \25011 );
buf \U$25009 ( \25013 , \25012 );
not \U$25010 ( \25014 , \25013 );
buf \U$25011 ( \25015 , \24667 );
not \U$25012 ( \25016 , \25015 );
or \U$25013 ( \25017 , \25014 , \25016 );
buf \U$25014 ( \25018 , \24664 );
not \U$25015 ( \25019 , \25018 );
buf \U$25016 ( \25020 , \24741 );
not \U$25017 ( \25021 , \25020 );
or \U$25018 ( \25022 , \25019 , \25021 );
buf \U$25019 ( \25023 , \24812 );
nand \U$25020 ( \25024 , \25022 , \25023 );
buf \U$25021 ( \25025 , \25024 );
buf \U$25022 ( \25026 , \25025 );
nand \U$25023 ( \25027 , \25017 , \25026 );
buf \U$25024 ( \25028 , \25027 );
buf \U$25025 ( \25029 , \25028 );
xor \U$25026 ( \25030 , \25009 , \25029 );
xor \U$25027 ( \25031 , \24089 , \24167 );
and \U$25028 ( \25032 , \25031 , \24224 );
and \U$25029 ( \25033 , \24089 , \24167 );
or \U$25030 ( \25034 , \25032 , \25033 );
buf \U$25031 ( \25035 , \25034 );
buf \U$25032 ( \25036 , \25035 );
xor \U$25033 ( \25037 , \25030 , \25036 );
buf \U$25034 ( \25038 , \25037 );
buf \U$25035 ( \25039 , \25038 );
not \U$25036 ( \25040 , \25039 );
buf \U$25037 ( \25041 , \25040 );
buf \U$25038 ( \25042 , \25041 );
and \U$25039 ( \25043 , \25003 , \25042 );
not \U$25040 ( \25044 , \25003 );
buf \U$25041 ( \25045 , \25038 );
and \U$25042 ( \25046 , \25044 , \25045 );
nor \U$25043 ( \25047 , \25043 , \25046 );
buf \U$25044 ( \25048 , \25047 );
buf \U$25045 ( \25049 , \25048 );
not \U$25046 ( \25050 , \25049 );
or \U$25047 ( \25051 , \24924 , \25050 );
buf \U$25048 ( \25052 , \25048 );
buf \U$25049 ( \25053 , \24922 );
or \U$25050 ( \25054 , \25052 , \25053 );
nand \U$25051 ( \25055 , \25051 , \25054 );
buf \U$25052 ( \25056 , \25055 );
buf \U$25053 ( \25057 , \25056 );
xor \U$25054 ( \25058 , \24238 , \24244 );
and \U$25055 ( \25059 , \25058 , \24281 );
and \U$25056 ( \25060 , \24238 , \24244 );
or \U$25057 ( \25061 , \25059 , \25060 );
buf \U$25058 ( \25062 , \25061 );
buf \U$25059 ( \25063 , \25062 );
xor \U$25060 ( \25064 , \25057 , \25063 );
buf \U$25061 ( \25065 , \23849 );
not \U$25062 ( \25066 , \25065 );
buf \U$25063 ( \25067 , \14825 );
not \U$25064 ( \25068 , \25067 );
or \U$25065 ( \25069 , \25066 , \25068 );
buf \U$25066 ( \25070 , \1588 );
buf \U$25067 ( \25071 , RIc0d8b18_45);
buf \U$25068 ( \25072 , RIc0d9a18_77);
xor \U$25069 ( \25073 , \25071 , \25072 );
buf \U$25070 ( \25074 , \25073 );
buf \U$25071 ( \25075 , \25074 );
nand \U$25072 ( \25076 , \25070 , \25075 );
buf \U$25073 ( \25077 , \25076 );
buf \U$25074 ( \25078 , \25077 );
nand \U$25075 ( \25079 , \25069 , \25078 );
buf \U$25076 ( \25080 , \25079 );
buf \U$25077 ( \25081 , \25080 );
not \U$25078 ( \25082 , \25081 );
buf \U$25079 ( \25083 , \25082 );
buf \U$25080 ( \25084 , \24117 );
not \U$25081 ( \25085 , \25084 );
buf \U$25082 ( \25086 , \13075 );
not \U$25083 ( \25087 , \25086 );
or \U$25084 ( \25088 , \25085 , \25087 );
buf \U$25085 ( \25089 , \1078 );
buf \U$25086 ( \25090 , RIc0d8938_41);
buf \U$25087 ( \25091 , RIc0d9bf8_81);
xor \U$25088 ( \25092 , \25090 , \25091 );
buf \U$25089 ( \25093 , \25092 );
buf \U$25090 ( \25094 , \25093 );
nand \U$25091 ( \25095 , \25089 , \25094 );
buf \U$25092 ( \25096 , \25095 );
buf \U$25093 ( \25097 , \25096 );
nand \U$25094 ( \25098 , \25088 , \25097 );
buf \U$25095 ( \25099 , \25098 );
xor \U$25096 ( \25100 , \25083 , \25099 );
buf \U$25097 ( \25101 , \24640 );
not \U$25098 ( \25102 , \25101 );
buf \U$25099 ( \25103 , \22350 );
not \U$25100 ( \25104 , \25103 );
or \U$25101 ( \25105 , \25102 , \25104 );
buf \U$25102 ( \25106 , RIc0dacd8_117);
buf \U$25103 ( \25107 , RIc0d7858_5);
xnor \U$25104 ( \25108 , \25106 , \25107 );
buf \U$25105 ( \25109 , \25108 );
buf \U$25106 ( \25110 , \25109 );
not \U$25107 ( \25111 , \25110 );
buf \U$25108 ( \25112 , \12937 );
nand \U$25109 ( \25113 , \25111 , \25112 );
buf \U$25110 ( \25114 , \25113 );
buf \U$25111 ( \25115 , \25114 );
nand \U$25112 ( \25116 , \25105 , \25115 );
buf \U$25113 ( \25117 , \25116 );
xnor \U$25114 ( \25118 , \25100 , \25117 );
buf \U$25115 ( \25119 , \25118 );
buf \U$25116 ( \25120 , \24099 );
not \U$25117 ( \25121 , \25120 );
buf \U$25118 ( \25122 , \279 );
not \U$25119 ( \25123 , \25122 );
or \U$25120 ( \25124 , \25121 , \25123 );
buf \U$25121 ( \25125 , \284 );
buf \U$25122 ( \25126 , RIc0d8ed8_53);
buf \U$25123 ( \25127 , RIc0d9658_69);
xor \U$25124 ( \25128 , \25126 , \25127 );
buf \U$25125 ( \25129 , \25128 );
buf \U$25126 ( \25130 , \25129 );
nand \U$25127 ( \25131 , \25125 , \25130 );
buf \U$25128 ( \25132 , \25131 );
buf \U$25129 ( \25133 , \25132 );
nand \U$25130 ( \25134 , \25124 , \25133 );
buf \U$25131 ( \25135 , \25134 );
buf \U$25132 ( \25136 , \25135 );
buf \U$25133 ( \25137 , \14275 );
not \U$25134 ( \25138 , \25137 );
buf \U$25135 ( \25139 , \16688 );
not \U$25136 ( \25140 , \25139 );
or \U$25137 ( \25141 , \25138 , \25140 );
buf \U$25138 ( \25142 , RIc0dafa8_123);
nand \U$25139 ( \25143 , \25141 , \25142 );
buf \U$25140 ( \25144 , \25143 );
buf \U$25141 ( \25145 , \25144 );
xor \U$25142 ( \25146 , \25136 , \25145 );
buf \U$25143 ( \25147 , \12331 );
buf \U$25144 ( \25148 , \24768 );
not \U$25145 ( \25149 , \25148 );
buf \U$25146 ( \25150 , \25149 );
buf \U$25147 ( \25151 , \25150 );
or \U$25148 ( \25152 , \25147 , \25151 );
buf \U$25149 ( \25153 , \13270 );
buf \U$25150 ( \25154 , RIc0da828_107);
buf \U$25151 ( \25155 , RIc0d7d08_15);
xor \U$25152 ( \25156 , \25154 , \25155 );
buf \U$25153 ( \25157 , \25156 );
buf \U$25154 ( \25158 , \25157 );
not \U$25155 ( \25159 , \25158 );
buf \U$25156 ( \25160 , \25159 );
buf \U$25157 ( \25161 , \25160 );
or \U$25158 ( \25162 , \25153 , \25161 );
nand \U$25159 ( \25163 , \25152 , \25162 );
buf \U$25160 ( \25164 , \25163 );
buf \U$25161 ( \25165 , \25164 );
xor \U$25162 ( \25166 , \25146 , \25165 );
buf \U$25163 ( \25167 , \25166 );
buf \U$25164 ( \25168 , \25167 );
xor \U$25165 ( \25169 , \25119 , \25168 );
buf \U$25166 ( \25170 , \23956 );
not \U$25167 ( \25171 , \25170 );
buf \U$25168 ( \25172 , \2269 );
not \U$25169 ( \25173 , \25172 );
or \U$25170 ( \25174 , \25171 , \25173 );
buf \U$25171 ( \25175 , \18277 );
xor \U$25172 ( \25176 , RIc0d9748_71, RIc0d8de8_51);
buf \U$25173 ( \25177 , \25176 );
nand \U$25174 ( \25178 , \25175 , \25177 );
buf \U$25175 ( \25179 , \25178 );
buf \U$25176 ( \25180 , \25179 );
nand \U$25177 ( \25181 , \25174 , \25180 );
buf \U$25178 ( \25182 , \25181 );
buf \U$25179 ( \25183 , \25182 );
buf \U$25180 ( \25184 , \23907 );
not \U$25181 ( \25185 , \25184 );
buf \U$25182 ( \25186 , \2066 );
not \U$25183 ( \25187 , \25186 );
or \U$25184 ( \25188 , \25185 , \25187 );
buf \U$25185 ( \25189 , \2070 );
buf \U$25186 ( \25190 , RIc0da378_97);
buf \U$25187 ( \25191 , RIc0d81b8_25);
xor \U$25188 ( \25192 , \25190 , \25191 );
buf \U$25189 ( \25193 , \25192 );
buf \U$25190 ( \25194 , \25193 );
nand \U$25191 ( \25195 , \25189 , \25194 );
buf \U$25192 ( \25196 , \25195 );
buf \U$25193 ( \25197 , \25196 );
nand \U$25194 ( \25198 , \25188 , \25197 );
buf \U$25195 ( \25199 , \25198 );
buf \U$25196 ( \25200 , \25199 );
xor \U$25197 ( \25201 , \25183 , \25200 );
buf \U$25198 ( \25202 , \989 );
buf \U$25199 ( \25203 , \23832 );
not \U$25200 ( \25204 , \25203 );
buf \U$25201 ( \25205 , \25204 );
buf \U$25202 ( \25206 , \25205 );
or \U$25203 ( \25207 , \25202 , \25206 );
buf \U$25204 ( \25208 , \996 );
buf \U$25205 ( \25209 , RIc0d8848_39);
buf \U$25206 ( \25210 , RIc0d9ce8_83);
xor \U$25207 ( \25211 , \25209 , \25210 );
buf \U$25208 ( \25212 , \25211 );
buf \U$25209 ( \25213 , \25212 );
not \U$25210 ( \25214 , \25213 );
buf \U$25211 ( \25215 , \25214 );
buf \U$25212 ( \25216 , \25215 );
or \U$25213 ( \25217 , \25208 , \25216 );
nand \U$25214 ( \25218 , \25207 , \25217 );
buf \U$25215 ( \25219 , \25218 );
buf \U$25216 ( \25220 , \25219 );
xor \U$25217 ( \25221 , \25201 , \25220 );
buf \U$25218 ( \25222 , \25221 );
buf \U$25219 ( \25223 , \25222 );
xor \U$25220 ( \25224 , \25169 , \25223 );
buf \U$25221 ( \25225 , \25224 );
buf \U$25222 ( \25226 , \25225 );
not \U$25223 ( \25227 , \25226 );
buf \U$25224 ( \25228 , \24079 );
not \U$25225 ( \25229 , \25228 );
buf \U$25226 ( \25230 , \12299 );
not \U$25227 ( \25231 , \25230 );
or \U$25228 ( \25232 , \25229 , \25231 );
buf \U$25229 ( \25233 , \12303 );
buf \U$25230 ( \25234 , RIc0d7948_7);
buf \U$25231 ( \25235 , RIc0dabe8_115);
xor \U$25232 ( \25236 , \25234 , \25235 );
buf \U$25233 ( \25237 , \25236 );
buf \U$25234 ( \25238 , \25237 );
nand \U$25235 ( \25239 , \25233 , \25238 );
buf \U$25236 ( \25240 , \25239 );
buf \U$25237 ( \25241 , \25240 );
nand \U$25238 ( \25242 , \25232 , \25241 );
buf \U$25239 ( \25243 , \25242 );
buf \U$25240 ( \25244 , \25243 );
buf \U$25241 ( \25245 , \24058 );
not \U$25242 ( \25246 , \25245 );
buf \U$25243 ( \25247 , \2607 );
not \U$25244 ( \25248 , \25247 );
or \U$25245 ( \25249 , \25246 , \25248 );
buf \U$25246 ( \25250 , RIc0d8668_35);
buf \U$25247 ( \25251 , RIc0d9ec8_87);
xnor \U$25248 ( \25252 , \25250 , \25251 );
buf \U$25249 ( \25253 , \25252 );
buf \U$25250 ( \25254 , \25253 );
not \U$25251 ( \25255 , \25254 );
buf \U$25252 ( \25256 , \816 );
nand \U$25253 ( \25257 , \25255 , \25256 );
buf \U$25254 ( \25258 , \25257 );
buf \U$25255 ( \25259 , \25258 );
nand \U$25256 ( \25260 , \25249 , \25259 );
buf \U$25257 ( \25261 , \25260 );
buf \U$25258 ( \25262 , \25261 );
xor \U$25259 ( \25263 , \25244 , \25262 );
buf \U$25260 ( \25264 , \24624 );
not \U$25261 ( \25265 , \25264 );
buf \U$25262 ( \25266 , \3534 );
not \U$25263 ( \25267 , \25266 );
or \U$25264 ( \25268 , \25265 , \25267 );
buf \U$25265 ( \25269 , \16676 );
buf \U$25266 ( \25270 , RIc0da558_101);
buf \U$25267 ( \25271 , RIc0d7fd8_21);
xor \U$25268 ( \25272 , \25270 , \25271 );
buf \U$25269 ( \25273 , \25272 );
buf \U$25270 ( \25274 , \25273 );
nand \U$25271 ( \25275 , \25269 , \25274 );
buf \U$25272 ( \25276 , \25275 );
buf \U$25273 ( \25277 , \25276 );
nand \U$25274 ( \25278 , \25268 , \25277 );
buf \U$25275 ( \25279 , \25278 );
buf \U$25276 ( \25280 , \25279 );
xor \U$25277 ( \25281 , \25263 , \25280 );
buf \U$25278 ( \25282 , \25281 );
buf \U$25279 ( \25283 , \25282 );
buf \U$25280 ( \25284 , \24041 );
not \U$25281 ( \25285 , \25284 );
buf \U$25282 ( \25286 , \1021 );
not \U$25283 ( \25287 , \25286 );
or \U$25284 ( \25288 , \25285 , \25287 );
buf \U$25285 ( \25289 , \402 );
xor \U$25286 ( \25290 , RIc0d9b08_79, RIc0d8a28_43);
buf \U$25287 ( \25291 , \25290 );
nand \U$25288 ( \25292 , \25289 , \25291 );
buf \U$25289 ( \25293 , \25292 );
buf \U$25290 ( \25294 , \25293 );
nand \U$25291 ( \25295 , \25288 , \25294 );
buf \U$25292 ( \25296 , \25295 );
buf \U$25293 ( \25297 , \25296 );
buf \U$25294 ( \25298 , \24178 );
not \U$25295 ( \25299 , \25298 );
buf \U$25296 ( \25300 , \951 );
not \U$25297 ( \25301 , \25300 );
or \U$25298 ( \25302 , \25299 , \25301 );
buf \U$25299 ( \25303 , \1401 );
buf \U$25300 ( \25304 , RIc0d8758_37);
buf \U$25301 ( \25305 , RIc0d9dd8_85);
xor \U$25302 ( \25306 , \25304 , \25305 );
buf \U$25303 ( \25307 , \25306 );
buf \U$25304 ( \25308 , \25307 );
nand \U$25305 ( \25309 , \25303 , \25308 );
buf \U$25306 ( \25310 , \25309 );
buf \U$25307 ( \25311 , \25310 );
nand \U$25308 ( \25312 , \25302 , \25311 );
buf \U$25309 ( \25313 , \25312 );
buf \U$25310 ( \25314 , \25313 );
xor \U$25311 ( \25315 , \25297 , \25314 );
buf \U$25312 ( \25316 , \23867 );
not \U$25313 ( \25317 , \25316 );
buf \U$25314 ( \25318 , \14210 );
not \U$25315 ( \25319 , \25318 );
or \U$25316 ( \25320 , \25317 , \25319 );
buf \U$25317 ( \25321 , \20211 );
buf \U$25318 ( \25322 , RIc0da918_109);
buf \U$25319 ( \25323 , RIc0d7c18_13);
xor \U$25320 ( \25324 , \25322 , \25323 );
buf \U$25321 ( \25325 , \25324 );
buf \U$25322 ( \25326 , \25325 );
nand \U$25323 ( \25327 , \25321 , \25326 );
buf \U$25324 ( \25328 , \25327 );
buf \U$25325 ( \25329 , \25328 );
nand \U$25326 ( \25330 , \25320 , \25329 );
buf \U$25327 ( \25331 , \25330 );
buf \U$25328 ( \25332 , \25331 );
xor \U$25329 ( \25333 , \25315 , \25332 );
buf \U$25330 ( \25334 , \25333 );
buf \U$25331 ( \25335 , \25334 );
xor \U$25332 ( \25336 , \25283 , \25335 );
buf \U$25333 ( \25337 , \24725 );
not \U$25334 ( \25338 , \25337 );
buf \U$25335 ( \25339 , \776 );
not \U$25336 ( \25340 , \25339 );
or \U$25337 ( \25341 , \25338 , \25340 );
buf \U$25338 ( \25342 , \791 );
xor \U$25339 ( \25343 , RIc0d9838_73, RIc0d8cf8_49);
buf \U$25340 ( \25344 , \25343 );
nand \U$25341 ( \25345 , \25342 , \25344 );
buf \U$25342 ( \25346 , \25345 );
buf \U$25343 ( \25347 , \25346 );
nand \U$25344 ( \25348 , \25341 , \25347 );
buf \U$25345 ( \25349 , \25348 );
buf \U$25346 ( \25350 , \25349 );
buf \U$25347 ( \25351 , \24214 );
not \U$25348 ( \25352 , \25351 );
buf \U$25349 ( \25353 , \14888 );
not \U$25350 ( \25354 , \25353 );
buf \U$25351 ( \25355 , \25354 );
buf \U$25352 ( \25356 , \25355 );
not \U$25353 ( \25357 , \25356 );
or \U$25354 ( \25358 , \25352 , \25357 );
buf \U$25355 ( \25359 , \14405 );
xor \U$25356 ( \25360 , RIc0daaf8_113, RIc0d7a38_9);
buf \U$25357 ( \25361 , \25360 );
nand \U$25358 ( \25362 , \25359 , \25361 );
buf \U$25359 ( \25363 , \25362 );
buf \U$25360 ( \25364 , \25363 );
nand \U$25361 ( \25365 , \25358 , \25364 );
buf \U$25362 ( \25366 , \25365 );
buf \U$25363 ( \25367 , \25366 );
xor \U$25364 ( \25368 , \25350 , \25367 );
buf \U$25365 ( \25369 , \2207 );
not \U$25366 ( \25370 , \25369 );
buf \U$25367 ( \25371 , \25370 );
buf \U$25368 ( \25372 , \25371 );
not \U$25369 ( \25373 , \25372 );
buf \U$25370 ( \25374 , \25373 );
buf \U$25371 ( \25375 , \25374 );
buf \U$25372 ( \25376 , \23971 );
or \U$25373 ( \25377 , \25375 , \25376 );
buf \U$25374 ( \25378 , \2199 );
buf \U$25375 ( \25379 , RIc0d80c8_23);
buf \U$25376 ( \25380 , RIc0da468_99);
xor \U$25377 ( \25381 , \25379 , \25380 );
buf \U$25378 ( \25382 , \25381 );
buf \U$25379 ( \25383 , \25382 );
not \U$25380 ( \25384 , \25383 );
buf \U$25381 ( \25385 , \25384 );
buf \U$25382 ( \25386 , \25385 );
or \U$25383 ( \25387 , \25378 , \25386 );
nand \U$25384 ( \25388 , \25377 , \25387 );
buf \U$25385 ( \25389 , \25388 );
buf \U$25386 ( \25390 , \25389 );
xor \U$25387 ( \25391 , \25368 , \25390 );
buf \U$25388 ( \25392 , \25391 );
buf \U$25389 ( \25393 , \25392 );
xor \U$25390 ( \25394 , \25336 , \25393 );
buf \U$25391 ( \25395 , \25394 );
buf \U$25392 ( \25396 , \25395 );
and \U$25393 ( \25397 , \23258 , \23259 );
buf \U$25394 ( \25398 , \25397 );
buf \U$25395 ( \25399 , \25398 );
buf \U$25396 ( \25400 , \24796 );
not \U$25397 ( \25401 , \25400 );
buf \U$25398 ( \25402 , \1823 );
not \U$25399 ( \25403 , \25402 );
or \U$25400 ( \25404 , \25401 , \25403 );
buf \U$25401 ( \25405 , \686 );
buf \U$25402 ( \25406 , RIc0d8fc8_55);
buf \U$25403 ( \25407 , RIc0d9568_67);
xor \U$25404 ( \25408 , \25406 , \25407 );
buf \U$25405 ( \25409 , \25408 );
buf \U$25406 ( \25410 , \25409 );
nand \U$25407 ( \25411 , \25405 , \25410 );
buf \U$25408 ( \25412 , \25411 );
buf \U$25409 ( \25413 , \25412 );
nand \U$25410 ( \25414 , \25404 , \25413 );
buf \U$25411 ( \25415 , \25414 );
buf \U$25412 ( \25416 , \25415 );
xor \U$25413 ( \25417 , \25399 , \25416 );
buf \U$25414 ( \25418 , \23891 );
not \U$25415 ( \25419 , \25418 );
buf \U$25416 ( \25420 , \2535 );
not \U$25417 ( \25421 , \25420 );
or \U$25418 ( \25422 , \25419 , \25421 );
buf \U$25419 ( \25423 , \533 );
buf \U$25420 ( \25424 , RIc0da0a8_91);
buf \U$25421 ( \25425 , RIc0d8488_31);
xor \U$25422 ( \25426 , \25424 , \25425 );
buf \U$25423 ( \25427 , \25426 );
buf \U$25424 ( \25428 , \25427 );
nand \U$25425 ( \25429 , \25423 , \25428 );
buf \U$25426 ( \25430 , \25429 );
buf \U$25427 ( \25431 , \25430 );
nand \U$25428 ( \25432 , \25422 , \25431 );
buf \U$25429 ( \25433 , \25432 );
buf \U$25430 ( \25434 , \25433 );
xor \U$25431 ( \25435 , \25417 , \25434 );
buf \U$25432 ( \25436 , \25435 );
buf \U$25433 ( \25437 , \25436 );
buf \U$25434 ( \25438 , \23924 );
not \U$25435 ( \25439 , \25438 );
buf \U$25436 ( \25440 , \3780 );
not \U$25437 ( \25441 , \25440 );
or \U$25438 ( \25442 , \25439 , \25441 );
buf \U$25439 ( \25443 , \1229 );
buf \U$25440 ( \25444 , RIc0d9478_65);
buf \U$25441 ( \25445 , RIc0d90b8_57);
xor \U$25442 ( \25446 , \25444 , \25445 );
buf \U$25443 ( \25447 , \25446 );
buf \U$25444 ( \25448 , \25447 );
nand \U$25445 ( \25449 , \25443 , \25448 );
buf \U$25446 ( \25450 , \25449 );
buf \U$25447 ( \25451 , \25450 );
nand \U$25448 ( \25452 , \25442 , \25451 );
buf \U$25449 ( \25453 , \25452 );
buf \U$25450 ( \25454 , \25453 );
buf \U$25451 ( \25455 , \24150 );
not \U$25452 ( \25456 , \25455 );
buf \U$25453 ( \25457 , \13860 );
not \U$25454 ( \25458 , \25457 );
or \U$25455 ( \25459 , \25456 , \25458 );
buf \U$25456 ( \25460 , \344 );
buf \U$25457 ( \25461 , RIc0d82a8_27);
buf \U$25458 ( \25462 , RIc0da288_95);
xor \U$25459 ( \25463 , \25461 , \25462 );
buf \U$25460 ( \25464 , \25463 );
buf \U$25461 ( \25465 , \25464 );
nand \U$25462 ( \25466 , \25460 , \25465 );
buf \U$25463 ( \25467 , \25466 );
buf \U$25464 ( \25468 , \25467 );
nand \U$25465 ( \25469 , \25459 , \25468 );
buf \U$25466 ( \25470 , \25469 );
buf \U$25467 ( \25471 , \25470 );
xor \U$25468 ( \25472 , \25454 , \25471 );
buf \U$25469 ( \25473 , \24750 );
not \U$25470 ( \25474 , \25473 );
buf \U$25471 ( \25475 , \15644 );
buf \U$25472 ( \25476 , \25475 );
not \U$25473 ( \25477 , \25476 );
or \U$25474 ( \25478 , \25474 , \25477 );
buf \U$25475 ( \25479 , \12744 );
buf \U$25476 ( \25480 , RIc0da738_105);
buf \U$25477 ( \25481 , RIc0d7df8_17);
and \U$25478 ( \25482 , \25480 , \25481 );
not \U$25479 ( \25483 , \25480 );
buf \U$25480 ( \25484 , \7834 );
and \U$25481 ( \25485 , \25483 , \25484 );
nor \U$25482 ( \25486 , \25482 , \25485 );
buf \U$25483 ( \25487 , \25486 );
buf \U$25484 ( \25488 , \25487 );
nand \U$25485 ( \25489 , \25479 , \25488 );
buf \U$25486 ( \25490 , \25489 );
buf \U$25487 ( \25491 , \25490 );
nand \U$25488 ( \25492 , \25478 , \25491 );
buf \U$25489 ( \25493 , \25492 );
buf \U$25490 ( \25494 , \25493 );
xor \U$25491 ( \25495 , \25472 , \25494 );
buf \U$25492 ( \25496 , \25495 );
buf \U$25493 ( \25497 , \25496 );
xor \U$25494 ( \25498 , \25437 , \25497 );
buf \U$25495 ( \25499 , \3387 );
not \U$25496 ( \25500 , \25499 );
buf \U$25497 ( \25501 , \24194 );
not \U$25498 ( \25502 , \25501 );
and \U$25499 ( \25503 , \25500 , \25502 );
buf \U$25500 ( \25504 , \13494 );
buf \U$25501 ( \25505 , RIc0d8578_33);
buf \U$25502 ( \25506 , RIc0d9fb8_89);
xnor \U$25503 ( \25507 , \25505 , \25506 );
buf \U$25504 ( \25508 , \25507 );
buf \U$25505 ( \25509 , \25508 );
nor \U$25506 ( \25510 , \25504 , \25509 );
buf \U$25507 ( \25511 , \25510 );
buf \U$25508 ( \25512 , \25511 );
nor \U$25509 ( \25513 , \25503 , \25512 );
buf \U$25510 ( \25514 , \25513 );
buf \U$25511 ( \25515 , \25514 );
not \U$25512 ( \25516 , \25515 );
buf \U$25513 ( \25517 , \24366 );
not \U$25514 ( \25518 , \25517 );
buf \U$25515 ( \25519 , \15397 );
not \U$25516 ( \25520 , \25519 );
or \U$25517 ( \25521 , \25518 , \25520 );
buf \U$25518 ( \25522 , \15403 );
buf \U$25519 ( \25523 , RIc0d7ee8_19);
buf \U$25520 ( \25524 , RIc0da648_103);
xor \U$25521 ( \25525 , \25523 , \25524 );
buf \U$25522 ( \25526 , \25525 );
buf \U$25523 ( \25527 , \25526 );
nand \U$25524 ( \25528 , \25522 , \25527 );
buf \U$25525 ( \25529 , \25528 );
buf \U$25526 ( \25530 , \25529 );
nand \U$25527 ( \25531 , \25521 , \25530 );
buf \U$25528 ( \25532 , \25531 );
buf \U$25529 ( \25533 , \25532 );
not \U$25530 ( \25534 , \25533 );
buf \U$25531 ( \25535 , \25534 );
buf \U$25532 ( \25536 , \25535 );
not \U$25533 ( \25537 , \25536 );
buf \U$25534 ( \25538 , \23993 );
not \U$25535 ( \25539 , \25538 );
buf \U$25536 ( \25540 , \13178 );
not \U$25537 ( \25541 , \25540 );
buf \U$25538 ( \25542 , \25541 );
buf \U$25539 ( \25543 , \25542 );
not \U$25540 ( \25544 , \25543 );
or \U$25541 ( \25545 , \25539 , \25544 );
buf \U$25542 ( \25546 , \13953 );
buf \U$25543 ( \25547 , RIc0dadc8_119);
buf \U$25544 ( \25548 , RIc0d7768_3);
xor \U$25545 ( \25549 , \25547 , \25548 );
buf \U$25546 ( \25550 , \25549 );
buf \U$25547 ( \25551 , \25550 );
nand \U$25548 ( \25552 , \25546 , \25551 );
buf \U$25549 ( \25553 , \25552 );
buf \U$25550 ( \25554 , \25553 );
nand \U$25551 ( \25555 , \25545 , \25554 );
buf \U$25552 ( \25556 , \25555 );
buf \U$25553 ( \25557 , \25556 );
not \U$25554 ( \25558 , \25557 );
or \U$25555 ( \25559 , \25537 , \25558 );
buf \U$25556 ( \25560 , \25556 );
buf \U$25557 ( \25561 , \25535 );
or \U$25558 ( \25562 , \25560 , \25561 );
nand \U$25559 ( \25563 , \25559 , \25562 );
buf \U$25560 ( \25564 , \25563 );
buf \U$25561 ( \25565 , \25564 );
not \U$25562 ( \25566 , \25565 );
or \U$25563 ( \25567 , \25516 , \25566 );
buf \U$25564 ( \25568 , \25564 );
buf \U$25565 ( \25569 , \25514 );
or \U$25566 ( \25570 , \25568 , \25569 );
nand \U$25567 ( \25571 , \25567 , \25570 );
buf \U$25568 ( \25572 , \25571 );
buf \U$25569 ( \25573 , \25572 );
xor \U$25570 ( \25574 , \25498 , \25573 );
buf \U$25571 ( \25575 , \25574 );
buf \U$25572 ( \25576 , \25575 );
xnor \U$25573 ( \25577 , \25396 , \25576 );
buf \U$25574 ( \25578 , \25577 );
buf \U$25575 ( \25579 , \25578 );
not \U$25576 ( \25580 , \25579 );
or \U$25577 ( \25581 , \25227 , \25580 );
buf \U$25578 ( \25582 , \25578 );
buf \U$25579 ( \25583 , \25225 );
or \U$25580 ( \25584 , \25582 , \25583 );
nand \U$25581 ( \25585 , \25581 , \25584 );
buf \U$25582 ( \25586 , \25585 );
buf \U$25583 ( \25587 , \25586 );
xor \U$25584 ( \25588 , \24251 , \24271 );
and \U$25585 ( \25589 , \25588 , \24278 );
and \U$25586 ( \25590 , \24251 , \24271 );
or \U$25587 ( \25591 , \25589 , \25590 );
buf \U$25588 ( \25592 , \25591 );
buf \U$25589 ( \25593 , \25592 );
xor \U$25590 ( \25594 , \25587 , \25593 );
xor \U$25591 ( \25595 , \24479 , \24585 );
and \U$25592 ( \25596 , \25595 , \24825 );
and \U$25593 ( \25597 , \24479 , \24585 );
or \U$25594 ( \25598 , \25596 , \25597 );
buf \U$25595 ( \25599 , \25598 );
buf \U$25596 ( \25600 , \25599 );
xor \U$25597 ( \25601 , \25594 , \25600 );
buf \U$25598 ( \25602 , \25601 );
buf \U$25599 ( \25603 , \25602 );
xor \U$25600 ( \25604 , \25064 , \25603 );
buf \U$25601 ( \25605 , \25604 );
buf \U$25602 ( \25606 , \25605 );
not \U$25603 ( \25607 , \25606 );
buf \U$25604 ( \25608 , \25607 );
buf \U$25605 ( \25609 , \25608 );
not \U$25606 ( \25610 , \25609 );
xor \U$25607 ( \25611 , \24308 , \24328 );
and \U$25608 ( \25612 , \25611 , \24828 );
and \U$25609 ( \25613 , \24308 , \24328 );
or \U$25610 ( \25614 , \25612 , \25613 );
buf \U$25611 ( \25615 , \25614 );
buf \U$25612 ( \25616 , \25615 );
not \U$25613 ( \25617 , \25616 );
buf \U$25614 ( \25618 , \23785 );
buf \U$25615 ( \25619 , \23802 );
or \U$25616 ( \25620 , \25618 , \25619 );
buf \U$25617 ( \25621 , \23762 );
nand \U$25618 ( \25622 , \25620 , \25621 );
buf \U$25619 ( \25623 , \25622 );
buf \U$25620 ( \25624 , \25623 );
buf \U$25621 ( \25625 , \23802 );
buf \U$25622 ( \25626 , \23785 );
nand \U$25623 ( \25627 , \25625 , \25626 );
buf \U$25624 ( \25628 , \25627 );
buf \U$25625 ( \25629 , \25628 );
nand \U$25626 ( \25630 , \25624 , \25629 );
buf \U$25627 ( \25631 , \25630 );
not \U$25628 ( \25632 , \16500 );
xor \U$25629 ( \25633 , RIc0d9928_75, RIc0d8c08_47);
not \U$25630 ( \25634 , \25633 );
or \U$25631 ( \25635 , \25632 , \25634 );
buf \U$25632 ( \25636 , \24655 );
not \U$25633 ( \25637 , \25636 );
buf \U$25634 ( \25638 , \25637 );
or \U$25635 ( \25639 , \18121 , \25638 );
nand \U$25636 ( \25640 , \25635 , \25639 );
buf \U$25637 ( \25641 , \25640 );
buf \U$25638 ( \25642 , \24381 );
not \U$25639 ( \25643 , \25642 );
buf \U$25640 ( \25644 , \12529 );
not \U$25641 ( \25645 , \25644 );
or \U$25642 ( \25646 , \25643 , \25645 );
buf \U$25643 ( \25647 , \12541 );
not \U$25644 ( \25648 , \25647 );
buf \U$25645 ( \25649 , \25648 );
buf \U$25646 ( \25650 , \25649 );
xor \U$25647 ( \25651 , RIc0daa08_111, RIc0d7b28_11);
buf \U$25648 ( \25652 , \25651 );
nand \U$25649 ( \25653 , \25650 , \25652 );
buf \U$25650 ( \25654 , \25653 );
buf \U$25651 ( \25655 , \25654 );
nand \U$25652 ( \25656 , \25646 , \25655 );
buf \U$25653 ( \25657 , \25656 );
buf \U$25654 ( \25658 , \25657 );
xor \U$25655 ( \25659 , \25641 , \25658 );
buf \U$25656 ( \25660 , \24698 );
not \U$25657 ( \25661 , \25660 );
buf \U$25658 ( \25662 , \1901 );
not \U$25659 ( \25663 , \25662 );
or \U$25660 ( \25664 , \25661 , \25663 );
buf \U$25661 ( \25665 , \481 );
buf \U$25662 ( \25666 , RIc0d8398_29);
buf \U$25663 ( \25667 , RIc0da198_93);
xor \U$25664 ( \25668 , \25666 , \25667 );
buf \U$25665 ( \25669 , \25668 );
buf \U$25666 ( \25670 , \25669 );
nand \U$25667 ( \25671 , \25665 , \25670 );
buf \U$25668 ( \25672 , \25671 );
buf \U$25669 ( \25673 , \25672 );
nand \U$25670 ( \25674 , \25664 , \25673 );
buf \U$25671 ( \25675 , \25674 );
buf \U$25672 ( \25676 , \25675 );
xor \U$25673 ( \25677 , \25659 , \25676 );
buf \U$25674 ( \25678 , \25677 );
buf \U$25675 ( \25679 , \25678 );
buf \U$25676 ( \25680 , \24494 );
buf \U$25677 ( \25681 , \24680 );
not \U$25678 ( \25682 , \25681 );
buf \U$25679 ( \25683 , \17089 );
not \U$25680 ( \25684 , \25683 );
or \U$25681 ( \25685 , \25682 , \25684 );
buf \U$25682 ( \25686 , RIc0daeb8_121);
buf \U$25683 ( \25687 , RIc0d7678_1);
xnor \U$25684 ( \25688 , \25686 , \25687 );
buf \U$25685 ( \25689 , \25688 );
buf \U$25686 ( \25690 , \25689 );
not \U$25687 ( \25691 , \25690 );
buf \U$25688 ( \25692 , \13314 );
nand \U$25689 ( \25693 , \25691 , \25692 );
buf \U$25690 ( \25694 , \25693 );
buf \U$25691 ( \25695 , \25694 );
nand \U$25692 ( \25696 , \25685 , \25695 );
buf \U$25693 ( \25697 , \25696 );
buf \U$25694 ( \25698 , \25697 );
not \U$25695 ( \25699 , \25698 );
buf \U$25696 ( \25700 , \25699 );
buf \U$25697 ( \25701 , \25700 );
and \U$25698 ( \25702 , \25680 , \25701 );
not \U$25699 ( \25703 , \25680 );
buf \U$25700 ( \25704 , \25697 );
and \U$25701 ( \25705 , \25703 , \25704 );
nor \U$25702 ( \25706 , \25702 , \25705 );
buf \U$25703 ( \25707 , \25706 );
buf \U$25704 ( \25708 , \25707 );
not \U$25705 ( \25709 , \25708 );
buf \U$25706 ( \25710 , \25709 );
buf \U$25707 ( \25711 , \25710 );
not \U$25708 ( \25712 , \25711 );
buf \U$25709 ( \25713 , \24731 );
buf \U$25710 ( \25714 , \24686 );
nor \U$25711 ( \25715 , \25713 , \25714 );
buf \U$25712 ( \25716 , \25715 );
buf \U$25713 ( \25717 , \25716 );
buf \U$25714 ( \25718 , \24711 );
or \U$25715 ( \25719 , \25717 , \25718 );
buf \U$25716 ( \25720 , \24731 );
buf \U$25717 ( \25721 , \24686 );
nand \U$25718 ( \25722 , \25720 , \25721 );
buf \U$25719 ( \25723 , \25722 );
buf \U$25720 ( \25724 , \25723 );
nand \U$25721 ( \25725 , \25719 , \25724 );
buf \U$25722 ( \25726 , \25725 );
buf \U$25723 ( \25727 , \25726 );
not \U$25724 ( \25728 , \25727 );
or \U$25725 ( \25729 , \25712 , \25728 );
buf \U$25726 ( \25730 , \25726 );
not \U$25727 ( \25731 , \25730 );
buf \U$25728 ( \25732 , \25707 );
nand \U$25729 ( \25733 , \25731 , \25732 );
buf \U$25730 ( \25734 , \25733 );
buf \U$25731 ( \25735 , \25734 );
nand \U$25732 ( \25736 , \25729 , \25735 );
buf \U$25733 ( \25737 , \25736 );
buf \U$25734 ( \25738 , \25737 );
xor \U$25735 ( \25739 , \25679 , \25738 );
not \U$25736 ( \25740 , \24435 );
not \U$25737 ( \25741 , \24464 );
or \U$25738 ( \25742 , \25740 , \25741 );
buf \U$25739 ( \25743 , \24464 );
not \U$25740 ( \25744 , \25743 );
buf \U$25741 ( \25745 , \25744 );
not \U$25742 ( \25746 , \25745 );
not \U$25743 ( \25747 , \24438 );
or \U$25744 ( \25748 , \25746 , \25747 );
nand \U$25745 ( \25749 , \25748 , \24414 );
nand \U$25746 ( \25750 , \25742 , \25749 );
buf \U$25747 ( \25751 , \25750 );
xor \U$25748 ( \25752 , \25739 , \25751 );
buf \U$25749 ( \25753 , \25752 );
buf \U$25750 ( \25754 , \25753 );
xor \U$25751 ( \25755 , \24535 , \24575 );
and \U$25752 ( \25756 , \25755 , \24582 );
and \U$25753 ( \25757 , \24535 , \24575 );
or \U$25754 ( \25758 , \25756 , \25757 );
buf \U$25755 ( \25759 , \25758 );
buf \U$25756 ( \25760 , \25759 );
xor \U$25757 ( \25761 , \25754 , \25760 );
buf \U$25758 ( \25762 , \24226 );
buf \U$25759 ( \25763 , \24030 );
or \U$25760 ( \25764 , \25762 , \25763 );
buf \U$25761 ( \25765 , \24010 );
nand \U$25762 ( \25766 , \25764 , \25765 );
buf \U$25763 ( \25767 , \25766 );
buf \U$25764 ( \25768 , \25767 );
buf \U$25765 ( \25769 , \24226 );
buf \U$25766 ( \25770 , \24030 );
nand \U$25767 ( \25771 , \25769 , \25770 );
buf \U$25768 ( \25772 , \25771 );
buf \U$25769 ( \25773 , \25772 );
nand \U$25770 ( \25774 , \25768 , \25773 );
buf \U$25771 ( \25775 , \25774 );
buf \U$25772 ( \25776 , \25775 );
xor \U$25773 ( \25777 , \25761 , \25776 );
buf \U$25774 ( \25778 , \25777 );
xor \U$25775 ( \25779 , \25631 , \25778 );
buf \U$25776 ( \25780 , \25779 );
xor \U$25777 ( \25781 , \23770 , \23776 );
and \U$25778 ( \25782 , \25781 , \23783 );
and \U$25779 ( \25783 , \23770 , \23776 );
or \U$25780 ( \25784 , \25782 , \25783 );
buf \U$25781 ( \25785 , \25784 );
buf \U$25782 ( \25786 , \25785 );
xor \U$25783 ( \25787 , \24335 , \24394 );
and \U$25784 ( \25788 , \25787 , \24476 );
and \U$25785 ( \25789 , \24335 , \24394 );
or \U$25786 ( \25790 , \25788 , \25789 );
buf \U$25787 ( \25791 , \25790 );
buf \U$25788 ( \25792 , \25791 );
xor \U$25789 ( \25793 , \25786 , \25792 );
xor \U$25790 ( \25794 , \24495 , \24516 );
and \U$25791 ( \25795 , \25794 , \24532 );
and \U$25792 ( \25796 , \24495 , \24516 );
or \U$25793 ( \25797 , \25795 , \25796 );
buf \U$25794 ( \25798 , \25797 );
buf \U$25795 ( \25799 , \25798 );
xor \U$25796 ( \25800 , \24550 , \24556 );
and \U$25797 ( \25801 , \25800 , \24572 );
and \U$25798 ( \25802 , \24550 , \24556 );
or \U$25799 ( \25803 , \25801 , \25802 );
buf \U$25800 ( \25804 , \25803 );
buf \U$25801 ( \25805 , \25804 );
xor \U$25802 ( \25806 , \25799 , \25805 );
buf \U$25803 ( \25807 , \24756 );
buf \U$25804 ( \25808 , \24802 );
nor \U$25805 ( \25809 , \25807 , \25808 );
buf \U$25806 ( \25810 , \25809 );
buf \U$25807 ( \25811 , \25810 );
buf \U$25808 ( \25812 , \24777 );
or \U$25809 ( \25813 , \25811 , \25812 );
buf \U$25810 ( \25814 , \24802 );
buf \U$25811 ( \25815 , \24756 );
nand \U$25812 ( \25816 , \25814 , \25815 );
buf \U$25813 ( \25817 , \25816 );
buf \U$25814 ( \25818 , \25817 );
nand \U$25815 ( \25819 , \25813 , \25818 );
buf \U$25816 ( \25820 , \25819 );
buf \U$25817 ( \25821 , \25820 );
buf \U$25818 ( \25822 , \24126 );
not \U$25819 ( \25823 , \25822 );
buf \U$25820 ( \25824 , \24132 );
not \U$25821 ( \25825 , \25824 );
or \U$25822 ( \25826 , \25823 , \25825 );
buf \U$25823 ( \25827 , \24156 );
nand \U$25824 ( \25828 , \25826 , \25827 );
buf \U$25825 ( \25829 , \25828 );
buf \U$25826 ( \25830 , \25829 );
buf \U$25827 ( \25831 , \24105 );
buf \U$25828 ( \25832 , \24123 );
nand \U$25829 ( \25833 , \25831 , \25832 );
buf \U$25830 ( \25834 , \25833 );
buf \U$25831 ( \25835 , \25834 );
nand \U$25832 ( \25836 , \25830 , \25835 );
buf \U$25833 ( \25837 , \25836 );
buf \U$25834 ( \25838 , \25837 );
xor \U$25835 ( \25839 , \25821 , \25838 );
xor \U$25836 ( \25840 , \24356 , \24373 );
and \U$25837 ( \25841 , \25840 , \24388 );
and \U$25838 ( \25842 , \24356 , \24373 );
or \U$25839 ( \25843 , \25841 , \25842 );
buf \U$25840 ( \25844 , \25843 );
buf \U$25841 ( \25845 , \25844 );
xor \U$25842 ( \25846 , \25839 , \25845 );
buf \U$25843 ( \25847 , \25846 );
buf \U$25844 ( \25848 , \25847 );
xor \U$25845 ( \25849 , \25806 , \25848 );
buf \U$25846 ( \25850 , \25849 );
buf \U$25847 ( \25851 , \25850 );
xor \U$25848 ( \25852 , \25793 , \25851 );
buf \U$25849 ( \25853 , \25852 );
buf \U$25850 ( \25854 , \25853 );
not \U$25851 ( \25855 , \25854 );
buf \U$25852 ( \25856 , \25855 );
buf \U$25853 ( \25857 , \25856 );
and \U$25854 ( \25858 , \25780 , \25857 );
not \U$25855 ( \25859 , \25780 );
buf \U$25856 ( \25860 , \25853 );
and \U$25857 ( \25861 , \25859 , \25860 );
nor \U$25858 ( \25862 , \25858 , \25861 );
buf \U$25859 ( \25863 , \25862 );
buf \U$25860 ( \25864 , \25863 );
not \U$25861 ( \25865 , \25864 );
or \U$25862 ( \25866 , \25617 , \25865 );
buf \U$25863 ( \25867 , \25615 );
buf \U$25864 ( \25868 , \25863 );
or \U$25865 ( \25869 , \25867 , \25868 );
nand \U$25866 ( \25870 , \25866 , \25869 );
buf \U$25867 ( \25871 , \25870 );
buf \U$25868 ( \25872 , \25871 );
not \U$25869 ( \25873 , \25872 );
buf \U$25870 ( \25874 , \23823 );
not \U$25871 ( \25875 , \25874 );
buf \U$25872 ( \25876 , \23817 );
not \U$25873 ( \25877 , \25876 );
buf \U$25874 ( \25878 , \25877 );
buf \U$25875 ( \25879 , \25878 );
nand \U$25876 ( \25880 , \25875 , \25879 );
buf \U$25877 ( \25881 , \25880 );
buf \U$25878 ( \25882 , \25881 );
buf \U$25879 ( \25883 , \24283 );
and \U$25880 ( \25884 , \25882 , \25883 );
buf \U$25881 ( \25885 , \23823 );
buf \U$25882 ( \25886 , \23817 );
and \U$25883 ( \25887 , \25885 , \25886 );
buf \U$25884 ( \25888 , \25887 );
buf \U$25885 ( \25889 , \25888 );
nor \U$25886 ( \25890 , \25884 , \25889 );
buf \U$25887 ( \25891 , \25890 );
buf \U$25888 ( \25892 , \25891 );
not \U$25889 ( \25893 , \25892 );
and \U$25890 ( \25894 , \25873 , \25893 );
buf \U$25891 ( \25895 , \25871 );
buf \U$25892 ( \25896 , \25891 );
and \U$25893 ( \25897 , \25895 , \25896 );
nor \U$25894 ( \25898 , \25894 , \25897 );
buf \U$25895 ( \25899 , \25898 );
not \U$25896 ( \25900 , \25899 );
buf \U$25897 ( \25901 , \25900 );
not \U$25898 ( \25902 , \25901 );
or \U$25899 ( \25903 , \25610 , \25902 );
buf \U$25900 ( \25904 , \25899 );
buf \U$25901 ( \25905 , \25605 );
nand \U$25902 ( \25906 , \25904 , \25905 );
buf \U$25903 ( \25907 , \25906 );
buf \U$25904 ( \25908 , \25907 );
nand \U$25905 ( \25909 , \25903 , \25908 );
buf \U$25906 ( \25910 , \25909 );
buf \U$25907 ( \25911 , \25910 );
xor \U$25908 ( \25912 , \24293 , \24831 );
and \U$25909 ( \25913 , \25912 , \24838 );
and \U$25910 ( \25914 , \24293 , \24831 );
or \U$25911 ( \25915 , \25913 , \25914 );
buf \U$25912 ( \25916 , \25915 );
buf \U$25913 ( \25917 , \25916 );
not \U$25914 ( \25918 , \25917 );
buf \U$25915 ( \25919 , \25918 );
buf \U$25916 ( \25920 , \25919 );
and \U$25917 ( \25921 , \25911 , \25920 );
not \U$25918 ( \25922 , \25911 );
buf \U$25919 ( \25923 , \25916 );
and \U$25920 ( \25924 , \25922 , \25923 );
nor \U$25921 ( \25925 , \25921 , \25924 );
buf \U$25922 ( \25926 , \25925 );
buf \U$25923 ( \25927 , \25926 );
nand \U$25924 ( \25928 , \24916 , \25927 );
buf \U$25925 ( \25929 , \25928 );
buf \U$25926 ( \25930 , \25929 );
nand \U$25927 ( \25931 , \24892 , \25930 );
buf \U$25928 ( \25932 , \25931 );
buf \U$25929 ( \25933 , \25932 );
xor \U$25930 ( \25934 , \25437 , \25497 );
and \U$25931 ( \25935 , \25934 , \25573 );
and \U$25932 ( \25936 , \25437 , \25497 );
or \U$25933 ( \25937 , \25935 , \25936 );
buf \U$25934 ( \25938 , \25937 );
xor \U$25935 ( \25939 , \25283 , \25335 );
and \U$25936 ( \25940 , \25939 , \25393 );
and \U$25937 ( \25941 , \25283 , \25335 );
or \U$25938 ( \25942 , \25940 , \25941 );
buf \U$25939 ( \25943 , \25942 );
xor \U$25940 ( \25944 , \25938 , \25943 );
xor \U$25941 ( \25945 , \25119 , \25168 );
and \U$25942 ( \25946 , \25945 , \25223 );
and \U$25943 ( \25947 , \25119 , \25168 );
or \U$25944 ( \25948 , \25946 , \25947 );
buf \U$25945 ( \25949 , \25948 );
xor \U$25946 ( \25950 , \25944 , \25949 );
buf \U$25947 ( \25951 , \25950 );
buf \U$25948 ( \25952 , \25575 );
not \U$25949 ( \25953 , \25952 );
buf \U$25950 ( \25954 , \25395 );
not \U$25951 ( \25955 , \25954 );
or \U$25952 ( \25956 , \25953 , \25955 );
buf \U$25953 ( \25957 , \25575 );
buf \U$25954 ( \25958 , \25395 );
or \U$25955 ( \25959 , \25957 , \25958 );
buf \U$25956 ( \25960 , \25225 );
nand \U$25957 ( \25961 , \25959 , \25960 );
buf \U$25958 ( \25962 , \25961 );
buf \U$25959 ( \25963 , \25962 );
nand \U$25960 ( \25964 , \25956 , \25963 );
buf \U$25961 ( \25965 , \25964 );
buf \U$25962 ( \25966 , \25965 );
not \U$25963 ( \25967 , \25966 );
buf \U$25964 ( \25968 , \25967 );
buf \U$25965 ( \25969 , \25968 );
and \U$25966 ( \25970 , \25951 , \25969 );
not \U$25967 ( \25971 , \25951 );
buf \U$25968 ( \25972 , \25965 );
and \U$25969 ( \25973 , \25971 , \25972 );
nor \U$25970 ( \25974 , \25970 , \25973 );
buf \U$25971 ( \25975 , \25974 );
buf \U$25972 ( \25976 , \25975 );
buf \U$25973 ( \25977 , \25083 );
not \U$25974 ( \25978 , \25977 );
buf \U$25975 ( \25979 , \25099 );
not \U$25976 ( \25980 , \25979 );
buf \U$25977 ( \25981 , \25980 );
buf \U$25978 ( \25982 , \25981 );
not \U$25979 ( \25983 , \25982 );
or \U$25980 ( \25984 , \25978 , \25983 );
buf \U$25981 ( \25985 , \25117 );
nand \U$25982 ( \25986 , \25984 , \25985 );
buf \U$25983 ( \25987 , \25986 );
buf \U$25984 ( \25988 , \25987 );
buf \U$25985 ( \25989 , \25099 );
buf \U$25986 ( \25990 , \25080 );
nand \U$25987 ( \25991 , \25989 , \25990 );
buf \U$25988 ( \25992 , \25991 );
buf \U$25989 ( \25993 , \25992 );
nand \U$25990 ( \25994 , \25988 , \25993 );
buf \U$25991 ( \25995 , \25994 );
buf \U$25992 ( \25996 , \25995 );
xor \U$25993 ( \25997 , \25244 , \25262 );
and \U$25994 ( \25998 , \25997 , \25280 );
and \U$25995 ( \25999 , \25244 , \25262 );
or \U$25996 ( \26000 , \25998 , \25999 );
buf \U$25997 ( \26001 , \26000 );
buf \U$25998 ( \26002 , \26001 );
xor \U$25999 ( \26003 , \25996 , \26002 );
xor \U$26000 ( \26004 , \25350 , \25367 );
and \U$26001 ( \26005 , \26004 , \25390 );
and \U$26002 ( \26006 , \25350 , \25367 );
or \U$26003 ( \26007 , \26005 , \26006 );
buf \U$26004 ( \26008 , \26007 );
buf \U$26005 ( \26009 , \26008 );
xor \U$26006 ( \26010 , \26003 , \26009 );
buf \U$26007 ( \26011 , \26010 );
buf \U$26008 ( \26012 , \26011 );
buf \U$26009 ( \26013 , \25535 );
not \U$26010 ( \26014 , \26013 );
buf \U$26011 ( \26015 , \25514 );
not \U$26012 ( \26016 , \26015 );
or \U$26013 ( \26017 , \26014 , \26016 );
buf \U$26014 ( \26018 , \25556 );
nand \U$26015 ( \26019 , \26017 , \26018 );
buf \U$26016 ( \26020 , \26019 );
buf \U$26017 ( \26021 , \26020 );
buf \U$26018 ( \26022 , \25514 );
not \U$26019 ( \26023 , \26022 );
buf \U$26020 ( \26024 , \25532 );
nand \U$26021 ( \26025 , \26023 , \26024 );
buf \U$26022 ( \26026 , \26025 );
buf \U$26023 ( \26027 , \26026 );
nand \U$26024 ( \26028 , \26021 , \26027 );
buf \U$26025 ( \26029 , \26028 );
buf \U$26026 ( \26030 , \26029 );
buf \U$26027 ( \26031 , \25182 );
buf \U$26028 ( \26032 , \25199 );
or \U$26029 ( \26033 , \26031 , \26032 );
buf \U$26030 ( \26034 , \25219 );
nand \U$26031 ( \26035 , \26033 , \26034 );
buf \U$26032 ( \26036 , \26035 );
buf \U$26033 ( \26037 , \26036 );
buf \U$26034 ( \26038 , \25199 );
buf \U$26035 ( \26039 , \25182 );
nand \U$26036 ( \26040 , \26038 , \26039 );
buf \U$26037 ( \26041 , \26040 );
buf \U$26038 ( \26042 , \26041 );
nand \U$26039 ( \26043 , \26037 , \26042 );
buf \U$26040 ( \26044 , \26043 );
buf \U$26041 ( \26045 , \26044 );
xor \U$26042 ( \26046 , \26030 , \26045 );
xor \U$26043 ( \26047 , \25454 , \25471 );
and \U$26044 ( \26048 , \26047 , \25494 );
and \U$26045 ( \26049 , \25454 , \25471 );
or \U$26046 ( \26050 , \26048 , \26049 );
buf \U$26047 ( \26051 , \26050 );
buf \U$26048 ( \26052 , \26051 );
xor \U$26049 ( \26053 , \26046 , \26052 );
buf \U$26050 ( \26054 , \26053 );
buf \U$26051 ( \26055 , \26054 );
xor \U$26052 ( \26056 , \26012 , \26055 );
xor \U$26053 ( \26057 , \25297 , \25314 );
and \U$26054 ( \26058 , \26057 , \25332 );
and \U$26055 ( \26059 , \25297 , \25314 );
or \U$26056 ( \26060 , \26058 , \26059 );
buf \U$26057 ( \26061 , \26060 );
buf \U$26058 ( \26062 , \26061 );
xor \U$26059 ( \26063 , \25641 , \25658 );
and \U$26060 ( \26064 , \26063 , \25676 );
and \U$26061 ( \26065 , \25641 , \25658 );
or \U$26062 ( \26066 , \26064 , \26065 );
buf \U$26063 ( \26067 , \26066 );
buf \U$26064 ( \26068 , \26067 );
xor \U$26065 ( \26069 , \26062 , \26068 );
xor \U$26066 ( \26070 , \25136 , \25145 );
and \U$26067 ( \26071 , \26070 , \25165 );
and \U$26068 ( \26072 , \25136 , \25145 );
or \U$26069 ( \26073 , \26071 , \26072 );
buf \U$26070 ( \26074 , \26073 );
buf \U$26071 ( \26075 , \26074 );
xor \U$26072 ( \26076 , \26069 , \26075 );
buf \U$26073 ( \26077 , \26076 );
buf \U$26074 ( \26078 , \26077 );
xor \U$26075 ( \26079 , \26056 , \26078 );
buf \U$26076 ( \26080 , \26079 );
buf \U$26077 ( \26081 , \26080 );
not \U$26078 ( \26082 , \26081 );
buf \U$26079 ( \26083 , \26082 );
buf \U$26080 ( \26084 , \26083 );
and \U$26081 ( \26085 , \25976 , \26084 );
not \U$26082 ( \26086 , \25976 );
buf \U$26083 ( \26087 , \26080 );
and \U$26084 ( \26088 , \26086 , \26087 );
nor \U$26085 ( \26089 , \26085 , \26088 );
buf \U$26086 ( \26090 , \26089 );
buf \U$26087 ( \26091 , \26090 );
buf \U$26090 ( \26092 , \25631 );
buf \U$26091 ( \26093 , \26092 );
not \U$26092 ( \26094 , \26093 );
buf \U$26095 ( \26095 , \25778 );
buf \U$26096 ( \26096 , \26095 );
not \U$26097 ( \26097 , \26096 );
or \U$26098 ( \26098 , \26094 , \26097 );
buf \U$26099 ( \26099 , \26095 );
buf \U$26100 ( \26100 , \26092 );
or \U$26101 ( \26101 , \26099 , \26100 );
buf \U$26102 ( \26102 , \25853 );
nand \U$26103 ( \26103 , \26101 , \26102 );
buf \U$26104 ( \26104 , \26103 );
buf \U$26105 ( \26105 , \26104 );
nand \U$26106 ( \26106 , \26098 , \26105 );
buf \U$26107 ( \26107 , \26106 );
buf \U$26108 ( \26108 , \26107 );
xor \U$26109 ( \26109 , \26091 , \26108 );
buf \U$26110 ( \26110 , \25343 );
not \U$26111 ( \26111 , \26110 );
buf \U$26112 ( \26112 , \12442 );
not \U$26113 ( \26113 , \26112 );
or \U$26114 ( \26114 , \26111 , \26113 );
buf \U$26115 ( \26115 , \1856 );
xor \U$26116 ( \26116 , RIc0d9838_73, RIc0d8c80_48);
buf \U$26117 ( \26117 , \26116 );
nand \U$26118 ( \26118 , \26115 , \26117 );
buf \U$26119 ( \26119 , \26118 );
buf \U$26120 ( \26120 , \26119 );
nand \U$26121 ( \26121 , \26114 , \26120 );
buf \U$26122 ( \26122 , \26121 );
buf \U$26123 ( \26123 , \26122 );
buf \U$26124 ( \26124 , \25464 );
not \U$26125 ( \26125 , \26124 );
buf \U$26126 ( \26126 , \330 );
not \U$26127 ( \26127 , \26126 );
or \U$26128 ( \26128 , \26125 , \26127 );
buf \U$26129 ( \26129 , \344 );
buf \U$26130 ( \26130 , RIc0da288_95);
buf \U$26131 ( \26131 , RIc0d8230_26);
xor \U$26132 ( \26132 , \26130 , \26131 );
buf \U$26133 ( \26133 , \26132 );
buf \U$26134 ( \26134 , \26133 );
nand \U$26135 ( \26135 , \26129 , \26134 );
buf \U$26136 ( \26136 , \26135 );
buf \U$26137 ( \26137 , \26136 );
nand \U$26138 ( \26138 , \26128 , \26137 );
buf \U$26139 ( \26139 , \26138 );
buf \U$26140 ( \26140 , \26139 );
xor \U$26141 ( \26141 , \26123 , \26140 );
buf \U$26142 ( \26142 , \25669 );
not \U$26143 ( \26143 , \26142 );
buf \U$26144 ( \26144 , \476 );
not \U$26145 ( \26145 , \26144 );
or \U$26146 ( \26146 , \26143 , \26145 );
buf \U$26147 ( \26147 , RIc0da198_93);
buf \U$26148 ( \26148 , RIc0d8320_28);
xnor \U$26149 ( \26149 , \26147 , \26148 );
buf \U$26150 ( \26150 , \26149 );
buf \U$26151 ( \26151 , \26150 );
not \U$26152 ( \26152 , \26151 );
buf \U$26153 ( \26153 , \4008 );
nand \U$26154 ( \26154 , \26152 , \26153 );
buf \U$26155 ( \26155 , \26154 );
buf \U$26156 ( \26156 , \26155 );
nand \U$26157 ( \26157 , \26146 , \26156 );
buf \U$26158 ( \26158 , \26157 );
buf \U$26159 ( \26159 , \26158 );
xor \U$26160 ( \26160 , \26141 , \26159 );
buf \U$26161 ( \26161 , \26160 );
buf \U$26162 ( \26162 , \26161 );
xor \U$26163 ( \26163 , \25399 , \25416 );
and \U$26164 ( \26164 , \26163 , \25434 );
and \U$26165 ( \26165 , \25399 , \25416 );
or \U$26166 ( \26166 , \26164 , \26165 );
buf \U$26167 ( \26167 , \26166 );
buf \U$26168 ( \26168 , \26167 );
xor \U$26169 ( \26169 , \26162 , \26168 );
buf \U$26170 ( \26170 , \26169 );
buf \U$26171 ( \26171 , \26170 );
buf \U$26172 ( \26172 , RIc0d87d0_38);
buf \U$26173 ( \26173 , RIc0d9ce8_83);
xor \U$26174 ( \26174 , \26172 , \26173 );
buf \U$26175 ( \26175 , \26174 );
buf \U$26176 ( \26176 , \26175 );
not \U$26177 ( \26177 , \26176 );
buf \U$26178 ( \26178 , \993 );
not \U$26179 ( \26179 , \26178 );
or \U$26180 ( \26180 , \26177 , \26179 );
buf \U$26181 ( \26181 , \1756 );
buf \U$26182 ( \26182 , \25212 );
buf \U$26183 ( \26183 , \566 );
nand \U$26184 ( \26184 , \26181 , \26182 , \26183 );
buf \U$26185 ( \26185 , \26184 );
buf \U$26186 ( \26186 , \26185 );
nand \U$26187 ( \26187 , \26180 , \26186 );
buf \U$26188 ( \26188 , \26187 );
buf \U$26189 ( \26189 , \26188 );
buf \U$26190 ( \26190 , \25157 );
not \U$26191 ( \26191 , \26190 );
buf \U$26192 ( \26192 , \17595 );
not \U$26193 ( \26193 , \26192 );
or \U$26194 ( \26194 , \26191 , \26193 );
buf \U$26195 ( \26195 , \12342 );
xor \U$26196 ( \26196 , RIc0da828_107, RIc0d7c90_14);
buf \U$26197 ( \26197 , \26196 );
nand \U$26198 ( \26198 , \26195 , \26197 );
buf \U$26199 ( \26199 , \26198 );
buf \U$26200 ( \26200 , \26199 );
nand \U$26201 ( \26201 , \26194 , \26200 );
buf \U$26202 ( \26202 , \26201 );
buf \U$26203 ( \26203 , \26202 );
xor \U$26204 ( \26204 , \26189 , \26203 );
buf \U$26205 ( \26205 , \25074 );
not \U$26206 ( \26206 , \26205 );
buf \U$26207 ( \26207 , \1183 );
not \U$26208 ( \26208 , \26207 );
or \U$26209 ( \26209 , \26206 , \26208 );
buf \U$26210 ( \26210 , \6141 );
xor \U$26211 ( \26211 , RIc0d9a18_77, RIc0d8aa0_44);
buf \U$26212 ( \26212 , \26211 );
nand \U$26213 ( \26213 , \26210 , \26212 );
buf \U$26214 ( \26214 , \26213 );
buf \U$26215 ( \26215 , \26214 );
nand \U$26216 ( \26216 , \26209 , \26215 );
buf \U$26217 ( \26217 , \26216 );
buf \U$26218 ( \26218 , \26217 );
xor \U$26219 ( \26219 , \26204 , \26218 );
buf \U$26220 ( \26220 , \26219 );
buf \U$26221 ( \26221 , \26220 );
and \U$26222 ( \26222 , \26171 , \26221 );
not \U$26223 ( \26223 , \26171 );
buf \U$26224 ( \26224 , \26220 );
not \U$26225 ( \26225 , \26224 );
buf \U$26226 ( \26226 , \26225 );
buf \U$26227 ( \26227 , \26226 );
and \U$26228 ( \26228 , \26223 , \26227 );
nor \U$26229 ( \26229 , \26222 , \26228 );
buf \U$26230 ( \26230 , \26229 );
buf \U$26231 ( \26231 , \26230 );
and \U$26232 ( \26232 , \23921 , \23922 );
buf \U$26233 ( \26233 , \26232 );
buf \U$26234 ( \26234 , \26233 );
buf \U$26235 ( \26235 , \284 );
buf \U$26236 ( \26236 , \272 );
buf \U$26237 ( \26237 , \25129 );
nand \U$26238 ( \26238 , \26236 , \26237 );
buf \U$26239 ( \26239 , \26238 );
buf \U$26240 ( \26240 , \26239 );
or \U$26241 ( \26241 , \26235 , \26240 );
buf \U$26242 ( \26242 , \21657 );
buf \U$26243 ( \26243 , RIc0d8e60_52);
buf \U$26244 ( \26244 , RIc0d9658_69);
xor \U$26245 ( \26245 , \26243 , \26244 );
buf \U$26246 ( \26246 , \26245 );
buf \U$26247 ( \26247 , \26246 );
nand \U$26248 ( \26248 , \26242 , \26247 );
buf \U$26249 ( \26249 , \26248 );
buf \U$26250 ( \26250 , \26249 );
nand \U$26251 ( \26251 , \26241 , \26250 );
buf \U$26252 ( \26252 , \26251 );
buf \U$26253 ( \26253 , \26252 );
xor \U$26254 ( \26254 , \26234 , \26253 );
buf \U$26255 ( \26255 , \25409 );
not \U$26256 ( \26256 , \26255 );
buf \U$26257 ( \26257 , \1414 );
not \U$26258 ( \26258 , \26257 );
or \U$26259 ( \26259 , \26256 , \26258 );
buf \U$26260 ( \26260 , \686 );
buf \U$26261 ( \26261 , RIc0d8f50_54);
buf \U$26262 ( \26262 , RIc0d9568_67);
xor \U$26263 ( \26263 , \26261 , \26262 );
buf \U$26264 ( \26264 , \26263 );
buf \U$26265 ( \26265 , \26264 );
nand \U$26266 ( \26266 , \26260 , \26265 );
buf \U$26267 ( \26267 , \26266 );
buf \U$26268 ( \26268 , \26267 );
nand \U$26269 ( \26269 , \26259 , \26268 );
buf \U$26270 ( \26270 , \26269 );
buf \U$26271 ( \26271 , \26270 );
xor \U$26272 ( \26272 , \26254 , \26271 );
buf \U$26273 ( \26273 , \26272 );
buf \U$26274 ( \26274 , \26273 );
buf \U$26275 ( \26275 , RIc0d88c0_40);
buf \U$26276 ( \26276 , RIc0d9bf8_81);
xor \U$26277 ( \26277 , \26275 , \26276 );
buf \U$26278 ( \26278 , \26277 );
buf \U$26279 ( \26279 , \26278 );
not \U$26280 ( \26280 , \26279 );
buf \U$26281 ( \26281 , \1078 );
not \U$26282 ( \26282 , \26281 );
or \U$26283 ( \26283 , \26280 , \26282 );
buf \U$26284 ( \26284 , \1056 );
buf \U$26285 ( \26285 , \25093 );
nand \U$26286 ( \26286 , \26284 , \26285 );
buf \U$26287 ( \26287 , \26286 );
buf \U$26288 ( \26288 , \26287 );
buf \U$26289 ( \26289 , \1078 );
or \U$26290 ( \26290 , \26288 , \26289 );
nand \U$26291 ( \26291 , \26283 , \26290 );
buf \U$26292 ( \26292 , \26291 );
buf \U$26293 ( \26293 , \26292 );
buf \U$26294 ( \26294 , \25487 );
not \U$26295 ( \26295 , \26294 );
buf \U$26296 ( \26296 , \12736 );
not \U$26297 ( \26297 , \26296 );
or \U$26298 ( \26298 , \26295 , \26297 );
buf \U$26299 ( \26299 , \15650 );
not \U$26300 ( \26300 , \26299 );
buf \U$26301 ( \26301 , \26300 );
buf \U$26302 ( \26302 , \26301 );
xor \U$26303 ( \26303 , RIc0da738_105, RIc0d7d80_16);
buf \U$26304 ( \26304 , \26303 );
nand \U$26305 ( \26305 , \26302 , \26304 );
buf \U$26306 ( \26306 , \26305 );
buf \U$26307 ( \26307 , \26306 );
nand \U$26308 ( \26308 , \26298 , \26307 );
buf \U$26309 ( \26309 , \26308 );
buf \U$26310 ( \26310 , \26309 );
xor \U$26311 ( \26311 , \26293 , \26310 );
buf \U$26312 ( \26312 , \25427 );
not \U$26313 ( \26313 , \26312 );
buf \U$26314 ( \26314 , \524 );
not \U$26315 ( \26315 , \26314 );
or \U$26316 ( \26316 , \26313 , \26315 );
buf \U$26317 ( \26317 , \714 );
buf \U$26318 ( \26318 , RIc0da0a8_91);
buf \U$26319 ( \26319 , RIc0d8410_30);
xor \U$26320 ( \26320 , \26318 , \26319 );
buf \U$26321 ( \26321 , \26320 );
buf \U$26322 ( \26322 , \26321 );
nand \U$26323 ( \26323 , \26317 , \26322 );
buf \U$26324 ( \26324 , \26323 );
buf \U$26325 ( \26325 , \26324 );
nand \U$26326 ( \26326 , \26316 , \26325 );
buf \U$26327 ( \26327 , \26326 );
buf \U$26328 ( \26328 , \26327 );
xor \U$26329 ( \26329 , \26311 , \26328 );
buf \U$26330 ( \26330 , \26329 );
buf \U$26331 ( \26331 , \26330 );
xor \U$26332 ( \26332 , \26274 , \26331 );
buf \U$26333 ( \26333 , \6270 );
buf \U$26334 ( \26334 , \25253 );
or \U$26335 ( \26335 , \26333 , \26334 );
buf \U$26336 ( \26336 , \634 );
buf \U$26337 ( \26337 , RIc0d85f0_34);
buf \U$26338 ( \26338 , RIc0d9ec8_87);
xor \U$26339 ( \26339 , \26337 , \26338 );
buf \U$26340 ( \26340 , \26339 );
buf \U$26341 ( \26341 , \26340 );
not \U$26342 ( \26342 , \26341 );
buf \U$26343 ( \26343 , \26342 );
buf \U$26344 ( \26344 , \26343 );
or \U$26345 ( \26345 , \26336 , \26344 );
nand \U$26346 ( \26346 , \26335 , \26345 );
buf \U$26347 ( \26347 , \26346 );
buf \U$26348 ( \26348 , \26347 );
buf \U$26349 ( \26349 , \25273 );
not \U$26350 ( \26350 , \26349 );
buf \U$26351 ( \26351 , \3535 );
not \U$26352 ( \26352 , \26351 );
or \U$26353 ( \26353 , \26350 , \26352 );
buf \U$26356 ( \26354 , \12839 );
buf \U$26357 ( \26355 , \26354 );
buf \U$26358 ( \26356 , RIc0da558_101);
buf \U$26359 ( \26357 , RIc0d7f60_20);
xor \U$26360 ( \26358 , \26356 , \26357 );
buf \U$26361 ( \26359 , \26358 );
buf \U$26362 ( \26360 , \26359 );
nand \U$26363 ( \26361 , \26355 , \26360 );
buf \U$26364 ( \26362 , \26361 );
buf \U$26365 ( \26363 , \26362 );
nand \U$26366 ( \26364 , \26353 , \26363 );
buf \U$26367 ( \26365 , \26364 );
buf \U$26368 ( \26366 , \26365 );
xor \U$26369 ( \26367 , \26348 , \26366 );
buf \U$26370 ( \26368 , \12968 );
buf \U$26371 ( \26369 , \25689 );
or \U$26372 ( \26370 , \26368 , \26369 );
buf \U$26373 ( \26371 , \16386 );
not \U$26374 ( \26372 , \26371 );
buf \U$26375 ( \26373 , \26372 );
buf \U$26376 ( \26374 , \26373 );
buf \U$26377 ( \26375 , \13166 );
or \U$26378 ( \26376 , \26374 , \26375 );
nand \U$26379 ( \26377 , \26370 , \26376 );
buf \U$26380 ( \26378 , \26377 );
buf \U$26381 ( \26379 , \26378 );
xor \U$26382 ( \26380 , \26367 , \26379 );
buf \U$26383 ( \26381 , \26380 );
buf \U$26384 ( \26382 , \26381 );
xor \U$26385 ( \26383 , \26332 , \26382 );
buf \U$26386 ( \26384 , \26383 );
buf \U$26387 ( \26385 , \26384 );
xor \U$26388 ( \26386 , \26231 , \26385 );
buf \U$26389 ( \26387 , \2812 );
buf \U$26390 ( \26388 , \25176 );
and \U$26391 ( \26389 , \26387 , \26388 );
buf \U$26392 ( \26390 , RIc0d8d70_50);
buf \U$26393 ( \26391 , RIc0d9748_71);
xor \U$26394 ( \26392 , \26390 , \26391 );
buf \U$26395 ( \26393 , \26392 );
buf \U$26396 ( \26394 , \26393 );
not \U$26397 ( \26395 , \26394 );
buf \U$26398 ( \26396 , \18274 );
nor \U$26399 ( \26397 , \26395 , \26396 );
buf \U$26400 ( \26398 , \26397 );
buf \U$26401 ( \26399 , \26398 );
nor \U$26402 ( \26400 , \26389 , \26399 );
buf \U$26403 ( \26401 , \26400 );
buf \U$26404 ( \26402 , \26401 );
not \U$26405 ( \26403 , \26402 );
buf \U$26406 ( \26404 , \26403 );
buf \U$26407 ( \26405 , \26404 );
not \U$26408 ( \26406 , \26405 );
buf \U$26409 ( \26407 , \25307 );
not \U$26410 ( \26408 , \26407 );
buf \U$26411 ( \26409 , \18767 );
not \U$26412 ( \26410 , \26409 );
buf \U$26413 ( \26411 , \26410 );
buf \U$26414 ( \26412 , \26411 );
nor \U$26415 ( \26413 , \26408 , \26412 );
buf \U$26416 ( \26414 , \26413 );
buf \U$26417 ( \26415 , \26414 );
buf \U$26418 ( \26416 , RIc0d86e0_36);
buf \U$26419 ( \26417 , RIc0d9dd8_85);
xor \U$26420 ( \26418 , \26416 , \26417 );
buf \U$26421 ( \26419 , \26418 );
buf \U$26422 ( \26420 , \26419 );
not \U$26423 ( \26421 , \26420 );
buf \U$26424 ( \26422 , \918 );
nor \U$26425 ( \26423 , \26421 , \26422 );
buf \U$26426 ( \26424 , \26423 );
buf \U$26427 ( \26425 , \26424 );
nor \U$26428 ( \26426 , \26415 , \26425 );
buf \U$26429 ( \26427 , \26426 );
buf \U$26430 ( \26428 , \26427 );
not \U$26431 ( \26429 , \26428 );
or \U$26432 ( \26430 , \26406 , \26429 );
buf \U$26433 ( \26431 , \26427 );
not \U$26434 ( \26432 , \26431 );
buf \U$26435 ( \26433 , \26432 );
buf \U$26436 ( \26434 , \26433 );
buf \U$26437 ( \26435 , \26401 );
nand \U$26438 ( \26436 , \26434 , \26435 );
buf \U$26439 ( \26437 , \26436 );
buf \U$26440 ( \26438 , \26437 );
nand \U$26441 ( \26439 , \26430 , \26438 );
buf \U$26442 ( \26440 , \26439 );
buf \U$26443 ( \26441 , \26440 );
buf \U$26444 ( \26442 , \25290 );
not \U$26445 ( \26443 , \26442 );
buf \U$26446 ( \26444 , \1351 );
not \U$26447 ( \26445 , \26444 );
or \U$26448 ( \26446 , \26443 , \26445 );
buf \U$26449 ( \26447 , \1025 );
buf \U$26450 ( \26448 , RIc0d89b0_42);
buf \U$26451 ( \26449 , RIc0d9b08_79);
xor \U$26452 ( \26450 , \26448 , \26449 );
buf \U$26453 ( \26451 , \26450 );
buf \U$26454 ( \26452 , \26451 );
nand \U$26455 ( \26453 , \26447 , \26452 );
buf \U$26456 ( \26454 , \26453 );
buf \U$26457 ( \26455 , \26454 );
nand \U$26458 ( \26456 , \26446 , \26455 );
buf \U$26459 ( \26457 , \26456 );
buf \U$26460 ( \26458 , \26457 );
xor \U$26461 ( \26459 , \26441 , \26458 );
buf \U$26462 ( \26460 , \26459 );
buf \U$26463 ( \26461 , \26460 );
buf \U$26464 ( \26462 , \25237 );
not \U$26465 ( \26463 , \26462 );
buf \U$26466 ( \26464 , \14681 );
not \U$26467 ( \26465 , \26464 );
buf \U$26468 ( \26466 , \26465 );
buf \U$26469 ( \26467 , \26466 );
not \U$26470 ( \26468 , \26467 );
or \U$26471 ( \26469 , \26463 , \26468 );
buf \U$26472 ( \26470 , \12303 );
xor \U$26473 ( \26471 , RIc0dabe8_115, RIc0d78d0_6);
buf \U$26474 ( \26472 , \26471 );
nand \U$26475 ( \26473 , \26470 , \26472 );
buf \U$26476 ( \26474 , \26473 );
buf \U$26477 ( \26475 , \26474 );
nand \U$26478 ( \26476 , \26469 , \26475 );
buf \U$26479 ( \26477 , \26476 );
buf \U$26480 ( \26478 , \26477 );
not \U$26481 ( \26479 , \26478 );
buf \U$26482 ( \26480 , \25360 );
not \U$26483 ( \26481 , \26480 );
buf \U$26484 ( \26482 , \14888 );
not \U$26485 ( \26483 , \26482 );
buf \U$26486 ( \26484 , \26483 );
buf \U$26487 ( \26485 , \26484 );
not \U$26488 ( \26486 , \26485 );
or \U$26489 ( \26487 , \26481 , \26486 );
buf \U$26490 ( \26488 , \12410 );
and \U$26491 ( \26489 , RIc0daaf8_113, \4448 );
not \U$26492 ( \26490 , RIc0daaf8_113);
and \U$26493 ( \26491 , \26490 , RIc0d79c0_8);
or \U$26494 ( \26492 , \26489 , \26491 );
buf \U$26495 ( \26493 , \26492 );
nand \U$26496 ( \26494 , \26488 , \26493 );
buf \U$26497 ( \26495 , \26494 );
buf \U$26498 ( \26496 , \26495 );
nand \U$26499 ( \26497 , \26487 , \26496 );
buf \U$26500 ( \26498 , \26497 );
buf \U$26501 ( \26499 , \26498 );
not \U$26502 ( \26500 , \26499 );
buf \U$26503 ( \26501 , \26500 );
buf \U$26504 ( \26502 , \26501 );
not \U$26505 ( \26503 , \26502 );
or \U$26506 ( \26504 , \26479 , \26503 );
buf \U$26507 ( \26505 , \26477 );
buf \U$26508 ( \26506 , \26501 );
or \U$26509 ( \26507 , \26505 , \26506 );
nand \U$26510 ( \26508 , \26504 , \26507 );
buf \U$26511 ( \26509 , \26508 );
buf \U$26512 ( \26510 , \26509 );
buf \U$26513 ( \26511 , \25508 );
not \U$26514 ( \26512 , \26511 );
buf \U$26515 ( \26513 , \26512 );
buf \U$26516 ( \26514 , \26513 );
not \U$26517 ( \26515 , \26514 );
buf \U$26518 ( \26516 , \437 );
not \U$26519 ( \26517 , \26516 );
or \U$26520 ( \26518 , \26515 , \26517 );
buf \U$26521 ( \26519 , \846 );
buf \U$26522 ( \26520 , RIc0d9fb8_89);
buf \U$26523 ( \26521 , RIc0d8500_32);
xor \U$26524 ( \26522 , \26520 , \26521 );
buf \U$26525 ( \26523 , \26522 );
buf \U$26526 ( \26524 , \26523 );
nand \U$26527 ( \26525 , \26519 , \26524 );
buf \U$26528 ( \26526 , \26525 );
buf \U$26529 ( \26527 , \26526 );
nand \U$26530 ( \26528 , \26518 , \26527 );
buf \U$26531 ( \26529 , \26528 );
buf \U$26532 ( \26530 , \26529 );
xor \U$26533 ( \26531 , \26510 , \26530 );
buf \U$26534 ( \26532 , \26531 );
buf \U$26535 ( \26533 , \26532 );
xor \U$26536 ( \26534 , \26461 , \26533 );
not \U$26537 ( \26535 , \13143 );
not \U$26538 ( \26536 , \25109 );
and \U$26539 ( \26537 , \26535 , \26536 );
buf \U$26540 ( \26538 , RIc0dacd8_117);
buf \U$26541 ( \26539 , RIc0d77e0_4);
and \U$26542 ( \26540 , \26538 , \26539 );
not \U$26543 ( \26541 , \26538 );
buf \U$26544 ( \26542 , \489 );
and \U$26545 ( \26543 , \26541 , \26542 );
nor \U$26546 ( \26544 , \26540 , \26543 );
buf \U$26547 ( \26545 , \26544 );
and \U$26548 ( \26546 , \12937 , \26545 );
nor \U$26549 ( \26547 , \26537 , \26546 );
buf \U$26550 ( \26548 , \26547 );
not \U$26551 ( \26549 , \26548 );
buf \U$26552 ( \26550 , \25651 );
not \U$26553 ( \26551 , \26550 );
buf \U$26554 ( \26552 , \18306 );
not \U$26555 ( \26553 , \26552 );
or \U$26556 ( \26554 , \26551 , \26553 );
buf \U$26557 ( \26555 , \18312 );
buf \U$26558 ( \26556 , RIc0daa08_111);
buf \U$26559 ( \26557 , RIc0d7ab0_10);
xor \U$26560 ( \26558 , \26556 , \26557 );
buf \U$26561 ( \26559 , \26558 );
buf \U$26562 ( \26560 , \26559 );
nand \U$26563 ( \26561 , \26555 , \26560 );
buf \U$26564 ( \26562 , \26561 );
buf \U$26565 ( \26563 , \26562 );
nand \U$26566 ( \26564 , \26554 , \26563 );
buf \U$26567 ( \26565 , \26564 );
buf \U$26568 ( \26566 , \26565 );
not \U$26569 ( \26567 , \26566 );
buf \U$26570 ( \26568 , \25193 );
not \U$26571 ( \26569 , \26568 );
buf \U$26572 ( \26570 , \2938 );
not \U$26573 ( \26571 , \26570 );
buf \U$26574 ( \26572 , \26571 );
buf \U$26575 ( \26573 , \26572 );
not \U$26576 ( \26574 , \26573 );
or \U$26577 ( \26575 , \26569 , \26574 );
buf \U$26578 ( \26576 , \734 );
buf \U$26579 ( \26577 , RIc0d8140_24);
buf \U$26580 ( \26578 , RIc0da378_97);
xor \U$26581 ( \26579 , \26577 , \26578 );
buf \U$26582 ( \26580 , \26579 );
buf \U$26583 ( \26581 , \26580 );
nand \U$26584 ( \26582 , \26576 , \26581 );
buf \U$26585 ( \26583 , \26582 );
buf \U$26586 ( \26584 , \26583 );
nand \U$26587 ( \26585 , \26575 , \26584 );
buf \U$26588 ( \26586 , \26585 );
buf \U$26589 ( \26587 , \26586 );
not \U$26590 ( \26588 , \26587 );
buf \U$26591 ( \26589 , \26588 );
buf \U$26592 ( \26590 , \26589 );
not \U$26593 ( \26591 , \26590 );
or \U$26594 ( \26592 , \26567 , \26591 );
buf \U$26595 ( \26593 , \26589 );
buf \U$26596 ( \26594 , \26565 );
or \U$26597 ( \26595 , \26593 , \26594 );
nand \U$26598 ( \26596 , \26592 , \26595 );
buf \U$26599 ( \26597 , \26596 );
buf \U$26600 ( \26598 , \26597 );
not \U$26601 ( \26599 , \26598 );
or \U$26602 ( \26600 , \26549 , \26599 );
buf \U$26603 ( \26601 , \26597 );
buf \U$26604 ( \26602 , \26547 );
or \U$26605 ( \26603 , \26601 , \26602 );
nand \U$26606 ( \26604 , \26600 , \26603 );
buf \U$26607 ( \26605 , \26604 );
buf \U$26608 ( \26606 , \26605 );
xor \U$26609 ( \26607 , \26534 , \26606 );
buf \U$26610 ( \26608 , \26607 );
buf \U$26611 ( \26609 , \26608 );
xor \U$26612 ( \26610 , \26386 , \26609 );
buf \U$26613 ( \26611 , \26610 );
buf \U$26614 ( \26612 , \26611 );
buf \U$26615 ( \26613 , \25447 );
not \U$26616 ( \26614 , \26613 );
buf \U$26617 ( \26615 , \12795 );
not \U$26618 ( \26616 , \26615 );
or \U$26619 ( \26617 , \26614 , \26616 );
buf \U$26620 ( \26618 , \1229 );
buf \U$26621 ( \26619 , RIc0d9478_65);
buf \U$26622 ( \26620 , RIc0d9040_56);
xor \U$26623 ( \26621 , \26619 , \26620 );
buf \U$26624 ( \26622 , \26621 );
buf \U$26625 ( \26623 , \26622 );
nand \U$26626 ( \26624 , \26618 , \26623 );
buf \U$26627 ( \26625 , \26624 );
buf \U$26628 ( \26626 , \26625 );
nand \U$26629 ( \26627 , \26617 , \26626 );
buf \U$26630 ( \26628 , \26627 );
buf \U$26631 ( \26629 , \26628 );
buf \U$26632 ( \26630 , \25633 );
not \U$26633 ( \26631 , \26630 );
buf \U$26634 ( \26632 , \2358 );
not \U$26635 ( \26633 , \26632 );
or \U$26636 ( \26634 , \26631 , \26633 );
buf \U$26637 ( \26635 , \1143 );
buf \U$26638 ( \26636 , RIc0d8b90_46);
buf \U$26639 ( \26637 , RIc0d9928_75);
xor \U$26640 ( \26638 , \26636 , \26637 );
buf \U$26641 ( \26639 , \26638 );
buf \U$26642 ( \26640 , \26639 );
nand \U$26643 ( \26641 , \26635 , \26640 );
buf \U$26644 ( \26642 , \26641 );
buf \U$26645 ( \26643 , \26642 );
nand \U$26646 ( \26644 , \26634 , \26643 );
buf \U$26647 ( \26645 , \26644 );
buf \U$26648 ( \26646 , \26645 );
xor \U$26649 ( \26647 , \26629 , \26646 );
buf \U$26650 ( \26648 , \25382 );
not \U$26651 ( \26649 , \26648 );
buf \U$26652 ( \26650 , \16744 );
not \U$26653 ( \26651 , \26650 );
or \U$26654 ( \26652 , \26649 , \26651 );
buf \U$26655 ( \26653 , \2476 );
buf \U$26656 ( \26654 , RIc0d8050_22);
buf \U$26657 ( \26655 , RIc0da468_99);
xor \U$26658 ( \26656 , \26654 , \26655 );
buf \U$26659 ( \26657 , \26656 );
buf \U$26660 ( \26658 , \26657 );
nand \U$26661 ( \26659 , \26653 , \26658 );
buf \U$26662 ( \26660 , \26659 );
buf \U$26663 ( \26661 , \26660 );
nand \U$26664 ( \26662 , \26652 , \26661 );
buf \U$26665 ( \26663 , \26662 );
buf \U$26666 ( \26664 , \26663 );
xor \U$26667 ( \26665 , \26647 , \26664 );
buf \U$26668 ( \26666 , \26665 );
buf \U$26669 ( \26667 , \26666 );
buf \U$26670 ( \26668 , \25550 );
not \U$26671 ( \26669 , \26668 );
buf \U$26672 ( \26670 , \14569 );
not \U$26673 ( \26671 , \26670 );
or \U$26674 ( \26672 , \26669 , \26671 );
buf \U$26675 ( \26673 , \13953 );
buf \U$26676 ( \26674 , RIc0dadc8_119);
buf \U$26677 ( \26675 , RIc0d76f0_2);
xor \U$26678 ( \26676 , \26674 , \26675 );
buf \U$26679 ( \26677 , \26676 );
buf \U$26680 ( \26678 , \26677 );
nand \U$26681 ( \26679 , \26673 , \26678 );
buf \U$26682 ( \26680 , \26679 );
buf \U$26683 ( \26681 , \26680 );
nand \U$26684 ( \26682 , \26672 , \26681 );
buf \U$26685 ( \26683 , \26682 );
buf \U$26686 ( \26684 , \26683 );
not \U$26687 ( \26685 , \26684 );
buf \U$26688 ( \26686 , \25325 );
not \U$26689 ( \26687 , \26686 );
buf \U$26690 ( \26688 , \13419 );
not \U$26691 ( \26689 , \26688 );
or \U$26692 ( \26690 , \26687 , \26689 );
buf \U$26693 ( \26691 , \14216 );
xor \U$26694 ( \26692 , RIc0da918_109, RIc0d7ba0_12);
buf \U$26695 ( \26693 , \26692 );
nand \U$26696 ( \26694 , \26691 , \26693 );
buf \U$26697 ( \26695 , \26694 );
buf \U$26698 ( \26696 , \26695 );
nand \U$26699 ( \26697 , \26690 , \26696 );
buf \U$26700 ( \26698 , \26697 );
buf \U$26701 ( \26699 , \26698 );
not \U$26702 ( \26700 , \26699 );
buf \U$26703 ( \26701 , \26700 );
buf \U$26704 ( \26702 , \26701 );
not \U$26705 ( \26703 , \26702 );
buf \U$26706 ( \26704 , \25526 );
not \U$26707 ( \26705 , \26704 );
buf \U$26708 ( \26706 , \17405 );
not \U$26709 ( \26707 , \26706 );
or \U$26710 ( \26708 , \26705 , \26707 );
buf \U$26711 ( \26709 , \15403 );
buf \U$26712 ( \26710 , RIc0da648_103);
buf \U$26713 ( \26711 , RIc0d7e70_18);
xor \U$26714 ( \26712 , \26710 , \26711 );
buf \U$26715 ( \26713 , \26712 );
buf \U$26716 ( \26714 , \26713 );
nand \U$26717 ( \26715 , \26709 , \26714 );
buf \U$26718 ( \26716 , \26715 );
buf \U$26719 ( \26717 , \26716 );
nand \U$26720 ( \26718 , \26708 , \26717 );
buf \U$26721 ( \26719 , \26718 );
buf \U$26722 ( \26720 , \26719 );
not \U$26723 ( \26721 , \26720 );
or \U$26724 ( \26722 , \26703 , \26721 );
buf \U$26725 ( \26723 , \26701 );
buf \U$26726 ( \26724 , \26719 );
or \U$26727 ( \26725 , \26723 , \26724 );
nand \U$26728 ( \26726 , \26722 , \26725 );
buf \U$26729 ( \26727 , \26726 );
buf \U$26730 ( \26728 , \26727 );
not \U$26731 ( \26729 , \26728 );
or \U$26732 ( \26730 , \26685 , \26729 );
buf \U$26733 ( \26731 , \26727 );
buf \U$26734 ( \26732 , \26683 );
or \U$26735 ( \26733 , \26731 , \26732 );
nand \U$26736 ( \26734 , \26730 , \26733 );
buf \U$26737 ( \26735 , \26734 );
buf \U$26738 ( \26736 , \26735 );
xor \U$26739 ( \26737 , \26667 , \26736 );
buf \U$26740 ( \26738 , \24952 );
buf \U$26741 ( \26739 , \24947 );
or \U$26742 ( \26740 , \26738 , \26739 );
buf \U$26743 ( \26741 , \24968 );
nand \U$26744 ( \26742 , \26740 , \26741 );
buf \U$26745 ( \26743 , \26742 );
buf \U$26746 ( \26744 , \26743 );
buf \U$26747 ( \26745 , \24952 );
buf \U$26748 ( \26746 , \24947 );
nand \U$26749 ( \26747 , \26745 , \26746 );
buf \U$26750 ( \26748 , \26747 );
buf \U$26751 ( \26749 , \26748 );
nand \U$26752 ( \26750 , \26744 , \26749 );
buf \U$26753 ( \26751 , \26750 );
buf \U$26754 ( \26752 , \26751 );
xor \U$26755 ( \26753 , \26737 , \26752 );
buf \U$26756 ( \26754 , \26753 );
buf \U$26757 ( \26755 , \26754 );
xor \U$26758 ( \26756 , \25679 , \25738 );
and \U$26759 ( \26757 , \26756 , \25751 );
and \U$26760 ( \26758 , \25679 , \25738 );
or \U$26761 ( \26759 , \26757 , \26758 );
buf \U$26762 ( \26760 , \26759 );
buf \U$26763 ( \26761 , \26760 );
xor \U$26764 ( \26762 , \26755 , \26761 );
buf \U$26765 ( \26763 , \24494 );
buf \U$26766 ( \26764 , \25700 );
nand \U$26767 ( \26765 , \26763 , \26764 );
buf \U$26768 ( \26766 , \26765 );
buf \U$26769 ( \26767 , \26766 );
not \U$26770 ( \26768 , \26767 );
buf \U$26771 ( \26769 , \25726 );
not \U$26772 ( \26770 , \26769 );
or \U$26773 ( \26771 , \26768 , \26770 );
buf \U$26774 ( \26772 , \24491 );
buf \U$26775 ( \26773 , \25697 );
nand \U$26776 ( \26774 , \26772 , \26773 );
buf \U$26777 ( \26775 , \26774 );
buf \U$26778 ( \26776 , \26775 );
nand \U$26779 ( \26777 , \26771 , \26776 );
buf \U$26780 ( \26778 , \26777 );
buf \U$26781 ( \26779 , \26778 );
xor \U$26782 ( \26780 , \25821 , \25838 );
and \U$26783 ( \26781 , \26780 , \25845 );
and \U$26784 ( \26782 , \25821 , \25838 );
or \U$26785 ( \26783 , \26781 , \26782 );
buf \U$26786 ( \26784 , \26783 );
buf \U$26787 ( \26785 , \26784 );
xor \U$26788 ( \26786 , \26779 , \26785 );
xor \U$26789 ( \26787 , \24987 , \24992 );
and \U$26790 ( \26788 , \26787 , \24998 );
and \U$26791 ( \26789 , \24987 , \24992 );
or \U$26792 ( \26790 , \26788 , \26789 );
buf \U$26793 ( \26791 , \26790 );
xor \U$26794 ( \26792 , \26786 , \26791 );
buf \U$26795 ( \26793 , \26792 );
buf \U$26796 ( \26794 , \26793 );
xor \U$26797 ( \26795 , \26762 , \26794 );
buf \U$26798 ( \26796 , \26795 );
buf \U$26799 ( \26797 , \26796 );
xor \U$26800 ( \26798 , \26612 , \26797 );
xor \U$26801 ( \26799 , \25786 , \25792 );
and \U$26802 ( \26800 , \26799 , \25851 );
and \U$26803 ( \26801 , \25786 , \25792 );
or \U$26804 ( \26802 , \26800 , \26801 );
buf \U$26805 ( \26803 , \26802 );
buf \U$26806 ( \26804 , \26803 );
xor \U$26807 ( \26805 , \26798 , \26804 );
buf \U$26808 ( \26806 , \26805 );
buf \U$26809 ( \26807 , \26806 );
xor \U$26810 ( \26808 , \26109 , \26807 );
buf \U$26811 ( \26809 , \26808 );
buf \U$26812 ( \26810 , \26809 );
not \U$26813 ( \26811 , \26810 );
xor \U$26814 ( \26812 , \25057 , \25063 );
and \U$26815 ( \26813 , \26812 , \25603 );
and \U$26816 ( \26814 , \25057 , \25063 );
or \U$26817 ( \26815 , \26813 , \26814 );
buf \U$26818 ( \26816 , \26815 );
buf \U$26819 ( \26817 , \26816 );
not \U$26820 ( \26818 , \26817 );
xor \U$26821 ( \26819 , \25754 , \25760 );
and \U$26822 ( \26820 , \26819 , \25776 );
and \U$26823 ( \26821 , \25754 , \25760 );
or \U$26824 ( \26822 , \26820 , \26821 );
buf \U$26825 ( \26823 , \26822 );
buf \U$26826 ( \26824 , \26823 );
buf \U$26827 ( \26825 , \24921 );
not \U$26828 ( \26826 , \26825 );
buf \U$26829 ( \26827 , \25038 );
not \U$26830 ( \26828 , \26827 );
or \U$26831 ( \26829 , \26826 , \26828 );
buf \U$26832 ( \26830 , \24921 );
buf \U$26833 ( \26831 , \25038 );
or \U$26834 ( \26832 , \26830 , \26831 );
buf \U$26835 ( \26833 , \25002 );
nand \U$26836 ( \26834 , \26832 , \26833 );
buf \U$26837 ( \26835 , \26834 );
buf \U$26838 ( \26836 , \26835 );
nand \U$26839 ( \26837 , \26829 , \26836 );
buf \U$26840 ( \26838 , \26837 );
buf \U$26841 ( \26839 , \26838 );
xor \U$26842 ( \26840 , \26824 , \26839 );
xor \U$26843 ( \26841 , \25799 , \25805 );
and \U$26844 ( \26842 , \26841 , \25848 );
and \U$26845 ( \26843 , \25799 , \25805 );
or \U$26846 ( \26844 , \26842 , \26843 );
buf \U$26847 ( \26845 , \26844 );
buf \U$26848 ( \26846 , \26845 );
xor \U$26849 ( \26847 , \25009 , \25029 );
and \U$26850 ( \26848 , \26847 , \25036 );
and \U$26851 ( \26849 , \25009 , \25029 );
or \U$26852 ( \26850 , \26848 , \26849 );
buf \U$26853 ( \26851 , \26850 );
buf \U$26854 ( \26852 , \26851 );
xor \U$26855 ( \26853 , \26846 , \26852 );
xor \U$26856 ( \26854 , \24933 , \24972 );
and \U$26857 ( \26855 , \26854 , \25000 );
and \U$26858 ( \26856 , \24933 , \24972 );
or \U$26859 ( \26857 , \26855 , \26856 );
buf \U$26860 ( \26858 , \26857 );
buf \U$26861 ( \26859 , \26858 );
xor \U$26862 ( \26860 , \26853 , \26859 );
buf \U$26863 ( \26861 , \26860 );
buf \U$26864 ( \26862 , \26861 );
xor \U$26865 ( \26863 , \26840 , \26862 );
buf \U$26866 ( \26864 , \26863 );
buf \U$26867 ( \26865 , \26864 );
not \U$26868 ( \26866 , \26865 );
xor \U$26869 ( \26867 , \25587 , \25593 );
and \U$26870 ( \26868 , \26867 , \25600 );
and \U$26871 ( \26869 , \25587 , \25593 );
or \U$26872 ( \26870 , \26868 , \26869 );
buf \U$26873 ( \26871 , \26870 );
buf \U$26874 ( \26872 , \26871 );
not \U$26875 ( \26873 , \26872 );
buf \U$26876 ( \26874 , \26873 );
buf \U$26877 ( \26875 , \26874 );
not \U$26878 ( \26876 , \26875 );
and \U$26879 ( \26877 , \26866 , \26876 );
buf \U$26880 ( \26878 , \26864 );
buf \U$26881 ( \26879 , \26874 );
and \U$26882 ( \26880 , \26878 , \26879 );
nor \U$26883 ( \26881 , \26877 , \26880 );
buf \U$26884 ( \26882 , \26881 );
buf \U$26885 ( \26883 , \26882 );
not \U$26886 ( \26884 , \26883 );
and \U$26887 ( \26885 , \26818 , \26884 );
buf \U$26888 ( \26886 , \26816 );
buf \U$26889 ( \26887 , \26882 );
and \U$26890 ( \26888 , \26886 , \26887 );
nor \U$26891 ( \26889 , \26885 , \26888 );
buf \U$26892 ( \26890 , \26889 );
buf \U$26893 ( \26891 , \26890 );
not \U$26894 ( \26892 , \26891 );
or \U$26895 ( \26893 , \26811 , \26892 );
buf \U$26896 ( \26894 , \26890 );
buf \U$26897 ( \26895 , \26809 );
or \U$26898 ( \26896 , \26894 , \26895 );
nand \U$26899 ( \26897 , \26893 , \26896 );
buf \U$26900 ( \26898 , \26897 );
buf \U$26901 ( \26899 , \26898 );
buf \U$26902 ( \26900 , \25615 );
not \U$26903 ( \26901 , \26900 );
buf \U$26904 ( \26902 , \25863 );
nand \U$26905 ( \26903 , \26901 , \26902 );
buf \U$26906 ( \26904 , \26903 );
buf \U$26907 ( \26905 , \26904 );
not \U$26908 ( \26906 , \26905 );
buf \U$26909 ( \26907 , \25891 );
not \U$26910 ( \26908 , \26907 );
buf \U$26911 ( \26909 , \26908 );
buf \U$26912 ( \26910 , \26909 );
not \U$26913 ( \26911 , \26910 );
or \U$26914 ( \26912 , \26906 , \26911 );
buf \U$26915 ( \26913 , \25863 );
not \U$26916 ( \26914 , \26913 );
buf \U$26917 ( \26915 , \25615 );
nand \U$26918 ( \26916 , \26914 , \26915 );
buf \U$26919 ( \26917 , \26916 );
buf \U$26920 ( \26918 , \26917 );
nand \U$26921 ( \26919 , \26912 , \26918 );
buf \U$26922 ( \26920 , \26919 );
buf \U$26923 ( \26921 , \26920 );
not \U$26924 ( \26922 , \26921 );
buf \U$26925 ( \26923 , \26922 );
buf \U$26926 ( \26924 , \26923 );
and \U$26927 ( \26925 , \26899 , \26924 );
not \U$26928 ( \26926 , \26899 );
buf \U$26929 ( \26927 , \26920 );
and \U$26930 ( \26928 , \26926 , \26927 );
nor \U$26931 ( \26929 , \26925 , \26928 );
buf \U$26932 ( \26930 , \26929 );
buf \U$26933 ( \26931 , \26930 );
buf \U$26934 ( \26932 , \25608 );
not \U$26935 ( \26933 , \26932 );
buf \U$26936 ( \26934 , \25919 );
not \U$26937 ( \26935 , \26934 );
or \U$26938 ( \26936 , \26933 , \26935 );
not \U$26939 ( \26937 , \25899 );
buf \U$26940 ( \26938 , \26937 );
nand \U$26941 ( \26939 , \26936 , \26938 );
buf \U$26942 ( \26940 , \26939 );
buf \U$26943 ( \26941 , \26940 );
buf \U$26944 ( \26942 , \25916 );
buf \U$26945 ( \26943 , \25605 );
nand \U$26946 ( \26944 , \26942 , \26943 );
buf \U$26947 ( \26945 , \26944 );
buf \U$26948 ( \26946 , \26945 );
nand \U$26949 ( \26947 , \26941 , \26946 );
buf \U$26950 ( \26948 , \26947 );
buf \U$26951 ( \26949 , \26948 );
not \U$26952 ( \26950 , \26949 );
buf \U$26953 ( \26951 , \26950 );
buf \U$26954 ( \26952 , \26951 );
nand \U$26955 ( \26953 , \26931 , \26952 );
buf \U$26956 ( \26954 , \26953 );
buf \U$26957 ( \26955 , \26954 );
buf \U$26958 ( \26956 , \26809 );
not \U$26959 ( \26957 , \26956 );
buf \U$26960 ( \26958 , \26957 );
buf \U$26961 ( \26959 , \26958 );
not \U$26962 ( \26960 , \26959 );
buf \U$26963 ( \26961 , \26890 );
not \U$26964 ( \26962 , \26961 );
or \U$26965 ( \26963 , \26960 , \26962 );
buf \U$26966 ( \26964 , \26920 );
nand \U$26967 ( \26965 , \26963 , \26964 );
buf \U$26968 ( \26966 , \26965 );
buf \U$26969 ( \26967 , \26966 );
buf \U$26970 ( \26968 , \26890 );
not \U$26971 ( \26969 , \26968 );
buf \U$26972 ( \26970 , \26809 );
nand \U$26973 ( \26971 , \26969 , \26970 );
buf \U$26974 ( \26972 , \26971 );
buf \U$26975 ( \26973 , \26972 );
nand \U$26976 ( \26974 , \26967 , \26973 );
buf \U$26977 ( \26975 , \26974 );
buf \U$26978 ( \26976 , \26975 );
not \U$26979 ( \26977 , \26976 );
xor \U$26980 ( \26978 , \26091 , \26108 );
and \U$26981 ( \26979 , \26978 , \26807 );
and \U$26982 ( \26980 , \26091 , \26108 );
or \U$26983 ( \26981 , \26979 , \26980 );
buf \U$26984 ( \26982 , \26981 );
buf \U$26985 ( \26983 , \26982 );
buf \U$26986 ( \26984 , \26864 );
not \U$26987 ( \26985 , \26984 );
buf \U$26988 ( \26986 , \26874 );
nand \U$26989 ( \26987 , \26985 , \26986 );
buf \U$26990 ( \26988 , \26987 );
buf \U$26991 ( \26989 , \26988 );
not \U$26992 ( \26990 , \26989 );
buf \U$26993 ( \26991 , \26816 );
not \U$26994 ( \26992 , \26991 );
or \U$26995 ( \26993 , \26990 , \26992 );
buf \U$26996 ( \26994 , \26864 );
buf \U$26997 ( \26995 , \26871 );
nand \U$26998 ( \26996 , \26994 , \26995 );
buf \U$26999 ( \26997 , \26996 );
buf \U$27000 ( \26998 , \26997 );
nand \U$27001 ( \26999 , \26993 , \26998 );
buf \U$27002 ( \27000 , \26999 );
buf \U$27003 ( \27001 , \27000 );
xor \U$27004 ( \27002 , \26983 , \27001 );
xor \U$27005 ( \27003 , \26846 , \26852 );
and \U$27006 ( \27004 , \27003 , \26859 );
and \U$27007 ( \27005 , \26846 , \26852 );
or \U$27008 ( \27006 , \27004 , \27005 );
buf \U$27009 ( \27007 , \27006 );
buf \U$27010 ( \27008 , \27007 );
buf \U$27011 ( \27009 , \25965 );
not \U$27012 ( \27010 , \27009 );
buf \U$27013 ( \27011 , \26080 );
not \U$27014 ( \27012 , \27011 );
or \U$27015 ( \27013 , \27010 , \27012 );
buf \U$27016 ( \27014 , \26080 );
buf \U$27017 ( \27015 , \25965 );
or \U$27018 ( \27016 , \27014 , \27015 );
buf \U$27019 ( \27017 , \25950 );
nand \U$27020 ( \27018 , \27016 , \27017 );
buf \U$27021 ( \27019 , \27018 );
buf \U$27022 ( \27020 , \27019 );
nand \U$27023 ( \27021 , \27013 , \27020 );
buf \U$27024 ( \27022 , \27021 );
buf \U$27025 ( \27023 , \27022 );
xor \U$27026 ( \27024 , \27008 , \27023 );
buf \U$27027 ( \27025 , \25943 );
buf \U$27028 ( \27026 , \25938 );
or \U$27029 ( \27027 , \27025 , \27026 );
buf \U$27030 ( \27028 , \25949 );
nand \U$27031 ( \27029 , \27027 , \27028 );
buf \U$27032 ( \27030 , \27029 );
buf \U$27033 ( \27031 , \27030 );
buf \U$27034 ( \27032 , \25943 );
buf \U$27035 ( \27033 , \25938 );
nand \U$27036 ( \27034 , \27032 , \27033 );
buf \U$27037 ( \27035 , \27034 );
buf \U$27038 ( \27036 , \27035 );
nand \U$27039 ( \27037 , \27031 , \27036 );
buf \U$27040 ( \27038 , \27037 );
buf \U$27041 ( \27039 , \27038 );
xor \U$27042 ( \27040 , \26012 , \26055 );
and \U$27043 ( \27041 , \27040 , \26078 );
and \U$27044 ( \27042 , \26012 , \26055 );
or \U$27045 ( \27043 , \27041 , \27042 );
buf \U$27046 ( \27044 , \27043 );
buf \U$27047 ( \27045 , \27044 );
xor \U$27048 ( \27046 , \27039 , \27045 );
xor \U$27049 ( \27047 , \25996 , \26002 );
and \U$27050 ( \27048 , \27047 , \26009 );
and \U$27051 ( \27049 , \25996 , \26002 );
or \U$27052 ( \27050 , \27048 , \27049 );
buf \U$27053 ( \27051 , \27050 );
xor \U$27054 ( \27052 , \26030 , \26045 );
and \U$27055 ( \27053 , \27052 , \26052 );
and \U$27056 ( \27054 , \26030 , \26045 );
or \U$27057 ( \27055 , \27053 , \27054 );
buf \U$27058 ( \27056 , \27055 );
xor \U$27059 ( \27057 , \27051 , \27056 );
xor \U$27060 ( \27058 , \26062 , \26068 );
and \U$27061 ( \27059 , \27058 , \26075 );
and \U$27062 ( \27060 , \26062 , \26068 );
or \U$27063 ( \27061 , \27059 , \27060 );
buf \U$27064 ( \27062 , \27061 );
xor \U$27065 ( \27063 , \27057 , \27062 );
buf \U$27066 ( \27064 , \27063 );
xor \U$27067 ( \27065 , \27046 , \27064 );
buf \U$27068 ( \27066 , \27065 );
buf \U$27069 ( \27067 , \27066 );
xor \U$27070 ( \27068 , \27024 , \27067 );
buf \U$27071 ( \27069 , \27068 );
buf \U$27072 ( \27070 , \27069 );
xor \U$27073 ( \27071 , \26824 , \26839 );
and \U$27074 ( \27072 , \27071 , \26862 );
and \U$27075 ( \27073 , \26824 , \26839 );
or \U$27076 ( \27074 , \27072 , \27073 );
buf \U$27077 ( \27075 , \27074 );
buf \U$27078 ( \27076 , \27075 );
xor \U$27079 ( \27077 , \27070 , \27076 );
buf \U$27080 ( \27078 , \26167 );
not \U$27081 ( \27079 , \27078 );
buf \U$27082 ( \27080 , \26220 );
not \U$27083 ( \27081 , \27080 );
or \U$27084 ( \27082 , \27079 , \27081 );
buf \U$27085 ( \27083 , \26220 );
buf \U$27086 ( \27084 , \26167 );
or \U$27087 ( \27085 , \27083 , \27084 );
buf \U$27088 ( \27086 , \26161 );
nand \U$27089 ( \27087 , \27085 , \27086 );
buf \U$27090 ( \27088 , \27087 );
buf \U$27091 ( \27089 , \27088 );
nand \U$27092 ( \27090 , \27082 , \27089 );
buf \U$27093 ( \27091 , \27090 );
buf \U$27094 ( \27092 , \27091 );
xor \U$27095 ( \27093 , \26274 , \26331 );
and \U$27096 ( \27094 , \27093 , \26382 );
and \U$27097 ( \27095 , \26274 , \26331 );
or \U$27098 ( \27096 , \27094 , \27095 );
buf \U$27099 ( \27097 , \27096 );
buf \U$27100 ( \27098 , \27097 );
xor \U$27101 ( \27099 , \27092 , \27098 );
xor \U$27102 ( \27100 , \26461 , \26533 );
and \U$27103 ( \27101 , \27100 , \26606 );
and \U$27104 ( \27102 , \26461 , \26533 );
or \U$27105 ( \27103 , \27101 , \27102 );
buf \U$27106 ( \27104 , \27103 );
buf \U$27107 ( \27105 , \27104 );
xor \U$27108 ( \27106 , \27099 , \27105 );
buf \U$27109 ( \27107 , \27106 );
buf \U$27110 ( \27108 , \27107 );
buf \U$27111 ( \27109 , \26683 );
xor \U$27112 ( \27110 , \26123 , \26140 );
and \U$27113 ( \27111 , \27110 , \26159 );
and \U$27114 ( \27112 , \26123 , \26140 );
or \U$27115 ( \27113 , \27111 , \27112 );
buf \U$27116 ( \27114 , \27113 );
buf \U$27117 ( \27115 , \27114 );
xor \U$27118 ( \27116 , \27109 , \27115 );
xor \U$27119 ( \27117 , \26348 , \26366 );
and \U$27120 ( \27118 , \27117 , \26379 );
and \U$27121 ( \27119 , \26348 , \26366 );
or \U$27122 ( \27120 , \27118 , \27119 );
buf \U$27123 ( \27121 , \27120 );
buf \U$27124 ( \27122 , \27121 );
xor \U$27125 ( \27123 , \27116 , \27122 );
buf \U$27126 ( \27124 , \27123 );
buf \U$27127 ( \27125 , \27124 );
xor \U$27128 ( \27126 , \26234 , \26253 );
and \U$27129 ( \27127 , \27126 , \26271 );
and \U$27130 ( \27128 , \26234 , \26253 );
or \U$27131 ( \27129 , \27127 , \27128 );
buf \U$27132 ( \27130 , \27129 );
buf \U$27133 ( \27131 , \27130 );
xor \U$27134 ( \27132 , \26293 , \26310 );
and \U$27135 ( \27133 , \27132 , \26328 );
and \U$27136 ( \27134 , \26293 , \26310 );
or \U$27137 ( \27135 , \27133 , \27134 );
buf \U$27138 ( \27136 , \27135 );
buf \U$27139 ( \27137 , \27136 );
xor \U$27140 ( \27138 , \27131 , \27137 );
xor \U$27141 ( \27139 , \26189 , \26203 );
and \U$27142 ( \27140 , \27139 , \26218 );
and \U$27143 ( \27141 , \26189 , \26203 );
or \U$27144 ( \27142 , \27140 , \27141 );
buf \U$27145 ( \27143 , \27142 );
buf \U$27146 ( \27144 , \27143 );
xor \U$27147 ( \27145 , \27138 , \27144 );
buf \U$27148 ( \27146 , \27145 );
buf \U$27149 ( \27147 , \27146 );
xor \U$27150 ( \27148 , \27125 , \27147 );
xor \U$27151 ( \27149 , \26629 , \26646 );
and \U$27152 ( \27150 , \27149 , \26664 );
and \U$27153 ( \27151 , \26629 , \26646 );
or \U$27154 ( \27152 , \27150 , \27151 );
buf \U$27155 ( \27153 , \27152 );
buf \U$27156 ( \27154 , \27153 );
buf \U$27157 ( \27155 , \26529 );
not \U$27158 ( \27156 , \27155 );
buf \U$27159 ( \27157 , \26498 );
not \U$27160 ( \27158 , \27157 );
or \U$27161 ( \27159 , \27156 , \27158 );
buf \U$27162 ( \27160 , \26529 );
not \U$27163 ( \27161 , \27160 );
buf \U$27164 ( \27162 , \27161 );
buf \U$27165 ( \27163 , \27162 );
not \U$27166 ( \27164 , \27163 );
buf \U$27167 ( \27165 , \26501 );
not \U$27168 ( \27166 , \27165 );
or \U$27169 ( \27167 , \27164 , \27166 );
buf \U$27170 ( \27168 , \26477 );
nand \U$27171 ( \27169 , \27167 , \27168 );
buf \U$27172 ( \27170 , \27169 );
buf \U$27173 ( \27171 , \27170 );
nand \U$27174 ( \27172 , \27159 , \27171 );
buf \U$27175 ( \27173 , \27172 );
buf \U$27176 ( \27174 , \27173 );
xor \U$27177 ( \27175 , \27154 , \27174 );
buf \U$27178 ( \27176 , \26547 );
not \U$27179 ( \27177 , \27176 );
buf \U$27180 ( \27178 , \26589 );
not \U$27181 ( \27179 , \27178 );
or \U$27182 ( \27180 , \27177 , \27179 );
buf \U$27183 ( \27181 , \26565 );
nand \U$27184 ( \27182 , \27180 , \27181 );
buf \U$27185 ( \27183 , \27182 );
buf \U$27186 ( \27184 , \27183 );
buf \U$27187 ( \27185 , \26547 );
not \U$27188 ( \27186 , \27185 );
buf \U$27189 ( \27187 , \26586 );
nand \U$27190 ( \27188 , \27186 , \27187 );
buf \U$27191 ( \27189 , \27188 );
buf \U$27192 ( \27190 , \27189 );
nand \U$27193 ( \27191 , \27184 , \27190 );
buf \U$27194 ( \27192 , \27191 );
buf \U$27195 ( \27193 , \27192 );
xor \U$27196 ( \27194 , \27175 , \27193 );
buf \U$27197 ( \27195 , \27194 );
buf \U$27198 ( \27196 , \27195 );
xor \U$27199 ( \27197 , \27148 , \27196 );
buf \U$27200 ( \27198 , \27197 );
buf \U$27201 ( \27199 , \27198 );
xor \U$27202 ( \27200 , \27108 , \27199 );
xor \U$27203 ( \27201 , \26231 , \26385 );
and \U$27204 ( \27202 , \27201 , \26609 );
and \U$27205 ( \27203 , \26231 , \26385 );
or \U$27206 ( \27204 , \27202 , \27203 );
buf \U$27207 ( \27205 , \27204 );
buf \U$27208 ( \27206 , \27205 );
xor \U$27209 ( \27207 , \27200 , \27206 );
buf \U$27210 ( \27208 , \27207 );
buf \U$27211 ( \27209 , \27208 );
buf \U$27212 ( \27210 , \26701 );
not \U$27213 ( \27211 , \27210 );
buf \U$27214 ( \27212 , \26683 );
not \U$27215 ( \27213 , \27212 );
or \U$27216 ( \27214 , \27211 , \27213 );
buf \U$27217 ( \27215 , \26719 );
nand \U$27218 ( \27216 , \27214 , \27215 );
buf \U$27219 ( \27217 , \27216 );
buf \U$27220 ( \27218 , \27217 );
buf \U$27221 ( \27219 , \26683 );
not \U$27222 ( \27220 , \27219 );
buf \U$27223 ( \27221 , \26698 );
nand \U$27224 ( \27222 , \27220 , \27221 );
buf \U$27225 ( \27223 , \27222 );
buf \U$27226 ( \27224 , \27223 );
nand \U$27227 ( \27225 , \27218 , \27224 );
buf \U$27228 ( \27226 , \27225 );
buf \U$27229 ( \27227 , \27226 );
buf \U$27230 ( \27228 , \26639 );
not \U$27231 ( \27229 , \27228 );
buf \U$27232 ( \27230 , \13991 );
not \U$27233 ( \27231 , \27230 );
or \U$27234 ( \27232 , \27229 , \27231 );
buf \U$27235 ( \27233 , \13998 );
buf \U$27236 ( \27234 , RIc0d8b18_45);
buf \U$27237 ( \27235 , RIc0d9928_75);
xor \U$27238 ( \27236 , \27234 , \27235 );
buf \U$27239 ( \27237 , \27236 );
buf \U$27240 ( \27238 , \27237 );
nand \U$27241 ( \27239 , \27233 , \27238 );
buf \U$27242 ( \27240 , \27239 );
buf \U$27243 ( \27241 , \27240 );
nand \U$27244 ( \27242 , \27232 , \27241 );
buf \U$27245 ( \27243 , \27242 );
buf \U$27246 ( \27244 , \27243 );
buf \U$27247 ( \27245 , \26492 );
not \U$27248 ( \27246 , \27245 );
buf \U$27249 ( \27247 , \16989 );
not \U$27250 ( \27248 , \27247 );
or \U$27251 ( \27249 , \27246 , \27248 );
buf \U$27252 ( \27250 , \16662 );
xor \U$27253 ( \27251 , RIc0daaf8_113, RIc0d7948_7);
buf \U$27254 ( \27252 , \27251 );
nand \U$27255 ( \27253 , \27250 , \27252 );
buf \U$27256 ( \27254 , \27253 );
buf \U$27257 ( \27255 , \27254 );
nand \U$27258 ( \27256 , \27249 , \27255 );
buf \U$27259 ( \27257 , \27256 );
buf \U$27260 ( \27258 , \27257 );
xor \U$27261 ( \27259 , \27244 , \27258 );
buf \U$27262 ( \27260 , \26211 );
not \U$27263 ( \27261 , \27260 );
buf \U$27264 ( \27262 , \1183 );
not \U$27265 ( \27263 , \27262 );
or \U$27266 ( \27264 , \27261 , \27263 );
buf \U$27267 ( \27265 , \1193 );
not \U$27268 ( \27266 , \27265 );
buf \U$27269 ( \27267 , \27266 );
buf \U$27270 ( \27268 , \27267 );
buf \U$27271 ( \27269 , RIc0d9a18_77);
buf \U$27272 ( \27270 , RIc0d8a28_43);
xor \U$27273 ( \27271 , \27269 , \27270 );
buf \U$27274 ( \27272 , \27271 );
buf \U$27275 ( \27273 , \27272 );
nand \U$27276 ( \27274 , \27268 , \27273 );
buf \U$27277 ( \27275 , \27274 );
buf \U$27278 ( \27276 , \27275 );
nand \U$27279 ( \27277 , \27264 , \27276 );
buf \U$27280 ( \27278 , \27277 );
buf \U$27281 ( \27279 , \27278 );
xor \U$27282 ( \27280 , \27259 , \27279 );
buf \U$27283 ( \27281 , \27280 );
buf \U$27284 ( \27282 , \27281 );
xor \U$27285 ( \27283 , \27227 , \27282 );
buf \U$27286 ( \27284 , \26559 );
not \U$27287 ( \27285 , \27284 );
buf \U$27288 ( \27286 , \12529 );
not \U$27289 ( \27287 , \27286 );
or \U$27290 ( \27288 , \27285 , \27287 );
buf \U$27291 ( \27289 , \18312 );
xor \U$27292 ( \27290 , RIc0daa08_111, RIc0d7a38_9);
buf \U$27293 ( \27291 , \27290 );
nand \U$27294 ( \27292 , \27289 , \27291 );
buf \U$27295 ( \27293 , \27292 );
buf \U$27296 ( \27294 , \27293 );
nand \U$27297 ( \27295 , \27288 , \27294 );
buf \U$27298 ( \27296 , \27295 );
buf \U$27299 ( \27297 , \27296 );
buf \U$27300 ( \27298 , \26419 );
not \U$27301 ( \27299 , \27298 );
buf \U$27302 ( \27300 , \6029 );
not \U$27303 ( \27301 , \27300 );
or \U$27304 ( \27302 , \27299 , \27301 );
buf \U$27305 ( \27303 , \921 );
xor \U$27306 ( \27304 , RIc0d9dd8_85, RIc0d8668_35);
buf \U$27307 ( \27305 , \27304 );
nand \U$27308 ( \27306 , \27303 , \27305 );
buf \U$27309 ( \27307 , \27306 );
buf \U$27310 ( \27308 , \27307 );
nand \U$27311 ( \27309 , \27302 , \27308 );
buf \U$27312 ( \27310 , \27309 );
buf \U$27313 ( \27311 , \27310 );
xor \U$27314 ( \27312 , \27297 , \27311 );
buf \U$27315 ( \27313 , \26657 );
not \U$27316 ( \27314 , \27313 );
buf \U$27317 ( \27315 , \25371 );
not \U$27318 ( \27316 , \27315 );
or \U$27319 ( \27317 , \27314 , \27316 );
buf \U$27320 ( \27318 , \16750 );
xor \U$27321 ( \27319 , RIc0da468_99, RIc0d7fd8_21);
buf \U$27322 ( \27320 , \27319 );
nand \U$27323 ( \27321 , \27318 , \27320 );
buf \U$27324 ( \27322 , \27321 );
buf \U$27325 ( \27323 , \27322 );
nand \U$27326 ( \27324 , \27317 , \27323 );
buf \U$27327 ( \27325 , \27324 );
buf \U$27328 ( \27326 , \27325 );
xor \U$27329 ( \27327 , \27312 , \27326 );
buf \U$27330 ( \27328 , \27327 );
buf \U$27331 ( \27329 , \27328 );
xor \U$27332 ( \27330 , \27283 , \27329 );
buf \U$27333 ( \27331 , \27330 );
buf \U$27334 ( \27332 , \27331 );
buf \U$27335 ( \27333 , \26404 );
not \U$27336 ( \27334 , \27333 );
buf \U$27337 ( \27335 , \26433 );
not \U$27338 ( \27336 , \27335 );
or \U$27339 ( \27337 , \27334 , \27336 );
not \U$27340 ( \27338 , \26427 );
not \U$27341 ( \27339 , \26401 );
or \U$27342 ( \27340 , \27338 , \27339 );
nand \U$27343 ( \27341 , \27340 , \26457 );
buf \U$27344 ( \27342 , \27341 );
nand \U$27345 ( \27343 , \27337 , \27342 );
buf \U$27346 ( \27344 , \27343 );
buf \U$27347 ( \27345 , \27344 );
and \U$27348 ( \27346 , \25444 , \25445 );
buf \U$27349 ( \27347 , \27346 );
buf \U$27350 ( \27348 , \27347 );
buf \U$27351 ( \27349 , \26264 );
not \U$27352 ( \27350 , \27349 );
buf \U$27353 ( \27351 , \1823 );
not \U$27354 ( \27352 , \27351 );
or \U$27355 ( \27353 , \27350 , \27352 );
buf \U$27356 ( \27354 , RIc0d8ed8_53);
buf \U$27357 ( \27355 , RIc0d9568_67);
xnor \U$27358 ( \27356 , \27354 , \27355 );
buf \U$27359 ( \27357 , \27356 );
buf \U$27360 ( \27358 , \27357 );
not \U$27361 ( \27359 , \27358 );
buf \U$27362 ( \27360 , \686 );
nand \U$27363 ( \27361 , \27359 , \27360 );
buf \U$27364 ( \27362 , \27361 );
buf \U$27365 ( \27363 , \27362 );
nand \U$27366 ( \27364 , \27353 , \27363 );
buf \U$27367 ( \27365 , \27364 );
buf \U$27368 ( \27366 , \27365 );
xor \U$27369 ( \27367 , \27348 , \27366 );
buf \U$27370 ( \27368 , \26321 );
not \U$27371 ( \27369 , \27368 );
buf \U$27372 ( \27370 , \2726 );
not \U$27373 ( \27371 , \27370 );
or \U$27374 ( \27372 , \27369 , \27371 );
buf \U$27375 ( \27373 , \714 );
buf \U$27376 ( \27374 , RIc0da0a8_91);
buf \U$27377 ( \27375 , RIc0d8398_29);
xor \U$27378 ( \27376 , \27374 , \27375 );
buf \U$27379 ( \27377 , \27376 );
buf \U$27380 ( \27378 , \27377 );
nand \U$27381 ( \27379 , \27373 , \27378 );
buf \U$27382 ( \27380 , \27379 );
buf \U$27383 ( \27381 , \27380 );
nand \U$27384 ( \27382 , \27372 , \27381 );
buf \U$27385 ( \27383 , \27382 );
buf \U$27386 ( \27384 , \27383 );
xor \U$27387 ( \27385 , \27367 , \27384 );
buf \U$27388 ( \27386 , \27385 );
buf \U$27389 ( \27387 , \27386 );
xor \U$27390 ( \27388 , \27345 , \27387 );
buf \U$27391 ( \27389 , \26622 );
not \U$27392 ( \27390 , \27389 );
buf \U$27393 ( \27391 , \12795 );
not \U$27394 ( \27392 , \27391 );
or \U$27395 ( \27393 , \27390 , \27392 );
buf \U$27396 ( \27394 , \1229 );
buf \U$27397 ( \27395 , RIc0d9478_65);
buf \U$27398 ( \27396 , RIc0d8fc8_55);
xor \U$27399 ( \27397 , \27395 , \27396 );
buf \U$27400 ( \27398 , \27397 );
buf \U$27401 ( \27399 , \27398 );
nand \U$27402 ( \27400 , \27394 , \27399 );
buf \U$27403 ( \27401 , \27400 );
buf \U$27404 ( \27402 , \27401 );
nand \U$27405 ( \27403 , \27393 , \27402 );
buf \U$27406 ( \27404 , \27403 );
buf \U$27407 ( \27405 , \27404 );
buf \U$27408 ( \27406 , \26393 );
not \U$27409 ( \27407 , \27406 );
buf \U$27410 ( \27408 , \2269 );
not \U$27411 ( \27409 , \27408 );
or \U$27412 ( \27410 , \27407 , \27409 );
buf \U$27413 ( \27411 , \2927 );
buf \U$27414 ( \27412 , RIc0d9748_71);
buf \U$27415 ( \27413 , RIc0d8cf8_49);
xor \U$27416 ( \27414 , \27412 , \27413 );
buf \U$27417 ( \27415 , \27414 );
buf \U$27418 ( \27416 , \27415 );
nand \U$27419 ( \27417 , \27411 , \27416 );
buf \U$27420 ( \27418 , \27417 );
buf \U$27421 ( \27419 , \27418 );
nand \U$27422 ( \27420 , \27410 , \27419 );
buf \U$27423 ( \27421 , \27420 );
buf \U$27424 ( \27422 , \27421 );
xor \U$27425 ( \27423 , \27405 , \27422 );
buf \U$27426 ( \27424 , \26580 );
not \U$27427 ( \27425 , \27424 );
buf \U$27428 ( \27426 , \16358 );
not \U$27429 ( \27427 , \27426 );
or \U$27430 ( \27428 , \27425 , \27427 );
buf \U$27431 ( \27429 , \734 );
buf \U$27432 ( \27430 , RIc0d80c8_23);
buf \U$27433 ( \27431 , RIc0da378_97);
xor \U$27434 ( \27432 , \27430 , \27431 );
buf \U$27435 ( \27433 , \27432 );
buf \U$27436 ( \27434 , \27433 );
nand \U$27437 ( \27435 , \27429 , \27434 );
buf \U$27438 ( \27436 , \27435 );
buf \U$27439 ( \27437 , \27436 );
nand \U$27440 ( \27438 , \27428 , \27437 );
buf \U$27441 ( \27439 , \27438 );
buf \U$27442 ( \27440 , \27439 );
xor \U$27443 ( \27441 , \27423 , \27440 );
buf \U$27444 ( \27442 , \27441 );
buf \U$27445 ( \27443 , \27442 );
xor \U$27446 ( \27444 , \27388 , \27443 );
buf \U$27447 ( \27445 , \27444 );
buf \U$27448 ( \27446 , \27445 );
xor \U$27449 ( \27447 , \27332 , \27446 );
buf \U$27450 ( \27448 , \26246 );
not \U$27451 ( \27449 , \27448 );
buf \U$27452 ( \27450 , \4691 );
not \U$27453 ( \27451 , \27450 );
or \U$27454 ( \27452 , \27449 , \27451 );
buf \U$27455 ( \27453 , \874 );
buf \U$27456 ( \27454 , RIc0d8de8_51);
buf \U$27457 ( \27455 , RIc0d9658_69);
xor \U$27458 ( \27456 , \27454 , \27455 );
buf \U$27459 ( \27457 , \27456 );
buf \U$27460 ( \27458 , \27457 );
nand \U$27461 ( \27459 , \27453 , \27458 );
buf \U$27462 ( \27460 , \27459 );
buf \U$27463 ( \27461 , \27460 );
nand \U$27464 ( \27462 , \27452 , \27461 );
buf \U$27465 ( \27463 , \27462 );
buf \U$27466 ( \27464 , \27463 );
not \U$27467 ( \27465 , \27464 );
buf \U$27468 ( \27466 , \26196 );
not \U$27469 ( \27467 , \27466 );
buf \U$27470 ( \27468 , \20741 );
not \U$27471 ( \27469 , \27468 );
or \U$27472 ( \27470 , \27467 , \27469 );
buf \U$27473 ( \27471 , \16071 );
xor \U$27474 ( \27472 , RIc0da828_107, RIc0d7c18_13);
buf \U$27475 ( \27473 , \27472 );
nand \U$27476 ( \27474 , \27471 , \27473 );
buf \U$27477 ( \27475 , \27474 );
buf \U$27478 ( \27476 , \27475 );
nand \U$27479 ( \27477 , \27470 , \27476 );
buf \U$27480 ( \27478 , \27477 );
buf \U$27481 ( \27479 , \27478 );
not \U$27482 ( \27480 , \27479 );
buf \U$27483 ( \27481 , \26175 );
not \U$27484 ( \27482 , \27481 );
buf \U$27485 ( \27483 , \12254 );
not \U$27486 ( \27484 , \27483 );
or \U$27487 ( \27485 , \27482 , \27484 );
buf \U$27488 ( \27486 , \993 );
buf \U$27489 ( \27487 , RIc0d8758_37);
buf \U$27490 ( \27488 , RIc0d9ce8_83);
xor \U$27491 ( \27489 , \27487 , \27488 );
buf \U$27492 ( \27490 , \27489 );
buf \U$27493 ( \27491 , \27490 );
nand \U$27494 ( \27492 , \27486 , \27491 );
buf \U$27495 ( \27493 , \27492 );
buf \U$27496 ( \27494 , \27493 );
nand \U$27497 ( \27495 , \27485 , \27494 );
buf \U$27498 ( \27496 , \27495 );
buf \U$27499 ( \27497 , \27496 );
not \U$27500 ( \27498 , \27497 );
buf \U$27501 ( \27499 , \27498 );
buf \U$27502 ( \27500 , \27499 );
not \U$27503 ( \27501 , \27500 );
and \U$27504 ( \27502 , \27480 , \27501 );
buf \U$27505 ( \27503 , \27478 );
buf \U$27506 ( \27504 , \27499 );
and \U$27507 ( \27505 , \27503 , \27504 );
nor \U$27508 ( \27506 , \27502 , \27505 );
buf \U$27509 ( \27507 , \27506 );
buf \U$27510 ( \27508 , \27507 );
not \U$27511 ( \27509 , \27508 );
or \U$27512 ( \27510 , \27465 , \27509 );
buf \U$27513 ( \27511 , \27507 );
buf \U$27514 ( \27512 , \27463 );
or \U$27515 ( \27513 , \27511 , \27512 );
nand \U$27516 ( \27514 , \27510 , \27513 );
buf \U$27517 ( \27515 , \27514 );
buf \U$27518 ( \27516 , \27515 );
buf \U$27519 ( \27517 , \26303 );
not \U$27520 ( \27518 , \27517 );
buf \U$27521 ( \27519 , \12736 );
not \U$27522 ( \27520 , \27519 );
or \U$27523 ( \27521 , \27518 , \27520 );
buf \U$27524 ( \27522 , \12744 );
buf \U$27525 ( \27523 , RIc0da738_105);
buf \U$27526 ( \27524 , RIc0d7d08_15);
xor \U$27527 ( \27525 , \27523 , \27524 );
buf \U$27528 ( \27526 , \27525 );
buf \U$27529 ( \27527 , \27526 );
nand \U$27530 ( \27528 , \27522 , \27527 );
buf \U$27531 ( \27529 , \27528 );
buf \U$27532 ( \27530 , \27529 );
nand \U$27533 ( \27531 , \27521 , \27530 );
buf \U$27534 ( \27532 , \27531 );
buf \U$27535 ( \27533 , \27532 );
buf \U$27536 ( \27534 , \26677 );
not \U$27537 ( \27535 , \27534 );
buf \U$27538 ( \27536 , \25542 );
not \U$27539 ( \27537 , \27536 );
or \U$27540 ( \27538 , \27535 , \27537 );
buf \U$27541 ( \27539 , \13953 );
buf \U$27542 ( \27540 , RIc0dadc8_119);
buf \U$27543 ( \27541 , RIc0d7678_1);
and \U$27544 ( \27542 , \27540 , \27541 );
not \U$27545 ( \27543 , \27540 );
buf \U$27546 ( \27544 , \974 );
and \U$27547 ( \27545 , \27543 , \27544 );
nor \U$27548 ( \27546 , \27542 , \27545 );
buf \U$27549 ( \27547 , \27546 );
buf \U$27550 ( \27548 , \27547 );
nand \U$27551 ( \27549 , \27539 , \27548 );
buf \U$27552 ( \27550 , \27549 );
buf \U$27553 ( \27551 , \27550 );
nand \U$27554 ( \27552 , \27538 , \27551 );
buf \U$27555 ( \27553 , \27552 );
buf \U$27556 ( \27554 , \27553 );
xor \U$27557 ( \27555 , \27533 , \27554 );
buf \U$27558 ( \27556 , \12975 );
not \U$27559 ( \27557 , \27556 );
buf \U$27560 ( \27558 , \27557 );
buf \U$27561 ( \27559 , \27558 );
not \U$27562 ( \27560 , \27559 );
buf \U$27563 ( \27561 , \12968 );
not \U$27564 ( \27562 , \27561 );
or \U$27565 ( \27563 , \27560 , \27562 );
buf \U$27566 ( \27564 , RIc0daeb8_121);
nand \U$27567 ( \27565 , \27563 , \27564 );
buf \U$27568 ( \27566 , \27565 );
buf \U$27569 ( \27567 , \27566 );
xor \U$27570 ( \27568 , \27555 , \27567 );
buf \U$27571 ( \27569 , \27568 );
buf \U$27572 ( \27570 , \27569 );
xor \U$27573 ( \27571 , \27516 , \27570 );
buf \U$27574 ( \27572 , \26523 );
not \U$27575 ( \27573 , \27572 );
buf \U$27576 ( \27574 , \18150 );
not \U$27577 ( \27575 , \27574 );
or \U$27578 ( \27576 , \27573 , \27575 );
buf \U$27579 ( \27577 , \442 );
buf \U$27580 ( \27578 , RIc0d8488_31);
buf \U$27581 ( \27579 , RIc0d9fb8_89);
xor \U$27582 ( \27580 , \27578 , \27579 );
buf \U$27583 ( \27581 , \27580 );
buf \U$27584 ( \27582 , \27581 );
nand \U$27585 ( \27583 , \27577 , \27582 );
buf \U$27586 ( \27584 , \27583 );
buf \U$27587 ( \27585 , \27584 );
nand \U$27588 ( \27586 , \27576 , \27585 );
buf \U$27589 ( \27587 , \27586 );
buf \U$27590 ( \27588 , \27587 );
buf \U$27591 ( \27589 , \26133 );
not \U$27592 ( \27590 , \27589 );
buf \U$27595 ( \27591 , \3714 );
buf \U$27596 ( \27592 , \27591 );
not \U$27597 ( \27593 , \27592 );
or \U$27598 ( \27594 , \27590 , \27593 );
buf \U$27599 ( \27595 , \344 );
xor \U$27600 ( \27596 , RIc0da288_95, RIc0d81b8_25);
buf \U$27601 ( \27597 , \27596 );
nand \U$27602 ( \27598 , \27595 , \27597 );
buf \U$27603 ( \27599 , \27598 );
buf \U$27604 ( \27600 , \27599 );
nand \U$27605 ( \27601 , \27594 , \27600 );
buf \U$27606 ( \27602 , \27601 );
buf \U$27607 ( \27603 , \27602 );
xor \U$27608 ( \27604 , \27588 , \27603 );
buf \U$27609 ( \27605 , \16575 );
buf \U$27610 ( \27606 , \26713 );
not \U$27611 ( \27607 , \27606 );
buf \U$27612 ( \27608 , \27607 );
buf \U$27613 ( \27609 , \27608 );
or \U$27614 ( \27610 , \27605 , \27609 );
buf \U$27615 ( \27611 , \4475 );
buf \U$27616 ( \27612 , RIc0da648_103);
buf \U$27617 ( \27613 , RIc0d7df8_17);
xor \U$27618 ( \27614 , \27612 , \27613 );
buf \U$27619 ( \27615 , \27614 );
buf \U$27620 ( \27616 , \27615 );
not \U$27621 ( \27617 , \27616 );
buf \U$27622 ( \27618 , \27617 );
buf \U$27623 ( \27619 , \27618 );
or \U$27624 ( \27620 , \27611 , \27619 );
nand \U$27625 ( \27621 , \27610 , \27620 );
buf \U$27626 ( \27622 , \27621 );
buf \U$27627 ( \27623 , \27622 );
xor \U$27628 ( \27624 , \27604 , \27623 );
buf \U$27629 ( \27625 , \27624 );
buf \U$27630 ( \27626 , \27625 );
xor \U$27631 ( \27627 , \27571 , \27626 );
buf \U$27632 ( \27628 , \27627 );
buf \U$27633 ( \27629 , \27628 );
xor \U$27634 ( \27630 , \27447 , \27629 );
buf \U$27635 ( \27631 , \27630 );
buf \U$27636 ( \27632 , \27631 );
xor \U$27637 ( \27633 , \26667 , \26736 );
and \U$27638 ( \27634 , \27633 , \26752 );
and \U$27639 ( \27635 , \26667 , \26736 );
or \U$27640 ( \27636 , \27634 , \27635 );
buf \U$27641 ( \27637 , \27636 );
buf \U$27642 ( \27638 , \27637 );
buf \U$27643 ( \27639 , \26451 );
not \U$27644 ( \27640 , \27639 );
buf \U$27645 ( \27641 , \12361 );
not \U$27646 ( \27642 , \27641 );
or \U$27647 ( \27643 , \27640 , \27642 );
buf \U$27648 ( \27644 , \3985 );
buf \U$27649 ( \27645 , RIc0d8938_41);
buf \U$27650 ( \27646 , RIc0d9b08_79);
xor \U$27651 ( \27647 , \27645 , \27646 );
buf \U$27652 ( \27648 , \27647 );
buf \U$27653 ( \27649 , \27648 );
nand \U$27654 ( \27650 , \27644 , \27649 );
buf \U$27655 ( \27651 , \27650 );
buf \U$27656 ( \27652 , \27651 );
nand \U$27657 ( \27653 , \27643 , \27652 );
buf \U$27658 ( \27654 , \27653 );
buf \U$27659 ( \27655 , \27654 );
buf \U$27660 ( \27656 , \26692 );
not \U$27661 ( \27657 , \27656 );
buf \U$27662 ( \27658 , \14207 );
not \U$27663 ( \27659 , \27658 );
buf \U$27664 ( \27660 , \27659 );
buf \U$27665 ( \27661 , \27660 );
not \U$27666 ( \27662 , \27661 );
or \U$27667 ( \27663 , \27657 , \27662 );
buf \U$27668 ( \27664 , \13426 );
xor \U$27669 ( \27665 , RIc0da918_109, RIc0d7b28_11);
buf \U$27670 ( \27666 , \27665 );
nand \U$27671 ( \27667 , \27664 , \27666 );
buf \U$27672 ( \27668 , \27667 );
buf \U$27673 ( \27669 , \27668 );
nand \U$27674 ( \27670 , \27663 , \27669 );
buf \U$27675 ( \27671 , \27670 );
buf \U$27676 ( \27672 , \27671 );
xor \U$27677 ( \27673 , \27655 , \27672 );
buf \U$27678 ( \27674 , \473 );
buf \U$27679 ( \27675 , \26150 );
or \U$27680 ( \27676 , \27674 , \27675 );
buf \U$27681 ( \27677 , \5886 );
buf \U$27682 ( \27678 , RIc0d82a8_27);
buf \U$27683 ( \27679 , RIc0da198_93);
xor \U$27684 ( \27680 , \27678 , \27679 );
buf \U$27685 ( \27681 , \27680 );
buf \U$27686 ( \27682 , \27681 );
not \U$27687 ( \27683 , \27682 );
buf \U$27688 ( \27684 , \27683 );
buf \U$27689 ( \27685 , \27684 );
or \U$27690 ( \27686 , \27677 , \27685 );
nand \U$27691 ( \27687 , \27676 , \27686 );
buf \U$27692 ( \27688 , \27687 );
buf \U$27693 ( \27689 , \27688 );
xor \U$27694 ( \27690 , \27673 , \27689 );
buf \U$27695 ( \27691 , \27690 );
buf \U$27696 ( \27692 , \27691 );
buf \U$27697 ( \27693 , \26340 );
not \U$27698 ( \27694 , \27693 );
buf \U$27699 ( \27695 , \4527 );
not \U$27700 ( \27696 , \27695 );
or \U$27701 ( \27697 , \27694 , \27696 );
buf \U$27702 ( \27698 , \14331 );
xor \U$27703 ( \27699 , RIc0d9ec8_87, RIc0d8578_33);
buf \U$27704 ( \27700 , \27699 );
nand \U$27705 ( \27701 , \27698 , \27700 );
buf \U$27706 ( \27702 , \27701 );
buf \U$27707 ( \27703 , \27702 );
nand \U$27708 ( \27704 , \27697 , \27703 );
buf \U$27709 ( \27705 , \27704 );
buf \U$27710 ( \27706 , \26359 );
not \U$27711 ( \27707 , \27706 );
buf \U$27712 ( \27708 , \3534 );
not \U$27713 ( \27709 , \27708 );
or \U$27714 ( \27710 , \27707 , \27709 );
buf \U$27715 ( \27711 , \16676 );
buf \U$27716 ( \27712 , RIc0da558_101);
buf \U$27717 ( \27713 , RIc0d7ee8_19);
xor \U$27718 ( \27714 , \27712 , \27713 );
buf \U$27719 ( \27715 , \27714 );
buf \U$27720 ( \27716 , \27715 );
nand \U$27721 ( \27717 , \27711 , \27716 );
buf \U$27722 ( \27718 , \27717 );
buf \U$27723 ( \27719 , \27718 );
nand \U$27724 ( \27720 , \27710 , \27719 );
buf \U$27725 ( \27721 , \27720 );
xor \U$27726 ( \27722 , \27705 , \27721 );
buf \U$27727 ( \27723 , \26116 );
not \U$27728 ( \27724 , \27723 );
buf \U$27729 ( \27725 , \18057 );
not \U$27730 ( \27726 , \27725 );
or \U$27731 ( \27727 , \27724 , \27726 );
buf \U$27732 ( \27728 , \791 );
xor \U$27733 ( \27729 , RIc0d9838_73, RIc0d8c08_47);
buf \U$27734 ( \27730 , \27729 );
nand \U$27735 ( \27731 , \27728 , \27730 );
buf \U$27736 ( \27732 , \27731 );
buf \U$27737 ( \27733 , \27732 );
nand \U$27738 ( \27734 , \27727 , \27733 );
buf \U$27739 ( \27735 , \27734 );
xor \U$27740 ( \27736 , \27722 , \27735 );
buf \U$27741 ( \27737 , \27736 );
xor \U$27742 ( \27738 , \27692 , \27737 );
buf \U$27743 ( \27739 , \26471 );
not \U$27744 ( \27740 , \27739 );
buf \U$27745 ( \27741 , \14681 );
not \U$27746 ( \27742 , \27741 );
buf \U$27747 ( \27743 , \27742 );
buf \U$27748 ( \27744 , \27743 );
not \U$27749 ( \27745 , \27744 );
or \U$27750 ( \27746 , \27740 , \27745 );
buf \U$27751 ( \27747 , \12303 );
buf \U$27752 ( \27748 , RIc0dabe8_115);
buf \U$27753 ( \27749 , RIc0d7858_5);
xor \U$27754 ( \27750 , \27748 , \27749 );
buf \U$27755 ( \27751 , \27750 );
buf \U$27756 ( \27752 , \27751 );
nand \U$27757 ( \27753 , \27747 , \27752 );
buf \U$27758 ( \27754 , \27753 );
buf \U$27759 ( \27755 , \27754 );
nand \U$27760 ( \27756 , \27746 , \27755 );
buf \U$27761 ( \27757 , \27756 );
buf \U$27762 ( \27758 , \26545 );
not \U$27763 ( \27759 , \27758 );
buf \U$27764 ( \27760 , \22350 );
not \U$27765 ( \27761 , \27760 );
or \U$27766 ( \27762 , \27759 , \27761 );
buf \U$27767 ( \27763 , \16559 );
buf \U$27768 ( \27764 , RIc0dacd8_117);
buf \U$27769 ( \27765 , RIc0d7768_3);
and \U$27770 ( \27766 , \27764 , \27765 );
not \U$27771 ( \27767 , \27764 );
buf \U$27772 ( \27768 , \304 );
and \U$27773 ( \27769 , \27767 , \27768 );
nor \U$27774 ( \27770 , \27766 , \27769 );
buf \U$27775 ( \27771 , \27770 );
buf \U$27776 ( \27772 , \27771 );
nand \U$27777 ( \27773 , \27763 , \27772 );
buf \U$27778 ( \27774 , \27773 );
buf \U$27779 ( \27775 , \27774 );
nand \U$27780 ( \27776 , \27762 , \27775 );
buf \U$27781 ( \27777 , \27776 );
xor \U$27782 ( \27778 , \27757 , \27777 );
buf \U$27783 ( \27779 , \26278 );
not \U$27784 ( \27780 , \27779 );
buf \U$27785 ( \27781 , \2766 );
not \U$27786 ( \27782 , \27781 );
or \U$27787 ( \27783 , \27780 , \27782 );
buf \U$27788 ( \27784 , \1078 );
buf \U$27789 ( \27785 , RIc0d9bf8_81);
buf \U$27790 ( \27786 , RIc0d8848_39);
xor \U$27791 ( \27787 , \27785 , \27786 );
buf \U$27792 ( \27788 , \27787 );
buf \U$27793 ( \27789 , \27788 );
nand \U$27794 ( \27790 , \27784 , \27789 );
buf \U$27795 ( \27791 , \27790 );
buf \U$27796 ( \27792 , \27791 );
nand \U$27797 ( \27793 , \27783 , \27792 );
buf \U$27798 ( \27794 , \27793 );
xor \U$27799 ( \27795 , \27778 , \27794 );
buf \U$27800 ( \27796 , \27795 );
xor \U$27801 ( \27797 , \27738 , \27796 );
buf \U$27802 ( \27798 , \27797 );
buf \U$27803 ( \27799 , \27798 );
xor \U$27804 ( \27800 , \27638 , \27799 );
xor \U$27805 ( \27801 , \26779 , \26785 );
and \U$27806 ( \27802 , \27801 , \26791 );
and \U$27807 ( \27803 , \26779 , \26785 );
or \U$27808 ( \27804 , \27802 , \27803 );
buf \U$27809 ( \27805 , \27804 );
buf \U$27810 ( \27806 , \27805 );
xor \U$27811 ( \27807 , \27800 , \27806 );
buf \U$27812 ( \27808 , \27807 );
buf \U$27813 ( \27809 , \27808 );
xor \U$27814 ( \27810 , \27632 , \27809 );
xor \U$27815 ( \27811 , \26755 , \26761 );
and \U$27816 ( \27812 , \27811 , \26794 );
and \U$27817 ( \27813 , \26755 , \26761 );
or \U$27818 ( \27814 , \27812 , \27813 );
buf \U$27819 ( \27815 , \27814 );
buf \U$27820 ( \27816 , \27815 );
xor \U$27821 ( \27817 , \27810 , \27816 );
buf \U$27822 ( \27818 , \27817 );
buf \U$27823 ( \27819 , \27818 );
xor \U$27824 ( \27820 , \27209 , \27819 );
xor \U$27825 ( \27821 , \26612 , \26797 );
and \U$27826 ( \27822 , \27821 , \26804 );
and \U$27827 ( \27823 , \26612 , \26797 );
or \U$27828 ( \27824 , \27822 , \27823 );
buf \U$27829 ( \27825 , \27824 );
buf \U$27830 ( \27826 , \27825 );
xor \U$27831 ( \27827 , \27820 , \27826 );
buf \U$27832 ( \27828 , \27827 );
buf \U$27833 ( \27829 , \27828 );
xor \U$27834 ( \27830 , \27077 , \27829 );
buf \U$27835 ( \27831 , \27830 );
buf \U$27836 ( \27832 , \27831 );
xor \U$27837 ( \27833 , \27002 , \27832 );
buf \U$27838 ( \27834 , \27833 );
buf \U$27839 ( \27835 , \27834 );
not \U$27840 ( \27836 , \27835 );
buf \U$27841 ( \27837 , \27836 );
buf \U$27842 ( \27838 , \27837 );
nand \U$27843 ( \27839 , \26977 , \27838 );
buf \U$27844 ( \27840 , \27839 );
buf \U$27845 ( \27841 , \27840 );
nand \U$27846 ( \27842 , \26955 , \27841 );
buf \U$27847 ( \27843 , \27842 );
buf \U$27848 ( \27844 , \27843 );
nor \U$27849 ( \27845 , \25933 , \27844 );
buf \U$27850 ( \27846 , \27845 );
buf \U$27851 ( \27847 , \27846 );
nand \U$27852 ( \27848 , \23757 , \27847 );
buf \U$27853 ( \27849 , \27848 );
buf \U$27854 ( \27850 , \27849 );
buf \U$27855 ( \27851 , RIc0d8758_37);
buf \U$27856 ( \27852 , RIc0d9bf8_81);
xor \U$27857 ( \27853 , \27851 , \27852 );
buf \U$27858 ( \27854 , \27853 );
buf \U$27859 ( \27855 , \27854 );
not \U$27860 ( \27856 , \27855 );
buf \U$27861 ( \27857 , \19544 );
not \U$27862 ( \27858 , \27857 );
or \U$27863 ( \27859 , \27856 , \27858 );
buf \U$27864 ( \27860 , \1078 );
buf \U$27865 ( \27861 , RIc0d86e0_36);
buf \U$27866 ( \27862 , RIc0d9bf8_81);
xor \U$27867 ( \27863 , \27861 , \27862 );
buf \U$27868 ( \27864 , \27863 );
buf \U$27869 ( \27865 , \27864 );
nand \U$27870 ( \27866 , \27860 , \27865 );
buf \U$27871 ( \27867 , \27866 );
buf \U$27872 ( \27868 , \27867 );
nand \U$27873 ( \27869 , \27859 , \27868 );
buf \U$27874 ( \27870 , \27869 );
not \U$27875 ( \27871 , \27870 );
buf \U$27876 ( \27872 , RIc0d8cf8_49);
buf \U$27877 ( \27873 , RIc0d9658_69);
xor \U$27878 ( \27874 , \27872 , \27873 );
buf \U$27879 ( \27875 , \27874 );
buf \U$27880 ( \27876 , \27875 );
not \U$27881 ( \27877 , \27876 );
buf \U$27882 ( \27878 , \13332 );
not \U$27883 ( \27879 , \27878 );
or \U$27884 ( \27880 , \27877 , \27879 );
buf \U$27885 ( \27881 , \283 );
buf \U$27886 ( \27882 , RIc0d8c80_48);
buf \U$27887 ( \27883 , RIc0d9658_69);
xor \U$27888 ( \27884 , \27882 , \27883 );
buf \U$27889 ( \27885 , \27884 );
buf \U$27890 ( \27886 , \27885 );
nand \U$27891 ( \27887 , \27881 , \27886 );
buf \U$27892 ( \27888 , \27887 );
buf \U$27893 ( \27889 , \27888 );
nand \U$27894 ( \27890 , \27880 , \27889 );
buf \U$27895 ( \27891 , \27890 );
not \U$27896 ( \27892 , \27891 );
or \U$27897 ( \27893 , \27871 , \27892 );
buf \U$27898 ( \27894 , \27870 );
buf \U$27899 ( \27895 , \27891 );
or \U$27900 ( \27896 , \27894 , \27895 );
buf \U$27901 ( \27897 , RIc0d8938_41);
buf \U$27902 ( \27898 , RIc0d9a18_77);
xor \U$27903 ( \27899 , \27897 , \27898 );
buf \U$27904 ( \27900 , \27899 );
buf \U$27905 ( \27901 , \27900 );
not \U$27906 ( \27902 , \27901 );
buf \U$27907 ( \27903 , \1431 );
not \U$27908 ( \27904 , \27903 );
or \U$27909 ( \27905 , \27902 , \27904 );
buf \U$27910 ( \27906 , \1196 );
buf \U$27911 ( \27907 , RIc0d88c0_40);
buf \U$27912 ( \27908 , RIc0d9a18_77);
xor \U$27913 ( \27909 , \27907 , \27908 );
buf \U$27914 ( \27910 , \27909 );
buf \U$27915 ( \27911 , \27910 );
nand \U$27916 ( \27912 , \27906 , \27911 );
buf \U$27917 ( \27913 , \27912 );
buf \U$27918 ( \27914 , \27913 );
nand \U$27919 ( \27915 , \27905 , \27914 );
buf \U$27920 ( \27916 , \27915 );
buf \U$27921 ( \27917 , \27916 );
nand \U$27922 ( \27918 , \27896 , \27917 );
buf \U$27923 ( \27919 , \27918 );
nand \U$27924 ( \27920 , \27893 , \27919 );
buf \U$27925 ( \27921 , \27920 );
buf \U$27926 ( \27922 , RIc0d8a28_43);
buf \U$27927 ( \27923 , RIc0d9928_75);
xor \U$27928 ( \27924 , \27922 , \27923 );
buf \U$27929 ( \27925 , \27924 );
buf \U$27930 ( \27926 , \27925 );
not \U$27931 ( \27927 , \27926 );
buf \U$27932 ( \27928 , \2358 );
not \U$27933 ( \27929 , \27928 );
or \U$27934 ( \27930 , \27927 , \27929 );
buf \U$27935 ( \27931 , \13998 );
xor \U$27936 ( \27932 , RIc0d9928_75, RIc0d89b0_42);
buf \U$27937 ( \27933 , \27932 );
nand \U$27938 ( \27934 , \27931 , \27933 );
buf \U$27939 ( \27935 , \27934 );
buf \U$27940 ( \27936 , \27935 );
nand \U$27941 ( \27937 , \27930 , \27936 );
buf \U$27942 ( \27938 , \27937 );
buf \U$27943 ( \27939 , \27938 );
not \U$27944 ( \27940 , \27939 );
buf \U$27945 ( \27941 , RIc0d7c18_13);
buf \U$27946 ( \27942 , RIc0da738_105);
xor \U$27947 ( \27943 , \27941 , \27942 );
buf \U$27948 ( \27944 , \27943 );
buf \U$27949 ( \27945 , \27944 );
not \U$27950 ( \27946 , \27945 );
buf \U$27951 ( \27947 , \14804 );
not \U$27952 ( \27948 , \27947 );
or \U$27953 ( \27949 , \27946 , \27948 );
buf \U$27954 ( \27950 , \26301 );
buf \U$27955 ( \27951 , RIc0d7ba0_12);
buf \U$27956 ( \27952 , RIc0da738_105);
xor \U$27957 ( \27953 , \27951 , \27952 );
buf \U$27958 ( \27954 , \27953 );
buf \U$27959 ( \27955 , \27954 );
nand \U$27960 ( \27956 , \27950 , \27955 );
buf \U$27961 ( \27957 , \27956 );
buf \U$27962 ( \27958 , \27957 );
nand \U$27963 ( \27959 , \27949 , \27958 );
buf \U$27964 ( \27960 , \27959 );
buf \U$27965 ( \27961 , \27960 );
not \U$27966 ( \27962 , \27961 );
or \U$27967 ( \27963 , \27940 , \27962 );
buf \U$27968 ( \27964 , \27938 );
buf \U$27969 ( \27965 , \27960 );
or \U$27970 ( \27966 , \27964 , \27965 );
buf \U$27971 ( \27967 , RIc0d7768_3);
buf \U$27972 ( \27968 , RIc0dabe8_115);
xor \U$27973 ( \27969 , \27967 , \27968 );
buf \U$27974 ( \27970 , \27969 );
buf \U$27975 ( \27971 , \27970 );
not \U$27976 ( \27972 , \27971 );
buf \U$27977 ( \27973 , \12299 );
not \U$27978 ( \27974 , \27973 );
or \U$27979 ( \27975 , \27972 , \27974 );
buf \U$27980 ( \27976 , \12303 );
buf \U$27981 ( \27977 , RIc0d76f0_2);
buf \U$27982 ( \27978 , RIc0dabe8_115);
xor \U$27983 ( \27979 , \27977 , \27978 );
buf \U$27984 ( \27980 , \27979 );
buf \U$27985 ( \27981 , \27980 );
nand \U$27986 ( \27982 , \27976 , \27981 );
buf \U$27987 ( \27983 , \27982 );
buf \U$27988 ( \27984 , \27983 );
nand \U$27989 ( \27985 , \27975 , \27984 );
buf \U$27990 ( \27986 , \27985 );
buf \U$27991 ( \27987 , \27986 );
nand \U$27992 ( \27988 , \27966 , \27987 );
buf \U$27993 ( \27989 , \27988 );
buf \U$27994 ( \27990 , \27989 );
nand \U$27995 ( \27991 , \27963 , \27990 );
buf \U$27996 ( \27992 , \27991 );
buf \U$27997 ( \27993 , \27992 );
xor \U$27998 ( \27994 , \27921 , \27993 );
buf \U$27999 ( \27995 , RIc0d9478_65);
buf \U$28000 ( \27996 , RIc0d8ed8_53);
and \U$28001 ( \27997 , \27995 , \27996 );
buf \U$28002 ( \27998 , \27997 );
buf \U$28003 ( \27999 , \27998 );
buf \U$28004 ( \28000 , RIc0d8d70_50);
buf \U$28005 ( \28001 , RIc0d9568_67);
xor \U$28006 ( \28002 , \28000 , \28001 );
buf \U$28007 ( \28003 , \28002 );
buf \U$28008 ( \28004 , \28003 );
not \U$28009 ( \28005 , \28004 );
buf \U$28010 ( \28006 , \2899 );
not \U$28011 ( \28007 , \28006 );
or \U$28012 ( \28008 , \28005 , \28007 );
buf \U$28013 ( \28009 , \686 );
buf \U$28014 ( \28010 , RIc0d8cf8_49);
buf \U$28015 ( \28011 , RIc0d9568_67);
xor \U$28016 ( \28012 , \28010 , \28011 );
buf \U$28017 ( \28013 , \28012 );
buf \U$28018 ( \28014 , \28013 );
nand \U$28019 ( \28015 , \28009 , \28014 );
buf \U$28020 ( \28016 , \28015 );
buf \U$28021 ( \28017 , \28016 );
nand \U$28022 ( \28018 , \28008 , \28017 );
buf \U$28023 ( \28019 , \28018 );
buf \U$28024 ( \28020 , \28019 );
xor \U$28025 ( \28021 , \27999 , \28020 );
xor \U$28026 ( \28022 , RIc0da0a8_91, RIc0d8230_26);
buf \U$28027 ( \28023 , \28022 );
not \U$28028 ( \28024 , \28023 );
buf \U$28029 ( \28025 , \704 );
not \U$28030 ( \28026 , \28025 );
or \U$28031 ( \28027 , \28024 , \28026 );
buf \U$28032 ( \28028 , \1933 );
xor \U$28033 ( \28029 , RIc0da0a8_91, RIc0d81b8_25);
buf \U$28034 ( \28030 , \28029 );
nand \U$28035 ( \28031 , \28028 , \28030 );
buf \U$28036 ( \28032 , \28031 );
buf \U$28037 ( \28033 , \28032 );
nand \U$28038 ( \28034 , \28027 , \28033 );
buf \U$28039 ( \28035 , \28034 );
buf \U$28040 ( \28036 , \28035 );
xor \U$28041 ( \28037 , \28021 , \28036 );
buf \U$28042 ( \28038 , \28037 );
buf \U$28043 ( \28039 , \28038 );
and \U$28044 ( \28040 , \27994 , \28039 );
and \U$28045 ( \28041 , \27921 , \27993 );
or \U$28046 ( \28042 , \28040 , \28041 );
buf \U$28047 ( \28043 , \28042 );
buf \U$28048 ( \28044 , \28043 );
buf \U$28049 ( \28045 , RIc0d9ce8_83);
buf \U$28050 ( \28046 , RIc0d85f0_34);
xor \U$28051 ( \28047 , \28045 , \28046 );
buf \U$28052 ( \28048 , \28047 );
buf \U$28053 ( \28049 , \28048 );
not \U$28054 ( \28050 , \28049 );
buf \U$28055 ( \28051 , \2088 );
not \U$28056 ( \28052 , \28051 );
or \U$28057 ( \28053 , \28050 , \28052 );
buf \U$28058 ( \28054 , \584 );
xor \U$28059 ( \28055 , RIc0d9ce8_83, RIc0d8578_33);
buf \U$28060 ( \28056 , \28055 );
nand \U$28061 ( \28057 , \28054 , \28056 );
buf \U$28062 ( \28058 , \28057 );
buf \U$28063 ( \28059 , \28058 );
nand \U$28064 ( \28060 , \28053 , \28059 );
buf \U$28065 ( \28061 , \28060 );
buf \U$28066 ( \28062 , \28061 );
buf \U$28067 ( \28063 , \27885 );
not \U$28068 ( \28064 , \28063 );
buf \U$28069 ( \28065 , \864 );
not \U$28070 ( \28066 , \28065 );
or \U$28071 ( \28067 , \28064 , \28066 );
buf \U$28072 ( \28068 , \21657 );
buf \U$28073 ( \28069 , RIc0d8c08_47);
buf \U$28074 ( \28070 , RIc0d9658_69);
xor \U$28075 ( \28071 , \28069 , \28070 );
buf \U$28076 ( \28072 , \28071 );
buf \U$28077 ( \28073 , \28072 );
nand \U$28078 ( \28074 , \28068 , \28073 );
buf \U$28079 ( \28075 , \28074 );
buf \U$28080 ( \28076 , \28075 );
nand \U$28081 ( \28077 , \28067 , \28076 );
buf \U$28082 ( \28078 , \28077 );
buf \U$28083 ( \28079 , \28078 );
xor \U$28084 ( \28080 , \28062 , \28079 );
buf \U$28085 ( \28081 , RIc0da828_107);
buf \U$28086 ( \28082 , RIc0d7ab0_10);
xnor \U$28087 ( \28083 , \28081 , \28082 );
buf \U$28088 ( \28084 , \28083 );
buf \U$28089 ( \28085 , \28084 );
not \U$28090 ( \28086 , \28085 );
buf \U$28091 ( \28087 , \28086 );
buf \U$28092 ( \28088 , \28087 );
not \U$28093 ( \28089 , \28088 );
buf \U$28094 ( \28090 , \17595 );
not \U$28095 ( \28091 , \28090 );
or \U$28096 ( \28092 , \28089 , \28091 );
buf \U$28097 ( \28093 , \12342 );
buf \U$28098 ( \28094 , RIc0d7a38_9);
buf \U$28099 ( \28095 , RIc0da828_107);
xor \U$28100 ( \28096 , \28094 , \28095 );
buf \U$28101 ( \28097 , \28096 );
buf \U$28102 ( \28098 , \28097 );
nand \U$28103 ( \28099 , \28093 , \28098 );
buf \U$28104 ( \28100 , \28099 );
buf \U$28105 ( \28101 , \28100 );
nand \U$28106 ( \28102 , \28092 , \28101 );
buf \U$28107 ( \28103 , \28102 );
buf \U$28108 ( \28104 , \28103 );
xor \U$28109 ( \28105 , \28080 , \28104 );
buf \U$28110 ( \28106 , \28105 );
not \U$28111 ( \28107 , \28106 );
buf \U$28112 ( \28108 , RIc0d9478_65);
buf \U$28113 ( \28109 , RIc0d8e60_52);
xor \U$28114 ( \28110 , \28108 , \28109 );
buf \U$28115 ( \28111 , \28110 );
buf \U$28116 ( \28112 , \28111 );
not \U$28117 ( \28113 , \28112 );
buf \U$28118 ( \28114 , \23253 );
not \U$28119 ( \28115 , \28114 );
or \U$28120 ( \28116 , \28113 , \28115 );
buf \U$28121 ( \28117 , \1229 );
buf \U$28122 ( \28118 , RIc0d9478_65);
buf \U$28123 ( \28119 , RIc0d8de8_51);
xor \U$28124 ( \28120 , \28118 , \28119 );
buf \U$28125 ( \28121 , \28120 );
buf \U$28126 ( \28122 , \28121 );
nand \U$28127 ( \28123 , \28117 , \28122 );
buf \U$28128 ( \28124 , \28123 );
buf \U$28129 ( \28125 , \28124 );
nand \U$28130 ( \28126 , \28116 , \28125 );
buf \U$28131 ( \28127 , \28126 );
buf \U$28132 ( \28128 , \28127 );
buf \U$28133 ( \28129 , RIc0d8b90_46);
buf \U$28134 ( \28130 , RIc0d9748_71);
xor \U$28135 ( \28131 , \28129 , \28130 );
buf \U$28136 ( \28132 , \28131 );
buf \U$28137 ( \28133 , \28132 );
not \U$28138 ( \28134 , \28133 );
buf \U$28139 ( \28135 , \12676 );
not \U$28140 ( \28136 , \28135 );
or \U$28141 ( \28137 , \28134 , \28136 );
buf \U$28142 ( \28138 , \2927 );
buf \U$28143 ( \28139 , RIc0d8b18_45);
buf \U$28144 ( \28140 , RIc0d9748_71);
xor \U$28145 ( \28141 , \28139 , \28140 );
buf \U$28146 ( \28142 , \28141 );
buf \U$28147 ( \28143 , \28142 );
nand \U$28148 ( \28144 , \28138 , \28143 );
buf \U$28149 ( \28145 , \28144 );
buf \U$28150 ( \28146 , \28145 );
nand \U$28151 ( \28147 , \28137 , \28146 );
buf \U$28152 ( \28148 , \28147 );
buf \U$28153 ( \28149 , \28148 );
xor \U$28154 ( \28150 , \28128 , \28149 );
buf \U$28155 ( \28151 , RIc0d7f60_20);
buf \U$28156 ( \28152 , RIc0da378_97);
xor \U$28157 ( \28153 , \28151 , \28152 );
buf \U$28158 ( \28154 , \28153 );
buf \U$28159 ( \28155 , \28154 );
not \U$28160 ( \28156 , \28155 );
buf \U$28161 ( \28157 , \15329 );
not \U$28162 ( \28158 , \28157 );
or \U$28163 ( \28159 , \28156 , \28158 );
buf \U$28164 ( \28160 , \2070 );
buf \U$28165 ( \28161 , RIc0d7ee8_19);
buf \U$28166 ( \28162 , RIc0da378_97);
xor \U$28167 ( \28163 , \28161 , \28162 );
buf \U$28168 ( \28164 , \28163 );
buf \U$28169 ( \28165 , \28164 );
nand \U$28170 ( \28166 , \28160 , \28165 );
buf \U$28171 ( \28167 , \28166 );
buf \U$28172 ( \28168 , \28167 );
nand \U$28173 ( \28169 , \28159 , \28168 );
buf \U$28174 ( \28170 , \28169 );
buf \U$28175 ( \28171 , \28170 );
xor \U$28176 ( \28172 , \28150 , \28171 );
buf \U$28177 ( \28173 , \28172 );
buf \U$28178 ( \28174 , \28173 );
not \U$28179 ( \28175 , \28174 );
buf \U$28180 ( \28176 , RIc0d7d80_16);
buf \U$28181 ( \28177 , RIc0da558_101);
xor \U$28182 ( \28178 , \28176 , \28177 );
buf \U$28183 ( \28179 , \28178 );
buf \U$28184 ( \28180 , \28179 );
not \U$28185 ( \28181 , \28180 );
buf \U$28186 ( \28182 , \20798 );
not \U$28187 ( \28183 , \28182 );
or \U$28188 ( \28184 , \28181 , \28183 );
buf \U$28189 ( \28185 , \15550 );
buf \U$28190 ( \28186 , RIc0d7d08_15);
buf \U$28191 ( \28187 , RIc0da558_101);
xor \U$28192 ( \28188 , \28186 , \28187 );
buf \U$28193 ( \28189 , \28188 );
buf \U$28194 ( \28190 , \28189 );
nand \U$28195 ( \28191 , \28185 , \28190 );
buf \U$28196 ( \28192 , \28191 );
buf \U$28197 ( \28193 , \28192 );
nand \U$28198 ( \28194 , \28184 , \28193 );
buf \U$28199 ( \28195 , \28194 );
buf \U$28200 ( \28196 , RIc0d8aa0_44);
buf \U$28201 ( \28197 , RIc0d9838_73);
xor \U$28202 ( \28198 , \28196 , \28197 );
buf \U$28203 ( \28199 , \28198 );
buf \U$28204 ( \28200 , \28199 );
not \U$28205 ( \28201 , \28200 );
buf \U$28206 ( \28202 , \14608 );
not \U$28207 ( \28203 , \28202 );
or \U$28208 ( \28204 , \28201 , \28203 );
buf \U$28209 ( \28205 , \791 );
buf \U$28210 ( \28206 , RIc0d8a28_43);
buf \U$28211 ( \28207 , RIc0d9838_73);
xor \U$28212 ( \28208 , \28206 , \28207 );
buf \U$28213 ( \28209 , \28208 );
buf \U$28214 ( \28210 , \28209 );
nand \U$28215 ( \28211 , \28205 , \28210 );
buf \U$28216 ( \28212 , \28211 );
buf \U$28217 ( \28213 , \28212 );
nand \U$28218 ( \28214 , \28204 , \28213 );
buf \U$28219 ( \28215 , \28214 );
buf \U$28220 ( \28216 , \28215 );
not \U$28221 ( \28217 , \28216 );
buf \U$28222 ( \28218 , \28217 );
and \U$28223 ( \28219 , \28195 , \28218 );
not \U$28224 ( \28220 , \28195 );
and \U$28225 ( \28221 , \28220 , \28215 );
or \U$28226 ( \28222 , \28219 , \28221 );
buf \U$28227 ( \28223 , \28222 );
buf \U$28228 ( \28224 , RIc0d8410_30);
buf \U$28229 ( \28225 , RIc0d9ec8_87);
xor \U$28230 ( \28226 , \28224 , \28225 );
buf \U$28231 ( \28227 , \28226 );
buf \U$28232 ( \28228 , \28227 );
not \U$28233 ( \28229 , \28228 );
buf \U$28234 ( \28230 , \14325 );
not \U$28235 ( \28231 , \28230 );
or \U$28236 ( \28232 , \28229 , \28231 );
buf \U$28237 ( \28233 , \14331 );
buf \U$28238 ( \28234 , RIc0d8398_29);
buf \U$28239 ( \28235 , RIc0d9ec8_87);
xor \U$28240 ( \28236 , \28234 , \28235 );
buf \U$28241 ( \28237 , \28236 );
buf \U$28242 ( \28238 , \28237 );
nand \U$28243 ( \28239 , \28233 , \28238 );
buf \U$28244 ( \28240 , \28239 );
buf \U$28245 ( \28241 , \28240 );
nand \U$28246 ( \28242 , \28232 , \28241 );
buf \U$28247 ( \28243 , \28242 );
buf \U$28248 ( \28244 , \28243 );
not \U$28249 ( \28245 , \28244 );
buf \U$28250 ( \28246 , \28245 );
buf \U$28251 ( \28247 , \28246 );
and \U$28252 ( \28248 , \28223 , \28247 );
not \U$28253 ( \28249 , \28223 );
buf \U$28254 ( \28250 , \28243 );
and \U$28255 ( \28251 , \28249 , \28250 );
nor \U$28256 ( \28252 , \28248 , \28251 );
buf \U$28257 ( \28253 , \28252 );
buf \U$28258 ( \28254 , \28253 );
nand \U$28259 ( \28255 , \28175 , \28254 );
buf \U$28260 ( \28256 , \28255 );
not \U$28261 ( \28257 , \28256 );
or \U$28262 ( \28258 , \28107 , \28257 );
buf \U$28263 ( \28259 , \28253 );
not \U$28264 ( \28260 , \28259 );
buf \U$28265 ( \28261 , \28173 );
nand \U$28266 ( \28262 , \28260 , \28261 );
buf \U$28267 ( \28263 , \28262 );
nand \U$28268 ( \28264 , \28258 , \28263 );
buf \U$28269 ( \28265 , \28264 );
xor \U$28270 ( \28266 , \28044 , \28265 );
buf \U$28271 ( \28267 , RIc0d8140_24);
buf \U$28272 ( \28268 , RIc0da198_93);
xor \U$28273 ( \28269 , \28267 , \28268 );
buf \U$28274 ( \28270 , \28269 );
buf \U$28275 ( \28271 , \28270 );
not \U$28276 ( \28272 , \28271 );
buf \U$28277 ( \28273 , \15995 );
not \U$28278 ( \28274 , \28273 );
or \U$28279 ( \28275 , \28272 , \28274 );
buf \U$28280 ( \28276 , \481 );
xor \U$28281 ( \28277 , RIc0da198_93, RIc0d80c8_23);
buf \U$28282 ( \28278 , \28277 );
nand \U$28283 ( \28279 , \28276 , \28278 );
buf \U$28284 ( \28280 , \28279 );
buf \U$28285 ( \28281 , \28280 );
nand \U$28286 ( \28282 , \28275 , \28281 );
buf \U$28287 ( \28283 , \28282 );
buf \U$28288 ( \28284 , \28283 );
xor \U$28289 ( \28285 , RIc0da918_109, RIc0d79c0_8);
buf \U$28290 ( \28286 , \28285 );
not \U$28291 ( \28287 , \28286 );
buf \U$28292 ( \28288 , \20759 );
not \U$28293 ( \28289 , \28288 );
or \U$28294 ( \28290 , \28287 , \28289 );
buf \U$28295 ( \28291 , \20211 );
xor \U$28296 ( \28292 , RIc0da918_109, RIc0d7948_7);
buf \U$28297 ( \28293 , \28292 );
nand \U$28298 ( \28294 , \28291 , \28293 );
buf \U$28299 ( \28295 , \28294 );
buf \U$28300 ( \28296 , \28295 );
nand \U$28301 ( \28297 , \28290 , \28296 );
buf \U$28302 ( \28298 , \28297 );
buf \U$28303 ( \28299 , \28298 );
xor \U$28304 ( \28300 , \28284 , \28299 );
buf \U$28305 ( \28301 , RIc0d9b08_79);
buf \U$28306 ( \28302 , RIc0d87d0_38);
xor \U$28307 ( \28303 , \28301 , \28302 );
buf \U$28308 ( \28304 , \28303 );
buf \U$28309 ( \28305 , \28304 );
not \U$28310 ( \28306 , \28305 );
buf \U$28311 ( \28307 , \1351 );
not \U$28312 ( \28308 , \28307 );
or \U$28313 ( \28309 , \28306 , \28308 );
buf \U$28314 ( \28310 , \1026 );
buf \U$28315 ( \28311 , RIc0d9b08_79);
buf \U$28316 ( \28312 , RIc0d8758_37);
xor \U$28317 ( \28313 , \28311 , \28312 );
buf \U$28318 ( \28314 , \28313 );
buf \U$28319 ( \28315 , \28314 );
nand \U$28320 ( \28316 , \28310 , \28315 );
buf \U$28321 ( \28317 , \28316 );
buf \U$28322 ( \28318 , \28317 );
nand \U$28323 ( \28319 , \28309 , \28318 );
buf \U$28324 ( \28320 , \28319 );
buf \U$28325 ( \28321 , \28320 );
xor \U$28326 ( \28322 , \28300 , \28321 );
buf \U$28327 ( \28323 , \28322 );
buf \U$28328 ( \28324 , \28323 );
buf \U$28329 ( \28325 , \27980 );
not \U$28330 ( \28326 , \28325 );
buf \U$28331 ( \28327 , \12299 );
not \U$28332 ( \28328 , \28327 );
or \U$28333 ( \28329 , \28326 , \28328 );
buf \U$28334 ( \28330 , \12303 );
buf \U$28335 ( \28331 , RIc0d7678_1);
buf \U$28336 ( \28332 , RIc0dabe8_115);
xor \U$28337 ( \28333 , \28331 , \28332 );
buf \U$28338 ( \28334 , \28333 );
buf \U$28339 ( \28335 , \28334 );
nand \U$28340 ( \28336 , \28330 , \28335 );
buf \U$28341 ( \28337 , \28336 );
buf \U$28342 ( \28338 , \28337 );
nand \U$28343 ( \28339 , \28329 , \28338 );
buf \U$28344 ( \28340 , \28339 );
buf \U$28345 ( \28341 , \28340 );
buf \U$28346 ( \28342 , \16556 );
not \U$28347 ( \28343 , \28342 );
buf \U$28348 ( \28344 , \12926 );
not \U$28349 ( \28345 , \28344 );
or \U$28350 ( \28346 , \28343 , \28345 );
buf \U$28351 ( \28347 , RIc0dacd8_117);
nand \U$28352 ( \28348 , \28346 , \28347 );
buf \U$28353 ( \28349 , \28348 );
buf \U$28354 ( \28350 , \28349 );
xor \U$28355 ( \28351 , \28341 , \28350 );
buf \U$28356 ( \28352 , \27864 );
not \U$28357 ( \28353 , \28352 );
buf \U$28358 ( \28354 , \17141 );
not \U$28359 ( \28355 , \28354 );
or \U$28360 ( \28356 , \28353 , \28355 );
buf \U$28361 ( \28357 , \1078 );
buf \U$28362 ( \28358 , RIc0d8668_35);
buf \U$28363 ( \28359 , RIc0d9bf8_81);
xor \U$28364 ( \28360 , \28358 , \28359 );
buf \U$28365 ( \28361 , \28360 );
buf \U$28366 ( \28362 , \28361 );
nand \U$28367 ( \28363 , \28357 , \28362 );
buf \U$28368 ( \28364 , \28363 );
buf \U$28369 ( \28365 , \28364 );
nand \U$28370 ( \28366 , \28356 , \28365 );
buf \U$28371 ( \28367 , \28366 );
buf \U$28372 ( \28368 , \28367 );
xor \U$28373 ( \28369 , \28351 , \28368 );
buf \U$28374 ( \28370 , \28369 );
buf \U$28375 ( \28371 , \28370 );
xor \U$28376 ( \28372 , \28324 , \28371 );
buf \U$28377 ( \28373 , \27932 );
not \U$28378 ( \28374 , \28373 );
buf \U$28379 ( \28375 , \2358 );
not \U$28380 ( \28376 , \28375 );
or \U$28381 ( \28377 , \28374 , \28376 );
buf \U$28382 ( \28378 , \16500 );
buf \U$28383 ( \28379 , RIc0d8938_41);
buf \U$28384 ( \28380 , RIc0d9928_75);
xor \U$28385 ( \28381 , \28379 , \28380 );
buf \U$28386 ( \28382 , \28381 );
buf \U$28387 ( \28383 , \28382 );
nand \U$28388 ( \28384 , \28378 , \28383 );
buf \U$28389 ( \28385 , \28384 );
buf \U$28390 ( \28386 , \28385 );
nand \U$28391 ( \28387 , \28377 , \28386 );
buf \U$28392 ( \28388 , \28387 );
buf \U$28393 ( \28389 , \28388 );
buf \U$28394 ( \28390 , \27910 );
not \U$28395 ( \28391 , \28390 );
buf \U$28396 ( \28392 , \1183 );
not \U$28397 ( \28393 , \28392 );
or \U$28398 ( \28394 , \28391 , \28393 );
buf \U$28399 ( \28395 , \3742 );
buf \U$28400 ( \28396 , RIc0d9a18_77);
buf \U$28401 ( \28397 , RIc0d8848_39);
xor \U$28402 ( \28398 , \28396 , \28397 );
buf \U$28403 ( \28399 , \28398 );
buf \U$28404 ( \28400 , \28399 );
nand \U$28405 ( \28401 , \28395 , \28400 );
buf \U$28406 ( \28402 , \28401 );
buf \U$28407 ( \28403 , \28402 );
nand \U$28408 ( \28404 , \28394 , \28403 );
buf \U$28409 ( \28405 , \28404 );
buf \U$28410 ( \28406 , \28405 );
xor \U$28411 ( \28407 , \28389 , \28406 );
xor \U$28412 ( \28408 , RIc0daaf8_113, RIc0d77e0_4);
buf \U$28413 ( \28409 , \28408 );
not \U$28414 ( \28410 , \28409 );
buf \U$28415 ( \28411 , \14888 );
not \U$28416 ( \28412 , \28411 );
buf \U$28417 ( \28413 , \28412 );
buf \U$28418 ( \28414 , \28413 );
not \U$28419 ( \28415 , \28414 );
or \U$28420 ( \28416 , \28410 , \28415 );
buf \U$28421 ( \28417 , \16662 );
buf \U$28422 ( \28418 , RIc0daaf8_113);
buf \U$28423 ( \28419 , RIc0d7768_3);
xor \U$28424 ( \28420 , \28418 , \28419 );
buf \U$28425 ( \28421 , \28420 );
buf \U$28426 ( \28422 , \28421 );
nand \U$28427 ( \28423 , \28417 , \28422 );
buf \U$28428 ( \28424 , \28423 );
buf \U$28429 ( \28425 , \28424 );
nand \U$28430 ( \28426 , \28416 , \28425 );
buf \U$28431 ( \28427 , \28426 );
buf \U$28432 ( \28428 , \28427 );
xor \U$28433 ( \28429 , \28407 , \28428 );
buf \U$28434 ( \28430 , \28429 );
buf \U$28435 ( \28431 , \28430 );
and \U$28436 ( \28432 , \28372 , \28431 );
and \U$28437 ( \28433 , \28324 , \28371 );
or \U$28438 ( \28434 , \28432 , \28433 );
buf \U$28439 ( \28435 , \28434 );
buf \U$28440 ( \28436 , \28435 );
and \U$28441 ( \28437 , \28266 , \28436 );
and \U$28442 ( \28438 , \28044 , \28265 );
or \U$28443 ( \28439 , \28437 , \28438 );
buf \U$28444 ( \28440 , \28439 );
buf \U$28445 ( \28441 , \28440 );
buf \U$28446 ( \28442 , \28218 );
not \U$28447 ( \28443 , \28442 );
buf \U$28448 ( \28444 , \28246 );
not \U$28449 ( \28445 , \28444 );
or \U$28450 ( \28446 , \28443 , \28445 );
buf \U$28451 ( \28447 , \28195 );
nand \U$28452 ( \28448 , \28446 , \28447 );
buf \U$28453 ( \28449 , \28448 );
buf \U$28454 ( \28450 , \28449 );
buf \U$28455 ( \28451 , \28243 );
buf \U$28456 ( \28452 , \28215 );
nand \U$28457 ( \28453 , \28451 , \28452 );
buf \U$28458 ( \28454 , \28453 );
buf \U$28459 ( \28455 , \28454 );
nand \U$28460 ( \28456 , \28450 , \28455 );
buf \U$28461 ( \28457 , \28456 );
buf \U$28462 ( \28458 , \28457 );
buf \U$28463 ( \28459 , \28367 );
buf \U$28464 ( \28460 , \28340 );
or \U$28465 ( \28461 , \28459 , \28460 );
buf \U$28466 ( \28462 , \28349 );
nand \U$28467 ( \28463 , \28461 , \28462 );
buf \U$28468 ( \28464 , \28463 );
buf \U$28469 ( \28465 , \28464 );
buf \U$28470 ( \28466 , \28367 );
buf \U$28471 ( \28467 , \28340 );
nand \U$28472 ( \28468 , \28466 , \28467 );
buf \U$28473 ( \28469 , \28468 );
buf \U$28474 ( \28470 , \28469 );
nand \U$28475 ( \28471 , \28465 , \28470 );
buf \U$28476 ( \28472 , \28471 );
buf \U$28477 ( \28473 , \28472 );
xor \U$28478 ( \28474 , \28458 , \28473 );
buf \U$28479 ( \28475 , RIc0d8320_28);
buf \U$28480 ( \28476 , RIc0d9fb8_89);
xor \U$28481 ( \28477 , \28475 , \28476 );
buf \U$28482 ( \28478 , \28477 );
buf \U$28483 ( \28479 , \28478 );
not \U$28484 ( \28480 , \28479 );
buf \U$28485 ( \28481 , \436 );
not \U$28486 ( \28482 , \28481 );
or \U$28487 ( \28483 , \28480 , \28482 );
buf \U$28488 ( \28484 , \442 );
buf \U$28489 ( \28485 , RIc0d82a8_27);
buf \U$28490 ( \28486 , RIc0d9fb8_89);
xor \U$28491 ( \28487 , \28485 , \28486 );
buf \U$28492 ( \28488 , \28487 );
buf \U$28493 ( \28489 , \28488 );
nand \U$28494 ( \28490 , \28484 , \28489 );
buf \U$28495 ( \28491 , \28490 );
buf \U$28496 ( \28492 , \28491 );
nand \U$28497 ( \28493 , \28483 , \28492 );
buf \U$28498 ( \28494 , \28493 );
buf \U$28499 ( \28495 , \28494 );
xor \U$28500 ( \28496 , RIc0da288_95, RIc0d8050_22);
buf \U$28501 ( \28497 , \28496 );
not \U$28502 ( \28498 , \28497 );
buf \U$28503 ( \28499 , \330 );
not \U$28504 ( \28500 , \28499 );
or \U$28505 ( \28501 , \28498 , \28500 );
buf \U$28506 ( \28502 , \14707 );
buf \U$28507 ( \28503 , RIc0da288_95);
buf \U$28508 ( \28504 , RIc0d7fd8_21);
xor \U$28509 ( \28505 , \28503 , \28504 );
buf \U$28510 ( \28506 , \28505 );
buf \U$28511 ( \28507 , \28506 );
nand \U$28512 ( \28508 , \28502 , \28507 );
buf \U$28513 ( \28509 , \28508 );
buf \U$28514 ( \28510 , \28509 );
nand \U$28515 ( \28511 , \28501 , \28510 );
buf \U$28516 ( \28512 , \28511 );
buf \U$28517 ( \28513 , \28512 );
xor \U$28518 ( \28514 , \28495 , \28513 );
buf \U$28519 ( \28515 , RIc0da648_103);
buf \U$28520 ( \28516 , RIc0d7c90_14);
xnor \U$28521 ( \28517 , \28515 , \28516 );
buf \U$28522 ( \28518 , \28517 );
buf \U$28523 ( \28519 , \28518 );
not \U$28524 ( \28520 , \28519 );
buf \U$28525 ( \28521 , \28520 );
buf \U$28526 ( \28522 , \28521 );
not \U$28527 ( \28523 , \28522 );
buf \U$28528 ( \28524 , \16578 );
not \U$28529 ( \28525 , \28524 );
or \U$28530 ( \28526 , \28523 , \28525 );
buf \U$28531 ( \28527 , \16584 );
buf \U$28532 ( \28528 , RIc0d7c18_13);
buf \U$28533 ( \28529 , RIc0da648_103);
xor \U$28534 ( \28530 , \28528 , \28529 );
buf \U$28535 ( \28531 , \28530 );
buf \U$28536 ( \28532 , \28531 );
nand \U$28537 ( \28533 , \28527 , \28532 );
buf \U$28538 ( \28534 , \28533 );
buf \U$28539 ( \28535 , \28534 );
nand \U$28540 ( \28536 , \28526 , \28535 );
buf \U$28541 ( \28537 , \28536 );
buf \U$28542 ( \28538 , \28537 );
and \U$28543 ( \28539 , \28514 , \28538 );
and \U$28544 ( \28540 , \28495 , \28513 );
or \U$28545 ( \28541 , \28539 , \28540 );
buf \U$28546 ( \28542 , \28541 );
buf \U$28547 ( \28543 , \28542 );
xor \U$28548 ( \28544 , \28474 , \28543 );
buf \U$28549 ( \28545 , \28544 );
buf \U$28550 ( \28546 , \28545 );
not \U$28551 ( \28547 , \28546 );
buf \U$28552 ( \28548 , \28547 );
buf \U$28553 ( \28549 , \28548 );
not \U$28554 ( \28550 , \28549 );
xor \U$28555 ( \28551 , \28284 , \28299 );
and \U$28556 ( \28552 , \28551 , \28321 );
and \U$28557 ( \28553 , \28284 , \28299 );
or \U$28558 ( \28554 , \28552 , \28553 );
buf \U$28559 ( \28555 , \28554 );
buf \U$28560 ( \28556 , RIc0d8500_32);
buf \U$28561 ( \28557 , RIc0d9dd8_85);
xor \U$28562 ( \28558 , \28556 , \28557 );
buf \U$28563 ( \28559 , \28558 );
buf \U$28564 ( \28560 , \28559 );
not \U$28565 ( \28561 , \28560 );
buf \U$28566 ( \28562 , \1389 );
not \U$28567 ( \28563 , \28562 );
or \U$28568 ( \28564 , \28561 , \28563 );
buf \U$28569 ( \28565 , \1401 );
buf \U$28570 ( \28566 , RIc0d9dd8_85);
buf \U$28571 ( \28567 , RIc0d8488_31);
xor \U$28572 ( \28568 , \28566 , \28567 );
buf \U$28573 ( \28569 , \28568 );
buf \U$28574 ( \28570 , \28569 );
nand \U$28575 ( \28571 , \28565 , \28570 );
buf \U$28576 ( \28572 , \28571 );
buf \U$28577 ( \28573 , \28572 );
nand \U$28578 ( \28574 , \28564 , \28573 );
buf \U$28579 ( \28575 , \28574 );
buf \U$28580 ( \28576 , \28575 );
not \U$28581 ( \28577 , \28576 );
buf \U$28582 ( \28578 , RIc0d78d0_6);
buf \U$28583 ( \28579 , RIc0daa08_111);
xor \U$28584 ( \28580 , \28578 , \28579 );
buf \U$28585 ( \28581 , \28580 );
buf \U$28586 ( \28582 , \28581 );
not \U$28587 ( \28583 , \28582 );
buf \U$28588 ( \28584 , \14100 );
not \U$28589 ( \28585 , \28584 );
or \U$28590 ( \28586 , \28583 , \28585 );
buf \U$28591 ( \28587 , \14353 );
buf \U$28592 ( \28588 , RIc0d7858_5);
buf \U$28593 ( \28589 , RIc0daa08_111);
xor \U$28594 ( \28590 , \28588 , \28589 );
buf \U$28595 ( \28591 , \28590 );
buf \U$28596 ( \28592 , \28591 );
nand \U$28597 ( \28593 , \28587 , \28592 );
buf \U$28598 ( \28594 , \28593 );
buf \U$28599 ( \28595 , \28594 );
nand \U$28600 ( \28596 , \28586 , \28595 );
buf \U$28601 ( \28597 , \28596 );
buf \U$28602 ( \28598 , \28597 );
not \U$28603 ( \28599 , \28598 );
or \U$28604 ( \28600 , \28577 , \28599 );
buf \U$28605 ( \28601 , \28575 );
buf \U$28606 ( \28602 , \28597 );
or \U$28607 ( \28603 , \28601 , \28602 );
xor \U$28608 ( \28604 , RIc0da468_99, RIc0d7e70_18);
buf \U$28609 ( \28605 , \28604 );
not \U$28610 ( \28606 , \28605 );
buf \U$28611 ( \28607 , \12578 );
not \U$28612 ( \28608 , \28607 );
or \U$28613 ( \28609 , \28606 , \28608 );
buf \U$28614 ( \28610 , \12584 );
xor \U$28615 ( \28611 , RIc0da468_99, RIc0d7df8_17);
buf \U$28616 ( \28612 , \28611 );
nand \U$28617 ( \28613 , \28610 , \28612 );
buf \U$28618 ( \28614 , \28613 );
buf \U$28619 ( \28615 , \28614 );
nand \U$28620 ( \28616 , \28609 , \28615 );
buf \U$28621 ( \28617 , \28616 );
buf \U$28622 ( \28618 , \28617 );
nand \U$28623 ( \28619 , \28603 , \28618 );
buf \U$28624 ( \28620 , \28619 );
buf \U$28625 ( \28621 , \28620 );
nand \U$28626 ( \28622 , \28600 , \28621 );
buf \U$28627 ( \28623 , \28622 );
xor \U$28628 ( \28624 , \28555 , \28623 );
xor \U$28629 ( \28625 , \28389 , \28406 );
and \U$28630 ( \28626 , \28625 , \28428 );
and \U$28631 ( \28627 , \28389 , \28406 );
or \U$28632 ( \28628 , \28626 , \28627 );
buf \U$28633 ( \28629 , \28628 );
xnor \U$28634 ( \28630 , \28624 , \28629 );
buf \U$28635 ( \28631 , \28630 );
not \U$28636 ( \28632 , \28631 );
or \U$28637 ( \28633 , \28550 , \28632 );
xor \U$28638 ( \28634 , \27999 , \28020 );
and \U$28639 ( \28635 , \28634 , \28036 );
and \U$28640 ( \28636 , \27999 , \28020 );
or \U$28641 ( \28637 , \28635 , \28636 );
buf \U$28642 ( \28638 , \28637 );
xor \U$28643 ( \28639 , \28128 , \28149 );
and \U$28644 ( \28640 , \28639 , \28171 );
and \U$28645 ( \28641 , \28128 , \28149 );
or \U$28646 ( \28642 , \28640 , \28641 );
buf \U$28647 ( \28643 , \28642 );
buf \U$28648 ( \28644 , \28643 );
not \U$28649 ( \28645 , \28644 );
buf \U$28650 ( \28646 , \28645 );
and \U$28651 ( \28647 , \28638 , \28646 );
not \U$28652 ( \28648 , \28638 );
and \U$28653 ( \28649 , \28648 , \28643 );
or \U$28654 ( \28650 , \28647 , \28649 );
buf \U$28655 ( \28651 , \28650 );
xor \U$28656 ( \28652 , \28062 , \28079 );
and \U$28657 ( \28653 , \28652 , \28104 );
and \U$28658 ( \28654 , \28062 , \28079 );
or \U$28659 ( \28655 , \28653 , \28654 );
buf \U$28660 ( \28656 , \28655 );
buf \U$28661 ( \28657 , \28656 );
not \U$28662 ( \28658 , \28657 );
buf \U$28663 ( \28659 , \28658 );
buf \U$28664 ( \28660 , \28659 );
and \U$28665 ( \28661 , \28651 , \28660 );
not \U$28666 ( \28662 , \28651 );
buf \U$28667 ( \28663 , \28656 );
and \U$28668 ( \28664 , \28662 , \28663 );
nor \U$28669 ( \28665 , \28661 , \28664 );
buf \U$28670 ( \28666 , \28665 );
buf \U$28671 ( \28667 , \28666 );
not \U$28672 ( \28668 , \28667 );
buf \U$28673 ( \28669 , \28668 );
buf \U$28674 ( \28670 , \28669 );
nand \U$28675 ( \28671 , \28633 , \28670 );
buf \U$28676 ( \28672 , \28671 );
buf \U$28677 ( \28673 , \28672 );
buf \U$28678 ( \28674 , \28630 );
not \U$28679 ( \28675 , \28674 );
buf \U$28680 ( \28676 , \28675 );
buf \U$28681 ( \28677 , \28676 );
buf \U$28682 ( \28678 , \28545 );
nand \U$28683 ( \28679 , \28677 , \28678 );
buf \U$28684 ( \28680 , \28679 );
buf \U$28685 ( \28681 , \28680 );
nand \U$28686 ( \28682 , \28673 , \28681 );
buf \U$28687 ( \28683 , \28682 );
buf \U$28688 ( \28684 , \28683 );
xor \U$28689 ( \28685 , \28441 , \28684 );
buf \U$28690 ( \28686 , \28591 );
not \U$28691 ( \28687 , \28686 );
buf \U$28692 ( \28688 , \14346 );
not \U$28693 ( \28689 , \28688 );
or \U$28694 ( \28690 , \28687 , \28689 );
buf \U$28695 ( \28691 , \14352 );
xor \U$28696 ( \28692 , RIc0daa08_111, RIc0d77e0_4);
buf \U$28697 ( \28693 , \28692 );
nand \U$28698 ( \28694 , \28691 , \28693 );
buf \U$28699 ( \28695 , \28694 );
buf \U$28700 ( \28696 , \28695 );
nand \U$28701 ( \28697 , \28690 , \28696 );
buf \U$28702 ( \28698 , \28697 );
buf \U$28703 ( \28699 , \28698 );
buf \U$28704 ( \28700 , \28611 );
not \U$28705 ( \28701 , \28700 );
buf \U$28706 ( \28702 , \14419 );
not \U$28707 ( \28703 , \28702 );
or \U$28708 ( \28704 , \28701 , \28703 );
buf \U$28709 ( \28705 , \12584 );
buf \U$28710 ( \28706 , RIc0d7d80_16);
buf \U$28711 ( \28707 , RIc0da468_99);
xor \U$28712 ( \28708 , \28706 , \28707 );
buf \U$28713 ( \28709 , \28708 );
buf \U$28714 ( \28710 , \28709 );
nand \U$28715 ( \28711 , \28705 , \28710 );
buf \U$28716 ( \28712 , \28711 );
buf \U$28717 ( \28713 , \28712 );
nand \U$28718 ( \28714 , \28704 , \28713 );
buf \U$28719 ( \28715 , \28714 );
buf \U$28720 ( \28716 , \28715 );
and \U$28721 ( \28717 , \28699 , \28716 );
not \U$28722 ( \28718 , \28699 );
buf \U$28723 ( \28719 , \28715 );
not \U$28724 ( \28720 , \28719 );
buf \U$28725 ( \28721 , \28720 );
buf \U$28726 ( \28722 , \28721 );
and \U$28727 ( \28723 , \28718 , \28722 );
nor \U$28728 ( \28724 , \28717 , \28723 );
buf \U$28729 ( \28725 , \28724 );
buf \U$28730 ( \28726 , \28725 );
buf \U$28731 ( \28727 , \28142 );
not \U$28732 ( \28728 , \28727 );
buf \U$28733 ( \28729 , \1263 );
not \U$28734 ( \28730 , \28729 );
or \U$28735 ( \28731 , \28728 , \28730 );
buf \U$28736 ( \28732 , \1282 );
xor \U$28737 ( \28733 , RIc0d9748_71, RIc0d8aa0_44);
buf \U$28738 ( \28734 , \28733 );
nand \U$28739 ( \28735 , \28732 , \28734 );
buf \U$28740 ( \28736 , \28735 );
buf \U$28741 ( \28737 , \28736 );
nand \U$28742 ( \28738 , \28731 , \28737 );
buf \U$28743 ( \28739 , \28738 );
buf \U$28744 ( \28740 , \28739 );
not \U$28745 ( \28741 , \28740 );
buf \U$28746 ( \28742 , \28741 );
buf \U$28747 ( \28743 , \28742 );
and \U$28748 ( \28744 , \28726 , \28743 );
not \U$28749 ( \28745 , \28726 );
buf \U$28750 ( \28746 , \28739 );
and \U$28751 ( \28747 , \28745 , \28746 );
nor \U$28752 ( \28748 , \28744 , \28747 );
buf \U$28753 ( \28749 , \28748 );
buf \U$28754 ( \28750 , \28749 );
not \U$28755 ( \28751 , \28750 );
buf \U$28756 ( \28752 , \28751 );
buf \U$28757 ( \28753 , \28752 );
not \U$28758 ( \28754 , \28753 );
buf \U$28759 ( \28755 , \28382 );
not \U$28760 ( \28756 , \28755 );
buf \U$28761 ( \28757 , \16494 );
not \U$28762 ( \28758 , \28757 );
or \U$28763 ( \28759 , \28756 , \28758 );
buf \U$28764 ( \28760 , \1565 );
buf \U$28765 ( \28761 , RIc0d88c0_40);
buf \U$28766 ( \28762 , RIc0d9928_75);
xor \U$28767 ( \28763 , \28761 , \28762 );
buf \U$28768 ( \28764 , \28763 );
buf \U$28769 ( \28765 , \28764 );
nand \U$28770 ( \28766 , \28760 , \28765 );
buf \U$28771 ( \28767 , \28766 );
buf \U$28772 ( \28768 , \28767 );
nand \U$28773 ( \28769 , \28759 , \28768 );
buf \U$28774 ( \28770 , \28769 );
buf \U$28775 ( \28771 , \28770 );
buf \U$28776 ( \28772 , \28421 );
not \U$28777 ( \28773 , \28772 );
buf \U$28778 ( \28774 , \14888 );
not \U$28779 ( \28775 , \28774 );
buf \U$28780 ( \28776 , \28775 );
buf \U$28781 ( \28777 , \28776 );
not \U$28782 ( \28778 , \28777 );
or \U$28783 ( \28779 , \28773 , \28778 );
buf \U$28784 ( \28780 , \14405 );
xor \U$28785 ( \28781 , RIc0daaf8_113, RIc0d76f0_2);
buf \U$28786 ( \28782 , \28781 );
nand \U$28787 ( \28783 , \28780 , \28782 );
buf \U$28788 ( \28784 , \28783 );
buf \U$28789 ( \28785 , \28784 );
nand \U$28790 ( \28786 , \28779 , \28785 );
buf \U$28791 ( \28787 , \28786 );
buf \U$28792 ( \28788 , \28787 );
xor \U$28793 ( \28789 , \28771 , \28788 );
buf \U$28794 ( \28790 , \28097 );
not \U$28795 ( \28791 , \28790 );
buf \U$28796 ( \28792 , \12331 );
not \U$28797 ( \28793 , \28792 );
buf \U$28798 ( \28794 , \28793 );
buf \U$28799 ( \28795 , \28794 );
not \U$28800 ( \28796 , \28795 );
or \U$28801 ( \28797 , \28791 , \28796 );
buf \U$28802 ( \28798 , \12342 );
buf \U$28803 ( \28799 , RIc0da828_107);
buf \U$28804 ( \28800 , RIc0d79c0_8);
xor \U$28805 ( \28801 , \28799 , \28800 );
buf \U$28806 ( \28802 , \28801 );
buf \U$28807 ( \28803 , \28802 );
nand \U$28808 ( \28804 , \28798 , \28803 );
buf \U$28809 ( \28805 , \28804 );
buf \U$28810 ( \28806 , \28805 );
nand \U$28811 ( \28807 , \28797 , \28806 );
buf \U$28812 ( \28808 , \28807 );
buf \U$28813 ( \28809 , \28808 );
not \U$28814 ( \28810 , \28809 );
buf \U$28815 ( \28811 , \28810 );
buf \U$28816 ( \28812 , \28811 );
xor \U$28817 ( \28813 , \28789 , \28812 );
buf \U$28818 ( \28814 , \28813 );
buf \U$28819 ( \28815 , \28814 );
not \U$28820 ( \28816 , \28815 );
buf \U$28821 ( \28817 , \28816 );
buf \U$28822 ( \28818 , \28817 );
not \U$28823 ( \28819 , \28818 );
or \U$28824 ( \28820 , \28754 , \28819 );
buf \U$28825 ( \28821 , \28749 );
not \U$28826 ( \28822 , \28821 );
buf \U$28827 ( \28823 , \28814 );
not \U$28828 ( \28824 , \28823 );
or \U$28829 ( \28825 , \28822 , \28824 );
buf \U$28830 ( \28826 , \28277 );
not \U$28831 ( \28827 , \28826 );
buf \U$28832 ( \28828 , \1901 );
not \U$28833 ( \28829 , \28828 );
or \U$28834 ( \28830 , \28827 , \28829 );
buf \U$28835 ( \28831 , \4008 );
buf \U$28836 ( \28832 , RIc0d8050_22);
buf \U$28837 ( \28833 , RIc0da198_93);
xor \U$28838 ( \28834 , \28832 , \28833 );
buf \U$28839 ( \28835 , \28834 );
buf \U$28840 ( \28836 , \28835 );
nand \U$28841 ( \28837 , \28831 , \28836 );
buf \U$28842 ( \28838 , \28837 );
buf \U$28843 ( \28839 , \28838 );
nand \U$28844 ( \28840 , \28830 , \28839 );
buf \U$28845 ( \28841 , \28840 );
buf \U$28846 ( \28842 , \28841 );
buf \U$28847 ( \28843 , \28029 );
not \U$28848 ( \28844 , \28843 );
buf \U$28849 ( \28845 , \2535 );
not \U$28850 ( \28846 , \28845 );
or \U$28851 ( \28847 , \28844 , \28846 );
buf \U$28852 ( \28848 , RIc0da0a8_91);
buf \U$28853 ( \28849 , RIc0d8140_24);
xnor \U$28854 ( \28850 , \28848 , \28849 );
buf \U$28855 ( \28851 , \28850 );
buf \U$28856 ( \28852 , \28851 );
not \U$28857 ( \28853 , \28852 );
buf \U$28858 ( \28854 , \714 );
nand \U$28859 ( \28855 , \28853 , \28854 );
buf \U$28860 ( \28856 , \28855 );
buf \U$28861 ( \28857 , \28856 );
nand \U$28862 ( \28858 , \28847 , \28857 );
buf \U$28863 ( \28859 , \28858 );
buf \U$28864 ( \28860 , \28859 );
xor \U$28865 ( \28861 , \28842 , \28860 );
buf \U$28866 ( \28862 , \28569 );
not \U$28867 ( \28863 , \28862 );
buf \U$28868 ( \28864 , \1389 );
not \U$28869 ( \28865 , \28864 );
or \U$28870 ( \28866 , \28863 , \28865 );
buf \U$28871 ( \28867 , RIc0d8410_30);
buf \U$28872 ( \28868 , RIc0d9dd8_85);
xnor \U$28873 ( \28869 , \28867 , \28868 );
buf \U$28874 ( \28870 , \28869 );
buf \U$28875 ( \28871 , \28870 );
not \U$28876 ( \28872 , \28871 );
buf \U$28877 ( \28873 , \2960 );
nand \U$28878 ( \28874 , \28872 , \28873 );
buf \U$28879 ( \28875 , \28874 );
buf \U$28880 ( \28876 , \28875 );
nand \U$28881 ( \28877 , \28866 , \28876 );
buf \U$28882 ( \28878 , \28877 );
buf \U$28883 ( \28879 , \28878 );
xor \U$28884 ( \28880 , \28861 , \28879 );
buf \U$28885 ( \28881 , \28880 );
buf \U$28886 ( \28882 , \28881 );
nand \U$28887 ( \28883 , \28825 , \28882 );
buf \U$28888 ( \28884 , \28883 );
buf \U$28889 ( \28885 , \28884 );
nand \U$28890 ( \28886 , \28820 , \28885 );
buf \U$28891 ( \28887 , \28886 );
buf \U$28892 ( \28888 , \28013 );
not \U$28893 ( \28889 , \28888 );
buf \U$28894 ( \28890 , \2899 );
not \U$28895 ( \28891 , \28890 );
or \U$28896 ( \28892 , \28889 , \28891 );
buf \U$28897 ( \28893 , \686 );
buf \U$28898 ( \28894 , RIc0d8c80_48);
buf \U$28899 ( \28895 , RIc0d9568_67);
xor \U$28900 ( \28896 , \28894 , \28895 );
buf \U$28901 ( \28897 , \28896 );
buf \U$28902 ( \28898 , \28897 );
nand \U$28903 ( \28899 , \28893 , \28898 );
buf \U$28904 ( \28900 , \28899 );
buf \U$28905 ( \28901 , \28900 );
nand \U$28906 ( \28902 , \28892 , \28901 );
buf \U$28907 ( \28903 , \28902 );
buf \U$28908 ( \28904 , \28903 );
buf \U$28909 ( \28905 , \28209 );
not \U$28910 ( \28906 , \28905 );
buf \U$28911 ( \28907 , \14608 );
not \U$28912 ( \28908 , \28907 );
or \U$28913 ( \28909 , \28906 , \28908 );
buf \U$28914 ( \28910 , \791 );
buf \U$28915 ( \28911 , RIc0d89b0_42);
buf \U$28916 ( \28912 , RIc0d9838_73);
xor \U$28917 ( \28913 , \28911 , \28912 );
buf \U$28918 ( \28914 , \28913 );
buf \U$28919 ( \28915 , \28914 );
nand \U$28920 ( \28916 , \28910 , \28915 );
buf \U$28921 ( \28917 , \28916 );
buf \U$28922 ( \28918 , \28917 );
nand \U$28923 ( \28919 , \28909 , \28918 );
buf \U$28924 ( \28920 , \28919 );
buf \U$28925 ( \28921 , \28920 );
xor \U$28926 ( \28922 , \28904 , \28921 );
buf \U$28927 ( \28923 , RIc0da738_105);
buf \U$28928 ( \28924 , RIc0d7b28_11);
xor \U$28929 ( \28925 , \28923 , \28924 );
buf \U$28930 ( \28926 , \28925 );
buf \U$28931 ( \28927 , \28926 );
not \U$28932 ( \28928 , \28927 );
buf \U$28933 ( \28929 , \15644 );
not \U$28934 ( \28930 , \28929 );
or \U$28935 ( \28931 , \28928 , \28930 );
buf \U$28936 ( \28932 , \15653 );
buf \U$28937 ( \28933 , RIc0da738_105);
buf \U$28938 ( \28934 , RIc0d7ab0_10);
xor \U$28939 ( \28935 , \28933 , \28934 );
buf \U$28940 ( \28936 , \28935 );
buf \U$28941 ( \28937 , \28936 );
nand \U$28942 ( \28938 , \28932 , \28937 );
buf \U$28943 ( \28939 , \28938 );
buf \U$28944 ( \28940 , \28939 );
nand \U$28945 ( \28941 , \28931 , \28940 );
buf \U$28946 ( \28942 , \28941 );
buf \U$28947 ( \28943 , \28942 );
xor \U$28948 ( \28944 , \28922 , \28943 );
buf \U$28949 ( \28945 , \28944 );
buf \U$28950 ( \28946 , \28945 );
not \U$28951 ( \28947 , \28946 );
buf \U$28952 ( \28948 , \28488 );
not \U$28953 ( \28949 , \28948 );
buf \U$28954 ( \28950 , \436 );
not \U$28955 ( \28951 , \28950 );
or \U$28956 ( \28952 , \28949 , \28951 );
buf \U$28957 ( \28953 , \846 );
xor \U$28958 ( \28954 , RIc0d9fb8_89, RIc0d8230_26);
buf \U$28959 ( \28955 , \28954 );
nand \U$28960 ( \28956 , \28953 , \28955 );
buf \U$28961 ( \28957 , \28956 );
buf \U$28962 ( \28958 , \28957 );
nand \U$28963 ( \28959 , \28952 , \28958 );
buf \U$28964 ( \28960 , \28959 );
buf \U$28965 ( \28961 , \28121 );
not \U$28966 ( \28962 , \28961 );
buf \U$28967 ( \28963 , \3780 );
not \U$28968 ( \28964 , \28963 );
or \U$28969 ( \28965 , \28962 , \28964 );
buf \U$28970 ( \28966 , \1229 );
buf \U$28971 ( \28967 , RIc0d9478_65);
buf \U$28972 ( \28968 , RIc0d8d70_50);
xor \U$28973 ( \28969 , \28967 , \28968 );
buf \U$28974 ( \28970 , \28969 );
buf \U$28975 ( \28971 , \28970 );
nand \U$28976 ( \28972 , \28966 , \28971 );
buf \U$28977 ( \28973 , \28972 );
buf \U$28978 ( \28974 , \28973 );
nand \U$28979 ( \28975 , \28965 , \28974 );
buf \U$28980 ( \28976 , \28975 );
xor \U$28981 ( \28977 , \28960 , \28976 );
buf \U$28982 ( \28978 , \28314 );
not \U$28983 ( \28979 , \28978 );
buf \U$28984 ( \28980 , \1351 );
not \U$28985 ( \28981 , \28980 );
or \U$28986 ( \28982 , \28979 , \28981 );
buf \U$28987 ( \28983 , \1025 );
buf \U$28988 ( \28984 , RIc0d86e0_36);
buf \U$28989 ( \28985 , RIc0d9b08_79);
xor \U$28990 ( \28986 , \28984 , \28985 );
buf \U$28991 ( \28987 , \28986 );
buf \U$28992 ( \28988 , \28987 );
nand \U$28993 ( \28989 , \28983 , \28988 );
buf \U$28994 ( \28990 , \28989 );
buf \U$28995 ( \28991 , \28990 );
nand \U$28996 ( \28992 , \28982 , \28991 );
buf \U$28997 ( \28993 , \28992 );
xnor \U$28998 ( \28994 , \28977 , \28993 );
buf \U$28999 ( \28995 , \28994 );
not \U$29000 ( \28996 , \28995 );
buf \U$29001 ( \28997 , \28996 );
buf \U$29002 ( \28998 , \28997 );
not \U$29003 ( \28999 , \28998 );
or \U$29004 ( \29000 , \28947 , \28999 );
buf \U$29005 ( \29001 , \28945 );
not \U$29006 ( \29002 , \29001 );
buf \U$29007 ( \29003 , \29002 );
buf \U$29008 ( \29004 , \29003 );
not \U$29009 ( \29005 , \29004 );
buf \U$29010 ( \29006 , \28994 );
not \U$29011 ( \29007 , \29006 );
or \U$29012 ( \29008 , \29005 , \29007 );
buf \U$29013 ( \29009 , \28072 );
not \U$29014 ( \29010 , \29009 );
buf \U$29015 ( \29011 , \4691 );
not \U$29016 ( \29012 , \29011 );
or \U$29017 ( \29013 , \29010 , \29012 );
buf \U$29018 ( \29014 , \284 );
buf \U$29019 ( \29015 , RIc0d8b90_46);
buf \U$29020 ( \29016 , RIc0d9658_69);
xor \U$29021 ( \29017 , \29015 , \29016 );
buf \U$29022 ( \29018 , \29017 );
buf \U$29023 ( \29019 , \29018 );
nand \U$29024 ( \29020 , \29014 , \29019 );
buf \U$29025 ( \29021 , \29020 );
buf \U$29026 ( \29022 , \29021 );
nand \U$29027 ( \29023 , \29013 , \29022 );
buf \U$29028 ( \29024 , \29023 );
buf \U$29029 ( \29025 , \28361 );
not \U$29030 ( \29026 , \29025 );
buf \U$29031 ( \29027 , \17141 );
not \U$29032 ( \29028 , \29027 );
or \U$29033 ( \29029 , \29026 , \29028 );
buf \U$29034 ( \29030 , \1078 );
xor \U$29035 ( \29031 , RIc0d9bf8_81, RIc0d85f0_34);
buf \U$29036 ( \29032 , \29031 );
nand \U$29037 ( \29033 , \29030 , \29032 );
buf \U$29038 ( \29034 , \29033 );
buf \U$29039 ( \29035 , \29034 );
nand \U$29040 ( \29036 , \29029 , \29035 );
buf \U$29041 ( \29037 , \29036 );
xor \U$29042 ( \29038 , \29024 , \29037 );
buf \U$29043 ( \29039 , \28399 );
not \U$29044 ( \29040 , \29039 );
buf \U$29045 ( \29041 , \1183 );
not \U$29046 ( \29042 , \29041 );
or \U$29047 ( \29043 , \29040 , \29042 );
buf \U$29048 ( \29044 , \3742 );
buf \U$29049 ( \29045 , RIc0d9a18_77);
buf \U$29050 ( \29046 , RIc0d87d0_38);
xor \U$29051 ( \29047 , \29045 , \29046 );
buf \U$29052 ( \29048 , \29047 );
buf \U$29053 ( \29049 , \29048 );
nand \U$29054 ( \29050 , \29044 , \29049 );
buf \U$29055 ( \29051 , \29050 );
buf \U$29056 ( \29052 , \29051 );
nand \U$29057 ( \29053 , \29043 , \29052 );
buf \U$29058 ( \29054 , \29053 );
xnor \U$29059 ( \29055 , \29038 , \29054 );
not \U$29060 ( \29056 , \29055 );
buf \U$29061 ( \29057 , \29056 );
nand \U$29062 ( \29058 , \29008 , \29057 );
buf \U$29063 ( \29059 , \29058 );
buf \U$29064 ( \29060 , \29059 );
nand \U$29065 ( \29061 , \29000 , \29060 );
buf \U$29066 ( \29062 , \29061 );
xor \U$29067 ( \29063 , \28887 , \29062 );
buf \U$29068 ( \29064 , \29063 );
buf \U$29069 ( \29065 , \28164 );
not \U$29070 ( \29066 , \29065 );
buf \U$29071 ( \29067 , \2938 );
not \U$29072 ( \29068 , \29067 );
buf \U$29073 ( \29069 , \29068 );
buf \U$29074 ( \29070 , \29069 );
not \U$29075 ( \29071 , \29070 );
or \U$29076 ( \29072 , \29066 , \29071 );
buf \U$29077 ( \29073 , \2070 );
xor \U$29078 ( \29074 , RIc0da378_97, RIc0d7e70_18);
buf \U$29079 ( \29075 , \29074 );
nand \U$29080 ( \29076 , \29073 , \29075 );
buf \U$29081 ( \29077 , \29076 );
buf \U$29082 ( \29078 , \29077 );
nand \U$29083 ( \29079 , \29072 , \29078 );
buf \U$29084 ( \29080 , \29079 );
buf \U$29085 ( \29081 , \29080 );
not \U$29086 ( \29082 , \29081 );
buf \U$29087 ( \29083 , \29082 );
buf \U$29088 ( \29084 , \29083 );
not \U$29089 ( \29085 , \29084 );
buf \U$29090 ( \29086 , \28292 );
not \U$29091 ( \29087 , \29086 );
buf \U$29092 ( \29088 , \20759 );
not \U$29093 ( \29089 , \29088 );
or \U$29094 ( \29090 , \29087 , \29089 );
buf \U$29095 ( \29091 , \13426 );
xor \U$29096 ( \29092 , RIc0da918_109, RIc0d78d0_6);
buf \U$29097 ( \29093 , \29092 );
nand \U$29098 ( \29094 , \29091 , \29093 );
buf \U$29099 ( \29095 , \29094 );
buf \U$29100 ( \29096 , \29095 );
nand \U$29101 ( \29097 , \29090 , \29096 );
buf \U$29102 ( \29098 , \29097 );
buf \U$29103 ( \29099 , \29098 );
not \U$29104 ( \29100 , \29099 );
buf \U$29105 ( \29101 , \29100 );
buf \U$29106 ( \29102 , \29101 );
not \U$29107 ( \29103 , \29102 );
or \U$29108 ( \29104 , \29085 , \29103 );
buf \U$29109 ( \29105 , \28055 );
not \U$29110 ( \29106 , \29105 );
buf \U$29111 ( \29107 , \1736 );
not \U$29112 ( \29108 , \29107 );
or \U$29113 ( \29109 , \29106 , \29108 );
buf \U$29114 ( \29110 , \584 );
buf \U$29115 ( \29111 , RIc0d9ce8_83);
buf \U$29116 ( \29112 , RIc0d8500_32);
xor \U$29117 ( \29113 , \29111 , \29112 );
buf \U$29118 ( \29114 , \29113 );
buf \U$29119 ( \29115 , \29114 );
nand \U$29120 ( \29116 , \29110 , \29115 );
buf \U$29121 ( \29117 , \29116 );
buf \U$29122 ( \29118 , \29117 );
nand \U$29123 ( \29119 , \29109 , \29118 );
buf \U$29124 ( \29120 , \29119 );
buf \U$29125 ( \29121 , \29120 );
nand \U$29126 ( \29122 , \29104 , \29121 );
buf \U$29127 ( \29123 , \29122 );
buf \U$29128 ( \29124 , \29123 );
buf \U$29129 ( \29125 , \29098 );
buf \U$29130 ( \29126 , \29080 );
nand \U$29131 ( \29127 , \29125 , \29126 );
buf \U$29132 ( \29128 , \29127 );
buf \U$29133 ( \29129 , \29128 );
nand \U$29134 ( \29130 , \29124 , \29129 );
buf \U$29135 ( \29131 , \29130 );
buf \U$29136 ( \29132 , \28739 );
not \U$29137 ( \29133 , \29132 );
buf \U$29138 ( \29134 , \28715 );
not \U$29139 ( \29135 , \29134 );
or \U$29140 ( \29136 , \29133 , \29135 );
buf \U$29141 ( \29137 , \28742 );
not \U$29142 ( \29138 , \29137 );
buf \U$29143 ( \29139 , \28721 );
not \U$29144 ( \29140 , \29139 );
or \U$29145 ( \29141 , \29138 , \29140 );
buf \U$29146 ( \29142 , \28698 );
nand \U$29147 ( \29143 , \29141 , \29142 );
buf \U$29148 ( \29144 , \29143 );
buf \U$29149 ( \29145 , \29144 );
nand \U$29150 ( \29146 , \29136 , \29145 );
buf \U$29151 ( \29147 , \29146 );
xor \U$29152 ( \29148 , \29131 , \29147 );
buf \U$29153 ( \29149 , \28787 );
buf \U$29154 ( \29150 , \28770 );
nor \U$29155 ( \29151 , \29149 , \29150 );
buf \U$29156 ( \29152 , \29151 );
buf \U$29157 ( \29153 , \29152 );
buf \U$29158 ( \29154 , \28811 );
or \U$29159 ( \29155 , \29153 , \29154 );
buf \U$29160 ( \29156 , \28787 );
buf \U$29161 ( \29157 , \28770 );
nand \U$29162 ( \29158 , \29156 , \29157 );
buf \U$29163 ( \29159 , \29158 );
buf \U$29164 ( \29160 , \29159 );
nand \U$29165 ( \29161 , \29155 , \29160 );
buf \U$29166 ( \29162 , \29161 );
xor \U$29167 ( \29163 , \29148 , \29162 );
buf \U$29168 ( \29164 , \29163 );
and \U$29169 ( \29165 , \29064 , \29164 );
not \U$29170 ( \29166 , \29064 );
buf \U$29171 ( \29167 , \29163 );
not \U$29172 ( \29168 , \29167 );
buf \U$29173 ( \29169 , \29168 );
buf \U$29174 ( \29170 , \29169 );
and \U$29175 ( \29171 , \29166 , \29170 );
nor \U$29176 ( \29172 , \29165 , \29171 );
buf \U$29177 ( \29173 , \29172 );
buf \U$29178 ( \29174 , \29173 );
xor \U$29179 ( \29175 , \28685 , \29174 );
buf \U$29180 ( \29176 , \29175 );
buf \U$29181 ( \29177 , \29176 );
xor \U$29182 ( \29178 , \28666 , \28545 );
and \U$29183 ( \29179 , \29178 , \28630 );
not \U$29184 ( \29180 , \29178 );
and \U$29185 ( \29181 , \29180 , \28676 );
nor \U$29186 ( \29182 , \29179 , \29181 );
buf \U$29187 ( \29183 , \29182 );
xor \U$29188 ( \29184 , \28173 , \28253 );
xnor \U$29189 ( \29185 , \29184 , \28106 );
buf \U$29190 ( \29186 , \29185 );
xor \U$29191 ( \29187 , \28324 , \28371 );
xor \U$29192 ( \29188 , \29187 , \28431 );
buf \U$29193 ( \29189 , \29188 );
buf \U$29194 ( \29190 , \29189 );
xor \U$29195 ( \29191 , \29186 , \29190 );
buf \U$29196 ( \29192 , \13953 );
buf \U$29197 ( \29193 , \23985 );
or \U$29198 ( \29194 , \29192 , \29193 );
buf \U$29199 ( \29195 , RIc0dadc8_119);
nand \U$29200 ( \29196 , \29194 , \29195 );
buf \U$29201 ( \29197 , \29196 );
buf \U$29202 ( \29198 , \29197 );
buf \U$29203 ( \29199 , \27547 );
not \U$29204 ( \29200 , \29199 );
buf \U$29205 ( \29201 , \25542 );
not \U$29206 ( \29202 , \29201 );
or \U$29207 ( \29203 , \29200 , \29202 );
buf \U$29208 ( \29204 , \13953 );
buf \U$29209 ( \29205 , RIc0dadc8_119);
nand \U$29210 ( \29206 , \29204 , \29205 );
buf \U$29211 ( \29207 , \29206 );
buf \U$29212 ( \29208 , \29207 );
nand \U$29213 ( \29209 , \29203 , \29208 );
buf \U$29214 ( \29210 , \29209 );
buf \U$29215 ( \29211 , \29210 );
nand \U$29216 ( \29212 , \29198 , \29211 );
buf \U$29217 ( \29213 , \29212 );
buf \U$29218 ( \29214 , \29213 );
buf \U$29219 ( \29215 , \29197 );
buf \U$29220 ( \29216 , \29210 );
or \U$29221 ( \29217 , \29215 , \29216 );
buf \U$29222 ( \29218 , RIc0da738_105);
buf \U$29223 ( \29219 , RIc0d7c90_14);
xor \U$29224 ( \29220 , \29218 , \29219 );
buf \U$29225 ( \29221 , \29220 );
buf \U$29226 ( \29222 , \29221 );
not \U$29227 ( \29223 , \29222 );
buf \U$29228 ( \29224 , \12736 );
not \U$29229 ( \29225 , \29224 );
or \U$29230 ( \29226 , \29223 , \29225 );
buf \U$29231 ( \29227 , \21880 );
buf \U$29232 ( \29228 , \27944 );
nand \U$29233 ( \29229 , \29227 , \29228 );
buf \U$29234 ( \29230 , \29229 );
buf \U$29235 ( \29231 , \29230 );
nand \U$29236 ( \29232 , \29226 , \29231 );
buf \U$29237 ( \29233 , \29232 );
buf \U$29238 ( \29234 , \29233 );
nand \U$29239 ( \29235 , \29217 , \29234 );
buf \U$29240 ( \29236 , \29235 );
buf \U$29241 ( \29237 , \29236 );
nand \U$29242 ( \29238 , \29214 , \29237 );
buf \U$29243 ( \29239 , \29238 );
buf \U$29244 ( \29240 , \29239 );
xor \U$29245 ( \29241 , RIc0d9748_71, RIc0d8c08_47);
and \U$29246 ( \29242 , \2923 , \29241 );
and \U$29247 ( \29243 , \1282 , \28132 );
nor \U$29248 ( \29244 , \29242 , \29243 );
buf \U$29249 ( \29245 , \29244 );
buf \U$29251 ( \29246 , \29245 );
buf \U$29252 ( \29247 , \29246 );
not \U$29253 ( \29248 , \29247 );
buf \U$29254 ( \29249 , RIc0daa08_111);
buf \U$29255 ( \29250 , RIc0d7948_7);
xor \U$29256 ( \29251 , \29249 , \29250 );
buf \U$29257 ( \29252 , \29251 );
buf \U$29258 ( \29253 , \29252 );
not \U$29259 ( \29254 , \29253 );
buf \U$29260 ( \29255 , \14346 );
not \U$29261 ( \29256 , \29255 );
or \U$29262 ( \29257 , \29254 , \29256 );
buf \U$29263 ( \29258 , \14106 );
buf \U$29264 ( \29259 , \28581 );
nand \U$29265 ( \29260 , \29258 , \29259 );
buf \U$29266 ( \29261 , \29260 );
buf \U$29267 ( \29262 , \29261 );
nand \U$29268 ( \29263 , \29257 , \29262 );
buf \U$29269 ( \29264 , \29263 );
buf \U$29270 ( \29265 , \29264 );
not \U$29271 ( \29266 , \29265 );
buf \U$29272 ( \29267 , \29266 );
buf \U$29273 ( \29268 , \29267 );
buf \U$29274 ( \29269 , RIc0da468_99);
buf \U$29275 ( \29270 , RIc0d7ee8_19);
xor \U$29276 ( \29271 , \29269 , \29270 );
buf \U$29277 ( \29272 , \29271 );
buf \U$29278 ( \29273 , \29272 );
not \U$29279 ( \29274 , \29273 );
buf \U$29280 ( \29275 , \16744 );
not \U$29281 ( \29276 , \29275 );
or \U$29282 ( \29277 , \29274 , \29276 );
buf \U$29283 ( \29278 , \16750 );
buf \U$29284 ( \29279 , \28604 );
nand \U$29285 ( \29280 , \29278 , \29279 );
buf \U$29286 ( \29281 , \29280 );
buf \U$29287 ( \29282 , \29281 );
nand \U$29288 ( \29283 , \29277 , \29282 );
buf \U$29289 ( \29284 , \29283 );
buf \U$29290 ( \29285 , \29284 );
xnor \U$29291 ( \29286 , \29268 , \29285 );
buf \U$29292 ( \29287 , \29286 );
buf \U$29293 ( \29288 , \29287 );
not \U$29294 ( \29289 , \29288 );
or \U$29295 ( \29290 , \29248 , \29289 );
buf \U$29296 ( \29291 , \29287 );
buf \U$29297 ( \29292 , \29246 );
or \U$29298 ( \29293 , \29291 , \29292 );
nand \U$29299 ( \29294 , \29290 , \29293 );
buf \U$29300 ( \29295 , \29294 );
buf \U$29301 ( \29296 , \29295 );
xor \U$29302 ( \29297 , \29240 , \29296 );
buf \U$29303 ( \29298 , \12361 );
buf \U$29304 ( \29299 , \27648 );
and \U$29305 ( \29300 , \29298 , \29299 );
buf \U$29306 ( \29301 , \402 );
xor \U$29307 ( \29302 , RIc0d9b08_79, RIc0d88c0_40);
buf \U$29308 ( \29303 , \29302 );
and \U$29309 ( \29304 , \29301 , \29303 );
nor \U$29310 ( \29305 , \29300 , \29304 );
buf \U$29311 ( \29306 , \29305 );
buf \U$29312 ( \29307 , \29306 );
not \U$29313 ( \29308 , \29307 );
buf \U$29314 ( \29309 , \29308 );
buf \U$29315 ( \29310 , \29309 );
not \U$29316 ( \29311 , \29310 );
buf \U$29317 ( \29312 , \27398 );
not \U$29318 ( \29313 , \29312 );
buf \U$29319 ( \29314 , \23253 );
not \U$29320 ( \29315 , \29314 );
or \U$29321 ( \29316 , \29313 , \29315 );
buf \U$29322 ( \29317 , \1229 );
buf \U$29323 ( \29318 , RIc0d9478_65);
buf \U$29324 ( \29319 , RIc0d8f50_54);
xor \U$29325 ( \29320 , \29318 , \29319 );
buf \U$29326 ( \29321 , \29320 );
buf \U$29327 ( \29322 , \29321 );
nand \U$29328 ( \29323 , \29317 , \29322 );
buf \U$29329 ( \29324 , \29323 );
buf \U$29330 ( \29325 , \29324 );
nand \U$29331 ( \29326 , \29316 , \29325 );
buf \U$29332 ( \29327 , \29326 );
buf \U$29333 ( \29328 , \29327 );
not \U$29334 ( \29329 , \29328 );
or \U$29335 ( \29330 , \29311 , \29329 );
buf \U$29336 ( \29331 , \29327 );
not \U$29337 ( \29332 , \29331 );
buf \U$29338 ( \29333 , \29306 );
nand \U$29339 ( \29334 , \29332 , \29333 );
buf \U$29340 ( \29335 , \29334 );
buf \U$29341 ( \29336 , \29335 );
buf \U$29342 ( \29337 , \27665 );
not \U$29343 ( \29338 , \29337 );
buf \U$29344 ( \29339 , \14210 );
not \U$29345 ( \29340 , \29339 );
or \U$29346 ( \29341 , \29338 , \29340 );
buf \U$29347 ( \29342 , \20211 );
buf \U$29348 ( \29343 , RIc0d7ab0_10);
buf \U$29349 ( \29344 , RIc0da918_109);
xor \U$29350 ( \29345 , \29343 , \29344 );
buf \U$29351 ( \29346 , \29345 );
buf \U$29352 ( \29347 , \29346 );
nand \U$29353 ( \29348 , \29342 , \29347 );
buf \U$29354 ( \29349 , \29348 );
buf \U$29355 ( \29350 , \29349 );
nand \U$29356 ( \29351 , \29341 , \29350 );
buf \U$29357 ( \29352 , \29351 );
buf \U$29358 ( \29353 , \29352 );
nand \U$29359 ( \29354 , \29336 , \29353 );
buf \U$29360 ( \29355 , \29354 );
buf \U$29361 ( \29356 , \29355 );
nand \U$29362 ( \29357 , \29330 , \29356 );
buf \U$29363 ( \29358 , \29357 );
buf \U$29364 ( \29359 , \29358 );
buf \U$29365 ( \29360 , \27415 );
not \U$29366 ( \29361 , \29360 );
buf \U$29367 ( \29362 , \1263 );
not \U$29368 ( \29363 , \29362 );
or \U$29369 ( \29364 , \29361 , \29363 );
buf \U$29370 ( \29365 , \1282 );
xor \U$29371 ( \29366 , RIc0d9748_71, RIc0d8c80_48);
buf \U$29372 ( \29367 , \29366 );
nand \U$29373 ( \29368 , \29365 , \29367 );
buf \U$29374 ( \29369 , \29368 );
buf \U$29375 ( \29370 , \29369 );
nand \U$29376 ( \29371 , \29364 , \29370 );
buf \U$29377 ( \29372 , \29371 );
not \U$29378 ( \29373 , \29372 );
buf \U$29379 ( \29374 , \27290 );
not \U$29380 ( \29375 , \29374 );
buf \U$29381 ( \29376 , \14346 );
not \U$29382 ( \29377 , \29376 );
or \U$29383 ( \29378 , \29375 , \29377 );
buf \U$29384 ( \29379 , \15864 );
buf \U$29385 ( \29380 , RIc0d79c0_8);
buf \U$29386 ( \29381 , RIc0daa08_111);
xor \U$29387 ( \29382 , \29380 , \29381 );
buf \U$29388 ( \29383 , \29382 );
buf \U$29389 ( \29384 , \29383 );
nand \U$29390 ( \29385 , \29379 , \29384 );
buf \U$29391 ( \29386 , \29385 );
buf \U$29392 ( \29387 , \29386 );
nand \U$29393 ( \29388 , \29378 , \29387 );
buf \U$29394 ( \29389 , \29388 );
buf \U$29395 ( \29390 , \29389 );
not \U$29396 ( \29391 , \29390 );
buf \U$29397 ( \29392 , \29391 );
nand \U$29398 ( \29393 , \29373 , \29392 );
not \U$29399 ( \29394 , \29393 );
buf \U$29400 ( \29395 , \27319 );
not \U$29401 ( \29396 , \29395 );
buf \U$29402 ( \29397 , \25371 );
not \U$29403 ( \29398 , \29397 );
or \U$29404 ( \29399 , \29396 , \29398 );
buf \U$29405 ( \29400 , \16750 );
buf \U$29406 ( \29401 , RIc0da468_99);
buf \U$29407 ( \29402 , RIc0d7f60_20);
xor \U$29408 ( \29403 , \29401 , \29402 );
buf \U$29409 ( \29404 , \29403 );
buf \U$29410 ( \29405 , \29404 );
nand \U$29411 ( \29406 , \29400 , \29405 );
buf \U$29412 ( \29407 , \29406 );
buf \U$29413 ( \29408 , \29407 );
nand \U$29414 ( \29409 , \29399 , \29408 );
buf \U$29415 ( \29410 , \29409 );
not \U$29416 ( \29411 , \29410 );
or \U$29417 ( \29412 , \29394 , \29411 );
buf \U$29418 ( \29413 , \29389 );
buf \U$29419 ( \29414 , \29372 );
nand \U$29420 ( \29415 , \29413 , \29414 );
buf \U$29421 ( \29416 , \29415 );
nand \U$29422 ( \29417 , \29412 , \29416 );
buf \U$29423 ( \29418 , \29417 );
xor \U$29424 ( \29419 , \29359 , \29418 );
buf \U$29425 ( \29420 , \27304 );
not \U$29426 ( \29421 , \29420 );
buf \U$29427 ( \29422 , \2399 );
not \U$29428 ( \29423 , \29422 );
or \U$29429 ( \29424 , \29421 , \29423 );
buf \U$29430 ( \29425 , \921 );
xor \U$29431 ( \29426 , RIc0d9dd8_85, RIc0d85f0_34);
buf \U$29432 ( \29427 , \29426 );
nand \U$29433 ( \29428 , \29425 , \29427 );
buf \U$29434 ( \29429 , \29428 );
buf \U$29435 ( \29430 , \29429 );
nand \U$29436 ( \29431 , \29424 , \29430 );
buf \U$29437 ( \29432 , \29431 );
buf \U$29438 ( \29433 , \29432 );
not \U$29439 ( \29434 , \29433 );
buf \U$29440 ( \29435 , \27251 );
not \U$29441 ( \29436 , \29435 );
buf \U$29442 ( \29437 , \25355 );
not \U$29443 ( \29438 , \29437 );
or \U$29444 ( \29439 , \29436 , \29438 );
buf \U$29445 ( \29440 , \16995 );
buf \U$29446 ( \29441 , RIc0d78d0_6);
buf \U$29447 ( \29442 , RIc0daaf8_113);
xor \U$29448 ( \29443 , \29441 , \29442 );
buf \U$29449 ( \29444 , \29443 );
buf \U$29450 ( \29445 , \29444 );
nand \U$29451 ( \29446 , \29440 , \29445 );
buf \U$29452 ( \29447 , \29446 );
buf \U$29453 ( \29448 , \29447 );
nand \U$29454 ( \29449 , \29439 , \29448 );
buf \U$29455 ( \29450 , \29449 );
buf \U$29456 ( \29451 , \29450 );
not \U$29457 ( \29452 , \29451 );
or \U$29458 ( \29453 , \29434 , \29452 );
buf \U$29459 ( \29454 , \29450 );
buf \U$29460 ( \29455 , \29432 );
or \U$29461 ( \29456 , \29454 , \29455 );
buf \U$29462 ( \29457 , \27715 );
not \U$29463 ( \29458 , \29457 );
buf \U$29464 ( \29459 , \4043 );
not \U$29465 ( \29460 , \29459 );
or \U$29466 ( \29461 , \29458 , \29460 );
buf \U$29467 ( \29462 , \4049 );
buf \U$29468 ( \29463 , RIc0d7e70_18);
buf \U$29469 ( \29464 , RIc0da558_101);
xor \U$29470 ( \29465 , \29463 , \29464 );
buf \U$29471 ( \29466 , \29465 );
buf \U$29472 ( \29467 , \29466 );
nand \U$29473 ( \29468 , \29462 , \29467 );
buf \U$29474 ( \29469 , \29468 );
buf \U$29475 ( \29470 , \29469 );
nand \U$29476 ( \29471 , \29461 , \29470 );
buf \U$29477 ( \29472 , \29471 );
buf \U$29478 ( \29473 , \29472 );
nand \U$29479 ( \29474 , \29456 , \29473 );
buf \U$29480 ( \29475 , \29474 );
buf \U$29481 ( \29476 , \29475 );
nand \U$29482 ( \29477 , \29453 , \29476 );
buf \U$29483 ( \29478 , \29477 );
buf \U$29484 ( \29479 , \29478 );
and \U$29485 ( \29480 , \29419 , \29479 );
and \U$29486 ( \29481 , \29359 , \29418 );
or \U$29487 ( \29482 , \29480 , \29481 );
buf \U$29488 ( \29483 , \29482 );
buf \U$29489 ( \29484 , \29483 );
and \U$29490 ( \29485 , \29297 , \29484 );
and \U$29491 ( \29486 , \29240 , \29296 );
or \U$29492 ( \29487 , \29485 , \29486 );
buf \U$29493 ( \29488 , \29487 );
buf \U$29494 ( \29489 , \29488 );
and \U$29495 ( \29490 , \29191 , \29489 );
and \U$29496 ( \29491 , \29186 , \29190 );
or \U$29497 ( \29492 , \29490 , \29491 );
buf \U$29498 ( \29493 , \29492 );
buf \U$29499 ( \29494 , \29493 );
xor \U$29500 ( \29495 , \29183 , \29494 );
buf \U$29501 ( \29496 , \29003 );
not \U$29502 ( \29497 , \29496 );
not \U$29503 ( \29498 , \29055 );
buf \U$29504 ( \29499 , \29498 );
not \U$29505 ( \29500 , \29499 );
or \U$29506 ( \29501 , \29497 , \29500 );
buf \U$29507 ( \29502 , \29055 );
buf \U$29508 ( \29503 , \28945 );
nand \U$29509 ( \29504 , \29502 , \29503 );
buf \U$29510 ( \29505 , \29504 );
buf \U$29511 ( \29506 , \29505 );
nand \U$29512 ( \29507 , \29501 , \29506 );
buf \U$29513 ( \29508 , \29507 );
buf \U$29514 ( \29509 , \29508 );
buf \U$29515 ( \29510 , \28997 );
and \U$29516 ( \29511 , \29509 , \29510 );
not \U$29517 ( \29512 , \29509 );
buf \U$29518 ( \29513 , \28994 );
and \U$29519 ( \29514 , \29512 , \29513 );
nor \U$29520 ( \29515 , \29511 , \29514 );
buf \U$29521 ( \29516 , \29515 );
buf \U$29522 ( \29517 , \29516 );
and \U$29523 ( \29518 , \28108 , \28109 );
buf \U$29524 ( \29519 , \29518 );
buf \U$29525 ( \29520 , \29519 );
buf \U$29526 ( \29521 , \28237 );
not \U$29527 ( \29522 , \29521 );
buf \U$29528 ( \29523 , \2607 );
not \U$29529 ( \29524 , \29523 );
or \U$29530 ( \29525 , \29522 , \29524 );
buf \U$29531 ( \29526 , \14331 );
buf \U$29532 ( \29527 , RIc0d9ec8_87);
buf \U$29533 ( \29528 , RIc0d8320_28);
xor \U$29534 ( \29529 , \29527 , \29528 );
buf \U$29535 ( \29530 , \29529 );
buf \U$29536 ( \29531 , \29530 );
nand \U$29537 ( \29532 , \29526 , \29531 );
buf \U$29538 ( \29533 , \29532 );
buf \U$29539 ( \29534 , \29533 );
nand \U$29540 ( \29535 , \29525 , \29534 );
buf \U$29541 ( \29536 , \29535 );
buf \U$29542 ( \29537 , \29536 );
not \U$29543 ( \29538 , \29537 );
buf \U$29544 ( \29539 , \29538 );
buf \U$29545 ( \29540 , \29539 );
xor \U$29546 ( \29541 , \29520 , \29540 );
buf \U$29547 ( \29542 , \28531 );
not \U$29548 ( \29543 , \29542 );
buf \U$29549 ( \29544 , \4483 );
not \U$29550 ( \29545 , \29544 );
buf \U$29551 ( \29546 , \29545 );
buf \U$29552 ( \29547 , \29546 );
not \U$29553 ( \29548 , \29547 );
or \U$29554 ( \29549 , \29543 , \29548 );
buf \U$29555 ( \29550 , \13712 );
buf \U$29556 ( \29551 , RIc0da648_103);
buf \U$29557 ( \29552 , RIc0d7ba0_12);
xor \U$29558 ( \29553 , \29551 , \29552 );
buf \U$29559 ( \29554 , \29553 );
buf \U$29560 ( \29555 , \29554 );
nand \U$29561 ( \29556 , \29550 , \29555 );
buf \U$29562 ( \29557 , \29556 );
buf \U$29563 ( \29558 , \29557 );
nand \U$29564 ( \29559 , \29549 , \29558 );
buf \U$29565 ( \29560 , \29559 );
buf \U$29566 ( \29561 , \29560 );
xor \U$29567 ( \29562 , \29541 , \29561 );
buf \U$29568 ( \29563 , \29562 );
buf \U$29569 ( \29564 , \29563 );
not \U$29570 ( \29565 , \29080 );
not \U$29571 ( \29566 , \29101 );
or \U$29572 ( \29567 , \29565 , \29566 );
buf \U$29573 ( \29568 , \29098 );
buf \U$29574 ( \29569 , \29083 );
nand \U$29575 ( \29570 , \29568 , \29569 );
buf \U$29576 ( \29571 , \29570 );
nand \U$29577 ( \29572 , \29567 , \29571 );
xor \U$29578 ( \29573 , \29572 , \29120 );
buf \U$29579 ( \29574 , \29573 );
xor \U$29580 ( \29575 , \29564 , \29574 );
buf \U$29581 ( \29576 , \28189 );
not \U$29582 ( \29577 , \29576 );
buf \U$29583 ( \29578 , \12833 );
not \U$29584 ( \29579 , \29578 );
or \U$29585 ( \29580 , \29577 , \29579 );
buf \U$29586 ( \29581 , \16676 );
xor \U$29587 ( \29582 , RIc0da558_101, RIc0d7c90_14);
buf \U$29588 ( \29583 , \29582 );
nand \U$29589 ( \29584 , \29581 , \29583 );
buf \U$29590 ( \29585 , \29584 );
buf \U$29591 ( \29586 , \29585 );
nand \U$29592 ( \29587 , \29580 , \29586 );
buf \U$29593 ( \29588 , \29587 );
buf \U$29594 ( \29589 , \28334 );
not \U$29595 ( \29590 , \29589 );
buf \U$29596 ( \29591 , \14186 );
not \U$29597 ( \29592 , \29591 );
or \U$29598 ( \29593 , \29590 , \29592 );
buf \U$29599 ( \29594 , \12303 );
buf \U$29600 ( \29595 , RIc0dabe8_115);
nand \U$29601 ( \29596 , \29594 , \29595 );
buf \U$29602 ( \29597 , \29596 );
buf \U$29603 ( \29598 , \29597 );
nand \U$29604 ( \29599 , \29593 , \29598 );
buf \U$29605 ( \29600 , \29599 );
buf \U$29606 ( \29601 , \29600 );
not \U$29607 ( \29602 , \29601 );
buf \U$29608 ( \29603 , \29602 );
and \U$29609 ( \29604 , \29588 , \29603 );
not \U$29610 ( \29605 , \29588 );
and \U$29611 ( \29606 , \29605 , \29600 );
or \U$29612 ( \29607 , \29604 , \29606 );
buf \U$29613 ( \29608 , \29607 );
buf \U$29614 ( \29609 , \28506 );
not \U$29615 ( \29610 , \29609 );
buf \U$29616 ( \29611 , \3714 );
not \U$29617 ( \29612 , \29611 );
or \U$29618 ( \29613 , \29610 , \29612 );
buf \U$29619 ( \29614 , \344 );
buf \U$29620 ( \29615 , RIc0da288_95);
buf \U$29621 ( \29616 , RIc0d7f60_20);
xor \U$29622 ( \29617 , \29615 , \29616 );
buf \U$29623 ( \29618 , \29617 );
buf \U$29624 ( \29619 , \29618 );
nand \U$29625 ( \29620 , \29614 , \29619 );
buf \U$29626 ( \29621 , \29620 );
buf \U$29627 ( \29622 , \29621 );
nand \U$29628 ( \29623 , \29613 , \29622 );
buf \U$29629 ( \29624 , \29623 );
buf \U$29630 ( \29625 , \29624 );
xor \U$29631 ( \29626 , \29608 , \29625 );
buf \U$29632 ( \29627 , \29626 );
buf \U$29633 ( \29628 , \29627 );
xor \U$29634 ( \29629 , \29575 , \29628 );
buf \U$29635 ( \29630 , \29629 );
buf \U$29636 ( \29631 , \29630 );
xor \U$29637 ( \29632 , \29517 , \29631 );
xor \U$29638 ( \29633 , \28814 , \28881 );
and \U$29639 ( \29634 , \29633 , \28749 );
not \U$29640 ( \29635 , \29633 );
and \U$29641 ( \29636 , \29635 , \28752 );
nor \U$29642 ( \29637 , \29634 , \29636 );
buf \U$29643 ( \29638 , \29637 );
xor \U$29644 ( \29639 , \29632 , \29638 );
buf \U$29645 ( \29640 , \29639 );
buf \U$29646 ( \29641 , \29640 );
and \U$29647 ( \29642 , \29495 , \29641 );
and \U$29648 ( \29643 , \29183 , \29494 );
or \U$29649 ( \29644 , \29642 , \29643 );
buf \U$29650 ( \29645 , \29644 );
buf \U$29651 ( \29646 , \29645 );
xor \U$29652 ( \29647 , \29177 , \29646 );
buf \U$29653 ( \29648 , \28638 );
not \U$29654 ( \29649 , \29648 );
buf \U$29655 ( \29650 , \29649 );
buf \U$29656 ( \29651 , \29650 );
not \U$29657 ( \29652 , \29651 );
buf \U$29658 ( \29653 , \28646 );
not \U$29659 ( \29654 , \29653 );
or \U$29660 ( \29655 , \29652 , \29654 );
buf \U$29661 ( \29656 , \28656 );
nand \U$29662 ( \29657 , \29655 , \29656 );
buf \U$29663 ( \29658 , \29657 );
buf \U$29664 ( \29659 , \29658 );
buf \U$29665 ( \29660 , \29650 );
not \U$29666 ( \29661 , \29660 );
buf \U$29667 ( \29662 , \28643 );
nand \U$29668 ( \29663 , \29661 , \29662 );
buf \U$29669 ( \29664 , \29663 );
buf \U$29670 ( \29665 , \29664 );
nand \U$29671 ( \29666 , \29659 , \29665 );
buf \U$29672 ( \29667 , \29666 );
buf \U$29673 ( \29668 , \29667 );
not \U$29674 ( \29669 , \29668 );
buf \U$29675 ( \29670 , \29669 );
buf \U$29676 ( \29671 , \29670 );
not \U$29677 ( \29672 , \29671 );
buf \U$29678 ( \29673 , \29536 );
buf \U$29679 ( \29674 , \28976 );
not \U$29680 ( \29675 , \29674 );
buf \U$29681 ( \29676 , \28960 );
not \U$29682 ( \29677 , \29676 );
or \U$29683 ( \29678 , \29675 , \29677 );
buf \U$29684 ( \29679 , \28960 );
buf \U$29685 ( \29680 , \28976 );
or \U$29686 ( \29681 , \29679 , \29680 );
buf \U$29687 ( \29682 , \28993 );
nand \U$29688 ( \29683 , \29681 , \29682 );
buf \U$29689 ( \29684 , \29683 );
buf \U$29690 ( \29685 , \29684 );
nand \U$29691 ( \29686 , \29678 , \29685 );
buf \U$29692 ( \29687 , \29686 );
buf \U$29693 ( \29688 , \29687 );
xor \U$29694 ( \29689 , \29673 , \29688 );
xor \U$29695 ( \29690 , \28842 , \28860 );
and \U$29696 ( \29691 , \29690 , \28879 );
and \U$29697 ( \29692 , \28842 , \28860 );
or \U$29698 ( \29693 , \29691 , \29692 );
buf \U$29699 ( \29694 , \29693 );
buf \U$29700 ( \29695 , \29694 );
xnor \U$29701 ( \29696 , \29689 , \29695 );
buf \U$29702 ( \29697 , \29696 );
buf \U$29703 ( \29698 , \29697 );
not \U$29704 ( \29699 , \29698 );
buf \U$29705 ( \29700 , \29699 );
buf \U$29706 ( \29701 , \29700 );
not \U$29707 ( \29702 , \29701 );
or \U$29708 ( \29703 , \29672 , \29702 );
buf \U$29709 ( \29704 , \29697 );
buf \U$29710 ( \29705 , \29667 );
nand \U$29711 ( \29706 , \29704 , \29705 );
buf \U$29712 ( \29707 , \29706 );
buf \U$29713 ( \29708 , \29707 );
nand \U$29714 ( \29709 , \29703 , \29708 );
buf \U$29715 ( \29710 , \29709 );
buf \U$29716 ( \29711 , \29037 );
not \U$29717 ( \29712 , \29711 );
buf \U$29718 ( \29713 , \29024 );
not \U$29719 ( \29714 , \29713 );
or \U$29720 ( \29715 , \29712 , \29714 );
buf \U$29721 ( \29716 , \29037 );
buf \U$29722 ( \29717 , \29024 );
or \U$29723 ( \29718 , \29716 , \29717 );
buf \U$29724 ( \29719 , \29054 );
nand \U$29725 ( \29720 , \29718 , \29719 );
buf \U$29726 ( \29721 , \29720 );
buf \U$29727 ( \29722 , \29721 );
nand \U$29728 ( \29723 , \29715 , \29722 );
buf \U$29729 ( \29724 , \29723 );
buf \U$29730 ( \29725 , \29724 );
buf \U$29731 ( \29726 , \28903 );
buf \U$29732 ( \29727 , \28920 );
or \U$29733 ( \29728 , \29726 , \29727 );
buf \U$29734 ( \29729 , \28942 );
nand \U$29735 ( \29730 , \29728 , \29729 );
buf \U$29736 ( \29731 , \29730 );
buf \U$29737 ( \29732 , \29731 );
buf \U$29738 ( \29733 , \28920 );
buf \U$29739 ( \29734 , \28903 );
nand \U$29740 ( \29735 , \29733 , \29734 );
buf \U$29741 ( \29736 , \29735 );
buf \U$29742 ( \29737 , \29736 );
nand \U$29743 ( \29738 , \29732 , \29737 );
buf \U$29744 ( \29739 , \29738 );
buf \U$29745 ( \29740 , \29739 );
xor \U$29746 ( \29741 , \29725 , \29740 );
buf \U$29747 ( \29742 , \29624 );
buf \U$29748 ( \29743 , \29588 );
nor \U$29749 ( \29744 , \29742 , \29743 );
buf \U$29750 ( \29745 , \29744 );
buf \U$29751 ( \29746 , \29745 );
buf \U$29752 ( \29747 , \29603 );
or \U$29753 ( \29748 , \29746 , \29747 );
buf \U$29754 ( \29749 , \29624 );
buf \U$29755 ( \29750 , \29588 );
nand \U$29756 ( \29751 , \29749 , \29750 );
buf \U$29757 ( \29752 , \29751 );
buf \U$29758 ( \29753 , \29752 );
nand \U$29759 ( \29754 , \29748 , \29753 );
buf \U$29760 ( \29755 , \29754 );
buf \U$29761 ( \29756 , \29755 );
xnor \U$29762 ( \29757 , \29741 , \29756 );
buf \U$29763 ( \29758 , \29757 );
not \U$29764 ( \29759 , \29758 );
and \U$29765 ( \29760 , \29710 , \29759 );
not \U$29766 ( \29761 , \29710 );
and \U$29767 ( \29762 , \29761 , \29758 );
nor \U$29768 ( \29763 , \29760 , \29762 );
buf \U$29769 ( \29764 , \29763 );
xor \U$29770 ( \29765 , \29517 , \29631 );
and \U$29771 ( \29766 , \29765 , \29638 );
and \U$29772 ( \29767 , \29517 , \29631 );
or \U$29773 ( \29768 , \29766 , \29767 );
buf \U$29774 ( \29769 , \29768 );
buf \U$29775 ( \29770 , \29769 );
xor \U$29776 ( \29771 , \29764 , \29770 );
buf \U$29777 ( \29772 , \28802 );
not \U$29778 ( \29773 , \29772 );
buf \U$29779 ( \29774 , \12334 );
not \U$29780 ( \29775 , \29774 );
or \U$29781 ( \29776 , \29773 , \29775 );
buf \U$29782 ( \29777 , \16071 );
buf \U$29783 ( \29778 , RIc0da828_107);
buf \U$29784 ( \29779 , RIc0d7948_7);
xor \U$29785 ( \29780 , \29778 , \29779 );
buf \U$29786 ( \29781 , \29780 );
buf \U$29787 ( \29782 , \29781 );
nand \U$29788 ( \29783 , \29777 , \29782 );
buf \U$29789 ( \29784 , \29783 );
buf \U$29790 ( \29785 , \29784 );
nand \U$29791 ( \29786 , \29776 , \29785 );
buf \U$29792 ( \29787 , \29786 );
buf \U$29793 ( \29788 , \29114 );
not \U$29794 ( \29789 , \29788 );
buf \U$29795 ( \29790 , \573 );
not \U$29796 ( \29791 , \29790 );
or \U$29797 ( \29792 , \29789 , \29791 );
buf \U$29798 ( \29793 , \584 );
xor \U$29799 ( \29794 , RIc0d9ce8_83, RIc0d8488_31);
buf \U$29800 ( \29795 , \29794 );
nand \U$29801 ( \29796 , \29793 , \29795 );
buf \U$29802 ( \29797 , \29796 );
buf \U$29803 ( \29798 , \29797 );
nand \U$29804 ( \29799 , \29792 , \29798 );
buf \U$29805 ( \29800 , \29799 );
buf \U$29806 ( \29801 , \29800 );
not \U$29807 ( \29802 , \29801 );
buf \U$29808 ( \29803 , \29802 );
xor \U$29809 ( \29804 , \29787 , \29803 );
buf \U$29810 ( \29805 , \29018 );
not \U$29811 ( \29806 , \29805 );
buf \U$29812 ( \29807 , \864 );
not \U$29813 ( \29808 , \29807 );
or \U$29814 ( \29809 , \29806 , \29808 );
buf \U$29815 ( \29810 , \284 );
buf \U$29816 ( \29811 , RIc0d9658_69);
buf \U$29817 ( \29812 , RIc0d8b18_45);
xor \U$29818 ( \29813 , \29811 , \29812 );
buf \U$29819 ( \29814 , \29813 );
buf \U$29820 ( \29815 , \29814 );
nand \U$29821 ( \29816 , \29810 , \29815 );
buf \U$29822 ( \29817 , \29816 );
buf \U$29823 ( \29818 , \29817 );
nand \U$29824 ( \29819 , \29809 , \29818 );
buf \U$29825 ( \29820 , \29819 );
xor \U$29826 ( \29821 , \29804 , \29820 );
buf \U$29827 ( \29822 , \29821 );
not \U$29828 ( \29823 , \29822 );
buf \U$29829 ( \29824 , \29823 );
buf \U$29830 ( \29825 , \29824 );
not \U$29831 ( \29826 , \29825 );
buf \U$29832 ( \29827 , \28954 );
not \U$29833 ( \29828 , \29827 );
buf \U$29834 ( \29829 , \2037 );
not \U$29835 ( \29830 , \29829 );
or \U$29836 ( \29831 , \29828 , \29830 );
buf \U$29837 ( \29832 , \16477 );
buf \U$29838 ( \29833 , RIc0d9fb8_89);
buf \U$29839 ( \29834 , RIc0d81b8_25);
xor \U$29840 ( \29835 , \29833 , \29834 );
buf \U$29841 ( \29836 , \29835 );
buf \U$29842 ( \29837 , \29836 );
nand \U$29843 ( \29838 , \29832 , \29837 );
buf \U$29844 ( \29839 , \29838 );
buf \U$29845 ( \29840 , \29839 );
nand \U$29846 ( \29841 , \29831 , \29840 );
buf \U$29847 ( \29842 , \29841 );
buf \U$29848 ( \29843 , \29842 );
buf \U$29849 ( \29844 , \29031 );
not \U$29850 ( \29845 , \29844 );
buf \U$29851 ( \29846 , \14532 );
not \U$29852 ( \29847 , \29846 );
or \U$29853 ( \29848 , \29845 , \29847 );
buf \U$29854 ( \29849 , RIc0d9bf8_81);
buf \U$29855 ( \29850 , RIc0d8578_33);
xnor \U$29856 ( \29851 , \29849 , \29850 );
buf \U$29857 ( \29852 , \29851 );
buf \U$29858 ( \29853 , \29852 );
not \U$29859 ( \29854 , \29853 );
buf \U$29860 ( \29855 , \1078 );
nand \U$29861 ( \29856 , \29854 , \29855 );
buf \U$29862 ( \29857 , \29856 );
buf \U$29863 ( \29858 , \29857 );
nand \U$29864 ( \29859 , \29848 , \29858 );
buf \U$29865 ( \29860 , \29859 );
buf \U$29866 ( \29861 , \29860 );
xor \U$29867 ( \29862 , \29843 , \29861 );
buf \U$29868 ( \29863 , \12303 );
not \U$29869 ( \29864 , \29863 );
buf \U$29870 ( \29865 , \29864 );
buf \U$29871 ( \29866 , \29865 );
not \U$29872 ( \29867 , \29866 );
buf \U$29873 ( \29868 , \14681 );
not \U$29874 ( \29869 , \29868 );
or \U$29875 ( \29870 , \29867 , \29869 );
buf \U$29876 ( \29871 , RIc0dabe8_115);
nand \U$29877 ( \29872 , \29870 , \29871 );
buf \U$29878 ( \29873 , \29872 );
buf \U$29879 ( \29874 , \29873 );
xor \U$29880 ( \29875 , \29862 , \29874 );
buf \U$29881 ( \29876 , \29875 );
buf \U$29882 ( \29877 , \29876 );
not \U$29883 ( \29878 , \29877 );
buf \U$29884 ( \29879 , \29878 );
buf \U$29885 ( \29880 , \29879 );
not \U$29886 ( \29881 , \29880 );
or \U$29887 ( \29882 , \29826 , \29881 );
buf \U$29888 ( \29883 , \29821 );
buf \U$29889 ( \29884 , \29876 );
nand \U$29890 ( \29885 , \29883 , \29884 );
buf \U$29891 ( \29886 , \29885 );
buf \U$29892 ( \29887 , \29886 );
nand \U$29893 ( \29888 , \29882 , \29887 );
buf \U$29894 ( \29889 , \29888 );
buf \U$29895 ( \29890 , \29889 );
buf \U$29896 ( \29891 , \28764 );
not \U$29897 ( \29892 , \29891 );
buf \U$29898 ( \29893 , \16494 );
not \U$29899 ( \29894 , \29893 );
or \U$29900 ( \29895 , \29892 , \29894 );
buf \U$29901 ( \29896 , \13389 );
buf \U$29902 ( \29897 , RIc0d9928_75);
buf \U$29903 ( \29898 , RIc0d8848_39);
xor \U$29904 ( \29899 , \29897 , \29898 );
buf \U$29905 ( \29900 , \29899 );
buf \U$29906 ( \29901 , \29900 );
nand \U$29907 ( \29902 , \29896 , \29901 );
buf \U$29908 ( \29903 , \29902 );
buf \U$29909 ( \29904 , \29903 );
nand \U$29910 ( \29905 , \29895 , \29904 );
buf \U$29911 ( \29906 , \29905 );
buf \U$29912 ( \29907 , \28781 );
not \U$29913 ( \29908 , \29907 );
buf \U$29914 ( \29909 , \16989 );
not \U$29915 ( \29910 , \29909 );
or \U$29916 ( \29911 , \29908 , \29910 );
buf \U$29917 ( \29912 , \12410 );
buf \U$29918 ( \29913 , RIc0daaf8_113);
buf \U$29919 ( \29914 , RIc0d7678_1);
xor \U$29920 ( \29915 , \29913 , \29914 );
buf \U$29921 ( \29916 , \29915 );
buf \U$29922 ( \29917 , \29916 );
nand \U$29923 ( \29918 , \29912 , \29917 );
buf \U$29924 ( \29919 , \29918 );
buf \U$29925 ( \29920 , \29919 );
nand \U$29926 ( \29921 , \29911 , \29920 );
buf \U$29927 ( \29922 , \29921 );
xor \U$29928 ( \29923 , \29906 , \29922 );
buf \U$29929 ( \29924 , \29048 );
not \U$29930 ( \29925 , \29924 );
buf \U$29931 ( \29926 , \1183 );
not \U$29932 ( \29927 , \29926 );
or \U$29933 ( \29928 , \29925 , \29927 );
buf \U$29934 ( \29929 , RIc0d9a18_77);
buf \U$29935 ( \29930 , RIc0d8758_37);
xnor \U$29936 ( \29931 , \29929 , \29930 );
buf \U$29937 ( \29932 , \29931 );
buf \U$29938 ( \29933 , \29932 );
not \U$29939 ( \29934 , \29933 );
buf \U$29940 ( \29935 , \6141 );
nand \U$29941 ( \29936 , \29934 , \29935 );
buf \U$29942 ( \29937 , \29936 );
buf \U$29943 ( \29938 , \29937 );
nand \U$29944 ( \29939 , \29928 , \29938 );
buf \U$29945 ( \29940 , \29939 );
xnor \U$29946 ( \29941 , \29923 , \29940 );
buf \U$29947 ( \29942 , \29941 );
not \U$29948 ( \29943 , \29942 );
buf \U$29949 ( \29944 , \29943 );
buf \U$29950 ( \29945 , \29944 );
and \U$29951 ( \29946 , \29890 , \29945 );
not \U$29952 ( \29947 , \29890 );
buf \U$29953 ( \29948 , \29941 );
and \U$29954 ( \29949 , \29947 , \29948 );
nor \U$29955 ( \29950 , \29946 , \29949 );
buf \U$29956 ( \29951 , \29950 );
buf \U$29957 ( \29952 , \29951 );
not \U$29958 ( \29953 , \29952 );
buf \U$29959 ( \29954 , \28987 );
not \U$29960 ( \29955 , \29954 );
buf \U$29961 ( \29956 , \14940 );
not \U$29962 ( \29957 , \29956 );
or \U$29963 ( \29958 , \29955 , \29957 );
buf \U$29964 ( \29959 , \402 );
buf \U$29965 ( \29960 , RIc0d8668_35);
buf \U$29966 ( \29961 , RIc0d9b08_79);
xor \U$29967 ( \29962 , \29960 , \29961 );
buf \U$29968 ( \29963 , \29962 );
buf \U$29969 ( \29964 , \29963 );
nand \U$29970 ( \29965 , \29959 , \29964 );
buf \U$29971 ( \29966 , \29965 );
buf \U$29972 ( \29967 , \29966 );
nand \U$29973 ( \29968 , \29958 , \29967 );
buf \U$29974 ( \29969 , \29968 );
buf \U$29975 ( \29970 , \29969 );
buf \U$29976 ( \29971 , \28835 );
not \U$29977 ( \29972 , \29971 );
buf \U$29978 ( \29973 , \476 );
not \U$29979 ( \29974 , \29973 );
or \U$29980 ( \29975 , \29972 , \29974 );
buf \U$29981 ( \29976 , \481 );
buf \U$29982 ( \29977 , RIc0da198_93);
buf \U$29983 ( \29978 , RIc0d7fd8_21);
xor \U$29984 ( \29979 , \29977 , \29978 );
buf \U$29985 ( \29980 , \29979 );
buf \U$29986 ( \29981 , \29980 );
nand \U$29987 ( \29982 , \29976 , \29981 );
buf \U$29988 ( \29983 , \29982 );
buf \U$29989 ( \29984 , \29983 );
nand \U$29990 ( \29985 , \29975 , \29984 );
buf \U$29991 ( \29986 , \29985 );
buf \U$29992 ( \29987 , \29986 );
xor \U$29993 ( \29988 , \29970 , \29987 );
buf \U$29994 ( \29989 , \29092 );
not \U$29995 ( \29990 , \29989 );
buf \U$29996 ( \29991 , \21959 );
not \U$29997 ( \29992 , \29991 );
or \U$29998 ( \29993 , \29990 , \29992 );
buf \U$29999 ( \29994 , \20211 );
buf \U$30000 ( \29995 , RIc0d7858_5);
buf \U$30001 ( \29996 , RIc0da918_109);
xor \U$30002 ( \29997 , \29995 , \29996 );
buf \U$30003 ( \29998 , \29997 );
buf \U$30004 ( \29999 , \29998 );
nand \U$30005 ( \30000 , \29994 , \29999 );
buf \U$30006 ( \30001 , \30000 );
buf \U$30007 ( \30002 , \30001 );
nand \U$30008 ( \30003 , \29993 , \30002 );
buf \U$30009 ( \30004 , \30003 );
buf \U$30010 ( \30005 , \30004 );
xor \U$30011 ( \30006 , \29988 , \30005 );
buf \U$30012 ( \30007 , \30006 );
buf \U$30013 ( \30008 , \30007 );
not \U$30014 ( \30009 , \30008 );
buf \U$30015 ( \30010 , \30009 );
buf \U$30016 ( \30011 , \30010 );
not \U$30017 ( \30012 , \30011 );
buf \U$30018 ( \30013 , \28709 );
not \U$30019 ( \30014 , \30013 );
buf \U$30020 ( \30015 , \21461 );
not \U$30021 ( \30016 , \30015 );
or \U$30022 ( \30017 , \30014 , \30016 );
buf \U$30023 ( \30018 , \22006 );
buf \U$30024 ( \30019 , RIc0da468_99);
buf \U$30025 ( \30020 , RIc0d7d08_15);
xor \U$30026 ( \30021 , \30019 , \30020 );
buf \U$30027 ( \30022 , \30021 );
buf \U$30028 ( \30023 , \30022 );
nand \U$30029 ( \30024 , \30018 , \30023 );
buf \U$30030 ( \30025 , \30024 );
buf \U$30031 ( \30026 , \30025 );
nand \U$30032 ( \30027 , \30017 , \30026 );
buf \U$30033 ( \30028 , \30027 );
buf \U$30034 ( \30029 , \30028 );
not \U$30035 ( \30030 , \30029 );
buf \U$30036 ( \30031 , \28692 );
not \U$30037 ( \30032 , \30031 );
buf \U$30038 ( \30033 , \14346 );
not \U$30039 ( \30034 , \30033 );
or \U$30040 ( \30035 , \30032 , \30034 );
buf \U$30041 ( \30036 , \14353 );
xor \U$30042 ( \30037 , RIc0daa08_111, RIc0d7768_3);
buf \U$30043 ( \30038 , \30037 );
nand \U$30044 ( \30039 , \30036 , \30038 );
buf \U$30045 ( \30040 , \30039 );
buf \U$30046 ( \30041 , \30040 );
nand \U$30047 ( \30042 , \30035 , \30041 );
buf \U$30048 ( \30043 , \30042 );
buf \U$30049 ( \30044 , \30043 );
not \U$30050 ( \30045 , \30044 );
buf \U$30051 ( \30046 , \30045 );
buf \U$30052 ( \30047 , \30046 );
not \U$30053 ( \30048 , \30047 );
or \U$30054 ( \30049 , \30030 , \30048 );
buf \U$30055 ( \30050 , \30028 );
buf \U$30056 ( \30051 , \30046 );
or \U$30057 ( \30052 , \30050 , \30051 );
nand \U$30058 ( \30053 , \30049 , \30052 );
buf \U$30059 ( \30054 , \30053 );
buf \U$30060 ( \30055 , \30054 );
buf \U$30061 ( \30056 , \26411 );
not \U$30062 ( \30057 , \30056 );
buf \U$30063 ( \30058 , \28870 );
not \U$30064 ( \30059 , \30058 );
and \U$30065 ( \30060 , \30057 , \30059 );
buf \U$30066 ( \30061 , \2960 );
buf \U$30067 ( \30062 , RIc0d9dd8_85);
buf \U$30068 ( \30063 , RIc0d8398_29);
xor \U$30069 ( \30064 , \30062 , \30063 );
buf \U$30070 ( \30065 , \30064 );
buf \U$30071 ( \30066 , \30065 );
and \U$30072 ( \30067 , \30061 , \30066 );
nor \U$30073 ( \30068 , \30060 , \30067 );
buf \U$30074 ( \30069 , \30068 );
buf \U$30075 ( \30070 , \30069 );
and \U$30076 ( \30071 , \30055 , \30070 );
not \U$30077 ( \30072 , \30055 );
buf \U$30078 ( \30073 , \30069 );
not \U$30079 ( \30074 , \30073 );
buf \U$30080 ( \30075 , \30074 );
buf \U$30081 ( \30076 , \30075 );
and \U$30082 ( \30077 , \30072 , \30076 );
nor \U$30083 ( \30078 , \30071 , \30077 );
buf \U$30084 ( \30079 , \30078 );
buf \U$30085 ( \30080 , \30079 );
not \U$30086 ( \30081 , \30080 );
buf \U$30087 ( \30082 , \30081 );
buf \U$30088 ( \30083 , \30082 );
not \U$30089 ( \30084 , \30083 );
or \U$30090 ( \30085 , \30012 , \30084 );
buf \U$30091 ( \30086 , \30079 );
buf \U$30092 ( \30087 , \30007 );
nand \U$30093 ( \30088 , \30086 , \30087 );
buf \U$30094 ( \30089 , \30088 );
buf \U$30095 ( \30090 , \30089 );
nand \U$30096 ( \30091 , \30085 , \30090 );
buf \U$30097 ( \30092 , \30091 );
buf \U$30098 ( \30093 , \30092 );
buf \U$30099 ( \30094 , \29582 );
not \U$30100 ( \30095 , \30094 );
buf \U$30101 ( \30096 , \3535 );
not \U$30102 ( \30097 , \30096 );
or \U$30103 ( \30098 , \30095 , \30097 );
buf \U$30104 ( \30099 , \15550 );
xor \U$30105 ( \30100 , RIc0da558_101, RIc0d7c18_13);
buf \U$30106 ( \30101 , \30100 );
nand \U$30107 ( \30102 , \30099 , \30101 );
buf \U$30108 ( \30103 , \30102 );
buf \U$30109 ( \30104 , \30103 );
nand \U$30110 ( \30105 , \30098 , \30104 );
buf \U$30111 ( \30106 , \30105 );
buf \U$30112 ( \30107 , \28914 );
not \U$30113 ( \30108 , \30107 );
buf \U$30114 ( \30109 , \776 );
not \U$30115 ( \30110 , \30109 );
or \U$30116 ( \30111 , \30108 , \30110 );
buf \U$30117 ( \30112 , \792 );
buf \U$30118 ( \30113 , RIc0d9838_73);
buf \U$30119 ( \30114 , RIc0d8938_41);
xor \U$30120 ( \30115 , \30113 , \30114 );
buf \U$30121 ( \30116 , \30115 );
buf \U$30122 ( \30117 , \30116 );
nand \U$30123 ( \30118 , \30112 , \30117 );
buf \U$30124 ( \30119 , \30118 );
buf \U$30125 ( \30120 , \30119 );
nand \U$30126 ( \30121 , \30111 , \30120 );
buf \U$30127 ( \30122 , \30121 );
buf \U$30128 ( \30123 , \30122 );
not \U$30129 ( \30124 , \30123 );
buf \U$30130 ( \30125 , \30124 );
xor \U$30131 ( \30126 , \30106 , \30125 );
buf \U$30132 ( \30127 , \615 );
not \U$30133 ( \30128 , \30127 );
buf \U$30134 ( \30129 , \29530 );
not \U$30135 ( \30130 , \30129 );
buf \U$30136 ( \30131 , \30130 );
buf \U$30137 ( \30132 , \30131 );
not \U$30138 ( \30133 , \30132 );
and \U$30139 ( \30134 , \30128 , \30133 );
buf \U$30140 ( \30135 , \634 );
xnor \U$30141 ( \30136 , RIc0d9ec8_87, RIc0d82a8_27);
buf \U$30142 ( \30137 , \30136 );
nor \U$30143 ( \30138 , \30135 , \30137 );
buf \U$30144 ( \30139 , \30138 );
buf \U$30145 ( \30140 , \30139 );
nor \U$30146 ( \30141 , \30134 , \30140 );
buf \U$30147 ( \30142 , \30141 );
buf \U$30148 ( \30143 , \30142 );
not \U$30149 ( \30144 , \30143 );
buf \U$30150 ( \30145 , \30144 );
xor \U$30151 ( \30146 , \30126 , \30145 );
buf \U$30152 ( \30147 , \30146 );
and \U$30153 ( \30148 , \30093 , \30147 );
not \U$30154 ( \30149 , \30093 );
buf \U$30155 ( \30150 , \30146 );
not \U$30156 ( \30151 , \30150 );
buf \U$30157 ( \30152 , \30151 );
buf \U$30158 ( \30153 , \30152 );
and \U$30159 ( \30154 , \30149 , \30153 );
nor \U$30160 ( \30155 , \30148 , \30154 );
buf \U$30161 ( \30156 , \30155 );
buf \U$30162 ( \30157 , \30156 );
not \U$30163 ( \30158 , \30157 );
or \U$30164 ( \30159 , \29953 , \30158 );
buf \U$30165 ( \30160 , \29951 );
buf \U$30166 ( \30161 , \30156 );
or \U$30167 ( \30162 , \30160 , \30161 );
nand \U$30168 ( \30163 , \30159 , \30162 );
buf \U$30169 ( \30164 , \30163 );
buf \U$30170 ( \30165 , \30164 );
buf \U$30171 ( \30166 , \28733 );
not \U$30172 ( \30167 , \30166 );
buf \U$30173 ( \30168 , \2923 );
not \U$30174 ( \30169 , \30168 );
or \U$30175 ( \30170 , \30167 , \30169 );
buf \U$30176 ( \30171 , \2927 );
xor \U$30177 ( \30172 , RIc0d9748_71, RIc0d8a28_43);
buf \U$30178 ( \30173 , \30172 );
nand \U$30179 ( \30174 , \30171 , \30173 );
buf \U$30180 ( \30175 , \30174 );
buf \U$30181 ( \30176 , \30175 );
nand \U$30182 ( \30177 , \30170 , \30176 );
buf \U$30183 ( \30178 , \30177 );
buf \U$30184 ( \30179 , \30178 );
buf \U$30185 ( \30180 , \28970 );
not \U$30186 ( \30181 , \30180 );
buf \U$30187 ( \30182 , \1224 );
not \U$30188 ( \30183 , \30182 );
or \U$30189 ( \30184 , \30181 , \30183 );
buf \U$30190 ( \30185 , \1229 );
buf \U$30191 ( \30186 , RIc0d9478_65);
buf \U$30192 ( \30187 , RIc0d8cf8_49);
xor \U$30193 ( \30188 , \30186 , \30187 );
buf \U$30194 ( \30189 , \30188 );
buf \U$30195 ( \30190 , \30189 );
nand \U$30196 ( \30191 , \30185 , \30190 );
buf \U$30197 ( \30192 , \30191 );
buf \U$30198 ( \30193 , \30192 );
nand \U$30199 ( \30194 , \30184 , \30193 );
buf \U$30200 ( \30195 , \30194 );
buf \U$30201 ( \30196 , \30195 );
xor \U$30202 ( \30197 , \30179 , \30196 );
buf \U$30203 ( \30198 , \749 );
buf \U$30204 ( \30199 , \29074 );
not \U$30205 ( \30200 , \30199 );
buf \U$30206 ( \30201 , \30200 );
buf \U$30207 ( \30202 , \30201 );
or \U$30208 ( \30203 , \30198 , \30202 );
buf \U$30209 ( \30204 , \737 );
buf \U$30210 ( \30205 , RIc0da378_97);
buf \U$30211 ( \30206 , RIc0d7df8_17);
xor \U$30212 ( \30207 , \30205 , \30206 );
buf \U$30213 ( \30208 , \30207 );
buf \U$30214 ( \30209 , \30208 );
not \U$30215 ( \30210 , \30209 );
buf \U$30216 ( \30211 , \30210 );
buf \U$30217 ( \30212 , \30211 );
or \U$30218 ( \30213 , \30204 , \30212 );
nand \U$30219 ( \30214 , \30203 , \30213 );
buf \U$30220 ( \30215 , \30214 );
buf \U$30221 ( \30216 , \30215 );
xor \U$30222 ( \30217 , \30197 , \30216 );
buf \U$30223 ( \30218 , \30217 );
buf \U$30224 ( \30219 , \30218 );
not \U$30225 ( \30220 , \30219 );
buf \U$30226 ( \30221 , \29618 );
not \U$30227 ( \30222 , \30221 );
buf \U$30228 ( \30223 , \330 );
not \U$30229 ( \30224 , \30223 );
or \U$30230 ( \30225 , \30222 , \30224 );
buf \U$30231 ( \30226 , \14707 );
buf \U$30232 ( \30227 , RIc0da288_95);
buf \U$30233 ( \30228 , RIc0d7ee8_19);
xor \U$30234 ( \30229 , \30227 , \30228 );
buf \U$30235 ( \30230 , \30229 );
buf \U$30236 ( \30231 , \30230 );
nand \U$30237 ( \30232 , \30226 , \30231 );
buf \U$30238 ( \30233 , \30232 );
buf \U$30239 ( \30234 , \30233 );
nand \U$30240 ( \30235 , \30225 , \30234 );
buf \U$30241 ( \30236 , \30235 );
buf \U$30242 ( \30237 , \29554 );
not \U$30243 ( \30238 , \30237 );
buf \U$30244 ( \30239 , \17405 );
not \U$30245 ( \30240 , \30239 );
or \U$30246 ( \30241 , \30238 , \30240 );
buf \U$30247 ( \30242 , \13048 );
buf \U$30248 ( \30243 , RIc0da648_103);
buf \U$30249 ( \30244 , RIc0d7b28_11);
xor \U$30250 ( \30245 , \30243 , \30244 );
buf \U$30251 ( \30246 , \30245 );
buf \U$30252 ( \30247 , \30246 );
nand \U$30253 ( \30248 , \30242 , \30247 );
buf \U$30254 ( \30249 , \30248 );
buf \U$30255 ( \30250 , \30249 );
nand \U$30256 ( \30251 , \30241 , \30250 );
buf \U$30257 ( \30252 , \30251 );
xor \U$30258 ( \30253 , \30236 , \30252 );
buf \U$30259 ( \30254 , \28936 );
not \U$30260 ( \30255 , \30254 );
buf \U$30261 ( \30256 , \12736 );
not \U$30262 ( \30257 , \30256 );
or \U$30263 ( \30258 , \30255 , \30257 );
buf \U$30264 ( \30259 , \21880 );
buf \U$30265 ( \30260 , RIc0d7a38_9);
buf \U$30266 ( \30261 , RIc0da738_105);
xor \U$30267 ( \30262 , \30260 , \30261 );
buf \U$30268 ( \30263 , \30262 );
buf \U$30269 ( \30264 , \30263 );
nand \U$30270 ( \30265 , \30259 , \30264 );
buf \U$30271 ( \30266 , \30265 );
buf \U$30272 ( \30267 , \30266 );
nand \U$30273 ( \30268 , \30258 , \30267 );
buf \U$30274 ( \30269 , \30268 );
xnor \U$30275 ( \30270 , \30253 , \30269 );
buf \U$30276 ( \30271 , \30270 );
not \U$30277 ( \30272 , \30271 );
or \U$30278 ( \30273 , \30220 , \30272 );
buf \U$30279 ( \30274 , \30270 );
buf \U$30280 ( \30275 , \30218 );
or \U$30281 ( \30276 , \30274 , \30275 );
nand \U$30282 ( \30277 , \30273 , \30276 );
buf \U$30283 ( \30278 , \30277 );
buf \U$30284 ( \30279 , \30278 );
and \U$30285 ( \30280 , \28118 , \28119 );
buf \U$30286 ( \30281 , \30280 );
buf \U$30287 ( \30282 , \30281 );
buf \U$30288 ( \30283 , \28897 );
not \U$30289 ( \30284 , \30283 );
buf \U$30290 ( \30285 , \678 );
not \U$30291 ( \30286 , \30285 );
or \U$30292 ( \30287 , \30284 , \30286 );
buf \U$30293 ( \30288 , \686 );
xor \U$30294 ( \30289 , RIc0d9568_67, RIc0d8c08_47);
buf \U$30295 ( \30290 , \30289 );
nand \U$30296 ( \30291 , \30288 , \30290 );
buf \U$30297 ( \30292 , \30291 );
buf \U$30298 ( \30293 , \30292 );
nand \U$30299 ( \30294 , \30287 , \30293 );
buf \U$30300 ( \30295 , \30294 );
buf \U$30301 ( \30296 , \30295 );
xor \U$30302 ( \30297 , \30282 , \30296 );
buf \U$30303 ( \30298 , \521 );
buf \U$30304 ( \30299 , \28851 );
or \U$30305 ( \30300 , \30298 , \30299 );
buf \U$30306 ( \30301 , \1933 );
not \U$30307 ( \30302 , \30301 );
buf \U$30308 ( \30303 , \30302 );
buf \U$30309 ( \30304 , \30303 );
buf \U$30310 ( \30305 , RIc0da0a8_91);
buf \U$30311 ( \30306 , RIc0d80c8_23);
xnor \U$30312 ( \30307 , \30305 , \30306 );
buf \U$30313 ( \30308 , \30307 );
buf \U$30314 ( \30309 , \30308 );
or \U$30315 ( \30310 , \30304 , \30309 );
nand \U$30316 ( \30311 , \30300 , \30310 );
buf \U$30317 ( \30312 , \30311 );
buf \U$30318 ( \30313 , \30312 );
xor \U$30319 ( \30314 , \30297 , \30313 );
buf \U$30320 ( \30315 , \30314 );
buf \U$30321 ( \30316 , \30315 );
not \U$30322 ( \30317 , \30316 );
buf \U$30323 ( \30318 , \30317 );
buf \U$30324 ( \30319 , \30318 );
and \U$30325 ( \30320 , \30279 , \30319 );
not \U$30326 ( \30321 , \30279 );
buf \U$30327 ( \30322 , \30315 );
and \U$30328 ( \30323 , \30321 , \30322 );
nor \U$30329 ( \30324 , \30320 , \30323 );
buf \U$30330 ( \30325 , \30324 );
buf \U$30331 ( \30326 , \30325 );
and \U$30332 ( \30327 , \30165 , \30326 );
not \U$30333 ( \30328 , \30165 );
buf \U$30334 ( \30329 , \30325 );
not \U$30335 ( \30330 , \30329 );
buf \U$30336 ( \30331 , \30330 );
buf \U$30337 ( \30332 , \30331 );
and \U$30338 ( \30333 , \30328 , \30332 );
or \U$30339 ( \30334 , \30327 , \30333 );
buf \U$30340 ( \30335 , \30334 );
buf \U$30341 ( \30336 , \30335 );
xor \U$30342 ( \30337 , \29771 , \30336 );
buf \U$30343 ( \30338 , \30337 );
buf \U$30344 ( \30339 , \30338 );
xor \U$30345 ( \30340 , \29647 , \30339 );
buf \U$30346 ( \30341 , \30340 );
buf \U$30347 ( \30342 , \30341 );
not \U$30348 ( \30343 , \30342 );
buf \U$30349 ( \30344 , \30343 );
buf \U$30350 ( \30345 , \30344 );
not \U$30351 ( \30346 , \30345 );
buf \U$30352 ( \30347 , \27954 );
not \U$30353 ( \30348 , \30347 );
buf \U$30354 ( \30349 , \15644 );
not \U$30355 ( \30350 , \30349 );
or \U$30356 ( \30351 , \30348 , \30350 );
buf \U$30357 ( \30352 , \12744 );
buf \U$30358 ( \30353 , \28926 );
nand \U$30359 ( \30354 , \30352 , \30353 );
buf \U$30360 ( \30355 , \30354 );
buf \U$30361 ( \30356 , \30355 );
nand \U$30362 ( \30357 , \30351 , \30356 );
buf \U$30363 ( \30358 , \30357 );
xor \U$30364 ( \30359 , RIc0dacd8_117, RIc0d7678_1);
buf \U$30365 ( \30360 , \30359 );
not \U$30366 ( \30361 , \30360 );
buf \U$30367 ( \30362 , \12923 );
not \U$30368 ( \30363 , \30362 );
or \U$30369 ( \30364 , \30361 , \30363 );
buf \U$30370 ( \30365 , \12936 );
buf \U$30371 ( \30366 , RIc0dacd8_117);
nand \U$30372 ( \30367 , \30365 , \30366 );
buf \U$30373 ( \30368 , \30367 );
buf \U$30374 ( \30369 , \30368 );
nand \U$30375 ( \30370 , \30364 , \30369 );
buf \U$30376 ( \30371 , \30370 );
buf \U$30377 ( \30372 , \30371 );
not \U$30378 ( \30373 , \30372 );
buf \U$30379 ( \30374 , \30373 );
xor \U$30380 ( \30375 , \30358 , \30374 );
buf \U$30381 ( \30376 , RIc0d7a38_9);
buf \U$30382 ( \30377 , RIc0da918_109);
xor \U$30383 ( \30378 , \30376 , \30377 );
buf \U$30384 ( \30379 , \30378 );
buf \U$30385 ( \30380 , \30379 );
not \U$30386 ( \30381 , \30380 );
buf \U$30387 ( \30382 , \13419 );
not \U$30388 ( \30383 , \30382 );
or \U$30389 ( \30384 , \30381 , \30383 );
buf \U$30390 ( \30385 , \20211 );
buf \U$30391 ( \30386 , \28285 );
nand \U$30392 ( \30387 , \30385 , \30386 );
buf \U$30393 ( \30388 , \30387 );
buf \U$30394 ( \30389 , \30388 );
nand \U$30395 ( \30390 , \30384 , \30389 );
buf \U$30396 ( \30391 , \30390 );
buf \U$30397 ( \30392 , \30391 );
buf \U$30398 ( \30393 , RIc0d7fd8_21);
buf \U$30399 ( \30394 , RIc0da378_97);
xor \U$30400 ( \30395 , \30393 , \30394 );
buf \U$30401 ( \30396 , \30395 );
buf \U$30402 ( \30397 , \30396 );
not \U$30403 ( \30398 , \30397 );
buf \U$30404 ( \30399 , \16086 );
not \U$30405 ( \30400 , \30399 );
or \U$30406 ( \30401 , \30398 , \30400 );
buf \U$30407 ( \30402 , \2070 );
buf \U$30408 ( \30403 , \28154 );
nand \U$30409 ( \30404 , \30402 , \30403 );
buf \U$30410 ( \30405 , \30404 );
buf \U$30411 ( \30406 , \30405 );
nand \U$30412 ( \30407 , \30401 , \30406 );
buf \U$30413 ( \30408 , \30407 );
buf \U$30414 ( \30409 , \30408 );
nor \U$30415 ( \30410 , \30392 , \30409 );
buf \U$30416 ( \30411 , \30410 );
buf \U$30417 ( \30412 , \30411 );
buf \U$30418 ( \30413 , \2091 );
not \U$30419 ( \30414 , \30413 );
buf \U$30420 ( \30415 , RIc0d8668_35);
buf \U$30421 ( \30416 , RIc0d9ce8_83);
xor \U$30422 ( \30417 , \30415 , \30416 );
buf \U$30423 ( \30418 , \30417 );
buf \U$30424 ( \30419 , \30418 );
not \U$30425 ( \30420 , \30419 );
buf \U$30426 ( \30421 , \30420 );
buf \U$30427 ( \30422 , \30421 );
not \U$30428 ( \30423 , \30422 );
and \U$30429 ( \30424 , \30414 , \30423 );
buf \U$30430 ( \30425 , \584 );
buf \U$30431 ( \30426 , \28048 );
and \U$30432 ( \30427 , \30425 , \30426 );
buf \U$30433 ( \30428 , \30427 );
buf \U$30434 ( \30429 , \30428 );
nor \U$30435 ( \30430 , \30424 , \30429 );
buf \U$30436 ( \30431 , \30430 );
buf \U$30437 ( \30432 , \30431 );
or \U$30438 ( \30433 , \30412 , \30432 );
buf \U$30439 ( \30434 , \30408 );
buf \U$30440 ( \30435 , \30391 );
nand \U$30441 ( \30436 , \30434 , \30435 );
buf \U$30442 ( \30437 , \30436 );
buf \U$30443 ( \30438 , \30437 );
nand \U$30444 ( \30439 , \30433 , \30438 );
buf \U$30445 ( \30440 , \30439 );
xnor \U$30446 ( \30441 , \30375 , \30440 );
buf \U$30447 ( \30442 , \30441 );
not \U$30448 ( \30443 , \30442 );
buf \U$30449 ( \30444 , \30443 );
buf \U$30450 ( \30445 , \30444 );
not \U$30451 ( \30446 , \30445 );
xor \U$30452 ( \30447 , \28597 , \28617 );
not \U$30453 ( \30448 , \28575 );
xor \U$30454 ( \30449 , \30447 , \30448 );
buf \U$30455 ( \30450 , \30449 );
not \U$30456 ( \30451 , \30450 );
xor \U$30457 ( \30452 , \28495 , \28513 );
xor \U$30458 ( \30453 , \30452 , \28538 );
buf \U$30459 ( \30454 , \30453 );
buf \U$30460 ( \30455 , \30454 );
not \U$30461 ( \30456 , \30455 );
or \U$30462 ( \30457 , \30451 , \30456 );
buf \U$30463 ( \30458 , \30449 );
buf \U$30464 ( \30459 , \30454 );
or \U$30465 ( \30460 , \30458 , \30459 );
nand \U$30466 ( \30461 , \30457 , \30460 );
buf \U$30467 ( \30462 , \30461 );
buf \U$30468 ( \30463 , \30462 );
not \U$30469 ( \30464 , \30463 );
or \U$30470 ( \30465 , \30446 , \30464 );
buf \U$30471 ( \30466 , \30462 );
buf \U$30472 ( \30467 , \30444 );
or \U$30473 ( \30468 , \30466 , \30467 );
nand \U$30474 ( \30469 , \30465 , \30468 );
buf \U$30475 ( \30470 , \30469 );
buf \U$30476 ( \30471 , \30470 );
buf \U$30477 ( \30472 , \30374 );
buf \U$30478 ( \30473 , \29444 );
not \U$30479 ( \30474 , \30473 );
buf \U$30480 ( \30475 , \12402 );
not \U$30481 ( \30476 , \30475 );
or \U$30482 ( \30477 , \30474 , \30476 );
buf \U$30483 ( \30478 , \16662 );
buf \U$30484 ( \30479 , RIc0d7858_5);
buf \U$30485 ( \30480 , RIc0daaf8_113);
xor \U$30486 ( \30481 , \30479 , \30480 );
buf \U$30487 ( \30482 , \30481 );
buf \U$30488 ( \30483 , \30482 );
nand \U$30489 ( \30484 , \30478 , \30483 );
buf \U$30490 ( \30485 , \30484 );
buf \U$30491 ( \30486 , \30485 );
nand \U$30492 ( \30487 , \30477 , \30486 );
buf \U$30493 ( \30488 , \30487 );
buf \U$30494 ( \30489 , \30488 );
not \U$30495 ( \30490 , \30489 );
buf \U$30496 ( \30491 , RIc0d8aa0_44);
buf \U$30497 ( \30492 , RIc0d9928_75);
xor \U$30498 ( \30493 , \30491 , \30492 );
buf \U$30499 ( \30494 , \30493 );
buf \U$30500 ( \30495 , \30494 );
not \U$30501 ( \30496 , \30495 );
buf \U$30502 ( \30497 , \2358 );
not \U$30503 ( \30498 , \30497 );
or \U$30504 ( \30499 , \30496 , \30498 );
buf \U$30505 ( \30500 , \1143 );
buf \U$30506 ( \30501 , \27925 );
nand \U$30507 ( \30502 , \30500 , \30501 );
buf \U$30508 ( \30503 , \30502 );
buf \U$30509 ( \30504 , \30503 );
nand \U$30510 ( \30505 , \30499 , \30504 );
buf \U$30511 ( \30506 , \30505 );
buf \U$30512 ( \30507 , \30506 );
not \U$30513 ( \30508 , \30507 );
or \U$30514 ( \30509 , \30490 , \30508 );
buf \U$30515 ( \30510 , \30506 );
buf \U$30516 ( \30511 , \30488 );
or \U$30517 ( \30512 , \30510 , \30511 );
buf \U$30518 ( \30513 , RIc0d9a18_77);
buf \U$30519 ( \30514 , RIc0d89b0_42);
xor \U$30520 ( \30515 , \30513 , \30514 );
buf \U$30521 ( \30516 , \30515 );
buf \U$30522 ( \30517 , \30516 );
not \U$30523 ( \30518 , \30517 );
buf \U$30524 ( \30519 , \1431 );
not \U$30525 ( \30520 , \30519 );
or \U$30526 ( \30521 , \30518 , \30520 );
buf \U$30527 ( \30522 , \3742 );
buf \U$30528 ( \30523 , \27900 );
nand \U$30529 ( \30524 , \30522 , \30523 );
buf \U$30530 ( \30525 , \30524 );
buf \U$30531 ( \30526 , \30525 );
nand \U$30532 ( \30527 , \30521 , \30526 );
buf \U$30533 ( \30528 , \30527 );
buf \U$30534 ( \30529 , \30528 );
nand \U$30535 ( \30530 , \30512 , \30529 );
buf \U$30536 ( \30531 , \30530 );
buf \U$30537 ( \30532 , \30531 );
nand \U$30538 ( \30533 , \30509 , \30532 );
buf \U$30539 ( \30534 , \30533 );
buf \U$30540 ( \30535 , \30534 );
xor \U$30541 ( \30536 , \30472 , \30535 );
buf \U$30542 ( \30537 , \29426 );
not \U$30543 ( \30538 , \30537 );
buf \U$30544 ( \30539 , \3292 );
not \U$30545 ( \30540 , \30539 );
or \U$30546 ( \30541 , \30538 , \30540 );
buf \U$30547 ( \30542 , \921 );
buf \U$30548 ( \30543 , RIc0d8578_33);
buf \U$30549 ( \30544 , RIc0d9dd8_85);
xor \U$30550 ( \30545 , \30543 , \30544 );
buf \U$30551 ( \30546 , \30545 );
buf \U$30552 ( \30547 , \30546 );
nand \U$30553 ( \30548 , \30542 , \30547 );
buf \U$30554 ( \30549 , \30548 );
buf \U$30555 ( \30550 , \30549 );
nand \U$30556 ( \30551 , \30541 , \30550 );
buf \U$30557 ( \30552 , \30551 );
buf \U$30558 ( \30553 , \30552 );
buf \U$30559 ( \30554 , \29404 );
not \U$30560 ( \30555 , \30554 );
buf \U$30561 ( \30556 , \2470 );
not \U$30562 ( \30557 , \30556 );
or \U$30563 ( \30558 , \30555 , \30557 );
buf \U$30564 ( \30559 , \14648 );
buf \U$30565 ( \30560 , \29272 );
nand \U$30566 ( \30561 , \30559 , \30560 );
buf \U$30567 ( \30562 , \30561 );
buf \U$30568 ( \30563 , \30562 );
nand \U$30569 ( \30564 , \30558 , \30563 );
buf \U$30570 ( \30565 , \30564 );
buf \U$30571 ( \30566 , \30565 );
xor \U$30572 ( \30567 , \30553 , \30566 );
buf \U$30573 ( \30568 , \29383 );
not \U$30574 ( \30569 , \30568 );
buf \U$30575 ( \30570 , \12529 );
not \U$30576 ( \30571 , \30570 );
or \U$30577 ( \30572 , \30569 , \30571 );
buf \U$30578 ( \30573 , \14353 );
buf \U$30579 ( \30574 , \29252 );
nand \U$30580 ( \30575 , \30573 , \30574 );
buf \U$30581 ( \30576 , \30575 );
buf \U$30582 ( \30577 , \30576 );
nand \U$30583 ( \30578 , \30572 , \30577 );
buf \U$30584 ( \30579 , \30578 );
buf \U$30585 ( \30580 , \30579 );
and \U$30586 ( \30581 , \30567 , \30580 );
and \U$30587 ( \30582 , \30553 , \30566 );
or \U$30588 ( \30583 , \30581 , \30582 );
buf \U$30589 ( \30584 , \30583 );
buf \U$30590 ( \30585 , \30584 );
xnor \U$30591 ( \30586 , \30536 , \30585 );
buf \U$30592 ( \30587 , \30586 );
buf \U$30593 ( \30588 , \30587 );
not \U$30594 ( \30589 , \30588 );
buf \U$30595 ( \30590 , \30589 );
buf \U$30596 ( \30591 , \30590 );
not \U$30597 ( \30592 , \30591 );
buf \U$30598 ( \30593 , RIc0d8500_32);
buf \U$30599 ( \30594 , RIc0d9ec8_87);
xor \U$30600 ( \30595 , \30593 , \30594 );
buf \U$30601 ( \30596 , \30595 );
buf \U$30602 ( \30597 , \30596 );
not \U$30603 ( \30598 , \30597 );
buf \U$30604 ( \30599 , \14325 );
not \U$30605 ( \30600 , \30599 );
or \U$30606 ( \30601 , \30598 , \30600 );
buf \U$30607 ( \30602 , \816 );
buf \U$30608 ( \30603 , RIc0d8488_31);
buf \U$30609 ( \30604 , RIc0d9ec8_87);
xor \U$30610 ( \30605 , \30603 , \30604 );
buf \U$30611 ( \30606 , \30605 );
buf \U$30612 ( \30607 , \30606 );
nand \U$30613 ( \30608 , \30602 , \30607 );
buf \U$30614 ( \30609 , \30608 );
buf \U$30615 ( \30610 , \30609 );
nand \U$30616 ( \30611 , \30601 , \30610 );
buf \U$30617 ( \30612 , \30611 );
buf \U$30618 ( \30613 , \30612 );
not \U$30619 ( \30614 , \30613 );
buf \U$30620 ( \30615 , RIc0d8b90_46);
buf \U$30621 ( \30616 , RIc0d9838_73);
xor \U$30622 ( \30617 , \30615 , \30616 );
buf \U$30623 ( \30618 , \30617 );
buf \U$30624 ( \30619 , \30618 );
not \U$30625 ( \30620 , \30619 );
buf \U$30626 ( \30621 , \14608 );
not \U$30627 ( \30622 , \30621 );
or \U$30628 ( \30623 , \30620 , \30622 );
buf \U$30629 ( \30624 , \1856 );
buf \U$30630 ( \30625 , RIc0d8b18_45);
buf \U$30631 ( \30626 , RIc0d9838_73);
xor \U$30632 ( \30627 , \30625 , \30626 );
buf \U$30633 ( \30628 , \30627 );
buf \U$30634 ( \30629 , \30628 );
nand \U$30635 ( \30630 , \30624 , \30629 );
buf \U$30636 ( \30631 , \30630 );
buf \U$30637 ( \30632 , \30631 );
nand \U$30638 ( \30633 , \30623 , \30632 );
buf \U$30639 ( \30634 , \30633 );
buf \U$30640 ( \30635 , \30634 );
not \U$30641 ( \30636 , \30635 );
or \U$30642 ( \30637 , \30614 , \30636 );
buf \U$30643 ( \30638 , \30612 );
buf \U$30644 ( \30639 , \30634 );
or \U$30645 ( \30640 , \30638 , \30639 );
buf \U$30646 ( \30641 , \29466 );
not \U$30647 ( \30642 , \30641 );
buf \U$30648 ( \30643 , \12833 );
not \U$30649 ( \30644 , \30643 );
or \U$30650 ( \30645 , \30642 , \30644 );
buf \U$30651 ( \30646 , \4049 );
buf \U$30652 ( \30647 , RIc0da558_101);
buf \U$30653 ( \30648 , RIc0d7df8_17);
xor \U$30654 ( \30649 , \30647 , \30648 );
buf \U$30655 ( \30650 , \30649 );
buf \U$30656 ( \30651 , \30650 );
nand \U$30657 ( \30652 , \30646 , \30651 );
buf \U$30658 ( \30653 , \30652 );
buf \U$30659 ( \30654 , \30653 );
nand \U$30660 ( \30655 , \30645 , \30654 );
buf \U$30661 ( \30656 , \30655 );
buf \U$30662 ( \30657 , \30656 );
nand \U$30663 ( \30658 , \30640 , \30657 );
buf \U$30664 ( \30659 , \30658 );
buf \U$30665 ( \30660 , \30659 );
nand \U$30666 ( \30661 , \30637 , \30660 );
buf \U$30667 ( \30662 , \30661 );
buf \U$30668 ( \30663 , RIc0d77e0_4);
buf \U$30669 ( \30664 , RIc0dabe8_115);
xor \U$30670 ( \30665 , \30663 , \30664 );
buf \U$30671 ( \30666 , \30665 );
buf \U$30672 ( \30667 , \30666 );
not \U$30673 ( \30668 , \30667 );
buf \U$30674 ( \30669 , \12299 );
not \U$30675 ( \30670 , \30669 );
or \U$30676 ( \30671 , \30668 , \30670 );
buf \U$30677 ( \30672 , \12303 );
buf \U$30678 ( \30673 , \27970 );
nand \U$30679 ( \30674 , \30672 , \30673 );
buf \U$30680 ( \30675 , \30674 );
buf \U$30681 ( \30676 , \30675 );
nand \U$30682 ( \30677 , \30671 , \30676 );
buf \U$30683 ( \30678 , \30677 );
buf \U$30684 ( \30679 , \30678 );
not \U$30685 ( \30680 , \30679 );
buf \U$30686 ( \30681 , \30680 );
buf \U$30687 ( \30682 , \30681 );
not \U$30688 ( \30683 , \30682 );
buf \U$30689 ( \30684 , RIc0d87d0_38);
buf \U$30690 ( \30685 , RIc0d9bf8_81);
xor \U$30691 ( \30686 , \30684 , \30685 );
buf \U$30692 ( \30687 , \30686 );
buf \U$30693 ( \30688 , \30687 );
not \U$30694 ( \30689 , \30688 );
buf \U$30695 ( \30690 , \13075 );
not \U$30696 ( \30691 , \30690 );
or \U$30697 ( \30692 , \30689 , \30691 );
buf \U$30698 ( \30693 , \1078 );
buf \U$30699 ( \30694 , \27854 );
nand \U$30700 ( \30695 , \30693 , \30694 );
buf \U$30701 ( \30696 , \30695 );
buf \U$30702 ( \30697 , \30696 );
nand \U$30703 ( \30698 , \30692 , \30697 );
buf \U$30704 ( \30699 , \30698 );
buf \U$30705 ( \30700 , \30699 );
not \U$30706 ( \30701 , \30700 );
buf \U$30707 ( \30702 , \30701 );
buf \U$30708 ( \30703 , \30702 );
not \U$30709 ( \30704 , \30703 );
or \U$30710 ( \30705 , \30683 , \30704 );
xor \U$30711 ( \30706 , RIc0dacd8_117, RIc0d76f0_2);
buf \U$30712 ( \30707 , \30706 );
not \U$30713 ( \30708 , \30707 );
buf \U$30714 ( \30709 , \13684 );
not \U$30715 ( \30710 , \30709 );
or \U$30716 ( \30711 , \30708 , \30710 );
buf \U$30717 ( \30712 , \16559 );
buf \U$30718 ( \30713 , \30359 );
nand \U$30719 ( \30714 , \30712 , \30713 );
buf \U$30720 ( \30715 , \30714 );
buf \U$30721 ( \30716 , \30715 );
nand \U$30722 ( \30717 , \30711 , \30716 );
buf \U$30723 ( \30718 , \30717 );
buf \U$30724 ( \30719 , \30718 );
nand \U$30725 ( \30720 , \30705 , \30719 );
buf \U$30726 ( \30721 , \30720 );
buf \U$30727 ( \30722 , \30721 );
buf \U$30728 ( \30723 , \30678 );
buf \U$30729 ( \30724 , \30699 );
nand \U$30730 ( \30725 , \30723 , \30724 );
buf \U$30731 ( \30726 , \30725 );
buf \U$30732 ( \30727 , \30726 );
nand \U$30733 ( \30728 , \30722 , \30727 );
buf \U$30734 ( \30729 , \30728 );
buf \U$30735 ( \30730 , \30729 );
not \U$30736 ( \30731 , \30730 );
buf \U$30737 ( \30732 , \30731 );
xor \U$30738 ( \30733 , \30662 , \30732 );
xor \U$30739 ( \30734 , RIc0da288_95, RIc0d8140_24);
buf \U$30740 ( \30735 , \30734 );
not \U$30741 ( \30736 , \30735 );
buf \U$30742 ( \30737 , \3714 );
not \U$30743 ( \30738 , \30737 );
or \U$30744 ( \30739 , \30736 , \30738 );
buf \U$30745 ( \30740 , \344 );
xor \U$30746 ( \30741 , RIc0da288_95, RIc0d80c8_23);
buf \U$30747 ( \30742 , \30741 );
nand \U$30748 ( \30743 , \30740 , \30742 );
buf \U$30749 ( \30744 , \30743 );
buf \U$30750 ( \30745 , \30744 );
nand \U$30751 ( \30746 , \30739 , \30745 );
buf \U$30752 ( \30747 , \30746 );
buf \U$30753 ( \30748 , \30747 );
not \U$30754 ( \30749 , \30748 );
buf \U$30755 ( \30750 , RIc0d8410_30);
buf \U$30756 ( \30751 , RIc0d9fb8_89);
xor \U$30757 ( \30752 , \30750 , \30751 );
buf \U$30758 ( \30753 , \30752 );
buf \U$30759 ( \30754 , \30753 );
not \U$30760 ( \30755 , \30754 );
buf \U$30761 ( \30756 , \2037 );
not \U$30762 ( \30757 , \30756 );
or \U$30763 ( \30758 , \30755 , \30757 );
buf \U$30764 ( \30759 , \846 );
buf \U$30765 ( \30760 , RIc0d9fb8_89);
buf \U$30766 ( \30761 , RIc0d8398_29);
xor \U$30767 ( \30762 , \30760 , \30761 );
buf \U$30768 ( \30763 , \30762 );
buf \U$30769 ( \30764 , \30763 );
nand \U$30770 ( \30765 , \30759 , \30764 );
buf \U$30771 ( \30766 , \30765 );
buf \U$30772 ( \30767 , \30766 );
nand \U$30773 ( \30768 , \30758 , \30767 );
buf \U$30774 ( \30769 , \30768 );
buf \U$30775 ( \30770 , \30769 );
not \U$30776 ( \30771 , \30770 );
or \U$30777 ( \30772 , \30749 , \30771 );
buf \U$30778 ( \30773 , \30747 );
buf \U$30779 ( \30774 , \30769 );
or \U$30780 ( \30775 , \30773 , \30774 );
buf \U$30781 ( \30776 , RIc0d7d80_16);
buf \U$30782 ( \30777 , RIc0da648_103);
xor \U$30783 ( \30778 , \30776 , \30777 );
buf \U$30784 ( \30779 , \30778 );
buf \U$30785 ( \30780 , \30779 );
not \U$30786 ( \30781 , \30780 );
buf \U$30787 ( \30782 , \15397 );
not \U$30788 ( \30783 , \30782 );
or \U$30789 ( \30784 , \30781 , \30783 );
buf \U$30790 ( \30785 , \15403 );
buf \U$30791 ( \30786 , RIc0d7d08_15);
buf \U$30792 ( \30787 , RIc0da648_103);
xor \U$30793 ( \30788 , \30786 , \30787 );
buf \U$30794 ( \30789 , \30788 );
buf \U$30795 ( \30790 , \30789 );
nand \U$30796 ( \30791 , \30785 , \30790 );
buf \U$30797 ( \30792 , \30791 );
buf \U$30798 ( \30793 , \30792 );
nand \U$30799 ( \30794 , \30784 , \30793 );
buf \U$30800 ( \30795 , \30794 );
buf \U$30801 ( \30796 , \30795 );
nand \U$30802 ( \30797 , \30775 , \30796 );
buf \U$30803 ( \30798 , \30797 );
buf \U$30804 ( \30799 , \30798 );
nand \U$30805 ( \30800 , \30772 , \30799 );
buf \U$30806 ( \30801 , \30800 );
xor \U$30807 ( \30802 , \30733 , \30801 );
buf \U$30808 ( \30803 , \30802 );
not \U$30809 ( \30804 , \30803 );
buf \U$30810 ( \30805 , \30804 );
buf \U$30811 ( \30806 , \30805 );
not \U$30812 ( \30807 , \30806 );
or \U$30813 ( \30808 , \30592 , \30807 );
buf \U$30814 ( \30809 , \30587 );
not \U$30815 ( \30810 , \30809 );
buf \U$30816 ( \30811 , \30802 );
not \U$30817 ( \30812 , \30811 );
or \U$30818 ( \30813 , \30810 , \30812 );
xor \U$30819 ( \30814 , \30553 , \30566 );
xor \U$30820 ( \30815 , \30814 , \30580 );
buf \U$30821 ( \30816 , \30815 );
buf \U$30822 ( \30817 , \30816 );
not \U$30823 ( \30818 , \30817 );
buf \U$30824 ( \30819 , \30634 );
buf \U$30825 ( \30820 , \30612 );
xor \U$30826 ( \30821 , \30819 , \30820 );
buf \U$30827 ( \30822 , \30656 );
xnor \U$30828 ( \30823 , \30821 , \30822 );
buf \U$30829 ( \30824 , \30823 );
buf \U$30830 ( \30825 , \30824 );
not \U$30831 ( \30826 , \30825 );
buf \U$30832 ( \30827 , \30826 );
buf \U$30833 ( \30828 , \30827 );
not \U$30834 ( \30829 , \30828 );
or \U$30835 ( \30830 , \30818 , \30829 );
buf \U$30836 ( \30831 , \30816 );
not \U$30837 ( \30832 , \30831 );
buf \U$30838 ( \30833 , \30832 );
buf \U$30839 ( \30834 , \30833 );
not \U$30840 ( \30835 , \30834 );
buf \U$30841 ( \30836 , \30824 );
not \U$30842 ( \30837 , \30836 );
or \U$30843 ( \30838 , \30835 , \30837 );
xor \U$30844 ( \30839 , \30506 , \30488 );
xor \U$30845 ( \30840 , \30839 , \30528 );
buf \U$30846 ( \30841 , \30840 );
nand \U$30847 ( \30842 , \30838 , \30841 );
buf \U$30848 ( \30843 , \30842 );
buf \U$30849 ( \30844 , \30843 );
nand \U$30850 ( \30845 , \30830 , \30844 );
buf \U$30851 ( \30846 , \30845 );
buf \U$30852 ( \30847 , \30846 );
nand \U$30853 ( \30848 , \30813 , \30847 );
buf \U$30854 ( \30849 , \30848 );
buf \U$30855 ( \30850 , \30849 );
nand \U$30856 ( \30851 , \30808 , \30850 );
buf \U$30857 ( \30852 , \30851 );
buf \U$30858 ( \30853 , \30852 );
xor \U$30859 ( \30854 , \30471 , \30853 );
buf \U$30860 ( \30855 , \30374 );
not \U$30861 ( \30856 , \30855 );
buf \U$30862 ( \30857 , \30534 );
not \U$30863 ( \30858 , \30857 );
or \U$30864 ( \30859 , \30856 , \30858 );
buf \U$30865 ( \30860 , \30371 );
not \U$30866 ( \30861 , \30860 );
buf \U$30867 ( \30862 , \30534 );
not \U$30868 ( \30863 , \30862 );
buf \U$30869 ( \30864 , \30863 );
buf \U$30870 ( \30865 , \30864 );
not \U$30871 ( \30866 , \30865 );
or \U$30872 ( \30867 , \30861 , \30866 );
buf \U$30873 ( \30868 , \30584 );
nand \U$30874 ( \30869 , \30867 , \30868 );
buf \U$30875 ( \30870 , \30869 );
buf \U$30876 ( \30871 , \30870 );
nand \U$30877 ( \30872 , \30859 , \30871 );
buf \U$30878 ( \30873 , \30872 );
buf \U$30879 ( \30874 , \30729 );
not \U$30880 ( \30875 , \30874 );
buf \U$30881 ( \30876 , \30662 );
not \U$30882 ( \30877 , \30876 );
or \U$30883 ( \30878 , \30875 , \30877 );
buf \U$30884 ( \30879 , \30732 );
not \U$30885 ( \30880 , \30879 );
buf \U$30886 ( \30881 , \30662 );
not \U$30887 ( \30882 , \30881 );
buf \U$30888 ( \30883 , \30882 );
buf \U$30889 ( \30884 , \30883 );
not \U$30890 ( \30885 , \30884 );
or \U$30891 ( \30886 , \30880 , \30885 );
buf \U$30892 ( \30887 , \30801 );
nand \U$30893 ( \30888 , \30886 , \30887 );
buf \U$30894 ( \30889 , \30888 );
buf \U$30895 ( \30890 , \30889 );
nand \U$30896 ( \30891 , \30878 , \30890 );
buf \U$30897 ( \30892 , \30891 );
xor \U$30898 ( \30893 , \30873 , \30892 );
and \U$30899 ( \30894 , \27395 , \27396 );
buf \U$30900 ( \30895 , \30894 );
buf \U$30901 ( \30896 , \30895 );
buf \U$30902 ( \30897 , \4904 );
buf \U$30903 ( \30898 , RIc0d8e60_52);
buf \U$30904 ( \30899 , RIc0d9568_67);
xor \U$30905 ( \30900 , \30898 , \30899 );
buf \U$30906 ( \30901 , \30900 );
buf \U$30907 ( \30902 , \30901 );
not \U$30908 ( \30903 , \30902 );
buf \U$30909 ( \30904 , \30903 );
buf \U$30910 ( \30905 , \30904 );
or \U$30911 ( \30906 , \30897 , \30905 );
buf \U$30912 ( \30907 , \685 );
xor \U$30913 ( \30908 , RIc0d9568_67, RIc0d8de8_51);
buf \U$30914 ( \30909 , \30908 );
nand \U$30915 ( \30910 , \30907 , \30909 );
buf \U$30916 ( \30911 , \30910 );
buf \U$30917 ( \30912 , \30911 );
nand \U$30918 ( \30913 , \30906 , \30912 );
buf \U$30919 ( \30914 , \30913 );
buf \U$30920 ( \30915 , \30914 );
xor \U$30921 ( \30916 , \30896 , \30915 );
buf \U$30922 ( \30917 , \16399 );
buf \U$30923 ( \30918 , RIc0d8320_28);
buf \U$30924 ( \30919 , RIc0da0a8_91);
xnor \U$30925 ( \30920 , \30918 , \30919 );
buf \U$30926 ( \30921 , \30920 );
buf \U$30927 ( \30922 , \30921 );
or \U$30928 ( \30923 , \30917 , \30922 );
buf \U$30929 ( \30924 , \530 );
buf \U$30930 ( \30925 , RIc0d82a8_27);
buf \U$30931 ( \30926 , RIc0da0a8_91);
xnor \U$30932 ( \30927 , \30925 , \30926 );
buf \U$30933 ( \30928 , \30927 );
buf \U$30934 ( \30929 , \30928 );
or \U$30935 ( \30930 , \30924 , \30929 );
nand \U$30936 ( \30931 , \30923 , \30930 );
buf \U$30937 ( \30932 , \30931 );
buf \U$30938 ( \30933 , \30932 );
and \U$30939 ( \30934 , \30916 , \30933 );
and \U$30940 ( \30935 , \30896 , \30915 );
or \U$30941 ( \30936 , \30934 , \30935 );
buf \U$30942 ( \30937 , \30936 );
buf \U$30943 ( \30938 , \30937 );
buf \U$30944 ( \30939 , \29321 );
not \U$30945 ( \30940 , \30939 );
buf \U$30946 ( \30941 , \23253 );
not \U$30947 ( \30942 , \30941 );
or \U$30948 ( \30943 , \30940 , \30942 );
buf \U$30949 ( \30944 , \1229 );
xor \U$30950 ( \30945 , \27995 , \27996 );
buf \U$30951 ( \30946 , \30945 );
buf \U$30952 ( \30947 , \30946 );
nand \U$30953 ( \30948 , \30944 , \30947 );
buf \U$30954 ( \30949 , \30948 );
buf \U$30955 ( \30950 , \30949 );
nand \U$30956 ( \30951 , \30943 , \30950 );
buf \U$30957 ( \30952 , \30951 );
buf \U$30958 ( \30953 , \30952 );
buf \U$30959 ( \30954 , \29366 );
not \U$30960 ( \30955 , \30954 );
buf \U$30961 ( \30956 , \1888 );
not \U$30962 ( \30957 , \30956 );
or \U$30963 ( \30958 , \30955 , \30957 );
buf \U$30964 ( \30959 , \2927 );
buf \U$30965 ( \30960 , \29241 );
nand \U$30966 ( \30961 , \30959 , \30960 );
buf \U$30967 ( \30962 , \30961 );
buf \U$30968 ( \30963 , \30962 );
nand \U$30969 ( \30964 , \30958 , \30963 );
buf \U$30970 ( \30965 , \30964 );
buf \U$30971 ( \30966 , \30965 );
xor \U$30972 ( \30967 , \30953 , \30966 );
buf \U$30973 ( \30968 , \2938 );
buf \U$30974 ( \30969 , RIc0d8050_22);
buf \U$30975 ( \30970 , RIc0da378_97);
xnor \U$30976 ( \30971 , \30969 , \30970 );
buf \U$30977 ( \30972 , \30971 );
buf \U$30978 ( \30973 , \30972 );
or \U$30979 ( \30974 , \30968 , \30973 );
buf \U$30980 ( \30975 , \737 );
buf \U$30981 ( \30976 , \30396 );
not \U$30982 ( \30977 , \30976 );
buf \U$30983 ( \30978 , \30977 );
buf \U$30984 ( \30979 , \30978 );
or \U$30985 ( \30980 , \30975 , \30979 );
nand \U$30986 ( \30981 , \30974 , \30980 );
buf \U$30987 ( \30982 , \30981 );
buf \U$30988 ( \30983 , \30982 );
and \U$30989 ( \30984 , \30967 , \30983 );
and \U$30990 ( \30985 , \30953 , \30966 );
or \U$30991 ( \30986 , \30984 , \30985 );
buf \U$30992 ( \30987 , \30986 );
buf \U$30993 ( \30988 , \30987 );
xor \U$30994 ( \30989 , \30938 , \30988 );
buf \U$30995 ( \30990 , RIc0d86e0_36);
buf \U$30996 ( \30991 , RIc0d9ce8_83);
xor \U$30997 ( \30992 , \30990 , \30991 );
buf \U$30998 ( \30993 , \30992 );
buf \U$30999 ( \30994 , \30993 );
not \U$31000 ( \30995 , \30994 );
buf \U$31001 ( \30996 , \12254 );
not \U$31002 ( \30997 , \30996 );
or \U$31003 ( \30998 , \30995 , \30997 );
buf \U$31004 ( \30999 , \584 );
buf \U$31005 ( \31000 , \30418 );
nand \U$31006 ( \31001 , \30999 , \31000 );
buf \U$31007 ( \31002 , \31001 );
buf \U$31008 ( \31003 , \31002 );
nand \U$31009 ( \31004 , \30998 , \31003 );
buf \U$31010 ( \31005 , \31004 );
buf \U$31011 ( \31006 , \31005 );
buf \U$31012 ( \31007 , RIc0d8d70_50);
buf \U$31013 ( \31008 , RIc0d9658_69);
xor \U$31014 ( \31009 , \31007 , \31008 );
buf \U$31015 ( \31010 , \31009 );
buf \U$31016 ( \31011 , \31010 );
not \U$31017 ( \31012 , \31011 );
buf \U$31018 ( \31013 , \279 );
not \U$31019 ( \31014 , \31013 );
or \U$31020 ( \31015 , \31012 , \31014 );
buf \U$31021 ( \31016 , \874 );
buf \U$31022 ( \31017 , \27875 );
nand \U$31023 ( \31018 , \31016 , \31017 );
buf \U$31024 ( \31019 , \31018 );
buf \U$31025 ( \31020 , \31019 );
nand \U$31026 ( \31021 , \31015 , \31020 );
buf \U$31027 ( \31022 , \31021 );
buf \U$31028 ( \31023 , \31022 );
xor \U$31029 ( \31024 , \31006 , \31023 );
buf \U$31030 ( \31025 , RIc0da828_107);
buf \U$31031 ( \31026 , RIc0d7ba0_12);
xor \U$31032 ( \31027 , \31025 , \31026 );
buf \U$31033 ( \31028 , \31027 );
buf \U$31034 ( \31029 , \31028 );
not \U$31035 ( \31030 , \31029 );
buf \U$31036 ( \31031 , \21898 );
not \U$31037 ( \31032 , \31031 );
or \U$31038 ( \31033 , \31030 , \31032 );
buf \U$31039 ( \31034 , \12342 );
xor \U$31040 ( \31035 , RIc0da828_107, RIc0d7b28_11);
buf \U$31041 ( \31036 , \31035 );
nand \U$31042 ( \31037 , \31034 , \31036 );
buf \U$31043 ( \31038 , \31037 );
buf \U$31044 ( \31039 , \31038 );
nand \U$31045 ( \31040 , \31033 , \31039 );
buf \U$31046 ( \31041 , \31040 );
buf \U$31047 ( \31042 , \31041 );
and \U$31048 ( \31043 , \31024 , \31042 );
and \U$31049 ( \31044 , \31006 , \31023 );
or \U$31050 ( \31045 , \31043 , \31044 );
buf \U$31051 ( \31046 , \31045 );
buf \U$31052 ( \31047 , \31046 );
and \U$31053 ( \31048 , \30989 , \31047 );
and \U$31054 ( \31049 , \30938 , \30988 );
or \U$31055 ( \31050 , \31048 , \31049 );
buf \U$31056 ( \31051 , \31050 );
xor \U$31057 ( \31052 , \30893 , \31051 );
buf \U$31058 ( \31053 , \31052 );
and \U$31059 ( \31054 , \30854 , \31053 );
and \U$31060 ( \31055 , \30471 , \30853 );
or \U$31061 ( \31056 , \31054 , \31055 );
buf \U$31062 ( \31057 , \31056 );
buf \U$31063 ( \31058 , \31051 );
buf \U$31064 ( \31059 , \30873 );
or \U$31065 ( \31060 , \31058 , \31059 );
buf \U$31066 ( \31061 , \30892 );
nand \U$31067 ( \31062 , \31060 , \31061 );
buf \U$31068 ( \31063 , \31062 );
buf \U$31069 ( \31064 , \30873 );
buf \U$31070 ( \31065 , \31051 );
nand \U$31071 ( \31066 , \31064 , \31065 );
buf \U$31072 ( \31067 , \31066 );
and \U$31073 ( \31068 , \31063 , \31067 );
buf \U$31074 ( \31069 , \31068 );
not \U$31075 ( \31070 , \31069 );
buf \U$31076 ( \31071 , \30454 );
not \U$31077 ( \31072 , \31071 );
buf \U$31078 ( \31073 , \30441 );
not \U$31079 ( \31074 , \31073 );
or \U$31080 ( \31075 , \31072 , \31074 );
buf \U$31081 ( \31076 , \30441 );
buf \U$31082 ( \31077 , \30454 );
or \U$31083 ( \31078 , \31076 , \31077 );
buf \U$31084 ( \31079 , \30449 );
not \U$31085 ( \31080 , \31079 );
buf \U$31086 ( \31081 , \31080 );
buf \U$31087 ( \31082 , \31081 );
nand \U$31088 ( \31083 , \31078 , \31082 );
buf \U$31089 ( \31084 , \31083 );
buf \U$31090 ( \31085 , \31084 );
nand \U$31091 ( \31086 , \31075 , \31085 );
buf \U$31092 ( \31087 , \31086 );
buf \U$31093 ( \31088 , \31087 );
not \U$31094 ( \31089 , \31088 );
and \U$31095 ( \31090 , \31070 , \31089 );
buf \U$31096 ( \31091 , \31087 );
buf \U$31097 ( \31092 , \31068 );
and \U$31098 ( \31093 , \31091 , \31092 );
nor \U$31099 ( \31094 , \31090 , \31093 );
buf \U$31100 ( \31095 , \31094 );
buf \U$31101 ( \31096 , \31095 );
buf \U$31102 ( \31097 , \30908 );
not \U$31103 ( \31098 , \31097 );
buf \U$31104 ( \31099 , \1822 );
not \U$31105 ( \31100 , \31099 );
or \U$31106 ( \31101 , \31098 , \31100 );
buf \U$31107 ( \31102 , \686 );
buf \U$31108 ( \31103 , \28003 );
nand \U$31109 ( \31104 , \31102 , \31103 );
buf \U$31110 ( \31105 , \31104 );
buf \U$31111 ( \31106 , \31105 );
nand \U$31112 ( \31107 , \31101 , \31106 );
buf \U$31113 ( \31108 , \31107 );
buf \U$31114 ( \31109 , \31108 );
buf \U$31115 ( \31110 , \30628 );
not \U$31116 ( \31111 , \31110 );
buf \U$31117 ( \31112 , \18057 );
not \U$31118 ( \31113 , \31112 );
or \U$31119 ( \31114 , \31111 , \31113 );
buf \U$31120 ( \31115 , \791 );
buf \U$31121 ( \31116 , \28199 );
nand \U$31122 ( \31117 , \31115 , \31116 );
buf \U$31123 ( \31118 , \31117 );
buf \U$31124 ( \31119 , \31118 );
nand \U$31125 ( \31120 , \31114 , \31119 );
buf \U$31126 ( \31121 , \31120 );
buf \U$31127 ( \31122 , \31121 );
xor \U$31128 ( \31123 , \31109 , \31122 );
buf \U$31129 ( \31124 , \12331 );
buf \U$31130 ( \31125 , \31035 );
not \U$31131 ( \31126 , \31125 );
buf \U$31132 ( \31127 , \31126 );
buf \U$31133 ( \31128 , \31127 );
or \U$31134 ( \31129 , \31124 , \31128 );
buf \U$31135 ( \31130 , \16064 );
buf \U$31136 ( \31131 , \28084 );
or \U$31137 ( \31132 , \31130 , \31131 );
nand \U$31138 ( \31133 , \31129 , \31132 );
buf \U$31139 ( \31134 , \31133 );
buf \U$31140 ( \31135 , \31134 );
and \U$31141 ( \31136 , \31123 , \31135 );
and \U$31142 ( \31137 , \31109 , \31122 );
or \U$31143 ( \31138 , \31136 , \31137 );
buf \U$31144 ( \31139 , \31138 );
buf \U$31145 ( \31140 , \31139 );
not \U$31146 ( \31141 , \31140 );
buf \U$31147 ( \31142 , \30606 );
not \U$31148 ( \31143 , \31142 );
buf \U$31149 ( \31144 , \2607 );
not \U$31150 ( \31145 , \31144 );
or \U$31151 ( \31146 , \31143 , \31145 );
buf \U$31152 ( \31147 , \816 );
buf \U$31153 ( \31148 , \28227 );
nand \U$31154 ( \31149 , \31147 , \31148 );
buf \U$31155 ( \31150 , \31149 );
buf \U$31156 ( \31151 , \31150 );
nand \U$31157 ( \31152 , \31146 , \31151 );
buf \U$31158 ( \31153 , \31152 );
buf \U$31159 ( \31154 , \31153 );
buf \U$31160 ( \31155 , \30763 );
not \U$31161 ( \31156 , \31155 );
buf \U$31162 ( \31157 , \3384 );
not \U$31163 ( \31158 , \31157 );
or \U$31164 ( \31159 , \31156 , \31158 );
buf \U$31165 ( \31160 , \846 );
buf \U$31166 ( \31161 , \28478 );
nand \U$31167 ( \31162 , \31160 , \31161 );
buf \U$31168 ( \31163 , \31162 );
buf \U$31169 ( \31164 , \31163 );
nand \U$31170 ( \31165 , \31159 , \31164 );
buf \U$31171 ( \31166 , \31165 );
buf \U$31172 ( \31167 , \31166 );
or \U$31173 ( \31168 , \31154 , \31167 );
buf \U$31174 ( \31169 , \30928 );
not \U$31175 ( \31170 , \31169 );
buf \U$31176 ( \31171 , \31170 );
buf \U$31177 ( \31172 , \31171 );
not \U$31178 ( \31173 , \31172 );
buf \U$31179 ( \31174 , \1927 );
not \U$31180 ( \31175 , \31174 );
or \U$31181 ( \31176 , \31173 , \31175 );
buf \U$31182 ( \31177 , \1933 );
buf \U$31183 ( \31178 , \28022 );
nand \U$31184 ( \31179 , \31177 , \31178 );
buf \U$31185 ( \31180 , \31179 );
buf \U$31186 ( \31181 , \31180 );
nand \U$31187 ( \31182 , \31176 , \31181 );
buf \U$31188 ( \31183 , \31182 );
buf \U$31189 ( \31184 , \31183 );
nand \U$31190 ( \31185 , \31168 , \31184 );
buf \U$31191 ( \31186 , \31185 );
buf \U$31192 ( \31187 , \31186 );
buf \U$31193 ( \31188 , \31153 );
buf \U$31194 ( \31189 , \31166 );
nand \U$31195 ( \31190 , \31188 , \31189 );
buf \U$31196 ( \31191 , \31190 );
buf \U$31197 ( \31192 , \31191 );
nand \U$31198 ( \31193 , \31187 , \31192 );
buf \U$31199 ( \31194 , \31193 );
buf \U$31200 ( \31195 , \31194 );
not \U$31201 ( \31196 , \31195 );
buf \U$31202 ( \31197 , \31196 );
buf \U$31203 ( \31198 , \31197 );
not \U$31204 ( \31199 , \31198 );
or \U$31205 ( \31200 , \31141 , \31199 );
buf \U$31206 ( \31201 , \31197 );
buf \U$31207 ( \31202 , \31139 );
or \U$31208 ( \31203 , \31201 , \31202 );
nand \U$31209 ( \31204 , \31200 , \31203 );
buf \U$31210 ( \31205 , \31204 );
buf \U$31211 ( \31206 , \31205 );
and \U$31212 ( \31207 , \29318 , \29319 );
buf \U$31213 ( \31208 , \31207 );
buf \U$31214 ( \31209 , \31208 );
buf \U$31215 ( \31210 , \30741 );
not \U$31216 ( \31211 , \31210 );
buf \U$31217 ( \31212 , \13860 );
not \U$31218 ( \31213 , \31212 );
or \U$31219 ( \31214 , \31211 , \31213 );
buf \U$31220 ( \31215 , \343 );
buf \U$31221 ( \31216 , \28496 );
nand \U$31222 ( \31217 , \31215 , \31216 );
buf \U$31223 ( \31218 , \31217 );
buf \U$31224 ( \31219 , \31218 );
nand \U$31225 ( \31220 , \31214 , \31219 );
buf \U$31226 ( \31221 , \31220 );
buf \U$31227 ( \31222 , \31221 );
xor \U$31228 ( \31223 , \31209 , \31222 );
buf \U$31229 ( \31224 , \4483 );
buf \U$31230 ( \31225 , \30789 );
not \U$31231 ( \31226 , \31225 );
buf \U$31232 ( \31227 , \31226 );
buf \U$31233 ( \31228 , \31227 );
or \U$31234 ( \31229 , \31224 , \31228 );
buf \U$31235 ( \31230 , \4475 );
buf \U$31236 ( \31231 , \28518 );
or \U$31237 ( \31232 , \31230 , \31231 );
nand \U$31238 ( \31233 , \31229 , \31232 );
buf \U$31239 ( \31234 , \31233 );
buf \U$31240 ( \31235 , \31234 );
and \U$31241 ( \31236 , \31223 , \31235 );
and \U$31242 ( \31237 , \31209 , \31222 );
or \U$31243 ( \31238 , \31236 , \31237 );
buf \U$31244 ( \31239 , \31238 );
buf \U$31245 ( \31240 , \31239 );
and \U$31246 ( \31241 , \31206 , \31240 );
not \U$31247 ( \31242 , \31206 );
buf \U$31248 ( \31243 , \31239 );
not \U$31249 ( \31244 , \31243 );
buf \U$31250 ( \31245 , \31244 );
buf \U$31251 ( \31246 , \31245 );
and \U$31252 ( \31247 , \31242 , \31246 );
nor \U$31253 ( \31248 , \31241 , \31247 );
buf \U$31254 ( \31249 , \31248 );
buf \U$31255 ( \31250 , \31249 );
xor \U$31256 ( \31251 , \31153 , \31183 );
buf \U$31257 ( \31252 , \31251 );
buf \U$31258 ( \31253 , \31166 );
and \U$31259 ( \31254 , \31252 , \31253 );
not \U$31260 ( \31255 , \31252 );
buf \U$31261 ( \31256 , \31166 );
not \U$31262 ( \31257 , \31256 );
buf \U$31263 ( \31258 , \31257 );
buf \U$31264 ( \31259 , \31258 );
and \U$31265 ( \31260 , \31255 , \31259 );
nor \U$31266 ( \31261 , \31254 , \31260 );
buf \U$31267 ( \31262 , \31261 );
buf \U$31268 ( \31263 , \31262 );
not \U$31269 ( \31264 , \31263 );
buf \U$31270 ( \31265 , \27870 );
not \U$31271 ( \31266 , \31265 );
buf \U$31272 ( \31267 , \31266 );
and \U$31273 ( \31268 , \27891 , \31267 );
not \U$31274 ( \31269 , \27891 );
and \U$31275 ( \31270 , \31269 , \27870 );
or \U$31276 ( \31271 , \31268 , \31270 );
and \U$31277 ( \31272 , \31271 , \27916 );
not \U$31278 ( \31273 , \31271 );
buf \U$31279 ( \31274 , \27916 );
not \U$31280 ( \31275 , \31274 );
buf \U$31281 ( \31276 , \31275 );
and \U$31282 ( \31277 , \31273 , \31276 );
nor \U$31283 ( \31278 , \31272 , \31277 );
buf \U$31284 ( \31279 , \31278 );
not \U$31285 ( \31280 , \31279 );
or \U$31286 ( \31281 , \31264 , \31280 );
buf \U$31287 ( \31282 , \31278 );
buf \U$31288 ( \31283 , \31262 );
or \U$31289 ( \31284 , \31282 , \31283 );
xor \U$31290 ( \31285 , \30408 , \30391 );
buf \U$31291 ( \31286 , \31285 );
buf \U$31292 ( \31287 , \30431 );
and \U$31293 ( \31288 , \31286 , \31287 );
not \U$31294 ( \31289 , \31286 );
buf \U$31295 ( \31290 , \30431 );
not \U$31296 ( \31291 , \31290 );
buf \U$31297 ( \31292 , \31291 );
buf \U$31298 ( \31293 , \31292 );
and \U$31299 ( \31294 , \31289 , \31293 );
nor \U$31300 ( \31295 , \31288 , \31294 );
buf \U$31301 ( \31296 , \31295 );
buf \U$31302 ( \31297 , \31296 );
not \U$31303 ( \31298 , \31297 );
buf \U$31304 ( \31299 , \31298 );
buf \U$31305 ( \31300 , \31299 );
nand \U$31306 ( \31301 , \31284 , \31300 );
buf \U$31307 ( \31302 , \31301 );
buf \U$31308 ( \31303 , \31302 );
nand \U$31309 ( \31304 , \31281 , \31303 );
buf \U$31310 ( \31305 , \31304 );
buf \U$31311 ( \31306 , \31305 );
or \U$31312 ( \31307 , \31250 , \31306 );
buf \U$31313 ( \31308 , \30946 );
not \U$31314 ( \31309 , \31308 );
buf \U$31315 ( \31310 , \23253 );
not \U$31316 ( \31311 , \31310 );
or \U$31317 ( \31312 , \31309 , \31311 );
buf \U$31318 ( \31313 , \1229 );
buf \U$31319 ( \31314 , \28111 );
nand \U$31320 ( \31315 , \31313 , \31314 );
buf \U$31321 ( \31316 , \31315 );
buf \U$31322 ( \31317 , \31316 );
nand \U$31323 ( \31318 , \31312 , \31317 );
buf \U$31324 ( \31319 , \31318 );
buf \U$31325 ( \31320 , \31319 );
not \U$31326 ( \31321 , \31320 );
buf \U$31327 ( \31322 , RIc0d9b08_79);
buf \U$31328 ( \31323 , RIc0d8848_39);
xor \U$31329 ( \31324 , \31322 , \31323 );
buf \U$31330 ( \31325 , \31324 );
buf \U$31331 ( \31326 , \31325 );
not \U$31332 ( \31327 , \31326 );
buf \U$31333 ( \31328 , \4509 );
not \U$31334 ( \31329 , \31328 );
or \U$31335 ( \31330 , \31327 , \31329 );
buf \U$31336 ( \31331 , \1025 );
buf \U$31337 ( \31332 , \28304 );
nand \U$31338 ( \31333 , \31331 , \31332 );
buf \U$31339 ( \31334 , \31333 );
buf \U$31340 ( \31335 , \31334 );
nand \U$31341 ( \31336 , \31330 , \31335 );
buf \U$31342 ( \31337 , \31336 );
buf \U$31343 ( \31338 , \31337 );
not \U$31344 ( \31339 , \31338 );
or \U$31345 ( \31340 , \31321 , \31339 );
buf \U$31346 ( \31341 , \31337 );
buf \U$31347 ( \31342 , \31319 );
or \U$31348 ( \31343 , \31341 , \31342 );
buf \U$31349 ( \31344 , RIc0d81b8_25);
buf \U$31350 ( \31345 , RIc0da198_93);
xor \U$31351 ( \31346 , \31344 , \31345 );
buf \U$31352 ( \31347 , \31346 );
buf \U$31353 ( \31348 , \31347 );
not \U$31354 ( \31349 , \31348 );
buf \U$31355 ( \31350 , \15995 );
not \U$31356 ( \31351 , \31350 );
or \U$31357 ( \31352 , \31349 , \31351 );
buf \U$31358 ( \31353 , \481 );
buf \U$31359 ( \31354 , \28270 );
nand \U$31360 ( \31355 , \31353 , \31354 );
buf \U$31361 ( \31356 , \31355 );
buf \U$31362 ( \31357 , \31356 );
nand \U$31363 ( \31358 , \31352 , \31357 );
buf \U$31364 ( \31359 , \31358 );
buf \U$31365 ( \31360 , \31359 );
nand \U$31366 ( \31361 , \31343 , \31360 );
buf \U$31367 ( \31362 , \31361 );
buf \U$31368 ( \31363 , \31362 );
nand \U$31369 ( \31364 , \31340 , \31363 );
buf \U$31370 ( \31365 , \31364 );
buf \U$31371 ( \31366 , \29244 );
not \U$31372 ( \31367 , \31366 );
buf \U$31373 ( \31368 , \29267 );
not \U$31374 ( \31369 , \31368 );
or \U$31375 ( \31370 , \31367 , \31369 );
buf \U$31376 ( \31371 , \29284 );
nand \U$31377 ( \31372 , \31370 , \31371 );
buf \U$31378 ( \31373 , \31372 );
buf \U$31379 ( \31374 , \31373 );
buf \U$31380 ( \31375 , \29244 );
not \U$31381 ( \31376 , \31375 );
buf \U$31382 ( \31377 , \29264 );
nand \U$31383 ( \31378 , \31376 , \31377 );
buf \U$31384 ( \31379 , \31378 );
buf \U$31385 ( \31380 , \31379 );
nand \U$31386 ( \31381 , \31374 , \31380 );
buf \U$31387 ( \31382 , \31381 );
xor \U$31388 ( \31383 , \31365 , \31382 );
buf \U$31389 ( \31384 , \30546 );
not \U$31390 ( \31385 , \31384 );
buf \U$31391 ( \31386 , \13737 );
not \U$31392 ( \31387 , \31386 );
or \U$31393 ( \31388 , \31385 , \31387 );
buf \U$31394 ( \31389 , \1401 );
buf \U$31395 ( \31390 , \28559 );
nand \U$31396 ( \31391 , \31389 , \31390 );
buf \U$31397 ( \31392 , \31391 );
buf \U$31398 ( \31393 , \31392 );
nand \U$31399 ( \31394 , \31388 , \31393 );
buf \U$31400 ( \31395 , \31394 );
buf \U$31401 ( \31396 , \31395 );
buf \U$31402 ( \31397 , \30650 );
not \U$31403 ( \31398 , \31397 );
buf \U$31404 ( \31399 , \3534 );
not \U$31405 ( \31400 , \31399 );
or \U$31406 ( \31401 , \31398 , \31400 );
buf \U$31407 ( \31402 , \16676 );
buf \U$31408 ( \31403 , \28179 );
nand \U$31409 ( \31404 , \31402 , \31403 );
buf \U$31410 ( \31405 , \31404 );
buf \U$31411 ( \31406 , \31405 );
nand \U$31412 ( \31407 , \31401 , \31406 );
buf \U$31413 ( \31408 , \31407 );
buf \U$31414 ( \31409 , \31408 );
xor \U$31415 ( \31410 , \31396 , \31409 );
buf \U$31416 ( \31411 , \30482 );
not \U$31417 ( \31412 , \31411 );
buf \U$31418 ( \31413 , \25355 );
not \U$31419 ( \31414 , \31413 );
or \U$31420 ( \31415 , \31412 , \31414 );
buf \U$31421 ( \31416 , \14405 );
buf \U$31422 ( \31417 , \28408 );
nand \U$31423 ( \31418 , \31416 , \31417 );
buf \U$31424 ( \31419 , \31418 );
buf \U$31425 ( \31420 , \31419 );
nand \U$31426 ( \31421 , \31415 , \31420 );
buf \U$31427 ( \31422 , \31421 );
buf \U$31428 ( \31423 , \31422 );
and \U$31429 ( \31424 , \31410 , \31423 );
and \U$31430 ( \31425 , \31396 , \31409 );
or \U$31431 ( \31426 , \31424 , \31425 );
buf \U$31432 ( \31427 , \31426 );
xnor \U$31433 ( \31428 , \31383 , \31427 );
buf \U$31434 ( \31429 , \31428 );
not \U$31435 ( \31430 , \31429 );
buf \U$31436 ( \31431 , \31430 );
buf \U$31437 ( \31432 , \31431 );
nand \U$31438 ( \31433 , \31307 , \31432 );
buf \U$31439 ( \31434 , \31433 );
buf \U$31440 ( \31435 , \31434 );
buf \U$31441 ( \31436 , \31249 );
buf \U$31442 ( \31437 , \31305 );
nand \U$31443 ( \31438 , \31436 , \31437 );
buf \U$31444 ( \31439 , \31438 );
buf \U$31445 ( \31440 , \31439 );
nand \U$31446 ( \31441 , \31435 , \31440 );
buf \U$31447 ( \31442 , \31441 );
buf \U$31448 ( \31443 , \31442 );
and \U$31449 ( \31444 , \31096 , \31443 );
not \U$31450 ( \31445 , \31096 );
buf \U$31451 ( \31446 , \31442 );
not \U$31452 ( \31447 , \31446 );
buf \U$31453 ( \31448 , \31447 );
buf \U$31454 ( \31449 , \31448 );
and \U$31455 ( \31450 , \31445 , \31449 );
nor \U$31456 ( \31451 , \31444 , \31450 );
buf \U$31457 ( \31452 , \31451 );
xor \U$31458 ( \31453 , \31057 , \31452 );
xor \U$31459 ( \31454 , \27921 , \27993 );
xor \U$31460 ( \31455 , \31454 , \28039 );
buf \U$31461 ( \31456 , \31455 );
buf \U$31462 ( \31457 , \31456 );
not \U$31463 ( \31458 , \31457 );
buf \U$31464 ( \31459 , \31319 );
buf \U$31465 ( \31460 , \31359 );
xor \U$31466 ( \31461 , \31459 , \31460 );
buf \U$31467 ( \31462 , \31337 );
xnor \U$31468 ( \31463 , \31461 , \31462 );
buf \U$31469 ( \31464 , \31463 );
buf \U$31470 ( \31465 , \31464 );
not \U$31471 ( \31466 , \31465 );
xor \U$31472 ( \31467 , \27986 , \27960 );
buf \U$31473 ( \31468 , \31467 );
buf \U$31474 ( \31469 , \27938 );
not \U$31475 ( \31470 , \31469 );
buf \U$31476 ( \31471 , \31470 );
buf \U$31477 ( \31472 , \31471 );
and \U$31478 ( \31473 , \31468 , \31472 );
not \U$31479 ( \31474 , \31468 );
buf \U$31480 ( \31475 , \27938 );
and \U$31481 ( \31476 , \31474 , \31475 );
nor \U$31482 ( \31477 , \31473 , \31476 );
buf \U$31483 ( \31478 , \31477 );
buf \U$31484 ( \31479 , \31478 );
not \U$31485 ( \31480 , \31479 );
or \U$31486 ( \31481 , \31466 , \31480 );
xor \U$31487 ( \31482 , \31396 , \31409 );
xor \U$31488 ( \31483 , \31482 , \31423 );
buf \U$31489 ( \31484 , \31483 );
buf \U$31490 ( \31485 , \31484 );
nand \U$31491 ( \31486 , \31481 , \31485 );
buf \U$31492 ( \31487 , \31486 );
buf \U$31493 ( \31488 , \31487 );
buf \U$31494 ( \31489 , \31478 );
not \U$31495 ( \31490 , \31489 );
buf \U$31496 ( \31491 , \31464 );
not \U$31497 ( \31492 , \31491 );
buf \U$31498 ( \31493 , \31492 );
buf \U$31499 ( \31494 , \31493 );
nand \U$31500 ( \31495 , \31490 , \31494 );
buf \U$31501 ( \31496 , \31495 );
buf \U$31502 ( \31497 , \31496 );
nand \U$31503 ( \31498 , \31488 , \31497 );
buf \U$31504 ( \31499 , \31498 );
buf \U$31505 ( \31500 , \31499 );
not \U$31506 ( \31501 , \31500 );
buf \U$31507 ( \31502 , \31501 );
buf \U$31508 ( \31503 , \31502 );
not \U$31509 ( \31504 , \31503 );
or \U$31510 ( \31505 , \31458 , \31504 );
buf \U$31511 ( \31506 , \31502 );
buf \U$31512 ( \31507 , \31456 );
or \U$31513 ( \31508 , \31506 , \31507 );
nand \U$31514 ( \31509 , \31505 , \31508 );
buf \U$31515 ( \31510 , \31509 );
buf \U$31516 ( \31511 , \31510 );
buf \U$31517 ( \31512 , \29302 );
not \U$31518 ( \31513 , \31512 );
buf \U$31519 ( \31514 , \396 );
not \U$31520 ( \31515 , \31514 );
or \U$31521 ( \31516 , \31513 , \31515 );
buf \U$31522 ( \31517 , \1025 );
buf \U$31523 ( \31518 , \31325 );
nand \U$31524 ( \31519 , \31517 , \31518 );
buf \U$31525 ( \31520 , \31519 );
buf \U$31526 ( \31521 , \31520 );
nand \U$31527 ( \31522 , \31516 , \31521 );
buf \U$31528 ( \31523 , \31522 );
buf \U$31529 ( \31524 , \31523 );
buf \U$31530 ( \31525 , \29346 );
not \U$31531 ( \31526 , \31525 );
buf \U$31532 ( \31527 , \13419 );
not \U$31533 ( \31528 , \31527 );
or \U$31534 ( \31529 , \31526 , \31528 );
buf \U$31535 ( \31530 , \13426 );
buf \U$31536 ( \31531 , \30379 );
nand \U$31537 ( \31532 , \31530 , \31531 );
buf \U$31538 ( \31533 , \31532 );
buf \U$31539 ( \31534 , \31533 );
nand \U$31540 ( \31535 , \31529 , \31534 );
buf \U$31541 ( \31536 , \31535 );
buf \U$31542 ( \31537 , \31536 );
nor \U$31543 ( \31538 , \31524 , \31537 );
buf \U$31544 ( \31539 , \31538 );
buf \U$31545 ( \31540 , \31539 );
buf \U$31546 ( \31541 , RIc0d8230_26);
buf \U$31547 ( \31542 , RIc0da198_93);
xor \U$31548 ( \31543 , \31541 , \31542 );
buf \U$31549 ( \31544 , \31543 );
buf \U$31550 ( \31545 , \31544 );
not \U$31551 ( \31546 , \31545 );
buf \U$31552 ( \31547 , \889 );
not \U$31553 ( \31548 , \31547 );
or \U$31554 ( \31549 , \31546 , \31548 );
buf \U$31555 ( \31550 , \481 );
buf \U$31556 ( \31551 , \31347 );
nand \U$31557 ( \31552 , \31550 , \31551 );
buf \U$31558 ( \31553 , \31552 );
buf \U$31559 ( \31554 , \31553 );
nand \U$31560 ( \31555 , \31549 , \31554 );
buf \U$31561 ( \31556 , \31555 );
buf \U$31562 ( \31557 , \31556 );
not \U$31563 ( \31558 , \31557 );
buf \U$31564 ( \31559 , \31558 );
buf \U$31565 ( \31560 , \31559 );
or \U$31566 ( \31561 , \31540 , \31560 );
buf \U$31567 ( \31562 , \31523 );
buf \U$31568 ( \31563 , \31536 );
nand \U$31569 ( \31564 , \31562 , \31563 );
buf \U$31570 ( \31565 , \31564 );
buf \U$31571 ( \31566 , \31565 );
nand \U$31572 ( \31567 , \31561 , \31566 );
buf \U$31573 ( \31568 , \31567 );
buf \U$31574 ( \31569 , \31568 );
xor \U$31575 ( \31570 , \31109 , \31122 );
xor \U$31576 ( \31571 , \31570 , \31135 );
buf \U$31577 ( \31572 , \31571 );
buf \U$31578 ( \31573 , \31572 );
xor \U$31579 ( \31574 , \31569 , \31573 );
xor \U$31580 ( \31575 , \31209 , \31222 );
xor \U$31581 ( \31576 , \31575 , \31235 );
buf \U$31582 ( \31577 , \31576 );
buf \U$31583 ( \31578 , \31577 );
and \U$31584 ( \31579 , \31574 , \31578 );
and \U$31585 ( \31580 , \31569 , \31573 );
or \U$31586 ( \31581 , \31579 , \31580 );
buf \U$31587 ( \31582 , \31581 );
buf \U$31588 ( \31583 , \31582 );
not \U$31589 ( \31584 , \31583 );
buf \U$31590 ( \31585 , \31584 );
buf \U$31591 ( \31586 , \31585 );
and \U$31592 ( \31587 , \31511 , \31586 );
not \U$31593 ( \31588 , \31511 );
buf \U$31594 ( \31589 , \31582 );
and \U$31595 ( \31590 , \31588 , \31589 );
nor \U$31596 ( \31591 , \31587 , \31590 );
buf \U$31597 ( \31592 , \31591 );
buf \U$31598 ( \31593 , \31592 );
xor \U$31599 ( \31594 , \30938 , \30988 );
xor \U$31600 ( \31595 , \31594 , \31047 );
buf \U$31601 ( \31596 , \31595 );
buf \U$31602 ( \31597 , \31596 );
buf \U$31603 ( \31598 , \27581 );
not \U$31604 ( \31599 , \31598 );
buf \U$31605 ( \31600 , \2037 );
not \U$31606 ( \31601 , \31600 );
or \U$31607 ( \31602 , \31599 , \31601 );
buf \U$31608 ( \31603 , \441 );
buf \U$31609 ( \31604 , \30753 );
nand \U$31610 ( \31605 , \31603 , \31604 );
buf \U$31611 ( \31606 , \31605 );
buf \U$31612 ( \31607 , \31606 );
nand \U$31613 ( \31608 , \31602 , \31607 );
buf \U$31614 ( \31609 , \31608 );
buf \U$31615 ( \31610 , \31609 );
buf \U$31616 ( \31611 , \27699 );
not \U$31617 ( \31612 , \31611 );
buf \U$31618 ( \31613 , \2607 );
not \U$31619 ( \31614 , \31613 );
or \U$31620 ( \31615 , \31612 , \31614 );
buf \U$31621 ( \31616 , \816 );
buf \U$31622 ( \31617 , \30596 );
nand \U$31623 ( \31618 , \31616 , \31617 );
buf \U$31624 ( \31619 , \31618 );
buf \U$31625 ( \31620 , \31619 );
nand \U$31626 ( \31621 , \31615 , \31620 );
buf \U$31627 ( \31622 , \31621 );
buf \U$31628 ( \31623 , \31622 );
or \U$31629 ( \31624 , \31610 , \31623 );
buf \U$31630 ( \31625 , \27751 );
not \U$31631 ( \31626 , \31625 );
buf \U$31632 ( \31627 , \14186 );
not \U$31633 ( \31628 , \31627 );
or \U$31634 ( \31629 , \31626 , \31628 );
buf \U$31635 ( \31630 , \12303 );
buf \U$31636 ( \31631 , \30666 );
nand \U$31637 ( \31632 , \31630 , \31631 );
buf \U$31638 ( \31633 , \31632 );
buf \U$31639 ( \31634 , \31633 );
nand \U$31640 ( \31635 , \31629 , \31634 );
buf \U$31641 ( \31636 , \31635 );
buf \U$31642 ( \31637 , \31636 );
nand \U$31643 ( \31638 , \31624 , \31637 );
buf \U$31644 ( \31639 , \31638 );
buf \U$31645 ( \31640 , \31639 );
buf \U$31646 ( \31641 , \31622 );
buf \U$31647 ( \31642 , \31609 );
nand \U$31648 ( \31643 , \31641 , \31642 );
buf \U$31649 ( \31644 , \31643 );
buf \U$31650 ( \31645 , \31644 );
nand \U$31651 ( \31646 , \31640 , \31645 );
buf \U$31652 ( \31647 , \31646 );
buf \U$31653 ( \31648 , \31647 );
not \U$31654 ( \31649 , \31648 );
not \U$31655 ( \31650 , \686 );
not \U$31656 ( \31651 , \30901 );
or \U$31657 ( \31652 , \31650 , \31651 );
or \U$31658 ( \31653 , \8209 , \27357 );
nand \U$31659 ( \31654 , \31652 , \31653 );
buf \U$31660 ( \31655 , \31654 );
buf \U$31661 ( \31656 , \27729 );
not \U$31662 ( \31657 , \31656 );
buf \U$31663 ( \31658 , \2871 );
not \U$31664 ( \31659 , \31658 );
or \U$31665 ( \31660 , \31657 , \31659 );
buf \U$31666 ( \31661 , \791 );
buf \U$31667 ( \31662 , \30618 );
nand \U$31668 ( \31663 , \31661 , \31662 );
buf \U$31669 ( \31664 , \31663 );
buf \U$31670 ( \31665 , \31664 );
nand \U$31671 ( \31666 , \31660 , \31665 );
buf \U$31672 ( \31667 , \31666 );
buf \U$31673 ( \31668 , \31667 );
xor \U$31674 ( \31669 , \31655 , \31668 );
buf \U$31675 ( \31670 , \27377 );
not \U$31676 ( \31671 , \31670 );
buf \U$31677 ( \31672 , \2535 );
not \U$31678 ( \31673 , \31672 );
or \U$31679 ( \31674 , \31671 , \31673 );
buf \U$31680 ( \31675 , \30921 );
not \U$31681 ( \31676 , \31675 );
buf \U$31682 ( \31677 , \1933 );
nand \U$31683 ( \31678 , \31676 , \31677 );
buf \U$31684 ( \31679 , \31678 );
buf \U$31685 ( \31680 , \31679 );
nand \U$31686 ( \31681 , \31674 , \31680 );
buf \U$31687 ( \31682 , \31681 );
buf \U$31688 ( \31683 , \31682 );
and \U$31689 ( \31684 , \31669 , \31683 );
and \U$31690 ( \31685 , \31655 , \31668 );
or \U$31691 ( \31686 , \31684 , \31685 );
buf \U$31692 ( \31687 , \31686 );
buf \U$31693 ( \31688 , \31687 );
not \U$31694 ( \31689 , \31688 );
or \U$31695 ( \31690 , \31649 , \31689 );
buf \U$31696 ( \31691 , \31687 );
buf \U$31697 ( \31692 , \31647 );
or \U$31698 ( \31693 , \31691 , \31692 );
buf \U$31699 ( \31694 , \27681 );
not \U$31700 ( \31695 , \31694 );
buf \U$31701 ( \31696 , \15995 );
not \U$31702 ( \31697 , \31696 );
or \U$31703 ( \31698 , \31695 , \31697 );
buf \U$31704 ( \31699 , \4008 );
buf \U$31705 ( \31700 , \31544 );
nand \U$31706 ( \31701 , \31699 , \31700 );
buf \U$31707 ( \31702 , \31701 );
buf \U$31708 ( \31703 , \31702 );
nand \U$31709 ( \31704 , \31698 , \31703 );
buf \U$31710 ( \31705 , \31704 );
buf \U$31711 ( \31706 , \31705 );
not \U$31712 ( \31707 , \31706 );
buf \U$31713 ( \31708 , \27596 );
not \U$31714 ( \31709 , \31708 );
buf \U$31715 ( \31710 , \330 );
not \U$31716 ( \31711 , \31710 );
or \U$31717 ( \31712 , \31709 , \31711 );
buf \U$31718 ( \31713 , \343 );
buf \U$31719 ( \31714 , \30734 );
nand \U$31720 ( \31715 , \31713 , \31714 );
buf \U$31721 ( \31716 , \31715 );
buf \U$31722 ( \31717 , \31716 );
nand \U$31723 ( \31718 , \31712 , \31717 );
buf \U$31724 ( \31719 , \31718 );
buf \U$31725 ( \31720 , \31719 );
not \U$31726 ( \31721 , \31720 );
or \U$31727 ( \31722 , \31707 , \31721 );
buf \U$31728 ( \31723 , \31719 );
buf \U$31729 ( \31724 , \31705 );
or \U$31730 ( \31725 , \31723 , \31724 );
buf \U$31731 ( \31726 , \27615 );
not \U$31732 ( \31727 , \31726 );
buf \U$31733 ( \31728 , \16578 );
not \U$31734 ( \31729 , \31728 );
or \U$31735 ( \31730 , \31727 , \31729 );
buf \U$31736 ( \31731 , \15403 );
buf \U$31737 ( \31732 , \30779 );
nand \U$31738 ( \31733 , \31731 , \31732 );
buf \U$31739 ( \31734 , \31733 );
buf \U$31740 ( \31735 , \31734 );
nand \U$31741 ( \31736 , \31730 , \31735 );
buf \U$31742 ( \31737 , \31736 );
buf \U$31743 ( \31738 , \31737 );
nand \U$31744 ( \31739 , \31725 , \31738 );
buf \U$31745 ( \31740 , \31739 );
buf \U$31746 ( \31741 , \31740 );
nand \U$31747 ( \31742 , \31722 , \31741 );
buf \U$31748 ( \31743 , \31742 );
buf \U$31749 ( \31744 , \31743 );
nand \U$31750 ( \31745 , \31693 , \31744 );
buf \U$31751 ( \31746 , \31745 );
buf \U$31752 ( \31747 , \31746 );
nand \U$31753 ( \31748 , \31690 , \31747 );
buf \U$31754 ( \31749 , \31748 );
buf \U$31755 ( \31750 , \31749 );
xor \U$31756 ( \31751 , \31597 , \31750 );
buf \U$31757 ( \31752 , \27457 );
not \U$31758 ( \31753 , \31752 );
buf \U$31759 ( \31754 , \279 );
not \U$31760 ( \31755 , \31754 );
or \U$31761 ( \31756 , \31753 , \31755 );
buf \U$31762 ( \31757 , \874 );
buf \U$31763 ( \31758 , \31010 );
nand \U$31764 ( \31759 , \31757 , \31758 );
buf \U$31765 ( \31760 , \31759 );
buf \U$31766 ( \31761 , \31760 );
nand \U$31767 ( \31762 , \31756 , \31761 );
buf \U$31768 ( \31763 , \31762 );
buf \U$31769 ( \31764 , \31763 );
buf \U$31770 ( \31765 , \27788 );
not \U$31771 ( \31766 , \31765 );
buf \U$31772 ( \31767 , \1063 );
not \U$31773 ( \31768 , \31767 );
or \U$31774 ( \31769 , \31766 , \31768 );
buf \U$31775 ( \31770 , \1078 );
buf \U$31776 ( \31771 , \30687 );
nand \U$31777 ( \31772 , \31770 , \31771 );
buf \U$31778 ( \31773 , \31772 );
buf \U$31779 ( \31774 , \31773 );
nand \U$31780 ( \31775 , \31769 , \31774 );
buf \U$31781 ( \31776 , \31775 );
buf \U$31782 ( \31777 , \31776 );
xor \U$31783 ( \31778 , \31764 , \31777 );
buf \U$31784 ( \31779 , \27272 );
not \U$31785 ( \31780 , \31779 );
buf \U$31786 ( \31781 , \1183 );
not \U$31787 ( \31782 , \31781 );
or \U$31788 ( \31783 , \31780 , \31782 );
buf \U$31789 ( \31784 , \1588 );
buf \U$31790 ( \31785 , \30516 );
nand \U$31791 ( \31786 , \31784 , \31785 );
buf \U$31792 ( \31787 , \31786 );
buf \U$31793 ( \31788 , \31787 );
nand \U$31794 ( \31789 , \31783 , \31788 );
buf \U$31795 ( \31790 , \31789 );
buf \U$31796 ( \31791 , \31790 );
and \U$31797 ( \31792 , \31778 , \31791 );
and \U$31798 ( \31793 , \31764 , \31777 );
or \U$31799 ( \31794 , \31792 , \31793 );
buf \U$31800 ( \31795 , \31794 );
buf \U$31801 ( \31796 , \31795 );
buf \U$31802 ( \31797 , \27237 );
not \U$31803 ( \31798 , \31797 );
buf \U$31804 ( \31799 , \2124 );
not \U$31805 ( \31800 , \31799 );
or \U$31806 ( \31801 , \31798 , \31800 );
buf \U$31807 ( \31802 , \16500 );
buf \U$31808 ( \31803 , \30494 );
nand \U$31809 ( \31804 , \31802 , \31803 );
buf \U$31810 ( \31805 , \31804 );
buf \U$31811 ( \31806 , \31805 );
nand \U$31812 ( \31807 , \31801 , \31806 );
buf \U$31813 ( \31808 , \31807 );
buf \U$31814 ( \31809 , \31808 );
buf \U$31815 ( \31810 , \27526 );
not \U$31816 ( \31811 , \31810 );
buf \U$31817 ( \31812 , \12736 );
not \U$31818 ( \31813 , \31812 );
or \U$31819 ( \31814 , \31811 , \31813 );
buf \U$31820 ( \31815 , \12744 );
buf \U$31821 ( \31816 , \29221 );
nand \U$31822 ( \31817 , \31815 , \31816 );
buf \U$31823 ( \31818 , \31817 );
buf \U$31824 ( \31819 , \31818 );
nand \U$31825 ( \31820 , \31814 , \31819 );
buf \U$31826 ( \31821 , \31820 );
buf \U$31827 ( \31822 , \31821 );
xor \U$31828 ( \31823 , \31809 , \31822 );
buf \U$31829 ( \31824 , \27472 );
not \U$31830 ( \31825 , \31824 );
buf \U$31831 ( \31826 , \17595 );
not \U$31832 ( \31827 , \31826 );
or \U$31833 ( \31828 , \31825 , \31827 );
buf \U$31834 ( \31829 , \16071 );
buf \U$31835 ( \31830 , \31028 );
nand \U$31836 ( \31831 , \31829 , \31830 );
buf \U$31837 ( \31832 , \31831 );
buf \U$31838 ( \31833 , \31832 );
nand \U$31839 ( \31834 , \31828 , \31833 );
buf \U$31840 ( \31835 , \31834 );
buf \U$31841 ( \31836 , \31835 );
and \U$31842 ( \31837 , \31823 , \31836 );
and \U$31843 ( \31838 , \31809 , \31822 );
or \U$31844 ( \31839 , \31837 , \31838 );
buf \U$31845 ( \31840 , \31839 );
buf \U$31846 ( \31841 , \31840 );
xor \U$31847 ( \31842 , \31796 , \31841 );
buf \U$31848 ( \31843 , \27771 );
not \U$31849 ( \31844 , \31843 );
buf \U$31850 ( \31845 , \12929 );
not \U$31851 ( \31846 , \31845 );
or \U$31852 ( \31847 , \31844 , \31846 );
buf \U$31853 ( \31848 , \12937 );
buf \U$31854 ( \31849 , \30706 );
nand \U$31855 ( \31850 , \31848 , \31849 );
buf \U$31856 ( \31851 , \31850 );
buf \U$31857 ( \31852 , \31851 );
nand \U$31858 ( \31853 , \31847 , \31852 );
buf \U$31859 ( \31854 , \31853 );
buf \U$31860 ( \31855 , \31854 );
buf \U$31861 ( \31856 , \27433 );
not \U$31862 ( \31857 , \31856 );
buf \U$31863 ( \31858 , \16358 );
not \U$31864 ( \31859 , \31858 );
or \U$31865 ( \31860 , \31857 , \31859 );
buf \U$31866 ( \31861 , \30972 );
not \U$31867 ( \31862 , \31861 );
buf \U$31868 ( \31863 , \2070 );
nand \U$31869 ( \31864 , \31862 , \31863 );
buf \U$31870 ( \31865 , \31864 );
buf \U$31871 ( \31866 , \31865 );
nand \U$31872 ( \31867 , \31860 , \31866 );
buf \U$31873 ( \31868 , \31867 );
buf \U$31874 ( \31869 , \31868 );
or \U$31875 ( \31870 , \31855 , \31869 );
buf \U$31876 ( \31871 , \27490 );
not \U$31877 ( \31872 , \31871 );
buf \U$31878 ( \31873 , \1736 );
not \U$31879 ( \31874 , \31873 );
or \U$31880 ( \31875 , \31872 , \31874 );
buf \U$31881 ( \31876 , \993 );
buf \U$31882 ( \31877 , \30993 );
nand \U$31883 ( \31878 , \31876 , \31877 );
buf \U$31884 ( \31879 , \31878 );
buf \U$31885 ( \31880 , \31879 );
nand \U$31886 ( \31881 , \31875 , \31880 );
buf \U$31887 ( \31882 , \31881 );
buf \U$31888 ( \31883 , \31882 );
nand \U$31889 ( \31884 , \31870 , \31883 );
buf \U$31890 ( \31885 , \31884 );
buf \U$31891 ( \31886 , \31885 );
buf \U$31892 ( \31887 , \31854 );
buf \U$31893 ( \31888 , \31868 );
nand \U$31894 ( \31889 , \31887 , \31888 );
buf \U$31895 ( \31890 , \31889 );
buf \U$31896 ( \31891 , \31890 );
nand \U$31897 ( \31892 , \31886 , \31891 );
buf \U$31898 ( \31893 , \31892 );
buf \U$31899 ( \31894 , \31893 );
and \U$31900 ( \31895 , \31842 , \31894 );
and \U$31901 ( \31896 , \31796 , \31841 );
or \U$31902 ( \31897 , \31895 , \31896 );
buf \U$31903 ( \31898 , \31897 );
buf \U$31904 ( \31899 , \31898 );
and \U$31905 ( \31900 , \31751 , \31899 );
and \U$31906 ( \31901 , \31597 , \31750 );
or \U$31907 ( \31902 , \31900 , \31901 );
buf \U$31908 ( \31903 , \31902 );
buf \U$31909 ( \31904 , \31903 );
not \U$31910 ( \31905 , \31904 );
buf \U$31911 ( \31906 , \31905 );
buf \U$31912 ( \31907 , \31906 );
nand \U$31913 ( \31908 , \31593 , \31907 );
buf \U$31914 ( \31909 , \31908 );
not \U$31915 ( \31910 , \31909 );
buf \U$31916 ( \31911 , \31249 );
not \U$31917 ( \31912 , \31911 );
buf \U$31918 ( \31913 , \31428 );
not \U$31919 ( \31914 , \31913 );
or \U$31920 ( \31915 , \31912 , \31914 );
buf \U$31921 ( \31916 , \31249 );
buf \U$31922 ( \31917 , \31428 );
or \U$31923 ( \31918 , \31916 , \31917 );
nand \U$31924 ( \31919 , \31915 , \31918 );
buf \U$31925 ( \31920 , \31919 );
buf \U$31926 ( \31921 , \31920 );
buf \U$31927 ( \31922 , \31305 );
not \U$31928 ( \31923 , \31922 );
buf \U$31929 ( \31924 , \31923 );
buf \U$31930 ( \31925 , \31924 );
xnor \U$31931 ( \31926 , \31921 , \31925 );
buf \U$31932 ( \31927 , \31926 );
not \U$31933 ( \31928 , \31927 );
or \U$31934 ( \31929 , \31910 , \31928 );
not \U$31935 ( \31930 , \31592 );
nand \U$31936 ( \31931 , \31930 , \31903 );
nand \U$31937 ( \31932 , \31929 , \31931 );
and \U$31938 ( \31933 , \31453 , \31932 );
not \U$31939 ( \31934 , \31453 );
buf \U$31940 ( \31935 , \31932 );
not \U$31941 ( \31936 , \31935 );
buf \U$31942 ( \31937 , \31936 );
and \U$31943 ( \31938 , \31934 , \31937 );
nor \U$31944 ( \31939 , \31933 , \31938 );
buf \U$31945 ( \31940 , \31939 );
not \U$31946 ( \31941 , \31940 );
xor \U$31947 ( \31942 , \29186 , \29190 );
xor \U$31948 ( \31943 , \31942 , \29489 );
buf \U$31949 ( \31944 , \31943 );
buf \U$31950 ( \31945 , \31944 );
xor \U$31951 ( \31946 , \31006 , \31023 );
xor \U$31952 ( \31947 , \31946 , \31042 );
buf \U$31953 ( \31948 , \31947 );
buf \U$31954 ( \31949 , \31948 );
xor \U$31955 ( \31950 , \30896 , \30915 );
xor \U$31956 ( \31951 , \31950 , \30933 );
buf \U$31957 ( \31952 , \31951 );
buf \U$31958 ( \31953 , \31952 );
or \U$31959 ( \31954 , \31949 , \31953 );
xor \U$31960 ( \31955 , \30953 , \30966 );
xor \U$31961 ( \31956 , \31955 , \30983 );
buf \U$31962 ( \31957 , \31956 );
buf \U$31963 ( \31958 , \31957 );
nand \U$31964 ( \31959 , \31954 , \31958 );
buf \U$31965 ( \31960 , \31959 );
buf \U$31966 ( \31961 , \31960 );
buf \U$31967 ( \31962 , \31948 );
buf \U$31968 ( \31963 , \31952 );
nand \U$31969 ( \31964 , \31962 , \31963 );
buf \U$31970 ( \31965 , \31964 );
buf \U$31971 ( \31966 , \31965 );
nand \U$31972 ( \31967 , \31961 , \31966 );
buf \U$31973 ( \31968 , \31967 );
buf \U$31974 ( \31969 , \31968 );
xor \U$31975 ( \31970 , \30681 , \30718 );
xor \U$31976 ( \31971 , \31970 , \30699 );
buf \U$31977 ( \31972 , \31971 );
not \U$31978 ( \31973 , \31972 );
buf \U$31979 ( \31974 , \30795 );
buf \U$31980 ( \31975 , \30747 );
xor \U$31981 ( \31976 , \31974 , \31975 );
buf \U$31982 ( \31977 , \30769 );
xnor \U$31983 ( \31978 , \31976 , \31977 );
buf \U$31984 ( \31979 , \31978 );
buf \U$31985 ( \31980 , \31979 );
not \U$31986 ( \31981 , \31980 );
or \U$31987 ( \31982 , \31973 , \31981 );
buf \U$31988 ( \31983 , \31536 );
buf \U$31989 ( \31984 , \31556 );
and \U$31990 ( \31985 , \31983 , \31984 );
not \U$31991 ( \31986 , \31983 );
buf \U$31992 ( \31987 , \31559 );
and \U$31993 ( \31988 , \31986 , \31987 );
nor \U$31994 ( \31989 , \31985 , \31988 );
buf \U$31995 ( \31990 , \31989 );
buf \U$31996 ( \31991 , \31990 );
buf \U$31997 ( \31992 , \31523 );
xor \U$31998 ( \31993 , \31991 , \31992 );
buf \U$31999 ( \31994 , \31993 );
buf \U$32000 ( \31995 , \31994 );
nand \U$32001 ( \31996 , \31982 , \31995 );
buf \U$32002 ( \31997 , \31996 );
buf \U$32003 ( \31998 , \31997 );
buf \U$32004 ( \31999 , \31979 );
not \U$32005 ( \32000 , \31999 );
buf \U$32006 ( \32001 , \31971 );
not \U$32007 ( \32002 , \32001 );
buf \U$32008 ( \32003 , \32002 );
buf \U$32009 ( \32004 , \32003 );
nand \U$32010 ( \32005 , \32000 , \32004 );
buf \U$32011 ( \32006 , \32005 );
buf \U$32012 ( \32007 , \32006 );
nand \U$32013 ( \32008 , \31998 , \32007 );
buf \U$32014 ( \32009 , \32008 );
buf \U$32015 ( \32010 , \32009 );
xor \U$32016 ( \32011 , \31969 , \32010 );
buf \U$32017 ( \32012 , \31478 );
not \U$32018 ( \32013 , \32012 );
buf \U$32019 ( \32014 , \31484 );
not \U$32020 ( \32015 , \32014 );
or \U$32021 ( \32016 , \32013 , \32015 );
buf \U$32022 ( \32017 , \31484 );
buf \U$32024 ( \32018 , \31478 );
or \U$32025 ( \32019 , \32017 , \32018 );
nand \U$32026 ( \32020 , \32016 , \32019 );
buf \U$32027 ( \32021 , \32020 );
buf \U$32028 ( \32022 , \32021 );
buf \U$32029 ( \32023 , \31493 );
xor \U$32030 ( \32024 , \32022 , \32023 );
buf \U$32031 ( \32025 , \32024 );
buf \U$32032 ( \32026 , \32025 );
and \U$32033 ( \32027 , \32011 , \32026 );
and \U$32034 ( \32028 , \31969 , \32010 );
or \U$32035 ( \32029 , \32027 , \32028 );
buf \U$32036 ( \32030 , \32029 );
not \U$32037 ( \32031 , \32030 );
not \U$32038 ( \32032 , \32031 );
buf \U$32039 ( \32033 , \32032 );
or \U$32040 ( \32034 , \31945 , \32033 );
xor \U$32041 ( \32035 , \31569 , \31573 );
xor \U$32042 ( \32036 , \32035 , \31578 );
buf \U$32043 ( \32037 , \32036 );
buf \U$32044 ( \32038 , \32037 );
not \U$32045 ( \32039 , \32038 );
buf \U$32046 ( \32040 , \31299 );
not \U$32047 ( \32041 , \32040 );
buf \U$32048 ( \32042 , \31278 );
not \U$32049 ( \32043 , \32042 );
buf \U$32050 ( \32044 , \32043 );
buf \U$32051 ( \32045 , \32044 );
not \U$32052 ( \32046 , \32045 );
or \U$32053 ( \32047 , \32041 , \32046 );
buf \U$32054 ( \32048 , \31296 );
buf \U$32055 ( \32049 , \31278 );
nand \U$32056 ( \32050 , \32048 , \32049 );
buf \U$32057 ( \32051 , \32050 );
buf \U$32058 ( \32052 , \32051 );
nand \U$32059 ( \32053 , \32047 , \32052 );
buf \U$32060 ( \32054 , \32053 );
buf \U$32061 ( \32055 , \32054 );
buf \U$32062 ( \32056 , \31262 );
xnor \U$32063 ( \32057 , \32055 , \32056 );
buf \U$32064 ( \32058 , \32057 );
buf \U$32065 ( \32059 , \32058 );
not \U$32066 ( \32060 , \32059 );
buf \U$32067 ( \32061 , \32060 );
buf \U$32068 ( \32062 , \32061 );
not \U$32069 ( \32063 , \32062 );
or \U$32070 ( \32064 , \32039 , \32063 );
buf \U$32071 ( \32065 , \32037 );
not \U$32072 ( \32066 , \32065 );
buf \U$32073 ( \32067 , \32066 );
buf \U$32074 ( \32068 , \32067 );
not \U$32075 ( \32069 , \32068 );
buf \U$32076 ( \32070 , \32058 );
not \U$32077 ( \32071 , \32070 );
or \U$32078 ( \32072 , \32069 , \32071 );
xor \U$32079 ( \32073 , \29233 , \29197 );
buf \U$32080 ( \32074 , \32073 );
buf \U$32081 ( \32075 , \29210 );
not \U$32082 ( \32076 , \32075 );
buf \U$32083 ( \32077 , \32076 );
buf \U$32084 ( \32078 , \32077 );
and \U$32085 ( \32079 , \32074 , \32078 );
not \U$32086 ( \32080 , \32074 );
buf \U$32087 ( \32081 , \29210 );
and \U$32088 ( \32082 , \32080 , \32081 );
nor \U$32089 ( \32083 , \32079 , \32082 );
buf \U$32090 ( \32084 , \32083 );
buf \U$32091 ( \32085 , \32084 );
not \U$32092 ( \32086 , \32085 );
and \U$32093 ( \32087 , \26619 , \26620 );
buf \U$32094 ( \32088 , \32087 );
buf \U$32095 ( \32089 , \32088 );
buf \U$32096 ( \32090 , \32077 );
xor \U$32097 ( \32091 , \32089 , \32090 );
buf \U$32098 ( \32092 , \27794 );
not \U$32099 ( \32093 , \32092 );
buf \U$32100 ( \32094 , \27757 );
not \U$32101 ( \32095 , \32094 );
or \U$32102 ( \32096 , \32093 , \32095 );
buf \U$32103 ( \32097 , \27757 );
buf \U$32104 ( \32098 , \27794 );
or \U$32105 ( \32099 , \32097 , \32098 );
buf \U$32106 ( \32100 , \27777 );
nand \U$32107 ( \32101 , \32099 , \32100 );
buf \U$32108 ( \32102 , \32101 );
buf \U$32109 ( \32103 , \32102 );
nand \U$32110 ( \32104 , \32096 , \32103 );
buf \U$32111 ( \32105 , \32104 );
buf \U$32112 ( \32106 , \32105 );
and \U$32113 ( \32107 , \32091 , \32106 );
and \U$32114 ( \32108 , \32089 , \32090 );
or \U$32115 ( \32109 , \32107 , \32108 );
buf \U$32116 ( \32110 , \32109 );
buf \U$32117 ( \32111 , \32110 );
not \U$32118 ( \32112 , \32111 );
buf \U$32119 ( \32113 , \32112 );
buf \U$32120 ( \32114 , \32113 );
not \U$32121 ( \32115 , \32114 );
or \U$32122 ( \32116 , \32086 , \32115 );
xor \U$32123 ( \32117 , \27348 , \27366 );
and \U$32124 ( \32118 , \32117 , \27384 );
and \U$32125 ( \32119 , \27348 , \27366 );
or \U$32126 ( \32120 , \32118 , \32119 );
buf \U$32127 ( \32121 , \32120 );
buf \U$32128 ( \32122 , \32121 );
xor \U$32129 ( \32123 , \27405 , \27422 );
and \U$32130 ( \32124 , \32123 , \27440 );
and \U$32131 ( \32125 , \27405 , \27422 );
or \U$32132 ( \32126 , \32124 , \32125 );
buf \U$32133 ( \32127 , \32126 );
buf \U$32134 ( \32128 , \32127 );
xor \U$32135 ( \32129 , \32122 , \32128 );
xor \U$32136 ( \32130 , \27533 , \27554 );
and \U$32137 ( \32131 , \32130 , \27567 );
and \U$32138 ( \32132 , \27533 , \27554 );
or \U$32139 ( \32133 , \32131 , \32132 );
buf \U$32140 ( \32134 , \32133 );
buf \U$32141 ( \32135 , \32134 );
and \U$32142 ( \32136 , \32129 , \32135 );
and \U$32143 ( \32137 , \32122 , \32128 );
or \U$32144 ( \32138 , \32136 , \32137 );
buf \U$32145 ( \32139 , \32138 );
buf \U$32146 ( \32140 , \32139 );
nand \U$32147 ( \32141 , \32116 , \32140 );
buf \U$32148 ( \32142 , \32141 );
buf \U$32149 ( \32143 , \32142 );
buf \U$32150 ( \32144 , \32084 );
not \U$32151 ( \32145 , \32144 );
buf \U$32152 ( \32146 , \32110 );
nand \U$32153 ( \32147 , \32145 , \32146 );
buf \U$32154 ( \32148 , \32147 );
buf \U$32155 ( \32149 , \32148 );
nand \U$32156 ( \32150 , \32143 , \32149 );
buf \U$32157 ( \32151 , \32150 );
buf \U$32158 ( \32152 , \32151 );
nand \U$32159 ( \32153 , \32072 , \32152 );
buf \U$32160 ( \32154 , \32153 );
buf \U$32161 ( \32155 , \32154 );
nand \U$32162 ( \32156 , \32064 , \32155 );
buf \U$32163 ( \32157 , \32156 );
buf \U$32164 ( \32158 , \32157 );
nand \U$32165 ( \32159 , \32034 , \32158 );
buf \U$32166 ( \32160 , \32159 );
buf \U$32167 ( \32161 , \32160 );
buf \U$32168 ( \32162 , \31944 );
buf \U$32169 ( \32163 , \32032 );
nand \U$32170 ( \32164 , \32162 , \32163 );
buf \U$32171 ( \32165 , \32164 );
buf \U$32172 ( \32166 , \32165 );
nand \U$32173 ( \32167 , \32161 , \32166 );
buf \U$32174 ( \32168 , \32167 );
buf \U$32175 ( \32169 , \32168 );
buf \U$32176 ( \32170 , \30358 );
not \U$32177 ( \32171 , \32170 );
buf \U$32178 ( \32172 , \30374 );
nand \U$32179 ( \32173 , \32171 , \32172 );
buf \U$32180 ( \32174 , \32173 );
buf \U$32181 ( \32175 , \32174 );
not \U$32182 ( \32176 , \32175 );
buf \U$32183 ( \32177 , \30440 );
not \U$32184 ( \32178 , \32177 );
or \U$32185 ( \32179 , \32176 , \32178 );
buf \U$32186 ( \32180 , \30358 );
buf \U$32187 ( \32181 , \30371 );
nand \U$32188 ( \32182 , \32180 , \32181 );
buf \U$32189 ( \32183 , \32182 );
buf \U$32190 ( \32184 , \32183 );
nand \U$32191 ( \32185 , \32179 , \32184 );
buf \U$32192 ( \32186 , \32185 );
buf \U$32193 ( \32187 , \32186 );
buf \U$32194 ( \32188 , \31245 );
not \U$32195 ( \32189 , \32188 );
buf \U$32196 ( \32190 , \31197 );
not \U$32197 ( \32191 , \32190 );
or \U$32198 ( \32192 , \32189 , \32191 );
buf \U$32199 ( \32193 , \31139 );
nand \U$32200 ( \32194 , \32192 , \32193 );
buf \U$32201 ( \32195 , \32194 );
buf \U$32202 ( \32196 , \32195 );
buf \U$32203 ( \32197 , \31194 );
buf \U$32204 ( \32198 , \31239 );
nand \U$32205 ( \32199 , \32197 , \32198 );
buf \U$32206 ( \32200 , \32199 );
buf \U$32207 ( \32201 , \32200 );
nand \U$32208 ( \32202 , \32196 , \32201 );
buf \U$32209 ( \32203 , \32202 );
buf \U$32210 ( \32204 , \32203 );
xor \U$32211 ( \32205 , \32187 , \32204 );
buf \U$32212 ( \32206 , \31427 );
not \U$32213 ( \32207 , \32206 );
buf \U$32214 ( \32208 , \31365 );
not \U$32215 ( \32209 , \32208 );
or \U$32216 ( \32210 , \32207 , \32209 );
not \U$32217 ( \32211 , \31373 );
not \U$32218 ( \32212 , \31379 );
or \U$32219 ( \32213 , \32211 , \32212 );
or \U$32220 ( \32214 , \31427 , \31365 );
nand \U$32221 ( \32215 , \32213 , \32214 );
buf \U$32222 ( \32216 , \32215 );
nand \U$32223 ( \32217 , \32210 , \32216 );
buf \U$32224 ( \32218 , \32217 );
buf \U$32225 ( \32219 , \32218 );
xor \U$32226 ( \32220 , \32205 , \32219 );
buf \U$32227 ( \32221 , \32220 );
buf \U$32228 ( \32222 , \32221 );
buf \U$32229 ( \32223 , \31456 );
not \U$32230 ( \32224 , \32223 );
buf \U$32231 ( \32225 , \31582 );
not \U$32232 ( \32226 , \32225 );
or \U$32233 ( \32227 , \32224 , \32226 );
buf \U$32234 ( \32228 , \31582 );
buf \U$32235 ( \32229 , \31456 );
or \U$32236 ( \32230 , \32228 , \32229 );
buf \U$32237 ( \32231 , \31499 );
nand \U$32238 ( \32232 , \32230 , \32231 );
buf \U$32239 ( \32233 , \32232 );
buf \U$32240 ( \32234 , \32233 );
nand \U$32241 ( \32235 , \32227 , \32234 );
buf \U$32242 ( \32236 , \32235 );
buf \U$32243 ( \32237 , \32236 );
xor \U$32244 ( \32238 , \32222 , \32237 );
xor \U$32245 ( \32239 , \28044 , \28265 );
xor \U$32246 ( \32240 , \32239 , \28436 );
buf \U$32247 ( \32241 , \32240 );
buf \U$32248 ( \32242 , \32241 );
xor \U$32249 ( \32243 , \32238 , \32242 );
buf \U$32250 ( \32244 , \32243 );
buf \U$32251 ( \32245 , \32244 );
xor \U$32252 ( \32246 , \32169 , \32245 );
xor \U$32253 ( \32247 , \29183 , \29494 );
xor \U$32254 ( \32248 , \32247 , \29641 );
buf \U$32255 ( \32249 , \32248 );
buf \U$32256 ( \32250 , \32249 );
xor \U$32257 ( \32251 , \32246 , \32250 );
buf \U$32258 ( \32252 , \32251 );
not \U$32259 ( \32253 , \32252 );
buf \U$32260 ( \32254 , \32253 );
not \U$32261 ( \32255 , \32254 );
or \U$32262 ( \32256 , \31941 , \32255 );
xor \U$32263 ( \32257 , \29240 , \29296 );
xor \U$32264 ( \32258 , \32257 , \29484 );
buf \U$32265 ( \32259 , \32258 );
buf \U$32266 ( \32260 , \32259 );
buf \U$32267 ( \32261 , \27705 );
not \U$32268 ( \32262 , \32261 );
buf \U$32269 ( \32263 , \27735 );
not \U$32270 ( \32264 , \32263 );
or \U$32271 ( \32265 , \32262 , \32264 );
buf \U$32272 ( \32266 , \27705 );
buf \U$32273 ( \32267 , \27735 );
or \U$32274 ( \32268 , \32266 , \32267 );
buf \U$32275 ( \32269 , \27721 );
nand \U$32276 ( \32270 , \32268 , \32269 );
buf \U$32277 ( \32271 , \32270 );
buf \U$32278 ( \32272 , \32271 );
nand \U$32279 ( \32273 , \32265 , \32272 );
buf \U$32280 ( \32274 , \32273 );
buf \U$32281 ( \32275 , \32274 );
not \U$32282 ( \32276 , \32275 );
buf \U$32283 ( \32277 , \32276 );
buf \U$32284 ( \32278 , \32277 );
not \U$32285 ( \32279 , \32278 );
xor \U$32286 ( \32280 , \27244 , \27258 );
and \U$32287 ( \32281 , \32280 , \27279 );
and \U$32288 ( \32282 , \27244 , \27258 );
or \U$32289 ( \32283 , \32281 , \32282 );
buf \U$32290 ( \32284 , \32283 );
buf \U$32291 ( \32285 , \32284 );
not \U$32292 ( \32286 , \32285 );
buf \U$32293 ( \32287 , \32286 );
buf \U$32294 ( \32288 , \32287 );
not \U$32295 ( \32289 , \32288 );
or \U$32296 ( \32290 , \32279 , \32289 );
xor \U$32297 ( \32291 , \27588 , \27603 );
and \U$32298 ( \32292 , \32291 , \27623 );
and \U$32299 ( \32293 , \27588 , \27603 );
or \U$32300 ( \32294 , \32292 , \32293 );
buf \U$32301 ( \32295 , \32294 );
buf \U$32302 ( \32296 , \32295 );
nand \U$32303 ( \32297 , \32290 , \32296 );
buf \U$32304 ( \32298 , \32297 );
buf \U$32305 ( \32299 , \32298 );
buf \U$32306 ( \32300 , \32284 );
buf \U$32307 ( \32301 , \32274 );
nand \U$32308 ( \32302 , \32300 , \32301 );
buf \U$32309 ( \32303 , \32302 );
buf \U$32310 ( \32304 , \32303 );
nand \U$32311 ( \32305 , \32299 , \32304 );
buf \U$32312 ( \32306 , \32305 );
buf \U$32313 ( \32307 , \32306 );
buf \U$32314 ( \32308 , \27496 );
not \U$32315 ( \32309 , \32308 );
buf \U$32316 ( \32310 , \27463 );
not \U$32317 ( \32311 , \32310 );
or \U$32318 ( \32312 , \32309 , \32311 );
or \U$32319 ( \32313 , \27463 , \27496 );
nand \U$32320 ( \32314 , \32313 , \27478 );
buf \U$32321 ( \32315 , \32314 );
nand \U$32322 ( \32316 , \32312 , \32315 );
buf \U$32323 ( \32317 , \32316 );
buf \U$32324 ( \32318 , \32317 );
not \U$32325 ( \32319 , \32318 );
xor \U$32326 ( \32320 , \27655 , \27672 );
and \U$32327 ( \32321 , \32320 , \27689 );
and \U$32328 ( \32322 , \27655 , \27672 );
or \U$32329 ( \32323 , \32321 , \32322 );
buf \U$32330 ( \32324 , \32323 );
buf \U$32331 ( \32325 , \32324 );
not \U$32332 ( \32326 , \32325 );
or \U$32333 ( \32327 , \32319 , \32326 );
buf \U$32334 ( \32328 , \32324 );
buf \U$32335 ( \32329 , \32317 );
or \U$32336 ( \32330 , \32328 , \32329 );
xor \U$32337 ( \32331 , \27297 , \27311 );
and \U$32338 ( \32332 , \32331 , \27326 );
and \U$32339 ( \32333 , \27297 , \27311 );
or \U$32340 ( \32334 , \32332 , \32333 );
buf \U$32341 ( \32335 , \32334 );
buf \U$32342 ( \32336 , \32335 );
nand \U$32343 ( \32337 , \32330 , \32336 );
buf \U$32344 ( \32338 , \32337 );
buf \U$32345 ( \32339 , \32338 );
nand \U$32346 ( \32340 , \32327 , \32339 );
buf \U$32347 ( \32341 , \32340 );
buf \U$32348 ( \32342 , \32341 );
xor \U$32349 ( \32343 , \32307 , \32342 );
xor \U$32350 ( \32344 , \29359 , \29418 );
xor \U$32351 ( \32345 , \32344 , \29479 );
buf \U$32352 ( \32346 , \32345 );
buf \U$32353 ( \32347 , \32346 );
and \U$32354 ( \32348 , \32343 , \32347 );
and \U$32355 ( \32349 , \32307 , \32342 );
or \U$32356 ( \32350 , \32348 , \32349 );
buf \U$32357 ( \32351 , \32350 );
buf \U$32358 ( \32352 , \32351 );
xor \U$32359 ( \32353 , \32260 , \32352 );
xor \U$32360 ( \32354 , \31597 , \31750 );
xor \U$32361 ( \32355 , \32354 , \31899 );
buf \U$32362 ( \32356 , \32355 );
buf \U$32363 ( \32357 , \32356 );
and \U$32364 ( \32358 , \32353 , \32357 );
and \U$32365 ( \32359 , \32260 , \32352 );
or \U$32366 ( \32360 , \32358 , \32359 );
buf \U$32367 ( \32361 , \32360 );
buf \U$32368 ( \32362 , \32361 );
xor \U$32369 ( \32363 , \30471 , \30853 );
xor \U$32370 ( \32364 , \32363 , \31053 );
buf \U$32371 ( \32365 , \32364 );
buf \U$32372 ( \32366 , \32365 );
xor \U$32373 ( \32367 , \32362 , \32366 );
xor \U$32374 ( \32368 , \31796 , \31841 );
xor \U$32375 ( \32369 , \32368 , \31894 );
buf \U$32376 ( \32370 , \32369 );
buf \U$32377 ( \32371 , \32370 );
not \U$32378 ( \32372 , \32371 );
xor \U$32379 ( \32373 , \31647 , \31743 );
xnor \U$32380 ( \32374 , \32373 , \31687 );
buf \U$32381 ( \32375 , \32374 );
not \U$32382 ( \32376 , \32375 );
buf \U$32383 ( \32377 , \32376 );
buf \U$32384 ( \32378 , \32377 );
not \U$32385 ( \32379 , \32378 );
or \U$32386 ( \32380 , \32372 , \32379 );
buf \U$32387 ( \32381 , \32370 );
not \U$32388 ( \32382 , \32381 );
buf \U$32389 ( \32383 , \32382 );
buf \U$32390 ( \32384 , \32383 );
not \U$32391 ( \32385 , \32384 );
buf \U$32392 ( \32386 , \32374 );
not \U$32393 ( \32387 , \32386 );
or \U$32394 ( \32388 , \32385 , \32387 );
xor \U$32395 ( \32389 , \29372 , \29392 );
xnor \U$32396 ( \32390 , \32389 , \29410 );
buf \U$32397 ( \32391 , \32390 );
buf \U$32398 ( \32392 , \29327 );
buf \U$32399 ( \32393 , \29309 );
xor \U$32400 ( \32394 , \32392 , \32393 );
buf \U$32401 ( \32395 , \29352 );
xor \U$32402 ( \32396 , \32394 , \32395 );
buf \U$32403 ( \32397 , \32396 );
buf \U$32404 ( \32398 , \32397 );
xor \U$32405 ( \32399 , \32391 , \32398 );
xor \U$32406 ( \32400 , \29472 , \29432 );
xor \U$32407 ( \32401 , \32400 , \29450 );
buf \U$32408 ( \32402 , \32401 );
and \U$32409 ( \32403 , \32399 , \32402 );
and \U$32410 ( \32404 , \32391 , \32398 );
or \U$32411 ( \32405 , \32403 , \32404 );
buf \U$32412 ( \32406 , \32405 );
buf \U$32413 ( \32407 , \32406 );
nand \U$32414 ( \32408 , \32388 , \32407 );
buf \U$32415 ( \32409 , \32408 );
buf \U$32416 ( \32410 , \32409 );
nand \U$32417 ( \32411 , \32380 , \32410 );
buf \U$32418 ( \32412 , \32411 );
buf \U$32419 ( \32413 , \32412 );
buf \U$32420 ( \32414 , \31609 );
buf \U$32421 ( \32415 , \31622 );
xor \U$32422 ( \32416 , \32414 , \32415 );
buf \U$32423 ( \32417 , \31636 );
xnor \U$32424 ( \32418 , \32416 , \32417 );
buf \U$32425 ( \32419 , \32418 );
buf \U$32426 ( \32420 , \32419 );
not \U$32427 ( \32421 , \32420 );
buf \U$32428 ( \32422 , \31705 );
buf \U$32429 ( \32423 , \31737 );
xor \U$32430 ( \32424 , \32422 , \32423 );
buf \U$32431 ( \32425 , \31719 );
xnor \U$32432 ( \32426 , \32424 , \32425 );
buf \U$32433 ( \32427 , \32426 );
buf \U$32434 ( \32428 , \32427 );
not \U$32435 ( \32429 , \32428 );
or \U$32436 ( \32430 , \32421 , \32429 );
xor \U$32437 ( \32431 , \31809 , \31822 );
xor \U$32438 ( \32432 , \32431 , \31836 );
buf \U$32439 ( \32433 , \32432 );
buf \U$32440 ( \32434 , \32433 );
nand \U$32441 ( \32435 , \32430 , \32434 );
buf \U$32442 ( \32436 , \32435 );
buf \U$32443 ( \32437 , \32436 );
buf \U$32444 ( \32438 , \32427 );
not \U$32445 ( \32439 , \32438 );
buf \U$32446 ( \32440 , \32419 );
not \U$32447 ( \32441 , \32440 );
buf \U$32448 ( \32442 , \32441 );
buf \U$32449 ( \32443 , \32442 );
nand \U$32450 ( \32444 , \32439 , \32443 );
buf \U$32451 ( \32445 , \32444 );
buf \U$32452 ( \32446 , \32445 );
nand \U$32453 ( \32447 , \32437 , \32446 );
buf \U$32454 ( \32448 , \32447 );
buf \U$32455 ( \32449 , \32448 );
xor \U$32456 ( \32450 , \31764 , \31777 );
xor \U$32457 ( \32451 , \32450 , \31791 );
buf \U$32458 ( \32452 , \32451 );
buf \U$32459 ( \32453 , \32452 );
xor \U$32460 ( \32454 , \31655 , \31668 );
xor \U$32461 ( \32455 , \32454 , \31683 );
buf \U$32462 ( \32456 , \32455 );
buf \U$32463 ( \32457 , \32456 );
xor \U$32464 ( \32458 , \32453 , \32457 );
xor \U$32465 ( \32459 , \31882 , \31854 );
xor \U$32466 ( \32460 , \32459 , \31868 );
buf \U$32467 ( \32461 , \32460 );
and \U$32468 ( \32462 , \32458 , \32461 );
and \U$32469 ( \32463 , \32453 , \32457 );
or \U$32470 ( \32464 , \32462 , \32463 );
buf \U$32471 ( \32465 , \32464 );
buf \U$32472 ( \32466 , \32465 );
xor \U$32473 ( \32467 , \32449 , \32466 );
buf \U$32474 ( \32468 , \30840 );
buf \U$32475 ( \32469 , \30816 );
xor \U$32476 ( \32470 , \32468 , \32469 );
buf \U$32477 ( \32471 , \30827 );
xor \U$32478 ( \32472 , \32470 , \32471 );
buf \U$32479 ( \32473 , \32472 );
buf \U$32480 ( \32474 , \32473 );
and \U$32481 ( \32475 , \32467 , \32474 );
and \U$32482 ( \32476 , \32449 , \32466 );
or \U$32483 ( \32477 , \32475 , \32476 );
buf \U$32484 ( \32478 , \32477 );
buf \U$32485 ( \32479 , \32478 );
xor \U$32486 ( \32480 , \32413 , \32479 );
xor \U$32487 ( \32481 , \31969 , \32010 );
xor \U$32488 ( \32482 , \32481 , \32026 );
buf \U$32489 ( \32483 , \32482 );
buf \U$32490 ( \32484 , \32483 );
and \U$32491 ( \32485 , \32480 , \32484 );
and \U$32492 ( \32486 , \32413 , \32479 );
or \U$32493 ( \32487 , \32485 , \32486 );
buf \U$32494 ( \32488 , \32487 );
buf \U$32495 ( \32489 , \32488 );
and \U$32496 ( \32490 , \32367 , \32489 );
and \U$32497 ( \32491 , \32362 , \32366 );
or \U$32498 ( \32492 , \32490 , \32491 );
buf \U$32499 ( \32493 , \32492 );
buf \U$32500 ( \32494 , \32493 );
nand \U$32501 ( \32495 , \32256 , \32494 );
buf \U$32502 ( \32496 , \32495 );
buf \U$32503 ( \32497 , \32496 );
buf \U$32504 ( \32498 , \31939 );
not \U$32505 ( \32499 , \32498 );
buf \U$32506 ( \32500 , \32252 );
nand \U$32507 ( \32501 , \32499 , \32500 );
buf \U$32508 ( \32502 , \32501 );
buf \U$32509 ( \32503 , \32502 );
nand \U$32510 ( \32504 , \32497 , \32503 );
buf \U$32511 ( \32505 , \32504 );
buf \U$32512 ( \32506 , \32505 );
not \U$32513 ( \32507 , \32506 );
buf \U$32514 ( \32508 , \32507 );
buf \U$32515 ( \32509 , \32508 );
not \U$32516 ( \32510 , \32509 );
or \U$32517 ( \32511 , \30346 , \32510 );
buf \U$32518 ( \32512 , \31452 );
not \U$32519 ( \32513 , \32512 );
buf \U$32520 ( \32514 , \32513 );
buf \U$32521 ( \32515 , \32514 );
not \U$32522 ( \32516 , \32515 );
buf \U$32523 ( \32517 , \31932 );
not \U$32524 ( \32518 , \32517 );
or \U$32525 ( \32519 , \32516 , \32518 );
buf \U$32526 ( \32520 , \31932 );
buf \U$32527 ( \32521 , \32514 );
or \U$32528 ( \32522 , \32520 , \32521 );
buf \U$32530 ( \32523 , \31057 );
nand \U$32531 ( \32524 , \32522 , \32523 );
buf \U$32532 ( \32525 , \32524 );
buf \U$32533 ( \32526 , \32525 );
nand \U$32534 ( \32527 , \32519 , \32526 );
buf \U$32535 ( \32528 , \32527 );
buf \U$32536 ( \32529 , \32528 );
not \U$32537 ( \32530 , \32529 );
buf \U$32538 ( \32531 , \31442 );
not \U$32539 ( \32532 , \32531 );
buf \U$32540 ( \32533 , \31087 );
not \U$32541 ( \32534 , \32533 );
buf \U$32542 ( \32535 , \31068 );
nand \U$32543 ( \32536 , \32534 , \32535 );
buf \U$32544 ( \32537 , \32536 );
buf \U$32545 ( \32538 , \32537 );
not \U$32546 ( \32539 , \32538 );
or \U$32547 ( \32540 , \32532 , \32539 );
buf \U$32548 ( \32541 , \31068 );
not \U$32549 ( \32542 , \32541 );
buf \U$32550 ( \32543 , \31087 );
nand \U$32551 ( \32544 , \32542 , \32543 );
buf \U$32552 ( \32545 , \32544 );
buf \U$32553 ( \32546 , \32545 );
nand \U$32554 ( \32547 , \32540 , \32546 );
buf \U$32555 ( \32548 , \32547 );
buf \U$32556 ( \32549 , \32548 );
xor \U$32557 ( \32550 , \29564 , \29574 );
and \U$32558 ( \32551 , \32550 , \29628 );
and \U$32559 ( \32552 , \29564 , \29574 );
or \U$32560 ( \32553 , \32551 , \32552 );
buf \U$32561 ( \32554 , \32553 );
buf \U$32562 ( \32555 , \32554 );
xor \U$32563 ( \32556 , \32187 , \32204 );
and \U$32564 ( \32557 , \32556 , \32219 );
and \U$32565 ( \32558 , \32187 , \32204 );
or \U$32566 ( \32559 , \32557 , \32558 );
buf \U$32567 ( \32560 , \32559 );
buf \U$32568 ( \32561 , \32560 );
xor \U$32569 ( \32562 , \32555 , \32561 );
xor \U$32570 ( \32563 , \29520 , \29540 );
and \U$32571 ( \32564 , \32563 , \29561 );
and \U$32572 ( \32565 , \29520 , \29540 );
or \U$32573 ( \32566 , \32564 , \32565 );
buf \U$32574 ( \32567 , \32566 );
buf \U$32575 ( \32568 , \32567 );
xor \U$32576 ( \32569 , \28458 , \28473 );
and \U$32577 ( \32570 , \32569 , \28543 );
and \U$32578 ( \32571 , \28458 , \28473 );
or \U$32579 ( \32572 , \32570 , \32571 );
buf \U$32580 ( \32573 , \32572 );
buf \U$32581 ( \32574 , \32573 );
xor \U$32582 ( \32575 , \32568 , \32574 );
not \U$32583 ( \32576 , \28629 );
not \U$32584 ( \32577 , \28623 );
or \U$32585 ( \32578 , \32576 , \32577 );
buf \U$32586 ( \32579 , \28629 );
buf \U$32587 ( \32580 , \28623 );
or \U$32588 ( \32581 , \32579 , \32580 );
buf \U$32589 ( \32582 , \28555 );
nand \U$32590 ( \32583 , \32581 , \32582 );
buf \U$32591 ( \32584 , \32583 );
nand \U$32592 ( \32585 , \32578 , \32584 );
buf \U$32593 ( \32586 , \32585 );
xor \U$32594 ( \32587 , \32575 , \32586 );
buf \U$32595 ( \32588 , \32587 );
buf \U$32596 ( \32589 , \32588 );
xor \U$32597 ( \32590 , \32562 , \32589 );
buf \U$32598 ( \32591 , \32590 );
not \U$32599 ( \32592 , \32591 );
buf \U$32600 ( \32593 , \32592 );
and \U$32601 ( \32594 , \32549 , \32593 );
not \U$32602 ( \32595 , \32549 );
buf \U$32603 ( \32596 , \32591 );
and \U$32604 ( \32597 , \32595 , \32596 );
nor \U$32605 ( \32598 , \32594 , \32597 );
buf \U$32606 ( \32599 , \32598 );
buf \U$32607 ( \32600 , \32599 );
not \U$32608 ( \32601 , \32600 );
xor \U$32609 ( \32602 , \32222 , \32237 );
and \U$32610 ( \32603 , \32602 , \32242 );
and \U$32611 ( \32604 , \32222 , \32237 );
or \U$32612 ( \32605 , \32603 , \32604 );
buf \U$32613 ( \32606 , \32605 );
buf \U$32614 ( \32607 , \32606 );
not \U$32615 ( \32608 , \32607 );
and \U$32616 ( \32609 , \32601 , \32608 );
buf \U$32617 ( \32610 , \32599 );
buf \U$32618 ( \32611 , \32606 );
and \U$32619 ( \32612 , \32610 , \32611 );
nor \U$32620 ( \32613 , \32609 , \32612 );
buf \U$32621 ( \32614 , \32613 );
buf \U$32622 ( \32615 , \32614 );
not \U$32623 ( \32616 , \32615 );
or \U$32624 ( \32617 , \32530 , \32616 );
buf \U$32625 ( \32618 , \32614 );
buf \U$32626 ( \32619 , \32528 );
or \U$32627 ( \32620 , \32618 , \32619 );
nand \U$32628 ( \32621 , \32617 , \32620 );
buf \U$32629 ( \32622 , \32621 );
buf \U$32630 ( \32623 , \32622 );
xor \U$32631 ( \32624 , \32169 , \32245 );
and \U$32632 ( \32625 , \32624 , \32250 );
and \U$32633 ( \32626 , \32169 , \32245 );
or \U$32634 ( \32627 , \32625 , \32626 );
buf \U$32635 ( \32628 , \32627 );
buf \U$32636 ( \32629 , \32628 );
xnor \U$32637 ( \32630 , \32623 , \32629 );
buf \U$32638 ( \32631 , \32630 );
buf \U$32639 ( \32632 , \32631 );
not \U$32640 ( \32633 , \32632 );
buf \U$32641 ( \32634 , \32633 );
buf \U$32642 ( \32635 , \32634 );
nand \U$32643 ( \32636 , \32511 , \32635 );
buf \U$32644 ( \32637 , \32636 );
buf \U$32645 ( \32638 , \32637 );
buf \U$32646 ( \32639 , \32505 );
buf \U$32647 ( \32640 , \30341 );
nand \U$32648 ( \32641 , \32639 , \32640 );
buf \U$32649 ( \32642 , \32641 );
buf \U$32650 ( \32643 , \32642 );
nand \U$32651 ( \32644 , \32638 , \32643 );
buf \U$32652 ( \32645 , \32644 );
buf \U$32653 ( \32646 , \32645 );
not \U$32654 ( \32647 , \32646 );
buf \U$32655 ( \32648 , \29667 );
not \U$32656 ( \32649 , \32648 );
buf \U$32657 ( \32650 , \29759 );
not \U$32658 ( \32651 , \32650 );
or \U$32659 ( \32652 , \32649 , \32651 );
buf \U$32660 ( \32653 , \29670 );
not \U$32661 ( \32654 , \32653 );
buf \U$32662 ( \32655 , \29758 );
not \U$32663 ( \32656 , \32655 );
or \U$32664 ( \32657 , \32654 , \32656 );
buf \U$32665 ( \32658 , \29700 );
nand \U$32666 ( \32659 , \32657 , \32658 );
buf \U$32667 ( \32660 , \32659 );
buf \U$32668 ( \32661 , \32660 );
nand \U$32669 ( \32662 , \32652 , \32661 );
buf \U$32670 ( \32663 , \32662 );
buf \U$32671 ( \32664 , \32663 );
not \U$32672 ( \32665 , \32664 );
or \U$32673 ( \32666 , \29724 , \29739 );
nand \U$32674 ( \32667 , \32666 , \29755 );
buf \U$32675 ( \32668 , \29739 );
buf \U$32676 ( \32669 , \29724 );
nand \U$32677 ( \32670 , \32668 , \32669 );
buf \U$32678 ( \32671 , \32670 );
nand \U$32679 ( \32672 , \32667 , \32671 );
buf \U$32680 ( \32673 , \32672 );
not \U$32681 ( \32674 , \32673 );
buf \U$32682 ( \32675 , \29162 );
not \U$32683 ( \32676 , \32675 );
buf \U$32684 ( \32677 , \29131 );
not \U$32685 ( \32678 , \32677 );
or \U$32686 ( \32679 , \32676 , \32678 );
buf \U$32687 ( \32680 , \29131 );
buf \U$32688 ( \32681 , \29162 );
or \U$32689 ( \32682 , \32680 , \32681 );
buf \U$32690 ( \32683 , \29147 );
nand \U$32691 ( \32684 , \32682 , \32683 );
buf \U$32692 ( \32685 , \32684 );
buf \U$32693 ( \32686 , \32685 );
nand \U$32694 ( \32687 , \32679 , \32686 );
buf \U$32695 ( \32688 , \32687 );
buf \U$32696 ( \32689 , \32688 );
not \U$32697 ( \32690 , \32689 );
buf \U$32698 ( \32691 , \32690 );
buf \U$32699 ( \32692 , \32691 );
not \U$32700 ( \32693 , \32692 );
or \U$32701 ( \32694 , \32674 , \32693 );
buf \U$32702 ( \32695 , \32672 );
not \U$32703 ( \32696 , \32695 );
buf \U$32704 ( \32697 , \32688 );
nand \U$32705 ( \32698 , \32696 , \32697 );
buf \U$32706 ( \32699 , \32698 );
buf \U$32707 ( \32700 , \32699 );
nand \U$32708 ( \32701 , \32694 , \32700 );
buf \U$32709 ( \32702 , \32701 );
buf \U$32710 ( \32703 , \32702 );
buf \U$32711 ( \32704 , \29820 );
not \U$32712 ( \32705 , \32704 );
buf \U$32713 ( \32706 , \29800 );
not \U$32714 ( \32707 , \32706 );
or \U$32715 ( \32708 , \32705 , \32707 );
buf \U$32716 ( \32709 , \29800 );
buf \U$32717 ( \32710 , \29820 );
or \U$32718 ( \32711 , \32709 , \32710 );
buf \U$32719 ( \32712 , \29787 );
nand \U$32720 ( \32713 , \32711 , \32712 );
buf \U$32721 ( \32714 , \32713 );
buf \U$32722 ( \32715 , \32714 );
nand \U$32723 ( \32716 , \32708 , \32715 );
buf \U$32724 ( \32717 , \32716 );
buf \U$32725 ( \32718 , \32717 );
not \U$32726 ( \32719 , \32718 );
xor \U$32727 ( \32720 , \30282 , \30296 );
and \U$32728 ( \32721 , \32720 , \30313 );
and \U$32729 ( \32722 , \30282 , \30296 );
or \U$32730 ( \32723 , \32721 , \32722 );
buf \U$32731 ( \32724 , \32723 );
buf \U$32732 ( \32725 , \32724 );
not \U$32733 ( \32726 , \32725 );
buf \U$32734 ( \32727 , \32726 );
buf \U$32735 ( \32728 , \32727 );
not \U$32736 ( \32729 , \32728 );
or \U$32737 ( \32730 , \32719 , \32729 );
buf \U$32738 ( \32731 , \32717 );
buf \U$32739 ( \32732 , \32727 );
or \U$32740 ( \32733 , \32731 , \32732 );
nand \U$32741 ( \32734 , \32730 , \32733 );
buf \U$32742 ( \32735 , \32734 );
buf \U$32743 ( \32736 , \32735 );
xor \U$32744 ( \32737 , \30179 , \30196 );
and \U$32745 ( \32738 , \32737 , \30216 );
and \U$32746 ( \32739 , \30179 , \30196 );
or \U$32747 ( \32740 , \32738 , \32739 );
buf \U$32748 ( \32741 , \32740 );
buf \U$32749 ( \32742 , \32741 );
not \U$32750 ( \32743 , \32742 );
buf \U$32751 ( \32744 , \32743 );
buf \U$32752 ( \32745 , \32744 );
and \U$32753 ( \32746 , \32736 , \32745 );
not \U$32754 ( \32747 , \32736 );
buf \U$32755 ( \32748 , \32741 );
and \U$32756 ( \32749 , \32747 , \32748 );
nor \U$32757 ( \32750 , \32746 , \32749 );
buf \U$32758 ( \32751 , \32750 );
buf \U$32759 ( \32752 , \32751 );
and \U$32760 ( \32753 , \32703 , \32752 );
not \U$32761 ( \32754 , \32703 );
buf \U$32762 ( \32755 , \32751 );
not \U$32763 ( \32756 , \32755 );
buf \U$32764 ( \32757 , \32756 );
buf \U$32765 ( \32758 , \32757 );
and \U$32766 ( \32759 , \32754 , \32758 );
nor \U$32767 ( \32760 , \32753 , \32759 );
buf \U$32768 ( \32761 , \32760 );
buf \U$32769 ( \32762 , \32761 );
not \U$32770 ( \32763 , \32762 );
and \U$32771 ( \32764 , \32665 , \32763 );
buf \U$32772 ( \32765 , \32761 );
buf \U$32773 ( \32766 , \32663 );
and \U$32774 ( \32767 , \32765 , \32766 );
nor \U$32775 ( \32768 , \32764 , \32767 );
buf \U$32776 ( \32769 , \32768 );
buf \U$32777 ( \32770 , \32769 );
buf \U$32778 ( \32771 , \30208 );
not \U$32779 ( \32772 , \32771 );
buf \U$32780 ( \32773 , \16358 );
not \U$32781 ( \32774 , \32773 );
or \U$32782 ( \32775 , \32772 , \32774 );
buf \U$32783 ( \32776 , \734 );
buf \U$32784 ( \32777 , RIc0da378_97);
buf \U$32785 ( \32778 , RIc0d7d80_16);
xor \U$32786 ( \32779 , \32777 , \32778 );
buf \U$32787 ( \32780 , \32779 );
buf \U$32788 ( \32781 , \32780 );
nand \U$32789 ( \32782 , \32776 , \32781 );
buf \U$32790 ( \32783 , \32782 );
buf \U$32791 ( \32784 , \32783 );
nand \U$32792 ( \32785 , \32775 , \32784 );
buf \U$32793 ( \32786 , \32785 );
buf \U$32794 ( \32787 , \29998 );
not \U$32795 ( \32788 , \32787 );
buf \U$32796 ( \32789 , \27660 );
not \U$32797 ( \32790 , \32789 );
or \U$32798 ( \32791 , \32788 , \32790 );
buf \U$32799 ( \32792 , \20211 );
buf \U$32800 ( \32793 , RIc0d77e0_4);
buf \U$32801 ( \32794 , RIc0da918_109);
xor \U$32802 ( \32795 , \32793 , \32794 );
buf \U$32803 ( \32796 , \32795 );
buf \U$32804 ( \32797 , \32796 );
nand \U$32805 ( \32798 , \32792 , \32797 );
buf \U$32806 ( \32799 , \32798 );
buf \U$32807 ( \32800 , \32799 );
nand \U$32808 ( \32801 , \32791 , \32800 );
buf \U$32809 ( \32802 , \32801 );
xor \U$32810 ( \32803 , \32786 , \32802 );
buf \U$32811 ( \32804 , \29794 );
not \U$32812 ( \32805 , \32804 );
buf \U$32813 ( \32806 , \2088 );
not \U$32814 ( \32807 , \32806 );
or \U$32815 ( \32808 , \32805 , \32807 );
buf \U$32816 ( \32809 , \993 );
buf \U$32817 ( \32810 , RIc0d8410_30);
buf \U$32818 ( \32811 , RIc0d9ce8_83);
xor \U$32819 ( \32812 , \32810 , \32811 );
buf \U$32820 ( \32813 , \32812 );
buf \U$32821 ( \32814 , \32813 );
nand \U$32822 ( \32815 , \32809 , \32814 );
buf \U$32823 ( \32816 , \32815 );
buf \U$32824 ( \32817 , \32816 );
nand \U$32825 ( \32818 , \32808 , \32817 );
buf \U$32826 ( \32819 , \32818 );
xor \U$32827 ( \32820 , \32803 , \32819 );
buf \U$32828 ( \32821 , \32820 );
and \U$32829 ( \32822 , \28967 , \28968 );
buf \U$32830 ( \32823 , \32822 );
buf \U$32831 ( \32824 , \32823 );
buf \U$32832 ( \32825 , \6270 );
not \U$32833 ( \32826 , \32825 );
buf \U$32834 ( \32827 , \30136 );
not \U$32835 ( \32828 , \32827 );
and \U$32836 ( \32829 , \32826 , \32828 );
xor \U$32837 ( \32830 , RIc0d9ec8_87, RIc0d8230_26);
buf \U$32838 ( \32831 , \32830 );
not \U$32839 ( \32832 , \32831 );
buf \U$32840 ( \32833 , \819 );
nor \U$32841 ( \32834 , \32832 , \32833 );
buf \U$32842 ( \32835 , \32834 );
buf \U$32843 ( \32836 , \32835 );
nor \U$32844 ( \32837 , \32829 , \32836 );
buf \U$32845 ( \32838 , \32837 );
buf \U$32846 ( \32839 , \32838 );
xor \U$32847 ( \32840 , \32824 , \32839 );
buf \U$32848 ( \32841 , \30252 );
not \U$32849 ( \32842 , \32841 );
buf \U$32850 ( \32843 , \30236 );
not \U$32851 ( \32844 , \32843 );
or \U$32852 ( \32845 , \32842 , \32844 );
buf \U$32853 ( \32846 , \30252 );
buf \U$32854 ( \32847 , \30236 );
or \U$32855 ( \32848 , \32846 , \32847 );
buf \U$32856 ( \32849 , \30269 );
nand \U$32857 ( \32850 , \32848 , \32849 );
buf \U$32858 ( \32851 , \32850 );
buf \U$32859 ( \32852 , \32851 );
nand \U$32860 ( \32853 , \32845 , \32852 );
buf \U$32861 ( \32854 , \32853 );
buf \U$32862 ( \32855 , \32854 );
xor \U$32863 ( \32856 , \32840 , \32855 );
buf \U$32864 ( \32857 , \32856 );
buf \U$32865 ( \32858 , \32857 );
xor \U$32866 ( \32859 , \32821 , \32858 );
buf \U$32867 ( \32860 , \29536 );
not \U$32868 ( \32861 , \32860 );
buf \U$32869 ( \32862 , \29687 );
not \U$32870 ( \32863 , \32862 );
or \U$32871 ( \32864 , \32861 , \32863 );
buf \U$32872 ( \32865 , \29687 );
buf \U$32873 ( \32866 , \29536 );
or \U$32874 ( \32867 , \32865 , \32866 );
buf \U$32875 ( \32868 , \29694 );
nand \U$32876 ( \32869 , \32867 , \32868 );
buf \U$32877 ( \32870 , \32869 );
buf \U$32878 ( \32871 , \32870 );
nand \U$32879 ( \32872 , \32864 , \32871 );
buf \U$32880 ( \32873 , \32872 );
buf \U$32881 ( \32874 , \32873 );
xor \U$32882 ( \32875 , \32859 , \32874 );
buf \U$32883 ( \32876 , \32875 );
buf \U$32884 ( \32877 , \32876 );
not \U$32885 ( \32878 , \32877 );
buf \U$32886 ( \32879 , \32878 );
buf \U$32887 ( \32880 , \32879 );
and \U$32888 ( \32881 , \32770 , \32880 );
not \U$32889 ( \32882 , \32770 );
buf \U$32890 ( \32883 , \32876 );
and \U$32891 ( \32884 , \32882 , \32883 );
nor \U$32892 ( \32885 , \32881 , \32884 );
buf \U$32893 ( \32886 , \32885 );
buf \U$32894 ( \32887 , \32886 );
xor \U$32895 ( \32888 , \29764 , \29770 );
and \U$32896 ( \32889 , \32888 , \30336 );
and \U$32897 ( \32890 , \29764 , \29770 );
or \U$32898 ( \32891 , \32889 , \32890 );
buf \U$32899 ( \32892 , \32891 );
buf \U$32900 ( \32893 , \32892 );
xor \U$32901 ( \32894 , \32887 , \32893 );
buf \U$32902 ( \32895 , \30325 );
not \U$32903 ( \32896 , \32895 );
buf \U$32904 ( \32897 , \30156 );
not \U$32905 ( \32898 , \32897 );
or \U$32906 ( \32899 , \32896 , \32898 );
buf \U$32907 ( \32900 , \29951 );
nand \U$32908 ( \32901 , \32899 , \32900 );
buf \U$32909 ( \32902 , \32901 );
buf \U$32910 ( \32903 , \32902 );
buf \U$32911 ( \32904 , \30156 );
not \U$32912 ( \32905 , \32904 );
buf \U$32913 ( \32906 , \30331 );
nand \U$32914 ( \32907 , \32905 , \32906 );
buf \U$32915 ( \32908 , \32907 );
buf \U$32916 ( \32909 , \32908 );
nand \U$32917 ( \32910 , \32903 , \32909 );
buf \U$32918 ( \32911 , \32910 );
buf \U$32919 ( \32912 , \32911 );
buf \U$32920 ( \32913 , \29944 );
not \U$32921 ( \32914 , \32913 );
buf \U$32922 ( \32915 , \29876 );
not \U$32923 ( \32916 , \32915 );
or \U$32924 ( \32917 , \32914 , \32916 );
not \U$32925 ( \32918 , \29941 );
not \U$32926 ( \32919 , \29879 );
or \U$32927 ( \32920 , \32918 , \32919 );
nand \U$32928 ( \32921 , \32920 , \29824 );
buf \U$32929 ( \32922 , \32921 );
nand \U$32930 ( \32923 , \32917 , \32922 );
buf \U$32931 ( \32924 , \32923 );
buf \U$32932 ( \32925 , \32924 );
buf \U$32933 ( \32926 , \30007 );
not \U$32934 ( \32927 , \32926 );
buf \U$32935 ( \32928 , \30152 );
not \U$32936 ( \32929 , \32928 );
or \U$32937 ( \32930 , \32927 , \32929 );
buf \U$32938 ( \32931 , \30010 );
not \U$32939 ( \32932 , \32931 );
buf \U$32940 ( \32933 , \30146 );
not \U$32941 ( \32934 , \32933 );
or \U$32942 ( \32935 , \32932 , \32934 );
buf \U$32943 ( \32936 , \30079 );
not \U$32944 ( \32937 , \32936 );
buf \U$32945 ( \32938 , \32937 );
buf \U$32946 ( \32939 , \32938 );
nand \U$32947 ( \32940 , \32935 , \32939 );
buf \U$32948 ( \32941 , \32940 );
buf \U$32949 ( \32942 , \32941 );
nand \U$32950 ( \32943 , \32930 , \32942 );
buf \U$32951 ( \32944 , \32943 );
buf \U$32952 ( \32945 , \32944 );
xor \U$32953 ( \32946 , \32925 , \32945 );
buf \U$32954 ( \32947 , \30315 );
not \U$32955 ( \32948 , \32947 );
buf \U$32956 ( \32949 , \30270 );
not \U$32957 ( \32950 , \32949 );
buf \U$32958 ( \32951 , \32950 );
buf \U$32959 ( \32952 , \32951 );
not \U$32960 ( \32953 , \32952 );
or \U$32961 ( \32954 , \32948 , \32953 );
buf \U$32962 ( \32955 , \30318 );
not \U$32963 ( \32956 , \32955 );
buf \U$32964 ( \32957 , \30270 );
not \U$32965 ( \32958 , \32957 );
or \U$32966 ( \32959 , \32956 , \32958 );
buf \U$32967 ( \32960 , \30218 );
nand \U$32968 ( \32961 , \32959 , \32960 );
buf \U$32969 ( \32962 , \32961 );
buf \U$32970 ( \32963 , \32962 );
nand \U$32971 ( \32964 , \32954 , \32963 );
buf \U$32972 ( \32965 , \32964 );
buf \U$32973 ( \32966 , \32965 );
xor \U$32974 ( \32967 , \32946 , \32966 );
buf \U$32975 ( \32968 , \32967 );
buf \U$32976 ( \32969 , \32968 );
xor \U$32977 ( \32970 , \32912 , \32969 );
xor \U$32978 ( \32971 , \29843 , \29861 );
and \U$32979 ( \32972 , \32971 , \29874 );
and \U$32980 ( \32973 , \29843 , \29861 );
or \U$32981 ( \32974 , \32972 , \32973 );
buf \U$32982 ( \32975 , \32974 );
buf \U$32983 ( \32976 , \30145 );
not \U$32984 ( \32977 , \32976 );
buf \U$32985 ( \32978 , \30122 );
not \U$32986 ( \32979 , \32978 );
or \U$32987 ( \32980 , \32977 , \32979 );
buf \U$32988 ( \32981 , \30142 );
not \U$32989 ( \32982 , \32981 );
buf \U$32990 ( \32983 , \30125 );
not \U$32991 ( \32984 , \32983 );
or \U$32992 ( \32985 , \32982 , \32984 );
buf \U$32993 ( \32986 , \30106 );
nand \U$32994 ( \32987 , \32985 , \32986 );
buf \U$32995 ( \32988 , \32987 );
buf \U$32996 ( \32989 , \32988 );
nand \U$32997 ( \32990 , \32980 , \32989 );
buf \U$32998 ( \32991 , \32990 );
xor \U$32999 ( \32992 , \32975 , \32991 );
buf \U$33000 ( \32993 , \32992 );
buf \U$33001 ( \32994 , \30289 );
not \U$33002 ( \32995 , \32994 );
buf \U$33003 ( \32996 , \4907 );
not \U$33004 ( \32997 , \32996 );
or \U$33005 ( \32998 , \32995 , \32997 );
buf \U$33006 ( \32999 , \686 );
xor \U$33007 ( \33000 , RIc0d9568_67, RIc0d8b90_46);
buf \U$33008 ( \33001 , \33000 );
nand \U$33009 ( \33002 , \32999 , \33001 );
buf \U$33010 ( \33003 , \33002 );
buf \U$33011 ( \33004 , \33003 );
nand \U$33012 ( \33005 , \32998 , \33004 );
buf \U$33013 ( \33006 , \33005 );
buf \U$33014 ( \33007 , \33006 );
buf \U$33015 ( \33008 , \30116 );
not \U$33016 ( \33009 , \33008 );
buf \U$33017 ( \33010 , \2871 );
not \U$33018 ( \33011 , \33010 );
or \U$33019 ( \33012 , \33009 , \33011 );
buf \U$33020 ( \33013 , \1856 );
buf \U$33021 ( \33014 , RIc0d9838_73);
buf \U$33022 ( \33015 , RIc0d88c0_40);
xor \U$33023 ( \33016 , \33014 , \33015 );
buf \U$33024 ( \33017 , \33016 );
buf \U$33025 ( \33018 , \33017 );
nand \U$33026 ( \33019 , \33013 , \33018 );
buf \U$33027 ( \33020 , \33019 );
buf \U$33028 ( \33021 , \33020 );
nand \U$33029 ( \33022 , \33012 , \33021 );
buf \U$33030 ( \33023 , \33022 );
buf \U$33031 ( \33024 , \33023 );
xor \U$33032 ( \33025 , \33007 , \33024 );
buf \U$33033 ( \33026 , \30308 );
not \U$33034 ( \33027 , \33026 );
buf \U$33035 ( \33028 , \33027 );
buf \U$33036 ( \33029 , \33028 );
not \U$33037 ( \33030 , \33029 );
buf \U$33038 ( \33031 , \2535 );
not \U$33039 ( \33032 , \33031 );
or \U$33040 ( \33033 , \33030 , \33032 );
buf \U$33041 ( \33034 , \714 );
buf \U$33042 ( \33035 , RIc0d8050_22);
buf \U$33043 ( \33036 , RIc0da0a8_91);
xor \U$33044 ( \33037 , \33035 , \33036 );
buf \U$33045 ( \33038 , \33037 );
buf \U$33046 ( \33039 , \33038 );
nand \U$33047 ( \33040 , \33034 , \33039 );
buf \U$33048 ( \33041 , \33040 );
buf \U$33049 ( \33042 , \33041 );
nand \U$33050 ( \33043 , \33033 , \33042 );
buf \U$33051 ( \33044 , \33043 );
buf \U$33052 ( \33045 , \33044 );
xor \U$33053 ( \33046 , \33025 , \33045 );
buf \U$33054 ( \33047 , \33046 );
buf \U$33055 ( \33048 , \33047 );
xnor \U$33056 ( \33049 , \32993 , \33048 );
buf \U$33057 ( \33050 , \33049 );
buf \U$33058 ( \33051 , \33050 );
not \U$33059 ( \33052 , \33051 );
xor \U$33060 ( \33053 , \29970 , \29987 );
and \U$33061 ( \33054 , \33053 , \30005 );
and \U$33062 ( \33055 , \29970 , \29987 );
or \U$33063 ( \33056 , \33054 , \33055 );
buf \U$33064 ( \33057 , \33056 );
buf \U$33065 ( \33058 , \30043 );
not \U$33066 ( \33059 , \33058 );
buf \U$33067 ( \33060 , \30075 );
not \U$33068 ( \33061 , \33060 );
or \U$33069 ( \33062 , \33059 , \33061 );
buf \U$33070 ( \33063 , \30069 );
not \U$33071 ( \33064 , \33063 );
buf \U$33072 ( \33065 , \30046 );
not \U$33073 ( \33066 , \33065 );
or \U$33074 ( \33067 , \33064 , \33066 );
buf \U$33075 ( \33068 , \30028 );
nand \U$33076 ( \33069 , \33067 , \33068 );
buf \U$33077 ( \33070 , \33069 );
buf \U$33078 ( \33071 , \33070 );
nand \U$33079 ( \33072 , \33062 , \33071 );
buf \U$33080 ( \33073 , \33072 );
buf \U$33081 ( \33074 , \33073 );
not \U$33082 ( \33075 , \33074 );
buf \U$33083 ( \33076 , \33075 );
xor \U$33084 ( \33077 , \33057 , \33076 );
buf \U$33085 ( \33078 , \29906 );
not \U$33086 ( \33079 , \33078 );
buf \U$33087 ( \33080 , \29922 );
not \U$33088 ( \33081 , \33080 );
or \U$33089 ( \33082 , \33079 , \33081 );
buf \U$33090 ( \33083 , \29922 );
buf \U$33091 ( \33084 , \29906 );
or \U$33092 ( \33085 , \33083 , \33084 );
buf \U$33093 ( \33086 , \29940 );
nand \U$33094 ( \33087 , \33085 , \33086 );
buf \U$33095 ( \33088 , \33087 );
buf \U$33096 ( \33089 , \33088 );
nand \U$33097 ( \33090 , \33082 , \33089 );
buf \U$33098 ( \33091 , \33090 );
xor \U$33099 ( \33092 , \33077 , \33091 );
buf \U$33100 ( \33093 , \33092 );
not \U$33101 ( \33094 , \33093 );
buf \U$33102 ( \33095 , \33094 );
buf \U$33103 ( \33096 , \33095 );
not \U$33104 ( \33097 , \33096 );
or \U$33105 ( \33098 , \33052 , \33097 );
buf \U$33106 ( \33099 , \33092 );
buf \U$33107 ( \33100 , \33050 );
not \U$33108 ( \33101 , \33100 );
buf \U$33109 ( \33102 , \33101 );
buf \U$33110 ( \33103 , \33102 );
nand \U$33111 ( \33104 , \33099 , \33103 );
buf \U$33112 ( \33105 , \33104 );
buf \U$33113 ( \33106 , \33105 );
nand \U$33114 ( \33107 , \33098 , \33106 );
buf \U$33115 ( \33108 , \33107 );
buf \U$33116 ( \33109 , \33108 );
buf \U$33117 ( \33110 , \29814 );
not \U$33118 ( \33111 , \33110 );
buf \U$33119 ( \33112 , \4692 );
not \U$33120 ( \33113 , \33112 );
or \U$33121 ( \33114 , \33111 , \33113 );
buf \U$33122 ( \33115 , \284 );
buf \U$33123 ( \33116 , RIc0d8aa0_44);
buf \U$33124 ( \33117 , RIc0d9658_69);
xor \U$33125 ( \33118 , \33116 , \33117 );
buf \U$33126 ( \33119 , \33118 );
buf \U$33127 ( \33120 , \33119 );
nand \U$33128 ( \33121 , \33115 , \33120 );
buf \U$33129 ( \33122 , \33121 );
buf \U$33130 ( \33123 , \33122 );
nand \U$33131 ( \33124 , \33114 , \33123 );
buf \U$33132 ( \33125 , \33124 );
buf \U$33133 ( \33126 , \33125 );
not \U$33134 ( \33127 , \33126 );
buf \U$33135 ( \33128 , \14532 );
not \U$33136 ( \33129 , \33128 );
buf \U$33137 ( \33130 , \33129 );
buf \U$33138 ( \33131 , \33130 );
not \U$33139 ( \33132 , \33131 );
buf \U$33140 ( \33133 , \29852 );
not \U$33141 ( \33134 , \33133 );
and \U$33142 ( \33135 , \33132 , \33134 );
buf \U$33143 ( \33136 , RIc0d9bf8_81);
buf \U$33144 ( \33137 , RIc0d8500_32);
xor \U$33145 ( \33138 , \33136 , \33137 );
buf \U$33146 ( \33139 , \33138 );
buf \U$33147 ( \33140 , \33139 );
not \U$33148 ( \33141 , \33140 );
buf \U$33149 ( \33142 , \2775 );
nor \U$33150 ( \33143 , \33141 , \33142 );
buf \U$33151 ( \33144 , \33143 );
buf \U$33152 ( \33145 , \33144 );
nor \U$33153 ( \33146 , \33135 , \33145 );
buf \U$33154 ( \33147 , \33146 );
buf \U$33155 ( \33148 , \33147 );
not \U$33156 ( \33149 , \33148 );
or \U$33157 ( \33150 , \33127 , \33149 );
buf \U$33158 ( \33151 , \33147 );
not \U$33159 ( \33152 , \33151 );
buf \U$33160 ( \33153 , \33152 );
buf \U$33161 ( \33154 , \33153 );
buf \U$33162 ( \33155 , \33125 );
not \U$33163 ( \33156 , \33155 );
buf \U$33164 ( \33157 , \33156 );
buf \U$33165 ( \33158 , \33157 );
nand \U$33166 ( \33159 , \33154 , \33158 );
buf \U$33167 ( \33160 , \33159 );
buf \U$33168 ( \33161 , \33160 );
nand \U$33169 ( \33162 , \33150 , \33161 );
buf \U$33170 ( \33163 , \33162 );
buf \U$33171 ( \33164 , \33163 );
buf \U$33172 ( \33165 , \1588 );
not \U$33173 ( \33166 , \33165 );
buf \U$33174 ( \33167 , RIc0d86e0_36);
buf \U$33175 ( \33168 , RIc0d9a18_77);
xor \U$33176 ( \33169 , \33167 , \33168 );
buf \U$33177 ( \33170 , \33169 );
buf \U$33178 ( \33171 , \33170 );
not \U$33179 ( \33172 , \33171 );
or \U$33180 ( \33173 , \33166 , \33172 );
buf \U$33181 ( \33174 , \5019 );
buf \U$33182 ( \33175 , \29932 );
or \U$33183 ( \33176 , \33174 , \33175 );
nand \U$33184 ( \33177 , \33173 , \33176 );
buf \U$33185 ( \33178 , \33177 );
buf \U$33186 ( \33179 , \33178 );
xnor \U$33187 ( \33180 , \33164 , \33179 );
buf \U$33188 ( \33181 , \33180 );
buf \U$33189 ( \33182 , \33181 );
not \U$33190 ( \33183 , \33182 );
buf \U$33191 ( \33184 , \30065 );
not \U$33192 ( \33185 , \33184 );
buf \U$33193 ( \33186 , \2399 );
not \U$33194 ( \33187 , \33186 );
or \U$33195 ( \33188 , \33185 , \33187 );
buf \U$33196 ( \33189 , \2960 );
buf \U$33197 ( \33190 , RIc0d8320_28);
buf \U$33198 ( \33191 , RIc0d9dd8_85);
xor \U$33199 ( \33192 , \33190 , \33191 );
buf \U$33200 ( \33193 , \33192 );
buf \U$33201 ( \33194 , \33193 );
nand \U$33202 ( \33195 , \33189 , \33194 );
buf \U$33203 ( \33196 , \33195 );
buf \U$33204 ( \33197 , \33196 );
nand \U$33205 ( \33198 , \33188 , \33197 );
buf \U$33206 ( \33199 , \33198 );
buf \U$33207 ( \33200 , \33199 );
not \U$33208 ( \33201 , \33200 );
buf \U$33209 ( \33202 , \33201 );
buf \U$33210 ( \33203 , \33202 );
not \U$33211 ( \33204 , \33203 );
buf \U$33212 ( \33205 , \29980 );
not \U$33213 ( \33206 , \33205 );
buf \U$33214 ( \33207 , \476 );
not \U$33215 ( \33208 , \33207 );
or \U$33216 ( \33209 , \33206 , \33208 );
buf \U$33217 ( \33210 , \4008 );
xor \U$33218 ( \33211 , RIc0da198_93, RIc0d7f60_20);
buf \U$33219 ( \33212 , \33211 );
nand \U$33220 ( \33213 , \33210 , \33212 );
buf \U$33221 ( \33214 , \33213 );
buf \U$33222 ( \33215 , \33214 );
nand \U$33223 ( \33216 , \33209 , \33215 );
buf \U$33224 ( \33217 , \33216 );
buf \U$33225 ( \33218 , \33217 );
not \U$33226 ( \33219 , \33218 );
buf \U$33227 ( \33220 , \29916 );
not \U$33228 ( \33221 , \33220 );
buf \U$33229 ( \33222 , \14888 );
not \U$33230 ( \33223 , \33222 );
buf \U$33231 ( \33224 , \33223 );
buf \U$33232 ( \33225 , \33224 );
not \U$33233 ( \33226 , \33225 );
or \U$33234 ( \33227 , \33221 , \33226 );
buf \U$33235 ( \33228 , \12410 );
buf \U$33236 ( \33229 , RIc0daaf8_113);
nand \U$33237 ( \33230 , \33228 , \33229 );
buf \U$33238 ( \33231 , \33230 );
buf \U$33239 ( \33232 , \33231 );
nand \U$33240 ( \33233 , \33227 , \33232 );
buf \U$33241 ( \33234 , \33233 );
buf \U$33242 ( \33235 , \33234 );
not \U$33243 ( \33236 , \33235 );
buf \U$33244 ( \33237 , \33236 );
buf \U$33245 ( \33238 , \33237 );
not \U$33246 ( \33239 , \33238 );
or \U$33247 ( \33240 , \33219 , \33239 );
buf \U$33248 ( \33241 , \33237 );
buf \U$33249 ( \33242 , \33217 );
or \U$33250 ( \33243 , \33241 , \33242 );
nand \U$33251 ( \33244 , \33240 , \33243 );
buf \U$33252 ( \33245 , \33244 );
buf \U$33253 ( \33246 , \33245 );
not \U$33254 ( \33247 , \33246 );
or \U$33255 ( \33248 , \33204 , \33247 );
buf \U$33256 ( \33249 , \33245 );
buf \U$33257 ( \33250 , \33202 );
or \U$33258 ( \33251 , \33249 , \33250 );
nand \U$33259 ( \33252 , \33248 , \33251 );
buf \U$33260 ( \33253 , \33252 );
buf \U$33261 ( \33254 , \33253 );
not \U$33262 ( \33255 , \33254 );
buf \U$33263 ( \33256 , \30100 );
not \U$33264 ( \33257 , \33256 );
buf \U$33267 ( \33258 , \12833 );
buf \U$33268 ( \33259 , \33258 );
not \U$33269 ( \33260 , \33259 );
or \U$33270 ( \33261 , \33257 , \33260 );
buf \U$33271 ( \33262 , \16676 );
xor \U$33272 ( \33263 , RIc0da558_101, RIc0d7ba0_12);
buf \U$33273 ( \33264 , \33263 );
nand \U$33274 ( \33265 , \33262 , \33264 );
buf \U$33275 ( \33266 , \33265 );
buf \U$33276 ( \33267 , \33266 );
nand \U$33277 ( \33268 , \33261 , \33267 );
buf \U$33278 ( \33269 , \33268 );
buf \U$33279 ( \33270 , \33269 );
not \U$33280 ( \33271 , \33270 );
buf \U$33281 ( \33272 , \30230 );
not \U$33282 ( \33273 , \33272 );
buf \U$33283 ( \33274 , \330 );
not \U$33284 ( \33275 , \33274 );
or \U$33285 ( \33276 , \33273 , \33275 );
buf \U$33286 ( \33277 , \14707 );
buf \U$33287 ( \33278 , RIc0da288_95);
buf \U$33288 ( \33279 , RIc0d7e70_18);
xor \U$33289 ( \33280 , \33278 , \33279 );
buf \U$33290 ( \33281 , \33280 );
buf \U$33291 ( \33282 , \33281 );
nand \U$33292 ( \33283 , \33277 , \33282 );
buf \U$33293 ( \33284 , \33283 );
buf \U$33294 ( \33285 , \33284 );
nand \U$33295 ( \33286 , \33276 , \33285 );
buf \U$33296 ( \33287 , \33286 );
buf \U$33297 ( \33288 , \33287 );
not \U$33298 ( \33289 , \33288 );
buf \U$33299 ( \33290 , \33289 );
buf \U$33300 ( \33291 , \33290 );
not \U$33301 ( \33292 , \33291 );
or \U$33302 ( \33293 , \33271 , \33292 );
buf \U$33303 ( \33294 , \33290 );
buf \U$33304 ( \33295 , \33269 );
or \U$33305 ( \33296 , \33294 , \33295 );
nand \U$33306 ( \33297 , \33293 , \33296 );
buf \U$33307 ( \33298 , \33297 );
buf \U$33308 ( \33299 , \33298 );
not \U$33309 ( \33300 , \33299 );
buf \U$33310 ( \33301 , \14346 );
not \U$33311 ( \33302 , \33301 );
buf \U$33312 ( \33303 , \33302 );
buf \U$33313 ( \33304 , \33303 );
not \U$33314 ( \33305 , \33304 );
buf \U$33315 ( \33306 , \30037 );
not \U$33316 ( \33307 , \33306 );
buf \U$33317 ( \33308 , \33307 );
buf \U$33318 ( \33309 , \33308 );
not \U$33319 ( \33310 , \33309 );
and \U$33320 ( \33311 , \33305 , \33310 );
buf \U$33321 ( \33312 , \14353 );
buf \U$33322 ( \33313 , RIc0d76f0_2);
buf \U$33323 ( \33314 , RIc0daa08_111);
xor \U$33324 ( \33315 , \33313 , \33314 );
buf \U$33325 ( \33316 , \33315 );
buf \U$33326 ( \33317 , \33316 );
and \U$33327 ( \33318 , \33312 , \33317 );
buf \U$33328 ( \33319 , \33318 );
buf \U$33329 ( \33320 , \33319 );
nor \U$33330 ( \33321 , \33311 , \33320 );
buf \U$33331 ( \33322 , \33321 );
buf \U$33334 ( \33323 , \33322 );
buf \U$33335 ( \33324 , \33323 );
not \U$33336 ( \33325 , \33324 );
and \U$33337 ( \33326 , \33300 , \33325 );
buf \U$33338 ( \33327 , \33298 );
buf \U$33339 ( \33328 , \33323 );
and \U$33340 ( \33329 , \33327 , \33328 );
nor \U$33341 ( \33330 , \33326 , \33329 );
buf \U$33342 ( \33331 , \33330 );
buf \U$33343 ( \33332 , \33331 );
not \U$33344 ( \33333 , \33332 );
or \U$33345 ( \33334 , \33255 , \33333 );
buf \U$33346 ( \33335 , \33331 );
buf \U$33347 ( \33336 , \33253 );
or \U$33348 ( \33337 , \33335 , \33336 );
nand \U$33349 ( \33338 , \33334 , \33337 );
buf \U$33350 ( \33339 , \33338 );
buf \U$33351 ( \33340 , \33339 );
not \U$33352 ( \33341 , \33340 );
or \U$33353 ( \33342 , \33183 , \33341 );
buf \U$33354 ( \33343 , \33339 );
buf \U$33355 ( \33344 , \33181 );
or \U$33356 ( \33345 , \33343 , \33344 );
nand \U$33357 ( \33346 , \33342 , \33345 );
buf \U$33358 ( \33347 , \33346 );
buf \U$33359 ( \33348 , \33347 );
xor \U$33360 ( \33349 , \33109 , \33348 );
buf \U$33361 ( \33350 , \33349 );
buf \U$33362 ( \33351 , \33350 );
xor \U$33363 ( \33352 , \32970 , \33351 );
buf \U$33364 ( \33353 , \33352 );
buf \U$33365 ( \33354 , \33353 );
xor \U$33366 ( \33355 , \32894 , \33354 );
buf \U$33367 ( \33356 , \33355 );
buf \U$33368 ( \33357 , \32548 );
not \U$33369 ( \33358 , \33357 );
buf \U$33370 ( \33359 , \32606 );
not \U$33371 ( \33360 , \33359 );
or \U$33372 ( \33361 , \33358 , \33360 );
buf \U$33373 ( \33362 , \32606 );
buf \U$33374 ( \33363 , \32548 );
or \U$33375 ( \33364 , \33362 , \33363 );
not \U$33376 ( \33365 , \32592 );
buf \U$33377 ( \33366 , \33365 );
nand \U$33378 ( \33367 , \33364 , \33366 );
buf \U$33379 ( \33368 , \33367 );
buf \U$33380 ( \33369 , \33368 );
nand \U$33381 ( \33370 , \33361 , \33369 );
buf \U$33382 ( \33371 , \33370 );
buf \U$33383 ( \33372 , \33371 );
not \U$33384 ( \33373 , \33372 );
xor \U$33385 ( \33374 , \32555 , \32561 );
and \U$33386 ( \33375 , \33374 , \32589 );
and \U$33387 ( \33376 , \32555 , \32561 );
or \U$33388 ( \33377 , \33375 , \33376 );
buf \U$33389 ( \33378 , \33377 );
buf \U$33390 ( \33379 , \33378 );
buf \U$33391 ( \33380 , \30189 );
not \U$33392 ( \33381 , \33380 );
buf \U$33393 ( \33382 , \12795 );
not \U$33394 ( \33383 , \33382 );
or \U$33395 ( \33384 , \33381 , \33383 );
buf \U$33396 ( \33385 , \1229 );
xor \U$33397 ( \33386 , RIc0d9478_65, RIc0d8c80_48);
buf \U$33398 ( \33387 , \33386 );
nand \U$33399 ( \33388 , \33385 , \33387 );
buf \U$33400 ( \33389 , \33388 );
buf \U$33401 ( \33390 , \33389 );
nand \U$33402 ( \33391 , \33384 , \33390 );
buf \U$33403 ( \33392 , \33391 );
buf \U$33404 ( \33393 , \33392 );
buf \U$33405 ( \33394 , \29963 );
not \U$33406 ( \33395 , \33394 );
buf \U$33407 ( \33396 , \1351 );
not \U$33408 ( \33397 , \33396 );
or \U$33409 ( \33398 , \33395 , \33397 );
buf \U$33410 ( \33399 , \1025 );
xor \U$33411 ( \33400 , RIc0d9b08_79, RIc0d85f0_34);
buf \U$33412 ( \33401 , \33400 );
nand \U$33413 ( \33402 , \33399 , \33401 );
buf \U$33414 ( \33403 , \33402 );
buf \U$33415 ( \33404 , \33403 );
nand \U$33416 ( \33405 , \33398 , \33404 );
buf \U$33417 ( \33406 , \33405 );
buf \U$33418 ( \33407 , \33406 );
xor \U$33419 ( \33408 , \33393 , \33407 );
buf \U$33420 ( \33409 , \30246 );
not \U$33421 ( \33410 , \33409 );
buf \U$33422 ( \33411 , \29546 );
not \U$33423 ( \33412 , \33411 );
or \U$33424 ( \33413 , \33410 , \33412 );
buf \U$33425 ( \33414 , \20243 );
buf \U$33426 ( \33415 , RIc0d7ab0_10);
buf \U$33427 ( \33416 , RIc0da648_103);
xor \U$33428 ( \33417 , \33415 , \33416 );
buf \U$33429 ( \33418 , \33417 );
buf \U$33430 ( \33419 , \33418 );
nand \U$33431 ( \33420 , \33414 , \33419 );
buf \U$33432 ( \33421 , \33420 );
buf \U$33433 ( \33422 , \33421 );
nand \U$33434 ( \33423 , \33413 , \33422 );
buf \U$33435 ( \33424 , \33423 );
buf \U$33436 ( \33425 , \33424 );
xor \U$33437 ( \33426 , \33408 , \33425 );
buf \U$33438 ( \33427 , \33426 );
buf \U$33439 ( \33428 , \33427 );
buf \U$33440 ( \33429 , \30022 );
not \U$33441 ( \33430 , \33429 );
buf \U$33442 ( \33431 , \2470 );
not \U$33443 ( \33432 , \33431 );
or \U$33444 ( \33433 , \33430 , \33432 );
buf \U$33445 ( \33434 , \14140 );
buf \U$33446 ( \33435 , RIc0da468_99);
buf \U$33447 ( \33436 , RIc0d7c90_14);
xor \U$33448 ( \33437 , \33435 , \33436 );
buf \U$33449 ( \33438 , \33437 );
buf \U$33450 ( \33439 , \33438 );
nand \U$33451 ( \33440 , \33434 , \33439 );
buf \U$33452 ( \33441 , \33440 );
buf \U$33453 ( \33442 , \33441 );
nand \U$33454 ( \33443 , \33433 , \33442 );
buf \U$33455 ( \33444 , \33443 );
buf \U$33456 ( \33445 , \29836 );
not \U$33457 ( \33446 , \33445 );
buf \U$33458 ( \33447 , \18150 );
not \U$33459 ( \33448 , \33447 );
or \U$33460 ( \33449 , \33446 , \33448 );
buf \U$33461 ( \33450 , \16477 );
buf \U$33462 ( \33451 , RIc0d9fb8_89);
buf \U$33463 ( \33452 , RIc0d8140_24);
xor \U$33464 ( \33453 , \33451 , \33452 );
buf \U$33465 ( \33454 , \33453 );
buf \U$33466 ( \33455 , \33454 );
nand \U$33467 ( \33456 , \33450 , \33455 );
buf \U$33468 ( \33457 , \33456 );
buf \U$33469 ( \33458 , \33457 );
nand \U$33470 ( \33459 , \33449 , \33458 );
buf \U$33471 ( \33460 , \33459 );
xor \U$33472 ( \33461 , \33444 , \33460 );
buf \U$33473 ( \33462 , \30172 );
not \U$33474 ( \33463 , \33462 );
buf \U$33475 ( \33464 , \1888 );
not \U$33476 ( \33465 , \33464 );
or \U$33477 ( \33466 , \33463 , \33465 );
buf \U$33478 ( \33467 , \1282 );
buf \U$33479 ( \33468 , RIc0d9748_71);
buf \U$33480 ( \33469 , RIc0d89b0_42);
xor \U$33481 ( \33470 , \33468 , \33469 );
buf \U$33482 ( \33471 , \33470 );
buf \U$33483 ( \33472 , \33471 );
nand \U$33484 ( \33473 , \33467 , \33472 );
buf \U$33485 ( \33474 , \33473 );
buf \U$33486 ( \33475 , \33474 );
nand \U$33487 ( \33476 , \33466 , \33475 );
buf \U$33488 ( \33477 , \33476 );
xor \U$33489 ( \33478 , \33461 , \33477 );
buf \U$33490 ( \33479 , \33478 );
xor \U$33491 ( \33480 , \33428 , \33479 );
buf \U$33492 ( \33481 , \30263 );
not \U$33493 ( \33482 , \33481 );
buf \U$33494 ( \33483 , \12736 );
not \U$33495 ( \33484 , \33483 );
or \U$33496 ( \33485 , \33482 , \33484 );
buf \U$33497 ( \33486 , \21880 );
buf \U$33498 ( \33487 , RIc0da738_105);
buf \U$33499 ( \33488 , RIc0d79c0_8);
xor \U$33500 ( \33489 , \33487 , \33488 );
buf \U$33501 ( \33490 , \33489 );
buf \U$33502 ( \33491 , \33490 );
nand \U$33503 ( \33492 , \33486 , \33491 );
buf \U$33504 ( \33493 , \33492 );
buf \U$33505 ( \33494 , \33493 );
nand \U$33506 ( \33495 , \33485 , \33494 );
buf \U$33507 ( \33496 , \33495 );
buf \U$33508 ( \33497 , \29781 );
not \U$33509 ( \33498 , \33497 );
buf \U$33510 ( \33499 , \28794 );
not \U$33511 ( \33500 , \33499 );
or \U$33512 ( \33501 , \33498 , \33500 );
buf \U$33513 ( \33502 , \16071 );
buf \U$33514 ( \33503 , RIc0d78d0_6);
buf \U$33515 ( \33504 , RIc0da828_107);
xor \U$33516 ( \33505 , \33503 , \33504 );
buf \U$33517 ( \33506 , \33505 );
buf \U$33518 ( \33507 , \33506 );
nand \U$33519 ( \33508 , \33502 , \33507 );
buf \U$33520 ( \33509 , \33508 );
buf \U$33521 ( \33510 , \33509 );
nand \U$33522 ( \33511 , \33501 , \33510 );
buf \U$33523 ( \33512 , \33511 );
xor \U$33524 ( \33513 , \33496 , \33512 );
buf \U$33525 ( \33514 , \10443 );
buf \U$33526 ( \33515 , \29900 );
not \U$33527 ( \33516 , \33515 );
buf \U$33528 ( \33517 , \33516 );
buf \U$33529 ( \33518 , \33517 );
or \U$33530 ( \33519 , \33514 , \33518 );
buf \U$33531 ( \33520 , \1370 );
xor \U$33532 ( \33521 , RIc0d9928_75, RIc0d87d0_38);
buf \U$33533 ( \33522 , \33521 );
not \U$33534 ( \33523 , \33522 );
buf \U$33535 ( \33524 , \33523 );
buf \U$33536 ( \33525 , \33524 );
or \U$33537 ( \33526 , \33520 , \33525 );
nand \U$33538 ( \33527 , \33519 , \33526 );
buf \U$33539 ( \33528 , \33527 );
xor \U$33540 ( \33529 , \33513 , \33528 );
buf \U$33541 ( \33530 , \33529 );
xor \U$33542 ( \33531 , \33480 , \33530 );
buf \U$33543 ( \33532 , \33531 );
buf \U$33544 ( \33533 , \33532 );
xor \U$33545 ( \33534 , \32568 , \32574 );
and \U$33546 ( \33535 , \33534 , \32586 );
and \U$33547 ( \33536 , \32568 , \32574 );
or \U$33548 ( \33537 , \33535 , \33536 );
buf \U$33549 ( \33538 , \33537 );
buf \U$33550 ( \33539 , \33538 );
xor \U$33551 ( \33540 , \33533 , \33539 );
buf \U$33552 ( \33541 , \28887 );
buf \U$33553 ( \33542 , \29163 );
or \U$33554 ( \33543 , \33541 , \33542 );
buf \U$33555 ( \33544 , \29062 );
nand \U$33556 ( \33545 , \33543 , \33544 );
buf \U$33557 ( \33546 , \33545 );
buf \U$33558 ( \33547 , \33546 );
buf \U$33559 ( \33548 , \29163 );
buf \U$33560 ( \33549 , \28887 );
nand \U$33561 ( \33550 , \33548 , \33549 );
buf \U$33562 ( \33551 , \33550 );
buf \U$33563 ( \33552 , \33551 );
nand \U$33564 ( \33553 , \33547 , \33552 );
buf \U$33565 ( \33554 , \33553 );
buf \U$33566 ( \33555 , \33554 );
xor \U$33567 ( \33556 , \33540 , \33555 );
buf \U$33568 ( \33557 , \33556 );
buf \U$33569 ( \33558 , \33557 );
xor \U$33570 ( \33559 , \33379 , \33558 );
xor \U$33571 ( \33560 , \28441 , \28684 );
and \U$33572 ( \33561 , \33560 , \29174 );
and \U$33573 ( \33562 , \28441 , \28684 );
or \U$33574 ( \33563 , \33561 , \33562 );
buf \U$33575 ( \33564 , \33563 );
buf \U$33576 ( \33565 , \33564 );
xor \U$33577 ( \33566 , \33559 , \33565 );
buf \U$33578 ( \33567 , \33566 );
buf \U$33579 ( \33568 , \33567 );
not \U$33580 ( \33569 , \33568 );
buf \U$33581 ( \33570 , \33569 );
buf \U$33582 ( \33571 , \33570 );
not \U$33583 ( \33572 , \33571 );
or \U$33584 ( \33573 , \33373 , \33572 );
buf \U$33585 ( \33574 , \33371 );
not \U$33586 ( \33575 , \33574 );
buf \U$33587 ( \33576 , \33567 );
nand \U$33588 ( \33577 , \33575 , \33576 );
buf \U$33589 ( \33578 , \33577 );
buf \U$33590 ( \33579 , \33578 );
nand \U$33591 ( \33580 , \33573 , \33579 );
buf \U$33592 ( \33581 , \33580 );
buf \U$33593 ( \33582 , \33581 );
xor \U$33594 ( \33583 , \29177 , \29646 );
and \U$33595 ( \33584 , \33583 , \30339 );
and \U$33596 ( \33585 , \29177 , \29646 );
or \U$33597 ( \33586 , \33584 , \33585 );
buf \U$33598 ( \33587 , \33586 );
buf \U$33599 ( \33588 , \33587 );
not \U$33600 ( \33589 , \33588 );
buf \U$33601 ( \33590 , \33589 );
buf \U$33602 ( \33591 , \33590 );
and \U$33603 ( \33592 , \33582 , \33591 );
not \U$33604 ( \33593 , \33582 );
buf \U$33605 ( \33594 , \33587 );
and \U$33606 ( \33595 , \33593 , \33594 );
nor \U$33607 ( \33596 , \33592 , \33595 );
buf \U$33608 ( \33597 , \33596 );
xor \U$33609 ( \33598 , \33356 , \33597 );
buf \U$33612 ( \33599 , \32528 );
buf \U$33613 ( \33600 , \33599 );
not \U$33614 ( \33601 , \33600 );
buf \U$33615 ( \33602 , \32628 );
not \U$33616 ( \33603 , \33602 );
or \U$33617 ( \33604 , \33601 , \33603 );
buf \U$33618 ( \33605 , \32628 );
buf \U$33619 ( \33606 , \33599 );
or \U$33620 ( \33607 , \33605 , \33606 );
buf \U$33621 ( \33608 , \32614 );
not \U$33622 ( \33609 , \33608 );
buf \U$33623 ( \33610 , \33609 );
buf \U$33624 ( \33611 , \33610 );
nand \U$33625 ( \33612 , \33607 , \33611 );
buf \U$33626 ( \33613 , \33612 );
buf \U$33627 ( \33614 , \33613 );
nand \U$33628 ( \33615 , \33604 , \33614 );
buf \U$33629 ( \33616 , \33615 );
xor \U$33630 ( \33617 , \33598 , \33616 );
buf \U$33631 ( \33618 , \33617 );
nand \U$33632 ( \33619 , \32647 , \33618 );
buf \U$33633 ( \33620 , \33619 );
buf \U$33634 ( \33621 , \33620 );
xor \U$33635 ( \33622 , \32912 , \32969 );
and \U$33636 ( \33623 , \33622 , \33351 );
and \U$33637 ( \33624 , \32912 , \32969 );
or \U$33638 ( \33625 , \33623 , \33624 );
buf \U$33639 ( \33626 , \33625 );
buf \U$33640 ( \33627 , \33626 );
not \U$33641 ( \33628 , \33627 );
buf \U$33642 ( \33629 , \32688 );
not \U$33643 ( \33630 , \33629 );
buf \U$33644 ( \33631 , \32757 );
not \U$33645 ( \33632 , \33631 );
or \U$33646 ( \33633 , \33630 , \33632 );
buf \U$33647 ( \33634 , \32691 );
not \U$33648 ( \33635 , \33634 );
buf \U$33649 ( \33636 , \32751 );
not \U$33650 ( \33637 , \33636 );
or \U$33651 ( \33638 , \33635 , \33637 );
buf \U$33652 ( \33639 , \32672 );
nand \U$33653 ( \33640 , \33638 , \33639 );
buf \U$33654 ( \33641 , \33640 );
buf \U$33655 ( \33642 , \33641 );
nand \U$33656 ( \33643 , \33633 , \33642 );
buf \U$33657 ( \33644 , \33643 );
buf \U$33658 ( \33645 , \33644 );
not \U$33659 ( \33646 , \33645 );
buf \U$33660 ( \33647 , \33646 );
buf \U$33661 ( \33648 , \33647 );
not \U$33662 ( \33649 , \33648 );
buf \U$33663 ( \33650 , \32727 );
not \U$33664 ( \33651 , \33650 );
buf \U$33665 ( \33652 , \32744 );
not \U$33666 ( \33653 , \33652 );
or \U$33667 ( \33654 , \33651 , \33653 );
buf \U$33668 ( \33655 , \32717 );
nand \U$33669 ( \33656 , \33654 , \33655 );
buf \U$33670 ( \33657 , \33656 );
buf \U$33671 ( \33658 , \33657 );
buf \U$33672 ( \33659 , \32724 );
buf \U$33673 ( \33660 , \32741 );
nand \U$33674 ( \33661 , \33659 , \33660 );
buf \U$33675 ( \33662 , \33661 );
buf \U$33676 ( \33663 , \33662 );
nand \U$33677 ( \33664 , \33658 , \33663 );
buf \U$33678 ( \33665 , \33664 );
buf \U$33679 ( \33666 , \33057 );
buf \U$33680 ( \33667 , \33091 );
or \U$33681 ( \33668 , \33666 , \33667 );
buf \U$33682 ( \33669 , \33073 );
nand \U$33683 ( \33670 , \33668 , \33669 );
buf \U$33684 ( \33671 , \33670 );
buf \U$33685 ( \33672 , \33671 );
buf \U$33686 ( \33673 , \33057 );
buf \U$33687 ( \33674 , \33091 );
nand \U$33688 ( \33675 , \33673 , \33674 );
buf \U$33689 ( \33676 , \33675 );
buf \U$33690 ( \33677 , \33676 );
nand \U$33691 ( \33678 , \33672 , \33677 );
buf \U$33692 ( \33679 , \33678 );
xor \U$33693 ( \33680 , \33665 , \33679 );
buf \U$33694 ( \33681 , \33680 );
not \U$33695 ( \33682 , \33681 );
buf \U$33696 ( \33683 , \33322 );
not \U$33697 ( \33684 , \33683 );
buf \U$33698 ( \33685 , \33290 );
not \U$33699 ( \33686 , \33685 );
or \U$33700 ( \33687 , \33684 , \33686 );
buf \U$33701 ( \33688 , \33269 );
nand \U$33702 ( \33689 , \33687 , \33688 );
buf \U$33703 ( \33690 , \33689 );
buf \U$33704 ( \33691 , \33690 );
buf \U$33705 ( \33692 , \33322 );
not \U$33706 ( \33693 , \33692 );
buf \U$33707 ( \33694 , \33287 );
nand \U$33708 ( \33695 , \33693 , \33694 );
buf \U$33709 ( \33696 , \33695 );
buf \U$33710 ( \33697 , \33696 );
nand \U$33711 ( \33698 , \33691 , \33697 );
buf \U$33712 ( \33699 , \33698 );
buf \U$33713 ( \33700 , \33699 );
buf \U$33714 ( \33701 , \33528 );
not \U$33715 ( \33702 , \33701 );
buf \U$33716 ( \33703 , \33496 );
not \U$33717 ( \33704 , \33703 );
or \U$33718 ( \33705 , \33702 , \33704 );
buf \U$33719 ( \33706 , \33496 );
buf \U$33720 ( \33707 , \33528 );
or \U$33721 ( \33708 , \33706 , \33707 );
buf \U$33722 ( \33709 , \33512 );
nand \U$33723 ( \33710 , \33708 , \33709 );
buf \U$33724 ( \33711 , \33710 );
buf \U$33725 ( \33712 , \33711 );
nand \U$33726 ( \33713 , \33705 , \33712 );
buf \U$33727 ( \33714 , \33713 );
buf \U$33728 ( \33715 , \33714 );
xor \U$33729 ( \33716 , \33700 , \33715 );
buf \U$33730 ( \33717 , \33716 );
buf \U$33731 ( \33718 , \33717 );
buf \U$33732 ( \33719 , \33023 );
buf \U$33733 ( \33720 , \33006 );
or \U$33734 ( \33721 , \33719 , \33720 );
buf \U$33735 ( \33722 , \33044 );
nand \U$33736 ( \33723 , \33721 , \33722 );
buf \U$33737 ( \33724 , \33723 );
buf \U$33738 ( \33725 , \33724 );
buf \U$33739 ( \33726 , \33023 );
buf \U$33740 ( \33727 , \33006 );
nand \U$33741 ( \33728 , \33726 , \33727 );
buf \U$33742 ( \33729 , \33728 );
buf \U$33743 ( \33730 , \33729 );
nand \U$33744 ( \33731 , \33725 , \33730 );
buf \U$33745 ( \33732 , \33731 );
buf \U$33746 ( \33733 , \33732 );
not \U$33747 ( \33734 , \33733 );
buf \U$33748 ( \33735 , \33734 );
buf \U$33749 ( \33736 , \33735 );
and \U$33750 ( \33737 , \33718 , \33736 );
not \U$33751 ( \33738 , \33718 );
buf \U$33752 ( \33739 , \33732 );
and \U$33753 ( \33740 , \33738 , \33739 );
nor \U$33754 ( \33741 , \33737 , \33740 );
buf \U$33755 ( \33742 , \33741 );
buf \U$33756 ( \33743 , \33742 );
not \U$33757 ( \33744 , \33743 );
and \U$33758 ( \33745 , \33682 , \33744 );
buf \U$33759 ( \33746 , \33680 );
buf \U$33760 ( \33747 , \33742 );
and \U$33761 ( \33748 , \33746 , \33747 );
nor \U$33762 ( \33749 , \33745 , \33748 );
buf \U$33763 ( \33750 , \33749 );
buf \U$33764 ( \33751 , \33750 );
not \U$33765 ( \33752 , \33751 );
buf \U$33766 ( \33753 , \33752 );
buf \U$33767 ( \33754 , \33753 );
not \U$33768 ( \33755 , \33754 );
or \U$33769 ( \33756 , \33649 , \33755 );
buf \U$33770 ( \33757 , \33750 );
buf \U$33771 ( \33758 , \33644 );
nand \U$33772 ( \33759 , \33757 , \33758 );
buf \U$33773 ( \33760 , \33759 );
buf \U$33774 ( \33761 , \33760 );
nand \U$33775 ( \33762 , \33756 , \33761 );
buf \U$33776 ( \33763 , \33762 );
buf \U$33777 ( \33764 , \33763 );
xor \U$33778 ( \33765 , \32925 , \32945 );
and \U$33779 ( \33766 , \33765 , \32966 );
and \U$33780 ( \33767 , \32925 , \32945 );
or \U$33781 ( \33768 , \33766 , \33767 );
buf \U$33782 ( \33769 , \33768 );
buf \U$33783 ( \33770 , \33769 );
xnor \U$33784 ( \33771 , \33764 , \33770 );
buf \U$33785 ( \33772 , \33771 );
buf \U$33786 ( \33773 , \33772 );
not \U$33787 ( \33774 , \33773 );
or \U$33788 ( \33775 , \33628 , \33774 );
buf \U$33789 ( \33776 , \33626 );
buf \U$33790 ( \33777 , \33772 );
or \U$33791 ( \33778 , \33776 , \33777 );
nand \U$33792 ( \33779 , \33775 , \33778 );
buf \U$33793 ( \33780 , \33779 );
buf \U$33794 ( \33781 , \33780 );
buf \U$33795 ( \33782 , \33102 );
not \U$33796 ( \33783 , \33782 );
buf \U$33797 ( \33784 , \33095 );
not \U$33798 ( \33785 , \33784 );
or \U$33799 ( \33786 , \33783 , \33785 );
buf \U$33800 ( \33787 , \33347 );
buf \U$33801 ( \33788 , \33092 );
buf \U$33802 ( \33789 , \33050 );
nand \U$33803 ( \33790 , \33788 , \33789 );
buf \U$33804 ( \33791 , \33790 );
buf \U$33805 ( \33792 , \33791 );
nand \U$33806 ( \33793 , \33787 , \33792 );
buf \U$33807 ( \33794 , \33793 );
buf \U$33808 ( \33795 , \33794 );
nand \U$33809 ( \33796 , \33786 , \33795 );
buf \U$33810 ( \33797 , \33796 );
buf \U$33811 ( \33798 , \33797 );
buf \U$33812 ( \33799 , \32991 );
not \U$33813 ( \33800 , \33799 );
buf \U$33814 ( \33801 , \32975 );
not \U$33815 ( \33802 , \33801 );
or \U$33816 ( \33803 , \33800 , \33802 );
buf \U$33817 ( \33804 , \32975 );
buf \U$33818 ( \33805 , \32991 );
or \U$33819 ( \33806 , \33804 , \33805 );
buf \U$33820 ( \33807 , \33047 );
nand \U$33821 ( \33808 , \33806 , \33807 );
buf \U$33822 ( \33809 , \33808 );
buf \U$33823 ( \33810 , \33809 );
nand \U$33824 ( \33811 , \33803 , \33810 );
buf \U$33825 ( \33812 , \33811 );
buf \U$33826 ( \33813 , \33812 );
buf \U$33827 ( \33814 , \32802 );
not \U$33828 ( \33815 , \33814 );
buf \U$33829 ( \33816 , \32786 );
not \U$33830 ( \33817 , \33816 );
or \U$33831 ( \33818 , \33815 , \33817 );
buf \U$33832 ( \33819 , \32802 );
buf \U$33833 ( \33820 , \32786 );
or \U$33834 ( \33821 , \33819 , \33820 );
buf \U$33835 ( \33822 , \32819 );
nand \U$33836 ( \33823 , \33821 , \33822 );
buf \U$33837 ( \33824 , \33823 );
buf \U$33838 ( \33825 , \33824 );
nand \U$33839 ( \33826 , \33818 , \33825 );
buf \U$33840 ( \33827 , \33826 );
xor \U$33841 ( \33828 , \33444 , \33460 );
and \U$33842 ( \33829 , \33828 , \33477 );
and \U$33843 ( \33830 , \33444 , \33460 );
or \U$33844 ( \33831 , \33829 , \33830 );
xor \U$33845 ( \33832 , \33827 , \33831 );
buf \U$33846 ( \33833 , \33147 );
not \U$33847 ( \33834 , \33833 );
buf \U$33848 ( \33835 , \33157 );
not \U$33849 ( \33836 , \33835 );
or \U$33850 ( \33837 , \33834 , \33836 );
buf \U$33851 ( \33838 , \33178 );
nand \U$33852 ( \33839 , \33837 , \33838 );
buf \U$33853 ( \33840 , \33839 );
buf \U$33854 ( \33841 , \33840 );
buf \U$33855 ( \33842 , \33153 );
buf \U$33856 ( \33843 , \33125 );
nand \U$33857 ( \33844 , \33842 , \33843 );
buf \U$33858 ( \33845 , \33844 );
buf \U$33859 ( \33846 , \33845 );
nand \U$33860 ( \33847 , \33841 , \33846 );
buf \U$33861 ( \33848 , \33847 );
xnor \U$33862 ( \33849 , \33832 , \33848 );
buf \U$33863 ( \33850 , \33849 );
not \U$33864 ( \33851 , \33850 );
buf \U$33865 ( \33852 , \33851 );
buf \U$33866 ( \33853 , \33852 );
xor \U$33867 ( \33854 , \33813 , \33853 );
buf \U$33868 ( \33855 , \33181 );
not \U$33869 ( \33856 , \33855 );
buf \U$33870 ( \33857 , \33331 );
not \U$33871 ( \33858 , \33857 );
or \U$33872 ( \33859 , \33856 , \33858 );
buf \U$33873 ( \33860 , \33253 );
nand \U$33874 ( \33861 , \33859 , \33860 );
buf \U$33875 ( \33862 , \33861 );
buf \U$33876 ( \33863 , \33862 );
buf \U$33877 ( \33864 , \33331 );
buf \U$33878 ( \33865 , \33181 );
or \U$33879 ( \33866 , \33864 , \33865 );
buf \U$33880 ( \33867 , \33866 );
buf \U$33881 ( \33868 , \33867 );
nand \U$33882 ( \33869 , \33863 , \33868 );
buf \U$33883 ( \33870 , \33869 );
buf \U$33884 ( \33871 , \33870 );
xor \U$33885 ( \33872 , \33854 , \33871 );
buf \U$33886 ( \33873 , \33872 );
buf \U$33887 ( \33874 , \33873 );
xor \U$33888 ( \33875 , \33798 , \33874 );
xor \U$33889 ( \33876 , \33428 , \33479 );
and \U$33890 ( \33877 , \33876 , \33530 );
and \U$33891 ( \33878 , \33428 , \33479 );
or \U$33892 ( \33879 , \33877 , \33878 );
buf \U$33893 ( \33880 , \33879 );
xor \U$33894 ( \33881 , \33393 , \33407 );
and \U$33895 ( \33882 , \33881 , \33425 );
and \U$33896 ( \33883 , \33393 , \33407 );
or \U$33897 ( \33884 , \33882 , \33883 );
buf \U$33898 ( \33885 , \33884 );
buf \U$33899 ( \33886 , \33885 );
not \U$33900 ( \33887 , \33886 );
buf \U$33901 ( \33888 , \33237 );
buf \U$33902 ( \33889 , \33202 );
nand \U$33903 ( \33890 , \33888 , \33889 );
buf \U$33904 ( \33891 , \33890 );
buf \U$33905 ( \33892 , \33891 );
buf \U$33906 ( \33893 , \33217 );
and \U$33907 ( \33894 , \33892 , \33893 );
buf \U$33908 ( \33895 , \33237 );
buf \U$33909 ( \33896 , \33202 );
nor \U$33910 ( \33897 , \33895 , \33896 );
buf \U$33911 ( \33898 , \33897 );
buf \U$33912 ( \33899 , \33898 );
nor \U$33913 ( \33900 , \33894 , \33899 );
buf \U$33914 ( \33901 , \33900 );
buf \U$33915 ( \33902 , \33901 );
not \U$33916 ( \33903 , \33902 );
or \U$33917 ( \33904 , \33887 , \33903 );
buf \U$33918 ( \33905 , \33901 );
not \U$33919 ( \33906 , \33905 );
buf \U$33920 ( \33907 , \33906 );
buf \U$33921 ( \33908 , \33907 );
buf \U$33922 ( \33909 , \33885 );
not \U$33923 ( \33910 , \33909 );
buf \U$33924 ( \33911 , \33910 );
buf \U$33925 ( \33912 , \33911 );
nand \U$33926 ( \33913 , \33908 , \33912 );
buf \U$33927 ( \33914 , \33913 );
buf \U$33928 ( \33915 , \33914 );
nand \U$33929 ( \33916 , \33904 , \33915 );
buf \U$33930 ( \33917 , \33916 );
buf \U$33931 ( \33918 , \33917 );
buf \U$33932 ( \33919 , \4868 );
not \U$33933 ( \33920 , \33919 );
buf \U$33934 ( \33921 , \33471 );
not \U$33935 ( \33922 , \33921 );
buf \U$33936 ( \33923 , \33922 );
buf \U$33937 ( \33924 , \33923 );
not \U$33938 ( \33925 , \33924 );
and \U$33939 ( \33926 , \33920 , \33925 );
buf \U$33940 ( \33927 , \1282 );
buf \U$33941 ( \33928 , RIc0d9748_71);
buf \U$33942 ( \33929 , RIc0d8938_41);
xor \U$33943 ( \33930 , \33928 , \33929 );
buf \U$33944 ( \33931 , \33930 );
buf \U$33945 ( \33932 , \33931 );
and \U$33946 ( \33933 , \33927 , \33932 );
nor \U$33947 ( \33934 , \33926 , \33933 );
buf \U$33948 ( \33935 , \33934 );
buf \U$33949 ( \33936 , \32780 );
not \U$33950 ( \33937 , \33936 );
buf \U$33951 ( \33938 , \2066 );
not \U$33952 ( \33939 , \33938 );
or \U$33953 ( \33940 , \33937 , \33939 );
buf \U$33954 ( \33941 , \734 );
xor \U$33955 ( \33942 , RIc0da378_97, RIc0d7d08_15);
buf \U$33956 ( \33943 , \33942 );
nand \U$33957 ( \33944 , \33941 , \33943 );
buf \U$33958 ( \33945 , \33944 );
buf \U$33959 ( \33946 , \33945 );
nand \U$33960 ( \33947 , \33940 , \33946 );
buf \U$33961 ( \33948 , \33947 );
xor \U$33962 ( \33949 , \33935 , \33948 );
buf \U$33963 ( \33950 , \33386 );
not \U$33964 ( \33951 , \33950 );
buf \U$33965 ( \33952 , \1224 );
not \U$33966 ( \33953 , \33952 );
or \U$33967 ( \33954 , \33951 , \33953 );
buf \U$33968 ( \33955 , \1229 );
buf \U$33969 ( \33956 , RIc0d9478_65);
buf \U$33970 ( \33957 , RIc0d8c08_47);
xor \U$33971 ( \33958 , \33956 , \33957 );
buf \U$33972 ( \33959 , \33958 );
buf \U$33973 ( \33960 , \33959 );
nand \U$33974 ( \33961 , \33955 , \33960 );
buf \U$33975 ( \33962 , \33961 );
buf \U$33976 ( \33963 , \33962 );
nand \U$33977 ( \33964 , \33954 , \33963 );
buf \U$33978 ( \33965 , \33964 );
buf \U$33979 ( \33966 , \33965 );
not \U$33980 ( \33967 , \33966 );
buf \U$33981 ( \33968 , \33967 );
xor \U$33982 ( \33969 , \33949 , \33968 );
buf \U$33983 ( \33970 , \33969 );
not \U$33984 ( \33971 , \33970 );
buf \U$33985 ( \33972 , \33971 );
buf \U$33986 ( \33973 , \33972 );
and \U$33987 ( \33974 , \33918 , \33973 );
not \U$33988 ( \33975 , \33918 );
buf \U$33989 ( \33976 , \33969 );
and \U$33990 ( \33977 , \33975 , \33976 );
nor \U$33991 ( \33978 , \33974 , \33977 );
buf \U$33992 ( \33979 , \33978 );
xor \U$33993 ( \33980 , \33880 , \33979 );
and \U$33994 ( \33981 , \30186 , \30187 );
buf \U$33995 ( \33982 , \33981 );
buf \U$33996 ( \33983 , \33982 );
buf \U$33997 ( \33984 , \33000 );
not \U$33998 ( \33985 , \33984 );
buf \U$33999 ( \33986 , \678 );
not \U$34000 ( \33987 , \33986 );
or \U$34001 ( \33988 , \33985 , \33987 );
buf \U$34002 ( \33989 , RIc0d9568_67);
buf \U$34003 ( \33990 , RIc0d8b18_45);
xnor \U$34004 ( \33991 , \33989 , \33990 );
buf \U$34005 ( \33992 , \33991 );
buf \U$34006 ( \33993 , \33992 );
not \U$34007 ( \33994 , \33993 );
buf \U$34008 ( \33995 , \686 );
nand \U$34009 ( \33996 , \33994 , \33995 );
buf \U$34010 ( \33997 , \33996 );
buf \U$34011 ( \33998 , \33997 );
nand \U$34012 ( \33999 , \33988 , \33998 );
buf \U$34013 ( \34000 , \33999 );
buf \U$34014 ( \34001 , \34000 );
xor \U$34015 ( \34002 , \33983 , \34001 );
buf \U$34016 ( \34003 , \33038 );
not \U$34017 ( \34004 , \34003 );
buf \U$34018 ( \34005 , \1927 );
not \U$34019 ( \34006 , \34005 );
or \U$34020 ( \34007 , \34004 , \34006 );
buf \U$34021 ( \34008 , RIc0da0a8_91);
buf \U$34022 ( \34009 , RIc0d7fd8_21);
xnor \U$34023 ( \34010 , \34008 , \34009 );
buf \U$34024 ( \34011 , \34010 );
buf \U$34025 ( \34012 , \34011 );
not \U$34026 ( \34013 , \34012 );
buf \U$34027 ( \34014 , \1933 );
nand \U$34028 ( \34015 , \34013 , \34014 );
buf \U$34029 ( \34016 , \34015 );
buf \U$34030 ( \34017 , \34016 );
nand \U$34031 ( \34018 , \34007 , \34017 );
buf \U$34032 ( \34019 , \34018 );
buf \U$34033 ( \34020 , \34019 );
xor \U$34034 ( \34021 , \34002 , \34020 );
buf \U$34035 ( \34022 , \34021 );
buf \U$34036 ( \34023 , \33139 );
not \U$34037 ( \34024 , \34023 );
buf \U$34038 ( \34025 , \1063 );
not \U$34039 ( \34026 , \34025 );
or \U$34040 ( \34027 , \34024 , \34026 );
buf \U$34041 ( \34028 , \1078 );
xor \U$34042 ( \34029 , RIc0d9bf8_81, RIc0d8488_31);
buf \U$34043 ( \34030 , \34029 );
nand \U$34044 ( \34031 , \34028 , \34030 );
buf \U$34045 ( \34032 , \34031 );
buf \U$34046 ( \34033 , \34032 );
nand \U$34047 ( \34034 , \34027 , \34033 );
buf \U$34048 ( \34035 , \34034 );
buf \U$34049 ( \34036 , \34035 );
buf \U$34050 ( \34037 , \33454 );
not \U$34051 ( \34038 , \34037 );
buf \U$34052 ( \34039 , \842 );
not \U$34053 ( \34040 , \34039 );
or \U$34054 ( \34041 , \34038 , \34040 );
xnor \U$34055 ( \34042 , RIc0d9fb8_89, RIc0d80c8_23);
buf \U$34056 ( \34043 , \34042 );
not \U$34057 ( \34044 , \34043 );
buf \U$34058 ( \34045 , \846 );
nand \U$34059 ( \34046 , \34044 , \34045 );
buf \U$34060 ( \34047 , \34046 );
buf \U$34061 ( \34048 , \34047 );
nand \U$34062 ( \34049 , \34041 , \34048 );
buf \U$34063 ( \34050 , \34049 );
buf \U$34064 ( \34051 , \34050 );
xor \U$34065 ( \34052 , \34036 , \34051 );
buf \U$34066 ( \34053 , \33281 );
not \U$34067 ( \34054 , \34053 );
buf \U$34068 ( \34055 , \27591 );
not \U$34069 ( \34056 , \34055 );
or \U$34070 ( \34057 , \34054 , \34056 );
buf \U$34071 ( \34058 , \344 );
buf \U$34072 ( \34059 , RIc0d7df8_17);
buf \U$34073 ( \34060 , RIc0da288_95);
xor \U$34074 ( \34061 , \34059 , \34060 );
buf \U$34075 ( \34062 , \34061 );
buf \U$34076 ( \34063 , \34062 );
nand \U$34077 ( \34064 , \34058 , \34063 );
buf \U$34078 ( \34065 , \34064 );
buf \U$34079 ( \34066 , \34065 );
nand \U$34080 ( \34067 , \34057 , \34066 );
buf \U$34081 ( \34068 , \34067 );
buf \U$34082 ( \34069 , \34068 );
xor \U$34083 ( \34070 , \34052 , \34069 );
buf \U$34084 ( \34071 , \34070 );
xor \U$34085 ( \34072 , \34022 , \34071 );
buf \U$34086 ( \34073 , \33017 );
not \U$34087 ( \34074 , \34073 );
buf \U$34088 ( \34075 , \14075 );
not \U$34089 ( \34076 , \34075 );
or \U$34090 ( \34077 , \34074 , \34076 );
buf \U$34091 ( \34078 , \792 );
buf \U$34092 ( \34079 , RIc0d9838_73);
buf \U$34093 ( \34080 , RIc0d8848_39);
xor \U$34094 ( \34081 , \34079 , \34080 );
buf \U$34095 ( \34082 , \34081 );
buf \U$34096 ( \34083 , \34082 );
nand \U$34097 ( \34084 , \34078 , \34083 );
buf \U$34098 ( \34085 , \34084 );
buf \U$34099 ( \34086 , \34085 );
nand \U$34100 ( \34087 , \34077 , \34086 );
buf \U$34101 ( \34088 , \34087 );
buf \U$34102 ( \34089 , \34088 );
buf \U$34103 ( \34090 , \32830 );
not \U$34104 ( \34091 , \34090 );
buf \U$34105 ( \34092 , \618 );
not \U$34106 ( \34093 , \34092 );
or \U$34107 ( \34094 , \34091 , \34093 );
buf \U$34108 ( \34095 , \14331 );
buf \U$34109 ( \34096 , RIc0d9ec8_87);
buf \U$34110 ( \34097 , RIc0d81b8_25);
xor \U$34111 ( \34098 , \34096 , \34097 );
buf \U$34112 ( \34099 , \34098 );
buf \U$34113 ( \34100 , \34099 );
nand \U$34114 ( \34101 , \34095 , \34100 );
buf \U$34115 ( \34102 , \34101 );
buf \U$34116 ( \34103 , \34102 );
nand \U$34117 ( \34104 , \34094 , \34103 );
buf \U$34118 ( \34105 , \34104 );
buf \U$34119 ( \34106 , \34105 );
xor \U$34120 ( \34107 , \34089 , \34106 );
buf \U$34121 ( \34108 , \33263 );
not \U$34122 ( \34109 , \34108 );
buf \U$34123 ( \34110 , \3535 );
not \U$34124 ( \34111 , \34110 );
or \U$34125 ( \34112 , \34109 , \34111 );
buf \U$34126 ( \34113 , \4049 );
buf \U$34127 ( \34114 , RIc0d7b28_11);
buf \U$34128 ( \34115 , RIc0da558_101);
xor \U$34129 ( \34116 , \34114 , \34115 );
buf \U$34130 ( \34117 , \34116 );
buf \U$34131 ( \34118 , \34117 );
nand \U$34132 ( \34119 , \34113 , \34118 );
buf \U$34133 ( \34120 , \34119 );
buf \U$34134 ( \34121 , \34120 );
nand \U$34135 ( \34122 , \34112 , \34121 );
buf \U$34136 ( \34123 , \34122 );
buf \U$34137 ( \34124 , \34123 );
xor \U$34138 ( \34125 , \34107 , \34124 );
buf \U$34139 ( \34126 , \34125 );
xor \U$34140 ( \34127 , \34072 , \34126 );
not \U$34141 ( \34128 , \34127 );
xor \U$34142 ( \34129 , \33980 , \34128 );
buf \U$34143 ( \34130 , \34129 );
xor \U$34144 ( \34131 , \33875 , \34130 );
buf \U$34145 ( \34132 , \34131 );
buf \U$34146 ( \34133 , \34132 );
xor \U$34147 ( \34134 , \33781 , \34133 );
buf \U$34148 ( \34135 , \34134 );
buf \U$34149 ( \34136 , \34135 );
not \U$34150 ( \34137 , \34136 );
xor \U$34151 ( \34138 , \33533 , \33539 );
and \U$34152 ( \34139 , \34138 , \33555 );
and \U$34153 ( \34140 , \33533 , \33539 );
or \U$34154 ( \34141 , \34139 , \34140 );
buf \U$34155 ( \34142 , \34141 );
buf \U$34156 ( \34143 , \34142 );
buf \U$34157 ( \34144 , \32876 );
not \U$34158 ( \34145 , \34144 );
buf \U$34159 ( \34146 , \32761 );
not \U$34160 ( \34147 , \34146 );
buf \U$34161 ( \34148 , \34147 );
buf \U$34162 ( \34149 , \34148 );
not \U$34163 ( \34150 , \34149 );
or \U$34164 ( \34151 , \34145 , \34150 );
buf \U$34165 ( \34152 , \34148 );
buf \U$34166 ( \34153 , \32876 );
or \U$34167 ( \34154 , \34152 , \34153 );
buf \U$34168 ( \34155 , \32663 );
nand \U$34169 ( \34156 , \34154 , \34155 );
buf \U$34170 ( \34157 , \34156 );
buf \U$34171 ( \34158 , \34157 );
nand \U$34172 ( \34159 , \34151 , \34158 );
buf \U$34173 ( \34160 , \34159 );
buf \U$34174 ( \34161 , \34160 );
xor \U$34175 ( \34162 , \34143 , \34161 );
buf \U$34176 ( \34163 , \33119 );
not \U$34177 ( \34164 , \34163 );
buf \U$34178 ( \34165 , \4692 );
not \U$34179 ( \34166 , \34165 );
or \U$34180 ( \34167 , \34164 , \34166 );
buf \U$34181 ( \34168 , \284 );
buf \U$34182 ( \34169 , RIc0d8a28_43);
buf \U$34183 ( \34170 , RIc0d9658_69);
xor \U$34184 ( \34171 , \34169 , \34170 );
buf \U$34185 ( \34172 , \34171 );
buf \U$34186 ( \34173 , \34172 );
nand \U$34187 ( \34174 , \34168 , \34173 );
buf \U$34188 ( \34175 , \34174 );
buf \U$34189 ( \34176 , \34175 );
nand \U$34190 ( \34177 , \34167 , \34176 );
buf \U$34191 ( \34178 , \34177 );
buf \U$34192 ( \34179 , \34178 );
buf \U$34193 ( \34180 , \32813 );
not \U$34194 ( \34181 , \34180 );
buf \U$34195 ( \34182 , \1736 );
not \U$34196 ( \34183 , \34182 );
or \U$34197 ( \34184 , \34181 , \34183 );
buf \U$34198 ( \34185 , \993 );
buf \U$34199 ( \34186 , RIc0d8398_29);
buf \U$34200 ( \34187 , RIc0d9ce8_83);
xor \U$34201 ( \34188 , \34186 , \34187 );
buf \U$34202 ( \34189 , \34188 );
buf \U$34203 ( \34190 , \34189 );
nand \U$34204 ( \34191 , \34185 , \34190 );
buf \U$34205 ( \34192 , \34191 );
buf \U$34206 ( \34193 , \34192 );
nand \U$34207 ( \34194 , \34184 , \34193 );
buf \U$34208 ( \34195 , \34194 );
buf \U$34209 ( \34196 , \34195 );
xor \U$34210 ( \34197 , \34179 , \34196 );
buf \U$34211 ( \34198 , \33506 );
not \U$34212 ( \34199 , \34198 );
buf \U$34213 ( \34200 , \12331 );
not \U$34214 ( \34201 , \34200 );
buf \U$34215 ( \34202 , \34201 );
buf \U$34216 ( \34203 , \34202 );
not \U$34217 ( \34204 , \34203 );
or \U$34218 ( \34205 , \34199 , \34204 );
buf \U$34219 ( \34206 , \12342 );
buf \U$34220 ( \34207 , RIc0da828_107);
buf \U$34221 ( \34208 , RIc0d7858_5);
xor \U$34222 ( \34209 , \34207 , \34208 );
buf \U$34223 ( \34210 , \34209 );
buf \U$34224 ( \34211 , \34210 );
nand \U$34225 ( \34212 , \34206 , \34211 );
buf \U$34226 ( \34213 , \34212 );
buf \U$34227 ( \34214 , \34213 );
nand \U$34228 ( \34215 , \34205 , \34214 );
buf \U$34229 ( \34216 , \34215 );
buf \U$34230 ( \34217 , \34216 );
xor \U$34231 ( \34218 , \34197 , \34217 );
buf \U$34232 ( \34219 , \34218 );
buf \U$34233 ( \34220 , \34219 );
not \U$34234 ( \34221 , \34220 );
buf \U$34235 ( \34222 , \34221 );
buf \U$34236 ( \34223 , \34222 );
not \U$34237 ( \34224 , \34223 );
buf \U$34238 ( \34225 , \33521 );
not \U$34239 ( \34226 , \34225 );
buf \U$34240 ( \34227 , \16494 );
not \U$34241 ( \34228 , \34227 );
or \U$34242 ( \34229 , \34226 , \34228 );
buf \U$34243 ( \34230 , \1143 );
buf \U$34244 ( \34231 , RIc0d8758_37);
buf \U$34245 ( \34232 , RIc0d9928_75);
xor \U$34246 ( \34233 , \34231 , \34232 );
buf \U$34247 ( \34234 , \34233 );
buf \U$34248 ( \34235 , \34234 );
nand \U$34249 ( \34236 , \34230 , \34235 );
buf \U$34250 ( \34237 , \34236 );
buf \U$34251 ( \34238 , \34237 );
nand \U$34252 ( \34239 , \34229 , \34238 );
buf \U$34253 ( \34240 , \34239 );
buf \U$34254 ( \34241 , \34240 );
buf \U$34255 ( \34242 , \12410 );
not \U$34256 ( \34243 , \34242 );
buf \U$34257 ( \34244 , \34243 );
buf \U$34258 ( \34245 , \34244 );
not \U$34259 ( \34246 , \34245 );
buf \U$34260 ( \34247 , \14888 );
not \U$34261 ( \34248 , \34247 );
or \U$34262 ( \34249 , \34246 , \34248 );
buf \U$34263 ( \34250 , RIc0daaf8_113);
nand \U$34264 ( \34251 , \34249 , \34250 );
buf \U$34265 ( \34252 , \34251 );
buf \U$34266 ( \34253 , \34252 );
xor \U$34267 ( \34254 , \34241 , \34253 );
buf \U$34268 ( \34255 , \33170 );
not \U$34269 ( \34256 , \34255 );
buf \U$34270 ( \34257 , \1183 );
not \U$34271 ( \34258 , \34257 );
or \U$34272 ( \34259 , \34256 , \34258 );
buf \U$34273 ( \34260 , \3742 );
buf \U$34274 ( \34261 , RIc0d8668_35);
buf \U$34275 ( \34262 , RIc0d9a18_77);
xor \U$34276 ( \34263 , \34261 , \34262 );
buf \U$34277 ( \34264 , \34263 );
buf \U$34278 ( \34265 , \34264 );
nand \U$34279 ( \34266 , \34260 , \34265 );
buf \U$34280 ( \34267 , \34266 );
buf \U$34281 ( \34268 , \34267 );
nand \U$34282 ( \34269 , \34259 , \34268 );
buf \U$34283 ( \34270 , \34269 );
buf \U$34284 ( \34271 , \34270 );
xor \U$34285 ( \34272 , \34254 , \34271 );
buf \U$34286 ( \34273 , \34272 );
buf \U$34287 ( \34274 , \34273 );
not \U$34288 ( \34275 , \34274 );
buf \U$34289 ( \34276 , \33438 );
not \U$34290 ( \34277 , \34276 );
buf \U$34291 ( \34278 , \19695 );
not \U$34292 ( \34279 , \34278 );
or \U$34293 ( \34280 , \34277 , \34279 );
buf \U$34294 ( \34281 , \14648 );
xor \U$34295 ( \34282 , RIc0da468_99, RIc0d7c18_13);
buf \U$34296 ( \34283 , \34282 );
nand \U$34297 ( \34284 , \34281 , \34283 );
buf \U$34298 ( \34285 , \34284 );
buf \U$34299 ( \34286 , \34285 );
nand \U$34300 ( \34287 , \34280 , \34286 );
buf \U$34301 ( \34288 , \34287 );
buf \U$34302 ( \34289 , \33316 );
not \U$34303 ( \34290 , \34289 );
buf \U$34304 ( \34291 , \14346 );
not \U$34305 ( \34292 , \34291 );
or \U$34306 ( \34293 , \34290 , \34292 );
buf \U$34307 ( \34294 , \14353 );
xor \U$34308 ( \34295 , RIc0daa08_111, RIc0d7678_1);
buf \U$34309 ( \34296 , \34295 );
nand \U$34310 ( \34297 , \34294 , \34296 );
buf \U$34311 ( \34298 , \34297 );
buf \U$34312 ( \34299 , \34298 );
nand \U$34313 ( \34300 , \34293 , \34299 );
buf \U$34314 ( \34301 , \34300 );
buf \U$34315 ( \34302 , \34301 );
not \U$34316 ( \34303 , \34302 );
buf \U$34317 ( \34304 , \34303 );
xor \U$34318 ( \34305 , \34288 , \34304 );
buf \U$34319 ( \34306 , \33193 );
not \U$34320 ( \34307 , \34306 );
buf \U$34321 ( \34308 , \5305 );
not \U$34322 ( \34309 , \34308 );
or \U$34323 ( \34310 , \34307 , \34309 );
buf \U$34324 ( \34311 , \921 );
buf \U$34325 ( \34312 , RIc0d82a8_27);
buf \U$34326 ( \34313 , RIc0d9dd8_85);
xor \U$34327 ( \34314 , \34312 , \34313 );
buf \U$34328 ( \34315 , \34314 );
buf \U$34329 ( \34316 , \34315 );
nand \U$34330 ( \34317 , \34311 , \34316 );
buf \U$34331 ( \34318 , \34317 );
buf \U$34332 ( \34319 , \34318 );
nand \U$34333 ( \34320 , \34310 , \34319 );
buf \U$34334 ( \34321 , \34320 );
buf \U$34335 ( \34322 , \34321 );
not \U$34336 ( \34323 , \34322 );
buf \U$34337 ( \34324 , \34323 );
xnor \U$34338 ( \34325 , \34305 , \34324 );
buf \U$34339 ( \34326 , \34325 );
not \U$34340 ( \34327 , \34326 );
or \U$34341 ( \34328 , \34275 , \34327 );
buf \U$34342 ( \34329 , \34325 );
buf \U$34343 ( \34330 , \34273 );
or \U$34344 ( \34331 , \34329 , \34330 );
nand \U$34345 ( \34332 , \34328 , \34331 );
buf \U$34346 ( \34333 , \34332 );
buf \U$34347 ( \34334 , \34333 );
not \U$34348 ( \34335 , \34334 );
or \U$34349 ( \34336 , \34224 , \34335 );
buf \U$34350 ( \34337 , \34333 );
buf \U$34351 ( \34338 , \34222 );
or \U$34352 ( \34339 , \34337 , \34338 );
nand \U$34353 ( \34340 , \34336 , \34339 );
buf \U$34354 ( \34341 , \34340 );
buf \U$34355 ( \34342 , \34341 );
buf \U$34356 ( \34343 , \33211 );
not \U$34357 ( \34344 , \34343 );
buf \U$34358 ( \34345 , \476 );
not \U$34359 ( \34346 , \34345 );
or \U$34360 ( \34347 , \34344 , \34346 );
buf \U$34361 ( \34348 , \481 );
xor \U$34362 ( \34349 , RIc0da198_93, RIc0d7ee8_19);
buf \U$34363 ( \34350 , \34349 );
nand \U$34364 ( \34351 , \34348 , \34350 );
buf \U$34365 ( \34352 , \34351 );
buf \U$34366 ( \34353 , \34352 );
nand \U$34367 ( \34354 , \34347 , \34353 );
buf \U$34368 ( \34355 , \34354 );
buf \U$34369 ( \34356 , \34355 );
buf \U$34370 ( \34357 , \33400 );
not \U$34371 ( \34358 , \34357 );
buf \U$34372 ( \34359 , \1021 );
not \U$34373 ( \34360 , \34359 );
or \U$34374 ( \34361 , \34358 , \34360 );
buf \U$34375 ( \34362 , \1026 );
buf \U$34376 ( \34363 , RIc0d8578_33);
buf \U$34377 ( \34364 , RIc0d9b08_79);
xor \U$34378 ( \34365 , \34363 , \34364 );
buf \U$34379 ( \34366 , \34365 );
buf \U$34380 ( \34367 , \34366 );
nand \U$34381 ( \34368 , \34362 , \34367 );
buf \U$34382 ( \34369 , \34368 );
buf \U$34383 ( \34370 , \34369 );
nand \U$34384 ( \34371 , \34361 , \34370 );
buf \U$34385 ( \34372 , \34371 );
buf \U$34386 ( \34373 , \34372 );
xor \U$34387 ( \34374 , \34356 , \34373 );
buf \U$34388 ( \34375 , \32796 );
not \U$34389 ( \34376 , \34375 );
buf \U$34390 ( \34377 , \21959 );
not \U$34391 ( \34378 , \34377 );
or \U$34392 ( \34379 , \34376 , \34378 );
buf \U$34393 ( \34380 , \20211 );
buf \U$34394 ( \34381 , RIc0da918_109);
buf \U$34395 ( \34382 , RIc0d7768_3);
and \U$34396 ( \34383 , \34381 , \34382 );
not \U$34397 ( \34384 , \34381 );
buf \U$34398 ( \34385 , \304 );
and \U$34399 ( \34386 , \34384 , \34385 );
nor \U$34400 ( \34387 , \34383 , \34386 );
buf \U$34401 ( \34388 , \34387 );
buf \U$34402 ( \34389 , \34388 );
nand \U$34403 ( \34390 , \34380 , \34389 );
buf \U$34404 ( \34391 , \34390 );
buf \U$34405 ( \34392 , \34391 );
nand \U$34406 ( \34393 , \34379 , \34392 );
buf \U$34407 ( \34394 , \34393 );
buf \U$34408 ( \34395 , \34394 );
xor \U$34409 ( \34396 , \34374 , \34395 );
buf \U$34410 ( \34397 , \34396 );
buf \U$34411 ( \34398 , \34397 );
not \U$34412 ( \34399 , \34398 );
buf \U$34413 ( \34400 , \33418 );
not \U$34414 ( \34401 , \34400 );
buf \U$34415 ( \34402 , \29546 );
not \U$34416 ( \34403 , \34402 );
or \U$34417 ( \34404 , \34401 , \34403 );
buf \U$34418 ( \34405 , \13048 );
buf \U$34419 ( \34406 , RIc0da648_103);
buf \U$34420 ( \34407 , RIc0d7a38_9);
xor \U$34421 ( \34408 , \34406 , \34407 );
buf \U$34422 ( \34409 , \34408 );
buf \U$34423 ( \34410 , \34409 );
nand \U$34424 ( \34411 , \34405 , \34410 );
buf \U$34425 ( \34412 , \34411 );
buf \U$34426 ( \34413 , \34412 );
nand \U$34427 ( \34414 , \34404 , \34413 );
buf \U$34428 ( \34415 , \34414 );
buf \U$34429 ( \34416 , \34415 );
not \U$34430 ( \34417 , \34416 );
buf \U$34431 ( \34418 , \33490 );
not \U$34432 ( \34419 , \34418 );
buf \U$34433 ( \34420 , \15644 );
not \U$34434 ( \34421 , \34420 );
or \U$34435 ( \34422 , \34419 , \34421 );
buf \U$34436 ( \34423 , \12744 );
buf \U$34437 ( \34424 , RIc0da738_105);
buf \U$34438 ( \34425 , RIc0d7948_7);
xor \U$34439 ( \34426 , \34424 , \34425 );
buf \U$34440 ( \34427 , \34426 );
buf \U$34441 ( \34428 , \34427 );
nand \U$34442 ( \34429 , \34423 , \34428 );
buf \U$34443 ( \34430 , \34429 );
buf \U$34444 ( \34431 , \34430 );
nand \U$34445 ( \34432 , \34422 , \34431 );
buf \U$34446 ( \34433 , \34432 );
buf \U$34447 ( \34434 , \34433 );
not \U$34448 ( \34435 , \34434 );
buf \U$34449 ( \34436 , \34435 );
buf \U$34450 ( \34437 , \34436 );
not \U$34451 ( \34438 , \34437 );
or \U$34452 ( \34439 , \34417 , \34438 );
buf \U$34453 ( \34440 , \34415 );
buf \U$34454 ( \34441 , \34436 );
or \U$34455 ( \34442 , \34440 , \34441 );
nand \U$34456 ( \34443 , \34439 , \34442 );
buf \U$34457 ( \34444 , \34443 );
buf \U$34458 ( \34445 , \34444 );
buf \U$34459 ( \34446 , \32838 );
and \U$34460 ( \34447 , \34445 , \34446 );
not \U$34461 ( \34448 , \34445 );
buf \U$34462 ( \34449 , \32838 );
not \U$34463 ( \34450 , \34449 );
buf \U$34464 ( \34451 , \34450 );
buf \U$34465 ( \34452 , \34451 );
and \U$34466 ( \34453 , \34448 , \34452 );
nor \U$34467 ( \34454 , \34447 , \34453 );
buf \U$34468 ( \34455 , \34454 );
buf \U$34469 ( \34456 , \34455 );
not \U$34470 ( \34457 , \34456 );
or \U$34471 ( \34458 , \34399 , \34457 );
buf \U$34472 ( \34459 , \34455 );
buf \U$34473 ( \34460 , \34397 );
or \U$34474 ( \34461 , \34459 , \34460 );
nand \U$34475 ( \34462 , \34458 , \34461 );
buf \U$34476 ( \34463 , \34462 );
buf \U$34477 ( \34464 , \34463 );
xor \U$34478 ( \34465 , \32824 , \32839 );
and \U$34479 ( \34466 , \34465 , \32855 );
and \U$34480 ( \34467 , \32824 , \32839 );
or \U$34481 ( \34468 , \34466 , \34467 );
buf \U$34482 ( \34469 , \34468 );
buf \U$34483 ( \34470 , \34469 );
xor \U$34484 ( \34471 , \34464 , \34470 );
buf \U$34485 ( \34472 , \34471 );
buf \U$34486 ( \34473 , \34472 );
xor \U$34487 ( \34474 , \34342 , \34473 );
xor \U$34488 ( \34475 , \32821 , \32858 );
and \U$34489 ( \34476 , \34475 , \32874 );
and \U$34490 ( \34477 , \32821 , \32858 );
or \U$34491 ( \34478 , \34476 , \34477 );
buf \U$34492 ( \34479 , \34478 );
buf \U$34493 ( \34480 , \34479 );
xor \U$34494 ( \34481 , \34474 , \34480 );
buf \U$34495 ( \34482 , \34481 );
buf \U$34496 ( \34483 , \34482 );
xor \U$34497 ( \34484 , \34162 , \34483 );
buf \U$34498 ( \34485 , \34484 );
buf \U$34499 ( \34486 , \34485 );
not \U$34500 ( \34487 , \34486 );
xor \U$34501 ( \34488 , \33379 , \33558 );
and \U$34502 ( \34489 , \34488 , \33565 );
and \U$34503 ( \34490 , \33379 , \33558 );
or \U$34504 ( \34491 , \34489 , \34490 );
buf \U$34505 ( \34492 , \34491 );
buf \U$34506 ( \34493 , \34492 );
not \U$34507 ( \34494 , \34493 );
buf \U$34508 ( \34495 , \34494 );
buf \U$34509 ( \34496 , \34495 );
not \U$34510 ( \34497 , \34496 );
or \U$34511 ( \34498 , \34487 , \34497 );
buf \U$34512 ( \34499 , \34485 );
buf \U$34513 ( \34500 , \34495 );
or \U$34514 ( \34501 , \34499 , \34500 );
nand \U$34515 ( \34502 , \34498 , \34501 );
buf \U$34516 ( \34503 , \34502 );
buf \U$34517 ( \34504 , \34503 );
xor \U$34518 ( \34505 , \32887 , \32893 );
and \U$34519 ( \34506 , \34505 , \33354 );
and \U$34520 ( \34507 , \32887 , \32893 );
or \U$34521 ( \34508 , \34506 , \34507 );
buf \U$34522 ( \34509 , \34508 );
buf \U$34523 ( \34510 , \34509 );
not \U$34524 ( \34511 , \34510 );
buf \U$34525 ( \34512 , \34511 );
buf \U$34526 ( \34513 , \34512 );
and \U$34527 ( \34514 , \34504 , \34513 );
not \U$34528 ( \34515 , \34504 );
buf \U$34529 ( \34516 , \34509 );
and \U$34530 ( \34517 , \34515 , \34516 );
nor \U$34531 ( \34518 , \34514 , \34517 );
buf \U$34532 ( \34519 , \34518 );
buf \U$34533 ( \34520 , \34519 );
not \U$34534 ( \34521 , \34520 );
or \U$34535 ( \34522 , \34137 , \34521 );
buf \U$34536 ( \34523 , \34135 );
buf \U$34537 ( \34524 , \34519 );
or \U$34538 ( \34525 , \34523 , \34524 );
nand \U$34539 ( \34526 , \34522 , \34525 );
buf \U$34540 ( \34527 , \34526 );
buf \U$34541 ( \34528 , \34527 );
buf \U$34542 ( \34529 , \33570 );
not \U$34543 ( \34530 , \34529 );
buf \U$34544 ( \34531 , \33590 );
not \U$34545 ( \34532 , \34531 );
or \U$34546 ( \34533 , \34530 , \34532 );
buf \U$34547 ( \34534 , \33371 );
nand \U$34548 ( \34535 , \34533 , \34534 );
buf \U$34549 ( \34536 , \34535 );
buf \U$34550 ( \34537 , \34536 );
buf \U$34551 ( \34538 , \33587 );
buf \U$34552 ( \34539 , \33567 );
nand \U$34553 ( \34540 , \34538 , \34539 );
buf \U$34554 ( \34541 , \34540 );
buf \U$34555 ( \34542 , \34541 );
nand \U$34556 ( \34543 , \34537 , \34542 );
buf \U$34557 ( \34544 , \34543 );
buf \U$34558 ( \34545 , \34544 );
not \U$34559 ( \34546 , \34545 );
buf \U$34560 ( \34547 , \34546 );
buf \U$34561 ( \34548 , \34547 );
and \U$34562 ( \34549 , \34528 , \34548 );
not \U$34563 ( \34550 , \34528 );
buf \U$34564 ( \34551 , \34544 );
and \U$34565 ( \34552 , \34550 , \34551 );
nor \U$34566 ( \34553 , \34549 , \34552 );
buf \U$34567 ( \34554 , \34553 );
buf \U$34568 ( \34555 , \34554 );
buf \U$34569 ( \34556 , \33356 );
not \U$34570 ( \34557 , \34556 );
buf \U$34571 ( \34558 , \34557 );
buf \U$34572 ( \34559 , \34558 );
not \U$34573 ( \34560 , \34559 );
buf \U$34574 ( \34561 , \33597 );
not \U$34575 ( \34562 , \34561 );
or \U$34576 ( \34563 , \34560 , \34562 );
buf \U$34577 ( \34564 , \33616 );
nand \U$34578 ( \34565 , \34563 , \34564 );
buf \U$34579 ( \34566 , \34565 );
buf \U$34580 ( \34567 , \34566 );
buf \U$34581 ( \34568 , \33597 );
not \U$34582 ( \34569 , \34568 );
buf \U$34583 ( \34570 , \33356 );
nand \U$34584 ( \34571 , \34569 , \34570 );
buf \U$34585 ( \34572 , \34571 );
buf \U$34586 ( \34573 , \34572 );
and \U$34587 ( \34574 , \34567 , \34573 );
buf \U$34588 ( \34575 , \34574 );
buf \U$34589 ( \34576 , \34575 );
nand \U$34590 ( \34577 , \34555 , \34576 );
buf \U$34591 ( \34578 , \34577 );
buf \U$34592 ( \34579 , \34578 );
nand \U$34593 ( \34580 , \33621 , \34579 );
buf \U$34594 ( \34581 , \34580 );
buf \U$34595 ( \34582 , \34581 );
not \U$34596 ( \34583 , \34582 );
buf \U$34597 ( \34584 , \31592 );
buf \U$34598 ( \34585 , \31906 );
and \U$34599 ( \34586 , \34584 , \34585 );
not \U$34600 ( \34587 , \34584 );
buf \U$34601 ( \34588 , \31903 );
and \U$34602 ( \34589 , \34587 , \34588 );
nor \U$34603 ( \34590 , \34586 , \34589 );
buf \U$34604 ( \34591 , \34590 );
buf \U$34605 ( \34592 , \34591 );
buf \U$34606 ( \34593 , \31927 );
not \U$34607 ( \34594 , \34593 );
buf \U$34608 ( \34595 , \34594 );
buf \U$34609 ( \34596 , \34595 );
and \U$34610 ( \34597 , \34592 , \34596 );
not \U$34611 ( \34598 , \34592 );
buf \U$34612 ( \34599 , \31927 );
and \U$34613 ( \34600 , \34598 , \34599 );
nor \U$34614 ( \34601 , \34597 , \34600 );
buf \U$34615 ( \34602 , \34601 );
buf \U$34616 ( \34603 , \34602 );
not \U$34617 ( \34604 , \34603 );
buf \U$34618 ( \34605 , \34604 );
buf \U$34619 ( \34606 , \34605 );
not \U$34620 ( \34607 , \34606 );
buf \U$34621 ( \34608 , \32157 );
not \U$34622 ( \34609 , \34608 );
buf \U$34623 ( \34610 , \32031 );
not \U$34624 ( \34611 , \34610 );
and \U$34625 ( \34612 , \34609 , \34611 );
buf \U$34626 ( \34613 , \32157 );
buf \U$34627 ( \34614 , \32031 );
and \U$34628 ( \34615 , \34613 , \34614 );
nor \U$34629 ( \34616 , \34612 , \34615 );
buf \U$34630 ( \34617 , \34616 );
buf \U$34631 ( \34618 , \34617 );
buf \U$34632 ( \34619 , \31944 );
xor \U$34633 ( \34620 , \34618 , \34619 );
buf \U$34634 ( \34621 , \34620 );
buf \U$34635 ( \34622 , \34621 );
not \U$34636 ( \34623 , \34622 );
buf \U$34637 ( \34624 , \34623 );
buf \U$34638 ( \34625 , \34624 );
not \U$34639 ( \34626 , \34625 );
or \U$34640 ( \34627 , \34607 , \34626 );
buf \U$34641 ( \34628 , \34602 );
not \U$34642 ( \34629 , \34628 );
buf \U$34643 ( \34630 , \34621 );
not \U$34644 ( \34631 , \34630 );
or \U$34645 ( \34632 , \34629 , \34631 );
xor \U$34646 ( \34633 , \30846 , \30587 );
and \U$34647 ( \34634 , \34633 , \30802 );
not \U$34648 ( \34635 , \34633 );
and \U$34649 ( \34636 , \34635 , \30805 );
nor \U$34650 ( \34637 , \34634 , \34636 );
buf \U$34651 ( \34638 , \34637 );
xor \U$34652 ( \34639 , \31957 , \31948 );
xor \U$34653 ( \34640 , \34639 , \31952 );
buf \U$34654 ( \34641 , \34640 );
buf \U$34655 ( \34642 , \31994 );
not \U$34656 ( \34643 , \34642 );
buf \U$34657 ( \34644 , \31979 );
not \U$34658 ( \34645 , \34644 );
and \U$34659 ( \34646 , \34643 , \34645 );
buf \U$34660 ( \34647 , \31979 );
buf \U$34661 ( \34648 , \31994 );
and \U$34662 ( \34649 , \34647 , \34648 );
nor \U$34663 ( \34650 , \34646 , \34649 );
buf \U$34664 ( \34651 , \34650 );
and \U$34665 ( \34652 , \34651 , \32003 );
not \U$34666 ( \34653 , \34651 );
and \U$34667 ( \34654 , \34653 , \31971 );
or \U$34668 ( \34655 , \34652 , \34654 );
buf \U$34669 ( \34656 , \34655 );
xor \U$34670 ( \34657 , \34641 , \34656 );
xor \U$34671 ( \34658 , \27109 , \27115 );
and \U$34672 ( \34659 , \34658 , \27122 );
and \U$34673 ( \34660 , \27109 , \27115 );
or \U$34674 ( \34661 , \34659 , \34660 );
buf \U$34675 ( \34662 , \34661 );
buf \U$34676 ( \34663 , \34662 );
not \U$34677 ( \34664 , \34663 );
xor \U$34678 ( \34665 , \32089 , \32090 );
xor \U$34679 ( \34666 , \34665 , \32106 );
buf \U$34680 ( \34667 , \34666 );
buf \U$34681 ( \34668 , \34667 );
not \U$34682 ( \34669 , \34668 );
or \U$34683 ( \34670 , \34664 , \34669 );
buf \U$34684 ( \34671 , \34667 );
buf \U$34685 ( \34672 , \34662 );
or \U$34686 ( \34673 , \34671 , \34672 );
xor \U$34687 ( \34674 , \27131 , \27137 );
and \U$34688 ( \34675 , \34674 , \27144 );
and \U$34689 ( \34676 , \27131 , \27137 );
or \U$34690 ( \34677 , \34675 , \34676 );
buf \U$34691 ( \34678 , \34677 );
buf \U$34692 ( \34679 , \34678 );
nand \U$34693 ( \34680 , \34673 , \34679 );
buf \U$34694 ( \34681 , \34680 );
buf \U$34695 ( \34682 , \34681 );
nand \U$34696 ( \34683 , \34670 , \34682 );
buf \U$34697 ( \34684 , \34683 );
buf \U$34698 ( \34685 , \34684 );
and \U$34699 ( \34686 , \34657 , \34685 );
and \U$34700 ( \34687 , \34641 , \34656 );
or \U$34701 ( \34688 , \34686 , \34687 );
buf \U$34702 ( \34689 , \34688 );
buf \U$34703 ( \34690 , \34689 );
xor \U$34704 ( \34691 , \34638 , \34690 );
buf \U$34705 ( \34692 , \32037 );
buf \U$34706 ( \34693 , \32061 );
xor \U$34707 ( \34694 , \34692 , \34693 );
buf \U$34708 ( \34695 , \32151 );
xor \U$34709 ( \34696 , \34694 , \34695 );
buf \U$34710 ( \34697 , \34696 );
buf \U$34711 ( \34698 , \34697 );
and \U$34712 ( \34699 , \34691 , \34698 );
and \U$34713 ( \34700 , \34638 , \34690 );
or \U$34714 ( \34701 , \34699 , \34700 );
buf \U$34715 ( \34702 , \34701 );
buf \U$34716 ( \34703 , \34702 );
nand \U$34717 ( \34704 , \34632 , \34703 );
buf \U$34718 ( \34705 , \34704 );
buf \U$34719 ( \34706 , \34705 );
nand \U$34720 ( \34707 , \34627 , \34706 );
buf \U$34721 ( \34708 , \34707 );
buf \U$34722 ( \34709 , \34708 );
buf \U$34723 ( \34710 , \32252 );
xor \U$34724 ( \34711 , \34709 , \34710 );
buf \U$34725 ( \34712 , \31939 );
not \U$34726 ( \34713 , \34712 );
buf \U$34727 ( \34714 , \32493 );
not \U$34728 ( \34715 , \34714 );
or \U$34729 ( \34716 , \34713 , \34715 );
buf \U$34730 ( \34717 , \32493 );
buf \U$34731 ( \34718 , \31939 );
or \U$34732 ( \34719 , \34717 , \34718 );
nand \U$34733 ( \34720 , \34716 , \34719 );
buf \U$34734 ( \34721 , \34720 );
buf \U$34735 ( \34722 , \34721 );
xor \U$34736 ( \34723 , \34711 , \34722 );
buf \U$34737 ( \34724 , \34723 );
buf \U$34738 ( \34725 , \34724 );
xor \U$34739 ( \34726 , \27345 , \27387 );
and \U$34740 ( \34727 , \34726 , \27443 );
and \U$34741 ( \34728 , \27345 , \27387 );
or \U$34742 ( \34729 , \34727 , \34728 );
buf \U$34743 ( \34730 , \34729 );
buf \U$34744 ( \34731 , \34730 );
not \U$34745 ( \34732 , \34731 );
xor \U$34746 ( \34733 , \32317 , \32324 );
buf \U$34747 ( \34734 , \34733 );
buf \U$34748 ( \34735 , \32335 );
not \U$34749 ( \34736 , \34735 );
buf \U$34750 ( \34737 , \34736 );
buf \U$34751 ( \34738 , \34737 );
and \U$34752 ( \34739 , \34734 , \34738 );
not \U$34753 ( \34740 , \34734 );
buf \U$34754 ( \34741 , \32335 );
and \U$34755 ( \34742 , \34740 , \34741 );
nor \U$34756 ( \34743 , \34739 , \34742 );
buf \U$34757 ( \34744 , \34743 );
buf \U$34758 ( \34745 , \34744 );
not \U$34759 ( \34746 , \34745 );
buf \U$34760 ( \34747 , \34746 );
buf \U$34761 ( \34748 , \34747 );
not \U$34762 ( \34749 , \34748 );
or \U$34763 ( \34750 , \34732 , \34749 );
buf \U$34764 ( \34751 , \34730 );
not \U$34765 ( \34752 , \34751 );
buf \U$34766 ( \34753 , \34744 );
nand \U$34767 ( \34754 , \34752 , \34753 );
buf \U$34768 ( \34755 , \34754 );
buf \U$34769 ( \34756 , \34755 );
xor \U$34770 ( \34757 , \27692 , \27737 );
and \U$34771 ( \34758 , \34757 , \27796 );
and \U$34772 ( \34759 , \27692 , \27737 );
or \U$34773 ( \34760 , \34758 , \34759 );
buf \U$34774 ( \34761 , \34760 );
buf \U$34775 ( \34762 , \34761 );
nand \U$34776 ( \34763 , \34756 , \34762 );
buf \U$34777 ( \34764 , \34763 );
buf \U$34778 ( \34765 , \34764 );
nand \U$34779 ( \34766 , \34750 , \34765 );
buf \U$34780 ( \34767 , \34766 );
buf \U$34781 ( \34768 , \34767 );
not \U$34782 ( \34769 , \34768 );
buf \U$34783 ( \34770 , \34769 );
buf \U$34784 ( \34771 , \34770 );
not \U$34785 ( \34772 , \34771 );
xor \U$34786 ( \34773 , \32307 , \32342 );
xor \U$34787 ( \34774 , \34773 , \32347 );
buf \U$34788 ( \34775 , \34774 );
buf \U$34789 ( \34776 , \34775 );
not \U$34790 ( \34777 , \34776 );
buf \U$34791 ( \34778 , \34777 );
buf \U$34792 ( \34779 , \34778 );
not \U$34793 ( \34780 , \34779 );
or \U$34794 ( \34781 , \34772 , \34780 );
buf \U$34795 ( \34782 , \27173 );
not \U$34796 ( \34783 , \34782 );
buf \U$34797 ( \34784 , \27153 );
not \U$34798 ( \34785 , \34784 );
or \U$34799 ( \34786 , \34783 , \34785 );
buf \U$34800 ( \34787 , \27173 );
buf \U$34801 ( \34788 , \27153 );
or \U$34802 ( \34789 , \34787 , \34788 );
buf \U$34803 ( \34790 , \27192 );
nand \U$34804 ( \34791 , \34789 , \34790 );
buf \U$34805 ( \34792 , \34791 );
buf \U$34806 ( \34793 , \34792 );
nand \U$34807 ( \34794 , \34786 , \34793 );
buf \U$34808 ( \34795 , \34794 );
buf \U$34809 ( \34796 , \34795 );
buf \U$34810 ( \34797 , \32295 );
not \U$34811 ( \34798 , \34797 );
buf \U$34812 ( \34799 , \34798 );
buf \U$34813 ( \34800 , \34799 );
not \U$34814 ( \34801 , \34800 );
buf \U$34815 ( \34802 , \32274 );
not \U$34816 ( \34803 , \34802 );
buf \U$34817 ( \34804 , \32287 );
not \U$34818 ( \34805 , \34804 );
or \U$34819 ( \34806 , \34803 , \34805 );
buf \U$34820 ( \34807 , \32287 );
buf \U$34821 ( \34808 , \32274 );
or \U$34822 ( \34809 , \34807 , \34808 );
nand \U$34823 ( \34810 , \34806 , \34809 );
buf \U$34824 ( \34811 , \34810 );
buf \U$34825 ( \34812 , \34811 );
not \U$34826 ( \34813 , \34812 );
or \U$34827 ( \34814 , \34801 , \34813 );
buf \U$34828 ( \34815 , \34811 );
buf \U$34829 ( \34816 , \34799 );
or \U$34830 ( \34817 , \34815 , \34816 );
nand \U$34831 ( \34818 , \34814 , \34817 );
buf \U$34832 ( \34819 , \34818 );
buf \U$34833 ( \34820 , \34819 );
xor \U$34834 ( \34821 , \34796 , \34820 );
xor \U$34835 ( \34822 , \32122 , \32128 );
xor \U$34836 ( \34823 , \34822 , \32135 );
buf \U$34837 ( \34824 , \34823 );
buf \U$34838 ( \34825 , \34824 );
and \U$34839 ( \34826 , \34821 , \34825 );
and \U$34840 ( \34827 , \34796 , \34820 );
or \U$34841 ( \34828 , \34826 , \34827 );
buf \U$34842 ( \34829 , \34828 );
buf \U$34843 ( \34830 , \34829 );
nand \U$34844 ( \34831 , \34781 , \34830 );
buf \U$34845 ( \34832 , \34831 );
buf \U$34846 ( \34833 , \34832 );
buf \U$34847 ( \34834 , \34775 );
buf \U$34848 ( \34835 , \34767 );
nand \U$34849 ( \34836 , \34834 , \34835 );
buf \U$34850 ( \34837 , \34836 );
buf \U$34851 ( \34838 , \34837 );
nand \U$34852 ( \34839 , \34833 , \34838 );
buf \U$34853 ( \34840 , \34839 );
buf \U$34854 ( \34841 , \34840 );
xor \U$34855 ( \34842 , \32260 , \32352 );
xor \U$34856 ( \34843 , \34842 , \32357 );
buf \U$34857 ( \34844 , \34843 );
buf \U$34858 ( \34845 , \34844 );
xor \U$34859 ( \34846 , \34841 , \34845 );
buf \U$34860 ( \34847 , \32383 );
not \U$34861 ( \34848 , \34847 );
buf \U$34862 ( \34849 , \32377 );
not \U$34863 ( \34850 , \34849 );
or \U$34864 ( \34851 , \34848 , \34850 );
buf \U$34865 ( \34852 , \32374 );
buf \U$34866 ( \34853 , \32370 );
nand \U$34867 ( \34854 , \34852 , \34853 );
buf \U$34868 ( \34855 , \34854 );
buf \U$34869 ( \34856 , \34855 );
nand \U$34870 ( \34857 , \34851 , \34856 );
buf \U$34871 ( \34858 , \34857 );
buf \U$34872 ( \34859 , \34858 );
buf \U$34873 ( \34860 , \32406 );
not \U$34874 ( \34861 , \34860 );
buf \U$34875 ( \34862 , \34861 );
buf \U$34876 ( \34863 , \34862 );
and \U$34877 ( \34864 , \34859 , \34863 );
not \U$34878 ( \34865 , \34859 );
buf \U$34879 ( \34866 , \32406 );
and \U$34880 ( \34867 , \34865 , \34866 );
nor \U$34881 ( \34868 , \34864 , \34867 );
buf \U$34882 ( \34869 , \34868 );
buf \U$34883 ( \34870 , \34869 );
not \U$34884 ( \34871 , \34870 );
buf \U$34885 ( \34872 , \34871 );
not \U$34886 ( \34873 , \34872 );
xnor \U$34887 ( \34874 , \32110 , \32084 );
buf \U$34888 ( \34875 , \34874 );
buf \U$34891 ( \34876 , \32139 );
buf \U$34892 ( \34877 , \34876 );
not \U$34893 ( \34878 , \34877 );
buf \U$34894 ( \34879 , \34878 );
buf \U$34895 ( \34880 , \34879 );
and \U$34896 ( \34881 , \34875 , \34880 );
not \U$34897 ( \34882 , \34875 );
buf \U$34898 ( \34883 , \34876 );
and \U$34899 ( \34884 , \34882 , \34883 );
nor \U$34900 ( \34885 , \34881 , \34884 );
buf \U$34901 ( \34886 , \34885 );
buf \U$34902 ( \34887 , \34886 );
not \U$34903 ( \34888 , \34887 );
buf \U$34904 ( \34889 , \34888 );
not \U$34905 ( \34890 , \34889 );
or \U$34906 ( \34891 , \34873 , \34890 );
not \U$34907 ( \34892 , \34869 );
not \U$34908 ( \34893 , \34886 );
or \U$34909 ( \34894 , \34892 , \34893 );
xor \U$34910 ( \34895 , \32449 , \32466 );
xor \U$34911 ( \34896 , \34895 , \32474 );
buf \U$34912 ( \34897 , \34896 );
nand \U$34913 ( \34898 , \34894 , \34897 );
nand \U$34914 ( \34899 , \34891 , \34898 );
buf \U$34915 ( \34900 , \34899 );
and \U$34916 ( \34901 , \34846 , \34900 );
and \U$34917 ( \34902 , \34841 , \34845 );
or \U$34918 ( \34903 , \34901 , \34902 );
buf \U$34919 ( \34904 , \34903 );
buf \U$34920 ( \34905 , \34904 );
xor \U$34921 ( \34906 , \32362 , \32366 );
xor \U$34922 ( \34907 , \34906 , \32489 );
buf \U$34923 ( \34908 , \34907 );
buf \U$34924 ( \34909 , \34908 );
xor \U$34925 ( \34910 , \34905 , \34909 );
xor \U$34926 ( \34911 , \32413 , \32479 );
xor \U$34927 ( \34912 , \34911 , \32484 );
buf \U$34928 ( \34913 , \34912 );
buf \U$34929 ( \34914 , \34913 );
not \U$34930 ( \34915 , \34914 );
xor \U$34931 ( \34916 , \27516 , \27570 );
and \U$34932 ( \34917 , \34916 , \27626 );
and \U$34933 ( \34918 , \27516 , \27570 );
or \U$34934 ( \34919 , \34917 , \34918 );
buf \U$34935 ( \34920 , \34919 );
buf \U$34936 ( \34921 , \34920 );
buf \U$34937 ( \34922 , \32442 );
not \U$34938 ( \34923 , \34922 );
buf \U$34939 ( \34924 , \34923 );
buf \U$34940 ( \34925 , \34924 );
not \U$34941 ( \34926 , \34925 );
buf \U$34942 ( \34927 , \32433 );
not \U$34943 ( \34928 , \34927 );
buf \U$34944 ( \34929 , \32427 );
not \U$34945 ( \34930 , \34929 );
or \U$34946 ( \34931 , \34928 , \34930 );
buf \U$34947 ( \34932 , \32427 );
buf \U$34948 ( \34933 , \32433 );
or \U$34949 ( \34934 , \34932 , \34933 );
nand \U$34950 ( \34935 , \34931 , \34934 );
buf \U$34951 ( \34936 , \34935 );
buf \U$34952 ( \34937 , \34936 );
not \U$34953 ( \34938 , \34937 );
or \U$34954 ( \34939 , \34926 , \34938 );
buf \U$34955 ( \34940 , \34936 );
buf \U$34956 ( \34941 , \34924 );
or \U$34957 ( \34942 , \34940 , \34941 );
nand \U$34958 ( \34943 , \34939 , \34942 );
buf \U$34959 ( \34944 , \34943 );
buf \U$34960 ( \34945 , \34944 );
xor \U$34961 ( \34946 , \34921 , \34945 );
xor \U$34962 ( \34947 , \32391 , \32398 );
xor \U$34963 ( \34948 , \34947 , \32402 );
buf \U$34964 ( \34949 , \34948 );
buf \U$34965 ( \34950 , \34949 );
and \U$34966 ( \34951 , \34946 , \34950 );
and \U$34967 ( \34952 , \34921 , \34945 );
or \U$34968 ( \34953 , \34951 , \34952 );
buf \U$34969 ( \34954 , \34953 );
buf \U$34970 ( \34955 , \34954 );
xor \U$34971 ( \34956 , \34641 , \34656 );
xor \U$34972 ( \34957 , \34956 , \34685 );
buf \U$34973 ( \34958 , \34957 );
buf \U$34974 ( \34959 , \34958 );
xor \U$34975 ( \34960 , \34955 , \34959 );
xor \U$34976 ( \34961 , \32453 , \32457 );
xor \U$34977 ( \34962 , \34961 , \32461 );
buf \U$34978 ( \34963 , \34962 );
buf \U$34979 ( \34964 , \34963 );
xor \U$34980 ( \34965 , \27227 , \27282 );
and \U$34981 ( \34966 , \34965 , \27329 );
and \U$34982 ( \34967 , \27227 , \27282 );
or \U$34983 ( \34968 , \34966 , \34967 );
buf \U$34984 ( \34969 , \34968 );
buf \U$34985 ( \34970 , \34969 );
xor \U$34986 ( \34971 , \34964 , \34970 );
xor \U$34987 ( \34972 , \27051 , \27056 );
and \U$34988 ( \34973 , \34972 , \27062 );
and \U$34989 ( \34974 , \27051 , \27056 );
or \U$34990 ( \34975 , \34973 , \34974 );
buf \U$34991 ( \34976 , \34975 );
and \U$34992 ( \34977 , \34971 , \34976 );
and \U$34993 ( \34978 , \34964 , \34970 );
or \U$34994 ( \34979 , \34977 , \34978 );
buf \U$34995 ( \34980 , \34979 );
buf \U$34996 ( \34981 , \34980 );
and \U$34997 ( \34982 , \34960 , \34981 );
and \U$34998 ( \34983 , \34955 , \34959 );
or \U$34999 ( \34984 , \34982 , \34983 );
buf \U$35000 ( \34985 , \34984 );
buf \U$35001 ( \34986 , \34985 );
not \U$35002 ( \34987 , \34986 );
or \U$35003 ( \34988 , \34915 , \34987 );
buf \U$35004 ( \34989 , \34985 );
buf \U$35005 ( \34990 , \34913 );
or \U$35006 ( \34991 , \34989 , \34990 );
xor \U$35007 ( \34992 , \34638 , \34690 );
xor \U$35008 ( \34993 , \34992 , \34698 );
buf \U$35009 ( \34994 , \34993 );
buf \U$35010 ( \34995 , \34994 );
nand \U$35011 ( \34996 , \34991 , \34995 );
buf \U$35012 ( \34997 , \34996 );
buf \U$35013 ( \34998 , \34997 );
nand \U$35014 ( \34999 , \34988 , \34998 );
buf \U$35015 ( \35000 , \34999 );
buf \U$35016 ( \35001 , \35000 );
and \U$35017 ( \35002 , \34910 , \35001 );
and \U$35018 ( \35003 , \34905 , \34909 );
or \U$35019 ( \35004 , \35002 , \35003 );
buf \U$35020 ( \35005 , \35004 );
buf \U$35021 ( \35006 , \35005 );
not \U$35022 ( \35007 , \35006 );
buf \U$35023 ( \35008 , \35007 );
buf \U$35024 ( \35009 , \35008 );
xor \U$35025 ( \35010 , \34725 , \35009 );
buf \U$35026 ( \35011 , \35010 );
buf \U$35027 ( \35012 , \35011 );
xor \U$35028 ( \35013 , \34905 , \34909 );
xor \U$35029 ( \35014 , \35013 , \35001 );
buf \U$35030 ( \35015 , \35014 );
buf \U$35031 ( \35016 , \35015 );
buf \U$35032 ( \35017 , \34621 );
buf \U$35033 ( \35018 , \34602 );
and \U$35034 ( \35019 , \35017 , \35018 );
not \U$35035 ( \35020 , \35017 );
buf \U$35036 ( \35021 , \34605 );
and \U$35037 ( \35022 , \35020 , \35021 );
nor \U$35038 ( \35023 , \35019 , \35022 );
buf \U$35039 ( \35024 , \35023 );
buf \U$35040 ( \35025 , \35024 );
buf \U$35041 ( \35026 , \34702 );
xor \U$35042 ( \35027 , \35025 , \35026 );
buf \U$35043 ( \35028 , \35027 );
buf \U$35044 ( \35029 , \35028 );
or \U$35045 ( \35030 , \35016 , \35029 );
xor \U$35046 ( \35031 , \27092 , \27098 );
and \U$35047 ( \35032 , \35031 , \27105 );
and \U$35048 ( \35033 , \27092 , \27098 );
or \U$35049 ( \35034 , \35032 , \35033 );
buf \U$35050 ( \35035 , \35034 );
buf \U$35051 ( \35036 , \35035 );
xor \U$35052 ( \35037 , \34662 , \34667 );
buf \U$35053 ( \35038 , \35037 );
buf \U$35054 ( \35039 , \34678 );
and \U$35055 ( \35040 , \35038 , \35039 );
not \U$35056 ( \35041 , \35038 );
buf \U$35057 ( \35042 , \34678 );
not \U$35058 ( \35043 , \35042 );
buf \U$35059 ( \35044 , \35043 );
buf \U$35060 ( \35045 , \35044 );
and \U$35061 ( \35046 , \35041 , \35045 );
nor \U$35062 ( \35047 , \35040 , \35046 );
buf \U$35063 ( \35048 , \35047 );
buf \U$35064 ( \35049 , \35048 );
xor \U$35065 ( \35050 , \35036 , \35049 );
xor \U$35066 ( \35051 , \27125 , \27147 );
and \U$35067 ( \35052 , \35051 , \27196 );
and \U$35068 ( \35053 , \27125 , \27147 );
or \U$35069 ( \35054 , \35052 , \35053 );
buf \U$35070 ( \35055 , \35054 );
buf \U$35071 ( \35056 , \35055 );
and \U$35072 ( \35057 , \35050 , \35056 );
and \U$35073 ( \35058 , \35036 , \35049 );
or \U$35074 ( \35059 , \35057 , \35058 );
buf \U$35075 ( \35060 , \35059 );
buf \U$35076 ( \35061 , \35060 );
buf \U$35077 ( \35062 , \34778 );
not \U$35078 ( \35063 , \35062 );
buf \U$35079 ( \35064 , \34829 );
not \U$35080 ( \35065 , \35064 );
or \U$35081 ( \35066 , \35063 , \35065 );
buf \U$35082 ( \35067 , \34778 );
buf \U$35083 ( \35068 , \34829 );
or \U$35084 ( \35069 , \35067 , \35068 );
nand \U$35085 ( \35070 , \35066 , \35069 );
buf \U$35086 ( \35071 , \35070 );
buf \U$35087 ( \35072 , \35071 );
buf \U$35088 ( \35073 , \34767 );
and \U$35089 ( \35074 , \35072 , \35073 );
not \U$35090 ( \35075 , \35072 );
buf \U$35091 ( \35076 , \34770 );
and \U$35092 ( \35077 , \35075 , \35076 );
nor \U$35093 ( \35078 , \35074 , \35077 );
buf \U$35094 ( \35079 , \35078 );
buf \U$35095 ( \35080 , \35079 );
xor \U$35096 ( \35081 , \35061 , \35080 );
buf \U$35097 ( \35082 , \34730 );
buf \U$35098 ( \35083 , \34747 );
xor \U$35099 ( \35084 , \35082 , \35083 );
buf \U$35100 ( \35085 , \34761 );
xor \U$35101 ( \35086 , \35084 , \35085 );
buf \U$35102 ( \35087 , \35086 );
buf \U$35103 ( \35088 , \35087 );
xor \U$35104 ( \35089 , \34796 , \34820 );
xor \U$35105 ( \35090 , \35089 , \34825 );
buf \U$35106 ( \35091 , \35090 );
buf \U$35107 ( \35092 , \35091 );
xor \U$35108 ( \35093 , \35088 , \35092 );
xor \U$35109 ( \35094 , \27332 , \27446 );
and \U$35110 ( \35095 , \35094 , \27629 );
and \U$35111 ( \35096 , \27332 , \27446 );
or \U$35112 ( \35097 , \35095 , \35096 );
buf \U$35113 ( \35098 , \35097 );
buf \U$35114 ( \35099 , \35098 );
and \U$35115 ( \35100 , \35093 , \35099 );
and \U$35116 ( \35101 , \35088 , \35092 );
or \U$35117 ( \35102 , \35100 , \35101 );
buf \U$35118 ( \35103 , \35102 );
buf \U$35119 ( \35104 , \35103 );
and \U$35120 ( \35105 , \35081 , \35104 );
and \U$35121 ( \35106 , \35061 , \35080 );
or \U$35122 ( \35107 , \35105 , \35106 );
buf \U$35123 ( \35108 , \35107 );
buf \U$35124 ( \35109 , \35108 );
xor \U$35125 ( \35110 , \34841 , \34845 );
xor \U$35126 ( \35111 , \35110 , \34900 );
buf \U$35127 ( \35112 , \35111 );
buf \U$35128 ( \35113 , \35112 );
xor \U$35129 ( \35114 , \35109 , \35113 );
buf \U$35130 ( \35115 , \34872 );
not \U$35131 ( \35116 , \35115 );
buf \U$35132 ( \35117 , \34897 );
buf \U$35133 ( \35118 , \34886 );
and \U$35134 ( \35119 , \35117 , \35118 );
not \U$35135 ( \35120 , \35117 );
buf \U$35136 ( \35121 , \34889 );
and \U$35137 ( \35122 , \35120 , \35121 );
nor \U$35138 ( \35123 , \35119 , \35122 );
buf \U$35139 ( \35124 , \35123 );
buf \U$35140 ( \35125 , \35124 );
not \U$35141 ( \35126 , \35125 );
or \U$35142 ( \35127 , \35116 , \35126 );
buf \U$35143 ( \35128 , \34872 );
buf \U$35144 ( \35129 , \35124 );
or \U$35145 ( \35130 , \35128 , \35129 );
nand \U$35146 ( \35131 , \35127 , \35130 );
buf \U$35147 ( \35132 , \35131 );
buf \U$35148 ( \35133 , \35132 );
xor \U$35149 ( \35134 , \34921 , \34945 );
xor \U$35150 ( \35135 , \35134 , \34950 );
buf \U$35151 ( \35136 , \35135 );
buf \U$35152 ( \35137 , \35136 );
xor \U$35153 ( \35138 , \27638 , \27799 );
and \U$35154 ( \35139 , \35138 , \27806 );
and \U$35155 ( \35140 , \27638 , \27799 );
or \U$35156 ( \35141 , \35139 , \35140 );
buf \U$35157 ( \35142 , \35141 );
buf \U$35158 ( \35143 , \35142 );
xor \U$35159 ( \35144 , \35137 , \35143 );
xor \U$35160 ( \35145 , \34964 , \34970 );
xor \U$35161 ( \35146 , \35145 , \34976 );
buf \U$35162 ( \35147 , \35146 );
buf \U$35163 ( \35148 , \35147 );
and \U$35164 ( \35149 , \35144 , \35148 );
and \U$35165 ( \35150 , \35137 , \35143 );
or \U$35166 ( \35151 , \35149 , \35150 );
buf \U$35167 ( \35152 , \35151 );
buf \U$35168 ( \35153 , \35152 );
xor \U$35169 ( \35154 , \35133 , \35153 );
xor \U$35170 ( \35155 , \34955 , \34959 );
xor \U$35171 ( \35156 , \35155 , \34981 );
buf \U$35172 ( \35157 , \35156 );
buf \U$35173 ( \35158 , \35157 );
and \U$35174 ( \35159 , \35154 , \35158 );
and \U$35175 ( \35160 , \35133 , \35153 );
or \U$35176 ( \35161 , \35159 , \35160 );
buf \U$35177 ( \35162 , \35161 );
buf \U$35178 ( \35163 , \35162 );
and \U$35179 ( \35164 , \35114 , \35163 );
and \U$35180 ( \35165 , \35109 , \35113 );
or \U$35181 ( \35166 , \35164 , \35165 );
buf \U$35182 ( \35167 , \35166 );
buf \U$35183 ( \35168 , \35167 );
nand \U$35184 ( \35169 , \35030 , \35168 );
buf \U$35185 ( \35170 , \35169 );
buf \U$35186 ( \35171 , \35170 );
buf \U$35187 ( \35172 , \35015 );
buf \U$35188 ( \35173 , \35028 );
nand \U$35189 ( \35174 , \35172 , \35173 );
buf \U$35190 ( \35175 , \35174 );
buf \U$35191 ( \35176 , \35175 );
and \U$35192 ( \35177 , \35171 , \35176 );
buf \U$35193 ( \35178 , \35177 );
buf \U$35194 ( \35179 , \35178 );
nor \U$35195 ( \35180 , \35012 , \35179 );
buf \U$35196 ( \35181 , \35180 );
buf \U$35197 ( \35182 , \35181 );
buf \U$35198 ( \35183 , \34708 );
not \U$35199 ( \35184 , \35183 );
buf \U$35200 ( \35185 , \35184 );
buf \U$35201 ( \35186 , \35185 );
not \U$35202 ( \35187 , \35186 );
buf \U$35203 ( \35188 , \35005 );
not \U$35204 ( \35189 , \35188 );
buf \U$35205 ( \35190 , \35189 );
buf \U$35206 ( \35191 , \35190 );
not \U$35207 ( \35192 , \35191 );
or \U$35208 ( \35193 , \35187 , \35192 );
buf \U$35209 ( \35194 , \32253 );
buf \U$35210 ( \35195 , \35194 );
not \U$35211 ( \35196 , \35195 );
buf \U$35214 ( \35197 , \34721 );
buf \U$35215 ( \35198 , \35197 );
not \U$35216 ( \35199 , \35198 );
or \U$35217 ( \35200 , \35196 , \35199 );
buf \U$35218 ( \35201 , \35197 );
buf \U$35219 ( \35202 , \35194 );
or \U$35220 ( \35203 , \35201 , \35202 );
nand \U$35221 ( \35204 , \35200 , \35203 );
buf \U$35222 ( \35205 , \35204 );
buf \U$35223 ( \35206 , \35205 );
nand \U$35224 ( \35207 , \35193 , \35206 );
buf \U$35225 ( \35208 , \35207 );
buf \U$35226 ( \35209 , \35208 );
buf \U$35227 ( \35210 , \35005 );
buf \U$35228 ( \35211 , \34708 );
nand \U$35229 ( \35212 , \35210 , \35211 );
buf \U$35230 ( \35213 , \35212 );
buf \U$35231 ( \35214 , \35213 );
nand \U$35232 ( \35215 , \35209 , \35214 );
buf \U$35233 ( \35216 , \35215 );
buf \U$35234 ( \35217 , \35216 );
not \U$35235 ( \35218 , \35217 );
buf \U$35236 ( \35219 , \35218 );
buf \U$35237 ( \35220 , \35219 );
buf \U$35238 ( \35221 , \30344 );
not \U$35239 ( \35222 , \35221 );
buf \U$35240 ( \35223 , \32634 );
not \U$35241 ( \35224 , \35223 );
or \U$35242 ( \35225 , \35222 , \35224 );
buf \U$35243 ( \35226 , \32631 );
buf \U$35244 ( \35227 , \30341 );
nand \U$35245 ( \35228 , \35226 , \35227 );
buf \U$35246 ( \35229 , \35228 );
buf \U$35247 ( \35230 , \35229 );
nand \U$35248 ( \35231 , \35225 , \35230 );
buf \U$35249 ( \35232 , \35231 );
buf \U$35250 ( \35233 , \35232 );
buf \U$35251 ( \35234 , \32508 );
and \U$35252 ( \35235 , \35233 , \35234 );
not \U$35253 ( \35236 , \35233 );
buf \U$35254 ( \35237 , \32505 );
and \U$35255 ( \35238 , \35236 , \35237 );
nor \U$35256 ( \35239 , \35235 , \35238 );
buf \U$35257 ( \35240 , \35239 );
buf \U$35258 ( \35241 , \35240 );
nand \U$35259 ( \35242 , \35220 , \35241 );
buf \U$35260 ( \35243 , \35242 );
buf \U$35261 ( \35244 , \35243 );
nand \U$35262 ( \35245 , \35182 , \35244 );
buf \U$35263 ( \35246 , \35245 );
buf \U$35264 ( \35247 , \35246 );
buf \U$35265 ( \35248 , \35240 );
not \U$35266 ( \35249 , \35248 );
buf \U$35267 ( \35250 , \35216 );
nand \U$35268 ( \35251 , \35249 , \35250 );
buf \U$35269 ( \35252 , \35251 );
buf \U$35270 ( \35253 , \35252 );
nand \U$35271 ( \35254 , \35247 , \35253 );
buf \U$35272 ( \35255 , \35254 );
buf \U$35273 ( \35256 , \35255 );
nand \U$35274 ( \35257 , \34583 , \35256 );
buf \U$35275 ( \35258 , \35257 );
buf \U$35276 ( \35259 , \35258 );
buf \U$35277 ( \35260 , \32645 );
not \U$35278 ( \35261 , \35260 );
buf \U$35279 ( \35262 , \33617 );
nor \U$35280 ( \35263 , \35261 , \35262 );
buf \U$35281 ( \35264 , \35263 );
buf \U$35282 ( \35265 , \35264 );
buf \U$35283 ( \35266 , \34578 );
nand \U$35284 ( \35267 , \35265 , \35266 );
buf \U$35285 ( \35268 , \35267 );
buf \U$35286 ( \35269 , \35268 );
nand \U$35287 ( \35270 , \35259 , \35269 );
buf \U$35288 ( \35271 , \35270 );
buf \U$35289 ( \35272 , \35271 );
buf \U$35291 ( \35273 , \34554 );
buf \U$35292 ( \35274 , \34575 );
nor \U$35293 ( \35275 , \35273 , \35274 );
buf \U$35294 ( \35276 , \35275 );
buf \U$35295 ( \35277 , \35276 );
nor \U$35296 ( \35278 , \35272 , \35277 );
buf \U$35297 ( \35279 , \35278 );
buf \U$35298 ( \35280 , \35279 );
not \U$35299 ( \35281 , \26930 );
buf \U$35300 ( \35282 , \35281 );
buf \U$35301 ( \35283 , \26948 );
nand \U$35302 ( \35284 , \35282 , \35283 );
buf \U$35303 ( \35285 , \35284 );
buf \U$35304 ( \35286 , \35285 );
buf \U$35305 ( \35287 , \25926 );
not \U$35306 ( \35288 , \35287 );
buf \U$35307 ( \35289 , \35288 );
buf \U$35308 ( \35290 , \35289 );
buf \U$35309 ( \35291 , \24914 );
nand \U$35310 ( \35292 , \35290 , \35291 );
buf \U$35311 ( \35293 , \35292 );
buf \U$35312 ( \35294 , \35293 );
buf \U$35313 ( \35295 , \27834 );
buf \U$35314 ( \35296 , \26975 );
nand \U$35315 ( \35297 , \35295 , \35296 );
buf \U$35316 ( \35298 , \35297 );
buf \U$35317 ( \35299 , \35298 );
and \U$35318 ( \35300 , \35286 , \35294 , \35299 );
buf \U$35319 ( \35301 , \35300 );
buf \U$35320 ( \35302 , \35301 );
not \U$35321 ( \35303 , \35302 );
buf \U$35322 ( \35304 , \25929 );
buf \U$35323 ( \35305 , \24862 );
buf \U$35324 ( \35306 , \24888 );
nor \U$35325 ( \35307 , \35305 , \35306 );
buf \U$35326 ( \35308 , \35307 );
buf \U$35327 ( \35309 , \35308 );
nand \U$35328 ( \35310 , \35304 , \35309 );
buf \U$35329 ( \35311 , \35310 );
buf \U$35330 ( \35312 , \35311 );
not \U$35331 ( \35313 , \35312 );
or \U$35332 ( \35314 , \35303 , \35313 );
buf \U$35333 ( \35315 , \26954 );
not \U$35334 ( \35316 , \35315 );
buf \U$35335 ( \35317 , \27840 );
not \U$35336 ( \35318 , \35317 );
or \U$35337 ( \35319 , \35316 , \35318 );
buf \U$35338 ( \35320 , \35298 );
nand \U$35339 ( \35321 , \35319 , \35320 );
buf \U$35340 ( \35322 , \35321 );
buf \U$35341 ( \35323 , \35322 );
nand \U$35342 ( \35324 , \35314 , \35323 );
buf \U$35343 ( \35325 , \35324 );
buf \U$35344 ( \35326 , \35325 );
nand \U$35345 ( \35327 , \27850 , \35280 , \35326 );
buf \U$35346 ( \35328 , \35327 );
buf \U$35347 ( \35329 , \35328 );
not \U$35348 ( \35330 , \35329 );
buf \U$35349 ( \35331 , \35243 );
buf \U$35350 ( \35332 , \35011 );
buf \U$35351 ( \35333 , \35178 );
nand \U$35352 ( \35334 , \35332 , \35333 );
buf \U$35353 ( \35335 , \35334 );
buf \U$35354 ( \35336 , \35335 );
nand \U$35355 ( \35337 , \35331 , \35336 );
buf \U$35356 ( \35338 , \35337 );
buf \U$35357 ( \35339 , \35338 );
buf \U$35358 ( \35340 , \34581 );
nor \U$35359 ( \35341 , \35339 , \35340 );
buf \U$35360 ( \35342 , \35341 );
buf \U$35361 ( \35343 , \35342 );
xor \U$35362 ( \35344 , \27209 , \27819 );
and \U$35363 ( \35345 , \35344 , \27826 );
and \U$35364 ( \35346 , \27209 , \27819 );
or \U$35365 ( \35347 , \35345 , \35346 );
buf \U$35366 ( \35348 , \35347 );
buf \U$35367 ( \35349 , \35348 );
xor \U$35368 ( \35350 , \27008 , \27023 );
and \U$35369 ( \35351 , \35350 , \27067 );
and \U$35370 ( \35352 , \27008 , \27023 );
or \U$35371 ( \35353 , \35351 , \35352 );
buf \U$35372 ( \35354 , \35353 );
buf \U$35373 ( \35355 , \35354 );
xor \U$35374 ( \35356 , \27039 , \27045 );
and \U$35375 ( \35357 , \35356 , \27064 );
and \U$35376 ( \35358 , \27039 , \27045 );
or \U$35377 ( \35359 , \35357 , \35358 );
buf \U$35378 ( \35360 , \35359 );
buf \U$35379 ( \35361 , \35360 );
xor \U$35380 ( \35362 , \35036 , \35049 );
xor \U$35381 ( \35363 , \35362 , \35056 );
buf \U$35382 ( \35364 , \35363 );
buf \U$35383 ( \35365 , \35364 );
xor \U$35384 ( \35366 , \35361 , \35365 );
xor \U$35385 ( \35367 , \27108 , \27199 );
and \U$35386 ( \35368 , \35367 , \27206 );
and \U$35387 ( \35369 , \27108 , \27199 );
or \U$35388 ( \35370 , \35368 , \35369 );
buf \U$35389 ( \35371 , \35370 );
buf \U$35390 ( \35372 , \35371 );
xor \U$35391 ( \35373 , \35366 , \35372 );
buf \U$35392 ( \35374 , \35373 );
buf \U$35393 ( \35375 , \35374 );
xor \U$35394 ( \35376 , \35355 , \35375 );
xor \U$35395 ( \35377 , \27632 , \27809 );
and \U$35396 ( \35378 , \35377 , \27816 );
and \U$35397 ( \35379 , \27632 , \27809 );
or \U$35398 ( \35380 , \35378 , \35379 );
buf \U$35399 ( \35381 , \35380 );
buf \U$35400 ( \35382 , \35381 );
xor \U$35401 ( \35383 , \35088 , \35092 );
xor \U$35402 ( \35384 , \35383 , \35099 );
buf \U$35403 ( \35385 , \35384 );
buf \U$35404 ( \35386 , \35385 );
xor \U$35405 ( \35387 , \35382 , \35386 );
xor \U$35406 ( \35388 , \35137 , \35143 );
xor \U$35407 ( \35389 , \35388 , \35148 );
buf \U$35408 ( \35390 , \35389 );
buf \U$35409 ( \35391 , \35390 );
xor \U$35410 ( \35392 , \35387 , \35391 );
buf \U$35411 ( \35393 , \35392 );
buf \U$35412 ( \35394 , \35393 );
xor \U$35413 ( \35395 , \35376 , \35394 );
buf \U$35414 ( \35396 , \35395 );
buf \U$35415 ( \35397 , \35396 );
xor \U$35416 ( \35398 , \35349 , \35397 );
xor \U$35417 ( \35399 , \27070 , \27076 );
and \U$35418 ( \35400 , \35399 , \27829 );
and \U$35419 ( \35401 , \27070 , \27076 );
or \U$35420 ( \35402 , \35400 , \35401 );
buf \U$35421 ( \35403 , \35402 );
buf \U$35422 ( \35404 , \35403 );
xor \U$35423 ( \35405 , \35398 , \35404 );
buf \U$35424 ( \35406 , \35405 );
buf \U$35425 ( \35407 , \35406 );
xor \U$35426 ( \35408 , \26983 , \27001 );
and \U$35427 ( \35409 , \35408 , \27832 );
and \U$35428 ( \35410 , \26983 , \27001 );
or \U$35429 ( \35411 , \35409 , \35410 );
buf \U$35430 ( \35412 , \35411 );
buf \U$35431 ( \35413 , \35412 );
or \U$35432 ( \35414 , \35407 , \35413 );
buf \U$35433 ( \35415 , \35414 );
buf \U$35434 ( \35416 , \35415 );
xor \U$35435 ( \35417 , \35349 , \35397 );
and \U$35436 ( \35418 , \35417 , \35404 );
and \U$35437 ( \35419 , \35349 , \35397 );
or \U$35438 ( \35420 , \35418 , \35419 );
buf \U$35439 ( \35421 , \35420 );
buf \U$35440 ( \35422 , \35421 );
not \U$35441 ( \35423 , \35422 );
buf \U$35442 ( \35424 , \35423 );
buf \U$35443 ( \35425 , \35424 );
xor \U$35444 ( \35426 , \35133 , \35153 );
xor \U$35445 ( \35427 , \35426 , \35158 );
buf \U$35446 ( \35428 , \35427 );
buf \U$35447 ( \35429 , \35428 );
xor \U$35448 ( \35430 , \35355 , \35375 );
and \U$35449 ( \35431 , \35430 , \35394 );
and \U$35450 ( \35432 , \35355 , \35375 );
or \U$35451 ( \35433 , \35431 , \35432 );
buf \U$35452 ( \35434 , \35433 );
buf \U$35453 ( \35435 , \35434 );
xor \U$35454 ( \35436 , \35429 , \35435 );
xor \U$35455 ( \35437 , \35361 , \35365 );
and \U$35456 ( \35438 , \35437 , \35372 );
and \U$35457 ( \35439 , \35361 , \35365 );
or \U$35458 ( \35440 , \35438 , \35439 );
buf \U$35459 ( \35441 , \35440 );
buf \U$35460 ( \35442 , \35441 );
xor \U$35461 ( \35443 , \35061 , \35080 );
xor \U$35462 ( \35444 , \35443 , \35104 );
buf \U$35463 ( \35445 , \35444 );
buf \U$35464 ( \35446 , \35445 );
xor \U$35465 ( \35447 , \35442 , \35446 );
xor \U$35466 ( \35448 , \35382 , \35386 );
and \U$35467 ( \35449 , \35448 , \35391 );
and \U$35468 ( \35450 , \35382 , \35386 );
or \U$35469 ( \35451 , \35449 , \35450 );
buf \U$35470 ( \35452 , \35451 );
buf \U$35471 ( \35453 , \35452 );
xor \U$35472 ( \35454 , \35447 , \35453 );
buf \U$35473 ( \35455 , \35454 );
buf \U$35474 ( \35456 , \35455 );
xor \U$35475 ( \35457 , \35436 , \35456 );
buf \U$35476 ( \35458 , \35457 );
buf \U$35477 ( \35459 , \35458 );
not \U$35478 ( \35460 , \35459 );
buf \U$35479 ( \35461 , \35460 );
buf \U$35480 ( \35462 , \35461 );
nand \U$35481 ( \35463 , \35425 , \35462 );
buf \U$35482 ( \35464 , \35463 );
buf \U$35483 ( \35465 , \35464 );
and \U$35484 ( \35466 , \35416 , \35465 );
buf \U$35485 ( \35467 , \35466 );
buf \U$35486 ( \35468 , \35467 );
xor \U$35487 ( \35469 , \34985 , \34913 );
xor \U$35488 ( \35470 , \35469 , \34994 );
buf \U$35489 ( \35471 , \35470 );
xor \U$35490 ( \35472 , \35442 , \35446 );
and \U$35491 ( \35473 , \35472 , \35453 );
and \U$35492 ( \35474 , \35442 , \35446 );
or \U$35493 ( \35475 , \35473 , \35474 );
buf \U$35494 ( \35476 , \35475 );
buf \U$35495 ( \35477 , \35476 );
xor \U$35496 ( \35478 , \35471 , \35477 );
xor \U$35497 ( \35479 , \35109 , \35113 );
xor \U$35498 ( \35480 , \35479 , \35163 );
buf \U$35499 ( \35481 , \35480 );
buf \U$35500 ( \35482 , \35481 );
xor \U$35501 ( \35483 , \35478 , \35482 );
buf \U$35502 ( \35484 , \35483 );
buf \U$35503 ( \35485 , \35484 );
not \U$35504 ( \35486 , \35485 );
xor \U$35505 ( \35487 , \35429 , \35435 );
and \U$35506 ( \35488 , \35487 , \35456 );
and \U$35507 ( \35489 , \35429 , \35435 );
or \U$35508 ( \35490 , \35488 , \35489 );
buf \U$35509 ( \35491 , \35490 );
buf \U$35510 ( \35492 , \35491 );
not \U$35511 ( \35493 , \35492 );
buf \U$35512 ( \35494 , \35493 );
buf \U$35513 ( \35495 , \35494 );
nand \U$35514 ( \35496 , \35486 , \35495 );
buf \U$35515 ( \35497 , \35496 );
buf \U$35516 ( \35498 , \35497 );
xor \U$35517 ( \35499 , \35471 , \35477 );
and \U$35518 ( \35500 , \35499 , \35482 );
and \U$35519 ( \35501 , \35471 , \35477 );
or \U$35520 ( \35502 , \35500 , \35501 );
buf \U$35521 ( \35503 , \35502 );
not \U$35522 ( \35504 , \35503 );
buf \U$35523 ( \35505 , \35015 );
buf \U$35524 ( \35506 , \35028 );
xor \U$35525 ( \35507 , \35505 , \35506 );
buf \U$35526 ( \35508 , \35507 );
buf \U$35527 ( \35509 , \35508 );
buf \U$35531 ( \35510 , \35167 );
xnor \U$35532 ( \35511 , \35509 , \35510 );
buf \U$35533 ( \35512 , \35511 );
nand \U$35534 ( \35513 , \35504 , \35512 );
buf \U$35535 ( \35514 , \35513 );
nand \U$35536 ( \35515 , \35343 , \35468 , \35498 , \35514 );
buf \U$35537 ( \35516 , \35515 );
buf \U$35538 ( \35517 , \35516 );
buf \U$35539 ( \35518 , \35279 );
nand \U$35540 ( \35519 , \35517 , \35518 );
buf \U$35541 ( \35520 , \35519 );
buf \U$35542 ( \35521 , \35520 );
not \U$35543 ( \35522 , \35521 );
or \U$35544 ( \35523 , \35330 , \35522 );
buf \U$35545 ( \35524 , \35513 );
not \U$35546 ( \35525 , \35524 );
buf \U$35547 ( \35526 , \35497 );
buf \U$35548 ( \35527 , \35406 );
buf \U$35549 ( \35528 , \35412 );
and \U$35550 ( \35529 , \35527 , \35528 );
buf \U$35551 ( \35530 , \35529 );
buf \U$35552 ( \35531 , \35530 );
buf \U$35553 ( \35532 , \35464 );
nand \U$35554 ( \35533 , \35526 , \35531 , \35532 );
buf \U$35555 ( \35534 , \35533 );
buf \U$35556 ( \35535 , \35534 );
buf \U$35557 ( \35536 , \35458 );
buf \U$35558 ( \35537 , \35421 );
nand \U$35559 ( \35538 , \35536 , \35537 );
buf \U$35560 ( \35539 , \35538 );
buf \U$35561 ( \35540 , \35539 );
not \U$35562 ( \35541 , \35540 );
buf \U$35563 ( \35542 , \35497 );
nand \U$35564 ( \35543 , \35541 , \35542 );
buf \U$35565 ( \35544 , \35543 );
buf \U$35566 ( \35545 , \35544 );
buf \U$35567 ( \35546 , \35484 );
buf \U$35568 ( \35547 , \35491 );
nand \U$35569 ( \35548 , \35546 , \35547 );
buf \U$35570 ( \35549 , \35548 );
buf \U$35571 ( \35550 , \35549 );
nand \U$35572 ( \35551 , \35535 , \35545 , \35550 );
buf \U$35573 ( \35552 , \35551 );
buf \U$35574 ( \35553 , \35552 );
not \U$35575 ( \35554 , \35553 );
or \U$35576 ( \35555 , \35525 , \35554 );
buf \U$35577 ( \35556 , \35512 );
not \U$35578 ( \35557 , \35556 );
buf \U$35579 ( \35558 , \35503 );
nand \U$35580 ( \35559 , \35557 , \35558 );
buf \U$35581 ( \35560 , \35559 );
buf \U$35582 ( \35561 , \35560 );
nand \U$35583 ( \35562 , \35555 , \35561 );
buf \U$35584 ( \35563 , \35562 );
buf \U$35585 ( \35564 , \35563 );
buf \U$35586 ( \35565 , \35342 );
nand \U$35587 ( \35566 , \35564 , \35565 );
buf \U$35588 ( \35567 , \35566 );
buf \U$35589 ( \35568 , \35567 );
nand \U$35590 ( \35569 , \35523 , \35568 );
buf \U$35591 ( \35570 , \35569 );
buf \U$35592 ( \35571 , \35570 );
xor \U$35593 ( \35572 , RIc0d9fb8_89, RIc0d7fd8_21);
buf \U$35594 ( \35573 , \35572 );
not \U$35595 ( \35574 , \35573 );
buf \U$35596 ( \35575 , \436 );
not \U$35597 ( \35576 , \35575 );
or \U$35598 ( \35577 , \35574 , \35576 );
buf \U$35599 ( \35578 , \442 );
buf \U$35600 ( \35579 , RIc0d7f60_20);
buf \U$35601 ( \35580 , RIc0d9fb8_89);
xor \U$35602 ( \35581 , \35579 , \35580 );
buf \U$35603 ( \35582 , \35581 );
buf \U$35604 ( \35583 , \35582 );
nand \U$35605 ( \35584 , \35578 , \35583 );
buf \U$35606 ( \35585 , \35584 );
buf \U$35607 ( \35586 , \35585 );
nand \U$35608 ( \35587 , \35577 , \35586 );
buf \U$35609 ( \35588 , \35587 );
not \U$35610 ( \35589 , \35588 );
buf \U$35611 ( \35590 , RIc0d9478_65);
buf \U$35612 ( \35591 , RIc0d8b18_45);
xor \U$35613 ( \35592 , \35590 , \35591 );
buf \U$35614 ( \35593 , \35592 );
buf \U$35615 ( \35594 , \35593 );
not \U$35616 ( \35595 , \35594 );
buf \U$35617 ( \35596 , \3780 );
not \U$35618 ( \35597 , \35596 );
or \U$35619 ( \35598 , \35595 , \35597 );
buf \U$35620 ( \35599 , \1229 );
buf \U$35621 ( \35600 , RIc0d9478_65);
buf \U$35622 ( \35601 , RIc0d8aa0_44);
xor \U$35623 ( \35602 , \35600 , \35601 );
buf \U$35624 ( \35603 , \35602 );
buf \U$35625 ( \35604 , \35603 );
nand \U$35626 ( \35605 , \35599 , \35604 );
buf \U$35627 ( \35606 , \35605 );
buf \U$35628 ( \35607 , \35606 );
nand \U$35629 ( \35608 , \35598 , \35607 );
buf \U$35630 ( \35609 , \35608 );
not \U$35631 ( \35610 , \35609 );
or \U$35632 ( \35611 , \35589 , \35610 );
buf \U$35633 ( \35612 , \35609 );
not \U$35634 ( \35613 , \35612 );
buf \U$35635 ( \35614 , \35613 );
not \U$35636 ( \35615 , \35614 );
buf \U$35637 ( \35616 , \35588 );
not \U$35638 ( \35617 , \35616 );
buf \U$35639 ( \35618 , \35617 );
not \U$35640 ( \35619 , \35618 );
or \U$35641 ( \35620 , \35615 , \35619 );
buf \U$35642 ( \35621 , RIc0da198_93);
buf \U$35643 ( \35622 , RIc0d7df8_17);
xor \U$35644 ( \35623 , \35621 , \35622 );
buf \U$35645 ( \35624 , \35623 );
buf \U$35646 ( \35625 , \35624 );
not \U$35647 ( \35626 , \35625 );
buf \U$35648 ( \35627 , \13569 );
not \U$35649 ( \35628 , \35627 );
or \U$35650 ( \35629 , \35626 , \35628 );
buf \U$35651 ( \35630 , \4008 );
buf \U$35652 ( \35631 , RIc0da198_93);
buf \U$35653 ( \35632 , RIc0d7d80_16);
xor \U$35654 ( \35633 , \35631 , \35632 );
buf \U$35655 ( \35634 , \35633 );
buf \U$35656 ( \35635 , \35634 );
nand \U$35657 ( \35636 , \35630 , \35635 );
buf \U$35658 ( \35637 , \35636 );
buf \U$35659 ( \35638 , \35637 );
nand \U$35660 ( \35639 , \35629 , \35638 );
buf \U$35661 ( \35640 , \35639 );
nand \U$35662 ( \35641 , \35620 , \35640 );
nand \U$35663 ( \35642 , \35611 , \35641 );
buf \U$35664 ( \35643 , \35642 );
buf \U$35665 ( \35644 , RIc0d9dd8_85);
buf \U$35666 ( \35645 , RIc0d81b8_25);
xor \U$35667 ( \35646 , \35644 , \35645 );
buf \U$35668 ( \35647 , \35646 );
buf \U$35669 ( \35648 , \35647 );
not \U$35670 ( \35649 , \35648 );
buf \U$35671 ( \35650 , \6029 );
not \U$35672 ( \35651 , \35650 );
or \U$35673 ( \35652 , \35649 , \35651 );
buf \U$35674 ( \35653 , \2960 );
buf \U$35675 ( \35654 , RIc0d8140_24);
buf \U$35676 ( \35655 , RIc0d9dd8_85);
xor \U$35677 ( \35656 , \35654 , \35655 );
buf \U$35678 ( \35657 , \35656 );
buf \U$35679 ( \35658 , \35657 );
nand \U$35680 ( \35659 , \35653 , \35658 );
buf \U$35681 ( \35660 , \35659 );
buf \U$35682 ( \35661 , \35660 );
nand \U$35683 ( \35662 , \35652 , \35661 );
buf \U$35684 ( \35663 , \35662 );
not \U$35685 ( \35664 , \35663 );
buf \U$35686 ( \35665 , RIc0d8848_39);
buf \U$35687 ( \35666 , RIc0d9748_71);
xor \U$35688 ( \35667 , \35665 , \35666 );
buf \U$35689 ( \35668 , \35667 );
buf \U$35690 ( \35669 , \35668 );
not \U$35691 ( \35670 , \35669 );
buf \U$35692 ( \35671 , \2923 );
not \U$35693 ( \35672 , \35671 );
or \U$35694 ( \35673 , \35670 , \35672 );
buf \U$35695 ( \35674 , \2927 );
buf \U$35696 ( \35675 , RIc0d87d0_38);
buf \U$35697 ( \35676 , RIc0d9748_71);
xor \U$35698 ( \35677 , \35675 , \35676 );
buf \U$35699 ( \35678 , \35677 );
buf \U$35700 ( \35679 , \35678 );
nand \U$35701 ( \35680 , \35674 , \35679 );
buf \U$35702 ( \35681 , \35680 );
buf \U$35703 ( \35682 , \35681 );
nand \U$35704 ( \35683 , \35673 , \35682 );
buf \U$35705 ( \35684 , \35683 );
buf \U$35706 ( \35685 , \35684 );
not \U$35707 ( \35686 , \35685 );
buf \U$35708 ( \35687 , \35686 );
nand \U$35709 ( \35688 , \35664 , \35687 );
not \U$35710 ( \35689 , \35688 );
buf \U$35711 ( \35690 , RIc0da468_99);
buf \U$35712 ( \35691 , RIc0d7b28_11);
xor \U$35713 ( \35692 , \35690 , \35691 );
buf \U$35714 ( \35693 , \35692 );
buf \U$35715 ( \35694 , \35693 );
not \U$35716 ( \35695 , \35694 );
buf \U$35717 ( \35696 , \14419 );
not \U$35718 ( \35697 , \35696 );
or \U$35719 ( \35698 , \35695 , \35697 );
buf \U$35720 ( \35699 , \22006 );
xor \U$35721 ( \35700 , RIc0da468_99, RIc0d7ab0_10);
buf \U$35722 ( \35701 , \35700 );
nand \U$35723 ( \35702 , \35699 , \35701 );
buf \U$35724 ( \35703 , \35702 );
buf \U$35725 ( \35704 , \35703 );
nand \U$35726 ( \35705 , \35698 , \35704 );
buf \U$35727 ( \35706 , \35705 );
not \U$35728 ( \35707 , \35706 );
or \U$35729 ( \35708 , \35689 , \35707 );
buf \U$35730 ( \35709 , \35663 );
buf \U$35731 ( \35710 , \35684 );
nand \U$35732 ( \35711 , \35709 , \35710 );
buf \U$35733 ( \35712 , \35711 );
nand \U$35734 ( \35713 , \35708 , \35712 );
buf \U$35735 ( \35714 , \35713 );
xor \U$35736 ( \35715 , \35643 , \35714 );
buf \U$35737 ( \35716 , RIc0d8488_31);
buf \U$35738 ( \35717 , RIc0d9b08_79);
xor \U$35739 ( \35718 , \35716 , \35717 );
buf \U$35740 ( \35719 , \35718 );
buf \U$35741 ( \35720 , \35719 );
not \U$35742 ( \35721 , \35720 );
buf \U$35743 ( \35722 , \396 );
not \U$35744 ( \35723 , \35722 );
or \U$35745 ( \35724 , \35721 , \35723 );
buf \U$35746 ( \35725 , \403 );
buf \U$35747 ( \35726 , RIc0d9b08_79);
buf \U$35748 ( \35727 , RIc0d8410_30);
xor \U$35749 ( \35728 , \35726 , \35727 );
buf \U$35750 ( \35729 , \35728 );
buf \U$35751 ( \35730 , \35729 );
nand \U$35752 ( \35731 , \35725 , \35730 );
buf \U$35753 ( \35732 , \35731 );
buf \U$35754 ( \35733 , \35732 );
nand \U$35755 ( \35734 , \35724 , \35733 );
buf \U$35756 ( \35735 , \35734 );
buf \U$35757 ( \35736 , \35735 );
buf \U$35758 ( \35737 , RIc0da828_107);
buf \U$35759 ( \35738 , RIc0d7768_3);
and \U$35760 ( \35739 , \35737 , \35738 );
not \U$35761 ( \35740 , \35737 );
buf \U$35762 ( \35741 , \304 );
and \U$35763 ( \35742 , \35740 , \35741 );
nor \U$35764 ( \35743 , \35739 , \35742 );
buf \U$35765 ( \35744 , \35743 );
buf \U$35766 ( \35745 , \35744 );
not \U$35767 ( \35746 , \35745 );
buf \U$35768 ( \35747 , \21898 );
not \U$35769 ( \35748 , \35747 );
or \U$35770 ( \35749 , \35746 , \35748 );
buf \U$35771 ( \35750 , \16071 );
xor \U$35772 ( \35751 , RIc0da828_107, RIc0d76f0_2);
buf \U$35773 ( \35752 , \35751 );
nand \U$35774 ( \35753 , \35750 , \35752 );
buf \U$35775 ( \35754 , \35753 );
buf \U$35776 ( \35755 , \35754 );
nand \U$35777 ( \35756 , \35749 , \35755 );
buf \U$35778 ( \35757 , \35756 );
buf \U$35779 ( \35758 , \35757 );
xor \U$35780 ( \35759 , \35736 , \35758 );
buf \U$35781 ( \35760 , RIc0da288_95);
buf \U$35782 ( \35761 , RIc0d7c90_14);
xor \U$35783 ( \35762 , \35760 , \35761 );
buf \U$35784 ( \35763 , \35762 );
buf \U$35785 ( \35764 , \35763 );
not \U$35786 ( \35765 , \35764 );
buf \U$35787 ( \35766 , \344 );
not \U$35788 ( \35767 , \35766 );
or \U$35789 ( \35768 , \35765 , \35767 );
buf \U$35790 ( \35769 , \14713 );
buf \U$35791 ( \35770 , RIc0da288_95);
buf \U$35792 ( \35771 , RIc0d7d08_15);
xor \U$35793 ( \35772 , \35770 , \35771 );
buf \U$35794 ( \35773 , \35772 );
buf \U$35795 ( \35774 , \35773 );
not \U$35796 ( \35775 , \35774 );
buf \U$35797 ( \35776 , \35775 );
buf \U$35798 ( \35777 , \35776 );
or \U$35799 ( \35778 , \35769 , \35777 );
nand \U$35800 ( \35779 , \35768 , \35778 );
buf \U$35801 ( \35780 , \35779 );
buf \U$35802 ( \35781 , \35780 );
and \U$35803 ( \35782 , \35759 , \35781 );
and \U$35804 ( \35783 , \35736 , \35758 );
or \U$35805 ( \35784 , \35782 , \35783 );
buf \U$35806 ( \35785 , \35784 );
buf \U$35807 ( \35786 , \35785 );
xor \U$35808 ( \35787 , \35715 , \35786 );
buf \U$35809 ( \35788 , \35787 );
buf \U$35810 ( \35789 , \35788 );
buf \U$35811 ( \35790 , RIc0d85f0_34);
buf \U$35812 ( \35791 , RIc0d9928_75);
xor \U$35813 ( \35792 , \35790 , \35791 );
buf \U$35814 ( \35793 , \35792 );
buf \U$35815 ( \35794 , \35793 );
not \U$35816 ( \35795 , \35794 );
buf \U$35817 ( \35796 , \16494 );
not \U$35818 ( \35797 , \35796 );
or \U$35819 ( \35798 , \35795 , \35797 );
buf \U$35820 ( \35799 , \1143 );
buf \U$35821 ( \35800 , RIc0d8578_33);
buf \U$35822 ( \35801 , RIc0d9928_75);
xor \U$35823 ( \35802 , \35800 , \35801 );
buf \U$35824 ( \35803 , \35802 );
buf \U$35825 ( \35804 , \35803 );
nand \U$35826 ( \35805 , \35799 , \35804 );
buf \U$35827 ( \35806 , \35805 );
buf \U$35828 ( \35807 , \35806 );
nand \U$35829 ( \35808 , \35798 , \35807 );
buf \U$35830 ( \35809 , \35808 );
buf \U$35831 ( \35810 , \35809 );
buf \U$35832 ( \35811 , RIc0d9a18_77);
buf \U$35833 ( \35812 , RIc0d8500_32);
xor \U$35834 ( \35813 , \35811 , \35812 );
buf \U$35835 ( \35814 , \35813 );
buf \U$35836 ( \35815 , \35814 );
not \U$35837 ( \35816 , \35815 );
buf \U$35838 ( \35817 , \1183 );
not \U$35839 ( \35818 , \35817 );
or \U$35840 ( \35819 , \35816 , \35818 );
buf \U$35841 ( \35820 , \6141 );
buf \U$35842 ( \35821 , RIc0d9a18_77);
buf \U$35843 ( \35822 , RIc0d8488_31);
xor \U$35844 ( \35823 , \35821 , \35822 );
buf \U$35845 ( \35824 , \35823 );
buf \U$35846 ( \35825 , \35824 );
nand \U$35847 ( \35826 , \35820 , \35825 );
buf \U$35848 ( \35827 , \35826 );
buf \U$35849 ( \35828 , \35827 );
nand \U$35850 ( \35829 , \35819 , \35828 );
buf \U$35851 ( \35830 , \35829 );
buf \U$35852 ( \35831 , \35830 );
xor \U$35853 ( \35832 , \35810 , \35831 );
buf \U$35854 ( \35833 , RIc0d9ec8_87);
buf \U$35855 ( \35834 , RIc0d8050_22);
xor \U$35856 ( \35835 , \35833 , \35834 );
buf \U$35857 ( \35836 , \35835 );
buf \U$35858 ( \35837 , \35836 );
not \U$35859 ( \35838 , \35837 );
buf \U$35860 ( \35839 , \1765 );
not \U$35861 ( \35840 , \35839 );
or \U$35862 ( \35841 , \35838 , \35840 );
buf \U$35863 ( \35842 , \14331 );
buf \U$35864 ( \35843 , RIc0d9ec8_87);
buf \U$35865 ( \35844 , RIc0d7fd8_21);
xor \U$35866 ( \35845 , \35843 , \35844 );
buf \U$35867 ( \35846 , \35845 );
buf \U$35868 ( \35847 , \35846 );
nand \U$35869 ( \35848 , \35842 , \35847 );
buf \U$35870 ( \35849 , \35848 );
buf \U$35871 ( \35850 , \35849 );
nand \U$35872 ( \35851 , \35841 , \35850 );
buf \U$35873 ( \35852 , \35851 );
buf \U$35874 ( \35853 , \35852 );
xor \U$35875 ( \35854 , \35832 , \35853 );
buf \U$35876 ( \35855 , \35854 );
buf \U$35877 ( \35856 , \35855 );
not \U$35878 ( \35857 , \35856 );
buf \U$35879 ( \35858 , \35857 );
buf \U$35880 ( \35859 , \35858 );
not \U$35881 ( \35860 , \35859 );
buf \U$35882 ( \35861 , \35700 );
not \U$35883 ( \35862 , \35861 );
buf \U$35884 ( \35863 , \14419 );
not \U$35885 ( \35864 , \35863 );
or \U$35886 ( \35865 , \35862 , \35864 );
buf \U$35887 ( \35866 , \22006 );
buf \U$35888 ( \35867 , RIc0d7a38_9);
buf \U$35889 ( \35868 , RIc0da468_99);
xor \U$35890 ( \35869 , \35867 , \35868 );
buf \U$35891 ( \35870 , \35869 );
buf \U$35892 ( \35871 , \35870 );
nand \U$35893 ( \35872 , \35866 , \35871 );
buf \U$35894 ( \35873 , \35872 );
buf \U$35895 ( \35874 , \35873 );
nand \U$35896 ( \35875 , \35865 , \35874 );
buf \U$35897 ( \35876 , \35875 );
buf \U$35898 ( \35877 , \35657 );
not \U$35899 ( \35878 , \35877 );
buf \U$35900 ( \35879 , \3292 );
not \U$35901 ( \35880 , \35879 );
or \U$35902 ( \35881 , \35878 , \35880 );
buf \U$35903 ( \35882 , \2960 );
xor \U$35904 ( \35883 , RIc0d9dd8_85, RIc0d80c8_23);
buf \U$35905 ( \35884 , \35883 );
nand \U$35906 ( \35885 , \35882 , \35884 );
buf \U$35907 ( \35886 , \35885 );
buf \U$35908 ( \35887 , \35886 );
nand \U$35909 ( \35888 , \35881 , \35887 );
buf \U$35910 ( \35889 , \35888 );
xor \U$35911 ( \35890 , \35876 , \35889 );
buf \U$35912 ( \35891 , \35890 );
buf \U$35913 ( \35892 , RIc0d86e0_36);
buf \U$35914 ( \35893 , RIc0d9838_73);
xor \U$35915 ( \35894 , \35892 , \35893 );
buf \U$35916 ( \35895 , \35894 );
buf \U$35917 ( \35896 , \35895 );
not \U$35918 ( \35897 , \35896 );
buf \U$35919 ( \35898 , \2871 );
not \U$35920 ( \35899 , \35898 );
or \U$35921 ( \35900 , \35897 , \35899 );
buf \U$35922 ( \35901 , \1856 );
buf \U$35923 ( \35902 , RIc0d8668_35);
buf \U$35924 ( \35903 , RIc0d9838_73);
xor \U$35925 ( \35904 , \35902 , \35903 );
buf \U$35926 ( \35905 , \35904 );
buf \U$35927 ( \35906 , \35905 );
nand \U$35928 ( \35907 , \35901 , \35906 );
buf \U$35929 ( \35908 , \35907 );
buf \U$35930 ( \35909 , \35908 );
nand \U$35931 ( \35910 , \35900 , \35909 );
buf \U$35932 ( \35911 , \35910 );
buf \U$35933 ( \35912 , \35911 );
not \U$35934 ( \35913 , \35912 );
buf \U$35935 ( \35914 , \35913 );
buf \U$35936 ( \35915 , \35914 );
and \U$35937 ( \35916 , \35891 , \35915 );
not \U$35938 ( \35917 , \35891 );
buf \U$35939 ( \35918 , \35911 );
and \U$35940 ( \35919 , \35917 , \35918 );
nor \U$35941 ( \35920 , \35916 , \35919 );
buf \U$35942 ( \35921 , \35920 );
buf \U$35943 ( \35922 , \35921 );
not \U$35944 ( \35923 , \35922 );
buf \U$35945 ( \35924 , \35923 );
buf \U$35946 ( \35925 , \35924 );
not \U$35947 ( \35926 , \35925 );
or \U$35948 ( \35927 , \35860 , \35926 );
buf \U$35949 ( \35928 , \35855 );
buf \U$35950 ( \35929 , \35921 );
nand \U$35951 ( \35930 , \35928 , \35929 );
buf \U$35952 ( \35931 , \35930 );
buf \U$35953 ( \35932 , \35931 );
nand \U$35954 ( \35933 , \35927 , \35932 );
buf \U$35955 ( \35934 , \35933 );
buf \U$35956 ( \35935 , \35934 );
xor \U$35957 ( \35936 , RIc0d9658_69, RIc0d88c0_40);
buf \U$35958 ( \35937 , \35936 );
not \U$35959 ( \35938 , \35937 );
buf \U$35960 ( \35939 , \4692 );
not \U$35961 ( \35940 , \35939 );
or \U$35962 ( \35941 , \35938 , \35940 );
buf \U$35963 ( \35942 , \284 );
xor \U$35964 ( \35943 , RIc0d9658_69, RIc0d8848_39);
buf \U$35965 ( \35944 , \35943 );
nand \U$35966 ( \35945 , \35942 , \35944 );
buf \U$35967 ( \35946 , \35945 );
buf \U$35968 ( \35947 , \35946 );
nand \U$35969 ( \35948 , \35941 , \35947 );
buf \U$35970 ( \35949 , \35948 );
buf \U$35971 ( \35950 , RIc0d9ce8_83);
buf \U$35972 ( \35951 , RIc0d8230_26);
xor \U$35973 ( \35952 , \35950 , \35951 );
buf \U$35974 ( \35953 , \35952 );
buf \U$35975 ( \35954 , \35953 );
not \U$35976 ( \35955 , \35954 );
buf \U$35977 ( \35956 , \1736 );
not \U$35978 ( \35957 , \35956 );
or \U$35979 ( \35958 , \35955 , \35957 );
buf \U$35980 ( \35959 , \584 );
buf \U$35981 ( \35960 , RIc0d9ce8_83);
buf \U$35982 ( \35961 , RIc0d81b8_25);
xor \U$35983 ( \35962 , \35960 , \35961 );
buf \U$35984 ( \35963 , \35962 );
buf \U$35985 ( \35964 , \35963 );
nand \U$35986 ( \35965 , \35959 , \35964 );
buf \U$35987 ( \35966 , \35965 );
buf \U$35988 ( \35967 , \35966 );
nand \U$35989 ( \35968 , \35958 , \35967 );
buf \U$35990 ( \35969 , \35968 );
buf \U$35991 ( \35970 , \35969 );
not \U$35992 ( \35971 , \35970 );
buf \U$35993 ( \35972 , \35971 );
xor \U$35994 ( \35973 , \35949 , \35972 );
buf \U$35995 ( \35974 , \35751 );
not \U$35996 ( \35975 , \35974 );
buf \U$35997 ( \35976 , \28794 );
not \U$35998 ( \35977 , \35976 );
or \U$35999 ( \35978 , \35975 , \35977 );
buf \U$36000 ( \35979 , \16071 );
xor \U$36001 ( \35980 , RIc0da828_107, RIc0d7678_1);
buf \U$36002 ( \35981 , \35980 );
nand \U$36003 ( \35982 , \35979 , \35981 );
buf \U$36004 ( \35983 , \35982 );
buf \U$36005 ( \35984 , \35983 );
nand \U$36006 ( \35985 , \35978 , \35984 );
buf \U$36007 ( \35986 , \35985 );
xnor \U$36008 ( \35987 , \35973 , \35986 );
buf \U$36009 ( \35988 , \35987 );
xor \U$36010 ( \35989 , \35935 , \35988 );
buf \U$36011 ( \35990 , \35989 );
buf \U$36012 ( \35991 , \35990 );
xor \U$36013 ( \35992 , \35789 , \35991 );
buf \U$36014 ( \35993 , \35582 );
not \U$36015 ( \35994 , \35993 );
buf \U$36016 ( \35995 , \18150 );
not \U$36017 ( \35996 , \35995 );
or \U$36018 ( \35997 , \35994 , \35996 );
buf \U$36019 ( \35998 , \16477 );
buf \U$36020 ( \35999 , RIc0d9fb8_89);
buf \U$36021 ( \36000 , RIc0d7ee8_19);
xor \U$36022 ( \36001 , \35999 , \36000 );
buf \U$36023 ( \36002 , \36001 );
buf \U$36024 ( \36003 , \36002 );
nand \U$36025 ( \36004 , \35998 , \36003 );
buf \U$36026 ( \36005 , \36004 );
buf \U$36027 ( \36006 , \36005 );
nand \U$36028 ( \36007 , \35997 , \36006 );
buf \U$36029 ( \36008 , \36007 );
xor \U$36030 ( \36009 , RIc0da558_101, RIc0d79c0_8);
buf \U$36031 ( \36010 , \36009 );
not \U$36032 ( \36011 , \36010 );
buf \U$36033 ( \36012 , \12833 );
not \U$36034 ( \36013 , \36012 );
or \U$36035 ( \36014 , \36011 , \36013 );
buf \U$36036 ( \36015 , \4049 );
buf \U$36037 ( \36016 , RIc0d7948_7);
buf \U$36038 ( \36017 , RIc0da558_101);
xor \U$36039 ( \36018 , \36016 , \36017 );
buf \U$36040 ( \36019 , \36018 );
buf \U$36041 ( \36020 , \36019 );
nand \U$36042 ( \36021 , \36015 , \36020 );
buf \U$36043 ( \36022 , \36021 );
buf \U$36044 ( \36023 , \36022 );
nand \U$36045 ( \36024 , \36014 , \36023 );
buf \U$36046 ( \36025 , \36024 );
xor \U$36047 ( \36026 , \36008 , \36025 );
xor \U$36048 ( \36027 , RIc0d9bf8_81, RIc0d8320_28);
buf \U$36049 ( \36028 , \36027 );
not \U$36050 ( \36029 , \36028 );
buf \U$36051 ( \36030 , \13075 );
not \U$36052 ( \36031 , \36030 );
or \U$36053 ( \36032 , \36029 , \36031 );
buf \U$36054 ( \36033 , \1078 );
xor \U$36055 ( \36034 , RIc0d9bf8_81, RIc0d82a8_27);
buf \U$36056 ( \36035 , \36034 );
nand \U$36057 ( \36036 , \36033 , \36035 );
buf \U$36058 ( \36037 , \36036 );
buf \U$36059 ( \36038 , \36037 );
nand \U$36060 ( \36039 , \36032 , \36038 );
buf \U$36061 ( \36040 , \36039 );
xor \U$36062 ( \36041 , \36026 , \36040 );
buf \U$36063 ( \36042 , \36041 );
not \U$36064 ( \36043 , \36042 );
buf \U$36065 ( \36044 , \36043 );
buf \U$36066 ( \36045 , \36044 );
not \U$36067 ( \36046 , \36045 );
buf \U$36068 ( \36047 , \35763 );
not \U$36069 ( \36048 , \36047 );
buf \U$36070 ( \36049 , \3714 );
not \U$36071 ( \36050 , \36049 );
or \U$36072 ( \36051 , \36048 , \36050 );
buf \U$36073 ( \36052 , \344 );
xor \U$36074 ( \36053 , RIc0da288_95, RIc0d7c18_13);
buf \U$36075 ( \36054 , \36053 );
nand \U$36076 ( \36055 , \36052 , \36054 );
buf \U$36077 ( \36056 , \36055 );
buf \U$36078 ( \36057 , \36056 );
nand \U$36079 ( \36058 , \36051 , \36057 );
buf \U$36080 ( \36059 , \36058 );
buf \U$36081 ( \36060 , \36059 );
buf \U$36082 ( \36061 , RIc0d78d0_6);
buf \U$36083 ( \36062 , RIc0da648_103);
xor \U$36084 ( \36063 , \36061 , \36062 );
buf \U$36085 ( \36064 , \36063 );
buf \U$36086 ( \36065 , \36064 );
not \U$36087 ( \36066 , \36065 );
buf \U$36088 ( \36067 , \15397 );
not \U$36089 ( \36068 , \36067 );
or \U$36090 ( \36069 , \36066 , \36068 );
buf \U$36091 ( \36070 , \20243 );
buf \U$36092 ( \36071 , RIc0d7858_5);
buf \U$36093 ( \36072 , RIc0da648_103);
xor \U$36094 ( \36073 , \36071 , \36072 );
buf \U$36095 ( \36074 , \36073 );
buf \U$36096 ( \36075 , \36074 );
nand \U$36097 ( \36076 , \36070 , \36075 );
buf \U$36098 ( \36077 , \36076 );
buf \U$36099 ( \36078 , \36077 );
nand \U$36100 ( \36079 , \36069 , \36078 );
buf \U$36101 ( \36080 , \36079 );
buf \U$36102 ( \36081 , \36080 );
and \U$36103 ( \36082 , \36060 , \36081 );
not \U$36104 ( \36083 , \36060 );
buf \U$36105 ( \36084 , \36080 );
not \U$36106 ( \36085 , \36084 );
buf \U$36107 ( \36086 , \36085 );
buf \U$36108 ( \36087 , \36086 );
and \U$36109 ( \36088 , \36083 , \36087 );
nor \U$36110 ( \36089 , \36082 , \36088 );
buf \U$36111 ( \36090 , \36089 );
buf \U$36112 ( \36091 , \36090 );
xor \U$36113 ( \36092 , RIc0da738_105, RIc0d77e0_4);
buf \U$36114 ( \36093 , \36092 );
not \U$36115 ( \36094 , \36093 );
buf \U$36116 ( \36095 , \12736 );
not \U$36117 ( \36096 , \36095 );
or \U$36118 ( \36097 , \36094 , \36096 );
buf \U$36119 ( \36098 , \15653 );
buf \U$36120 ( \36099 , RIc0da738_105);
buf \U$36121 ( \36100 , RIc0d7768_3);
xor \U$36122 ( \36101 , \36099 , \36100 );
buf \U$36123 ( \36102 , \36101 );
buf \U$36124 ( \36103 , \36102 );
nand \U$36125 ( \36104 , \36098 , \36103 );
buf \U$36126 ( \36105 , \36104 );
buf \U$36127 ( \36106 , \36105 );
nand \U$36128 ( \36107 , \36097 , \36106 );
buf \U$36129 ( \36108 , \36107 );
buf \U$36130 ( \36109 , \36108 );
xnor \U$36131 ( \36110 , \36091 , \36109 );
buf \U$36132 ( \36111 , \36110 );
buf \U$36133 ( \36112 , \36111 );
not \U$36134 ( \36113 , \36112 );
buf \U$36135 ( \36114 , \36113 );
buf \U$36136 ( \36115 , \36114 );
not \U$36137 ( \36116 , \36115 );
or \U$36138 ( \36117 , \36046 , \36116 );
buf \U$36139 ( \36118 , \36111 );
buf \U$36140 ( \36119 , \36041 );
nand \U$36141 ( \36120 , \36118 , \36119 );
buf \U$36142 ( \36121 , \36120 );
buf \U$36143 ( \36122 , \36121 );
nand \U$36144 ( \36123 , \36117 , \36122 );
buf \U$36145 ( \36124 , \36123 );
buf \U$36146 ( \36125 , \36124 );
and \U$36147 ( \36126 , \35590 , \35591 );
buf \U$36148 ( \36127 , \36126 );
buf \U$36149 ( \36128 , \36127 );
buf \U$36150 ( \36129 , RIc0d9568_67);
buf \U$36151 ( \36130 , RIc0d89b0_42);
xor \U$36152 ( \36131 , \36129 , \36130 );
buf \U$36153 ( \36132 , \36131 );
buf \U$36154 ( \36133 , \36132 );
not \U$36155 ( \36134 , \36133 );
buf \U$36156 ( \36135 , \2900 );
not \U$36157 ( \36136 , \36135 );
or \U$36158 ( \36137 , \36134 , \36136 );
buf \U$36159 ( \36138 , \686 );
buf \U$36160 ( \36139 , RIc0d8938_41);
buf \U$36161 ( \36140 , RIc0d9568_67);
xor \U$36162 ( \36141 , \36139 , \36140 );
buf \U$36163 ( \36142 , \36141 );
buf \U$36164 ( \36143 , \36142 );
nand \U$36165 ( \36144 , \36138 , \36143 );
buf \U$36166 ( \36145 , \36144 );
buf \U$36167 ( \36146 , \36145 );
nand \U$36168 ( \36147 , \36137 , \36146 );
buf \U$36169 ( \36148 , \36147 );
buf \U$36170 ( \36149 , \36148 );
xor \U$36171 ( \36150 , \36128 , \36149 );
buf \U$36172 ( \36151 , RIc0d7e70_18);
buf \U$36173 ( \36152 , RIc0da0a8_91);
xor \U$36174 ( \36153 , \36151 , \36152 );
buf \U$36175 ( \36154 , \36153 );
buf \U$36176 ( \36155 , \36154 );
not \U$36177 ( \36156 , \36155 );
buf \U$36178 ( \36157 , \2535 );
not \U$36179 ( \36158 , \36157 );
or \U$36180 ( \36159 , \36156 , \36158 );
buf \U$36181 ( \36160 , \1933 );
buf \U$36182 ( \36161 , RIc0da0a8_91);
buf \U$36183 ( \36162 , RIc0d7df8_17);
xor \U$36184 ( \36163 , \36161 , \36162 );
buf \U$36185 ( \36164 , \36163 );
buf \U$36186 ( \36165 , \36164 );
nand \U$36187 ( \36166 , \36160 , \36165 );
buf \U$36188 ( \36167 , \36166 );
buf \U$36189 ( \36168 , \36167 );
nand \U$36190 ( \36169 , \36159 , \36168 );
buf \U$36191 ( \36170 , \36169 );
buf \U$36192 ( \36171 , \36170 );
xor \U$36193 ( \36172 , \36150 , \36171 );
buf \U$36194 ( \36173 , \36172 );
buf \U$36195 ( \36174 , \36173 );
xor \U$36196 ( \36175 , \36125 , \36174 );
buf \U$36197 ( \36176 , \36175 );
buf \U$36198 ( \36177 , \36176 );
and \U$36199 ( \36178 , \35992 , \36177 );
and \U$36200 ( \36179 , \35789 , \35991 );
or \U$36201 ( \36180 , \36178 , \36179 );
buf \U$36202 ( \36181 , \36180 );
buf \U$36203 ( \36182 , \36181 );
not \U$36204 ( \36183 , \36182 );
buf \U$36205 ( \36184 , \36183 );
buf \U$36206 ( \36185 , \36184 );
not \U$36207 ( \36186 , \36185 );
buf \U$36208 ( \36187 , \35634 );
not \U$36209 ( \36188 , \36187 );
buf \U$36210 ( \36189 , \889 );
not \U$36211 ( \36190 , \36189 );
or \U$36212 ( \36191 , \36188 , \36190 );
buf \U$36213 ( \36192 , \481 );
xor \U$36214 ( \36193 , RIc0da198_93, RIc0d7d08_15);
buf \U$36215 ( \36194 , \36193 );
nand \U$36216 ( \36195 , \36192 , \36194 );
buf \U$36217 ( \36196 , \36195 );
buf \U$36218 ( \36197 , \36196 );
nand \U$36219 ( \36198 , \36191 , \36197 );
buf \U$36220 ( \36199 , \36198 );
buf \U$36221 ( \36200 , \36199 );
buf \U$36222 ( \36201 , \20211 );
not \U$36223 ( \36202 , \36201 );
buf \U$36224 ( \36203 , \36202 );
buf \U$36225 ( \36204 , \36203 );
not \U$36226 ( \36205 , \36204 );
buf \U$36227 ( \36206 , \14207 );
not \U$36228 ( \36207 , \36206 );
or \U$36229 ( \36208 , \36205 , \36207 );
buf \U$36230 ( \36209 , RIc0da918_109);
nand \U$36231 ( \36210 , \36208 , \36209 );
buf \U$36232 ( \36211 , \36210 );
buf \U$36233 ( \36212 , \36211 );
or \U$36234 ( \36213 , \36200 , \36212 );
buf \U$36235 ( \36214 , \36213 );
buf \U$36236 ( \36215 , \36214 );
buf \U$36237 ( \36216 , \35729 );
not \U$36238 ( \36217 , \36216 );
buf \U$36239 ( \36218 , \4509 );
not \U$36240 ( \36219 , \36218 );
or \U$36241 ( \36220 , \36217 , \36219 );
buf \U$36242 ( \36221 , \402 );
buf \U$36243 ( \36222 , RIc0d9b08_79);
buf \U$36244 ( \36223 , RIc0d8398_29);
xor \U$36245 ( \36224 , \36222 , \36223 );
buf \U$36246 ( \36225 , \36224 );
buf \U$36247 ( \36226 , \36225 );
nand \U$36248 ( \36227 , \36221 , \36226 );
buf \U$36249 ( \36228 , \36227 );
buf \U$36250 ( \36229 , \36228 );
nand \U$36251 ( \36230 , \36220 , \36229 );
buf \U$36252 ( \36231 , \36230 );
buf \U$36253 ( \36232 , \36231 );
and \U$36254 ( \36233 , \36215 , \36232 );
buf \U$36255 ( \36234 , \36199 );
buf \U$36256 ( \36235 , \36211 );
and \U$36257 ( \36236 , \36234 , \36235 );
buf \U$36258 ( \36237 , \36236 );
buf \U$36259 ( \36238 , \36237 );
nor \U$36260 ( \36239 , \36233 , \36238 );
buf \U$36261 ( \36240 , \36239 );
buf \U$36262 ( \36241 , \36240 );
not \U$36263 ( \36242 , \36241 );
not \U$36264 ( \36243 , \36059 );
nand \U$36265 ( \36244 , \36243 , \36086 );
not \U$36266 ( \36245 , \36244 );
not \U$36267 ( \36246 , \36108 );
or \U$36268 ( \36247 , \36245 , \36246 );
buf \U$36269 ( \36248 , \36059 );
buf \U$36270 ( \36249 , \36080 );
nand \U$36271 ( \36250 , \36248 , \36249 );
buf \U$36272 ( \36251 , \36250 );
nand \U$36273 ( \36252 , \36247 , \36251 );
buf \U$36274 ( \36253 , \36252 );
not \U$36275 ( \36254 , \36253 );
or \U$36276 ( \36255 , \36242 , \36254 );
buf \U$36277 ( \36256 , \36252 );
buf \U$36278 ( \36257 , \36240 );
or \U$36279 ( \36258 , \36256 , \36257 );
nand \U$36280 ( \36259 , \36255 , \36258 );
buf \U$36281 ( \36260 , \36259 );
buf \U$36282 ( \36261 , \36260 );
not \U$36283 ( \36262 , \36261 );
xor \U$36284 ( \36263 , \36008 , \36025 );
and \U$36285 ( \36264 , \36263 , \36040 );
and \U$36286 ( \36265 , \36008 , \36025 );
or \U$36287 ( \36266 , \36264 , \36265 );
buf \U$36288 ( \36267 , \36266 );
not \U$36289 ( \36268 , \36267 );
buf \U$36290 ( \36269 , \36268 );
buf \U$36291 ( \36270 , \36269 );
not \U$36292 ( \36271 , \36270 );
and \U$36293 ( \36272 , \36262 , \36271 );
buf \U$36294 ( \36273 , \36260 );
buf \U$36295 ( \36274 , \36269 );
and \U$36296 ( \36275 , \36273 , \36274 );
nor \U$36297 ( \36276 , \36272 , \36275 );
buf \U$36298 ( \36277 , \36276 );
buf \U$36299 ( \36278 , \36277 );
not \U$36300 ( \36279 , \36278 );
buf \U$36301 ( \36280 , \35883 );
not \U$36302 ( \36281 , \36280 );
buf \U$36303 ( \36282 , \1388 );
not \U$36304 ( \36283 , \36282 );
or \U$36305 ( \36284 , \36281 , \36283 );
buf \U$36306 ( \36285 , \17010 );
xor \U$36307 ( \36286 , RIc0d9dd8_85, RIc0d8050_22);
buf \U$36308 ( \36287 , \36286 );
nand \U$36309 ( \36288 , \36285 , \36287 );
buf \U$36310 ( \36289 , \36288 );
buf \U$36311 ( \36290 , \36289 );
nand \U$36312 ( \36291 , \36284 , \36290 );
buf \U$36313 ( \36292 , \36291 );
buf \U$36314 ( \36293 , \36292 );
buf \U$36315 ( \36294 , \35803 );
not \U$36316 ( \36295 , \36294 );
buf \U$36317 ( \36296 , \13383 );
not \U$36318 ( \36297 , \36296 );
or \U$36319 ( \36298 , \36295 , \36297 );
buf \U$36320 ( \36299 , \1143 );
xor \U$36321 ( \36300 , RIc0d9928_75, RIc0d8500_32);
buf \U$36322 ( \36301 , \36300 );
nand \U$36323 ( \36302 , \36299 , \36301 );
buf \U$36324 ( \36303 , \36302 );
buf \U$36325 ( \36304 , \36303 );
nand \U$36326 ( \36305 , \36298 , \36304 );
buf \U$36327 ( \36306 , \36305 );
buf \U$36328 ( \36307 , \36306 );
xor \U$36329 ( \36308 , \36293 , \36307 );
buf \U$36330 ( \36309 , \36102 );
not \U$36331 ( \36310 , \36309 );
buf \U$36332 ( \36311 , \12736 );
not \U$36333 ( \36312 , \36311 );
or \U$36334 ( \36313 , \36310 , \36312 );
buf \U$36335 ( \36314 , \12744 );
buf \U$36336 ( \36315 , RIc0da738_105);
buf \U$36337 ( \36316 , RIc0d76f0_2);
xor \U$36338 ( \36317 , \36315 , \36316 );
buf \U$36339 ( \36318 , \36317 );
buf \U$36340 ( \36319 , \36318 );
nand \U$36341 ( \36320 , \36314 , \36319 );
buf \U$36342 ( \36321 , \36320 );
buf \U$36343 ( \36322 , \36321 );
nand \U$36344 ( \36323 , \36313 , \36322 );
buf \U$36345 ( \36324 , \36323 );
buf \U$36346 ( \36325 , \36324 );
xor \U$36347 ( \36326 , \36308 , \36325 );
buf \U$36348 ( \36327 , \36326 );
buf \U$36349 ( \36328 , \36327 );
buf \U$36350 ( \36329 , RIc0d8758_37);
buf \U$36351 ( \36330 , RIc0d9748_71);
xor \U$36352 ( \36331 , \36329 , \36330 );
buf \U$36353 ( \36332 , \36331 );
buf \U$36354 ( \36333 , \36332 );
not \U$36355 ( \36334 , \36333 );
buf \U$36356 ( \36335 , \12676 );
not \U$36357 ( \36336 , \36335 );
or \U$36358 ( \36337 , \36334 , \36336 );
buf \U$36359 ( \36338 , \12683 );
buf \U$36360 ( \36339 , RIc0d86e0_36);
buf \U$36361 ( \36340 , RIc0d9748_71);
xor \U$36362 ( \36341 , \36339 , \36340 );
buf \U$36363 ( \36342 , \36341 );
buf \U$36364 ( \36343 , \36342 );
nand \U$36365 ( \36344 , \36338 , \36343 );
buf \U$36366 ( \36345 , \36344 );
buf \U$36367 ( \36346 , \36345 );
nand \U$36368 ( \36347 , \36337 , \36346 );
buf \U$36369 ( \36348 , \36347 );
buf \U$36370 ( \36349 , \36348 );
buf \U$36371 ( \36350 , \35963 );
not \U$36372 ( \36351 , \36350 );
buf \U$36373 ( \36352 , \2088 );
not \U$36374 ( \36353 , \36352 );
or \U$36375 ( \36354 , \36351 , \36353 );
buf \U$36376 ( \36355 , \993 );
xor \U$36377 ( \36356 , RIc0d9ce8_83, RIc0d8140_24);
buf \U$36378 ( \36357 , \36356 );
nand \U$36379 ( \36358 , \36355 , \36357 );
buf \U$36380 ( \36359 , \36358 );
buf \U$36381 ( \36360 , \36359 );
nand \U$36382 ( \36361 , \36354 , \36360 );
buf \U$36383 ( \36362 , \36361 );
buf \U$36384 ( \36363 , \36362 );
xor \U$36385 ( \36364 , \36349 , \36363 );
buf \U$36386 ( \36365 , RIc0da378_97);
buf \U$36387 ( \36366 , RIc0d7b28_11);
xor \U$36388 ( \36367 , \36365 , \36366 );
buf \U$36389 ( \36368 , \36367 );
buf \U$36390 ( \36369 , \36368 );
not \U$36391 ( \36370 , \36369 );
buf \U$36392 ( \36371 , \2066 );
not \U$36393 ( \36372 , \36371 );
or \U$36394 ( \36373 , \36370 , \36372 );
buf \U$36395 ( \36374 , \2070 );
buf \U$36396 ( \36375 , RIc0d7ab0_10);
buf \U$36397 ( \36376 , RIc0da378_97);
xor \U$36398 ( \36377 , \36375 , \36376 );
buf \U$36399 ( \36378 , \36377 );
buf \U$36400 ( \36379 , \36378 );
nand \U$36401 ( \36380 , \36374 , \36379 );
buf \U$36402 ( \36381 , \36380 );
buf \U$36403 ( \36382 , \36381 );
nand \U$36404 ( \36383 , \36373 , \36382 );
buf \U$36405 ( \36384 , \36383 );
buf \U$36406 ( \36385 , \36384 );
xor \U$36407 ( \36386 , \36364 , \36385 );
buf \U$36408 ( \36387 , \36386 );
buf \U$36409 ( \36388 , \36387 );
xor \U$36410 ( \36389 , \36328 , \36388 );
buf \U$36411 ( \36390 , \36019 );
not \U$36412 ( \36391 , \36390 );
buf \U$36413 ( \36392 , \4042 );
not \U$36414 ( \36393 , \36392 );
or \U$36415 ( \36394 , \36391 , \36393 );
buf \U$36416 ( \36395 , \12839 );
xor \U$36417 ( \36396 , RIc0da558_101, RIc0d78d0_6);
buf \U$36418 ( \36397 , \36396 );
nand \U$36419 ( \36398 , \36395 , \36397 );
buf \U$36420 ( \36399 , \36398 );
buf \U$36421 ( \36400 , \36399 );
nand \U$36422 ( \36401 , \36394 , \36400 );
buf \U$36423 ( \36402 , \36401 );
buf \U$36424 ( \36403 , \36402 );
buf \U$36425 ( \36404 , \36053 );
not \U$36426 ( \36405 , \36404 );
buf \U$36427 ( \36406 , \330 );
not \U$36428 ( \36407 , \36406 );
or \U$36429 ( \36408 , \36405 , \36407 );
buf \U$36430 ( \36409 , \14707 );
xor \U$36431 ( \36410 , RIc0da288_95, RIc0d7ba0_12);
buf \U$36432 ( \36411 , \36410 );
nand \U$36433 ( \36412 , \36409 , \36411 );
buf \U$36434 ( \36413 , \36412 );
buf \U$36435 ( \36414 , \36413 );
nand \U$36436 ( \36415 , \36408 , \36414 );
buf \U$36437 ( \36416 , \36415 );
buf \U$36438 ( \36417 , \36416 );
xor \U$36439 ( \36418 , \36403 , \36417 );
buf \U$36440 ( \36419 , \36074 );
not \U$36441 ( \36420 , \36419 );
buf \U$36442 ( \36421 , \16578 );
not \U$36443 ( \36422 , \36421 );
or \U$36444 ( \36423 , \36420 , \36422 );
buf \U$36445 ( \36424 , \18416 );
buf \U$36446 ( \36425 , RIc0da648_103);
buf \U$36447 ( \36426 , RIc0d77e0_4);
and \U$36448 ( \36427 , \36425 , \36426 );
not \U$36449 ( \36428 , \36425 );
buf \U$36450 ( \36429 , \489 );
and \U$36451 ( \36430 , \36428 , \36429 );
nor \U$36452 ( \36431 , \36427 , \36430 );
buf \U$36453 ( \36432 , \36431 );
buf \U$36454 ( \36433 , \36432 );
nand \U$36455 ( \36434 , \36424 , \36433 );
buf \U$36456 ( \36435 , \36434 );
buf \U$36457 ( \36436 , \36435 );
nand \U$36458 ( \36437 , \36423 , \36436 );
buf \U$36459 ( \36438 , \36437 );
buf \U$36460 ( \36439 , \36438 );
xor \U$36461 ( \36440 , \36418 , \36439 );
buf \U$36462 ( \36441 , \36440 );
buf \U$36463 ( \36442 , \36441 );
xor \U$36464 ( \36443 , \36389 , \36442 );
buf \U$36465 ( \36444 , \36443 );
buf \U$36466 ( \36445 , \36444 );
not \U$36467 ( \36446 , \36445 );
or \U$36468 ( \36447 , \36279 , \36446 );
buf \U$36469 ( \36448 , \36444 );
buf \U$36470 ( \36449 , \36277 );
or \U$36471 ( \36450 , \36448 , \36449 );
nand \U$36472 ( \36451 , \36447 , \36450 );
buf \U$36473 ( \36452 , \36451 );
buf \U$36474 ( \36453 , \36452 );
buf \U$36475 ( \36454 , \35949 );
not \U$36476 ( \36455 , \36454 );
buf \U$36477 ( \36456 , \36455 );
buf \U$36478 ( \36457 , \36456 );
not \U$36479 ( \36458 , \36457 );
buf \U$36480 ( \36459 , \35972 );
not \U$36481 ( \36460 , \36459 );
or \U$36482 ( \36461 , \36458 , \36460 );
buf \U$36483 ( \36462 , \35986 );
nand \U$36484 ( \36463 , \36461 , \36462 );
buf \U$36485 ( \36464 , \36463 );
buf \U$36486 ( \36465 , \36464 );
buf \U$36487 ( \36466 , \35969 );
buf \U$36488 ( \36467 , \35949 );
nand \U$36489 ( \36468 , \36466 , \36467 );
buf \U$36490 ( \36469 , \36468 );
buf \U$36491 ( \36470 , \36469 );
nand \U$36492 ( \36471 , \36465 , \36470 );
buf \U$36493 ( \36472 , \36471 );
buf \U$36494 ( \36473 , \36472 );
buf \U$36495 ( \36474 , \36164 );
not \U$36496 ( \36475 , \36474 );
buf \U$36497 ( \36476 , \1927 );
not \U$36498 ( \36477 , \36476 );
or \U$36499 ( \36478 , \36475 , \36477 );
buf \U$36500 ( \36479 , \533 );
xor \U$36501 ( \36480 , RIc0da0a8_91, RIc0d7d80_16);
buf \U$36502 ( \36481 , \36480 );
nand \U$36503 ( \36482 , \36479 , \36481 );
buf \U$36504 ( \36483 , \36482 );
buf \U$36505 ( \36484 , \36483 );
nand \U$36506 ( \36485 , \36478 , \36484 );
buf \U$36507 ( \36486 , \36485 );
buf \U$36508 ( \36487 , RIc0d9478_65);
buf \U$36509 ( \36488 , RIc0d8a28_43);
xor \U$36510 ( \36489 , \36487 , \36488 );
buf \U$36511 ( \36490 , \36489 );
buf \U$36512 ( \36491 , \36490 );
not \U$36513 ( \36492 , \36491 );
buf \U$36514 ( \36493 , \1224 );
not \U$36515 ( \36494 , \36493 );
or \U$36516 ( \36495 , \36492 , \36494 );
buf \U$36517 ( \36496 , \1229 );
buf \U$36518 ( \36497 , RIc0d9478_65);
buf \U$36519 ( \36498 , RIc0d89b0_42);
xor \U$36520 ( \36499 , \36497 , \36498 );
buf \U$36521 ( \36500 , \36499 );
buf \U$36522 ( \36501 , \36500 );
nand \U$36523 ( \36502 , \36496 , \36501 );
buf \U$36524 ( \36503 , \36502 );
buf \U$36525 ( \36504 , \36503 );
nand \U$36526 ( \36505 , \36495 , \36504 );
buf \U$36527 ( \36506 , \36505 );
buf \U$36528 ( \36507 , \36506 );
not \U$36529 ( \36508 , \36507 );
buf \U$36530 ( \36509 , \36508 );
xor \U$36531 ( \36510 , \36486 , \36509 );
buf \U$36532 ( \36511 , \36142 );
not \U$36533 ( \36512 , \36511 );
buf \U$36534 ( \36513 , \4904 );
nor \U$36535 ( \36514 , \36512 , \36513 );
buf \U$36536 ( \36515 , \36514 );
buf \U$36537 ( \36516 , \36515 );
buf \U$36538 ( \36517 , \686 );
buf \U$36539 ( \36518 , RIc0d88c0_40);
buf \U$36540 ( \36519 , RIc0d9568_67);
xor \U$36541 ( \36520 , \36518 , \36519 );
buf \U$36542 ( \36521 , \36520 );
buf \U$36543 ( \36522 , \36521 );
and \U$36544 ( \36523 , \36517 , \36522 );
buf \U$36545 ( \36524 , \36523 );
buf \U$36546 ( \36525 , \36524 );
nor \U$36547 ( \36526 , \36516 , \36525 );
buf \U$36548 ( \36527 , \36526 );
xor \U$36549 ( \36528 , \36510 , \36527 );
buf \U$36550 ( \36529 , \36528 );
xor \U$36551 ( \36530 , \36473 , \36529 );
buf \U$36552 ( \36531 , \36193 );
not \U$36553 ( \36532 , \36531 );
buf \U$36554 ( \36533 , \13569 );
not \U$36555 ( \36534 , \36533 );
or \U$36556 ( \36535 , \36532 , \36534 );
buf \U$36557 ( \36536 , \4008 );
xor \U$36558 ( \36537 , RIc0da198_93, RIc0d7c90_14);
buf \U$36559 ( \36538 , \36537 );
nand \U$36560 ( \36539 , \36536 , \36538 );
buf \U$36561 ( \36540 , \36539 );
buf \U$36562 ( \36541 , \36540 );
nand \U$36563 ( \36542 , \36535 , \36541 );
buf \U$36564 ( \36543 , \36542 );
buf \U$36565 ( \36544 , \36002 );
not \U$36566 ( \36545 , \36544 );
buf \U$36567 ( \36546 , \18150 );
not \U$36568 ( \36547 , \36546 );
or \U$36569 ( \36548 , \36545 , \36547 );
buf \U$36570 ( \36549 , \846 );
xor \U$36571 ( \36550 , RIc0d9fb8_89, RIc0d7e70_18);
buf \U$36572 ( \36551 , \36550 );
nand \U$36573 ( \36552 , \36549 , \36551 );
buf \U$36574 ( \36553 , \36552 );
buf \U$36575 ( \36554 , \36553 );
nand \U$36576 ( \36555 , \36548 , \36554 );
buf \U$36577 ( \36556 , \36555 );
xor \U$36578 ( \36557 , \36543 , \36556 );
buf \U$36579 ( \36558 , \36225 );
not \U$36580 ( \36559 , \36558 );
buf \U$36581 ( \36560 , \4509 );
not \U$36582 ( \36561 , \36560 );
or \U$36583 ( \36562 , \36559 , \36561 );
buf \U$36584 ( \36563 , \3985 );
buf \U$36585 ( \36564 , RIc0d9b08_79);
buf \U$36586 ( \36565 , RIc0d8320_28);
xor \U$36587 ( \36566 , \36564 , \36565 );
buf \U$36588 ( \36567 , \36566 );
buf \U$36589 ( \36568 , \36567 );
nand \U$36590 ( \36569 , \36563 , \36568 );
buf \U$36591 ( \36570 , \36569 );
buf \U$36592 ( \36571 , \36570 );
nand \U$36593 ( \36572 , \36562 , \36571 );
buf \U$36594 ( \36573 , \36572 );
xor \U$36595 ( \36574 , \36557 , \36573 );
buf \U$36596 ( \36575 , \36574 );
xor \U$36597 ( \36576 , \36530 , \36575 );
buf \U$36598 ( \36577 , \36576 );
buf \U$36599 ( \36578 , \36577 );
not \U$36600 ( \36579 , \36578 );
buf \U$36601 ( \36580 , \36579 );
buf \U$36602 ( \36581 , \36580 );
and \U$36603 ( \36582 , \36453 , \36581 );
not \U$36604 ( \36583 , \36453 );
buf \U$36605 ( \36584 , \36577 );
and \U$36606 ( \36585 , \36583 , \36584 );
nor \U$36607 ( \36586 , \36582 , \36585 );
buf \U$36608 ( \36587 , \36586 );
buf \U$36609 ( \36588 , \36587 );
not \U$36610 ( \36589 , \36588 );
buf \U$36611 ( \36590 , \36589 );
buf \U$36612 ( \36591 , \36590 );
not \U$36613 ( \36592 , \36591 );
or \U$36614 ( \36593 , \36186 , \36592 );
buf \U$36615 ( \36594 , \36587 );
buf \U$36616 ( \36595 , \36181 );
nand \U$36617 ( \36596 , \36594 , \36595 );
buf \U$36618 ( \36597 , \36596 );
buf \U$36619 ( \36598 , \36597 );
nand \U$36620 ( \36599 , \36593 , \36598 );
buf \U$36621 ( \36600 , \36599 );
buf \U$36622 ( \36601 , RIc0d9478_65);
buf \U$36623 ( \36602 , RIc0d8b90_46);
and \U$36624 ( \36603 , \36601 , \36602 );
buf \U$36625 ( \36604 , \36603 );
buf \U$36626 ( \36605 , \36604 );
buf \U$36627 ( \36606 , RIc0d7948_7);
buf \U$36628 ( \36607 , RIc0da648_103);
xor \U$36629 ( \36608 , \36606 , \36607 );
buf \U$36630 ( \36609 , \36608 );
buf \U$36631 ( \36610 , \36609 );
not \U$36632 ( \36611 , \36610 );
buf \U$36633 ( \36612 , \13042 );
not \U$36634 ( \36613 , \36612 );
or \U$36635 ( \36614 , \36611 , \36613 );
buf \U$36636 ( \36615 , \13048 );
buf \U$36637 ( \36616 , \36064 );
nand \U$36638 ( \36617 , \36615 , \36616 );
buf \U$36639 ( \36618 , \36617 );
buf \U$36640 ( \36619 , \36618 );
nand \U$36641 ( \36620 , \36614 , \36619 );
buf \U$36642 ( \36621 , \36620 );
buf \U$36643 ( \36622 , \36621 );
xor \U$36644 ( \36623 , \36605 , \36622 );
buf \U$36645 ( \36624 , \22631 );
not \U$36646 ( \36625 , \36624 );
buf \U$36647 ( \36626 , \36625 );
buf \U$36648 ( \36627 , \36626 );
not \U$36649 ( \36628 , \36627 );
buf \U$36650 ( \36629 , RIc0d7a38_9);
buf \U$36651 ( \36630 , RIc0da558_101);
xnor \U$36652 ( \36631 , \36629 , \36630 );
buf \U$36653 ( \36632 , \36631 );
buf \U$36654 ( \36633 , \36632 );
not \U$36655 ( \36634 , \36633 );
and \U$36656 ( \36635 , \36628 , \36634 );
not \U$36657 ( \36636 , \36009 );
buf \U$36658 ( \36637 , \26354 );
not \U$36659 ( \36638 , \36637 );
buf \U$36660 ( \36639 , \36638 );
nor \U$36661 ( \36640 , \36636 , \36639 );
buf \U$36662 ( \36641 , \36640 );
nor \U$36663 ( \36642 , \36635 , \36641 );
buf \U$36664 ( \36643 , \36642 );
buf \U$36665 ( \36644 , \36643 );
and \U$36666 ( \36645 , \36623 , \36644 );
and \U$36667 ( \36646 , \36605 , \36622 );
or \U$36668 ( \36647 , \36645 , \36646 );
buf \U$36669 ( \36648 , \36647 );
buf \U$36670 ( \36649 , \36648 );
buf \U$36671 ( \36650 , \36237 );
not \U$36672 ( \36651 , \36650 );
buf \U$36673 ( \36652 , \36214 );
nand \U$36674 ( \36653 , \36651 , \36652 );
buf \U$36675 ( \36654 , \36653 );
buf \U$36676 ( \36655 , \36654 );
buf \U$36677 ( \36656 , \36231 );
xnor \U$36678 ( \36657 , \36655 , \36656 );
buf \U$36679 ( \36658 , \36657 );
buf \U$36680 ( \36659 , \36658 );
xor \U$36681 ( \36660 , \36649 , \36659 );
buf \U$36682 ( \36661 , RIc0d8500_32);
buf \U$36683 ( \36662 , RIc0d9b08_79);
xor \U$36684 ( \36663 , \36661 , \36662 );
buf \U$36685 ( \36664 , \36663 );
buf \U$36686 ( \36665 , \36664 );
not \U$36687 ( \36666 , \36665 );
buf \U$36688 ( \36667 , \14940 );
not \U$36689 ( \36668 , \36667 );
or \U$36690 ( \36669 , \36666 , \36668 );
buf \U$36691 ( \36670 , \1025 );
buf \U$36692 ( \36671 , \35719 );
nand \U$36693 ( \36672 , \36670 , \36671 );
buf \U$36694 ( \36673 , \36672 );
buf \U$36695 ( \36674 , \36673 );
nand \U$36696 ( \36675 , \36669 , \36674 );
buf \U$36697 ( \36676 , \36675 );
buf \U$36698 ( \36677 , \36676 );
xor \U$36699 ( \36678 , RIc0da198_93, RIc0d7e70_18);
buf \U$36700 ( \36679 , \36678 );
not \U$36701 ( \36680 , \36679 );
buf \U$36702 ( \36681 , \889 );
not \U$36703 ( \36682 , \36681 );
or \U$36704 ( \36683 , \36680 , \36682 );
buf \U$36705 ( \36684 , \4008 );
buf \U$36706 ( \36685 , \35624 );
nand \U$36707 ( \36686 , \36684 , \36685 );
buf \U$36708 ( \36687 , \36686 );
buf \U$36709 ( \36688 , \36687 );
nand \U$36710 ( \36689 , \36683 , \36688 );
buf \U$36711 ( \36690 , \36689 );
buf \U$36712 ( \36691 , \36690 );
xor \U$36713 ( \36692 , \36677 , \36691 );
buf \U$36714 ( \36693 , RIc0d76f0_2);
buf \U$36715 ( \36694 , RIc0da918_109);
xor \U$36716 ( \36695 , \36693 , \36694 );
buf \U$36717 ( \36696 , \36695 );
buf \U$36718 ( \36697 , \36696 );
not \U$36719 ( \36698 , \36697 );
buf \U$36720 ( \36699 , \14210 );
not \U$36721 ( \36700 , \36699 );
or \U$36722 ( \36701 , \36698 , \36700 );
buf \U$36723 ( \36702 , \20211 );
buf \U$36724 ( \36703 , RIc0d7678_1);
buf \U$36725 ( \36704 , RIc0da918_109);
xor \U$36726 ( \36705 , \36703 , \36704 );
buf \U$36727 ( \36706 , \36705 );
buf \U$36728 ( \36707 , \36706 );
nand \U$36729 ( \36708 , \36702 , \36707 );
buf \U$36730 ( \36709 , \36708 );
buf \U$36731 ( \36710 , \36709 );
nand \U$36732 ( \36711 , \36701 , \36710 );
buf \U$36733 ( \36712 , \36711 );
buf \U$36734 ( \36713 , \36712 );
and \U$36735 ( \36714 , \36692 , \36713 );
and \U$36736 ( \36715 , \36677 , \36691 );
or \U$36737 ( \36716 , \36714 , \36715 );
buf \U$36738 ( \36717 , \36716 );
buf \U$36739 ( \36718 , \36717 );
not \U$36740 ( \36719 , \36718 );
buf \U$36741 ( \36720 , RIc0d8410_30);
buf \U$36742 ( \36721 , RIc0d9bf8_81);
xor \U$36743 ( \36722 , \36720 , \36721 );
buf \U$36744 ( \36723 , \36722 );
buf \U$36745 ( \36724 , \36723 );
not \U$36746 ( \36725 , \36724 );
buf \U$36747 ( \36726 , \13075 );
not \U$36748 ( \36727 , \36726 );
or \U$36749 ( \36728 , \36725 , \36727 );
buf \U$36750 ( \36729 , \1078 );
xor \U$36751 ( \36730 , RIc0d9bf8_81, RIc0d8398_29);
buf \U$36752 ( \36731 , \36730 );
nand \U$36753 ( \36732 , \36729 , \36731 );
buf \U$36754 ( \36733 , \36732 );
buf \U$36755 ( \36734 , \36733 );
nand \U$36756 ( \36735 , \36728 , \36734 );
buf \U$36757 ( \36736 , \36735 );
buf \U$36758 ( \36737 , \36736 );
not \U$36759 ( \36738 , \36737 );
xor \U$36760 ( \36739 , RIc0da288_95, RIc0d7d80_16);
buf \U$36761 ( \36740 , \36739 );
not \U$36762 ( \36741 , \36740 );
buf \U$36763 ( \36742 , \330 );
not \U$36764 ( \36743 , \36742 );
or \U$36765 ( \36744 , \36741 , \36743 );
buf \U$36766 ( \36745 , \344 );
buf \U$36767 ( \36746 , \35773 );
nand \U$36768 ( \36747 , \36745 , \36746 );
buf \U$36769 ( \36748 , \36747 );
buf \U$36770 ( \36749 , \36748 );
nand \U$36771 ( \36750 , \36744 , \36749 );
buf \U$36772 ( \36751 , \36750 );
buf \U$36773 ( \36752 , \36751 );
not \U$36774 ( \36753 , \36752 );
or \U$36775 ( \36754 , \36738 , \36753 );
buf \U$36776 ( \36755 , \36751 );
buf \U$36777 ( \36756 , \36736 );
or \U$36778 ( \36757 , \36755 , \36756 );
xor \U$36779 ( \36758 , RIc0da648_103, RIc0d79c0_8);
buf \U$36780 ( \36759 , \36758 );
not \U$36781 ( \36760 , \36759 );
buf \U$36782 ( \36761 , \16578 );
not \U$36783 ( \36762 , \36761 );
or \U$36784 ( \36763 , \36760 , \36762 );
buf \U$36785 ( \36764 , \16584 );
buf \U$36786 ( \36765 , \36609 );
nand \U$36787 ( \36766 , \36764 , \36765 );
buf \U$36788 ( \36767 , \36766 );
buf \U$36789 ( \36768 , \36767 );
nand \U$36790 ( \36769 , \36763 , \36768 );
buf \U$36791 ( \36770 , \36769 );
buf \U$36792 ( \36771 , \36770 );
nand \U$36793 ( \36772 , \36757 , \36771 );
buf \U$36794 ( \36773 , \36772 );
buf \U$36795 ( \36774 , \36773 );
nand \U$36796 ( \36775 , \36754 , \36774 );
buf \U$36797 ( \36776 , \36775 );
buf \U$36798 ( \36777 , \36776 );
not \U$36799 ( \36778 , \36777 );
or \U$36800 ( \36779 , \36719 , \36778 );
buf \U$36801 ( \36780 , \36717 );
not \U$36802 ( \36781 , \36780 );
buf \U$36803 ( \36782 , \36781 );
buf \U$36804 ( \36783 , \36782 );
not \U$36805 ( \36784 , \36783 );
buf \U$36806 ( \36785 , \36776 );
not \U$36807 ( \36786 , \36785 );
buf \U$36808 ( \36787 , \36786 );
buf \U$36809 ( \36788 , \36787 );
not \U$36810 ( \36789 , \36788 );
or \U$36811 ( \36790 , \36784 , \36789 );
buf \U$36812 ( \36791 , \615 );
buf \U$36813 ( \36792 , RIc0d8140_24);
buf \U$36814 ( \36793 , RIc0d9ec8_87);
xnor \U$36815 ( \36794 , \36792 , \36793 );
buf \U$36816 ( \36795 , \36794 );
buf \U$36817 ( \36796 , \36795 );
or \U$36818 ( \36797 , \36791 , \36796 );
buf \U$36819 ( \36798 , \819 );
buf \U$36820 ( \36799 , RIc0d80c8_23);
buf \U$36821 ( \36800 , RIc0d9ec8_87);
xnor \U$36822 ( \36801 , \36799 , \36800 );
buf \U$36823 ( \36802 , \36801 );
buf \U$36824 ( \36803 , \36802 );
or \U$36825 ( \36804 , \36798 , \36803 );
nand \U$36826 ( \36805 , \36797 , \36804 );
buf \U$36827 ( \36806 , \36805 );
buf \U$36828 ( \36807 , \36806 );
xor \U$36829 ( \36808 , RIc0da558_101, RIc0d7ab0_10);
buf \U$36830 ( \36809 , \36808 );
not \U$36831 ( \36810 , \36809 );
buf \U$36832 ( \36811 , \33258 );
not \U$36833 ( \36812 , \36811 );
or \U$36834 ( \36813 , \36810 , \36812 );
buf \U$36835 ( \36814 , \36632 );
not \U$36836 ( \36815 , \36814 );
buf \U$36837 ( \36816 , \16676 );
nand \U$36838 ( \36817 , \36815 , \36816 );
buf \U$36839 ( \36818 , \36817 );
buf \U$36840 ( \36819 , \36818 );
nand \U$36841 ( \36820 , \36813 , \36819 );
buf \U$36842 ( \36821 , \36820 );
buf \U$36843 ( \36822 , \36821 );
xor \U$36844 ( \36823 , \36807 , \36822 );
buf \U$36845 ( \36824 , RIc0d9fb8_89);
buf \U$36846 ( \36825 , RIc0d8050_22);
xnor \U$36847 ( \36826 , \36824 , \36825 );
buf \U$36848 ( \36827 , \36826 );
buf \U$36849 ( \36828 , \36827 );
not \U$36850 ( \36829 , \36828 );
buf \U$36851 ( \36830 , \36829 );
buf \U$36852 ( \36831 , \36830 );
not \U$36853 ( \36832 , \36831 );
buf \U$36854 ( \36833 , \3384 );
not \U$36855 ( \36834 , \36833 );
or \U$36856 ( \36835 , \36832 , \36834 );
buf \U$36857 ( \36836 , \846 );
buf \U$36858 ( \36837 , \35572 );
nand \U$36859 ( \36838 , \36836 , \36837 );
buf \U$36860 ( \36839 , \36838 );
buf \U$36861 ( \36840 , \36839 );
nand \U$36862 ( \36841 , \36835 , \36840 );
buf \U$36863 ( \36842 , \36841 );
buf \U$36864 ( \36843 , \36842 );
and \U$36865 ( \36844 , \36823 , \36843 );
and \U$36866 ( \36845 , \36807 , \36822 );
or \U$36867 ( \36846 , \36844 , \36845 );
buf \U$36868 ( \36847 , \36846 );
buf \U$36869 ( \36848 , \36847 );
nand \U$36870 ( \36849 , \36790 , \36848 );
buf \U$36871 ( \36850 , \36849 );
buf \U$36872 ( \36851 , \36850 );
nand \U$36873 ( \36852 , \36779 , \36851 );
buf \U$36874 ( \36853 , \36852 );
buf \U$36875 ( \36854 , \36853 );
and \U$36876 ( \36855 , \36660 , \36854 );
and \U$36877 ( \36856 , \36649 , \36659 );
or \U$36878 ( \36857 , \36855 , \36856 );
buf \U$36879 ( \36858 , \36857 );
buf \U$36880 ( \36859 , \36858 );
buf \U$36881 ( \36860 , \35943 );
not \U$36882 ( \36861 , \36860 );
buf \U$36883 ( \36862 , \864 );
not \U$36884 ( \36863 , \36862 );
or \U$36885 ( \36864 , \36861 , \36863 );
buf \U$36886 ( \36865 , \874 );
buf \U$36887 ( \36866 , RIc0d9658_69);
buf \U$36888 ( \36867 , RIc0d87d0_38);
xor \U$36889 ( \36868 , \36866 , \36867 );
buf \U$36890 ( \36869 , \36868 );
buf \U$36891 ( \36870 , \36869 );
nand \U$36892 ( \36871 , \36865 , \36870 );
buf \U$36893 ( \36872 , \36871 );
buf \U$36894 ( \36873 , \36872 );
nand \U$36895 ( \36874 , \36864 , \36873 );
buf \U$36896 ( \36875 , \36874 );
buf \U$36897 ( \36876 , \36034 );
not \U$36898 ( \36877 , \36876 );
buf \U$36899 ( \36878 , \1063 );
not \U$36900 ( \36879 , \36878 );
or \U$36901 ( \36880 , \36877 , \36879 );
buf \U$36902 ( \36881 , \1078 );
buf \U$36903 ( \36882 , RIc0d9bf8_81);
buf \U$36904 ( \36883 , RIc0d8230_26);
xor \U$36905 ( \36884 , \36882 , \36883 );
buf \U$36906 ( \36885 , \36884 );
buf \U$36907 ( \36886 , \36885 );
nand \U$36908 ( \36887 , \36881 , \36886 );
buf \U$36909 ( \36888 , \36887 );
buf \U$36910 ( \36889 , \36888 );
nand \U$36911 ( \36890 , \36880 , \36889 );
buf \U$36912 ( \36891 , \36890 );
xor \U$36913 ( \36892 , \36875 , \36891 );
buf \U$36914 ( \36893 , \35824 );
not \U$36915 ( \36894 , \36893 );
buf \U$36916 ( \36895 , \1183 );
not \U$36917 ( \36896 , \36895 );
or \U$36918 ( \36897 , \36894 , \36896 );
buf \U$36919 ( \36898 , \6141 );
xor \U$36920 ( \36899 , RIc0d9a18_77, RIc0d8410_30);
buf \U$36921 ( \36900 , \36899 );
nand \U$36922 ( \36901 , \36898 , \36900 );
buf \U$36923 ( \36902 , \36901 );
buf \U$36924 ( \36903 , \36902 );
nand \U$36925 ( \36904 , \36897 , \36903 );
buf \U$36926 ( \36905 , \36904 );
xor \U$36927 ( \36906 , \36892 , \36905 );
buf \U$36928 ( \36907 , \36906 );
buf \U$36929 ( \36908 , \35846 );
not \U$36930 ( \36909 , \36908 );
buf \U$36931 ( \36910 , \809 );
not \U$36932 ( \36911 , \36910 );
or \U$36933 ( \36912 , \36909 , \36911 );
buf \U$36934 ( \36913 , \816 );
buf \U$36935 ( \36914 , RIc0d9ec8_87);
buf \U$36936 ( \36915 , RIc0d7f60_20);
xor \U$36937 ( \36916 , \36914 , \36915 );
buf \U$36938 ( \36917 , \36916 );
buf \U$36939 ( \36918 , \36917 );
nand \U$36940 ( \36919 , \36913 , \36918 );
buf \U$36941 ( \36920 , \36919 );
buf \U$36942 ( \36921 , \36920 );
nand \U$36943 ( \36922 , \36912 , \36921 );
buf \U$36944 ( \36923 , \36922 );
buf \U$36945 ( \36924 , \35980 );
not \U$36946 ( \36925 , \36924 );
buf \U$36947 ( \36926 , \28794 );
not \U$36948 ( \36927 , \36926 );
or \U$36949 ( \36928 , \36925 , \36927 );
buf \U$36950 ( \36929 , \12342 );
buf \U$36951 ( \36930 , RIc0da828_107);
nand \U$36952 ( \36931 , \36929 , \36930 );
buf \U$36953 ( \36932 , \36931 );
buf \U$36954 ( \36933 , \36932 );
nand \U$36955 ( \36934 , \36928 , \36933 );
buf \U$36956 ( \36935 , \36934 );
xor \U$36957 ( \36936 , \36923 , \36935 );
buf \U$36958 ( \36937 , \35905 );
not \U$36959 ( \36938 , \36937 );
buf \U$36960 ( \36939 , \2871 );
not \U$36961 ( \36940 , \36939 );
or \U$36962 ( \36941 , \36938 , \36940 );
buf \U$36963 ( \36942 , \792 );
buf \U$36964 ( \36943 , RIc0d9838_73);
buf \U$36965 ( \36944 , RIc0d85f0_34);
xor \U$36966 ( \36945 , \36943 , \36944 );
buf \U$36967 ( \36946 , \36945 );
buf \U$36968 ( \36947 , \36946 );
nand \U$36969 ( \36948 , \36942 , \36947 );
buf \U$36970 ( \36949 , \36948 );
buf \U$36971 ( \36950 , \36949 );
nand \U$36972 ( \36951 , \36941 , \36950 );
buf \U$36973 ( \36952 , \36951 );
xor \U$36974 ( \36953 , \36936 , \36952 );
buf \U$36975 ( \36954 , \36953 );
xor \U$36976 ( \36955 , \36907 , \36954 );
xor \U$36977 ( \36956 , \35643 , \35714 );
and \U$36978 ( \36957 , \36956 , \35786 );
and \U$36979 ( \36958 , \35643 , \35714 );
or \U$36980 ( \36959 , \36957 , \36958 );
buf \U$36981 ( \36960 , \36959 );
buf \U$36982 ( \36961 , \36960 );
xor \U$36983 ( \36962 , \36955 , \36961 );
buf \U$36984 ( \36963 , \36962 );
buf \U$36985 ( \36964 , \36963 );
xor \U$36986 ( \36965 , \36859 , \36964 );
buf \U$36987 ( \36966 , \36643 );
not \U$36988 ( \36967 , \36966 );
buf \U$36989 ( \36968 , \36967 );
buf \U$36990 ( \36969 , \36968 );
xor \U$36991 ( \36970 , RIc0d9928_75, RIc0d8668_35);
buf \U$36992 ( \36971 , \36970 );
not \U$36993 ( \36972 , \36971 );
buf \U$36994 ( \36973 , \1125 );
not \U$36995 ( \36974 , \36973 );
buf \U$36996 ( \36975 , \36974 );
buf \U$36997 ( \36976 , \36975 );
not \U$36998 ( \36977 , \36976 );
or \U$36999 ( \36978 , \36972 , \36977 );
buf \U$37000 ( \36979 , \1143 );
buf \U$37001 ( \36980 , \35793 );
nand \U$37002 ( \36981 , \36979 , \36980 );
buf \U$37003 ( \36982 , \36981 );
buf \U$37004 ( \36983 , \36982 );
nand \U$37005 ( \36984 , \36978 , \36983 );
buf \U$37006 ( \36985 , \36984 );
buf \U$37007 ( \36986 , \36985 );
not \U$37008 ( \36987 , \36986 );
buf \U$37009 ( \36988 , \36802 );
not \U$37010 ( \36989 , \36988 );
buf \U$37011 ( \36990 , \36989 );
buf \U$37012 ( \36991 , \36990 );
not \U$37013 ( \36992 , \36991 );
buf \U$37014 ( \36993 , \1765 );
not \U$37015 ( \36994 , \36993 );
or \U$37016 ( \36995 , \36992 , \36994 );
buf \U$37017 ( \36996 , \3631 );
buf \U$37018 ( \36997 , \35836 );
nand \U$37019 ( \36998 , \36996 , \36997 );
buf \U$37020 ( \36999 , \36998 );
buf \U$37021 ( \37000 , \36999 );
nand \U$37022 ( \37001 , \36995 , \37000 );
buf \U$37023 ( \37002 , \37001 );
buf \U$37024 ( \37003 , \37002 );
not \U$37025 ( \37004 , \37003 );
or \U$37026 ( \37005 , \36987 , \37004 );
buf \U$37027 ( \37006 , \37002 );
buf \U$37028 ( \37007 , \36985 );
or \U$37029 ( \37008 , \37006 , \37007 );
buf \U$37030 ( \37009 , RIc0d7858_5);
buf \U$37031 ( \37010 , RIc0da738_105);
xor \U$37032 ( \37011 , \37009 , \37010 );
buf \U$37033 ( \37012 , \37011 );
buf \U$37034 ( \37013 , \37012 );
not \U$37035 ( \37014 , \37013 );
buf \U$37036 ( \37015 , \25475 );
not \U$37037 ( \37016 , \37015 );
or \U$37038 ( \37017 , \37014 , \37016 );
buf \U$37039 ( \37018 , \12744 );
buf \U$37040 ( \37019 , \36092 );
nand \U$37041 ( \37020 , \37018 , \37019 );
buf \U$37042 ( \37021 , \37020 );
buf \U$37043 ( \37022 , \37021 );
nand \U$37044 ( \37023 , \37017 , \37022 );
buf \U$37045 ( \37024 , \37023 );
buf \U$37046 ( \37025 , \37024 );
nand \U$37047 ( \37026 , \37008 , \37025 );
buf \U$37048 ( \37027 , \37026 );
buf \U$37049 ( \37028 , \37027 );
nand \U$37050 ( \37029 , \37005 , \37028 );
buf \U$37051 ( \37030 , \37029 );
buf \U$37052 ( \37031 , \37030 );
xor \U$37053 ( \37032 , \36969 , \37031 );
buf \U$37054 ( \37033 , RIc0d8938_41);
buf \U$37055 ( \37034 , RIc0d9658_69);
xor \U$37056 ( \37035 , \37033 , \37034 );
buf \U$37057 ( \37036 , \37035 );
buf \U$37058 ( \37037 , \37036 );
not \U$37059 ( \37038 , \37037 );
buf \U$37060 ( \37039 , \864 );
not \U$37061 ( \37040 , \37039 );
or \U$37062 ( \37041 , \37038 , \37040 );
buf \U$37063 ( \37042 , \284 );
buf \U$37064 ( \37043 , \35936 );
nand \U$37065 ( \37044 , \37042 , \37043 );
buf \U$37066 ( \37045 , \37044 );
buf \U$37067 ( \37046 , \37045 );
nand \U$37068 ( \37047 , \37041 , \37046 );
buf \U$37069 ( \37048 , \37047 );
buf \U$37070 ( \37049 , \37048 );
not \U$37071 ( \37050 , \37049 );
buf \U$37072 ( \37051 , \36730 );
not \U$37073 ( \37052 , \37051 );
buf \U$37074 ( \37053 , \13075 );
not \U$37075 ( \37054 , \37053 );
or \U$37076 ( \37055 , \37052 , \37054 );
buf \U$37077 ( \37056 , \1078 );
buf \U$37078 ( \37057 , \36027 );
nand \U$37079 ( \37058 , \37056 , \37057 );
buf \U$37080 ( \37059 , \37058 );
buf \U$37081 ( \37060 , \37059 );
nand \U$37082 ( \37061 , \37055 , \37060 );
buf \U$37083 ( \37062 , \37061 );
buf \U$37084 ( \37063 , \37062 );
not \U$37085 ( \37064 , \37063 );
or \U$37086 ( \37065 , \37050 , \37064 );
buf \U$37087 ( \37066 , \37062 );
buf \U$37088 ( \37067 , \37048 );
or \U$37089 ( \37068 , \37066 , \37067 );
buf \U$37090 ( \37069 , RIc0d8578_33);
buf \U$37091 ( \37070 , RIc0d9a18_77);
xor \U$37092 ( \37071 , \37069 , \37070 );
buf \U$37093 ( \37072 , \37071 );
buf \U$37094 ( \37073 , \37072 );
not \U$37095 ( \37074 , \37073 );
buf \U$37096 ( \37075 , \1183 );
not \U$37097 ( \37076 , \37075 );
or \U$37098 ( \37077 , \37074 , \37076 );
buf \U$37099 ( \37078 , \27267 );
buf \U$37100 ( \37079 , \35814 );
nand \U$37101 ( \37080 , \37078 , \37079 );
buf \U$37102 ( \37081 , \37080 );
buf \U$37103 ( \37082 , \37081 );
nand \U$37104 ( \37083 , \37077 , \37082 );
buf \U$37105 ( \37084 , \37083 );
buf \U$37106 ( \37085 , \37084 );
nand \U$37107 ( \37086 , \37068 , \37085 );
buf \U$37108 ( \37087 , \37086 );
buf \U$37109 ( \37088 , \37087 );
nand \U$37110 ( \37089 , \37065 , \37088 );
buf \U$37111 ( \37090 , \37089 );
buf \U$37112 ( \37091 , \37090 );
xnor \U$37113 ( \37092 , \37032 , \37091 );
buf \U$37114 ( \37093 , \37092 );
buf \U$37115 ( \37094 , \37093 );
not \U$37116 ( \37095 , \37094 );
buf \U$37117 ( \37096 , RIc0d7c18_13);
buf \U$37118 ( \37097 , RIc0da378_97);
xor \U$37119 ( \37098 , \37096 , \37097 );
buf \U$37120 ( \37099 , \37098 );
buf \U$37121 ( \37100 , \37099 );
not \U$37122 ( \37101 , \37100 );
buf \U$37123 ( \37102 , \15329 );
not \U$37124 ( \37103 , \37102 );
or \U$37125 ( \37104 , \37101 , \37103 );
buf \U$37126 ( \37105 , \2070 );
buf \U$37127 ( \37106 , RIc0d7ba0_12);
buf \U$37128 ( \37107 , RIc0da378_97);
xor \U$37129 ( \37108 , \37106 , \37107 );
buf \U$37130 ( \37109 , \37108 );
buf \U$37131 ( \37110 , \37109 );
nand \U$37132 ( \37111 , \37105 , \37110 );
buf \U$37133 ( \37112 , \37111 );
buf \U$37134 ( \37113 , \37112 );
nand \U$37135 ( \37114 , \37104 , \37113 );
buf \U$37136 ( \37115 , \37114 );
buf \U$37137 ( \37116 , \37115 );
buf \U$37138 ( \37117 , \36706 );
not \U$37139 ( \37118 , \37117 );
buf \U$37140 ( \37119 , \13419 );
not \U$37141 ( \37120 , \37119 );
or \U$37142 ( \37121 , \37118 , \37120 );
buf \U$37143 ( \37122 , \13426 );
buf \U$37144 ( \37123 , RIc0da918_109);
nand \U$37145 ( \37124 , \37122 , \37123 );
buf \U$37146 ( \37125 , \37124 );
buf \U$37147 ( \37126 , \37125 );
nand \U$37148 ( \37127 , \37121 , \37126 );
buf \U$37149 ( \37128 , \37127 );
buf \U$37150 ( \37129 , \37128 );
nor \U$37151 ( \37130 , \37116 , \37129 );
buf \U$37152 ( \37131 , \37130 );
buf \U$37153 ( \37132 , \37131 );
xor \U$37154 ( \37133 , RIc0d9ce8_83, RIc0d82a8_27);
buf \U$37155 ( \37134 , \37133 );
not \U$37156 ( \37135 , \37134 );
buf \U$37157 ( \37136 , \1736 );
not \U$37158 ( \37137 , \37136 );
or \U$37159 ( \37138 , \37135 , \37137 );
buf \U$37160 ( \37139 , \993 );
buf \U$37161 ( \37140 , \35953 );
nand \U$37162 ( \37141 , \37139 , \37140 );
buf \U$37163 ( \37142 , \37141 );
buf \U$37164 ( \37143 , \37142 );
nand \U$37165 ( \37144 , \37138 , \37143 );
buf \U$37166 ( \37145 , \37144 );
buf \U$37167 ( \37146 , \37145 );
not \U$37168 ( \37147 , \37146 );
buf \U$37169 ( \37148 , \37147 );
buf \U$37170 ( \37149 , \37148 );
or \U$37171 ( \37150 , \37132 , \37149 );
buf \U$37172 ( \37151 , \37115 );
buf \U$37173 ( \37152 , \37128 );
nand \U$37174 ( \37153 , \37151 , \37152 );
buf \U$37175 ( \37154 , \37153 );
buf \U$37176 ( \37155 , \37154 );
nand \U$37177 ( \37156 , \37150 , \37155 );
buf \U$37178 ( \37157 , \37156 );
buf \U$37179 ( \37158 , \37157 );
not \U$37180 ( \37159 , \37158 );
buf \U$37181 ( \37160 , RIc0d8758_37);
buf \U$37182 ( \37161 , RIc0d9838_73);
xor \U$37183 ( \37162 , \37160 , \37161 );
buf \U$37184 ( \37163 , \37162 );
buf \U$37185 ( \37164 , \37163 );
not \U$37186 ( \37165 , \37164 );
buf \U$37187 ( \37166 , \1677 );
not \U$37188 ( \37167 , \37166 );
or \U$37189 ( \37168 , \37165 , \37167 );
buf \U$37190 ( \37169 , \791 );
buf \U$37191 ( \37170 , \35895 );
nand \U$37192 ( \37171 , \37169 , \37170 );
buf \U$37193 ( \37172 , \37171 );
buf \U$37194 ( \37173 , \37172 );
nand \U$37195 ( \37174 , \37168 , \37173 );
buf \U$37196 ( \37175 , \37174 );
buf \U$37197 ( \37176 , \37175 );
xor \U$37198 ( \37177 , RIc0d9568_67, RIc0d8a28_43);
buf \U$37199 ( \37178 , \37177 );
not \U$37200 ( \37179 , \37178 );
buf \U$37201 ( \37180 , \4907 );
not \U$37202 ( \37181 , \37180 );
or \U$37203 ( \37182 , \37179 , \37181 );
buf \U$37204 ( \37183 , \686 );
buf \U$37205 ( \37184 , \36132 );
nand \U$37206 ( \37185 , \37183 , \37184 );
buf \U$37207 ( \37186 , \37185 );
buf \U$37208 ( \37187 , \37186 );
nand \U$37209 ( \37188 , \37182 , \37187 );
buf \U$37210 ( \37189 , \37188 );
buf \U$37211 ( \37190 , \37189 );
or \U$37212 ( \37191 , \37176 , \37190 );
buf \U$37213 ( \37192 , RIc0d7ee8_19);
buf \U$37214 ( \37193 , RIc0da0a8_91);
xor \U$37215 ( \37194 , \37192 , \37193 );
buf \U$37216 ( \37195 , \37194 );
buf \U$37217 ( \37196 , \37195 );
not \U$37218 ( \37197 , \37196 );
buf \U$37219 ( \37198 , \16402 );
not \U$37220 ( \37199 , \37198 );
or \U$37221 ( \37200 , \37197 , \37199 );
buf \U$37222 ( \37201 , \1933 );
buf \U$37223 ( \37202 , \36154 );
nand \U$37224 ( \37203 , \37201 , \37202 );
buf \U$37225 ( \37204 , \37203 );
buf \U$37226 ( \37205 , \37204 );
nand \U$37227 ( \37206 , \37200 , \37205 );
buf \U$37228 ( \37207 , \37206 );
buf \U$37229 ( \37208 , \37207 );
nand \U$37230 ( \37209 , \37191 , \37208 );
buf \U$37231 ( \37210 , \37209 );
buf \U$37232 ( \37211 , \37210 );
buf \U$37233 ( \37212 , \37175 );
buf \U$37234 ( \37213 , \37189 );
nand \U$37235 ( \37214 , \37212 , \37213 );
buf \U$37236 ( \37215 , \37214 );
buf \U$37237 ( \37216 , \37215 );
nand \U$37238 ( \37217 , \37211 , \37216 );
buf \U$37239 ( \37218 , \37217 );
buf \U$37240 ( \37219 , \37218 );
not \U$37241 ( \37220 , \37219 );
buf \U$37242 ( \37221 , \37220 );
buf \U$37243 ( \37222 , \37221 );
not \U$37244 ( \37223 , \37222 );
or \U$37245 ( \37224 , \37159 , \37223 );
buf \U$37246 ( \37225 , \37221 );
buf \U$37247 ( \37226 , \37157 );
or \U$37248 ( \37227 , \37225 , \37226 );
nand \U$37249 ( \37228 , \37224 , \37227 );
buf \U$37250 ( \37229 , \37228 );
buf \U$37251 ( \37230 , \37229 );
not \U$37252 ( \37231 , \37230 );
buf \U$37253 ( \37232 , \37109 );
not \U$37254 ( \37233 , \37232 );
buf \U$37255 ( \37234 , \2941 );
not \U$37256 ( \37235 , \37234 );
or \U$37257 ( \37236 , \37233 , \37235 );
buf \U$37258 ( \37237 , \2070 );
buf \U$37259 ( \37238 , \36368 );
nand \U$37260 ( \37239 , \37237 , \37238 );
buf \U$37261 ( \37240 , \37239 );
buf \U$37262 ( \37241 , \37240 );
nand \U$37263 ( \37242 , \37236 , \37241 );
buf \U$37264 ( \37243 , \37242 );
buf \U$37265 ( \37244 , \35603 );
not \U$37266 ( \37245 , \37244 );
buf \U$37267 ( \37246 , \12795 );
not \U$37268 ( \37247 , \37246 );
or \U$37269 ( \37248 , \37245 , \37247 );
buf \U$37270 ( \37249 , \1229 );
buf \U$37271 ( \37250 , \36490 );
nand \U$37272 ( \37251 , \37249 , \37250 );
buf \U$37273 ( \37252 , \37251 );
buf \U$37274 ( \37253 , \37252 );
nand \U$37275 ( \37254 , \37248 , \37253 );
buf \U$37276 ( \37255 , \37254 );
xor \U$37277 ( \37256 , \37243 , \37255 );
buf \U$37278 ( \37257 , \37256 );
not \U$37279 ( \37258 , \37257 );
buf \U$37280 ( \37259 , \2815 );
not \U$37281 ( \37260 , \37259 );
buf \U$37282 ( \37261 , \35678 );
not \U$37283 ( \37262 , \37261 );
buf \U$37284 ( \37263 , \37262 );
buf \U$37285 ( \37264 , \37263 );
not \U$37286 ( \37265 , \37264 );
and \U$37287 ( \37266 , \37260 , \37265 );
buf \U$37288 ( \37267 , \36332 );
not \U$37289 ( \37268 , \37267 );
buf \U$37290 ( \37269 , \18274 );
nor \U$37291 ( \37270 , \37268 , \37269 );
buf \U$37292 ( \37271 , \37270 );
buf \U$37293 ( \37272 , \37271 );
nor \U$37294 ( \37273 , \37266 , \37272 );
buf \U$37295 ( \37274 , \37273 );
buf \U$37296 ( \37275 , \37274 );
not \U$37297 ( \37276 , \37275 );
and \U$37298 ( \37277 , \37258 , \37276 );
buf \U$37299 ( \37278 , \37256 );
buf \U$37300 ( \37279 , \37274 );
and \U$37301 ( \37280 , \37278 , \37279 );
nor \U$37302 ( \37281 , \37277 , \37280 );
buf \U$37303 ( \37282 , \37281 );
buf \U$37304 ( \37283 , \37282 );
not \U$37305 ( \37284 , \37283 );
and \U$37306 ( \37285 , \37231 , \37284 );
buf \U$37307 ( \37286 , \37229 );
buf \U$37308 ( \37287 , \37282 );
and \U$37309 ( \37288 , \37286 , \37287 );
nor \U$37310 ( \37289 , \37285 , \37288 );
buf \U$37311 ( \37290 , \37289 );
buf \U$37312 ( \37291 , \37290 );
not \U$37313 ( \37292 , \37291 );
or \U$37314 ( \37293 , \37095 , \37292 );
xor \U$37315 ( \37294 , \35687 , \35706 );
xor \U$37316 ( \37295 , \37294 , \35663 );
buf \U$37317 ( \37296 , \37295 );
not \U$37318 ( \37297 , \37296 );
buf \U$37319 ( \37298 , \37297 );
buf \U$37320 ( \37299 , \37298 );
not \U$37321 ( \37300 , \37299 );
and \U$37322 ( \37301 , \35618 , \35614 );
not \U$37323 ( \37302 , \35618 );
and \U$37324 ( \37303 , \37302 , \35609 );
or \U$37325 ( \37304 , \37301 , \37303 );
xor \U$37326 ( \37305 , \37304 , \35640 );
buf \U$37327 ( \37306 , \37305 );
not \U$37328 ( \37307 , \37306 );
buf \U$37329 ( \37308 , \37307 );
buf \U$37330 ( \37309 , \37308 );
not \U$37331 ( \37310 , \37309 );
or \U$37332 ( \37311 , \37300 , \37310 );
buf \U$37333 ( \37312 , \37295 );
not \U$37334 ( \37313 , \37312 );
buf \U$37335 ( \37314 , \37305 );
not \U$37336 ( \37315 , \37314 );
or \U$37337 ( \37316 , \37313 , \37315 );
xor \U$37338 ( \37317 , \37207 , \37175 );
buf \U$37339 ( \37318 , \37317 );
buf \U$37340 ( \37319 , \37189 );
and \U$37341 ( \37320 , \37318 , \37319 );
not \U$37342 ( \37321 , \37318 );
buf \U$37343 ( \37322 , \37189 );
not \U$37344 ( \37323 , \37322 );
buf \U$37345 ( \37324 , \37323 );
buf \U$37346 ( \37325 , \37324 );
and \U$37347 ( \37326 , \37321 , \37325 );
nor \U$37348 ( \37327 , \37320 , \37326 );
buf \U$37349 ( \37328 , \37327 );
buf \U$37350 ( \37329 , \37328 );
nand \U$37351 ( \37330 , \37316 , \37329 );
buf \U$37352 ( \37331 , \37330 );
buf \U$37353 ( \37332 , \37331 );
nand \U$37354 ( \37333 , \37311 , \37332 );
buf \U$37355 ( \37334 , \37333 );
buf \U$37356 ( \37335 , \37334 );
nand \U$37357 ( \37336 , \37293 , \37335 );
buf \U$37358 ( \37337 , \37336 );
buf \U$37359 ( \37338 , \37337 );
not \U$37360 ( \37339 , \37290 );
buf \U$37361 ( \37340 , \37093 );
not \U$37362 ( \37341 , \37340 );
buf \U$37363 ( \37342 , \37341 );
nand \U$37364 ( \37343 , \37339 , \37342 );
buf \U$37365 ( \37344 , \37343 );
nand \U$37366 ( \37345 , \37338 , \37344 );
buf \U$37367 ( \37346 , \37345 );
buf \U$37368 ( \37347 , \37346 );
xor \U$37369 ( \37348 , \36965 , \37347 );
buf \U$37370 ( \37349 , \37348 );
xnor \U$37371 ( \37350 , \36600 , \37349 );
buf \U$37372 ( \37351 , \37350 );
not \U$37373 ( \37352 , \37351 );
buf \U$37374 ( \37353 , RIc0d86e0_36);
buf \U$37375 ( \37354 , RIc0d9928_75);
xor \U$37376 ( \37355 , \37353 , \37354 );
buf \U$37377 ( \37356 , \37355 );
buf \U$37378 ( \37357 , \37356 );
not \U$37379 ( \37358 , \37357 );
buf \U$37380 ( \37359 , \2358 );
not \U$37381 ( \37360 , \37359 );
or \U$37382 ( \37361 , \37358 , \37360 );
buf \U$37383 ( \37362 , \16500 );
buf \U$37384 ( \37363 , \36970 );
nand \U$37385 ( \37364 , \37362 , \37363 );
buf \U$37386 ( \37365 , \37364 );
buf \U$37387 ( \37366 , \37365 );
nand \U$37388 ( \37367 , \37361 , \37366 );
buf \U$37389 ( \37368 , \37367 );
buf \U$37390 ( \37369 , \37368 );
not \U$37391 ( \37370 , \37369 );
buf \U$37392 ( \37371 , RIc0d9838_73);
buf \U$37393 ( \37372 , RIc0d87d0_38);
xor \U$37394 ( \37373 , \37371 , \37372 );
buf \U$37395 ( \37374 , \37373 );
buf \U$37396 ( \37375 , \37374 );
not \U$37397 ( \37376 , \37375 );
buf \U$37398 ( \37377 , \12442 );
not \U$37399 ( \37378 , \37377 );
or \U$37400 ( \37379 , \37376 , \37378 );
buf \U$37401 ( \37380 , \791 );
buf \U$37402 ( \37381 , \37163 );
nand \U$37403 ( \37382 , \37380 , \37381 );
buf \U$37404 ( \37383 , \37382 );
buf \U$37405 ( \37384 , \37383 );
nand \U$37406 ( \37385 , \37379 , \37384 );
buf \U$37407 ( \37386 , \37385 );
buf \U$37408 ( \37387 , \37386 );
not \U$37409 ( \37388 , \37387 );
or \U$37410 ( \37389 , \37370 , \37388 );
buf \U$37411 ( \37390 , \37386 );
buf \U$37412 ( \37391 , \37368 );
or \U$37413 ( \37392 , \37390 , \37391 );
buf \U$37414 ( \37393 , RIc0d9a18_77);
buf \U$37415 ( \37394 , RIc0d85f0_34);
xor \U$37416 ( \37395 , \37393 , \37394 );
buf \U$37417 ( \37396 , \37395 );
buf \U$37418 ( \37397 , \37396 );
not \U$37419 ( \37398 , \37397 );
buf \U$37420 ( \37399 , \1432 );
not \U$37421 ( \37400 , \37399 );
or \U$37422 ( \37401 , \37398 , \37400 );
buf \U$37423 ( \37402 , \1196 );
buf \U$37424 ( \37403 , \37072 );
nand \U$37425 ( \37404 , \37402 , \37403 );
buf \U$37426 ( \37405 , \37404 );
buf \U$37427 ( \37406 , \37405 );
nand \U$37428 ( \37407 , \37401 , \37406 );
buf \U$37429 ( \37408 , \37407 );
buf \U$37430 ( \37409 , \37408 );
nand \U$37431 ( \37410 , \37392 , \37409 );
buf \U$37432 ( \37411 , \37410 );
buf \U$37433 ( \37412 , \37411 );
nand \U$37434 ( \37413 , \37389 , \37412 );
buf \U$37435 ( \37414 , \37413 );
buf \U$37436 ( \37415 , \37414 );
not \U$37437 ( \37416 , \37415 );
buf \U$37438 ( \37417 , \37416 );
buf \U$37439 ( \37418 , \37417 );
not \U$37440 ( \37419 , \37418 );
buf \U$37441 ( \37420 , RIc0d9748_71);
buf \U$37442 ( \37421 , RIc0d88c0_40);
xor \U$37443 ( \37422 , \37420 , \37421 );
buf \U$37444 ( \37423 , \37422 );
buf \U$37445 ( \37424 , \37423 );
not \U$37446 ( \37425 , \37424 );
buf \U$37447 ( \37426 , \2269 );
not \U$37448 ( \37427 , \37426 );
or \U$37449 ( \37428 , \37425 , \37427 );
buf \U$37450 ( \37429 , \1282 );
buf \U$37451 ( \37430 , \35668 );
nand \U$37452 ( \37431 , \37429 , \37430 );
buf \U$37453 ( \37432 , \37431 );
buf \U$37454 ( \37433 , \37432 );
nand \U$37455 ( \37434 , \37428 , \37433 );
buf \U$37456 ( \37435 , \37434 );
buf \U$37457 ( \37436 , \37435 );
not \U$37458 ( \37437 , \37436 );
xor \U$37459 ( \37438 , \36601 , \36602 );
buf \U$37460 ( \37439 , \37438 );
buf \U$37461 ( \37440 , \37439 );
not \U$37462 ( \37441 , \37440 );
buf \U$37463 ( \37442 , \12795 );
not \U$37464 ( \37443 , \37442 );
or \U$37465 ( \37444 , \37441 , \37443 );
buf \U$37466 ( \37445 , \1229 );
buf \U$37467 ( \37446 , \35593 );
nand \U$37468 ( \37447 , \37445 , \37446 );
buf \U$37469 ( \37448 , \37447 );
buf \U$37470 ( \37449 , \37448 );
nand \U$37471 ( \37450 , \37444 , \37449 );
buf \U$37472 ( \37451 , \37450 );
buf \U$37473 ( \37452 , \37451 );
not \U$37474 ( \37453 , \37452 );
or \U$37475 ( \37454 , \37437 , \37453 );
buf \U$37476 ( \37455 , \37435 );
not \U$37477 ( \37456 , \37455 );
buf \U$37478 ( \37457 , \37456 );
buf \U$37479 ( \37458 , \37457 );
not \U$37480 ( \37459 , \37458 );
buf \U$37481 ( \37460 , \37451 );
not \U$37482 ( \37461 , \37460 );
buf \U$37483 ( \37462 , \37461 );
buf \U$37484 ( \37463 , \37462 );
not \U$37485 ( \37464 , \37463 );
or \U$37486 ( \37465 , \37459 , \37464 );
buf \U$37487 ( \37466 , RIc0da378_97);
buf \U$37488 ( \37467 , RIc0d7c90_14);
xor \U$37489 ( \37468 , \37466 , \37467 );
buf \U$37490 ( \37469 , \37468 );
buf \U$37491 ( \37470 , \37469 );
not \U$37492 ( \37471 , \37470 );
buf \U$37493 ( \37472 , \2941 );
not \U$37494 ( \37473 , \37472 );
or \U$37495 ( \37474 , \37471 , \37473 );
buf \U$37496 ( \37475 , \734 );
buf \U$37497 ( \37476 , \37099 );
nand \U$37498 ( \37477 , \37475 , \37476 );
buf \U$37499 ( \37478 , \37477 );
buf \U$37500 ( \37479 , \37478 );
nand \U$37501 ( \37480 , \37474 , \37479 );
buf \U$37502 ( \37481 , \37480 );
buf \U$37503 ( \37482 , \37481 );
nand \U$37504 ( \37483 , \37465 , \37482 );
buf \U$37505 ( \37484 , \37483 );
buf \U$37506 ( \37485 , \37484 );
nand \U$37507 ( \37486 , \37454 , \37485 );
buf \U$37508 ( \37487 , \37486 );
buf \U$37509 ( \37488 , \37487 );
not \U$37510 ( \37489 , \37488 );
buf \U$37511 ( \37490 , \37489 );
buf \U$37512 ( \37491 , \37490 );
not \U$37513 ( \37492 , \37491 );
or \U$37514 ( \37493 , \37419 , \37492 );
buf \U$37515 ( \37494 , RIc0d9ce8_83);
buf \U$37516 ( \37495 , RIc0d8320_28);
xor \U$37517 ( \37496 , \37494 , \37495 );
buf \U$37518 ( \37497 , \37496 );
buf \U$37519 ( \37498 , \37497 );
not \U$37520 ( \37499 , \37498 );
buf \U$37521 ( \37500 , \1736 );
not \U$37522 ( \37501 , \37500 );
or \U$37523 ( \37502 , \37499 , \37501 );
buf \U$37524 ( \37503 , \584 );
buf \U$37525 ( \37504 , \37133 );
nand \U$37526 ( \37505 , \37503 , \37504 );
buf \U$37527 ( \37506 , \37505 );
buf \U$37528 ( \37507 , \37506 );
nand \U$37529 ( \37508 , \37502 , \37507 );
buf \U$37530 ( \37509 , \37508 );
buf \U$37531 ( \37510 , \37509 );
buf \U$37532 ( \37511 , RIc0d89b0_42);
buf \U$37533 ( \37512 , RIc0d9658_69);
xor \U$37534 ( \37513 , \37511 , \37512 );
buf \U$37535 ( \37514 , \37513 );
buf \U$37536 ( \37515 , \37514 );
not \U$37537 ( \37516 , \37515 );
buf \U$37538 ( \37517 , \864 );
not \U$37539 ( \37518 , \37517 );
or \U$37540 ( \37519 , \37516 , \37518 );
buf \U$37541 ( \37520 , \284 );
buf \U$37542 ( \37521 , \37036 );
nand \U$37543 ( \37522 , \37520 , \37521 );
buf \U$37544 ( \37523 , \37522 );
buf \U$37545 ( \37524 , \37523 );
nand \U$37546 ( \37525 , \37519 , \37524 );
buf \U$37547 ( \37526 , \37525 );
buf \U$37548 ( \37527 , \37526 );
xor \U$37549 ( \37528 , \37510 , \37527 );
xor \U$37550 ( \37529 , RIc0da828_107, RIc0d77e0_4);
buf \U$37551 ( \37530 , \37529 );
not \U$37552 ( \37531 , \37530 );
buf \U$37553 ( \37532 , \12331 );
not \U$37554 ( \37533 , \37532 );
buf \U$37555 ( \37534 , \37533 );
buf \U$37556 ( \37535 , \37534 );
not \U$37557 ( \37536 , \37535 );
or \U$37558 ( \37537 , \37531 , \37536 );
buf \U$37559 ( \37538 , \12342 );
buf \U$37560 ( \37539 , \35744 );
nand \U$37561 ( \37540 , \37538 , \37539 );
buf \U$37562 ( \37541 , \37540 );
buf \U$37563 ( \37542 , \37541 );
nand \U$37564 ( \37543 , \37537 , \37542 );
buf \U$37565 ( \37544 , \37543 );
buf \U$37566 ( \37545 , \37544 );
and \U$37567 ( \37546 , \37528 , \37545 );
and \U$37568 ( \37547 , \37510 , \37527 );
or \U$37569 ( \37548 , \37546 , \37547 );
buf \U$37570 ( \37549 , \37548 );
buf \U$37571 ( \37550 , \37549 );
nand \U$37572 ( \37551 , \37493 , \37550 );
buf \U$37573 ( \37552 , \37551 );
buf \U$37574 ( \37553 , \37552 );
buf \U$37575 ( \37554 , \37414 );
buf \U$37576 ( \37555 , \37487 );
nand \U$37577 ( \37556 , \37554 , \37555 );
buf \U$37578 ( \37557 , \37556 );
buf \U$37579 ( \37558 , \37557 );
nand \U$37580 ( \37559 , \37553 , \37558 );
buf \U$37581 ( \37560 , \37559 );
buf \U$37582 ( \37561 , \37560 );
buf \U$37583 ( \37562 , \37115 );
buf \U$37584 ( \37563 , \37128 );
xor \U$37585 ( \37564 , \37562 , \37563 );
buf \U$37586 ( \37565 , \37564 );
buf \U$37587 ( \37566 , \37565 );
buf \U$37588 ( \37567 , \37145 );
and \U$37589 ( \37568 , \37566 , \37567 );
not \U$37590 ( \37569 , \37566 );
buf \U$37591 ( \37570 , \37148 );
and \U$37592 ( \37571 , \37569 , \37570 );
nor \U$37593 ( \37572 , \37568 , \37571 );
buf \U$37594 ( \37573 , \37572 );
buf \U$37595 ( \37574 , \37573 );
not \U$37596 ( \37575 , \37574 );
xor \U$37597 ( \37576 , \37048 , \37062 );
buf \U$37598 ( \37577 , \37576 );
buf \U$37599 ( \37578 , \37084 );
xor \U$37600 ( \37579 , \37577 , \37578 );
buf \U$37601 ( \37580 , \37579 );
buf \U$37602 ( \37581 , \37580 );
not \U$37603 ( \37582 , \37581 );
or \U$37604 ( \37583 , \37575 , \37582 );
buf \U$37605 ( \37584 , \37580 );
buf \U$37606 ( \37585 , \37573 );
or \U$37607 ( \37586 , \37584 , \37585 );
buf \U$37608 ( \37587 , \37002 );
not \U$37609 ( \37588 , \37587 );
buf \U$37610 ( \37589 , \37024 );
not \U$37611 ( \37590 , \37589 );
buf \U$37612 ( \37591 , \37590 );
buf \U$37613 ( \37592 , \37591 );
not \U$37614 ( \37593 , \37592 );
or \U$37615 ( \37594 , \37588 , \37593 );
buf \U$37616 ( \37595 , \37002 );
not \U$37617 ( \37596 , \37595 );
buf \U$37618 ( \37597 , \37024 );
nand \U$37619 ( \37598 , \37596 , \37597 );
buf \U$37620 ( \37599 , \37598 );
buf \U$37621 ( \37600 , \37599 );
nand \U$37622 ( \37601 , \37594 , \37600 );
buf \U$37623 ( \37602 , \37601 );
buf \U$37624 ( \37603 , \37602 );
buf \U$37625 ( \37604 , \36985 );
not \U$37626 ( \37605 , \37604 );
buf \U$37627 ( \37606 , \37605 );
buf \U$37628 ( \37607 , \37606 );
and \U$37629 ( \37608 , \37603 , \37607 );
not \U$37630 ( \37609 , \37603 );
buf \U$37631 ( \37610 , \36985 );
and \U$37632 ( \37611 , \37609 , \37610 );
nor \U$37633 ( \37612 , \37608 , \37611 );
buf \U$37634 ( \37613 , \37612 );
buf \U$37635 ( \37614 , \37613 );
not \U$37636 ( \37615 , \37614 );
buf \U$37637 ( \37616 , \37615 );
buf \U$37638 ( \37617 , \37616 );
nand \U$37639 ( \37618 , \37586 , \37617 );
buf \U$37640 ( \37619 , \37618 );
buf \U$37641 ( \37620 , \37619 );
nand \U$37642 ( \37621 , \37583 , \37620 );
buf \U$37643 ( \37622 , \37621 );
buf \U$37644 ( \37623 , \37622 );
xor \U$37645 ( \37624 , \37561 , \37623 );
and \U$37646 ( \37625 , \33956 , \33957 );
buf \U$37647 ( \37626 , \37625 );
buf \U$37648 ( \37627 , \37626 );
xor \U$37649 ( \37628 , RIc0d9568_67, RIc0d8aa0_44);
buf \U$37650 ( \37629 , \37628 );
not \U$37651 ( \37630 , \37629 );
buf \U$37652 ( \37631 , \1823 );
not \U$37653 ( \37632 , \37631 );
or \U$37654 ( \37633 , \37630 , \37632 );
buf \U$37655 ( \37634 , \686 );
buf \U$37656 ( \37635 , \37177 );
nand \U$37657 ( \37636 , \37634 , \37635 );
buf \U$37658 ( \37637 , \37636 );
buf \U$37659 ( \37638 , \37637 );
nand \U$37660 ( \37639 , \37633 , \37638 );
buf \U$37661 ( \37640 , \37639 );
buf \U$37662 ( \37641 , \37640 );
xor \U$37663 ( \37642 , \37627 , \37641 );
buf \U$37664 ( \37643 , RIc0d7f60_20);
buf \U$37665 ( \37644 , RIc0da0a8_91);
xnor \U$37666 ( \37645 , \37643 , \37644 );
buf \U$37667 ( \37646 , \37645 );
buf \U$37668 ( \37647 , \37646 );
not \U$37669 ( \37648 , \37647 );
buf \U$37670 ( \37649 , \37648 );
buf \U$37671 ( \37650 , \37649 );
not \U$37672 ( \37651 , \37650 );
buf \U$37673 ( \37652 , \704 );
not \U$37674 ( \37653 , \37652 );
or \U$37675 ( \37654 , \37651 , \37653 );
buf \U$37676 ( \37655 , \13293 );
buf \U$37677 ( \37656 , \37195 );
nand \U$37678 ( \37657 , \37655 , \37656 );
buf \U$37679 ( \37658 , \37657 );
buf \U$37680 ( \37659 , \37658 );
nand \U$37681 ( \37660 , \37654 , \37659 );
buf \U$37682 ( \37661 , \37660 );
buf \U$37683 ( \37662 , \37661 );
and \U$37684 ( \37663 , \37642 , \37662 );
and \U$37685 ( \37664 , \37627 , \37641 );
or \U$37686 ( \37665 , \37663 , \37664 );
buf \U$37687 ( \37666 , \37665 );
buf \U$37688 ( \37667 , \37666 );
xor \U$37689 ( \37668 , RIc0da468_99, RIc0d7ba0_12);
buf \U$37690 ( \37669 , \37668 );
not \U$37691 ( \37670 , \37669 );
buf \U$37692 ( \37671 , \21461 );
not \U$37693 ( \37672 , \37671 );
or \U$37694 ( \37673 , \37670 , \37672 );
buf \U$37695 ( \37674 , \14648 );
buf \U$37696 ( \37675 , \35693 );
nand \U$37697 ( \37676 , \37674 , \37675 );
buf \U$37698 ( \37677 , \37676 );
buf \U$37699 ( \37678 , \37677 );
nand \U$37700 ( \37679 , \37673 , \37678 );
buf \U$37701 ( \37680 , \37679 );
buf \U$37702 ( \37681 , \37680 );
buf \U$37703 ( \37682 , RIc0d8230_26);
buf \U$37704 ( \37683 , RIc0d9dd8_85);
xor \U$37705 ( \37684 , \37682 , \37683 );
buf \U$37706 ( \37685 , \37684 );
buf \U$37707 ( \37686 , \37685 );
not \U$37708 ( \37687 , \37686 );
buf \U$37709 ( \37688 , \6029 );
not \U$37710 ( \37689 , \37688 );
or \U$37711 ( \37690 , \37687 , \37689 );
buf \U$37712 ( \37691 , \2960 );
buf \U$37713 ( \37692 , \35647 );
nand \U$37714 ( \37693 , \37691 , \37692 );
buf \U$37715 ( \37694 , \37693 );
buf \U$37716 ( \37695 , \37694 );
nand \U$37717 ( \37696 , \37690 , \37695 );
buf \U$37718 ( \37697 , \37696 );
buf \U$37719 ( \37698 , \37697 );
xor \U$37720 ( \37699 , \37681 , \37698 );
buf \U$37721 ( \37700 , \12541 );
not \U$37722 ( \37701 , \37700 );
buf \U$37723 ( \37702 , \18306 );
not \U$37724 ( \37703 , \37702 );
buf \U$37725 ( \37704 , \37703 );
buf \U$37726 ( \37705 , \37704 );
not \U$37727 ( \37706 , \37705 );
or \U$37728 ( \37707 , \37701 , \37706 );
buf \U$37729 ( \37708 , RIc0daa08_111);
nand \U$37730 ( \37709 , \37707 , \37708 );
buf \U$37731 ( \37710 , \37709 );
buf \U$37732 ( \37711 , \37710 );
and \U$37733 ( \37712 , \37699 , \37711 );
and \U$37734 ( \37713 , \37681 , \37698 );
or \U$37735 ( \37714 , \37712 , \37713 );
buf \U$37736 ( \37715 , \37714 );
buf \U$37737 ( \37716 , \37715 );
xor \U$37738 ( \37717 , \37667 , \37716 );
xor \U$37739 ( \37718 , \35736 , \35758 );
xor \U$37740 ( \37719 , \37718 , \35781 );
buf \U$37741 ( \37720 , \37719 );
buf \U$37742 ( \37721 , \37720 );
and \U$37743 ( \37722 , \37717 , \37721 );
and \U$37744 ( \37723 , \37667 , \37716 );
or \U$37745 ( \37724 , \37722 , \37723 );
buf \U$37746 ( \37725 , \37724 );
buf \U$37747 ( \37726 , \37725 );
xor \U$37748 ( \37727 , \37624 , \37726 );
buf \U$37749 ( \37728 , \37727 );
buf \U$37750 ( \37729 , \37728 );
xor \U$37751 ( \37730 , \35789 , \35991 );
xor \U$37752 ( \37731 , \37730 , \36177 );
buf \U$37753 ( \37732 , \37731 );
buf \U$37754 ( \37733 , \37732 );
xor \U$37755 ( \37734 , \37729 , \37733 );
xor \U$37756 ( \37735 , \36605 , \36622 );
xor \U$37757 ( \37736 , \37735 , \36644 );
buf \U$37758 ( \37737 , \37736 );
buf \U$37759 ( \37738 , \37737 );
buf \U$37760 ( \37739 , \34099 );
not \U$37761 ( \37740 , \37739 );
buf \U$37762 ( \37741 , \4527 );
not \U$37763 ( \37742 , \37741 );
or \U$37764 ( \37743 , \37740 , \37742 );
buf \U$37765 ( \37744 , \36795 );
not \U$37766 ( \37745 , \37744 );
buf \U$37767 ( \37746 , \816 );
nand \U$37768 ( \37747 , \37745 , \37746 );
buf \U$37769 ( \37748 , \37747 );
buf \U$37770 ( \37749 , \37748 );
nand \U$37771 ( \37750 , \37743 , \37749 );
buf \U$37772 ( \37751 , \37750 );
buf \U$37773 ( \37752 , \37751 );
buf \U$37774 ( \37753 , RIc0da738_105);
buf \U$37775 ( \37754 , RIc0d78d0_6);
xor \U$37776 ( \37755 , \37753 , \37754 );
buf \U$37777 ( \37756 , \37755 );
buf \U$37778 ( \37757 , \37756 );
not \U$37779 ( \37758 , \37757 );
buf \U$37780 ( \37759 , \12736 );
not \U$37781 ( \37760 , \37759 );
or \U$37782 ( \37761 , \37758 , \37760 );
buf \U$37783 ( \37762 , \12744 );
buf \U$37784 ( \37763 , \37012 );
nand \U$37785 ( \37764 , \37762 , \37763 );
buf \U$37786 ( \37765 , \37764 );
buf \U$37787 ( \37766 , \37765 );
nand \U$37788 ( \37767 , \37761 , \37766 );
buf \U$37789 ( \37768 , \37767 );
buf \U$37790 ( \37769 , \37768 );
xor \U$37791 ( \37770 , \37752 , \37769 );
buf \U$37792 ( \37771 , \8209 );
not \U$37793 ( \37772 , \37771 );
buf \U$37794 ( \37773 , \33992 );
not \U$37795 ( \37774 , \37773 );
and \U$37796 ( \37775 , \37772 , \37774 );
buf \U$37797 ( \37776 , \686 );
buf \U$37798 ( \37777 , \37628 );
and \U$37799 ( \37778 , \37776 , \37777 );
nor \U$37800 ( \37779 , \37775 , \37778 );
buf \U$37801 ( \37780 , \37779 );
buf \U$37802 ( \37781 , \37780 );
not \U$37803 ( \37782 , \37781 );
buf \U$37804 ( \37783 , \34082 );
not \U$37805 ( \37784 , \37783 );
buf \U$37806 ( \37785 , \12442 );
not \U$37807 ( \37786 , \37785 );
or \U$37808 ( \37787 , \37784 , \37786 );
buf \U$37809 ( \37788 , \2882 );
buf \U$37810 ( \37789 , \37374 );
nand \U$37811 ( \37790 , \37788 , \37789 );
buf \U$37812 ( \37791 , \37790 );
buf \U$37813 ( \37792 , \37791 );
nand \U$37814 ( \37793 , \37787 , \37792 );
buf \U$37815 ( \37794 , \37793 );
buf \U$37816 ( \37795 , \37794 );
not \U$37817 ( \37796 , \37795 );
buf \U$37818 ( \37797 , \37796 );
buf \U$37819 ( \37798 , \37797 );
not \U$37820 ( \37799 , \37798 );
or \U$37821 ( \37800 , \37782 , \37799 );
buf \U$37822 ( \37801 , \521 );
not \U$37823 ( \37802 , \37801 );
buf \U$37824 ( \37803 , \34011 );
not \U$37825 ( \37804 , \37803 );
and \U$37826 ( \37805 , \37802 , \37804 );
buf \U$37827 ( \37806 , \711 );
buf \U$37828 ( \37807 , \37646 );
nor \U$37829 ( \37808 , \37806 , \37807 );
buf \U$37830 ( \37809 , \37808 );
buf \U$37831 ( \37810 , \37809 );
nor \U$37832 ( \37811 , \37805 , \37810 );
buf \U$37833 ( \37812 , \37811 );
buf \U$37834 ( \37813 , \37812 );
not \U$37835 ( \37814 , \37813 );
buf \U$37836 ( \37815 , \37814 );
buf \U$37837 ( \37816 , \37815 );
nand \U$37838 ( \37817 , \37800 , \37816 );
buf \U$37839 ( \37818 , \37817 );
buf \U$37840 ( \37819 , \37818 );
buf \U$37841 ( \37820 , \37794 );
buf \U$37842 ( \37821 , \37780 );
not \U$37843 ( \37822 , \37821 );
buf \U$37844 ( \37823 , \37822 );
buf \U$37845 ( \37824 , \37823 );
nand \U$37846 ( \37825 , \37820 , \37824 );
buf \U$37847 ( \37826 , \37825 );
buf \U$37848 ( \37827 , \37826 );
nand \U$37849 ( \37828 , \37819 , \37827 );
buf \U$37850 ( \37829 , \37828 );
buf \U$37851 ( \37830 , \37829 );
and \U$37852 ( \37831 , \37770 , \37830 );
and \U$37853 ( \37832 , \37752 , \37769 );
or \U$37854 ( \37833 , \37831 , \37832 );
buf \U$37855 ( \37834 , \37833 );
buf \U$37856 ( \37835 , \37834 );
xor \U$37857 ( \37836 , \37738 , \37835 );
buf \U$37858 ( \37837 , \34315 );
not \U$37859 ( \37838 , \37837 );
buf \U$37860 ( \37839 , \13737 );
not \U$37861 ( \37840 , \37839 );
or \U$37862 ( \37841 , \37838 , \37840 );
buf \U$37863 ( \37842 , \1401 );
buf \U$37864 ( \37843 , \37685 );
nand \U$37865 ( \37844 , \37842 , \37843 );
buf \U$37866 ( \37845 , \37844 );
buf \U$37867 ( \37846 , \37845 );
nand \U$37868 ( \37847 , \37841 , \37846 );
buf \U$37869 ( \37848 , \37847 );
buf \U$37870 ( \37849 , \37848 );
not \U$37871 ( \37850 , \37849 );
buf \U$37872 ( \37851 , \34366 );
not \U$37873 ( \37852 , \37851 );
buf \U$37874 ( \37853 , \14940 );
not \U$37875 ( \37854 , \37853 );
or \U$37876 ( \37855 , \37852 , \37854 );
buf \U$37877 ( \37856 , \1025 );
buf \U$37878 ( \37857 , \36664 );
nand \U$37879 ( \37858 , \37856 , \37857 );
buf \U$37880 ( \37859 , \37858 );
buf \U$37881 ( \37860 , \37859 );
nand \U$37882 ( \37861 , \37855 , \37860 );
buf \U$37883 ( \37862 , \37861 );
buf \U$37884 ( \37863 , \37862 );
not \U$37885 ( \37864 , \37863 );
or \U$37886 ( \37865 , \37850 , \37864 );
buf \U$37887 ( \37866 , \37862 );
buf \U$37888 ( \37867 , \37848 );
or \U$37889 ( \37868 , \37866 , \37867 );
buf \U$37890 ( \37869 , \34117 );
not \U$37891 ( \37870 , \37869 );
buf \U$37892 ( \37871 , \4042 );
not \U$37893 ( \37872 , \37871 );
or \U$37894 ( \37873 , \37870 , \37872 );
buf \U$37895 ( \37874 , \4049 );
buf \U$37896 ( \37875 , \36808 );
nand \U$37897 ( \37876 , \37874 , \37875 );
buf \U$37898 ( \37877 , \37876 );
buf \U$37899 ( \37878 , \37877 );
nand \U$37900 ( \37879 , \37873 , \37878 );
buf \U$37901 ( \37880 , \37879 );
buf \U$37902 ( \37881 , \37880 );
nand \U$37903 ( \37882 , \37868 , \37881 );
buf \U$37904 ( \37883 , \37882 );
buf \U$37905 ( \37884 , \37883 );
nand \U$37906 ( \37885 , \37865 , \37884 );
buf \U$37907 ( \37886 , \37885 );
buf \U$37908 ( \37887 , \37886 );
buf \U$37909 ( \37888 , \33931 );
not \U$37910 ( \37889 , \37888 );
buf \U$37911 ( \37890 , \2269 );
not \U$37912 ( \37891 , \37890 );
or \U$37913 ( \37892 , \37889 , \37891 );
buf \U$37914 ( \37893 , \1282 );
buf \U$37915 ( \37894 , \37423 );
nand \U$37916 ( \37895 , \37893 , \37894 );
buf \U$37917 ( \37896 , \37895 );
buf \U$37918 ( \37897 , \37896 );
nand \U$37919 ( \37898 , \37892 , \37897 );
buf \U$37920 ( \37899 , \37898 );
buf \U$37921 ( \37900 , \37899 );
not \U$37922 ( \37901 , \37900 );
buf \U$37923 ( \37902 , \34295 );
not \U$37924 ( \37903 , \37902 );
buf \U$37925 ( \37904 , \14346 );
not \U$37926 ( \37905 , \37904 );
or \U$37927 ( \37906 , \37903 , \37905 );
buf \U$37928 ( \37907 , \14352 );
buf \U$37929 ( \37908 , RIc0daa08_111);
nand \U$37930 ( \37909 , \37907 , \37908 );
buf \U$37931 ( \37910 , \37909 );
buf \U$37932 ( \37911 , \37910 );
nand \U$37933 ( \37912 , \37906 , \37911 );
buf \U$37934 ( \37913 , \37912 );
buf \U$37935 ( \37914 , \37913 );
not \U$37936 ( \37915 , \37914 );
or \U$37937 ( \37916 , \37901 , \37915 );
buf \U$37938 ( \37917 , \37899 );
not \U$37939 ( \37918 , \37917 );
buf \U$37940 ( \37919 , \37918 );
buf \U$37941 ( \37920 , \37919 );
not \U$37942 ( \37921 , \37920 );
buf \U$37943 ( \37922 , \37913 );
not \U$37944 ( \37923 , \37922 );
buf \U$37945 ( \37924 , \37923 );
buf \U$37946 ( \37925 , \37924 );
not \U$37947 ( \37926 , \37925 );
or \U$37948 ( \37927 , \37921 , \37926 );
buf \U$37949 ( \37928 , \34282 );
not \U$37950 ( \37929 , \37928 );
buf \U$37951 ( \37930 , \14419 );
not \U$37952 ( \37931 , \37930 );
or \U$37953 ( \37932 , \37929 , \37931 );
buf \U$37954 ( \37933 , \12584 );
buf \U$37955 ( \37934 , \37668 );
nand \U$37956 ( \37935 , \37933 , \37934 );
buf \U$37957 ( \37936 , \37935 );
buf \U$37958 ( \37937 , \37936 );
nand \U$37959 ( \37938 , \37932 , \37937 );
buf \U$37960 ( \37939 , \37938 );
buf \U$37961 ( \37940 , \37939 );
nand \U$37962 ( \37941 , \37927 , \37940 );
buf \U$37963 ( \37942 , \37941 );
buf \U$37964 ( \37943 , \37942 );
nand \U$37965 ( \37944 , \37916 , \37943 );
buf \U$37966 ( \37945 , \37944 );
buf \U$37967 ( \37946 , \37945 );
xor \U$37968 ( \37947 , \37887 , \37946 );
buf \U$37969 ( \37948 , \33959 );
not \U$37970 ( \37949 , \37948 );
buf \U$37971 ( \37950 , \3780 );
not \U$37972 ( \37951 , \37950 );
or \U$37973 ( \37952 , \37949 , \37951 );
buf \U$37974 ( \37953 , \4427 );
buf \U$37975 ( \37954 , \37439 );
nand \U$37976 ( \37955 , \37953 , \37954 );
buf \U$37977 ( \37956 , \37955 );
buf \U$37978 ( \37957 , \37956 );
nand \U$37979 ( \37958 , \37952 , \37957 );
buf \U$37980 ( \37959 , \37958 );
buf \U$37981 ( \37960 , \37959 );
not \U$37982 ( \37961 , \37960 );
buf \U$37983 ( \37962 , \37961 );
buf \U$37984 ( \37963 , \37962 );
not \U$37985 ( \37964 , \37963 );
buf \U$37986 ( \37965 , \34409 );
not \U$37987 ( \37966 , \37965 );
buf \U$37988 ( \37967 , \18220 );
not \U$37989 ( \37968 , \37967 );
or \U$37990 ( \37969 , \37966 , \37968 );
buf \U$37991 ( \37970 , \18416 );
buf \U$37992 ( \37971 , \36758 );
nand \U$37993 ( \37972 , \37970 , \37971 );
buf \U$37994 ( \37973 , \37972 );
buf \U$37995 ( \37974 , \37973 );
nand \U$37996 ( \37975 , \37969 , \37974 );
buf \U$37997 ( \37976 , \37975 );
buf \U$37998 ( \37977 , \37976 );
not \U$37999 ( \37978 , \37977 );
buf \U$38000 ( \37979 , \37978 );
buf \U$38001 ( \37980 , \37979 );
not \U$38002 ( \37981 , \37980 );
or \U$38003 ( \37982 , \37964 , \37981 );
buf \U$38004 ( \37983 , \34349 );
not \U$38005 ( \37984 , \37983 );
buf \U$38006 ( \37985 , \13569 );
not \U$38007 ( \37986 , \37985 );
or \U$38008 ( \37987 , \37984 , \37986 );
buf \U$38009 ( \37988 , \481 );
buf \U$38010 ( \37989 , \36678 );
nand \U$38011 ( \37990 , \37988 , \37989 );
buf \U$38012 ( \37991 , \37990 );
buf \U$38013 ( \37992 , \37991 );
nand \U$38014 ( \37993 , \37987 , \37992 );
buf \U$38015 ( \37994 , \37993 );
buf \U$38016 ( \37995 , \37994 );
nand \U$38017 ( \37996 , \37982 , \37995 );
buf \U$38018 ( \37997 , \37996 );
buf \U$38019 ( \37998 , \37997 );
buf \U$38020 ( \37999 , \37976 );
buf \U$38021 ( \38000 , \37959 );
nand \U$38022 ( \38001 , \37999 , \38000 );
buf \U$38023 ( \38002 , \38001 );
buf \U$38024 ( \38003 , \38002 );
nand \U$38025 ( \38004 , \37998 , \38003 );
buf \U$38026 ( \38005 , \38004 );
buf \U$38027 ( \38006 , \38005 );
and \U$38028 ( \38007 , \37947 , \38006 );
and \U$38029 ( \38008 , \37887 , \37946 );
or \U$38030 ( \38009 , \38007 , \38008 );
buf \U$38031 ( \38010 , \38009 );
buf \U$38032 ( \38011 , \38010 );
and \U$38033 ( \38012 , \37836 , \38011 );
and \U$38034 ( \38013 , \37738 , \37835 );
or \U$38035 ( \38014 , \38012 , \38013 );
buf \U$38036 ( \38015 , \38014 );
buf \U$38037 ( \38016 , \38015 );
xor \U$38038 ( \38017 , \36649 , \36659 );
xor \U$38039 ( \38018 , \38017 , \36854 );
buf \U$38040 ( \38019 , \38018 );
buf \U$38041 ( \38020 , \38019 );
xor \U$38042 ( \38021 , \38016 , \38020 );
buf \U$38043 ( \38022 , \34189 );
not \U$38044 ( \38023 , \38022 );
buf \U$38045 ( \38024 , \1736 );
not \U$38046 ( \38025 , \38024 );
or \U$38047 ( \38026 , \38023 , \38025 );
buf \U$38048 ( \38027 , \584 );
buf \U$38049 ( \38028 , \37497 );
nand \U$38050 ( \38029 , \38027 , \38028 );
buf \U$38051 ( \38030 , \38029 );
buf \U$38052 ( \38031 , \38030 );
nand \U$38053 ( \38032 , \38026 , \38031 );
buf \U$38054 ( \38033 , \38032 );
not \U$38055 ( \38034 , \38033 );
not \U$38056 ( \38035 , \5368 );
not \U$38057 ( \38036 , \36827 );
and \U$38058 ( \38037 , \38035 , \38036 );
not \U$38059 ( \38038 , \3384 );
nor \U$38060 ( \38039 , \38038 , \34042 );
nor \U$38061 ( \38040 , \38037 , \38039 );
buf \U$38062 ( \38041 , \38040 );
not \U$38063 ( \38042 , \38041 );
buf \U$38064 ( \38043 , \38042 );
not \U$38065 ( \38044 , \38043 );
or \U$38066 ( \38045 , \38034 , \38044 );
not \U$38067 ( \38046 , \38040 );
buf \U$38068 ( \38047 , \38033 );
not \U$38069 ( \38048 , \38047 );
buf \U$38070 ( \38049 , \38048 );
not \U$38071 ( \38050 , \38049 );
or \U$38072 ( \38051 , \38046 , \38050 );
buf \U$38073 ( \38052 , \33942 );
not \U$38074 ( \38053 , \38052 );
buf \U$38075 ( \38054 , \26572 );
not \U$38076 ( \38055 , \38054 );
or \U$38077 ( \38056 , \38053 , \38055 );
buf \U$38078 ( \38057 , \2070 );
buf \U$38079 ( \38058 , \37469 );
nand \U$38080 ( \38059 , \38057 , \38058 );
buf \U$38081 ( \38060 , \38059 );
buf \U$38082 ( \38061 , \38060 );
nand \U$38083 ( \38062 , \38056 , \38061 );
buf \U$38084 ( \38063 , \38062 );
nand \U$38085 ( \38064 , \38051 , \38063 );
nand \U$38086 ( \38065 , \38045 , \38064 );
buf \U$38087 ( \38066 , \38065 );
not \U$38088 ( \38067 , \38066 );
buf \U$38089 ( \38068 , \38067 );
buf \U$38090 ( \38069 , \38068 );
not \U$38091 ( \38070 , \38069 );
buf \U$38092 ( \38071 , \34172 );
not \U$38093 ( \38072 , \38071 );
buf \U$38094 ( \38073 , \4691 );
not \U$38095 ( \38074 , \38073 );
or \U$38096 ( \38075 , \38072 , \38074 );
buf \U$38097 ( \38076 , \284 );
buf \U$38098 ( \38077 , \37514 );
nand \U$38099 ( \38078 , \38076 , \38077 );
buf \U$38100 ( \38079 , \38078 );
buf \U$38101 ( \38080 , \38079 );
nand \U$38102 ( \38081 , \38075 , \38080 );
buf \U$38103 ( \38082 , \38081 );
buf \U$38104 ( \38083 , \34029 );
not \U$38105 ( \38084 , \38083 );
buf \U$38106 ( \38085 , \17141 );
not \U$38107 ( \38086 , \38085 );
or \U$38108 ( \38087 , \38084 , \38086 );
buf \U$38109 ( \38088 , \1078 );
buf \U$38110 ( \38089 , \36723 );
nand \U$38111 ( \38090 , \38088 , \38089 );
buf \U$38112 ( \38091 , \38090 );
buf \U$38113 ( \38092 , \38091 );
nand \U$38114 ( \38093 , \38087 , \38092 );
buf \U$38115 ( \38094 , \38093 );
xor \U$38116 ( \38095 , \38082 , \38094 );
buf \U$38117 ( \38096 , \34264 );
not \U$38118 ( \38097 , \38096 );
buf \U$38119 ( \38098 , \1431 );
not \U$38120 ( \38099 , \38098 );
or \U$38121 ( \38100 , \38097 , \38099 );
buf \U$38122 ( \38101 , \1588 );
buf \U$38123 ( \38102 , \37396 );
nand \U$38124 ( \38103 , \38101 , \38102 );
buf \U$38125 ( \38104 , \38103 );
buf \U$38126 ( \38105 , \38104 );
nand \U$38127 ( \38106 , \38100 , \38105 );
buf \U$38128 ( \38107 , \38106 );
and \U$38129 ( \38108 , \38095 , \38107 );
and \U$38130 ( \38109 , \38082 , \38094 );
or \U$38131 ( \38110 , \38108 , \38109 );
buf \U$38132 ( \38111 , \38110 );
not \U$38133 ( \38112 , \38111 );
buf \U$38134 ( \38113 , \38112 );
buf \U$38135 ( \38114 , \38113 );
not \U$38136 ( \38115 , \38114 );
or \U$38137 ( \38116 , \38070 , \38115 );
buf \U$38138 ( \38117 , \34210 );
not \U$38139 ( \38118 , \38117 );
buf \U$38140 ( \38119 , \20741 );
not \U$38141 ( \38120 , \38119 );
or \U$38142 ( \38121 , \38118 , \38120 );
buf \U$38143 ( \38122 , \12342 );
buf \U$38144 ( \38123 , \37529 );
nand \U$38145 ( \38124 , \38122 , \38123 );
buf \U$38146 ( \38125 , \38124 );
buf \U$38147 ( \38126 , \38125 );
nand \U$38148 ( \38127 , \38121 , \38126 );
buf \U$38149 ( \38128 , \38127 );
not \U$38150 ( \38129 , \38128 );
buf \U$38151 ( \38130 , \1124 );
not \U$38152 ( \38131 , \38130 );
buf \U$38153 ( \38132 , \34234 );
not \U$38154 ( \38133 , \38132 );
buf \U$38155 ( \38134 , \38133 );
buf \U$38156 ( \38135 , \38134 );
not \U$38157 ( \38136 , \38135 );
and \U$38158 ( \38137 , \38131 , \38136 );
buf \U$38159 ( \38138 , \37356 );
not \U$38160 ( \38139 , \38138 );
buf \U$38161 ( \38140 , \2372 );
nor \U$38162 ( \38141 , \38139 , \38140 );
buf \U$38163 ( \38142 , \38141 );
buf \U$38164 ( \38143 , \38142 );
nor \U$38165 ( \38144 , \38137 , \38143 );
buf \U$38166 ( \38145 , \38144 );
buf \U$38167 ( \38146 , \38145 );
not \U$38168 ( \38147 , \38146 );
buf \U$38169 ( \38148 , \38147 );
not \U$38170 ( \38149 , \38148 );
or \U$38171 ( \38150 , \38129 , \38149 );
not \U$38172 ( \38151 , \38145 );
buf \U$38173 ( \38152 , \38128 );
not \U$38174 ( \38153 , \38152 );
buf \U$38175 ( \38154 , \38153 );
not \U$38176 ( \38155 , \38154 );
or \U$38177 ( \38156 , \38151 , \38155 );
buf \U$38178 ( \38157 , \34427 );
not \U$38179 ( \38158 , \38157 );
buf \U$38180 ( \38159 , \12736 );
not \U$38181 ( \38160 , \38159 );
or \U$38182 ( \38161 , \38158 , \38160 );
buf \U$38183 ( \38162 , \12744 );
buf \U$38184 ( \38163 , \37756 );
nand \U$38185 ( \38164 , \38162 , \38163 );
buf \U$38186 ( \38165 , \38164 );
buf \U$38187 ( \38166 , \38165 );
nand \U$38188 ( \38167 , \38161 , \38166 );
buf \U$38189 ( \38168 , \38167 );
nand \U$38190 ( \38169 , \38156 , \38168 );
nand \U$38191 ( \38170 , \38150 , \38169 );
buf \U$38192 ( \38171 , \38170 );
nand \U$38193 ( \38172 , \38116 , \38171 );
buf \U$38194 ( \38173 , \38172 );
buf \U$38195 ( \38174 , \38173 );
buf \U$38196 ( \38175 , \38110 );
buf \U$38197 ( \38176 , \38065 );
nand \U$38198 ( \38177 , \38175 , \38176 );
buf \U$38199 ( \38178 , \38177 );
buf \U$38200 ( \38179 , \38178 );
nand \U$38201 ( \38180 , \38174 , \38179 );
buf \U$38202 ( \38181 , \38180 );
buf \U$38203 ( \38182 , \38181 );
xor \U$38204 ( \38183 , \37386 , \37368 );
xnor \U$38205 ( \38184 , \38183 , \37408 );
buf \U$38206 ( \38185 , \38184 );
xor \U$38207 ( \38186 , \37627 , \37641 );
xor \U$38208 ( \38187 , \38186 , \37662 );
buf \U$38209 ( \38188 , \38187 );
buf \U$38210 ( \38189 , \38188 );
not \U$38211 ( \38190 , \38189 );
buf \U$38212 ( \38191 , \38190 );
buf \U$38213 ( \38192 , \38191 );
nand \U$38214 ( \38193 , \38185 , \38192 );
buf \U$38215 ( \38194 , \38193 );
not \U$38216 ( \38195 , \38194 );
xor \U$38217 ( \38196 , \36807 , \36822 );
xor \U$38218 ( \38197 , \38196 , \36843 );
buf \U$38219 ( \38198 , \38197 );
not \U$38220 ( \38199 , \38198 );
or \U$38221 ( \38200 , \38195 , \38199 );
buf \U$38222 ( \38201 , \38191 );
not \U$38223 ( \38202 , \38201 );
buf \U$38224 ( \38203 , \38184 );
not \U$38225 ( \38204 , \38203 );
buf \U$38226 ( \38205 , \38204 );
buf \U$38227 ( \38206 , \38205 );
nand \U$38228 ( \38207 , \38202 , \38206 );
buf \U$38229 ( \38208 , \38207 );
nand \U$38230 ( \38209 , \38200 , \38208 );
buf \U$38231 ( \38210 , \38209 );
xor \U$38232 ( \38211 , \38182 , \38210 );
xor \U$38233 ( \38212 , \37667 , \37716 );
xor \U$38234 ( \38213 , \38212 , \37721 );
buf \U$38235 ( \38214 , \38213 );
buf \U$38236 ( \38215 , \38214 );
and \U$38237 ( \38216 , \38211 , \38215 );
and \U$38238 ( \38217 , \38182 , \38210 );
or \U$38239 ( \38218 , \38216 , \38217 );
buf \U$38240 ( \38219 , \38218 );
buf \U$38241 ( \38220 , \38219 );
xor \U$38242 ( \38221 , \38021 , \38220 );
buf \U$38243 ( \38222 , \38221 );
buf \U$38244 ( \38223 , \38222 );
and \U$38245 ( \38224 , \37734 , \38223 );
and \U$38246 ( \38225 , \37729 , \37733 );
or \U$38247 ( \38226 , \38224 , \38225 );
buf \U$38248 ( \38227 , \38226 );
buf \U$38249 ( \38228 , \38227 );
not \U$38250 ( \38229 , \38228 );
and \U$38251 ( \38230 , \37352 , \38229 );
buf \U$38252 ( \38231 , \38227 );
buf \U$38253 ( \38232 , \37350 );
and \U$38254 ( \38233 , \38231 , \38232 );
nor \U$38255 ( \38234 , \38230 , \38233 );
buf \U$38256 ( \38235 , \38234 );
buf \U$38257 ( \38236 , \38235 );
not \U$38258 ( \38237 , \38236 );
xor \U$38259 ( \38238 , \37738 , \37835 );
xor \U$38260 ( \38239 , \38238 , \38011 );
buf \U$38261 ( \38240 , \38239 );
buf \U$38262 ( \38241 , \38240 );
xor \U$38263 ( \38242 , \37752 , \37769 );
xor \U$38264 ( \38243 , \38242 , \37830 );
buf \U$38265 ( \38244 , \38243 );
buf \U$38266 ( \38245 , \38244 );
buf \U$38267 ( \38246 , \37751 );
not \U$38268 ( \38247 , \38246 );
buf \U$38269 ( \38248 , \38247 );
buf \U$38270 ( \38249 , \38248 );
buf \U$38271 ( \38250 , \33935 );
not \U$38272 ( \38251 , \38250 );
buf \U$38273 ( \38252 , \33968 );
not \U$38274 ( \38253 , \38252 );
or \U$38275 ( \38254 , \38251 , \38253 );
buf \U$38276 ( \38255 , \33948 );
nand \U$38277 ( \38256 , \38254 , \38255 );
buf \U$38278 ( \38257 , \38256 );
buf \U$38279 ( \38258 , \38257 );
buf \U$38280 ( \38259 , \33935 );
not \U$38281 ( \38260 , \38259 );
buf \U$38282 ( \38261 , \33965 );
nand \U$38283 ( \38262 , \38260 , \38261 );
buf \U$38284 ( \38263 , \38262 );
buf \U$38285 ( \38264 , \38263 );
nand \U$38286 ( \38265 , \38258 , \38264 );
buf \U$38287 ( \38266 , \38265 );
buf \U$38288 ( \38267 , \38266 );
xor \U$38289 ( \38268 , \38249 , \38267 );
xor \U$38290 ( \38269 , \34179 , \34196 );
and \U$38291 ( \38270 , \38269 , \34217 );
and \U$38292 ( \38271 , \34179 , \34196 );
or \U$38293 ( \38272 , \38270 , \38271 );
buf \U$38294 ( \38273 , \38272 );
buf \U$38295 ( \38274 , \38273 );
and \U$38296 ( \38275 , \38268 , \38274 );
and \U$38297 ( \38276 , \38249 , \38267 );
or \U$38298 ( \38277 , \38275 , \38276 );
buf \U$38299 ( \38278 , \38277 );
buf \U$38300 ( \38279 , \38278 );
xor \U$38301 ( \38280 , \38245 , \38279 );
xor \U$38302 ( \38281 , \34089 , \34106 );
and \U$38303 ( \38282 , \38281 , \34124 );
and \U$38304 ( \38283 , \34089 , \34106 );
or \U$38305 ( \38284 , \38282 , \38283 );
buf \U$38306 ( \38285 , \38284 );
buf \U$38307 ( \38286 , \38285 );
xor \U$38308 ( \38287 , \34036 , \34051 );
and \U$38309 ( \38288 , \38287 , \34069 );
and \U$38310 ( \38289 , \34036 , \34051 );
or \U$38311 ( \38290 , \38288 , \38289 );
buf \U$38312 ( \38291 , \38290 );
buf \U$38313 ( \38292 , \38291 );
xor \U$38314 ( \38293 , \38286 , \38292 );
xor \U$38315 ( \38294 , \34356 , \34373 );
and \U$38316 ( \38295 , \38294 , \34395 );
and \U$38317 ( \38296 , \34356 , \34373 );
or \U$38318 ( \38297 , \38295 , \38296 );
buf \U$38319 ( \38298 , \38297 );
buf \U$38320 ( \38299 , \38298 );
and \U$38321 ( \38300 , \38293 , \38299 );
and \U$38322 ( \38301 , \38286 , \38292 );
or \U$38323 ( \38302 , \38300 , \38301 );
buf \U$38324 ( \38303 , \38302 );
buf \U$38325 ( \38304 , \38303 );
and \U$38326 ( \38305 , \38280 , \38304 );
and \U$38327 ( \38306 , \38245 , \38279 );
or \U$38328 ( \38307 , \38305 , \38306 );
buf \U$38329 ( \38308 , \38307 );
buf \U$38330 ( \38309 , \38308 );
xor \U$38331 ( \38310 , \38241 , \38309 );
xor \U$38332 ( \38311 , \34241 , \34253 );
and \U$38333 ( \38312 , \38311 , \34271 );
and \U$38334 ( \38313 , \34241 , \34253 );
or \U$38335 ( \38314 , \38312 , \38313 );
buf \U$38336 ( \38315 , \38314 );
buf \U$38337 ( \38316 , \38315 );
xor \U$38338 ( \38317 , \33983 , \34001 );
and \U$38339 ( \38318 , \38317 , \34020 );
and \U$38340 ( \38319 , \33983 , \34001 );
or \U$38341 ( \38320 , \38318 , \38319 );
buf \U$38342 ( \38321 , \38320 );
buf \U$38343 ( \38322 , \38321 );
xor \U$38344 ( \38323 , \38316 , \38322 );
buf \U$38345 ( \38324 , \34324 );
not \U$38346 ( \38325 , \38324 );
buf \U$38347 ( \38326 , \34288 );
not \U$38348 ( \38327 , \38326 );
buf \U$38349 ( \38328 , \38327 );
buf \U$38350 ( \38329 , \38328 );
not \U$38351 ( \38330 , \38329 );
or \U$38352 ( \38331 , \38325 , \38330 );
buf \U$38353 ( \38332 , \34301 );
nand \U$38354 ( \38333 , \38331 , \38332 );
buf \U$38355 ( \38334 , \38333 );
buf \U$38356 ( \38335 , \38334 );
buf \U$38357 ( \38336 , \34288 );
buf \U$38358 ( \38337 , \34321 );
nand \U$38359 ( \38338 , \38336 , \38337 );
buf \U$38360 ( \38339 , \38338 );
buf \U$38361 ( \38340 , \38339 );
nand \U$38362 ( \38341 , \38335 , \38340 );
buf \U$38363 ( \38342 , \38341 );
buf \U$38364 ( \38343 , \38342 );
and \U$38365 ( \38344 , \38323 , \38343 );
and \U$38366 ( \38345 , \38316 , \38322 );
or \U$38367 ( \38346 , \38344 , \38345 );
buf \U$38368 ( \38347 , \38346 );
buf \U$38369 ( \38348 , \38347 );
xor \U$38370 ( \38349 , \37880 , \37862 );
xor \U$38371 ( \38350 , \38349 , \37848 );
buf \U$38372 ( \38351 , \38350 );
buf \U$38373 ( \38352 , \37794 );
not \U$38374 ( \38353 , \38352 );
buf \U$38375 ( \38354 , \37812 );
not \U$38376 ( \38355 , \38354 );
and \U$38377 ( \38356 , \38353 , \38355 );
buf \U$38378 ( \38357 , \37794 );
buf \U$38379 ( \38358 , \37812 );
and \U$38380 ( \38359 , \38357 , \38358 );
nor \U$38381 ( \38360 , \38356 , \38359 );
buf \U$38382 ( \38361 , \38360 );
buf \U$38383 ( \38362 , \38361 );
buf \U$38384 ( \38363 , \37780 );
and \U$38385 ( \38364 , \38362 , \38363 );
not \U$38386 ( \38365 , \38362 );
buf \U$38387 ( \38366 , \37823 );
and \U$38388 ( \38367 , \38365 , \38366 );
nor \U$38389 ( \38368 , \38364 , \38367 );
buf \U$38390 ( \38369 , \38368 );
buf \U$38391 ( \38370 , \38369 );
xor \U$38392 ( \38371 , \38351 , \38370 );
buf \U$38393 ( \38372 , RIc0d8c80_48);
buf \U$38394 ( \38373 , RIc0d9478_65);
nand \U$38395 ( \38374 , \38372 , \38373 );
buf \U$38396 ( \38375 , \38374 );
buf \U$38397 ( \38376 , \38375 );
buf \U$38398 ( \38377 , \34388 );
not \U$38399 ( \38378 , \38377 );
buf \U$38400 ( \38379 , \27660 );
not \U$38401 ( \38380 , \38379 );
or \U$38402 ( \38381 , \38378 , \38380 );
buf \U$38403 ( \38382 , \20211 );
buf \U$38404 ( \38383 , \36696 );
nand \U$38405 ( \38384 , \38382 , \38383 );
buf \U$38406 ( \38385 , \38384 );
buf \U$38407 ( \38386 , \38385 );
nand \U$38408 ( \38387 , \38381 , \38386 );
buf \U$38409 ( \38388 , \38387 );
buf \U$38410 ( \38389 , \38388 );
xor \U$38411 ( \38390 , \38376 , \38389 );
buf \U$38412 ( \38391 , \34062 );
not \U$38413 ( \38392 , \38391 );
buf \U$38414 ( \38393 , \330 );
not \U$38415 ( \38394 , \38393 );
or \U$38416 ( \38395 , \38392 , \38394 );
buf \U$38417 ( \38396 , \344 );
buf \U$38418 ( \38397 , \36739 );
nand \U$38419 ( \38398 , \38396 , \38397 );
buf \U$38420 ( \38399 , \38398 );
buf \U$38421 ( \38400 , \38399 );
nand \U$38422 ( \38401 , \38395 , \38400 );
buf \U$38423 ( \38402 , \38401 );
buf \U$38424 ( \38403 , \38402 );
xnor \U$38425 ( \38404 , \38390 , \38403 );
buf \U$38426 ( \38405 , \38404 );
buf \U$38427 ( \38406 , \38405 );
and \U$38428 ( \38407 , \38371 , \38406 );
and \U$38429 ( \38408 , \38351 , \38370 );
or \U$38430 ( \38409 , \38407 , \38408 );
buf \U$38431 ( \38410 , \38409 );
buf \U$38432 ( \38411 , \38410 );
xor \U$38433 ( \38412 , \38348 , \38411 );
xor \U$38434 ( \38413 , \38049 , \38063 );
xnor \U$38435 ( \38414 , \38413 , \38043 );
buf \U$38436 ( \38415 , \38414 );
xor \U$38437 ( \38416 , \38082 , \38094 );
xor \U$38438 ( \38417 , \38416 , \38107 );
buf \U$38439 ( \38418 , \38417 );
or \U$38440 ( \38419 , \38415 , \38418 );
and \U$38441 ( \38420 , \37994 , \37979 );
not \U$38442 ( \38421 , \37994 );
and \U$38443 ( \38422 , \38421 , \37976 );
or \U$38444 ( \38423 , \38420 , \38422 );
and \U$38445 ( \38424 , \38423 , \37962 );
not \U$38446 ( \38425 , \38423 );
and \U$38447 ( \38426 , \38425 , \37959 );
nor \U$38448 ( \38427 , \38424 , \38426 );
buf \U$38449 ( \38428 , \38427 );
not \U$38450 ( \38429 , \38428 );
buf \U$38451 ( \38430 , \38429 );
buf \U$38452 ( \38431 , \38430 );
nand \U$38453 ( \38432 , \38419 , \38431 );
buf \U$38454 ( \38433 , \38432 );
buf \U$38455 ( \38434 , \38433 );
buf \U$38456 ( \38435 , \38414 );
buf \U$38457 ( \38436 , \38417 );
nand \U$38458 ( \38437 , \38435 , \38436 );
buf \U$38459 ( \38438 , \38437 );
buf \U$38460 ( \38439 , \38438 );
nand \U$38461 ( \38440 , \38434 , \38439 );
buf \U$38462 ( \38441 , \38440 );
buf \U$38463 ( \38442 , \38441 );
and \U$38464 ( \38443 , \38412 , \38442 );
and \U$38465 ( \38444 , \38348 , \38411 );
or \U$38466 ( \38445 , \38443 , \38444 );
buf \U$38467 ( \38446 , \38445 );
buf \U$38468 ( \38447 , \38446 );
and \U$38469 ( \38448 , \38310 , \38447 );
and \U$38470 ( \38449 , \38241 , \38309 );
or \U$38471 ( \38450 , \38448 , \38449 );
buf \U$38472 ( \38451 , \38450 );
buf \U$38473 ( \38452 , \38451 );
xor \U$38474 ( \38453 , \37887 , \37946 );
xor \U$38475 ( \38454 , \38453 , \38006 );
buf \U$38476 ( \38455 , \38454 );
not \U$38477 ( \38456 , \38455 );
buf \U$38478 ( \38457 , \38170 );
not \U$38479 ( \38458 , \38457 );
buf \U$38480 ( \38459 , \38113 );
not \U$38481 ( \38460 , \38459 );
or \U$38482 ( \38461 , \38458 , \38460 );
buf \U$38483 ( \38462 , \38113 );
buf \U$38484 ( \38463 , \38170 );
or \U$38485 ( \38464 , \38462 , \38463 );
nand \U$38486 ( \38465 , \38461 , \38464 );
buf \U$38487 ( \38466 , \38465 );
buf \U$38488 ( \38467 , \38466 );
buf \U$38489 ( \38468 , \38065 );
xnor \U$38490 ( \38469 , \38467 , \38468 );
buf \U$38491 ( \38470 , \38469 );
nand \U$38492 ( \38471 , \38456 , \38470 );
not \U$38493 ( \38472 , \38471 );
xor \U$38494 ( \38473 , \36770 , \36751 );
xor \U$38495 ( \38474 , \38473 , \36736 );
buf \U$38496 ( \38475 , \38402 );
buf \U$38497 ( \38476 , \38375 );
not \U$38498 ( \38477 , \38476 );
buf \U$38499 ( \38478 , \38477 );
buf \U$38500 ( \38479 , \38478 );
or \U$38501 ( \38480 , \38475 , \38479 );
buf \U$38502 ( \38481 , \38388 );
nand \U$38503 ( \38482 , \38480 , \38481 );
buf \U$38504 ( \38483 , \38482 );
buf \U$38505 ( \38484 , \38483 );
buf \U$38506 ( \38485 , \38402 );
buf \U$38507 ( \38486 , \38478 );
nand \U$38508 ( \38487 , \38485 , \38486 );
buf \U$38509 ( \38488 , \38487 );
buf \U$38510 ( \38489 , \38488 );
nand \U$38511 ( \38490 , \38484 , \38489 );
buf \U$38512 ( \38491 , \38490 );
buf \U$38513 ( \38492 , \38491 );
not \U$38514 ( \38493 , \38492 );
buf \U$38515 ( \38494 , \37462 );
not \U$38516 ( \38495 , \38494 );
buf \U$38517 ( \38496 , \37481 );
not \U$38518 ( \38497 , \38496 );
or \U$38519 ( \38498 , \38495 , \38497 );
buf \U$38520 ( \38499 , \37481 );
buf \U$38521 ( \38500 , \37462 );
or \U$38522 ( \38501 , \38499 , \38500 );
nand \U$38523 ( \38502 , \38498 , \38501 );
buf \U$38524 ( \38503 , \38502 );
buf \U$38525 ( \38504 , \38503 );
buf \U$38526 ( \38505 , \37457 );
and \U$38527 ( \38506 , \38504 , \38505 );
not \U$38528 ( \38507 , \38504 );
buf \U$38529 ( \38508 , \37435 );
and \U$38530 ( \38509 , \38507 , \38508 );
nor \U$38531 ( \38510 , \38506 , \38509 );
buf \U$38532 ( \38511 , \38510 );
buf \U$38533 ( \38512 , \38511 );
not \U$38534 ( \38513 , \38512 );
or \U$38535 ( \38514 , \38493 , \38513 );
buf \U$38536 ( \38515 , \38511 );
buf \U$38537 ( \38516 , \38491 );
or \U$38538 ( \38517 , \38515 , \38516 );
nand \U$38539 ( \38518 , \38514 , \38517 );
buf \U$38540 ( \38519 , \38518 );
xor \U$38541 ( \38520 , \38474 , \38519 );
not \U$38542 ( \38521 , \38520 );
or \U$38543 ( \38522 , \38472 , \38521 );
buf \U$38544 ( \38523 , \38470 );
not \U$38545 ( \38524 , \38523 );
buf \U$38546 ( \38525 , \38455 );
nand \U$38547 ( \38526 , \38524 , \38525 );
buf \U$38548 ( \38527 , \38526 );
nand \U$38549 ( \38528 , \38522 , \38527 );
buf \U$38550 ( \38529 , \38528 );
xor \U$38551 ( \38530 , \37939 , \37924 );
xnor \U$38552 ( \38531 , \38530 , \37919 );
buf \U$38553 ( \38532 , \38531 );
not \U$38554 ( \38533 , \38532 );
buf \U$38555 ( \38534 , \38533 );
buf \U$38556 ( \38535 , \38534 );
not \U$38557 ( \38536 , \38535 );
buf \U$38558 ( \38537 , \34433 );
not \U$38559 ( \38538 , \38537 );
buf \U$38560 ( \38539 , \34451 );
not \U$38561 ( \38540 , \38539 );
or \U$38562 ( \38541 , \38538 , \38540 );
buf \U$38563 ( \38542 , \34436 );
not \U$38564 ( \38543 , \38542 );
buf \U$38565 ( \38544 , \32838 );
not \U$38566 ( \38545 , \38544 );
or \U$38567 ( \38546 , \38543 , \38545 );
buf \U$38568 ( \38547 , \34415 );
nand \U$38569 ( \38548 , \38546 , \38547 );
buf \U$38570 ( \38549 , \38548 );
buf \U$38571 ( \38550 , \38549 );
nand \U$38572 ( \38551 , \38541 , \38550 );
buf \U$38573 ( \38552 , \38551 );
buf \U$38574 ( \38553 , \38552 );
not \U$38575 ( \38554 , \38553 );
or \U$38576 ( \38555 , \38536 , \38554 );
buf \U$38577 ( \38556 , \38531 );
not \U$38578 ( \38557 , \38556 );
buf \U$38579 ( \38558 , \38552 );
not \U$38580 ( \38559 , \38558 );
buf \U$38581 ( \38560 , \38559 );
buf \U$38582 ( \38561 , \38560 );
not \U$38583 ( \38562 , \38561 );
or \U$38584 ( \38563 , \38557 , \38562 );
buf \U$38585 ( \38564 , \38168 );
not \U$38586 ( \38565 , \38564 );
buf \U$38587 ( \38566 , \38154 );
not \U$38588 ( \38567 , \38566 );
or \U$38589 ( \38568 , \38565 , \38567 );
buf \U$38590 ( \38569 , \38154 );
buf \U$38591 ( \38570 , \38168 );
or \U$38592 ( \38571 , \38569 , \38570 );
nand \U$38593 ( \38572 , \38568 , \38571 );
buf \U$38594 ( \38573 , \38572 );
buf \U$38595 ( \38574 , \38573 );
buf \U$38596 ( \38575 , \38148 );
and \U$38597 ( \38576 , \38574 , \38575 );
not \U$38598 ( \38577 , \38574 );
buf \U$38599 ( \38578 , \38145 );
and \U$38600 ( \38579 , \38577 , \38578 );
nor \U$38601 ( \38580 , \38576 , \38579 );
buf \U$38602 ( \38581 , \38580 );
buf \U$38603 ( \38582 , \38581 );
nand \U$38604 ( \38583 , \38563 , \38582 );
buf \U$38605 ( \38584 , \38583 );
buf \U$38606 ( \38585 , \38584 );
nand \U$38607 ( \38586 , \38555 , \38585 );
buf \U$38608 ( \38587 , \38586 );
buf \U$38609 ( \38588 , \38587 );
xor \U$38610 ( \38589 , \36677 , \36691 );
xor \U$38611 ( \38590 , \38589 , \36713 );
buf \U$38612 ( \38591 , \38590 );
buf \U$38613 ( \38592 , \38591 );
xor \U$38614 ( \38593 , \37681 , \37698 );
xor \U$38615 ( \38594 , \38593 , \37711 );
buf \U$38616 ( \38595 , \38594 );
buf \U$38617 ( \38596 , \38595 );
xor \U$38618 ( \38597 , \38592 , \38596 );
xor \U$38619 ( \38598 , \37510 , \37527 );
xor \U$38620 ( \38599 , \38598 , \37545 );
buf \U$38621 ( \38600 , \38599 );
buf \U$38622 ( \38601 , \38600 );
xor \U$38623 ( \38602 , \38597 , \38601 );
buf \U$38624 ( \38603 , \38602 );
buf \U$38625 ( \38604 , \38603 );
xor \U$38626 ( \38605 , \38588 , \38604 );
buf \U$38627 ( \38606 , \38188 );
buf \U$38628 ( \38607 , \38198 );
xor \U$38629 ( \38608 , \38606 , \38607 );
buf \U$38630 ( \38609 , \38205 );
xor \U$38631 ( \38610 , \38608 , \38609 );
buf \U$38632 ( \38611 , \38610 );
buf \U$38633 ( \38612 , \38611 );
and \U$38634 ( \38613 , \38605 , \38612 );
and \U$38635 ( \38614 , \38588 , \38604 );
or \U$38636 ( \38615 , \38613 , \38614 );
buf \U$38637 ( \38616 , \38615 );
buf \U$38638 ( \38617 , \38616 );
xor \U$38639 ( \38618 , \38529 , \38617 );
xor \U$38640 ( \38619 , \36782 , \36847 );
xor \U$38641 ( \38620 , \38619 , \36787 );
buf \U$38642 ( \38621 , \38620 );
not \U$38643 ( \38622 , \38621 );
buf \U$38644 ( \38623 , \38622 );
buf \U$38645 ( \38624 , \38623 );
not \U$38646 ( \38625 , \38624 );
buf \U$38647 ( \38626 , \38491 );
not \U$38648 ( \38627 , \38626 );
buf \U$38649 ( \38628 , \38627 );
buf \U$38650 ( \38629 , \38628 );
not \U$38651 ( \38630 , \38629 );
buf \U$38652 ( \38631 , \38511 );
not \U$38653 ( \38632 , \38631 );
or \U$38654 ( \38633 , \38630 , \38632 );
buf \U$38655 ( \38634 , \38474 );
nand \U$38656 ( \38635 , \38633 , \38634 );
buf \U$38657 ( \38636 , \38635 );
buf \U$38658 ( \38637 , \38636 );
buf \U$38659 ( \38638 , \38511 );
not \U$38660 ( \38639 , \38638 );
buf \U$38661 ( \38640 , \38491 );
nand \U$38662 ( \38641 , \38639 , \38640 );
buf \U$38663 ( \38642 , \38641 );
buf \U$38664 ( \38643 , \38642 );
nand \U$38665 ( \38644 , \38637 , \38643 );
buf \U$38666 ( \38645 , \38644 );
xor \U$38667 ( \38646 , \38592 , \38596 );
and \U$38668 ( \38647 , \38646 , \38601 );
and \U$38669 ( \38648 , \38592 , \38596 );
or \U$38670 ( \38649 , \38647 , \38648 );
buf \U$38671 ( \38650 , \38649 );
xor \U$38672 ( \38651 , \38645 , \38650 );
buf \U$38673 ( \38652 , \38651 );
not \U$38674 ( \38653 , \38652 );
or \U$38675 ( \38654 , \38625 , \38653 );
buf \U$38676 ( \38655 , \38651 );
buf \U$38677 ( \38656 , \38623 );
or \U$38678 ( \38657 , \38655 , \38656 );
nand \U$38679 ( \38658 , \38654 , \38657 );
buf \U$38680 ( \38659 , \38658 );
buf \U$38681 ( \38660 , \38659 );
and \U$38682 ( \38661 , \38618 , \38660 );
and \U$38683 ( \38662 , \38529 , \38617 );
or \U$38684 ( \38663 , \38661 , \38662 );
buf \U$38685 ( \38664 , \38663 );
buf \U$38686 ( \38665 , \38664 );
xor \U$38687 ( \38666 , \38452 , \38665 );
buf \U$38688 ( \38667 , \38650 );
buf \U$38689 ( \38668 , \38620 );
or \U$38690 ( \38669 , \38667 , \38668 );
buf \U$38691 ( \38670 , \38645 );
nand \U$38692 ( \38671 , \38669 , \38670 );
buf \U$38693 ( \38672 , \38671 );
buf \U$38694 ( \38673 , \38672 );
buf \U$38695 ( \38674 , \38650 );
buf \U$38696 ( \38675 , \38620 );
nand \U$38697 ( \38676 , \38674 , \38675 );
buf \U$38698 ( \38677 , \38676 );
buf \U$38699 ( \38678 , \38677 );
nand \U$38700 ( \38679 , \38673 , \38678 );
buf \U$38701 ( \38680 , \38679 );
buf \U$38702 ( \38681 , \38680 );
buf \U$38703 ( \38682 , \37573 );
not \U$38704 ( \38683 , \38682 );
buf \U$38705 ( \38684 , \37613 );
not \U$38706 ( \38685 , \38684 );
or \U$38707 ( \38686 , \38683 , \38685 );
buf \U$38708 ( \38687 , \37613 );
buf \U$38709 ( \38688 , \37573 );
or \U$38710 ( \38689 , \38687 , \38688 );
nand \U$38711 ( \38690 , \38686 , \38689 );
buf \U$38712 ( \38691 , \38690 );
buf \U$38713 ( \38692 , \38691 );
buf \U$38714 ( \38693 , \37580 );
xor \U$38715 ( \38694 , \38692 , \38693 );
buf \U$38716 ( \38695 , \38694 );
buf \U$38717 ( \38696 , \38695 );
buf \U$38718 ( \38697 , \37549 );
buf \U$38719 ( \38698 , \37487 );
not \U$38720 ( \38699 , \38698 );
buf \U$38721 ( \38700 , \37417 );
not \U$38722 ( \38701 , \38700 );
or \U$38723 ( \38702 , \38699 , \38701 );
buf \U$38724 ( \38703 , \37490 );
buf \U$38725 ( \38704 , \37414 );
nand \U$38726 ( \38705 , \38703 , \38704 );
buf \U$38727 ( \38706 , \38705 );
buf \U$38728 ( \38707 , \38706 );
nand \U$38729 ( \38708 , \38702 , \38707 );
buf \U$38730 ( \38709 , \38708 );
buf \U$38731 ( \38710 , \38709 );
xor \U$38732 ( \38711 , \38697 , \38710 );
buf \U$38733 ( \38712 , \38711 );
buf \U$38734 ( \38713 , \38712 );
or \U$38735 ( \38714 , \38696 , \38713 );
buf \U$38736 ( \38715 , \37305 );
not \U$38737 ( \38716 , \38715 );
buf \U$38738 ( \38717 , \37328 );
not \U$38739 ( \38718 , \38717 );
or \U$38740 ( \38719 , \38716 , \38718 );
buf \U$38741 ( \38720 , \37305 );
buf \U$38742 ( \38721 , \37328 );
or \U$38743 ( \38722 , \38720 , \38721 );
nand \U$38744 ( \38723 , \38719 , \38722 );
buf \U$38745 ( \38724 , \38723 );
buf \U$38746 ( \38725 , \38724 );
buf \U$38747 ( \38726 , \37298 );
and \U$38748 ( \38727 , \38725 , \38726 );
not \U$38749 ( \38728 , \38725 );
buf \U$38750 ( \38729 , \37295 );
and \U$38751 ( \38730 , \38728 , \38729 );
nor \U$38752 ( \38731 , \38727 , \38730 );
buf \U$38753 ( \38732 , \38731 );
buf \U$38754 ( \38733 , \38732 );
nand \U$38755 ( \38734 , \38714 , \38733 );
buf \U$38756 ( \38735 , \38734 );
buf \U$38757 ( \38736 , \38735 );
buf \U$38758 ( \38737 , \38695 );
buf \U$38759 ( \38738 , \38712 );
nand \U$38760 ( \38739 , \38737 , \38738 );
buf \U$38761 ( \38740 , \38739 );
buf \U$38762 ( \38741 , \38740 );
nand \U$38763 ( \38742 , \38736 , \38741 );
buf \U$38764 ( \38743 , \38742 );
buf \U$38765 ( \38744 , \38743 );
xor \U$38766 ( \38745 , \38681 , \38744 );
buf \U$38767 ( \38746 , \37334 );
not \U$38768 ( \38747 , \38746 );
buf \U$38769 ( \38748 , \37290 );
not \U$38770 ( \38749 , \38748 );
or \U$38771 ( \38750 , \38747 , \38749 );
buf \U$38772 ( \38751 , \37290 );
buf \U$38773 ( \38752 , \37334 );
or \U$38774 ( \38753 , \38751 , \38752 );
nand \U$38775 ( \38754 , \38750 , \38753 );
buf \U$38776 ( \38755 , \38754 );
buf \U$38777 ( \38756 , \38755 );
buf \U$38778 ( \38757 , \37342 );
and \U$38779 ( \38758 , \38756 , \38757 );
not \U$38780 ( \38759 , \38756 );
buf \U$38781 ( \38760 , \37093 );
and \U$38782 ( \38761 , \38759 , \38760 );
nor \U$38783 ( \38762 , \38758 , \38761 );
buf \U$38784 ( \38763 , \38762 );
buf \U$38785 ( \38764 , \38763 );
xor \U$38786 ( \38765 , \38745 , \38764 );
buf \U$38787 ( \38766 , \38765 );
buf \U$38788 ( \38767 , \38766 );
and \U$38789 ( \38768 , \38666 , \38767 );
and \U$38790 ( \38769 , \38452 , \38665 );
or \U$38791 ( \38770 , \38768 , \38769 );
buf \U$38792 ( \38771 , \38770 );
buf \U$38793 ( \38772 , \38771 );
not \U$38794 ( \38773 , \38772 );
and \U$38795 ( \38774 , \38237 , \38773 );
buf \U$38796 ( \38775 , \38771 );
buf \U$38797 ( \38776 , \38235 );
and \U$38798 ( \38777 , \38775 , \38776 );
nor \U$38799 ( \38778 , \38774 , \38777 );
buf \U$38800 ( \38779 , \38778 );
buf \U$38801 ( \38780 , \38779 );
not \U$38802 ( \38781 , \38780 );
buf \U$38803 ( \38782 , \38781 );
buf \U$38804 ( \38783 , \38782 );
xor \U$38805 ( \38784 , \38016 , \38020 );
and \U$38806 ( \38785 , \38784 , \38220 );
and \U$38807 ( \38786 , \38016 , \38020 );
or \U$38808 ( \38787 , \38785 , \38786 );
buf \U$38809 ( \38788 , \38787 );
buf \U$38810 ( \38789 , \38788 );
buf \U$38811 ( \38790 , \35870 );
not \U$38812 ( \38791 , \38790 );
buf \U$38813 ( \38792 , \16744 );
not \U$38814 ( \38793 , \38792 );
or \U$38815 ( \38794 , \38791 , \38793 );
buf \U$38816 ( \38795 , \2476 );
buf \U$38817 ( \38796 , RIc0da468_99);
buf \U$38818 ( \38797 , RIc0d79c0_8);
xor \U$38819 ( \38798 , \38796 , \38797 );
buf \U$38820 ( \38799 , \38798 );
buf \U$38821 ( \38800 , \38799 );
nand \U$38822 ( \38801 , \38795 , \38800 );
buf \U$38823 ( \38802 , \38801 );
buf \U$38824 ( \38803 , \38802 );
nand \U$38825 ( \38804 , \38794 , \38803 );
buf \U$38826 ( \38805 , \38804 );
buf \U$38827 ( \38806 , \38805 );
not \U$38828 ( \38807 , \38806 );
and \U$38829 ( \38808 , \35600 , \35601 );
buf \U$38830 ( \38809 , \38808 );
buf \U$38831 ( \38810 , \38809 );
not \U$38832 ( \38811 , \38810 );
and \U$38833 ( \38812 , \38807 , \38811 );
buf \U$38834 ( \38813 , \38805 );
buf \U$38835 ( \38814 , \38809 );
and \U$38836 ( \38815 , \38813 , \38814 );
nor \U$38837 ( \38816 , \38812 , \38815 );
buf \U$38838 ( \38817 , \38816 );
buf \U$38839 ( \38818 , \38817 );
not \U$38840 ( \38819 , \38818 );
not \U$38841 ( \38820 , \37255 );
buf \U$38842 ( \38821 , \38820 );
not \U$38843 ( \38822 , \38821 );
buf \U$38844 ( \38823 , \37274 );
not \U$38845 ( \38824 , \38823 );
or \U$38846 ( \38825 , \38822 , \38824 );
buf \U$38847 ( \38826 , \37243 );
nand \U$38848 ( \38827 , \38825 , \38826 );
buf \U$38849 ( \38828 , \38827 );
buf \U$38850 ( \38829 , \38828 );
or \U$38851 ( \38830 , \37274 , \38820 );
buf \U$38852 ( \38831 , \38830 );
nand \U$38853 ( \38832 , \38829 , \38831 );
buf \U$38854 ( \38833 , \38832 );
buf \U$38855 ( \38834 , \38833 );
not \U$38856 ( \38835 , \38834 );
or \U$38857 ( \38836 , \38819 , \38835 );
buf \U$38858 ( \38837 , \38833 );
buf \U$38859 ( \38838 , \38817 );
or \U$38860 ( \38839 , \38837 , \38838 );
nand \U$38861 ( \38840 , \38836 , \38839 );
buf \U$38862 ( \38841 , \38840 );
buf \U$38863 ( \38842 , \38841 );
buf \U$38864 ( \38843 , \36968 );
not \U$38865 ( \38844 , \38843 );
buf \U$38866 ( \38845 , \37090 );
not \U$38867 ( \38846 , \38845 );
or \U$38868 ( \38847 , \38844 , \38846 );
buf \U$38869 ( \38848 , \37090 );
buf \U$38870 ( \38849 , \36968 );
or \U$38871 ( \38850 , \38848 , \38849 );
buf \U$38872 ( \38851 , \37030 );
nand \U$38873 ( \38852 , \38850 , \38851 );
buf \U$38874 ( \38853 , \38852 );
buf \U$38875 ( \38854 , \38853 );
nand \U$38876 ( \38855 , \38847 , \38854 );
buf \U$38877 ( \38856 , \38855 );
buf \U$38878 ( \38857 , \38856 );
xor \U$38879 ( \38858 , \38842 , \38857 );
xor \U$38880 ( \38859 , \36128 , \36149 );
and \U$38881 ( \38860 , \38859 , \36171 );
and \U$38882 ( \38861 , \36128 , \36149 );
or \U$38883 ( \38862 , \38860 , \38861 );
buf \U$38884 ( \38863 , \38862 );
buf \U$38885 ( \38864 , \38863 );
xor \U$38886 ( \38865 , \35810 , \35831 );
and \U$38887 ( \38866 , \38865 , \35853 );
and \U$38888 ( \38867 , \35810 , \35831 );
or \U$38889 ( \38868 , \38866 , \38867 );
buf \U$38890 ( \38869 , \38868 );
buf \U$38891 ( \38870 , \38869 );
xor \U$38892 ( \38871 , \38864 , \38870 );
buf \U$38893 ( \38872 , \35889 );
not \U$38894 ( \38873 , \38872 );
buf \U$38895 ( \38874 , \35911 );
not \U$38896 ( \38875 , \38874 );
or \U$38897 ( \38876 , \38873 , \38875 );
buf \U$38898 ( \38877 , \35911 );
buf \U$38899 ( \38878 , \35889 );
or \U$38900 ( \38879 , \38877 , \38878 );
buf \U$38901 ( \38880 , \35876 );
nand \U$38902 ( \38881 , \38879 , \38880 );
buf \U$38903 ( \38882 , \38881 );
buf \U$38904 ( \38883 , \38882 );
nand \U$38905 ( \38884 , \38876 , \38883 );
buf \U$38906 ( \38885 , \38884 );
buf \U$38907 ( \38886 , \38885 );
xor \U$38908 ( \38887 , \38871 , \38886 );
buf \U$38909 ( \38888 , \38887 );
buf \U$38910 ( \38889 , \38888 );
xor \U$38911 ( \38890 , \38858 , \38889 );
buf \U$38912 ( \38891 , \38890 );
buf \U$38913 ( \38892 , \38891 );
xor \U$38914 ( \38893 , \37561 , \37623 );
and \U$38915 ( \38894 , \38893 , \37726 );
and \U$38916 ( \38895 , \37561 , \37623 );
or \U$38917 ( \38896 , \38894 , \38895 );
buf \U$38918 ( \38897 , \38896 );
buf \U$38919 ( \38898 , \38897 );
xor \U$38920 ( \38899 , \38892 , \38898 );
buf \U$38921 ( \38900 , \35921 );
not \U$38922 ( \38901 , \38900 );
buf \U$38923 ( \38902 , \35858 );
not \U$38924 ( \38903 , \38902 );
or \U$38925 ( \38904 , \38901 , \38903 );
buf \U$38926 ( \38905 , \35987 );
nand \U$38927 ( \38906 , \38904 , \38905 );
buf \U$38928 ( \38907 , \38906 );
buf \U$38929 ( \38908 , \38907 );
buf \U$38930 ( \38909 , \35921 );
not \U$38931 ( \38910 , \38909 );
buf \U$38932 ( \38911 , \35855 );
nand \U$38933 ( \38912 , \38910 , \38911 );
buf \U$38934 ( \38913 , \38912 );
buf \U$38935 ( \38914 , \38913 );
nand \U$38936 ( \38915 , \38908 , \38914 );
buf \U$38937 ( \38916 , \38915 );
buf \U$38938 ( \38917 , \36173 );
not \U$38939 ( \38918 , \38917 );
buf \U$38940 ( \38919 , \36041 );
not \U$38941 ( \38920 , \38919 );
or \U$38942 ( \38921 , \38918 , \38920 );
buf \U$38943 ( \38922 , \36173 );
buf \U$38944 ( \38923 , \36041 );
or \U$38945 ( \38924 , \38922 , \38923 );
buf \U$38946 ( \38925 , \36114 );
nand \U$38947 ( \38926 , \38924 , \38925 );
buf \U$38948 ( \38927 , \38926 );
buf \U$38949 ( \38928 , \38927 );
nand \U$38950 ( \38929 , \38921 , \38928 );
buf \U$38951 ( \38930 , \38929 );
xor \U$38952 ( \38931 , \38916 , \38930 );
buf \U$38953 ( \38932 , \37221 );
not \U$38954 ( \38933 , \38932 );
buf \U$38955 ( \38934 , \37282 );
not \U$38956 ( \38935 , \38934 );
or \U$38957 ( \38936 , \38933 , \38935 );
buf \U$38958 ( \38937 , \37157 );
nand \U$38959 ( \38938 , \38936 , \38937 );
buf \U$38960 ( \38939 , \38938 );
buf \U$38961 ( \38940 , \38939 );
buf \U$38962 ( \38941 , \37282 );
not \U$38963 ( \38942 , \38941 );
buf \U$38964 ( \38943 , \37218 );
nand \U$38965 ( \38944 , \38942 , \38943 );
buf \U$38966 ( \38945 , \38944 );
buf \U$38967 ( \38946 , \38945 );
nand \U$38968 ( \38947 , \38940 , \38946 );
buf \U$38969 ( \38948 , \38947 );
xor \U$38970 ( \38949 , \38931 , \38948 );
buf \U$38971 ( \38950 , \38949 );
xor \U$38972 ( \38951 , \38899 , \38950 );
buf \U$38973 ( \38952 , \38951 );
buf \U$38974 ( \38953 , \38952 );
xor \U$38975 ( \38954 , \38789 , \38953 );
xor \U$38976 ( \38955 , \38681 , \38744 );
and \U$38977 ( \38956 , \38955 , \38764 );
and \U$38978 ( \38957 , \38681 , \38744 );
or \U$38979 ( \38958 , \38956 , \38957 );
buf \U$38980 ( \38959 , \38958 );
buf \U$38981 ( \38960 , \38959 );
xor \U$38982 ( \38961 , \38954 , \38960 );
buf \U$38983 ( \38962 , \38961 );
buf \U$38984 ( \38963 , \38962 );
or \U$38985 ( \38964 , \38783 , \38963 );
buf \U$38986 ( \38965 , \38732 );
buf \U$38987 ( \38966 , \38712 );
and \U$38988 ( \38967 , \38965 , \38966 );
not \U$38989 ( \38968 , \38965 );
buf \U$38990 ( \38969 , \38712 );
not \U$38991 ( \38970 , \38969 );
buf \U$38992 ( \38971 , \38970 );
buf \U$38993 ( \38972 , \38971 );
and \U$38994 ( \38973 , \38968 , \38972 );
nor \U$38995 ( \38974 , \38967 , \38973 );
buf \U$38996 ( \38975 , \38974 );
buf \U$38997 ( \38976 , \38975 );
buf \U$38998 ( \38977 , \38695 );
and \U$38999 ( \38978 , \38976 , \38977 );
not \U$39000 ( \38979 , \38976 );
buf \U$39001 ( \38980 , \38695 );
not \U$39002 ( \38981 , \38980 );
buf \U$39003 ( \38982 , \38981 );
buf \U$39004 ( \38983 , \38982 );
and \U$39005 ( \38984 , \38979 , \38983 );
nor \U$39006 ( \38985 , \38978 , \38984 );
buf \U$39007 ( \38986 , \38985 );
buf \U$39008 ( \38987 , \38986 );
xor \U$39009 ( \38988 , \38182 , \38210 );
xor \U$39010 ( \38989 , \38988 , \38215 );
buf \U$39011 ( \38990 , \38989 );
buf \U$39012 ( \38991 , \38990 );
xor \U$39013 ( \38992 , \38987 , \38991 );
not \U$39014 ( \38993 , \33699 );
nand \U$39015 ( \38994 , \38993 , \33735 );
not \U$39016 ( \38995 , \38994 );
not \U$39017 ( \38996 , \33714 );
or \U$39018 ( \38997 , \38995 , \38996 );
buf \U$39019 ( \38998 , \33699 );
buf \U$39020 ( \38999 , \33732 );
nand \U$39021 ( \39000 , \38998 , \38999 );
buf \U$39022 ( \39001 , \39000 );
nand \U$39023 ( \39002 , \38997 , \39001 );
buf \U$39024 ( \39003 , \39002 );
buf \U$39025 ( \39004 , \33848 );
not \U$39026 ( \39005 , \39004 );
buf \U$39027 ( \39006 , \33827 );
not \U$39028 ( \39007 , \39006 );
or \U$39029 ( \39008 , \39005 , \39007 );
buf \U$39030 ( \39009 , \33848 );
buf \U$39031 ( \39010 , \33827 );
or \U$39032 ( \39011 , \39009 , \39010 );
buf \U$39033 ( \39012 , \33831 );
nand \U$39034 ( \39013 , \39011 , \39012 );
buf \U$39035 ( \39014 , \39013 );
buf \U$39036 ( \39015 , \39014 );
nand \U$39037 ( \39016 , \39008 , \39015 );
buf \U$39038 ( \39017 , \39016 );
buf \U$39039 ( \39018 , \39017 );
xor \U$39040 ( \39019 , \39003 , \39018 );
xor \U$39041 ( \39020 , \38249 , \38267 );
xor \U$39042 ( \39021 , \39020 , \38274 );
buf \U$39043 ( \39022 , \39021 );
buf \U$39044 ( \39023 , \39022 );
and \U$39045 ( \39024 , \39019 , \39023 );
and \U$39046 ( \39025 , \39003 , \39018 );
or \U$39047 ( \39026 , \39024 , \39025 );
buf \U$39048 ( \39027 , \39026 );
buf \U$39049 ( \39028 , \39027 );
xor \U$39050 ( \39029 , \38245 , \38279 );
xor \U$39051 ( \39030 , \39029 , \38304 );
buf \U$39052 ( \39031 , \39030 );
buf \U$39053 ( \39032 , \39031 );
xor \U$39054 ( \39033 , \39028 , \39032 );
buf \U$39055 ( \39034 , \34071 );
buf \U$39056 ( \39035 , \34126 );
or \U$39057 ( \39036 , \39034 , \39035 );
buf \U$39058 ( \39037 , \34022 );
nand \U$39059 ( \39038 , \39036 , \39037 );
buf \U$39060 ( \39039 , \39038 );
buf \U$39061 ( \39040 , \39039 );
buf \U$39062 ( \39041 , \34126 );
buf \U$39063 ( \39042 , \34071 );
nand \U$39064 ( \39043 , \39041 , \39042 );
buf \U$39065 ( \39044 , \39043 );
buf \U$39066 ( \39045 , \39044 );
nand \U$39067 ( \39046 , \39040 , \39045 );
buf \U$39068 ( \39047 , \39046 );
buf \U$39069 ( \39048 , \39047 );
buf \U$39070 ( \39049 , \34273 );
not \U$39071 ( \39050 , \39049 );
buf \U$39072 ( \39051 , \34219 );
not \U$39073 ( \39052 , \39051 );
or \U$39074 ( \39053 , \39050 , \39052 );
buf \U$39075 ( \39054 , \34219 );
buf \U$39076 ( \39055 , \34273 );
or \U$39077 ( \39056 , \39054 , \39055 );
buf \U$39078 ( \39057 , \34325 );
not \U$39079 ( \39058 , \39057 );
buf \U$39080 ( \39059 , \39058 );
buf \U$39081 ( \39060 , \39059 );
nand \U$39082 ( \39061 , \39056 , \39060 );
buf \U$39083 ( \39062 , \39061 );
buf \U$39084 ( \39063 , \39062 );
nand \U$39085 ( \39064 , \39053 , \39063 );
buf \U$39086 ( \39065 , \39064 );
buf \U$39087 ( \39066 , \39065 );
xor \U$39088 ( \39067 , \39048 , \39066 );
xor \U$39089 ( \39068 , \38286 , \38292 );
xor \U$39090 ( \39069 , \39068 , \38299 );
buf \U$39091 ( \39070 , \39069 );
buf \U$39092 ( \39071 , \39070 );
and \U$39093 ( \39072 , \39067 , \39071 );
and \U$39094 ( \39073 , \39048 , \39066 );
or \U$39095 ( \39074 , \39072 , \39073 );
buf \U$39096 ( \39075 , \39074 );
buf \U$39097 ( \39076 , \39075 );
and \U$39098 ( \39077 , \39033 , \39076 );
and \U$39099 ( \39078 , \39028 , \39032 );
or \U$39100 ( \39079 , \39077 , \39078 );
buf \U$39101 ( \39080 , \39079 );
buf \U$39102 ( \39081 , \39080 );
and \U$39103 ( \39082 , \38992 , \39081 );
and \U$39104 ( \39083 , \38987 , \38991 );
or \U$39105 ( \39084 , \39082 , \39083 );
buf \U$39106 ( \39085 , \39084 );
buf \U$39107 ( \39086 , \39085 );
xor \U$39108 ( \39087 , \37729 , \37733 );
xor \U$39109 ( \39088 , \39087 , \38223 );
buf \U$39110 ( \39089 , \39088 );
buf \U$39111 ( \39090 , \39089 );
xor \U$39112 ( \39091 , \39086 , \39090 );
xor \U$39113 ( \39092 , \38452 , \38665 );
xor \U$39114 ( \39093 , \39092 , \38767 );
buf \U$39115 ( \39094 , \39093 );
buf \U$39116 ( \39095 , \39094 );
and \U$39117 ( \39096 , \39091 , \39095 );
and \U$39118 ( \39097 , \39086 , \39090 );
or \U$39119 ( \39098 , \39096 , \39097 );
buf \U$39120 ( \39099 , \39098 );
buf \U$39121 ( \39100 , \39099 );
nand \U$39122 ( \39101 , \38964 , \39100 );
buf \U$39123 ( \39102 , \39101 );
buf \U$39124 ( \39103 , \39102 );
buf \U$39125 ( \39104 , \38782 );
buf \U$39126 ( \39105 , \38962 );
nand \U$39127 ( \39106 , \39104 , \39105 );
buf \U$39128 ( \39107 , \39106 );
buf \U$39129 ( \39108 , \39107 );
nand \U$39130 ( \39109 , \39103 , \39108 );
buf \U$39131 ( \39110 , \39109 );
buf \U$39132 ( \39111 , \39110 );
not \U$39133 ( \39112 , \39111 );
buf \U$39134 ( \39113 , \39112 );
buf \U$39135 ( \39114 , \39113 );
buf \U$39136 ( \39115 , \36356 );
not \U$39137 ( \39116 , \39115 );
buf \U$39138 ( \39117 , \1736 );
not \U$39139 ( \39118 , \39117 );
or \U$39140 ( \39119 , \39116 , \39118 );
xnor \U$39141 ( \39120 , RIc0d9ce8_83, RIc0d80c8_23);
buf \U$39142 ( \39121 , \39120 );
not \U$39143 ( \39122 , \39121 );
buf \U$39144 ( \39123 , \993 );
nand \U$39145 ( \39124 , \39122 , \39123 );
buf \U$39146 ( \39125 , \39124 );
buf \U$39147 ( \39126 , \39125 );
nand \U$39148 ( \39127 , \39119 , \39126 );
buf \U$39149 ( \39128 , \39127 );
buf \U$39150 ( \39129 , \13270 );
not \U$39151 ( \39130 , \39129 );
buf \U$39152 ( \39131 , \12331 );
not \U$39153 ( \39132 , \39131 );
or \U$39154 ( \39133 , \39130 , \39132 );
buf \U$39155 ( \39134 , RIc0da828_107);
nand \U$39156 ( \39135 , \39133 , \39134 );
buf \U$39157 ( \39136 , \39135 );
xor \U$39158 ( \39137 , \39128 , \39136 );
buf \U$39159 ( \39138 , \36869 );
not \U$39160 ( \39139 , \39138 );
buf \U$39161 ( \39140 , \4692 );
not \U$39162 ( \39141 , \39140 );
or \U$39163 ( \39142 , \39139 , \39141 );
buf \U$39164 ( \39143 , \874 );
buf \U$39165 ( \39144 , RIc0d9658_69);
buf \U$39166 ( \39145 , RIc0d8758_37);
xor \U$39167 ( \39146 , \39144 , \39145 );
buf \U$39168 ( \39147 , \39146 );
buf \U$39169 ( \39148 , \39147 );
nand \U$39170 ( \39149 , \39143 , \39148 );
buf \U$39171 ( \39150 , \39149 );
buf \U$39172 ( \39151 , \39150 );
nand \U$39173 ( \39152 , \39142 , \39151 );
buf \U$39174 ( \39153 , \39152 );
xnor \U$39175 ( \39154 , \39137 , \39153 );
buf \U$39176 ( \39155 , \38799 );
not \U$39177 ( \39156 , \39155 );
buf \U$39178 ( \39157 , \21461 );
not \U$39179 ( \39158 , \39157 );
or \U$39180 ( \39159 , \39156 , \39158 );
buf \U$39181 ( \39160 , \22006 );
buf \U$39182 ( \39161 , RIc0da468_99);
buf \U$39183 ( \39162 , RIc0d7948_7);
xor \U$39184 ( \39163 , \39161 , \39162 );
buf \U$39185 ( \39164 , \39163 );
buf \U$39186 ( \39165 , \39164 );
nand \U$39187 ( \39166 , \39160 , \39165 );
buf \U$39188 ( \39167 , \39166 );
buf \U$39189 ( \39168 , \39167 );
nand \U$39190 ( \39169 , \39159 , \39168 );
buf \U$39191 ( \39170 , \39169 );
buf \U$39192 ( \39171 , \39170 );
buf \U$39193 ( \39172 , \36917 );
not \U$39194 ( \39173 , \39172 );
buf \U$39195 ( \39174 , \4527 );
not \U$39196 ( \39175 , \39174 );
or \U$39197 ( \39176 , \39173 , \39175 );
buf \U$39198 ( \39177 , \14331 );
xor \U$39199 ( \39178 , RIc0d9ec8_87, RIc0d7ee8_19);
buf \U$39200 ( \39179 , \39178 );
nand \U$39201 ( \39180 , \39177 , \39179 );
buf \U$39202 ( \39181 , \39180 );
buf \U$39203 ( \39182 , \39181 );
nand \U$39204 ( \39183 , \39176 , \39182 );
buf \U$39205 ( \39184 , \39183 );
buf \U$39206 ( \39185 , \39184 );
xor \U$39207 ( \39186 , \39171 , \39185 );
buf \U$39208 ( \39187 , \39186 );
buf \U$39209 ( \39188 , \39187 );
buf \U$39210 ( \39189 , \36946 );
not \U$39211 ( \39190 , \39189 );
buf \U$39212 ( \39191 , \12442 );
not \U$39213 ( \39192 , \39191 );
or \U$39214 ( \39193 , \39190 , \39192 );
buf \U$39215 ( \39194 , \791 );
buf \U$39216 ( \39195 , RIc0d9838_73);
buf \U$39217 ( \39196 , RIc0d8578_33);
xor \U$39218 ( \39197 , \39195 , \39196 );
buf \U$39219 ( \39198 , \39197 );
buf \U$39220 ( \39199 , \39198 );
nand \U$39221 ( \39200 , \39194 , \39199 );
buf \U$39222 ( \39201 , \39200 );
buf \U$39223 ( \39202 , \39201 );
nand \U$39224 ( \39203 , \39193 , \39202 );
buf \U$39225 ( \39204 , \39203 );
buf \U$39226 ( \39205 , \39204 );
and \U$39227 ( \39206 , \39188 , \39205 );
not \U$39228 ( \39207 , \39188 );
buf \U$39229 ( \39208 , \39204 );
not \U$39230 ( \39209 , \39208 );
buf \U$39231 ( \39210 , \39209 );
buf \U$39232 ( \39211 , \39210 );
and \U$39233 ( \39212 , \39207 , \39211 );
nor \U$39234 ( \39213 , \39206 , \39212 );
buf \U$39235 ( \39214 , \39213 );
xor \U$39236 ( \39215 , \39154 , \39214 );
buf \U$39237 ( \39216 , \36432 );
not \U$39238 ( \39217 , \39216 );
buf \U$39239 ( \39218 , \13042 );
not \U$39240 ( \39219 , \39218 );
or \U$39241 ( \39220 , \39217 , \39219 );
buf \U$39242 ( \39221 , \20243 );
buf \U$39243 ( \39222 , RIc0d7768_3);
buf \U$39244 ( \39223 , RIc0da648_103);
xor \U$39245 ( \39224 , \39222 , \39223 );
buf \U$39246 ( \39225 , \39224 );
buf \U$39247 ( \39226 , \39225 );
nand \U$39248 ( \39227 , \39221 , \39226 );
buf \U$39249 ( \39228 , \39227 );
buf \U$39250 ( \39229 , \39228 );
nand \U$39251 ( \39230 , \39220 , \39229 );
buf \U$39252 ( \39231 , \39230 );
buf \U$39253 ( \39232 , \36318 );
not \U$39254 ( \39233 , \39232 );
buf \U$39255 ( \39234 , \15644 );
not \U$39256 ( \39235 , \39234 );
or \U$39257 ( \39236 , \39233 , \39235 );
buf \U$39258 ( \39237 , \15653 );
buf \U$39259 ( \39238 , RIc0da738_105);
buf \U$39260 ( \39239 , RIc0d7678_1);
and \U$39261 ( \39240 , \39238 , \39239 );
not \U$39262 ( \39241 , \39238 );
buf \U$39263 ( \39242 , \974 );
and \U$39264 ( \39243 , \39241 , \39242 );
nor \U$39265 ( \39244 , \39240 , \39243 );
buf \U$39266 ( \39245 , \39244 );
buf \U$39267 ( \39246 , \39245 );
nand \U$39268 ( \39247 , \39237 , \39246 );
buf \U$39269 ( \39248 , \39247 );
buf \U$39270 ( \39249 , \39248 );
nand \U$39271 ( \39250 , \39236 , \39249 );
buf \U$39272 ( \39251 , \39250 );
xor \U$39273 ( \39252 , \39231 , \39251 );
buf \U$39274 ( \39253 , \39252 );
buf \U$39275 ( \39254 , \38805 );
and \U$39276 ( \39255 , \39253 , \39254 );
not \U$39277 ( \39256 , \39253 );
buf \U$39278 ( \39257 , \38805 );
not \U$39279 ( \39258 , \39257 );
buf \U$39280 ( \39259 , \39258 );
buf \U$39281 ( \39260 , \39259 );
and \U$39282 ( \39261 , \39256 , \39260 );
nor \U$39283 ( \39262 , \39255 , \39261 );
buf \U$39284 ( \39263 , \39262 );
xnor \U$39285 ( \39264 , \39215 , \39263 );
buf \U$39286 ( \39265 , \39264 );
xor \U$39287 ( \39266 , \36907 , \36954 );
and \U$39288 ( \39267 , \39266 , \36961 );
and \U$39289 ( \39268 , \36907 , \36954 );
or \U$39290 ( \39269 , \39267 , \39268 );
buf \U$39291 ( \39270 , \39269 );
buf \U$39292 ( \39271 , \39270 );
xor \U$39293 ( \39272 , \39265 , \39271 );
buf \U$39294 ( \39273 , \38930 );
buf \U$39295 ( \39274 , \38948 );
or \U$39296 ( \39275 , \39273 , \39274 );
buf \U$39297 ( \39276 , \38916 );
nand \U$39298 ( \39277 , \39275 , \39276 );
buf \U$39299 ( \39278 , \39277 );
buf \U$39300 ( \39279 , \39278 );
buf \U$39301 ( \39280 , \38930 );
buf \U$39302 ( \39281 , \38948 );
nand \U$39303 ( \39282 , \39280 , \39281 );
buf \U$39304 ( \39283 , \39282 );
buf \U$39305 ( \39284 , \39283 );
nand \U$39306 ( \39285 , \39279 , \39284 );
buf \U$39307 ( \39286 , \39285 );
buf \U$39308 ( \39287 , \39286 );
xor \U$39309 ( \39288 , \39272 , \39287 );
buf \U$39310 ( \39289 , \39288 );
buf \U$39311 ( \39290 , \39289 );
xor \U$39312 ( \39291 , \38892 , \38898 );
and \U$39313 ( \39292 , \39291 , \38950 );
and \U$39314 ( \39293 , \38892 , \38898 );
or \U$39315 ( \39294 , \39292 , \39293 );
buf \U$39316 ( \39295 , \39294 );
buf \U$39317 ( \39296 , \39295 );
xor \U$39318 ( \39297 , \39290 , \39296 );
xor \U$39319 ( \39298 , \36328 , \36388 );
and \U$39320 ( \39299 , \39298 , \36442 );
and \U$39321 ( \39300 , \36328 , \36388 );
or \U$39322 ( \39301 , \39299 , \39300 );
buf \U$39323 ( \39302 , \39301 );
buf \U$39324 ( \39303 , \39302 );
not \U$39325 ( \39304 , \39303 );
xor \U$39326 ( \39305 , \36349 , \36363 );
and \U$39327 ( \39306 , \39305 , \36385 );
and \U$39328 ( \39307 , \36349 , \36363 );
or \U$39329 ( \39308 , \39306 , \39307 );
buf \U$39330 ( \39309 , \39308 );
xor \U$39331 ( \39310 , \36293 , \36307 );
and \U$39332 ( \39311 , \39310 , \36325 );
and \U$39333 ( \39312 , \36293 , \36307 );
or \U$39334 ( \39313 , \39311 , \39312 );
buf \U$39335 ( \39314 , \39313 );
xor \U$39336 ( \39315 , \39309 , \39314 );
buf \U$39337 ( \39316 , \36527 );
not \U$39338 ( \39317 , \39316 );
buf \U$39339 ( \39318 , \39317 );
buf \U$39340 ( \39319 , \39318 );
not \U$39341 ( \39320 , \39319 );
buf \U$39342 ( \39321 , \36506 );
not \U$39343 ( \39322 , \39321 );
or \U$39344 ( \39323 , \39320 , \39322 );
buf \U$39345 ( \39324 , \36527 );
not \U$39346 ( \39325 , \39324 );
buf \U$39347 ( \39326 , \36509 );
not \U$39348 ( \39327 , \39326 );
or \U$39349 ( \39328 , \39325 , \39327 );
buf \U$39350 ( \39329 , \36486 );
nand \U$39351 ( \39330 , \39328 , \39329 );
buf \U$39352 ( \39331 , \39330 );
buf \U$39353 ( \39332 , \39331 );
nand \U$39354 ( \39333 , \39323 , \39332 );
buf \U$39355 ( \39334 , \39333 );
xnor \U$39356 ( \39335 , \39315 , \39334 );
buf \U$39357 ( \39336 , \39335 );
not \U$39358 ( \39337 , \39336 );
or \U$39359 ( \39338 , \39304 , \39337 );
buf \U$39360 ( \39339 , \39302 );
buf \U$39361 ( \39340 , \39335 );
or \U$39362 ( \39341 , \39339 , \39340 );
nand \U$39363 ( \39342 , \39338 , \39341 );
buf \U$39364 ( \39343 , \39342 );
buf \U$39365 ( \39344 , \39343 );
xor \U$39366 ( \39345 , \36473 , \36529 );
and \U$39367 ( \39346 , \39345 , \36575 );
and \U$39368 ( \39347 , \36473 , \36529 );
or \U$39369 ( \39348 , \39346 , \39347 );
buf \U$39370 ( \39349 , \39348 );
buf \U$39371 ( \39350 , \39349 );
not \U$39372 ( \39351 , \39350 );
buf \U$39373 ( \39352 , \39351 );
buf \U$39374 ( \39353 , \39352 );
and \U$39375 ( \39354 , \39344 , \39353 );
not \U$39376 ( \39355 , \39344 );
buf \U$39377 ( \39356 , \39349 );
and \U$39378 ( \39357 , \39355 , \39356 );
nor \U$39379 ( \39358 , \39354 , \39357 );
buf \U$39380 ( \39359 , \39358 );
buf \U$39381 ( \39360 , \39359 );
not \U$39382 ( \39361 , \39360 );
xor \U$39383 ( \39362 , \38842 , \38857 );
and \U$39384 ( \39363 , \39362 , \38889 );
and \U$39385 ( \39364 , \38842 , \38857 );
or \U$39386 ( \39365 , \39363 , \39364 );
buf \U$39387 ( \39366 , \39365 );
buf \U$39388 ( \39367 , \39366 );
not \U$39389 ( \39368 , \39367 );
buf \U$39390 ( \39369 , \38809 );
not \U$39391 ( \39370 , \39369 );
buf \U$39392 ( \39371 , \38805 );
nand \U$39393 ( \39372 , \39370 , \39371 );
buf \U$39394 ( \39373 , \39372 );
buf \U$39395 ( \39374 , \39373 );
not \U$39396 ( \39375 , \39374 );
buf \U$39397 ( \39376 , \38833 );
not \U$39398 ( \39377 , \39376 );
or \U$39399 ( \39378 , \39375 , \39377 );
buf \U$39400 ( \39379 , \39259 );
buf \U$39401 ( \39380 , \38809 );
nand \U$39402 ( \39381 , \39379 , \39380 );
buf \U$39403 ( \39382 , \39381 );
buf \U$39404 ( \39383 , \39382 );
nand \U$39405 ( \39384 , \39378 , \39383 );
buf \U$39406 ( \39385 , \39384 );
buf \U$39407 ( \39386 , \39385 );
buf \U$39408 ( \39387 , \36266 );
not \U$39409 ( \39388 , \39387 );
buf \U$39410 ( \39389 , \36252 );
not \U$39411 ( \39390 , \39389 );
or \U$39412 ( \39391 , \39388 , \39390 );
buf \U$39413 ( \39392 , \36266 );
buf \U$39414 ( \39393 , \36252 );
or \U$39415 ( \39394 , \39392 , \39393 );
buf \U$39416 ( \39395 , \36240 );
not \U$39417 ( \39396 , \39395 );
buf \U$39418 ( \39397 , \39396 );
buf \U$39419 ( \39398 , \39397 );
nand \U$39420 ( \39399 , \39394 , \39398 );
buf \U$39421 ( \39400 , \39399 );
buf \U$39422 ( \39401 , \39400 );
nand \U$39423 ( \39402 , \39391 , \39401 );
buf \U$39424 ( \39403 , \39402 );
buf \U$39425 ( \39404 , \39403 );
xor \U$39426 ( \39405 , \39386 , \39404 );
xor \U$39427 ( \39406 , \38864 , \38870 );
and \U$39428 ( \39407 , \39406 , \38886 );
and \U$39429 ( \39408 , \38864 , \38870 );
or \U$39430 ( \39409 , \39407 , \39408 );
buf \U$39431 ( \39410 , \39409 );
buf \U$39432 ( \39411 , \39410 );
xnor \U$39433 ( \39412 , \39405 , \39411 );
buf \U$39434 ( \39413 , \39412 );
buf \U$39435 ( \39414 , \39413 );
not \U$39436 ( \39415 , \39414 );
or \U$39437 ( \39416 , \39368 , \39415 );
buf \U$39438 ( \39417 , \39413 );
buf \U$39439 ( \39418 , \39366 );
or \U$39440 ( \39419 , \39417 , \39418 );
nand \U$39441 ( \39420 , \39416 , \39419 );
buf \U$39442 ( \39421 , \39420 );
buf \U$39443 ( \39422 , \39421 );
not \U$39444 ( \39423 , \39422 );
or \U$39445 ( \39424 , \39361 , \39423 );
buf \U$39446 ( \39425 , \39421 );
buf \U$39447 ( \39426 , \39359 );
or \U$39448 ( \39427 , \39425 , \39426 );
nand \U$39449 ( \39428 , \39424 , \39427 );
buf \U$39450 ( \39429 , \39428 );
buf \U$39451 ( \39430 , \39429 );
xor \U$39452 ( \39431 , \39297 , \39430 );
buf \U$39453 ( \39432 , \39431 );
buf \U$39454 ( \39433 , \36277 );
not \U$39455 ( \39434 , \39433 );
buf \U$39456 ( \39435 , \39434 );
buf \U$39457 ( \39436 , \39435 );
not \U$39458 ( \39437 , \39436 );
buf \U$39459 ( \39438 , \36577 );
not \U$39460 ( \39439 , \39438 );
or \U$39461 ( \39440 , \39437 , \39439 );
buf \U$39462 ( \39441 , \36577 );
buf \U$39463 ( \39442 , \39435 );
or \U$39464 ( \39443 , \39441 , \39442 );
buf \U$39465 ( \39444 , \36444 );
nand \U$39466 ( \39445 , \39443 , \39444 );
buf \U$39467 ( \39446 , \39445 );
buf \U$39468 ( \39447 , \39446 );
nand \U$39469 ( \39448 , \39440 , \39447 );
buf \U$39470 ( \39449 , \39448 );
buf \U$39471 ( \39450 , \36573 );
buf \U$39472 ( \39451 , \36556 );
or \U$39473 ( \39452 , \39450 , \39451 );
buf \U$39474 ( \39453 , \36543 );
nand \U$39475 ( \39454 , \39452 , \39453 );
buf \U$39476 ( \39455 , \39454 );
buf \U$39477 ( \39456 , \39455 );
buf \U$39478 ( \39457 , \36573 );
buf \U$39479 ( \39458 , \36556 );
nand \U$39480 ( \39459 , \39457 , \39458 );
buf \U$39481 ( \39460 , \39459 );
buf \U$39482 ( \39461 , \39460 );
nand \U$39483 ( \39462 , \39456 , \39461 );
buf \U$39484 ( \39463 , \39462 );
buf \U$39485 ( \39464 , \39463 );
buf \U$39486 ( \39465 , \36875 );
not \U$39487 ( \39466 , \39465 );
buf \U$39488 ( \39467 , \36891 );
not \U$39489 ( \39468 , \39467 );
or \U$39490 ( \39469 , \39466 , \39468 );
buf \U$39491 ( \39470 , \36875 );
buf \U$39492 ( \39471 , \36891 );
or \U$39493 ( \39472 , \39470 , \39471 );
buf \U$39494 ( \39473 , \36905 );
nand \U$39495 ( \39474 , \39472 , \39473 );
buf \U$39496 ( \39475 , \39474 );
buf \U$39497 ( \39476 , \39475 );
nand \U$39498 ( \39477 , \39469 , \39476 );
buf \U$39499 ( \39478 , \39477 );
buf \U$39500 ( \39479 , \39478 );
xor \U$39501 ( \39480 , \39464 , \39479 );
xor \U$39502 ( \39481 , \36403 , \36417 );
and \U$39503 ( \39482 , \39481 , \36439 );
and \U$39504 ( \39483 , \36403 , \36417 );
or \U$39505 ( \39484 , \39482 , \39483 );
buf \U$39506 ( \39485 , \39484 );
buf \U$39507 ( \39486 , \39485 );
xor \U$39508 ( \39487 , \39480 , \39486 );
buf \U$39509 ( \39488 , \39487 );
and \U$39510 ( \39489 , \36487 , \36488 );
buf \U$39511 ( \39490 , \39489 );
buf \U$39512 ( \39491 , \39490 );
buf \U$39513 ( \39492 , \36521 );
not \U$39514 ( \39493 , \39492 );
buf \U$39515 ( \39494 , \1823 );
not \U$39516 ( \39495 , \39494 );
or \U$39517 ( \39496 , \39493 , \39495 );
buf \U$39518 ( \39497 , \686 );
buf \U$39519 ( \39498 , RIc0d8848_39);
buf \U$39520 ( \39499 , RIc0d9568_67);
xor \U$39521 ( \39500 , \39498 , \39499 );
buf \U$39522 ( \39501 , \39500 );
buf \U$39523 ( \39502 , \39501 );
nand \U$39524 ( \39503 , \39497 , \39502 );
buf \U$39525 ( \39504 , \39503 );
buf \U$39526 ( \39505 , \39504 );
nand \U$39527 ( \39506 , \39496 , \39505 );
buf \U$39528 ( \39507 , \39506 );
buf \U$39529 ( \39508 , \39507 );
xor \U$39530 ( \39509 , \39491 , \39508 );
buf \U$39531 ( \39510 , \36480 );
not \U$39532 ( \39511 , \39510 );
buf \U$39533 ( \39512 , \2535 );
not \U$39534 ( \39513 , \39512 );
or \U$39535 ( \39514 , \39511 , \39513 );
buf \U$39536 ( \39515 , \533 );
xor \U$39537 ( \39516 , RIc0da0a8_91, RIc0d7d08_15);
buf \U$39538 ( \39517 , \39516 );
nand \U$39539 ( \39518 , \39515 , \39517 );
buf \U$39540 ( \39519 , \39518 );
buf \U$39541 ( \39520 , \39519 );
nand \U$39542 ( \39521 , \39514 , \39520 );
buf \U$39543 ( \39522 , \39521 );
buf \U$39544 ( \39523 , \39522 );
xor \U$39545 ( \39524 , \39509 , \39523 );
buf \U$39546 ( \39525 , \39524 );
buf \U$39547 ( \39526 , \39525 );
buf \U$39548 ( \39527 , \36952 );
not \U$39549 ( \39528 , \39527 );
buf \U$39550 ( \39529 , \36923 );
not \U$39551 ( \39530 , \39529 );
or \U$39552 ( \39531 , \39528 , \39530 );
buf \U$39553 ( \39532 , \36923 );
buf \U$39554 ( \39533 , \36952 );
or \U$39555 ( \39534 , \39532 , \39533 );
buf \U$39556 ( \39535 , \36935 );
nand \U$39557 ( \39536 , \39534 , \39535 );
buf \U$39558 ( \39537 , \39536 );
buf \U$39559 ( \39538 , \39537 );
nand \U$39560 ( \39539 , \39531 , \39538 );
buf \U$39561 ( \39540 , \39539 );
buf \U$39562 ( \39541 , \39540 );
xor \U$39563 ( \39542 , \39526 , \39541 );
buf \U$39564 ( \39543 , \36500 );
not \U$39565 ( \39544 , \39543 );
buf \U$39566 ( \39545 , \12795 );
not \U$39567 ( \39546 , \39545 );
or \U$39568 ( \39547 , \39544 , \39546 );
buf \U$39569 ( \39548 , \1229 );
buf \U$39570 ( \39549 , RIc0d9478_65);
buf \U$39571 ( \39550 , RIc0d8938_41);
xor \U$39572 ( \39551 , \39549 , \39550 );
buf \U$39573 ( \39552 , \39551 );
buf \U$39574 ( \39553 , \39552 );
nand \U$39575 ( \39554 , \39548 , \39553 );
buf \U$39576 ( \39555 , \39554 );
buf \U$39577 ( \39556 , \39555 );
nand \U$39578 ( \39557 , \39547 , \39556 );
buf \U$39579 ( \39558 , \39557 );
buf \U$39580 ( \39559 , \39558 );
buf \U$39581 ( \39560 , \36342 );
not \U$39582 ( \39561 , \39560 );
buf \U$39583 ( \39562 , \2269 );
not \U$39584 ( \39563 , \39562 );
or \U$39585 ( \39564 , \39561 , \39563 );
buf \U$39586 ( \39565 , \18277 );
buf \U$39587 ( \39566 , RIc0d9748_71);
buf \U$39588 ( \39567 , RIc0d8668_35);
xor \U$39589 ( \39568 , \39566 , \39567 );
buf \U$39590 ( \39569 , \39568 );
buf \U$39591 ( \39570 , \39569 );
nand \U$39592 ( \39571 , \39565 , \39570 );
buf \U$39593 ( \39572 , \39571 );
buf \U$39594 ( \39573 , \39572 );
nand \U$39595 ( \39574 , \39564 , \39573 );
buf \U$39596 ( \39575 , \39574 );
buf \U$39597 ( \39576 , \39575 );
xor \U$39598 ( \39577 , \39559 , \39576 );
buf \U$39599 ( \39578 , \36378 );
not \U$39600 ( \39579 , \39578 );
buf \U$39601 ( \39580 , \29069 );
not \U$39602 ( \39581 , \39580 );
or \U$39603 ( \39582 , \39579 , \39581 );
buf \U$39604 ( \39583 , \734 );
buf \U$39605 ( \39584 , RIc0da378_97);
buf \U$39606 ( \39585 , RIc0d7a38_9);
and \U$39607 ( \39586 , \39584 , \39585 );
not \U$39608 ( \39587 , \39584 );
buf \U$39609 ( \39588 , \5976 );
and \U$39610 ( \39589 , \39587 , \39588 );
nor \U$39611 ( \39590 , \39586 , \39589 );
buf \U$39612 ( \39591 , \39590 );
buf \U$39613 ( \39592 , \39591 );
nand \U$39614 ( \39593 , \39583 , \39592 );
buf \U$39615 ( \39594 , \39593 );
buf \U$39616 ( \39595 , \39594 );
nand \U$39617 ( \39596 , \39582 , \39595 );
buf \U$39618 ( \39597 , \39596 );
buf \U$39619 ( \39598 , \39597 );
xor \U$39620 ( \39599 , \39577 , \39598 );
buf \U$39621 ( \39600 , \39599 );
buf \U$39622 ( \39601 , \39600 );
xor \U$39623 ( \39602 , \39542 , \39601 );
buf \U$39624 ( \39603 , \39602 );
xor \U$39625 ( \39604 , \39488 , \39603 );
buf \U$39626 ( \39605 , \36885 );
not \U$39627 ( \39606 , \39605 );
buf \U$39628 ( \39607 , \14532 );
not \U$39629 ( \39608 , \39607 );
or \U$39630 ( \39609 , \39606 , \39608 );
buf \U$39631 ( \39610 , \1078 );
buf \U$39632 ( \39611 , RIc0d9bf8_81);
buf \U$39633 ( \39612 , RIc0d81b8_25);
xor \U$39634 ( \39613 , \39611 , \39612 );
buf \U$39635 ( \39614 , \39613 );
buf \U$39636 ( \39615 , \39614 );
nand \U$39637 ( \39616 , \39610 , \39615 );
buf \U$39638 ( \39617 , \39616 );
buf \U$39639 ( \39618 , \39617 );
nand \U$39640 ( \39619 , \39609 , \39618 );
buf \U$39641 ( \39620 , \39619 );
buf \U$39642 ( \39621 , \39620 );
buf \U$39643 ( \39622 , \36396 );
not \U$39644 ( \39623 , \39622 );
buf \U$39645 ( \39624 , \3535 );
not \U$39646 ( \39625 , \39624 );
or \U$39647 ( \39626 , \39623 , \39625 );
buf \U$39648 ( \39627 , \16676 );
buf \U$39649 ( \39628 , RIc0d7858_5);
buf \U$39650 ( \39629 , RIc0da558_101);
xor \U$39651 ( \39630 , \39628 , \39629 );
buf \U$39652 ( \39631 , \39630 );
buf \U$39653 ( \39632 , \39631 );
nand \U$39654 ( \39633 , \39627 , \39632 );
buf \U$39655 ( \39634 , \39633 );
buf \U$39656 ( \39635 , \39634 );
nand \U$39657 ( \39636 , \39626 , \39635 );
buf \U$39658 ( \39637 , \39636 );
buf \U$39659 ( \39638 , \39637 );
xor \U$39660 ( \39639 , \39621 , \39638 );
buf \U$39661 ( \39640 , \36410 );
not \U$39662 ( \39641 , \39640 );
buf \U$39663 ( \39642 , \330 );
not \U$39664 ( \39643 , \39642 );
or \U$39665 ( \39644 , \39641 , \39643 );
buf \U$39666 ( \39645 , RIc0da288_95);
buf \U$39667 ( \39646 , RIc0d7b28_11);
xnor \U$39668 ( \39647 , \39645 , \39646 );
buf \U$39669 ( \39648 , \39647 );
buf \U$39670 ( \39649 , \39648 );
not \U$39671 ( \39650 , \39649 );
buf \U$39672 ( \39651 , \344 );
nand \U$39673 ( \39652 , \39650 , \39651 );
buf \U$39674 ( \39653 , \39652 );
buf \U$39675 ( \39654 , \39653 );
nand \U$39676 ( \39655 , \39644 , \39654 );
buf \U$39677 ( \39656 , \39655 );
buf \U$39678 ( \39657 , \39656 );
xor \U$39679 ( \39658 , \39639 , \39657 );
buf \U$39680 ( \39659 , \39658 );
buf \U$39681 ( \39660 , \36550 );
not \U$39682 ( \39661 , \39660 );
buf \U$39683 ( \39662 , \3384 );
not \U$39684 ( \39663 , \39662 );
or \U$39685 ( \39664 , \39661 , \39663 );
buf \U$39686 ( \39665 , \442 );
buf \U$39687 ( \39666 , RIc0d7df8_17);
buf \U$39688 ( \39667 , RIc0d9fb8_89);
xor \U$39689 ( \39668 , \39666 , \39667 );
buf \U$39690 ( \39669 , \39668 );
buf \U$39691 ( \39670 , \39669 );
nand \U$39692 ( \39671 , \39665 , \39670 );
buf \U$39693 ( \39672 , \39671 );
buf \U$39694 ( \39673 , \39672 );
nand \U$39695 ( \39674 , \39664 , \39673 );
buf \U$39696 ( \39675 , \39674 );
buf \U$39697 ( \39676 , \36300 );
not \U$39698 ( \39677 , \39676 );
buf \U$39699 ( \39678 , \13383 );
not \U$39700 ( \39679 , \39678 );
or \U$39701 ( \39680 , \39677 , \39679 );
buf \U$39702 ( \39681 , \1143 );
xor \U$39703 ( \39682 , RIc0d9928_75, RIc0d8488_31);
buf \U$39704 ( \39683 , \39682 );
nand \U$39705 ( \39684 , \39681 , \39683 );
buf \U$39706 ( \39685 , \39684 );
buf \U$39707 ( \39686 , \39685 );
nand \U$39708 ( \39687 , \39680 , \39686 );
buf \U$39709 ( \39688 , \39687 );
xor \U$39710 ( \39689 , \39675 , \39688 );
buf \U$39711 ( \39690 , \36899 );
not \U$39712 ( \39691 , \39690 );
buf \U$39713 ( \39692 , \1183 );
not \U$39714 ( \39693 , \39692 );
or \U$39715 ( \39694 , \39691 , \39693 );
buf \U$39716 ( \39695 , \6141 );
buf \U$39717 ( \39696 , RIc0d8398_29);
buf \U$39718 ( \39697 , RIc0d9a18_77);
xor \U$39719 ( \39698 , \39696 , \39697 );
buf \U$39720 ( \39699 , \39698 );
buf \U$39721 ( \39700 , \39699 );
nand \U$39722 ( \39701 , \39695 , \39700 );
buf \U$39723 ( \39702 , \39701 );
buf \U$39724 ( \39703 , \39702 );
nand \U$39725 ( \39704 , \39694 , \39703 );
buf \U$39726 ( \39705 , \39704 );
xor \U$39727 ( \39706 , \39689 , \39705 );
buf \U$39728 ( \39707 , \39706 );
not \U$39729 ( \39708 , \39707 );
buf \U$39730 ( \39709 , \39708 );
and \U$39731 ( \39710 , \39659 , \39709 );
not \U$39732 ( \39711 , \39659 );
and \U$39733 ( \39712 , \39711 , \39706 );
or \U$39734 ( \39713 , \39710 , \39712 );
buf \U$39735 ( \39714 , \39713 );
buf \U$39736 ( \39715 , \36286 );
not \U$39737 ( \39716 , \39715 );
buf \U$39738 ( \39717 , \951 );
not \U$39739 ( \39718 , \39717 );
or \U$39740 ( \39719 , \39716 , \39718 );
buf \U$39741 ( \39720 , \921 );
buf \U$39742 ( \39721 , RIc0d9dd8_85);
buf \U$39743 ( \39722 , RIc0d7fd8_21);
xor \U$39744 ( \39723 , \39721 , \39722 );
buf \U$39745 ( \39724 , \39723 );
buf \U$39746 ( \39725 , \39724 );
nand \U$39747 ( \39726 , \39720 , \39725 );
buf \U$39748 ( \39727 , \39726 );
buf \U$39749 ( \39728 , \39727 );
nand \U$39750 ( \39729 , \39719 , \39728 );
buf \U$39751 ( \39730 , \39729 );
buf \U$39752 ( \39731 , \39730 );
buf \U$39753 ( \39732 , \36567 );
not \U$39754 ( \39733 , \39732 );
buf \U$39755 ( \39734 , \1021 );
not \U$39756 ( \39735 , \39734 );
or \U$39757 ( \39736 , \39733 , \39735 );
buf \U$39758 ( \39737 , \1026 );
buf \U$39759 ( \39738 , RIc0d9b08_79);
buf \U$39760 ( \39739 , RIc0d82a8_27);
xor \U$39761 ( \39740 , \39738 , \39739 );
buf \U$39762 ( \39741 , \39740 );
buf \U$39763 ( \39742 , \39741 );
nand \U$39764 ( \39743 , \39737 , \39742 );
buf \U$39765 ( \39744 , \39743 );
buf \U$39766 ( \39745 , \39744 );
nand \U$39767 ( \39746 , \39736 , \39745 );
buf \U$39768 ( \39747 , \39746 );
buf \U$39769 ( \39748 , \39747 );
xor \U$39770 ( \39749 , \39731 , \39748 );
buf \U$39771 ( \39750 , \36537 );
not \U$39772 ( \39751 , \39750 );
buf \U$39773 ( \39752 , \1901 );
not \U$39774 ( \39753 , \39752 );
or \U$39775 ( \39754 , \39751 , \39753 );
buf \U$39776 ( \39755 , \4008 );
buf \U$39777 ( \39756 , RIc0d7c18_13);
buf \U$39778 ( \39757 , RIc0da198_93);
xor \U$39779 ( \39758 , \39756 , \39757 );
buf \U$39780 ( \39759 , \39758 );
buf \U$39781 ( \39760 , \39759 );
nand \U$39782 ( \39761 , \39755 , \39760 );
buf \U$39783 ( \39762 , \39761 );
buf \U$39784 ( \39763 , \39762 );
nand \U$39785 ( \39764 , \39754 , \39763 );
buf \U$39786 ( \39765 , \39764 );
buf \U$39787 ( \39766 , \39765 );
xor \U$39788 ( \39767 , \39749 , \39766 );
buf \U$39789 ( \39768 , \39767 );
buf \U$39790 ( \39769 , \39768 );
not \U$39791 ( \39770 , \39769 );
buf \U$39792 ( \39771 , \39770 );
buf \U$39793 ( \39772 , \39771 );
and \U$39794 ( \39773 , \39714 , \39772 );
not \U$39795 ( \39774 , \39714 );
buf \U$39796 ( \39775 , \39768 );
and \U$39797 ( \39776 , \39774 , \39775 );
nor \U$39798 ( \39777 , \39773 , \39776 );
buf \U$39799 ( \39778 , \39777 );
and \U$39800 ( \39779 , \39604 , \39778 );
not \U$39801 ( \39780 , \39604 );
buf \U$39802 ( \39781 , \39778 );
not \U$39803 ( \39782 , \39781 );
buf \U$39804 ( \39783 , \39782 );
and \U$39805 ( \39784 , \39780 , \39783 );
nor \U$39806 ( \39785 , \39779 , \39784 );
xor \U$39807 ( \39786 , \39449 , \39785 );
xor \U$39808 ( \39787 , \36859 , \36964 );
and \U$39809 ( \39788 , \39787 , \37347 );
and \U$39810 ( \39789 , \36859 , \36964 );
or \U$39811 ( \39790 , \39788 , \39789 );
buf \U$39812 ( \39791 , \39790 );
xor \U$39813 ( \39792 , \39786 , \39791 );
buf \U$39814 ( \39793 , \39792 );
not \U$39815 ( \39794 , \39793 );
buf \U$39816 ( \39795 , \36181 );
not \U$39817 ( \39796 , \39795 );
buf \U$39818 ( \39797 , \37349 );
not \U$39819 ( \39798 , \39797 );
or \U$39820 ( \39799 , \39796 , \39798 );
buf \U$39821 ( \39800 , \37349 );
buf \U$39822 ( \39801 , \36181 );
or \U$39823 ( \39802 , \39800 , \39801 );
buf \U$39824 ( \39803 , \36590 );
nand \U$39825 ( \39804 , \39802 , \39803 );
buf \U$39826 ( \39805 , \39804 );
buf \U$39827 ( \39806 , \39805 );
nand \U$39828 ( \39807 , \39799 , \39806 );
buf \U$39829 ( \39808 , \39807 );
buf \U$39830 ( \39809 , \39808 );
not \U$39831 ( \39810 , \39809 );
or \U$39832 ( \39811 , \39794 , \39810 );
buf \U$39833 ( \39812 , \39808 );
buf \U$39834 ( \39813 , \39792 );
or \U$39835 ( \39814 , \39812 , \39813 );
nand \U$39836 ( \39815 , \39811 , \39814 );
buf \U$39837 ( \39816 , \39815 );
buf \U$39838 ( \39817 , \39816 );
xor \U$39839 ( \39818 , \38789 , \38953 );
and \U$39840 ( \39819 , \39818 , \38960 );
and \U$39841 ( \39820 , \38789 , \38953 );
or \U$39842 ( \39821 , \39819 , \39820 );
buf \U$39843 ( \39822 , \39821 );
buf \U$39844 ( \39823 , \39822 );
not \U$39845 ( \39824 , \39823 );
buf \U$39846 ( \39825 , \39824 );
buf \U$39847 ( \39826 , \39825 );
and \U$39848 ( \39827 , \39817 , \39826 );
not \U$39849 ( \39828 , \39817 );
buf \U$39850 ( \39829 , \39822 );
and \U$39851 ( \39830 , \39828 , \39829 );
nor \U$39852 ( \39831 , \39827 , \39830 );
buf \U$39853 ( \39832 , \39831 );
xor \U$39854 ( \39833 , \39432 , \39832 );
buf \U$39855 ( \39834 , \38771 );
not \U$39856 ( \39835 , \39834 );
buf \U$39857 ( \39836 , \38227 );
not \U$39858 ( \39837 , \39836 );
buf \U$39859 ( \39838 , \37350 );
nand \U$39860 ( \39839 , \39837 , \39838 );
buf \U$39861 ( \39840 , \39839 );
buf \U$39862 ( \39841 , \39840 );
not \U$39863 ( \39842 , \39841 );
or \U$39864 ( \39843 , \39835 , \39842 );
buf \U$39865 ( \39844 , \37350 );
not \U$39866 ( \39845 , \39844 );
buf \U$39867 ( \39846 , \38227 );
nand \U$39868 ( \39847 , \39845 , \39846 );
buf \U$39869 ( \39848 , \39847 );
buf \U$39870 ( \39849 , \39848 );
nand \U$39871 ( \39850 , \39843 , \39849 );
buf \U$39872 ( \39851 , \39850 );
xor \U$39873 ( \39852 , \39833 , \39851 );
buf \U$39874 ( \39853 , \39852 );
nand \U$39875 ( \39854 , \39114 , \39853 );
buf \U$39876 ( \39855 , \39854 );
buf \U$39877 ( \39856 , \39855 );
xor \U$39878 ( \39857 , \38962 , \38779 );
xor \U$39879 ( \39858 , \39857 , \39099 );
buf \U$39880 ( \39859 , \39858 );
xor \U$39881 ( \39860 , \39086 , \39090 );
xor \U$39882 ( \39861 , \39860 , \39095 );
buf \U$39883 ( \39862 , \39861 );
buf \U$39884 ( \39863 , \39862 );
xor \U$39885 ( \39864 , \38241 , \38309 );
xor \U$39886 ( \39865 , \39864 , \38447 );
buf \U$39887 ( \39866 , \39865 );
buf \U$39888 ( \39867 , \39866 );
buf \U$39889 ( \39868 , \33911 );
not \U$39890 ( \39869 , \39868 );
buf \U$39891 ( \39870 , \33901 );
not \U$39892 ( \39871 , \39870 );
or \U$39893 ( \39872 , \39869 , \39871 );
buf \U$39894 ( \39873 , \33969 );
nand \U$39895 ( \39874 , \39872 , \39873 );
buf \U$39896 ( \39875 , \39874 );
buf \U$39897 ( \39876 , \39875 );
buf \U$39898 ( \39877 , \33907 );
buf \U$39899 ( \39878 , \33885 );
nand \U$39900 ( \39879 , \39877 , \39878 );
buf \U$39901 ( \39880 , \39879 );
buf \U$39902 ( \39881 , \39880 );
nand \U$39903 ( \39882 , \39876 , \39881 );
buf \U$39904 ( \39883 , \39882 );
buf \U$39905 ( \39884 , \39883 );
xor \U$39906 ( \39885 , \38316 , \38322 );
xor \U$39907 ( \39886 , \39885 , \38343 );
buf \U$39908 ( \39887 , \39886 );
buf \U$39909 ( \39888 , \39887 );
xor \U$39910 ( \39889 , \39884 , \39888 );
xor \U$39911 ( \39890 , \38351 , \38370 );
xor \U$39912 ( \39891 , \39890 , \38406 );
buf \U$39913 ( \39892 , \39891 );
buf \U$39914 ( \39893 , \39892 );
and \U$39915 ( \39894 , \39889 , \39893 );
and \U$39916 ( \39895 , \39884 , \39888 );
or \U$39917 ( \39896 , \39894 , \39895 );
buf \U$39918 ( \39897 , \39896 );
buf \U$39919 ( \39898 , \39897 );
xor \U$39920 ( \39899 , \38348 , \38411 );
xor \U$39921 ( \39900 , \39899 , \38442 );
buf \U$39922 ( \39901 , \39900 );
buf \U$39923 ( \39902 , \39901 );
xor \U$39924 ( \39903 , \39898 , \39902 );
xor \U$39925 ( \39904 , \38455 , \38470 );
xnor \U$39926 ( \39905 , \39904 , \38520 );
buf \U$39927 ( \39906 , \39905 );
and \U$39928 ( \39907 , \39903 , \39906 );
and \U$39929 ( \39908 , \39898 , \39902 );
or \U$39930 ( \39909 , \39907 , \39908 );
buf \U$39931 ( \39910 , \39909 );
buf \U$39932 ( \39911 , \39910 );
xor \U$39933 ( \39912 , \39867 , \39911 );
xor \U$39934 ( \39913 , \38529 , \38617 );
xor \U$39935 ( \39914 , \39913 , \38660 );
buf \U$39936 ( \39915 , \39914 );
buf \U$39937 ( \39916 , \39915 );
and \U$39938 ( \39917 , \39912 , \39916 );
and \U$39939 ( \39918 , \39867 , \39911 );
or \U$39940 ( \39919 , \39917 , \39918 );
buf \U$39941 ( \39920 , \39919 );
buf \U$39942 ( \39921 , \39920 );
or \U$39943 ( \39922 , \39863 , \39921 );
xor \U$39944 ( \39923 , \38987 , \38991 );
xor \U$39945 ( \39924 , \39923 , \39081 );
buf \U$39946 ( \39925 , \39924 );
buf \U$39947 ( \39926 , \39925 );
xor \U$39948 ( \39927 , \38588 , \38604 );
xor \U$39949 ( \39928 , \39927 , \38612 );
buf \U$39950 ( \39929 , \39928 );
buf \U$39951 ( \39930 , \39929 );
xor \U$39952 ( \39931 , \38417 , \38427 );
xor \U$39953 ( \39932 , \39931 , \38414 );
buf \U$39954 ( \39933 , \39932 );
not \U$39955 ( \39934 , \39933 );
buf \U$39956 ( \39935 , \34469 );
not \U$39957 ( \39936 , \39935 );
not \U$39958 ( \39937 , \34397 );
nand \U$39959 ( \39938 , \39937 , \34455 );
buf \U$39960 ( \39939 , \39938 );
not \U$39961 ( \39940 , \39939 );
or \U$39962 ( \39941 , \39936 , \39940 );
buf \U$39963 ( \39942 , \34455 );
not \U$39964 ( \39943 , \39942 );
buf \U$39965 ( \39944 , \34397 );
nand \U$39966 ( \39945 , \39943 , \39944 );
buf \U$39967 ( \39946 , \39945 );
buf \U$39968 ( \39947 , \39946 );
nand \U$39969 ( \39948 , \39941 , \39947 );
buf \U$39970 ( \39949 , \39948 );
buf \U$39971 ( \39950 , \39949 );
not \U$39972 ( \39951 , \39950 );
buf \U$39973 ( \39952 , \39951 );
buf \U$39974 ( \39953 , \39952 );
not \U$39975 ( \39954 , \39953 );
or \U$39976 ( \39955 , \39934 , \39954 );
buf \U$39977 ( \39956 , \38531 );
not \U$39978 ( \39957 , \39956 );
buf \U$39979 ( \39958 , \38581 );
not \U$39980 ( \39959 , \39958 );
or \U$39981 ( \39960 , \39957 , \39959 );
buf \U$39982 ( \39961 , \38531 );
buf \U$39983 ( \39962 , \38581 );
or \U$39984 ( \39963 , \39961 , \39962 );
nand \U$39985 ( \39964 , \39960 , \39963 );
buf \U$39986 ( \39965 , \39964 );
buf \U$39987 ( \39966 , \39965 );
buf \U$39988 ( \39967 , \38552 );
and \U$39989 ( \39968 , \39966 , \39967 );
not \U$39990 ( \39969 , \39966 );
buf \U$39991 ( \39970 , \38560 );
and \U$39992 ( \39971 , \39969 , \39970 );
nor \U$39993 ( \39972 , \39968 , \39971 );
buf \U$39994 ( \39973 , \39972 );
buf \U$39995 ( \39974 , \39973 );
nand \U$39996 ( \39975 , \39955 , \39974 );
buf \U$39997 ( \39976 , \39975 );
buf \U$39998 ( \39977 , \39976 );
buf \U$39999 ( \39978 , \39932 );
not \U$40000 ( \39979 , \39978 );
buf \U$40001 ( \39980 , \39979 );
buf \U$40002 ( \39981 , \39980 );
buf \U$40003 ( \39982 , \39949 );
nand \U$40004 ( \39983 , \39981 , \39982 );
buf \U$40005 ( \39984 , \39983 );
buf \U$40006 ( \39985 , \39984 );
and \U$40007 ( \39986 , \39977 , \39985 );
buf \U$40008 ( \39987 , \39986 );
buf \U$40009 ( \39988 , \39987 );
not \U$40010 ( \39989 , \39988 );
buf \U$40011 ( \39990 , \39989 );
buf \U$40012 ( \39991 , \39990 );
or \U$40013 ( \39992 , \39930 , \39991 );
buf \U$40014 ( \39993 , \39992 );
buf \U$40015 ( \39994 , \39993 );
not \U$40016 ( \39995 , \39994 );
buf \U$40017 ( \39996 , \33812 );
not \U$40018 ( \39997 , \39996 );
buf \U$40019 ( \39998 , \33852 );
not \U$40020 ( \39999 , \39998 );
or \U$40021 ( \40000 , \39997 , \39999 );
buf \U$40022 ( \40001 , \33812 );
not \U$40023 ( \40002 , \40001 );
buf \U$40024 ( \40003 , \33849 );
nand \U$40025 ( \40004 , \40002 , \40003 );
buf \U$40026 ( \40005 , \40004 );
buf \U$40027 ( \40006 , \40005 );
buf \U$40028 ( \40007 , \33870 );
nand \U$40029 ( \40008 , \40006 , \40007 );
buf \U$40030 ( \40009 , \40008 );
buf \U$40031 ( \40010 , \40009 );
nand \U$40032 ( \40011 , \40000 , \40010 );
buf \U$40033 ( \40012 , \40011 );
buf \U$40034 ( \40013 , \40012 );
not \U$40035 ( \40014 , \40013 );
buf \U$40036 ( \40015 , \40014 );
buf \U$40037 ( \40016 , \40015 );
not \U$40038 ( \40017 , \40016 );
xor \U$40039 ( \40018 , \39003 , \39018 );
xor \U$40040 ( \40019 , \40018 , \39023 );
buf \U$40041 ( \40020 , \40019 );
buf \U$40042 ( \40021 , \40020 );
not \U$40043 ( \40022 , \40021 );
buf \U$40044 ( \40023 , \40022 );
buf \U$40045 ( \40024 , \40023 );
not \U$40046 ( \40025 , \40024 );
or \U$40047 ( \40026 , \40017 , \40025 );
buf \U$40048 ( \40027 , \33665 );
not \U$40049 ( \40028 , \40027 );
buf \U$40050 ( \40029 , \33742 );
not \U$40051 ( \40030 , \40029 );
buf \U$40052 ( \40031 , \40030 );
buf \U$40053 ( \40032 , \40031 );
not \U$40054 ( \40033 , \40032 );
or \U$40055 ( \40034 , \40028 , \40033 );
buf \U$40056 ( \40035 , \33665 );
not \U$40057 ( \40036 , \40035 );
buf \U$40058 ( \40037 , \40036 );
buf \U$40059 ( \40038 , \40037 );
not \U$40060 ( \40039 , \40038 );
buf \U$40061 ( \40040 , \33742 );
not \U$40062 ( \40041 , \40040 );
or \U$40063 ( \40042 , \40039 , \40041 );
buf \U$40064 ( \40043 , \33679 );
nand \U$40065 ( \40044 , \40042 , \40043 );
buf \U$40066 ( \40045 , \40044 );
buf \U$40067 ( \40046 , \40045 );
nand \U$40068 ( \40047 , \40034 , \40046 );
buf \U$40069 ( \40048 , \40047 );
buf \U$40070 ( \40049 , \40048 );
nand \U$40071 ( \40050 , \40026 , \40049 );
buf \U$40072 ( \40051 , \40050 );
buf \U$40073 ( \40052 , \40051 );
buf \U$40074 ( \40053 , \40020 );
buf \U$40075 ( \40054 , \40012 );
nand \U$40076 ( \40055 , \40053 , \40054 );
buf \U$40077 ( \40056 , \40055 );
buf \U$40078 ( \40057 , \40056 );
nand \U$40079 ( \40058 , \40052 , \40057 );
buf \U$40080 ( \40059 , \40058 );
buf \U$40081 ( \40060 , \40059 );
not \U$40082 ( \40061 , \40060 );
or \U$40083 ( \40062 , \39995 , \40061 );
buf \U$40084 ( \40063 , \39929 );
buf \U$40085 ( \40064 , \39990 );
nand \U$40086 ( \40065 , \40063 , \40064 );
buf \U$40087 ( \40066 , \40065 );
buf \U$40088 ( \40067 , \40066 );
nand \U$40089 ( \40068 , \40062 , \40067 );
buf \U$40090 ( \40069 , \40068 );
buf \U$40091 ( \40070 , \40069 );
xor \U$40092 ( \40071 , \39926 , \40070 );
xor \U$40093 ( \40072 , \39048 , \39066 );
xor \U$40094 ( \40073 , \40072 , \39071 );
buf \U$40095 ( \40074 , \40073 );
buf \U$40096 ( \40075 , \40074 );
xor \U$40097 ( \40076 , \39884 , \39888 );
xor \U$40098 ( \40077 , \40076 , \39893 );
buf \U$40099 ( \40078 , \40077 );
buf \U$40100 ( \40079 , \40078 );
or \U$40101 ( \40080 , \40075 , \40079 );
buf \U$40102 ( \40081 , \33979 );
not \U$40103 ( \40082 , \40081 );
buf \U$40104 ( \40083 , \40082 );
buf \U$40105 ( \40084 , \40083 );
not \U$40106 ( \40085 , \40084 );
buf \U$40107 ( \40086 , \34127 );
not \U$40108 ( \40087 , \40086 );
or \U$40109 ( \40088 , \40085 , \40087 );
buf \U$40110 ( \40089 , \34127 );
buf \U$40111 ( \40090 , \40083 );
or \U$40112 ( \40091 , \40089 , \40090 );
buf \U$40113 ( \40092 , \33880 );
nand \U$40114 ( \40093 , \40091 , \40092 );
buf \U$40115 ( \40094 , \40093 );
buf \U$40116 ( \40095 , \40094 );
nand \U$40117 ( \40096 , \40088 , \40095 );
buf \U$40118 ( \40097 , \40096 );
buf \U$40119 ( \40098 , \40097 );
nand \U$40120 ( \40099 , \40080 , \40098 );
buf \U$40121 ( \40100 , \40099 );
buf \U$40122 ( \40101 , \40100 );
buf \U$40123 ( \40102 , \40074 );
buf \U$40124 ( \40103 , \40078 );
nand \U$40125 ( \40104 , \40102 , \40103 );
buf \U$40126 ( \40105 , \40104 );
buf \U$40127 ( \40106 , \40105 );
nand \U$40128 ( \40107 , \40101 , \40106 );
buf \U$40129 ( \40108 , \40107 );
buf \U$40130 ( \40109 , \40108 );
xor \U$40131 ( \40110 , \39028 , \39032 );
xor \U$40132 ( \40111 , \40110 , \39076 );
buf \U$40133 ( \40112 , \40111 );
buf \U$40134 ( \40113 , \40112 );
xor \U$40135 ( \40114 , \40109 , \40113 );
xor \U$40136 ( \40115 , \39898 , \39902 );
xor \U$40137 ( \40116 , \40115 , \39906 );
buf \U$40138 ( \40117 , \40116 );
buf \U$40139 ( \40118 , \40117 );
and \U$40140 ( \40119 , \40114 , \40118 );
and \U$40141 ( \40120 , \40109 , \40113 );
or \U$40142 ( \40121 , \40119 , \40120 );
buf \U$40143 ( \40122 , \40121 );
buf \U$40144 ( \40123 , \40122 );
and \U$40145 ( \40124 , \40071 , \40123 );
and \U$40146 ( \40125 , \39926 , \40070 );
or \U$40147 ( \40126 , \40124 , \40125 );
buf \U$40148 ( \40127 , \40126 );
buf \U$40149 ( \40128 , \40127 );
nand \U$40150 ( \40129 , \39922 , \40128 );
buf \U$40151 ( \40130 , \40129 );
buf \U$40152 ( \40131 , \40130 );
buf \U$40153 ( \40132 , \39862 );
buf \U$40154 ( \40133 , \39920 );
nand \U$40155 ( \40134 , \40132 , \40133 );
buf \U$40156 ( \40135 , \40134 );
buf \U$40157 ( \40136 , \40135 );
nand \U$40158 ( \40137 , \40131 , \40136 );
buf \U$40159 ( \40138 , \40137 );
buf \U$40160 ( \40139 , \40138 );
not \U$40161 ( \40140 , \40139 );
buf \U$40162 ( \40141 , \40140 );
buf \U$40163 ( \40142 , \40141 );
nand \U$40164 ( \40143 , \39859 , \40142 );
buf \U$40165 ( \40144 , \40143 );
buf \U$40166 ( \40145 , \40144 );
nand \U$40167 ( \40146 , \39856 , \40145 );
buf \U$40168 ( \40147 , \40146 );
buf \U$40169 ( \40148 , \40147 );
buf \U$40170 ( \40149 , RIc0d8320_28);
buf \U$40171 ( \40150 , RIc0d9a18_77);
xor \U$40172 ( \40151 , \40149 , \40150 );
buf \U$40173 ( \40152 , \40151 );
buf \U$40174 ( \40153 , \40152 );
not \U$40175 ( \40154 , \40153 );
buf \U$40176 ( \40155 , \1431 );
not \U$40177 ( \40156 , \40155 );
or \U$40178 ( \40157 , \40154 , \40156 );
buf \U$40179 ( \40158 , RIc0d9a18_77);
buf \U$40180 ( \40159 , RIc0d82a8_27);
xnor \U$40181 ( \40160 , \40158 , \40159 );
buf \U$40182 ( \40161 , \40160 );
buf \U$40183 ( \40162 , \40161 );
not \U$40184 ( \40163 , \40162 );
buf \U$40185 ( \40164 , \14374 );
nand \U$40186 ( \40165 , \40163 , \40164 );
buf \U$40187 ( \40166 , \40165 );
buf \U$40188 ( \40167 , \40166 );
nand \U$40189 ( \40168 , \40157 , \40167 );
buf \U$40190 ( \40169 , \40168 );
xor \U$40191 ( \40170 , RIc0d9928_75, RIc0d8410_30);
buf \U$40192 ( \40171 , \40170 );
not \U$40193 ( \40172 , \40171 );
buf \U$40194 ( \40173 , \2358 );
not \U$40195 ( \40174 , \40173 );
or \U$40196 ( \40175 , \40172 , \40174 );
buf \U$40197 ( \40176 , \16500 );
buf \U$40198 ( \40177 , RIc0d9928_75);
buf \U$40199 ( \40178 , RIc0d8398_29);
xor \U$40200 ( \40179 , \40177 , \40178 );
buf \U$40201 ( \40180 , \40179 );
buf \U$40202 ( \40181 , \40180 );
nand \U$40203 ( \40182 , \40176 , \40181 );
buf \U$40204 ( \40183 , \40182 );
buf \U$40205 ( \40184 , \40183 );
nand \U$40206 ( \40185 , \40175 , \40184 );
buf \U$40207 ( \40186 , \40185 );
xor \U$40208 ( \40187 , \40169 , \40186 );
buf \U$40209 ( \40188 , RIc0da558_101);
buf \U$40210 ( \40189 , RIc0d77e0_4);
and \U$40211 ( \40190 , \40188 , \40189 );
not \U$40212 ( \40191 , \40188 );
buf \U$40213 ( \40192 , \489 );
and \U$40214 ( \40193 , \40191 , \40192 );
nor \U$40215 ( \40194 , \40190 , \40193 );
buf \U$40216 ( \40195 , \40194 );
buf \U$40217 ( \40196 , \40195 );
not \U$40218 ( \40197 , \40196 );
buf \U$40219 ( \40198 , \4043 );
not \U$40220 ( \40199 , \40198 );
or \U$40221 ( \40200 , \40197 , \40199 );
buf \U$40222 ( \40201 , RIc0d7768_3);
buf \U$40223 ( \40202 , RIc0da558_101);
xnor \U$40224 ( \40203 , \40201 , \40202 );
buf \U$40225 ( \40204 , \40203 );
buf \U$40226 ( \40205 , \40204 );
not \U$40227 ( \40206 , \40205 );
buf \U$40228 ( \40207 , \26354 );
nand \U$40229 ( \40208 , \40206 , \40207 );
buf \U$40230 ( \40209 , \40208 );
buf \U$40231 ( \40210 , \40209 );
nand \U$40232 ( \40211 , \40200 , \40210 );
buf \U$40233 ( \40212 , \40211 );
not \U$40234 ( \40213 , \40212 );
xor \U$40235 ( \40214 , \40187 , \40213 );
buf \U$40236 ( \40215 , \40214 );
not \U$40237 ( \40216 , \40215 );
buf \U$40238 ( \40217 , \40216 );
buf \U$40239 ( \40218 , \40217 );
and \U$40240 ( \40219 , \39549 , \39550 );
buf \U$40241 ( \40220 , \40219 );
buf \U$40242 ( \40221 , \40220 );
xor \U$40243 ( \40222 , RIc0d9568_67, RIc0d87d0_38);
buf \U$40244 ( \40223 , \40222 );
not \U$40245 ( \40224 , \40223 );
buf \U$40246 ( \40225 , \1414 );
not \U$40247 ( \40226 , \40225 );
or \U$40248 ( \40227 , \40224 , \40226 );
buf \U$40249 ( \40228 , \686 );
buf \U$40250 ( \40229 , RIc0d9568_67);
buf \U$40251 ( \40230 , RIc0d8758_37);
xor \U$40252 ( \40231 , \40229 , \40230 );
buf \U$40253 ( \40232 , \40231 );
buf \U$40254 ( \40233 , \40232 );
nand \U$40255 ( \40234 , \40228 , \40233 );
buf \U$40256 ( \40235 , \40234 );
buf \U$40257 ( \40236 , \40235 );
nand \U$40258 ( \40237 , \40227 , \40236 );
buf \U$40259 ( \40238 , \40237 );
buf \U$40260 ( \40239 , \40238 );
xor \U$40261 ( \40240 , \40221 , \40239 );
buf \U$40262 ( \40241 , RIc0da0a8_91);
buf \U$40263 ( \40242 , RIc0d7c90_14);
and \U$40264 ( \40243 , \40241 , \40242 );
not \U$40265 ( \40244 , \40241 );
buf \U$40266 ( \40245 , RIc0d7c90_14);
not \U$40267 ( \40246 , \40245 );
buf \U$40268 ( \40247 , \40246 );
buf \U$40269 ( \40248 , \40247 );
and \U$40270 ( \40249 , \40244 , \40248 );
nor \U$40271 ( \40250 , \40243 , \40249 );
buf \U$40272 ( \40251 , \40250 );
buf \U$40273 ( \40252 , \40251 );
not \U$40274 ( \40253 , \40252 );
buf \U$40275 ( \40254 , \2535 );
not \U$40276 ( \40255 , \40254 );
or \U$40277 ( \40256 , \40253 , \40255 );
buf \U$40278 ( \40257 , RIc0da0a8_91);
buf \U$40279 ( \40258 , RIc0d7c18_13);
xnor \U$40280 ( \40259 , \40257 , \40258 );
buf \U$40281 ( \40260 , \40259 );
buf \U$40282 ( \40261 , \40260 );
not \U$40283 ( \40262 , \40261 );
buf \U$40284 ( \40263 , \1933 );
nand \U$40285 ( \40264 , \40262 , \40263 );
buf \U$40286 ( \40265 , \40264 );
buf \U$40287 ( \40266 , \40265 );
nand \U$40288 ( \40267 , \40256 , \40266 );
buf \U$40289 ( \40268 , \40267 );
buf \U$40290 ( \40269 , \40268 );
xnor \U$40291 ( \40270 , \40240 , \40269 );
buf \U$40292 ( \40271 , \40270 );
buf \U$40293 ( \40272 , \40271 );
not \U$40294 ( \40273 , \40272 );
buf \U$40295 ( \40274 , \40273 );
buf \U$40296 ( \40275 , \40274 );
and \U$40297 ( \40276 , \40218 , \40275 );
not \U$40298 ( \40277 , \40218 );
buf \U$40299 ( \40278 , \40271 );
and \U$40300 ( \40279 , \40277 , \40278 );
nor \U$40301 ( \40280 , \40276 , \40279 );
buf \U$40302 ( \40281 , \40280 );
buf \U$40303 ( \40282 , \40281 );
buf \U$40304 ( \40283 , RIc0d8500_32);
buf \U$40305 ( \40284 , RIc0d9838_73);
xor \U$40306 ( \40285 , \40283 , \40284 );
buf \U$40307 ( \40286 , \40285 );
buf \U$40308 ( \40287 , \40286 );
not \U$40309 ( \40288 , \40287 );
buf \U$40310 ( \40289 , \1677 );
not \U$40311 ( \40290 , \40289 );
or \U$40312 ( \40291 , \40288 , \40290 );
buf \U$40313 ( \40292 , \1856 );
buf \U$40314 ( \40293 , RIc0d8488_31);
buf \U$40315 ( \40294 , RIc0d9838_73);
xor \U$40316 ( \40295 , \40293 , \40294 );
buf \U$40317 ( \40296 , \40295 );
buf \U$40318 ( \40297 , \40296 );
nand \U$40319 ( \40298 , \40292 , \40297 );
buf \U$40320 ( \40299 , \40298 );
buf \U$40321 ( \40300 , \40299 );
nand \U$40322 ( \40301 , \40291 , \40300 );
buf \U$40323 ( \40302 , \40301 );
buf \U$40324 ( \40303 , \40302 );
buf \U$40325 ( \40304 , RIc0d9b08_79);
buf \U$40326 ( \40305 , RIc0d8230_26);
xor \U$40327 ( \40306 , \40304 , \40305 );
buf \U$40328 ( \40307 , \40306 );
buf \U$40329 ( \40308 , \40307 );
not \U$40330 ( \40309 , \40308 );
buf \U$40331 ( \40310 , \1021 );
not \U$40332 ( \40311 , \40310 );
or \U$40333 ( \40312 , \40309 , \40311 );
buf \U$40334 ( \40313 , RIc0d9b08_79);
buf \U$40335 ( \40314 , RIc0d81b8_25);
xnor \U$40336 ( \40315 , \40313 , \40314 );
buf \U$40337 ( \40316 , \40315 );
buf \U$40338 ( \40317 , \40316 );
not \U$40339 ( \40318 , \40317 );
buf \U$40340 ( \40319 , \1025 );
nand \U$40341 ( \40320 , \40318 , \40319 );
buf \U$40342 ( \40321 , \40320 );
buf \U$40343 ( \40322 , \40321 );
nand \U$40344 ( \40323 , \40312 , \40322 );
buf \U$40345 ( \40324 , \40323 );
buf \U$40346 ( \40325 , \40324 );
xor \U$40347 ( \40326 , \40303 , \40325 );
buf \U$40348 ( \40327 , \473 );
buf \U$40349 ( \40328 , RIc0d7ba0_12);
buf \U$40350 ( \40329 , RIc0da198_93);
xor \U$40351 ( \40330 , \40328 , \40329 );
buf \U$40352 ( \40331 , \40330 );
buf \U$40353 ( \40332 , \40331 );
not \U$40354 ( \40333 , \40332 );
buf \U$40355 ( \40334 , \40333 );
buf \U$40356 ( \40335 , \40334 );
or \U$40357 ( \40336 , \40327 , \40335 );
buf \U$40358 ( \40337 , \481 );
not \U$40359 ( \40338 , \40337 );
buf \U$40360 ( \40339 , \40338 );
buf \U$40361 ( \40340 , \40339 );
buf \U$40362 ( \40341 , RIc0da198_93);
buf \U$40363 ( \40342 , RIc0d7b28_11);
xor \U$40364 ( \40343 , \40341 , \40342 );
buf \U$40365 ( \40344 , \40343 );
buf \U$40366 ( \40345 , \40344 );
not \U$40367 ( \40346 , \40345 );
buf \U$40368 ( \40347 , \40346 );
buf \U$40369 ( \40348 , \40347 );
or \U$40370 ( \40349 , \40340 , \40348 );
nand \U$40371 ( \40350 , \40336 , \40349 );
buf \U$40372 ( \40351 , \40350 );
buf \U$40373 ( \40352 , \40351 );
xor \U$40374 ( \40353 , \40326 , \40352 );
buf \U$40375 ( \40354 , \40353 );
buf \U$40376 ( \40355 , \40354 );
xor \U$40377 ( \40356 , \40282 , \40355 );
buf \U$40378 ( \40357 , \40356 );
buf \U$40379 ( \40358 , \40357 );
buf \U$40380 ( \40359 , RIc0d9748_71);
buf \U$40381 ( \40360 , RIc0d85f0_34);
xor \U$40382 ( \40361 , \40359 , \40360 );
buf \U$40383 ( \40362 , \40361 );
buf \U$40384 ( \40363 , \40362 );
not \U$40385 ( \40364 , \40363 );
buf \U$40386 ( \40365 , \2812 );
not \U$40387 ( \40366 , \40365 );
or \U$40388 ( \40367 , \40364 , \40366 );
buf \U$40389 ( \40368 , \1282 );
buf \U$40390 ( \40369 , RIc0d8578_33);
buf \U$40391 ( \40370 , RIc0d9748_71);
xor \U$40392 ( \40371 , \40369 , \40370 );
buf \U$40393 ( \40372 , \40371 );
buf \U$40394 ( \40373 , \40372 );
nand \U$40395 ( \40374 , \40368 , \40373 );
buf \U$40396 ( \40375 , \40374 );
buf \U$40397 ( \40376 , \40375 );
nand \U$40398 ( \40377 , \40367 , \40376 );
buf \U$40399 ( \40378 , \40377 );
buf \U$40400 ( \40379 , \40378 );
not \U$40401 ( \40380 , \40379 );
buf \U$40402 ( \40381 , \40380 );
buf \U$40403 ( \40382 , RIc0d9478_65);
buf \U$40404 ( \40383 , RIc0d88c0_40);
xor \U$40405 ( \40384 , \40382 , \40383 );
buf \U$40406 ( \40385 , \40384 );
buf \U$40407 ( \40386 , \40385 );
not \U$40408 ( \40387 , \40386 );
buf \U$40409 ( \40388 , \1224 );
not \U$40410 ( \40389 , \40388 );
or \U$40411 ( \40390 , \40387 , \40389 );
buf \U$40412 ( \40391 , \1229 );
xor \U$40413 ( \40392 , \4379 , \4380 );
buf \U$40414 ( \40393 , \40392 );
buf \U$40415 ( \40394 , \40393 );
nand \U$40416 ( \40395 , \40391 , \40394 );
buf \U$40417 ( \40396 , \40395 );
buf \U$40418 ( \40397 , \40396 );
nand \U$40419 ( \40398 , \40390 , \40397 );
buf \U$40420 ( \40399 , \40398 );
buf \U$40421 ( \40400 , \40399 );
not \U$40422 ( \40401 , \40400 );
buf \U$40423 ( \40402 , \40401 );
xor \U$40424 ( \40403 , \40381 , \40402 );
buf \U$40425 ( \40404 , RIc0d79c0_8);
buf \U$40426 ( \40405 , RIc0da378_97);
xor \U$40427 ( \40406 , \40404 , \40405 );
buf \U$40428 ( \40407 , \40406 );
buf \U$40429 ( \40408 , \40407 );
not \U$40430 ( \40409 , \40408 );
buf \U$40431 ( \40410 , \16358 );
not \U$40432 ( \40411 , \40410 );
or \U$40433 ( \40412 , \40409 , \40411 );
buf \U$40434 ( \40413 , \734 );
buf \U$40435 ( \40414 , RIc0d7948_7);
buf \U$40436 ( \40415 , RIc0da378_97);
xor \U$40437 ( \40416 , \40414 , \40415 );
buf \U$40438 ( \40417 , \40416 );
buf \U$40439 ( \40418 , \40417 );
nand \U$40440 ( \40419 , \40413 , \40418 );
buf \U$40441 ( \40420 , \40419 );
buf \U$40442 ( \40421 , \40420 );
nand \U$40443 ( \40422 , \40412 , \40421 );
buf \U$40444 ( \40423 , \40422 );
xor \U$40445 ( \40424 , \40403 , \40423 );
buf \U$40446 ( \40425 , \40424 );
buf \U$40447 ( \40426 , RIc0d7d80_16);
buf \U$40448 ( \40427 , RIc0d9fb8_89);
xor \U$40449 ( \40428 , \40426 , \40427 );
buf \U$40450 ( \40429 , \40428 );
buf \U$40451 ( \40430 , \40429 );
not \U$40452 ( \40431 , \40430 );
buf \U$40453 ( \40432 , \2038 );
not \U$40454 ( \40433 , \40432 );
or \U$40455 ( \40434 , \40431 , \40433 );
buf \U$40456 ( \40435 , RIc0d9fb8_89);
buf \U$40457 ( \40436 , RIc0d7d08_15);
xnor \U$40458 ( \40437 , \40435 , \40436 );
buf \U$40459 ( \40438 , \40437 );
buf \U$40460 ( \40439 , \40438 );
not \U$40461 ( \40440 , \40439 );
buf \U$40462 ( \40441 , \846 );
nand \U$40463 ( \40442 , \40440 , \40441 );
buf \U$40464 ( \40443 , \40442 );
buf \U$40465 ( \40444 , \40443 );
nand \U$40466 ( \40445 , \40434 , \40444 );
buf \U$40467 ( \40446 , \40445 );
buf \U$40468 ( \40447 , \40446 );
buf \U$40469 ( \40448 , RIc0d9ec8_87);
buf \U$40470 ( \40449 , RIc0d7e70_18);
and \U$40471 ( \40450 , \40448 , \40449 );
not \U$40472 ( \40451 , \40448 );
buf \U$40473 ( \40452 , \7820 );
and \U$40474 ( \40453 , \40451 , \40452 );
nor \U$40475 ( \40454 , \40450 , \40453 );
buf \U$40476 ( \40455 , \40454 );
buf \U$40477 ( \40456 , \40455 );
not \U$40478 ( \40457 , \40456 );
buf \U$40479 ( \40458 , \4527 );
not \U$40480 ( \40459 , \40458 );
or \U$40481 ( \40460 , \40457 , \40459 );
buf \U$40482 ( \40461 , RIc0d7df8_17);
buf \U$40483 ( \40462 , RIc0d9ec8_87);
xnor \U$40484 ( \40463 , \40461 , \40462 );
buf \U$40485 ( \40464 , \40463 );
buf \U$40486 ( \40465 , \40464 );
not \U$40487 ( \40466 , \40465 );
buf \U$40488 ( \40467 , \3631 );
nand \U$40489 ( \40468 , \40466 , \40467 );
buf \U$40490 ( \40469 , \40468 );
buf \U$40491 ( \40470 , \40469 );
nand \U$40492 ( \40471 , \40460 , \40470 );
buf \U$40493 ( \40472 , \40471 );
buf \U$40494 ( \40473 , \40472 );
xor \U$40495 ( \40474 , \40447 , \40473 );
buf \U$40496 ( \40475 , \25374 );
buf \U$40497 ( \40476 , RIc0da468_99);
buf \U$40498 ( \40477 , RIc0d78d0_6);
xnor \U$40499 ( \40478 , \40476 , \40477 );
buf \U$40500 ( \40479 , \40478 );
buf \U$40501 ( \40480 , \40479 );
or \U$40502 ( \40481 , \40475 , \40480 );
buf \U$40503 ( \40482 , \2198 );
buf \U$40504 ( \40483 , RIc0da468_99);
buf \U$40505 ( \40484 , RIc0d7858_5);
and \U$40506 ( \40485 , \40483 , \40484 );
not \U$40507 ( \40486 , \40483 );
buf \U$40508 ( \40487 , \1990 );
and \U$40509 ( \40488 , \40486 , \40487 );
nor \U$40510 ( \40489 , \40485 , \40488 );
buf \U$40511 ( \40490 , \40489 );
buf \U$40512 ( \40491 , \40490 );
not \U$40513 ( \40492 , \40491 );
buf \U$40514 ( \40493 , \40492 );
buf \U$40515 ( \40494 , \40493 );
or \U$40516 ( \40495 , \40482 , \40494 );
nand \U$40517 ( \40496 , \40481 , \40495 );
buf \U$40518 ( \40497 , \40496 );
buf \U$40519 ( \40498 , \40497 );
xor \U$40520 ( \40499 , \40474 , \40498 );
buf \U$40521 ( \40500 , \40499 );
buf \U$40522 ( \40501 , \40500 );
xor \U$40523 ( \40502 , \40425 , \40501 );
buf \U$40524 ( \40503 , \2769 );
buf \U$40525 ( \40504 , RIc0d8140_24);
buf \U$40526 ( \40505 , RIc0d9bf8_81);
xnor \U$40527 ( \40506 , \40504 , \40505 );
buf \U$40528 ( \40507 , \40506 );
buf \U$40529 ( \40508 , \40507 );
or \U$40530 ( \40509 , \40503 , \40508 );
buf \U$40531 ( \40510 , \2775 );
buf \U$40532 ( \40511 , RIc0d80c8_23);
buf \U$40533 ( \40512 , RIc0d9bf8_81);
xnor \U$40534 ( \40513 , \40511 , \40512 );
buf \U$40535 ( \40514 , \40513 );
buf \U$40536 ( \40515 , \40514 );
or \U$40537 ( \40516 , \40510 , \40515 );
nand \U$40538 ( \40517 , \40509 , \40516 );
buf \U$40539 ( \40518 , \40517 );
buf \U$40540 ( \40519 , \40518 );
buf \U$40541 ( \40520 , \17405 );
not \U$40542 ( \40521 , \40520 );
buf \U$40543 ( \40522 , \40521 );
buf \U$40544 ( \40523 , \40522 );
buf \U$40545 ( \40524 , RIc0da648_103);
buf \U$40546 ( \40525 , RIc0d76f0_2);
xnor \U$40547 ( \40526 , \40524 , \40525 );
buf \U$40548 ( \40527 , \40526 );
buf \U$40549 ( \40528 , \40527 );
or \U$40550 ( \40529 , \40523 , \40528 );
buf \U$40551 ( \40530 , \4475 );
buf \U$40552 ( \40531 , RIc0da648_103);
buf \U$40553 ( \40532 , RIc0d7678_1);
and \U$40554 ( \40533 , \40531 , \40532 );
not \U$40555 ( \40534 , \40531 );
buf \U$40556 ( \40535 , \974 );
and \U$40557 ( \40536 , \40534 , \40535 );
nor \U$40558 ( \40537 , \40533 , \40536 );
buf \U$40559 ( \40538 , \40537 );
buf \U$40560 ( \40539 , \40538 );
not \U$40561 ( \40540 , \40539 );
buf \U$40562 ( \40541 , \40540 );
buf \U$40563 ( \40542 , \40541 );
or \U$40564 ( \40543 , \40530 , \40542 );
nand \U$40565 ( \40544 , \40529 , \40543 );
buf \U$40566 ( \40545 , \40544 );
buf \U$40567 ( \40546 , \40545 );
xor \U$40568 ( \40547 , \40519 , \40546 );
buf \U$40569 ( \40548 , \333 );
buf \U$40570 ( \40549 , RIc0da288_95);
not \U$40571 ( \40550 , \40549 );
buf \U$40572 ( \40551 , \40550 );
buf \U$40573 ( \40552 , \40551 );
buf \U$40574 ( \40553 , RIc0d7ab0_10);
and \U$40575 ( \40554 , \40552 , \40553 );
buf \U$40576 ( \40555 , \4546 );
buf \U$40577 ( \40556 , RIc0da288_95);
and \U$40578 ( \40557 , \40555 , \40556 );
nor \U$40579 ( \40558 , \40554 , \40557 );
buf \U$40580 ( \40559 , \40558 );
buf \U$40581 ( \40560 , \40559 );
or \U$40582 ( \40561 , \40548 , \40560 );
buf \U$40583 ( \40562 , \4849 );
buf \U$40584 ( \40563 , \40551 );
buf \U$40585 ( \40564 , RIc0d7a38_9);
and \U$40586 ( \40565 , \40563 , \40564 );
buf \U$40587 ( \40566 , \5976 );
buf \U$40588 ( \40567 , RIc0da288_95);
and \U$40589 ( \40568 , \40566 , \40567 );
nor \U$40590 ( \40569 , \40565 , \40568 );
buf \U$40591 ( \40570 , \40569 );
buf \U$40592 ( \40571 , \40570 );
or \U$40593 ( \40572 , \40562 , \40571 );
nand \U$40594 ( \40573 , \40561 , \40572 );
buf \U$40595 ( \40574 , \40573 );
buf \U$40596 ( \40575 , \40574 );
xor \U$40597 ( \40576 , \40547 , \40575 );
buf \U$40598 ( \40577 , \40576 );
buf \U$40599 ( \40578 , \40577 );
xor \U$40600 ( \40579 , \40502 , \40578 );
buf \U$40601 ( \40580 , \40579 );
buf \U$40602 ( \40581 , \40580 );
xor \U$40603 ( \40582 , \40358 , \40581 );
or \U$40604 ( \40583 , \39314 , \39334 );
nand \U$40605 ( \40584 , \40583 , \39309 );
buf \U$40606 ( \40585 , \40584 );
buf \U$40607 ( \40586 , \39314 );
buf \U$40608 ( \40587 , \39334 );
nand \U$40609 ( \40588 , \40586 , \40587 );
buf \U$40610 ( \40589 , \40588 );
buf \U$40611 ( \40590 , \40589 );
nand \U$40612 ( \40591 , \40585 , \40590 );
buf \U$40613 ( \40592 , \40591 );
buf \U$40614 ( \40593 , \40592 );
buf \U$40615 ( \40594 , \39251 );
buf \U$40616 ( \40595 , \38805 );
or \U$40617 ( \40596 , \40594 , \40595 );
buf \U$40618 ( \40597 , \39231 );
nand \U$40619 ( \40598 , \40596 , \40597 );
buf \U$40620 ( \40599 , \40598 );
buf \U$40621 ( \40600 , \40599 );
buf \U$40622 ( \40601 , \39251 );
buf \U$40623 ( \40602 , \38805 );
nand \U$40624 ( \40603 , \40601 , \40602 );
buf \U$40625 ( \40604 , \40603 );
buf \U$40626 ( \40605 , \40604 );
and \U$40627 ( \40606 , \40600 , \40605 );
buf \U$40628 ( \40607 , \40606 );
buf \U$40629 ( \40608 , \40607 );
not \U$40630 ( \40609 , \40608 );
buf \U$40631 ( \40610 , \40609 );
buf \U$40632 ( \40611 , \40610 );
or \U$40633 ( \40612 , \40593 , \40611 );
xor \U$40634 ( \40613 , \39464 , \39479 );
and \U$40635 ( \40614 , \40613 , \39486 );
and \U$40636 ( \40615 , \39464 , \39479 );
or \U$40637 ( \40616 , \40614 , \40615 );
buf \U$40638 ( \40617 , \40616 );
buf \U$40639 ( \40618 , \40617 );
nand \U$40640 ( \40619 , \40612 , \40618 );
buf \U$40641 ( \40620 , \40619 );
buf \U$40642 ( \40621 , \40620 );
buf \U$40643 ( \40622 , \40592 );
buf \U$40644 ( \40623 , \40610 );
nand \U$40645 ( \40624 , \40622 , \40623 );
buf \U$40646 ( \40625 , \40624 );
buf \U$40647 ( \40626 , \40625 );
nand \U$40648 ( \40627 , \40621 , \40626 );
buf \U$40649 ( \40628 , \40627 );
buf \U$40650 ( \40629 , \40628 );
xor \U$40651 ( \40630 , \40582 , \40629 );
buf \U$40652 ( \40631 , \40630 );
buf \U$40653 ( \40632 , \40631 );
buf \U$40654 ( \40633 , \40592 );
not \U$40655 ( \40634 , \40633 );
buf \U$40656 ( \40635 , \40607 );
not \U$40657 ( \40636 , \40635 );
and \U$40658 ( \40637 , \40634 , \40636 );
buf \U$40659 ( \40638 , \40592 );
buf \U$40660 ( \40639 , \40607 );
and \U$40661 ( \40640 , \40638 , \40639 );
nor \U$40662 ( \40641 , \40637 , \40640 );
buf \U$40663 ( \40642 , \40641 );
buf \U$40664 ( \40643 , \40642 );
buf \U$40665 ( \40644 , \40617 );
xor \U$40666 ( \40645 , \40643 , \40644 );
buf \U$40667 ( \40646 , \40645 );
buf \U$40668 ( \40647 , \40646 );
not \U$40669 ( \40648 , \40647 );
buf \U$40670 ( \40649 , \39349 );
not \U$40671 ( \40650 , \40649 );
buf \U$40672 ( \40651 , \39335 );
not \U$40673 ( \40652 , \40651 );
buf \U$40674 ( \40653 , \40652 );
buf \U$40675 ( \40654 , \40653 );
not \U$40676 ( \40655 , \40654 );
or \U$40677 ( \40656 , \40650 , \40655 );
buf \U$40678 ( \40657 , \40653 );
buf \U$40679 ( \40658 , \39349 );
or \U$40680 ( \40659 , \40657 , \40658 );
buf \U$40681 ( \40660 , \39302 );
nand \U$40682 ( \40661 , \40659 , \40660 );
buf \U$40683 ( \40662 , \40661 );
buf \U$40684 ( \40663 , \40662 );
nand \U$40685 ( \40664 , \40656 , \40663 );
buf \U$40686 ( \40665 , \40664 );
buf \U$40687 ( \40666 , \40665 );
not \U$40688 ( \40667 , \40666 );
buf \U$40689 ( \40668 , \40667 );
buf \U$40690 ( \40669 , \40668 );
not \U$40691 ( \40670 , \40669 );
or \U$40692 ( \40671 , \40648 , \40670 );
buf \U$40693 ( \40672 , \39783 );
buf \U$40694 ( \40673 , \39488 );
or \U$40695 ( \40674 , \40672 , \40673 );
buf \U$40696 ( \40675 , \39603 );
nand \U$40697 ( \40676 , \40674 , \40675 );
buf \U$40698 ( \40677 , \40676 );
buf \U$40699 ( \40678 , \40677 );
buf \U$40700 ( \40679 , \39783 );
buf \U$40701 ( \40680 , \39488 );
nand \U$40702 ( \40681 , \40679 , \40680 );
buf \U$40703 ( \40682 , \40681 );
buf \U$40704 ( \40683 , \40682 );
nand \U$40705 ( \40684 , \40678 , \40683 );
buf \U$40706 ( \40685 , \40684 );
buf \U$40707 ( \40686 , \40685 );
nand \U$40708 ( \40687 , \40671 , \40686 );
buf \U$40709 ( \40688 , \40687 );
buf \U$40710 ( \40689 , \40688 );
buf \U$40711 ( \40690 , \40646 );
not \U$40712 ( \40691 , \40690 );
buf \U$40713 ( \40692 , \40665 );
nand \U$40714 ( \40693 , \40691 , \40692 );
buf \U$40715 ( \40694 , \40693 );
buf \U$40716 ( \40695 , \40694 );
nand \U$40717 ( \40696 , \40689 , \40695 );
buf \U$40718 ( \40697 , \40696 );
buf \U$40719 ( \40698 , \40697 );
xor \U$40720 ( \40699 , \40632 , \40698 );
buf \U$40721 ( \40700 , RIc0d7f60_20);
buf \U$40722 ( \40701 , RIc0d9dd8_85);
xor \U$40723 ( \40702 , \40700 , \40701 );
buf \U$40724 ( \40703 , \40702 );
buf \U$40725 ( \40704 , \40703 );
not \U$40726 ( \40705 , \40704 );
buf \U$40727 ( \40706 , \6029 );
not \U$40728 ( \40707 , \40706 );
or \U$40729 ( \40708 , \40705 , \40707 );
buf \U$40730 ( \40709 , RIc0d7ee8_19);
buf \U$40731 ( \40710 , RIc0d9dd8_85);
xnor \U$40732 ( \40711 , \40709 , \40710 );
buf \U$40733 ( \40712 , \40711 );
buf \U$40734 ( \40713 , \40712 );
not \U$40735 ( \40714 , \40713 );
buf \U$40736 ( \40715 , \2960 );
nand \U$40737 ( \40716 , \40714 , \40715 );
buf \U$40738 ( \40717 , \40716 );
buf \U$40739 ( \40718 , \40717 );
nand \U$40740 ( \40719 , \40708 , \40718 );
buf \U$40741 ( \40720 , \40719 );
buf \U$40742 ( \40721 , \40720 );
buf \U$40743 ( \40722 , RIc0d86e0_36);
buf \U$40744 ( \40723 , RIc0d9658_69);
xor \U$40745 ( \40724 , \40722 , \40723 );
buf \U$40746 ( \40725 , \40724 );
buf \U$40747 ( \40726 , \40725 );
not \U$40748 ( \40727 , \40726 );
buf \U$40749 ( \40728 , \864 );
not \U$40750 ( \40729 , \40728 );
or \U$40751 ( \40730 , \40727 , \40729 );
buf \U$40752 ( \40731 , \284 );
buf \U$40753 ( \40732 , RIc0d8668_35);
buf \U$40754 ( \40733 , RIc0d9658_69);
xor \U$40755 ( \40734 , \40732 , \40733 );
buf \U$40756 ( \40735 , \40734 );
buf \U$40757 ( \40736 , \40735 );
nand \U$40758 ( \40737 , \40731 , \40736 );
buf \U$40759 ( \40738 , \40737 );
buf \U$40760 ( \40739 , \40738 );
nand \U$40761 ( \40740 , \40730 , \40739 );
buf \U$40762 ( \40741 , \40740 );
buf \U$40763 ( \40742 , \40741 );
xor \U$40764 ( \40743 , \40721 , \40742 );
buf \U$40765 ( \40744 , \989 );
buf \U$40766 ( \40745 , RIc0d8050_22);
buf \U$40767 ( \40746 , RIc0d9ce8_83);
xnor \U$40768 ( \40747 , \40745 , \40746 );
buf \U$40769 ( \40748 , \40747 );
buf \U$40770 ( \40749 , \40748 );
or \U$40771 ( \40750 , \40744 , \40749 );
buf \U$40772 ( \40751 , \996 );
buf \U$40773 ( \40752 , \1050 );
buf \U$40774 ( \40753 , RIc0d7fd8_21);
and \U$40775 ( \40754 , \40752 , \40753 );
buf \U$40776 ( \40755 , \16240 );
buf \U$40777 ( \40756 , RIc0d9ce8_83);
and \U$40778 ( \40757 , \40755 , \40756 );
nor \U$40779 ( \40758 , \40754 , \40757 );
buf \U$40780 ( \40759 , \40758 );
buf \U$40781 ( \40760 , \40759 );
or \U$40782 ( \40761 , \40751 , \40760 );
nand \U$40783 ( \40762 , \40750 , \40761 );
buf \U$40784 ( \40763 , \40762 );
buf \U$40785 ( \40764 , \40763 );
xor \U$40786 ( \40765 , \40743 , \40764 );
buf \U$40787 ( \40766 , \40765 );
buf \U$40788 ( \40767 , \40766 );
buf \U$40789 ( \40768 , \39178 );
not \U$40790 ( \40769 , \40768 );
buf \U$40791 ( \40770 , \2607 );
not \U$40792 ( \40771 , \40770 );
or \U$40793 ( \40772 , \40769 , \40771 );
buf \U$40794 ( \40773 , \3631 );
buf \U$40795 ( \40774 , \40455 );
nand \U$40796 ( \40775 , \40773 , \40774 );
buf \U$40797 ( \40776 , \40775 );
buf \U$40798 ( \40777 , \40776 );
nand \U$40799 ( \40778 , \40772 , \40777 );
buf \U$40800 ( \40779 , \40778 );
buf \U$40801 ( \40780 , \12744 );
not \U$40802 ( \40781 , \40780 );
buf \U$40803 ( \40782 , \40781 );
buf \U$40804 ( \40783 , \40782 );
not \U$40805 ( \40784 , \40783 );
buf \U$40806 ( \40785 , \12736 );
not \U$40807 ( \40786 , \40785 );
buf \U$40808 ( \40787 , \40786 );
buf \U$40809 ( \40788 , \40787 );
not \U$40810 ( \40789 , \40788 );
or \U$40811 ( \40790 , \40784 , \40789 );
buf \U$40812 ( \40791 , RIc0da738_105);
nand \U$40813 ( \40792 , \40790 , \40791 );
buf \U$40814 ( \40793 , \40792 );
buf \U$40815 ( \40794 , \40793 );
not \U$40816 ( \40795 , \40794 );
buf \U$40817 ( \40796 , \40795 );
xor \U$40818 ( \40797 , \40779 , \40796 );
and \U$40819 ( \40798 , \36497 , \36498 );
buf \U$40820 ( \40799 , \40798 );
buf \U$40821 ( \40800 , \40799 );
buf \U$40822 ( \40801 , \39724 );
not \U$40823 ( \40802 , \40801 );
buf \U$40824 ( \40803 , \6029 );
not \U$40825 ( \40804 , \40803 );
or \U$40826 ( \40805 , \40802 , \40804 );
buf \U$40827 ( \40806 , \921 );
buf \U$40828 ( \40807 , \40703 );
nand \U$40829 ( \40808 , \40806 , \40807 );
buf \U$40830 ( \40809 , \40808 );
buf \U$40831 ( \40810 , \40809 );
nand \U$40832 ( \40811 , \40805 , \40810 );
buf \U$40833 ( \40812 , \40811 );
buf \U$40834 ( \40813 , \40812 );
xor \U$40835 ( \40814 , \40800 , \40813 );
buf \U$40836 ( \40815 , \27591 );
not \U$40837 ( \40816 , \40815 );
buf \U$40838 ( \40817 , \40816 );
buf \U$40839 ( \40818 , \40817 );
buf \U$40840 ( \40819 , \39648 );
or \U$40841 ( \40820 , \40818 , \40819 );
buf \U$40842 ( \40821 , \14704 );
buf \U$40843 ( \40822 , \40559 );
or \U$40844 ( \40823 , \40821 , \40822 );
nand \U$40845 ( \40824 , \40820 , \40823 );
buf \U$40846 ( \40825 , \40824 );
buf \U$40847 ( \40826 , \40825 );
and \U$40848 ( \40827 , \40814 , \40826 );
and \U$40849 ( \40828 , \40800 , \40813 );
or \U$40850 ( \40829 , \40827 , \40828 );
buf \U$40851 ( \40830 , \40829 );
xnor \U$40852 ( \40831 , \40797 , \40830 );
buf \U$40853 ( \40832 , \40831 );
xor \U$40854 ( \40833 , \40767 , \40832 );
buf \U$40855 ( \40834 , \39688 );
not \U$40856 ( \40835 , \40834 );
buf \U$40857 ( \40836 , \39675 );
not \U$40858 ( \40837 , \40836 );
or \U$40859 ( \40838 , \40835 , \40837 );
buf \U$40860 ( \40839 , \39675 );
buf \U$40861 ( \40840 , \39688 );
or \U$40862 ( \40841 , \40839 , \40840 );
buf \U$40863 ( \40842 , \39705 );
nand \U$40864 ( \40843 , \40841 , \40842 );
buf \U$40865 ( \40844 , \40843 );
buf \U$40866 ( \40845 , \40844 );
nand \U$40867 ( \40846 , \40838 , \40845 );
buf \U$40868 ( \40847 , \40846 );
buf \U$40869 ( \40848 , \40847 );
xor \U$40870 ( \40849 , \39491 , \39508 );
and \U$40871 ( \40850 , \40849 , \39523 );
and \U$40872 ( \40851 , \39491 , \39508 );
or \U$40873 ( \40852 , \40850 , \40851 );
buf \U$40874 ( \40853 , \40852 );
buf \U$40875 ( \40854 , \40853 );
or \U$40876 ( \40855 , \40848 , \40854 );
buf \U$40877 ( \40856 , \39204 );
not \U$40878 ( \40857 , \40856 );
buf \U$40879 ( \40858 , \39184 );
not \U$40880 ( \40859 , \40858 );
or \U$40881 ( \40860 , \40857 , \40859 );
buf \U$40882 ( \40861 , \39184 );
buf \U$40883 ( \40862 , \39204 );
or \U$40884 ( \40863 , \40861 , \40862 );
buf \U$40885 ( \40864 , \39170 );
nand \U$40886 ( \40865 , \40863 , \40864 );
buf \U$40887 ( \40866 , \40865 );
buf \U$40888 ( \40867 , \40866 );
nand \U$40889 ( \40868 , \40860 , \40867 );
buf \U$40890 ( \40869 , \40868 );
buf \U$40891 ( \40870 , \40869 );
nand \U$40892 ( \40871 , \40855 , \40870 );
buf \U$40893 ( \40872 , \40871 );
buf \U$40894 ( \40873 , \40872 );
buf \U$40895 ( \40874 , \40847 );
buf \U$40896 ( \40875 , \40853 );
nand \U$40897 ( \40876 , \40874 , \40875 );
buf \U$40898 ( \40877 , \40876 );
buf \U$40899 ( \40878 , \40877 );
nand \U$40900 ( \40879 , \40873 , \40878 );
buf \U$40901 ( \40880 , \40879 );
buf \U$40902 ( \40881 , \40880 );
xor \U$40903 ( \40882 , \40833 , \40881 );
buf \U$40904 ( \40883 , \40882 );
buf \U$40905 ( \40884 , \40883 );
xor \U$40906 ( \40885 , \39526 , \39541 );
and \U$40907 ( \40886 , \40885 , \39601 );
and \U$40908 ( \40887 , \39526 , \39541 );
or \U$40909 ( \40888 , \40886 , \40887 );
buf \U$40910 ( \40889 , \40888 );
buf \U$40911 ( \40890 , \40889 );
buf \U$40912 ( \40891 , \39153 );
not \U$40913 ( \40892 , \40891 );
buf \U$40914 ( \40893 , \39128 );
not \U$40915 ( \40894 , \40893 );
or \U$40916 ( \40895 , \40892 , \40894 );
buf \U$40917 ( \40896 , \39128 );
buf \U$40918 ( \40897 , \39153 );
or \U$40919 ( \40898 , \40896 , \40897 );
buf \U$40920 ( \40899 , \39136 );
nand \U$40921 ( \40900 , \40898 , \40899 );
buf \U$40922 ( \40901 , \40900 );
buf \U$40923 ( \40902 , \40901 );
nand \U$40924 ( \40903 , \40895 , \40902 );
buf \U$40925 ( \40904 , \40903 );
buf \U$40926 ( \40905 , \40904 );
xor \U$40927 ( \40906 , \39559 , \39576 );
and \U$40928 ( \40907 , \40906 , \39598 );
and \U$40929 ( \40908 , \39559 , \39576 );
or \U$40930 ( \40909 , \40907 , \40908 );
buf \U$40931 ( \40910 , \40909 );
buf \U$40932 ( \40911 , \40910 );
xor \U$40933 ( \40912 , \40905 , \40911 );
buf \U$40934 ( \40913 , \39501 );
not \U$40935 ( \40914 , \40913 );
buf \U$40936 ( \40915 , \1823 );
not \U$40937 ( \40916 , \40915 );
or \U$40938 ( \40917 , \40914 , \40916 );
buf \U$40939 ( \40918 , \686 );
buf \U$40940 ( \40919 , \40222 );
nand \U$40941 ( \40920 , \40918 , \40919 );
buf \U$40942 ( \40921 , \40920 );
buf \U$40943 ( \40922 , \40921 );
nand \U$40944 ( \40923 , \40917 , \40922 );
buf \U$40945 ( \40924 , \40923 );
buf \U$40946 ( \40925 , \40924 );
buf \U$40947 ( \40926 , \39552 );
not \U$40948 ( \40927 , \40926 );
buf \U$40949 ( \40928 , \1224 );
not \U$40950 ( \40929 , \40928 );
or \U$40951 ( \40930 , \40927 , \40929 );
buf \U$40952 ( \40931 , \1229 );
buf \U$40953 ( \40932 , \40385 );
nand \U$40954 ( \40933 , \40931 , \40932 );
buf \U$40955 ( \40934 , \40933 );
buf \U$40956 ( \40935 , \40934 );
nand \U$40957 ( \40936 , \40930 , \40935 );
buf \U$40958 ( \40937 , \40936 );
buf \U$40959 ( \40938 , \40937 );
xor \U$40960 ( \40939 , \40925 , \40938 );
buf \U$40961 ( \40940 , \39516 );
not \U$40962 ( \40941 , \40940 );
buf \U$40963 ( \40942 , \1927 );
not \U$40964 ( \40943 , \40942 );
or \U$40965 ( \40944 , \40941 , \40943 );
buf \U$40966 ( \40945 , \1933 );
buf \U$40967 ( \40946 , \40251 );
nand \U$40968 ( \40947 , \40945 , \40946 );
buf \U$40969 ( \40948 , \40947 );
buf \U$40970 ( \40949 , \40948 );
nand \U$40971 ( \40950 , \40944 , \40949 );
buf \U$40972 ( \40951 , \40950 );
buf \U$40973 ( \40952 , \40951 );
xor \U$40974 ( \40953 , \40939 , \40952 );
buf \U$40975 ( \40954 , \40953 );
buf \U$40976 ( \40955 , \40954 );
xor \U$40977 ( \40956 , \40912 , \40955 );
buf \U$40978 ( \40957 , \40956 );
buf \U$40979 ( \40958 , \40957 );
xor \U$40980 ( \40959 , \40890 , \40958 );
buf \U$40981 ( \40960 , \40779 );
not \U$40982 ( \40961 , \40960 );
buf \U$40983 ( \40962 , \40961 );
buf \U$40984 ( \40963 , \40962 );
xor \U$40985 ( \40964 , \39731 , \39748 );
and \U$40986 ( \40965 , \40964 , \39766 );
and \U$40987 ( \40966 , \39731 , \39748 );
or \U$40988 ( \40967 , \40965 , \40966 );
buf \U$40989 ( \40968 , \40967 );
buf \U$40990 ( \40969 , \40968 );
xor \U$40991 ( \40970 , \40963 , \40969 );
xor \U$40992 ( \40971 , \39621 , \39638 );
and \U$40993 ( \40972 , \40971 , \39657 );
and \U$40994 ( \40973 , \39621 , \39638 );
or \U$40995 ( \40974 , \40972 , \40973 );
buf \U$40996 ( \40975 , \40974 );
buf \U$40997 ( \40976 , \40975 );
xor \U$40998 ( \40977 , \40970 , \40976 );
buf \U$40999 ( \40978 , \40977 );
buf \U$41000 ( \40979 , \40978 );
and \U$41001 ( \40980 , \40959 , \40979 );
and \U$41002 ( \40981 , \40890 , \40958 );
or \U$41003 ( \40982 , \40980 , \40981 );
buf \U$41004 ( \40983 , \40982 );
buf \U$41005 ( \40984 , \40983 );
xor \U$41006 ( \40985 , \40884 , \40984 );
xor \U$41007 ( \40986 , \40963 , \40969 );
and \U$41008 ( \40987 , \40986 , \40976 );
and \U$41009 ( \40988 , \40963 , \40969 );
or \U$41010 ( \40989 , \40987 , \40988 );
buf \U$41011 ( \40990 , \40989 );
buf \U$41012 ( \40991 , \40990 );
xor \U$41013 ( \40992 , \40925 , \40938 );
and \U$41014 ( \40993 , \40992 , \40952 );
and \U$41015 ( \40994 , \40925 , \40938 );
or \U$41016 ( \40995 , \40993 , \40994 );
buf \U$41017 ( \40996 , \40995 );
buf \U$41018 ( \40997 , \40996 );
buf \U$41019 ( \40998 , \39198 );
not \U$41020 ( \40999 , \40998 );
buf \U$41021 ( \41000 , \2871 );
not \U$41022 ( \41001 , \41000 );
or \U$41023 ( \41002 , \40999 , \41001 );
buf \U$41024 ( \41003 , \792 );
buf \U$41025 ( \41004 , \40286 );
nand \U$41026 ( \41005 , \41003 , \41004 );
buf \U$41027 ( \41006 , \41005 );
buf \U$41028 ( \41007 , \41006 );
nand \U$41029 ( \41008 , \41002 , \41007 );
buf \U$41030 ( \41009 , \41008 );
buf \U$41031 ( \41010 , \41009 );
not \U$41032 ( \41011 , \41010 );
buf \U$41033 ( \41012 , \39245 );
not \U$41034 ( \41013 , \41012 );
buf \U$41035 ( \41014 , \12736 );
not \U$41036 ( \41015 , \41014 );
or \U$41037 ( \41016 , \41013 , \41015 );
buf \U$41038 ( \41017 , \21880 );
buf \U$41039 ( \41018 , RIc0da738_105);
nand \U$41040 ( \41019 , \41017 , \41018 );
buf \U$41041 ( \41020 , \41019 );
buf \U$41042 ( \41021 , \41020 );
nand \U$41043 ( \41022 , \41016 , \41021 );
buf \U$41044 ( \41023 , \41022 );
buf \U$41045 ( \41024 , \41023 );
not \U$41046 ( \41025 , \41024 );
or \U$41047 ( \41026 , \41011 , \41025 );
buf \U$41048 ( \41027 , \41023 );
buf \U$41049 ( \41028 , \41009 );
or \U$41050 ( \41029 , \41027 , \41028 );
buf \U$41051 ( \41030 , \1739 );
not \U$41052 ( \41031 , \41030 );
buf \U$41053 ( \41032 , \39120 );
not \U$41054 ( \41033 , \41032 );
and \U$41055 ( \41034 , \41031 , \41033 );
buf \U$41056 ( \41035 , \996 );
buf \U$41057 ( \41036 , \40748 );
nor \U$41058 ( \41037 , \41035 , \41036 );
buf \U$41059 ( \41038 , \41037 );
buf \U$41060 ( \41039 , \41038 );
nor \U$41061 ( \41040 , \41034 , \41039 );
buf \U$41062 ( \41041 , \41040 );
buf \U$41063 ( \41042 , \41041 );
not \U$41064 ( \41043 , \41042 );
buf \U$41065 ( \41044 , \41043 );
buf \U$41066 ( \41045 , \41044 );
nand \U$41067 ( \41046 , \41029 , \41045 );
buf \U$41068 ( \41047 , \41046 );
buf \U$41069 ( \41048 , \41047 );
nand \U$41070 ( \41049 , \41026 , \41048 );
buf \U$41071 ( \41050 , \41049 );
buf \U$41072 ( \41051 , \41050 );
xor \U$41073 ( \41052 , \40997 , \41051 );
buf \U$41074 ( \41053 , \39147 );
not \U$41075 ( \41054 , \41053 );
buf \U$41076 ( \41055 , \864 );
not \U$41077 ( \41056 , \41055 );
or \U$41078 ( \41057 , \41054 , \41056 );
buf \U$41079 ( \41058 , \284 );
buf \U$41080 ( \41059 , \40725 );
nand \U$41081 ( \41060 , \41058 , \41059 );
buf \U$41082 ( \41061 , \41060 );
buf \U$41083 ( \41062 , \41061 );
nand \U$41084 ( \41063 , \41057 , \41062 );
buf \U$41085 ( \41064 , \41063 );
buf \U$41086 ( \41065 , \41064 );
not \U$41087 ( \41066 , \41065 );
buf \U$41088 ( \41067 , \39614 );
not \U$41089 ( \41068 , \41067 );
buf \U$41090 ( \41069 , \1064 );
not \U$41091 ( \41070 , \41069 );
or \U$41092 ( \41071 , \41068 , \41070 );
buf \U$41093 ( \41072 , \40507 );
not \U$41094 ( \41073 , \41072 );
buf \U$41095 ( \41074 , \1078 );
nand \U$41096 ( \41075 , \41073 , \41074 );
buf \U$41097 ( \41076 , \41075 );
buf \U$41098 ( \41077 , \41076 );
nand \U$41099 ( \41078 , \41071 , \41077 );
buf \U$41100 ( \41079 , \41078 );
buf \U$41101 ( \41080 , \41079 );
not \U$41102 ( \41081 , \41080 );
or \U$41103 ( \41082 , \41066 , \41081 );
buf \U$41104 ( \41083 , \41079 );
buf \U$41105 ( \41084 , \41064 );
or \U$41106 ( \41085 , \41083 , \41084 );
buf \U$41107 ( \41086 , \39699 );
not \U$41108 ( \41087 , \41086 );
buf \U$41109 ( \41088 , \1432 );
not \U$41110 ( \41089 , \41088 );
or \U$41111 ( \41090 , \41087 , \41089 );
buf \U$41112 ( \41091 , \3742 );
buf \U$41113 ( \41092 , \40152 );
nand \U$41114 ( \41093 , \41091 , \41092 );
buf \U$41115 ( \41094 , \41093 );
buf \U$41116 ( \41095 , \41094 );
nand \U$41117 ( \41096 , \41090 , \41095 );
buf \U$41118 ( \41097 , \41096 );
buf \U$41119 ( \41098 , \41097 );
nand \U$41120 ( \41099 , \41085 , \41098 );
buf \U$41121 ( \41100 , \41099 );
buf \U$41122 ( \41101 , \41100 );
nand \U$41123 ( \41102 , \41082 , \41101 );
buf \U$41124 ( \41103 , \41102 );
buf \U$41125 ( \41104 , \41103 );
xor \U$41126 ( \41105 , \41052 , \41104 );
buf \U$41127 ( \41106 , \41105 );
buf \U$41128 ( \41107 , \41106 );
xor \U$41129 ( \41108 , \40991 , \41107 );
buf \U$41130 ( \41109 , \39569 );
not \U$41131 ( \41110 , \41109 );
buf \U$41132 ( \41111 , \2812 );
not \U$41133 ( \41112 , \41111 );
or \U$41134 ( \41113 , \41110 , \41112 );
buf \U$41135 ( \41114 , \1276 );
buf \U$41136 ( \41115 , \40362 );
nand \U$41137 ( \41116 , \41114 , \41115 );
buf \U$41138 ( \41117 , \41116 );
buf \U$41139 ( \41118 , \41117 );
nand \U$41140 ( \41119 , \41113 , \41118 );
buf \U$41141 ( \41120 , \41119 );
buf \U$41142 ( \41121 , \41120 );
buf \U$41143 ( \41122 , \39225 );
not \U$41144 ( \41123 , \41122 );
buf \U$41145 ( \41124 , \18220 );
not \U$41146 ( \41125 , \41124 );
or \U$41147 ( \41126 , \41123 , \41125 );
buf \U$41148 ( \41127 , \40527 );
not \U$41149 ( \41128 , \41127 );
buf \U$41150 ( \41129 , \13048 );
nand \U$41151 ( \41130 , \41128 , \41129 );
buf \U$41152 ( \41131 , \41130 );
buf \U$41153 ( \41132 , \41131 );
nand \U$41154 ( \41133 , \41126 , \41132 );
buf \U$41155 ( \41134 , \41133 );
buf \U$41156 ( \41135 , \41134 );
xor \U$41157 ( \41136 , \41121 , \41135 );
buf \U$41158 ( \41137 , \39591 );
not \U$41159 ( \41138 , \41137 );
buf \U$41160 ( \41139 , \29069 );
not \U$41161 ( \41140 , \41139 );
or \U$41162 ( \41141 , \41138 , \41140 );
buf \U$41163 ( \41142 , \2070 );
buf \U$41164 ( \41143 , \40407 );
nand \U$41165 ( \41144 , \41142 , \41143 );
buf \U$41166 ( \41145 , \41144 );
buf \U$41167 ( \41146 , \41145 );
nand \U$41168 ( \41147 , \41141 , \41146 );
buf \U$41169 ( \41148 , \41147 );
buf \U$41170 ( \41149 , \41148 );
xor \U$41171 ( \41150 , \41136 , \41149 );
buf \U$41172 ( \41151 , \41150 );
buf \U$41173 ( \41152 , \41151 );
buf \U$41174 ( \41153 , \39741 );
not \U$41175 ( \41154 , \41153 );
buf \U$41176 ( \41155 , \396 );
not \U$41177 ( \41156 , \41155 );
or \U$41178 ( \41157 , \41154 , \41156 );
buf \U$41179 ( \41158 , \402 );
buf \U$41180 ( \41159 , \40307 );
nand \U$41181 ( \41160 , \41158 , \41159 );
buf \U$41182 ( \41161 , \41160 );
buf \U$41183 ( \41162 , \41161 );
nand \U$41184 ( \41163 , \41157 , \41162 );
buf \U$41185 ( \41164 , \41163 );
buf \U$41186 ( \41165 , \41164 );
buf \U$41187 ( \41166 , \39759 );
not \U$41188 ( \41167 , \41166 );
buf \U$41189 ( \41168 , \1901 );
not \U$41190 ( \41169 , \41168 );
or \U$41191 ( \41170 , \41167 , \41169 );
buf \U$41192 ( \41171 , \4008 );
buf \U$41193 ( \41172 , \40331 );
nand \U$41194 ( \41173 , \41171 , \41172 );
buf \U$41195 ( \41174 , \41173 );
buf \U$41196 ( \41175 , \41174 );
nand \U$41197 ( \41176 , \41170 , \41175 );
buf \U$41198 ( \41177 , \41176 );
buf \U$41199 ( \41178 , \41177 );
xor \U$41200 ( \41179 , \41165 , \41178 );
buf \U$41201 ( \41180 , \39631 );
not \U$41202 ( \41181 , \41180 );
buf \U$41203 ( \41182 , \22631 );
not \U$41204 ( \41183 , \41182 );
or \U$41205 ( \41184 , \41181 , \41183 );
buf \U$41206 ( \41185 , \16676 );
buf \U$41207 ( \41186 , \40195 );
nand \U$41208 ( \41187 , \41185 , \41186 );
buf \U$41209 ( \41188 , \41187 );
buf \U$41210 ( \41189 , \41188 );
nand \U$41211 ( \41190 , \41184 , \41189 );
buf \U$41212 ( \41191 , \41190 );
buf \U$41213 ( \41192 , \41191 );
xor \U$41214 ( \41193 , \41179 , \41192 );
buf \U$41215 ( \41194 , \41193 );
buf \U$41216 ( \41195 , \41194 );
xor \U$41217 ( \41196 , \41152 , \41195 );
buf \U$41218 ( \41197 , \39682 );
not \U$41219 ( \41198 , \41197 );
buf \U$41220 ( \41199 , \36975 );
not \U$41221 ( \41200 , \41199 );
or \U$41222 ( \41201 , \41198 , \41200 );
buf \U$41223 ( \41202 , \1143 );
buf \U$41224 ( \41203 , \40170 );
nand \U$41225 ( \41204 , \41202 , \41203 );
buf \U$41226 ( \41205 , \41204 );
buf \U$41227 ( \41206 , \41205 );
nand \U$41228 ( \41207 , \41201 , \41206 );
buf \U$41229 ( \41208 , \41207 );
buf \U$41230 ( \41209 , \41208 );
buf \U$41231 ( \41210 , \39164 );
not \U$41232 ( \41211 , \41210 );
buf \U$41233 ( \41212 , \19695 );
not \U$41234 ( \41213 , \41212 );
or \U$41235 ( \41214 , \41211 , \41213 );
buf \U$41236 ( \41215 , \40479 );
not \U$41237 ( \41216 , \41215 );
buf \U$41238 ( \41217 , \14140 );
nand \U$41239 ( \41218 , \41216 , \41217 );
buf \U$41240 ( \41219 , \41218 );
buf \U$41241 ( \41220 , \41219 );
nand \U$41242 ( \41221 , \41214 , \41220 );
buf \U$41243 ( \41222 , \41221 );
buf \U$41244 ( \41223 , \41222 );
xor \U$41245 ( \41224 , \41209 , \41223 );
buf \U$41246 ( \41225 , \39669 );
not \U$41247 ( \41226 , \41225 );
buf \U$41248 ( \41227 , \2038 );
not \U$41249 ( \41228 , \41227 );
or \U$41250 ( \41229 , \41226 , \41228 );
buf \U$41251 ( \41230 , \442 );
buf \U$41252 ( \41231 , \40429 );
nand \U$41253 ( \41232 , \41230 , \41231 );
buf \U$41254 ( \41233 , \41232 );
buf \U$41255 ( \41234 , \41233 );
nand \U$41256 ( \41235 , \41229 , \41234 );
buf \U$41257 ( \41236 , \41235 );
buf \U$41258 ( \41237 , \41236 );
xor \U$41259 ( \41238 , \41224 , \41237 );
buf \U$41260 ( \41239 , \41238 );
buf \U$41261 ( \41240 , \41239 );
and \U$41262 ( \41241 , \41196 , \41240 );
and \U$41263 ( \41242 , \41152 , \41195 );
or \U$41264 ( \41243 , \41241 , \41242 );
buf \U$41265 ( \41244 , \41243 );
buf \U$41266 ( \41245 , \41244 );
xor \U$41267 ( \41246 , \41108 , \41245 );
buf \U$41268 ( \41247 , \41246 );
buf \U$41269 ( \41248 , \41247 );
xor \U$41270 ( \41249 , \40985 , \41248 );
buf \U$41271 ( \41250 , \41249 );
buf \U$41272 ( \41251 , \41250 );
xor \U$41273 ( \41252 , \40699 , \41251 );
buf \U$41274 ( \41253 , \41252 );
buf \U$41275 ( \41254 , \41253 );
buf \U$41276 ( \41255 , \39768 );
not \U$41277 ( \41256 , \41255 );
buf \U$41278 ( \41257 , \39706 );
not \U$41279 ( \41258 , \41257 );
or \U$41280 ( \41259 , \41256 , \41258 );
buf \U$41281 ( \41260 , \39706 );
buf \U$41282 ( \41261 , \39768 );
or \U$41283 ( \41262 , \41260 , \41261 );
buf \U$41284 ( \41263 , \39659 );
nand \U$41285 ( \41264 , \41262 , \41263 );
buf \U$41286 ( \41265 , \41264 );
buf \U$41287 ( \41266 , \41265 );
nand \U$41288 ( \41267 , \41259 , \41266 );
buf \U$41289 ( \41268 , \41267 );
buf \U$41290 ( \41269 , \41268 );
not \U$41291 ( \41270 , \41269 );
buf \U$41292 ( \41271 , \40869 );
buf \U$41293 ( \41272 , \40847 );
xor \U$41294 ( \41273 , \41271 , \41272 );
buf \U$41295 ( \41274 , \41273 );
buf \U$41296 ( \41275 , \41274 );
not \U$41297 ( \41276 , \41275 );
buf \U$41298 ( \41277 , \40853 );
not \U$41299 ( \41278 , \41277 );
buf \U$41300 ( \41279 , \41278 );
buf \U$41301 ( \41280 , \41279 );
not \U$41302 ( \41281 , \41280 );
and \U$41303 ( \41282 , \41276 , \41281 );
buf \U$41304 ( \41283 , \41274 );
buf \U$41305 ( \41284 , \41279 );
and \U$41306 ( \41285 , \41283 , \41284 );
nor \U$41307 ( \41286 , \41282 , \41285 );
buf \U$41308 ( \41287 , \41286 );
buf \U$41309 ( \41288 , \41287 );
not \U$41310 ( \41289 , \41288 );
buf \U$41311 ( \41290 , \41289 );
buf \U$41312 ( \41291 , \41290 );
not \U$41313 ( \41292 , \41291 );
or \U$41314 ( \41293 , \41270 , \41292 );
buf \U$41315 ( \41294 , \41290 );
buf \U$41316 ( \41295 , \41268 );
or \U$41317 ( \41296 , \41294 , \41295 );
buf \U$41318 ( \41297 , \39263 );
buf \U$41319 ( \41298 , \39214 );
or \U$41320 ( \41299 , \41297 , \41298 );
buf \U$41321 ( \41300 , \39154 );
not \U$41322 ( \41301 , \41300 );
buf \U$41323 ( \41302 , \41301 );
buf \U$41324 ( \41303 , \41302 );
nand \U$41325 ( \41304 , \41299 , \41303 );
buf \U$41326 ( \41305 , \41304 );
buf \U$41327 ( \41306 , \41305 );
buf \U$41328 ( \41307 , \39263 );
buf \U$41329 ( \41308 , \39214 );
nand \U$41330 ( \41309 , \41307 , \41308 );
buf \U$41331 ( \41310 , \41309 );
buf \U$41332 ( \41311 , \41310 );
nand \U$41333 ( \41312 , \41306 , \41311 );
buf \U$41334 ( \41313 , \41312 );
buf \U$41335 ( \41314 , \41313 );
nand \U$41336 ( \41315 , \41296 , \41314 );
buf \U$41337 ( \41316 , \41315 );
buf \U$41338 ( \41317 , \41316 );
nand \U$41339 ( \41318 , \41293 , \41317 );
buf \U$41340 ( \41319 , \41318 );
buf \U$41341 ( \41320 , \41319 );
xor \U$41342 ( \41321 , \40905 , \40911 );
and \U$41343 ( \41322 , \41321 , \40955 );
and \U$41344 ( \41323 , \40905 , \40911 );
or \U$41345 ( \41324 , \41322 , \41323 );
buf \U$41346 ( \41325 , \41324 );
buf \U$41347 ( \41326 , \41325 );
xor \U$41348 ( \41327 , \41165 , \41178 );
and \U$41349 ( \41328 , \41327 , \41192 );
and \U$41350 ( \41329 , \41165 , \41178 );
or \U$41351 ( \41330 , \41328 , \41329 );
buf \U$41352 ( \41331 , \41330 );
buf \U$41353 ( \41332 , \41331 );
xor \U$41354 ( \41333 , \41121 , \41135 );
and \U$41355 ( \41334 , \41333 , \41149 );
and \U$41356 ( \41335 , \41121 , \41135 );
or \U$41357 ( \41336 , \41334 , \41335 );
buf \U$41358 ( \41337 , \41336 );
buf \U$41359 ( \41338 , \41337 );
xor \U$41360 ( \41339 , \41332 , \41338 );
xor \U$41361 ( \41340 , \41209 , \41223 );
and \U$41362 ( \41341 , \41340 , \41237 );
and \U$41363 ( \41342 , \41209 , \41223 );
or \U$41364 ( \41343 , \41341 , \41342 );
buf \U$41365 ( \41344 , \41343 );
buf \U$41366 ( \41345 , \41344 );
xor \U$41367 ( \41346 , \41339 , \41345 );
buf \U$41368 ( \41347 , \41346 );
buf \U$41369 ( \41348 , \41347 );
xor \U$41370 ( \41349 , \41326 , \41348 );
xor \U$41371 ( \41350 , \40800 , \40813 );
xor \U$41372 ( \41351 , \41350 , \40826 );
buf \U$41373 ( \41352 , \41351 );
buf \U$41374 ( \41353 , \41352 );
xor \U$41375 ( \41354 , \41009 , \41023 );
xnor \U$41376 ( \41355 , \41354 , \41041 );
buf \U$41377 ( \41356 , \41355 );
xor \U$41378 ( \41357 , \41353 , \41356 );
buf \U$41379 ( \41358 , \41079 );
buf \U$41380 ( \41359 , \41064 );
xor \U$41381 ( \41360 , \41358 , \41359 );
buf \U$41382 ( \41361 , \41360 );
buf \U$41383 ( \41362 , \41361 );
buf \U$41384 ( \41363 , \41097 );
xor \U$41385 ( \41364 , \41362 , \41363 );
buf \U$41386 ( \41365 , \41364 );
buf \U$41387 ( \41366 , \41365 );
and \U$41388 ( \41367 , \41357 , \41366 );
and \U$41389 ( \41368 , \41353 , \41356 );
or \U$41390 ( \41369 , \41367 , \41368 );
buf \U$41391 ( \41370 , \41369 );
buf \U$41392 ( \41371 , \41370 );
xor \U$41393 ( \41372 , \41349 , \41371 );
buf \U$41394 ( \41373 , \41372 );
buf \U$41395 ( \41374 , \41373 );
xor \U$41396 ( \41375 , \41320 , \41374 );
xor \U$41397 ( \41376 , \41152 , \41195 );
xor \U$41398 ( \41377 , \41376 , \41240 );
buf \U$41399 ( \41378 , \41377 );
buf \U$41400 ( \41379 , \41378 );
xor \U$41401 ( \41380 , \41353 , \41356 );
xor \U$41402 ( \41381 , \41380 , \41366 );
buf \U$41403 ( \41382 , \41381 );
buf \U$41404 ( \41383 , \41382 );
xor \U$41405 ( \41384 , \41379 , \41383 );
buf \U$41406 ( \41385 , \39410 );
buf \U$41407 ( \41386 , \39385 );
or \U$41408 ( \41387 , \41385 , \41386 );
buf \U$41409 ( \41388 , \39403 );
nand \U$41410 ( \41389 , \41387 , \41388 );
buf \U$41411 ( \41390 , \41389 );
buf \U$41412 ( \41391 , \41390 );
buf \U$41413 ( \41392 , \39410 );
buf \U$41414 ( \41393 , \39385 );
nand \U$41415 ( \41394 , \41392 , \41393 );
buf \U$41416 ( \41395 , \41394 );
buf \U$41417 ( \41396 , \41395 );
nand \U$41418 ( \41397 , \41391 , \41396 );
buf \U$41419 ( \41398 , \41397 );
buf \U$41420 ( \41399 , \41398 );
and \U$41421 ( \41400 , \41384 , \41399 );
and \U$41422 ( \41401 , \41379 , \41383 );
or \U$41423 ( \41402 , \41400 , \41401 );
buf \U$41424 ( \41403 , \41402 );
buf \U$41425 ( \41404 , \41403 );
xor \U$41426 ( \41405 , \41375 , \41404 );
buf \U$41427 ( \41406 , \41405 );
buf \U$41428 ( \41407 , \41406 );
xor \U$41429 ( \41408 , \40890 , \40958 );
xor \U$41430 ( \41409 , \41408 , \40979 );
buf \U$41431 ( \41410 , \41409 );
buf \U$41432 ( \41411 , \41410 );
not \U$41433 ( \41412 , \41411 );
xor \U$41434 ( \41413 , \41287 , \41268 );
xor \U$41435 ( \41414 , \41413 , \41313 );
buf \U$41436 ( \41415 , \41414 );
not \U$41437 ( \41416 , \41415 );
buf \U$41438 ( \41417 , \41416 );
buf \U$41439 ( \41418 , \41417 );
not \U$41440 ( \41419 , \41418 );
or \U$41441 ( \41420 , \41412 , \41419 );
buf \U$41442 ( \41421 , \41417 );
buf \U$41443 ( \41422 , \41410 );
or \U$41444 ( \41423 , \41421 , \41422 );
xor \U$41445 ( \41424 , \41379 , \41383 );
xor \U$41446 ( \41425 , \41424 , \41399 );
buf \U$41447 ( \41426 , \41425 );
buf \U$41448 ( \41427 , \41426 );
nand \U$41449 ( \41428 , \41423 , \41427 );
buf \U$41450 ( \41429 , \41428 );
buf \U$41451 ( \41430 , \41429 );
nand \U$41452 ( \41431 , \41420 , \41430 );
buf \U$41453 ( \41432 , \41431 );
buf \U$41454 ( \41433 , \41432 );
xor \U$41455 ( \41434 , \41407 , \41433 );
xor \U$41456 ( \41435 , \39265 , \39271 );
and \U$41457 ( \41436 , \41435 , \39287 );
and \U$41458 ( \41437 , \39265 , \39271 );
or \U$41459 ( \41438 , \41436 , \41437 );
buf \U$41460 ( \41439 , \41438 );
buf \U$41461 ( \41440 , \41439 );
buf \U$41462 ( \41441 , \39359 );
not \U$41463 ( \41442 , \41441 );
buf \U$41464 ( \41443 , \41442 );
not \U$41465 ( \41444 , \41443 );
buf \U$41466 ( \41445 , \39413 );
not \U$41467 ( \41446 , \41445 );
buf \U$41468 ( \41447 , \41446 );
not \U$41469 ( \41448 , \41447 );
or \U$41470 ( \41449 , \41444 , \41448 );
not \U$41471 ( \41450 , \39413 );
not \U$41472 ( \41451 , \39359 );
or \U$41473 ( \41452 , \41450 , \41451 );
nand \U$41474 ( \41453 , \41452 , \39366 );
nand \U$41475 ( \41454 , \41449 , \41453 );
buf \U$41476 ( \41455 , \41454 );
xor \U$41477 ( \41456 , \41440 , \41455 );
buf \U$41478 ( \41457 , \40685 );
not \U$41479 ( \41458 , \41457 );
buf \U$41480 ( \41459 , \41458 );
buf \U$41481 ( \41460 , \41459 );
not \U$41482 ( \41461 , \41460 );
buf \U$41483 ( \41462 , \40646 );
not \U$41484 ( \41463 , \41462 );
buf \U$41485 ( \41464 , \40665 );
not \U$41486 ( \41465 , \41464 );
or \U$41487 ( \41466 , \41463 , \41465 );
buf \U$41488 ( \41467 , \40665 );
buf \U$41489 ( \41468 , \40646 );
or \U$41490 ( \41469 , \41467 , \41468 );
nand \U$41491 ( \41470 , \41466 , \41469 );
buf \U$41492 ( \41471 , \41470 );
buf \U$41493 ( \41472 , \41471 );
not \U$41494 ( \41473 , \41472 );
or \U$41495 ( \41474 , \41461 , \41473 );
buf \U$41496 ( \41475 , \41471 );
buf \U$41497 ( \41476 , \41459 );
or \U$41498 ( \41477 , \41475 , \41476 );
nand \U$41499 ( \41478 , \41474 , \41477 );
buf \U$41500 ( \41479 , \41478 );
buf \U$41501 ( \41480 , \41479 );
and \U$41502 ( \41481 , \41456 , \41480 );
and \U$41503 ( \41482 , \41440 , \41455 );
or \U$41504 ( \41483 , \41481 , \41482 );
buf \U$41505 ( \41484 , \41483 );
buf \U$41506 ( \41485 , \41484 );
xor \U$41507 ( \41486 , \41434 , \41485 );
buf \U$41508 ( \41487 , \41486 );
buf \U$41509 ( \41488 , \41487 );
xor \U$41510 ( \41489 , \41254 , \41488 );
and \U$41511 ( \41490 , \41410 , \41414 );
not \U$41512 ( \41491 , \41410 );
and \U$41513 ( \41492 , \41491 , \41417 );
nor \U$41514 ( \41493 , \41490 , \41492 );
xor \U$41515 ( \41494 , \41493 , \41426 );
buf \U$41516 ( \41495 , \41494 );
not \U$41517 ( \41496 , \41495 );
buf \U$41518 ( \41497 , \41496 );
buf \U$41519 ( \41498 , \41497 );
not \U$41520 ( \41499 , \41498 );
xor \U$41521 ( \41500 , \39290 , \39296 );
and \U$41522 ( \41501 , \41500 , \39430 );
and \U$41523 ( \41502 , \39290 , \39296 );
or \U$41524 ( \41503 , \41501 , \41502 );
buf \U$41525 ( \41504 , \41503 );
buf \U$41526 ( \41505 , \41504 );
not \U$41527 ( \41506 , \41505 );
or \U$41528 ( \41507 , \41499 , \41506 );
buf \U$41529 ( \41508 , \41504 );
buf \U$41530 ( \41509 , \41497 );
or \U$41531 ( \41510 , \41508 , \41509 );
buf \U$41532 ( \41511 , \39449 );
not \U$41533 ( \41512 , \41511 );
buf \U$41534 ( \41513 , \41512 );
buf \U$41535 ( \41514 , \41513 );
not \U$41536 ( \41515 , \41514 );
buf \U$41537 ( \41516 , \39785 );
not \U$41538 ( \41517 , \41516 );
or \U$41539 ( \41518 , \41515 , \41517 );
buf \U$41540 ( \41519 , \39791 );
nand \U$41541 ( \41520 , \41518 , \41519 );
buf \U$41542 ( \41521 , \41520 );
buf \U$41543 ( \41522 , \41521 );
buf \U$41544 ( \41523 , \39785 );
not \U$41545 ( \41524 , \41523 );
buf \U$41546 ( \41525 , \39449 );
nand \U$41547 ( \41526 , \41524 , \41525 );
buf \U$41548 ( \41527 , \41526 );
buf \U$41549 ( \41528 , \41527 );
nand \U$41550 ( \41529 , \41522 , \41528 );
buf \U$41551 ( \41530 , \41529 );
buf \U$41552 ( \41531 , \41530 );
nand \U$41553 ( \41532 , \41510 , \41531 );
buf \U$41554 ( \41533 , \41532 );
buf \U$41555 ( \41534 , \41533 );
nand \U$41556 ( \41535 , \41507 , \41534 );
buf \U$41557 ( \41536 , \41535 );
buf \U$41558 ( \41537 , \41536 );
xor \U$41559 ( \41538 , \41489 , \41537 );
buf \U$41560 ( \41539 , \41538 );
buf \U$41561 ( \41540 , \41539 );
buf \U$41562 ( \41541 , \41494 );
not \U$41563 ( \41542 , \41541 );
buf \U$41564 ( \41543 , \41530 );
not \U$41565 ( \41544 , \41543 );
and \U$41566 ( \41545 , \41542 , \41544 );
buf \U$41567 ( \41546 , \41494 );
buf \U$41568 ( \41547 , \41530 );
and \U$41569 ( \41548 , \41546 , \41547 );
nor \U$41570 ( \41549 , \41545 , \41548 );
buf \U$41571 ( \41550 , \41549 );
buf \U$41572 ( \41551 , \41550 );
not \U$41573 ( \41552 , \41551 );
buf \U$41574 ( \41553 , \41504 );
not \U$41575 ( \41554 , \41553 );
and \U$41576 ( \41555 , \41552 , \41554 );
buf \U$41577 ( \41556 , \41504 );
buf \U$41578 ( \41557 , \41550 );
and \U$41579 ( \41558 , \41556 , \41557 );
nor \U$41580 ( \41559 , \41555 , \41558 );
buf \U$41581 ( \41560 , \41559 );
buf \U$41582 ( \41561 , \41560 );
not \U$41583 ( \41562 , \41561 );
buf \U$41584 ( \41563 , \41562 );
buf \U$41585 ( \41564 , \41563 );
xor \U$41586 ( \41565 , \41440 , \41455 );
xor \U$41587 ( \41566 , \41565 , \41480 );
buf \U$41588 ( \41567 , \41566 );
buf \U$41589 ( \41568 , \41567 );
or \U$41590 ( \41569 , \41564 , \41568 );
buf \U$41591 ( \41570 , \39792 );
not \U$41592 ( \41571 , \41570 );
buf \U$41593 ( \41572 , \41571 );
buf \U$41594 ( \41573 , \41572 );
not \U$41595 ( \41574 , \41573 );
buf \U$41596 ( \41575 , \39808 );
not \U$41597 ( \41576 , \41575 );
or \U$41598 ( \41577 , \41574 , \41576 );
buf \U$41599 ( \41578 , \39792 );
not \U$41600 ( \41579 , \41578 );
buf \U$41601 ( \41580 , \39808 );
not \U$41602 ( \41581 , \41580 );
buf \U$41603 ( \41582 , \41581 );
buf \U$41604 ( \41583 , \41582 );
not \U$41605 ( \41584 , \41583 );
or \U$41606 ( \41585 , \41579 , \41584 );
buf \U$41607 ( \41586 , \39822 );
nand \U$41608 ( \41587 , \41585 , \41586 );
buf \U$41609 ( \41588 , \41587 );
buf \U$41610 ( \41589 , \41588 );
nand \U$41611 ( \41590 , \41577 , \41589 );
buf \U$41612 ( \41591 , \41590 );
buf \U$41613 ( \41592 , \41591 );
nand \U$41614 ( \41593 , \41569 , \41592 );
buf \U$41615 ( \41594 , \41593 );
buf \U$41616 ( \41595 , \41594 );
buf \U$41617 ( \41596 , \41563 );
buf \U$41618 ( \41597 , \41567 );
nand \U$41619 ( \41598 , \41596 , \41597 );
buf \U$41620 ( \41599 , \41598 );
buf \U$41621 ( \41600 , \41599 );
nand \U$41622 ( \41601 , \41595 , \41600 );
buf \U$41623 ( \41602 , \41601 );
buf \U$41624 ( \41603 , \41602 );
nor \U$41625 ( \41604 , \41540 , \41603 );
buf \U$41626 ( \41605 , \41604 );
buf \U$41627 ( \41606 , \41605 );
not \U$41628 ( \41607 , \41606 );
buf \U$41629 ( \41608 , \39832 );
not \U$41630 ( \41609 , \41608 );
buf \U$41631 ( \41610 , \41609 );
buf \U$41632 ( \41611 , \41610 );
buf \U$41633 ( \41612 , \39432 );
or \U$41634 ( \41613 , \41611 , \41612 );
buf \U$41635 ( \41614 , \39851 );
nand \U$41636 ( \41615 , \41613 , \41614 );
buf \U$41637 ( \41616 , \41615 );
buf \U$41638 ( \41617 , \41616 );
buf \U$41639 ( \41618 , \41610 );
buf \U$41640 ( \41619 , \39432 );
nand \U$41641 ( \41620 , \41618 , \41619 );
buf \U$41642 ( \41621 , \41620 );
buf \U$41643 ( \41622 , \41621 );
nand \U$41644 ( \41623 , \41617 , \41622 );
buf \U$41645 ( \41624 , \41623 );
buf \U$41646 ( \41625 , \41624 );
not \U$41647 ( \41626 , \41625 );
xor \U$41648 ( \41627 , \41567 , \41560 );
xor \U$41649 ( \41628 , \41627 , \41591 );
buf \U$41650 ( \41629 , \41628 );
nand \U$41651 ( \41630 , \41626 , \41629 );
buf \U$41652 ( \41631 , \41630 );
buf \U$41653 ( \41632 , \41631 );
nand \U$41654 ( \41633 , \41607 , \41632 );
buf \U$41655 ( \41634 , \41633 );
buf \U$41656 ( \41635 , \41634 );
nor \U$41657 ( \41636 , \40148 , \41635 );
buf \U$41658 ( \41637 , \41636 );
buf \U$41659 ( \41638 , \41637 );
xor \U$41660 ( \41639 , \40109 , \40113 );
xor \U$41661 ( \41640 , \41639 , \40118 );
buf \U$41662 ( \41641 , \41640 );
xor \U$41663 ( \41642 , \34342 , \34473 );
and \U$41664 ( \41643 , \41642 , \34480 );
and \U$41665 ( \41644 , \34342 , \34473 );
or \U$41666 ( \41645 , \41643 , \41644 );
buf \U$41667 ( \41646 , \41645 );
buf \U$41668 ( \41647 , \41646 );
not \U$41669 ( \41648 , \41647 );
not \U$41670 ( \41649 , \33753 );
not \U$41671 ( \41650 , \33644 );
or \U$41672 ( \41651 , \41649 , \41650 );
not \U$41673 ( \41652 , \33647 );
not \U$41674 ( \41653 , \33750 );
or \U$41675 ( \41654 , \41652 , \41653 );
nand \U$41676 ( \41655 , \41654 , \33769 );
nand \U$41677 ( \41656 , \41651 , \41655 );
buf \U$41678 ( \41657 , \41656 );
not \U$41679 ( \41658 , \41657 );
or \U$41680 ( \41659 , \41648 , \41658 );
buf \U$41681 ( \41660 , \41656 );
buf \U$41682 ( \41661 , \41646 );
or \U$41683 ( \41662 , \41660 , \41661 );
and \U$41684 ( \41663 , \39973 , \39952 );
not \U$41685 ( \41664 , \39973 );
and \U$41686 ( \41665 , \41664 , \39949 );
or \U$41687 ( \41666 , \41663 , \41665 );
buf \U$41688 ( \41667 , \41666 );
buf \U$41689 ( \41668 , \39980 );
and \U$41690 ( \41669 , \41667 , \41668 );
not \U$41691 ( \41670 , \41667 );
buf \U$41692 ( \41671 , \39932 );
and \U$41693 ( \41672 , \41670 , \41671 );
nor \U$41694 ( \41673 , \41669 , \41672 );
buf \U$41695 ( \41674 , \41673 );
buf \U$41696 ( \41675 , \41674 );
nand \U$41697 ( \41676 , \41662 , \41675 );
buf \U$41698 ( \41677 , \41676 );
buf \U$41699 ( \41678 , \41677 );
nand \U$41700 ( \41679 , \41659 , \41678 );
buf \U$41701 ( \41680 , \41679 );
xor \U$41702 ( \41681 , \39987 , \39929 );
buf \U$41703 ( \41682 , \41681 );
not \U$41704 ( \41683 , \41682 );
buf \U$41705 ( \41684 , \40059 );
not \U$41706 ( \41685 , \41684 );
and \U$41707 ( \41686 , \41683 , \41685 );
buf \U$41708 ( \41687 , \40059 );
buf \U$41709 ( \41688 , \41681 );
and \U$41710 ( \41689 , \41687 , \41688 );
nor \U$41711 ( \41690 , \41686 , \41689 );
buf \U$41712 ( \41691 , \41690 );
xor \U$41713 ( \41692 , \41680 , \41691 );
xor \U$41714 ( \41693 , \33798 , \33874 );
and \U$41715 ( \41694 , \41693 , \34130 );
and \U$41716 ( \41695 , \33798 , \33874 );
or \U$41717 ( \41696 , \41694 , \41695 );
buf \U$41718 ( \41697 , \41696 );
buf \U$41719 ( \41698 , \41697 );
not \U$41720 ( \41699 , \41698 );
buf \U$41721 ( \41700 , \40015 );
not \U$41722 ( \41701 , \41700 );
buf \U$41723 ( \41702 , \40020 );
not \U$41724 ( \41703 , \41702 );
or \U$41725 ( \41704 , \41701 , \41703 );
buf \U$41726 ( \41705 , \40015 );
buf \U$41727 ( \41706 , \40020 );
or \U$41728 ( \41707 , \41705 , \41706 );
nand \U$41729 ( \41708 , \41704 , \41707 );
buf \U$41730 ( \41709 , \41708 );
buf \U$41731 ( \41710 , \41709 );
buf \U$41732 ( \41711 , \40048 );
xor \U$41733 ( \41712 , \41710 , \41711 );
buf \U$41734 ( \41713 , \41712 );
buf \U$41735 ( \41714 , \41713 );
not \U$41736 ( \41715 , \41714 );
or \U$41737 ( \41716 , \41699 , \41715 );
buf \U$41738 ( \41717 , \41697 );
buf \U$41739 ( \41718 , \41713 );
or \U$41740 ( \41719 , \41717 , \41718 );
xor \U$41741 ( \41720 , \40097 , \40078 );
xor \U$41742 ( \41721 , \41720 , \40074 );
buf \U$41743 ( \41722 , \41721 );
nand \U$41744 ( \41723 , \41719 , \41722 );
buf \U$41745 ( \41724 , \41723 );
buf \U$41746 ( \41725 , \41724 );
nand \U$41747 ( \41726 , \41716 , \41725 );
buf \U$41748 ( \41727 , \41726 );
xor \U$41749 ( \41728 , \41692 , \41727 );
xor \U$41750 ( \41729 , \41641 , \41728 );
buf \U$41751 ( \41730 , \41674 );
not \U$41752 ( \41731 , \41730 );
buf \U$41753 ( \41732 , \41646 );
not \U$41754 ( \41733 , \41732 );
buf \U$41755 ( \41734 , \41733 );
buf \U$41756 ( \41735 , \41734 );
not \U$41757 ( \41736 , \41735 );
or \U$41758 ( \41737 , \41731 , \41736 );
buf \U$41759 ( \41738 , \41646 );
buf \U$41760 ( \41739 , \41674 );
not \U$41761 ( \41740 , \41739 );
buf \U$41762 ( \41741 , \41740 );
buf \U$41763 ( \41742 , \41741 );
nand \U$41764 ( \41743 , \41738 , \41742 );
buf \U$41765 ( \41744 , \41743 );
buf \U$41766 ( \41745 , \41744 );
nand \U$41767 ( \41746 , \41737 , \41745 );
buf \U$41768 ( \41747 , \41746 );
buf \U$41769 ( \41748 , \41747 );
buf \U$41770 ( \41749 , \41656 );
not \U$41771 ( \41750 , \41749 );
buf \U$41772 ( \41751 , \41750 );
buf \U$41773 ( \41752 , \41751 );
and \U$41774 ( \41753 , \41748 , \41752 );
not \U$41775 ( \41754 , \41748 );
buf \U$41776 ( \41755 , \41656 );
and \U$41777 ( \41756 , \41754 , \41755 );
nor \U$41778 ( \41757 , \41753 , \41756 );
buf \U$41779 ( \41758 , \41757 );
buf \U$41780 ( \41759 , \41758 );
not \U$41781 ( \41760 , \41759 );
buf \U$41782 ( \41761 , \41760 );
buf \U$41783 ( \41762 , \41761 );
not \U$41784 ( \41763 , \41762 );
buf \U$41785 ( \41764 , \33626 );
not \U$41786 ( \41765 , \41764 );
buf \U$41787 ( \41766 , \33772 );
not \U$41788 ( \41767 , \41766 );
buf \U$41789 ( \41768 , \41767 );
buf \U$41790 ( \41769 , \41768 );
not \U$41791 ( \41770 , \41769 );
or \U$41792 ( \41771 , \41765 , \41770 );
buf \U$41793 ( \41772 , \41768 );
buf \U$41794 ( \41773 , \33626 );
or \U$41795 ( \41774 , \41772 , \41773 );
buf \U$41796 ( \41775 , \34132 );
nand \U$41797 ( \41776 , \41774 , \41775 );
buf \U$41798 ( \41777 , \41776 );
buf \U$41799 ( \41778 , \41777 );
nand \U$41800 ( \41779 , \41771 , \41778 );
buf \U$41801 ( \41780 , \41779 );
buf \U$41802 ( \41781 , \41780 );
not \U$41803 ( \41782 , \41781 );
or \U$41804 ( \41783 , \41763 , \41782 );
buf \U$41805 ( \41784 , \41780 );
buf \U$41806 ( \41785 , \41761 );
or \U$41807 ( \41786 , \41784 , \41785 );
xor \U$41808 ( \41787 , \34143 , \34161 );
and \U$41809 ( \41788 , \41787 , \34483 );
and \U$41810 ( \41789 , \34143 , \34161 );
or \U$41811 ( \41790 , \41788 , \41789 );
buf \U$41812 ( \41791 , \41790 );
buf \U$41813 ( \41792 , \41791 );
nand \U$41814 ( \41793 , \41786 , \41792 );
buf \U$41815 ( \41794 , \41793 );
buf \U$41816 ( \41795 , \41794 );
nand \U$41817 ( \41796 , \41783 , \41795 );
buf \U$41818 ( \41797 , \41796 );
xor \U$41819 ( \41798 , \41729 , \41797 );
buf \U$41820 ( \41799 , \41798 );
xor \U$41821 ( \41800 , \41697 , \41713 );
buf \U$41822 ( \41801 , \41800 );
buf \U$41823 ( \41802 , \41721 );
not \U$41824 ( \41803 , \41802 );
buf \U$41825 ( \41804 , \41803 );
buf \U$41826 ( \41805 , \41804 );
and \U$41827 ( \41806 , \41801 , \41805 );
not \U$41828 ( \41807 , \41801 );
buf \U$41829 ( \41808 , \41721 );
and \U$41830 ( \41809 , \41807 , \41808 );
nor \U$41831 ( \41810 , \41806 , \41809 );
buf \U$41832 ( \41811 , \41810 );
buf \U$41833 ( \41812 , \41811 );
buf \U$41834 ( \41813 , \34495 );
not \U$41835 ( \41814 , \41813 );
buf \U$41836 ( \41815 , \34485 );
not \U$41837 ( \41816 , \41815 );
buf \U$41838 ( \41817 , \41816 );
buf \U$41839 ( \41818 , \41817 );
not \U$41840 ( \41819 , \41818 );
or \U$41841 ( \41820 , \41814 , \41819 );
buf \U$41842 ( \41821 , \34509 );
nand \U$41843 ( \41822 , \41820 , \41821 );
buf \U$41844 ( \41823 , \41822 );
buf \U$41845 ( \41824 , \41823 );
buf \U$41846 ( \41825 , \41817 );
not \U$41847 ( \41826 , \41825 );
buf \U$41848 ( \41827 , \34492 );
nand \U$41849 ( \41828 , \41826 , \41827 );
buf \U$41850 ( \41829 , \41828 );
buf \U$41851 ( \41830 , \41829 );
and \U$41852 ( \41831 , \41824 , \41830 );
buf \U$41853 ( \41832 , \41831 );
buf \U$41854 ( \41833 , \41832 );
xor \U$41855 ( \41834 , \41812 , \41833 );
buf \U$41856 ( \41835 , \41791 );
not \U$41857 ( \41836 , \41835 );
buf \U$41858 ( \41837 , \41758 );
not \U$41859 ( \41838 , \41837 );
or \U$41860 ( \41839 , \41836 , \41838 );
buf \U$41861 ( \41840 , \41758 );
buf \U$41862 ( \41841 , \41791 );
or \U$41863 ( \41842 , \41840 , \41841 );
nand \U$41864 ( \41843 , \41839 , \41842 );
buf \U$41865 ( \41844 , \41843 );
buf \U$41866 ( \41845 , \41844 );
buf \U$41867 ( \41846 , \41780 );
not \U$41868 ( \41847 , \41846 );
buf \U$41869 ( \41848 , \41847 );
buf \U$41870 ( \41849 , \41848 );
and \U$41871 ( \41850 , \41845 , \41849 );
not \U$41872 ( \41851 , \41845 );
buf \U$41873 ( \41852 , \41780 );
and \U$41874 ( \41853 , \41851 , \41852 );
nor \U$41875 ( \41854 , \41850 , \41853 );
buf \U$41876 ( \41855 , \41854 );
buf \U$41877 ( \41856 , \41855 );
and \U$41878 ( \41857 , \41834 , \41856 );
and \U$41879 ( \41858 , \41812 , \41833 );
or \U$41880 ( \41859 , \41857 , \41858 );
buf \U$41881 ( \41860 , \41859 );
buf \U$41882 ( \41861 , \41860 );
nand \U$41883 ( \41862 , \41799 , \41861 );
buf \U$41884 ( \41863 , \41862 );
buf \U$41885 ( \41864 , \41863 );
buf \U$41886 ( \41865 , \34135 );
not \U$41887 ( \41866 , \41865 );
buf \U$41888 ( \41867 , \41866 );
buf \U$41889 ( \41868 , \41867 );
not \U$41890 ( \41869 , \41868 );
buf \U$41891 ( \41870 , \34519 );
not \U$41892 ( \41871 , \41870 );
or \U$41893 ( \41872 , \41869 , \41871 );
buf \U$41894 ( \41873 , \34544 );
nand \U$41895 ( \41874 , \41872 , \41873 );
buf \U$41896 ( \41875 , \41874 );
buf \U$41897 ( \41876 , \41875 );
buf \U$41898 ( \41877 , \34519 );
not \U$41899 ( \41878 , \41877 );
buf \U$41900 ( \41879 , \34135 );
nand \U$41901 ( \41880 , \41878 , \41879 );
buf \U$41902 ( \41881 , \41880 );
buf \U$41903 ( \41882 , \41881 );
nand \U$41904 ( \41883 , \41876 , \41882 );
buf \U$41905 ( \41884 , \41883 );
buf \U$41906 ( \41885 , \41884 );
not \U$41907 ( \41886 , \41885 );
xor \U$41908 ( \41887 , \41812 , \41833 );
xor \U$41909 ( \41888 , \41887 , \41856 );
buf \U$41910 ( \41889 , \41888 );
buf \U$41911 ( \41890 , \41889 );
nand \U$41912 ( \41891 , \41886 , \41890 );
buf \U$41913 ( \41892 , \41891 );
buf \U$41914 ( \41893 , \41892 );
and \U$41915 ( \41894 , \41864 , \41893 );
buf \U$41916 ( \41895 , \41894 );
buf \U$41917 ( \41896 , \41895 );
xor \U$41918 ( \41897 , \39867 , \39911 );
xor \U$41919 ( \41898 , \41897 , \39916 );
buf \U$41920 ( \41899 , \41898 );
xor \U$41921 ( \41900 , \39926 , \40070 );
xor \U$41922 ( \41901 , \41900 , \40123 );
buf \U$41923 ( \41902 , \41901 );
or \U$41924 ( \41903 , \41899 , \41902 );
buf \U$41925 ( \41904 , \41691 );
not \U$41926 ( \41905 , \41904 );
buf \U$41927 ( \41906 , \41905 );
buf \U$41928 ( \41907 , \41906 );
not \U$41929 ( \41908 , \41907 );
buf \U$41930 ( \41909 , \41680 );
not \U$41931 ( \41910 , \41909 );
or \U$41932 ( \41911 , \41908 , \41910 );
buf \U$41933 ( \41912 , \41691 );
not \U$41934 ( \41913 , \41912 );
buf \U$41935 ( \41914 , \41680 );
not \U$41936 ( \41915 , \41914 );
buf \U$41937 ( \41916 , \41915 );
buf \U$41938 ( \41917 , \41916 );
not \U$41939 ( \41918 , \41917 );
or \U$41940 ( \41919 , \41913 , \41918 );
buf \U$41941 ( \41920 , \41727 );
nand \U$41942 ( \41921 , \41919 , \41920 );
buf \U$41943 ( \41922 , \41921 );
buf \U$41944 ( \41923 , \41922 );
nand \U$41945 ( \41924 , \41911 , \41923 );
buf \U$41946 ( \41925 , \41924 );
nand \U$41947 ( \41926 , \41903 , \41925 );
buf \U$41948 ( \41927 , \41926 );
buf \U$41949 ( \41928 , \41902 );
buf \U$41950 ( \41929 , \41899 );
nand \U$41951 ( \41930 , \41928 , \41929 );
buf \U$41952 ( \41931 , \41930 );
buf \U$41953 ( \41932 , \41931 );
nand \U$41954 ( \41933 , \41927 , \41932 );
buf \U$41955 ( \41934 , \41933 );
buf \U$41956 ( \41935 , \41934 );
not \U$41957 ( \41936 , \41935 );
buf \U$41958 ( \41937 , \39920 );
buf \U$41959 ( \41938 , \40127 );
xor \U$41960 ( \41939 , \41937 , \41938 );
buf \U$41961 ( \41940 , \39862 );
xnor \U$41962 ( \41941 , \41939 , \41940 );
buf \U$41963 ( \41942 , \41941 );
buf \U$41964 ( \41943 , \41942 );
nand \U$41965 ( \41944 , \41936 , \41943 );
buf \U$41966 ( \41945 , \41944 );
buf \U$41967 ( \41946 , \41945 );
not \U$41968 ( \41947 , \41641 );
nand \U$41969 ( \41948 , \41947 , \41728 );
not \U$41970 ( \41949 , \41948 );
not \U$41971 ( \41950 , \41797 );
or \U$41972 ( \41951 , \41949 , \41950 );
buf \U$41973 ( \41952 , \41728 );
not \U$41974 ( \41953 , \41952 );
buf \U$41975 ( \41954 , \41641 );
nand \U$41976 ( \41955 , \41953 , \41954 );
buf \U$41977 ( \41956 , \41955 );
nand \U$41978 ( \41957 , \41951 , \41956 );
buf \U$41979 ( \41958 , \41957 );
not \U$41980 ( \41959 , \41958 );
buf \U$41981 ( \41960 , \41899 );
buf \U$41982 ( \41961 , \41925 );
xor \U$41983 ( \41962 , \41960 , \41961 );
buf \U$41984 ( \41963 , \41902 );
xnor \U$41985 ( \41964 , \41962 , \41963 );
buf \U$41986 ( \41965 , \41964 );
buf \U$41987 ( \41966 , \41965 );
nand \U$41988 ( \41967 , \41959 , \41966 );
buf \U$41989 ( \41968 , \41967 );
buf \U$41990 ( \41969 , \41968 );
and \U$41991 ( \41970 , \41638 , \41896 , \41946 , \41969 );
buf \U$41992 ( \41971 , \41970 );
buf \U$41993 ( \41972 , \41971 );
xor \U$41994 ( \41973 , \41254 , \41488 );
and \U$41995 ( \41974 , \41973 , \41537 );
and \U$41996 ( \41975 , \41254 , \41488 );
or \U$41997 ( \41976 , \41974 , \41975 );
buf \U$41998 ( \41977 , \41976 );
buf \U$41999 ( \41978 , \41977 );
not \U$42000 ( \41979 , \41978 );
xor \U$42001 ( \41980 , \40358 , \40581 );
and \U$42002 ( \41981 , \41980 , \40629 );
and \U$42003 ( \41982 , \40358 , \40581 );
or \U$42004 ( \41983 , \41981 , \41982 );
buf \U$42005 ( \41984 , \41983 );
buf \U$42006 ( \41985 , \41984 );
and \U$42007 ( \41986 , \40382 , \40383 );
buf \U$42008 ( \41987 , \41986 );
buf \U$42009 ( \41988 , \41987 );
buf \U$42010 ( \41989 , \812 );
not \U$42011 ( \41990 , \41989 );
buf \U$42012 ( \41991 , \40464 );
not \U$42013 ( \41992 , \41991 );
and \U$42014 ( \41993 , \41990 , \41992 );
buf \U$42015 ( \41994 , \816 );
buf \U$42016 ( \41995 , \4524 );
and \U$42017 ( \41996 , \41994 , \41995 );
buf \U$42018 ( \41997 , \41996 );
buf \U$42019 ( \41998 , \41997 );
nor \U$42020 ( \41999 , \41993 , \41998 );
buf \U$42021 ( \42000 , \41999 );
buf \U$42022 ( \42001 , \42000 );
xor \U$42023 ( \42002 , \41988 , \42001 );
buf \U$42024 ( \42003 , \954 );
buf \U$42025 ( \42004 , \40712 );
or \U$42026 ( \42005 , \42003 , \42004 );
buf \U$42027 ( \42006 , \2963 );
buf \U$42028 ( \42007 , RIc0d9dd8_85);
buf \U$42029 ( \42008 , RIc0d7e70_18);
and \U$42030 ( \42009 , \42007 , \42008 );
not \U$42031 ( \42010 , \42007 );
buf \U$42032 ( \42011 , \7820 );
and \U$42033 ( \42012 , \42010 , \42011 );
nor \U$42034 ( \42013 , \42009 , \42012 );
buf \U$42035 ( \42014 , \42013 );
buf \U$42036 ( \42015 , \42014 );
not \U$42037 ( \42016 , \42015 );
buf \U$42038 ( \42017 , \42016 );
buf \U$42039 ( \42018 , \42017 );
or \U$42040 ( \42019 , \42006 , \42018 );
nand \U$42041 ( \42020 , \42005 , \42019 );
buf \U$42042 ( \42021 , \42020 );
buf \U$42043 ( \42022 , \42021 );
xor \U$42044 ( \42023 , \42002 , \42022 );
buf \U$42045 ( \42024 , \42023 );
buf \U$42046 ( \42025 , \42024 );
buf \U$42047 ( \42026 , \397 );
not \U$42048 ( \42027 , \42026 );
buf \U$42049 ( \42028 , \42027 );
buf \U$42050 ( \42029 , \42028 );
buf \U$42051 ( \42030 , \40316 );
or \U$42052 ( \42031 , \42029 , \42030 );
buf \U$42053 ( \42032 , \8178 );
buf \U$42054 ( \42033 , \4501 );
or \U$42055 ( \42034 , \42032 , \42033 );
nand \U$42056 ( \42035 , \42031 , \42034 );
buf \U$42057 ( \42036 , \42035 );
buf \U$42058 ( \42037 , \42036 );
buf \U$42059 ( \42038 , \4043 );
not \U$42060 ( \42039 , \42038 );
buf \U$42061 ( \42040 , \42039 );
buf \U$42062 ( \42041 , \42040 );
buf \U$42063 ( \42042 , \40204 );
or \U$42064 ( \42043 , \42041 , \42042 );
buf \U$42065 ( \42044 , \36639 );
buf \U$42066 ( \42045 , RIc0d76f0_2);
buf \U$42067 ( \42046 , RIc0da558_101);
xor \U$42068 ( \42047 , \42045 , \42046 );
buf \U$42069 ( \42048 , \42047 );
buf \U$42070 ( \42049 , \42048 );
not \U$42071 ( \42050 , \42049 );
buf \U$42072 ( \42051 , \42050 );
buf \U$42073 ( \42052 , \42051 );
or \U$42074 ( \42053 , \42044 , \42052 );
nand \U$42075 ( \42054 , \42043 , \42053 );
buf \U$42076 ( \42055 , \42054 );
buf \U$42077 ( \42056 , \42055 );
xor \U$42078 ( \42057 , \42037 , \42056 );
buf \U$42079 ( \42058 , \333 );
buf \U$42080 ( \42059 , \40570 );
or \U$42081 ( \42060 , \42058 , \42059 );
buf \U$42082 ( \42061 , \4849 );
buf \U$42083 ( \42062 , \4452 );
not \U$42084 ( \42063 , \42062 );
buf \U$42085 ( \42064 , \42063 );
buf \U$42086 ( \42065 , \42064 );
or \U$42087 ( \42066 , \42061 , \42065 );
nand \U$42088 ( \42067 , \42060 , \42066 );
buf \U$42089 ( \42068 , \42067 );
buf \U$42090 ( \42069 , \42068 );
xor \U$42091 ( \42070 , \42057 , \42069 );
buf \U$42092 ( \42071 , \42070 );
buf \U$42093 ( \42072 , \42071 );
xor \U$42094 ( \42073 , \42025 , \42072 );
xor \U$42095 ( \42074 , \40997 , \41051 );
and \U$42096 ( \42075 , \42074 , \41104 );
and \U$42097 ( \42076 , \40997 , \41051 );
or \U$42098 ( \42077 , \42075 , \42076 );
buf \U$42099 ( \42078 , \42077 );
buf \U$42100 ( \42079 , \42078 );
xor \U$42101 ( \42080 , \42073 , \42079 );
buf \U$42102 ( \42081 , \42080 );
buf \U$42103 ( \42082 , \42081 );
xor \U$42104 ( \42083 , \41326 , \41348 );
and \U$42105 ( \42084 , \42083 , \41371 );
and \U$42106 ( \42085 , \41326 , \41348 );
or \U$42107 ( \42086 , \42084 , \42085 );
buf \U$42108 ( \42087 , \42086 );
buf \U$42109 ( \42088 , \42087 );
xor \U$42110 ( \42089 , \42082 , \42088 );
buf \U$42111 ( \42090 , \40962 );
buf \U$42112 ( \42091 , \40796 );
or \U$42113 ( \42092 , \42090 , \42091 );
buf \U$42114 ( \42093 , \40962 );
not \U$42115 ( \42094 , \42093 );
buf \U$42116 ( \42095 , \40796 );
not \U$42117 ( \42096 , \42095 );
or \U$42118 ( \42097 , \42094 , \42096 );
buf \U$42119 ( \42098 , \40830 );
nand \U$42120 ( \42099 , \42097 , \42098 );
buf \U$42121 ( \42100 , \42099 );
buf \U$42122 ( \42101 , \42100 );
nand \U$42123 ( \42102 , \42092 , \42101 );
buf \U$42124 ( \42103 , \42102 );
buf \U$42125 ( \42104 , \42103 );
xor \U$42126 ( \42105 , \41332 , \41338 );
and \U$42127 ( \42106 , \42105 , \41345 );
and \U$42128 ( \42107 , \41332 , \41338 );
or \U$42129 ( \42108 , \42106 , \42107 );
buf \U$42130 ( \42109 , \42108 );
buf \U$42131 ( \42110 , \42109 );
xor \U$42132 ( \42111 , \42104 , \42110 );
xor \U$42133 ( \42112 , \40425 , \40501 );
and \U$42134 ( \42113 , \42112 , \40578 );
and \U$42135 ( \42114 , \40425 , \40501 );
or \U$42136 ( \42115 , \42113 , \42114 );
buf \U$42137 ( \42116 , \42115 );
buf \U$42138 ( \42117 , \42116 );
xor \U$42139 ( \42118 , \42111 , \42117 );
buf \U$42140 ( \42119 , \42118 );
buf \U$42141 ( \42120 , \42119 );
xor \U$42142 ( \42121 , \42089 , \42120 );
buf \U$42143 ( \42122 , \42121 );
buf \U$42144 ( \42123 , \42122 );
xor \U$42145 ( \42124 , \41985 , \42123 );
xor \U$42146 ( \42125 , \40884 , \40984 );
and \U$42147 ( \42126 , \42125 , \41248 );
and \U$42148 ( \42127 , \40884 , \40984 );
or \U$42149 ( \42128 , \42126 , \42127 );
buf \U$42150 ( \42129 , \42128 );
buf \U$42151 ( \42130 , \42129 );
xor \U$42152 ( \42131 , \42124 , \42130 );
buf \U$42153 ( \42132 , \42131 );
buf \U$42154 ( \42133 , \42132 );
xor \U$42155 ( \42134 , \41320 , \41374 );
and \U$42156 ( \42135 , \42134 , \41404 );
and \U$42157 ( \42136 , \41320 , \41374 );
or \U$42158 ( \42137 , \42135 , \42136 );
buf \U$42159 ( \42138 , \42137 );
buf \U$42160 ( \42139 , \42138 );
xor \U$42161 ( \42140 , \40991 , \41107 );
and \U$42162 ( \42141 , \42140 , \41245 );
and \U$42163 ( \42142 , \40991 , \41107 );
or \U$42164 ( \42143 , \42141 , \42142 );
buf \U$42165 ( \42144 , \42143 );
buf \U$42166 ( \42145 , \42144 );
buf \U$42167 ( \42146 , \40274 );
not \U$42168 ( \42147 , \42146 );
buf \U$42169 ( \42148 , \40217 );
not \U$42170 ( \42149 , \42148 );
or \U$42171 ( \42150 , \42147 , \42149 );
not \U$42172 ( \42151 , \40214 );
not \U$42173 ( \42152 , \40271 );
or \U$42174 ( \42153 , \42151 , \42152 );
nand \U$42175 ( \42154 , \42153 , \40354 );
buf \U$42176 ( \42155 , \42154 );
nand \U$42177 ( \42156 , \42150 , \42155 );
buf \U$42178 ( \42157 , \42156 );
buf \U$42179 ( \42158 , \42157 );
buf \U$42180 ( \42159 , \40238 );
buf \U$42181 ( \42160 , \40220 );
or \U$42182 ( \42161 , \42159 , \42160 );
buf \U$42183 ( \42162 , \40268 );
nand \U$42184 ( \42163 , \42161 , \42162 );
buf \U$42185 ( \42164 , \42163 );
buf \U$42186 ( \42165 , \42164 );
buf \U$42187 ( \42166 , \40238 );
buf \U$42188 ( \42167 , \40220 );
nand \U$42189 ( \42168 , \42166 , \42167 );
buf \U$42190 ( \42169 , \42168 );
buf \U$42191 ( \42170 , \42169 );
nand \U$42192 ( \42171 , \42165 , \42170 );
buf \U$42193 ( \42172 , \42171 );
buf \U$42194 ( \42173 , \42172 );
buf \U$42195 ( \42174 , \40186 );
not \U$42196 ( \42175 , \42174 );
buf \U$42197 ( \42176 , \40169 );
not \U$42198 ( \42177 , \42176 );
or \U$42199 ( \42178 , \42175 , \42177 );
buf \U$42200 ( \42179 , \40169 );
buf \U$42201 ( \42180 , \40186 );
or \U$42202 ( \42181 , \42179 , \42180 );
buf \U$42203 ( \42182 , \40212 );
nand \U$42204 ( \42183 , \42181 , \42182 );
buf \U$42205 ( \42184 , \42183 );
buf \U$42206 ( \42185 , \42184 );
nand \U$42207 ( \42186 , \42178 , \42185 );
buf \U$42208 ( \42187 , \42186 );
buf \U$42209 ( \42188 , \42187 );
xor \U$42210 ( \42189 , \42173 , \42188 );
xor \U$42211 ( \42190 , \40447 , \40473 );
and \U$42212 ( \42191 , \42190 , \40498 );
and \U$42213 ( \42192 , \40447 , \40473 );
or \U$42214 ( \42193 , \42191 , \42192 );
buf \U$42215 ( \42194 , \42193 );
buf \U$42216 ( \42195 , \42194 );
xor \U$42217 ( \42196 , \42189 , \42195 );
buf \U$42218 ( \42197 , \42196 );
buf \U$42219 ( \42198 , \42197 );
xor \U$42220 ( \42199 , \42158 , \42198 );
xor \U$42221 ( \42200 , \40303 , \40325 );
and \U$42222 ( \42201 , \42200 , \40352 );
and \U$42223 ( \42202 , \40303 , \40325 );
or \U$42224 ( \42203 , \42201 , \42202 );
buf \U$42225 ( \42204 , \42203 );
buf \U$42226 ( \42205 , \42204 );
xor \U$42227 ( \42206 , \40721 , \40742 );
and \U$42228 ( \42207 , \42206 , \40764 );
and \U$42229 ( \42208 , \40721 , \40742 );
or \U$42230 ( \42209 , \42207 , \42208 );
buf \U$42231 ( \42210 , \42209 );
buf \U$42232 ( \42211 , \42210 );
xor \U$42233 ( \42212 , \42205 , \42211 );
xor \U$42234 ( \42213 , \40519 , \40546 );
and \U$42235 ( \42214 , \42213 , \40575 );
and \U$42236 ( \42215 , \40519 , \40546 );
or \U$42237 ( \42216 , \42214 , \42215 );
buf \U$42238 ( \42217 , \42216 );
buf \U$42239 ( \42218 , \42217 );
xor \U$42240 ( \42219 , \42212 , \42218 );
buf \U$42241 ( \42220 , \42219 );
buf \U$42242 ( \42221 , \42220 );
xor \U$42243 ( \42222 , \42199 , \42221 );
buf \U$42244 ( \42223 , \42222 );
buf \U$42245 ( \42224 , \42223 );
xor \U$42246 ( \42225 , \42145 , \42224 );
buf \U$42247 ( \42226 , \40381 );
not \U$42248 ( \42227 , \42226 );
buf \U$42249 ( \42228 , \40402 );
not \U$42250 ( \42229 , \42228 );
or \U$42251 ( \42230 , \42227 , \42229 );
buf \U$42252 ( \42231 , \40423 );
nand \U$42253 ( \42232 , \42230 , \42231 );
buf \U$42254 ( \42233 , \42232 );
buf \U$42255 ( \42234 , \42233 );
buf \U$42256 ( \42235 , \40399 );
buf \U$42257 ( \42236 , \40378 );
nand \U$42258 ( \42237 , \42235 , \42236 );
buf \U$42259 ( \42238 , \42237 );
buf \U$42260 ( \42239 , \42238 );
nand \U$42261 ( \42240 , \42234 , \42239 );
buf \U$42262 ( \42241 , \42240 );
buf \U$42263 ( \42242 , \42241 );
buf \U$42264 ( \42243 , \40393 );
not \U$42265 ( \42244 , \42243 );
buf \U$42266 ( \42245 , \1224 );
not \U$42267 ( \42246 , \42245 );
or \U$42268 ( \42247 , \42244 , \42246 );
buf \U$42269 ( \42248 , \1229 );
buf \U$42270 ( \42249 , \4433 );
nand \U$42271 ( \42250 , \42248 , \42249 );
buf \U$42272 ( \42251 , \42250 );
buf \U$42273 ( \42252 , \42251 );
nand \U$42274 ( \42253 , \42247 , \42252 );
buf \U$42275 ( \42254 , \42253 );
buf \U$42276 ( \42255 , \42254 );
buf \U$42277 ( \42256 , \40232 );
not \U$42278 ( \42257 , \42256 );
buf \U$42279 ( \42258 , \1823 );
not \U$42280 ( \42259 , \42258 );
or \U$42281 ( \42260 , \42257 , \42259 );
buf \U$42282 ( \42261 , \686 );
buf \U$42283 ( \42262 , \4387 );
nand \U$42284 ( \42263 , \42261 , \42262 );
buf \U$42285 ( \42264 , \42263 );
buf \U$42286 ( \42265 , \42264 );
nand \U$42287 ( \42266 , \42260 , \42265 );
buf \U$42288 ( \42267 , \42266 );
buf \U$42289 ( \42268 , \42267 );
xor \U$42290 ( \42269 , \42255 , \42268 );
buf \U$42291 ( \42270 , \521 );
buf \U$42292 ( \42271 , \40260 );
or \U$42293 ( \42272 , \42270 , \42271 );
buf \U$42294 ( \42273 , \710 );
buf \U$42295 ( \42274 , \4406 );
or \U$42296 ( \42275 , \42273 , \42274 );
nand \U$42297 ( \42276 , \42272 , \42275 );
buf \U$42298 ( \42277 , \42276 );
buf \U$42299 ( \42278 , \42277 );
xor \U$42300 ( \42279 , \42269 , \42278 );
buf \U$42301 ( \42280 , \42279 );
buf \U$42302 ( \42281 , \42280 );
xor \U$42303 ( \42282 , \42242 , \42281 );
buf \U$42304 ( \42283 , \40417 );
not \U$42305 ( \42284 , \42283 );
buf \U$42306 ( \42285 , \26572 );
not \U$42307 ( \42286 , \42285 );
or \U$42308 ( \42287 , \42284 , \42286 );
buf \U$42309 ( \42288 , \734 );
buf \U$42310 ( \42289 , \4326 );
nand \U$42311 ( \42290 , \42288 , \42289 );
buf \U$42312 ( \42291 , \42290 );
buf \U$42313 ( \42292 , \42291 );
nand \U$42314 ( \42293 , \42287 , \42292 );
buf \U$42315 ( \42294 , \42293 );
buf \U$42316 ( \42295 , \40538 );
not \U$42317 ( \42296 , \42295 );
buf \U$42318 ( \42297 , \29546 );
not \U$42319 ( \42298 , \42297 );
or \U$42320 ( \42299 , \42296 , \42298 );
buf \U$42321 ( \42300 , \16584 );
buf \U$42322 ( \42301 , RIc0da648_103);
nand \U$42323 ( \42302 , \42300 , \42301 );
buf \U$42324 ( \42303 , \42302 );
buf \U$42325 ( \42304 , \42303 );
nand \U$42326 ( \42305 , \42299 , \42304 );
buf \U$42327 ( \42306 , \42305 );
xor \U$42328 ( \42307 , \42294 , \42306 );
buf \U$42329 ( \42308 , \3816 );
buf \U$42330 ( \42309 , \40180 );
not \U$42331 ( \42310 , \42309 );
buf \U$42332 ( \42311 , \42310 );
buf \U$42333 ( \42312 , \42311 );
or \U$42334 ( \42313 , \42308 , \42312 );
buf \U$42335 ( \42314 , RIc0d8320_28);
buf \U$42336 ( \42315 , RIc0d9928_75);
xor \U$42337 ( \42316 , \42314 , \42315 );
buf \U$42338 ( \42317 , \42316 );
buf \U$42339 ( \42318 , \42317 );
not \U$42340 ( \42319 , \42318 );
buf \U$42341 ( \42320 , \42319 );
buf \U$42342 ( \42321 , \42320 );
buf \U$42343 ( \42322 , \1562 );
or \U$42344 ( \42323 , \42321 , \42322 );
nand \U$42345 ( \42324 , \42313 , \42323 );
buf \U$42346 ( \42325 , \42324 );
xnor \U$42347 ( \42326 , \42307 , \42325 );
buf \U$42348 ( \42327 , \42326 );
not \U$42349 ( \42328 , \42327 );
buf \U$42350 ( \42329 , \42328 );
buf \U$42351 ( \42330 , \42329 );
xor \U$42352 ( \42331 , \42282 , \42330 );
buf \U$42353 ( \42332 , \42331 );
buf \U$42354 ( \42333 , \42332 );
buf \U$42355 ( \42334 , \40490 );
not \U$42356 ( \42335 , \42334 );
buf \U$42357 ( \42336 , \25371 );
not \U$42358 ( \42337 , \42336 );
or \U$42359 ( \42338 , \42335 , \42337 );
buf \U$42360 ( \42339 , RIc0d77e0_4);
buf \U$42361 ( \42340 , RIc0da468_99);
xnor \U$42362 ( \42341 , \42339 , \42340 );
buf \U$42363 ( \42342 , \42341 );
buf \U$42364 ( \42343 , \42342 );
not \U$42365 ( \42344 , \42343 );
buf \U$42366 ( \42345 , \14648 );
nand \U$42367 ( \42346 , \42344 , \42345 );
buf \U$42368 ( \42347 , \42346 );
buf \U$42369 ( \42348 , \42347 );
nand \U$42370 ( \42349 , \42338 , \42348 );
buf \U$42371 ( \42350 , \42349 );
buf \U$42372 ( \42351 , \42350 );
buf \U$42373 ( \42352 , \40344 );
not \U$42374 ( \42353 , \42352 );
buf \U$42375 ( \42354 , \3415 );
not \U$42376 ( \42355 , \42354 );
or \U$42377 ( \42356 , \42353 , \42355 );
buf \U$42378 ( \42357 , \481 );
buf \U$42379 ( \42358 , \4550 );
nand \U$42380 ( \42359 , \42357 , \42358 );
buf \U$42381 ( \42360 , \42359 );
buf \U$42382 ( \42361 , \42360 );
nand \U$42383 ( \42362 , \42356 , \42361 );
buf \U$42384 ( \42363 , \42362 );
buf \U$42385 ( \42364 , \42363 );
xor \U$42386 ( \42365 , \42351 , \42364 );
buf \U$42387 ( \42366 , \5362 );
buf \U$42388 ( \42367 , \40438 );
or \U$42389 ( \42368 , \42366 , \42367 );
buf \U$42390 ( \42369 , \5368 );
and \U$42391 ( \42370 , RIc0d9fb8_89, \40247 );
not \U$42392 ( \42371 , RIc0d9fb8_89);
and \U$42393 ( \42372 , \42371 , RIc0d7c90_14);
nor \U$42394 ( \42373 , \42370 , \42372 );
buf \U$42395 ( \42374 , \42373 );
or \U$42396 ( \42375 , \42369 , \42374 );
nand \U$42397 ( \42376 , \42368 , \42375 );
buf \U$42398 ( \42377 , \42376 );
buf \U$42399 ( \42378 , \42377 );
xor \U$42400 ( \42379 , \42365 , \42378 );
buf \U$42401 ( \42380 , \42379 );
buf \U$42402 ( \42381 , \42380 );
buf \U$42403 ( \42382 , \40372 );
not \U$42404 ( \42383 , \42382 );
buf \U$42405 ( \42384 , \2812 );
not \U$42406 ( \42385 , \42384 );
or \U$42407 ( \42386 , \42383 , \42385 );
buf \U$42408 ( \42387 , \1282 );
buf \U$42409 ( \42388 , \4311 );
nand \U$42410 ( \42389 , \42387 , \42388 );
buf \U$42411 ( \42390 , \42389 );
buf \U$42412 ( \42391 , \42390 );
nand \U$42413 ( \42392 , \42386 , \42391 );
buf \U$42414 ( \42393 , \42392 );
buf \U$42415 ( \42394 , \42393 );
buf \U$42416 ( \42395 , \40296 );
not \U$42417 ( \42396 , \42395 );
buf \U$42418 ( \42397 , \2871 );
not \U$42419 ( \42398 , \42397 );
or \U$42420 ( \42399 , \42396 , \42398 );
buf \U$42421 ( \42400 , RIc0d8410_30);
buf \U$42422 ( \42401 , RIc0d9838_73);
xnor \U$42423 ( \42402 , \42400 , \42401 );
buf \U$42424 ( \42403 , \42402 );
buf \U$42425 ( \42404 , \42403 );
not \U$42426 ( \42405 , \42404 );
buf \U$42427 ( \42406 , \791 );
nand \U$42428 ( \42407 , \42405 , \42406 );
buf \U$42429 ( \42408 , \42407 );
buf \U$42430 ( \42409 , \42408 );
nand \U$42431 ( \42410 , \42399 , \42409 );
buf \U$42432 ( \42411 , \42410 );
buf \U$42433 ( \42412 , \42411 );
xor \U$42434 ( \42413 , \42394 , \42412 );
buf \U$42435 ( \42414 , \989 );
buf \U$42436 ( \42415 , \40759 );
or \U$42437 ( \42416 , \42414 , \42415 );
buf \U$42438 ( \42417 , \996 );
buf \U$42439 ( \42418 , \4349 );
or \U$42440 ( \42419 , \42417 , \42418 );
nand \U$42441 ( \42420 , \42416 , \42419 );
buf \U$42442 ( \42421 , \42420 );
buf \U$42443 ( \42422 , \42421 );
xor \U$42444 ( \42423 , \42413 , \42422 );
buf \U$42445 ( \42424 , \42423 );
buf \U$42446 ( \42425 , \42424 );
xor \U$42447 ( \42426 , \42381 , \42425 );
buf \U$42448 ( \42427 , \40735 );
not \U$42449 ( \42428 , \42427 );
buf \U$42450 ( \42429 , \4692 );
not \U$42451 ( \42430 , \42429 );
or \U$42452 ( \42431 , \42428 , \42430 );
buf \U$42453 ( \42432 , \284 );
buf \U$42454 ( \42433 , RIc0d85f0_34);
buf \U$42455 ( \42434 , RIc0d9658_69);
xor \U$42456 ( \42435 , \42433 , \42434 );
buf \U$42457 ( \42436 , \42435 );
buf \U$42458 ( \42437 , \42436 );
nand \U$42459 ( \42438 , \42432 , \42437 );
buf \U$42460 ( \42439 , \42438 );
buf \U$42461 ( \42440 , \42439 );
nand \U$42462 ( \42441 , \42431 , \42440 );
buf \U$42463 ( \42442 , \42441 );
buf \U$42464 ( \42443 , \42442 );
buf \U$42465 ( \42444 , \40514 );
not \U$42466 ( \42445 , \42444 );
buf \U$42467 ( \42446 , \42445 );
buf \U$42468 ( \42447 , \42446 );
not \U$42469 ( \42448 , \42447 );
buf \U$42470 ( \42449 , \1063 );
not \U$42471 ( \42450 , \42449 );
or \U$42472 ( \42451 , \42448 , \42450 );
buf \U$42473 ( \42452 , RIc0d9bf8_81);
buf \U$42474 ( \42453 , RIc0d8050_22);
xnor \U$42475 ( \42454 , \42452 , \42453 );
buf \U$42476 ( \42455 , \42454 );
buf \U$42477 ( \42456 , \42455 );
not \U$42478 ( \42457 , \42456 );
buf \U$42479 ( \42458 , \1078 );
nand \U$42480 ( \42459 , \42457 , \42458 );
buf \U$42481 ( \42460 , \42459 );
buf \U$42482 ( \42461 , \42460 );
nand \U$42483 ( \42462 , \42451 , \42461 );
buf \U$42484 ( \42463 , \42462 );
buf \U$42485 ( \42464 , \42463 );
xor \U$42486 ( \42465 , \42443 , \42464 );
buf \U$42487 ( \42466 , \7753 );
buf \U$42488 ( \42467 , \40161 );
or \U$42489 ( \42468 , \42466 , \42467 );
buf \U$42490 ( \42469 , \1193 );
buf \U$42491 ( \42470 , RIc0d8230_26);
buf \U$42492 ( \42471 , RIc0d9a18_77);
xor \U$42493 ( \42472 , \42470 , \42471 );
buf \U$42494 ( \42473 , \42472 );
buf \U$42495 ( \42474 , \42473 );
not \U$42496 ( \42475 , \42474 );
buf \U$42497 ( \42476 , \42475 );
buf \U$42498 ( \42477 , \42476 );
or \U$42499 ( \42478 , \42469 , \42477 );
nand \U$42500 ( \42479 , \42468 , \42478 );
buf \U$42501 ( \42480 , \42479 );
buf \U$42502 ( \42481 , \42480 );
xor \U$42503 ( \42482 , \42465 , \42481 );
buf \U$42504 ( \42483 , \42482 );
buf \U$42505 ( \42484 , \42483 );
xor \U$42506 ( \42485 , \42426 , \42484 );
buf \U$42507 ( \42486 , \42485 );
buf \U$42508 ( \42487 , \42486 );
xor \U$42509 ( \42488 , \42333 , \42487 );
xor \U$42510 ( \42489 , \40767 , \40832 );
and \U$42511 ( \42490 , \42489 , \40881 );
and \U$42512 ( \42491 , \40767 , \40832 );
or \U$42513 ( \42492 , \42490 , \42491 );
buf \U$42514 ( \42493 , \42492 );
buf \U$42515 ( \42494 , \42493 );
xor \U$42516 ( \42495 , \42488 , \42494 );
buf \U$42517 ( \42496 , \42495 );
buf \U$42518 ( \42497 , \42496 );
xor \U$42519 ( \42498 , \42225 , \42497 );
buf \U$42520 ( \42499 , \42498 );
buf \U$42521 ( \42500 , \42499 );
xor \U$42522 ( \42501 , \42139 , \42500 );
xor \U$42523 ( \42502 , \40632 , \40698 );
and \U$42524 ( \42503 , \42502 , \41251 );
and \U$42525 ( \42504 , \40632 , \40698 );
or \U$42526 ( \42505 , \42503 , \42504 );
buf \U$42527 ( \42506 , \42505 );
buf \U$42528 ( \42507 , \42506 );
xor \U$42529 ( \42508 , \42501 , \42507 );
buf \U$42530 ( \42509 , \42508 );
buf \U$42531 ( \42510 , \42509 );
xor \U$42532 ( \42511 , \42133 , \42510 );
xor \U$42533 ( \42512 , \41407 , \41433 );
and \U$42534 ( \42513 , \42512 , \41485 );
and \U$42535 ( \42514 , \41407 , \41433 );
or \U$42536 ( \42515 , \42513 , \42514 );
buf \U$42537 ( \42516 , \42515 );
buf \U$42538 ( \42517 , \42516 );
xor \U$42539 ( \42518 , \42511 , \42517 );
buf \U$42540 ( \42519 , \42518 );
buf \U$42541 ( \42520 , \42519 );
not \U$42542 ( \42521 , \42520 );
buf \U$42543 ( \42522 , \42521 );
buf \U$42544 ( \42523 , \42522 );
nand \U$42545 ( \42524 , \41979 , \42523 );
buf \U$42546 ( \42525 , \42524 );
buf \U$42547 ( \42526 , \42525 );
xor \U$42548 ( \42527 , \42133 , \42510 );
and \U$42549 ( \42528 , \42527 , \42517 );
and \U$42550 ( \42529 , \42133 , \42510 );
or \U$42551 ( \42530 , \42528 , \42529 );
buf \U$42552 ( \42531 , \42530 );
not \U$42553 ( \42532 , \42531 );
xor \U$42554 ( \42533 , \41985 , \42123 );
and \U$42555 ( \42534 , \42533 , \42130 );
and \U$42556 ( \42535 , \41985 , \42123 );
or \U$42557 ( \42536 , \42534 , \42535 );
buf \U$42558 ( \42537 , \42536 );
buf \U$42559 ( \42538 , \42537 );
not \U$42560 ( \42539 , \42538 );
buf \U$42561 ( \42540 , \42539 );
buf \U$42562 ( \42541 , \42540 );
xor \U$42563 ( \42542 , \42139 , \42500 );
and \U$42564 ( \42543 , \42542 , \42507 );
and \U$42565 ( \42544 , \42139 , \42500 );
or \U$42566 ( \42545 , \42543 , \42544 );
buf \U$42567 ( \42546 , \42545 );
buf \U$42568 ( \42547 , \42546 );
not \U$42569 ( \42548 , \42547 );
buf \U$42570 ( \42549 , \42548 );
buf \U$42571 ( \42550 , \42549 );
xor \U$42572 ( \42551 , \42541 , \42550 );
xor \U$42573 ( \42552 , \42145 , \42224 );
and \U$42574 ( \42553 , \42552 , \42497 );
and \U$42575 ( \42554 , \42145 , \42224 );
or \U$42576 ( \42555 , \42553 , \42554 );
buf \U$42577 ( \42556 , \42555 );
xor \U$42578 ( \42557 , \42104 , \42110 );
and \U$42579 ( \42558 , \42557 , \42117 );
and \U$42580 ( \42559 , \42104 , \42110 );
or \U$42581 ( \42560 , \42558 , \42559 );
buf \U$42582 ( \42561 , \42560 );
buf \U$42583 ( \42562 , \42561 );
buf \U$42584 ( \42563 , \42241 );
not \U$42585 ( \42564 , \42563 );
buf \U$42586 ( \42565 , \42329 );
not \U$42587 ( \42566 , \42565 );
or \U$42588 ( \42567 , \42564 , \42566 );
buf \U$42589 ( \42568 , \42241 );
not \U$42590 ( \42569 , \42568 );
buf \U$42591 ( \42570 , \42326 );
nand \U$42592 ( \42571 , \42569 , \42570 );
buf \U$42593 ( \42572 , \42571 );
buf \U$42594 ( \42573 , \42572 );
buf \U$42595 ( \42574 , \42280 );
nand \U$42596 ( \42575 , \42573 , \42574 );
buf \U$42597 ( \42576 , \42575 );
buf \U$42598 ( \42577 , \42576 );
nand \U$42599 ( \42578 , \42567 , \42577 );
buf \U$42600 ( \42579 , \42578 );
buf \U$42601 ( \42580 , \42579 );
buf \U$42602 ( \42581 , \42000 );
not \U$42603 ( \42582 , \42581 );
buf \U$42604 ( \42583 , \42582 );
buf \U$42605 ( \42584 , \42583 );
xor \U$42606 ( \42585 , \42394 , \42412 );
and \U$42607 ( \42586 , \42585 , \42422 );
and \U$42608 ( \42587 , \42394 , \42412 );
or \U$42609 ( \42588 , \42586 , \42587 );
buf \U$42610 ( \42589 , \42588 );
buf \U$42611 ( \42590 , \42589 );
xor \U$42612 ( \42591 , \42584 , \42590 );
buf \U$42613 ( \42592 , \42325 );
buf \U$42614 ( \42593 , \42294 );
or \U$42615 ( \42594 , \42592 , \42593 );
buf \U$42616 ( \42595 , \42306 );
nand \U$42617 ( \42596 , \42594 , \42595 );
buf \U$42618 ( \42597 , \42596 );
buf \U$42619 ( \42598 , \42597 );
buf \U$42620 ( \42599 , \42325 );
buf \U$42621 ( \42600 , \42294 );
nand \U$42622 ( \42601 , \42599 , \42600 );
buf \U$42623 ( \42602 , \42601 );
buf \U$42624 ( \42603 , \42602 );
nand \U$42625 ( \42604 , \42598 , \42603 );
buf \U$42626 ( \42605 , \42604 );
buf \U$42627 ( \42606 , \42605 );
xor \U$42628 ( \42607 , \42591 , \42606 );
buf \U$42629 ( \42608 , \42607 );
buf \U$42630 ( \42609 , \42608 );
xor \U$42631 ( \42610 , \42580 , \42609 );
xor \U$42632 ( \42611 , \42381 , \42425 );
and \U$42633 ( \42612 , \42611 , \42484 );
and \U$42634 ( \42613 , \42381 , \42425 );
or \U$42635 ( \42614 , \42612 , \42613 );
buf \U$42636 ( \42615 , \42614 );
buf \U$42637 ( \42616 , \42615 );
xor \U$42638 ( \42617 , \42610 , \42616 );
buf \U$42639 ( \42618 , \42617 );
buf \U$42640 ( \42619 , \42618 );
xor \U$42641 ( \42620 , \42562 , \42619 );
xor \U$42642 ( \42621 , \42443 , \42464 );
and \U$42643 ( \42622 , \42621 , \42481 );
and \U$42644 ( \42623 , \42443 , \42464 );
or \U$42645 ( \42624 , \42622 , \42623 );
buf \U$42646 ( \42625 , \42624 );
buf \U$42647 ( \42626 , \42625 );
xor \U$42648 ( \42627 , \4383 , \4400 );
xor \U$42649 ( \42628 , \42627 , \4417 );
buf \U$42650 ( \42629 , \42628 );
buf \U$42651 ( \42630 , \42629 );
xor \U$42652 ( \42631 , \42626 , \42630 );
xor \U$42653 ( \42632 , \4537 , \4562 );
buf \U$42654 ( \42633 , \42632 );
buf \U$42655 ( \42634 , \4519 );
xor \U$42656 ( \42635 , \42633 , \42634 );
buf \U$42657 ( \42636 , \42635 );
buf \U$42658 ( \42637 , \42636 );
xor \U$42659 ( \42638 , \42631 , \42637 );
buf \U$42660 ( \42639 , \42638 );
buf \U$42661 ( \42640 , \42639 );
xor \U$42662 ( \42641 , \41988 , \42001 );
and \U$42663 ( \42642 , \42641 , \42022 );
and \U$42664 ( \42643 , \41988 , \42001 );
or \U$42665 ( \42644 , \42642 , \42643 );
buf \U$42666 ( \42645 , \42644 );
buf \U$42667 ( \42646 , \42645 );
buf \U$42668 ( \42647 , \3566 );
buf \U$42669 ( \42648 , \42455 );
or \U$42670 ( \42649 , \42647 , \42648 );
buf \U$42671 ( \42650 , \1610 );
buf \U$42672 ( \42651 , \3692 );
not \U$42673 ( \42652 , \42651 );
buf \U$42674 ( \42653 , \42652 );
buf \U$42675 ( \42654 , \42653 );
or \U$42676 ( \42655 , \42650 , \42654 );
nand \U$42677 ( \42656 , \42649 , \42655 );
buf \U$42678 ( \42657 , \42656 );
buf \U$42679 ( \42658 , \42657 );
not \U$42680 ( \42659 , \42658 );
buf \U$42681 ( \42660 , \42473 );
not \U$42682 ( \42661 , \42660 );
buf \U$42683 ( \42662 , \1432 );
not \U$42684 ( \42663 , \42662 );
or \U$42685 ( \42664 , \42661 , \42663 );
buf \U$42686 ( \42665 , \6141 );
buf \U$42687 ( \42666 , \3734 );
nand \U$42688 ( \42667 , \42665 , \42666 );
buf \U$42689 ( \42668 , \42667 );
buf \U$42690 ( \42669 , \42668 );
nand \U$42691 ( \42670 , \42664 , \42669 );
buf \U$42692 ( \42671 , \42670 );
buf \U$42693 ( \42672 , \42671 );
not \U$42694 ( \42673 , \42672 );
buf \U$42695 ( \42674 , \42673 );
buf \U$42696 ( \42675 , \42674 );
not \U$42697 ( \42676 , \42675 );
buf \U$42698 ( \42677 , \42048 );
not \U$42699 ( \42678 , \42677 );
buf \U$42700 ( \42679 , \22631 );
not \U$42701 ( \42680 , \42679 );
or \U$42702 ( \42681 , \42678 , \42680 );
buf \U$42703 ( \42682 , \4049 );
buf \U$42704 ( \42683 , \4039 );
nand \U$42705 ( \42684 , \42682 , \42683 );
buf \U$42706 ( \42685 , \42684 );
buf \U$42707 ( \42686 , \42685 );
nand \U$42708 ( \42687 , \42681 , \42686 );
buf \U$42709 ( \42688 , \42687 );
buf \U$42710 ( \42689 , \42688 );
not \U$42711 ( \42690 , \42689 );
and \U$42712 ( \42691 , \42676 , \42690 );
buf \U$42713 ( \42692 , \42674 );
buf \U$42714 ( \42693 , \42688 );
and \U$42715 ( \42694 , \42692 , \42693 );
nor \U$42716 ( \42695 , \42691 , \42694 );
buf \U$42717 ( \42696 , \42695 );
buf \U$42718 ( \42697 , \42696 );
not \U$42719 ( \42698 , \42697 );
or \U$42720 ( \42699 , \42659 , \42698 );
buf \U$42721 ( \42700 , \42696 );
buf \U$42722 ( \42701 , \42657 );
or \U$42723 ( \42702 , \42700 , \42701 );
nand \U$42724 ( \42703 , \42699 , \42702 );
buf \U$42725 ( \42704 , \42703 );
buf \U$42726 ( \42705 , \42704 );
xor \U$42727 ( \42706 , \42646 , \42705 );
xor \U$42728 ( \42707 , \4489 , \4464 );
xor \U$42729 ( \42708 , \42707 , \4439 );
buf \U$42730 ( \42709 , \42708 );
xor \U$42731 ( \42710 , \42706 , \42709 );
buf \U$42732 ( \42711 , \42710 );
buf \U$42733 ( \42712 , \42711 );
xor \U$42734 ( \42713 , \42640 , \42712 );
buf \U$42735 ( \42714 , \42317 );
not \U$42736 ( \42715 , \42714 );
buf \U$42737 ( \42716 , \2124 );
not \U$42738 ( \42717 , \42716 );
or \U$42739 ( \42718 , \42715 , \42717 );
buf \U$42740 ( \42719 , \3821 );
not \U$42741 ( \42720 , \42719 );
buf \U$42742 ( \42721 , \1143 );
nand \U$42743 ( \42722 , \42720 , \42721 );
buf \U$42744 ( \42723 , \42722 );
buf \U$42745 ( \42724 , \42723 );
nand \U$42746 ( \42725 , \42718 , \42724 );
buf \U$42747 ( \42726 , \42725 );
buf \U$42748 ( \42727 , \42726 );
buf \U$42749 ( \42728 , \3957 );
not \U$42750 ( \42729 , \42728 );
buf \U$42751 ( \42730 , \846 );
not \U$42752 ( \42731 , \42730 );
or \U$42753 ( \42732 , \42729 , \42731 );
buf \U$42754 ( \42733 , \42373 );
not \U$42755 ( \42734 , \42733 );
buf \U$42756 ( \42735 , \2038 );
nand \U$42757 ( \42736 , \42734 , \42735 );
buf \U$42758 ( \42737 , \42736 );
buf \U$42759 ( \42738 , \42737 );
nand \U$42760 ( \42739 , \42732 , \42738 );
buf \U$42761 ( \42740 , \42739 );
buf \U$42762 ( \42741 , \42740 );
xor \U$42763 ( \42742 , \42727 , \42741 );
buf \U$42764 ( \42743 , \25374 );
buf \U$42765 ( \42744 , \42342 );
or \U$42766 ( \42745 , \42743 , \42744 );
buf \U$42767 ( \42746 , \2198 );
buf \U$42768 ( \42747 , \3837 );
or \U$42769 ( \42748 , \42746 , \42747 );
nand \U$42770 ( \42749 , \42745 , \42748 );
buf \U$42771 ( \42750 , \42749 );
buf \U$42772 ( \42751 , \42750 );
xor \U$42773 ( \42752 , \42742 , \42751 );
buf \U$42774 ( \42753 , \42752 );
xor \U$42775 ( \42754 , \4365 , \4339 );
xor \U$42776 ( \42755 , \42754 , \4323 );
xor \U$42777 ( \42756 , \42753 , \42755 );
buf \U$42778 ( \42757 , \42014 );
not \U$42779 ( \42758 , \42757 );
buf \U$42780 ( \42759 , \2399 );
not \U$42781 ( \42760 , \42759 );
or \U$42782 ( \42761 , \42758 , \42760 );
buf \U$42783 ( \42762 , \1401 );
buf \U$42784 ( \42763 , \4083 );
nand \U$42785 ( \42764 , \42762 , \42763 );
buf \U$42786 ( \42765 , \42764 );
buf \U$42787 ( \42766 , \42765 );
nand \U$42788 ( \42767 , \42761 , \42766 );
buf \U$42789 ( \42768 , \42767 );
buf \U$42790 ( \42769 , \42768 );
buf \U$42791 ( \42770 , \42436 );
not \U$42792 ( \42771 , \42770 );
buf \U$42793 ( \42772 , \279 );
not \U$42794 ( \42773 , \42772 );
or \U$42795 ( \42774 , \42771 , \42773 );
buf \U$42796 ( \42775 , \4292 );
not \U$42797 ( \42776 , \42775 );
buf \U$42798 ( \42777 , \874 );
nand \U$42799 ( \42778 , \42776 , \42777 );
buf \U$42800 ( \42779 , \42778 );
buf \U$42801 ( \42780 , \42779 );
nand \U$42802 ( \42781 , \42774 , \42780 );
buf \U$42803 ( \42782 , \42781 );
buf \U$42804 ( \42783 , \42782 );
xor \U$42805 ( \42784 , \42769 , \42783 );
buf \U$42806 ( \42785 , \779 );
buf \U$42807 ( \42786 , \42403 );
or \U$42808 ( \42787 , \42785 , \42786 );
buf \U$42809 ( \42788 , \9493 );
buf \U$42810 ( \42789 , \4123 );
or \U$42811 ( \42790 , \42788 , \42789 );
nand \U$42812 ( \42791 , \42787 , \42790 );
buf \U$42813 ( \42792 , \42791 );
buf \U$42814 ( \42793 , \42792 );
xor \U$42815 ( \42794 , \42784 , \42793 );
buf \U$42816 ( \42795 , \42794 );
xor \U$42817 ( \42796 , \42756 , \42795 );
buf \U$42818 ( \42797 , \42796 );
xor \U$42819 ( \42798 , \42713 , \42797 );
buf \U$42820 ( \42799 , \42798 );
buf \U$42821 ( \42800 , \42799 );
xor \U$42822 ( \42801 , \42620 , \42800 );
buf \U$42823 ( \42802 , \42801 );
xnor \U$42824 ( \42803 , \42556 , \42802 );
buf \U$42825 ( \42804 , \42803 );
not \U$42826 ( \42805 , \42804 );
xor \U$42827 ( \42806 , \42333 , \42487 );
and \U$42828 ( \42807 , \42806 , \42494 );
and \U$42829 ( \42808 , \42333 , \42487 );
or \U$42830 ( \42809 , \42807 , \42808 );
buf \U$42831 ( \42810 , \42809 );
buf \U$42832 ( \42811 , \42810 );
xor \U$42833 ( \42812 , \42082 , \42088 );
and \U$42834 ( \42813 , \42812 , \42120 );
and \U$42835 ( \42814 , \42082 , \42088 );
or \U$42836 ( \42815 , \42813 , \42814 );
buf \U$42837 ( \42816 , \42815 );
buf \U$42838 ( \42817 , \42816 );
xor \U$42839 ( \42818 , \42811 , \42817 );
xor \U$42840 ( \42819 , \42025 , \42072 );
and \U$42841 ( \42820 , \42819 , \42079 );
and \U$42842 ( \42821 , \42025 , \42072 );
or \U$42843 ( \42822 , \42820 , \42821 );
buf \U$42844 ( \42823 , \42822 );
buf \U$42845 ( \42824 , \42823 );
xor \U$42846 ( \42825 , \42158 , \42198 );
and \U$42847 ( \42826 , \42825 , \42221 );
and \U$42848 ( \42827 , \42158 , \42198 );
or \U$42849 ( \42828 , \42826 , \42827 );
buf \U$42850 ( \42829 , \42828 );
buf \U$42851 ( \42830 , \42829 );
xor \U$42852 ( \42831 , \42824 , \42830 );
xor \U$42853 ( \42832 , \42173 , \42188 );
and \U$42854 ( \42833 , \42832 , \42195 );
and \U$42855 ( \42834 , \42173 , \42188 );
or \U$42856 ( \42835 , \42833 , \42834 );
buf \U$42857 ( \42836 , \42835 );
buf \U$42858 ( \42837 , \42836 );
xor \U$42859 ( \42838 , \42205 , \42211 );
and \U$42860 ( \42839 , \42838 , \42218 );
and \U$42861 ( \42840 , \42205 , \42211 );
or \U$42862 ( \42841 , \42839 , \42840 );
buf \U$42863 ( \42842 , \42841 );
buf \U$42864 ( \42843 , \42842 );
xor \U$42865 ( \42844 , \42837 , \42843 );
xor \U$42866 ( \42845 , \42255 , \42268 );
and \U$42867 ( \42846 , \42845 , \42278 );
and \U$42868 ( \42847 , \42255 , \42268 );
or \U$42869 ( \42848 , \42846 , \42847 );
buf \U$42870 ( \42849 , \42848 );
buf \U$42871 ( \42850 , \42849 );
xor \U$42872 ( \42851 , \42351 , \42364 );
and \U$42873 ( \42852 , \42851 , \42378 );
and \U$42874 ( \42853 , \42351 , \42364 );
or \U$42875 ( \42854 , \42852 , \42853 );
buf \U$42876 ( \42855 , \42854 );
buf \U$42877 ( \42856 , \42855 );
xor \U$42878 ( \42857 , \42850 , \42856 );
xor \U$42879 ( \42858 , \42037 , \42056 );
and \U$42880 ( \42859 , \42858 , \42069 );
and \U$42881 ( \42860 , \42037 , \42056 );
or \U$42882 ( \42861 , \42859 , \42860 );
buf \U$42883 ( \42862 , \42861 );
buf \U$42884 ( \42863 , \42862 );
xor \U$42885 ( \42864 , \42857 , \42863 );
buf \U$42886 ( \42865 , \42864 );
buf \U$42887 ( \42866 , \42865 );
xor \U$42888 ( \42867 , \42844 , \42866 );
buf \U$42889 ( \42868 , \42867 );
buf \U$42890 ( \42869 , \42868 );
xor \U$42891 ( \42870 , \42831 , \42869 );
buf \U$42892 ( \42871 , \42870 );
buf \U$42893 ( \42872 , \42871 );
xor \U$42894 ( \42873 , \42818 , \42872 );
buf \U$42895 ( \42874 , \42873 );
buf \U$42896 ( \42875 , \42874 );
not \U$42897 ( \42876 , \42875 );
and \U$42898 ( \42877 , \42805 , \42876 );
buf \U$42899 ( \42878 , \42803 );
buf \U$42900 ( \42879 , \42874 );
and \U$42901 ( \42880 , \42878 , \42879 );
nor \U$42902 ( \42881 , \42877 , \42880 );
buf \U$42903 ( \42882 , \42881 );
buf \U$42904 ( \42883 , \42882 );
xor \U$42905 ( \42884 , \42551 , \42883 );
buf \U$42906 ( \42885 , \42884 );
nand \U$42907 ( \42886 , \42532 , \42885 );
buf \U$42908 ( \42887 , \42886 );
nand \U$42909 ( \42888 , \42526 , \42887 );
buf \U$42910 ( \42889 , \42888 );
buf \U$42911 ( \42890 , \42889 );
not \U$42912 ( \42891 , \42890 );
buf \U$42913 ( \42892 , \42891 );
buf \U$42914 ( \42893 , \42892 );
xor \U$42915 ( \42894 , \42811 , \42817 );
and \U$42916 ( \42895 , \42894 , \42872 );
and \U$42917 ( \42896 , \42811 , \42817 );
or \U$42918 ( \42897 , \42895 , \42896 );
buf \U$42919 ( \42898 , \42897 );
buf \U$42920 ( \42899 , \42898 );
not \U$42921 ( \42900 , \42899 );
buf \U$42922 ( \42901 , \42900 );
buf \U$42923 ( \42902 , \42901 );
not \U$42924 ( \42903 , \42902 );
xor \U$42925 ( \42904 , \42562 , \42619 );
and \U$42926 ( \42905 , \42904 , \42800 );
and \U$42927 ( \42906 , \42562 , \42619 );
or \U$42928 ( \42907 , \42905 , \42906 );
buf \U$42929 ( \42908 , \42907 );
xor \U$42930 ( \42909 , \42580 , \42609 );
and \U$42931 ( \42910 , \42909 , \42616 );
and \U$42932 ( \42911 , \42580 , \42609 );
or \U$42933 ( \42912 , \42910 , \42911 );
buf \U$42934 ( \42913 , \42912 );
xor \U$42935 ( \42914 , \4422 , \4496 );
xor \U$42936 ( \42915 , \42914 , \4574 );
buf \U$42937 ( \42916 , \42915 );
buf \U$42938 ( \42917 , \42916 );
buf \U$42939 ( \42918 , \42671 );
not \U$42940 ( \42919 , \42918 );
buf \U$42941 ( \42920 , \42657 );
not \U$42942 ( \42921 , \42920 );
or \U$42943 ( \42922 , \42919 , \42921 );
buf \U$42944 ( \42923 , \42657 );
buf \U$42945 ( \42924 , \42671 );
or \U$42946 ( \42925 , \42923 , \42924 );
buf \U$42947 ( \42926 , \42688 );
nand \U$42948 ( \42927 , \42925 , \42926 );
buf \U$42949 ( \42928 , \42927 );
buf \U$42950 ( \42929 , \42928 );
nand \U$42951 ( \42930 , \42922 , \42929 );
buf \U$42952 ( \42931 , \42930 );
buf \U$42953 ( \42932 , \42931 );
xor \U$42954 ( \42933 , \42769 , \42783 );
and \U$42955 ( \42934 , \42933 , \42793 );
and \U$42956 ( \42935 , \42769 , \42783 );
or \U$42957 ( \42936 , \42934 , \42935 );
buf \U$42958 ( \42937 , \42936 );
buf \U$42959 ( \42938 , \42937 );
xor \U$42960 ( \42939 , \42932 , \42938 );
xor \U$42961 ( \42940 , \42727 , \42741 );
and \U$42962 ( \42941 , \42940 , \42751 );
and \U$42963 ( \42942 , \42727 , \42741 );
or \U$42964 ( \42943 , \42941 , \42942 );
buf \U$42965 ( \42944 , \42943 );
buf \U$42966 ( \42945 , \42944 );
xor \U$42967 ( \42946 , \42939 , \42945 );
buf \U$42968 ( \42947 , \42946 );
buf \U$42969 ( \42948 , \42947 );
xor \U$42970 ( \42949 , \42917 , \42948 );
buf \U$42971 ( \42950 , \42795 );
not \U$42972 ( \42951 , \42950 );
buf \U$42973 ( \42952 , \42753 );
not \U$42974 ( \42953 , \42952 );
or \U$42975 ( \42954 , \42951 , \42953 );
buf \U$42976 ( \42955 , \42753 );
buf \U$42977 ( \42956 , \42795 );
or \U$42978 ( \42957 , \42955 , \42956 );
buf \U$42979 ( \42958 , \42755 );
nand \U$42980 ( \42959 , \42957 , \42958 );
buf \U$42981 ( \42960 , \42959 );
buf \U$42982 ( \42961 , \42960 );
nand \U$42983 ( \42962 , \42954 , \42961 );
buf \U$42984 ( \42963 , \42962 );
buf \U$42985 ( \42964 , \42963 );
xor \U$42986 ( \42965 , \42949 , \42964 );
buf \U$42987 ( \42966 , \42965 );
xor \U$42988 ( \42967 , \42913 , \42966 );
xor \U$42989 ( \42968 , \42640 , \42712 );
and \U$42990 ( \42969 , \42968 , \42797 );
and \U$42991 ( \42970 , \42640 , \42712 );
or \U$42992 ( \42971 , \42969 , \42970 );
buf \U$42993 ( \42972 , \42971 );
xnor \U$42994 ( \42973 , \42967 , \42972 );
xnor \U$42995 ( \42974 , \42908 , \42973 );
buf \U$42996 ( \42975 , \42974 );
not \U$42997 ( \42976 , \42975 );
xor \U$42998 ( \42977 , \42646 , \42705 );
and \U$42999 ( \42978 , \42977 , \42709 );
and \U$43000 ( \42979 , \42646 , \42705 );
or \U$43001 ( \42980 , \42978 , \42979 );
buf \U$43002 ( \42981 , \42980 );
buf \U$43003 ( \42982 , \42981 );
xor \U$43004 ( \42983 , \42626 , \42630 );
and \U$43005 ( \42984 , \42983 , \42637 );
and \U$43006 ( \42985 , \42626 , \42630 );
or \U$43007 ( \42986 , \42984 , \42985 );
buf \U$43008 ( \42987 , \42986 );
buf \U$43009 ( \42988 , \42987 );
xor \U$43010 ( \42989 , \42982 , \42988 );
xor \U$43011 ( \42990 , \4031 , \4057 );
xor \U$43012 ( \42991 , \42990 , \4074 );
buf \U$43013 ( \42992 , \42991 );
buf \U$43014 ( \42993 , \42992 );
xor \U$43015 ( \42994 , \3705 , \3749 );
xor \U$43016 ( \42995 , \42994 , \3724 );
buf \U$43017 ( \42996 , \42995 );
xor \U$43018 ( \42997 , \42993 , \42996 );
and \U$43019 ( \42998 , \4015 , \3973 );
not \U$43020 ( \42999 , \4015 );
and \U$43021 ( \43000 , \42999 , \3970 );
or \U$43022 ( \43001 , \42998 , \43000 );
buf \U$43023 ( \43002 , \43001 );
buf \U$43024 ( \43003 , \3992 );
and \U$43025 ( \43004 , \43002 , \43003 );
not \U$43026 ( \43005 , \43002 );
buf \U$43027 ( \43006 , \3995 );
and \U$43028 ( \43007 , \43005 , \43006 );
nor \U$43029 ( \43008 , \43004 , \43007 );
buf \U$43030 ( \43009 , \43008 );
buf \U$43031 ( \43010 , \43009 );
xor \U$43032 ( \43011 , \42997 , \43010 );
buf \U$43033 ( \43012 , \43011 );
buf \U$43034 ( \43013 , \43012 );
xor \U$43035 ( \43014 , \42989 , \43013 );
buf \U$43036 ( \43015 , \43014 );
buf \U$43037 ( \43016 , \43015 );
xor \U$43038 ( \43017 , \42824 , \42830 );
and \U$43039 ( \43018 , \43017 , \42869 );
and \U$43040 ( \43019 , \42824 , \42830 );
or \U$43041 ( \43020 , \43018 , \43019 );
buf \U$43042 ( \43021 , \43020 );
buf \U$43043 ( \43022 , \43021 );
xor \U$43044 ( \43023 , \43016 , \43022 );
xor \U$43045 ( \43024 , \3773 , \3791 );
xor \U$43046 ( \43025 , \43024 , \3808 );
buf \U$43047 ( \43026 , \43025 );
buf \U$43048 ( \43027 , \4096 );
buf \U$43049 ( \43028 , \4113 );
and \U$43050 ( \43029 , \43027 , \43028 );
not \U$43051 ( \43030 , \43027 );
buf \U$43052 ( \43031 , \4116 );
and \U$43053 ( \43032 , \43030 , \43031 );
nor \U$43054 ( \43033 , \43029 , \43032 );
buf \U$43055 ( \43034 , \43033 );
buf \U$43056 ( \43035 , \43034 );
buf \U$43057 ( \43036 , \4133 );
xor \U$43058 ( \43037 , \43035 , \43036 );
buf \U$43059 ( \43038 , \43037 );
buf \U$43060 ( \43039 , \43038 );
xor \U$43061 ( \43040 , \43026 , \43039 );
buf \U$43062 ( \43041 , \3828 );
not \U$43063 ( \43042 , \43041 );
buf \U$43064 ( \43043 , \3871 );
buf \U$43065 ( \43044 , \3852 );
xnor \U$43066 ( \43045 , \43043 , \43044 );
buf \U$43067 ( \43046 , \43045 );
buf \U$43068 ( \43047 , \43046 );
not \U$43069 ( \43048 , \43047 );
or \U$43070 ( \43049 , \43042 , \43048 );
buf \U$43071 ( \43050 , \43046 );
buf \U$43072 ( \43051 , \3828 );
or \U$43073 ( \43052 , \43050 , \43051 );
nand \U$43074 ( \43053 , \43049 , \43052 );
buf \U$43075 ( \43054 , \43053 );
buf \U$43076 ( \43055 , \43054 );
xor \U$43077 ( \43056 , \43040 , \43055 );
buf \U$43078 ( \43057 , \43056 );
buf \U$43079 ( \43058 , \43057 );
xor \U$43080 ( \43059 , \4287 , \4306 );
xor \U$43081 ( \43060 , \43059 , \4372 );
buf \U$43082 ( \43061 , \43060 );
buf \U$43083 ( \43062 , \43061 );
xor \U$43084 ( \43063 , \42584 , \42590 );
and \U$43085 ( \43064 , \43063 , \42606 );
and \U$43086 ( \43065 , \42584 , \42590 );
or \U$43087 ( \43066 , \43064 , \43065 );
buf \U$43088 ( \43067 , \43066 );
buf \U$43089 ( \43068 , \43067 );
xor \U$43090 ( \43069 , \43062 , \43068 );
xor \U$43091 ( \43070 , \42850 , \42856 );
and \U$43092 ( \43071 , \43070 , \42863 );
and \U$43093 ( \43072 , \42850 , \42856 );
or \U$43094 ( \43073 , \43071 , \43072 );
buf \U$43095 ( \43074 , \43073 );
buf \U$43096 ( \43075 , \43074 );
xor \U$43097 ( \43076 , \43069 , \43075 );
buf \U$43098 ( \43077 , \43076 );
buf \U$43099 ( \43078 , \43077 );
xor \U$43100 ( \43079 , \43058 , \43078 );
xor \U$43101 ( \43080 , \42837 , \42843 );
and \U$43102 ( \43081 , \43080 , \42866 );
and \U$43103 ( \43082 , \42837 , \42843 );
or \U$43104 ( \43083 , \43081 , \43082 );
buf \U$43105 ( \43084 , \43083 );
buf \U$43106 ( \43085 , \43084 );
xor \U$43107 ( \43086 , \43079 , \43085 );
buf \U$43108 ( \43087 , \43086 );
buf \U$43109 ( \43088 , \43087 );
xnor \U$43110 ( \43089 , \43023 , \43088 );
buf \U$43111 ( \43090 , \43089 );
buf \U$43112 ( \43091 , \43090 );
not \U$43113 ( \43092 , \43091 );
or \U$43114 ( \43093 , \42976 , \43092 );
buf \U$43115 ( \43094 , \43090 );
buf \U$43116 ( \43095 , \42974 );
or \U$43117 ( \43096 , \43094 , \43095 );
nand \U$43118 ( \43097 , \43093 , \43096 );
buf \U$43119 ( \43098 , \43097 );
buf \U$43120 ( \43099 , \43098 );
not \U$43121 ( \43100 , \43099 );
or \U$43122 ( \43101 , \42903 , \43100 );
not \U$43123 ( \43102 , \43098 );
buf \U$43124 ( \43103 , \43102 );
buf \U$43125 ( \43104 , \42898 );
nand \U$43126 ( \43105 , \43103 , \43104 );
buf \U$43127 ( \43106 , \43105 );
buf \U$43128 ( \43107 , \43106 );
nand \U$43129 ( \43108 , \43101 , \43107 );
buf \U$43130 ( \43109 , \43108 );
buf \U$43131 ( \43110 , \43109 );
buf \U$43132 ( \43111 , \42802 );
not \U$43133 ( \43112 , \43111 );
buf \U$43134 ( \43113 , \42874 );
not \U$43135 ( \43114 , \43113 );
or \U$43136 ( \43115 , \43112 , \43114 );
or \U$43137 ( \43116 , \42874 , \42802 );
nand \U$43138 ( \43117 , \43116 , \42556 );
buf \U$43139 ( \43118 , \43117 );
nand \U$43140 ( \43119 , \43115 , \43118 );
buf \U$43141 ( \43120 , \43119 );
buf \U$43142 ( \43121 , \43120 );
not \U$43143 ( \43122 , \43121 );
buf \U$43144 ( \43123 , \43122 );
buf \U$43145 ( \43124 , \43123 );
and \U$43146 ( \43125 , \43110 , \43124 );
not \U$43147 ( \43126 , \43110 );
buf \U$43148 ( \43127 , \43120 );
and \U$43149 ( \43128 , \43126 , \43127 );
nor \U$43150 ( \43129 , \43125 , \43128 );
buf \U$43151 ( \43130 , \43129 );
buf \U$43152 ( \43131 , \43130 );
xor \U$43153 ( \43132 , \42541 , \42550 );
and \U$43154 ( \43133 , \43132 , \42883 );
and \U$43155 ( \43134 , \42541 , \42550 );
or \U$43156 ( \43135 , \43133 , \43134 );
buf \U$43157 ( \43136 , \43135 );
buf \U$43158 ( \43137 , \43136 );
nand \U$43159 ( \43138 , \43131 , \43137 );
buf \U$43160 ( \43139 , \43138 );
buf \U$43161 ( \43140 , \43139 );
buf \U$43162 ( \43141 , \42898 );
not \U$43163 ( \43142 , \43141 );
not \U$43164 ( \43143 , \43098 );
not \U$43165 ( \43144 , \43143 );
buf \U$43166 ( \43145 , \43144 );
not \U$43167 ( \43146 , \43145 );
or \U$43168 ( \43147 , \43142 , \43146 );
buf \U$43169 ( \43148 , \42901 );
not \U$43170 ( \43149 , \43148 );
buf \U$43171 ( \43150 , \43143 );
not \U$43172 ( \43151 , \43150 );
or \U$43173 ( \43152 , \43149 , \43151 );
buf \U$43174 ( \43153 , \43120 );
nand \U$43175 ( \43154 , \43152 , \43153 );
buf \U$43176 ( \43155 , \43154 );
buf \U$43177 ( \43156 , \43155 );
nand \U$43178 ( \43157 , \43147 , \43156 );
buf \U$43179 ( \43158 , \43157 );
buf \U$43180 ( \43159 , \43158 );
not \U$43181 ( \43160 , \43159 );
buf \U$43182 ( \43161 , \43015 );
not \U$43183 ( \43162 , \43161 );
buf \U$43184 ( \43163 , \43087 );
not \U$43185 ( \43164 , \43163 );
or \U$43186 ( \43165 , \43162 , \43164 );
buf \U$43187 ( \43166 , \43087 );
buf \U$43188 ( \43167 , \43015 );
or \U$43189 ( \43168 , \43166 , \43167 );
buf \U$43190 ( \43169 , \43021 );
nand \U$43191 ( \43170 , \43168 , \43169 );
buf \U$43192 ( \43171 , \43170 );
buf \U$43193 ( \43172 , \43171 );
nand \U$43194 ( \43173 , \43165 , \43172 );
buf \U$43195 ( \43174 , \43173 );
buf \U$43196 ( \43175 , \43174 );
not \U$43197 ( \43176 , \43175 );
buf \U$43198 ( \43177 , \43176 );
buf \U$43199 ( \43178 , \43177 );
xor \U$43200 ( \43179 , \42982 , \42988 );
and \U$43201 ( \43180 , \43179 , \43013 );
and \U$43202 ( \43181 , \42982 , \42988 );
or \U$43203 ( \43182 , \43180 , \43181 );
buf \U$43204 ( \43183 , \43182 );
buf \U$43205 ( \43184 , \43183 );
xor \U$43206 ( \43185 , \43058 , \43078 );
and \U$43207 ( \43186 , \43185 , \43085 );
and \U$43208 ( \43187 , \43058 , \43078 );
or \U$43209 ( \43188 , \43186 , \43187 );
buf \U$43210 ( \43189 , \43188 );
buf \U$43211 ( \43190 , \43189 );
xor \U$43212 ( \43191 , \43184 , \43190 );
xor \U$43213 ( \43192 , \4188 , \4206 );
xor \U$43214 ( \43193 , \43192 , \4184 );
buf \U$43215 ( \43194 , \43193 );
xor \U$43216 ( \43195 , \43062 , \43068 );
and \U$43217 ( \43196 , \43195 , \43075 );
and \U$43218 ( \43197 , \43062 , \43068 );
or \U$43219 ( \43198 , \43196 , \43197 );
buf \U$43220 ( \43199 , \43198 );
buf \U$43221 ( \43200 , \43199 );
xor \U$43222 ( \43201 , \43194 , \43200 );
xor \U$43223 ( \43202 , \42917 , \42948 );
and \U$43224 ( \43203 , \43202 , \42964 );
and \U$43225 ( \43204 , \42917 , \42948 );
or \U$43226 ( \43205 , \43203 , \43204 );
buf \U$43227 ( \43206 , \43205 );
buf \U$43228 ( \43207 , \43206 );
xor \U$43229 ( \43208 , \43201 , \43207 );
buf \U$43230 ( \43209 , \43208 );
buf \U$43231 ( \43210 , \43209 );
xor \U$43232 ( \43211 , \43191 , \43210 );
buf \U$43233 ( \43212 , \43211 );
buf \U$43234 ( \43213 , \43212 );
not \U$43235 ( \43214 , \43213 );
buf \U$43236 ( \43215 , \43214 );
buf \U$43237 ( \43216 , \43215 );
not \U$43238 ( \43217 , \43216 );
buf \U$43239 ( \43218 , \42913 );
not \U$43240 ( \43219 , \43218 );
buf \U$43241 ( \43220 , \42966 );
not \U$43242 ( \43221 , \43220 );
or \U$43243 ( \43222 , \43219 , \43221 );
buf \U$43244 ( \43223 , \42966 );
buf \U$43245 ( \43224 , \42913 );
or \U$43246 ( \43225 , \43223 , \43224 );
buf \U$43247 ( \43226 , \42972 );
nand \U$43248 ( \43227 , \43225 , \43226 );
buf \U$43249 ( \43228 , \43227 );
buf \U$43250 ( \43229 , \43228 );
nand \U$43251 ( \43230 , \43222 , \43229 );
buf \U$43252 ( \43231 , \43230 );
buf \U$43253 ( \43232 , \43231 );
not \U$43254 ( \43233 , \43232 );
xor \U$43255 ( \43234 , \4286 , \4377 );
xor \U$43256 ( \43235 , \43234 , \4579 );
buf \U$43257 ( \43236 , \43235 );
buf \U$43258 ( \43237 , \43236 );
xor \U$43259 ( \43238 , \42932 , \42938 );
and \U$43260 ( \43239 , \43238 , \42945 );
and \U$43261 ( \43240 , \42932 , \42938 );
or \U$43262 ( \43241 , \43239 , \43240 );
buf \U$43263 ( \43242 , \43241 );
buf \U$43264 ( \43243 , \43242 );
xor \U$43265 ( \43244 , \4026 , \4078 );
xor \U$43266 ( \43245 , \43244 , \4140 );
buf \U$43267 ( \43246 , \43245 );
xor \U$43268 ( \43247 , \43243 , \43246 );
xor \U$43269 ( \43248 , \42993 , \42996 );
and \U$43270 ( \43249 , \43248 , \43010 );
and \U$43271 ( \43250 , \42993 , \42996 );
or \U$43272 ( \43251 , \43249 , \43250 );
buf \U$43273 ( \43252 , \43251 );
buf \U$43274 ( \43253 , \43252 );
xor \U$43275 ( \43254 , \43247 , \43253 );
buf \U$43276 ( \43255 , \43254 );
buf \U$43277 ( \43256 , \43255 );
xor \U$43278 ( \43257 , \43237 , \43256 );
xor \U$43279 ( \43258 , \3756 , \3812 );
xor \U$43280 ( \43259 , \43258 , \3883 );
buf \U$43281 ( \43260 , \43259 );
buf \U$43282 ( \43261 , \43260 );
xor \U$43283 ( \43262 , \43026 , \43039 );
and \U$43284 ( \43263 , \43262 , \43055 );
and \U$43285 ( \43264 , \43026 , \43039 );
or \U$43286 ( \43265 , \43263 , \43264 );
buf \U$43287 ( \43266 , \43265 );
buf \U$43288 ( \43267 , \43266 );
xor \U$43289 ( \43268 , \43261 , \43267 );
buf \U$43290 ( \43269 , \4246 );
buf \U$43291 ( \43270 , \4235 );
and \U$43292 ( \43271 , \43269 , \43270 );
not \U$43293 ( \43272 , \43269 );
buf \U$43294 ( \43273 , \4232 );
and \U$43295 ( \43274 , \43272 , \43273 );
nor \U$43296 ( \43275 , \43271 , \43274 );
buf \U$43297 ( \43276 , \43275 );
buf \U$43298 ( \43277 , \43276 );
buf \U$43299 ( \43278 , \4228 );
and \U$43300 ( \43279 , \43277 , \43278 );
not \U$43301 ( \43280 , \43277 );
buf \U$43302 ( \43281 , \4225 );
and \U$43303 ( \43282 , \43280 , \43281 );
nor \U$43304 ( \43283 , \43279 , \43282 );
buf \U$43305 ( \43284 , \43283 );
buf \U$43306 ( \43285 , \43284 );
xor \U$43307 ( \43286 , \43268 , \43285 );
buf \U$43308 ( \43287 , \43286 );
buf \U$43309 ( \43288 , \43287 );
xor \U$43310 ( \43289 , \43257 , \43288 );
buf \U$43311 ( \43290 , \43289 );
buf \U$43312 ( \43291 , \43290 );
not \U$43313 ( \43292 , \43291 );
buf \U$43314 ( \43293 , \43292 );
buf \U$43315 ( \43294 , \43293 );
not \U$43316 ( \43295 , \43294 );
or \U$43317 ( \43296 , \43233 , \43295 );
buf \U$43318 ( \43297 , \43231 );
not \U$43319 ( \43298 , \43297 );
buf \U$43320 ( \43299 , \43290 );
nand \U$43321 ( \43300 , \43298 , \43299 );
buf \U$43322 ( \43301 , \43300 );
buf \U$43323 ( \43302 , \43301 );
nand \U$43324 ( \43303 , \43296 , \43302 );
buf \U$43325 ( \43304 , \43303 );
buf \U$43326 ( \43305 , \43304 );
not \U$43327 ( \43306 , \43305 );
and \U$43328 ( \43307 , \43217 , \43306 );
buf \U$43329 ( \43308 , \43215 );
buf \U$43330 ( \43309 , \43304 );
and \U$43331 ( \43310 , \43308 , \43309 );
nor \U$43332 ( \43311 , \43307 , \43310 );
buf \U$43333 ( \43312 , \43311 );
buf \U$43334 ( \43313 , \43312 );
xor \U$43335 ( \43314 , \43178 , \43313 );
buf \U$43336 ( \43315 , \42973 );
not \U$43337 ( \43316 , \43315 );
buf \U$43338 ( \43317 , \43090 );
not \U$43339 ( \43318 , \43317 );
or \U$43340 ( \43319 , \43316 , \43318 );
buf \U$43341 ( \43320 , \42908 );
nand \U$43342 ( \43321 , \43319 , \43320 );
buf \U$43343 ( \43322 , \43321 );
buf \U$43344 ( \43323 , \43322 );
or \U$43345 ( \43324 , \43090 , \42973 );
buf \U$43346 ( \43325 , \43324 );
and \U$43347 ( \43326 , \43323 , \43325 );
buf \U$43348 ( \43327 , \43326 );
buf \U$43349 ( \43328 , \43327 );
xor \U$43350 ( \43329 , \43314 , \43328 );
buf \U$43351 ( \43330 , \43329 );
buf \U$43352 ( \43331 , \43330 );
nand \U$43353 ( \43332 , \43160 , \43331 );
buf \U$43354 ( \43333 , \43332 );
buf \U$43355 ( \43334 , \43333 );
and \U$43356 ( \43335 , \42893 , \43140 , \43334 );
buf \U$43357 ( \43336 , \43335 );
buf \U$43358 ( \43337 , \43336 );
and \U$43359 ( \43338 , \41972 , \43337 );
buf \U$43360 ( \43339 , \43338 );
buf \U$43361 ( \43340 , \43339 );
xor \U$43362 ( \43341 , \43261 , \43267 );
and \U$43363 ( \43342 , \43341 , \43285 );
and \U$43364 ( \43343 , \43261 , \43267 );
or \U$43365 ( \43344 , \43342 , \43343 );
buf \U$43366 ( \43345 , \43344 );
buf \U$43367 ( \43346 , \43345 );
xor \U$43368 ( \43347 , \4266 , \4270 );
xor \U$43369 ( \43348 , \43347 , \4584 );
buf \U$43370 ( \43349 , \43348 );
buf \U$43371 ( \43350 , \43349 );
xor \U$43372 ( \43351 , \43346 , \43350 );
xor \U$43373 ( \43352 , \43194 , \43200 );
and \U$43374 ( \43353 , \43352 , \43207 );
and \U$43375 ( \43354 , \43194 , \43200 );
or \U$43376 ( \43355 , \43353 , \43354 );
buf \U$43377 ( \43356 , \43355 );
buf \U$43378 ( \43357 , \43356 );
xor \U$43379 ( \43358 , \43351 , \43357 );
buf \U$43380 ( \43359 , \43358 );
xor \U$43381 ( \43360 , \43237 , \43256 );
and \U$43382 ( \43361 , \43360 , \43288 );
and \U$43383 ( \43362 , \43237 , \43256 );
or \U$43384 ( \43363 , \43361 , \43362 );
buf \U$43385 ( \43364 , \43363 );
buf \U$43386 ( \43365 , \43364 );
xor \U$43387 ( \43366 , \43243 , \43246 );
and \U$43388 ( \43367 , \43366 , \43253 );
and \U$43389 ( \43368 , \43243 , \43246 );
or \U$43390 ( \43369 , \43367 , \43368 );
buf \U$43391 ( \43370 , \43369 );
buf \U$43392 ( \43371 , \43370 );
xor \U$43393 ( \43372 , \4144 , \4148 );
xor \U$43394 ( \43373 , \43372 , \4153 );
buf \U$43395 ( \43374 , \43373 );
buf \U$43396 ( \43375 , \43374 );
xor \U$43397 ( \43376 , \43371 , \43375 );
xor \U$43398 ( \43377 , \4213 , \4253 );
xor \U$43399 ( \43378 , \43377 , \4257 );
buf \U$43400 ( \43379 , \43378 );
buf \U$43401 ( \43380 , \43379 );
xor \U$43402 ( \43381 , \43376 , \43380 );
buf \U$43403 ( \43382 , \43381 );
buf \U$43404 ( \43383 , \43382 );
xor \U$43405 ( \43384 , \43365 , \43383 );
xor \U$43406 ( \43385 , \43184 , \43190 );
and \U$43407 ( \43386 , \43385 , \43210 );
and \U$43408 ( \43387 , \43184 , \43190 );
or \U$43409 ( \43388 , \43386 , \43387 );
buf \U$43410 ( \43389 , \43388 );
buf \U$43411 ( \43390 , \43389 );
xor \U$43412 ( \43391 , \43384 , \43390 );
buf \U$43413 ( \43392 , \43391 );
xor \U$43414 ( \43393 , \43359 , \43392 );
buf \U$43415 ( \43394 , \43231 );
not \U$43416 ( \43395 , \43394 );
buf \U$43417 ( \43396 , \43290 );
not \U$43418 ( \43397 , \43396 );
or \U$43419 ( \43398 , \43395 , \43397 );
buf \U$43420 ( \43399 , \43290 );
buf \U$43421 ( \43400 , \43231 );
or \U$43422 ( \43401 , \43399 , \43400 );
buf \U$43423 ( \43402 , \43212 );
nand \U$43424 ( \43403 , \43401 , \43402 );
buf \U$43425 ( \43404 , \43403 );
buf \U$43426 ( \43405 , \43404 );
nand \U$43427 ( \43406 , \43398 , \43405 );
buf \U$43428 ( \43407 , \43406 );
xnor \U$43429 ( \43408 , \43393 , \43407 );
buf \U$43430 ( \43409 , \43408 );
xor \U$43431 ( \43410 , \43178 , \43313 );
and \U$43432 ( \43411 , \43410 , \43328 );
and \U$43433 ( \43412 , \43178 , \43313 );
or \U$43434 ( \43413 , \43411 , \43412 );
buf \U$43435 ( \43414 , \43413 );
buf \U$43436 ( \43415 , \43414 );
nand \U$43437 ( \43416 , \43409 , \43415 );
buf \U$43438 ( \43417 , \43416 );
buf \U$43439 ( \43418 , \43417 );
xor \U$43440 ( \43419 , \43359 , \43392 );
and \U$43441 ( \43420 , \43419 , \43407 );
and \U$43442 ( \43421 , \43359 , \43392 );
or \U$43443 ( \43422 , \43420 , \43421 );
buf \U$43444 ( \43423 , \43422 );
xor \U$43445 ( \43424 , \4262 , \4589 );
xor \U$43446 ( \43425 , \43424 , \4594 );
buf \U$43447 ( \43426 , \43425 );
buf \U$43448 ( \43427 , \43426 );
xor \U$43449 ( \43428 , \43365 , \43383 );
and \U$43450 ( \43429 , \43428 , \43390 );
and \U$43451 ( \43430 , \43365 , \43383 );
or \U$43452 ( \43431 , \43429 , \43430 );
buf \U$43453 ( \43432 , \43431 );
buf \U$43454 ( \43433 , \43432 );
xor \U$43455 ( \43434 , \43427 , \43433 );
xor \U$43456 ( \43435 , \43371 , \43375 );
and \U$43457 ( \43436 , \43435 , \43380 );
and \U$43458 ( \43437 , \43371 , \43375 );
or \U$43459 ( \43438 , \43436 , \43437 );
buf \U$43460 ( \43439 , \43438 );
buf \U$43461 ( \43440 , \43439 );
xor \U$43462 ( \43441 , \4158 , \4162 );
xor \U$43463 ( \43442 , \43441 , \4166 );
buf \U$43464 ( \43443 , \43442 );
buf \U$43465 ( \43444 , \43443 );
xor \U$43466 ( \43445 , \43440 , \43444 );
xor \U$43467 ( \43446 , \43346 , \43350 );
and \U$43468 ( \43447 , \43446 , \43357 );
and \U$43469 ( \43448 , \43346 , \43350 );
or \U$43470 ( \43449 , \43447 , \43448 );
buf \U$43471 ( \43450 , \43449 );
buf \U$43472 ( \43451 , \43450 );
xor \U$43473 ( \43452 , \43445 , \43451 );
buf \U$43474 ( \43453 , \43452 );
buf \U$43475 ( \43454 , \43453 );
xor \U$43476 ( \43455 , \43434 , \43454 );
buf \U$43477 ( \43456 , \43455 );
buf \U$43478 ( \43457 , \43456 );
or \U$43479 ( \43458 , \43423 , \43457 );
buf \U$43480 ( \43459 , \43458 );
buf \U$43481 ( \43460 , \43459 );
nand \U$43482 ( \43461 , \43418 , \43460 );
buf \U$43483 ( \43462 , \43461 );
buf \U$43484 ( \43463 , \43462 );
xor \U$43485 ( \43464 , \43440 , \43444 );
and \U$43486 ( \43465 , \43464 , \43451 );
and \U$43487 ( \43466 , \43440 , \43444 );
or \U$43488 ( \43467 , \43465 , \43466 );
buf \U$43489 ( \43468 , \43467 );
buf \U$43490 ( \43469 , \43468 );
xor \U$43491 ( \43470 , \3903 , \3922 );
xor \U$43492 ( \43471 , \43470 , \3932 );
buf \U$43493 ( \43472 , \43471 );
buf \U$43494 ( \43473 , \43472 );
xor \U$43495 ( \43474 , \43469 , \43473 );
buf \U$43496 ( \43475 , \4598 );
not \U$43497 ( \43476 , \43475 );
xnor \U$43498 ( \43477 , \4170 , \4175 );
buf \U$43499 ( \43478 , \43477 );
not \U$43500 ( \43479 , \43478 );
or \U$43501 ( \43480 , \43476 , \43479 );
buf \U$43502 ( \43481 , \43477 );
buf \U$43503 ( \43482 , \4598 );
or \U$43504 ( \43483 , \43481 , \43482 );
nand \U$43505 ( \43484 , \43480 , \43483 );
buf \U$43506 ( \43485 , \43484 );
buf \U$43507 ( \43486 , \43485 );
xor \U$43508 ( \43487 , \43474 , \43486 );
buf \U$43509 ( \43488 , \43487 );
buf \U$43510 ( \43489 , \43488 );
xor \U$43511 ( \43490 , \43427 , \43433 );
and \U$43512 ( \43491 , \43490 , \43454 );
and \U$43513 ( \43492 , \43427 , \43433 );
or \U$43514 ( \43493 , \43491 , \43492 );
buf \U$43515 ( \43494 , \43493 );
buf \U$43516 ( \43495 , \43494 );
nor \U$43517 ( \43496 , \43489 , \43495 );
buf \U$43518 ( \43497 , \43496 );
buf \U$43519 ( \43498 , \43497 );
nor \U$43520 ( \43499 , \43463 , \43498 );
buf \U$43521 ( \43500 , \43499 );
buf \U$43522 ( \43501 , \43500 );
xor \U$43523 ( \43502 , \3949 , \4605 );
xor \U$43524 ( \43503 , \43502 , \4610 );
buf \U$43525 ( \43504 , \43503 );
buf \U$43526 ( \43505 , \43504 );
xor \U$43527 ( \43506 , \43469 , \43473 );
and \U$43528 ( \43507 , \43506 , \43486 );
and \U$43529 ( \43508 , \43469 , \43473 );
or \U$43530 ( \43509 , \43507 , \43508 );
buf \U$43531 ( \43510 , \43509 );
buf \U$43532 ( \43511 , \43510 );
or \U$43533 ( \43512 , \43505 , \43511 );
buf \U$43534 ( \43513 , \43512 );
buf \U$43535 ( \43514 , \43513 );
and \U$43536 ( \43515 , \43501 , \43514 );
buf \U$43537 ( \43516 , \43515 );
buf \U$43538 ( \43517 , \43516 );
nand \U$43539 ( \43518 , \43340 , \43517 );
buf \U$43540 ( \43519 , \43518 );
buf \U$43541 ( \43520 , \43519 );
not \U$43542 ( \43521 , \43520 );
buf \U$43543 ( \43522 , \43521 );
buf \U$43544 ( \43523 , \43522 );
nand \U$43545 ( \43524 , \35571 , \43523 );
buf \U$43546 ( \43525 , \43524 );
buf \U$43547 ( \43526 , \43525 );
buf \U$43548 ( \43527 , \43139 );
not \U$43549 ( \43528 , \43527 );
buf \U$43550 ( \43529 , \42886 );
not \U$43551 ( \43530 , \43529 );
buf \U$43552 ( \43531 , \43530 );
buf \U$43553 ( \43532 , \43531 );
buf \U$43554 ( \43533 , \42519 );
buf \U$43555 ( \43534 , \41977 );
nand \U$43556 ( \43535 , \43533 , \43534 );
buf \U$43557 ( \43536 , \43535 );
buf \U$43558 ( \43537 , \43536 );
or \U$43559 ( \43538 , \43532 , \43537 );
buf \U$43560 ( \43539 , \42885 );
not \U$43561 ( \43540 , \43539 );
buf \U$43562 ( \43541 , \42531 );
nand \U$43563 ( \43542 , \43540 , \43541 );
buf \U$43564 ( \43543 , \43542 );
buf \U$43565 ( \43544 , \43543 );
nand \U$43566 ( \43545 , \43538 , \43544 );
buf \U$43567 ( \43546 , \43545 );
buf \U$43568 ( \43547 , \43546 );
not \U$43569 ( \43548 , \43547 );
or \U$43570 ( \43549 , \43528 , \43548 );
buf \U$43571 ( \43550 , \43130 );
buf \U$43572 ( \43551 , \43136 );
or \U$43573 ( \43552 , \43550 , \43551 );
buf \U$43574 ( \43553 , \43552 );
buf \U$43575 ( \43554 , \43553 );
nand \U$43576 ( \43555 , \43549 , \43554 );
buf \U$43577 ( \43556 , \43555 );
buf \U$43578 ( \43557 , \43556 );
buf \U$43579 ( \43558 , \43333 );
buf \U$43580 ( \43559 , \43558 );
nand \U$43581 ( \43560 , \43557 , \43559 );
buf \U$43582 ( \43561 , \43560 );
buf \U$43583 ( \43562 , \43561 );
buf \U$43584 ( \43563 , \43330 );
not \U$43585 ( \43564 , \43563 );
buf \U$43586 ( \43565 , \43158 );
nand \U$43587 ( \43566 , \43564 , \43565 );
buf \U$43588 ( \43567 , \43566 );
buf \U$43589 ( \43568 , \43567 );
nand \U$43590 ( \43569 , \43562 , \43568 );
buf \U$43591 ( \43570 , \43569 );
buf \U$43592 ( \43571 , \43570 );
not \U$43593 ( \43572 , \43571 );
buf \U$43594 ( \43573 , \43139 );
buf \U$43595 ( \43574 , \43333 );
and \U$43596 ( \43575 , \43573 , \43574 );
buf \U$43597 ( \43576 , \43575 );
buf \U$43598 ( \43577 , \43576 );
buf \U$43599 ( \43578 , \41634 );
not \U$43600 ( \43579 , \43578 );
buf \U$43601 ( \43580 , \43579 );
buf \U$43602 ( \43581 , \43580 );
and \U$43603 ( \43582 , \43577 , \43581 );
buf \U$43604 ( \43583 , \43582 );
buf \U$43605 ( \43584 , \43583 );
buf \U$43606 ( \43585 , \40147 );
buf \U$43607 ( \43586 , \42889 );
nor \U$43608 ( \43587 , \43585 , \43586 );
buf \U$43609 ( \43588 , \43587 );
buf \U$43610 ( \43589 , \43588 );
buf \U$43611 ( \43590 , \41889 );
not \U$43612 ( \43591 , \43590 );
buf \U$43613 ( \43592 , \41884 );
nand \U$43614 ( \43593 , \43591 , \43592 );
buf \U$43615 ( \43594 , \43593 );
buf \U$43616 ( \43595 , \43594 );
not \U$43617 ( \43596 , \43595 );
buf \U$43620 ( \43597 , \41863 );
buf \U$43621 ( \43598 , \43597 );
nand \U$43622 ( \43599 , \43596 , \43598 );
buf \U$43623 ( \43600 , \43599 );
buf \U$43624 ( \43601 , \43600 );
buf \U$43625 ( \43602 , \41798 );
buf \U$43626 ( \43603 , \41860 );
or \U$43627 ( \43604 , \43602 , \43603 );
buf \U$43628 ( \43605 , \43604 );
buf \U$43629 ( \43606 , \43605 );
nand \U$43630 ( \43607 , \43601 , \43606 );
buf \U$43631 ( \43608 , \43607 );
buf \U$43632 ( \43609 , \43608 );
buf \U$43633 ( \43610 , \41945 );
buf \U$43634 ( \43611 , \41968 );
and \U$43635 ( \43612 , \43610 , \43611 );
buf \U$43636 ( \43613 , \43612 );
buf \U$43637 ( \43614 , \43613 );
nand \U$43638 ( \43615 , \43584 , \43589 , \43609 , \43614 );
buf \U$43639 ( \43616 , \43615 );
buf \U$43640 ( \43617 , \43616 );
buf \U$43641 ( \43618 , \43583 );
buf \U$43642 ( \43619 , \43588 );
buf \U$43643 ( \43620 , \41965 );
not \U$43644 ( \43621 , \43620 );
buf \U$43645 ( \43622 , \41957 );
nand \U$43646 ( \43623 , \43621 , \43622 );
buf \U$43647 ( \43624 , \43623 );
buf \U$43648 ( \43625 , \43624 );
not \U$43649 ( \43626 , \43625 );
buf \U$43650 ( \43627 , \41945 );
nand \U$43651 ( \43628 , \43626 , \43627 );
buf \U$43652 ( \43629 , \43628 );
buf \U$43653 ( \43630 , \43629 );
buf \U$43654 ( \43631 , \41942 );
not \U$43655 ( \43632 , \43631 );
buf \U$43656 ( \43633 , \41934 );
nand \U$43657 ( \43634 , \43632 , \43633 );
buf \U$43658 ( \43635 , \43634 );
buf \U$43659 ( \43636 , \43635 );
nand \U$43660 ( \43637 , \43630 , \43636 );
buf \U$43661 ( \43638 , \43637 );
buf \U$43662 ( \43639 , \43638 );
nand \U$43663 ( \43640 , \43618 , \43619 , \43639 );
buf \U$43664 ( \43641 , \43640 );
buf \U$43665 ( \43642 , \43641 );
buf \U$43666 ( \43643 , \43580 );
not \U$43667 ( \43644 , \43643 );
buf \U$43668 ( \43645 , \39855 );
not \U$43669 ( \43646 , \43645 );
buf \U$43670 ( \43647 , \43646 );
buf \U$43671 ( \43648 , \43647 );
buf \U$43672 ( \43649 , \39858 );
not \U$43673 ( \43650 , \43649 );
buf \U$43674 ( \43651 , \43650 );
buf \U$43675 ( \43652 , \43651 );
buf \U$43676 ( \43653 , \40138 );
nand \U$43677 ( \43654 , \43652 , \43653 );
buf \U$43678 ( \43655 , \43654 );
buf \U$43679 ( \43656 , \43655 );
or \U$43680 ( \43657 , \43648 , \43656 );
buf \U$43681 ( \43658 , \39852 );
not \U$43682 ( \43659 , \43658 );
buf \U$43683 ( \43660 , \39110 );
nand \U$43684 ( \43661 , \43659 , \43660 );
buf \U$43685 ( \43662 , \43661 );
buf \U$43686 ( \43663 , \43662 );
nand \U$43687 ( \43664 , \43657 , \43663 );
buf \U$43688 ( \43665 , \43664 );
buf \U$43689 ( \43666 , \43665 );
not \U$43690 ( \43667 , \43666 );
or \U$43691 ( \43668 , \43644 , \43667 );
not \U$43692 ( \43669 , \41605 );
buf \U$43693 ( \43670 , \41628 );
not \U$43694 ( \43671 , \43670 );
buf \U$43695 ( \43672 , \41624 );
nand \U$43696 ( \43673 , \43671 , \43672 );
buf \U$43697 ( \43674 , \43673 );
not \U$43698 ( \43675 , \43674 );
and \U$43699 ( \43676 , \43669 , \43675 );
buf \U$43700 ( \43677 , \41539 );
buf \U$43701 ( \43678 , \41602 );
and \U$43702 ( \43679 , \43677 , \43678 );
buf \U$43703 ( \43680 , \43679 );
nor \U$43704 ( \43681 , \43676 , \43680 );
buf \U$43705 ( \43682 , \43681 );
nand \U$43706 ( \43683 , \43668 , \43682 );
buf \U$43707 ( \43684 , \43683 );
buf \U$43708 ( \43685 , \43684 );
buf \U$43709 ( \43686 , \43336 );
nand \U$43710 ( \43687 , \43685 , \43686 );
buf \U$43711 ( \43688 , \43687 );
buf \U$43712 ( \43689 , \43688 );
nand \U$43713 ( \43690 , \43572 , \43617 , \43642 , \43689 );
buf \U$43714 ( \43691 , \43690 );
buf \U$43715 ( \43692 , \43691 );
buf \U$43716 ( \43693 , \43516 );
and \U$43717 ( \43694 , \43692 , \43693 );
buf \U$43718 ( \43695 , \43513 );
not \U$43719 ( \43696 , \43695 );
buf \U$43720 ( \43697 , \43497 );
not \U$43721 ( \43698 , \43697 );
buf \U$43722 ( \43699 , \43698 );
buf \U$43723 ( \43700 , \43699 );
not \U$43724 ( \43701 , \43700 );
buf \U$43725 ( \43702 , \43459 );
not \U$43726 ( \43703 , \43702 );
buf \U$43727 ( \43704 , \43408 );
buf \U$43728 ( \43705 , \43414 );
nor \U$43729 ( \43706 , \43704 , \43705 );
buf \U$43730 ( \43707 , \43706 );
buf \U$43731 ( \43708 , \43707 );
not \U$43732 ( \43709 , \43708 );
or \U$43733 ( \43710 , \43703 , \43709 );
buf \U$43734 ( \43711 , \43456 );
buf \U$43735 ( \43712 , \43422 );
nand \U$43736 ( \43713 , \43711 , \43712 );
buf \U$43737 ( \43714 , \43713 );
buf \U$43738 ( \43715 , \43714 );
nand \U$43739 ( \43716 , \43710 , \43715 );
buf \U$43740 ( \43717 , \43716 );
buf \U$43741 ( \43718 , \43717 );
not \U$43742 ( \43719 , \43718 );
or \U$43743 ( \43720 , \43701 , \43719 );
buf \U$43744 ( \43721 , \43488 );
buf \U$43745 ( \43722 , \43494 );
nand \U$43746 ( \43723 , \43721 , \43722 );
buf \U$43747 ( \43724 , \43723 );
buf \U$43748 ( \43725 , \43724 );
nand \U$43749 ( \43726 , \43720 , \43725 );
buf \U$43750 ( \43727 , \43726 );
buf \U$43751 ( \43728 , \43727 );
not \U$43752 ( \43729 , \43728 );
or \U$43753 ( \43730 , \43696 , \43729 );
buf \U$43754 ( \43731 , \43504 );
buf \U$43755 ( \43732 , \43510 );
nand \U$43756 ( \43733 , \43731 , \43732 );
buf \U$43757 ( \43734 , \43733 );
buf \U$43758 ( \43735 , \43734 );
nand \U$43759 ( \43736 , \43730 , \43735 );
buf \U$43760 ( \43737 , \43736 );
buf \U$43761 ( \43738 , \43737 );
nor \U$43762 ( \43739 , \43694 , \43738 );
buf \U$43763 ( \43740 , \43739 );
buf \U$43764 ( \43741 , \43740 );
nand \U$43765 ( \43742 , \43526 , \43741 );
buf \U$43766 ( \43743 , \43742 );
buf \U$43767 ( \43744 , \43743 );
not \U$43768 ( \43745 , \43744 );
buf \U$43769 ( \43746 , \43745 );
buf \U$43770 ( \43747 , \43746 );
buf \U$43771 ( \43748 , \25932 );
not \U$43772 ( \43749 , \43748 );
buf \U$43773 ( \43750 , \43749 );
buf \U$43774 ( \43751 , \43750 );
buf \U$43775 ( \43752 , \27843 );
not \U$43776 ( \43753 , \43752 );
buf \U$43777 ( \43754 , \43753 );
buf \U$43778 ( \43755 , \43754 );
buf \U$43779 ( \43756 , \23729 );
buf \U$43780 ( \43757 , \21568 );
buf \U$43781 ( \43758 , \19303 );
buf \U$43782 ( \43759 , \20361 );
or \U$43783 ( \43760 , \43758 , \43759 );
buf \U$43784 ( \43761 , \43760 );
buf \U$43785 ( \43762 , \43761 );
and \U$43786 ( \43763 , \43757 , \43762 );
buf \U$43787 ( \43764 , \43763 );
buf \U$43788 ( \43765 , \43764 );
and \U$43789 ( \43766 , \43751 , \43755 , \43756 , \43765 );
buf \U$43790 ( \43767 , \43766 );
buf \U$43791 ( \43768 , \43767 );
not \U$43792 ( \43769 , \43768 );
buf \U$43793 ( \43770 , \35516 );
nor \U$43794 ( \43771 , \43769 , \43770 );
buf \U$43795 ( \43772 , \43771 );
buf \U$43796 ( \43773 , \43772 );
not \U$43797 ( \43774 , \43773 );
buf \U$43798 ( \43775 , \43519 );
nor \U$43799 ( \43776 , \43774 , \43775 );
buf \U$43800 ( \43777 , \43776 );
buf \U$43801 ( \43778 , \43777 );
not \U$43802 ( \43779 , \15608 );
not \U$43803 ( \43780 , \43779 );
buf \U$43804 ( \43781 , \43780 );
not \U$43805 ( \43782 , \43781 );
buf \U$43806 ( \43783 , RIc0d8230_26);
buf \U$43807 ( \43784 , RIc0db188_127);
xor \U$43808 ( \43785 , \43783 , \43784 );
buf \U$43809 ( \43786 , \43785 );
not \U$43810 ( \43787 , \43786 );
or \U$43811 ( \43788 , \43782 , \43787 );
buf \U$43812 ( \43789 , RIc0d81b8_25);
buf \U$43813 ( \43790 , RIc0db188_127);
xnor \U$43814 ( \43791 , \43789 , \43790 );
buf \U$43815 ( \43792 , \43791 );
or \U$43816 ( \43793 , \12647 , \43792 );
nand \U$43817 ( \43794 , \43788 , \43793 );
buf \U$43818 ( \43795 , \43794 );
buf \U$43819 ( \43796 , RIc0d9130_58);
buf \U$43820 ( \43797 , RIc0da288_95);
xor \U$43821 ( \43798 , \43796 , \43797 );
buf \U$43822 ( \43799 , \43798 );
buf \U$43823 ( \43800 , \43799 );
not \U$43824 ( \43801 , \43800 );
buf \U$43825 ( \43802 , \330 );
not \U$43826 ( \43803 , \43802 );
or \U$43827 ( \43804 , \43801 , \43803 );
buf \U$43828 ( \43805 , \344 );
xor \U$43829 ( \43806 , RIc0da288_95, RIc0d90b8_57);
buf \U$43830 ( \43807 , \43806 );
nand \U$43831 ( \43808 , \43805 , \43807 );
buf \U$43832 ( \43809 , \43808 );
buf \U$43833 ( \43810 , \43809 );
nand \U$43834 ( \43811 , \43804 , \43810 );
buf \U$43835 ( \43812 , \43811 );
buf \U$43836 ( \43813 , \43812 );
xor \U$43837 ( \43814 , \43795 , \43813 );
buf \U$43838 ( \43815 , \22595 );
buf \U$43839 ( \43816 , RIc0d87d0_38);
buf \U$43840 ( \43817 , RIc0dabe8_115);
xnor \U$43841 ( \43818 , \43816 , \43817 );
buf \U$43842 ( \43819 , \43818 );
buf \U$43843 ( \43820 , \43819 );
or \U$43844 ( \43821 , \43815 , \43820 );
buf \U$43845 ( \43822 , \29865 );
buf \U$43846 ( \43823 , RIc0d8758_37);
buf \U$43847 ( \43824 , RIc0dabe8_115);
xor \U$43848 ( \43825 , \43823 , \43824 );
buf \U$43849 ( \43826 , \43825 );
buf \U$43850 ( \43827 , \43826 );
not \U$43851 ( \43828 , \43827 );
buf \U$43852 ( \43829 , \43828 );
buf \U$43853 ( \43830 , \43829 );
or \U$43854 ( \43831 , \43822 , \43830 );
nand \U$43855 ( \43832 , \43821 , \43831 );
buf \U$43856 ( \43833 , \43832 );
buf \U$43857 ( \43834 , \43833 );
and \U$43858 ( \43835 , \43814 , \43834 );
and \U$43859 ( \43836 , \43795 , \43813 );
or \U$43860 ( \43837 , \43835 , \43836 );
buf \U$43861 ( \43838 , \43837 );
buf \U$43862 ( \43839 , \43838 );
buf \U$43863 ( \43840 , \634 );
buf \U$43864 ( \43841 , RIc0d9400_64);
not \U$43865 ( \43842 , \43841 );
buf \U$43866 ( \43843 , \43842 );
buf \U$43867 ( \43844 , \43843 );
nor \U$43868 ( \43845 , \43840 , \43844 );
buf \U$43869 ( \43846 , \43845 );
buf \U$43870 ( \43847 , \43846 );
buf \U$43871 ( \43848 , \43826 );
not \U$43872 ( \43849 , \43848 );
buf \U$43873 ( \43850 , \14186 );
not \U$43874 ( \43851 , \43850 );
or \U$43875 ( \43852 , \43849 , \43851 );
buf \U$43876 ( \43853 , \14690 );
xor \U$43877 ( \43854 , RIc0dabe8_115, RIc0d86e0_36);
buf \U$43878 ( \43855 , \43854 );
nand \U$43879 ( \43856 , \43853 , \43855 );
buf \U$43880 ( \43857 , \43856 );
buf \U$43881 ( \43858 , \43857 );
nand \U$43882 ( \43859 , \43852 , \43858 );
buf \U$43883 ( \43860 , \43859 );
buf \U$43884 ( \43861 , \43860 );
xor \U$43885 ( \43862 , \43847 , \43861 );
buf \U$43886 ( \43863 , \521 );
buf \U$43887 ( \43864 , RIc0da0a8_91);
buf \U$43888 ( \43865 , RIc0d9298_61);
xnor \U$43889 ( \43866 , \43864 , \43865 );
buf \U$43890 ( \43867 , \43866 );
buf \U$43891 ( \43868 , \43867 );
or \U$43892 ( \43869 , \43863 , \43868 );
buf \U$43893 ( \43870 , \530 );
buf \U$43894 ( \43871 , RIc0d9220_60);
buf \U$43895 ( \43872 , RIc0da0a8_91);
xnor \U$43896 ( \43873 , \43871 , \43872 );
buf \U$43897 ( \43874 , \43873 );
buf \U$43898 ( \43875 , \43874 );
or \U$43899 ( \43876 , \43870 , \43875 );
nand \U$43900 ( \43877 , \43869 , \43876 );
buf \U$43901 ( \43878 , \43877 );
buf \U$43902 ( \43879 , \43878 );
xor \U$43903 ( \43880 , \43862 , \43879 );
buf \U$43904 ( \43881 , \43880 );
buf \U$43905 ( \43882 , \43881 );
xor \U$43906 ( \43883 , \43839 , \43882 );
xor \U$43907 ( \43884 , RIc0dadc8_119, RIc0d8578_33);
buf \U$43908 ( \43885 , \43884 );
not \U$43909 ( \43886 , \43885 );
buf \U$43910 ( \43887 , \13181 );
not \U$43911 ( \43888 , \43887 );
or \U$43912 ( \43889 , \43886 , \43888 );
buf \U$43913 ( \43890 , \13005 );
buf \U$43914 ( \43891 , RIc0d8500_32);
buf \U$43915 ( \43892 , RIc0dadc8_119);
xor \U$43916 ( \43893 , \43891 , \43892 );
buf \U$43917 ( \43894 , \43893 );
buf \U$43918 ( \43895 , \43894 );
nand \U$43919 ( \43896 , \43890 , \43895 );
buf \U$43920 ( \43897 , \43896 );
buf \U$43921 ( \43898 , \43897 );
nand \U$43922 ( \43899 , \43889 , \43898 );
buf \U$43923 ( \43900 , \43899 );
buf \U$43924 ( \43901 , \43900 );
not \U$43925 ( \43902 , \43901 );
buf \U$43926 ( \43903 , \21959 );
not \U$43927 ( \43904 , \43903 );
buf \U$43928 ( \43905 , \43904 );
buf \U$43929 ( \43906 , \43905 );
not \U$43930 ( \43907 , \43906 );
buf \U$43931 ( \43908 , RIc0da918_109);
buf \U$43932 ( \43909 , RIc0d8a28_43);
xnor \U$43933 ( \43910 , \43908 , \43909 );
buf \U$43934 ( \43911 , \43910 );
buf \U$43935 ( \43912 , \43911 );
not \U$43936 ( \43913 , \43912 );
and \U$43937 ( \43914 , \43907 , \43913 );
buf \U$43938 ( \43915 , \20211 );
not \U$43939 ( \43916 , \43915 );
xnor \U$43940 ( \43917 , RIc0da918_109, RIc0d89b0_42);
buf \U$43941 ( \43918 , \43917 );
nor \U$43942 ( \43919 , \43916 , \43918 );
buf \U$43943 ( \43920 , \43919 );
buf \U$43944 ( \43921 , \43920 );
nor \U$43945 ( \43922 , \43914 , \43921 );
buf \U$43946 ( \43923 , \43922 );
buf \U$43947 ( \43924 , \43923 );
not \U$43948 ( \43925 , \43924 );
or \U$43949 ( \43926 , \43902 , \43925 );
buf \U$43950 ( \43927 , \43900 );
buf \U$43951 ( \43928 , \43923 );
or \U$43952 ( \43929 , \43927 , \43928 );
nand \U$43953 ( \43930 , \43926 , \43929 );
buf \U$43954 ( \43931 , \43930 );
buf \U$43955 ( \43932 , \43931 );
buf \U$43956 ( \43933 , RIc0d9fb8_89);
buf \U$43957 ( \43934 , RIc0d9388_63);
and \U$43958 ( \43935 , \43933 , \43934 );
not \U$43959 ( \43936 , \43933 );
buf \U$43960 ( \43937 , RIc0d9388_63);
not \U$43961 ( \43938 , \43937 );
buf \U$43962 ( \43939 , \43938 );
buf \U$43963 ( \43940 , \43939 );
and \U$43964 ( \43941 , \43936 , \43940 );
nor \U$43965 ( \43942 , \43935 , \43941 );
buf \U$43966 ( \43943 , \43942 );
buf \U$43967 ( \43944 , \43943 );
not \U$43968 ( \43945 , \43944 );
buf \U$43969 ( \43946 , \2038 );
not \U$43970 ( \43947 , \43946 );
or \U$43971 ( \43948 , \43945 , \43947 );
buf \U$43972 ( \43949 , \846 );
buf \U$43973 ( \43950 , RIc0d9310_62);
buf \U$43974 ( \43951 , RIc0d9fb8_89);
xor \U$43975 ( \43952 , \43950 , \43951 );
buf \U$43976 ( \43953 , \43952 );
buf \U$43977 ( \43954 , \43953 );
nand \U$43978 ( \43955 , \43949 , \43954 );
buf \U$43979 ( \43956 , \43955 );
buf \U$43980 ( \43957 , \43956 );
nand \U$43981 ( \43958 , \43948 , \43957 );
buf \U$43982 ( \43959 , \43958 );
buf \U$43983 ( \43960 , \43959 );
xor \U$43984 ( \43961 , \43932 , \43960 );
buf \U$43985 ( \43962 , \43961 );
buf \U$43986 ( \43963 , \43962 );
and \U$43987 ( \43964 , \43883 , \43963 );
and \U$43988 ( \43965 , \43839 , \43882 );
or \U$43989 ( \43966 , \43964 , \43965 );
buf \U$43990 ( \43967 , \43966 );
buf \U$43991 ( \43968 , \43806 );
not \U$43992 ( \43969 , \43968 );
buf \U$43993 ( \43970 , \3714 );
not \U$43994 ( \43971 , \43970 );
or \U$43995 ( \43972 , \43969 , \43971 );
buf \U$43996 ( \43973 , \343 );
buf \U$43997 ( \43974 , RIc0da288_95);
buf \U$43998 ( \43975 , RIc0d9040_56);
xor \U$43999 ( \43976 , \43974 , \43975 );
buf \U$44000 ( \43977 , \43976 );
buf \U$44001 ( \43978 , \43977 );
nand \U$44002 ( \43979 , \43973 , \43978 );
buf \U$44003 ( \43980 , \43979 );
buf \U$44004 ( \43981 , \43980 );
nand \U$44005 ( \43982 , \43972 , \43981 );
buf \U$44006 ( \43983 , \43982 );
buf \U$44007 ( \43984 , \43792 );
not \U$44008 ( \43985 , \43984 );
buf \U$44009 ( \43986 , \43985 );
buf \U$44010 ( \43987 , \43986 );
not \U$44011 ( \43988 , \43987 );
buf \U$44012 ( \43989 , \43780 );
not \U$44013 ( \43990 , \43989 );
or \U$44014 ( \43991 , \43988 , \43990 );
buf \U$44015 ( \43992 , RIc0d8140_24);
buf \U$44016 ( \43993 , RIc0db188_127);
xnor \U$44017 ( \43994 , \43992 , \43993 );
buf \U$44018 ( \43995 , \43994 );
buf \U$44019 ( \43996 , \43995 );
buf \U$44020 ( \43997 , \12647 );
or \U$44021 ( \43998 , \43996 , \43997 );
buf \U$44022 ( \43999 , \43998 );
buf \U$44023 ( \44000 , \43999 );
nand \U$44024 ( \44001 , \43991 , \44000 );
buf \U$44025 ( \44002 , \44001 );
xor \U$44026 ( \44003 , \43983 , \44002 );
buf \U$44027 ( \44004 , RIc0d8b18_45);
buf \U$44028 ( \44005 , RIc0da828_107);
xor \U$44029 ( \44006 , \44004 , \44005 );
buf \U$44030 ( \44007 , \44006 );
buf \U$44031 ( \44008 , \44007 );
not \U$44032 ( \44009 , \44008 );
buf \U$44033 ( \44010 , \20741 );
not \U$44034 ( \44011 , \44010 );
or \U$44035 ( \44012 , \44009 , \44011 );
buf \U$44036 ( \44013 , \16071 );
buf \U$44037 ( \44014 , RIc0d8aa0_44);
buf \U$44038 ( \44015 , RIc0da828_107);
xor \U$44039 ( \44016 , \44014 , \44015 );
buf \U$44040 ( \44017 , \44016 );
buf \U$44041 ( \44018 , \44017 );
nand \U$44042 ( \44019 , \44013 , \44018 );
buf \U$44043 ( \44020 , \44019 );
buf \U$44044 ( \44021 , \44020 );
nand \U$44045 ( \44022 , \44012 , \44021 );
buf \U$44046 ( \44023 , \44022 );
xor \U$44047 ( \44024 , \44003 , \44023 );
buf \U$44048 ( \44025 , \44024 );
not \U$44049 ( \44026 , \44025 );
not \U$44050 ( \44027 , \4483 );
buf \U$44051 ( \44028 , RIc0d8cf8_49);
buf \U$44052 ( \44029 , RIc0da648_103);
xnor \U$44053 ( \44030 , \44028 , \44029 );
buf \U$44054 ( \44031 , \44030 );
not \U$44055 ( \44032 , \44031 );
and \U$44056 ( \44033 , \44027 , \44032 );
xor \U$44057 ( \44034 , RIc0da648_103, RIc0d8c80_48);
and \U$44058 ( \44035 , \20243 , \44034 );
nor \U$44059 ( \44036 , \44033 , \44035 );
buf \U$44060 ( \44037 , \44036 );
not \U$44061 ( \44038 , \44037 );
buf \U$44062 ( \44039 , \44038 );
buf \U$44063 ( \44040 , \44039 );
not \U$44064 ( \44041 , \44040 );
xnor \U$44065 ( \44042 , RIc0dacd8_117, RIc0d8668_35);
buf \U$44066 ( \44043 , \44042 );
not \U$44067 ( \44044 , \44043 );
buf \U$44068 ( \44045 , \44044 );
buf \U$44069 ( \44046 , \44045 );
not \U$44070 ( \44047 , \44046 );
buf \U$44071 ( \44048 , \12929 );
not \U$44072 ( \44049 , \44048 );
or \U$44073 ( \44050 , \44047 , \44049 );
buf \U$44074 ( \44051 , \22356 );
xor \U$44075 ( \44052 , RIc0dacd8_117, RIc0d85f0_34);
buf \U$44076 ( \44053 , \44052 );
nand \U$44077 ( \44054 , \44051 , \44053 );
buf \U$44078 ( \44055 , \44054 );
buf \U$44079 ( \44056 , \44055 );
nand \U$44080 ( \44057 , \44050 , \44056 );
buf \U$44081 ( \44058 , \44057 );
buf \U$44082 ( \44059 , \44058 );
not \U$44083 ( \44060 , \44059 );
buf \U$44084 ( \44061 , \44060 );
buf \U$44085 ( \44062 , \44061 );
not \U$44086 ( \44063 , \44062 );
or \U$44087 ( \44064 , \44041 , \44063 );
buf \U$44088 ( \44065 , \44058 );
buf \U$44089 ( \44066 , \44036 );
nand \U$44090 ( \44067 , \44065 , \44066 );
buf \U$44091 ( \44068 , \44067 );
buf \U$44092 ( \44069 , \44068 );
nand \U$44093 ( \44070 , \44064 , \44069 );
buf \U$44094 ( \44071 , \44070 );
buf \U$44095 ( \44072 , \44071 );
buf \U$44096 ( \44073 , RIc0d8938_41);
buf \U$44097 ( \44074 , RIc0daa08_111);
xor \U$44098 ( \44075 , \44073 , \44074 );
buf \U$44099 ( \44076 , \44075 );
buf \U$44100 ( \44077 , \44076 );
not \U$44101 ( \44078 , \44077 );
buf \U$44102 ( \44079 , \18306 );
not \U$44103 ( \44080 , \44079 );
or \U$44104 ( \44081 , \44078 , \44080 );
buf \U$44105 ( \44082 , \14353 );
xor \U$44106 ( \44083 , RIc0daa08_111, RIc0d88c0_40);
buf \U$44107 ( \44084 , \44083 );
nand \U$44108 ( \44085 , \44082 , \44084 );
buf \U$44109 ( \44086 , \44085 );
buf \U$44110 ( \44087 , \44086 );
nand \U$44111 ( \44088 , \44081 , \44087 );
buf \U$44112 ( \44089 , \44088 );
buf \U$44113 ( \44090 , \44089 );
xnor \U$44114 ( \44091 , \44072 , \44090 );
buf \U$44115 ( \44092 , \44091 );
buf \U$44116 ( \44093 , \44092 );
not \U$44117 ( \44094 , \44093 );
buf \U$44118 ( \44095 , \44094 );
buf \U$44119 ( \44096 , \44095 );
not \U$44120 ( \44097 , \44096 );
or \U$44121 ( \44098 , \44026 , \44097 );
buf \U$44122 ( \44099 , \44024 );
not \U$44123 ( \44100 , \44099 );
buf \U$44124 ( \44101 , \44100 );
buf \U$44125 ( \44102 , \44101 );
not \U$44126 ( \44103 , \44102 );
buf \U$44127 ( \44104 , \44092 );
not \U$44128 ( \44105 , \44104 );
or \U$44129 ( \44106 , \44103 , \44105 );
buf \U$44130 ( \44107 , RIc0daeb8_121);
buf \U$44131 ( \44108 , RIc0d8488_31);
xor \U$44132 ( \44109 , \44107 , \44108 );
buf \U$44133 ( \44110 , \44109 );
buf \U$44134 ( \44111 , \44110 );
not \U$44135 ( \44112 , \44111 );
buf \U$44136 ( \44113 , \13310 );
not \U$44137 ( \44114 , \44113 );
or \U$44138 ( \44115 , \44112 , \44114 );
buf \U$44139 ( \44116 , \13314 );
buf \U$44140 ( \44117 , RIc0d8410_30);
buf \U$44141 ( \44118 , RIc0daeb8_121);
xor \U$44142 ( \44119 , \44117 , \44118 );
buf \U$44143 ( \44120 , \44119 );
buf \U$44144 ( \44121 , \44120 );
nand \U$44145 ( \44122 , \44116 , \44121 );
buf \U$44146 ( \44123 , \44122 );
buf \U$44147 ( \44124 , \44123 );
nand \U$44148 ( \44125 , \44115 , \44124 );
buf \U$44149 ( \44126 , \44125 );
buf \U$44150 ( \44127 , RIc0da378_97);
buf \U$44151 ( \44128 , RIc0d8fc8_55);
xor \U$44152 ( \44129 , \44127 , \44128 );
buf \U$44153 ( \44130 , \44129 );
buf \U$44154 ( \44131 , \44130 );
not \U$44155 ( \44132 , \44131 );
buf \U$44156 ( \44133 , \16358 );
not \U$44157 ( \44134 , \44133 );
or \U$44158 ( \44135 , \44132 , \44134 );
buf \U$44159 ( \44136 , \2070 );
buf \U$44160 ( \44137 , RIc0da378_97);
buf \U$44161 ( \44138 , RIc0d8f50_54);
xor \U$44162 ( \44139 , \44137 , \44138 );
buf \U$44163 ( \44140 , \44139 );
buf \U$44164 ( \44141 , \44140 );
nand \U$44165 ( \44142 , \44136 , \44141 );
buf \U$44166 ( \44143 , \44142 );
buf \U$44167 ( \44144 , \44143 );
nand \U$44168 ( \44145 , \44135 , \44144 );
buf \U$44169 ( \44146 , \44145 );
xor \U$44170 ( \44147 , \44126 , \44146 );
buf \U$44171 ( \44148 , RIc0d91a8_59);
buf \U$44172 ( \44149 , RIc0da198_93);
xor \U$44173 ( \44150 , \44148 , \44149 );
buf \U$44174 ( \44151 , \44150 );
buf \U$44175 ( \44152 , \44151 );
not \U$44176 ( \44153 , \44152 );
buf \U$44177 ( \44154 , \1901 );
not \U$44178 ( \44155 , \44154 );
or \U$44179 ( \44156 , \44153 , \44155 );
buf \U$44180 ( \44157 , \4008 );
xor \U$44181 ( \44158 , RIc0da198_93, RIc0d9130_58);
buf \U$44182 ( \44159 , \44158 );
nand \U$44183 ( \44160 , \44157 , \44159 );
buf \U$44184 ( \44161 , \44160 );
buf \U$44185 ( \44162 , \44161 );
nand \U$44186 ( \44163 , \44156 , \44162 );
buf \U$44187 ( \44164 , \44163 );
xor \U$44188 ( \44165 , \44147 , \44164 );
buf \U$44189 ( \44166 , \44165 );
nand \U$44190 ( \44167 , \44106 , \44166 );
buf \U$44191 ( \44168 , \44167 );
buf \U$44192 ( \44169 , \44168 );
nand \U$44193 ( \44170 , \44098 , \44169 );
buf \U$44194 ( \44171 , \44170 );
xor \U$44195 ( \44172 , \43967 , \44171 );
buf \U$44196 ( \44173 , RIc0da738_105);
buf \U$44197 ( \44174 , RIc0d8c80_48);
xor \U$44198 ( \44175 , \44173 , \44174 );
buf \U$44199 ( \44176 , \44175 );
buf \U$44200 ( \44177 , \44176 );
not \U$44201 ( \44178 , \44177 );
buf \U$44202 ( \44179 , \15644 );
not \U$44203 ( \44180 , \44179 );
or \U$44204 ( \44181 , \44178 , \44180 );
buf \U$44205 ( \44182 , \12744 );
buf \U$44206 ( \44183 , RIc0d8c08_47);
buf \U$44207 ( \44184 , RIc0da738_105);
xor \U$44208 ( \44185 , \44183 , \44184 );
buf \U$44209 ( \44186 , \44185 );
buf \U$44210 ( \44187 , \44186 );
nand \U$44211 ( \44188 , \44182 , \44187 );
buf \U$44212 ( \44189 , \44188 );
buf \U$44213 ( \44190 , \44189 );
nand \U$44214 ( \44191 , \44181 , \44190 );
buf \U$44215 ( \44192 , \44191 );
buf \U$44216 ( \44193 , \44192 );
not \U$44217 ( \44194 , \44193 );
buf \U$44218 ( \44195 , RIc0d8aa0_44);
buf \U$44219 ( \44196 , RIc0da918_109);
xor \U$44220 ( \44197 , \44195 , \44196 );
buf \U$44221 ( \44198 , \44197 );
buf \U$44222 ( \44199 , \44198 );
not \U$44223 ( \44200 , \44199 );
buf \U$44224 ( \44201 , \27660 );
not \U$44225 ( \44202 , \44201 );
or \U$44226 ( \44203 , \44200 , \44202 );
buf \U$44227 ( \44204 , \43911 );
not \U$44228 ( \44205 , \44204 );
buf \U$44229 ( \44206 , \20211 );
nand \U$44230 ( \44207 , \44205 , \44206 );
buf \U$44231 ( \44208 , \44207 );
buf \U$44232 ( \44209 , \44208 );
nand \U$44233 ( \44210 , \44203 , \44209 );
buf \U$44234 ( \44211 , \44210 );
buf \U$44235 ( \44212 , \44211 );
not \U$44236 ( \44213 , \44212 );
or \U$44237 ( \44214 , \44194 , \44213 );
buf \U$44238 ( \44215 , \44211 );
buf \U$44239 ( \44216 , \44192 );
or \U$44240 ( \44217 , \44215 , \44216 );
xor \U$44241 ( \44218 , RIc0dadc8_119, RIc0d85f0_34);
buf \U$44242 ( \44219 , \44218 );
not \U$44243 ( \44220 , \44219 );
buf \U$44244 ( \44221 , \13949 );
not \U$44245 ( \44222 , \44221 );
or \U$44246 ( \44223 , \44220 , \44222 );
buf \U$44247 ( \44224 , \13953 );
buf \U$44248 ( \44225 , \43884 );
nand \U$44249 ( \44226 , \44224 , \44225 );
buf \U$44250 ( \44227 , \44226 );
buf \U$44251 ( \44228 , \44227 );
nand \U$44252 ( \44229 , \44223 , \44228 );
buf \U$44253 ( \44230 , \44229 );
buf \U$44254 ( \44231 , \44230 );
nand \U$44255 ( \44232 , \44217 , \44231 );
buf \U$44256 ( \44233 , \44232 );
buf \U$44257 ( \44234 , \44233 );
nand \U$44258 ( \44235 , \44214 , \44234 );
buf \U$44259 ( \44236 , \44235 );
buf \U$44260 ( \44237 , \44236 );
not \U$44261 ( \44238 , \44237 );
buf \U$44262 ( \44239 , RIc0d89b0_42);
buf \U$44263 ( \44240 , RIc0daa08_111);
xor \U$44264 ( \44241 , \44239 , \44240 );
buf \U$44265 ( \44242 , \44241 );
buf \U$44266 ( \44243 , \44242 );
not \U$44267 ( \44244 , \44243 );
buf \U$44268 ( \44245 , \12529 );
not \U$44269 ( \44246 , \44245 );
or \U$44270 ( \44247 , \44244 , \44246 );
buf \U$44271 ( \44248 , \14353 );
buf \U$44272 ( \44249 , \44076 );
nand \U$44273 ( \44250 , \44248 , \44249 );
buf \U$44274 ( \44251 , \44250 );
buf \U$44275 ( \44252 , \44251 );
nand \U$44276 ( \44253 , \44247 , \44252 );
buf \U$44277 ( \44254 , \44253 );
buf \U$44278 ( \44255 , \44254 );
not \U$44279 ( \44256 , \44255 );
buf \U$44280 ( \44257 , \25355 );
not \U$44281 ( \44258 , \44257 );
buf \U$44282 ( \44259 , \44258 );
buf \U$44283 ( \44260 , \44259 );
buf \U$44284 ( \44261 , RIc0d88c0_40);
buf \U$44285 ( \44262 , RIc0daaf8_113);
xnor \U$44286 ( \44263 , \44261 , \44262 );
buf \U$44287 ( \44264 , \44263 );
buf \U$44288 ( \44265 , \44264 );
or \U$44289 ( \44266 , \44260 , \44265 );
buf \U$44290 ( \44267 , \14402 );
buf \U$44291 ( \44268 , RIc0d8848_39);
buf \U$44292 ( \44269 , RIc0daaf8_113);
xor \U$44293 ( \44270 , \44268 , \44269 );
buf \U$44294 ( \44271 , \44270 );
buf \U$44295 ( \44272 , \44271 );
not \U$44296 ( \44273 , \44272 );
buf \U$44297 ( \44274 , \44273 );
buf \U$44298 ( \44275 , \44274 );
or \U$44299 ( \44276 , \44267 , \44275 );
nand \U$44300 ( \44277 , \44266 , \44276 );
buf \U$44301 ( \44278 , \44277 );
buf \U$44302 ( \44279 , \44278 );
not \U$44303 ( \44280 , \44279 );
or \U$44304 ( \44281 , \44256 , \44280 );
buf \U$44305 ( \44282 , \44278 );
buf \U$44306 ( \44283 , \44254 );
or \U$44307 ( \44284 , \44282 , \44283 );
buf \U$44308 ( \44285 , \14982 );
not \U$44309 ( \44286 , \44285 );
buf \U$44310 ( \44287 , RIc0d8410_30);
buf \U$44311 ( \44288 , RIc0dafa8_123);
xor \U$44312 ( \44289 , \44287 , \44288 );
buf \U$44313 ( \44290 , \44289 );
buf \U$44314 ( \44291 , \44290 );
not \U$44315 ( \44292 , \44291 );
or \U$44316 ( \44293 , \44286 , \44292 );
buf \U$44317 ( \44294 , \16695 );
buf \U$44318 ( \44295 , RIc0d8398_29);
buf \U$44319 ( \44296 , RIc0dafa8_123);
xnor \U$44320 ( \44297 , \44295 , \44296 );
buf \U$44321 ( \44298 , \44297 );
buf \U$44322 ( \44299 , \44298 );
or \U$44323 ( \44300 , \44294 , \44299 );
nand \U$44324 ( \44301 , \44293 , \44300 );
buf \U$44325 ( \44302 , \44301 );
buf \U$44326 ( \44303 , \44302 );
nand \U$44327 ( \44304 , \44284 , \44303 );
buf \U$44328 ( \44305 , \44304 );
buf \U$44329 ( \44306 , \44305 );
nand \U$44330 ( \44307 , \44281 , \44306 );
buf \U$44331 ( \44308 , \44307 );
buf \U$44332 ( \44309 , \44308 );
not \U$44333 ( \44310 , \44309 );
or \U$44334 ( \44311 , \44238 , \44310 );
buf \U$44335 ( \44312 , \44308 );
buf \U$44336 ( \44313 , \44236 );
or \U$44337 ( \44314 , \44312 , \44313 );
xor \U$44338 ( \44315 , RIc0daeb8_121, RIc0d8500_32);
buf \U$44339 ( \44316 , \44315 );
not \U$44340 ( \44317 , \44316 );
buf \U$44341 ( \44318 , \19487 );
not \U$44342 ( \44319 , \44318 );
or \U$44343 ( \44320 , \44317 , \44319 );
buf \U$44344 ( \44321 , \13314 );
buf \U$44345 ( \44322 , \44110 );
nand \U$44346 ( \44323 , \44321 , \44322 );
buf \U$44347 ( \44324 , \44323 );
buf \U$44348 ( \44325 , \44324 );
nand \U$44349 ( \44326 , \44320 , \44325 );
buf \U$44350 ( \44327 , \44326 );
buf \U$44351 ( \44328 , \44327 );
buf \U$44352 ( \44329 , RIc0d9220_60);
buf \U$44353 ( \44330 , RIc0da198_93);
xor \U$44354 ( \44331 , \44329 , \44330 );
buf \U$44355 ( \44332 , \44331 );
buf \U$44356 ( \44333 , \44332 );
not \U$44357 ( \44334 , \44333 );
buf \U$44358 ( \44335 , \889 );
not \U$44359 ( \44336 , \44335 );
or \U$44360 ( \44337 , \44334 , \44336 );
buf \U$44361 ( \44338 , \4008 );
buf \U$44362 ( \44339 , \44151 );
nand \U$44363 ( \44340 , \44338 , \44339 );
buf \U$44364 ( \44341 , \44340 );
buf \U$44365 ( \44342 , \44341 );
nand \U$44366 ( \44343 , \44337 , \44342 );
buf \U$44367 ( \44344 , \44343 );
buf \U$44368 ( \44345 , \44344 );
xor \U$44369 ( \44346 , \44328 , \44345 );
buf \U$44370 ( \44347 , RIc0d8b90_46);
buf \U$44371 ( \44348 , RIc0da828_107);
xor \U$44372 ( \44349 , \44347 , \44348 );
buf \U$44373 ( \44350 , \44349 );
buf \U$44374 ( \44351 , \44350 );
not \U$44375 ( \44352 , \44351 );
buf \U$44376 ( \44353 , \37534 );
not \U$44377 ( \44354 , \44353 );
or \U$44378 ( \44355 , \44352 , \44354 );
buf \U$44379 ( \44356 , \12342 );
buf \U$44380 ( \44357 , \44007 );
nand \U$44381 ( \44358 , \44356 , \44357 );
buf \U$44382 ( \44359 , \44358 );
buf \U$44383 ( \44360 , \44359 );
nand \U$44384 ( \44361 , \44355 , \44360 );
buf \U$44385 ( \44362 , \44361 );
buf \U$44386 ( \44363 , \44362 );
and \U$44387 ( \44364 , \44346 , \44363 );
and \U$44388 ( \44365 , \44328 , \44345 );
or \U$44389 ( \44366 , \44364 , \44365 );
buf \U$44390 ( \44367 , \44366 );
buf \U$44391 ( \44368 , \44367 );
nand \U$44392 ( \44369 , \44314 , \44368 );
buf \U$44393 ( \44370 , \44369 );
buf \U$44394 ( \44371 , \44370 );
nand \U$44395 ( \44372 , \44311 , \44371 );
buf \U$44396 ( \44373 , \44372 );
xor \U$44397 ( \44374 , \44172 , \44373 );
buf \U$44398 ( \44375 , \44374 );
buf \U$44399 ( \44376 , RIc0d82a8_27);
buf \U$44400 ( \44377 , RIc0db098_125);
xor \U$44401 ( \44378 , \44376 , \44377 );
buf \U$44402 ( \44379 , \44378 );
buf \U$44403 ( \44380 , \44379 );
not \U$44404 ( \44381 , \44380 );
buf \U$44407 ( \44382 , \15789 );
buf \U$44408 ( \44383 , \44382 );
not \U$44409 ( \44384 , \44383 );
or \U$44410 ( \44385 , \44381 , \44384 );
buf \U$44411 ( \44386 , \13465 );
buf \U$44412 ( \44387 , RIc0d8230_26);
buf \U$44413 ( \44388 , RIc0db098_125);
xor \U$44414 ( \44389 , \44387 , \44388 );
buf \U$44415 ( \44390 , \44389 );
buf \U$44416 ( \44391 , \44390 );
nand \U$44417 ( \44392 , \44386 , \44391 );
buf \U$44418 ( \44393 , \44392 );
buf \U$44419 ( \44394 , \44393 );
nand \U$44420 ( \44395 , \44385 , \44394 );
buf \U$44421 ( \44396 , \44395 );
buf \U$44422 ( \44397 , RIc0d8de8_51);
buf \U$44423 ( \44398 , RIc0da558_101);
xor \U$44424 ( \44399 , \44397 , \44398 );
buf \U$44425 ( \44400 , \44399 );
buf \U$44426 ( \44401 , \44400 );
not \U$44427 ( \44402 , \44401 );
buf \U$44428 ( \44403 , \33258 );
not \U$44429 ( \44404 , \44403 );
or \U$44430 ( \44405 , \44402 , \44404 );
buf \U$44431 ( \44406 , \16676 );
xor \U$44432 ( \44407 , RIc0da558_101, RIc0d8d70_50);
buf \U$44433 ( \44408 , \44407 );
nand \U$44434 ( \44409 , \44406 , \44408 );
buf \U$44435 ( \44410 , \44409 );
buf \U$44436 ( \44411 , \44410 );
nand \U$44437 ( \44412 , \44405 , \44411 );
buf \U$44438 ( \44413 , \44412 );
xor \U$44439 ( \44414 , \44396 , \44413 );
buf \U$44440 ( \44415 , \44186 );
not \U$44441 ( \44416 , \44415 );
buf \U$44442 ( \44417 , \12736 );
not \U$44443 ( \44418 , \44417 );
or \U$44444 ( \44419 , \44416 , \44418 );
buf \U$44445 ( \44420 , \12744 );
buf \U$44446 ( \44421 , RIc0d8b90_46);
buf \U$44447 ( \44422 , RIc0da738_105);
xor \U$44448 ( \44423 , \44421 , \44422 );
buf \U$44449 ( \44424 , \44423 );
buf \U$44450 ( \44425 , \44424 );
nand \U$44451 ( \44426 , \44420 , \44425 );
buf \U$44452 ( \44427 , \44426 );
buf \U$44453 ( \44428 , \44427 );
nand \U$44454 ( \44429 , \44419 , \44428 );
buf \U$44455 ( \44430 , \44429 );
xor \U$44456 ( \44431 , \44414 , \44430 );
buf \U$44457 ( \44432 , \44431 );
not \U$44458 ( \44433 , \44432 );
buf \U$44459 ( \44434 , RIc0d8ed8_53);
buf \U$44460 ( \44435 , RIc0da468_99);
xor \U$44461 ( \44436 , \44434 , \44435 );
buf \U$44462 ( \44437 , \44436 );
buf \U$44463 ( \44438 , \44437 );
not \U$44464 ( \44439 , \44438 );
buf \U$44465 ( \44440 , \19695 );
not \U$44466 ( \44441 , \44440 );
or \U$44467 ( \44442 , \44439 , \44441 );
buf \U$44468 ( \44443 , \2476 );
xor \U$44469 ( \44444 , RIc0da468_99, RIc0d8e60_52);
buf \U$44470 ( \44445 , \44444 );
nand \U$44471 ( \44446 , \44443 , \44445 );
buf \U$44472 ( \44447 , \44446 );
buf \U$44473 ( \44448 , \44447 );
nand \U$44474 ( \44449 , \44442 , \44448 );
buf \U$44475 ( \44450 , \44449 );
buf \U$44476 ( \44451 , \44450 );
buf \U$44477 ( \44452 , \44271 );
not \U$44478 ( \44453 , \44452 );
buf \U$44479 ( \44454 , \26484 );
not \U$44480 ( \44455 , \44454 );
or \U$44481 ( \44456 , \44453 , \44455 );
buf \U$44482 ( \44457 , \12410 );
buf \U$44483 ( \44458 , RIc0d87d0_38);
buf \U$44484 ( \44459 , RIc0daaf8_113);
xor \U$44485 ( \44460 , \44458 , \44459 );
buf \U$44486 ( \44461 , \44460 );
buf \U$44487 ( \44462 , \44461 );
nand \U$44488 ( \44463 , \44457 , \44462 );
buf \U$44489 ( \44464 , \44463 );
buf \U$44490 ( \44465 , \44464 );
nand \U$44491 ( \44466 , \44456 , \44465 );
buf \U$44492 ( \44467 , \44466 );
buf \U$44493 ( \44468 , \44467 );
xor \U$44494 ( \44469 , \44451 , \44468 );
buf \U$44495 ( \44470 , \16688 );
buf \U$44496 ( \44471 , \44298 );
or \U$44497 ( \44472 , \44470 , \44471 );
buf \U$44498 ( \44473 , \16695 );
buf \U$44499 ( \44474 , RIc0dafa8_123);
buf \U$44500 ( \44475 , RIc0d8320_28);
xnor \U$44501 ( \44476 , \44474 , \44475 );
buf \U$44502 ( \44477 , \44476 );
buf \U$44503 ( \44478 , \44477 );
or \U$44504 ( \44479 , \44473 , \44478 );
nand \U$44505 ( \44480 , \44472 , \44479 );
buf \U$44506 ( \44481 , \44480 );
buf \U$44507 ( \44482 , \44481 );
xor \U$44508 ( \44483 , \44469 , \44482 );
buf \U$44509 ( \44484 , \44483 );
buf \U$44510 ( \44485 , \44484 );
not \U$44511 ( \44486 , \44485 );
or \U$44512 ( \44487 , \44433 , \44486 );
buf \U$44513 ( \44488 , \44484 );
buf \U$44514 ( \44489 , \44431 );
or \U$44515 ( \44490 , \44488 , \44489 );
buf \U$44516 ( \44491 , RIc0d9400_64);
buf \U$44517 ( \44492 , RIc0d9fb8_89);
xor \U$44518 ( \44493 , \44491 , \44492 );
buf \U$44519 ( \44494 , \44493 );
buf \U$44520 ( \44495 , \44494 );
not \U$44521 ( \44496 , \44495 );
buf \U$44522 ( \44497 , \3384 );
not \U$44523 ( \44498 , \44497 );
or \U$44524 ( \44499 , \44496 , \44498 );
buf \U$44525 ( \44500 , \442 );
buf \U$44526 ( \44501 , \43943 );
nand \U$44527 ( \44502 , \44500 , \44501 );
buf \U$44528 ( \44503 , \44502 );
buf \U$44529 ( \44504 , \44503 );
nand \U$44530 ( \44505 , \44499 , \44504 );
buf \U$44531 ( \44506 , \44505 );
buf \U$44532 ( \44507 , \44506 );
buf \U$44533 ( \44508 , RIc0d9400_64);
buf \U$44534 ( \44509 , RIc0da030_90);
or \U$44535 ( \44510 , \44508 , \44509 );
buf \U$44536 ( \44511 , RIc0da0a8_91);
nand \U$44537 ( \44512 , \44510 , \44511 );
buf \U$44538 ( \44513 , \44512 );
buf \U$44539 ( \44514 , \44513 );
buf \U$44540 ( \44515 , RIc0d9400_64);
buf \U$44541 ( \44516 , RIc0da030_90);
nand \U$44542 ( \44517 , \44515 , \44516 );
buf \U$44543 ( \44518 , \44517 );
buf \U$44544 ( \44519 , \44518 );
buf \U$44545 ( \44520 , RIc0d9fb8_89);
and \U$44546 ( \44521 , \44514 , \44519 , \44520 );
buf \U$44547 ( \44522 , \44521 );
buf \U$44548 ( \44523 , \44522 );
buf \U$44549 ( \44524 , RIc0d9310_62);
buf \U$44550 ( \44525 , RIc0da0a8_91);
xor \U$44551 ( \44526 , \44524 , \44525 );
buf \U$44552 ( \44527 , \44526 );
buf \U$44553 ( \44528 , \44527 );
not \U$44554 ( \44529 , \44528 );
buf \U$44555 ( \44530 , \2726 );
not \U$44556 ( \44531 , \44530 );
or \U$44557 ( \44532 , \44529 , \44531 );
buf \U$44558 ( \44533 , \43867 );
not \U$44559 ( \44534 , \44533 );
buf \U$44560 ( \44535 , \714 );
nand \U$44561 ( \44536 , \44534 , \44535 );
buf \U$44562 ( \44537 , \44536 );
buf \U$44563 ( \44538 , \44537 );
nand \U$44564 ( \44539 , \44532 , \44538 );
buf \U$44565 ( \44540 , \44539 );
buf \U$44566 ( \44541 , \44540 );
xor \U$44567 ( \44542 , \44523 , \44541 );
buf \U$44568 ( \44543 , \44542 );
buf \U$44569 ( \44544 , \44543 );
xor \U$44570 ( \44545 , \44507 , \44544 );
buf \U$44571 ( \44546 , RIc0db098_125);
buf \U$44572 ( \44547 , RIc0d8398_29);
xor \U$44573 ( \44548 , \44546 , \44547 );
buf \U$44574 ( \44549 , \44548 );
buf \U$44575 ( \44550 , \44549 );
not \U$44576 ( \44551 , \44550 );
buf \U$44577 ( \44552 , \13461 );
not \U$44578 ( \44553 , \44552 );
or \U$44579 ( \44554 , \44551 , \44553 );
buf \U$44580 ( \44555 , RIc0db098_125);
buf \U$44581 ( \44556 , RIc0d8320_28);
xnor \U$44582 ( \44557 , \44555 , \44556 );
buf \U$44583 ( \44558 , \44557 );
buf \U$44584 ( \44559 , \44558 );
not \U$44585 ( \44560 , \44559 );
buf \U$44586 ( \44561 , \13465 );
nand \U$44587 ( \44562 , \44560 , \44561 );
buf \U$44588 ( \44563 , \44562 );
buf \U$44589 ( \44564 , \44563 );
nand \U$44590 ( \44565 , \44554 , \44564 );
buf \U$44591 ( \44566 , \44565 );
buf \U$44592 ( \44567 , \44566 );
not \U$44593 ( \44568 , \44567 );
buf \U$44594 ( \44569 , RIc0da558_101);
buf \U$44595 ( \44570 , RIc0d8ed8_53);
xor \U$44596 ( \44571 , \44569 , \44570 );
buf \U$44597 ( \44572 , \44571 );
buf \U$44598 ( \44573 , \44572 );
not \U$44599 ( \44574 , \44573 );
buf \U$44600 ( \44575 , \22631 );
not \U$44601 ( \44576 , \44575 );
or \U$44602 ( \44577 , \44574 , \44576 );
buf \U$44603 ( \44578 , \15550 );
buf \U$44604 ( \44579 , RIc0d8e60_52);
buf \U$44605 ( \44580 , RIc0da558_101);
xor \U$44606 ( \44581 , \44579 , \44580 );
buf \U$44607 ( \44582 , \44581 );
buf \U$44608 ( \44583 , \44582 );
nand \U$44609 ( \44584 , \44578 , \44583 );
buf \U$44610 ( \44585 , \44584 );
buf \U$44611 ( \44586 , \44585 );
nand \U$44612 ( \44587 , \44577 , \44586 );
buf \U$44613 ( \44588 , \44587 );
buf \U$44614 ( \44589 , \44588 );
not \U$44615 ( \44590 , \44589 );
or \U$44616 ( \44591 , \44568 , \44590 );
buf \U$44617 ( \44592 , \44588 );
buf \U$44618 ( \44593 , \44566 );
or \U$44619 ( \44594 , \44592 , \44593 );
buf \U$44620 ( \44595 , RIc0d8de8_51);
buf \U$44621 ( \44596 , RIc0da648_103);
xor \U$44622 ( \44597 , \44595 , \44596 );
buf \U$44623 ( \44598 , \44597 );
buf \U$44624 ( \44599 , \44598 );
not \U$44625 ( \44600 , \44599 );
buf \U$44626 ( \44601 , \13706 );
not \U$44627 ( \44602 , \44601 );
or \U$44628 ( \44603 , \44600 , \44602 );
buf \U$44629 ( \44604 , \13048 );
buf \U$44630 ( \44605 , RIc0d8d70_50);
buf \U$44631 ( \44606 , RIc0da648_103);
xor \U$44632 ( \44607 , \44605 , \44606 );
buf \U$44633 ( \44608 , \44607 );
buf \U$44634 ( \44609 , \44608 );
nand \U$44635 ( \44610 , \44604 , \44609 );
buf \U$44636 ( \44611 , \44610 );
buf \U$44637 ( \44612 , \44611 );
nand \U$44638 ( \44613 , \44603 , \44612 );
buf \U$44639 ( \44614 , \44613 );
buf \U$44640 ( \44615 , \44614 );
nand \U$44641 ( \44616 , \44594 , \44615 );
buf \U$44642 ( \44617 , \44616 );
buf \U$44643 ( \44618 , \44617 );
nand \U$44644 ( \44619 , \44591 , \44618 );
buf \U$44645 ( \44620 , \44619 );
buf \U$44646 ( \44621 , \44620 );
and \U$44647 ( \44622 , \44545 , \44621 );
and \U$44648 ( \44623 , \44507 , \44544 );
or \U$44649 ( \44624 , \44622 , \44623 );
buf \U$44650 ( \44625 , \44624 );
buf \U$44651 ( \44626 , \44625 );
nand \U$44652 ( \44627 , \44490 , \44626 );
buf \U$44653 ( \44628 , \44627 );
buf \U$44654 ( \44629 , \44628 );
nand \U$44655 ( \44630 , \44487 , \44629 );
buf \U$44656 ( \44631 , \44630 );
buf \U$44657 ( \44632 , \44631 );
xor \U$44658 ( \44633 , \43847 , \43861 );
and \U$44659 ( \44634 , \44633 , \43879 );
and \U$44660 ( \44635 , \43847 , \43861 );
or \U$44661 ( \44636 , \44634 , \44635 );
buf \U$44662 ( \44637 , \44636 );
buf \U$44663 ( \44638 , \44637 );
buf \U$44664 ( \44639 , \15608 );
not \U$44665 ( \44640 , \44639 );
buf \U$44666 ( \44641 , \44640 );
buf \U$44667 ( \44642 , \43995 );
or \U$44668 ( \44643 , \44641 , \44642 );
buf \U$44669 ( \44644 , \12647 );
buf \U$44670 ( \44645 , RIc0d80c8_23);
buf \U$44671 ( \44646 , RIc0db188_127);
xnor \U$44672 ( \44647 , \44645 , \44646 );
buf \U$44673 ( \44648 , \44647 );
buf \U$44674 ( \44649 , \44648 );
or \U$44675 ( \44650 , \44644 , \44649 );
nand \U$44676 ( \44651 , \44643 , \44650 );
buf \U$44677 ( \44652 , \44651 );
buf \U$44678 ( \44653 , \44652 );
buf \U$44679 ( \44654 , \44120 );
not \U$44680 ( \44655 , \44654 );
buf \U$44681 ( \44656 , \17089 );
not \U$44682 ( \44657 , \44656 );
or \U$44683 ( \44658 , \44655 , \44657 );
buf \U$44684 ( \44659 , \13314 );
xor \U$44685 ( \44660 , RIc0daeb8_121, RIc0d8398_29);
buf \U$44686 ( \44661 , \44660 );
nand \U$44687 ( \44662 , \44659 , \44661 );
buf \U$44688 ( \44663 , \44662 );
buf \U$44689 ( \44664 , \44663 );
nand \U$44690 ( \44665 , \44658 , \44664 );
buf \U$44691 ( \44666 , \44665 );
buf \U$44692 ( \44667 , \44666 );
xor \U$44693 ( \44668 , \44653 , \44667 );
buf \U$44694 ( \44669 , \333 );
buf \U$44695 ( \44670 , \43977 );
not \U$44696 ( \44671 , \44670 );
buf \U$44697 ( \44672 , \44671 );
buf \U$44698 ( \44673 , \44672 );
or \U$44699 ( \44674 , \44669 , \44673 );
buf \U$44700 ( \44675 , \14704 );
buf \U$44701 ( \44676 , RIc0da288_95);
buf \U$44702 ( \44677 , RIc0d8fc8_55);
xor \U$44703 ( \44678 , \44676 , \44677 );
buf \U$44704 ( \44679 , \44678 );
buf \U$44705 ( \44680 , \44679 );
not \U$44706 ( \44681 , \44680 );
buf \U$44707 ( \44682 , \44681 );
buf \U$44708 ( \44683 , \44682 );
or \U$44709 ( \44684 , \44675 , \44683 );
nand \U$44710 ( \44685 , \44674 , \44684 );
buf \U$44711 ( \44686 , \44685 );
buf \U$44712 ( \44687 , \44686 );
xor \U$44713 ( \44688 , \44668 , \44687 );
buf \U$44714 ( \44689 , \44688 );
buf \U$44715 ( \44690 , \44689 );
xor \U$44716 ( \44691 , \44638 , \44690 );
buf \U$44717 ( \44692 , \44407 );
not \U$44718 ( \44693 , \44692 );
buf \U$44719 ( \44694 , \3535 );
not \U$44720 ( \44695 , \44694 );
or \U$44721 ( \44696 , \44693 , \44695 );
buf \U$44722 ( \44697 , \16676 );
buf \U$44723 ( \44698 , RIc0d8cf8_49);
buf \U$44724 ( \44699 , RIc0da558_101);
xor \U$44725 ( \44700 , \44698 , \44699 );
buf \U$44726 ( \44701 , \44700 );
buf \U$44727 ( \44702 , \44701 );
nand \U$44728 ( \44703 , \44697 , \44702 );
buf \U$44729 ( \44704 , \44703 );
buf \U$44730 ( \44705 , \44704 );
nand \U$44731 ( \44706 , \44696 , \44705 );
buf \U$44732 ( \44707 , \44706 );
buf \U$44733 ( \44708 , \44017 );
not \U$44734 ( \44709 , \44708 );
buf \U$44735 ( \44710 , \17595 );
not \U$44736 ( \44711 , \44710 );
or \U$44737 ( \44712 , \44709 , \44711 );
buf \U$44738 ( \44713 , \12342 );
xor \U$44739 ( \44714 , RIc0da828_107, RIc0d8a28_43);
buf \U$44740 ( \44715 , \44714 );
nand \U$44741 ( \44716 , \44713 , \44715 );
buf \U$44742 ( \44717 , \44716 );
buf \U$44743 ( \44718 , \44717 );
nand \U$44744 ( \44719 , \44712 , \44718 );
buf \U$44745 ( \44720 , \44719 );
buf \U$44746 ( \44721 , \43854 );
not \U$44747 ( \44722 , \44721 );
buf \U$44748 ( \44723 , \14186 );
not \U$44749 ( \44724 , \44723 );
or \U$44750 ( \44725 , \44722 , \44724 );
buf \U$44751 ( \44726 , \14690 );
buf \U$44752 ( \44727 , RIc0d8668_35);
buf \U$44753 ( \44728 , RIc0dabe8_115);
xor \U$44754 ( \44729 , \44727 , \44728 );
buf \U$44755 ( \44730 , \44729 );
buf \U$44756 ( \44731 , \44730 );
nand \U$44757 ( \44732 , \44726 , \44731 );
buf \U$44758 ( \44733 , \44732 );
buf \U$44759 ( \44734 , \44733 );
nand \U$44760 ( \44735 , \44725 , \44734 );
buf \U$44761 ( \44736 , \44735 );
xor \U$44762 ( \44737 , \44720 , \44736 );
xor \U$44763 ( \44738 , \44707 , \44737 );
buf \U$44764 ( \44739 , \44738 );
xor \U$44765 ( \44740 , \44691 , \44739 );
buf \U$44766 ( \44741 , \44740 );
buf \U$44767 ( \44742 , \44741 );
xor \U$44768 ( \44743 , \44632 , \44742 );
buf \U$44769 ( \44744 , \44444 );
not \U$44770 ( \44745 , \44744 );
buf \U$44771 ( \44746 , \25371 );
not \U$44772 ( \44747 , \44746 );
or \U$44773 ( \44748 , \44745 , \44747 );
buf \U$44774 ( \44749 , \14648 );
xor \U$44775 ( \44750 , RIc0da468_99, RIc0d8de8_51);
buf \U$44776 ( \44751 , \44750 );
nand \U$44777 ( \44752 , \44749 , \44751 );
buf \U$44778 ( \44753 , \44752 );
buf \U$44779 ( \44754 , \44753 );
nand \U$44780 ( \44755 , \44748 , \44754 );
buf \U$44781 ( \44756 , \44755 );
buf \U$44782 ( \44757 , \44083 );
not \U$44783 ( \44758 , \44757 );
buf \U$44784 ( \44759 , \12529 );
not \U$44785 ( \44760 , \44759 );
or \U$44786 ( \44761 , \44758 , \44760 );
buf \U$44787 ( \44762 , \15864 );
xor \U$44788 ( \44763 , RIc0daa08_111, RIc0d8848_39);
buf \U$44789 ( \44764 , \44763 );
nand \U$44790 ( \44765 , \44762 , \44764 );
buf \U$44791 ( \44766 , \44765 );
buf \U$44792 ( \44767 , \44766 );
nand \U$44793 ( \44768 , \44761 , \44767 );
buf \U$44794 ( \44769 , \44768 );
xor \U$44795 ( \44770 , \44756 , \44769 );
buf \U$44796 ( \44771 , \44140 );
not \U$44797 ( \44772 , \44771 );
buf \U$44798 ( \44773 , \2066 );
not \U$44799 ( \44774 , \44773 );
or \U$44800 ( \44775 , \44772 , \44774 );
buf \U$44801 ( \44776 , \2070 );
buf \U$44802 ( \44777 , RIc0da378_97);
buf \U$44803 ( \44778 , RIc0d8ed8_53);
xor \U$44804 ( \44779 , \44777 , \44778 );
buf \U$44805 ( \44780 , \44779 );
buf \U$44806 ( \44781 , \44780 );
nand \U$44807 ( \44782 , \44776 , \44781 );
buf \U$44808 ( \44783 , \44782 );
buf \U$44809 ( \44784 , \44783 );
nand \U$44810 ( \44785 , \44775 , \44784 );
buf \U$44811 ( \44786 , \44785 );
xor \U$44812 ( \44787 , \44770 , \44786 );
buf \U$44813 ( \44788 , \44787 );
buf \U$44814 ( \44789 , \43917 );
not \U$44815 ( \44790 , \44789 );
buf \U$44816 ( \44791 , \44790 );
buf \U$44817 ( \44792 , \44791 );
not \U$44818 ( \44793 , \44792 );
buf \U$44819 ( \44794 , \27660 );
not \U$44820 ( \44795 , \44794 );
or \U$44821 ( \44796 , \44793 , \44795 );
buf \U$44822 ( \44797 , \20211 );
buf \U$44823 ( \44798 , RIc0d8938_41);
buf \U$44824 ( \44799 , RIc0da918_109);
xor \U$44825 ( \44800 , \44798 , \44799 );
buf \U$44826 ( \44801 , \44800 );
buf \U$44827 ( \44802 , \44801 );
nand \U$44828 ( \44803 , \44797 , \44802 );
buf \U$44829 ( \44804 , \44803 );
buf \U$44830 ( \44805 , \44804 );
nand \U$44831 ( \44806 , \44796 , \44805 );
buf \U$44832 ( \44807 , \44806 );
buf \U$44833 ( \44808 , \44807 );
buf \U$44834 ( \44809 , \44390 );
not \U$44835 ( \44810 , \44809 );
buf \U$44836 ( \44811 , \17992 );
not \U$44837 ( \44812 , \44811 );
buf \U$44838 ( \44813 , \44812 );
buf \U$44839 ( \44814 , \44813 );
not \U$44840 ( \44815 , \44814 );
or \U$44841 ( \44816 , \44810 , \44815 );
buf \U$44842 ( \44817 , RIc0db098_125);
buf \U$44843 ( \44818 , RIc0d81b8_25);
xnor \U$44844 ( \44819 , \44817 , \44818 );
buf \U$44845 ( \44820 , \44819 );
buf \U$44846 ( \44821 , \44820 );
not \U$44847 ( \44822 , \44821 );
buf \U$44848 ( \44823 , \15793 );
nand \U$44849 ( \44824 , \44822 , \44823 );
buf \U$44850 ( \44825 , \44824 );
buf \U$44851 ( \44826 , \44825 );
nand \U$44852 ( \44827 , \44816 , \44826 );
buf \U$44853 ( \44828 , \44827 );
buf \U$44854 ( \44829 , \44828 );
and \U$44855 ( \44830 , \44808 , \44829 );
not \U$44856 ( \44831 , \44808 );
buf \U$44857 ( \44832 , \44828 );
not \U$44858 ( \44833 , \44832 );
buf \U$44859 ( \44834 , \44833 );
buf \U$44860 ( \44835 , \44834 );
and \U$44861 ( \44836 , \44831 , \44835 );
nor \U$44862 ( \44837 , \44830 , \44836 );
buf \U$44863 ( \44838 , \44837 );
buf \U$44864 ( \44839 , RIc0d9400_64);
buf \U$44865 ( \44840 , RIc0d9f40_88);
or \U$44866 ( \44841 , \44839 , \44840 );
buf \U$44867 ( \44842 , RIc0d9fb8_89);
nand \U$44868 ( \44843 , \44841 , \44842 );
buf \U$44869 ( \44844 , \44843 );
buf \U$44870 ( \44845 , \44844 );
buf \U$44871 ( \44846 , RIc0d9400_64);
buf \U$44872 ( \44847 , RIc0d9f40_88);
nand \U$44873 ( \44848 , \44846 , \44847 );
buf \U$44874 ( \44849 , \44848 );
buf \U$44875 ( \44850 , \44849 );
buf \U$44876 ( \44851 , RIc0d9ec8_87);
and \U$44877 ( \44852 , \44845 , \44850 , \44851 );
buf \U$44878 ( \44853 , \44852 );
buf \U$44879 ( \44854 , \44853 );
buf \U$44880 ( \44855 , \43953 );
not \U$44881 ( \44856 , \44855 );
buf \U$44882 ( \44857 , \2038 );
not \U$44883 ( \44858 , \44857 );
or \U$44884 ( \44859 , \44856 , \44858 );
buf \U$44885 ( \44860 , \442 );
buf \U$44886 ( \44861 , RIc0d9fb8_89);
buf \U$44887 ( \44862 , RIc0d9298_61);
xor \U$44888 ( \44863 , \44861 , \44862 );
buf \U$44889 ( \44864 , \44863 );
buf \U$44890 ( \44865 , \44864 );
nand \U$44891 ( \44866 , \44860 , \44865 );
buf \U$44892 ( \44867 , \44866 );
buf \U$44893 ( \44868 , \44867 );
nand \U$44894 ( \44869 , \44859 , \44868 );
buf \U$44895 ( \44870 , \44869 );
buf \U$44896 ( \44871 , \44870 );
xor \U$44897 ( \44872 , \44854 , \44871 );
buf \U$44898 ( \44873 , \44872 );
xor \U$44899 ( \44874 , \44838 , \44873 );
buf \U$44900 ( \44875 , \44874 );
xor \U$44901 ( \44876 , \44788 , \44875 );
and \U$44902 ( \44877 , \44523 , \44541 );
buf \U$44903 ( \44878 , \44877 );
buf \U$44904 ( \44879 , \44878 );
buf \U$44905 ( \44880 , \22350 );
not \U$44906 ( \44881 , \44880 );
buf \U$44907 ( \44882 , \44881 );
buf \U$44908 ( \44883 , \44882 );
not \U$44909 ( \44884 , \44883 );
buf \U$44910 ( \44885 , RIc0dacd8_117);
buf \U$44911 ( \44886 , RIc0d86e0_36);
xnor \U$44912 ( \44887 , \44885 , \44886 );
buf \U$44913 ( \44888 , \44887 );
buf \U$44914 ( \44889 , \44888 );
not \U$44915 ( \44890 , \44889 );
and \U$44916 ( \44891 , \44884 , \44890 );
buf \U$44917 ( \44892 , \12937 );
not \U$44918 ( \44893 , \44892 );
buf \U$44919 ( \44894 , \44893 );
buf \U$44920 ( \44895 , \44894 );
buf \U$44921 ( \44896 , \44042 );
nor \U$44922 ( \44897 , \44895 , \44896 );
buf \U$44923 ( \44898 , \44897 );
buf \U$44924 ( \44899 , \44898 );
nor \U$44925 ( \44900 , \44891 , \44899 );
buf \U$44926 ( \44901 , \44900 );
buf \U$44927 ( \44902 , \44901 );
not \U$44928 ( \44903 , \44902 );
not \U$44929 ( \44904 , \2938 );
buf \U$44930 ( \44905 , RIc0d9040_56);
buf \U$44931 ( \44906 , RIc0da378_97);
xnor \U$44932 ( \44907 , \44905 , \44906 );
buf \U$44933 ( \44908 , \44907 );
not \U$44934 ( \44909 , \44908 );
and \U$44935 ( \44910 , \44904 , \44909 );
and \U$44936 ( \44911 , \2070 , \44130 );
nor \U$44937 ( \44912 , \44910 , \44911 );
buf \U$44938 ( \44913 , \44912 );
not \U$44939 ( \44914 , \44913 );
or \U$44940 ( \44915 , \44903 , \44914 );
buf \U$44941 ( \44916 , \44608 );
not \U$44942 ( \44917 , \44916 );
buf \U$44943 ( \44918 , \13706 );
not \U$44944 ( \44919 , \44918 );
or \U$44945 ( \44920 , \44917 , \44919 );
buf \U$44946 ( \44921 , \44031 );
not \U$44947 ( \44922 , \44921 );
buf \U$44948 ( \44923 , \16584 );
nand \U$44949 ( \44924 , \44922 , \44923 );
buf \U$44950 ( \44925 , \44924 );
buf \U$44951 ( \44926 , \44925 );
nand \U$44952 ( \44927 , \44920 , \44926 );
buf \U$44953 ( \44928 , \44927 );
buf \U$44954 ( \44929 , \44928 );
nand \U$44955 ( \44930 , \44915 , \44929 );
buf \U$44956 ( \44931 , \44930 );
buf \U$44957 ( \44932 , \44931 );
buf \U$44958 ( \44933 , \44912 );
not \U$44959 ( \44934 , \44933 );
buf \U$44960 ( \44935 , \44934 );
buf \U$44961 ( \44936 , \44935 );
buf \U$44962 ( \44937 , \44901 );
not \U$44963 ( \44938 , \44937 );
buf \U$44964 ( \44939 , \44938 );
buf \U$44965 ( \44940 , \44939 );
nand \U$44966 ( \44941 , \44936 , \44940 );
buf \U$44967 ( \44942 , \44941 );
buf \U$44968 ( \44943 , \44942 );
nand \U$44969 ( \44944 , \44932 , \44943 );
buf \U$44970 ( \44945 , \44944 );
buf \U$44971 ( \44946 , \44945 );
xor \U$44972 ( \44947 , \44879 , \44946 );
buf \U$44973 ( \44948 , \44582 );
not \U$44974 ( \44949 , \44948 );
buf \U$44975 ( \44950 , \4043 );
not \U$44976 ( \44951 , \44950 );
or \U$44977 ( \44952 , \44949 , \44951 );
buf \U$44978 ( \44953 , \4049 );
buf \U$44979 ( \44954 , \44400 );
nand \U$44980 ( \44955 , \44953 , \44954 );
buf \U$44981 ( \44956 , \44955 );
buf \U$44982 ( \44957 , \44956 );
nand \U$44983 ( \44958 , \44952 , \44957 );
buf \U$44984 ( \44959 , \44958 );
buf \U$44985 ( \44960 , \44959 );
not \U$44986 ( \44961 , \44960 );
buf \U$44987 ( \44962 , RIc0d8f50_54);
buf \U$44988 ( \44963 , RIc0da468_99);
xor \U$44989 ( \44964 , \44962 , \44963 );
buf \U$44990 ( \44965 , \44964 );
buf \U$44991 ( \44966 , \44965 );
not \U$44992 ( \44967 , \44966 );
buf \U$44993 ( \44968 , \2470 );
not \U$44994 ( \44969 , \44968 );
or \U$44995 ( \44970 , \44967 , \44969 );
buf \U$44996 ( \44971 , \2476 );
buf \U$44997 ( \44972 , \44437 );
nand \U$44998 ( \44973 , \44971 , \44972 );
buf \U$44999 ( \44974 , \44973 );
buf \U$45000 ( \44975 , \44974 );
nand \U$45001 ( \44976 , \44970 , \44975 );
buf \U$45002 ( \44977 , \44976 );
buf \U$45003 ( \44978 , \44977 );
not \U$45004 ( \44979 , \44978 );
or \U$45005 ( \44980 , \44961 , \44979 );
buf \U$45006 ( \44981 , \44977 );
buf \U$45007 ( \44982 , \44959 );
or \U$45008 ( \44983 , \44981 , \44982 );
buf \U$45009 ( \44984 , \14468 );
buf \U$45010 ( \44985 , \44558 );
or \U$45011 ( \44986 , \44984 , \44985 );
buf \U$45012 ( \44987 , \22744 );
buf \U$45013 ( \44988 , \44379 );
not \U$45014 ( \44989 , \44988 );
buf \U$45015 ( \44990 , \44989 );
buf \U$45016 ( \44991 , \44990 );
or \U$45017 ( \44992 , \44987 , \44991 );
nand \U$45018 ( \44993 , \44986 , \44992 );
buf \U$45019 ( \44994 , \44993 );
buf \U$45020 ( \44995 , \44994 );
nand \U$45021 ( \44996 , \44983 , \44995 );
buf \U$45022 ( \44997 , \44996 );
buf \U$45023 ( \44998 , \44997 );
nand \U$45024 ( \44999 , \44980 , \44998 );
buf \U$45025 ( \45000 , \44999 );
buf \U$45026 ( \45001 , \45000 );
and \U$45027 ( \45002 , \44947 , \45001 );
and \U$45028 ( \45003 , \44879 , \44946 );
or \U$45029 ( \45004 , \45002 , \45003 );
buf \U$45030 ( \45005 , \45004 );
buf \U$45031 ( \45006 , \45005 );
xor \U$45032 ( \45007 , \44876 , \45006 );
buf \U$45033 ( \45008 , \45007 );
buf \U$45034 ( \45009 , \45008 );
xor \U$45035 ( \45010 , \44743 , \45009 );
buf \U$45036 ( \45011 , \45010 );
buf \U$45037 ( \45012 , \45011 );
xor \U$45038 ( \45013 , \44375 , \45012 );
xor \U$45039 ( \45014 , \43839 , \43882 );
xor \U$45040 ( \45015 , \45014 , \43963 );
buf \U$45041 ( \45016 , \45015 );
buf \U$45042 ( \45017 , \45016 );
buf \U$45043 ( \45018 , \44024 );
not \U$45044 ( \45019 , \45018 );
buf \U$45045 ( \45020 , \44165 );
buf \U$45046 ( \45021 , \44095 );
and \U$45047 ( \45022 , \45020 , \45021 );
not \U$45048 ( \45023 , \45020 );
buf \U$45049 ( \45024 , \44092 );
and \U$45050 ( \45025 , \45023 , \45024 );
nor \U$45051 ( \45026 , \45022 , \45025 );
buf \U$45052 ( \45027 , \45026 );
buf \U$45053 ( \45028 , \45027 );
not \U$45054 ( \45029 , \45028 );
buf \U$45055 ( \45030 , \45029 );
buf \U$45056 ( \45031 , \45030 );
not \U$45057 ( \45032 , \45031 );
or \U$45058 ( \45033 , \45019 , \45032 );
buf \U$45059 ( \45034 , \44024 );
not \U$45060 ( \45035 , \45034 );
buf \U$45061 ( \45036 , \45027 );
nand \U$45062 ( \45037 , \45035 , \45036 );
buf \U$45063 ( \45038 , \45037 );
buf \U$45064 ( \45039 , \45038 );
nand \U$45065 ( \45040 , \45033 , \45039 );
buf \U$45066 ( \45041 , \45040 );
buf \U$45067 ( \45042 , \45041 );
xor \U$45068 ( \45043 , \45017 , \45042 );
xor \U$45069 ( \45044 , RIc0da918_109, RIc0d8b90_46);
buf \U$45070 ( \45045 , \45044 );
not \U$45071 ( \45046 , \45045 );
buf \U$45072 ( \45047 , \13419 );
not \U$45073 ( \45048 , \45047 );
or \U$45074 ( \45049 , \45046 , \45048 );
buf \U$45075 ( \45050 , \14216 );
xor \U$45076 ( \45051 , RIc0da918_109, RIc0d8b18_45);
buf \U$45077 ( \45052 , \45051 );
nand \U$45078 ( \45053 , \45050 , \45052 );
buf \U$45079 ( \45054 , \45053 );
buf \U$45080 ( \45055 , \45054 );
nand \U$45081 ( \45056 , \45049 , \45055 );
buf \U$45082 ( \45057 , \45056 );
buf \U$45083 ( \45058 , \45057 );
xor \U$45084 ( \45059 , RIc0dacd8_117, RIc0d87d0_38);
buf \U$45085 ( \45060 , \45059 );
not \U$45086 ( \45061 , \45060 );
buf \U$45087 ( \45062 , \13146 );
not \U$45088 ( \45063 , \45062 );
or \U$45089 ( \45064 , \45061 , \45063 );
buf \U$45090 ( \45065 , \12937 );
buf \U$45091 ( \45066 , RIc0dacd8_117);
buf \U$45092 ( \45067 , RIc0d8758_37);
xor \U$45093 ( \45068 , \45066 , \45067 );
buf \U$45094 ( \45069 , \45068 );
buf \U$45095 ( \45070 , \45069 );
nand \U$45096 ( \45071 , \45065 , \45070 );
buf \U$45097 ( \45072 , \45071 );
buf \U$45098 ( \45073 , \45072 );
nand \U$45099 ( \45074 , \45064 , \45073 );
buf \U$45100 ( \45075 , \45074 );
buf \U$45101 ( \45076 , \45075 );
xor \U$45102 ( \45077 , \45058 , \45076 );
buf \U$45103 ( \45078 , RIc0d8488_31);
buf \U$45104 ( \45079 , RIc0dafa8_123);
xor \U$45105 ( \45080 , \45078 , \45079 );
buf \U$45106 ( \45081 , \45080 );
buf \U$45107 ( \45082 , \45081 );
not \U$45108 ( \45083 , \45082 );
buf \U$45109 ( \45084 , \16692 );
not \U$45110 ( \45085 , \45084 );
or \U$45111 ( \45086 , \45083 , \45085 );
buf \U$45112 ( \45087 , \14982 );
not \U$45113 ( \45088 , \45087 );
buf \U$45114 ( \45089 , \45088 );
buf \U$45115 ( \45090 , \45089 );
buf \U$45116 ( \45091 , RIc0d8500_32);
buf \U$45117 ( \45092 , RIc0dafa8_123);
xnor \U$45118 ( \45093 , \45091 , \45092 );
buf \U$45119 ( \45094 , \45093 );
buf \U$45120 ( \45095 , \45094 );
or \U$45121 ( \45096 , \45090 , \45095 );
nand \U$45122 ( \45097 , \45086 , \45096 );
buf \U$45123 ( \45098 , \45097 );
buf \U$45124 ( \45099 , \45098 );
and \U$45125 ( \45100 , \45077 , \45099 );
and \U$45126 ( \45101 , \45058 , \45076 );
or \U$45127 ( \45102 , \45100 , \45101 );
buf \U$45128 ( \45103 , \45102 );
buf \U$45129 ( \45104 , \45103 );
buf \U$45130 ( \45105 , RIc0db098_125);
buf \U$45131 ( \45106 , RIc0d8410_30);
xor \U$45132 ( \45107 , \45105 , \45106 );
buf \U$45133 ( \45108 , \45107 );
buf \U$45134 ( \45109 , \45108 );
not \U$45135 ( \45110 , \45109 );
buf \U$45136 ( \45111 , \17995 );
not \U$45137 ( \45112 , \45111 );
or \U$45138 ( \45113 , \45110 , \45112 );
buf \U$45139 ( \45114 , \13465 );
buf \U$45140 ( \45115 , \44549 );
nand \U$45141 ( \45116 , \45114 , \45115 );
buf \U$45142 ( \45117 , \45116 );
buf \U$45143 ( \45118 , \45117 );
nand \U$45144 ( \45119 , \45113 , \45118 );
buf \U$45145 ( \45120 , \45119 );
buf \U$45146 ( \45121 , \45120 );
xor \U$45147 ( \45122 , RIc0da558_101, RIc0d8f50_54);
buf \U$45148 ( \45123 , \45122 );
not \U$45149 ( \45124 , \45123 );
buf \U$45150 ( \45125 , \22631 );
not \U$45151 ( \45126 , \45125 );
or \U$45152 ( \45127 , \45124 , \45126 );
buf \U$45153 ( \45128 , \12839 );
buf \U$45154 ( \45129 , \44572 );
nand \U$45155 ( \45130 , \45128 , \45129 );
buf \U$45156 ( \45131 , \45130 );
buf \U$45157 ( \45132 , \45131 );
nand \U$45158 ( \45133 , \45127 , \45132 );
buf \U$45159 ( \45134 , \45133 );
buf \U$45160 ( \45135 , \45134 );
xor \U$45161 ( \45136 , \45121 , \45135 );
buf \U$45162 ( \45137 , RIc0dabe8_115);
buf \U$45163 ( \45138 , RIc0d88c0_40);
xor \U$45164 ( \45139 , \45137 , \45138 );
buf \U$45165 ( \45140 , \45139 );
buf \U$45166 ( \45141 , \45140 );
not \U$45167 ( \45142 , \45141 );
buf \U$45168 ( \45143 , \14186 );
not \U$45169 ( \45144 , \45143 );
or \U$45170 ( \45145 , \45142 , \45144 );
buf \U$45171 ( \45146 , RIc0dabe8_115);
buf \U$45172 ( \45147 , RIc0d8848_39);
xnor \U$45173 ( \45148 , \45146 , \45147 );
buf \U$45174 ( \45149 , \45148 );
buf \U$45175 ( \45150 , \45149 );
not \U$45176 ( \45151 , \45150 );
buf \U$45177 ( \45152 , \14690 );
nand \U$45178 ( \45153 , \45151 , \45152 );
buf \U$45179 ( \45154 , \45153 );
buf \U$45180 ( \45155 , \45154 );
nand \U$45181 ( \45156 , \45145 , \45155 );
buf \U$45182 ( \45157 , \45156 );
buf \U$45183 ( \45158 , \45157 );
and \U$45184 ( \45159 , \45136 , \45158 );
and \U$45185 ( \45160 , \45121 , \45135 );
or \U$45186 ( \45161 , \45159 , \45160 );
buf \U$45187 ( \45162 , \45161 );
buf \U$45188 ( \45163 , \45162 );
xor \U$45189 ( \45164 , \45104 , \45163 );
buf \U$45190 ( \45165 , RIc0da738_105);
buf \U$45191 ( \45166 , RIc0d8d70_50);
xor \U$45192 ( \45167 , \45165 , \45166 );
buf \U$45193 ( \45168 , \45167 );
buf \U$45194 ( \45169 , \45168 );
not \U$45195 ( \45170 , \45169 );
buf \U$45196 ( \45171 , \12736 );
not \U$45197 ( \45172 , \45171 );
or \U$45198 ( \45173 , \45170 , \45172 );
buf \U$45199 ( \45174 , \26301 );
buf \U$45200 ( \45175 , RIc0d8cf8_49);
buf \U$45201 ( \45176 , RIc0da738_105);
xor \U$45202 ( \45177 , \45175 , \45176 );
buf \U$45203 ( \45178 , \45177 );
buf \U$45204 ( \45179 , \45178 );
nand \U$45205 ( \45180 , \45174 , \45179 );
buf \U$45206 ( \45181 , \45180 );
buf \U$45207 ( \45182 , \45181 );
nand \U$45208 ( \45183 , \45173 , \45182 );
buf \U$45209 ( \45184 , \45183 );
buf \U$45210 ( \45185 , \45184 );
buf \U$45211 ( \45186 , RIc0daaf8_113);
buf \U$45212 ( \45187 , RIc0d89b0_42);
and \U$45213 ( \45188 , \45186 , \45187 );
not \U$45214 ( \45189 , \45186 );
buf \U$45215 ( \45190 , RIc0d89b0_42);
not \U$45216 ( \45191 , \45190 );
buf \U$45217 ( \45192 , \45191 );
buf \U$45218 ( \45193 , \45192 );
and \U$45219 ( \45194 , \45189 , \45193 );
nor \U$45220 ( \45195 , \45188 , \45194 );
buf \U$45221 ( \45196 , \45195 );
buf \U$45222 ( \45197 , \45196 );
not \U$45223 ( \45198 , \45197 );
buf \U$45224 ( \45199 , \26484 );
not \U$45225 ( \45200 , \45199 );
or \U$45226 ( \45201 , \45198 , \45200 );
buf \U$45227 ( \45202 , RIc0daaf8_113);
buf \U$45228 ( \45203 , RIc0d8938_41);
xnor \U$45229 ( \45204 , \45202 , \45203 );
buf \U$45230 ( \45205 , \45204 );
buf \U$45231 ( \45206 , \45205 );
not \U$45232 ( \45207 , \45206 );
buf \U$45233 ( \45208 , \12410 );
nand \U$45234 ( \45209 , \45207 , \45208 );
buf \U$45235 ( \45210 , \45209 );
buf \U$45236 ( \45211 , \45210 );
nand \U$45237 ( \45212 , \45201 , \45211 );
buf \U$45238 ( \45213 , \45212 );
buf \U$45239 ( \45214 , \45213 );
xor \U$45240 ( \45215 , \45185 , \45214 );
buf \U$45241 ( \45216 , \13178 );
buf \U$45242 ( \45217 , RIc0d86e0_36);
buf \U$45243 ( \45218 , RIc0dadc8_119);
xnor \U$45244 ( \45219 , \45217 , \45218 );
buf \U$45245 ( \45220 , \45219 );
buf \U$45246 ( \45221 , \45220 );
or \U$45247 ( \45222 , \45216 , \45221 );
buf \U$45248 ( \45223 , \13005 );
not \U$45249 ( \45224 , \45223 );
buf \U$45250 ( \45225 , \45224 );
buf \U$45251 ( \45226 , \45225 );
xor \U$45252 ( \45227 , RIc0dadc8_119, RIc0d8668_35);
buf \U$45253 ( \45228 , \45227 );
not \U$45254 ( \45229 , \45228 );
buf \U$45255 ( \45230 , \45229 );
buf \U$45256 ( \45231 , \45230 );
or \U$45257 ( \45232 , \45226 , \45231 );
nand \U$45258 ( \45233 , \45222 , \45232 );
buf \U$45259 ( \45234 , \45233 );
buf \U$45260 ( \45235 , \45234 );
and \U$45261 ( \45236 , \45215 , \45235 );
and \U$45262 ( \45237 , \45185 , \45214 );
or \U$45263 ( \45238 , \45236 , \45237 );
buf \U$45264 ( \45239 , \45238 );
buf \U$45265 ( \45240 , \45239 );
and \U$45266 ( \45241 , \45164 , \45240 );
and \U$45267 ( \45242 , \45104 , \45163 );
or \U$45268 ( \45243 , \45241 , \45242 );
buf \U$45269 ( \45244 , \45243 );
buf \U$45270 ( \45245 , \45244 );
xor \U$45271 ( \45246 , \44507 , \44544 );
xor \U$45272 ( \45247 , \45246 , \44621 );
buf \U$45273 ( \45248 , \45247 );
buf \U$45274 ( \45249 , \45248 );
xor \U$45275 ( \45250 , \45245 , \45249 );
buf \U$45276 ( \45251 , RIc0d8aa0_44);
buf \U$45277 ( \45252 , RIc0daa08_111);
xor \U$45278 ( \45253 , \45251 , \45252 );
buf \U$45279 ( \45254 , \45253 );
buf \U$45280 ( \45255 , \45254 );
not \U$45281 ( \45256 , \45255 );
buf \U$45282 ( \45257 , \18306 );
not \U$45283 ( \45258 , \45257 );
or \U$45284 ( \45259 , \45256 , \45258 );
buf \U$45285 ( \45260 , \18312 );
buf \U$45286 ( \45261 , RIc0d8a28_43);
buf \U$45287 ( \45262 , RIc0daa08_111);
xor \U$45288 ( \45263 , \45261 , \45262 );
buf \U$45289 ( \45264 , \45263 );
buf \U$45290 ( \45265 , \45264 );
nand \U$45291 ( \45266 , \45260 , \45265 );
buf \U$45292 ( \45267 , \45266 );
buf \U$45293 ( \45268 , \45267 );
nand \U$45294 ( \45269 , \45259 , \45268 );
buf \U$45295 ( \45270 , \45269 );
buf \U$45296 ( \45271 , \45270 );
not \U$45297 ( \45272 , \45271 );
buf \U$45298 ( \45273 , RIc0d8e60_52);
buf \U$45299 ( \45274 , RIc0da648_103);
xor \U$45300 ( \45275 , \45273 , \45274 );
buf \U$45301 ( \45276 , \45275 );
buf \U$45302 ( \45277 , \45276 );
not \U$45303 ( \45278 , \45277 );
buf \U$45304 ( \45279 , \13042 );
not \U$45305 ( \45280 , \45279 );
or \U$45306 ( \45281 , \45278 , \45280 );
buf \U$45307 ( \45282 , \16584 );
buf \U$45308 ( \45283 , \44598 );
nand \U$45309 ( \45284 , \45282 , \45283 );
buf \U$45310 ( \45285 , \45284 );
buf \U$45311 ( \45286 , \45285 );
nand \U$45312 ( \45287 , \45281 , \45286 );
buf \U$45313 ( \45288 , \45287 );
buf \U$45314 ( \45289 , \45288 );
not \U$45315 ( \45290 , \45289 );
or \U$45316 ( \45291 , \45272 , \45290 );
buf \U$45317 ( \45292 , \45288 );
buf \U$45318 ( \45293 , \45270 );
or \U$45319 ( \45294 , \45292 , \45293 );
xor \U$45320 ( \45295 , RIc0da828_107, RIc0d8c80_48);
buf \U$45321 ( \45296 , \45295 );
not \U$45322 ( \45297 , \45296 );
buf \U$45323 ( \45298 , \34202 );
not \U$45324 ( \45299 , \45298 );
or \U$45325 ( \45300 , \45297 , \45299 );
buf \U$45326 ( \45301 , \16071 );
buf \U$45327 ( \45302 , RIc0d8c08_47);
buf \U$45328 ( \45303 , RIc0da828_107);
xor \U$45329 ( \45304 , \45302 , \45303 );
buf \U$45330 ( \45305 , \45304 );
buf \U$45331 ( \45306 , \45305 );
nand \U$45332 ( \45307 , \45301 , \45306 );
buf \U$45333 ( \45308 , \45307 );
buf \U$45334 ( \45309 , \45308 );
nand \U$45335 ( \45310 , \45300 , \45309 );
buf \U$45336 ( \45311 , \45310 );
buf \U$45337 ( \45312 , \45311 );
nand \U$45338 ( \45313 , \45294 , \45312 );
buf \U$45339 ( \45314 , \45313 );
buf \U$45340 ( \45315 , \45314 );
nand \U$45341 ( \45316 , \45291 , \45315 );
buf \U$45342 ( \45317 , \45316 );
buf \U$45343 ( \45318 , \45317 );
buf \U$45344 ( \45319 , RIc0d8320_28);
buf \U$45345 ( \45320 , RIc0db188_127);
xor \U$45346 ( \45321 , \45319 , \45320 );
buf \U$45347 ( \45322 , \45321 );
buf \U$45348 ( \45323 , \45322 );
not \U$45349 ( \45324 , \45323 );
buf \U$45350 ( \45325 , \15609 );
not \U$45351 ( \45326 , \45325 );
or \U$45352 ( \45327 , \45324 , \45326 );
buf \U$45353 ( \45328 , RIc0d82a8_27);
buf \U$45354 ( \45329 , RIc0db188_127);
xor \U$45355 ( \45330 , \45328 , \45329 );
buf \U$45356 ( \45331 , \45330 );
buf \U$45357 ( \45332 , \45331 );
buf \U$45358 ( \45333 , RIc0db200_128);
nand \U$45359 ( \45334 , \45332 , \45333 );
buf \U$45360 ( \45335 , \45334 );
buf \U$45361 ( \45336 , \45335 );
nand \U$45362 ( \45337 , \45327 , \45336 );
buf \U$45363 ( \45338 , \45337 );
buf \U$45364 ( \45339 , \45338 );
buf \U$45365 ( \45340 , RIc0d9400_64);
buf \U$45366 ( \45341 , RIc0da0a8_91);
xor \U$45367 ( \45342 , \45340 , \45341 );
buf \U$45368 ( \45343 , \45342 );
buf \U$45369 ( \45344 , \45343 );
not \U$45370 ( \45345 , \45344 );
buf \U$45371 ( \45346 , \2535 );
not \U$45372 ( \45347 , \45346 );
or \U$45373 ( \45348 , \45345 , \45347 );
buf \U$45374 ( \45349 , \533 );
xor \U$45375 ( \45350 , RIc0da0a8_91, RIc0d9388_63);
buf \U$45376 ( \45351 , \45350 );
nand \U$45377 ( \45352 , \45349 , \45351 );
buf \U$45378 ( \45353 , \45352 );
buf \U$45379 ( \45354 , \45353 );
nand \U$45380 ( \45355 , \45348 , \45354 );
buf \U$45381 ( \45356 , \45355 );
buf \U$45382 ( \45357 , \45356 );
xor \U$45383 ( \45358 , \45339 , \45357 );
buf \U$45384 ( \45359 , RIc0da378_97);
buf \U$45385 ( \45360 , RIc0d9130_58);
xor \U$45386 ( \45361 , \45359 , \45360 );
buf \U$45387 ( \45362 , \45361 );
buf \U$45388 ( \45363 , \45362 );
not \U$45389 ( \45364 , \45363 );
buf \U$45390 ( \45365 , \2066 );
not \U$45391 ( \45366 , \45365 );
or \U$45392 ( \45367 , \45364 , \45366 );
buf \U$45393 ( \45368 , \734 );
xor \U$45394 ( \45369 , RIc0da378_97, RIc0d90b8_57);
buf \U$45395 ( \45370 , \45369 );
nand \U$45396 ( \45371 , \45368 , \45370 );
buf \U$45397 ( \45372 , \45371 );
buf \U$45398 ( \45373 , \45372 );
nand \U$45399 ( \45374 , \45367 , \45373 );
buf \U$45400 ( \45375 , \45374 );
buf \U$45401 ( \45376 , \45375 );
and \U$45402 ( \45377 , \45358 , \45376 );
and \U$45403 ( \45378 , \45339 , \45357 );
or \U$45404 ( \45379 , \45377 , \45378 );
buf \U$45405 ( \45380 , \45379 );
buf \U$45406 ( \45381 , \45380 );
xor \U$45407 ( \45382 , \45318 , \45381 );
buf \U$45408 ( \45383 , RIc0daeb8_121);
buf \U$45409 ( \45384 , RIc0d85f0_34);
xor \U$45410 ( \45385 , \45383 , \45384 );
buf \U$45411 ( \45386 , \45385 );
buf \U$45412 ( \45387 , \45386 );
not \U$45413 ( \45388 , \45387 );
buf \U$45414 ( \45389 , \19487 );
not \U$45415 ( \45390 , \45389 );
or \U$45416 ( \45391 , \45388 , \45390 );
buf \U$45417 ( \45392 , RIc0d8578_33);
buf \U$45418 ( \45393 , RIc0daeb8_121);
xnor \U$45419 ( \45394 , \45392 , \45393 );
buf \U$45420 ( \45395 , \45394 );
buf \U$45421 ( \45396 , \45395 );
not \U$45422 ( \45397 , \45396 );
buf \U$45423 ( \45398 , \13314 );
nand \U$45424 ( \45399 , \45397 , \45398 );
buf \U$45425 ( \45400 , \45399 );
buf \U$45426 ( \45401 , \45400 );
nand \U$45427 ( \45402 , \45391 , \45401 );
buf \U$45428 ( \45403 , \45402 );
buf \U$45429 ( \45404 , \45403 );
buf \U$45430 ( \45405 , RIc0da468_99);
buf \U$45431 ( \45406 , RIc0d9040_56);
xor \U$45432 ( \45407 , \45405 , \45406 );
buf \U$45433 ( \45408 , \45407 );
buf \U$45434 ( \45409 , \45408 );
not \U$45435 ( \45410 , \45409 );
buf \U$45436 ( \45411 , \2470 );
not \U$45437 ( \45412 , \45411 );
or \U$45438 ( \45413 , \45410 , \45412 );
buf \U$45439 ( \45414 , \16750 );
buf \U$45440 ( \45415 , RIc0da468_99);
buf \U$45441 ( \45416 , RIc0d8fc8_55);
xor \U$45442 ( \45417 , \45415 , \45416 );
buf \U$45443 ( \45418 , \45417 );
buf \U$45444 ( \45419 , \45418 );
nand \U$45445 ( \45420 , \45414 , \45419 );
buf \U$45446 ( \45421 , \45420 );
buf \U$45447 ( \45422 , \45421 );
nand \U$45448 ( \45423 , \45413 , \45422 );
buf \U$45449 ( \45424 , \45423 );
buf \U$45450 ( \45425 , \45424 );
xor \U$45451 ( \45426 , \45404 , \45425 );
xor \U$45452 ( \45427 , RIc0da288_95, RIc0d91a8_59);
buf \U$45453 ( \45428 , \45427 );
not \U$45454 ( \45429 , \45428 );
buf \U$45455 ( \45430 , \14707 );
not \U$45456 ( \45431 , \45430 );
or \U$45457 ( \45432 , \45429 , \45431 );
buf \U$45458 ( \45433 , \14713 );
buf \U$45459 ( \45434 , RIc0da288_95);
buf \U$45460 ( \45435 , RIc0d9220_60);
xnor \U$45461 ( \45436 , \45434 , \45435 );
buf \U$45462 ( \45437 , \45436 );
buf \U$45463 ( \45438 , \45437 );
or \U$45464 ( \45439 , \45433 , \45438 );
nand \U$45465 ( \45440 , \45432 , \45439 );
buf \U$45466 ( \45441 , \45440 );
buf \U$45467 ( \45442 , \45441 );
and \U$45468 ( \45443 , \45426 , \45442 );
and \U$45469 ( \45444 , \45404 , \45425 );
or \U$45470 ( \45445 , \45443 , \45444 );
buf \U$45471 ( \45446 , \45445 );
buf \U$45472 ( \45447 , \45446 );
and \U$45473 ( \45448 , \45382 , \45447 );
and \U$45474 ( \45449 , \45318 , \45381 );
or \U$45475 ( \45450 , \45448 , \45449 );
buf \U$45476 ( \45451 , \45450 );
buf \U$45477 ( \45452 , \45451 );
and \U$45478 ( \45453 , \45250 , \45452 );
and \U$45479 ( \45454 , \45245 , \45249 );
or \U$45480 ( \45455 , \45453 , \45454 );
buf \U$45481 ( \45456 , \45455 );
buf \U$45482 ( \45457 , \45456 );
and \U$45483 ( \45458 , \45043 , \45457 );
and \U$45484 ( \45459 , \45017 , \45042 );
or \U$45485 ( \45460 , \45458 , \45459 );
buf \U$45486 ( \45461 , \45460 );
buf \U$45487 ( \45462 , \45461 );
and \U$45488 ( \45463 , \45013 , \45462 );
and \U$45489 ( \45464 , \44375 , \45012 );
or \U$45490 ( \45465 , \45463 , \45464 );
buf \U$45491 ( \45466 , \45465 );
buf \U$45492 ( \45467 , \45466 );
buf \U$45493 ( \45468 , \44625 );
not \U$45494 ( \45469 , \45468 );
buf \U$45495 ( \45470 , \44431 );
buf \U$45496 ( \45471 , \44484 );
not \U$45497 ( \45472 , \45471 );
buf \U$45498 ( \45473 , \45472 );
buf \U$45499 ( \45474 , \45473 );
and \U$45500 ( \45475 , \45470 , \45474 );
not \U$45501 ( \45476 , \45470 );
buf \U$45502 ( \45477 , \44484 );
and \U$45503 ( \45478 , \45476 , \45477 );
nor \U$45504 ( \45479 , \45475 , \45478 );
buf \U$45505 ( \45480 , \45479 );
buf \U$45506 ( \45481 , \45480 );
not \U$45507 ( \45482 , \45481 );
or \U$45508 ( \45483 , \45469 , \45482 );
buf \U$45509 ( \45484 , \45480 );
buf \U$45510 ( \45485 , \44625 );
or \U$45511 ( \45486 , \45484 , \45485 );
nand \U$45512 ( \45487 , \45483 , \45486 );
buf \U$45513 ( \45488 , \45487 );
buf \U$45514 ( \45489 , \45488 );
buf \U$45515 ( \45490 , \16477 );
buf \U$45516 ( \45491 , RIc0d9400_64);
and \U$45517 ( \45492 , \45490 , \45491 );
buf \U$45518 ( \45493 , \45492 );
buf \U$45519 ( \45494 , \45493 );
buf \U$45520 ( \45495 , RIc0d9298_61);
buf \U$45521 ( \45496 , RIc0da198_93);
xor \U$45522 ( \45497 , \45495 , \45496 );
buf \U$45523 ( \45498 , \45497 );
buf \U$45524 ( \45499 , \45498 );
not \U$45525 ( \45500 , \45499 );
buf \U$45526 ( \45501 , \1901 );
not \U$45527 ( \45502 , \45501 );
or \U$45528 ( \45503 , \45500 , \45502 );
buf \U$45529 ( \45504 , \4008 );
buf \U$45530 ( \45505 , \44332 );
nand \U$45531 ( \45506 , \45504 , \45505 );
buf \U$45532 ( \45507 , \45506 );
buf \U$45533 ( \45508 , \45507 );
nand \U$45534 ( \45509 , \45503 , \45508 );
buf \U$45535 ( \45510 , \45509 );
buf \U$45536 ( \45511 , \45510 );
xor \U$45537 ( \45512 , \45494 , \45511 );
buf \U$45538 ( \45513 , \45069 );
not \U$45539 ( \45514 , \45513 );
buf \U$45540 ( \45515 , \22350 );
not \U$45541 ( \45516 , \45515 );
or \U$45542 ( \45517 , \45514 , \45516 );
buf \U$45543 ( \45518 , \44888 );
not \U$45544 ( \45519 , \45518 );
buf \U$45545 ( \45520 , \12937 );
nand \U$45546 ( \45521 , \45519 , \45520 );
buf \U$45547 ( \45522 , \45521 );
buf \U$45548 ( \45523 , \45522 );
nand \U$45549 ( \45524 , \45517 , \45523 );
buf \U$45550 ( \45525 , \45524 );
buf \U$45551 ( \45526 , \45525 );
xnor \U$45552 ( \45527 , \45512 , \45526 );
buf \U$45553 ( \45528 , \45527 );
buf \U$45554 ( \45529 , \45528 );
not \U$45555 ( \45530 , \45529 );
buf \U$45556 ( \45531 , \45530 );
buf \U$45557 ( \45532 , \45531 );
not \U$45558 ( \45533 , \45532 );
buf \U$45559 ( \45534 , \45051 );
not \U$45560 ( \45535 , \45534 );
buf \U$45561 ( \45536 , \21959 );
not \U$45562 ( \45537 , \45536 );
or \U$45563 ( \45538 , \45535 , \45537 );
buf \U$45564 ( \45539 , \16232 );
buf \U$45565 ( \45540 , \44198 );
nand \U$45566 ( \45541 , \45539 , \45540 );
buf \U$45567 ( \45542 , \45541 );
buf \U$45568 ( \45543 , \45542 );
nand \U$45569 ( \45544 , \45538 , \45543 );
buf \U$45570 ( \45545 , \45544 );
buf \U$45571 ( \45546 , \13310 );
not \U$45572 ( \45547 , \45546 );
buf \U$45573 ( \45548 , \45547 );
buf \U$45574 ( \45549 , \45548 );
not \U$45575 ( \45550 , \45549 );
buf \U$45576 ( \45551 , \45395 );
not \U$45577 ( \45552 , \45551 );
and \U$45578 ( \45553 , \45550 , \45552 );
buf \U$45579 ( \45554 , \44315 );
not \U$45580 ( \45555 , \45554 );
buf \U$45581 ( \45556 , \13314 );
not \U$45582 ( \45557 , \45556 );
buf \U$45583 ( \45558 , \45557 );
buf \U$45584 ( \45559 , \45558 );
nor \U$45585 ( \45560 , \45555 , \45559 );
buf \U$45586 ( \45561 , \45560 );
buf \U$45587 ( \45562 , \45561 );
nor \U$45588 ( \45563 , \45553 , \45562 );
buf \U$45589 ( \45564 , \45563 );
xor \U$45590 ( \45565 , \45545 , \45564 );
buf \U$45591 ( \45566 , \45081 );
not \U$45592 ( \45567 , \45566 );
buf \U$45593 ( \45568 , \16688 );
not \U$45594 ( \45569 , \45568 );
buf \U$45595 ( \45570 , \45569 );
buf \U$45596 ( \45571 , \45570 );
not \U$45597 ( \45572 , \45571 );
or \U$45598 ( \45573 , \45567 , \45572 );
buf \U$45599 ( \45574 , \14278 );
buf \U$45600 ( \45575 , \44290 );
nand \U$45601 ( \45576 , \45574 , \45575 );
buf \U$45602 ( \45577 , \45576 );
buf \U$45603 ( \45578 , \45577 );
nand \U$45604 ( \45579 , \45573 , \45578 );
buf \U$45605 ( \45580 , \45579 );
xor \U$45606 ( \45581 , \45565 , \45580 );
buf \U$45607 ( \45582 , \45581 );
not \U$45608 ( \45583 , \45582 );
buf \U$45609 ( \45584 , \45583 );
buf \U$45610 ( \45585 , \45584 );
not \U$45611 ( \45586 , \45585 );
or \U$45612 ( \45587 , \45533 , \45586 );
buf \U$45613 ( \45588 , \45528 );
not \U$45614 ( \45589 , \45588 );
buf \U$45615 ( \45590 , \45581 );
not \U$45616 ( \45591 , \45590 );
or \U$45617 ( \45592 , \45589 , \45591 );
not \U$45618 ( \45593 , \14888 );
not \U$45619 ( \45594 , \45205 );
and \U$45620 ( \45595 , \45593 , \45594 );
buf \U$45621 ( \45596 , \34244 );
buf \U$45622 ( \45597 , \44264 );
nor \U$45623 ( \45598 , \45596 , \45597 );
buf \U$45624 ( \45599 , \45598 );
nor \U$45625 ( \45600 , \45595 , \45599 );
buf \U$45626 ( \45601 , \45418 );
not \U$45627 ( \45602 , \45601 );
buf \U$45628 ( \45603 , \14419 );
not \U$45629 ( \45604 , \45603 );
or \U$45630 ( \45605 , \45602 , \45604 );
buf \U$45631 ( \45606 , \2476 );
buf \U$45632 ( \45607 , \44965 );
nand \U$45633 ( \45608 , \45606 , \45607 );
buf \U$45634 ( \45609 , \45608 );
buf \U$45635 ( \45610 , \45609 );
nand \U$45636 ( \45611 , \45605 , \45610 );
buf \U$45637 ( \45612 , \45611 );
xor \U$45638 ( \45613 , \45600 , \45612 );
buf \U$45639 ( \45614 , \45427 );
not \U$45640 ( \45615 , \45614 );
buf \U$45641 ( \45616 , \27591 );
not \U$45642 ( \45617 , \45616 );
or \U$45643 ( \45618 , \45615 , \45617 );
buf \U$45644 ( \45619 , \344 );
buf \U$45645 ( \45620 , \43799 );
nand \U$45646 ( \45621 , \45619 , \45620 );
buf \U$45647 ( \45622 , \45621 );
buf \U$45648 ( \45623 , \45622 );
nand \U$45649 ( \45624 , \45618 , \45623 );
buf \U$45650 ( \45625 , \45624 );
xnor \U$45651 ( \45626 , \45613 , \45625 );
buf \U$45652 ( \45627 , \45626 );
nand \U$45653 ( \45628 , \45592 , \45627 );
buf \U$45654 ( \45629 , \45628 );
buf \U$45655 ( \45630 , \45629 );
nand \U$45656 ( \45631 , \45587 , \45630 );
buf \U$45657 ( \45632 , \45631 );
buf \U$45658 ( \45633 , \45632 );
buf \U$45659 ( \45634 , \44218 );
not \U$45660 ( \45635 , \45634 );
buf \U$45661 ( \45636 , \13005 );
not \U$45662 ( \45637 , \45636 );
or \U$45663 ( \45638 , \45635 , \45637 );
buf \U$45664 ( \45639 , \45225 );
buf \U$45665 ( \45640 , \45227 );
buf \U$45666 ( \45641 , \12995 );
nand \U$45667 ( \45642 , \45639 , \45640 , \45641 );
buf \U$45668 ( \45643 , \45642 );
buf \U$45669 ( \45644 , \45643 );
nand \U$45670 ( \45645 , \45638 , \45644 );
buf \U$45671 ( \45646 , \45645 );
buf \U$45672 ( \45647 , \45646 );
buf \U$45673 ( \45648 , \45178 );
not \U$45674 ( \45649 , \45648 );
buf \U$45675 ( \45650 , \25475 );
not \U$45676 ( \45651 , \45650 );
or \U$45677 ( \45652 , \45649 , \45651 );
buf \U$45678 ( \45653 , \15653 );
buf \U$45679 ( \45654 , \44176 );
nand \U$45680 ( \45655 , \45653 , \45654 );
buf \U$45681 ( \45656 , \45655 );
buf \U$45682 ( \45657 , \45656 );
nand \U$45683 ( \45658 , \45652 , \45657 );
buf \U$45684 ( \45659 , \45658 );
buf \U$45685 ( \45660 , \45659 );
xor \U$45686 ( \45661 , \45647 , \45660 );
buf \U$45687 ( \45662 , \14681 );
buf \U$45688 ( \45663 , \45149 );
or \U$45689 ( \45664 , \45662 , \45663 );
buf \U$45690 ( \45665 , \29865 );
buf \U$45691 ( \45666 , \43819 );
or \U$45692 ( \45667 , \45665 , \45666 );
nand \U$45693 ( \45668 , \45664 , \45667 );
buf \U$45694 ( \45669 , \45668 );
buf \U$45695 ( \45670 , \45669 );
xor \U$45696 ( \45671 , \45661 , \45670 );
buf \U$45697 ( \45672 , \45671 );
buf \U$45698 ( \45673 , \45672 );
not \U$45699 ( \45674 , \45673 );
xor \U$45700 ( \45675 , \44566 , \44588 );
xnor \U$45701 ( \45676 , \45675 , \44614 );
buf \U$45702 ( \45677 , \45676 );
not \U$45703 ( \45678 , \45677 );
buf \U$45704 ( \45679 , \45678 );
buf \U$45705 ( \45680 , \45679 );
not \U$45706 ( \45681 , \45680 );
or \U$45707 ( \45682 , \45674 , \45681 );
buf \U$45708 ( \45683 , \45672 );
not \U$45709 ( \45684 , \45683 );
buf \U$45710 ( \45685 , \45684 );
buf \U$45711 ( \45686 , \45685 );
not \U$45712 ( \45687 , \45686 );
buf \U$45713 ( \45688 , \45676 );
not \U$45714 ( \45689 , \45688 );
or \U$45715 ( \45690 , \45687 , \45689 );
buf \U$45716 ( \45691 , \45331 );
not \U$45717 ( \45692 , \45691 );
buf \U$45718 ( \45693 , \44639 );
not \U$45719 ( \45694 , \45693 );
or \U$45720 ( \45695 , \45692 , \45694 );
buf \U$45721 ( \45696 , \43786 );
buf \U$45722 ( \45697 , RIc0db200_128);
nand \U$45723 ( \45698 , \45696 , \45697 );
buf \U$45724 ( \45699 , \45698 );
buf \U$45725 ( \45700 , \45699 );
nand \U$45726 ( \45701 , \45695 , \45700 );
buf \U$45727 ( \45702 , \45701 );
buf \U$45728 ( \45703 , \45702 );
buf \U$45729 ( \45704 , \45305 );
not \U$45730 ( \45705 , \45704 );
buf \U$45731 ( \45706 , \19414 );
not \U$45732 ( \45707 , \45706 );
or \U$45733 ( \45708 , \45705 , \45707 );
buf \U$45734 ( \45709 , \16071 );
buf \U$45735 ( \45710 , \44350 );
nand \U$45736 ( \45711 , \45709 , \45710 );
buf \U$45737 ( \45712 , \45711 );
buf \U$45738 ( \45713 , \45712 );
nand \U$45739 ( \45714 , \45708 , \45713 );
buf \U$45740 ( \45715 , \45714 );
buf \U$45741 ( \45716 , \45715 );
xor \U$45742 ( \45717 , \45703 , \45716 );
buf \U$45743 ( \45718 , \45264 );
not \U$45744 ( \45719 , \45718 );
buf \U$45745 ( \45720 , \18306 );
not \U$45746 ( \45721 , \45720 );
or \U$45747 ( \45722 , \45719 , \45721 );
buf \U$45748 ( \45723 , \14352 );
not \U$45749 ( \45724 , \45723 );
buf \U$45750 ( \45725 , \45724 );
buf \U$45751 ( \45726 , \45725 );
not \U$45752 ( \45727 , \45726 );
buf \U$45753 ( \45728 , \45727 );
buf \U$45754 ( \45729 , \45728 );
buf \U$45755 ( \45730 , \44242 );
nand \U$45756 ( \45731 , \45729 , \45730 );
buf \U$45757 ( \45732 , \45731 );
buf \U$45758 ( \45733 , \45732 );
nand \U$45759 ( \45734 , \45722 , \45733 );
buf \U$45760 ( \45735 , \45734 );
buf \U$45761 ( \45736 , \45735 );
xnor \U$45762 ( \45737 , \45717 , \45736 );
buf \U$45763 ( \45738 , \45737 );
buf \U$45764 ( \45739 , \45738 );
not \U$45765 ( \45740 , \45739 );
buf \U$45766 ( \45741 , \45740 );
buf \U$45767 ( \45742 , \45741 );
nand \U$45768 ( \45743 , \45690 , \45742 );
buf \U$45769 ( \45744 , \45743 );
buf \U$45770 ( \45745 , \45744 );
nand \U$45771 ( \45746 , \45682 , \45745 );
buf \U$45772 ( \45747 , \45746 );
buf \U$45773 ( \45748 , \45747 );
xor \U$45774 ( \45749 , \45633 , \45748 );
xor \U$45775 ( \45750 , \45647 , \45660 );
and \U$45776 ( \45751 , \45750 , \45670 );
and \U$45777 ( \45752 , \45647 , \45660 );
or \U$45778 ( \45753 , \45751 , \45752 );
buf \U$45779 ( \45754 , \45753 );
buf \U$45780 ( \45755 , \45754 );
buf \U$45781 ( \45756 , \45625 );
buf \U$45782 ( \45757 , \45612 );
nor \U$45783 ( \45758 , \45756 , \45757 );
buf \U$45784 ( \45759 , \45758 );
buf \U$45785 ( \45760 , \45759 );
buf \U$45786 ( \45761 , \45600 );
or \U$45787 ( \45762 , \45760 , \45761 );
buf \U$45788 ( \45763 , \45625 );
buf \U$45789 ( \45764 , \45612 );
nand \U$45790 ( \45765 , \45763 , \45764 );
buf \U$45791 ( \45766 , \45765 );
buf \U$45792 ( \45767 , \45766 );
nand \U$45793 ( \45768 , \45762 , \45767 );
buf \U$45794 ( \45769 , \45768 );
buf \U$45795 ( \45770 , \45769 );
xor \U$45796 ( \45771 , \45755 , \45770 );
xor \U$45797 ( \45772 , \44328 , \44345 );
xor \U$45798 ( \45773 , \45772 , \44363 );
buf \U$45799 ( \45774 , \45773 );
buf \U$45800 ( \45775 , \45774 );
xor \U$45801 ( \45776 , \45771 , \45775 );
buf \U$45802 ( \45777 , \45776 );
buf \U$45803 ( \45778 , \45777 );
and \U$45804 ( \45779 , \45749 , \45778 );
and \U$45805 ( \45780 , \45633 , \45748 );
or \U$45806 ( \45781 , \45779 , \45780 );
buf \U$45807 ( \45782 , \45781 );
buf \U$45808 ( \45783 , \45782 );
xor \U$45809 ( \45784 , \45489 , \45783 );
buf \U$45810 ( \45785 , \45525 );
buf \U$45811 ( \45786 , \45493 );
nor \U$45812 ( \45787 , \45785 , \45786 );
buf \U$45813 ( \45788 , \45787 );
buf \U$45814 ( \45789 , \45788 );
buf \U$45815 ( \45790 , \45510 );
not \U$45816 ( \45791 , \45790 );
buf \U$45817 ( \45792 , \45791 );
buf \U$45818 ( \45793 , \45792 );
or \U$45819 ( \45794 , \45789 , \45793 );
buf \U$45820 ( \45795 , \45525 );
buf \U$45821 ( \45796 , \45493 );
nand \U$45822 ( \45797 , \45795 , \45796 );
buf \U$45823 ( \45798 , \45797 );
buf \U$45824 ( \45799 , \45798 );
nand \U$45825 ( \45800 , \45794 , \45799 );
buf \U$45826 ( \45801 , \45800 );
buf \U$45827 ( \45802 , \45801 );
not \U$45828 ( \45803 , \45802 );
buf \U$45829 ( \45804 , \45803 );
buf \U$45830 ( \45805 , \45804 );
not \U$45831 ( \45806 , \45805 );
buf \U$45832 ( \45807 , \45702 );
buf \U$45833 ( \45808 , \45715 );
or \U$45834 ( \45809 , \45807 , \45808 );
buf \U$45835 ( \45810 , \45735 );
nand \U$45836 ( \45811 , \45809 , \45810 );
buf \U$45837 ( \45812 , \45811 );
buf \U$45838 ( \45813 , \45812 );
buf \U$45839 ( \45814 , \45715 );
buf \U$45840 ( \45815 , \45702 );
nand \U$45841 ( \45816 , \45814 , \45815 );
buf \U$45842 ( \45817 , \45816 );
buf \U$45843 ( \45818 , \45817 );
nand \U$45844 ( \45819 , \45813 , \45818 );
buf \U$45845 ( \45820 , \45819 );
buf \U$45846 ( \45821 , \45564 );
not \U$45847 ( \45822 , \45821 );
buf \U$45848 ( \45823 , \45545 );
not \U$45849 ( \45824 , \45823 );
buf \U$45850 ( \45825 , \45824 );
buf \U$45851 ( \45826 , \45825 );
not \U$45852 ( \45827 , \45826 );
or \U$45853 ( \45828 , \45822 , \45827 );
buf \U$45854 ( \45829 , \45580 );
nand \U$45855 ( \45830 , \45828 , \45829 );
buf \U$45856 ( \45831 , \45830 );
buf \U$45857 ( \45832 , \45831 );
buf \U$45858 ( \45833 , \45564 );
not \U$45859 ( \45834 , \45833 );
buf \U$45860 ( \45835 , \45545 );
nand \U$45861 ( \45836 , \45834 , \45835 );
buf \U$45862 ( \45837 , \45836 );
buf \U$45863 ( \45838 , \45837 );
nand \U$45864 ( \45839 , \45832 , \45838 );
buf \U$45865 ( \45840 , \45839 );
xor \U$45866 ( \45841 , \45820 , \45840 );
buf \U$45867 ( \45842 , \45841 );
not \U$45868 ( \45843 , \45842 );
or \U$45869 ( \45844 , \45806 , \45843 );
buf \U$45870 ( \45845 , \45841 );
buf \U$45871 ( \45846 , \45804 );
or \U$45872 ( \45847 , \45845 , \45846 );
nand \U$45873 ( \45848 , \45844 , \45847 );
buf \U$45874 ( \45849 , \45848 );
buf \U$45875 ( \45850 , \45849 );
xor \U$45876 ( \45851 , \44192 , \44230 );
xor \U$45877 ( \45852 , \45851 , \44211 );
buf \U$45878 ( \45853 , \45852 );
buf \U$45879 ( \45854 , \44939 );
not \U$45880 ( \45855 , \45854 );
buf \U$45881 ( \45856 , \44912 );
not \U$45882 ( \45857 , \45856 );
or \U$45883 ( \45858 , \45855 , \45857 );
buf \U$45884 ( \45859 , \44935 );
buf \U$45885 ( \45860 , \44901 );
nand \U$45886 ( \45861 , \45859 , \45860 );
buf \U$45887 ( \45862 , \45861 );
buf \U$45888 ( \45863 , \45862 );
nand \U$45889 ( \45864 , \45858 , \45863 );
buf \U$45890 ( \45865 , \45864 );
xor \U$45891 ( \45866 , \44928 , \45865 );
buf \U$45892 ( \45867 , \45866 );
xor \U$45893 ( \45868 , \45853 , \45867 );
xor \U$45894 ( \45869 , \43795 , \43813 );
xor \U$45895 ( \45870 , \45869 , \43834 );
buf \U$45896 ( \45871 , \45870 );
buf \U$45897 ( \45872 , \45871 );
xor \U$45898 ( \45873 , \45868 , \45872 );
buf \U$45899 ( \45874 , \45873 );
buf \U$45900 ( \45875 , \45874 );
xor \U$45901 ( \45876 , \45850 , \45875 );
buf \U$45902 ( \45877 , \521 );
buf \U$45903 ( \45878 , \45350 );
not \U$45904 ( \45879 , \45878 );
buf \U$45905 ( \45880 , \45879 );
buf \U$45906 ( \45881 , \45880 );
or \U$45907 ( \45882 , \45877 , \45881 );
buf \U$45908 ( \45883 , \13293 );
not \U$45909 ( \45884 , \45883 );
buf \U$45910 ( \45885 , \45884 );
buf \U$45911 ( \45886 , \45885 );
buf \U$45912 ( \45887 , \44527 );
not \U$45913 ( \45888 , \45887 );
buf \U$45914 ( \45889 , \45888 );
buf \U$45915 ( \45890 , \45889 );
or \U$45916 ( \45891 , \45886 , \45890 );
nand \U$45917 ( \45892 , \45882 , \45891 );
buf \U$45918 ( \45893 , \45892 );
buf \U$45919 ( \45894 , \45893 );
buf \U$45920 ( \45895 , \45369 );
not \U$45921 ( \45896 , \45895 );
buf \U$45922 ( \45897 , \2066 );
not \U$45923 ( \45898 , \45897 );
or \U$45924 ( \45899 , \45896 , \45898 );
buf \U$45925 ( \45900 , \44908 );
not \U$45926 ( \45901 , \45900 );
buf \U$45927 ( \45902 , \2070 );
nand \U$45928 ( \45903 , \45901 , \45902 );
buf \U$45929 ( \45904 , \45903 );
buf \U$45930 ( \45905 , \45904 );
nand \U$45931 ( \45906 , \45899 , \45905 );
buf \U$45932 ( \45907 , \45906 );
buf \U$45933 ( \45908 , \45907 );
xor \U$45934 ( \45909 , \45894 , \45908 );
buf \U$45935 ( \45910 , RIc0d9400_64);
buf \U$45936 ( \45911 , RIc0da120_92);
or \U$45937 ( \45912 , \45910 , \45911 );
buf \U$45938 ( \45913 , RIc0da198_93);
nand \U$45939 ( \45914 , \45912 , \45913 );
buf \U$45940 ( \45915 , \45914 );
buf \U$45941 ( \45916 , \45915 );
buf \U$45942 ( \45917 , RIc0d9400_64);
buf \U$45943 ( \45918 , RIc0da120_92);
nand \U$45944 ( \45919 , \45917 , \45918 );
buf \U$45945 ( \45920 , \45919 );
buf \U$45946 ( \45921 , \45920 );
buf \U$45947 ( \45922 , RIc0da0a8_91);
and \U$45948 ( \45923 , \45916 , \45921 , \45922 );
buf \U$45949 ( \45924 , \45923 );
buf \U$45950 ( \45925 , \45924 );
buf \U$45951 ( \45926 , RIc0d9310_62);
buf \U$45952 ( \45927 , RIc0da198_93);
xor \U$45953 ( \45928 , \45926 , \45927 );
buf \U$45954 ( \45929 , \45928 );
buf \U$45955 ( \45930 , \45929 );
not \U$45956 ( \45931 , \45930 );
buf \U$45957 ( \45932 , \3415 );
not \U$45958 ( \45933 , \45932 );
or \U$45959 ( \45934 , \45931 , \45933 );
buf \U$45960 ( \45935 , \4008 );
buf \U$45961 ( \45936 , \45498 );
nand \U$45962 ( \45937 , \45935 , \45936 );
buf \U$45963 ( \45938 , \45937 );
buf \U$45964 ( \45939 , \45938 );
nand \U$45965 ( \45940 , \45934 , \45939 );
buf \U$45966 ( \45941 , \45940 );
buf \U$45967 ( \45942 , \45941 );
and \U$45968 ( \45943 , \45925 , \45942 );
buf \U$45969 ( \45944 , \45943 );
buf \U$45970 ( \45945 , \45944 );
and \U$45971 ( \45946 , \45909 , \45945 );
and \U$45972 ( \45947 , \45894 , \45908 );
or \U$45973 ( \45948 , \45946 , \45947 );
buf \U$45974 ( \45949 , \45948 );
buf \U$45975 ( \45950 , \45949 );
xor \U$45976 ( \45951 , \44994 , \44977 );
xor \U$45977 ( \45952 , \45951 , \44959 );
buf \U$45978 ( \45953 , \45952 );
xor \U$45979 ( \45954 , \45950 , \45953 );
buf \U$45980 ( \45955 , \44278 );
not \U$45981 ( \45956 , \45955 );
xnor \U$45982 ( \45957 , \44302 , \44254 );
buf \U$45983 ( \45958 , \45957 );
not \U$45984 ( \45959 , \45958 );
or \U$45985 ( \45960 , \45956 , \45959 );
buf \U$45986 ( \45961 , \45957 );
buf \U$45987 ( \45962 , \44278 );
or \U$45988 ( \45963 , \45961 , \45962 );
nand \U$45989 ( \45964 , \45960 , \45963 );
buf \U$45990 ( \45965 , \45964 );
buf \U$45991 ( \45966 , \45965 );
xor \U$45992 ( \45967 , \45954 , \45966 );
buf \U$45993 ( \45968 , \45967 );
buf \U$45994 ( \45969 , \45968 );
and \U$45995 ( \45970 , \45876 , \45969 );
and \U$45996 ( \45971 , \45850 , \45875 );
or \U$45997 ( \45972 , \45970 , \45971 );
buf \U$45998 ( \45973 , \45972 );
buf \U$45999 ( \45974 , \45973 );
and \U$46000 ( \45975 , \45784 , \45974 );
and \U$46001 ( \45976 , \45489 , \45783 );
or \U$46002 ( \45977 , \45975 , \45976 );
buf \U$46003 ( \45978 , \45977 );
buf \U$46004 ( \45979 , \45978 );
buf \U$46005 ( \45980 , \45820 );
not \U$46006 ( \45981 , \45980 );
buf \U$46007 ( \45982 , \45801 );
not \U$46008 ( \45983 , \45982 );
or \U$46009 ( \45984 , \45981 , \45983 );
buf \U$46010 ( \45985 , \45820 );
buf \U$46011 ( \45986 , \45801 );
or \U$46012 ( \45987 , \45985 , \45986 );
buf \U$46013 ( \45988 , \45840 );
nand \U$46014 ( \45989 , \45987 , \45988 );
buf \U$46015 ( \45990 , \45989 );
buf \U$46016 ( \45991 , \45990 );
nand \U$46017 ( \45992 , \45984 , \45991 );
buf \U$46018 ( \45993 , \45992 );
buf \U$46019 ( \45994 , \45993 );
not \U$46020 ( \45995 , \45994 );
xor \U$46021 ( \45996 , \44236 , \44367 );
xnor \U$46022 ( \45997 , \45996 , \44308 );
buf \U$46023 ( \45998 , \45997 );
not \U$46024 ( \45999 , \45998 );
buf \U$46025 ( \46000 , \45999 );
buf \U$46026 ( \46001 , \46000 );
not \U$46027 ( \46002 , \46001 );
or \U$46028 ( \46003 , \45995 , \46002 );
buf \U$46029 ( \46004 , \45993 );
not \U$46030 ( \46005 , \46004 );
buf \U$46031 ( \46006 , \46005 );
buf \U$46032 ( \46007 , \46006 );
not \U$46033 ( \46008 , \46007 );
buf \U$46034 ( \46009 , \45997 );
not \U$46035 ( \46010 , \46009 );
or \U$46036 ( \46011 , \46008 , \46010 );
xor \U$46037 ( \46012 , \45853 , \45867 );
and \U$46038 ( \46013 , \46012 , \45872 );
and \U$46039 ( \46014 , \45853 , \45867 );
or \U$46040 ( \46015 , \46013 , \46014 );
buf \U$46041 ( \46016 , \46015 );
buf \U$46042 ( \46017 , \46016 );
nand \U$46043 ( \46018 , \46011 , \46017 );
buf \U$46044 ( \46019 , \46018 );
buf \U$46045 ( \46020 , \46019 );
nand \U$46046 ( \46021 , \46003 , \46020 );
buf \U$46047 ( \46022 , \46021 );
buf \U$46048 ( \46023 , \46022 );
xor \U$46049 ( \46024 , \45755 , \45770 );
and \U$46050 ( \46025 , \46024 , \45775 );
and \U$46051 ( \46026 , \45755 , \45770 );
or \U$46052 ( \46027 , \46025 , \46026 );
buf \U$46053 ( \46028 , \46027 );
buf \U$46054 ( \46029 , \46028 );
xor \U$46055 ( \46030 , \44879 , \44946 );
xor \U$46056 ( \46031 , \46030 , \45001 );
buf \U$46057 ( \46032 , \46031 );
buf \U$46058 ( \46033 , \46032 );
xor \U$46059 ( \46034 , \46029 , \46033 );
xor \U$46060 ( \46035 , \45950 , \45953 );
and \U$46061 ( \46036 , \46035 , \45966 );
and \U$46062 ( \46037 , \45950 , \45953 );
or \U$46063 ( \46038 , \46036 , \46037 );
buf \U$46064 ( \46039 , \46038 );
buf \U$46065 ( \46040 , \46039 );
and \U$46066 ( \46041 , \46034 , \46040 );
and \U$46067 ( \46042 , \46029 , \46033 );
or \U$46068 ( \46043 , \46041 , \46042 );
buf \U$46069 ( \46044 , \46043 );
buf \U$46070 ( \46045 , \46044 );
xor \U$46071 ( \46046 , \46023 , \46045 );
buf \U$46072 ( \46047 , \44002 );
not \U$46073 ( \46048 , \46047 );
buf \U$46074 ( \46049 , \43983 );
not \U$46075 ( \46050 , \46049 );
or \U$46076 ( \46051 , \46048 , \46050 );
buf \U$46077 ( \46052 , \43983 );
buf \U$46078 ( \46053 , \44002 );
or \U$46079 ( \46054 , \46052 , \46053 );
buf \U$46080 ( \46055 , \44023 );
nand \U$46081 ( \46056 , \46054 , \46055 );
buf \U$46082 ( \46057 , \46056 );
buf \U$46083 ( \46058 , \46057 );
nand \U$46084 ( \46059 , \46051 , \46058 );
buf \U$46085 ( \46060 , \46059 );
buf \U$46086 ( \46061 , \44164 );
not \U$46087 ( \46062 , \46061 );
buf \U$46088 ( \46063 , \44146 );
not \U$46089 ( \46064 , \46063 );
or \U$46090 ( \46065 , \46062 , \46064 );
buf \U$46091 ( \46066 , \44146 );
buf \U$46092 ( \46067 , \44164 );
or \U$46093 ( \46068 , \46066 , \46067 );
buf \U$46094 ( \46069 , \44126 );
nand \U$46095 ( \46070 , \46068 , \46069 );
buf \U$46096 ( \46071 , \46070 );
buf \U$46097 ( \46072 , \46071 );
nand \U$46098 ( \46073 , \46065 , \46072 );
buf \U$46099 ( \46074 , \46073 );
xor \U$46100 ( \46075 , \46060 , \46074 );
buf \U$46101 ( \46076 , \43959 );
not \U$46102 ( \46077 , \46076 );
buf \U$46103 ( \46078 , \43900 );
not \U$46104 ( \46079 , \46078 );
or \U$46105 ( \46080 , \46077 , \46079 );
buf \U$46106 ( \46081 , \43900 );
buf \U$46107 ( \46082 , \43959 );
or \U$46108 ( \46083 , \46081 , \46082 );
buf \U$46109 ( \46084 , \43923 );
not \U$46110 ( \46085 , \46084 );
buf \U$46111 ( \46086 , \46085 );
buf \U$46112 ( \46087 , \46086 );
nand \U$46113 ( \46088 , \46083 , \46087 );
buf \U$46114 ( \46089 , \46088 );
buf \U$46115 ( \46090 , \46089 );
nand \U$46116 ( \46091 , \46080 , \46090 );
buf \U$46117 ( \46092 , \46091 );
xor \U$46118 ( \46093 , \46075 , \46092 );
buf \U$46119 ( \46094 , \46093 );
buf \U$46120 ( \46095 , \44413 );
not \U$46121 ( \46096 , \46095 );
buf \U$46122 ( \46097 , \44430 );
not \U$46123 ( \46098 , \46097 );
or \U$46124 ( \46099 , \46096 , \46098 );
buf \U$46125 ( \46100 , \44430 );
buf \U$46126 ( \46101 , \44413 );
or \U$46127 ( \46102 , \46100 , \46101 );
buf \U$46128 ( \46103 , \44396 );
nand \U$46129 ( \46104 , \46102 , \46103 );
buf \U$46130 ( \46105 , \46104 );
buf \U$46131 ( \46106 , \46105 );
nand \U$46132 ( \46107 , \46099 , \46106 );
buf \U$46133 ( \46108 , \46107 );
buf \U$46134 ( \46109 , \46108 );
not \U$46135 ( \46110 , \44039 );
not \U$46136 ( \46111 , \44058 );
or \U$46137 ( \46112 , \46110 , \46111 );
not \U$46138 ( \46113 , \44036 );
not \U$46139 ( \46114 , \44061 );
or \U$46140 ( \46115 , \46113 , \46114 );
nand \U$46141 ( \46116 , \46115 , \44089 );
nand \U$46142 ( \46117 , \46112 , \46116 );
buf \U$46143 ( \46118 , \46117 );
xor \U$46144 ( \46119 , \46109 , \46118 );
xor \U$46145 ( \46120 , \44451 , \44468 );
and \U$46146 ( \46121 , \46120 , \44482 );
and \U$46147 ( \46122 , \44451 , \44468 );
or \U$46148 ( \46123 , \46121 , \46122 );
buf \U$46149 ( \46124 , \46123 );
buf \U$46150 ( \46125 , \46124 );
xor \U$46151 ( \46126 , \46119 , \46125 );
buf \U$46152 ( \46127 , \46126 );
buf \U$46153 ( \46128 , \46127 );
xor \U$46154 ( \46129 , \46094 , \46128 );
buf \U$46155 ( \46130 , \44034 );
not \U$46156 ( \46131 , \46130 );
buf \U$46157 ( \46132 , \29546 );
not \U$46158 ( \46133 , \46132 );
or \U$46159 ( \46134 , \46131 , \46133 );
buf \U$46160 ( \46135 , \20243 );
buf \U$46161 ( \46136 , RIc0d8c08_47);
buf \U$46162 ( \46137 , RIc0da648_103);
xor \U$46163 ( \46138 , \46136 , \46137 );
buf \U$46164 ( \46139 , \46138 );
buf \U$46165 ( \46140 , \46139 );
nand \U$46166 ( \46141 , \46135 , \46140 );
buf \U$46167 ( \46142 , \46141 );
buf \U$46168 ( \46143 , \46142 );
nand \U$46169 ( \46144 , \46134 , \46143 );
buf \U$46170 ( \46145 , \46144 );
buf \U$46171 ( \46146 , \46145 );
buf \U$46172 ( \46147 , \44052 );
not \U$46173 ( \46148 , \46147 );
buf \U$46174 ( \46149 , \22350 );
not \U$46175 ( \46150 , \46149 );
or \U$46176 ( \46151 , \46148 , \46150 );
buf \U$46177 ( \46152 , \22356 );
buf \U$46178 ( \46153 , RIc0dacd8_117);
buf \U$46179 ( \46154 , RIc0d8578_33);
and \U$46180 ( \46155 , \46153 , \46154 );
not \U$46181 ( \46156 , \46153 );
buf \U$46182 ( \46157 , RIc0d8578_33);
not \U$46183 ( \46158 , \46157 );
buf \U$46184 ( \46159 , \46158 );
buf \U$46185 ( \46160 , \46159 );
and \U$46186 ( \46161 , \46156 , \46160 );
nor \U$46187 ( \46162 , \46155 , \46161 );
buf \U$46188 ( \46163 , \46162 );
buf \U$46189 ( \46164 , \46163 );
nand \U$46190 ( \46165 , \46152 , \46164 );
buf \U$46191 ( \46166 , \46165 );
buf \U$46192 ( \46167 , \46166 );
nand \U$46193 ( \46168 , \46151 , \46167 );
buf \U$46194 ( \46169 , \46168 );
buf \U$46195 ( \46170 , \46169 );
xor \U$46196 ( \46171 , \46146 , \46170 );
buf \U$46197 ( \46172 , RIc0dafa8_123);
buf \U$46198 ( \46173 , RIc0d82a8_27);
xor \U$46199 ( \46174 , \46172 , \46173 );
buf \U$46200 ( \46175 , \46174 );
buf \U$46201 ( \46176 , \46175 );
not \U$46202 ( \46177 , \46176 );
buf \U$46203 ( \46178 , \14278 );
not \U$46204 ( \46179 , \46178 );
or \U$46205 ( \46180 , \46177 , \46179 );
buf \U$46206 ( \46181 , \14982 );
not \U$46207 ( \46182 , \46181 );
buf \U$46208 ( \46183 , \46182 );
buf \U$46209 ( \46184 , \46183 );
buf \U$46210 ( \46185 , \44477 );
or \U$46211 ( \46186 , \46184 , \46185 );
nand \U$46212 ( \46187 , \46180 , \46186 );
buf \U$46213 ( \46188 , \46187 );
buf \U$46214 ( \46189 , \46188 );
xor \U$46215 ( \46190 , \46171 , \46189 );
buf \U$46216 ( \46191 , \46190 );
buf \U$46217 ( \46192 , \46191 );
not \U$46218 ( \46193 , \46192 );
buf \U$46219 ( \46194 , \44158 );
not \U$46220 ( \46195 , \46194 );
buf \U$46221 ( \46196 , \13569 );
not \U$46222 ( \46197 , \46196 );
or \U$46223 ( \46198 , \46195 , \46197 );
buf \U$46224 ( \46199 , \4008 );
xor \U$46225 ( \46200 , RIc0da198_93, RIc0d90b8_57);
buf \U$46226 ( \46201 , \46200 );
nand \U$46227 ( \46202 , \46199 , \46201 );
buf \U$46228 ( \46203 , \46202 );
buf \U$46229 ( \46204 , \46203 );
nand \U$46230 ( \46205 , \46198 , \46204 );
buf \U$46231 ( \46206 , \46205 );
buf \U$46232 ( \46207 , \46206 );
buf \U$46233 ( \46208 , \43874 );
not \U$46234 ( \46209 , \46208 );
buf \U$46235 ( \46210 , \46209 );
buf \U$46236 ( \46211 , \46210 );
not \U$46237 ( \46212 , \46211 );
buf \U$46238 ( \46213 , \2535 );
not \U$46239 ( \46214 , \46213 );
or \U$46240 ( \46215 , \46212 , \46214 );
buf \U$46241 ( \46216 , \714 );
buf \U$46242 ( \46217 , RIc0da0a8_91);
buf \U$46243 ( \46218 , RIc0d91a8_59);
xor \U$46244 ( \46219 , \46217 , \46218 );
buf \U$46245 ( \46220 , \46219 );
buf \U$46246 ( \46221 , \46220 );
nand \U$46247 ( \46222 , \46216 , \46221 );
buf \U$46248 ( \46223 , \46222 );
buf \U$46249 ( \46224 , \46223 );
nand \U$46250 ( \46225 , \46215 , \46224 );
buf \U$46251 ( \46226 , \46225 );
buf \U$46252 ( \46227 , \46226 );
xor \U$46253 ( \46228 , \46207 , \46227 );
buf \U$46254 ( \46229 , \44424 );
not \U$46255 ( \46230 , \46229 );
buf \U$46256 ( \46231 , \12736 );
not \U$46257 ( \46232 , \46231 );
or \U$46258 ( \46233 , \46230 , \46232 );
buf \U$46259 ( \46234 , \15653 );
buf \U$46260 ( \46235 , RIc0d8b18_45);
buf \U$46261 ( \46236 , RIc0da738_105);
xor \U$46262 ( \46237 , \46235 , \46236 );
buf \U$46263 ( \46238 , \46237 );
buf \U$46264 ( \46239 , \46238 );
nand \U$46265 ( \46240 , \46234 , \46239 );
buf \U$46266 ( \46241 , \46240 );
buf \U$46267 ( \46242 , \46241 );
nand \U$46268 ( \46243 , \46233 , \46242 );
buf \U$46269 ( \46244 , \46243 );
buf \U$46270 ( \46245 , \46244 );
xor \U$46271 ( \46246 , \46228 , \46245 );
buf \U$46272 ( \46247 , \46246 );
buf \U$46273 ( \46248 , \44461 );
not \U$46274 ( \46249 , \46248 );
buf \U$46275 ( \46250 , \25355 );
not \U$46276 ( \46251 , \46250 );
or \U$46277 ( \46252 , \46249 , \46251 );
buf \U$46278 ( \46253 , \14405 );
xor \U$46279 ( \46254 , RIc0daaf8_113, RIc0d8758_37);
buf \U$46280 ( \46255 , \46254 );
nand \U$46281 ( \46256 , \46253 , \46255 );
buf \U$46282 ( \46257 , \46256 );
buf \U$46283 ( \46258 , \46257 );
nand \U$46284 ( \46259 , \46252 , \46258 );
buf \U$46285 ( \46260 , \46259 );
buf \U$46286 ( \46261 , \43894 );
not \U$46287 ( \46262 , \46261 );
buf \U$46288 ( \46263 , \13949 );
not \U$46289 ( \46264 , \46263 );
or \U$46290 ( \46265 , \46262 , \46264 );
buf \U$46291 ( \46266 , \13953 );
buf \U$46292 ( \46267 , RIc0d8488_31);
buf \U$46293 ( \46268 , RIc0dadc8_119);
xor \U$46294 ( \46269 , \46267 , \46268 );
buf \U$46295 ( \46270 , \46269 );
buf \U$46296 ( \46271 , \46270 );
nand \U$46297 ( \46272 , \46266 , \46271 );
buf \U$46298 ( \46273 , \46272 );
buf \U$46299 ( \46274 , \46273 );
nand \U$46300 ( \46275 , \46265 , \46274 );
buf \U$46301 ( \46276 , \46275 );
xor \U$46302 ( \46277 , \46260 , \46276 );
buf \U$46303 ( \46278 , \46277 );
buf \U$46304 ( \46279 , RIc0d9ec8_87);
buf \U$46305 ( \46280 , RIc0d9400_64);
and \U$46306 ( \46281 , \46279 , \46280 );
not \U$46307 ( \46282 , \46279 );
buf \U$46308 ( \46283 , \43843 );
and \U$46309 ( \46284 , \46282 , \46283 );
nor \U$46310 ( \46285 , \46281 , \46284 );
buf \U$46311 ( \46286 , \46285 );
buf \U$46312 ( \46287 , \46286 );
not \U$46313 ( \46288 , \46287 );
buf \U$46314 ( \46289 , \2607 );
not \U$46315 ( \46290 , \46289 );
or \U$46316 ( \46291 , \46288 , \46290 );
buf \U$46317 ( \46292 , \816 );
xor \U$46318 ( \46293 , RIc0d9ec8_87, RIc0d9388_63);
buf \U$46319 ( \46294 , \46293 );
nand \U$46320 ( \46295 , \46292 , \46294 );
buf \U$46321 ( \46296 , \46295 );
buf \U$46322 ( \46297 , \46296 );
nand \U$46323 ( \46298 , \46291 , \46297 );
buf \U$46324 ( \46299 , \46298 );
buf \U$46325 ( \46300 , \46299 );
xnor \U$46326 ( \46301 , \46278 , \46300 );
buf \U$46327 ( \46302 , \46301 );
xor \U$46328 ( \46303 , \46247 , \46302 );
buf \U$46329 ( \46304 , \46303 );
not \U$46330 ( \46305 , \46304 );
or \U$46331 ( \46306 , \46193 , \46305 );
buf \U$46332 ( \46307 , \46303 );
buf \U$46333 ( \46308 , \46191 );
or \U$46334 ( \46309 , \46307 , \46308 );
nand \U$46335 ( \46310 , \46306 , \46309 );
buf \U$46336 ( \46311 , \46310 );
buf \U$46337 ( \46312 , \46311 );
xor \U$46338 ( \46313 , \46129 , \46312 );
buf \U$46339 ( \46314 , \46313 );
buf \U$46340 ( \46315 , \46314 );
xor \U$46341 ( \46316 , \46046 , \46315 );
buf \U$46342 ( \46317 , \46316 );
buf \U$46343 ( \46318 , \46317 );
xor \U$46344 ( \46319 , \45979 , \46318 );
buf \U$46345 ( \46320 , \45993 );
buf \U$46346 ( \46321 , \46000 );
xor \U$46347 ( \46322 , \46320 , \46321 );
buf \U$46348 ( \46323 , \46016 );
xor \U$46349 ( \46324 , \46322 , \46323 );
buf \U$46350 ( \46325 , \46324 );
buf \U$46351 ( \46326 , \46325 );
xor \U$46352 ( \46327 , \46029 , \46033 );
xor \U$46353 ( \46328 , \46327 , \46040 );
buf \U$46354 ( \46329 , \46328 );
buf \U$46355 ( \46330 , \46329 );
xor \U$46356 ( \46331 , \46326 , \46330 );
xor \U$46357 ( \46332 , \45017 , \45042 );
xor \U$46358 ( \46333 , \46332 , \45457 );
buf \U$46359 ( \46334 , \46333 );
buf \U$46360 ( \46335 , \46334 );
and \U$46361 ( \46336 , \46331 , \46335 );
and \U$46362 ( \46337 , \46326 , \46330 );
or \U$46363 ( \46338 , \46336 , \46337 );
buf \U$46364 ( \46339 , \46338 );
buf \U$46365 ( \46340 , \46339 );
and \U$46366 ( \46341 , \46319 , \46340 );
and \U$46367 ( \46342 , \45979 , \46318 );
or \U$46368 ( \46343 , \46341 , \46342 );
buf \U$46369 ( \46344 , \46343 );
buf \U$46370 ( \46345 , \46344 );
xor \U$46371 ( \46346 , \45467 , \46345 );
xor \U$46372 ( \46347 , \46023 , \46045 );
and \U$46373 ( \46348 , \46347 , \46315 );
and \U$46374 ( \46349 , \46023 , \46045 );
or \U$46375 ( \46350 , \46348 , \46349 );
buf \U$46376 ( \46351 , \46350 );
buf \U$46377 ( \46352 , \46351 );
buf \U$46378 ( \46353 , \43967 );
not \U$46379 ( \46354 , \46353 );
buf \U$46380 ( \46355 , \44171 );
not \U$46381 ( \46356 , \46355 );
or \U$46382 ( \46357 , \46354 , \46356 );
buf \U$46383 ( \46358 , \44171 );
buf \U$46384 ( \46359 , \43967 );
or \U$46385 ( \46360 , \46358 , \46359 );
buf \U$46386 ( \46361 , \44373 );
nand \U$46387 ( \46362 , \46360 , \46361 );
buf \U$46388 ( \46363 , \46362 );
buf \U$46389 ( \46364 , \46363 );
nand \U$46390 ( \46365 , \46357 , \46364 );
buf \U$46391 ( \46366 , \46365 );
buf \U$46392 ( \46367 , \46366 );
xor \U$46393 ( \46368 , \46094 , \46128 );
and \U$46394 ( \46369 , \46368 , \46312 );
and \U$46395 ( \46370 , \46094 , \46128 );
or \U$46396 ( \46371 , \46369 , \46370 );
buf \U$46397 ( \46372 , \46371 );
buf \U$46398 ( \46373 , \46372 );
xor \U$46399 ( \46374 , \46367 , \46373 );
buf \U$46400 ( \46375 , \44801 );
not \U$46401 ( \46376 , \46375 );
buf \U$46402 ( \46377 , \14210 );
not \U$46403 ( \46378 , \46377 );
or \U$46404 ( \46379 , \46376 , \46378 );
buf \U$46405 ( \46380 , \20211 );
buf \U$46406 ( \46381 , RIc0da918_109);
buf \U$46407 ( \46382 , RIc0d88c0_40);
xor \U$46408 ( \46383 , \46381 , \46382 );
buf \U$46409 ( \46384 , \46383 );
buf \U$46410 ( \46385 , \46384 );
nand \U$46411 ( \46386 , \46380 , \46385 );
buf \U$46412 ( \46387 , \46386 );
buf \U$46413 ( \46388 , \46387 );
nand \U$46414 ( \46389 , \46379 , \46388 );
buf \U$46415 ( \46390 , \46389 );
buf \U$46416 ( \46391 , \46390 );
and \U$46417 ( \46392 , \44854 , \44871 );
buf \U$46418 ( \46393 , \46392 );
buf \U$46419 ( \46394 , \46393 );
xor \U$46420 ( \46395 , \46391 , \46394 );
buf \U$46421 ( \46396 , \44736 );
buf \U$46422 ( \46397 , \44720 );
or \U$46423 ( \46398 , \46396 , \46397 );
buf \U$46424 ( \46399 , \44707 );
nand \U$46425 ( \46400 , \46398 , \46399 );
buf \U$46426 ( \46401 , \46400 );
buf \U$46427 ( \46402 , \46401 );
buf \U$46428 ( \46403 , \44720 );
buf \U$46429 ( \46404 , \44736 );
nand \U$46430 ( \46405 , \46403 , \46404 );
buf \U$46431 ( \46406 , \46405 );
buf \U$46432 ( \46407 , \46406 );
nand \U$46433 ( \46408 , \46402 , \46407 );
buf \U$46434 ( \46409 , \46408 );
buf \U$46435 ( \46410 , \46409 );
xor \U$46436 ( \46411 , \46395 , \46410 );
buf \U$46437 ( \46412 , \46411 );
buf \U$46438 ( \46413 , \46412 );
xor \U$46439 ( \46414 , \44638 , \44690 );
and \U$46440 ( \46415 , \46414 , \44739 );
and \U$46441 ( \46416 , \44638 , \44690 );
or \U$46442 ( \46417 , \46415 , \46416 );
buf \U$46443 ( \46418 , \46417 );
buf \U$46444 ( \46419 , \46418 );
xor \U$46445 ( \46420 , \46413 , \46419 );
buf \U$46446 ( \46421 , \46139 );
not \U$46447 ( \46422 , \46421 );
buf \U$46448 ( \46423 , \29546 );
not \U$46449 ( \46424 , \46423 );
or \U$46450 ( \46425 , \46422 , \46424 );
buf \U$46451 ( \46426 , RIc0da648_103);
buf \U$46452 ( \46427 , RIc0d8b90_46);
xnor \U$46453 ( \46428 , \46426 , \46427 );
buf \U$46454 ( \46429 , \46428 );
buf \U$46455 ( \46430 , \46429 );
not \U$46456 ( \46431 , \46430 );
buf \U$46457 ( \46432 , \16584 );
nand \U$46458 ( \46433 , \46431 , \46432 );
buf \U$46459 ( \46434 , \46433 );
buf \U$46460 ( \46435 , \46434 );
nand \U$46461 ( \46436 , \46425 , \46435 );
buf \U$46462 ( \46437 , \46436 );
buf \U$46463 ( \46438 , \46437 );
buf \U$46464 ( \46439 , \46163 );
not \U$46465 ( \46440 , \46439 );
buf \U$46466 ( \46441 , \13146 );
not \U$46467 ( \46442 , \46441 );
or \U$46468 ( \46443 , \46440 , \46442 );
buf \U$46469 ( \46444 , \12937 );
buf \U$46470 ( \46445 , RIc0d8500_32);
buf \U$46471 ( \46446 , RIc0dacd8_117);
xor \U$46472 ( \46447 , \46445 , \46446 );
buf \U$46473 ( \46448 , \46447 );
buf \U$46474 ( \46449 , \46448 );
nand \U$46475 ( \46450 , \46444 , \46449 );
buf \U$46476 ( \46451 , \46450 );
buf \U$46477 ( \46452 , \46451 );
nand \U$46478 ( \46453 , \46443 , \46452 );
buf \U$46479 ( \46454 , \46453 );
buf \U$46480 ( \46455 , \46454 );
xor \U$46481 ( \46456 , \46438 , \46455 );
buf \U$46482 ( \46457 , \13461 );
not \U$46483 ( \46458 , \46457 );
buf \U$46484 ( \46459 , \46458 );
buf \U$46485 ( \46460 , \46459 );
buf \U$46486 ( \46461 , \44820 );
or \U$46487 ( \46462 , \46460 , \46461 );
buf \U$46488 ( \46463 , \22744 );
buf \U$46489 ( \46464 , RIc0d8140_24);
buf \U$46490 ( \46465 , RIc0db098_125);
xor \U$46491 ( \46466 , \46464 , \46465 );
buf \U$46492 ( \46467 , \46466 );
buf \U$46493 ( \46468 , \46467 );
not \U$46494 ( \46469 , \46468 );
buf \U$46495 ( \46470 , \46469 );
buf \U$46496 ( \46471 , \46470 );
or \U$46497 ( \46472 , \46463 , \46471 );
nand \U$46498 ( \46473 , \46462 , \46472 );
buf \U$46499 ( \46474 , \46473 );
buf \U$46500 ( \46475 , \46474 );
xor \U$46501 ( \46476 , \46456 , \46475 );
buf \U$46502 ( \46477 , \46476 );
buf \U$46503 ( \46478 , \46477 );
not \U$46504 ( \46479 , \46478 );
buf \U$46505 ( \46480 , \46479 );
buf \U$46506 ( \46481 , \46480 );
not \U$46507 ( \46482 , \46481 );
xor \U$46508 ( \46483 , \44653 , \44667 );
and \U$46509 ( \46484 , \46483 , \44687 );
and \U$46510 ( \46485 , \44653 , \44667 );
or \U$46511 ( \46486 , \46484 , \46485 );
buf \U$46512 ( \46487 , \46486 );
buf \U$46513 ( \46488 , \46487 );
not \U$46514 ( \46489 , \46488 );
buf \U$46515 ( \46490 , \46299 );
not \U$46516 ( \46491 , \46490 );
buf \U$46517 ( \46492 , \46260 );
not \U$46518 ( \46493 , \46492 );
or \U$46519 ( \46494 , \46491 , \46493 );
buf \U$46520 ( \46495 , \46260 );
buf \U$46521 ( \46496 , \46299 );
or \U$46522 ( \46497 , \46495 , \46496 );
buf \U$46523 ( \46498 , \46276 );
nand \U$46524 ( \46499 , \46497 , \46498 );
buf \U$46525 ( \46500 , \46499 );
buf \U$46526 ( \46501 , \46500 );
nand \U$46527 ( \46502 , \46494 , \46501 );
buf \U$46528 ( \46503 , \46502 );
buf \U$46529 ( \46504 , \46503 );
not \U$46530 ( \46505 , \46504 );
buf \U$46531 ( \46506 , \46505 );
buf \U$46532 ( \46507 , \46506 );
not \U$46533 ( \46508 , \46507 );
or \U$46534 ( \46509 , \46489 , \46508 );
buf \U$46535 ( \46510 , \46506 );
buf \U$46536 ( \46511 , \46487 );
or \U$46537 ( \46512 , \46510 , \46511 );
nand \U$46538 ( \46513 , \46509 , \46512 );
buf \U$46539 ( \46514 , \46513 );
buf \U$46540 ( \46515 , \46514 );
not \U$46541 ( \46516 , \46515 );
or \U$46542 ( \46517 , \46482 , \46516 );
buf \U$46543 ( \46518 , \46514 );
buf \U$46544 ( \46519 , \46480 );
or \U$46545 ( \46520 , \46518 , \46519 );
nand \U$46546 ( \46521 , \46517 , \46520 );
buf \U$46547 ( \46522 , \46521 );
buf \U$46548 ( \46523 , \46522 );
xor \U$46549 ( \46524 , \46420 , \46523 );
buf \U$46550 ( \46525 , \46524 );
buf \U$46551 ( \46526 , \46525 );
xor \U$46552 ( \46527 , \46374 , \46526 );
buf \U$46553 ( \46528 , \46527 );
buf \U$46554 ( \46529 , \46528 );
xor \U$46555 ( \46530 , \46352 , \46529 );
xor \U$46556 ( \46531 , \44632 , \44742 );
and \U$46557 ( \46532 , \46531 , \45009 );
and \U$46558 ( \46533 , \44632 , \44742 );
or \U$46559 ( \46534 , \46532 , \46533 );
buf \U$46560 ( \46535 , \46534 );
buf \U$46561 ( \46536 , \46535 );
buf \U$46562 ( \46537 , \46191 );
not \U$46563 ( \46538 , \46537 );
buf \U$46564 ( \46539 , \46247 );
not \U$46565 ( \46540 , \46539 );
or \U$46566 ( \46541 , \46538 , \46540 );
buf \U$46567 ( \46542 , \46247 );
buf \U$46568 ( \46543 , \46191 );
or \U$46569 ( \46544 , \46542 , \46543 );
buf \U$46570 ( \46545 , \46302 );
not \U$46571 ( \46546 , \46545 );
buf \U$46572 ( \46547 , \46546 );
buf \U$46573 ( \46548 , \46547 );
nand \U$46574 ( \46549 , \46544 , \46548 );
buf \U$46575 ( \46550 , \46549 );
buf \U$46576 ( \46551 , \46550 );
nand \U$46577 ( \46552 , \46541 , \46551 );
buf \U$46578 ( \46553 , \46552 );
buf \U$46579 ( \46554 , \46553 );
not \U$46580 ( \46555 , \46554 );
buf \U$46581 ( \46556 , \44769 );
buf \U$46582 ( \46557 , \44786 );
or \U$46583 ( \46558 , \46556 , \46557 );
buf \U$46584 ( \46559 , \44756 );
nand \U$46585 ( \46560 , \46558 , \46559 );
buf \U$46586 ( \46561 , \46560 );
buf \U$46587 ( \46562 , \46561 );
buf \U$46588 ( \46563 , \44786 );
buf \U$46589 ( \46564 , \44769 );
nand \U$46590 ( \46565 , \46563 , \46564 );
buf \U$46591 ( \46566 , \46565 );
buf \U$46592 ( \46567 , \46566 );
nand \U$46593 ( \46568 , \46562 , \46567 );
buf \U$46594 ( \46569 , \46568 );
buf \U$46595 ( \46570 , \46569 );
xor \U$46596 ( \46571 , \46207 , \46227 );
and \U$46597 ( \46572 , \46571 , \46245 );
and \U$46598 ( \46573 , \46207 , \46227 );
or \U$46599 ( \46574 , \46572 , \46573 );
buf \U$46600 ( \46575 , \46574 );
buf \U$46601 ( \46576 , \46575 );
xor \U$46602 ( \46577 , \46570 , \46576 );
xor \U$46603 ( \46578 , \46146 , \46170 );
and \U$46604 ( \46579 , \46578 , \46189 );
and \U$46605 ( \46580 , \46146 , \46170 );
or \U$46606 ( \46581 , \46579 , \46580 );
buf \U$46607 ( \46582 , \46581 );
buf \U$46608 ( \46583 , \46582 );
xor \U$46609 ( \46584 , \46577 , \46583 );
buf \U$46610 ( \46585 , \46584 );
buf \U$46611 ( \46586 , \46585 );
not \U$46612 ( \46587 , \46586 );
buf \U$46613 ( \46588 , \46587 );
buf \U$46614 ( \46589 , \46588 );
not \U$46615 ( \46590 , \46589 );
or \U$46616 ( \46591 , \46555 , \46590 );
buf \U$46617 ( \46592 , \46585 );
buf \U$46618 ( \46593 , \46553 );
not \U$46619 ( \46594 , \46593 );
buf \U$46620 ( \46595 , \46594 );
buf \U$46621 ( \46596 , \46595 );
nand \U$46622 ( \46597 , \46592 , \46596 );
buf \U$46623 ( \46598 , \46597 );
buf \U$46624 ( \46599 , \46598 );
nand \U$46625 ( \46600 , \46591 , \46599 );
buf \U$46626 ( \46601 , \46600 );
buf \U$46627 ( \46602 , \46601 );
buf \U$46628 ( \46603 , \46220 );
not \U$46629 ( \46604 , \46603 );
buf \U$46630 ( \46605 , \2726 );
not \U$46631 ( \46606 , \46605 );
or \U$46632 ( \46607 , \46604 , \46606 );
buf \U$46633 ( \46608 , \533 );
buf \U$46634 ( \46609 , RIc0da0a8_91);
buf \U$46635 ( \46610 , RIc0d9130_58);
xor \U$46636 ( \46611 , \46609 , \46610 );
buf \U$46637 ( \46612 , \46611 );
buf \U$46638 ( \46613 , \46612 );
nand \U$46639 ( \46614 , \46608 , \46613 );
buf \U$46640 ( \46615 , \46614 );
buf \U$46641 ( \46616 , \46615 );
nand \U$46642 ( \46617 , \46607 , \46616 );
buf \U$46643 ( \46618 , \46617 );
buf \U$46644 ( \46619 , \46618 );
buf \U$46645 ( \46620 , \46238 );
not \U$46646 ( \46621 , \46620 );
buf \U$46647 ( \46622 , \15644 );
not \U$46648 ( \46623 , \46622 );
or \U$46649 ( \46624 , \46621 , \46623 );
buf \U$46650 ( \46625 , \21880 );
buf \U$46651 ( \46626 , RIc0da738_105);
buf \U$46652 ( \46627 , RIc0d8aa0_44);
xor \U$46653 ( \46628 , \46626 , \46627 );
buf \U$46654 ( \46629 , \46628 );
buf \U$46655 ( \46630 , \46629 );
nand \U$46656 ( \46631 , \46625 , \46630 );
buf \U$46657 ( \46632 , \46631 );
buf \U$46658 ( \46633 , \46632 );
nand \U$46659 ( \46634 , \46624 , \46633 );
buf \U$46660 ( \46635 , \46634 );
buf \U$46661 ( \46636 , \46635 );
xor \U$46662 ( \46637 , \46619 , \46636 );
buf \U$46663 ( \46638 , \44714 );
not \U$46664 ( \46639 , \46638 );
buf \U$46665 ( \46640 , \28794 );
not \U$46666 ( \46641 , \46640 );
or \U$46667 ( \46642 , \46639 , \46641 );
buf \U$46668 ( \46643 , \16071 );
buf \U$46669 ( \46644 , RIc0d89b0_42);
buf \U$46670 ( \46645 , RIc0da828_107);
xor \U$46671 ( \46646 , \46644 , \46645 );
buf \U$46672 ( \46647 , \46646 );
buf \U$46673 ( \46648 , \46647 );
nand \U$46674 ( \46649 , \46643 , \46648 );
buf \U$46675 ( \46650 , \46649 );
buf \U$46676 ( \46651 , \46650 );
nand \U$46677 ( \46652 , \46642 , \46651 );
buf \U$46678 ( \46653 , \46652 );
buf \U$46679 ( \46654 , \46653 );
xor \U$46680 ( \46655 , \46637 , \46654 );
buf \U$46681 ( \46656 , \46655 );
buf \U$46682 ( \46657 , \46656 );
buf \U$46683 ( \46658 , \44780 );
not \U$46684 ( \46659 , \46658 );
buf \U$46685 ( \46660 , \13092 );
not \U$46686 ( \46661 , \46660 );
or \U$46687 ( \46662 , \46659 , \46661 );
buf \U$46688 ( \46663 , \2070 );
buf \U$46689 ( \46664 , RIc0da378_97);
buf \U$46690 ( \46665 , RIc0d8e60_52);
xor \U$46691 ( \46666 , \46664 , \46665 );
buf \U$46692 ( \46667 , \46666 );
buf \U$46693 ( \46668 , \46667 );
nand \U$46694 ( \46669 , \46663 , \46668 );
buf \U$46695 ( \46670 , \46669 );
buf \U$46696 ( \46671 , \46670 );
nand \U$46697 ( \46672 , \46662 , \46671 );
buf \U$46698 ( \46673 , \46672 );
buf \U$46699 ( \46674 , \44750 );
not \U$46700 ( \46675 , \46674 );
buf \U$46701 ( \46676 , \16744 );
not \U$46702 ( \46677 , \46676 );
or \U$46703 ( \46678 , \46675 , \46677 );
buf \U$46704 ( \46679 , \2476 );
buf \U$46705 ( \46680 , RIc0da468_99);
buf \U$46706 ( \46681 , RIc0d8d70_50);
xor \U$46707 ( \46682 , \46680 , \46681 );
buf \U$46708 ( \46683 , \46682 );
buf \U$46709 ( \46684 , \46683 );
nand \U$46710 ( \46685 , \46679 , \46684 );
buf \U$46711 ( \46686 , \46685 );
buf \U$46712 ( \46687 , \46686 );
nand \U$46713 ( \46688 , \46678 , \46687 );
buf \U$46714 ( \46689 , \46688 );
xor \U$46715 ( \46690 , \46673 , \46689 );
buf \U$46716 ( \46691 , \46175 );
not \U$46717 ( \46692 , \46691 );
buf \U$46718 ( \46693 , \14982 );
not \U$46719 ( \46694 , \46693 );
or \U$46720 ( \46695 , \46692 , \46694 );
buf \U$46721 ( \46696 , \14278 );
buf \U$46722 ( \46697 , RIc0dafa8_123);
buf \U$46723 ( \46698 , RIc0d8230_26);
xor \U$46724 ( \46699 , \46697 , \46698 );
buf \U$46725 ( \46700 , \46699 );
buf \U$46726 ( \46701 , \46700 );
nand \U$46727 ( \46702 , \46696 , \46701 );
buf \U$46728 ( \46703 , \46702 );
buf \U$46729 ( \46704 , \46703 );
nand \U$46730 ( \46705 , \46695 , \46704 );
buf \U$46731 ( \46706 , \46705 );
xor \U$46732 ( \46707 , \46690 , \46706 );
buf \U$46733 ( \46708 , \46707 );
xor \U$46734 ( \46709 , \46657 , \46708 );
buf \U$46735 ( \46710 , \46293 );
not \U$46736 ( \46711 , \46710 );
buf \U$46737 ( \46712 , \1765 );
not \U$46738 ( \46713 , \46712 );
or \U$46739 ( \46714 , \46711 , \46713 );
buf \U$46740 ( \46715 , \816 );
buf \U$46741 ( \46716 , RIc0d9ec8_87);
buf \U$46742 ( \46717 , RIc0d9310_62);
xor \U$46743 ( \46718 , \46716 , \46717 );
buf \U$46744 ( \46719 , \46718 );
buf \U$46745 ( \46720 , \46719 );
nand \U$46746 ( \46721 , \46715 , \46720 );
buf \U$46747 ( \46722 , \46721 );
buf \U$46748 ( \46723 , \46722 );
nand \U$46749 ( \46724 , \46714 , \46723 );
buf \U$46750 ( \46725 , \46724 );
buf \U$46751 ( \46726 , \46725 );
buf \U$46752 ( \46727 , \46200 );
not \U$46753 ( \46728 , \46727 );
buf \U$46754 ( \46729 , \1901 );
not \U$46755 ( \46730 , \46729 );
or \U$46756 ( \46731 , \46728 , \46730 );
buf \U$46757 ( \46732 , \4008 );
buf \U$46758 ( \46733 , RIc0da198_93);
buf \U$46759 ( \46734 , RIc0d9040_56);
xor \U$46760 ( \46735 , \46733 , \46734 );
buf \U$46761 ( \46736 , \46735 );
buf \U$46762 ( \46737 , \46736 );
nand \U$46763 ( \46738 , \46732 , \46737 );
buf \U$46764 ( \46739 , \46738 );
buf \U$46765 ( \46740 , \46739 );
nand \U$46766 ( \46741 , \46731 , \46740 );
buf \U$46767 ( \46742 , \46741 );
buf \U$46768 ( \46743 , \46742 );
xor \U$46769 ( \46744 , \46726 , \46743 );
buf \U$46770 ( \46745 , \46270 );
not \U$46771 ( \46746 , \46745 );
buf \U$46772 ( \46747 , \14569 );
not \U$46773 ( \46748 , \46747 );
or \U$46774 ( \46749 , \46746 , \46748 );
buf \U$46775 ( \46750 , \13005 );
buf \U$46776 ( \46751 , RIc0dadc8_119);
buf \U$46777 ( \46752 , RIc0d8410_30);
xor \U$46778 ( \46753 , \46751 , \46752 );
buf \U$46779 ( \46754 , \46753 );
buf \U$46780 ( \46755 , \46754 );
nand \U$46781 ( \46756 , \46750 , \46755 );
buf \U$46782 ( \46757 , \46756 );
buf \U$46783 ( \46758 , \46757 );
nand \U$46784 ( \46759 , \46749 , \46758 );
buf \U$46785 ( \46760 , \46759 );
buf \U$46786 ( \46761 , \46760 );
xor \U$46787 ( \46762 , \46744 , \46761 );
buf \U$46788 ( \46763 , \46762 );
buf \U$46789 ( \46764 , \46763 );
xor \U$46790 ( \46765 , \46709 , \46764 );
buf \U$46791 ( \46766 , \46765 );
buf \U$46792 ( \46767 , \46766 );
xor \U$46793 ( \46768 , \46602 , \46767 );
buf \U$46794 ( \46769 , \46768 );
buf \U$46795 ( \46770 , \46769 );
xor \U$46796 ( \46771 , \46536 , \46770 );
buf \U$46797 ( \46772 , \2960 );
buf \U$46798 ( \46773 , RIc0d9400_64);
and \U$46799 ( \46774 , \46772 , \46773 );
buf \U$46800 ( \46775 , \46774 );
buf \U$46801 ( \46776 , \46775 );
buf \U$46802 ( \46777 , \44864 );
not \U$46803 ( \46778 , \46777 );
buf \U$46804 ( \46779 , \3384 );
not \U$46805 ( \46780 , \46779 );
or \U$46806 ( \46781 , \46778 , \46780 );
buf \U$46807 ( \46782 , \16477 );
xor \U$46808 ( \46783 , RIc0d9fb8_89, RIc0d9220_60);
buf \U$46809 ( \46784 , \46783 );
nand \U$46810 ( \46785 , \46782 , \46784 );
buf \U$46811 ( \46786 , \46785 );
buf \U$46812 ( \46787 , \46786 );
nand \U$46813 ( \46788 , \46781 , \46787 );
buf \U$46814 ( \46789 , \46788 );
buf \U$46815 ( \46790 , \46789 );
xor \U$46816 ( \46791 , \46776 , \46790 );
buf \U$46817 ( \46792 , \46254 );
not \U$46818 ( \46793 , \46792 );
buf \U$46819 ( \46794 , \33224 );
not \U$46820 ( \46795 , \46794 );
or \U$46821 ( \46796 , \46793 , \46795 );
buf \U$46822 ( \46797 , \14405 );
xor \U$46823 ( \46798 , RIc0daaf8_113, RIc0d86e0_36);
buf \U$46824 ( \46799 , \46798 );
nand \U$46825 ( \46800 , \46797 , \46799 );
buf \U$46826 ( \46801 , \46800 );
buf \U$46827 ( \46802 , \46801 );
nand \U$46828 ( \46803 , \46796 , \46802 );
buf \U$46829 ( \46804 , \46803 );
buf \U$46830 ( \46805 , \46804 );
xor \U$46831 ( \46806 , \46791 , \46805 );
buf \U$46832 ( \46807 , \46806 );
buf \U$46833 ( \46808 , \46807 );
xor \U$46834 ( \46809 , RIc0db188_127, RIc0d8050_22);
not \U$46835 ( \46810 , \46809 );
not \U$46836 ( \46811 , RIc0db200_128);
or \U$46837 ( \46812 , \46810 , \46811 );
buf \U$46838 ( \46813 , \44639 );
not \U$46839 ( \46814 , \46813 );
or \U$46840 ( \46815 , \46814 , \44648 );
nand \U$46841 ( \46816 , \46812 , \46815 );
buf \U$46842 ( \46817 , \46816 );
buf \U$46843 ( \46818 , \44763 );
not \U$46844 ( \46819 , \46818 );
buf \U$46845 ( \46820 , \14346 );
not \U$46846 ( \46821 , \46820 );
or \U$46847 ( \46822 , \46819 , \46821 );
buf \U$46848 ( \46823 , \14353 );
xor \U$46849 ( \46824 , RIc0daa08_111, RIc0d87d0_38);
buf \U$46850 ( \46825 , \46824 );
nand \U$46851 ( \46826 , \46823 , \46825 );
buf \U$46852 ( \46827 , \46826 );
buf \U$46853 ( \46828 , \46827 );
nand \U$46854 ( \46829 , \46822 , \46828 );
buf \U$46855 ( \46830 , \46829 );
buf \U$46856 ( \46831 , \46830 );
xor \U$46857 ( \46832 , \46817 , \46831 );
buf \U$46858 ( \46833 , \45548 );
buf \U$46859 ( \46834 , \44660 );
not \U$46860 ( \46835 , \46834 );
buf \U$46861 ( \46836 , \46835 );
buf \U$46862 ( \46837 , \46836 );
or \U$46863 ( \46838 , \46833 , \46837 );
buf \U$46864 ( \46839 , \27558 );
buf \U$46865 ( \46840 , RIc0d8320_28);
buf \U$46866 ( \46841 , RIc0daeb8_121);
xnor \U$46867 ( \46842 , \46840 , \46841 );
buf \U$46868 ( \46843 , \46842 );
buf \U$46869 ( \46844 , \46843 );
or \U$46870 ( \46845 , \46839 , \46844 );
nand \U$46871 ( \46846 , \46838 , \46845 );
buf \U$46872 ( \46847 , \46846 );
buf \U$46873 ( \46848 , \46847 );
xor \U$46874 ( \46849 , \46832 , \46848 );
buf \U$46875 ( \46850 , \46849 );
buf \U$46876 ( \46851 , \46850 );
xor \U$46877 ( \46852 , \46808 , \46851 );
buf \U$46878 ( \46853 , \44701 );
not \U$46879 ( \46854 , \46853 );
buf \U$46880 ( \46855 , \22631 );
not \U$46881 ( \46856 , \46855 );
or \U$46882 ( \46857 , \46854 , \46856 );
buf \U$46883 ( \46858 , \12839 );
buf \U$46884 ( \46859 , RIc0da558_101);
buf \U$46885 ( \46860 , RIc0d8c80_48);
xor \U$46886 ( \46861 , \46859 , \46860 );
buf \U$46887 ( \46862 , \46861 );
buf \U$46888 ( \46863 , \46862 );
nand \U$46889 ( \46864 , \46858 , \46863 );
buf \U$46890 ( \46865 , \46864 );
buf \U$46891 ( \46866 , \46865 );
nand \U$46892 ( \46867 , \46857 , \46866 );
buf \U$46893 ( \46868 , \46867 );
buf \U$46894 ( \46869 , \44730 );
not \U$46895 ( \46870 , \46869 );
buf \U$46896 ( \46871 , \22595 );
not \U$46897 ( \46872 , \46871 );
buf \U$46898 ( \46873 , \46872 );
buf \U$46899 ( \46874 , \46873 );
not \U$46900 ( \46875 , \46874 );
or \U$46901 ( \46876 , \46870 , \46875 );
buf \U$46902 ( \46877 , RIc0dabe8_115);
buf \U$46903 ( \46878 , RIc0d85f0_34);
xnor \U$46904 ( \46879 , \46877 , \46878 );
buf \U$46905 ( \46880 , \46879 );
buf \U$46906 ( \46881 , \46880 );
not \U$46907 ( \46882 , \46881 );
buf \U$46908 ( \46883 , \12303 );
nand \U$46909 ( \46884 , \46882 , \46883 );
buf \U$46910 ( \46885 , \46884 );
buf \U$46911 ( \46886 , \46885 );
nand \U$46912 ( \46887 , \46876 , \46886 );
buf \U$46913 ( \46888 , \46887 );
xor \U$46914 ( \46889 , \46868 , \46888 );
buf \U$46915 ( \46890 , \44679 );
not \U$46916 ( \46891 , \46890 );
buf \U$46917 ( \46892 , \27591 );
not \U$46918 ( \46893 , \46892 );
or \U$46919 ( \46894 , \46891 , \46893 );
buf \U$46920 ( \46895 , \344 );
buf \U$46921 ( \46896 , RIc0da288_95);
buf \U$46922 ( \46897 , RIc0d8f50_54);
xor \U$46923 ( \46898 , \46896 , \46897 );
buf \U$46924 ( \46899 , \46898 );
buf \U$46925 ( \46900 , \46899 );
nand \U$46926 ( \46901 , \46895 , \46900 );
buf \U$46927 ( \46902 , \46901 );
buf \U$46928 ( \46903 , \46902 );
nand \U$46929 ( \46904 , \46894 , \46903 );
buf \U$46930 ( \46905 , \46904 );
xor \U$46931 ( \46906 , \46889 , \46905 );
buf \U$46932 ( \46907 , \46906 );
xor \U$46933 ( \46908 , \46852 , \46907 );
buf \U$46934 ( \46909 , \46908 );
buf \U$46935 ( \46910 , \46909 );
xor \U$46936 ( \46911 , \44788 , \44875 );
and \U$46937 ( \46912 , \46911 , \45006 );
and \U$46938 ( \46913 , \44788 , \44875 );
or \U$46939 ( \46914 , \46912 , \46913 );
buf \U$46940 ( \46915 , \46914 );
buf \U$46941 ( \46916 , \46915 );
xor \U$46942 ( \46917 , \46910 , \46916 );
buf \U$46943 ( \46918 , \44828 );
not \U$46944 ( \46919 , \46918 );
buf \U$46945 ( \46920 , \44807 );
not \U$46946 ( \46921 , \46920 );
or \U$46947 ( \46922 , \46919 , \46921 );
buf \U$46948 ( \46923 , \44873 );
buf \U$46949 ( \46924 , \44807 );
not \U$46950 ( \46925 , \46924 );
buf \U$46951 ( \46926 , \44834 );
nand \U$46952 ( \46927 , \46925 , \46926 );
buf \U$46953 ( \46928 , \46927 );
buf \U$46954 ( \46929 , \46928 );
nand \U$46955 ( \46930 , \46923 , \46929 );
buf \U$46956 ( \46931 , \46930 );
buf \U$46957 ( \46932 , \46931 );
nand \U$46958 ( \46933 , \46922 , \46932 );
buf \U$46959 ( \46934 , \46933 );
buf \U$46960 ( \46935 , \46934 );
buf \U$46961 ( \46936 , \46060 );
buf \U$46962 ( \46937 , \46074 );
or \U$46963 ( \46938 , \46936 , \46937 );
buf \U$46964 ( \46939 , \46092 );
nand \U$46965 ( \46940 , \46938 , \46939 );
buf \U$46966 ( \46941 , \46940 );
buf \U$46967 ( \46942 , \46941 );
buf \U$46968 ( \46943 , \46060 );
buf \U$46969 ( \46944 , \46074 );
nand \U$46970 ( \46945 , \46943 , \46944 );
buf \U$46971 ( \46946 , \46945 );
buf \U$46972 ( \46947 , \46946 );
nand \U$46973 ( \46948 , \46942 , \46947 );
buf \U$46974 ( \46949 , \46948 );
buf \U$46975 ( \46950 , \46949 );
xor \U$46976 ( \46951 , \46935 , \46950 );
xor \U$46977 ( \46952 , \46109 , \46118 );
and \U$46978 ( \46953 , \46952 , \46125 );
and \U$46979 ( \46954 , \46109 , \46118 );
or \U$46980 ( \46955 , \46953 , \46954 );
buf \U$46981 ( \46956 , \46955 );
buf \U$46982 ( \46957 , \46956 );
xor \U$46983 ( \46958 , \46951 , \46957 );
buf \U$46984 ( \46959 , \46958 );
buf \U$46985 ( \46960 , \46959 );
xor \U$46986 ( \46961 , \46917 , \46960 );
buf \U$46987 ( \46962 , \46961 );
buf \U$46988 ( \46963 , \46962 );
xor \U$46989 ( \46964 , \46771 , \46963 );
buf \U$46990 ( \46965 , \46964 );
buf \U$46991 ( \46966 , \46965 );
xor \U$46992 ( \46967 , \46530 , \46966 );
buf \U$46993 ( \46968 , \46967 );
buf \U$46994 ( \46969 , \46968 );
xor \U$46995 ( \46970 , \46346 , \46969 );
buf \U$46996 ( \46971 , \46970 );
buf \U$46997 ( \46972 , \46971 );
xor \U$46998 ( \46973 , \45979 , \46318 );
xor \U$46999 ( \46974 , \46973 , \46340 );
buf \U$47000 ( \46975 , \46974 );
buf \U$47001 ( \46976 , \46975 );
xor \U$47002 ( \46977 , \44375 , \45012 );
xor \U$47003 ( \46978 , \46977 , \45462 );
buf \U$47004 ( \46979 , \46978 );
buf \U$47005 ( \46980 , \46979 );
or \U$47006 ( \46981 , \46976 , \46980 );
xor \U$47007 ( \46982 , \45894 , \45908 );
xor \U$47008 ( \46983 , \46982 , \45945 );
buf \U$47009 ( \46984 , \46983 );
buf \U$47010 ( \46985 , \46984 );
xor \U$47011 ( \46986 , \45925 , \45942 );
buf \U$47012 ( \46987 , \46986 );
buf \U$47013 ( \46988 , \46987 );
buf \U$47014 ( \46989 , RIc0d90b8_57);
buf \U$47015 ( \46990 , RIc0da468_99);
xor \U$47016 ( \46991 , \46989 , \46990 );
buf \U$47017 ( \46992 , \46991 );
buf \U$47018 ( \46993 , \46992 );
not \U$47019 ( \46994 , \46993 );
buf \U$47020 ( \46995 , \19695 );
not \U$47021 ( \46996 , \46995 );
or \U$47022 ( \46997 , \46994 , \46996 );
buf \U$47023 ( \46998 , \14140 );
buf \U$47024 ( \46999 , \45408 );
nand \U$47025 ( \47000 , \46998 , \46999 );
buf \U$47026 ( \47001 , \47000 );
buf \U$47027 ( \47002 , \47001 );
nand \U$47028 ( \47003 , \46997 , \47002 );
buf \U$47029 ( \47004 , \47003 );
buf \U$47030 ( \47005 , \47004 );
not \U$47031 ( \47006 , \47005 );
buf \U$47032 ( \47007 , RIc0da198_93);
buf \U$47033 ( \47008 , RIc0d9388_63);
xor \U$47034 ( \47009 , \47007 , \47008 );
buf \U$47035 ( \47010 , \47009 );
buf \U$47036 ( \47011 , \47010 );
not \U$47037 ( \47012 , \47011 );
buf \U$47038 ( \47013 , \13569 );
not \U$47039 ( \47014 , \47013 );
or \U$47040 ( \47015 , \47012 , \47014 );
buf \U$47041 ( \47016 , \4008 );
buf \U$47042 ( \47017 , \45929 );
nand \U$47043 ( \47018 , \47016 , \47017 );
buf \U$47044 ( \47019 , \47018 );
buf \U$47045 ( \47020 , \47019 );
nand \U$47046 ( \47021 , \47015 , \47020 );
buf \U$47047 ( \47022 , \47021 );
buf \U$47048 ( \47023 , \47022 );
not \U$47049 ( \47024 , \47023 );
or \U$47050 ( \47025 , \47006 , \47024 );
buf \U$47051 ( \47026 , \47022 );
buf \U$47052 ( \47027 , \47004 );
or \U$47053 ( \47028 , \47026 , \47027 );
buf \U$47054 ( \47029 , RIc0d8578_33);
buf \U$47055 ( \47030 , RIc0dafa8_123);
xor \U$47056 ( \47031 , \47029 , \47030 );
buf \U$47057 ( \47032 , \47031 );
buf \U$47058 ( \47033 , \47032 );
not \U$47059 ( \47034 , \47033 );
buf \U$47060 ( \47035 , \46183 );
not \U$47061 ( \47036 , \47035 );
buf \U$47062 ( \47037 , \47036 );
buf \U$47063 ( \47038 , \47037 );
not \U$47064 ( \47039 , \47038 );
or \U$47065 ( \47040 , \47034 , \47039 );
buf \U$47066 ( \47041 , \45094 );
not \U$47067 ( \47042 , \47041 );
buf \U$47068 ( \47043 , \16692 );
nand \U$47069 ( \47044 , \47042 , \47043 );
buf \U$47070 ( \47045 , \47044 );
buf \U$47071 ( \47046 , \47045 );
nand \U$47072 ( \47047 , \47040 , \47046 );
buf \U$47073 ( \47048 , \47047 );
buf \U$47074 ( \47049 , \47048 );
nand \U$47075 ( \47050 , \47028 , \47049 );
buf \U$47076 ( \47051 , \47050 );
buf \U$47077 ( \47052 , \47051 );
nand \U$47078 ( \47053 , \47025 , \47052 );
buf \U$47079 ( \47054 , \47053 );
buf \U$47080 ( \47055 , \47054 );
xor \U$47081 ( \47056 , \46988 , \47055 );
xnor \U$47082 ( \47057 , RIc0da918_109, RIc0d8c08_47);
buf \U$47083 ( \47058 , \47057 );
not \U$47084 ( \47059 , \47058 );
buf \U$47085 ( \47060 , \47059 );
buf \U$47086 ( \47061 , \47060 );
not \U$47087 ( \47062 , \47061 );
buf \U$47088 ( \47063 , \21959 );
not \U$47089 ( \47064 , \47063 );
or \U$47090 ( \47065 , \47062 , \47064 );
buf \U$47091 ( \47066 , \16232 );
buf \U$47092 ( \47067 , \45044 );
nand \U$47093 ( \47068 , \47066 , \47067 );
buf \U$47094 ( \47069 , \47068 );
buf \U$47095 ( \47070 , \47069 );
nand \U$47096 ( \47071 , \47065 , \47070 );
buf \U$47097 ( \47072 , \47071 );
buf \U$47098 ( \47073 , \47072 );
not \U$47099 ( \47074 , \47073 );
buf \U$47100 ( \47075 , RIc0d8de8_51);
buf \U$47101 ( \47076 , RIc0da738_105);
xor \U$47102 ( \47077 , \47075 , \47076 );
buf \U$47103 ( \47078 , \47077 );
buf \U$47104 ( \47079 , \47078 );
not \U$47105 ( \47080 , \47079 );
buf \U$47106 ( \47081 , \15644 );
not \U$47107 ( \47082 , \47081 );
or \U$47108 ( \47083 , \47080 , \47082 );
buf \U$47109 ( \47084 , \12744 );
buf \U$47110 ( \47085 , \45168 );
nand \U$47111 ( \47086 , \47084 , \47085 );
buf \U$47112 ( \47087 , \47086 );
buf \U$47113 ( \47088 , \47087 );
nand \U$47114 ( \47089 , \47083 , \47088 );
buf \U$47115 ( \47090 , \47089 );
buf \U$47116 ( \47091 , \47090 );
not \U$47117 ( \47092 , \47091 );
or \U$47118 ( \47093 , \47074 , \47092 );
buf \U$47119 ( \47094 , \47090 );
buf \U$47120 ( \47095 , \47072 );
or \U$47121 ( \47096 , \47094 , \47095 );
buf \U$47122 ( \47097 , RIc0d8ed8_53);
buf \U$47123 ( \47098 , RIc0da648_103);
xor \U$47124 ( \47099 , \47097 , \47098 );
buf \U$47125 ( \47100 , \47099 );
buf \U$47126 ( \47101 , \47100 );
not \U$47127 ( \47102 , \47101 );
buf \U$47128 ( \47103 , \13042 );
not \U$47129 ( \47104 , \47103 );
or \U$47130 ( \47105 , \47102 , \47104 );
buf \U$47131 ( \47106 , \18416 );
buf \U$47132 ( \47107 , \45276 );
nand \U$47133 ( \47108 , \47106 , \47107 );
buf \U$47134 ( \47109 , \47108 );
buf \U$47135 ( \47110 , \47109 );
nand \U$47136 ( \47111 , \47105 , \47110 );
buf \U$47137 ( \47112 , \47111 );
buf \U$47138 ( \47113 , \47112 );
nand \U$47139 ( \47114 , \47096 , \47113 );
buf \U$47140 ( \47115 , \47114 );
buf \U$47141 ( \47116 , \47115 );
nand \U$47142 ( \47117 , \47093 , \47116 );
buf \U$47143 ( \47118 , \47117 );
buf \U$47144 ( \47119 , \47118 );
and \U$47145 ( \47120 , \47056 , \47119 );
and \U$47146 ( \47121 , \46988 , \47055 );
or \U$47147 ( \47122 , \47120 , \47121 );
buf \U$47148 ( \47123 , \47122 );
buf \U$47149 ( \47124 , \47123 );
xor \U$47150 ( \47125 , \46985 , \47124 );
buf \U$47151 ( \47126 , RIc0d8398_29);
buf \U$47152 ( \47127 , RIc0db188_127);
xor \U$47153 ( \47128 , \47126 , \47127 );
buf \U$47154 ( \47129 , \47128 );
buf \U$47155 ( \47130 , \47129 );
not \U$47156 ( \47131 , \47130 );
buf \U$47157 ( \47132 , \15609 );
not \U$47158 ( \47133 , \47132 );
or \U$47159 ( \47134 , \47131 , \47133 );
buf \U$47160 ( \47135 , \45322 );
buf \U$47161 ( \47136 , RIc0db200_128);
nand \U$47162 ( \47137 , \47135 , \47136 );
buf \U$47163 ( \47138 , \47137 );
buf \U$47164 ( \47139 , \47138 );
nand \U$47165 ( \47140 , \47134 , \47139 );
buf \U$47166 ( \47141 , \47140 );
buf \U$47167 ( \47142 , \47141 );
buf \U$47168 ( \47143 , \45295 );
not \U$47169 ( \47144 , \47143 );
buf \U$47170 ( \47145 , \12342 );
not \U$47171 ( \47146 , \47145 );
or \U$47172 ( \47147 , \47144 , \47146 );
buf \U$47173 ( \47148 , RIc0d8cf8_49);
buf \U$47174 ( \47149 , RIc0da828_107);
xnor \U$47175 ( \47150 , \47148 , \47149 );
buf \U$47176 ( \47151 , \47150 );
buf \U$47177 ( \47152 , \47151 );
not \U$47178 ( \47153 , \47152 );
buf \U$47179 ( \47154 , \16064 );
buf \U$47180 ( \47155 , \12327 );
nand \U$47181 ( \47156 , \47153 , \47154 , \47155 );
buf \U$47182 ( \47157 , \47156 );
buf \U$47183 ( \47158 , \47157 );
nand \U$47184 ( \47159 , \47147 , \47158 );
buf \U$47185 ( \47160 , \47159 );
buf \U$47186 ( \47161 , \47160 );
xor \U$47187 ( \47162 , \47142 , \47161 );
buf \U$47188 ( \47163 , RIc0d8b18_45);
buf \U$47189 ( \47164 , RIc0daa08_111);
xor \U$47190 ( \47165 , \47163 , \47164 );
buf \U$47191 ( \47166 , \47165 );
buf \U$47192 ( \47167 , \47166 );
not \U$47193 ( \47168 , \47167 );
buf \U$47194 ( \47169 , \14346 );
not \U$47195 ( \47170 , \47169 );
or \U$47196 ( \47171 , \47168 , \47170 );
buf \U$47197 ( \47172 , \14106 );
buf \U$47198 ( \47173 , \45254 );
nand \U$47199 ( \47174 , \47172 , \47173 );
buf \U$47200 ( \47175 , \47174 );
buf \U$47201 ( \47176 , \47175 );
nand \U$47202 ( \47177 , \47171 , \47176 );
buf \U$47203 ( \47178 , \47177 );
buf \U$47204 ( \47179 , \47178 );
and \U$47205 ( \47180 , \47162 , \47179 );
and \U$47206 ( \47181 , \47142 , \47161 );
or \U$47207 ( \47182 , \47180 , \47181 );
buf \U$47208 ( \47183 , \47182 );
buf \U$47209 ( \47184 , \47183 );
buf \U$47210 ( \47185 , \533 );
buf \U$47211 ( \47186 , RIc0d9400_64);
and \U$47212 ( \47187 , \47185 , \47186 );
buf \U$47213 ( \47188 , \47187 );
buf \U$47214 ( \47189 , \47188 );
buf \U$47215 ( \47190 , RIc0dadc8_119);
buf \U$47216 ( \47191 , RIc0d8758_37);
xor \U$47217 ( \47192 , \47190 , \47191 );
buf \U$47218 ( \47193 , \47192 );
buf \U$47219 ( \47194 , \47193 );
not \U$47220 ( \47195 , \47194 );
buf \U$47221 ( \47196 , \23985 );
not \U$47222 ( \47197 , \47196 );
or \U$47223 ( \47198 , \47195 , \47197 );
buf \U$47224 ( \47199 , \45220 );
not \U$47225 ( \47200 , \47199 );
buf \U$47226 ( \47201 , \13005 );
nand \U$47227 ( \47202 , \47200 , \47201 );
buf \U$47228 ( \47203 , \47202 );
buf \U$47229 ( \47204 , \47203 );
nand \U$47230 ( \47205 , \47198 , \47204 );
buf \U$47231 ( \47206 , \47205 );
buf \U$47232 ( \47207 , \47206 );
xor \U$47233 ( \47208 , \47189 , \47207 );
buf \U$47234 ( \47209 , \14713 );
buf \U$47235 ( \47210 , RIc0da288_95);
buf \U$47236 ( \47211 , RIc0d9298_61);
xor \U$47237 ( \47212 , \47210 , \47211 );
buf \U$47238 ( \47213 , \47212 );
buf \U$47239 ( \47214 , \47213 );
not \U$47240 ( \47215 , \47214 );
buf \U$47241 ( \47216 , \47215 );
buf \U$47242 ( \47217 , \47216 );
or \U$47243 ( \47218 , \47209 , \47217 );
buf \U$47244 ( \47219 , \4849 );
buf \U$47245 ( \47220 , \45437 );
or \U$47246 ( \47221 , \47219 , \47220 );
nand \U$47247 ( \47222 , \47218 , \47221 );
buf \U$47248 ( \47223 , \47222 );
buf \U$47249 ( \47224 , \47223 );
and \U$47250 ( \47225 , \47208 , \47224 );
and \U$47251 ( \47226 , \47189 , \47207 );
or \U$47252 ( \47227 , \47225 , \47226 );
buf \U$47253 ( \47228 , \47227 );
buf \U$47254 ( \47229 , \47228 );
xor \U$47255 ( \47230 , \47184 , \47229 );
buf \U$47256 ( \47231 , RIc0da558_101);
buf \U$47257 ( \47232 , RIc0d8fc8_55);
xor \U$47258 ( \47233 , \47231 , \47232 );
buf \U$47259 ( \47234 , \47233 );
buf \U$47260 ( \47235 , \47234 );
not \U$47261 ( \47236 , \47235 );
buf \U$47262 ( \47237 , \33258 );
not \U$47263 ( \47238 , \47237 );
or \U$47264 ( \47239 , \47236 , \47238 );
buf \U$47265 ( \47240 , \26354 );
buf \U$47266 ( \47241 , \45122 );
nand \U$47267 ( \47242 , \47240 , \47241 );
buf \U$47268 ( \47243 , \47242 );
buf \U$47269 ( \47244 , \47243 );
nand \U$47270 ( \47245 , \47239 , \47244 );
buf \U$47271 ( \47246 , \47245 );
buf \U$47272 ( \47247 , \47246 );
buf \U$47273 ( \47248 , RIc0d8a28_43);
buf \U$47274 ( \47249 , RIc0daaf8_113);
xor \U$47275 ( \47250 , \47248 , \47249 );
buf \U$47276 ( \47251 , \47250 );
buf \U$47277 ( \47252 , \47251 );
not \U$47278 ( \47253 , \47252 );
buf \U$47279 ( \47254 , \25355 );
not \U$47280 ( \47255 , \47254 );
or \U$47281 ( \47256 , \47253 , \47255 );
buf \U$47282 ( \47257 , \16995 );
buf \U$47283 ( \47258 , \45196 );
nand \U$47284 ( \47259 , \47257 , \47258 );
buf \U$47285 ( \47260 , \47259 );
buf \U$47286 ( \47261 , \47260 );
nand \U$47287 ( \47262 , \47256 , \47261 );
buf \U$47288 ( \47263 , \47262 );
buf \U$47289 ( \47264 , \47263 );
xor \U$47290 ( \47265 , \47247 , \47264 );
buf \U$47291 ( \47266 , RIc0db098_125);
buf \U$47292 ( \47267 , RIc0d8488_31);
xnor \U$47293 ( \47268 , \47266 , \47267 );
buf \U$47294 ( \47269 , \47268 );
buf \U$47295 ( \47270 , \47269 );
not \U$47296 ( \47271 , \47270 );
buf \U$47297 ( \47272 , \47271 );
buf \U$47298 ( \47273 , \47272 );
not \U$47299 ( \47274 , \47273 );
buf \U$47300 ( \47275 , \44813 );
not \U$47301 ( \47276 , \47275 );
or \U$47302 ( \47277 , \47274 , \47276 );
buf \U$47303 ( \47278 , \13465 );
buf \U$47304 ( \47279 , \45108 );
nand \U$47305 ( \47280 , \47278 , \47279 );
buf \U$47306 ( \47281 , \47280 );
buf \U$47307 ( \47282 , \47281 );
nand \U$47308 ( \47283 , \47277 , \47282 );
buf \U$47309 ( \47284 , \47283 );
buf \U$47310 ( \47285 , \47284 );
and \U$47311 ( \47286 , \47265 , \47285 );
and \U$47312 ( \47287 , \47247 , \47264 );
or \U$47313 ( \47288 , \47286 , \47287 );
buf \U$47314 ( \47289 , \47288 );
buf \U$47315 ( \47290 , \47289 );
and \U$47316 ( \47291 , \47230 , \47290 );
and \U$47317 ( \47292 , \47184 , \47229 );
or \U$47318 ( \47293 , \47291 , \47292 );
buf \U$47319 ( \47294 , \47293 );
buf \U$47320 ( \47295 , \47294 );
and \U$47321 ( \47296 , \47125 , \47295 );
and \U$47322 ( \47297 , \46985 , \47124 );
or \U$47323 ( \47298 , \47296 , \47297 );
buf \U$47324 ( \47299 , \47298 );
buf \U$47325 ( \47300 , \47299 );
xor \U$47326 ( \47301 , \45121 , \45135 );
xor \U$47327 ( \47302 , \47301 , \45158 );
buf \U$47328 ( \47303 , \47302 );
buf \U$47329 ( \47304 , \47303 );
xor \U$47330 ( \47305 , \45339 , \45357 );
xor \U$47331 ( \47306 , \47305 , \45376 );
buf \U$47332 ( \47307 , \47306 );
buf \U$47333 ( \47308 , \47307 );
or \U$47334 ( \47309 , \47304 , \47308 );
xor \U$47335 ( \47310 , \45404 , \45425 );
xor \U$47336 ( \47311 , \47310 , \45442 );
buf \U$47337 ( \47312 , \47311 );
buf \U$47338 ( \47313 , \47312 );
nand \U$47339 ( \47314 , \47309 , \47313 );
buf \U$47340 ( \47315 , \47314 );
buf \U$47341 ( \47316 , \47315 );
buf \U$47342 ( \47317 , \47303 );
buf \U$47343 ( \47318 , \47307 );
nand \U$47344 ( \47319 , \47317 , \47318 );
buf \U$47345 ( \47320 , \47319 );
buf \U$47346 ( \47321 , \47320 );
nand \U$47347 ( \47322 , \47316 , \47321 );
buf \U$47348 ( \47323 , \47322 );
buf \U$47349 ( \47324 , \47323 );
xor \U$47350 ( \47325 , \45058 , \45076 );
xor \U$47351 ( \47326 , \47325 , \45099 );
buf \U$47352 ( \47327 , \47326 );
buf \U$47353 ( \47328 , \47327 );
buf \U$47354 ( \47329 , RIc0da378_97);
buf \U$47355 ( \47330 , RIc0d91a8_59);
xor \U$47356 ( \47331 , \47329 , \47330 );
buf \U$47357 ( \47332 , \47331 );
buf \U$47358 ( \47333 , \47332 );
not \U$47359 ( \47334 , \47333 );
buf \U$47360 ( \47335 , \2066 );
not \U$47361 ( \47336 , \47335 );
or \U$47362 ( \47337 , \47334 , \47336 );
buf \U$47363 ( \47338 , \734 );
buf \U$47364 ( \47339 , \45362 );
nand \U$47365 ( \47340 , \47338 , \47339 );
buf \U$47366 ( \47341 , \47340 );
buf \U$47367 ( \47342 , \47341 );
nand \U$47368 ( \47343 , \47337 , \47342 );
buf \U$47369 ( \47344 , \47343 );
buf \U$47370 ( \47345 , \47344 );
buf \U$47371 ( \47346 , RIc0dacd8_117);
buf \U$47372 ( \47347 , RIc0d8848_39);
xor \U$47373 ( \47348 , \47346 , \47347 );
buf \U$47374 ( \47349 , \47348 );
buf \U$47375 ( \47350 , \47349 );
not \U$47376 ( \47351 , \47350 );
buf \U$47377 ( \47352 , \12929 );
not \U$47378 ( \47353 , \47352 );
or \U$47379 ( \47354 , \47351 , \47353 );
buf \U$47380 ( \47355 , \22356 );
buf \U$47381 ( \47356 , \45059 );
nand \U$47382 ( \47357 , \47355 , \47356 );
buf \U$47383 ( \47358 , \47357 );
buf \U$47384 ( \47359 , \47358 );
nand \U$47385 ( \47360 , \47354 , \47359 );
buf \U$47386 ( \47361 , \47360 );
buf \U$47387 ( \47362 , \47361 );
xor \U$47388 ( \47363 , \47345 , \47362 );
buf \U$47389 ( \47364 , RIc0d8938_41);
buf \U$47390 ( \47365 , RIc0dabe8_115);
xor \U$47391 ( \47366 , \47364 , \47365 );
buf \U$47392 ( \47367 , \47366 );
buf \U$47393 ( \47368 , \47367 );
not \U$47394 ( \47369 , \47368 );
buf \U$47395 ( \47370 , \27743 );
not \U$47396 ( \47371 , \47370 );
or \U$47397 ( \47372 , \47369 , \47371 );
buf \U$47398 ( \47373 , \12303 );
buf \U$47399 ( \47374 , \45140 );
nand \U$47400 ( \47375 , \47373 , \47374 );
buf \U$47401 ( \47376 , \47375 );
buf \U$47402 ( \47377 , \47376 );
nand \U$47403 ( \47378 , \47372 , \47377 );
buf \U$47404 ( \47379 , \47378 );
buf \U$47405 ( \47380 , \47379 );
and \U$47406 ( \47381 , \47363 , \47380 );
and \U$47407 ( \47382 , \47345 , \47362 );
or \U$47408 ( \47383 , \47381 , \47382 );
buf \U$47409 ( \47384 , \47383 );
buf \U$47410 ( \47385 , \47384 );
xor \U$47411 ( \47386 , \47328 , \47385 );
xor \U$47412 ( \47387 , \45185 , \45214 );
xor \U$47413 ( \47388 , \47387 , \45235 );
buf \U$47414 ( \47389 , \47388 );
buf \U$47415 ( \47390 , \47389 );
and \U$47416 ( \47391 , \47386 , \47390 );
and \U$47417 ( \47392 , \47328 , \47385 );
or \U$47418 ( \47393 , \47391 , \47392 );
buf \U$47419 ( \47394 , \47393 );
buf \U$47420 ( \47395 , \47394 );
xor \U$47421 ( \47396 , \47324 , \47395 );
xor \U$47422 ( \47397 , \45104 , \45163 );
xor \U$47423 ( \47398 , \47397 , \45240 );
buf \U$47424 ( \47399 , \47398 );
buf \U$47425 ( \47400 , \47399 );
and \U$47426 ( \47401 , \47396 , \47400 );
and \U$47427 ( \47402 , \47324 , \47395 );
or \U$47428 ( \47403 , \47401 , \47402 );
buf \U$47429 ( \47404 , \47403 );
buf \U$47430 ( \47405 , \47404 );
xor \U$47431 ( \47406 , \47300 , \47405 );
xor \U$47432 ( \47407 , \45245 , \45249 );
xor \U$47433 ( \47408 , \47407 , \45452 );
buf \U$47434 ( \47409 , \47408 );
buf \U$47435 ( \47410 , \47409 );
and \U$47436 ( \47411 , \47406 , \47410 );
and \U$47437 ( \47412 , \47300 , \47405 );
or \U$47438 ( \47413 , \47411 , \47412 );
buf \U$47439 ( \47414 , \47413 );
buf \U$47440 ( \47415 , \47414 );
xor \U$47441 ( \47416 , \45489 , \45783 );
xor \U$47442 ( \47417 , \47416 , \45974 );
buf \U$47443 ( \47418 , \47417 );
buf \U$47444 ( \47419 , \47418 );
xor \U$47445 ( \47420 , \47415 , \47419 );
xor \U$47446 ( \47421 , \46326 , \46330 );
xor \U$47447 ( \47422 , \47421 , \46335 );
buf \U$47448 ( \47423 , \47422 );
buf \U$47449 ( \47424 , \47423 );
and \U$47450 ( \47425 , \47420 , \47424 );
and \U$47451 ( \47426 , \47415 , \47419 );
or \U$47452 ( \47427 , \47425 , \47426 );
buf \U$47453 ( \47428 , \47427 );
buf \U$47454 ( \47429 , \47428 );
nand \U$47455 ( \47430 , \46981 , \47429 );
buf \U$47456 ( \47431 , \47430 );
buf \U$47457 ( \47432 , \47431 );
buf \U$47458 ( \47433 , \46975 );
buf \U$47459 ( \47434 , \46979 );
nand \U$47460 ( \47435 , \47433 , \47434 );
buf \U$47461 ( \47436 , \47435 );
buf \U$47462 ( \47437 , \47436 );
nand \U$47463 ( \47438 , \47432 , \47437 );
buf \U$47464 ( \47439 , \47438 );
buf \U$47465 ( \47440 , \47439 );
or \U$47466 ( \47441 , \46972 , \47440 );
buf \U$47467 ( \47442 , \47441 );
buf \U$47468 ( \47443 , \47442 );
xor \U$47469 ( \47444 , \47415 , \47419 );
xor \U$47470 ( \47445 , \47444 , \47424 );
buf \U$47471 ( \47446 , \47445 );
not \U$47472 ( \47447 , \47446 );
xor \U$47473 ( \47448 , \45318 , \45381 );
xor \U$47474 ( \47449 , \47448 , \45447 );
buf \U$47475 ( \47450 , \47449 );
buf \U$47476 ( \47451 , \47450 );
buf \U$47477 ( \47452 , \45741 );
not \U$47478 ( \47453 , \47452 );
buf \U$47479 ( \47454 , \45685 );
not \U$47480 ( \47455 , \47454 );
or \U$47481 ( \47456 , \47453 , \47455 );
buf \U$47482 ( \47457 , \45672 );
buf \U$47483 ( \47458 , \45738 );
nand \U$47484 ( \47459 , \47457 , \47458 );
buf \U$47485 ( \47460 , \47459 );
buf \U$47486 ( \47461 , \47460 );
nand \U$47487 ( \47462 , \47456 , \47461 );
buf \U$47488 ( \47463 , \47462 );
buf \U$47489 ( \47464 , \47463 );
buf \U$47490 ( \47465 , \45679 );
and \U$47491 ( \47466 , \47464 , \47465 );
not \U$47492 ( \47467 , \47464 );
buf \U$47493 ( \47468 , \45676 );
and \U$47494 ( \47469 , \47467 , \47468 );
nor \U$47495 ( \47470 , \47466 , \47469 );
buf \U$47496 ( \47471 , \47470 );
buf \U$47497 ( \47472 , \47471 );
xor \U$47498 ( \47473 , \47451 , \47472 );
buf \U$47499 ( \47474 , \45581 );
not \U$47500 ( \47475 , \47474 );
buf \U$47501 ( \47476 , \45626 );
not \U$47502 ( \47477 , \47476 );
or \U$47503 ( \47478 , \47475 , \47477 );
buf \U$47504 ( \47479 , \45626 );
buf \U$47505 ( \47480 , \45581 );
or \U$47506 ( \47481 , \47479 , \47480 );
nand \U$47507 ( \47482 , \47478 , \47481 );
buf \U$47508 ( \47483 , \47482 );
buf \U$47509 ( \47484 , \47483 );
buf \U$47510 ( \47485 , \45531 );
and \U$47511 ( \47486 , \47484 , \47485 );
not \U$47512 ( \47487 , \47484 );
buf \U$47513 ( \47488 , \45528 );
and \U$47514 ( \47489 , \47487 , \47488 );
nor \U$47515 ( \47490 , \47486 , \47489 );
buf \U$47516 ( \47491 , \47490 );
buf \U$47517 ( \47492 , \47491 );
and \U$47518 ( \47493 , \47473 , \47492 );
and \U$47519 ( \47494 , \47451 , \47472 );
or \U$47520 ( \47495 , \47493 , \47494 );
buf \U$47521 ( \47496 , \47495 );
buf \U$47522 ( \47497 , \47496 );
not \U$47523 ( \47498 , \47497 );
xor \U$47524 ( \47499 , \45633 , \45748 );
xor \U$47525 ( \47500 , \47499 , \45778 );
buf \U$47526 ( \47501 , \47500 );
buf \U$47527 ( \47502 , \47501 );
not \U$47528 ( \47503 , \47502 );
or \U$47529 ( \47504 , \47498 , \47503 );
buf \U$47530 ( \47505 , \47501 );
buf \U$47531 ( \47506 , \47496 );
or \U$47532 ( \47507 , \47505 , \47506 );
xor \U$47533 ( \47508 , \45850 , \45875 );
xor \U$47534 ( \47509 , \47508 , \45969 );
buf \U$47535 ( \47510 , \47509 );
buf \U$47536 ( \47511 , \47510 );
nand \U$47537 ( \47512 , \47507 , \47511 );
buf \U$47538 ( \47513 , \47512 );
buf \U$47539 ( \47514 , \47513 );
nand \U$47540 ( \47515 , \47504 , \47514 );
buf \U$47541 ( \47516 , \47515 );
buf \U$47542 ( \47517 , \47516 );
not \U$47543 ( \47518 , \47517 );
xor \U$47544 ( \47519 , \47300 , \47405 );
xor \U$47545 ( \47520 , \47519 , \47410 );
buf \U$47546 ( \47521 , \47520 );
buf \U$47547 ( \47522 , \47521 );
not \U$47548 ( \47523 , \47522 );
xor \U$47549 ( \47524 , \46988 , \47055 );
xor \U$47550 ( \47525 , \47524 , \47119 );
buf \U$47551 ( \47526 , \47525 );
buf \U$47552 ( \47527 , \47526 );
xor \U$47553 ( \47528 , \47312 , \47307 );
xor \U$47554 ( \47529 , \47528 , \47303 );
buf \U$47555 ( \47530 , \47529 );
xor \U$47556 ( \47531 , \47527 , \47530 );
xor \U$47557 ( \47532 , \47328 , \47385 );
xor \U$47558 ( \47533 , \47532 , \47390 );
buf \U$47559 ( \47534 , \47533 );
buf \U$47560 ( \47535 , \47534 );
and \U$47561 ( \47536 , \47531 , \47535 );
and \U$47562 ( \47537 , \47527 , \47530 );
or \U$47563 ( \47538 , \47536 , \47537 );
buf \U$47564 ( \47539 , \47538 );
buf \U$47565 ( \47540 , \47539 );
xor \U$47566 ( \47541 , \47324 , \47395 );
xor \U$47567 ( \47542 , \47541 , \47400 );
buf \U$47568 ( \47543 , \47542 );
buf \U$47569 ( \47544 , \47543 );
xor \U$47570 ( \47545 , \47540 , \47544 );
xor \U$47571 ( \47546 , \47451 , \47472 );
xor \U$47572 ( \47547 , \47546 , \47492 );
buf \U$47573 ( \47548 , \47547 );
buf \U$47574 ( \47549 , \47548 );
and \U$47575 ( \47550 , \47545 , \47549 );
and \U$47576 ( \47551 , \47540 , \47544 );
or \U$47577 ( \47552 , \47550 , \47551 );
buf \U$47578 ( \47553 , \47552 );
buf \U$47579 ( \47554 , \47553 );
not \U$47580 ( \47555 , \47554 );
or \U$47581 ( \47556 , \47523 , \47555 );
buf \U$47582 ( \47557 , \47553 );
buf \U$47583 ( \47558 , \47521 );
or \U$47584 ( \47559 , \47557 , \47558 );
xor \U$47585 ( \47560 , \45288 , \45311 );
xor \U$47586 ( \47561 , \47560 , \45270 );
buf \U$47587 ( \47562 , \47561 );
buf \U$47588 ( \47563 , \16386 );
not \U$47589 ( \47564 , \47563 );
buf \U$47590 ( \47565 , \45386 );
not \U$47591 ( \47566 , \47565 );
or \U$47592 ( \47567 , \47564 , \47566 );
buf \U$47593 ( \47568 , \13310 );
not \U$47594 ( \47569 , \47568 );
buf \U$47595 ( \47570 , \47569 );
buf \U$47596 ( \47571 , \47570 );
buf \U$47597 ( \47572 , RIc0d8668_35);
buf \U$47598 ( \47573 , RIc0daeb8_121);
xnor \U$47599 ( \47574 , \47572 , \47573 );
buf \U$47600 ( \47575 , \47574 );
buf \U$47601 ( \47576 , \47575 );
or \U$47602 ( \47577 , \47571 , \47576 );
nand \U$47603 ( \47578 , \47567 , \47577 );
buf \U$47604 ( \47579 , \47578 );
buf \U$47605 ( \47580 , \47579 );
xor \U$47606 ( \47581 , RIc0da288_95, RIc0d9310_62);
buf \U$47607 ( \47582 , \47581 );
not \U$47608 ( \47583 , \47582 );
buf \U$47609 ( \47584 , \330 );
not \U$47610 ( \47585 , \47584 );
or \U$47611 ( \47586 , \47583 , \47585 );
buf \U$47612 ( \47587 , \344 );
buf \U$47613 ( \47588 , \47213 );
nand \U$47614 ( \47589 , \47587 , \47588 );
buf \U$47615 ( \47590 , \47589 );
buf \U$47616 ( \47591 , \47590 );
nand \U$47617 ( \47592 , \47586 , \47591 );
buf \U$47618 ( \47593 , \47592 );
buf \U$47619 ( \47594 , \47593 );
not \U$47620 ( \47595 , \47594 );
buf \U$47621 ( \47596 , RIc0d9400_64);
buf \U$47622 ( \47597 , RIc0da210_94);
or \U$47623 ( \47598 , \47596 , \47597 );
buf \U$47624 ( \47599 , RIc0da288_95);
nand \U$47625 ( \47600 , \47598 , \47599 );
buf \U$47626 ( \47601 , \47600 );
buf \U$47627 ( \47602 , \47601 );
buf \U$47628 ( \47603 , RIc0d9400_64);
buf \U$47629 ( \47604 , RIc0da210_94);
nand \U$47630 ( \47605 , \47603 , \47604 );
buf \U$47631 ( \47606 , \47605 );
buf \U$47632 ( \47607 , \47606 );
buf \U$47633 ( \47608 , RIc0da198_93);
nand \U$47634 ( \47609 , \47602 , \47607 , \47608 );
buf \U$47635 ( \47610 , \47609 );
buf \U$47636 ( \47611 , \47610 );
nor \U$47637 ( \47612 , \47595 , \47611 );
buf \U$47638 ( \47613 , \47612 );
buf \U$47639 ( \47614 , \47613 );
xor \U$47640 ( \47615 , \47580 , \47614 );
buf \U$47641 ( \47616 , \14207 );
not \U$47642 ( \47617 , \47616 );
buf \U$47643 ( \47618 , RIc0da918_109);
buf \U$47644 ( \47619 , RIc0d8c80_48);
xnor \U$47645 ( \47620 , \47618 , \47619 );
buf \U$47646 ( \47621 , \47620 );
buf \U$47647 ( \47622 , \47621 );
not \U$47648 ( \47623 , \47622 );
and \U$47649 ( \47624 , \47617 , \47623 );
buf \U$47650 ( \47625 , \36203 );
buf \U$47651 ( \47626 , \47057 );
nor \U$47652 ( \47627 , \47625 , \47626 );
buf \U$47653 ( \47628 , \47627 );
buf \U$47654 ( \47629 , \47628 );
nor \U$47655 ( \47630 , \47624 , \47629 );
buf \U$47656 ( \47631 , \47630 );
buf \U$47657 ( \47632 , \47631 );
not \U$47658 ( \47633 , \47632 );
buf \U$47659 ( \47634 , \47633 );
buf \U$47660 ( \47635 , \47634 );
buf \U$47661 ( \47636 , RIc0d9400_64);
buf \U$47662 ( \47637 , RIc0da198_93);
xor \U$47663 ( \47638 , \47636 , \47637 );
buf \U$47664 ( \47639 , \47638 );
buf \U$47665 ( \47640 , \47639 );
not \U$47666 ( \47641 , \47640 );
buf \U$47667 ( \47642 , \13569 );
not \U$47668 ( \47643 , \47642 );
or \U$47669 ( \47644 , \47641 , \47643 );
buf \U$47670 ( \47645 , \4008 );
buf \U$47671 ( \47646 , \47010 );
nand \U$47672 ( \47647 , \47645 , \47646 );
buf \U$47673 ( \47648 , \47647 );
buf \U$47674 ( \47649 , \47648 );
nand \U$47675 ( \47650 , \47644 , \47649 );
buf \U$47676 ( \47651 , \47650 );
buf \U$47677 ( \47652 , \47651 );
or \U$47678 ( \47653 , \47635 , \47652 );
buf \U$47679 ( \47654 , RIc0d85f0_34);
buf \U$47680 ( \47655 , RIc0dafa8_123);
xor \U$47681 ( \47656 , \47654 , \47655 );
buf \U$47682 ( \47657 , \47656 );
buf \U$47683 ( \47658 , \47657 );
not \U$47684 ( \47659 , \47658 );
buf \U$47685 ( \47660 , \47037 );
not \U$47686 ( \47661 , \47660 );
or \U$47687 ( \47662 , \47659 , \47661 );
buf \U$47688 ( \47663 , \16692 );
buf \U$47689 ( \47664 , \47032 );
nand \U$47690 ( \47665 , \47663 , \47664 );
buf \U$47691 ( \47666 , \47665 );
buf \U$47692 ( \47667 , \47666 );
nand \U$47693 ( \47668 , \47662 , \47667 );
buf \U$47694 ( \47669 , \47668 );
buf \U$47695 ( \47670 , \47669 );
nand \U$47696 ( \47671 , \47653 , \47670 );
buf \U$47697 ( \47672 , \47671 );
buf \U$47698 ( \47673 , \47672 );
buf \U$47699 ( \47674 , \47634 );
buf \U$47700 ( \47675 , \47651 );
nand \U$47701 ( \47676 , \47674 , \47675 );
buf \U$47702 ( \47677 , \47676 );
buf \U$47703 ( \47678 , \47677 );
nand \U$47704 ( \47679 , \47673 , \47678 );
buf \U$47705 ( \47680 , \47679 );
buf \U$47706 ( \47681 , \47680 );
and \U$47707 ( \47682 , \47615 , \47681 );
and \U$47708 ( \47683 , \47580 , \47614 );
or \U$47709 ( \47684 , \47682 , \47683 );
buf \U$47710 ( \47685 , \47684 );
buf \U$47711 ( \47686 , \47685 );
xor \U$47712 ( \47687 , \47562 , \47686 );
buf \U$47713 ( \47688 , RIc0daa08_111);
buf \U$47714 ( \47689 , RIc0d8b90_46);
xor \U$47715 ( \47690 , \47688 , \47689 );
buf \U$47716 ( \47691 , \47690 );
buf \U$47717 ( \47692 , \47691 );
not \U$47718 ( \47693 , \47692 );
buf \U$47719 ( \47694 , \12529 );
not \U$47720 ( \47695 , \47694 );
or \U$47721 ( \47696 , \47693 , \47695 );
buf \U$47722 ( \47697 , \18312 );
buf \U$47723 ( \47698 , \47166 );
nand \U$47724 ( \47699 , \47697 , \47698 );
buf \U$47725 ( \47700 , \47699 );
buf \U$47726 ( \47701 , \47700 );
nand \U$47727 ( \47702 , \47696 , \47701 );
buf \U$47728 ( \47703 , \47702 );
buf \U$47729 ( \47704 , \47703 );
buf \U$47730 ( \47705 , RIc0d8e60_52);
buf \U$47731 ( \47706 , RIc0da738_105);
xor \U$47732 ( \47707 , \47705 , \47706 );
buf \U$47733 ( \47708 , \47707 );
buf \U$47734 ( \47709 , \47708 );
not \U$47735 ( \47710 , \47709 );
buf \U$47736 ( \47711 , \12736 );
not \U$47737 ( \47712 , \47711 );
or \U$47738 ( \47713 , \47710 , \47712 );
buf \U$47739 ( \47714 , \12744 );
buf \U$47740 ( \47715 , \47078 );
nand \U$47741 ( \47716 , \47714 , \47715 );
buf \U$47742 ( \47717 , \47716 );
buf \U$47743 ( \47718 , \47717 );
nand \U$47744 ( \47719 , \47713 , \47718 );
buf \U$47745 ( \47720 , \47719 );
buf \U$47746 ( \47721 , \47720 );
or \U$47747 ( \47722 , \47704 , \47721 );
xor \U$47748 ( \47723 , RIc0da648_103, RIc0d8f50_54);
buf \U$47749 ( \47724 , \47723 );
not \U$47750 ( \47725 , \47724 );
buf \U$47751 ( \47726 , \29546 );
not \U$47752 ( \47727 , \47726 );
or \U$47753 ( \47728 , \47725 , \47727 );
buf \U$47754 ( \47729 , \13712 );
buf \U$47755 ( \47730 , \47100 );
nand \U$47756 ( \47731 , \47729 , \47730 );
buf \U$47757 ( \47732 , \47731 );
buf \U$47758 ( \47733 , \47732 );
nand \U$47759 ( \47734 , \47728 , \47733 );
buf \U$47760 ( \47735 , \47734 );
buf \U$47761 ( \47736 , \47735 );
nand \U$47762 ( \47737 , \47722 , \47736 );
buf \U$47763 ( \47738 , \47737 );
buf \U$47764 ( \47739 , \47738 );
buf \U$47765 ( \47740 , \47703 );
buf \U$47766 ( \47741 , \47720 );
nand \U$47767 ( \47742 , \47740 , \47741 );
buf \U$47768 ( \47743 , \47742 );
buf \U$47769 ( \47744 , \47743 );
nand \U$47770 ( \47745 , \47739 , \47744 );
buf \U$47771 ( \47746 , \47745 );
buf \U$47772 ( \47747 , \47746 );
buf \U$47773 ( \47748 , RIc0d8aa0_44);
buf \U$47774 ( \47749 , RIc0daaf8_113);
xor \U$47775 ( \47750 , \47748 , \47749 );
buf \U$47776 ( \47751 , \47750 );
buf \U$47777 ( \47752 , \47751 );
not \U$47778 ( \47753 , \47752 );
buf \U$47779 ( \47754 , \28413 );
not \U$47780 ( \47755 , \47754 );
or \U$47781 ( \47756 , \47753 , \47755 );
buf \U$47782 ( \47757 , \16662 );
buf \U$47783 ( \47758 , \47251 );
nand \U$47784 ( \47759 , \47757 , \47758 );
buf \U$47785 ( \47760 , \47759 );
buf \U$47786 ( \47761 , \47760 );
nand \U$47787 ( \47762 , \47756 , \47761 );
buf \U$47788 ( \47763 , \47762 );
buf \U$47789 ( \47764 , \47763 );
not \U$47790 ( \47765 , \47764 );
buf \U$47791 ( \47766 , RIc0dadc8_119);
buf \U$47792 ( \47767 , RIc0d87d0_38);
xor \U$47793 ( \47768 , \47766 , \47767 );
buf \U$47794 ( \47769 , \47768 );
buf \U$47795 ( \47770 , \47769 );
not \U$47796 ( \47771 , \47770 );
buf \U$47797 ( \47772 , \13181 );
not \U$47798 ( \47773 , \47772 );
or \U$47799 ( \47774 , \47771 , \47773 );
buf \U$47800 ( \47775 , \13953 );
buf \U$47801 ( \47776 , \47193 );
nand \U$47802 ( \47777 , \47775 , \47776 );
buf \U$47803 ( \47778 , \47777 );
buf \U$47804 ( \47779 , \47778 );
nand \U$47805 ( \47780 , \47774 , \47779 );
buf \U$47806 ( \47781 , \47780 );
buf \U$47807 ( \47782 , \47781 );
not \U$47808 ( \47783 , \47782 );
or \U$47809 ( \47784 , \47765 , \47783 );
buf \U$47810 ( \47785 , \47781 );
buf \U$47811 ( \47786 , \47763 );
or \U$47812 ( \47787 , \47785 , \47786 );
buf \U$47813 ( \47788 , \14468 );
not \U$47814 ( \47789 , \47788 );
buf \U$47815 ( \47790 , RIc0d8500_32);
buf \U$47816 ( \47791 , RIc0db098_125);
xnor \U$47817 ( \47792 , \47790 , \47791 );
buf \U$47818 ( \47793 , \47792 );
buf \U$47819 ( \47794 , \47793 );
not \U$47820 ( \47795 , \47794 );
and \U$47821 ( \47796 , \47789 , \47795 );
buf \U$47822 ( \47797 , \18699 );
buf \U$47823 ( \47798 , \47269 );
nor \U$47824 ( \47799 , \47797 , \47798 );
buf \U$47825 ( \47800 , \47799 );
buf \U$47826 ( \47801 , \47800 );
nor \U$47827 ( \47802 , \47796 , \47801 );
buf \U$47828 ( \47803 , \47802 );
not \U$47829 ( \47804 , \47803 );
buf \U$47830 ( \47805 , \47804 );
nand \U$47831 ( \47806 , \47787 , \47805 );
buf \U$47832 ( \47807 , \47806 );
buf \U$47833 ( \47808 , \47807 );
nand \U$47834 ( \47809 , \47784 , \47808 );
buf \U$47835 ( \47810 , \47809 );
buf \U$47836 ( \47811 , \47810 );
xor \U$47837 ( \47812 , \47747 , \47811 );
buf \U$47838 ( \47813 , \3518 );
xor \U$47839 ( \47814 , RIc0da558_101, RIc0d9040_56);
buf \U$47840 ( \47815 , \47814 );
buf \U$47841 ( \47816 , \3521 );
nand \U$47842 ( \47817 , \47813 , \47815 , \47816 );
buf \U$47843 ( \47818 , \47817 );
buf \U$47844 ( \47819 , \47818 );
buf \U$47845 ( \47820 , \15550 );
buf \U$47846 ( \47821 , \47234 );
nand \U$47847 ( \47822 , \47820 , \47821 );
buf \U$47848 ( \47823 , \47822 );
buf \U$47849 ( \47824 , \47823 );
nand \U$47850 ( \47825 , \47819 , \47824 );
buf \U$47851 ( \47826 , \47825 );
buf \U$47852 ( \47827 , \47826 );
buf \U$47853 ( \47828 , RIc0d9220_60);
buf \U$47854 ( \47829 , RIc0da378_97);
xor \U$47855 ( \47830 , \47828 , \47829 );
buf \U$47856 ( \47831 , \47830 );
buf \U$47857 ( \47832 , \47831 );
not \U$47858 ( \47833 , \47832 );
buf \U$47859 ( \47834 , \2066 );
not \U$47860 ( \47835 , \47834 );
or \U$47861 ( \47836 , \47833 , \47835 );
buf \U$47862 ( \47837 , \734 );
buf \U$47863 ( \47838 , \47332 );
nand \U$47864 ( \47839 , \47837 , \47838 );
buf \U$47865 ( \47840 , \47839 );
buf \U$47866 ( \47841 , \47840 );
nand \U$47867 ( \47842 , \47836 , \47841 );
buf \U$47868 ( \47843 , \47842 );
buf \U$47869 ( \47844 , \47843 );
xor \U$47870 ( \47845 , \47827 , \47844 );
buf \U$47871 ( \47846 , RIc0d89b0_42);
buf \U$47872 ( \47847 , RIc0dabe8_115);
xor \U$47873 ( \47848 , \47846 , \47847 );
buf \U$47874 ( \47849 , \47848 );
buf \U$47875 ( \47850 , \47849 );
not \U$47876 ( \47851 , \47850 );
buf \U$47877 ( \47852 , \14186 );
not \U$47878 ( \47853 , \47852 );
or \U$47879 ( \47854 , \47851 , \47853 );
buf \U$47880 ( \47855 , \12303 );
buf \U$47881 ( \47856 , \47367 );
nand \U$47882 ( \47857 , \47855 , \47856 );
buf \U$47883 ( \47858 , \47857 );
buf \U$47884 ( \47859 , \47858 );
nand \U$47885 ( \47860 , \47854 , \47859 );
buf \U$47886 ( \47861 , \47860 );
buf \U$47887 ( \47862 , \47861 );
and \U$47888 ( \47863 , \47845 , \47862 );
and \U$47889 ( \47864 , \47827 , \47844 );
or \U$47890 ( \47865 , \47863 , \47864 );
buf \U$47891 ( \47866 , \47865 );
buf \U$47892 ( \47867 , \47866 );
and \U$47893 ( \47868 , \47812 , \47867 );
and \U$47894 ( \47869 , \47747 , \47811 );
or \U$47895 ( \47870 , \47868 , \47869 );
buf \U$47896 ( \47871 , \47870 );
buf \U$47897 ( \47872 , \47871 );
and \U$47898 ( \47873 , \47687 , \47872 );
and \U$47899 ( \47874 , \47562 , \47686 );
or \U$47900 ( \47875 , \47873 , \47874 );
buf \U$47901 ( \47876 , \47875 );
buf \U$47902 ( \47877 , \47876 );
not \U$47903 ( \47878 , \15609 );
buf \U$47904 ( \47879 , \47878 );
buf \U$47905 ( \47880 , RIc0d8410_30);
buf \U$47906 ( \47881 , RIc0db188_127);
xor \U$47907 ( \47882 , \47880 , \47881 );
buf \U$47908 ( \47883 , \47882 );
buf \U$47909 ( \47884 , \47883 );
not \U$47910 ( \47885 , \47884 );
buf \U$47911 ( \47886 , \47885 );
buf \U$47912 ( \47887 , \47886 );
or \U$47913 ( \47888 , \47879 , \47887 );
buf \U$47914 ( \47889 , \12647 );
buf \U$47915 ( \47890 , \47129 );
not \U$47916 ( \47891 , \47890 );
buf \U$47917 ( \47892 , \47891 );
buf \U$47918 ( \47893 , \47892 );
or \U$47919 ( \47894 , \47889 , \47893 );
nand \U$47920 ( \47895 , \47888 , \47894 );
buf \U$47921 ( \47896 , \47895 );
buf \U$47922 ( \47897 , \47896 );
xor \U$47923 ( \47898 , RIc0dacd8_117, RIc0d88c0_40);
buf \U$47924 ( \47899 , \47898 );
not \U$47925 ( \47900 , \47899 );
buf \U$47926 ( \47901 , \12923 );
not \U$47927 ( \47902 , \47901 );
or \U$47928 ( \47903 , \47900 , \47902 );
buf \U$47929 ( \47904 , \16559 );
buf \U$47930 ( \47905 , \47349 );
nand \U$47931 ( \47906 , \47904 , \47905 );
buf \U$47932 ( \47907 , \47906 );
buf \U$47933 ( \47908 , \47907 );
nand \U$47934 ( \47909 , \47903 , \47908 );
buf \U$47935 ( \47910 , \47909 );
buf \U$47936 ( \47911 , \47910 );
xor \U$47937 ( \47912 , \47897 , \47911 );
buf \U$47938 ( \47913 , \12331 );
buf \U$47939 ( \47914 , RIc0da828_107);
buf \U$47940 ( \47915 , RIc0d8d70_50);
xor \U$47941 ( \47916 , \47914 , \47915 );
buf \U$47942 ( \47917 , \47916 );
buf \U$47943 ( \47918 , \47917 );
not \U$47944 ( \47919 , \47918 );
buf \U$47945 ( \47920 , \47919 );
buf \U$47946 ( \47921 , \47920 );
or \U$47947 ( \47922 , \47913 , \47921 );
buf \U$47948 ( \47923 , \16064 );
buf \U$47949 ( \47924 , \47151 );
or \U$47950 ( \47925 , \47923 , \47924 );
nand \U$47951 ( \47926 , \47922 , \47925 );
buf \U$47952 ( \47927 , \47926 );
buf \U$47953 ( \47928 , \47927 );
and \U$47954 ( \47929 , \47912 , \47928 );
and \U$47955 ( \47930 , \47897 , \47911 );
or \U$47956 ( \47931 , \47929 , \47930 );
buf \U$47957 ( \47932 , \47931 );
buf \U$47958 ( \47933 , \47932 );
xor \U$47959 ( \47934 , \47189 , \47207 );
xor \U$47960 ( \47935 , \47934 , \47224 );
buf \U$47961 ( \47936 , \47935 );
buf \U$47962 ( \47937 , \47936 );
xor \U$47963 ( \47938 , \47933 , \47937 );
xor \U$47964 ( \47939 , \47247 , \47264 );
xor \U$47965 ( \47940 , \47939 , \47285 );
buf \U$47966 ( \47941 , \47940 );
buf \U$47967 ( \47942 , \47941 );
and \U$47968 ( \47943 , \47938 , \47942 );
and \U$47969 ( \47944 , \47933 , \47937 );
or \U$47970 ( \47945 , \47943 , \47944 );
buf \U$47971 ( \47946 , \47945 );
buf \U$47972 ( \47947 , \47946 );
xor \U$47973 ( \47948 , \47142 , \47161 );
xor \U$47974 ( \47949 , \47948 , \47179 );
buf \U$47975 ( \47950 , \47949 );
buf \U$47976 ( \47951 , \47950 );
xor \U$47977 ( \47952 , \47345 , \47362 );
xor \U$47978 ( \47953 , \47952 , \47380 );
buf \U$47979 ( \47954 , \47953 );
buf \U$47980 ( \47955 , \47954 );
xor \U$47981 ( \47956 , \47951 , \47955 );
xor \U$47982 ( \47957 , \47004 , \47022 );
xor \U$47983 ( \47958 , \47957 , \47048 );
buf \U$47984 ( \47959 , \47958 );
and \U$47985 ( \47960 , \47956 , \47959 );
and \U$47986 ( \47961 , \47951 , \47955 );
or \U$47987 ( \47962 , \47960 , \47961 );
buf \U$47988 ( \47963 , \47962 );
buf \U$47989 ( \47964 , \47963 );
xor \U$47990 ( \47965 , \47947 , \47964 );
xor \U$47991 ( \47966 , \47184 , \47229 );
xor \U$47992 ( \47967 , \47966 , \47290 );
buf \U$47993 ( \47968 , \47967 );
buf \U$47994 ( \47969 , \47968 );
and \U$47995 ( \47970 , \47965 , \47969 );
and \U$47996 ( \47971 , \47947 , \47964 );
or \U$47997 ( \47972 , \47970 , \47971 );
buf \U$47998 ( \47973 , \47972 );
buf \U$47999 ( \47974 , \47973 );
xor \U$48000 ( \47975 , \47877 , \47974 );
xor \U$48001 ( \47976 , \46985 , \47124 );
xor \U$48002 ( \47977 , \47976 , \47295 );
buf \U$48003 ( \47978 , \47977 );
buf \U$48004 ( \47979 , \47978 );
and \U$48005 ( \47980 , \47975 , \47979 );
and \U$48006 ( \47981 , \47877 , \47974 );
or \U$48007 ( \47982 , \47980 , \47981 );
buf \U$48008 ( \47983 , \47982 );
buf \U$48009 ( \47984 , \47983 );
nand \U$48010 ( \47985 , \47559 , \47984 );
buf \U$48011 ( \47986 , \47985 );
buf \U$48012 ( \47987 , \47986 );
nand \U$48013 ( \47988 , \47556 , \47987 );
buf \U$48014 ( \47989 , \47988 );
buf \U$48015 ( \47990 , \47989 );
not \U$48016 ( \47991 , \47990 );
buf \U$48017 ( \47992 , \47991 );
buf \U$48018 ( \47993 , \47992 );
nand \U$48019 ( \47994 , \47518 , \47993 );
buf \U$48020 ( \47995 , \47994 );
not \U$48021 ( \47996 , \47995 );
or \U$48022 ( \47997 , \47447 , \47996 );
buf \U$48023 ( \47998 , \47989 );
buf \U$48024 ( \47999 , \47516 );
nand \U$48025 ( \48000 , \47998 , \47999 );
buf \U$48026 ( \48001 , \48000 );
nand \U$48027 ( \48002 , \47997 , \48001 );
buf \U$48028 ( \48003 , \48002 );
not \U$48029 ( \48004 , \48003 );
buf \U$48030 ( \48005 , \46979 );
buf \U$48031 ( \48006 , \47428 );
xor \U$48032 ( \48007 , \48005 , \48006 );
buf \U$48033 ( \48008 , \46975 );
xnor \U$48034 ( \48009 , \48007 , \48008 );
buf \U$48035 ( \48010 , \48009 );
buf \U$48036 ( \48011 , \48010 );
nand \U$48037 ( \48012 , \48004 , \48011 );
buf \U$48038 ( \48013 , \48012 );
buf \U$48039 ( \48014 , \48013 );
buf \U$48040 ( \48015 , \46503 );
not \U$48041 ( \48016 , \48015 );
buf \U$48042 ( \48017 , \46487 );
not \U$48043 ( \48018 , \48017 );
or \U$48044 ( \48019 , \48016 , \48018 );
buf \U$48045 ( \48020 , \46487 );
buf \U$48046 ( \48021 , \46503 );
or \U$48047 ( \48022 , \48020 , \48021 );
buf \U$48048 ( \48023 , \46477 );
nand \U$48049 ( \48024 , \48022 , \48023 );
buf \U$48050 ( \48025 , \48024 );
buf \U$48051 ( \48026 , \48025 );
nand \U$48052 ( \48027 , \48019 , \48026 );
buf \U$48053 ( \48028 , \48027 );
xor \U$48054 ( \48029 , \46776 , \46790 );
and \U$48055 ( \48030 , \48029 , \46805 );
and \U$48056 ( \48031 , \46776 , \46790 );
or \U$48057 ( \48032 , \48030 , \48031 );
buf \U$48058 ( \48033 , \48032 );
xor \U$48059 ( \48034 , \46817 , \46831 );
and \U$48060 ( \48035 , \48034 , \46848 );
and \U$48061 ( \48036 , \46817 , \46831 );
or \U$48062 ( \48037 , \48035 , \48036 );
buf \U$48063 ( \48038 , \48037 );
xor \U$48064 ( \48039 , \48033 , \48038 );
buf \U$48065 ( \48040 , \48039 );
buf \U$48066 ( \48041 , \46736 );
not \U$48067 ( \48042 , \48041 );
buf \U$48068 ( \48043 , \3415 );
not \U$48069 ( \48044 , \48043 );
or \U$48070 ( \48045 , \48042 , \48044 );
buf \U$48071 ( \48046 , \4008 );
xor \U$48072 ( \48047 , RIc0da198_93, RIc0d8fc8_55);
buf \U$48073 ( \48048 , \48047 );
nand \U$48074 ( \48049 , \48046 , \48048 );
buf \U$48075 ( \48050 , \48049 );
buf \U$48076 ( \48051 , \48050 );
nand \U$48077 ( \48052 , \48045 , \48051 );
buf \U$48078 ( \48053 , \48052 );
buf \U$48079 ( \48054 , \46629 );
not \U$48080 ( \48055 , \48054 );
buf \U$48081 ( \48056 , \25475 );
not \U$48082 ( \48057 , \48056 );
or \U$48083 ( \48058 , \48055 , \48057 );
buf \U$48084 ( \48059 , \12744 );
buf \U$48085 ( \48060 , RIc0da738_105);
buf \U$48086 ( \48061 , RIc0d8a28_43);
xor \U$48087 ( \48062 , \48060 , \48061 );
buf \U$48088 ( \48063 , \48062 );
buf \U$48089 ( \48064 , \48063 );
nand \U$48090 ( \48065 , \48059 , \48064 );
buf \U$48091 ( \48066 , \48065 );
buf \U$48092 ( \48067 , \48066 );
nand \U$48093 ( \48068 , \48058 , \48067 );
buf \U$48094 ( \48069 , \48068 );
xor \U$48095 ( \48070 , \48053 , \48069 );
buf \U$48096 ( \48071 , \46467 );
not \U$48097 ( \48072 , \48071 );
buf \U$48098 ( \48073 , \13460 );
not \U$48099 ( \48074 , \48073 );
or \U$48100 ( \48075 , \48072 , \48074 );
buf \U$48101 ( \48076 , RIc0db098_125);
buf \U$48102 ( \48077 , RIc0d80c8_23);
xnor \U$48103 ( \48078 , \48076 , \48077 );
buf \U$48104 ( \48079 , \48078 );
buf \U$48105 ( \48080 , \48079 );
not \U$48106 ( \48081 , \48080 );
buf \U$48107 ( \48082 , \15793 );
nand \U$48108 ( \48083 , \48081 , \48082 );
buf \U$48109 ( \48084 , \48083 );
buf \U$48110 ( \48085 , \48084 );
nand \U$48111 ( \48086 , \48075 , \48085 );
buf \U$48112 ( \48087 , \48086 );
xnor \U$48113 ( \48088 , \48070 , \48087 );
buf \U$48114 ( \48089 , \48088 );
not \U$48115 ( \48090 , \48089 );
buf \U$48116 ( \48091 , \48090 );
buf \U$48117 ( \48092 , \48091 );
and \U$48118 ( \48093 , \48040 , \48092 );
not \U$48119 ( \48094 , \48040 );
buf \U$48120 ( \48095 , \48088 );
and \U$48121 ( \48096 , \48094 , \48095 );
nor \U$48122 ( \48097 , \48093 , \48096 );
buf \U$48123 ( \48098 , \48097 );
xor \U$48124 ( \48099 , \48028 , \48098 );
xor \U$48125 ( \48100 , \46808 , \46851 );
and \U$48126 ( \48101 , \48100 , \46907 );
and \U$48127 ( \48102 , \46808 , \46851 );
or \U$48128 ( \48103 , \48101 , \48102 );
buf \U$48129 ( \48104 , \48103 );
xor \U$48130 ( \48105 , \48099 , \48104 );
buf \U$48131 ( \48106 , \48105 );
xor \U$48132 ( \48107 , \46910 , \46916 );
and \U$48133 ( \48108 , \48107 , \46960 );
and \U$48134 ( \48109 , \46910 , \46916 );
or \U$48135 ( \48110 , \48108 , \48109 );
buf \U$48136 ( \48111 , \48110 );
buf \U$48137 ( \48112 , \48111 );
xor \U$48138 ( \48113 , \48106 , \48112 );
buf \U$48139 ( \48114 , \26411 );
not \U$48140 ( \48115 , \48114 );
buf \U$48141 ( \48116 , RIc0d9dd8_85);
buf \U$48142 ( \48117 , \43843 );
and \U$48143 ( \48118 , \48116 , \48117 );
not \U$48144 ( \48119 , \48116 );
buf \U$48145 ( \48120 , RIc0d9400_64);
and \U$48146 ( \48121 , \48119 , \48120 );
nor \U$48147 ( \48122 , \48118 , \48121 );
buf \U$48148 ( \48123 , \48122 );
buf \U$48149 ( \48124 , \48123 );
not \U$48150 ( \48125 , \48124 );
and \U$48151 ( \48126 , \48115 , \48125 );
buf \U$48152 ( \48127 , \2960 );
buf \U$48153 ( \48128 , RIc0d9dd8_85);
buf \U$48154 ( \48129 , RIc0d9388_63);
xor \U$48155 ( \48130 , \48128 , \48129 );
buf \U$48156 ( \48131 , \48130 );
buf \U$48157 ( \48132 , \48131 );
and \U$48158 ( \48133 , \48127 , \48132 );
nor \U$48159 ( \48134 , \48126 , \48133 );
buf \U$48160 ( \48135 , \48134 );
buf \U$48161 ( \48136 , \46824 );
not \U$48162 ( \48137 , \48136 );
buf \U$48163 ( \48138 , \12529 );
not \U$48164 ( \48139 , \48138 );
or \U$48165 ( \48140 , \48137 , \48139 );
buf \U$48166 ( \48141 , \14353 );
buf \U$48167 ( \48142 , RIc0daa08_111);
buf \U$48168 ( \48143 , RIc0d8758_37);
xor \U$48169 ( \48144 , \48142 , \48143 );
buf \U$48170 ( \48145 , \48144 );
buf \U$48171 ( \48146 , \48145 );
nand \U$48172 ( \48147 , \48141 , \48146 );
buf \U$48173 ( \48148 , \48147 );
buf \U$48174 ( \48149 , \48148 );
nand \U$48175 ( \48150 , \48140 , \48149 );
buf \U$48176 ( \48151 , \48150 );
buf \U$48177 ( \48152 , \48151 );
not \U$48178 ( \48153 , \48152 );
buf \U$48179 ( \48154 , \48153 );
xor \U$48180 ( \48155 , \48135 , \48154 );
buf \U$48181 ( \48156 , \46448 );
not \U$48182 ( \48157 , \48156 );
buf \U$48183 ( \48158 , \22350 );
not \U$48184 ( \48159 , \48158 );
or \U$48185 ( \48160 , \48157 , \48159 );
buf \U$48186 ( \48161 , \22356 );
xor \U$48187 ( \48162 , RIc0dacd8_117, RIc0d8488_31);
buf \U$48188 ( \48163 , \48162 );
nand \U$48189 ( \48164 , \48161 , \48163 );
buf \U$48190 ( \48165 , \48164 );
buf \U$48191 ( \48166 , \48165 );
nand \U$48192 ( \48167 , \48160 , \48166 );
buf \U$48193 ( \48168 , \48167 );
xor \U$48194 ( \48169 , \48155 , \48168 );
buf \U$48195 ( \48170 , \48169 );
not \U$48196 ( \48171 , \48170 );
buf \U$48197 ( \48172 , \46754 );
not \U$48198 ( \48173 , \48172 );
buf \U$48199 ( \48174 , \25542 );
not \U$48200 ( \48175 , \48174 );
or \U$48201 ( \48176 , \48173 , \48175 );
buf \U$48202 ( \48177 , \13005 );
buf \U$48203 ( \48178 , RIc0dadc8_119);
buf \U$48204 ( \48179 , RIc0d8398_29);
xor \U$48205 ( \48180 , \48178 , \48179 );
buf \U$48206 ( \48181 , \48180 );
buf \U$48207 ( \48182 , \48181 );
nand \U$48208 ( \48183 , \48177 , \48182 );
buf \U$48209 ( \48184 , \48183 );
buf \U$48210 ( \48185 , \48184 );
nand \U$48211 ( \48186 , \48176 , \48185 );
buf \U$48212 ( \48187 , \48186 );
buf \U$48213 ( \48188 , \48187 );
not \U$48214 ( \48189 , \48188 );
buf \U$48215 ( \48190 , \48189 );
buf \U$48216 ( \48191 , \46384 );
not \U$48217 ( \48192 , \48191 );
buf \U$48218 ( \48193 , \14210 );
not \U$48219 ( \48194 , \48193 );
or \U$48220 ( \48195 , \48192 , \48194 );
buf \U$48221 ( \48196 , \20211 );
xor \U$48222 ( \48197 , RIc0da918_109, RIc0d8848_39);
buf \U$48223 ( \48198 , \48197 );
nand \U$48224 ( \48199 , \48196 , \48198 );
buf \U$48225 ( \48200 , \48199 );
buf \U$48226 ( \48201 , \48200 );
nand \U$48227 ( \48202 , \48195 , \48201 );
buf \U$48228 ( \48203 , \48202 );
xor \U$48229 ( \48204 , \48190 , \48203 );
buf \U$48230 ( \48205 , \46899 );
not \U$48231 ( \48206 , \48205 );
buf \U$48232 ( \48207 , \3714 );
not \U$48233 ( \48208 , \48207 );
or \U$48234 ( \48209 , \48206 , \48208 );
buf \U$48235 ( \48210 , \344 );
buf \U$48236 ( \48211 , RIc0da288_95);
buf \U$48237 ( \48212 , RIc0d8ed8_53);
xor \U$48238 ( \48213 , \48211 , \48212 );
buf \U$48239 ( \48214 , \48213 );
buf \U$48240 ( \48215 , \48214 );
nand \U$48241 ( \48216 , \48210 , \48215 );
buf \U$48242 ( \48217 , \48216 );
buf \U$48243 ( \48218 , \48217 );
nand \U$48244 ( \48219 , \48209 , \48218 );
buf \U$48245 ( \48220 , \48219 );
xor \U$48246 ( \48221 , \48204 , \48220 );
buf \U$48247 ( \48222 , \48221 );
not \U$48248 ( \48223 , \48222 );
or \U$48249 ( \48224 , \48171 , \48223 );
buf \U$48250 ( \48225 , \48221 );
not \U$48251 ( \48226 , \48225 );
buf \U$48252 ( \48227 , \48226 );
buf \U$48253 ( \48228 , \48227 );
buf \U$48254 ( \48229 , \48169 );
not \U$48255 ( \48230 , \48229 );
buf \U$48256 ( \48231 , \48230 );
buf \U$48257 ( \48232 , \48231 );
nand \U$48258 ( \48233 , \48228 , \48232 );
buf \U$48259 ( \48234 , \48233 );
buf \U$48260 ( \48235 , \48234 );
nand \U$48261 ( \48236 , \48224 , \48235 );
buf \U$48262 ( \48237 , \48236 );
buf \U$48263 ( \48238 , \48237 );
buf \U$48264 ( \48239 , \46809 );
not \U$48265 ( \48240 , \48239 );
buf \U$48266 ( \48241 , \15609 );
not \U$48267 ( \48242 , \48241 );
or \U$48268 ( \48243 , \48240 , \48242 );
buf \U$48269 ( \48244 , RIc0d7fd8_21);
buf \U$48270 ( \48245 , RIc0db188_127);
xor \U$48271 ( \48246 , \48244 , \48245 );
buf \U$48272 ( \48247 , \48246 );
buf \U$48273 ( \48248 , \48247 );
buf \U$48274 ( \48249 , RIc0db200_128);
nand \U$48275 ( \48250 , \48248 , \48249 );
buf \U$48276 ( \48251 , \48250 );
buf \U$48277 ( \48252 , \48251 );
nand \U$48278 ( \48253 , \48243 , \48252 );
buf \U$48279 ( \48254 , \48253 );
buf \U$48280 ( \48255 , \48254 );
buf \U$48281 ( \48256 , \46798 );
not \U$48282 ( \48257 , \48256 );
buf \U$48283 ( \48258 , \33224 );
not \U$48284 ( \48259 , \48258 );
or \U$48285 ( \48260 , \48257 , \48259 );
buf \U$48286 ( \48261 , RIc0daaf8_113);
buf \U$48287 ( \48262 , RIc0d8668_35);
xnor \U$48288 ( \48263 , \48261 , \48262 );
buf \U$48289 ( \48264 , \48263 );
buf \U$48290 ( \48265 , \48264 );
not \U$48291 ( \48266 , \48265 );
buf \U$48292 ( \48267 , \12410 );
nand \U$48293 ( \48268 , \48266 , \48267 );
buf \U$48294 ( \48269 , \48268 );
buf \U$48295 ( \48270 , \48269 );
nand \U$48296 ( \48271 , \48260 , \48270 );
buf \U$48297 ( \48272 , \48271 );
buf \U$48298 ( \48273 , \48272 );
xor \U$48299 ( \48274 , \48255 , \48273 );
buf \U$48300 ( \48275 , \46683 );
not \U$48301 ( \48276 , \48275 );
buf \U$48302 ( \48277 , \25371 );
not \U$48303 ( \48278 , \48277 );
or \U$48304 ( \48279 , \48276 , \48278 );
buf \U$48305 ( \48280 , \14648 );
buf \U$48306 ( \48281 , RIc0da468_99);
buf \U$48307 ( \48282 , RIc0d8cf8_49);
xor \U$48308 ( \48283 , \48281 , \48282 );
buf \U$48309 ( \48284 , \48283 );
buf \U$48310 ( \48285 , \48284 );
nand \U$48311 ( \48286 , \48280 , \48285 );
buf \U$48312 ( \48287 , \48286 );
buf \U$48313 ( \48288 , \48287 );
nand \U$48314 ( \48289 , \48279 , \48288 );
buf \U$48315 ( \48290 , \48289 );
buf \U$48316 ( \48291 , \48290 );
xnor \U$48317 ( \48292 , \48274 , \48291 );
buf \U$48318 ( \48293 , \48292 );
buf \U$48319 ( \48294 , \48293 );
not \U$48320 ( \48295 , \48294 );
buf \U$48321 ( \48296 , \48295 );
buf \U$48322 ( \48297 , \48296 );
and \U$48323 ( \48298 , \48238 , \48297 );
not \U$48324 ( \48299 , \48238 );
buf \U$48325 ( \48300 , \48293 );
and \U$48326 ( \48301 , \48299 , \48300 );
nor \U$48327 ( \48302 , \48298 , \48301 );
buf \U$48328 ( \48303 , \48302 );
buf \U$48329 ( \48304 , \48303 );
xor \U$48330 ( \48305 , \46935 , \46950 );
and \U$48331 ( \48306 , \48305 , \46957 );
and \U$48332 ( \48307 , \46935 , \46950 );
or \U$48333 ( \48308 , \48306 , \48307 );
buf \U$48334 ( \48309 , \48308 );
buf \U$48335 ( \48310 , \48309 );
xor \U$48336 ( \48311 , \48304 , \48310 );
xor \U$48337 ( \48312 , \46391 , \46394 );
and \U$48338 ( \48313 , \48312 , \46410 );
and \U$48339 ( \48314 , \46391 , \46394 );
or \U$48340 ( \48315 , \48313 , \48314 );
buf \U$48341 ( \48316 , \48315 );
buf \U$48342 ( \48317 , \48316 );
xor \U$48343 ( \48318 , \46570 , \46576 );
and \U$48344 ( \48319 , \48318 , \46583 );
and \U$48345 ( \48320 , \46570 , \46576 );
or \U$48346 ( \48321 , \48319 , \48320 );
buf \U$48347 ( \48322 , \48321 );
buf \U$48348 ( \48323 , \48322 );
xor \U$48349 ( \48324 , \48317 , \48323 );
xor \U$48350 ( \48325 , \46657 , \46708 );
and \U$48351 ( \48326 , \48325 , \46764 );
and \U$48352 ( \48327 , \46657 , \46708 );
or \U$48353 ( \48328 , \48326 , \48327 );
buf \U$48354 ( \48329 , \48328 );
buf \U$48355 ( \48330 , \48329 );
xor \U$48356 ( \48331 , \48324 , \48330 );
buf \U$48357 ( \48332 , \48331 );
buf \U$48358 ( \48333 , \48332 );
xor \U$48359 ( \48334 , \48311 , \48333 );
buf \U$48360 ( \48335 , \48334 );
buf \U$48361 ( \48336 , \48335 );
xor \U$48362 ( \48337 , \48113 , \48336 );
buf \U$48363 ( \48338 , \48337 );
buf \U$48364 ( \48339 , \48338 );
xor \U$48365 ( \48340 , \46352 , \46529 );
and \U$48366 ( \48341 , \48340 , \46966 );
and \U$48367 ( \48342 , \46352 , \46529 );
or \U$48368 ( \48343 , \48341 , \48342 );
buf \U$48369 ( \48344 , \48343 );
buf \U$48370 ( \48345 , \48344 );
xor \U$48371 ( \48346 , \48339 , \48345 );
xor \U$48372 ( \48347 , \46367 , \46373 );
and \U$48373 ( \48348 , \48347 , \46526 );
and \U$48374 ( \48349 , \46367 , \46373 );
or \U$48375 ( \48350 , \48348 , \48349 );
buf \U$48376 ( \48351 , \48350 );
buf \U$48377 ( \48352 , \48351 );
xor \U$48378 ( \48353 , \46413 , \46419 );
and \U$48379 ( \48354 , \48353 , \46523 );
and \U$48380 ( \48355 , \46413 , \46419 );
or \U$48381 ( \48356 , \48354 , \48355 );
buf \U$48382 ( \48357 , \48356 );
buf \U$48383 ( \48358 , \48357 );
buf \U$48384 ( \48359 , \46595 );
not \U$48385 ( \48360 , \48359 );
buf \U$48386 ( \48361 , \46588 );
not \U$48387 ( \48362 , \48361 );
or \U$48388 ( \48363 , \48360 , \48362 );
buf \U$48389 ( \48364 , \46766 );
nand \U$48390 ( \48365 , \48363 , \48364 );
buf \U$48391 ( \48366 , \48365 );
buf \U$48392 ( \48367 , \48366 );
buf \U$48393 ( \48368 , \46585 );
buf \U$48394 ( \48369 , \46553 );
nand \U$48395 ( \48370 , \48368 , \48369 );
buf \U$48396 ( \48371 , \48370 );
buf \U$48397 ( \48372 , \48371 );
nand \U$48398 ( \48373 , \48367 , \48372 );
buf \U$48399 ( \48374 , \48373 );
buf \U$48400 ( \48375 , \48374 );
xor \U$48401 ( \48376 , \48358 , \48375 );
buf \U$48402 ( \48377 , \46843 );
not \U$48403 ( \48378 , \48377 );
buf \U$48404 ( \48379 , \48378 );
buf \U$48405 ( \48380 , \48379 );
not \U$48406 ( \48381 , \48380 );
buf \U$48407 ( \48382 , \19487 );
not \U$48408 ( \48383 , \48382 );
or \U$48409 ( \48384 , \48381 , \48383 );
buf \U$48410 ( \48385 , \13314 );
buf \U$48411 ( \48386 , RIc0daeb8_121);
buf \U$48412 ( \48387 , RIc0d82a8_27);
xor \U$48413 ( \48388 , \48386 , \48387 );
buf \U$48414 ( \48389 , \48388 );
buf \U$48415 ( \48390 , \48389 );
nand \U$48416 ( \48391 , \48385 , \48390 );
buf \U$48417 ( \48392 , \48391 );
buf \U$48418 ( \48393 , \48392 );
nand \U$48419 ( \48394 , \48384 , \48393 );
buf \U$48420 ( \48395 , \48394 );
buf \U$48421 ( \48396 , \46667 );
not \U$48422 ( \48397 , \48396 );
buf \U$48423 ( \48398 , \2066 );
not \U$48424 ( \48399 , \48398 );
or \U$48425 ( \48400 , \48397 , \48399 );
buf \U$48426 ( \48401 , \734 );
xor \U$48427 ( \48402 , RIc0da378_97, RIc0d8de8_51);
buf \U$48428 ( \48403 , \48402 );
nand \U$48429 ( \48404 , \48401 , \48403 );
buf \U$48430 ( \48405 , \48404 );
buf \U$48431 ( \48406 , \48405 );
nand \U$48432 ( \48407 , \48400 , \48406 );
buf \U$48433 ( \48408 , \48407 );
xor \U$48434 ( \48409 , \48395 , \48408 );
buf \U$48435 ( \48410 , \48409 );
buf \U$48436 ( \48411 , \46862 );
not \U$48437 ( \48412 , \48411 );
buf \U$48438 ( \48413 , \4042 );
not \U$48439 ( \48414 , \48413 );
or \U$48440 ( \48415 , \48412 , \48414 );
buf \U$48441 ( \48416 , \12839 );
xor \U$48442 ( \48417 , RIc0da558_101, RIc0d8c08_47);
buf \U$48443 ( \48418 , \48417 );
nand \U$48444 ( \48419 , \48416 , \48418 );
buf \U$48445 ( \48420 , \48419 );
buf \U$48446 ( \48421 , \48420 );
nand \U$48447 ( \48422 , \48415 , \48421 );
buf \U$48448 ( \48423 , \48422 );
buf \U$48449 ( \48424 , \48423 );
xnor \U$48450 ( \48425 , \48410 , \48424 );
buf \U$48451 ( \48426 , \48425 );
buf \U$48452 ( \48427 , \48426 );
not \U$48453 ( \48428 , \48427 );
buf \U$48454 ( \48429 , \46612 );
not \U$48455 ( \48430 , \48429 );
buf \U$48456 ( \48431 , \2535 );
not \U$48457 ( \48432 , \48431 );
or \U$48458 ( \48433 , \48430 , \48432 );
buf \U$48459 ( \48434 , \13293 );
buf \U$48460 ( \48435 , RIc0da0a8_91);
buf \U$48461 ( \48436 , RIc0d90b8_57);
xor \U$48462 ( \48437 , \48435 , \48436 );
buf \U$48463 ( \48438 , \48437 );
buf \U$48464 ( \48439 , \48438 );
nand \U$48465 ( \48440 , \48434 , \48439 );
buf \U$48466 ( \48441 , \48440 );
buf \U$48467 ( \48442 , \48441 );
nand \U$48468 ( \48443 , \48433 , \48442 );
buf \U$48469 ( \48444 , \48443 );
buf \U$48470 ( \48445 , \48444 );
buf \U$48471 ( \48446 , \46783 );
not \U$48472 ( \48447 , \48446 );
buf \U$48473 ( \48448 , \2038 );
not \U$48474 ( \48449 , \48448 );
or \U$48475 ( \48450 , \48447 , \48449 );
buf \U$48476 ( \48451 , \846 );
buf \U$48477 ( \48452 , RIc0d91a8_59);
buf \U$48478 ( \48453 , RIc0d9fb8_89);
xor \U$48479 ( \48454 , \48452 , \48453 );
buf \U$48480 ( \48455 , \48454 );
buf \U$48481 ( \48456 , \48455 );
nand \U$48482 ( \48457 , \48451 , \48456 );
buf \U$48483 ( \48458 , \48457 );
buf \U$48484 ( \48459 , \48458 );
nand \U$48485 ( \48460 , \48450 , \48459 );
buf \U$48486 ( \48461 , \48460 );
buf \U$48487 ( \48462 , \48461 );
xor \U$48488 ( \48463 , \48445 , \48462 );
buf \U$48489 ( \48464 , \4483 );
buf \U$48490 ( \48465 , \46429 );
or \U$48491 ( \48466 , \48464 , \48465 );
buf \U$48492 ( \48467 , \4475 );
buf \U$48493 ( \48468 , RIc0d8b18_45);
buf \U$48494 ( \48469 , RIc0da648_103);
xnor \U$48495 ( \48470 , \48468 , \48469 );
buf \U$48496 ( \48471 , \48470 );
buf \U$48497 ( \48472 , \48471 );
or \U$48498 ( \48473 , \48467 , \48472 );
nand \U$48499 ( \48474 , \48466 , \48473 );
buf \U$48500 ( \48475 , \48474 );
buf \U$48501 ( \48476 , \48475 );
xor \U$48502 ( \48477 , \48463 , \48476 );
buf \U$48503 ( \48478 , \48477 );
buf \U$48504 ( \48479 , \48478 );
not \U$48505 ( \48480 , \48479 );
or \U$48506 ( \48481 , \48428 , \48480 );
buf \U$48507 ( \48482 , \48478 );
not \U$48508 ( \48483 , \48482 );
buf \U$48509 ( \48484 , \48426 );
not \U$48510 ( \48485 , \48484 );
buf \U$48511 ( \48486 , \48485 );
buf \U$48512 ( \48487 , \48486 );
nand \U$48513 ( \48488 , \48483 , \48487 );
buf \U$48514 ( \48489 , \48488 );
buf \U$48515 ( \48490 , \48489 );
nand \U$48516 ( \48491 , \48481 , \48490 );
buf \U$48517 ( \48492 , \48491 );
buf \U$48518 ( \48493 , \48492 );
buf \U$48519 ( \48494 , \46647 );
not \U$48520 ( \48495 , \48494 );
buf \U$48521 ( \48496 , \34202 );
not \U$48522 ( \48497 , \48496 );
or \U$48523 ( \48498 , \48495 , \48497 );
buf \U$48524 ( \48499 , \12342 );
buf \U$48525 ( \48500 , RIc0d8938_41);
buf \U$48526 ( \48501 , RIc0da828_107);
xor \U$48527 ( \48502 , \48500 , \48501 );
buf \U$48528 ( \48503 , \48502 );
buf \U$48529 ( \48504 , \48503 );
nand \U$48530 ( \48505 , \48499 , \48504 );
buf \U$48531 ( \48506 , \48505 );
buf \U$48532 ( \48507 , \48506 );
nand \U$48533 ( \48508 , \48498 , \48507 );
buf \U$48534 ( \48509 , \48508 );
buf \U$48535 ( \48510 , \48509 );
buf \U$48536 ( \48511 , \14681 );
not \U$48537 ( \48512 , \48511 );
buf \U$48538 ( \48513 , \46880 );
not \U$48539 ( \48514 , \48513 );
and \U$48540 ( \48515 , \48512 , \48514 );
buf \U$48541 ( \48516 , \29865 );
buf \U$48542 ( \48517 , RIc0dabe8_115);
buf \U$48543 ( \48518 , RIc0d8578_33);
xnor \U$48544 ( \48519 , \48517 , \48518 );
buf \U$48545 ( \48520 , \48519 );
buf \U$48546 ( \48521 , \48520 );
nor \U$48547 ( \48522 , \48516 , \48521 );
buf \U$48548 ( \48523 , \48522 );
buf \U$48549 ( \48524 , \48523 );
nor \U$48550 ( \48525 , \48515 , \48524 );
buf \U$48551 ( \48526 , \48525 );
buf \U$48552 ( \48527 , \48526 );
not \U$48553 ( \48528 , \48527 );
buf \U$48554 ( \48529 , \46700 );
not \U$48555 ( \48530 , \48529 );
buf \U$48556 ( \48531 , \14982 );
not \U$48557 ( \48532 , \48531 );
or \U$48558 ( \48533 , \48530 , \48532 );
buf \U$48559 ( \48534 , \16692 );
xor \U$48560 ( \48535 , RIc0dafa8_123, RIc0d81b8_25);
buf \U$48561 ( \48536 , \48535 );
nand \U$48562 ( \48537 , \48534 , \48536 );
buf \U$48563 ( \48538 , \48537 );
buf \U$48564 ( \48539 , \48538 );
nand \U$48565 ( \48540 , \48533 , \48539 );
buf \U$48566 ( \48541 , \48540 );
buf \U$48567 ( \48542 , \48541 );
not \U$48568 ( \48543 , \48542 );
or \U$48569 ( \48544 , \48528 , \48543 );
buf \U$48570 ( \48545 , \48541 );
buf \U$48571 ( \48546 , \48526 );
or \U$48572 ( \48547 , \48545 , \48546 );
nand \U$48573 ( \48548 , \48544 , \48547 );
buf \U$48574 ( \48549 , \48548 );
buf \U$48575 ( \48550 , \48549 );
xnor \U$48576 ( \48551 , \48510 , \48550 );
buf \U$48577 ( \48552 , \48551 );
buf \U$48578 ( \48553 , \48552 );
not \U$48579 ( \48554 , \48553 );
buf \U$48580 ( \48555 , \48554 );
buf \U$48581 ( \48556 , \48555 );
and \U$48582 ( \48557 , \48493 , \48556 );
not \U$48583 ( \48558 , \48493 );
buf \U$48584 ( \48559 , \48552 );
and \U$48585 ( \48560 , \48558 , \48559 );
nor \U$48586 ( \48561 , \48557 , \48560 );
buf \U$48587 ( \48562 , \48561 );
buf \U$48588 ( \48563 , \48562 );
not \U$48589 ( \48564 , \48563 );
buf \U$48590 ( \48565 , \48564 );
buf \U$48591 ( \48566 , \48565 );
not \U$48592 ( \48567 , \48566 );
buf \U$48593 ( \48568 , \6270 );
buf \U$48594 ( \48569 , \46719 );
not \U$48595 ( \48570 , \48569 );
buf \U$48596 ( \48571 , \48570 );
buf \U$48597 ( \48572 , \48571 );
or \U$48598 ( \48573 , \48568 , \48572 );
buf \U$48599 ( \48574 , \634 );
buf \U$48600 ( \48575 , RIc0d9298_61);
buf \U$48601 ( \48576 , RIc0d9ec8_87);
xor \U$48602 ( \48577 , \48575 , \48576 );
buf \U$48603 ( \48578 , \48577 );
buf \U$48604 ( \48579 , \48578 );
not \U$48605 ( \48580 , \48579 );
buf \U$48606 ( \48581 , \48580 );
buf \U$48607 ( \48582 , \48581 );
or \U$48608 ( \48583 , \48574 , \48582 );
nand \U$48609 ( \48584 , \48573 , \48583 );
buf \U$48610 ( \48585 , \48584 );
buf \U$48611 ( \48586 , RIc0d9400_64);
buf \U$48612 ( \48587 , RIc0d9e50_86);
or \U$48613 ( \48588 , \48586 , \48587 );
buf \U$48614 ( \48589 , RIc0d9ec8_87);
nand \U$48615 ( \48590 , \48588 , \48589 );
buf \U$48616 ( \48591 , \48590 );
buf \U$48617 ( \48592 , \48591 );
buf \U$48618 ( \48593 , RIc0d9400_64);
buf \U$48619 ( \48594 , RIc0d9e50_86);
nand \U$48620 ( \48595 , \48593 , \48594 );
buf \U$48621 ( \48596 , \48595 );
buf \U$48622 ( \48597 , \48596 );
buf \U$48623 ( \48598 , RIc0d9dd8_85);
nand \U$48624 ( \48599 , \48592 , \48597 , \48598 );
buf \U$48625 ( \48600 , \48599 );
xor \U$48626 ( \48601 , \48585 , \48600 );
buf \U$48627 ( \48602 , \48601 );
not \U$48628 ( \48603 , \48602 );
xor \U$48629 ( \48604 , \46673 , \46689 );
and \U$48630 ( \48605 , \48604 , \46706 );
and \U$48631 ( \48606 , \46673 , \46689 );
or \U$48632 ( \48607 , \48605 , \48606 );
buf \U$48633 ( \48608 , \48607 );
not \U$48634 ( \48609 , \48608 );
or \U$48635 ( \48610 , \48603 , \48609 );
buf \U$48636 ( \48611 , \48607 );
buf \U$48637 ( \48612 , \48601 );
or \U$48638 ( \48613 , \48611 , \48612 );
nand \U$48639 ( \48614 , \48610 , \48613 );
buf \U$48640 ( \48615 , \48614 );
buf \U$48641 ( \48616 , \48615 );
not \U$48642 ( \48617 , \48616 );
xor \U$48643 ( \48618 , \46438 , \46455 );
and \U$48644 ( \48619 , \48618 , \46475 );
and \U$48645 ( \48620 , \46438 , \46455 );
or \U$48646 ( \48621 , \48619 , \48620 );
buf \U$48647 ( \48622 , \48621 );
buf \U$48648 ( \48623 , \48622 );
not \U$48649 ( \48624 , \48623 );
buf \U$48650 ( \48625 , \48624 );
buf \U$48651 ( \48626 , \48625 );
not \U$48652 ( \48627 , \48626 );
and \U$48653 ( \48628 , \48617 , \48627 );
buf \U$48654 ( \48629 , \48615 );
buf \U$48655 ( \48630 , \48625 );
and \U$48656 ( \48631 , \48629 , \48630 );
nor \U$48657 ( \48632 , \48628 , \48631 );
buf \U$48658 ( \48633 , \48632 );
buf \U$48659 ( \48634 , \48633 );
not \U$48660 ( \48635 , \48634 );
xor \U$48661 ( \48636 , \46619 , \46636 );
and \U$48662 ( \48637 , \48636 , \46654 );
and \U$48663 ( \48638 , \46619 , \46636 );
or \U$48664 ( \48639 , \48637 , \48638 );
buf \U$48665 ( \48640 , \48639 );
buf \U$48666 ( \48641 , \48640 );
not \U$48667 ( \48642 , \48641 );
buf \U$48668 ( \48643 , \46905 );
buf \U$48669 ( \48644 , \46868 );
or \U$48670 ( \48645 , \48643 , \48644 );
buf \U$48671 ( \48646 , \46888 );
nand \U$48672 ( \48647 , \48645 , \48646 );
buf \U$48673 ( \48648 , \48647 );
buf \U$48674 ( \48649 , \48648 );
buf \U$48675 ( \48650 , \46905 );
buf \U$48676 ( \48651 , \46868 );
nand \U$48677 ( \48652 , \48650 , \48651 );
buf \U$48678 ( \48653 , \48652 );
buf \U$48679 ( \48654 , \48653 );
nand \U$48680 ( \48655 , \48649 , \48654 );
buf \U$48681 ( \48656 , \48655 );
buf \U$48682 ( \48657 , \48656 );
not \U$48683 ( \48658 , \48657 );
buf \U$48684 ( \48659 , \48658 );
buf \U$48685 ( \48660 , \48659 );
not \U$48686 ( \48661 , \48660 );
and \U$48687 ( \48662 , \48642 , \48661 );
buf \U$48688 ( \48663 , \48640 );
buf \U$48689 ( \48664 , \48659 );
and \U$48690 ( \48665 , \48663 , \48664 );
nor \U$48691 ( \48666 , \48662 , \48665 );
buf \U$48692 ( \48667 , \48666 );
buf \U$48693 ( \48668 , \48667 );
xor \U$48694 ( \48669 , \46726 , \46743 );
and \U$48695 ( \48670 , \48669 , \46761 );
and \U$48696 ( \48671 , \46726 , \46743 );
or \U$48697 ( \48672 , \48670 , \48671 );
buf \U$48698 ( \48673 , \48672 );
buf \U$48699 ( \48674 , \48673 );
and \U$48700 ( \48675 , \48668 , \48674 );
not \U$48701 ( \48676 , \48668 );
buf \U$48702 ( \48677 , \48673 );
not \U$48703 ( \48678 , \48677 );
buf \U$48704 ( \48679 , \48678 );
buf \U$48705 ( \48680 , \48679 );
and \U$48706 ( \48681 , \48676 , \48680 );
nor \U$48707 ( \48682 , \48675 , \48681 );
buf \U$48708 ( \48683 , \48682 );
buf \U$48709 ( \48684 , \48683 );
not \U$48710 ( \48685 , \48684 );
buf \U$48711 ( \48686 , \48685 );
buf \U$48712 ( \48687 , \48686 );
not \U$48713 ( \48688 , \48687 );
or \U$48714 ( \48689 , \48635 , \48688 );
buf \U$48715 ( \48690 , \48686 );
buf \U$48716 ( \48691 , \48633 );
or \U$48717 ( \48692 , \48690 , \48691 );
nand \U$48718 ( \48693 , \48689 , \48692 );
buf \U$48719 ( \48694 , \48693 );
buf \U$48720 ( \48695 , \48694 );
not \U$48721 ( \48696 , \48695 );
or \U$48722 ( \48697 , \48567 , \48696 );
buf \U$48723 ( \48698 , \48694 );
buf \U$48724 ( \48699 , \48565 );
or \U$48725 ( \48700 , \48698 , \48699 );
nand \U$48726 ( \48701 , \48697 , \48700 );
buf \U$48727 ( \48702 , \48701 );
buf \U$48728 ( \48703 , \48702 );
xor \U$48729 ( \48704 , \48376 , \48703 );
buf \U$48730 ( \48705 , \48704 );
buf \U$48731 ( \48706 , \48705 );
xor \U$48732 ( \48707 , \48352 , \48706 );
xor \U$48733 ( \48708 , \46536 , \46770 );
and \U$48734 ( \48709 , \48708 , \46963 );
and \U$48735 ( \48710 , \46536 , \46770 );
or \U$48736 ( \48711 , \48709 , \48710 );
buf \U$48737 ( \48712 , \48711 );
buf \U$48738 ( \48713 , \48712 );
xor \U$48739 ( \48714 , \48707 , \48713 );
buf \U$48740 ( \48715 , \48714 );
buf \U$48741 ( \48716 , \48715 );
xor \U$48742 ( \48717 , \48346 , \48716 );
buf \U$48743 ( \48718 , \48717 );
buf \U$48744 ( \48719 , \48718 );
xor \U$48745 ( \48720 , \45467 , \46345 );
and \U$48746 ( \48721 , \48720 , \46969 );
and \U$48747 ( \48722 , \45467 , \46345 );
or \U$48748 ( \48723 , \48721 , \48722 );
buf \U$48749 ( \48724 , \48723 );
buf \U$48750 ( \48725 , \48724 );
or \U$48751 ( \48726 , \48719 , \48725 );
buf \U$48752 ( \48727 , \48726 );
buf \U$48753 ( \48728 , \48727 );
buf \U$48754 ( \48729 , \47516 );
buf \U$48755 ( \48730 , \47989 );
xor \U$48756 ( \48731 , \48729 , \48730 );
buf \U$48757 ( \48732 , \47446 );
xnor \U$48758 ( \48733 , \48731 , \48732 );
buf \U$48759 ( \48734 , \48733 );
buf \U$48760 ( \48735 , \48734 );
buf \U$48761 ( \48736 , \47496 );
buf \U$48762 ( \48737 , \47501 );
and \U$48763 ( \48738 , \48736 , \48737 );
not \U$48764 ( \48739 , \48736 );
buf \U$48765 ( \48740 , \47501 );
not \U$48766 ( \48741 , \48740 );
buf \U$48767 ( \48742 , \48741 );
buf \U$48768 ( \48743 , \48742 );
and \U$48769 ( \48744 , \48739 , \48743 );
nor \U$48770 ( \48745 , \48738 , \48744 );
buf \U$48771 ( \48746 , \48745 );
buf \U$48772 ( \48747 , \48746 );
buf \U$48773 ( \48748 , \47510 );
not \U$48774 ( \48749 , \48748 );
buf \U$48775 ( \48750 , \48749 );
buf \U$48776 ( \48751 , \48750 );
and \U$48777 ( \48752 , \48747 , \48751 );
not \U$48778 ( \48753 , \48747 );
buf \U$48779 ( \48754 , \47510 );
and \U$48780 ( \48755 , \48753 , \48754 );
nor \U$48781 ( \48756 , \48752 , \48755 );
buf \U$48782 ( \48757 , \48756 );
buf \U$48783 ( \48758 , \48757 );
xor \U$48784 ( \48759 , \47112 , \47072 );
xor \U$48785 ( \48760 , \48759 , \47090 );
buf \U$48786 ( \48761 , \48760 );
buf \U$48787 ( \48762 , RIc0d86e0_36);
buf \U$48788 ( \48763 , RIc0daeb8_121);
xor \U$48789 ( \48764 , \48762 , \48763 );
buf \U$48790 ( \48765 , \48764 );
buf \U$48791 ( \48766 , \48765 );
not \U$48792 ( \48767 , \48766 );
buf \U$48793 ( \48768 , \16382 );
not \U$48794 ( \48769 , \48768 );
or \U$48795 ( \48770 , \48767 , \48769 );
buf \U$48796 ( \48771 , \47575 );
not \U$48797 ( \48772 , \48771 );
buf \U$48798 ( \48773 , \12975 );
nand \U$48799 ( \48774 , \48772 , \48773 );
buf \U$48800 ( \48775 , \48774 );
buf \U$48801 ( \48776 , \48775 );
nand \U$48802 ( \48777 , \48770 , \48776 );
buf \U$48803 ( \48778 , \48777 );
buf \U$48804 ( \48779 , \48778 );
not \U$48805 ( \48780 , \48779 );
buf \U$48806 ( \48781 , RIc0d9130_58);
buf \U$48807 ( \48782 , RIc0da468_99);
xor \U$48808 ( \48783 , \48781 , \48782 );
buf \U$48809 ( \48784 , \48783 );
buf \U$48810 ( \48785 , \48784 );
not \U$48811 ( \48786 , \48785 );
buf \U$48812 ( \48787 , \2470 );
not \U$48813 ( \48788 , \48787 );
or \U$48814 ( \48789 , \48786 , \48788 );
buf \U$48815 ( \48790 , \14648 );
buf \U$48816 ( \48791 , \46992 );
nand \U$48817 ( \48792 , \48790 , \48791 );
buf \U$48818 ( \48793 , \48792 );
buf \U$48819 ( \48794 , \48793 );
nand \U$48820 ( \48795 , \48789 , \48794 );
buf \U$48821 ( \48796 , \48795 );
buf \U$48822 ( \48797 , \48796 );
not \U$48823 ( \48798 , \48797 );
or \U$48824 ( \48799 , \48780 , \48798 );
buf \U$48825 ( \48800 , \47610 );
not \U$48826 ( \48801 , \48800 );
buf \U$48827 ( \48802 , \47593 );
not \U$48828 ( \48803 , \48802 );
or \U$48829 ( \48804 , \48801 , \48803 );
buf \U$48830 ( \48805 , \47593 );
buf \U$48831 ( \48806 , \47610 );
or \U$48832 ( \48807 , \48805 , \48806 );
nand \U$48833 ( \48808 , \48804 , \48807 );
buf \U$48834 ( \48809 , \48808 );
buf \U$48835 ( \48810 , \48809 );
buf \U$48836 ( \48811 , \48778 );
not \U$48837 ( \48812 , \48811 );
buf \U$48838 ( \48813 , \48796 );
not \U$48839 ( \48814 , \48813 );
buf \U$48840 ( \48815 , \48814 );
buf \U$48841 ( \48816 , \48815 );
nand \U$48842 ( \48817 , \48812 , \48816 );
buf \U$48843 ( \48818 , \48817 );
buf \U$48844 ( \48819 , \48818 );
nand \U$48845 ( \48820 , \48810 , \48819 );
buf \U$48846 ( \48821 , \48820 );
buf \U$48847 ( \48822 , \48821 );
nand \U$48848 ( \48823 , \48799 , \48822 );
buf \U$48849 ( \48824 , \48823 );
buf \U$48850 ( \48825 , \48824 );
xor \U$48851 ( \48826 , \48761 , \48825 );
xor \U$48852 ( \48827 , \47580 , \47614 );
xor \U$48853 ( \48828 , \48827 , \47681 );
buf \U$48854 ( \48829 , \48828 );
buf \U$48855 ( \48830 , \48829 );
and \U$48856 ( \48831 , \48826 , \48830 );
and \U$48857 ( \48832 , \48761 , \48825 );
or \U$48858 ( \48833 , \48831 , \48832 );
buf \U$48859 ( \48834 , \48833 );
buf \U$48860 ( \48835 , \48834 );
xor \U$48861 ( \48836 , \47562 , \47686 );
xor \U$48862 ( \48837 , \48836 , \47872 );
buf \U$48863 ( \48838 , \48837 );
buf \U$48864 ( \48839 , \48838 );
xor \U$48865 ( \48840 , \48835 , \48839 );
buf \U$48866 ( \48841 , RIc0daaf8_113);
buf \U$48867 ( \48842 , RIc0d8b18_45);
xnor \U$48868 ( \48843 , \48841 , \48842 );
buf \U$48869 ( \48844 , \48843 );
buf \U$48870 ( \48845 , \48844 );
not \U$48871 ( \48846 , \48845 );
buf \U$48872 ( \48847 , \48846 );
buf \U$48873 ( \48848 , \48847 );
not \U$48874 ( \48849 , \48848 );
buf \U$48875 ( \48850 , \16656 );
not \U$48876 ( \48851 , \48850 );
or \U$48877 ( \48852 , \48849 , \48851 );
buf \U$48878 ( \48853 , \16662 );
buf \U$48879 ( \48854 , \47751 );
nand \U$48880 ( \48855 , \48853 , \48854 );
buf \U$48881 ( \48856 , \48855 );
buf \U$48882 ( \48857 , \48856 );
nand \U$48883 ( \48858 , \48852 , \48857 );
buf \U$48884 ( \48859 , \48858 );
buf \U$48885 ( \48860 , \48859 );
not \U$48886 ( \48861 , \48860 );
buf \U$48887 ( \48862 , \48861 );
buf \U$48888 ( \48863 , \48862 );
not \U$48889 ( \48864 , \48863 );
buf \U$48890 ( \48865 , \12926 );
not \U$48891 ( \48866 , \48865 );
xor \U$48892 ( \48867 , RIc0dacd8_117, RIc0d8938_41);
buf \U$48893 ( \48868 , \48867 );
not \U$48894 ( \48869 , \48868 );
buf \U$48895 ( \48870 , \48869 );
buf \U$48896 ( \48871 , \48870 );
not \U$48897 ( \48872 , \48871 );
and \U$48898 ( \48873 , \48866 , \48872 );
buf \U$48899 ( \48874 , \47898 );
not \U$48900 ( \48875 , \48874 );
buf \U$48901 ( \48876 , \16556 );
nor \U$48902 ( \48877 , \48875 , \48876 );
buf \U$48903 ( \48878 , \48877 );
buf \U$48904 ( \48879 , \48878 );
nor \U$48905 ( \48880 , \48873 , \48879 );
buf \U$48906 ( \48881 , \48880 );
buf \U$48907 ( \48882 , \48881 );
not \U$48908 ( \48883 , \48882 );
or \U$48909 ( \48884 , \48864 , \48883 );
buf \U$48910 ( \48885 , RIc0d8fc8_55);
buf \U$48911 ( \48886 , RIc0da648_103);
xor \U$48912 ( \48887 , \48885 , \48886 );
buf \U$48913 ( \48888 , \48887 );
buf \U$48914 ( \48889 , \48888 );
not \U$48915 ( \48890 , \48889 );
buf \U$48916 ( \48891 , \16578 );
not \U$48917 ( \48892 , \48891 );
or \U$48918 ( \48893 , \48890 , \48892 );
buf \U$48919 ( \48894 , \13048 );
buf \U$48920 ( \48895 , \47723 );
nand \U$48921 ( \48896 , \48894 , \48895 );
buf \U$48922 ( \48897 , \48896 );
buf \U$48923 ( \48898 , \48897 );
nand \U$48924 ( \48899 , \48893 , \48898 );
buf \U$48925 ( \48900 , \48899 );
buf \U$48926 ( \48901 , \48900 );
nand \U$48927 ( \48902 , \48884 , \48901 );
buf \U$48928 ( \48903 , \48902 );
buf \U$48929 ( \48904 , \48903 );
buf \U$48930 ( \48905 , \48881 );
not \U$48931 ( \48906 , \48905 );
buf \U$48932 ( \48907 , \48859 );
nand \U$48933 ( \48908 , \48906 , \48907 );
buf \U$48934 ( \48909 , \48908 );
buf \U$48935 ( \48910 , \48909 );
nand \U$48936 ( \48911 , \48904 , \48910 );
buf \U$48937 ( \48912 , \48911 );
buf \U$48938 ( \48913 , \48912 );
not \U$48939 ( \48914 , \48913 );
buf \U$48940 ( \48915 , RIc0da828_107);
buf \U$48941 ( \48916 , RIc0d8de8_51);
xor \U$48942 ( \48917 , \48915 , \48916 );
buf \U$48943 ( \48918 , \48917 );
buf \U$48944 ( \48919 , \48918 );
not \U$48945 ( \48920 , \48919 );
buf \U$48946 ( \48921 , \12334 );
not \U$48947 ( \48922 , \48921 );
or \U$48948 ( \48923 , \48920 , \48922 );
buf \U$48949 ( \48924 , \12342 );
buf \U$48950 ( \48925 , \47917 );
nand \U$48951 ( \48926 , \48924 , \48925 );
buf \U$48952 ( \48927 , \48926 );
buf \U$48953 ( \48928 , \48927 );
nand \U$48954 ( \48929 , \48923 , \48928 );
buf \U$48955 ( \48930 , \48929 );
xor \U$48956 ( \48931 , RIc0da288_95, RIc0d9388_63);
buf \U$48957 ( \48932 , \48931 );
not \U$48958 ( \48933 , \48932 );
buf \U$48959 ( \48934 , \330 );
not \U$48960 ( \48935 , \48934 );
or \U$48961 ( \48936 , \48933 , \48935 );
buf \U$48962 ( \48937 , \14707 );
buf \U$48963 ( \48938 , \47581 );
nand \U$48964 ( \48939 , \48937 , \48938 );
buf \U$48965 ( \48940 , \48939 );
buf \U$48966 ( \48941 , \48940 );
nand \U$48967 ( \48942 , \48936 , \48941 );
buf \U$48968 ( \48943 , \48942 );
xor \U$48969 ( \48944 , \48930 , \48943 );
buf \U$48970 ( \48945 , RIc0da558_101);
buf \U$48971 ( \48946 , RIc0d90b8_57);
xor \U$48972 ( \48947 , \48945 , \48946 );
buf \U$48973 ( \48948 , \48947 );
buf \U$48974 ( \48949 , \48948 );
not \U$48975 ( \48950 , \48949 );
buf \U$48976 ( \48951 , \3535 );
not \U$48977 ( \48952 , \48951 );
or \U$48978 ( \48953 , \48950 , \48952 );
buf \U$48979 ( \48954 , \15550 );
buf \U$48980 ( \48955 , \47814 );
nand \U$48981 ( \48956 , \48954 , \48955 );
buf \U$48982 ( \48957 , \48956 );
buf \U$48983 ( \48958 , \48957 );
nand \U$48984 ( \48959 , \48953 , \48958 );
buf \U$48985 ( \48960 , \48959 );
and \U$48986 ( \48961 , \48944 , \48960 );
and \U$48987 ( \48962 , \48930 , \48943 );
or \U$48988 ( \48963 , \48961 , \48962 );
buf \U$48989 ( \48964 , \48963 );
not \U$48990 ( \48965 , \48964 );
or \U$48991 ( \48966 , \48914 , \48965 );
buf \U$48992 ( \48967 , \48963 );
buf \U$48993 ( \48968 , \48912 );
or \U$48994 ( \48969 , \48967 , \48968 );
buf \U$48995 ( \48970 , RIc0db098_125);
buf \U$48996 ( \48971 , RIc0d8578_33);
and \U$48997 ( \48972 , \48970 , \48971 );
not \U$48998 ( \48973 , \48970 );
buf \U$48999 ( \48974 , \46159 );
and \U$49000 ( \48975 , \48973 , \48974 );
nor \U$49001 ( \48976 , \48972 , \48975 );
buf \U$49002 ( \48977 , \48976 );
buf \U$49003 ( \48978 , \48977 );
not \U$49004 ( \48979 , \48978 );
buf \U$49005 ( \48980 , \15789 );
not \U$49006 ( \48981 , \48980 );
or \U$49007 ( \48982 , \48979 , \48981 );
buf \U$49008 ( \48983 , \47793 );
not \U$49009 ( \48984 , \48983 );
buf \U$49010 ( \48985 , \15793 );
nand \U$49011 ( \48986 , \48984 , \48985 );
buf \U$49012 ( \48987 , \48986 );
buf \U$49013 ( \48988 , \48987 );
nand \U$49014 ( \48989 , \48982 , \48988 );
buf \U$49015 ( \48990 , \48989 );
buf \U$49016 ( \48991 , \48990 );
not \U$49017 ( \48992 , \48991 );
buf \U$49018 ( \48993 , RIc0d8a28_43);
buf \U$49019 ( \48994 , RIc0dabe8_115);
xor \U$49020 ( \48995 , \48993 , \48994 );
buf \U$49021 ( \48996 , \48995 );
buf \U$49022 ( \48997 , \48996 );
not \U$49023 ( \48998 , \48997 );
buf \U$49024 ( \48999 , \14186 );
not \U$49025 ( \49000 , \48999 );
or \U$49026 ( \49001 , \48998 , \49000 );
buf \U$49027 ( \49002 , \12303 );
buf \U$49028 ( \49003 , \47849 );
nand \U$49029 ( \49004 , \49002 , \49003 );
buf \U$49030 ( \49005 , \49004 );
buf \U$49031 ( \49006 , \49005 );
nand \U$49032 ( \49007 , \49001 , \49006 );
buf \U$49033 ( \49008 , \49007 );
buf \U$49034 ( \49009 , \49008 );
not \U$49035 ( \49010 , \49009 );
or \U$49036 ( \49011 , \48992 , \49010 );
buf \U$49037 ( \49012 , \49008 );
buf \U$49038 ( \49013 , \48990 );
or \U$49039 ( \49014 , \49012 , \49013 );
buf \U$49040 ( \49015 , RIc0d8668_35);
buf \U$49041 ( \49016 , RIc0dafa8_123);
xor \U$49042 ( \49017 , \49015 , \49016 );
buf \U$49043 ( \49018 , \49017 );
buf \U$49044 ( \49019 , \49018 );
not \U$49045 ( \49020 , \49019 );
buf \U$49046 ( \49021 , \14982 );
not \U$49047 ( \49022 , \49021 );
or \U$49048 ( \49023 , \49020 , \49022 );
buf \U$49049 ( \49024 , \16692 );
buf \U$49050 ( \49025 , \47657 );
nand \U$49051 ( \49026 , \49024 , \49025 );
buf \U$49052 ( \49027 , \49026 );
buf \U$49053 ( \49028 , \49027 );
nand \U$49054 ( \49029 , \49023 , \49028 );
buf \U$49055 ( \49030 , \49029 );
buf \U$49056 ( \49031 , \49030 );
nand \U$49057 ( \49032 , \49014 , \49031 );
buf \U$49058 ( \49033 , \49032 );
buf \U$49059 ( \49034 , \49033 );
nand \U$49060 ( \49035 , \49011 , \49034 );
buf \U$49061 ( \49036 , \49035 );
buf \U$49062 ( \49037 , \49036 );
nand \U$49063 ( \49038 , \48969 , \49037 );
buf \U$49064 ( \49039 , \49038 );
buf \U$49065 ( \49040 , \49039 );
nand \U$49066 ( \49041 , \48966 , \49040 );
buf \U$49067 ( \49042 , \49041 );
buf \U$49068 ( \49043 , \49042 );
xor \U$49069 ( \49044 , RIc0db188_127, RIc0d8488_31);
buf \U$49070 ( \49045 , \49044 );
not \U$49071 ( \49046 , \49045 );
buf \U$49072 ( \49047 , \15609 );
not \U$49073 ( \49048 , \49047 );
or \U$49074 ( \49049 , \49046 , \49048 );
buf \U$49075 ( \49050 , \47883 );
buf \U$49076 ( \49051 , RIc0db200_128);
nand \U$49077 ( \49052 , \49050 , \49051 );
buf \U$49078 ( \49053 , \49052 );
buf \U$49079 ( \49054 , \49053 );
nand \U$49080 ( \49055 , \49049 , \49054 );
buf \U$49081 ( \49056 , \49055 );
buf \U$49082 ( \49057 , \49056 );
not \U$49083 ( \49058 , \49057 );
buf \U$49084 ( \49059 , RIc0d8848_39);
buf \U$49085 ( \49060 , RIc0dadc8_119);
xor \U$49086 ( \49061 , \49059 , \49060 );
buf \U$49087 ( \49062 , \49061 );
buf \U$49088 ( \49063 , \49062 );
not \U$49089 ( \49064 , \49063 );
buf \U$49090 ( \49065 , \14569 );
not \U$49091 ( \49066 , \49065 );
or \U$49092 ( \49067 , \49064 , \49066 );
buf \U$49093 ( \49068 , \13953 );
buf \U$49094 ( \49069 , \47769 );
nand \U$49095 ( \49070 , \49068 , \49069 );
buf \U$49096 ( \49071 , \49070 );
buf \U$49097 ( \49072 , \49071 );
nand \U$49098 ( \49073 , \49067 , \49072 );
buf \U$49099 ( \49074 , \49073 );
buf \U$49100 ( \49075 , \49074 );
not \U$49101 ( \49076 , \49075 );
or \U$49102 ( \49077 , \49058 , \49076 );
buf \U$49103 ( \49078 , \49074 );
buf \U$49104 ( \49079 , \49056 );
or \U$49105 ( \49080 , \49078 , \49079 );
buf \U$49106 ( \49081 , RIc0d91a8_59);
buf \U$49107 ( \49082 , RIc0da468_99);
xor \U$49108 ( \49083 , \49081 , \49082 );
buf \U$49109 ( \49084 , \49083 );
buf \U$49110 ( \49085 , \49084 );
not \U$49111 ( \49086 , \49085 );
buf \U$49112 ( \49087 , \2470 );
not \U$49113 ( \49088 , \49087 );
or \U$49114 ( \49089 , \49086 , \49088 );
buf \U$49115 ( \49090 , \14648 );
buf \U$49116 ( \49091 , \48784 );
nand \U$49117 ( \49092 , \49090 , \49091 );
buf \U$49118 ( \49093 , \49092 );
buf \U$49119 ( \49094 , \49093 );
nand \U$49120 ( \49095 , \49089 , \49094 );
buf \U$49121 ( \49096 , \49095 );
buf \U$49122 ( \49097 , \49096 );
nand \U$49123 ( \49098 , \49080 , \49097 );
buf \U$49124 ( \49099 , \49098 );
buf \U$49125 ( \49100 , \49099 );
nand \U$49126 ( \49101 , \49077 , \49100 );
buf \U$49127 ( \49102 , \49101 );
buf \U$49128 ( \49103 , \49102 );
not \U$49129 ( \49104 , \49103 );
buf \U$49130 ( \49105 , \4008 );
buf \U$49131 ( \49106 , RIc0d9400_64);
and \U$49132 ( \49107 , \49105 , \49106 );
buf \U$49133 ( \49108 , \49107 );
buf \U$49134 ( \49109 , \49108 );
not \U$49135 ( \49110 , \49109 );
xor \U$49136 ( \49111 , RIc0da378_97, RIc0d9298_61);
buf \U$49137 ( \49112 , \49111 );
not \U$49138 ( \49113 , \49112 );
buf \U$49139 ( \49114 , \2941 );
not \U$49140 ( \49115 , \49114 );
or \U$49141 ( \49116 , \49113 , \49115 );
buf \U$49142 ( \49117 , \734 );
buf \U$49143 ( \49118 , \47831 );
nand \U$49144 ( \49119 , \49117 , \49118 );
buf \U$49145 ( \49120 , \49119 );
buf \U$49146 ( \49121 , \49120 );
nand \U$49147 ( \49122 , \49116 , \49121 );
buf \U$49148 ( \49123 , \49122 );
buf \U$49149 ( \49124 , \49123 );
not \U$49150 ( \49125 , \49124 );
or \U$49151 ( \49126 , \49110 , \49125 );
buf \U$49152 ( \49127 , \49123 );
buf \U$49153 ( \49128 , \49108 );
or \U$49154 ( \49129 , \49127 , \49128 );
buf \U$49155 ( \49130 , RIc0daeb8_121);
buf \U$49156 ( \49131 , RIc0d8758_37);
xnor \U$49157 ( \49132 , \49130 , \49131 );
buf \U$49158 ( \49133 , \49132 );
buf \U$49159 ( \49134 , \49133 );
not \U$49160 ( \49135 , \49134 );
buf \U$49161 ( \49136 , \49135 );
buf \U$49162 ( \49137 , \49136 );
not \U$49163 ( \49138 , \49137 );
buf \U$49164 ( \49139 , \16382 );
not \U$49165 ( \49140 , \49139 );
or \U$49166 ( \49141 , \49138 , \49140 );
buf \U$49167 ( \49142 , \16386 );
buf \U$49168 ( \49143 , \48765 );
nand \U$49169 ( \49144 , \49142 , \49143 );
buf \U$49170 ( \49145 , \49144 );
buf \U$49171 ( \49146 , \49145 );
nand \U$49172 ( \49147 , \49141 , \49146 );
buf \U$49173 ( \49148 , \49147 );
buf \U$49174 ( \49149 , \49148 );
nand \U$49175 ( \49150 , \49129 , \49149 );
buf \U$49176 ( \49151 , \49150 );
buf \U$49177 ( \49152 , \49151 );
nand \U$49178 ( \49153 , \49126 , \49152 );
buf \U$49179 ( \49154 , \49153 );
buf \U$49180 ( \49155 , \49154 );
not \U$49181 ( \49156 , \49155 );
or \U$49182 ( \49157 , \49104 , \49156 );
buf \U$49183 ( \49158 , \49154 );
buf \U$49184 ( \49159 , \49102 );
or \U$49185 ( \49160 , \49158 , \49159 );
xor \U$49186 ( \49161 , RIc0da918_109, RIc0d8cf8_49);
buf \U$49187 ( \49162 , \49161 );
not \U$49188 ( \49163 , \49162 );
buf \U$49189 ( \49164 , \14210 );
not \U$49190 ( \49165 , \49164 );
or \U$49191 ( \49166 , \49163 , \49165 );
buf \U$49192 ( \49167 , \47621 );
not \U$49193 ( \49168 , \49167 );
buf \U$49194 ( \49169 , \15909 );
nand \U$49195 ( \49170 , \49168 , \49169 );
buf \U$49196 ( \49171 , \49170 );
buf \U$49197 ( \49172 , \49171 );
nand \U$49198 ( \49173 , \49166 , \49172 );
buf \U$49199 ( \49174 , \49173 );
buf \U$49200 ( \49175 , \49174 );
buf \U$49201 ( \49176 , RIc0da738_105);
buf \U$49202 ( \49177 , RIc0d8ed8_53);
xnor \U$49203 ( \49178 , \49176 , \49177 );
buf \U$49204 ( \49179 , \49178 );
buf \U$49205 ( \49180 , \49179 );
not \U$49206 ( \49181 , \49180 );
buf \U$49207 ( \49182 , \49181 );
buf \U$49208 ( \49183 , \49182 );
not \U$49209 ( \49184 , \49183 );
buf \U$49210 ( \49185 , \12736 );
not \U$49211 ( \49186 , \49185 );
or \U$49212 ( \49187 , \49184 , \49186 );
buf \U$49213 ( \49188 , \12744 );
buf \U$49214 ( \49189 , \47708 );
nand \U$49215 ( \49190 , \49188 , \49189 );
buf \U$49216 ( \49191 , \49190 );
buf \U$49217 ( \49192 , \49191 );
nand \U$49218 ( \49193 , \49187 , \49192 );
buf \U$49219 ( \49194 , \49193 );
buf \U$49220 ( \49195 , \49194 );
xor \U$49221 ( \49196 , \49175 , \49195 );
buf \U$49222 ( \49197 , RIc0daa08_111);
buf \U$49223 ( \49198 , RIc0d8c08_47);
xor \U$49224 ( \49199 , \49197 , \49198 );
buf \U$49225 ( \49200 , \49199 );
buf \U$49226 ( \49201 , \49200 );
not \U$49227 ( \49202 , \49201 );
buf \U$49228 ( \49203 , \12529 );
not \U$49229 ( \49204 , \49203 );
or \U$49230 ( \49205 , \49202 , \49204 );
buf \U$49231 ( \49206 , \15864 );
buf \U$49232 ( \49207 , \47691 );
nand \U$49233 ( \49208 , \49206 , \49207 );
buf \U$49234 ( \49209 , \49208 );
buf \U$49235 ( \49210 , \49209 );
nand \U$49236 ( \49211 , \49205 , \49210 );
buf \U$49237 ( \49212 , \49211 );
buf \U$49238 ( \49213 , \49212 );
and \U$49239 ( \49214 , \49196 , \49213 );
and \U$49240 ( \49215 , \49175 , \49195 );
or \U$49241 ( \49216 , \49214 , \49215 );
buf \U$49242 ( \49217 , \49216 );
buf \U$49243 ( \49218 , \49217 );
nand \U$49244 ( \49219 , \49160 , \49218 );
buf \U$49245 ( \49220 , \49219 );
buf \U$49246 ( \49221 , \49220 );
nand \U$49247 ( \49222 , \49157 , \49221 );
buf \U$49248 ( \49223 , \49222 );
buf \U$49249 ( \49224 , \49223 );
xor \U$49250 ( \49225 , \49043 , \49224 );
xor \U$49251 ( \49226 , \47747 , \47811 );
xor \U$49252 ( \49227 , \49226 , \47867 );
buf \U$49253 ( \49228 , \49227 );
buf \U$49254 ( \49229 , \49228 );
and \U$49255 ( \49230 , \49225 , \49229 );
and \U$49256 ( \49231 , \49043 , \49224 );
or \U$49257 ( \49232 , \49230 , \49231 );
buf \U$49258 ( \49233 , \49232 );
buf \U$49259 ( \49234 , \49233 );
and \U$49260 ( \49235 , \48840 , \49234 );
and \U$49261 ( \49236 , \48835 , \48839 );
or \U$49262 ( \49237 , \49235 , \49236 );
buf \U$49263 ( \49238 , \49237 );
buf \U$49264 ( \49239 , \49238 );
xor \U$49265 ( \49240 , \47877 , \47974 );
xor \U$49266 ( \49241 , \49240 , \47979 );
buf \U$49267 ( \49242 , \49241 );
buf \U$49268 ( \49243 , \49242 );
xor \U$49269 ( \49244 , \49239 , \49243 );
xor \U$49270 ( \49245 , \47933 , \47937 );
xor \U$49271 ( \49246 , \49245 , \47942 );
buf \U$49272 ( \49247 , \49246 );
buf \U$49273 ( \49248 , \49247 );
xor \U$49274 ( \49249 , \47951 , \47955 );
xor \U$49275 ( \49250 , \49249 , \47959 );
buf \U$49276 ( \49251 , \49250 );
buf \U$49277 ( \49252 , \49251 );
or \U$49278 ( \49253 , \49248 , \49252 );
xor \U$49279 ( \49254 , \47827 , \47844 );
xor \U$49280 ( \49255 , \49254 , \47862 );
buf \U$49281 ( \49256 , \49255 );
buf \U$49282 ( \49257 , \49256 );
not \U$49283 ( \49258 , \49257 );
buf \U$49284 ( \49259 , \49258 );
buf \U$49285 ( \49260 , \49259 );
not \U$49286 ( \49261 , \49260 );
buf \U$49287 ( \49262 , \47803 );
not \U$49288 ( \49263 , \49262 );
buf \U$49289 ( \49264 , \47781 );
not \U$49290 ( \49265 , \49264 );
or \U$49291 ( \49266 , \49263 , \49265 );
buf \U$49292 ( \49267 , \47781 );
buf \U$49293 ( \49268 , \47803 );
or \U$49294 ( \49269 , \49267 , \49268 );
nand \U$49295 ( \49270 , \49266 , \49269 );
buf \U$49296 ( \49271 , \49270 );
buf \U$49297 ( \49272 , \49271 );
buf \U$49298 ( \49273 , \47763 );
not \U$49299 ( \49274 , \49273 );
buf \U$49300 ( \49275 , \49274 );
buf \U$49301 ( \49276 , \49275 );
and \U$49302 ( \49277 , \49272 , \49276 );
not \U$49303 ( \49278 , \49272 );
buf \U$49304 ( \49279 , \47763 );
and \U$49305 ( \49280 , \49278 , \49279 );
nor \U$49306 ( \49281 , \49277 , \49280 );
buf \U$49307 ( \49282 , \49281 );
buf \U$49308 ( \49283 , \49282 );
not \U$49309 ( \49284 , \49283 );
or \U$49310 ( \49285 , \49261 , \49284 );
xor \U$49311 ( \49286 , \47651 , \47631 );
xor \U$49312 ( \49287 , \49286 , \47669 );
buf \U$49313 ( \49288 , \49287 );
not \U$49314 ( \49289 , \49288 );
buf \U$49315 ( \49290 , \49289 );
buf \U$49316 ( \49291 , \49290 );
nand \U$49317 ( \49292 , \49285 , \49291 );
buf \U$49318 ( \49293 , \49292 );
buf \U$49319 ( \49294 , \49293 );
buf \U$49320 ( \49295 , \49282 );
not \U$49321 ( \49296 , \49295 );
buf \U$49322 ( \49297 , \49296 );
buf \U$49323 ( \49298 , \49297 );
buf \U$49324 ( \49299 , \49256 );
nand \U$49325 ( \49300 , \49298 , \49299 );
buf \U$49326 ( \49301 , \49300 );
buf \U$49327 ( \49302 , \49301 );
nand \U$49328 ( \49303 , \49294 , \49302 );
buf \U$49329 ( \49304 , \49303 );
buf \U$49330 ( \49305 , \49304 );
nand \U$49331 ( \49306 , \49253 , \49305 );
buf \U$49332 ( \49307 , \49306 );
buf \U$49333 ( \49308 , \49307 );
buf \U$49334 ( \49309 , \49247 );
buf \U$49335 ( \49310 , \49251 );
nand \U$49336 ( \49311 , \49309 , \49310 );
buf \U$49337 ( \49312 , \49311 );
buf \U$49338 ( \49313 , \49312 );
nand \U$49339 ( \49314 , \49308 , \49313 );
buf \U$49340 ( \49315 , \49314 );
buf \U$49341 ( \49316 , \49315 );
xor \U$49342 ( \49317 , \47947 , \47964 );
xor \U$49343 ( \49318 , \49317 , \47969 );
buf \U$49344 ( \49319 , \49318 );
buf \U$49345 ( \49320 , \49319 );
xor \U$49346 ( \49321 , \49316 , \49320 );
xor \U$49347 ( \49322 , \47527 , \47530 );
xor \U$49348 ( \49323 , \49322 , \47535 );
buf \U$49349 ( \49324 , \49323 );
buf \U$49350 ( \49325 , \49324 );
and \U$49351 ( \49326 , \49321 , \49325 );
and \U$49352 ( \49327 , \49316 , \49320 );
or \U$49353 ( \49328 , \49326 , \49327 );
buf \U$49354 ( \49329 , \49328 );
buf \U$49355 ( \49330 , \49329 );
and \U$49356 ( \49331 , \49244 , \49330 );
and \U$49357 ( \49332 , \49239 , \49243 );
or \U$49358 ( \49333 , \49331 , \49332 );
buf \U$49359 ( \49334 , \49333 );
buf \U$49360 ( \49335 , \49334 );
not \U$49361 ( \49336 , \49335 );
buf \U$49362 ( \49337 , \49336 );
buf \U$49363 ( \49338 , \49337 );
xor \U$49364 ( \49339 , \48758 , \49338 );
buf \U$49365 ( \49340 , \47521 );
not \U$49366 ( \49341 , \49340 );
buf \U$49367 ( \49342 , \47983 );
not \U$49368 ( \49343 , \49342 );
buf \U$49369 ( \49344 , \49343 );
buf \U$49370 ( \49345 , \49344 );
not \U$49371 ( \49346 , \49345 );
and \U$49372 ( \49347 , \49341 , \49346 );
buf \U$49373 ( \49348 , \47521 );
buf \U$49374 ( \49349 , \49344 );
and \U$49375 ( \49350 , \49348 , \49349 );
nor \U$49376 ( \49351 , \49347 , \49350 );
buf \U$49377 ( \49352 , \49351 );
buf \U$49378 ( \49353 , \49352 );
buf \U$49379 ( \49354 , \47553 );
and \U$49380 ( \49355 , \49353 , \49354 );
not \U$49381 ( \49356 , \49353 );
buf \U$49382 ( \49357 , \47553 );
not \U$49383 ( \49358 , \49357 );
buf \U$49384 ( \49359 , \49358 );
buf \U$49385 ( \49360 , \49359 );
and \U$49386 ( \49361 , \49356 , \49360 );
nor \U$49387 ( \49362 , \49355 , \49361 );
buf \U$49388 ( \49363 , \49362 );
buf \U$49389 ( \49364 , \49363 );
and \U$49390 ( \49365 , \49339 , \49364 );
and \U$49391 ( \49366 , \48758 , \49338 );
or \U$49392 ( \49367 , \49365 , \49366 );
buf \U$49393 ( \49368 , \49367 );
buf \U$49394 ( \49369 , \49368 );
nand \U$49395 ( \49370 , \48735 , \49369 );
buf \U$49396 ( \49371 , \49370 );
buf \U$49397 ( \49372 , \49371 );
and \U$49398 ( \49373 , \47443 , \48014 , \48728 , \49372 );
buf \U$49399 ( \49374 , \49373 );
buf \U$49400 ( \49375 , \49374 );
not \U$49401 ( \49376 , \49375 );
buf \U$49402 ( \49377 , \49056 );
buf \U$49403 ( \49378 , \49074 );
xor \U$49404 ( \49379 , \49377 , \49378 );
buf \U$49405 ( \49380 , \49096 );
xnor \U$49406 ( \49381 , \49379 , \49380 );
buf \U$49407 ( \49382 , \49381 );
buf \U$49408 ( \49383 , \49382 );
not \U$49409 ( \49384 , \49383 );
buf \U$49410 ( \49385 , \49108 );
buf \U$49411 ( \49386 , \49148 );
xor \U$49412 ( \49387 , \49385 , \49386 );
buf \U$49413 ( \49388 , \49123 );
xnor \U$49414 ( \49389 , \49387 , \49388 );
buf \U$49415 ( \49390 , \49389 );
buf \U$49416 ( \49391 , \49390 );
not \U$49417 ( \49392 , \49391 );
or \U$49418 ( \49393 , \49384 , \49392 );
xor \U$49419 ( \49394 , \48859 , \48881 );
not \U$49420 ( \49395 , \48900 );
xor \U$49421 ( \49396 , \49394 , \49395 );
buf \U$49422 ( \49397 , \49396 );
nand \U$49423 ( \49398 , \49393 , \49397 );
buf \U$49424 ( \49399 , \49398 );
buf \U$49425 ( \49400 , \49399 );
buf \U$49426 ( \49401 , \49390 );
not \U$49427 ( \49402 , \49401 );
buf \U$49428 ( \49403 , \49402 );
buf \U$49429 ( \49404 , \49403 );
buf \U$49430 ( \49405 , \49382 );
not \U$49431 ( \49406 , \49405 );
buf \U$49432 ( \49407 , \49406 );
buf \U$49433 ( \49408 , \49407 );
nand \U$49434 ( \49409 , \49404 , \49408 );
buf \U$49435 ( \49410 , \49409 );
buf \U$49436 ( \49411 , \49410 );
nand \U$49437 ( \49412 , \49400 , \49411 );
buf \U$49438 ( \49413 , \49412 );
buf \U$49439 ( \49414 , \49413 );
xor \U$49440 ( \49415 , \48963 , \49036 );
xor \U$49441 ( \49416 , \49415 , \48912 );
buf \U$49442 ( \49417 , \49416 );
xor \U$49443 ( \49418 , \49414 , \49417 );
buf \U$49444 ( \49419 , \49154 );
buf \U$49445 ( \49420 , \49102 );
xor \U$49446 ( \49421 , \49419 , \49420 );
buf \U$49447 ( \49422 , \49421 );
buf \U$49448 ( \49423 , \49422 );
buf \U$49449 ( \49424 , \49217 );
xor \U$49450 ( \49425 , \49423 , \49424 );
buf \U$49451 ( \49426 , \49425 );
buf \U$49452 ( \49427 , \49426 );
and \U$49453 ( \49428 , \49418 , \49427 );
and \U$49454 ( \49429 , \49414 , \49417 );
or \U$49455 ( \49430 , \49428 , \49429 );
buf \U$49456 ( \49431 , \49430 );
buf \U$49457 ( \49432 , \49431 );
buf \U$49458 ( \49433 , \48867 );
not \U$49459 ( \49434 , \49433 );
buf \U$49460 ( \49435 , \12937 );
not \U$49461 ( \49436 , \49435 );
or \U$49462 ( \49437 , \49434 , \49436 );
buf \U$49463 ( \49438 , \16556 );
buf \U$49464 ( \49439 , RIc0d89b0_42);
buf \U$49465 ( \49440 , RIc0dacd8_117);
xor \U$49466 ( \49441 , \49439 , \49440 );
buf \U$49467 ( \49442 , \49441 );
buf \U$49468 ( \49443 , \49442 );
buf \U$49469 ( \49444 , \12917 );
nand \U$49470 ( \49445 , \49438 , \49443 , \49444 );
buf \U$49471 ( \49446 , \49445 );
buf \U$49472 ( \49447 , \49446 );
nand \U$49473 ( \49448 , \49437 , \49447 );
buf \U$49474 ( \49449 , \49448 );
buf \U$49475 ( \49450 , \49449 );
not \U$49476 ( \49451 , \49450 );
buf \U$49477 ( \49452 , \49084 );
not \U$49478 ( \49453 , \49452 );
buf \U$49479 ( \49454 , \16750 );
not \U$49480 ( \49455 , \49454 );
or \U$49481 ( \49456 , \49453 , \49455 );
buf \U$49482 ( \49457 , \2199 );
buf \U$49483 ( \49458 , RIc0d9220_60);
buf \U$49484 ( \49459 , RIc0da468_99);
xor \U$49485 ( \49460 , \49458 , \49459 );
buf \U$49486 ( \49461 , \49460 );
buf \U$49487 ( \49462 , \49461 );
buf \U$49488 ( \49463 , \2203 );
nand \U$49489 ( \49464 , \49457 , \49462 , \49463 );
buf \U$49490 ( \49465 , \49464 );
buf \U$49491 ( \49466 , \49465 );
nand \U$49492 ( \49467 , \49456 , \49466 );
buf \U$49493 ( \49468 , \49467 );
buf \U$49494 ( \49469 , \49468 );
not \U$49495 ( \49470 , \49469 );
buf \U$49496 ( \49471 , \49470 );
buf \U$49497 ( \49472 , \49471 );
nand \U$49498 ( \49473 , \49451 , \49472 );
buf \U$49499 ( \49474 , \49473 );
buf \U$49500 ( \49475 , \49474 );
not \U$49501 ( \49476 , \49475 );
buf \U$49502 ( \49477 , RIc0d88c0_40);
buf \U$49503 ( \49478 , RIc0dadc8_119);
xor \U$49504 ( \49479 , \49477 , \49478 );
buf \U$49505 ( \49480 , \49479 );
buf \U$49506 ( \49481 , \49480 );
not \U$49507 ( \49482 , \49481 );
buf \U$49508 ( \49483 , \13949 );
not \U$49509 ( \49484 , \49483 );
or \U$49510 ( \49485 , \49482 , \49484 );
buf \U$49511 ( \49486 , \13953 );
buf \U$49512 ( \49487 , \49062 );
nand \U$49513 ( \49488 , \49486 , \49487 );
buf \U$49514 ( \49489 , \49488 );
buf \U$49515 ( \49490 , \49489 );
nand \U$49516 ( \49491 , \49485 , \49490 );
buf \U$49517 ( \49492 , \49491 );
buf \U$49518 ( \49493 , \49492 );
not \U$49519 ( \49494 , \49493 );
or \U$49520 ( \49495 , \49476 , \49494 );
buf \U$49521 ( \49496 , \49449 );
buf \U$49522 ( \49497 , \49468 );
nand \U$49523 ( \49498 , \49496 , \49497 );
buf \U$49524 ( \49499 , \49498 );
buf \U$49525 ( \49500 , \49499 );
nand \U$49526 ( \49501 , \49495 , \49500 );
buf \U$49527 ( \49502 , \49501 );
buf \U$49528 ( \49503 , \49502 );
buf \U$49529 ( \49504 , \49161 );
not \U$49530 ( \49505 , \49504 );
buf \U$49531 ( \49506 , \14216 );
not \U$49532 ( \49507 , \49506 );
or \U$49533 ( \49508 , \49505 , \49507 );
buf \U$49534 ( \49509 , \13423 );
xor \U$49535 ( \49510 , RIc0da918_109, RIc0d8d70_50);
buf \U$49536 ( \49511 , \49510 );
buf \U$49537 ( \49512 , \13413 );
nand \U$49538 ( \49513 , \49509 , \49511 , \49512 );
buf \U$49539 ( \49514 , \49513 );
buf \U$49540 ( \49515 , \49514 );
nand \U$49541 ( \49516 , \49508 , \49515 );
buf \U$49542 ( \49517 , \49516 );
buf \U$49543 ( \49518 , \49517 );
not \U$49544 ( \49519 , \49044 );
not \U$49545 ( \49520 , RIc0db200_128);
or \U$49546 ( \49521 , \49519 , \49520 );
buf \U$49547 ( \49522 , RIc0d8500_32);
buf \U$49548 ( \49523 , RIc0db188_127);
xnor \U$49549 ( \49524 , \49522 , \49523 );
buf \U$49550 ( \49525 , \49524 );
or \U$49551 ( \49526 , \18008 , \49525 );
nand \U$49552 ( \49527 , \49521 , \49526 );
buf \U$49553 ( \49528 , \49527 );
xor \U$49554 ( \49529 , \49518 , \49528 );
buf \U$49555 ( \49530 , \12532 );
buf \U$49556 ( \49531 , RIc0daa08_111);
buf \U$49557 ( \49532 , RIc0d8c80_48);
xor \U$49558 ( \49533 , \49531 , \49532 );
buf \U$49559 ( \49534 , \49533 );
buf \U$49560 ( \49535 , \49534 );
not \U$49561 ( \49536 , \49535 );
buf \U$49562 ( \49537 , \49536 );
buf \U$49563 ( \49538 , \49537 );
or \U$49564 ( \49539 , \49530 , \49538 );
buf \U$49565 ( \49540 , \14353 );
not \U$49566 ( \49541 , \49540 );
buf \U$49567 ( \49542 , \49541 );
buf \U$49568 ( \49543 , \49542 );
buf \U$49569 ( \49544 , \49200 );
not \U$49570 ( \49545 , \49544 );
buf \U$49571 ( \49546 , \49545 );
buf \U$49572 ( \49547 , \49546 );
or \U$49573 ( \49548 , \49543 , \49547 );
nand \U$49574 ( \49549 , \49539 , \49548 );
buf \U$49575 ( \49550 , \49549 );
buf \U$49576 ( \49551 , \49550 );
and \U$49577 ( \49552 , \49529 , \49551 );
and \U$49578 ( \49553 , \49518 , \49528 );
or \U$49579 ( \49554 , \49552 , \49553 );
buf \U$49580 ( \49555 , \49554 );
buf \U$49581 ( \49556 , \49555 );
or \U$49582 ( \49557 , \49503 , \49556 );
buf \U$49583 ( \49558 , RIc0da828_107);
buf \U$49584 ( \49559 , RIc0d8e60_52);
xor \U$49585 ( \49560 , \49558 , \49559 );
buf \U$49586 ( \49561 , \49560 );
buf \U$49587 ( \49562 , \49561 );
not \U$49588 ( \49563 , \49562 );
buf \U$49589 ( \49564 , \28794 );
not \U$49590 ( \49565 , \49564 );
or \U$49591 ( \49566 , \49563 , \49565 );
buf \U$49592 ( \49567 , \16071 );
buf \U$49593 ( \49568 , \48918 );
nand \U$49594 ( \49569 , \49567 , \49568 );
buf \U$49595 ( \49570 , \49569 );
buf \U$49596 ( \49571 , \49570 );
nand \U$49597 ( \49572 , \49566 , \49571 );
buf \U$49598 ( \49573 , \49572 );
buf \U$49599 ( \49574 , \49573 );
not \U$49600 ( \49575 , \49574 );
buf \U$49601 ( \49576 , \40787 );
buf \U$49602 ( \49577 , RIc0da738_105);
buf \U$49603 ( \49578 , RIc0d8f50_54);
xnor \U$49604 ( \49579 , \49577 , \49578 );
buf \U$49605 ( \49580 , \49579 );
buf \U$49606 ( \49581 , \49580 );
or \U$49607 ( \49582 , \49576 , \49581 );
buf \U$49608 ( \49583 , \15650 );
buf \U$49609 ( \49584 , \49179 );
or \U$49610 ( \49585 , \49583 , \49584 );
nand \U$49611 ( \49586 , \49582 , \49585 );
buf \U$49612 ( \49587 , \49586 );
buf \U$49613 ( \49588 , \49587 );
not \U$49614 ( \49589 , \49588 );
or \U$49615 ( \49590 , \49575 , \49589 );
buf \U$49616 ( \49591 , \49573 );
buf \U$49617 ( \49592 , \49587 );
or \U$49618 ( \49593 , \49591 , \49592 );
buf \U$49619 ( \49594 , RIc0da288_95);
buf \U$49620 ( \49595 , RIc0d9400_64);
and \U$49621 ( \49596 , \49594 , \49595 );
not \U$49622 ( \49597 , \49594 );
buf \U$49623 ( \49598 , \43843 );
and \U$49624 ( \49599 , \49597 , \49598 );
nor \U$49625 ( \49600 , \49596 , \49599 );
buf \U$49626 ( \49601 , \49600 );
buf \U$49627 ( \49602 , \49601 );
not \U$49628 ( \49603 , \49602 );
buf \U$49629 ( \49604 , \330 );
not \U$49630 ( \49605 , \49604 );
or \U$49631 ( \49606 , \49603 , \49605 );
buf \U$49632 ( \49607 , \344 );
buf \U$49633 ( \49608 , \48931 );
nand \U$49634 ( \49609 , \49607 , \49608 );
buf \U$49635 ( \49610 , \49609 );
buf \U$49636 ( \49611 , \49610 );
nand \U$49637 ( \49612 , \49606 , \49611 );
buf \U$49638 ( \49613 , \49612 );
buf \U$49639 ( \49614 , \49613 );
nand \U$49640 ( \49615 , \49593 , \49614 );
buf \U$49641 ( \49616 , \49615 );
buf \U$49642 ( \49617 , \49616 );
nand \U$49643 ( \49618 , \49590 , \49617 );
buf \U$49644 ( \49619 , \49618 );
buf \U$49645 ( \49620 , \49619 );
nand \U$49646 ( \49621 , \49557 , \49620 );
buf \U$49647 ( \49622 , \49621 );
buf \U$49648 ( \49623 , \49622 );
buf \U$49649 ( \49624 , \49502 );
buf \U$49650 ( \49625 , \49555 );
nand \U$49651 ( \49626 , \49624 , \49625 );
buf \U$49652 ( \49627 , \49626 );
buf \U$49653 ( \49628 , \49627 );
nand \U$49654 ( \49629 , \49623 , \49628 );
buf \U$49655 ( \49630 , \49629 );
buf \U$49656 ( \49631 , \49630 );
buf \U$49657 ( \49632 , RIc0d9310_62);
buf \U$49658 ( \49633 , RIc0da378_97);
xor \U$49659 ( \49634 , \49632 , \49633 );
buf \U$49660 ( \49635 , \49634 );
buf \U$49661 ( \49636 , \49635 );
not \U$49662 ( \49637 , \49636 );
buf \U$49663 ( \49638 , \29069 );
not \U$49664 ( \49639 , \49638 );
or \U$49665 ( \49640 , \49637 , \49639 );
buf \U$49666 ( \49641 , \2070 );
buf \U$49667 ( \49642 , \49111 );
nand \U$49668 ( \49643 , \49641 , \49642 );
buf \U$49669 ( \49644 , \49643 );
buf \U$49670 ( \49645 , \49644 );
nand \U$49671 ( \49646 , \49640 , \49645 );
buf \U$49672 ( \49647 , \49646 );
buf \U$49673 ( \49648 , \49647 );
not \U$49674 ( \49649 , \49648 );
buf \U$49675 ( \49650 , RIc0d9400_64);
buf \U$49676 ( \49651 , RIc0da300_96);
or \U$49677 ( \49652 , \49650 , \49651 );
buf \U$49678 ( \49653 , RIc0da378_97);
nand \U$49679 ( \49654 , \49652 , \49653 );
buf \U$49680 ( \49655 , \49654 );
buf \U$49681 ( \49656 , \49655 );
buf \U$49682 ( \49657 , RIc0d9400_64);
buf \U$49683 ( \49658 , RIc0da300_96);
nand \U$49684 ( \49659 , \49657 , \49658 );
buf \U$49685 ( \49660 , \49659 );
buf \U$49686 ( \49661 , \49660 );
buf \U$49687 ( \49662 , RIc0da288_95);
nand \U$49688 ( \49663 , \49656 , \49661 , \49662 );
buf \U$49689 ( \49664 , \49663 );
buf \U$49690 ( \49665 , \49664 );
nor \U$49691 ( \49666 , \49649 , \49665 );
buf \U$49692 ( \49667 , \49666 );
buf \U$49693 ( \49668 , \49667 );
not \U$49694 ( \49669 , \49668 );
buf \U$49695 ( \49670 , \19487 );
not \U$49696 ( \49671 , \49670 );
buf \U$49697 ( \49672 , \49671 );
buf \U$49698 ( \49673 , \49672 );
not \U$49699 ( \49674 , \49673 );
buf \U$49700 ( \49675 , RIc0daeb8_121);
buf \U$49701 ( \49676 , RIc0d87d0_38);
xnor \U$49702 ( \49677 , \49675 , \49676 );
buf \U$49703 ( \49678 , \49677 );
buf \U$49704 ( \49679 , \49678 );
not \U$49705 ( \49680 , \49679 );
and \U$49706 ( \49681 , \49674 , \49680 );
buf \U$49707 ( \49682 , \26373 );
buf \U$49708 ( \49683 , \49133 );
nor \U$49709 ( \49684 , \49682 , \49683 );
buf \U$49710 ( \49685 , \49684 );
buf \U$49711 ( \49686 , \49685 );
nor \U$49712 ( \49687 , \49681 , \49686 );
buf \U$49713 ( \49688 , \49687 );
buf \U$49714 ( \49689 , \49688 );
not \U$49715 ( \49690 , \49689 );
buf \U$49716 ( \49691 , \14888 );
not \U$49717 ( \49692 , \49691 );
buf \U$49718 ( \49693 , RIc0daaf8_113);
buf \U$49719 ( \49694 , RIc0d8b90_46);
xnor \U$49720 ( \49695 , \49693 , \49694 );
buf \U$49721 ( \49696 , \49695 );
buf \U$49722 ( \49697 , \49696 );
not \U$49723 ( \49698 , \49697 );
and \U$49724 ( \49699 , \49692 , \49698 );
buf \U$49725 ( \49700 , \34244 );
buf \U$49726 ( \49701 , \48844 );
nor \U$49727 ( \49702 , \49700 , \49701 );
buf \U$49728 ( \49703 , \49702 );
buf \U$49729 ( \49704 , \49703 );
nor \U$49730 ( \49705 , \49699 , \49704 );
buf \U$49731 ( \49706 , \49705 );
buf \U$49732 ( \49707 , \49706 );
not \U$49733 ( \49708 , \49707 );
or \U$49734 ( \49709 , \49690 , \49708 );
buf \U$49735 ( \49710 , RIc0da648_103);
buf \U$49736 ( \49711 , RIc0d9040_56);
xnor \U$49737 ( \49712 , \49710 , \49711 );
buf \U$49738 ( \49713 , \49712 );
buf \U$49739 ( \49714 , \49713 );
not \U$49740 ( \49715 , \49714 );
buf \U$49741 ( \49716 , \49715 );
buf \U$49742 ( \49717 , \49716 );
not \U$49743 ( \49718 , \49717 );
buf \U$49744 ( \49719 , \13042 );
not \U$49745 ( \49720 , \49719 );
or \U$49746 ( \49721 , \49718 , \49720 );
buf \U$49747 ( \49722 , \20243 );
buf \U$49748 ( \49723 , \48888 );
nand \U$49749 ( \49724 , \49722 , \49723 );
buf \U$49750 ( \49725 , \49724 );
buf \U$49751 ( \49726 , \49725 );
nand \U$49752 ( \49727 , \49721 , \49726 );
buf \U$49753 ( \49728 , \49727 );
buf \U$49754 ( \49729 , \49728 );
nand \U$49755 ( \49730 , \49709 , \49729 );
buf \U$49756 ( \49731 , \49730 );
buf \U$49757 ( \49732 , \49731 );
buf \U$49758 ( \49733 , \49688 );
not \U$49759 ( \49734 , \49733 );
buf \U$49760 ( \49735 , \49734 );
buf \U$49761 ( \49736 , \49735 );
buf \U$49762 ( \49737 , \49706 );
not \U$49763 ( \49738 , \49737 );
buf \U$49764 ( \49739 , \49738 );
buf \U$49765 ( \49740 , \49739 );
nand \U$49766 ( \49741 , \49736 , \49740 );
buf \U$49767 ( \49742 , \49741 );
buf \U$49768 ( \49743 , \49742 );
nand \U$49769 ( \49744 , \49732 , \49743 );
buf \U$49770 ( \49745 , \49744 );
buf \U$49771 ( \49746 , \49745 );
not \U$49772 ( \49747 , \49746 );
or \U$49773 ( \49748 , \49669 , \49747 );
buf \U$49774 ( \49749 , \49745 );
buf \U$49775 ( \49750 , \49667 );
or \U$49776 ( \49751 , \49749 , \49750 );
buf \U$49777 ( \49752 , RIc0db098_125);
buf \U$49778 ( \49753 , RIc0d85f0_34);
xor \U$49779 ( \49754 , \49752 , \49753 );
buf \U$49780 ( \49755 , \49754 );
buf \U$49781 ( \49756 , \49755 );
not \U$49782 ( \49757 , \49756 );
buf \U$49783 ( \49758 , \13460 );
not \U$49784 ( \49759 , \49758 );
or \U$49785 ( \49760 , \49757 , \49759 );
buf \U$49786 ( \49761 , \13465 );
buf \U$49787 ( \49762 , \48977 );
nand \U$49788 ( \49763 , \49761 , \49762 );
buf \U$49789 ( \49764 , \49763 );
buf \U$49790 ( \49765 , \49764 );
nand \U$49791 ( \49766 , \49760 , \49765 );
buf \U$49792 ( \49767 , \49766 );
buf \U$49793 ( \49768 , \49767 );
not \U$49794 ( \49769 , \49768 );
buf \U$49795 ( \49770 , RIc0d86e0_36);
buf \U$49796 ( \49771 , RIc0dafa8_123);
xnor \U$49797 ( \49772 , \49770 , \49771 );
buf \U$49798 ( \49773 , \49772 );
buf \U$49799 ( \49774 , \49773 );
not \U$49800 ( \49775 , \49774 );
buf \U$49801 ( \49776 , \49775 );
buf \U$49802 ( \49777 , \49776 );
not \U$49803 ( \49778 , \49777 );
buf \U$49804 ( \49779 , \47037 );
not \U$49805 ( \49780 , \49779 );
or \U$49806 ( \49781 , \49778 , \49780 );
buf \U$49807 ( \49782 , \16692 );
buf \U$49808 ( \49783 , \49018 );
nand \U$49809 ( \49784 , \49782 , \49783 );
buf \U$49810 ( \49785 , \49784 );
buf \U$49811 ( \49786 , \49785 );
nand \U$49812 ( \49787 , \49781 , \49786 );
buf \U$49813 ( \49788 , \49787 );
buf \U$49814 ( \49789 , \49788 );
not \U$49815 ( \49790 , \49789 );
or \U$49816 ( \49791 , \49769 , \49790 );
buf \U$49817 ( \49792 , \49788 );
buf \U$49818 ( \49793 , \49767 );
or \U$49819 ( \49794 , \49792 , \49793 );
buf \U$49820 ( \49795 , RIc0da558_101);
buf \U$49821 ( \49796 , RIc0d9130_58);
xnor \U$49822 ( \49797 , \49795 , \49796 );
buf \U$49823 ( \49798 , \49797 );
buf \U$49824 ( \49799 , \49798 );
not \U$49825 ( \49800 , \49799 );
buf \U$49826 ( \49801 , \49800 );
buf \U$49827 ( \49802 , \49801 );
not \U$49828 ( \49803 , \49802 );
buf \U$49829 ( \49804 , \4042 );
not \U$49830 ( \49805 , \49804 );
or \U$49831 ( \49806 , \49803 , \49805 );
buf \U$49832 ( \49807 , \26354 );
buf \U$49833 ( \49808 , \48948 );
nand \U$49834 ( \49809 , \49807 , \49808 );
buf \U$49835 ( \49810 , \49809 );
buf \U$49836 ( \49811 , \49810 );
nand \U$49837 ( \49812 , \49806 , \49811 );
buf \U$49838 ( \49813 , \49812 );
buf \U$49839 ( \49814 , \49813 );
nand \U$49840 ( \49815 , \49794 , \49814 );
buf \U$49841 ( \49816 , \49815 );
buf \U$49842 ( \49817 , \49816 );
nand \U$49843 ( \49818 , \49791 , \49817 );
buf \U$49844 ( \49819 , \49818 );
buf \U$49845 ( \49820 , \49819 );
nand \U$49846 ( \49821 , \49751 , \49820 );
buf \U$49847 ( \49822 , \49821 );
buf \U$49848 ( \49823 , \49822 );
nand \U$49849 ( \49824 , \49748 , \49823 );
buf \U$49850 ( \49825 , \49824 );
buf \U$49851 ( \49826 , \49825 );
xor \U$49852 ( \49827 , \49631 , \49826 );
xor \U$49853 ( \49828 , \48930 , \48943 );
xor \U$49854 ( \49829 , \49828 , \48960 );
buf \U$49855 ( \49830 , \49829 );
xor \U$49856 ( \49831 , \49175 , \49195 );
xor \U$49857 ( \49832 , \49831 , \49213 );
buf \U$49858 ( \49833 , \49832 );
buf \U$49859 ( \49834 , \49833 );
or \U$49860 ( \49835 , \49830 , \49834 );
xor \U$49861 ( \49836 , \49030 , \48990 );
xor \U$49862 ( \49837 , \49836 , \49008 );
buf \U$49863 ( \49838 , \49837 );
nand \U$49864 ( \49839 , \49835 , \49838 );
buf \U$49865 ( \49840 , \49839 );
buf \U$49866 ( \49841 , \49840 );
buf \U$49867 ( \49842 , \49829 );
buf \U$49868 ( \49843 , \49833 );
nand \U$49869 ( \49844 , \49842 , \49843 );
buf \U$49870 ( \49845 , \49844 );
buf \U$49871 ( \49846 , \49845 );
nand \U$49872 ( \49847 , \49841 , \49846 );
buf \U$49873 ( \49848 , \49847 );
buf \U$49874 ( \49849 , \49848 );
and \U$49875 ( \49850 , \49827 , \49849 );
and \U$49876 ( \49851 , \49631 , \49826 );
or \U$49877 ( \49852 , \49850 , \49851 );
buf \U$49878 ( \49853 , \49852 );
buf \U$49879 ( \49854 , \49853 );
xor \U$49880 ( \49855 , \49432 , \49854 );
buf \U$49881 ( \49856 , \49304 );
not \U$49882 ( \49857 , \49856 );
buf \U$49883 ( \49858 , \49857 );
buf \U$49884 ( \49859 , \49858 );
not \U$49885 ( \49860 , \49859 );
buf \U$49886 ( \49861 , \49247 );
not \U$49887 ( \49862 , \49861 );
or \U$49888 ( \49863 , \49860 , \49862 );
buf \U$49889 ( \49864 , \49858 );
buf \U$49890 ( \49865 , \49247 );
or \U$49891 ( \49866 , \49864 , \49865 );
nand \U$49892 ( \49867 , \49863 , \49866 );
buf \U$49893 ( \49868 , \49867 );
buf \U$49894 ( \49869 , \49868 );
buf \U$49895 ( \49870 , \49251 );
and \U$49896 ( \49871 , \49869 , \49870 );
not \U$49897 ( \49872 , \49869 );
buf \U$49898 ( \49873 , \49251 );
not \U$49899 ( \49874 , \49873 );
buf \U$49900 ( \49875 , \49874 );
buf \U$49901 ( \49876 , \49875 );
and \U$49902 ( \49877 , \49872 , \49876 );
nor \U$49903 ( \49878 , \49871 , \49877 );
buf \U$49904 ( \49879 , \49878 );
buf \U$49905 ( \49880 , \49879 );
and \U$49906 ( \49881 , \49855 , \49880 );
and \U$49907 ( \49882 , \49432 , \49854 );
or \U$49908 ( \49883 , \49881 , \49882 );
buf \U$49909 ( \49884 , \49883 );
buf \U$49910 ( \49885 , \49884 );
not \U$49911 ( \49886 , \49885 );
buf \U$49912 ( \49887 , \49886 );
buf \U$49913 ( \49888 , \49259 );
not \U$49914 ( \49889 , \49888 );
buf \U$49915 ( \49890 , \49290 );
not \U$49916 ( \49891 , \49890 );
or \U$49917 ( \49892 , \49889 , \49891 );
buf \U$49918 ( \49893 , \49287 );
buf \U$49919 ( \49894 , \49256 );
nand \U$49920 ( \49895 , \49893 , \49894 );
buf \U$49921 ( \49896 , \49895 );
buf \U$49922 ( \49897 , \49896 );
nand \U$49923 ( \49898 , \49892 , \49897 );
buf \U$49924 ( \49899 , \49898 );
buf \U$49925 ( \49900 , \49899 );
buf \U$49926 ( \49901 , \49297 );
and \U$49927 ( \49902 , \49900 , \49901 );
not \U$49928 ( \49903 , \49900 );
buf \U$49929 ( \49904 , \49282 );
and \U$49930 ( \49905 , \49903 , \49904 );
nor \U$49931 ( \49906 , \49902 , \49905 );
buf \U$49932 ( \49907 , \49906 );
buf \U$49933 ( \49908 , \49907 );
xor \U$49934 ( \49909 , \47897 , \47911 );
xor \U$49935 ( \49910 , \49909 , \47928 );
buf \U$49936 ( \49911 , \49910 );
buf \U$49937 ( \49912 , \49911 );
xor \U$49938 ( \49913 , \47735 , \47703 );
xor \U$49939 ( \49914 , \49913 , \47720 );
buf \U$49940 ( \49915 , \49914 );
xor \U$49941 ( \49916 , \49912 , \49915 );
xor \U$49942 ( \49917 , \48778 , \48815 );
xnor \U$49943 ( \49918 , \49917 , \48809 );
buf \U$49944 ( \49919 , \49918 );
xor \U$49945 ( \49920 , \49916 , \49919 );
buf \U$49946 ( \49921 , \49920 );
buf \U$49947 ( \49922 , \49921 );
xor \U$49948 ( \49923 , \49908 , \49922 );
xor \U$49949 ( \49924 , \49631 , \49826 );
xor \U$49950 ( \49925 , \49924 , \49849 );
buf \U$49951 ( \49926 , \49925 );
buf \U$49952 ( \49927 , \49926 );
and \U$49953 ( \49928 , \49923 , \49927 );
and \U$49954 ( \49929 , \49908 , \49922 );
or \U$49955 ( \49930 , \49928 , \49929 );
buf \U$49956 ( \49931 , \49930 );
buf \U$49957 ( \49932 , \49931 );
xor \U$49958 ( \49933 , \49912 , \49915 );
and \U$49959 ( \49934 , \49933 , \49919 );
and \U$49960 ( \49935 , \49912 , \49915 );
or \U$49961 ( \49936 , \49934 , \49935 );
buf \U$49962 ( \49937 , \49936 );
buf \U$49963 ( \49938 , \49937 );
xor \U$49964 ( \49939 , \48761 , \48825 );
xor \U$49965 ( \49940 , \49939 , \48830 );
buf \U$49966 ( \49941 , \49940 );
buf \U$49967 ( \49942 , \49941 );
xor \U$49968 ( \49943 , \49938 , \49942 );
xor \U$49969 ( \49944 , \49043 , \49224 );
xor \U$49970 ( \49945 , \49944 , \49229 );
buf \U$49971 ( \49946 , \49945 );
buf \U$49972 ( \49947 , \49946 );
xor \U$49973 ( \49948 , \49943 , \49947 );
buf \U$49974 ( \49949 , \49948 );
buf \U$49975 ( \49950 , \49949 );
xor \U$49976 ( \49951 , \49932 , \49950 );
buf \U$49977 ( \49952 , \14681 );
xor \U$49978 ( \49953 , RIc0dabe8_115, RIc0d8aa0_44);
buf \U$49979 ( \49954 , \49953 );
not \U$49980 ( \49955 , \49954 );
buf \U$49981 ( \49956 , \49955 );
buf \U$49982 ( \49957 , \49956 );
or \U$49983 ( \49958 , \49952 , \49957 );
buf \U$49984 ( \49959 , \29865 );
buf \U$49985 ( \49960 , \48996 );
not \U$49986 ( \49961 , \49960 );
buf \U$49987 ( \49962 , \49961 );
buf \U$49988 ( \49963 , \49962 );
or \U$49989 ( \49964 , \49959 , \49963 );
nand \U$49990 ( \49965 , \49958 , \49964 );
buf \U$49991 ( \49966 , \49965 );
buf \U$49992 ( \49967 , \49966 );
buf \U$49993 ( \49968 , \49664 );
not \U$49994 ( \49969 , \49968 );
buf \U$49995 ( \49970 , \49647 );
not \U$49996 ( \49971 , \49970 );
or \U$49997 ( \49972 , \49969 , \49971 );
buf \U$49998 ( \49973 , \49647 );
buf \U$49999 ( \49974 , \49664 );
or \U$50000 ( \49975 , \49973 , \49974 );
nand \U$50001 ( \49976 , \49972 , \49975 );
buf \U$50002 ( \49977 , \49976 );
buf \U$50003 ( \49978 , \49977 );
xor \U$50004 ( \49979 , \49967 , \49978 );
xor \U$50005 ( \49980 , RIc0dabe8_115, RIc0d8b18_45);
buf \U$50006 ( \49981 , \49980 );
not \U$50007 ( \49982 , \49981 );
buf \U$50008 ( \49983 , \14186 );
not \U$50009 ( \49984 , \49983 );
or \U$50010 ( \49985 , \49982 , \49984 );
buf \U$50011 ( \49986 , \12303 );
buf \U$50012 ( \49987 , \49953 );
nand \U$50013 ( \49988 , \49986 , \49987 );
buf \U$50014 ( \49989 , \49988 );
buf \U$50015 ( \49990 , \49989 );
nand \U$50016 ( \49991 , \49985 , \49990 );
buf \U$50017 ( \49992 , \49991 );
buf \U$50018 ( \49993 , \49992 );
buf \U$50019 ( \49994 , RIc0d8c08_47);
buf \U$50020 ( \49995 , RIc0daaf8_113);
xor \U$50021 ( \49996 , \49994 , \49995 );
buf \U$50022 ( \49997 , \49996 );
buf \U$50023 ( \49998 , \49997 );
not \U$50024 ( \49999 , \49998 );
buf \U$50025 ( \50000 , \28413 );
not \U$50026 ( \50001 , \50000 );
or \U$50027 ( \50002 , \49999 , \50001 );
buf \U$50028 ( \50003 , \49696 );
not \U$50029 ( \50004 , \50003 );
buf \U$50030 ( \50005 , \16662 );
nand \U$50031 ( \50006 , \50004 , \50005 );
buf \U$50032 ( \50007 , \50006 );
buf \U$50033 ( \50008 , \50007 );
nand \U$50034 ( \50009 , \50002 , \50008 );
buf \U$50035 ( \50010 , \50009 );
buf \U$50036 ( \50011 , \50010 );
nor \U$50037 ( \50012 , \49993 , \50011 );
buf \U$50038 ( \50013 , \50012 );
buf \U$50039 ( \50014 , \50013 );
buf \U$50040 ( \50015 , \4483 );
not \U$50041 ( \50016 , \50015 );
buf \U$50042 ( \50017 , RIc0da648_103);
buf \U$50043 ( \50018 , RIc0d90b8_57);
xnor \U$50044 ( \50019 , \50017 , \50018 );
buf \U$50045 ( \50020 , \50019 );
buf \U$50046 ( \50021 , \50020 );
not \U$50047 ( \50022 , \50021 );
and \U$50048 ( \50023 , \50016 , \50022 );
buf \U$50049 ( \50024 , \4475 );
buf \U$50050 ( \50025 , \49713 );
nor \U$50051 ( \50026 , \50024 , \50025 );
buf \U$50052 ( \50027 , \50026 );
buf \U$50053 ( \50028 , \50027 );
nor \U$50054 ( \50029 , \50023 , \50028 );
buf \U$50055 ( \50030 , \50029 );
buf \U$50056 ( \50031 , \50030 );
or \U$50057 ( \50032 , \50014 , \50031 );
buf \U$50058 ( \50033 , \50010 );
buf \U$50059 ( \50034 , \49992 );
nand \U$50060 ( \50035 , \50033 , \50034 );
buf \U$50061 ( \50036 , \50035 );
buf \U$50062 ( \50037 , \50036 );
nand \U$50063 ( \50038 , \50032 , \50037 );
buf \U$50064 ( \50039 , \50038 );
buf \U$50065 ( \50040 , \50039 );
and \U$50066 ( \50041 , \49979 , \50040 );
and \U$50067 ( \50042 , \49967 , \49978 );
or \U$50068 ( \50043 , \50041 , \50042 );
buf \U$50069 ( \50044 , \50043 );
buf \U$50070 ( \50045 , \50044 );
not \U$50071 ( \50046 , \50045 );
buf \U$50072 ( \50047 , \12651 );
buf \U$50073 ( \50048 , RIc0d8578_33);
buf \U$50074 ( \50049 , RIc0db188_127);
xor \U$50075 ( \50050 , \50048 , \50049 );
buf \U$50076 ( \50051 , \50050 );
buf \U$50077 ( \50052 , \50051 );
not \U$50078 ( \50053 , \50052 );
buf \U$50079 ( \50054 , \50053 );
buf \U$50080 ( \50055 , \50054 );
or \U$50081 ( \50056 , \50047 , \50055 );
buf \U$50082 ( \50057 , \12647 );
buf \U$50083 ( \50058 , \49525 );
or \U$50084 ( \50059 , \50057 , \50058 );
nand \U$50085 ( \50060 , \50056 , \50059 );
buf \U$50086 ( \50061 , \50060 );
buf \U$50087 ( \50062 , \50061 );
buf \U$50088 ( \50063 , \343 );
buf \U$50089 ( \50064 , RIc0d9400_64);
and \U$50090 ( \50065 , \50063 , \50064 );
buf \U$50091 ( \50066 , \50065 );
buf \U$50092 ( \50067 , \50066 );
xor \U$50093 ( \50068 , \50062 , \50067 );
xor \U$50094 ( \50069 , RIc0da468_99, RIc0d9298_61);
buf \U$50095 ( \50070 , \50069 );
not \U$50096 ( \50071 , \50070 );
buf \U$50097 ( \50072 , \16744 );
not \U$50098 ( \50073 , \50072 );
or \U$50099 ( \50074 , \50071 , \50073 );
buf \U$50100 ( \50075 , \12584 );
buf \U$50101 ( \50076 , \49461 );
nand \U$50102 ( \50077 , \50075 , \50076 );
buf \U$50103 ( \50078 , \50077 );
buf \U$50104 ( \50079 , \50078 );
nand \U$50105 ( \50080 , \50074 , \50079 );
buf \U$50106 ( \50081 , \50080 );
buf \U$50107 ( \50082 , \50081 );
and \U$50108 ( \50083 , \50068 , \50082 );
and \U$50109 ( \50084 , \50062 , \50067 );
or \U$50110 ( \50085 , \50083 , \50084 );
buf \U$50111 ( \50086 , \50085 );
buf \U$50112 ( \50087 , \50086 );
buf \U$50113 ( \50088 , RIc0db098_125);
buf \U$50114 ( \50089 , RIc0d8668_35);
xor \U$50115 ( \50090 , \50088 , \50089 );
buf \U$50116 ( \50091 , \50090 );
buf \U$50117 ( \50092 , \50091 );
not \U$50118 ( \50093 , \50092 );
buf \U$50119 ( \50094 , \14471 );
not \U$50120 ( \50095 , \50094 );
or \U$50121 ( \50096 , \50093 , \50095 );
buf \U$50122 ( \50097 , \15793 );
buf \U$50123 ( \50098 , \49755 );
nand \U$50124 ( \50099 , \50097 , \50098 );
buf \U$50125 ( \50100 , \50099 );
buf \U$50126 ( \50101 , \50100 );
nand \U$50127 ( \50102 , \50096 , \50101 );
buf \U$50128 ( \50103 , \50102 );
buf \U$50129 ( \50104 , \50103 );
xor \U$50130 ( \50105 , RIc0daa08_111, RIc0d8cf8_49);
buf \U$50131 ( \50106 , \50105 );
not \U$50132 ( \50107 , \50106 );
buf \U$50133 ( \50108 , \12529 );
not \U$50134 ( \50109 , \50108 );
or \U$50135 ( \50110 , \50107 , \50109 );
buf \U$50136 ( \50111 , \14106 );
buf \U$50137 ( \50112 , \49534 );
nand \U$50138 ( \50113 , \50111 , \50112 );
buf \U$50139 ( \50114 , \50113 );
buf \U$50140 ( \50115 , \50114 );
nand \U$50141 ( \50116 , \50110 , \50115 );
buf \U$50142 ( \50117 , \50116 );
buf \U$50143 ( \50118 , \50117 );
nor \U$50144 ( \50119 , \50104 , \50118 );
buf \U$50145 ( \50120 , \50119 );
buf \U$50146 ( \50121 , \50120 );
buf \U$50147 ( \50122 , \46183 );
not \U$50148 ( \50123 , \50122 );
buf \U$50149 ( \50124 , RIc0dafa8_123);
buf \U$50150 ( \50125 , RIc0d8758_37);
xor \U$50151 ( \50126 , \50124 , \50125 );
buf \U$50152 ( \50127 , \50126 );
buf \U$50153 ( \50128 , \50127 );
not \U$50154 ( \50129 , \50128 );
buf \U$50155 ( \50130 , \50129 );
buf \U$50156 ( \50131 , \50130 );
not \U$50157 ( \50132 , \50131 );
and \U$50158 ( \50133 , \50123 , \50132 );
buf \U$50159 ( \50134 , \16692 );
not \U$50160 ( \50135 , \50134 );
buf \U$50161 ( \50136 , \49773 );
nor \U$50162 ( \50137 , \50135 , \50136 );
buf \U$50163 ( \50138 , \50137 );
buf \U$50164 ( \50139 , \50138 );
nor \U$50165 ( \50140 , \50133 , \50139 );
buf \U$50166 ( \50141 , \50140 );
buf \U$50167 ( \50142 , \50141 );
or \U$50168 ( \50143 , \50121 , \50142 );
buf \U$50169 ( \50144 , \50117 );
buf \U$50170 ( \50145 , \50103 );
nand \U$50171 ( \50146 , \50144 , \50145 );
buf \U$50172 ( \50147 , \50146 );
buf \U$50173 ( \50148 , \50147 );
nand \U$50174 ( \50149 , \50143 , \50148 );
buf \U$50175 ( \50150 , \50149 );
buf \U$50176 ( \50151 , \50150 );
xor \U$50177 ( \50152 , \50087 , \50151 );
buf \U$50178 ( \50153 , \36626 );
buf \U$50179 ( \50154 , RIc0da558_101);
buf \U$50180 ( \50155 , RIc0d91a8_59);
xor \U$50181 ( \50156 , \50154 , \50155 );
buf \U$50182 ( \50157 , \50156 );
buf \U$50183 ( \50158 , \50157 );
not \U$50184 ( \50159 , \50158 );
buf \U$50185 ( \50160 , \50159 );
buf \U$50186 ( \50161 , \50160 );
or \U$50187 ( \50162 , \50153 , \50161 );
buf \U$50188 ( \50163 , \16676 );
not \U$50189 ( \50164 , \50163 );
buf \U$50190 ( \50165 , \50164 );
buf \U$50191 ( \50166 , \50165 );
buf \U$50192 ( \50167 , \49798 );
or \U$50193 ( \50168 , \50166 , \50167 );
nand \U$50194 ( \50169 , \50162 , \50168 );
buf \U$50195 ( \50170 , \50169 );
buf \U$50196 ( \50171 , \50170 );
xor \U$50197 ( \50172 , RIc0daeb8_121, RIc0d8848_39);
buf \U$50198 ( \50173 , \50172 );
not \U$50199 ( \50174 , \50173 );
buf \U$50200 ( \50175 , \19487 );
not \U$50201 ( \50176 , \50175 );
or \U$50202 ( \50177 , \50174 , \50176 );
buf \U$50203 ( \50178 , \49678 );
not \U$50204 ( \50179 , \50178 );
buf \U$50205 ( \50180 , \13314 );
nand \U$50206 ( \50181 , \50179 , \50180 );
buf \U$50207 ( \50182 , \50181 );
buf \U$50208 ( \50183 , \50182 );
nand \U$50209 ( \50184 , \50177 , \50183 );
buf \U$50210 ( \50185 , \50184 );
buf \U$50211 ( \50186 , \50185 );
xor \U$50212 ( \50187 , \50171 , \50186 );
buf \U$50213 ( \50188 , \13178 );
buf \U$50214 ( \50189 , RIc0dadc8_119);
buf \U$50215 ( \50190 , RIc0d8938_41);
xnor \U$50216 ( \50191 , \50189 , \50190 );
buf \U$50217 ( \50192 , \50191 );
buf \U$50218 ( \50193 , \50192 );
or \U$50219 ( \50194 , \50188 , \50193 );
buf \U$50220 ( \50195 , \45225 );
buf \U$50221 ( \50196 , \49480 );
not \U$50222 ( \50197 , \50196 );
buf \U$50223 ( \50198 , \50197 );
buf \U$50224 ( \50199 , \50198 );
or \U$50225 ( \50200 , \50195 , \50199 );
nand \U$50226 ( \50201 , \50194 , \50200 );
buf \U$50227 ( \50202 , \50201 );
buf \U$50228 ( \50203 , \50202 );
and \U$50229 ( \50204 , \50187 , \50203 );
and \U$50230 ( \50205 , \50171 , \50186 );
or \U$50231 ( \50206 , \50204 , \50205 );
buf \U$50232 ( \50207 , \50206 );
buf \U$50233 ( \50208 , \50207 );
and \U$50234 ( \50209 , \50152 , \50208 );
and \U$50235 ( \50210 , \50087 , \50151 );
or \U$50236 ( \50211 , \50209 , \50210 );
buf \U$50237 ( \50212 , \50211 );
buf \U$50238 ( \50213 , \50212 );
not \U$50239 ( \50214 , \50213 );
or \U$50240 ( \50215 , \50046 , \50214 );
buf \U$50241 ( \50216 , \50212 );
buf \U$50242 ( \50217 , \50044 );
or \U$50243 ( \50218 , \50216 , \50217 );
xor \U$50244 ( \50219 , \49619 , \49502 );
xor \U$50245 ( \50220 , \50219 , \49555 );
buf \U$50246 ( \50221 , \50220 );
nand \U$50247 ( \50222 , \50218 , \50221 );
buf \U$50248 ( \50223 , \50222 );
buf \U$50249 ( \50224 , \50223 );
nand \U$50250 ( \50225 , \50215 , \50224 );
buf \U$50251 ( \50226 , \50225 );
buf \U$50252 ( \50227 , \50226 );
xor \U$50253 ( \50228 , \49767 , \49813 );
xnor \U$50254 ( \50229 , \50228 , \49788 );
buf \U$50255 ( \50230 , \50229 );
not \U$50256 ( \50231 , \50230 );
buf \U$50257 ( \50232 , \50231 );
buf \U$50258 ( \50233 , \50232 );
not \U$50259 ( \50234 , \50233 );
buf \U$50260 ( \50235 , \49735 );
not \U$50261 ( \50236 , \50235 );
buf \U$50262 ( \50237 , \49706 );
not \U$50263 ( \50238 , \50237 );
or \U$50264 ( \50239 , \50236 , \50238 );
buf \U$50265 ( \50240 , \49739 );
buf \U$50266 ( \50241 , \49688 );
nand \U$50267 ( \50242 , \50240 , \50241 );
buf \U$50268 ( \50243 , \50242 );
buf \U$50269 ( \50244 , \50243 );
nand \U$50270 ( \50245 , \50239 , \50244 );
buf \U$50271 ( \50246 , \50245 );
buf \U$50272 ( \50247 , \50246 );
buf \U$50273 ( \50248 , \49728 );
xnor \U$50274 ( \50249 , \50247 , \50248 );
buf \U$50275 ( \50250 , \50249 );
buf \U$50276 ( \50251 , \50250 );
not \U$50277 ( \50252 , \50251 );
buf \U$50278 ( \50253 , \50252 );
buf \U$50279 ( \50254 , \50253 );
not \U$50280 ( \50255 , \50254 );
or \U$50281 ( \50256 , \50234 , \50255 );
buf \U$50282 ( \50257 , \50250 );
not \U$50283 ( \50258 , \50257 );
buf \U$50284 ( \50259 , \50229 );
not \U$50285 ( \50260 , \50259 );
or \U$50286 ( \50261 , \50258 , \50260 );
buf \U$50287 ( \50262 , RIc0da828_107);
buf \U$50288 ( \50263 , RIc0d8ed8_53);
xor \U$50289 ( \50264 , \50262 , \50263 );
buf \U$50290 ( \50265 , \50264 );
buf \U$50291 ( \50266 , \50265 );
not \U$50292 ( \50267 , \50266 );
buf \U$50293 ( \50268 , \17595 );
not \U$50294 ( \50269 , \50268 );
or \U$50295 ( \50270 , \50267 , \50269 );
buf \U$50296 ( \50271 , \12342 );
buf \U$50297 ( \50272 , \49561 );
nand \U$50298 ( \50273 , \50271 , \50272 );
buf \U$50299 ( \50274 , \50273 );
buf \U$50300 ( \50275 , \50274 );
nand \U$50301 ( \50276 , \50270 , \50275 );
buf \U$50302 ( \50277 , \50276 );
buf \U$50303 ( \50278 , \50277 );
xor \U$50304 ( \50279 , RIc0da918_109, RIc0d8de8_51);
buf \U$50305 ( \50280 , \50279 );
not \U$50306 ( \50281 , \50280 );
buf \U$50307 ( \50282 , \21959 );
not \U$50308 ( \50283 , \50282 );
or \U$50309 ( \50284 , \50281 , \50283 );
buf \U$50310 ( \50285 , \20211 );
buf \U$50311 ( \50286 , \49510 );
nand \U$50312 ( \50287 , \50285 , \50286 );
buf \U$50313 ( \50288 , \50287 );
buf \U$50314 ( \50289 , \50288 );
nand \U$50315 ( \50290 , \50284 , \50289 );
buf \U$50316 ( \50291 , \50290 );
buf \U$50317 ( \50292 , \50291 );
xor \U$50318 ( \50293 , \50278 , \50292 );
buf \U$50319 ( \50294 , RIc0da378_97);
buf \U$50320 ( \50295 , RIc0d9388_63);
and \U$50321 ( \50296 , \50294 , \50295 );
not \U$50322 ( \50297 , \50294 );
buf \U$50323 ( \50298 , \43939 );
and \U$50324 ( \50299 , \50297 , \50298 );
nor \U$50325 ( \50300 , \50296 , \50299 );
buf \U$50326 ( \50301 , \50300 );
buf \U$50327 ( \50302 , \50301 );
not \U$50328 ( \50303 , \50302 );
buf \U$50329 ( \50304 , \2066 );
not \U$50330 ( \50305 , \50304 );
or \U$50331 ( \50306 , \50303 , \50305 );
buf \U$50332 ( \50307 , \2070 );
buf \U$50333 ( \50308 , \49635 );
nand \U$50334 ( \50309 , \50307 , \50308 );
buf \U$50335 ( \50310 , \50309 );
buf \U$50336 ( \50311 , \50310 );
nand \U$50337 ( \50312 , \50306 , \50311 );
buf \U$50338 ( \50313 , \50312 );
buf \U$50339 ( \50314 , \50313 );
and \U$50340 ( \50315 , \50293 , \50314 );
and \U$50341 ( \50316 , \50278 , \50292 );
or \U$50342 ( \50317 , \50315 , \50316 );
buf \U$50343 ( \50318 , \50317 );
buf \U$50344 ( \50319 , \50318 );
nand \U$50345 ( \50320 , \50261 , \50319 );
buf \U$50346 ( \50321 , \50320 );
buf \U$50347 ( \50322 , \50321 );
nand \U$50348 ( \50323 , \50256 , \50322 );
buf \U$50349 ( \50324 , \50323 );
buf \U$50350 ( \50325 , \50324 );
xor \U$50351 ( \50326 , \49449 , \49471 );
xnor \U$50352 ( \50327 , \50326 , \49492 );
buf \U$50353 ( \50328 , \50327 );
xor \U$50354 ( \50329 , \49518 , \49528 );
xor \U$50355 ( \50330 , \50329 , \49551 );
buf \U$50356 ( \50331 , \50330 );
buf \U$50357 ( \50332 , \50331 );
xor \U$50358 ( \50333 , \50328 , \50332 );
xor \U$50359 ( \50334 , \49573 , \49613 );
xor \U$50360 ( \50335 , \50334 , \49587 );
buf \U$50361 ( \50336 , \50335 );
and \U$50362 ( \50337 , \50333 , \50336 );
and \U$50363 ( \50338 , \50328 , \50332 );
or \U$50364 ( \50339 , \50337 , \50338 );
buf \U$50365 ( \50340 , \50339 );
buf \U$50366 ( \50341 , \50340 );
nor \U$50367 ( \50342 , \50325 , \50341 );
buf \U$50368 ( \50343 , \50342 );
buf \U$50369 ( \50344 , \50343 );
buf \U$50370 ( \50345 , \49667 );
buf \U$50371 ( \50346 , \49745 );
xor \U$50372 ( \50347 , \50345 , \50346 );
buf \U$50373 ( \50348 , \49819 );
xnor \U$50374 ( \50349 , \50347 , \50348 );
buf \U$50375 ( \50350 , \50349 );
buf \U$50376 ( \50351 , \50350 );
or \U$50377 ( \50352 , \50344 , \50351 );
buf \U$50378 ( \50353 , \50324 );
buf \U$50379 ( \50354 , \50340 );
nand \U$50380 ( \50355 , \50353 , \50354 );
buf \U$50381 ( \50356 , \50355 );
buf \U$50382 ( \50357 , \50356 );
nand \U$50383 ( \50358 , \50352 , \50357 );
buf \U$50384 ( \50359 , \50358 );
buf \U$50385 ( \50360 , \50359 );
xor \U$50386 ( \50361 , \50227 , \50360 );
xor \U$50387 ( \50362 , \49414 , \49417 );
xor \U$50388 ( \50363 , \50362 , \49427 );
buf \U$50389 ( \50364 , \50363 );
buf \U$50390 ( \50365 , \50364 );
and \U$50391 ( \50366 , \50361 , \50365 );
and \U$50392 ( \50367 , \50227 , \50360 );
or \U$50393 ( \50368 , \50366 , \50367 );
buf \U$50394 ( \50369 , \50368 );
buf \U$50395 ( \50370 , \50369 );
and \U$50396 ( \50371 , \49951 , \50370 );
and \U$50397 ( \50372 , \49932 , \49950 );
or \U$50398 ( \50373 , \50371 , \50372 );
buf \U$50399 ( \50374 , \50373 );
xor \U$50400 ( \50375 , \49887 , \50374 );
xor \U$50401 ( \50376 , \49938 , \49942 );
and \U$50402 ( \50377 , \50376 , \49947 );
and \U$50403 ( \50378 , \49938 , \49942 );
or \U$50404 ( \50379 , \50377 , \50378 );
buf \U$50405 ( \50380 , \50379 );
buf \U$50406 ( \50381 , \50380 );
xor \U$50407 ( \50382 , \48835 , \48839 );
xor \U$50408 ( \50383 , \50382 , \49234 );
buf \U$50409 ( \50384 , \50383 );
buf \U$50410 ( \50385 , \50384 );
xor \U$50411 ( \50386 , \50381 , \50385 );
xor \U$50412 ( \50387 , \49316 , \49320 );
xor \U$50413 ( \50388 , \50387 , \49325 );
buf \U$50414 ( \50389 , \50388 );
buf \U$50415 ( \50390 , \50389 );
xor \U$50416 ( \50391 , \50386 , \50390 );
buf \U$50417 ( \50392 , \50391 );
xor \U$50418 ( \50393 , \50375 , \50392 );
buf \U$50419 ( \50394 , \50393 );
xor \U$50420 ( \50395 , \49432 , \49854 );
xor \U$50421 ( \50396 , \50395 , \49880 );
buf \U$50422 ( \50397 , \50396 );
buf \U$50423 ( \50398 , \50397 );
xor \U$50424 ( \50399 , \49908 , \49922 );
xor \U$50425 ( \50400 , \50399 , \49927 );
buf \U$50426 ( \50401 , \50400 );
buf \U$50427 ( \50402 , \50401 );
not \U$50428 ( \50403 , \50402 );
buf \U$50429 ( \50404 , \49382 );
not \U$50430 ( \50405 , \50404 );
buf \U$50431 ( \50406 , \49403 );
not \U$50432 ( \50407 , \50406 );
or \U$50433 ( \50408 , \50405 , \50407 );
buf \U$50434 ( \50409 , \49390 );
buf \U$50435 ( \50410 , \49407 );
nand \U$50436 ( \50411 , \50409 , \50410 );
buf \U$50437 ( \50412 , \50411 );
buf \U$50438 ( \50413 , \50412 );
nand \U$50439 ( \50414 , \50408 , \50413 );
buf \U$50440 ( \50415 , \50414 );
buf \U$50441 ( \50416 , \50415 );
buf \U$50442 ( \50417 , \49396 );
xor \U$50443 ( \50418 , \50416 , \50417 );
buf \U$50444 ( \50419 , \50418 );
buf \U$50445 ( \50420 , \50419 );
xor \U$50446 ( \50421 , \49837 , \49829 );
buf \U$50447 ( \50422 , \50421 );
buf \U$50448 ( \50423 , \49833 );
xor \U$50449 ( \50424 , \50422 , \50423 );
buf \U$50450 ( \50425 , \50424 );
buf \U$50451 ( \50426 , \50425 );
xor \U$50452 ( \50427 , \50420 , \50426 );
xor \U$50453 ( \50428 , RIc0da738_105, RIc0d8fc8_55);
buf \U$50454 ( \50429 , \50428 );
not \U$50455 ( \50430 , \50429 );
buf \U$50456 ( \50431 , \12736 );
not \U$50457 ( \50432 , \50431 );
or \U$50458 ( \50433 , \50430 , \50432 );
buf \U$50459 ( \50434 , \49580 );
not \U$50460 ( \50435 , \50434 );
buf \U$50461 ( \50436 , \15653 );
nand \U$50462 ( \50437 , \50435 , \50436 );
buf \U$50463 ( \50438 , \50437 );
buf \U$50464 ( \50439 , \50438 );
nand \U$50465 ( \50440 , \50433 , \50439 );
buf \U$50466 ( \50441 , \50440 );
buf \U$50467 ( \50442 , \50441 );
xor \U$50468 ( \50443 , RIc0dacd8_117, RIc0d8a28_43);
buf \U$50469 ( \50444 , \50443 );
not \U$50470 ( \50445 , \50444 );
buf \U$50471 ( \50446 , \12929 );
not \U$50472 ( \50447 , \50446 );
or \U$50473 ( \50448 , \50445 , \50447 );
buf \U$50474 ( \50449 , \12937 );
buf \U$50475 ( \50450 , \49442 );
nand \U$50476 ( \50451 , \50449 , \50450 );
buf \U$50477 ( \50452 , \50451 );
buf \U$50478 ( \50453 , \50452 );
nand \U$50479 ( \50454 , \50448 , \50453 );
buf \U$50480 ( \50455 , \50454 );
buf \U$50481 ( \50456 , \50455 );
xor \U$50482 ( \50457 , \50442 , \50456 );
buf \U$50483 ( \50458 , RIc0d9400_64);
buf \U$50484 ( \50459 , RIc0da3f0_98);
or \U$50485 ( \50460 , \50458 , \50459 );
buf \U$50486 ( \50461 , RIc0da468_99);
nand \U$50487 ( \50462 , \50460 , \50461 );
buf \U$50488 ( \50463 , \50462 );
buf \U$50489 ( \50464 , \50463 );
buf \U$50490 ( \50465 , RIc0d9400_64);
buf \U$50491 ( \50466 , RIc0da3f0_98);
nand \U$50492 ( \50467 , \50465 , \50466 );
buf \U$50493 ( \50468 , \50467 );
buf \U$50494 ( \50469 , \50468 );
buf \U$50495 ( \50470 , RIc0da378_97);
and \U$50496 ( \50471 , \50464 , \50469 , \50470 );
buf \U$50497 ( \50472 , \50471 );
buf \U$50498 ( \50473 , \50472 );
buf \U$50499 ( \50474 , RIc0da468_99);
buf \U$50500 ( \50475 , RIc0d9310_62);
xor \U$50501 ( \50476 , \50474 , \50475 );
buf \U$50502 ( \50477 , \50476 );
buf \U$50503 ( \50478 , \50477 );
not \U$50504 ( \50479 , \50478 );
buf \U$50505 ( \50480 , \16744 );
not \U$50506 ( \50481 , \50480 );
or \U$50507 ( \50482 , \50479 , \50481 );
buf \U$50508 ( \50483 , \12584 );
buf \U$50509 ( \50484 , \50069 );
nand \U$50510 ( \50485 , \50483 , \50484 );
buf \U$50511 ( \50486 , \50485 );
buf \U$50512 ( \50487 , \50486 );
nand \U$50513 ( \50488 , \50482 , \50487 );
buf \U$50514 ( \50489 , \50488 );
buf \U$50515 ( \50490 , \50489 );
and \U$50516 ( \50491 , \50473 , \50490 );
buf \U$50517 ( \50492 , \50491 );
buf \U$50518 ( \50493 , \50492 );
and \U$50519 ( \50494 , \50457 , \50493 );
and \U$50520 ( \50495 , \50442 , \50456 );
or \U$50521 ( \50496 , \50494 , \50495 );
buf \U$50522 ( \50497 , \50496 );
buf \U$50523 ( \50498 , \50497 );
buf \U$50524 ( \50499 , RIc0daeb8_121);
buf \U$50525 ( \50500 , RIc0d88c0_40);
xor \U$50526 ( \50501 , \50499 , \50500 );
buf \U$50527 ( \50502 , \50501 );
buf \U$50528 ( \50503 , \50502 );
not \U$50529 ( \50504 , \50503 );
buf \U$50530 ( \50505 , \15420 );
not \U$50531 ( \50506 , \50505 );
or \U$50532 ( \50507 , \50504 , \50506 );
buf \U$50533 ( \50508 , \12975 );
buf \U$50534 ( \50509 , \50172 );
nand \U$50535 ( \50510 , \50508 , \50509 );
buf \U$50536 ( \50511 , \50510 );
buf \U$50537 ( \50512 , \50511 );
nand \U$50538 ( \50513 , \50507 , \50512 );
buf \U$50539 ( \50514 , \50513 );
not \U$50540 ( \50515 , \50514 );
xor \U$50541 ( \50516 , RIc0daa08_111, RIc0d8d70_50);
buf \U$50542 ( \50517 , \50516 );
not \U$50543 ( \50518 , \50517 );
buf \U$50544 ( \50519 , \14346 );
not \U$50545 ( \50520 , \50519 );
or \U$50546 ( \50521 , \50518 , \50520 );
buf \U$50547 ( \50522 , \14106 );
buf \U$50548 ( \50523 , \50105 );
nand \U$50549 ( \50524 , \50522 , \50523 );
buf \U$50550 ( \50525 , \50524 );
buf \U$50551 ( \50526 , \50525 );
nand \U$50552 ( \50527 , \50521 , \50526 );
buf \U$50553 ( \50528 , \50527 );
not \U$50554 ( \50529 , \50528 );
or \U$50555 ( \50530 , \50515 , \50529 );
buf \U$50556 ( \50531 , \50528 );
not \U$50557 ( \50532 , \50531 );
buf \U$50558 ( \50533 , \50532 );
not \U$50559 ( \50534 , \50533 );
buf \U$50560 ( \50535 , \50514 );
not \U$50561 ( \50536 , \50535 );
buf \U$50562 ( \50537 , \50536 );
not \U$50563 ( \50538 , \50537 );
or \U$50564 ( \50539 , \50534 , \50538 );
buf \U$50565 ( \50540 , RIc0d86e0_36);
buf \U$50566 ( \50541 , RIc0db098_125);
xor \U$50567 ( \50542 , \50540 , \50541 );
buf \U$50568 ( \50543 , \50542 );
buf \U$50569 ( \50544 , \50543 );
not \U$50570 ( \50545 , \50544 );
buf \U$50571 ( \50546 , \13461 );
not \U$50572 ( \50547 , \50546 );
or \U$50573 ( \50548 , \50545 , \50547 );
buf \U$50574 ( \50549 , \13465 );
buf \U$50575 ( \50550 , \50091 );
nand \U$50576 ( \50551 , \50549 , \50550 );
buf \U$50577 ( \50552 , \50551 );
buf \U$50578 ( \50553 , \50552 );
nand \U$50579 ( \50554 , \50548 , \50553 );
buf \U$50580 ( \50555 , \50554 );
nand \U$50581 ( \50556 , \50539 , \50555 );
nand \U$50582 ( \50557 , \50530 , \50556 );
buf \U$50583 ( \50558 , \50557 );
buf \U$50584 ( \50559 , RIc0d85f0_34);
buf \U$50585 ( \50560 , RIc0db188_127);
xor \U$50586 ( \50561 , \50559 , \50560 );
buf \U$50587 ( \50562 , \50561 );
buf \U$50588 ( \50563 , \50562 );
not \U$50589 ( \50564 , \50563 );
buf \U$50590 ( \50565 , \46813 );
not \U$50591 ( \50566 , \50565 );
or \U$50592 ( \50567 , \50564 , \50566 );
buf \U$50593 ( \50568 , \50051 );
buf \U$50594 ( \50569 , RIc0db200_128);
nand \U$50595 ( \50570 , \50568 , \50569 );
buf \U$50596 ( \50571 , \50570 );
buf \U$50597 ( \50572 , \50571 );
nand \U$50598 ( \50573 , \50567 , \50572 );
buf \U$50599 ( \50574 , \50573 );
buf \U$50600 ( \50575 , \50574 );
xor \U$50601 ( \50576 , RIc0da558_101, RIc0d9220_60);
buf \U$50602 ( \50577 , \50576 );
not \U$50603 ( \50578 , \50577 );
buf \U$50604 ( \50579 , \12833 );
not \U$50605 ( \50580 , \50579 );
or \U$50606 ( \50581 , \50578 , \50580 );
buf \U$50607 ( \50582 , \16676 );
buf \U$50608 ( \50583 , \50157 );
nand \U$50609 ( \50584 , \50582 , \50583 );
buf \U$50610 ( \50585 , \50584 );
buf \U$50611 ( \50586 , \50585 );
nand \U$50612 ( \50587 , \50581 , \50586 );
buf \U$50613 ( \50588 , \50587 );
buf \U$50614 ( \50589 , \50588 );
xor \U$50615 ( \50590 , \50575 , \50589 );
buf \U$50616 ( \50591 , RIc0dadc8_119);
buf \U$50617 ( \50592 , RIc0d89b0_42);
xor \U$50618 ( \50593 , \50591 , \50592 );
buf \U$50619 ( \50594 , \50593 );
buf \U$50620 ( \50595 , \50594 );
not \U$50621 ( \50596 , \50595 );
buf \U$50622 ( \50597 , \14569 );
not \U$50623 ( \50598 , \50597 );
or \U$50624 ( \50599 , \50596 , \50598 );
buf \U$50625 ( \50600 , \50192 );
not \U$50626 ( \50601 , \50600 );
buf \U$50627 ( \50602 , \13953 );
nand \U$50628 ( \50603 , \50601 , \50602 );
buf \U$50629 ( \50604 , \50603 );
buf \U$50630 ( \50605 , \50604 );
nand \U$50631 ( \50606 , \50599 , \50605 );
buf \U$50632 ( \50607 , \50606 );
buf \U$50633 ( \50608 , \50607 );
and \U$50634 ( \50609 , \50590 , \50608 );
and \U$50635 ( \50610 , \50575 , \50589 );
or \U$50636 ( \50611 , \50609 , \50610 );
buf \U$50637 ( \50612 , \50611 );
buf \U$50638 ( \50613 , \50612 );
xor \U$50639 ( \50614 , \50558 , \50613 );
xor \U$50640 ( \50615 , RIc0daaf8_113, RIc0d8c80_48);
buf \U$50641 ( \50616 , \50615 );
not \U$50642 ( \50617 , \50616 );
buf \U$50643 ( \50618 , \26484 );
not \U$50644 ( \50619 , \50618 );
or \U$50645 ( \50620 , \50617 , \50619 );
buf \U$50646 ( \50621 , \12410 );
buf \U$50647 ( \50622 , \49997 );
nand \U$50648 ( \50623 , \50621 , \50622 );
buf \U$50649 ( \50624 , \50623 );
buf \U$50650 ( \50625 , \50624 );
nand \U$50651 ( \50626 , \50620 , \50625 );
buf \U$50652 ( \50627 , \50626 );
buf \U$50653 ( \50628 , \50627 );
buf \U$50654 ( \50629 , RIc0d8aa0_44);
buf \U$50655 ( \50630 , RIc0dacd8_117);
xor \U$50656 ( \50631 , \50629 , \50630 );
buf \U$50657 ( \50632 , \50631 );
buf \U$50658 ( \50633 , \50632 );
not \U$50659 ( \50634 , \50633 );
buf \U$50660 ( \50635 , \13146 );
not \U$50661 ( \50636 , \50635 );
or \U$50662 ( \50637 , \50634 , \50636 );
buf \U$50663 ( \50638 , \22356 );
buf \U$50664 ( \50639 , \50443 );
nand \U$50665 ( \50640 , \50638 , \50639 );
buf \U$50666 ( \50641 , \50640 );
buf \U$50667 ( \50642 , \50641 );
nand \U$50668 ( \50643 , \50637 , \50642 );
buf \U$50669 ( \50644 , \50643 );
buf \U$50670 ( \50645 , \50644 );
nor \U$50671 ( \50646 , \50628 , \50645 );
buf \U$50672 ( \50647 , \50646 );
buf \U$50673 ( \50648 , \50647 );
buf \U$50674 ( \50649 , RIc0da738_105);
buf \U$50675 ( \50650 , RIc0d9040_56);
xor \U$50676 ( \50651 , \50649 , \50650 );
buf \U$50677 ( \50652 , \50651 );
buf \U$50678 ( \50653 , \50652 );
not \U$50679 ( \50654 , \50653 );
buf \U$50680 ( \50655 , \12736 );
not \U$50681 ( \50656 , \50655 );
or \U$50682 ( \50657 , \50654 , \50656 );
buf \U$50683 ( \50658 , \12744 );
buf \U$50684 ( \50659 , \50428 );
nand \U$50685 ( \50660 , \50658 , \50659 );
buf \U$50686 ( \50661 , \50660 );
buf \U$50687 ( \50662 , \50661 );
nand \U$50688 ( \50663 , \50657 , \50662 );
buf \U$50689 ( \50664 , \50663 );
buf \U$50690 ( \50665 , \50664 );
not \U$50691 ( \50666 , \50665 );
buf \U$50692 ( \50667 , \50666 );
buf \U$50693 ( \50668 , \50667 );
or \U$50694 ( \50669 , \50648 , \50668 );
buf \U$50695 ( \50670 , \50627 );
buf \U$50696 ( \50671 , \50644 );
nand \U$50697 ( \50672 , \50670 , \50671 );
buf \U$50698 ( \50673 , \50672 );
buf \U$50699 ( \50674 , \50673 );
nand \U$50700 ( \50675 , \50669 , \50674 );
buf \U$50701 ( \50676 , \50675 );
buf \U$50702 ( \50677 , \50676 );
and \U$50703 ( \50678 , \50614 , \50677 );
and \U$50704 ( \50679 , \50558 , \50613 );
or \U$50705 ( \50680 , \50678 , \50679 );
buf \U$50706 ( \50681 , \50680 );
buf \U$50707 ( \50682 , \50681 );
xor \U$50708 ( \50683 , \50498 , \50682 );
xor \U$50709 ( \50684 , \49967 , \49978 );
xor \U$50710 ( \50685 , \50684 , \50040 );
buf \U$50711 ( \50686 , \50685 );
buf \U$50712 ( \50687 , \50686 );
and \U$50713 ( \50688 , \50683 , \50687 );
and \U$50714 ( \50689 , \50498 , \50682 );
or \U$50715 ( \50690 , \50688 , \50689 );
buf \U$50716 ( \50691 , \50690 );
buf \U$50717 ( \50692 , \50691 );
and \U$50718 ( \50693 , \50427 , \50692 );
and \U$50719 ( \50694 , \50420 , \50426 );
or \U$50720 ( \50695 , \50693 , \50694 );
buf \U$50721 ( \50696 , \50695 );
buf \U$50722 ( \50697 , \50696 );
not \U$50723 ( \50698 , \50697 );
or \U$50724 ( \50699 , \50403 , \50698 );
buf \U$50725 ( \50700 , \50696 );
buf \U$50726 ( \50701 , \50401 );
or \U$50727 ( \50702 , \50700 , \50701 );
xor \U$50728 ( \50703 , \50044 , \50212 );
xnor \U$50729 ( \50704 , \50703 , \50220 );
buf \U$50730 ( \50705 , \50704 );
not \U$50731 ( \50706 , \50705 );
buf \U$50732 ( \50707 , RIc0d8b90_46);
buf \U$50733 ( \50708 , RIc0dabe8_115);
xor \U$50734 ( \50709 , \50707 , \50708 );
buf \U$50735 ( \50710 , \50709 );
buf \U$50736 ( \50711 , \50710 );
not \U$50737 ( \50712 , \50711 );
buf \U$50738 ( \50713 , \14684 );
not \U$50739 ( \50714 , \50713 );
or \U$50740 ( \50715 , \50712 , \50714 );
buf \U$50741 ( \50716 , \14690 );
buf \U$50742 ( \50717 , \49980 );
nand \U$50743 ( \50718 , \50716 , \50717 );
buf \U$50744 ( \50719 , \50718 );
buf \U$50745 ( \50720 , \50719 );
nand \U$50746 ( \50721 , \50715 , \50720 );
buf \U$50747 ( \50722 , \50721 );
buf \U$50748 ( \50723 , \50722 );
buf \U$50749 ( \50724 , RIc0d8e60_52);
buf \U$50750 ( \50725 , RIc0da918_109);
xor \U$50751 ( \50726 , \50724 , \50725 );
buf \U$50752 ( \50727 , \50726 );
buf \U$50753 ( \50728 , \50727 );
not \U$50754 ( \50729 , \50728 );
buf \U$50755 ( \50730 , \21959 );
not \U$50756 ( \50731 , \50730 );
or \U$50757 ( \50732 , \50729 , \50731 );
buf \U$50758 ( \50733 , \20211 );
buf \U$50759 ( \50734 , \50279 );
nand \U$50760 ( \50735 , \50733 , \50734 );
buf \U$50761 ( \50736 , \50735 );
buf \U$50762 ( \50737 , \50736 );
nand \U$50763 ( \50738 , \50732 , \50737 );
buf \U$50764 ( \50739 , \50738 );
buf \U$50765 ( \50740 , \50739 );
nor \U$50766 ( \50741 , \50723 , \50740 );
buf \U$50767 ( \50742 , \50741 );
buf \U$50768 ( \50743 , \50742 );
buf \U$50769 ( \50744 , RIc0d9130_58);
buf \U$50770 ( \50745 , RIc0da648_103);
xor \U$50771 ( \50746 , \50744 , \50745 );
buf \U$50772 ( \50747 , \50746 );
buf \U$50773 ( \50748 , \50747 );
not \U$50774 ( \50749 , \50748 );
buf \U$50775 ( \50750 , \29546 );
not \U$50776 ( \50751 , \50750 );
or \U$50777 ( \50752 , \50749 , \50751 );
buf \U$50778 ( \50753 , \50020 );
not \U$50779 ( \50754 , \50753 );
buf \U$50780 ( \50755 , \13048 );
nand \U$50781 ( \50756 , \50754 , \50755 );
buf \U$50782 ( \50757 , \50756 );
buf \U$50783 ( \50758 , \50757 );
nand \U$50784 ( \50759 , \50752 , \50758 );
buf \U$50785 ( \50760 , \50759 );
buf \U$50786 ( \50761 , \50760 );
not \U$50787 ( \50762 , \50761 );
buf \U$50788 ( \50763 , \50762 );
buf \U$50789 ( \50764 , \50763 );
or \U$50790 ( \50765 , \50743 , \50764 );
buf \U$50791 ( \50766 , \50722 );
buf \U$50792 ( \50767 , \50739 );
nand \U$50793 ( \50768 , \50766 , \50767 );
buf \U$50794 ( \50769 , \50768 );
buf \U$50795 ( \50770 , \50769 );
nand \U$50796 ( \50771 , \50765 , \50770 );
buf \U$50797 ( \50772 , \50771 );
buf \U$50798 ( \50773 , \50772 );
xor \U$50799 ( \50774 , \50062 , \50067 );
xor \U$50800 ( \50775 , \50774 , \50082 );
buf \U$50801 ( \50776 , \50775 );
buf \U$50802 ( \50777 , \50776 );
or \U$50803 ( \50778 , \50773 , \50777 );
xor \U$50804 ( \50779 , RIc0dafa8_123, RIc0d87d0_38);
buf \U$50805 ( \50780 , \50779 );
not \U$50806 ( \50781 , \50780 );
buf \U$50807 ( \50782 , \14982 );
not \U$50808 ( \50783 , \50782 );
or \U$50809 ( \50784 , \50781 , \50783 );
buf \U$50810 ( \50785 , \16692 );
buf \U$50811 ( \50786 , \50127 );
nand \U$50812 ( \50787 , \50785 , \50786 );
buf \U$50813 ( \50788 , \50787 );
buf \U$50814 ( \50789 , \50788 );
nand \U$50815 ( \50790 , \50784 , \50789 );
buf \U$50816 ( \50791 , \50790 );
buf \U$50817 ( \50792 , \50791 );
not \U$50818 ( \50793 , \50792 );
buf \U$50819 ( \50794 , \50793 );
buf \U$50820 ( \50795 , \50794 );
not \U$50821 ( \50796 , \50795 );
buf \U$50822 ( \50797 , RIc0da828_107);
buf \U$50823 ( \50798 , RIc0d8f50_54);
xor \U$50824 ( \50799 , \50797 , \50798 );
buf \U$50825 ( \50800 , \50799 );
buf \U$50826 ( \50801 , \50800 );
not \U$50827 ( \50802 , \50801 );
buf \U$50828 ( \50803 , \21898 );
not \U$50829 ( \50804 , \50803 );
or \U$50830 ( \50805 , \50802 , \50804 );
buf \U$50831 ( \50806 , \12342 );
buf \U$50832 ( \50807 , \50265 );
nand \U$50833 ( \50808 , \50806 , \50807 );
buf \U$50834 ( \50809 , \50808 );
buf \U$50835 ( \50810 , \50809 );
nand \U$50836 ( \50811 , \50805 , \50810 );
buf \U$50837 ( \50812 , \50811 );
buf \U$50838 ( \50813 , \50812 );
not \U$50839 ( \50814 , \50813 );
buf \U$50840 ( \50815 , \50814 );
buf \U$50841 ( \50816 , \50815 );
not \U$50842 ( \50817 , \50816 );
or \U$50843 ( \50818 , \50796 , \50817 );
buf \U$50844 ( \50819 , RIc0d9400_64);
buf \U$50845 ( \50820 , RIc0da378_97);
xor \U$50846 ( \50821 , \50819 , \50820 );
buf \U$50847 ( \50822 , \50821 );
buf \U$50848 ( \50823 , \50822 );
not \U$50849 ( \50824 , \50823 );
buf \U$50850 ( \50825 , \2941 );
not \U$50851 ( \50826 , \50825 );
or \U$50852 ( \50827 , \50824 , \50826 );
buf \U$50853 ( \50828 , \734 );
buf \U$50854 ( \50829 , \50301 );
nand \U$50855 ( \50830 , \50828 , \50829 );
buf \U$50856 ( \50831 , \50830 );
buf \U$50857 ( \50832 , \50831 );
nand \U$50858 ( \50833 , \50827 , \50832 );
buf \U$50859 ( \50834 , \50833 );
buf \U$50860 ( \50835 , \50834 );
nand \U$50861 ( \50836 , \50818 , \50835 );
buf \U$50862 ( \50837 , \50836 );
buf \U$50863 ( \50838 , \50837 );
buf \U$50864 ( \50839 , \50812 );
buf \U$50865 ( \50840 , \50791 );
nand \U$50866 ( \50841 , \50839 , \50840 );
buf \U$50867 ( \50842 , \50841 );
buf \U$50868 ( \50843 , \50842 );
nand \U$50869 ( \50844 , \50838 , \50843 );
buf \U$50870 ( \50845 , \50844 );
buf \U$50871 ( \50846 , \50845 );
nand \U$50872 ( \50847 , \50778 , \50846 );
buf \U$50873 ( \50848 , \50847 );
buf \U$50874 ( \50849 , \50848 );
buf \U$50875 ( \50850 , \50776 );
buf \U$50876 ( \50851 , \50772 );
nand \U$50877 ( \50852 , \50850 , \50851 );
buf \U$50878 ( \50853 , \50852 );
buf \U$50879 ( \50854 , \50853 );
nand \U$50880 ( \50855 , \50849 , \50854 );
buf \U$50881 ( \50856 , \50855 );
buf \U$50882 ( \50857 , \50856 );
xor \U$50883 ( \50858 , \50278 , \50292 );
xor \U$50884 ( \50859 , \50858 , \50314 );
buf \U$50885 ( \50860 , \50859 );
buf \U$50886 ( \50861 , \50860 );
buf \U$50887 ( \50862 , \50010 );
not \U$50888 ( \50863 , \50862 );
buf \U$50889 ( \50864 , \50863 );
buf \U$50890 ( \50865 , \50864 );
not \U$50891 ( \50866 , \50865 );
buf \U$50892 ( \50867 , \49992 );
not \U$50893 ( \50868 , \50867 );
buf \U$50894 ( \50869 , \50030 );
not \U$50895 ( \50870 , \50869 );
or \U$50896 ( \50871 , \50868 , \50870 );
buf \U$50897 ( \50872 , \49992 );
buf \U$50898 ( \50873 , \50030 );
or \U$50899 ( \50874 , \50872 , \50873 );
nand \U$50900 ( \50875 , \50871 , \50874 );
buf \U$50901 ( \50876 , \50875 );
buf \U$50902 ( \50877 , \50876 );
not \U$50903 ( \50878 , \50877 );
or \U$50904 ( \50879 , \50866 , \50878 );
buf \U$50905 ( \50880 , \50876 );
buf \U$50906 ( \50881 , \50864 );
or \U$50907 ( \50882 , \50880 , \50881 );
nand \U$50908 ( \50883 , \50879 , \50882 );
buf \U$50909 ( \50884 , \50883 );
buf \U$50910 ( \50885 , \50884 );
or \U$50911 ( \50886 , \50861 , \50885 );
xor \U$50912 ( \50887 , \50117 , \50103 );
xnor \U$50913 ( \50888 , \50887 , \50141 );
buf \U$50914 ( \50889 , \50888 );
nand \U$50915 ( \50890 , \50886 , \50889 );
buf \U$50916 ( \50891 , \50890 );
buf \U$50917 ( \50892 , \50891 );
buf \U$50918 ( \50893 , \50860 );
buf \U$50919 ( \50894 , \50884 );
nand \U$50920 ( \50895 , \50893 , \50894 );
buf \U$50921 ( \50896 , \50895 );
buf \U$50922 ( \50897 , \50896 );
nand \U$50923 ( \50898 , \50892 , \50897 );
buf \U$50924 ( \50899 , \50898 );
buf \U$50925 ( \50900 , \50899 );
xor \U$50926 ( \50901 , \50857 , \50900 );
xor \U$50927 ( \50902 , \50087 , \50151 );
xor \U$50928 ( \50903 , \50902 , \50208 );
buf \U$50929 ( \50904 , \50903 );
buf \U$50930 ( \50905 , \50904 );
and \U$50931 ( \50906 , \50901 , \50905 );
and \U$50932 ( \50907 , \50857 , \50900 );
or \U$50933 ( \50908 , \50906 , \50907 );
buf \U$50934 ( \50909 , \50908 );
buf \U$50935 ( \50910 , \50909 );
not \U$50936 ( \50911 , \50910 );
buf \U$50937 ( \50912 , \50911 );
buf \U$50938 ( \50913 , \50912 );
not \U$50939 ( \50914 , \50913 );
or \U$50940 ( \50915 , \50706 , \50914 );
buf \U$50941 ( \50916 , \50350 );
not \U$50942 ( \50917 , \50916 );
buf \U$50943 ( \50918 , \50324 );
not \U$50944 ( \50919 , \50918 );
or \U$50945 ( \50920 , \50917 , \50919 );
buf \U$50946 ( \50921 , \50324 );
buf \U$50947 ( \50922 , \50350 );
or \U$50948 ( \50923 , \50921 , \50922 );
nand \U$50949 ( \50924 , \50920 , \50923 );
buf \U$50950 ( \50925 , \50924 );
buf \U$50951 ( \50926 , \50925 );
buf \U$50952 ( \50927 , \50340 );
and \U$50953 ( \50928 , \50926 , \50927 );
not \U$50954 ( \50929 , \50926 );
buf \U$50955 ( \50930 , \50340 );
not \U$50956 ( \50931 , \50930 );
buf \U$50957 ( \50932 , \50931 );
buf \U$50958 ( \50933 , \50932 );
and \U$50959 ( \50934 , \50929 , \50933 );
nor \U$50960 ( \50935 , \50928 , \50934 );
buf \U$50961 ( \50936 , \50935 );
buf \U$50962 ( \50937 , \50936 );
nand \U$50963 ( \50938 , \50915 , \50937 );
buf \U$50964 ( \50939 , \50938 );
buf \U$50965 ( \50940 , \50939 );
buf \U$50966 ( \50941 , \50704 );
not \U$50967 ( \50942 , \50941 );
buf \U$50968 ( \50943 , \50909 );
nand \U$50969 ( \50944 , \50942 , \50943 );
buf \U$50970 ( \50945 , \50944 );
buf \U$50971 ( \50946 , \50945 );
nand \U$50972 ( \50947 , \50940 , \50946 );
buf \U$50973 ( \50948 , \50947 );
buf \U$50974 ( \50949 , \50948 );
nand \U$50975 ( \50950 , \50702 , \50949 );
buf \U$50976 ( \50951 , \50950 );
buf \U$50977 ( \50952 , \50951 );
nand \U$50978 ( \50953 , \50699 , \50952 );
buf \U$50979 ( \50954 , \50953 );
buf \U$50980 ( \50955 , \50954 );
or \U$50981 ( \50956 , \50398 , \50955 );
xor \U$50982 ( \50957 , \49932 , \49950 );
xor \U$50983 ( \50958 , \50957 , \50370 );
buf \U$50984 ( \50959 , \50958 );
buf \U$50985 ( \50960 , \50959 );
nand \U$50986 ( \50961 , \50956 , \50960 );
buf \U$50987 ( \50962 , \50961 );
buf \U$50988 ( \50963 , \50962 );
buf \U$50989 ( \50964 , \50954 );
buf \U$50990 ( \50965 , \50397 );
nand \U$50991 ( \50966 , \50964 , \50965 );
buf \U$50992 ( \50967 , \50966 );
buf \U$50993 ( \50968 , \50967 );
nand \U$50994 ( \50969 , \50963 , \50968 );
buf \U$50995 ( \50970 , \50969 );
buf \U$50996 ( \50971 , \50970 );
not \U$50997 ( \50972 , \50971 );
buf \U$50998 ( \50973 , \50972 );
buf \U$50999 ( \50974 , \50973 );
nand \U$51000 ( \50975 , \50394 , \50974 );
buf \U$51001 ( \50976 , \50975 );
buf \U$51002 ( \50977 , \50976 );
xor \U$51003 ( \50978 , \50227 , \50360 );
xor \U$51004 ( \50979 , \50978 , \50365 );
buf \U$51005 ( \50980 , \50979 );
buf \U$51006 ( \50981 , \50980 );
xor \U$51007 ( \50982 , \50328 , \50332 );
xor \U$51008 ( \50983 , \50982 , \50336 );
buf \U$51009 ( \50984 , \50983 );
buf \U$51010 ( \50985 , \50984 );
xor \U$51011 ( \50986 , \50171 , \50186 );
xor \U$51012 ( \50987 , \50986 , \50203 );
buf \U$51013 ( \50988 , \50987 );
buf \U$51014 ( \50989 , \50988 );
xor \U$51015 ( \50990 , \50442 , \50456 );
xor \U$51016 ( \50991 , \50990 , \50493 );
buf \U$51017 ( \50992 , \50991 );
buf \U$51018 ( \50993 , \50992 );
xor \U$51019 ( \50994 , \50989 , \50993 );
xor \U$51020 ( \50995 , \50473 , \50490 );
buf \U$51021 ( \50996 , \50995 );
buf \U$51022 ( \50997 , \50996 );
buf \U$51023 ( \50998 , RIc0dadc8_119);
buf \U$51024 ( \50999 , RIc0d8a28_43);
xor \U$51025 ( \51000 , \50998 , \50999 );
buf \U$51026 ( \51001 , \51000 );
buf \U$51027 ( \51002 , \51001 );
not \U$51028 ( \51003 , \51002 );
buf \U$51029 ( \51004 , \23985 );
not \U$51030 ( \51005 , \51004 );
or \U$51031 ( \51006 , \51003 , \51005 );
buf \U$51032 ( \51007 , \13005 );
buf \U$51033 ( \51008 , \50594 );
nand \U$51034 ( \51009 , \51007 , \51008 );
buf \U$51035 ( \51010 , \51009 );
buf \U$51036 ( \51011 , \51010 );
nand \U$51037 ( \51012 , \51006 , \51011 );
buf \U$51038 ( \51013 , \51012 );
buf \U$51039 ( \51014 , \51013 );
not \U$51040 ( \51015 , \51014 );
buf \U$51041 ( \51016 , \51015 );
buf \U$51042 ( \51017 , \51016 );
not \U$51043 ( \51018 , \51017 );
buf \U$51044 ( \51019 , RIc0d8fc8_55);
buf \U$51045 ( \51020 , RIc0da828_107);
xor \U$51046 ( \51021 , \51019 , \51020 );
buf \U$51047 ( \51022 , \51021 );
buf \U$51048 ( \51023 , \51022 );
not \U$51049 ( \51024 , \51023 );
buf \U$51050 ( \51025 , \19414 );
not \U$51051 ( \51026 , \51025 );
or \U$51052 ( \51027 , \51024 , \51026 );
buf \U$51053 ( \51028 , \12342 );
buf \U$51054 ( \51029 , \50800 );
nand \U$51055 ( \51030 , \51028 , \51029 );
buf \U$51056 ( \51031 , \51030 );
buf \U$51057 ( \51032 , \51031 );
nand \U$51058 ( \51033 , \51027 , \51032 );
buf \U$51059 ( \51034 , \51033 );
buf \U$51060 ( \51035 , \51034 );
not \U$51061 ( \51036 , \51035 );
buf \U$51062 ( \51037 , \51036 );
buf \U$51063 ( \51038 , \51037 );
not \U$51064 ( \51039 , \51038 );
or \U$51065 ( \51040 , \51018 , \51039 );
buf \U$51066 ( \51041 , RIc0d91a8_59);
buf \U$51067 ( \51042 , RIc0da648_103);
xor \U$51068 ( \51043 , \51041 , \51042 );
buf \U$51069 ( \51044 , \51043 );
buf \U$51070 ( \51045 , \51044 );
not \U$51071 ( \51046 , \51045 );
buf \U$51072 ( \51047 , \17405 );
not \U$51073 ( \51048 , \51047 );
or \U$51074 ( \51049 , \51046 , \51048 );
buf \U$51075 ( \51050 , \18416 );
buf \U$51076 ( \51051 , \50747 );
nand \U$51077 ( \51052 , \51050 , \51051 );
buf \U$51078 ( \51053 , \51052 );
buf \U$51079 ( \51054 , \51053 );
nand \U$51080 ( \51055 , \51049 , \51054 );
buf \U$51081 ( \51056 , \51055 );
buf \U$51082 ( \51057 , \51056 );
nand \U$51083 ( \51058 , \51040 , \51057 );
buf \U$51084 ( \51059 , \51058 );
buf \U$51085 ( \51060 , \51059 );
buf \U$51086 ( \51061 , \51034 );
buf \U$51087 ( \51062 , \51013 );
nand \U$51088 ( \51063 , \51061 , \51062 );
buf \U$51089 ( \51064 , \51063 );
buf \U$51090 ( \51065 , \51064 );
nand \U$51091 ( \51066 , \51060 , \51065 );
buf \U$51092 ( \51067 , \51066 );
buf \U$51093 ( \51068 , \51067 );
xor \U$51094 ( \51069 , \50997 , \51068 );
buf \U$51095 ( \51070 , \734 );
buf \U$51096 ( \51071 , RIc0d9400_64);
and \U$51097 ( \51072 , \51070 , \51071 );
buf \U$51098 ( \51073 , \51072 );
buf \U$51099 ( \51074 , \51073 );
xor \U$51100 ( \51075 , RIc0da558_101, RIc0d9298_61);
buf \U$51101 ( \51076 , \51075 );
not \U$51102 ( \51077 , \51076 );
buf \U$51103 ( \51078 , \3535 );
not \U$51104 ( \51079 , \51078 );
or \U$51105 ( \51080 , \51077 , \51079 );
buf \U$51106 ( \51081 , \16676 );
buf \U$51107 ( \51082 , \50576 );
nand \U$51108 ( \51083 , \51081 , \51082 );
buf \U$51109 ( \51084 , \51083 );
buf \U$51110 ( \51085 , \51084 );
nand \U$51111 ( \51086 , \51080 , \51085 );
buf \U$51112 ( \51087 , \51086 );
buf \U$51113 ( \51088 , \51087 );
xor \U$51114 ( \51089 , \51074 , \51088 );
xor \U$51115 ( \51090 , RIc0db098_125, RIc0d8758_37);
buf \U$51116 ( \51091 , \51090 );
not \U$51117 ( \51092 , \51091 );
buf \U$51118 ( \51093 , \17992 );
not \U$51119 ( \51094 , \51093 );
buf \U$51120 ( \51095 , \51094 );
buf \U$51121 ( \51096 , \51095 );
not \U$51122 ( \51097 , \51096 );
or \U$51123 ( \51098 , \51092 , \51097 );
buf \U$51124 ( \51099 , \15793 );
buf \U$51125 ( \51100 , \50543 );
nand \U$51126 ( \51101 , \51099 , \51100 );
buf \U$51127 ( \51102 , \51101 );
buf \U$51128 ( \51103 , \51102 );
nand \U$51129 ( \51104 , \51098 , \51103 );
buf \U$51130 ( \51105 , \51104 );
buf \U$51131 ( \51106 , \51105 );
and \U$51132 ( \51107 , \51089 , \51106 );
and \U$51133 ( \51108 , \51074 , \51088 );
or \U$51134 ( \51109 , \51107 , \51108 );
buf \U$51135 ( \51110 , \51109 );
buf \U$51136 ( \51111 , \51110 );
and \U$51137 ( \51112 , \51069 , \51111 );
and \U$51138 ( \51113 , \50997 , \51068 );
or \U$51139 ( \51114 , \51112 , \51113 );
buf \U$51140 ( \51115 , \51114 );
buf \U$51141 ( \51116 , \51115 );
and \U$51142 ( \51117 , \50994 , \51116 );
and \U$51143 ( \51118 , \50989 , \50993 );
or \U$51144 ( \51119 , \51117 , \51118 );
buf \U$51145 ( \51120 , \51119 );
buf \U$51146 ( \51121 , \51120 );
xor \U$51147 ( \51122 , \50985 , \51121 );
buf \U$51148 ( \51123 , \50318 );
not \U$51149 ( \51124 , \51123 );
buf \U$51150 ( \51125 , \50229 );
not \U$51151 ( \51126 , \51125 );
or \U$51152 ( \51127 , \51124 , \51126 );
buf \U$51153 ( \51128 , \50318 );
buf \U$51154 ( \51129 , \50229 );
or \U$51155 ( \51130 , \51128 , \51129 );
nand \U$51156 ( \51131 , \51127 , \51130 );
buf \U$51157 ( \51132 , \51131 );
buf \U$51158 ( \51133 , \51132 );
buf \U$51159 ( \51134 , \50253 );
and \U$51160 ( \51135 , \51133 , \51134 );
not \U$51161 ( \51136 , \51133 );
buf \U$51162 ( \51137 , \50250 );
and \U$51163 ( \51138 , \51136 , \51137 );
nor \U$51164 ( \51139 , \51135 , \51138 );
buf \U$51165 ( \51140 , \51139 );
buf \U$51166 ( \51141 , \51140 );
and \U$51167 ( \51142 , \51122 , \51141 );
and \U$51168 ( \51143 , \50985 , \51121 );
or \U$51169 ( \51144 , \51142 , \51143 );
buf \U$51170 ( \51145 , \51144 );
buf \U$51171 ( \51146 , \51145 );
xor \U$51172 ( \51147 , \50420 , \50426 );
xor \U$51173 ( \51148 , \51147 , \50692 );
buf \U$51174 ( \51149 , \51148 );
buf \U$51175 ( \51150 , \51149 );
xor \U$51176 ( \51151 , \51146 , \51150 );
xor \U$51177 ( \51152 , \50498 , \50682 );
xor \U$51178 ( \51153 , \51152 , \50687 );
buf \U$51179 ( \51154 , \51153 );
buf \U$51180 ( \51155 , \51154 );
buf \U$51181 ( \51156 , RIc0d8668_35);
buf \U$51182 ( \51157 , RIc0db188_127);
xor \U$51183 ( \51158 , \51156 , \51157 );
buf \U$51184 ( \51159 , \51158 );
buf \U$51185 ( \51160 , \51159 );
not \U$51186 ( \51161 , \51160 );
buf \U$51187 ( \51162 , \15609 );
not \U$51188 ( \51163 , \51162 );
or \U$51189 ( \51164 , \51161 , \51163 );
buf \U$51190 ( \51165 , \50562 );
buf \U$51191 ( \51166 , RIc0db200_128);
nand \U$51192 ( \51167 , \51165 , \51166 );
buf \U$51193 ( \51168 , \51167 );
buf \U$51194 ( \51169 , \51168 );
nand \U$51195 ( \51170 , \51164 , \51169 );
buf \U$51196 ( \51171 , \51170 );
buf \U$51197 ( \51172 , \51171 );
buf \U$51198 ( \51173 , RIc0d8cf8_49);
buf \U$51199 ( \51174 , RIc0daaf8_113);
xor \U$51200 ( \51175 , \51173 , \51174 );
buf \U$51201 ( \51176 , \51175 );
buf \U$51202 ( \51177 , \51176 );
not \U$51203 ( \51178 , \51177 );
buf \U$51204 ( \51179 , \28413 );
not \U$51205 ( \51180 , \51179 );
or \U$51206 ( \51181 , \51178 , \51180 );
buf \U$51207 ( \51182 , \14405 );
buf \U$51208 ( \51183 , \50615 );
nand \U$51209 ( \51184 , \51182 , \51183 );
buf \U$51210 ( \51185 , \51184 );
buf \U$51211 ( \51186 , \51185 );
nand \U$51212 ( \51187 , \51181 , \51186 );
buf \U$51213 ( \51188 , \51187 );
buf \U$51214 ( \51189 , \51188 );
xor \U$51215 ( \51190 , \51172 , \51189 );
buf \U$51216 ( \51191 , \50779 );
not \U$51217 ( \51192 , \51191 );
buf \U$51218 ( \51193 , \16692 );
not \U$51219 ( \51194 , \51193 );
or \U$51220 ( \51195 , \51192 , \51194 );
buf \U$51221 ( \51196 , \46183 );
buf \U$51222 ( \51197 , RIc0dafa8_123);
buf \U$51223 ( \51198 , RIc0d8848_39);
xnor \U$51224 ( \51199 , \51197 , \51198 );
buf \U$51225 ( \51200 , \51199 );
buf \U$51226 ( \51201 , \51200 );
or \U$51227 ( \51202 , \51196 , \51201 );
nand \U$51228 ( \51203 , \51195 , \51202 );
buf \U$51229 ( \51204 , \51203 );
buf \U$51230 ( \51205 , \51204 );
and \U$51231 ( \51206 , \51190 , \51205 );
and \U$51232 ( \51207 , \51172 , \51189 );
or \U$51233 ( \51208 , \51206 , \51207 );
buf \U$51234 ( \51209 , \51208 );
buf \U$51235 ( \51210 , \51209 );
buf \U$51236 ( \51211 , RIc0d90b8_57);
buf \U$51237 ( \51212 , RIc0da738_105);
xor \U$51238 ( \51213 , \51211 , \51212 );
buf \U$51239 ( \51214 , \51213 );
buf \U$51240 ( \51215 , \51214 );
not \U$51241 ( \51216 , \51215 );
buf \U$51242 ( \51217 , \25475 );
not \U$51243 ( \51218 , \51217 );
or \U$51244 ( \51219 , \51216 , \51218 );
buf \U$51245 ( \51220 , \12744 );
buf \U$51246 ( \51221 , \50652 );
nand \U$51247 ( \51222 , \51220 , \51221 );
buf \U$51248 ( \51223 , \51222 );
buf \U$51249 ( \51224 , \51223 );
nand \U$51250 ( \51225 , \51219 , \51224 );
buf \U$51251 ( \51226 , \51225 );
buf \U$51252 ( \51227 , \51226 );
not \U$51253 ( \51228 , \51227 );
buf \U$51254 ( \51229 , \51228 );
buf \U$51255 ( \51230 , \51229 );
not \U$51256 ( \51231 , \51230 );
buf \U$51257 ( \51232 , RIc0da468_99);
buf \U$51258 ( \51233 , RIc0d9388_63);
xor \U$51259 ( \51234 , \51232 , \51233 );
buf \U$51260 ( \51235 , \51234 );
buf \U$51261 ( \51236 , \51235 );
not \U$51262 ( \51237 , \51236 );
buf \U$51263 ( \51238 , \21461 );
not \U$51264 ( \51239 , \51238 );
or \U$51265 ( \51240 , \51237 , \51239 );
buf \U$51266 ( \51241 , \14140 );
buf \U$51267 ( \51242 , \50477 );
nand \U$51268 ( \51243 , \51241 , \51242 );
buf \U$51269 ( \51244 , \51243 );
buf \U$51270 ( \51245 , \51244 );
nand \U$51271 ( \51246 , \51240 , \51245 );
buf \U$51272 ( \51247 , \51246 );
buf \U$51273 ( \51248 , \51247 );
not \U$51274 ( \51249 , \51248 );
buf \U$51275 ( \51250 , \51249 );
buf \U$51276 ( \51251 , \51250 );
not \U$51277 ( \51252 , \51251 );
or \U$51278 ( \51253 , \51231 , \51252 );
buf \U$51279 ( \51254 , RIc0d8c08_47);
buf \U$51280 ( \51255 , RIc0dabe8_115);
xor \U$51281 ( \51256 , \51254 , \51255 );
buf \U$51282 ( \51257 , \51256 );
buf \U$51283 ( \51258 , \51257 );
not \U$51284 ( \51259 , \51258 );
buf \U$51285 ( \51260 , \14186 );
not \U$51286 ( \51261 , \51260 );
or \U$51287 ( \51262 , \51259 , \51261 );
buf \U$51288 ( \51263 , \12303 );
buf \U$51289 ( \51264 , \50710 );
nand \U$51290 ( \51265 , \51263 , \51264 );
buf \U$51291 ( \51266 , \51265 );
buf \U$51292 ( \51267 , \51266 );
nand \U$51293 ( \51268 , \51262 , \51267 );
buf \U$51294 ( \51269 , \51268 );
buf \U$51295 ( \51270 , \51269 );
nand \U$51296 ( \51271 , \51253 , \51270 );
buf \U$51297 ( \51272 , \51271 );
buf \U$51298 ( \51273 , \51272 );
buf \U$51299 ( \51274 , \51247 );
buf \U$51300 ( \51275 , \51226 );
nand \U$51301 ( \51276 , \51274 , \51275 );
buf \U$51302 ( \51277 , \51276 );
buf \U$51303 ( \51278 , \51277 );
nand \U$51304 ( \51279 , \51273 , \51278 );
buf \U$51305 ( \51280 , \51279 );
buf \U$51306 ( \51281 , \51280 );
xor \U$51307 ( \51282 , \51210 , \51281 );
buf \U$51308 ( \51283 , RIc0d8ed8_53);
buf \U$51309 ( \51284 , RIc0da918_109);
xor \U$51310 ( \51285 , \51283 , \51284 );
buf \U$51311 ( \51286 , \51285 );
buf \U$51312 ( \51287 , \51286 );
not \U$51313 ( \51288 , \51287 );
buf \U$51314 ( \51289 , \21959 );
not \U$51315 ( \51290 , \51289 );
or \U$51316 ( \51291 , \51288 , \51290 );
buf \U$51317 ( \51292 , \15909 );
buf \U$51318 ( \51293 , \50727 );
nand \U$51319 ( \51294 , \51292 , \51293 );
buf \U$51320 ( \51295 , \51294 );
buf \U$51321 ( \51296 , \51295 );
nand \U$51322 ( \51297 , \51291 , \51296 );
buf \U$51323 ( \51298 , \51297 );
buf \U$51324 ( \51299 , RIc0daa08_111);
buf \U$51325 ( \51300 , RIc0d8de8_51);
xor \U$51326 ( \51301 , \51299 , \51300 );
buf \U$51327 ( \51302 , \51301 );
buf \U$51328 ( \51303 , \51302 );
not \U$51329 ( \51304 , \51303 );
buf \U$51330 ( \51305 , \12529 );
not \U$51331 ( \51306 , \51305 );
or \U$51332 ( \51307 , \51304 , \51306 );
buf \U$51333 ( \51308 , \14353 );
buf \U$51334 ( \51309 , \50516 );
nand \U$51335 ( \51310 , \51308 , \51309 );
buf \U$51336 ( \51311 , \51310 );
buf \U$51337 ( \51312 , \51311 );
nand \U$51338 ( \51313 , \51307 , \51312 );
buf \U$51339 ( \51314 , \51313 );
xor \U$51340 ( \51315 , \51298 , \51314 );
xor \U$51341 ( \51316 , RIc0dacd8_117, RIc0d8b18_45);
buf \U$51342 ( \51317 , \51316 );
not \U$51343 ( \51318 , \51317 );
buf \U$51344 ( \51319 , \22350 );
not \U$51345 ( \51320 , \51319 );
or \U$51346 ( \51321 , \51318 , \51320 );
buf \U$51347 ( \51322 , \22356 );
buf \U$51348 ( \51323 , \50632 );
nand \U$51349 ( \51324 , \51322 , \51323 );
buf \U$51350 ( \51325 , \51324 );
buf \U$51351 ( \51326 , \51325 );
nand \U$51352 ( \51327 , \51321 , \51326 );
buf \U$51353 ( \51328 , \51327 );
and \U$51354 ( \51329 , \51315 , \51328 );
and \U$51355 ( \51330 , \51298 , \51314 );
or \U$51356 ( \51331 , \51329 , \51330 );
buf \U$51357 ( \51332 , \51331 );
and \U$51358 ( \51333 , \51282 , \51332 );
and \U$51359 ( \51334 , \51210 , \51281 );
or \U$51360 ( \51335 , \51333 , \51334 );
buf \U$51361 ( \51336 , \51335 );
buf \U$51362 ( \51337 , \51336 );
xor \U$51363 ( \51338 , \50644 , \50667 );
xor \U$51364 ( \51339 , \51338 , \50627 );
buf \U$51365 ( \51340 , \51339 );
not \U$51366 ( \51341 , \51340 );
buf \U$51367 ( \51342 , \51341 );
not \U$51368 ( \51343 , \51342 );
xor \U$51369 ( \51344 , \50575 , \50589 );
xor \U$51370 ( \51345 , \51344 , \50608 );
buf \U$51371 ( \51346 , \51345 );
not \U$51372 ( \51347 , \51346 );
or \U$51373 ( \51348 , \51343 , \51347 );
buf \U$51374 ( \51349 , \51346 );
not \U$51375 ( \51350 , \51349 );
buf \U$51376 ( \51351 , \51350 );
not \U$51377 ( \51352 , \51351 );
not \U$51378 ( \51353 , \51339 );
or \U$51379 ( \51354 , \51352 , \51353 );
buf \U$51380 ( \51355 , \50528 );
not \U$51381 ( \51356 , \51355 );
buf \U$51382 ( \51357 , \50537 );
not \U$51383 ( \51358 , \51357 );
or \U$51384 ( \51359 , \51356 , \51358 );
not \U$51385 ( \51360 , \50528 );
nand \U$51386 ( \51361 , \51360 , \50514 );
buf \U$51387 ( \51362 , \51361 );
nand \U$51388 ( \51363 , \51359 , \51362 );
buf \U$51389 ( \51364 , \51363 );
buf \U$51390 ( \51365 , \51364 );
buf \U$51391 ( \51366 , \50555 );
xnor \U$51392 ( \51367 , \51365 , \51366 );
buf \U$51393 ( \51368 , \51367 );
buf \U$51394 ( \51369 , \51368 );
not \U$51395 ( \51370 , \51369 );
buf \U$51396 ( \51371 , \51370 );
nand \U$51397 ( \51372 , \51354 , \51371 );
nand \U$51398 ( \51373 , \51348 , \51372 );
buf \U$51399 ( \51374 , \51373 );
xor \U$51400 ( \51375 , \51337 , \51374 );
xor \U$51401 ( \51376 , \50772 , \50845 );
xor \U$51402 ( \51377 , \51376 , \50776 );
buf \U$51403 ( \51378 , \51377 );
and \U$51404 ( \51379 , \51375 , \51378 );
and \U$51405 ( \51380 , \51337 , \51374 );
or \U$51406 ( \51381 , \51379 , \51380 );
buf \U$51407 ( \51382 , \51381 );
buf \U$51408 ( \51383 , \51382 );
xor \U$51409 ( \51384 , \51155 , \51383 );
xor \U$51410 ( \51385 , \50857 , \50900 );
xor \U$51411 ( \51386 , \51385 , \50905 );
buf \U$51412 ( \51387 , \51386 );
buf \U$51413 ( \51388 , \51387 );
and \U$51414 ( \51389 , \51384 , \51388 );
and \U$51415 ( \51390 , \51155 , \51383 );
or \U$51416 ( \51391 , \51389 , \51390 );
buf \U$51417 ( \51392 , \51391 );
buf \U$51418 ( \51393 , \51392 );
and \U$51419 ( \51394 , \51151 , \51393 );
and \U$51420 ( \51395 , \51146 , \51150 );
or \U$51421 ( \51396 , \51394 , \51395 );
buf \U$51422 ( \51397 , \51396 );
buf \U$51423 ( \51398 , \51397 );
xor \U$51424 ( \51399 , \50981 , \51398 );
buf \U$51425 ( \51400 , \50696 );
buf \U$51426 ( \51401 , \50401 );
xor \U$51427 ( \51402 , \51400 , \51401 );
buf \U$51428 ( \51403 , \51402 );
buf \U$51429 ( \51404 , \51403 );
buf \U$51430 ( \51405 , \50948 );
and \U$51431 ( \51406 , \51404 , \51405 );
not \U$51432 ( \51407 , \51404 );
buf \U$51433 ( \51408 , \50948 );
not \U$51434 ( \51409 , \51408 );
buf \U$51435 ( \51410 , \51409 );
buf \U$51436 ( \51411 , \51410 );
and \U$51437 ( \51412 , \51407 , \51411 );
nor \U$51438 ( \51413 , \51406 , \51412 );
buf \U$51439 ( \51414 , \51413 );
buf \U$51440 ( \51415 , \51414 );
and \U$51441 ( \51416 , \51399 , \51415 );
and \U$51442 ( \51417 , \50981 , \51398 );
or \U$51443 ( \51418 , \51416 , \51417 );
buf \U$51444 ( \51419 , \51418 );
buf \U$51445 ( \51420 , \51419 );
not \U$51446 ( \51421 , \51420 );
buf \U$51447 ( \51422 , \50397 );
buf \U$51448 ( \51423 , \50954 );
xor \U$51449 ( \51424 , \51422 , \51423 );
buf \U$51450 ( \51425 , \50959 );
xnor \U$51451 ( \51426 , \51424 , \51425 );
buf \U$51452 ( \51427 , \51426 );
buf \U$51453 ( \51428 , \51427 );
nand \U$51454 ( \51429 , \51421 , \51428 );
buf \U$51455 ( \51430 , \51429 );
buf \U$51456 ( \51431 , \51430 );
and \U$51457 ( \51432 , \50977 , \51431 );
buf \U$51458 ( \51433 , \51432 );
buf \U$51459 ( \51434 , \51433 );
not \U$51460 ( \51435 , \50392 );
buf \U$51461 ( \51436 , \50374 );
not \U$51462 ( \51437 , \51436 );
buf \U$51463 ( \51438 , \49887 );
nand \U$51464 ( \51439 , \51437 , \51438 );
buf \U$51465 ( \51440 , \51439 );
not \U$51466 ( \51441 , \51440 );
or \U$51467 ( \51442 , \51435 , \51441 );
buf \U$51468 ( \51443 , \50374 );
buf \U$51469 ( \51444 , \49884 );
nand \U$51470 ( \51445 , \51443 , \51444 );
buf \U$51471 ( \51446 , \51445 );
nand \U$51472 ( \51447 , \51442 , \51446 );
buf \U$51473 ( \51448 , \51447 );
not \U$51474 ( \51449 , \51448 );
xor \U$51475 ( \51450 , \47540 , \47544 );
xor \U$51476 ( \51451 , \51450 , \47549 );
buf \U$51477 ( \51452 , \51451 );
buf \U$51478 ( \51453 , \51452 );
xor \U$51479 ( \51454 , \50381 , \50385 );
and \U$51480 ( \51455 , \51454 , \50390 );
and \U$51481 ( \51456 , \50381 , \50385 );
or \U$51482 ( \51457 , \51455 , \51456 );
buf \U$51483 ( \51458 , \51457 );
buf \U$51484 ( \51459 , \51458 );
xor \U$51485 ( \51460 , \51453 , \51459 );
xor \U$51486 ( \51461 , \49239 , \49243 );
xor \U$51487 ( \51462 , \51461 , \49330 );
buf \U$51488 ( \51463 , \51462 );
buf \U$51489 ( \51464 , \51463 );
xnor \U$51490 ( \51465 , \51460 , \51464 );
buf \U$51491 ( \51466 , \51465 );
buf \U$51492 ( \51467 , \51466 );
nand \U$51493 ( \51468 , \51449 , \51467 );
buf \U$51494 ( \51469 , \51468 );
buf \U$51495 ( \51470 , \51469 );
buf \U$51496 ( \51471 , \51452 );
buf \U$51497 ( \51472 , \51458 );
or \U$51498 ( \51473 , \51471 , \51472 );
buf \U$51499 ( \51474 , \51463 );
nand \U$51500 ( \51475 , \51473 , \51474 );
buf \U$51501 ( \51476 , \51475 );
buf \U$51502 ( \51477 , \51476 );
buf \U$51503 ( \51478 , \51458 );
buf \U$51504 ( \51479 , \51452 );
nand \U$51505 ( \51480 , \51478 , \51479 );
buf \U$51506 ( \51481 , \51480 );
buf \U$51507 ( \51482 , \51481 );
nand \U$51508 ( \51483 , \51477 , \51482 );
buf \U$51509 ( \51484 , \51483 );
not \U$51510 ( \51485 , \51484 );
xor \U$51511 ( \51486 , \48758 , \49338 );
xor \U$51512 ( \51487 , \51486 , \49364 );
buf \U$51513 ( \51488 , \51487 );
nand \U$51514 ( \51489 , \51485 , \51488 );
buf \U$51515 ( \51490 , \51489 );
nand \U$51516 ( \51491 , \51434 , \51470 , \51490 );
buf \U$51517 ( \51492 , \51491 );
buf \U$51518 ( \51493 , \51492 );
xor \U$51519 ( \51494 , \51155 , \51383 );
xor \U$51520 ( \51495 , \51494 , \51388 );
buf \U$51521 ( \51496 , \51495 );
buf \U$51522 ( \51497 , \51496 );
buf \U$51523 ( \51498 , \16386 );
not \U$51524 ( \51499 , \51498 );
buf \U$51525 ( \51500 , \50502 );
not \U$51526 ( \51501 , \51500 );
or \U$51527 ( \51502 , \51499 , \51501 );
buf \U$51528 ( \51503 , \12968 );
buf \U$51529 ( \51504 , RIc0daeb8_121);
buf \U$51530 ( \51505 , RIc0d8938_41);
xnor \U$51531 ( \51506 , \51504 , \51505 );
buf \U$51532 ( \51507 , \51506 );
buf \U$51533 ( \51508 , \51507 );
or \U$51534 ( \51509 , \51503 , \51508 );
nand \U$51535 ( \51510 , \51502 , \51509 );
buf \U$51536 ( \51511 , \51510 );
buf \U$51537 ( \51512 , \51511 );
buf \U$51538 ( \51513 , \14405 );
buf \U$51539 ( \51514 , \12396 );
buf \U$51540 ( \51515 , RIc0d8d70_50);
buf \U$51541 ( \51516 , RIc0daaf8_113);
xor \U$51542 ( \51517 , \51515 , \51516 );
buf \U$51543 ( \51518 , \51517 );
buf \U$51544 ( \51519 , \51518 );
nand \U$51545 ( \51520 , \51514 , \51519 );
buf \U$51546 ( \51521 , \51520 );
buf \U$51547 ( \51522 , \51521 );
nor \U$51548 ( \51523 , \51513 , \51522 );
buf \U$51549 ( \51524 , \51523 );
buf \U$51550 ( \51525 , \51524 );
not \U$51551 ( \51526 , \51525 );
buf \U$51552 ( \51527 , \12410 );
buf \U$51553 ( \51528 , \51176 );
nand \U$51554 ( \51529 , \51527 , \51528 );
buf \U$51555 ( \51530 , \51529 );
buf \U$51556 ( \51531 , \51530 );
nand \U$51557 ( \51532 , \51526 , \51531 );
buf \U$51558 ( \51533 , \51532 );
buf \U$51559 ( \51534 , \51533 );
buf \U$51560 ( \51535 , RIc0d86e0_36);
buf \U$51561 ( \51536 , RIc0db188_127);
xor \U$51562 ( \51537 , \51535 , \51536 );
buf \U$51563 ( \51538 , \51537 );
buf \U$51564 ( \51539 , \51538 );
not \U$51565 ( \51540 , \51539 );
buf \U$51566 ( \51541 , \15609 );
not \U$51567 ( \51542 , \51541 );
or \U$51568 ( \51543 , \51540 , \51542 );
buf \U$51569 ( \51544 , \51159 );
buf \U$51570 ( \51545 , RIc0db200_128);
nand \U$51571 ( \51546 , \51544 , \51545 );
buf \U$51572 ( \51547 , \51546 );
buf \U$51573 ( \51548 , \51547 );
nand \U$51574 ( \51549 , \51543 , \51548 );
buf \U$51575 ( \51550 , \51549 );
buf \U$51576 ( \51551 , \51550 );
or \U$51577 ( \51552 , \51534 , \51551 );
xor \U$51578 ( \51553 , RIc0db098_125, RIc0d87d0_38);
buf \U$51579 ( \51554 , \51553 );
not \U$51580 ( \51555 , \51554 );
buf \U$51581 ( \51556 , \13461 );
not \U$51582 ( \51557 , \51556 );
or \U$51583 ( \51558 , \51555 , \51557 );
buf \U$51584 ( \51559 , \13465 );
buf \U$51585 ( \51560 , \51090 );
nand \U$51586 ( \51561 , \51559 , \51560 );
buf \U$51587 ( \51562 , \51561 );
buf \U$51588 ( \51563 , \51562 );
nand \U$51589 ( \51564 , \51558 , \51563 );
buf \U$51590 ( \51565 , \51564 );
buf \U$51591 ( \51566 , \51565 );
nand \U$51592 ( \51567 , \51552 , \51566 );
buf \U$51593 ( \51568 , \51567 );
buf \U$51594 ( \51569 , \51568 );
buf \U$51595 ( \51570 , \51550 );
buf \U$51596 ( \51571 , \51533 );
nand \U$51597 ( \51572 , \51570 , \51571 );
buf \U$51598 ( \51573 , \51572 );
buf \U$51599 ( \51574 , \51573 );
nand \U$51600 ( \51575 , \51569 , \51574 );
buf \U$51601 ( \51576 , \51575 );
buf \U$51602 ( \51577 , \51576 );
xor \U$51603 ( \51578 , \51512 , \51577 );
buf \U$51604 ( \51579 , RIc0d9310_62);
buf \U$51605 ( \51580 , RIc0da558_101);
xor \U$51606 ( \51581 , \51579 , \51580 );
buf \U$51607 ( \51582 , \51581 );
buf \U$51608 ( \51583 , \51582 );
not \U$51609 ( \51584 , \51583 );
buf \U$51610 ( \51585 , \3535 );
not \U$51611 ( \51586 , \51585 );
or \U$51612 ( \51587 , \51584 , \51586 );
buf \U$51613 ( \51588 , \4049 );
buf \U$51614 ( \51589 , \51075 );
nand \U$51615 ( \51590 , \51588 , \51589 );
buf \U$51616 ( \51591 , \51590 );
buf \U$51617 ( \51592 , \51591 );
nand \U$51618 ( \51593 , \51587 , \51592 );
buf \U$51619 ( \51594 , \51593 );
buf \U$51620 ( \51595 , \51594 );
not \U$51621 ( \51596 , \51595 );
buf \U$51622 ( \51597 , RIc0d9400_64);
buf \U$51623 ( \51598 , RIc0da4e0_100);
or \U$51624 ( \51599 , \51597 , \51598 );
buf \U$51625 ( \51600 , RIc0da558_101);
nand \U$51626 ( \51601 , \51599 , \51600 );
buf \U$51627 ( \51602 , \51601 );
buf \U$51628 ( \51603 , \51602 );
buf \U$51629 ( \51604 , RIc0d9400_64);
buf \U$51630 ( \51605 , RIc0da4e0_100);
nand \U$51631 ( \51606 , \51604 , \51605 );
buf \U$51632 ( \51607 , \51606 );
buf \U$51633 ( \51608 , \51607 );
buf \U$51634 ( \51609 , RIc0da468_99);
nand \U$51635 ( \51610 , \51603 , \51608 , \51609 );
buf \U$51636 ( \51611 , \51610 );
buf \U$51637 ( \51612 , \51611 );
nor \U$51638 ( \51613 , \51596 , \51612 );
buf \U$51639 ( \51614 , \51613 );
buf \U$51640 ( \51615 , \51614 );
and \U$51641 ( \51616 , \51578 , \51615 );
and \U$51642 ( \51617 , \51512 , \51577 );
or \U$51643 ( \51618 , \51616 , \51617 );
buf \U$51644 ( \51619 , \51618 );
buf \U$51645 ( \51620 , \51619 );
not \U$51646 ( \51621 , \51620 );
xor \U$51647 ( \51622 , \50739 , \50763 );
xnor \U$51648 ( \51623 , \51622 , \50722 );
buf \U$51649 ( \51624 , \51623 );
not \U$51650 ( \51625 , \51624 );
or \U$51651 ( \51626 , \51621 , \51625 );
buf \U$51652 ( \51627 , \51623 );
buf \U$51653 ( \51628 , \51619 );
or \U$51654 ( \51629 , \51627 , \51628 );
buf \U$51655 ( \51630 , \50834 );
not \U$51656 ( \51631 , \51630 );
buf \U$51657 ( \51632 , \50815 );
not \U$51658 ( \51633 , \51632 );
or \U$51659 ( \51634 , \51631 , \51633 );
buf \U$51660 ( \51635 , \50815 );
buf \U$51661 ( \51636 , \50834 );
or \U$51662 ( \51637 , \51635 , \51636 );
nand \U$51663 ( \51638 , \51634 , \51637 );
buf \U$51664 ( \51639 , \51638 );
buf \U$51665 ( \51640 , \51639 );
buf \U$51666 ( \51641 , \50791 );
and \U$51667 ( \51642 , \51640 , \51641 );
not \U$51668 ( \51643 , \51640 );
buf \U$51669 ( \51644 , \50794 );
and \U$51670 ( \51645 , \51643 , \51644 );
nor \U$51671 ( \51646 , \51642 , \51645 );
buf \U$51672 ( \51647 , \51646 );
buf \U$51673 ( \51648 , \51647 );
nand \U$51674 ( \51649 , \51629 , \51648 );
buf \U$51675 ( \51650 , \51649 );
buf \U$51676 ( \51651 , \51650 );
nand \U$51677 ( \51652 , \51626 , \51651 );
buf \U$51678 ( \51653 , \51652 );
buf \U$51679 ( \51654 , \51653 );
xor \U$51680 ( \51655 , \50558 , \50613 );
xor \U$51681 ( \51656 , \51655 , \50677 );
buf \U$51682 ( \51657 , \51656 );
buf \U$51683 ( \51658 , \51657 );
xor \U$51684 ( \51659 , \51654 , \51658 );
xor \U$51685 ( \51660 , \50860 , \50888 );
xor \U$51686 ( \51661 , \51660 , \50884 );
buf \U$51687 ( \51662 , \51661 );
and \U$51688 ( \51663 , \51659 , \51662 );
and \U$51689 ( \51664 , \51654 , \51658 );
or \U$51690 ( \51665 , \51663 , \51664 );
buf \U$51691 ( \51666 , \51665 );
buf \U$51692 ( \51667 , \51666 );
xor \U$51693 ( \51668 , \50985 , \51121 );
xor \U$51694 ( \51669 , \51668 , \51141 );
buf \U$51695 ( \51670 , \51669 );
buf \U$51696 ( \51671 , \51670 );
xor \U$51697 ( \51672 , \51667 , \51671 );
xor \U$51698 ( \51673 , \50989 , \50993 );
xor \U$51699 ( \51674 , \51673 , \51116 );
buf \U$51700 ( \51675 , \51674 );
buf \U$51701 ( \51676 , \51675 );
xor \U$51702 ( \51677 , \50997 , \51068 );
xor \U$51703 ( \51678 , \51677 , \51111 );
buf \U$51704 ( \51679 , \51678 );
buf \U$51705 ( \51680 , \51679 );
xor \U$51706 ( \51681 , \51210 , \51281 );
xor \U$51707 ( \51682 , \51681 , \51332 );
buf \U$51708 ( \51683 , \51682 );
buf \U$51709 ( \51684 , \51683 );
or \U$51710 ( \51685 , \51680 , \51684 );
xor \U$51711 ( \51686 , RIc0daa08_111, RIc0d8e60_52);
buf \U$51712 ( \51687 , \51686 );
not \U$51713 ( \51688 , \51687 );
buf \U$51714 ( \51689 , \12529 );
not \U$51715 ( \51690 , \51689 );
or \U$51716 ( \51691 , \51688 , \51690 );
buf \U$51717 ( \51692 , \14106 );
buf \U$51718 ( \51693 , \51302 );
nand \U$51719 ( \51694 , \51692 , \51693 );
buf \U$51720 ( \51695 , \51694 );
buf \U$51721 ( \51696 , \51695 );
nand \U$51722 ( \51697 , \51691 , \51696 );
buf \U$51723 ( \51698 , \51697 );
buf \U$51724 ( \51699 , \51698 );
buf \U$51725 ( \51700 , RIc0d9130_58);
buf \U$51726 ( \51701 , RIc0da738_105);
xor \U$51727 ( \51702 , \51700 , \51701 );
buf \U$51728 ( \51703 , \51702 );
buf \U$51729 ( \51704 , \51703 );
not \U$51730 ( \51705 , \51704 );
buf \U$51731 ( \51706 , \12736 );
not \U$51732 ( \51707 , \51706 );
or \U$51733 ( \51708 , \51705 , \51707 );
buf \U$51734 ( \51709 , \21880 );
buf \U$51735 ( \51710 , \51214 );
nand \U$51736 ( \51711 , \51709 , \51710 );
buf \U$51737 ( \51712 , \51711 );
buf \U$51738 ( \51713 , \51712 );
nand \U$51739 ( \51714 , \51708 , \51713 );
buf \U$51740 ( \51715 , \51714 );
buf \U$51741 ( \51716 , \51715 );
xor \U$51742 ( \51717 , \51699 , \51716 );
buf \U$51743 ( \51718 , \14207 );
buf \U$51744 ( \51719 , RIc0da918_109);
buf \U$51745 ( \51720 , RIc0d8f50_54);
xnor \U$51746 ( \51721 , \51719 , \51720 );
buf \U$51747 ( \51722 , \51721 );
buf \U$51748 ( \51723 , \51722 );
or \U$51749 ( \51724 , \51718 , \51723 );
buf \U$51750 ( \51725 , \36203 );
buf \U$51751 ( \51726 , \51286 );
not \U$51752 ( \51727 , \51726 );
buf \U$51753 ( \51728 , \51727 );
buf \U$51754 ( \51729 , \51728 );
or \U$51755 ( \51730 , \51725 , \51729 );
nand \U$51756 ( \51731 , \51724 , \51730 );
buf \U$51757 ( \51732 , \51731 );
buf \U$51758 ( \51733 , \51732 );
and \U$51759 ( \51734 , \51717 , \51733 );
and \U$51760 ( \51735 , \51699 , \51716 );
or \U$51761 ( \51736 , \51734 , \51735 );
buf \U$51762 ( \51737 , \51736 );
buf \U$51763 ( \51738 , \51737 );
buf \U$51764 ( \51739 , RIc0dacd8_117);
buf \U$51765 ( \51740 , RIc0d8b90_46);
xor \U$51766 ( \51741 , \51739 , \51740 );
buf \U$51767 ( \51742 , \51741 );
buf \U$51768 ( \51743 , \51742 );
not \U$51769 ( \51744 , \51743 );
buf \U$51770 ( \51745 , \22350 );
not \U$51771 ( \51746 , \51745 );
or \U$51772 ( \51747 , \51744 , \51746 );
buf \U$51773 ( \51748 , \16559 );
buf \U$51774 ( \51749 , \51316 );
nand \U$51775 ( \51750 , \51748 , \51749 );
buf \U$51776 ( \51751 , \51750 );
buf \U$51777 ( \51752 , \51751 );
nand \U$51778 ( \51753 , \51747 , \51752 );
buf \U$51779 ( \51754 , \51753 );
buf \U$51780 ( \51755 , \51754 );
xor \U$51781 ( \51756 , RIc0dadc8_119, RIc0d8aa0_44);
buf \U$51782 ( \51757 , \51756 );
not \U$51783 ( \51758 , \51757 );
buf \U$51784 ( \51759 , \14569 );
not \U$51785 ( \51760 , \51759 );
or \U$51786 ( \51761 , \51758 , \51760 );
buf \U$51787 ( \51762 , \13953 );
buf \U$51788 ( \51763 , \51001 );
nand \U$51789 ( \51764 , \51762 , \51763 );
buf \U$51790 ( \51765 , \51764 );
buf \U$51791 ( \51766 , \51765 );
nand \U$51792 ( \51767 , \51761 , \51766 );
buf \U$51793 ( \51768 , \51767 );
buf \U$51794 ( \51769 , \51768 );
xor \U$51795 ( \51770 , \51755 , \51769 );
xor \U$51796 ( \51771 , RIc0da648_103, RIc0d9220_60);
buf \U$51797 ( \51772 , \51771 );
not \U$51798 ( \51773 , \51772 );
buf \U$51799 ( \51774 , \16578 );
not \U$51800 ( \51775 , \51774 );
or \U$51801 ( \51776 , \51773 , \51775 );
buf \U$51802 ( \51777 , \13712 );
buf \U$51803 ( \51778 , \51044 );
nand \U$51804 ( \51779 , \51777 , \51778 );
buf \U$51805 ( \51780 , \51779 );
buf \U$51806 ( \51781 , \51780 );
nand \U$51807 ( \51782 , \51776 , \51781 );
buf \U$51808 ( \51783 , \51782 );
buf \U$51809 ( \51784 , \51783 );
and \U$51810 ( \51785 , \51770 , \51784 );
and \U$51811 ( \51786 , \51755 , \51769 );
or \U$51812 ( \51787 , \51785 , \51786 );
buf \U$51813 ( \51788 , \51787 );
buf \U$51814 ( \51789 , \51788 );
xor \U$51815 ( \51790 , \51738 , \51789 );
buf \U$51816 ( \51791 , RIc0d8c80_48);
buf \U$51817 ( \51792 , RIc0dabe8_115);
xor \U$51818 ( \51793 , \51791 , \51792 );
buf \U$51819 ( \51794 , \51793 );
buf \U$51820 ( \51795 , \51794 );
not \U$51821 ( \51796 , \51795 );
buf \U$51822 ( \51797 , \14186 );
not \U$51823 ( \51798 , \51797 );
or \U$51824 ( \51799 , \51796 , \51798 );
buf \U$51825 ( \51800 , \12303 );
buf \U$51826 ( \51801 , \51257 );
nand \U$51827 ( \51802 , \51800 , \51801 );
buf \U$51828 ( \51803 , \51802 );
buf \U$51829 ( \51804 , \51803 );
nand \U$51830 ( \51805 , \51799 , \51804 );
buf \U$51831 ( \51806 , \51805 );
buf \U$51832 ( \51807 , \51806 );
buf \U$51833 ( \51808 , RIc0d9400_64);
buf \U$51834 ( \51809 , RIc0da468_99);
xor \U$51835 ( \51810 , \51808 , \51809 );
buf \U$51836 ( \51811 , \51810 );
buf \U$51837 ( \51812 , \51811 );
not \U$51838 ( \51813 , \51812 );
buf \U$51839 ( \51814 , \2470 );
not \U$51840 ( \51815 , \51814 );
or \U$51841 ( \51816 , \51813 , \51815 );
buf \U$51842 ( \51817 , \14648 );
buf \U$51843 ( \51818 , \51235 );
nand \U$51844 ( \51819 , \51817 , \51818 );
buf \U$51845 ( \51820 , \51819 );
buf \U$51846 ( \51821 , \51820 );
nand \U$51847 ( \51822 , \51816 , \51821 );
buf \U$51848 ( \51823 , \51822 );
buf \U$51849 ( \51824 , \51823 );
xor \U$51850 ( \51825 , \51807 , \51824 );
buf \U$51851 ( \51826 , RIc0dafa8_123);
buf \U$51852 ( \51827 , RIc0d88c0_40);
xor \U$51853 ( \51828 , \51826 , \51827 );
buf \U$51854 ( \51829 , \51828 );
buf \U$51855 ( \51830 , \51829 );
not \U$51856 ( \51831 , \51830 );
buf \U$51857 ( \51832 , \14982 );
not \U$51858 ( \51833 , \51832 );
or \U$51859 ( \51834 , \51831 , \51833 );
buf \U$51860 ( \51835 , \51200 );
not \U$51861 ( \51836 , \51835 );
buf \U$51862 ( \51837 , \14278 );
nand \U$51863 ( \51838 , \51836 , \51837 );
buf \U$51864 ( \51839 , \51838 );
buf \U$51865 ( \51840 , \51839 );
nand \U$51866 ( \51841 , \51834 , \51840 );
buf \U$51867 ( \51842 , \51841 );
buf \U$51868 ( \51843 , \51842 );
and \U$51869 ( \51844 , \51825 , \51843 );
and \U$51870 ( \51845 , \51807 , \51824 );
or \U$51871 ( \51846 , \51844 , \51845 );
buf \U$51872 ( \51847 , \51846 );
buf \U$51873 ( \51848 , \51847 );
and \U$51874 ( \51849 , \51790 , \51848 );
and \U$51875 ( \51850 , \51738 , \51789 );
or \U$51876 ( \51851 , \51849 , \51850 );
buf \U$51877 ( \51852 , \51851 );
buf \U$51878 ( \51853 , \51852 );
nand \U$51879 ( \51854 , \51685 , \51853 );
buf \U$51880 ( \51855 , \51854 );
buf \U$51881 ( \51856 , \51855 );
buf \U$51882 ( \51857 , \51679 );
buf \U$51883 ( \51858 , \51683 );
nand \U$51884 ( \51859 , \51857 , \51858 );
buf \U$51885 ( \51860 , \51859 );
buf \U$51886 ( \51861 , \51860 );
nand \U$51887 ( \51862 , \51856 , \51861 );
buf \U$51888 ( \51863 , \51862 );
buf \U$51889 ( \51864 , \51863 );
xor \U$51890 ( \51865 , \51676 , \51864 );
xor \U$51891 ( \51866 , \51172 , \51189 );
xor \U$51892 ( \51867 , \51866 , \51205 );
buf \U$51893 ( \51868 , \51867 );
buf \U$51894 ( \51869 , \51868 );
buf \U$51895 ( \51870 , \51229 );
not \U$51896 ( \51871 , \51870 );
buf \U$51897 ( \51872 , \51250 );
not \U$51898 ( \51873 , \51872 );
buf \U$51899 ( \51874 , \51269 );
not \U$51900 ( \51875 , \51874 );
or \U$51901 ( \51876 , \51873 , \51875 );
buf \U$51902 ( \51877 , \51269 );
buf \U$51903 ( \51878 , \51250 );
or \U$51904 ( \51879 , \51877 , \51878 );
nand \U$51905 ( \51880 , \51876 , \51879 );
buf \U$51906 ( \51881 , \51880 );
buf \U$51907 ( \51882 , \51881 );
not \U$51908 ( \51883 , \51882 );
or \U$51909 ( \51884 , \51871 , \51883 );
buf \U$51910 ( \51885 , \51881 );
buf \U$51911 ( \51886 , \51229 );
or \U$51912 ( \51887 , \51885 , \51886 );
nand \U$51913 ( \51888 , \51884 , \51887 );
buf \U$51914 ( \51889 , \51888 );
buf \U$51915 ( \51890 , \51889 );
xor \U$51916 ( \51891 , \51869 , \51890 );
and \U$51917 ( \51892 , RIc0daeb8_121, \45192 );
not \U$51918 ( \51893 , RIc0daeb8_121);
and \U$51919 ( \51894 , \51893 , RIc0d89b0_42);
or \U$51920 ( \51895 , \51892 , \51894 );
buf \U$51921 ( \51896 , \51895 );
not \U$51922 ( \51897 , \51896 );
buf \U$51923 ( \51898 , \19487 );
not \U$51924 ( \51899 , \51898 );
or \U$51925 ( \51900 , \51897 , \51899 );
buf \U$51926 ( \51901 , \51507 );
not \U$51927 ( \51902 , \51901 );
buf \U$51928 ( \51903 , \13314 );
nand \U$51929 ( \51904 , \51902 , \51903 );
buf \U$51930 ( \51905 , \51904 );
buf \U$51931 ( \51906 , \51905 );
nand \U$51932 ( \51907 , \51900 , \51906 );
buf \U$51933 ( \51908 , \51907 );
buf \U$51934 ( \51909 , \51908 );
not \U$51935 ( \51910 , \51909 );
buf \U$51936 ( \51911 , RIc0da828_107);
buf \U$51937 ( \51912 , RIc0d9040_56);
xnor \U$51938 ( \51913 , \51911 , \51912 );
buf \U$51939 ( \51914 , \51913 );
buf \U$51940 ( \51915 , \51914 );
not \U$51941 ( \51916 , \51915 );
buf \U$51942 ( \51917 , \51916 );
buf \U$51943 ( \51918 , \51917 );
not \U$51944 ( \51919 , \51918 );
buf \U$51945 ( \51920 , \21898 );
not \U$51946 ( \51921 , \51920 );
or \U$51947 ( \51922 , \51919 , \51921 );
buf \U$51948 ( \51923 , \16071 );
buf \U$51949 ( \51924 , \51022 );
nand \U$51950 ( \51925 , \51923 , \51924 );
buf \U$51951 ( \51926 , \51925 );
buf \U$51952 ( \51927 , \51926 );
nand \U$51953 ( \51928 , \51922 , \51927 );
buf \U$51954 ( \51929 , \51928 );
buf \U$51955 ( \51930 , \51929 );
not \U$51956 ( \51931 , \51930 );
or \U$51957 ( \51932 , \51910 , \51931 );
xor \U$51958 ( \51933 , \51594 , \51611 );
buf \U$51959 ( \51934 , \51933 );
not \U$51960 ( \51935 , \51934 );
buf \U$51961 ( \51936 , \51908 );
not \U$51962 ( \51937 , \51936 );
buf \U$51963 ( \51938 , \51929 );
not \U$51964 ( \51939 , \51938 );
buf \U$51965 ( \51940 , \51939 );
buf \U$51966 ( \51941 , \51940 );
nand \U$51967 ( \51942 , \51937 , \51941 );
buf \U$51968 ( \51943 , \51942 );
buf \U$51969 ( \51944 , \51943 );
nand \U$51970 ( \51945 , \51935 , \51944 );
buf \U$51971 ( \51946 , \51945 );
buf \U$51972 ( \51947 , \51946 );
nand \U$51973 ( \51948 , \51932 , \51947 );
buf \U$51974 ( \51949 , \51948 );
buf \U$51975 ( \51950 , \51949 );
and \U$51976 ( \51951 , \51891 , \51950 );
and \U$51977 ( \51952 , \51869 , \51890 );
or \U$51978 ( \51953 , \51951 , \51952 );
buf \U$51979 ( \51954 , \51953 );
buf \U$51980 ( \51955 , \51954 );
not \U$51981 ( \51956 , \51955 );
buf \U$51982 ( \51957 , \51351 );
not \U$51983 ( \51958 , \51957 );
buf \U$51984 ( \51959 , \51371 );
not \U$51985 ( \51960 , \51959 );
or \U$51986 ( \51961 , \51958 , \51960 );
buf \U$51987 ( \51962 , \51368 );
buf \U$51988 ( \51963 , \51346 );
nand \U$51989 ( \51964 , \51962 , \51963 );
buf \U$51990 ( \51965 , \51964 );
buf \U$51991 ( \51966 , \51965 );
nand \U$51992 ( \51967 , \51961 , \51966 );
buf \U$51993 ( \51968 , \51967 );
buf \U$51994 ( \51969 , \51968 );
buf \U$51995 ( \51970 , \51342 );
and \U$51996 ( \51971 , \51969 , \51970 );
not \U$51997 ( \51972 , \51969 );
buf \U$51998 ( \51973 , \51339 );
and \U$51999 ( \51974 , \51972 , \51973 );
nor \U$52000 ( \51975 , \51971 , \51974 );
buf \U$52001 ( \51976 , \51975 );
buf \U$52002 ( \51977 , \51976 );
not \U$52003 ( \51978 , \51977 );
or \U$52004 ( \51979 , \51956 , \51978 );
buf \U$52005 ( \51980 , \51976 );
buf \U$52006 ( \51981 , \51954 );
or \U$52007 ( \51982 , \51980 , \51981 );
buf \U$52008 ( \51983 , \51013 );
not \U$52009 ( \51984 , \51983 );
buf \U$52010 ( \51985 , \51037 );
not \U$52011 ( \51986 , \51985 );
or \U$52012 ( \51987 , \51984 , \51986 );
buf \U$52013 ( \51988 , \51034 );
buf \U$52014 ( \51989 , \51016 );
nand \U$52015 ( \51990 , \51988 , \51989 );
buf \U$52016 ( \51991 , \51990 );
buf \U$52017 ( \51992 , \51991 );
nand \U$52018 ( \51993 , \51987 , \51992 );
buf \U$52019 ( \51994 , \51993 );
buf \U$52020 ( \51995 , \51994 );
buf \U$52021 ( \51996 , \51056 );
xor \U$52022 ( \51997 , \51995 , \51996 );
buf \U$52023 ( \51998 , \51997 );
buf \U$52024 ( \51999 , \51998 );
xor \U$52025 ( \52000 , \51074 , \51088 );
xor \U$52026 ( \52001 , \52000 , \51106 );
buf \U$52027 ( \52002 , \52001 );
buf \U$52028 ( \52003 , \52002 );
xor \U$52029 ( \52004 , \51999 , \52003 );
xor \U$52030 ( \52005 , \51298 , \51314 );
xor \U$52031 ( \52006 , \52005 , \51328 );
buf \U$52032 ( \52007 , \52006 );
and \U$52033 ( \52008 , \52004 , \52007 );
and \U$52034 ( \52009 , \51999 , \52003 );
or \U$52035 ( \52010 , \52008 , \52009 );
buf \U$52036 ( \52011 , \52010 );
buf \U$52037 ( \52012 , \52011 );
nand \U$52038 ( \52013 , \51982 , \52012 );
buf \U$52039 ( \52014 , \52013 );
buf \U$52040 ( \52015 , \52014 );
nand \U$52041 ( \52016 , \51979 , \52015 );
buf \U$52042 ( \52017 , \52016 );
buf \U$52043 ( \52018 , \52017 );
and \U$52044 ( \52019 , \51865 , \52018 );
and \U$52045 ( \52020 , \51676 , \51864 );
or \U$52046 ( \52021 , \52019 , \52020 );
buf \U$52047 ( \52022 , \52021 );
buf \U$52048 ( \52023 , \52022 );
xor \U$52049 ( \52024 , \51672 , \52023 );
buf \U$52050 ( \52025 , \52024 );
buf \U$52051 ( \52026 , \52025 );
xor \U$52052 ( \52027 , \51497 , \52026 );
xor \U$52053 ( \52028 , \51654 , \51658 );
xor \U$52054 ( \52029 , \52028 , \51662 );
buf \U$52055 ( \52030 , \52029 );
buf \U$52056 ( \52031 , \52030 );
xor \U$52057 ( \52032 , \51337 , \51374 );
xor \U$52058 ( \52033 , \52032 , \51378 );
buf \U$52059 ( \52034 , \52033 );
buf \U$52060 ( \52035 , \52034 );
xor \U$52061 ( \52036 , \52031 , \52035 );
xor \U$52062 ( \52037 , \51676 , \51864 );
xor \U$52063 ( \52038 , \52037 , \52018 );
buf \U$52064 ( \52039 , \52038 );
buf \U$52065 ( \52040 , \52039 );
and \U$52066 ( \52041 , \52036 , \52040 );
and \U$52067 ( \52042 , \52031 , \52035 );
or \U$52068 ( \52043 , \52041 , \52042 );
buf \U$52069 ( \52044 , \52043 );
buf \U$52070 ( \52045 , \52044 );
xor \U$52071 ( \52046 , \52027 , \52045 );
buf \U$52072 ( \52047 , \52046 );
buf \U$52073 ( \52048 , \52047 );
xor \U$52074 ( \52049 , \51647 , \51623 );
xor \U$52075 ( \52050 , \52049 , \51619 );
buf \U$52076 ( \52051 , \52050 );
xor \U$52077 ( \52052 , \51512 , \51577 );
xor \U$52078 ( \52053 , \52052 , \51615 );
buf \U$52079 ( \52054 , \52053 );
buf \U$52080 ( \52055 , \52054 );
buf \U$52081 ( \52056 , \51703 );
not \U$52082 ( \52057 , \52056 );
buf \U$52083 ( \52058 , \12744 );
not \U$52084 ( \52059 , \52058 );
or \U$52085 ( \52060 , \52057 , \52059 );
buf \U$52086 ( \52061 , \40782 );
buf \U$52087 ( \52062 , RIc0d91a8_59);
buf \U$52088 ( \52063 , RIc0da738_105);
xor \U$52089 ( \52064 , \52062 , \52063 );
buf \U$52090 ( \52065 , \52064 );
buf \U$52091 ( \52066 , \52065 );
buf \U$52092 ( \52067 , \12731 );
nand \U$52093 ( \52068 , \52061 , \52066 , \52067 );
buf \U$52094 ( \52069 , \52068 );
buf \U$52095 ( \52070 , \52069 );
nand \U$52096 ( \52071 , \52060 , \52070 );
buf \U$52097 ( \52072 , \52071 );
buf \U$52098 ( \52073 , \52072 );
buf \U$52099 ( \52074 , \51895 );
not \U$52100 ( \52075 , \52074 );
buf \U$52101 ( \52076 , \12975 );
not \U$52102 ( \52077 , \52076 );
or \U$52103 ( \52078 , \52075 , \52077 );
buf \U$52104 ( \52079 , \12975 );
not \U$52105 ( \52080 , \52079 );
buf \U$52106 ( \52081 , \52080 );
buf \U$52107 ( \52082 , \52081 );
xor \U$52108 ( \52083 , RIc0daeb8_121, RIc0d8a28_43);
buf \U$52109 ( \52084 , \52083 );
buf \U$52110 ( \52085 , \12964 );
nand \U$52111 ( \52086 , \52082 , \52084 , \52085 );
buf \U$52112 ( \52087 , \52086 );
buf \U$52113 ( \52088 , \52087 );
nand \U$52114 ( \52089 , \52078 , \52088 );
buf \U$52115 ( \52090 , \52089 );
buf \U$52116 ( \52091 , \52090 );
xor \U$52117 ( \52092 , \52073 , \52091 );
buf \U$52118 ( \52093 , \14207 );
xor \U$52119 ( \52094 , RIc0da918_109, RIc0d8fc8_55);
buf \U$52120 ( \52095 , \52094 );
not \U$52121 ( \52096 , \52095 );
buf \U$52122 ( \52097 , \52096 );
buf \U$52123 ( \52098 , \52097 );
or \U$52124 ( \52099 , \52093 , \52098 );
buf \U$52125 ( \52100 , \13423 );
buf \U$52126 ( \52101 , \51722 );
or \U$52127 ( \52102 , \52100 , \52101 );
nand \U$52128 ( \52103 , \52099 , \52102 );
buf \U$52129 ( \52104 , \52103 );
buf \U$52130 ( \52105 , \52104 );
and \U$52131 ( \52106 , \52092 , \52105 );
and \U$52132 ( \52107 , \52073 , \52091 );
or \U$52133 ( \52108 , \52106 , \52107 );
buf \U$52134 ( \52109 , \52108 );
buf \U$52135 ( \52110 , \52109 );
not \U$52136 ( \52111 , \52110 );
buf \U$52137 ( \52112 , \51533 );
buf \U$52138 ( \52113 , \51550 );
xor \U$52139 ( \52114 , \52112 , \52113 );
buf \U$52140 ( \52115 , \51565 );
xor \U$52141 ( \52116 , \52114 , \52115 );
buf \U$52142 ( \52117 , \52116 );
buf \U$52143 ( \52118 , \52117 );
not \U$52144 ( \52119 , \52118 );
or \U$52145 ( \52120 , \52111 , \52119 );
buf \U$52146 ( \52121 , \52117 );
buf \U$52147 ( \52122 , \52109 );
or \U$52148 ( \52123 , \52121 , \52122 );
buf \U$52149 ( \52124 , RIc0d8758_37);
buf \U$52150 ( \52125 , RIc0db188_127);
xor \U$52151 ( \52126 , \52124 , \52125 );
buf \U$52152 ( \52127 , \52126 );
buf \U$52153 ( \52128 , \52127 );
not \U$52154 ( \52129 , \52128 );
buf \U$52155 ( \52130 , \43780 );
not \U$52156 ( \52131 , \52130 );
or \U$52157 ( \52132 , \52129 , \52131 );
buf \U$52158 ( \52133 , \51538 );
buf \U$52159 ( \52134 , RIc0db200_128);
nand \U$52160 ( \52135 , \52133 , \52134 );
buf \U$52161 ( \52136 , \52135 );
buf \U$52162 ( \52137 , \52136 );
nand \U$52163 ( \52138 , \52132 , \52137 );
buf \U$52164 ( \52139 , \52138 );
buf \U$52165 ( \52140 , \52139 );
not \U$52166 ( \52141 , \52140 );
buf \U$52167 ( \52142 , RIc0dafa8_123);
buf \U$52168 ( \52143 , RIc0d8938_41);
xor \U$52169 ( \52144 , \52142 , \52143 );
buf \U$52170 ( \52145 , \52144 );
buf \U$52171 ( \52146 , \52145 );
not \U$52172 ( \52147 , \52146 );
buf \U$52173 ( \52148 , \14982 );
not \U$52174 ( \52149 , \52148 );
or \U$52175 ( \52150 , \52147 , \52149 );
buf \U$52176 ( \52151 , \16692 );
buf \U$52177 ( \52152 , \51829 );
nand \U$52178 ( \52153 , \52151 , \52152 );
buf \U$52179 ( \52154 , \52153 );
buf \U$52180 ( \52155 , \52154 );
nand \U$52181 ( \52156 , \52150 , \52155 );
buf \U$52182 ( \52157 , \52156 );
buf \U$52183 ( \52158 , \52157 );
not \U$52184 ( \52159 , \52158 );
or \U$52185 ( \52160 , \52141 , \52159 );
buf \U$52186 ( \52161 , \52157 );
buf \U$52187 ( \52162 , \52139 );
or \U$52188 ( \52163 , \52161 , \52162 );
buf \U$52189 ( \52164 , RIc0d8848_39);
buf \U$52190 ( \52165 , RIc0db098_125);
xor \U$52191 ( \52166 , \52164 , \52165 );
buf \U$52192 ( \52167 , \52166 );
buf \U$52193 ( \52168 , \52167 );
not \U$52194 ( \52169 , \52168 );
buf \U$52195 ( \52170 , \15789 );
not \U$52196 ( \52171 , \52170 );
or \U$52197 ( \52172 , \52169 , \52171 );
buf \U$52198 ( \52173 , \15793 );
buf \U$52199 ( \52174 , \51553 );
nand \U$52200 ( \52175 , \52173 , \52174 );
buf \U$52201 ( \52176 , \52175 );
buf \U$52202 ( \52177 , \52176 );
nand \U$52203 ( \52178 , \52172 , \52177 );
buf \U$52204 ( \52179 , \52178 );
buf \U$52205 ( \52180 , \52179 );
nand \U$52206 ( \52181 , \52163 , \52180 );
buf \U$52207 ( \52182 , \52181 );
buf \U$52208 ( \52183 , \52182 );
nand \U$52209 ( \52184 , \52160 , \52183 );
buf \U$52210 ( \52185 , \52184 );
buf \U$52211 ( \52186 , \52185 );
nand \U$52212 ( \52187 , \52123 , \52186 );
buf \U$52213 ( \52188 , \52187 );
buf \U$52214 ( \52189 , \52188 );
nand \U$52215 ( \52190 , \52120 , \52189 );
buf \U$52216 ( \52191 , \52190 );
buf \U$52217 ( \52192 , \52191 );
xor \U$52218 ( \52193 , \52055 , \52192 );
buf \U$52219 ( \52194 , RIc0daaf8_113);
buf \U$52220 ( \52195 , RIc0d8de8_51);
xor \U$52221 ( \52196 , \52194 , \52195 );
buf \U$52222 ( \52197 , \52196 );
buf \U$52223 ( \52198 , \52197 );
not \U$52224 ( \52199 , \52198 );
buf \U$52225 ( \52200 , \14891 );
not \U$52226 ( \52201 , \52200 );
or \U$52227 ( \52202 , \52199 , \52201 );
buf \U$52228 ( \52203 , \12410 );
buf \U$52229 ( \52204 , \51518 );
nand \U$52230 ( \52205 , \52203 , \52204 );
buf \U$52231 ( \52206 , \52205 );
buf \U$52232 ( \52207 , \52206 );
nand \U$52233 ( \52208 , \52202 , \52207 );
buf \U$52234 ( \52209 , \52208 );
buf \U$52235 ( \52210 , \52209 );
xor \U$52236 ( \52211 , RIc0dacd8_117, RIc0d8c08_47);
buf \U$52237 ( \52212 , \52211 );
not \U$52238 ( \52213 , \52212 );
buf \U$52239 ( \52214 , \22350 );
not \U$52240 ( \52215 , \52214 );
or \U$52241 ( \52216 , \52213 , \52215 );
buf \U$52242 ( \52217 , \16559 );
buf \U$52243 ( \52218 , \51742 );
nand \U$52244 ( \52219 , \52217 , \52218 );
buf \U$52245 ( \52220 , \52219 );
buf \U$52246 ( \52221 , \52220 );
nand \U$52247 ( \52222 , \52216 , \52221 );
buf \U$52248 ( \52223 , \52222 );
buf \U$52249 ( \52224 , \52223 );
xor \U$52250 ( \52225 , \52210 , \52224 );
buf \U$52251 ( \52226 , RIc0da558_101);
buf \U$52252 ( \52227 , RIc0d9388_63);
and \U$52253 ( \52228 , \52226 , \52227 );
not \U$52254 ( \52229 , \52226 );
buf \U$52255 ( \52230 , \43939 );
and \U$52256 ( \52231 , \52229 , \52230 );
nor \U$52257 ( \52232 , \52228 , \52231 );
buf \U$52258 ( \52233 , \52232 );
buf \U$52259 ( \52234 , \52233 );
not \U$52260 ( \52235 , \52234 );
buf \U$52261 ( \52236 , \3535 );
not \U$52262 ( \52237 , \52236 );
or \U$52263 ( \52238 , \52235 , \52237 );
buf \U$52264 ( \52239 , \4049 );
buf \U$52265 ( \52240 , \51582 );
nand \U$52266 ( \52241 , \52239 , \52240 );
buf \U$52267 ( \52242 , \52241 );
buf \U$52268 ( \52243 , \52242 );
nand \U$52269 ( \52244 , \52238 , \52243 );
buf \U$52270 ( \52245 , \52244 );
buf \U$52271 ( \52246 , \52245 );
and \U$52272 ( \52247 , \52225 , \52246 );
and \U$52273 ( \52248 , \52210 , \52224 );
or \U$52274 ( \52249 , \52247 , \52248 );
buf \U$52275 ( \52250 , \52249 );
buf \U$52276 ( \52251 , \52250 );
buf \U$52277 ( \52252 , \51794 );
not \U$52278 ( \52253 , \52252 );
buf \U$52279 ( \52254 , \12303 );
not \U$52280 ( \52255 , \52254 );
or \U$52281 ( \52256 , \52253 , \52255 );
buf \U$52282 ( \52257 , \12278 );
buf \U$52283 ( \52258 , RIc0d8cf8_49);
buf \U$52284 ( \52259 , RIc0dabe8_115);
xor \U$52285 ( \52260 , \52258 , \52259 );
buf \U$52286 ( \52261 , \52260 );
buf \U$52287 ( \52262 , \52261 );
buf \U$52288 ( \52263 , \12293 );
nand \U$52289 ( \52264 , \52257 , \52262 , \52263 );
buf \U$52290 ( \52265 , \52264 );
buf \U$52291 ( \52266 , \52265 );
nand \U$52292 ( \52267 , \52256 , \52266 );
buf \U$52293 ( \52268 , \52267 );
buf \U$52294 ( \52269 , \52268 );
buf \U$52295 ( \52270 , \12584 );
buf \U$52296 ( \52271 , RIc0d9400_64);
and \U$52297 ( \52272 , \52270 , \52271 );
buf \U$52298 ( \52273 , \52272 );
buf \U$52299 ( \52274 , \52273 );
xor \U$52300 ( \52275 , \52269 , \52274 );
buf \U$52301 ( \52276 , RIc0da648_103);
buf \U$52302 ( \52277 , RIc0d9298_61);
xor \U$52303 ( \52278 , \52276 , \52277 );
buf \U$52304 ( \52279 , \52278 );
buf \U$52305 ( \52280 , \52279 );
not \U$52306 ( \52281 , \52280 );
buf \U$52307 ( \52282 , \17405 );
not \U$52308 ( \52283 , \52282 );
or \U$52309 ( \52284 , \52281 , \52283 );
buf \U$52310 ( \52285 , \13712 );
buf \U$52311 ( \52286 , \51771 );
nand \U$52312 ( \52287 , \52285 , \52286 );
buf \U$52313 ( \52288 , \52287 );
buf \U$52314 ( \52289 , \52288 );
nand \U$52315 ( \52290 , \52284 , \52289 );
buf \U$52316 ( \52291 , \52290 );
buf \U$52317 ( \52292 , \52291 );
and \U$52318 ( \52293 , \52275 , \52292 );
and \U$52319 ( \52294 , \52269 , \52274 );
or \U$52320 ( \52295 , \52293 , \52294 );
buf \U$52321 ( \52296 , \52295 );
buf \U$52322 ( \52297 , \52296 );
or \U$52323 ( \52298 , \52251 , \52297 );
buf \U$52324 ( \52299 , \51686 );
not \U$52325 ( \52300 , \52299 );
buf \U$52326 ( \52301 , \14352 );
not \U$52327 ( \52302 , \52301 );
or \U$52328 ( \52303 , \52300 , \52302 );
buf \U$52329 ( \52304 , \12540 );
and \U$52330 ( \52305 , RIc0daa08_111, \23372 );
not \U$52331 ( \52306 , RIc0daa08_111);
and \U$52332 ( \52307 , \52306 , RIc0d8ed8_53);
or \U$52333 ( \52308 , \52305 , \52307 );
buf \U$52334 ( \52309 , \52308 );
buf \U$52335 ( \52310 , \12517 );
nand \U$52336 ( \52311 , \52304 , \52309 , \52310 );
buf \U$52337 ( \52312 , \52311 );
buf \U$52338 ( \52313 , \52312 );
nand \U$52339 ( \52314 , \52303 , \52313 );
buf \U$52340 ( \52315 , \52314 );
buf \U$52341 ( \52316 , \52315 );
buf \U$52342 ( \52317 , \51756 );
not \U$52343 ( \52318 , \52317 );
buf \U$52344 ( \52319 , \13005 );
not \U$52345 ( \52320 , \52319 );
or \U$52346 ( \52321 , \52318 , \52320 );
buf \U$52347 ( \52322 , \45225 );
xor \U$52348 ( \52323 , RIc0dadc8_119, RIc0d8b18_45);
buf \U$52349 ( \52324 , \52323 );
buf \U$52350 ( \52325 , \12995 );
nand \U$52351 ( \52326 , \52322 , \52324 , \52325 );
buf \U$52352 ( \52327 , \52326 );
buf \U$52353 ( \52328 , \52327 );
nand \U$52354 ( \52329 , \52321 , \52328 );
buf \U$52355 ( \52330 , \52329 );
buf \U$52356 ( \52331 , \52330 );
xor \U$52357 ( \52332 , \52316 , \52331 );
buf \U$52358 ( \52333 , \12331 );
buf \U$52359 ( \52334 , RIc0d90b8_57);
buf \U$52360 ( \52335 , RIc0da828_107);
xnor \U$52361 ( \52336 , \52334 , \52335 );
buf \U$52362 ( \52337 , \52336 );
buf \U$52363 ( \52338 , \52337 );
or \U$52364 ( \52339 , \52333 , \52338 );
buf \U$52365 ( \52340 , \13270 );
buf \U$52366 ( \52341 , \51914 );
or \U$52367 ( \52342 , \52340 , \52341 );
nand \U$52368 ( \52343 , \52339 , \52342 );
buf \U$52369 ( \52344 , \52343 );
buf \U$52370 ( \52345 , \52344 );
and \U$52371 ( \52346 , \52332 , \52345 );
and \U$52372 ( \52347 , \52316 , \52331 );
or \U$52373 ( \52348 , \52346 , \52347 );
buf \U$52374 ( \52349 , \52348 );
buf \U$52375 ( \52350 , \52349 );
nand \U$52376 ( \52351 , \52298 , \52350 );
buf \U$52377 ( \52352 , \52351 );
buf \U$52378 ( \52353 , \52352 );
buf \U$52379 ( \52354 , \52250 );
buf \U$52380 ( \52355 , \52296 );
nand \U$52381 ( \52356 , \52354 , \52355 );
buf \U$52382 ( \52357 , \52356 );
buf \U$52383 ( \52358 , \52357 );
nand \U$52384 ( \52359 , \52353 , \52358 );
buf \U$52385 ( \52360 , \52359 );
buf \U$52386 ( \52361 , \52360 );
and \U$52387 ( \52362 , \52193 , \52361 );
and \U$52388 ( \52363 , \52055 , \52192 );
or \U$52389 ( \52364 , \52362 , \52363 );
buf \U$52390 ( \52365 , \52364 );
buf \U$52391 ( \52366 , \52365 );
xor \U$52392 ( \52367 , \52051 , \52366 );
xor \U$52393 ( \52368 , \51755 , \51769 );
xor \U$52394 ( \52369 , \52368 , \51784 );
buf \U$52395 ( \52370 , \52369 );
buf \U$52396 ( \52371 , \52370 );
not \U$52397 ( \52372 , \52371 );
xor \U$52398 ( \52373 , \51807 , \51824 );
xor \U$52399 ( \52374 , \52373 , \51843 );
buf \U$52400 ( \52375 , \52374 );
buf \U$52401 ( \52376 , \52375 );
not \U$52402 ( \52377 , \52376 );
or \U$52403 ( \52378 , \52372 , \52377 );
buf \U$52404 ( \52379 , \52375 );
buf \U$52405 ( \52380 , \52370 );
or \U$52406 ( \52381 , \52379 , \52380 );
xor \U$52407 ( \52382 , \51699 , \51716 );
xor \U$52408 ( \52383 , \52382 , \51733 );
buf \U$52409 ( \52384 , \52383 );
buf \U$52410 ( \52385 , \52384 );
nand \U$52411 ( \52386 , \52381 , \52385 );
buf \U$52412 ( \52387 , \52386 );
buf \U$52413 ( \52388 , \52387 );
nand \U$52414 ( \52389 , \52378 , \52388 );
buf \U$52415 ( \52390 , \52389 );
buf \U$52416 ( \52391 , \52390 );
xor \U$52417 ( \52392 , \51738 , \51789 );
xor \U$52418 ( \52393 , \52392 , \51848 );
buf \U$52419 ( \52394 , \52393 );
buf \U$52420 ( \52395 , \52394 );
xor \U$52421 ( \52396 , \52391 , \52395 );
xor \U$52422 ( \52397 , \51869 , \51890 );
xor \U$52423 ( \52398 , \52397 , \51950 );
buf \U$52424 ( \52399 , \52398 );
buf \U$52425 ( \52400 , \52399 );
and \U$52426 ( \52401 , \52396 , \52400 );
and \U$52427 ( \52402 , \52391 , \52395 );
or \U$52428 ( \52403 , \52401 , \52402 );
buf \U$52429 ( \52404 , \52403 );
buf \U$52430 ( \52405 , \52404 );
and \U$52431 ( \52406 , \52367 , \52405 );
and \U$52432 ( \52407 , \52051 , \52366 );
or \U$52433 ( \52408 , \52406 , \52407 );
buf \U$52434 ( \52409 , \52408 );
buf \U$52435 ( \52410 , \52409 );
xor \U$52436 ( \52411 , \51999 , \52003 );
xor \U$52437 ( \52412 , \52411 , \52007 );
buf \U$52438 ( \52413 , \52412 );
buf \U$52439 ( \52414 , \52413 );
not \U$52440 ( \52415 , \52414 );
buf \U$52441 ( \52416 , \52349 );
not \U$52442 ( \52417 , \52416 );
buf \U$52443 ( \52418 , \52296 );
not \U$52444 ( \52419 , \52418 );
buf \U$52445 ( \52420 , \52419 );
buf \U$52446 ( \52421 , \52420 );
not \U$52447 ( \52422 , \52421 );
and \U$52448 ( \52423 , \52417 , \52422 );
buf \U$52449 ( \52424 , \52349 );
buf \U$52450 ( \52425 , \52420 );
and \U$52451 ( \52426 , \52424 , \52425 );
nor \U$52452 ( \52427 , \52423 , \52426 );
buf \U$52453 ( \52428 , \52427 );
buf \U$52454 ( \52429 , \52428 );
buf \U$52455 ( \52430 , \52250 );
and \U$52456 ( \52431 , \52429 , \52430 );
not \U$52457 ( \52432 , \52429 );
buf \U$52458 ( \52433 , \52250 );
not \U$52459 ( \52434 , \52433 );
buf \U$52460 ( \52435 , \52434 );
buf \U$52461 ( \52436 , \52435 );
and \U$52462 ( \52437 , \52432 , \52436 );
nor \U$52463 ( \52438 , \52431 , \52437 );
buf \U$52464 ( \52439 , \52438 );
not \U$52465 ( \52440 , \52439 );
buf \U$52466 ( \52441 , \52109 );
not \U$52467 ( \52442 , \52441 );
buf \U$52468 ( \52443 , \52185 );
not \U$52469 ( \52444 , \52443 );
buf \U$52470 ( \52445 , \52444 );
buf \U$52471 ( \52446 , \52445 );
not \U$52472 ( \52447 , \52446 );
or \U$52473 ( \52448 , \52442 , \52447 );
buf \U$52474 ( \52449 , \52109 );
buf \U$52475 ( \52450 , \52445 );
or \U$52476 ( \52451 , \52449 , \52450 );
nand \U$52477 ( \52452 , \52448 , \52451 );
buf \U$52478 ( \52453 , \52452 );
buf \U$52479 ( \52454 , \52453 );
buf \U$52480 ( \52455 , \52117 );
not \U$52481 ( \52456 , \52455 );
buf \U$52482 ( \52457 , \52456 );
buf \U$52483 ( \52458 , \52457 );
and \U$52484 ( \52459 , \52454 , \52458 );
not \U$52485 ( \52460 , \52454 );
buf \U$52486 ( \52461 , \52117 );
and \U$52487 ( \52462 , \52460 , \52461 );
nor \U$52488 ( \52463 , \52459 , \52462 );
buf \U$52489 ( \52464 , \52463 );
not \U$52490 ( \52465 , \52464 );
or \U$52491 ( \52466 , \52440 , \52465 );
buf \U$52492 ( \52467 , RIc0d87d0_38);
buf \U$52493 ( \52468 , RIc0db188_127);
xor \U$52494 ( \52469 , \52467 , \52468 );
buf \U$52495 ( \52470 , \52469 );
buf \U$52496 ( \52471 , \52470 );
not \U$52497 ( \52472 , \52471 );
buf \U$52498 ( \52473 , \44639 );
not \U$52499 ( \52474 , \52473 );
or \U$52500 ( \52475 , \52472 , \52474 );
buf \U$52501 ( \52476 , \52127 );
buf \U$52502 ( \52477 , RIc0db200_128);
nand \U$52503 ( \52478 , \52476 , \52477 );
buf \U$52504 ( \52479 , \52478 );
buf \U$52505 ( \52480 , \52479 );
nand \U$52506 ( \52481 , \52475 , \52480 );
buf \U$52507 ( \52482 , \52481 );
buf \U$52508 ( \52483 , \52482 );
buf \U$52509 ( \52484 , RIc0da918_109);
buf \U$52510 ( \52485 , RIc0d9040_56);
xor \U$52511 ( \52486 , \52484 , \52485 );
buf \U$52512 ( \52487 , \52486 );
buf \U$52513 ( \52488 , \52487 );
not \U$52514 ( \52489 , \52488 );
buf \U$52515 ( \52490 , \27660 );
not \U$52516 ( \52491 , \52490 );
or \U$52517 ( \52492 , \52489 , \52491 );
buf \U$52518 ( \52493 , \13426 );
buf \U$52519 ( \52494 , \52094 );
nand \U$52520 ( \52495 , \52493 , \52494 );
buf \U$52521 ( \52496 , \52495 );
buf \U$52522 ( \52497 , \52496 );
nand \U$52523 ( \52498 , \52492 , \52497 );
buf \U$52524 ( \52499 , \52498 );
buf \U$52525 ( \52500 , \52499 );
xor \U$52526 ( \52501 , \52483 , \52500 );
buf \U$52527 ( \52502 , RIc0d89b0_42);
buf \U$52528 ( \52503 , RIc0dafa8_123);
xor \U$52529 ( \52504 , \52502 , \52503 );
buf \U$52530 ( \52505 , \52504 );
buf \U$52531 ( \52506 , \52505 );
not \U$52532 ( \52507 , \52506 );
buf \U$52533 ( \52508 , \14982 );
not \U$52534 ( \52509 , \52508 );
or \U$52535 ( \52510 , \52507 , \52509 );
buf \U$52536 ( \52511 , \16692 );
buf \U$52537 ( \52512 , \52145 );
nand \U$52538 ( \52513 , \52511 , \52512 );
buf \U$52539 ( \52514 , \52513 );
buf \U$52540 ( \52515 , \52514 );
nand \U$52541 ( \52516 , \52510 , \52515 );
buf \U$52542 ( \52517 , \52516 );
buf \U$52543 ( \52518 , \52517 );
and \U$52544 ( \52519 , \52501 , \52518 );
and \U$52545 ( \52520 , \52483 , \52500 );
or \U$52546 ( \52521 , \52519 , \52520 );
buf \U$52547 ( \52522 , \52521 );
buf \U$52548 ( \52523 , \52522 );
not \U$52549 ( \52524 , \40787 );
buf \U$52550 ( \52525 , RIc0da738_105);
buf \U$52551 ( \52526 , RIc0d9220_60);
xnor \U$52552 ( \52527 , \52525 , \52526 );
buf \U$52553 ( \52528 , \52527 );
not \U$52554 ( \52529 , \52528 );
and \U$52555 ( \52530 , \52524 , \52529 );
buf \U$52556 ( \52531 , \52065 );
not \U$52557 ( \52532 , \52531 );
buf \U$52558 ( \52533 , \15650 );
nor \U$52559 ( \52534 , \52532 , \52533 );
buf \U$52560 ( \52535 , \52534 );
nor \U$52561 ( \52536 , \52530 , \52535 );
buf \U$52562 ( \52537 , \52536 );
not \U$52563 ( \52538 , \52537 );
xor \U$52564 ( \52539 , RIc0daeb8_121, RIc0d8aa0_44);
buf \U$52565 ( \52540 , \52539 );
not \U$52566 ( \52541 , \52540 );
buf \U$52567 ( \52542 , \16382 );
not \U$52568 ( \52543 , \52542 );
or \U$52569 ( \52544 , \52541 , \52543 );
buf \U$52570 ( \52545 , \13314 );
buf \U$52571 ( \52546 , \52083 );
nand \U$52572 ( \52547 , \52545 , \52546 );
buf \U$52573 ( \52548 , \52547 );
buf \U$52574 ( \52549 , \52548 );
nand \U$52575 ( \52550 , \52544 , \52549 );
buf \U$52576 ( \52551 , \52550 );
buf \U$52577 ( \52552 , \52551 );
not \U$52578 ( \52553 , \52552 );
buf \U$52579 ( \52554 , \52553 );
buf \U$52580 ( \52555 , \52554 );
not \U$52581 ( \52556 , \52555 );
or \U$52582 ( \52557 , \52538 , \52556 );
buf \U$52583 ( \52558 , RIc0d8f50_54);
buf \U$52584 ( \52559 , RIc0daa08_111);
xnor \U$52585 ( \52560 , \52558 , \52559 );
buf \U$52586 ( \52561 , \52560 );
buf \U$52587 ( \52562 , \52561 );
not \U$52588 ( \52563 , \52562 );
buf \U$52589 ( \52564 , \52563 );
buf \U$52590 ( \52565 , \52564 );
not \U$52591 ( \52566 , \52565 );
buf \U$52592 ( \52567 , \14346 );
not \U$52593 ( \52568 , \52567 );
or \U$52594 ( \52569 , \52566 , \52568 );
buf \U$52595 ( \52570 , \14106 );
buf \U$52596 ( \52571 , \52308 );
nand \U$52597 ( \52572 , \52570 , \52571 );
buf \U$52598 ( \52573 , \52572 );
buf \U$52599 ( \52574 , \52573 );
nand \U$52600 ( \52575 , \52569 , \52574 );
buf \U$52601 ( \52576 , \52575 );
buf \U$52602 ( \52577 , \52576 );
nand \U$52603 ( \52578 , \52557 , \52577 );
buf \U$52604 ( \52579 , \52578 );
buf \U$52605 ( \52580 , \52579 );
buf \U$52606 ( \52581 , \52536 );
not \U$52607 ( \52582 , \52581 );
buf \U$52608 ( \52583 , \52551 );
nand \U$52609 ( \52584 , \52582 , \52583 );
buf \U$52610 ( \52585 , \52584 );
buf \U$52611 ( \52586 , \52585 );
nand \U$52612 ( \52587 , \52580 , \52586 );
buf \U$52613 ( \52588 , \52587 );
buf \U$52614 ( \52589 , \52588 );
xor \U$52615 ( \52590 , \52523 , \52589 );
xor \U$52616 ( \52591 , \52210 , \52224 );
xor \U$52617 ( \52592 , \52591 , \52246 );
buf \U$52618 ( \52593 , \52592 );
buf \U$52619 ( \52594 , \52593 );
and \U$52620 ( \52595 , \52590 , \52594 );
and \U$52621 ( \52596 , \52523 , \52589 );
or \U$52622 ( \52597 , \52595 , \52596 );
buf \U$52623 ( \52598 , \52597 );
nand \U$52624 ( \52599 , \52466 , \52598 );
buf \U$52625 ( \52600 , \52599 );
buf \U$52626 ( \52601 , \52439 );
not \U$52627 ( \52602 , \52601 );
buf \U$52628 ( \52603 , \52464 );
not \U$52629 ( \52604 , \52603 );
buf \U$52630 ( \52605 , \52604 );
buf \U$52631 ( \52606 , \52605 );
nand \U$52632 ( \52607 , \52602 , \52606 );
buf \U$52633 ( \52608 , \52607 );
buf \U$52634 ( \52609 , \52608 );
nand \U$52635 ( \52610 , \52600 , \52609 );
buf \U$52636 ( \52611 , \52610 );
buf \U$52637 ( \52612 , \52611 );
not \U$52638 ( \52613 , \52612 );
or \U$52639 ( \52614 , \52415 , \52613 );
buf \U$52640 ( \52615 , \52611 );
buf \U$52641 ( \52616 , \52413 );
or \U$52642 ( \52617 , \52615 , \52616 );
and \U$52643 ( \52618 , \51908 , \51940 );
not \U$52644 ( \52619 , \51908 );
and \U$52645 ( \52620 , \52619 , \51929 );
nor \U$52646 ( \52621 , \52618 , \52620 );
xor \U$52647 ( \52622 , \52621 , \51933 );
buf \U$52648 ( \52623 , \52622 );
xor \U$52649 ( \52624 , \52269 , \52274 );
xor \U$52650 ( \52625 , \52624 , \52292 );
buf \U$52651 ( \52626 , \52625 );
buf \U$52652 ( \52627 , \52626 );
not \U$52653 ( \52628 , \52627 );
buf \U$52654 ( \52629 , \52157 );
buf \U$52655 ( \52630 , \52139 );
xor \U$52656 ( \52631 , \52629 , \52630 );
buf \U$52657 ( \52632 , \52631 );
buf \U$52658 ( \52633 , \52632 );
buf \U$52659 ( \52634 , \52179 );
xor \U$52660 ( \52635 , \52633 , \52634 );
buf \U$52661 ( \52636 , \52635 );
buf \U$52662 ( \52637 , \52636 );
not \U$52663 ( \52638 , \52637 );
or \U$52664 ( \52639 , \52628 , \52638 );
buf \U$52665 ( \52640 , \52636 );
buf \U$52666 ( \52641 , \52626 );
or \U$52667 ( \52642 , \52640 , \52641 );
xor \U$52668 ( \52643 , \52316 , \52331 );
xor \U$52669 ( \52644 , \52643 , \52345 );
buf \U$52670 ( \52645 , \52644 );
buf \U$52671 ( \52646 , \52645 );
nand \U$52672 ( \52647 , \52642 , \52646 );
buf \U$52673 ( \52648 , \52647 );
buf \U$52674 ( \52649 , \52648 );
nand \U$52675 ( \52650 , \52639 , \52649 );
buf \U$52676 ( \52651 , \52650 );
buf \U$52677 ( \52652 , \52651 );
xor \U$52678 ( \52653 , \52623 , \52652 );
buf \U$52679 ( \52654 , RIc0da648_103);
buf \U$52680 ( \52655 , RIc0d9310_62);
xor \U$52681 ( \52656 , \52654 , \52655 );
buf \U$52682 ( \52657 , \52656 );
buf \U$52683 ( \52658 , \52657 );
not \U$52684 ( \52659 , \52658 );
buf \U$52685 ( \52660 , \13042 );
not \U$52686 ( \52661 , \52660 );
or \U$52687 ( \52662 , \52659 , \52661 );
buf \U$52688 ( \52663 , \13048 );
buf \U$52689 ( \52664 , \52279 );
nand \U$52690 ( \52665 , \52663 , \52664 );
buf \U$52691 ( \52666 , \52665 );
buf \U$52692 ( \52667 , \52666 );
nand \U$52693 ( \52668 , \52662 , \52667 );
buf \U$52694 ( \52669 , \52668 );
buf \U$52695 ( \52670 , \52669 );
not \U$52696 ( \52671 , \52670 );
buf \U$52697 ( \52672 , RIc0d9400_64);
buf \U$52698 ( \52673 , RIc0da5d0_102);
nand \U$52699 ( \52674 , \52672 , \52673 );
buf \U$52700 ( \52675 , \52674 );
buf \U$52701 ( \52676 , \52675 );
buf \U$52702 ( \52677 , RIc0da558_101);
and \U$52703 ( \52678 , \52676 , \52677 );
buf \U$52704 ( \52679 , \52678 );
buf \U$52705 ( \52680 , \52679 );
buf \U$52706 ( \52681 , RIc0d9400_64);
buf \U$52707 ( \52682 , RIc0da5d0_102);
or \U$52708 ( \52683 , \52681 , \52682 );
buf \U$52709 ( \52684 , RIc0da648_103);
nand \U$52710 ( \52685 , \52683 , \52684 );
buf \U$52711 ( \52686 , \52685 );
buf \U$52712 ( \52687 , \52686 );
nand \U$52713 ( \52688 , \52680 , \52687 );
buf \U$52714 ( \52689 , \52688 );
buf \U$52715 ( \52690 , \52689 );
nor \U$52716 ( \52691 , \52671 , \52690 );
buf \U$52717 ( \52692 , \52691 );
buf \U$52718 ( \52693 , \52692 );
xor \U$52719 ( \52694 , RIc0daaf8_113, RIc0d8e60_52);
buf \U$52720 ( \52695 , \52694 );
not \U$52721 ( \52696 , \52695 );
buf \U$52722 ( \52697 , \33224 );
not \U$52723 ( \52698 , \52697 );
or \U$52724 ( \52699 , \52696 , \52698 );
buf \U$52725 ( \52700 , \12410 );
buf \U$52726 ( \52701 , \52197 );
nand \U$52727 ( \52702 , \52700 , \52701 );
buf \U$52728 ( \52703 , \52702 );
buf \U$52729 ( \52704 , \52703 );
nand \U$52730 ( \52705 , \52699 , \52704 );
buf \U$52731 ( \52706 , \52705 );
buf \U$52732 ( \52707 , \52706 );
not \U$52733 ( \52708 , \52707 );
xor \U$52734 ( \52709 , RIc0da828_107, RIc0d9130_58);
buf \U$52735 ( \52710 , \52709 );
not \U$52736 ( \52711 , \52710 );
buf \U$52737 ( \52712 , \34202 );
not \U$52738 ( \52713 , \52712 );
or \U$52739 ( \52714 , \52711 , \52713 );
buf \U$52740 ( \52715 , \52337 );
not \U$52741 ( \52716 , \52715 );
buf \U$52742 ( \52717 , \16071 );
nand \U$52743 ( \52718 , \52716 , \52717 );
buf \U$52744 ( \52719 , \52718 );
buf \U$52745 ( \52720 , \52719 );
nand \U$52746 ( \52721 , \52714 , \52720 );
buf \U$52747 ( \52722 , \52721 );
buf \U$52748 ( \52723 , \52722 );
not \U$52749 ( \52724 , \52723 );
or \U$52750 ( \52725 , \52708 , \52724 );
buf \U$52751 ( \52726 , \52722 );
buf \U$52752 ( \52727 , \52706 );
or \U$52753 ( \52728 , \52726 , \52727 );
buf \U$52754 ( \52729 , RIc0dadc8_119);
buf \U$52755 ( \52730 , RIc0d8b90_46);
xor \U$52756 ( \52731 , \52729 , \52730 );
buf \U$52757 ( \52732 , \52731 );
buf \U$52758 ( \52733 , \52732 );
not \U$52759 ( \52734 , \52733 );
buf \U$52760 ( \52735 , \25542 );
not \U$52761 ( \52736 , \52735 );
or \U$52762 ( \52737 , \52734 , \52736 );
buf \U$52763 ( \52738 , \13953 );
buf \U$52764 ( \52739 , \52323 );
nand \U$52765 ( \52740 , \52738 , \52739 );
buf \U$52766 ( \52741 , \52740 );
buf \U$52767 ( \52742 , \52741 );
nand \U$52768 ( \52743 , \52737 , \52742 );
buf \U$52769 ( \52744 , \52743 );
buf \U$52770 ( \52745 , \52744 );
nand \U$52771 ( \52746 , \52728 , \52745 );
buf \U$52772 ( \52747 , \52746 );
buf \U$52773 ( \52748 , \52747 );
nand \U$52774 ( \52749 , \52725 , \52748 );
buf \U$52775 ( \52750 , \52749 );
buf \U$52776 ( \52751 , \52750 );
xor \U$52777 ( \52752 , \52693 , \52751 );
buf \U$52778 ( \52753 , RIc0d8c80_48);
buf \U$52779 ( \52754 , RIc0dacd8_117);
xor \U$52780 ( \52755 , \52753 , \52754 );
buf \U$52781 ( \52756 , \52755 );
buf \U$52782 ( \52757 , \52756 );
not \U$52783 ( \52758 , \52757 );
buf \U$52784 ( \52759 , \22350 );
not \U$52785 ( \52760 , \52759 );
or \U$52786 ( \52761 , \52758 , \52760 );
buf \U$52787 ( \52762 , \22356 );
buf \U$52788 ( \52763 , \52211 );
nand \U$52789 ( \52764 , \52762 , \52763 );
buf \U$52790 ( \52765 , \52764 );
buf \U$52791 ( \52766 , \52765 );
nand \U$52792 ( \52767 , \52761 , \52766 );
buf \U$52793 ( \52768 , \52767 );
buf \U$52794 ( \52769 , \52768 );
buf \U$52795 ( \52770 , RIc0d8d70_50);
buf \U$52796 ( \52771 , RIc0dabe8_115);
xor \U$52797 ( \52772 , \52770 , \52771 );
buf \U$52798 ( \52773 , \52772 );
buf \U$52799 ( \52774 , \52773 );
not \U$52800 ( \52775 , \52774 );
buf \U$52801 ( \52776 , \26466 );
not \U$52802 ( \52777 , \52776 );
or \U$52803 ( \52778 , \52775 , \52777 );
buf \U$52804 ( \52779 , \12303 );
buf \U$52805 ( \52780 , \52261 );
nand \U$52806 ( \52781 , \52779 , \52780 );
buf \U$52807 ( \52782 , \52781 );
buf \U$52808 ( \52783 , \52782 );
nand \U$52809 ( \52784 , \52778 , \52783 );
buf \U$52810 ( \52785 , \52784 );
buf \U$52811 ( \52786 , \52785 );
or \U$52812 ( \52787 , \52769 , \52786 );
buf \U$52813 ( \52788 , RIc0d9400_64);
buf \U$52814 ( \52789 , RIc0da558_101);
xor \U$52815 ( \52790 , \52788 , \52789 );
buf \U$52816 ( \52791 , \52790 );
buf \U$52817 ( \52792 , \52791 );
not \U$52818 ( \52793 , \52792 );
buf \U$52819 ( \52794 , \22631 );
not \U$52820 ( \52795 , \52794 );
or \U$52821 ( \52796 , \52793 , \52795 );
buf \U$52822 ( \52797 , \4049 );
buf \U$52823 ( \52798 , \52233 );
nand \U$52824 ( \52799 , \52797 , \52798 );
buf \U$52825 ( \52800 , \52799 );
buf \U$52826 ( \52801 , \52800 );
nand \U$52827 ( \52802 , \52796 , \52801 );
buf \U$52828 ( \52803 , \52802 );
buf \U$52829 ( \52804 , \52803 );
nand \U$52830 ( \52805 , \52787 , \52804 );
buf \U$52831 ( \52806 , \52805 );
buf \U$52832 ( \52807 , \52806 );
buf \U$52833 ( \52808 , \52785 );
buf \U$52834 ( \52809 , \52768 );
nand \U$52835 ( \52810 , \52808 , \52809 );
buf \U$52836 ( \52811 , \52810 );
buf \U$52837 ( \52812 , \52811 );
nand \U$52838 ( \52813 , \52807 , \52812 );
buf \U$52839 ( \52814 , \52813 );
buf \U$52840 ( \52815 , \52814 );
and \U$52841 ( \52816 , \52752 , \52815 );
and \U$52842 ( \52817 , \52693 , \52751 );
or \U$52843 ( \52818 , \52816 , \52817 );
buf \U$52844 ( \52819 , \52818 );
buf \U$52845 ( \52820 , \52819 );
and \U$52846 ( \52821 , \52653 , \52820 );
and \U$52847 ( \52822 , \52623 , \52652 );
or \U$52848 ( \52823 , \52821 , \52822 );
buf \U$52849 ( \52824 , \52823 );
buf \U$52850 ( \52825 , \52824 );
nand \U$52851 ( \52826 , \52617 , \52825 );
buf \U$52852 ( \52827 , \52826 );
buf \U$52853 ( \52828 , \52827 );
nand \U$52854 ( \52829 , \52614 , \52828 );
buf \U$52855 ( \52830 , \52829 );
buf \U$52856 ( \52831 , \52830 );
buf \U$52857 ( \52832 , \51683 );
not \U$52858 ( \52833 , \52832 );
buf \U$52859 ( \52834 , \51852 );
buf \U$52860 ( \52835 , \51679 );
xnor \U$52861 ( \52836 , \52834 , \52835 );
buf \U$52862 ( \52837 , \52836 );
buf \U$52863 ( \52838 , \52837 );
not \U$52864 ( \52839 , \52838 );
or \U$52865 ( \52840 , \52833 , \52839 );
buf \U$52866 ( \52841 , \51683 );
buf \U$52867 ( \52842 , \52837 );
or \U$52868 ( \52843 , \52841 , \52842 );
nand \U$52869 ( \52844 , \52840 , \52843 );
buf \U$52870 ( \52845 , \52844 );
buf \U$52871 ( \52846 , \52845 );
xor \U$52872 ( \52847 , \52831 , \52846 );
xor \U$52873 ( \52848 , \51976 , \51954 );
xor \U$52874 ( \52849 , \52848 , \52011 );
buf \U$52875 ( \52850 , \52849 );
and \U$52876 ( \52851 , \52847 , \52850 );
and \U$52877 ( \52852 , \52831 , \52846 );
or \U$52878 ( \52853 , \52851 , \52852 );
buf \U$52879 ( \52854 , \52853 );
buf \U$52880 ( \52855 , \52854 );
xor \U$52881 ( \52856 , \52410 , \52855 );
xor \U$52882 ( \52857 , \52031 , \52035 );
xor \U$52883 ( \52858 , \52857 , \52040 );
buf \U$52884 ( \52859 , \52858 );
buf \U$52885 ( \52860 , \52859 );
and \U$52886 ( \52861 , \52856 , \52860 );
and \U$52887 ( \52862 , \52410 , \52855 );
or \U$52888 ( \52863 , \52861 , \52862 );
buf \U$52889 ( \52864 , \52863 );
buf \U$52890 ( \52865 , \52864 );
nand \U$52891 ( \52866 , \52048 , \52865 );
buf \U$52892 ( \52867 , \52866 );
not \U$52893 ( \52868 , \52867 );
xor \U$52894 ( \52869 , \52410 , \52855 );
xor \U$52895 ( \52870 , \52869 , \52860 );
buf \U$52896 ( \52871 , \52870 );
buf \U$52897 ( \52872 , \52871 );
xor \U$52898 ( \52873 , \52055 , \52192 );
xor \U$52899 ( \52874 , \52873 , \52361 );
buf \U$52900 ( \52875 , \52874 );
buf \U$52901 ( \52876 , \52875 );
xor \U$52902 ( \52877 , \52391 , \52395 );
xor \U$52903 ( \52878 , \52877 , \52400 );
buf \U$52904 ( \52879 , \52878 );
buf \U$52905 ( \52880 , \52879 );
xor \U$52906 ( \52881 , \52876 , \52880 );
xor \U$52907 ( \52882 , \52375 , \52370 );
xor \U$52908 ( \52883 , \52882 , \52384 );
buf \U$52909 ( \52884 , \52883 );
xor \U$52910 ( \52885 , \52073 , \52091 );
xor \U$52911 ( \52886 , \52885 , \52105 );
buf \U$52912 ( \52887 , \52886 );
buf \U$52913 ( \52888 , \52887 );
buf \U$52914 ( \52889 , \17992 );
buf \U$52915 ( \52890 , RIc0db098_125);
buf \U$52916 ( \52891 , RIc0d88c0_40);
xor \U$52917 ( \52892 , \52890 , \52891 );
buf \U$52918 ( \52893 , \52892 );
buf \U$52919 ( \52894 , \52893 );
not \U$52920 ( \52895 , \52894 );
buf \U$52921 ( \52896 , \52895 );
buf \U$52922 ( \52897 , \52896 );
or \U$52923 ( \52898 , \52889 , \52897 );
buf \U$52924 ( \52899 , \22744 );
buf \U$52925 ( \52900 , \52167 );
not \U$52926 ( \52901 , \52900 );
buf \U$52927 ( \52902 , \52901 );
buf \U$52928 ( \52903 , \52902 );
or \U$52929 ( \52904 , \52899 , \52903 );
nand \U$52930 ( \52905 , \52898 , \52904 );
buf \U$52931 ( \52906 , \52905 );
buf \U$52932 ( \52907 , \52906 );
buf \U$52933 ( \52908 , \52689 );
not \U$52934 ( \52909 , \52908 );
buf \U$52935 ( \52910 , \52669 );
not \U$52936 ( \52911 , \52910 );
or \U$52937 ( \52912 , \52909 , \52911 );
buf \U$52938 ( \52913 , \52669 );
buf \U$52939 ( \52914 , \52689 );
or \U$52940 ( \52915 , \52913 , \52914 );
nand \U$52941 ( \52916 , \52912 , \52915 );
buf \U$52942 ( \52917 , \52916 );
buf \U$52943 ( \52918 , \52917 );
xor \U$52944 ( \52919 , \52907 , \52918 );
buf \U$52945 ( \52920 , \16676 );
buf \U$52946 ( \52921 , RIc0d9400_64);
and \U$52947 ( \52922 , \52920 , \52921 );
buf \U$52948 ( \52923 , \52922 );
buf \U$52949 ( \52924 , \52923 );
xor \U$52950 ( \52925 , RIc0da738_105, RIc0d9298_61);
buf \U$52951 ( \52926 , \52925 );
not \U$52952 ( \52927 , \52926 );
buf \U$52953 ( \52928 , \12736 );
not \U$52954 ( \52929 , \52928 );
or \U$52955 ( \52930 , \52927 , \52929 );
buf \U$52956 ( \52931 , \52528 );
not \U$52957 ( \52932 , \52931 );
buf \U$52958 ( \52933 , \12744 );
nand \U$52959 ( \52934 , \52932 , \52933 );
buf \U$52960 ( \52935 , \52934 );
buf \U$52961 ( \52936 , \52935 );
nand \U$52962 ( \52937 , \52930 , \52936 );
buf \U$52963 ( \52938 , \52937 );
buf \U$52964 ( \52939 , \52938 );
xor \U$52965 ( \52940 , \52924 , \52939 );
buf \U$52966 ( \52941 , RIc0d8de8_51);
buf \U$52967 ( \52942 , RIc0dabe8_115);
xor \U$52968 ( \52943 , \52941 , \52942 );
buf \U$52969 ( \52944 , \52943 );
buf \U$52970 ( \52945 , \52944 );
not \U$52971 ( \52946 , \52945 );
buf \U$52972 ( \52947 , \26466 );
not \U$52973 ( \52948 , \52947 );
or \U$52974 ( \52949 , \52946 , \52948 );
buf \U$52975 ( \52950 , \12303 );
buf \U$52976 ( \52951 , \52773 );
nand \U$52977 ( \52952 , \52950 , \52951 );
buf \U$52978 ( \52953 , \52952 );
buf \U$52979 ( \52954 , \52953 );
nand \U$52980 ( \52955 , \52949 , \52954 );
buf \U$52981 ( \52956 , \52955 );
buf \U$52982 ( \52957 , \52956 );
and \U$52983 ( \52958 , \52940 , \52957 );
and \U$52984 ( \52959 , \52924 , \52939 );
or \U$52985 ( \52960 , \52958 , \52959 );
buf \U$52986 ( \52961 , \52960 );
buf \U$52987 ( \52962 , \52961 );
and \U$52988 ( \52963 , \52919 , \52962 );
and \U$52989 ( \52964 , \52907 , \52918 );
or \U$52990 ( \52965 , \52963 , \52964 );
buf \U$52991 ( \52966 , \52965 );
buf \U$52992 ( \52967 , \52966 );
xor \U$52993 ( \52968 , \52888 , \52967 );
xor \U$52994 ( \52969 , RIc0db098_125, RIc0d8938_41);
buf \U$52995 ( \52970 , \52969 );
not \U$52996 ( \52971 , \52970 );
buf \U$52997 ( \52972 , \17995 );
not \U$52998 ( \52973 , \52972 );
or \U$52999 ( \52974 , \52971 , \52973 );
buf \U$53000 ( \52975 , \15793 );
buf \U$53001 ( \52976 , \52893 );
nand \U$53002 ( \52977 , \52975 , \52976 );
buf \U$53003 ( \52978 , \52977 );
buf \U$53004 ( \52979 , \52978 );
nand \U$53005 ( \52980 , \52974 , \52979 );
buf \U$53006 ( \52981 , \52980 );
not \U$53007 ( \52982 , \52981 );
buf \U$53008 ( \52983 , \12532 );
not \U$53009 ( \52984 , \52983 );
buf \U$53010 ( \52985 , RIc0daa08_111);
buf \U$53011 ( \52986 , RIc0d8fc8_55);
xnor \U$53012 ( \52987 , \52985 , \52986 );
buf \U$53013 ( \52988 , \52987 );
buf \U$53014 ( \52989 , \52988 );
not \U$53015 ( \52990 , \52989 );
and \U$53016 ( \52991 , \52984 , \52990 );
buf \U$53017 ( \52992 , \14353 );
not \U$53018 ( \52993 , \52992 );
buf \U$53019 ( \52994 , \52561 );
nor \U$53020 ( \52995 , \52993 , \52994 );
buf \U$53021 ( \52996 , \52995 );
buf \U$53022 ( \52997 , \52996 );
nor \U$53023 ( \52998 , \52991 , \52997 );
buf \U$53024 ( \52999 , \52998 );
nand \U$53025 ( \53000 , \52982 , \52999 );
not \U$53026 ( \53001 , \53000 );
buf \U$53027 ( \53002 , RIc0d8cf8_49);
buf \U$53028 ( \53003 , RIc0dacd8_117);
xor \U$53029 ( \53004 , \53002 , \53003 );
buf \U$53030 ( \53005 , \53004 );
buf \U$53031 ( \53006 , \53005 );
not \U$53032 ( \53007 , \53006 );
buf \U$53033 ( \53008 , \22350 );
not \U$53034 ( \53009 , \53008 );
or \U$53035 ( \53010 , \53007 , \53009 );
buf \U$53036 ( \53011 , \12937 );
buf \U$53037 ( \53012 , \52756 );
nand \U$53038 ( \53013 , \53011 , \53012 );
buf \U$53039 ( \53014 , \53013 );
buf \U$53040 ( \53015 , \53014 );
nand \U$53041 ( \53016 , \53010 , \53015 );
buf \U$53042 ( \53017 , \53016 );
not \U$53043 ( \53018 , \53017 );
or \U$53044 ( \53019 , \53001 , \53018 );
buf \U$53045 ( \53020 , \52999 );
not \U$53046 ( \53021 , \53020 );
buf \U$53047 ( \53022 , \52981 );
nand \U$53048 ( \53023 , \53021 , \53022 );
buf \U$53049 ( \53024 , \53023 );
nand \U$53050 ( \53025 , \53019 , \53024 );
buf \U$53051 ( \53026 , \53025 );
not \U$53052 ( \53027 , \53026 );
xor \U$53053 ( \53028 , RIc0da918_109, RIc0d90b8_57);
buf \U$53054 ( \53029 , \53028 );
not \U$53055 ( \53030 , \53029 );
buf \U$53056 ( \53031 , \21959 );
not \U$53057 ( \53032 , \53031 );
or \U$53058 ( \53033 , \53030 , \53032 );
buf \U$53059 ( \53034 , \20211 );
buf \U$53060 ( \53035 , \52487 );
nand \U$53061 ( \53036 , \53034 , \53035 );
buf \U$53062 ( \53037 , \53036 );
buf \U$53063 ( \53038 , \53037 );
nand \U$53064 ( \53039 , \53033 , \53038 );
buf \U$53065 ( \53040 , \53039 );
buf \U$53066 ( \53041 , \53040 );
buf \U$53067 ( \53042 , RIc0d9388_63);
buf \U$53068 ( \53043 , RIc0da648_103);
xor \U$53069 ( \53044 , \53042 , \53043 );
buf \U$53070 ( \53045 , \53044 );
buf \U$53071 ( \53046 , \53045 );
not \U$53072 ( \53047 , \53046 );
buf \U$53073 ( \53048 , \16578 );
not \U$53074 ( \53049 , \53048 );
or \U$53075 ( \53050 , \53047 , \53049 );
buf \U$53076 ( \53051 , \18416 );
buf \U$53077 ( \53052 , \52657 );
nand \U$53078 ( \53053 , \53051 , \53052 );
buf \U$53079 ( \53054 , \53053 );
buf \U$53080 ( \53055 , \53054 );
nand \U$53081 ( \53056 , \53050 , \53055 );
buf \U$53082 ( \53057 , \53056 );
buf \U$53083 ( \53058 , \53057 );
xor \U$53084 ( \53059 , \53041 , \53058 );
buf \U$53085 ( \53060 , RIc0d91a8_59);
buf \U$53086 ( \53061 , RIc0da828_107);
xor \U$53087 ( \53062 , \53060 , \53061 );
buf \U$53088 ( \53063 , \53062 );
buf \U$53089 ( \53064 , \53063 );
not \U$53090 ( \53065 , \53064 );
buf \U$53091 ( \53066 , \37534 );
not \U$53092 ( \53067 , \53066 );
or \U$53093 ( \53068 , \53065 , \53067 );
buf \U$53094 ( \53069 , \16071 );
buf \U$53095 ( \53070 , \52709 );
nand \U$53096 ( \53071 , \53069 , \53070 );
buf \U$53097 ( \53072 , \53071 );
buf \U$53098 ( \53073 , \53072 );
nand \U$53099 ( \53074 , \53068 , \53073 );
buf \U$53100 ( \53075 , \53074 );
buf \U$53101 ( \53076 , \53075 );
and \U$53102 ( \53077 , \53059 , \53076 );
and \U$53103 ( \53078 , \53041 , \53058 );
or \U$53104 ( \53079 , \53077 , \53078 );
buf \U$53105 ( \53080 , \53079 );
buf \U$53106 ( \53081 , \53080 );
not \U$53107 ( \53082 , \53081 );
or \U$53108 ( \53083 , \53027 , \53082 );
buf \U$53109 ( \53084 , \53080 );
buf \U$53110 ( \53085 , \53025 );
or \U$53111 ( \53086 , \53084 , \53085 );
buf \U$53112 ( \53087 , RIc0d8a28_43);
buf \U$53113 ( \53088 , RIc0dafa8_123);
xor \U$53114 ( \53089 , \53087 , \53088 );
buf \U$53115 ( \53090 , \53089 );
buf \U$53116 ( \53091 , \53090 );
not \U$53117 ( \53092 , \53091 );
buf \U$53118 ( \53093 , \14982 );
not \U$53119 ( \53094 , \53093 );
or \U$53120 ( \53095 , \53092 , \53094 );
buf \U$53121 ( \53096 , \14278 );
buf \U$53122 ( \53097 , \52505 );
nand \U$53123 ( \53098 , \53096 , \53097 );
buf \U$53124 ( \53099 , \53098 );
buf \U$53125 ( \53100 , \53099 );
nand \U$53126 ( \53101 , \53095 , \53100 );
buf \U$53127 ( \53102 , \53101 );
buf \U$53128 ( \53103 , \53102 );
buf \U$53129 ( \53104 , RIc0daaf8_113);
buf \U$53130 ( \53105 , RIc0d8ed8_53);
xor \U$53131 ( \53106 , \53104 , \53105 );
buf \U$53132 ( \53107 , \53106 );
buf \U$53133 ( \53108 , \53107 );
not \U$53134 ( \53109 , \53108 );
buf \U$53135 ( \53110 , \33224 );
not \U$53136 ( \53111 , \53110 );
or \U$53137 ( \53112 , \53109 , \53111 );
buf \U$53138 ( \53113 , \12410 );
buf \U$53139 ( \53114 , \52694 );
nand \U$53140 ( \53115 , \53113 , \53114 );
buf \U$53141 ( \53116 , \53115 );
buf \U$53142 ( \53117 , \53116 );
nand \U$53143 ( \53118 , \53112 , \53117 );
buf \U$53144 ( \53119 , \53118 );
buf \U$53145 ( \53120 , \53119 );
or \U$53146 ( \53121 , \53103 , \53120 );
buf \U$53147 ( \53122 , \49672 );
not \U$53148 ( \53123 , \53122 );
buf \U$53149 ( \53124 , RIc0daeb8_121);
buf \U$53150 ( \53125 , RIc0d8b18_45);
xnor \U$53151 ( \53126 , \53124 , \53125 );
buf \U$53152 ( \53127 , \53126 );
buf \U$53153 ( \53128 , \53127 );
not \U$53154 ( \53129 , \53128 );
and \U$53155 ( \53130 , \53123 , \53129 );
buf \U$53156 ( \53131 , \52539 );
not \U$53157 ( \53132 , \53131 );
buf \U$53158 ( \53133 , \26373 );
nor \U$53159 ( \53134 , \53132 , \53133 );
buf \U$53160 ( \53135 , \53134 );
buf \U$53161 ( \53136 , \53135 );
nor \U$53162 ( \53137 , \53130 , \53136 );
buf \U$53163 ( \53138 , \53137 );
buf \U$53164 ( \53139 , \53138 );
not \U$53165 ( \53140 , \53139 );
buf \U$53166 ( \53141 , \53140 );
buf \U$53167 ( \53142 , \53141 );
nand \U$53168 ( \53143 , \53121 , \53142 );
buf \U$53169 ( \53144 , \53143 );
buf \U$53170 ( \53145 , \53144 );
buf \U$53171 ( \53146 , \53102 );
buf \U$53172 ( \53147 , \53119 );
nand \U$53173 ( \53148 , \53146 , \53147 );
buf \U$53174 ( \53149 , \53148 );
buf \U$53175 ( \53150 , \53149 );
nand \U$53176 ( \53151 , \53145 , \53150 );
buf \U$53177 ( \53152 , \53151 );
buf \U$53178 ( \53153 , \53152 );
nand \U$53179 ( \53154 , \53086 , \53153 );
buf \U$53180 ( \53155 , \53154 );
buf \U$53181 ( \53156 , \53155 );
nand \U$53182 ( \53157 , \53083 , \53156 );
buf \U$53183 ( \53158 , \53157 );
buf \U$53184 ( \53159 , \53158 );
and \U$53185 ( \53160 , \52968 , \53159 );
and \U$53186 ( \53161 , \52888 , \52967 );
or \U$53187 ( \53162 , \53160 , \53161 );
buf \U$53188 ( \53163 , \53162 );
buf \U$53189 ( \53164 , \53163 );
xor \U$53190 ( \53165 , \52884 , \53164 );
xor \U$53191 ( \53166 , \52693 , \52751 );
xor \U$53192 ( \53167 , \53166 , \52815 );
buf \U$53193 ( \53168 , \53167 );
buf \U$53194 ( \53169 , \53168 );
xor \U$53195 ( \53170 , \52523 , \52589 );
xor \U$53196 ( \53171 , \53170 , \52594 );
buf \U$53197 ( \53172 , \53171 );
buf \U$53198 ( \53173 , \53172 );
xor \U$53199 ( \53174 , \53169 , \53173 );
xor \U$53200 ( \53175 , \52483 , \52500 );
xor \U$53201 ( \53176 , \53175 , \52518 );
buf \U$53202 ( \53177 , \53176 );
buf \U$53203 ( \53178 , \53177 );
buf \U$53204 ( \53179 , \52536 );
not \U$53205 ( \53180 , \53179 );
buf \U$53206 ( \53181 , \52576 );
not \U$53207 ( \53182 , \53181 );
buf \U$53208 ( \53183 , \52554 );
not \U$53209 ( \53184 , \53183 );
or \U$53210 ( \53185 , \53182 , \53184 );
buf \U$53211 ( \53186 , \52554 );
buf \U$53212 ( \53187 , \52576 );
or \U$53213 ( \53188 , \53186 , \53187 );
nand \U$53214 ( \53189 , \53185 , \53188 );
buf \U$53215 ( \53190 , \53189 );
buf \U$53216 ( \53191 , \53190 );
not \U$53217 ( \53192 , \53191 );
or \U$53218 ( \53193 , \53180 , \53192 );
buf \U$53219 ( \53194 , \53190 );
buf \U$53220 ( \53195 , \52536 );
or \U$53221 ( \53196 , \53194 , \53195 );
nand \U$53222 ( \53197 , \53193 , \53196 );
buf \U$53223 ( \53198 , \53197 );
buf \U$53224 ( \53199 , \53198 );
xor \U$53225 ( \53200 , \53178 , \53199 );
xor \U$53226 ( \53201 , \52803 , \52785 );
xor \U$53227 ( \53202 , \53201 , \52768 );
buf \U$53228 ( \53203 , \53202 );
and \U$53229 ( \53204 , \53200 , \53203 );
and \U$53230 ( \53205 , \53178 , \53199 );
or \U$53231 ( \53206 , \53204 , \53205 );
buf \U$53232 ( \53207 , \53206 );
buf \U$53233 ( \53208 , \53207 );
and \U$53234 ( \53209 , \53174 , \53208 );
and \U$53235 ( \53210 , \53169 , \53173 );
or \U$53236 ( \53211 , \53209 , \53210 );
buf \U$53237 ( \53212 , \53211 );
buf \U$53238 ( \53213 , \53212 );
and \U$53239 ( \53214 , \53165 , \53213 );
and \U$53240 ( \53215 , \52884 , \53164 );
or \U$53241 ( \53216 , \53214 , \53215 );
buf \U$53242 ( \53217 , \53216 );
buf \U$53243 ( \53218 , \53217 );
and \U$53244 ( \53219 , \52881 , \53218 );
and \U$53245 ( \53220 , \52876 , \52880 );
or \U$53246 ( \53221 , \53219 , \53220 );
buf \U$53247 ( \53222 , \53221 );
buf \U$53248 ( \53223 , \53222 );
xor \U$53249 ( \53224 , \52051 , \52366 );
xor \U$53250 ( \53225 , \53224 , \52405 );
buf \U$53251 ( \53226 , \53225 );
buf \U$53252 ( \53227 , \53226 );
or \U$53253 ( \53228 , \53223 , \53227 );
xor \U$53254 ( \53229 , \52831 , \52846 );
xor \U$53255 ( \53230 , \53229 , \52850 );
buf \U$53256 ( \53231 , \53230 );
buf \U$53257 ( \53232 , \53231 );
nand \U$53258 ( \53233 , \53228 , \53232 );
buf \U$53259 ( \53234 , \53233 );
buf \U$53260 ( \53235 , \53234 );
buf \U$53261 ( \53236 , \53222 );
buf \U$53262 ( \53237 , \53226 );
nand \U$53263 ( \53238 , \53236 , \53237 );
buf \U$53264 ( \53239 , \53238 );
buf \U$53265 ( \53240 , \53239 );
nand \U$53266 ( \53241 , \53235 , \53240 );
buf \U$53267 ( \53242 , \53241 );
buf \U$53268 ( \53243 , \53242 );
nand \U$53269 ( \53244 , \52872 , \53243 );
buf \U$53270 ( \53245 , \53244 );
not \U$53271 ( \53246 , \53245 );
or \U$53272 ( \53247 , \52868 , \53246 );
buf \U$53273 ( \53248 , \52047 );
not \U$53274 ( \53249 , \53248 );
buf \U$53275 ( \53250 , \53249 );
buf \U$53276 ( \53251 , \53250 );
buf \U$53277 ( \53252 , \52864 );
not \U$53278 ( \53253 , \53252 );
buf \U$53279 ( \53254 , \53253 );
buf \U$53280 ( \53255 , \53254 );
nand \U$53281 ( \53256 , \53251 , \53255 );
buf \U$53282 ( \53257 , \53256 );
nand \U$53283 ( \53258 , \53247 , \53257 );
buf \U$53284 ( \53259 , \53258 );
xor \U$53285 ( \53260 , \50909 , \50704 );
xnor \U$53286 ( \53261 , \53260 , \50936 );
buf \U$53287 ( \53262 , \53261 );
xor \U$53288 ( \53263 , \51667 , \51671 );
and \U$53289 ( \53264 , \53263 , \52023 );
and \U$53290 ( \53265 , \51667 , \51671 );
or \U$53291 ( \53266 , \53264 , \53265 );
buf \U$53292 ( \53267 , \53266 );
buf \U$53293 ( \53268 , \53267 );
xor \U$53294 ( \53269 , \53262 , \53268 );
xor \U$53295 ( \53270 , \51146 , \51150 );
xor \U$53296 ( \53271 , \53270 , \51393 );
buf \U$53297 ( \53272 , \53271 );
buf \U$53298 ( \53273 , \53272 );
xor \U$53299 ( \53274 , \53269 , \53273 );
buf \U$53300 ( \53275 , \53274 );
buf \U$53301 ( \53276 , \53275 );
not \U$53302 ( \53277 , \53276 );
buf \U$53303 ( \53278 , \53277 );
buf \U$53304 ( \53279 , \53278 );
xor \U$53305 ( \53280 , \51497 , \52026 );
and \U$53306 ( \53281 , \53280 , \52045 );
and \U$53307 ( \53282 , \51497 , \52026 );
or \U$53308 ( \53283 , \53281 , \53282 );
buf \U$53309 ( \53284 , \53283 );
buf \U$53310 ( \53285 , \53284 );
not \U$53311 ( \53286 , \53285 );
buf \U$53312 ( \53287 , \53286 );
buf \U$53313 ( \53288 , \53287 );
nand \U$53314 ( \53289 , \53279 , \53288 );
buf \U$53315 ( \53290 , \53289 );
buf \U$53316 ( \53291 , \53290 );
not \U$53317 ( \53292 , \53291 );
buf \U$53318 ( \53293 , \53292 );
buf \U$53319 ( \53294 , \53293 );
or \U$53320 ( \53295 , \53259 , \53294 );
xor \U$53321 ( \53296 , \50981 , \51398 );
xor \U$53322 ( \53297 , \53296 , \51415 );
buf \U$53323 ( \53298 , \53297 );
buf \U$53324 ( \53299 , \53298 );
xor \U$53325 ( \53300 , \53262 , \53268 );
and \U$53326 ( \53301 , \53300 , \53273 );
and \U$53327 ( \53302 , \53262 , \53268 );
or \U$53328 ( \53303 , \53301 , \53302 );
buf \U$53329 ( \53304 , \53303 );
buf \U$53330 ( \53305 , \53304 );
nand \U$53331 ( \53306 , \53299 , \53305 );
buf \U$53332 ( \53307 , \53306 );
buf \U$53333 ( \53308 , \53307 );
buf \U$53334 ( \53309 , \53275 );
buf \U$53335 ( \53310 , \53284 );
nand \U$53336 ( \53311 , \53309 , \53310 );
buf \U$53337 ( \53312 , \53311 );
buf \U$53338 ( \53313 , \53312 );
and \U$53339 ( \53314 , \53308 , \53313 );
buf \U$53340 ( \53315 , \53314 );
buf \U$53341 ( \53316 , \53315 );
nand \U$53342 ( \53317 , \53295 , \53316 );
buf \U$53343 ( \53318 , \53317 );
buf \U$53344 ( \53319 , \53318 );
buf \U$53345 ( \53320 , \53298 );
buf \U$53346 ( \53321 , \53304 );
or \U$53347 ( \53322 , \53320 , \53321 );
buf \U$53348 ( \53323 , \53322 );
buf \U$53349 ( \53324 , \53323 );
nand \U$53350 ( \53325 , \53319 , \53324 );
buf \U$53351 ( \53326 , \53325 );
buf \U$53352 ( \53327 , \53326 );
or \U$53353 ( \53328 , \51493 , \53327 );
buf \U$53354 ( \53329 , \51488 );
not \U$53355 ( \53330 , \53329 );
buf \U$53356 ( \53331 , \51484 );
nand \U$53357 ( \53332 , \53330 , \53331 );
buf \U$53358 ( \53333 , \53332 );
buf \U$53359 ( \53334 , \53333 );
nand \U$53360 ( \53335 , \53328 , \53334 );
buf \U$53361 ( \53336 , \53335 );
buf \U$53362 ( \53337 , \53336 );
buf \U$53363 ( \53338 , \50976 );
buf \U$53364 ( \53339 , \51419 );
not \U$53365 ( \53340 , \53339 );
buf \U$53366 ( \53341 , \51427 );
nor \U$53367 ( \53342 , \53340 , \53341 );
buf \U$53368 ( \53343 , \53342 );
buf \U$53369 ( \53344 , \53343 );
nand \U$53370 ( \53345 , \53338 , \53344 );
buf \U$53371 ( \53346 , \53345 );
buf \U$53372 ( \53347 , \53346 );
buf \U$53373 ( \53348 , \50393 );
not \U$53374 ( \53349 , \53348 );
buf \U$53375 ( \53350 , \50970 );
nand \U$53376 ( \53351 , \53349 , \53350 );
buf \U$53377 ( \53352 , \53351 );
buf \U$53378 ( \53353 , \53352 );
nand \U$53379 ( \53354 , \53347 , \53353 );
buf \U$53380 ( \53355 , \53354 );
buf \U$53381 ( \53356 , \53355 );
buf \U$53382 ( \53357 , \51469 );
nand \U$53383 ( \53358 , \53356 , \53357 );
buf \U$53384 ( \53359 , \53358 );
buf \U$53385 ( \53360 , \53359 );
buf \U$53386 ( \53361 , \51466 );
not \U$53387 ( \53362 , \53361 );
buf \U$53388 ( \53363 , \53362 );
buf \U$53389 ( \53364 , \53363 );
buf \U$53390 ( \53365 , \51447 );
nand \U$53391 ( \53366 , \53364 , \53365 );
buf \U$53392 ( \53367 , \53366 );
buf \U$53393 ( \53368 , \53367 );
and \U$53394 ( \53369 , \53360 , \53368 );
buf \U$53395 ( \53370 , \51489 );
not \U$53396 ( \53371 , \53370 );
buf \U$53397 ( \53372 , \53371 );
buf \U$53398 ( \53373 , \53372 );
nor \U$53399 ( \53374 , \53369 , \53373 );
buf \U$53400 ( \53375 , \53374 );
buf \U$53401 ( \53376 , \53375 );
nor \U$53402 ( \53377 , \53337 , \53376 );
buf \U$53403 ( \53378 , \53377 );
not \U$53404 ( \53379 , \53378 );
buf \U$53405 ( \53380 , \53379 );
not \U$53406 ( \53381 , \53380 );
or \U$53407 ( \53382 , \49376 , \53381 );
not \U$53408 ( \53383 , \48727 );
buf \U$53409 ( \53384 , \48718 );
buf \U$53410 ( \53385 , \48724 );
nand \U$53411 ( \53386 , \53384 , \53385 );
buf \U$53412 ( \53387 , \53386 );
not \U$53413 ( \53388 , \53387 );
nor \U$53414 ( \53389 , \53388 , \47442 );
nor \U$53415 ( \53390 , \53383 , \53389 );
buf \U$53416 ( \53391 , \53390 );
buf \U$53417 ( \53392 , \53387 );
buf \U$53418 ( \53393 , \46971 );
buf \U$53419 ( \53394 , \47439 );
nand \U$53420 ( \53395 , \53393 , \53394 );
buf \U$53421 ( \53396 , \53395 );
buf \U$53422 ( \53397 , \53396 );
and \U$53423 ( \53398 , \53392 , \53397 );
buf \U$53424 ( \53399 , \53398 );
buf \U$53425 ( \53400 , \53399 );
buf \U$53426 ( \53401 , \48013 );
buf \U$53427 ( \53402 , \48734 );
buf \U$53428 ( \53403 , \49368 );
nor \U$53429 ( \53404 , \53402 , \53403 );
buf \U$53430 ( \53405 , \53404 );
buf \U$53431 ( \53406 , \53405 );
nand \U$53432 ( \53407 , \53401 , \53406 );
buf \U$53433 ( \53408 , \53407 );
buf \U$53434 ( \53409 , \53408 );
buf \U$53435 ( \53410 , \48010 );
not \U$53436 ( \53411 , \53410 );
buf \U$53437 ( \53412 , \48002 );
nand \U$53438 ( \53413 , \53411 , \53412 );
buf \U$53439 ( \53414 , \53413 );
buf \U$53440 ( \53415 , \53414 );
nand \U$53441 ( \53416 , \53400 , \53409 , \53415 );
buf \U$53442 ( \53417 , \53416 );
buf \U$53443 ( \53418 , \53417 );
nand \U$53444 ( \53419 , \53391 , \53418 );
buf \U$53445 ( \53420 , \53419 );
buf \U$53446 ( \53421 , \53420 );
nand \U$53447 ( \53422 , \53382 , \53421 );
buf \U$53448 ( \53423 , \53422 );
buf \U$53449 ( \53424 , \53423 );
buf \U$53450 ( \53425 , RIc0d7e70_18);
buf \U$53451 ( \53426 , RIc0db188_127);
xor \U$53452 ( \53427 , \53425 , \53426 );
buf \U$53453 ( \53428 , \53427 );
buf \U$53454 ( \53429 , \53428 );
not \U$53455 ( \53430 , \53429 );
buf \U$53456 ( \53431 , \15609 );
not \U$53457 ( \53432 , \53431 );
or \U$53458 ( \53433 , \53430 , \53432 );
buf \U$53459 ( \53434 , RIc0d7df8_17);
buf \U$53460 ( \53435 , RIc0db188_127);
xor \U$53461 ( \53436 , \53434 , \53435 );
buf \U$53462 ( \53437 , \53436 );
buf \U$53463 ( \53438 , \53437 );
buf \U$53464 ( \53439 , RIc0db200_128);
nand \U$53465 ( \53440 , \53438 , \53439 );
buf \U$53466 ( \53441 , \53440 );
buf \U$53467 ( \53442 , \53441 );
nand \U$53468 ( \53443 , \53433 , \53442 );
buf \U$53469 ( \53444 , \53443 );
buf \U$53470 ( \53445 , \53444 );
buf \U$53471 ( \53446 , RIc0d9fb8_89);
buf \U$53472 ( \53447 , RIc0d9040_56);
xor \U$53473 ( \53448 , \53446 , \53447 );
buf \U$53474 ( \53449 , \53448 );
buf \U$53475 ( \53450 , \53449 );
not \U$53476 ( \53451 , \53450 );
buf \U$53477 ( \53452 , \842 );
not \U$53478 ( \53453 , \53452 );
or \U$53479 ( \53454 , \53451 , \53453 );
buf \U$53480 ( \53455 , \16477 );
buf \U$53481 ( \53456 , RIc0d9fb8_89);
buf \U$53482 ( \53457 , RIc0d8fc8_55);
xor \U$53483 ( \53458 , \53456 , \53457 );
buf \U$53484 ( \53459 , \53458 );
buf \U$53485 ( \53460 , \53459 );
nand \U$53486 ( \53461 , \53455 , \53460 );
buf \U$53487 ( \53462 , \53461 );
buf \U$53488 ( \53463 , \53462 );
nand \U$53489 ( \53464 , \53454 , \53463 );
buf \U$53490 ( \53465 , \53464 );
buf \U$53491 ( \53466 , \53465 );
xor \U$53492 ( \53467 , \53445 , \53466 );
buf \U$53493 ( \53468 , RIc0d8f50_54);
buf \U$53494 ( \53469 , RIc0da0a8_91);
xor \U$53495 ( \53470 , \53468 , \53469 );
buf \U$53496 ( \53471 , \53470 );
buf \U$53497 ( \53472 , \53471 );
not \U$53498 ( \53473 , \53472 );
buf \U$53499 ( \53474 , \1927 );
not \U$53500 ( \53475 , \53474 );
or \U$53501 ( \53476 , \53473 , \53475 );
buf \U$53502 ( \53477 , \1933 );
buf \U$53503 ( \53478 , RIc0d8ed8_53);
buf \U$53504 ( \53479 , RIc0da0a8_91);
xor \U$53505 ( \53480 , \53478 , \53479 );
buf \U$53506 ( \53481 , \53480 );
buf \U$53507 ( \53482 , \53481 );
nand \U$53508 ( \53483 , \53477 , \53482 );
buf \U$53509 ( \53484 , \53483 );
buf \U$53510 ( \53485 , \53484 );
nand \U$53511 ( \53486 , \53476 , \53485 );
buf \U$53512 ( \53487 , \53486 );
buf \U$53513 ( \53488 , \53487 );
xnor \U$53514 ( \53489 , \53467 , \53488 );
buf \U$53515 ( \53490 , \53489 );
buf \U$53516 ( \53491 , RIc0d9bf8_81);
buf \U$53517 ( \53492 , RIc0d9400_64);
xor \U$53518 ( \53493 , \53491 , \53492 );
buf \U$53519 ( \53494 , \53493 );
buf \U$53520 ( \53495 , \53494 );
not \U$53521 ( \53496 , \53495 );
buf \U$53522 ( \53497 , \13075 );
not \U$53523 ( \53498 , \53497 );
or \U$53524 ( \53499 , \53496 , \53498 );
buf \U$53525 ( \53500 , \1078 );
buf \U$53526 ( \53501 , RIc0d9388_63);
buf \U$53527 ( \53502 , RIc0d9bf8_81);
xor \U$53528 ( \53503 , \53501 , \53502 );
buf \U$53529 ( \53504 , \53503 );
buf \U$53530 ( \53505 , \53504 );
nand \U$53531 ( \53506 , \53500 , \53505 );
buf \U$53532 ( \53507 , \53506 );
buf \U$53533 ( \53508 , \53507 );
nand \U$53534 ( \53509 , \53499 , \53508 );
buf \U$53535 ( \53510 , \53509 );
buf \U$53536 ( \53511 , \53510 );
buf \U$53537 ( \53512 , RIc0d8500_32);
buf \U$53538 ( \53513 , RIc0daaf8_113);
xor \U$53539 ( \53514 , \53512 , \53513 );
buf \U$53540 ( \53515 , \53514 );
buf \U$53541 ( \53516 , \53515 );
not \U$53542 ( \53517 , \53516 );
buf \U$53543 ( \53518 , \28413 );
not \U$53544 ( \53519 , \53518 );
or \U$53545 ( \53520 , \53517 , \53519 );
buf \U$53546 ( \53521 , \12410 );
buf \U$53547 ( \53522 , RIc0daaf8_113);
buf \U$53548 ( \53523 , RIc0d8488_31);
xor \U$53549 ( \53524 , \53522 , \53523 );
buf \U$53550 ( \53525 , \53524 );
buf \U$53551 ( \53526 , \53525 );
nand \U$53552 ( \53527 , \53521 , \53526 );
buf \U$53553 ( \53528 , \53527 );
buf \U$53554 ( \53529 , \53528 );
nand \U$53555 ( \53530 , \53520 , \53529 );
buf \U$53556 ( \53531 , \53530 );
buf \U$53557 ( \53532 , \53531 );
xor \U$53558 ( \53533 , \53511 , \53532 );
buf \U$53559 ( \53534 , RIc0d87d0_38);
buf \U$53560 ( \53535 , RIc0da828_107);
xor \U$53561 ( \53536 , \53534 , \53535 );
buf \U$53562 ( \53537 , \53536 );
buf \U$53563 ( \53538 , \53537 );
not \U$53564 ( \53539 , \53538 );
buf \U$53565 ( \53540 , \17595 );
not \U$53566 ( \53541 , \53540 );
or \U$53567 ( \53542 , \53539 , \53541 );
buf \U$53568 ( \53543 , \12342 );
buf \U$53569 ( \53544 , RIc0d8758_37);
buf \U$53570 ( \53545 , RIc0da828_107);
xor \U$53571 ( \53546 , \53544 , \53545 );
buf \U$53572 ( \53547 , \53546 );
buf \U$53573 ( \53548 , \53547 );
nand \U$53574 ( \53549 , \53543 , \53548 );
buf \U$53575 ( \53550 , \53549 );
buf \U$53576 ( \53551 , \53550 );
nand \U$53577 ( \53552 , \53542 , \53551 );
buf \U$53578 ( \53553 , \53552 );
buf \U$53579 ( \53554 , \53553 );
xor \U$53580 ( \53555 , \53533 , \53554 );
buf \U$53581 ( \53556 , \53555 );
buf \U$53582 ( \53557 , \53556 );
not \U$53583 ( \53558 , \53557 );
buf \U$53584 ( \53559 , RIc0d8320_28);
buf \U$53585 ( \53560 , RIc0dacd8_117);
xor \U$53586 ( \53561 , \53559 , \53560 );
buf \U$53587 ( \53562 , \53561 );
buf \U$53588 ( \53563 , \53562 );
not \U$53589 ( \53564 , \53563 );
buf \U$53590 ( \53565 , \13684 );
not \U$53591 ( \53566 , \53565 );
or \U$53592 ( \53567 , \53564 , \53566 );
buf \U$53593 ( \53568 , \12937 );
buf \U$53594 ( \53569 , RIc0d82a8_27);
buf \U$53595 ( \53570 , RIc0dacd8_117);
xor \U$53596 ( \53571 , \53569 , \53570 );
buf \U$53597 ( \53572 , \53571 );
buf \U$53598 ( \53573 , \53572 );
nand \U$53599 ( \53574 , \53568 , \53573 );
buf \U$53600 ( \53575 , \53574 );
buf \U$53601 ( \53576 , \53575 );
nand \U$53602 ( \53577 , \53567 , \53576 );
buf \U$53603 ( \53578 , \53577 );
buf \U$53604 ( \53579 , RIc0d8e60_52);
buf \U$53605 ( \53580 , RIc0da198_93);
xor \U$53606 ( \53581 , \53579 , \53580 );
buf \U$53607 ( \53582 , \53581 );
buf \U$53608 ( \53583 , \53582 );
not \U$53609 ( \53584 , \53583 );
buf \U$53610 ( \53585 , \15995 );
not \U$53611 ( \53586 , \53585 );
or \U$53612 ( \53587 , \53584 , \53586 );
buf \U$53613 ( \53588 , \4008 );
buf \U$53614 ( \53589 , RIc0d8de8_51);
buf \U$53615 ( \53590 , RIc0da198_93);
xor \U$53616 ( \53591 , \53589 , \53590 );
buf \U$53617 ( \53592 , \53591 );
buf \U$53618 ( \53593 , \53592 );
nand \U$53619 ( \53594 , \53588 , \53593 );
buf \U$53620 ( \53595 , \53594 );
buf \U$53621 ( \53596 , \53595 );
nand \U$53622 ( \53597 , \53587 , \53596 );
buf \U$53623 ( \53598 , \53597 );
xor \U$53624 ( \53599 , \53578 , \53598 );
buf \U$53625 ( \53600 , \53599 );
xor \U$53626 ( \53601 , RIc0da648_103, RIc0d89b0_42);
buf \U$53627 ( \53602 , \53601 );
not \U$53628 ( \53603 , \53602 );
buf \U$53629 ( \53604 , \29546 );
not \U$53630 ( \53605 , \53604 );
or \U$53631 ( \53606 , \53603 , \53605 );
buf \U$53632 ( \53607 , \16584 );
xor \U$53633 ( \53608 , RIc0da648_103, RIc0d8938_41);
buf \U$53634 ( \53609 , \53608 );
nand \U$53635 ( \53610 , \53607 , \53609 );
buf \U$53636 ( \53611 , \53610 );
buf \U$53637 ( \53612 , \53611 );
nand \U$53638 ( \53613 , \53606 , \53612 );
buf \U$53639 ( \53614 , \53613 );
buf \U$53640 ( \53615 , \53614 );
not \U$53641 ( \53616 , \53615 );
buf \U$53642 ( \53617 , \53616 );
buf \U$53643 ( \53618 , \53617 );
and \U$53644 ( \53619 , \53600 , \53618 );
not \U$53645 ( \53620 , \53600 );
buf \U$53646 ( \53621 , \53614 );
and \U$53647 ( \53622 , \53620 , \53621 );
nor \U$53648 ( \53623 , \53619 , \53622 );
buf \U$53649 ( \53624 , \53623 );
buf \U$53650 ( \53625 , \53624 );
not \U$53651 ( \53626 , \53625 );
and \U$53652 ( \53627 , \53558 , \53626 );
buf \U$53653 ( \53628 , \53556 );
buf \U$53654 ( \53629 , \53624 );
and \U$53655 ( \53630 , \53628 , \53629 );
nor \U$53656 ( \53631 , \53627 , \53630 );
buf \U$53657 ( \53632 , \53631 );
xor \U$53658 ( \53633 , \53490 , \53632 );
buf \U$53659 ( \53634 , \53633 );
buf \U$53660 ( \53635 , RIc0da918_109);
buf \U$53661 ( \53636 , RIc0d86e0_36);
xor \U$53662 ( \53637 , \53635 , \53636 );
buf \U$53663 ( \53638 , \53637 );
buf \U$53664 ( \53639 , \53638 );
not \U$53665 ( \53640 , \53639 );
buf \U$53666 ( \53641 , \20759 );
not \U$53667 ( \53642 , \53641 );
or \U$53668 ( \53643 , \53640 , \53642 );
buf \U$53669 ( \53644 , \14216 );
buf \U$53670 ( \53645 , RIc0da918_109);
buf \U$53671 ( \53646 , RIc0d8668_35);
xor \U$53672 ( \53647 , \53645 , \53646 );
buf \U$53673 ( \53648 , \53647 );
buf \U$53674 ( \53649 , \53648 );
nand \U$53675 ( \53650 , \53644 , \53649 );
buf \U$53676 ( \53651 , \53650 );
buf \U$53677 ( \53652 , \53651 );
nand \U$53678 ( \53653 , \53643 , \53652 );
buf \U$53679 ( \53654 , \53653 );
buf \U$53680 ( \53655 , \53654 );
buf \U$53681 ( \53656 , RIc0dafa8_123);
buf \U$53682 ( \53657 , RIc0d8050_22);
xor \U$53683 ( \53658 , \53656 , \53657 );
buf \U$53684 ( \53659 , \53658 );
buf \U$53685 ( \53660 , \53659 );
not \U$53686 ( \53661 , \53660 );
buf \U$53687 ( \53662 , \14982 );
not \U$53688 ( \53663 , \53662 );
or \U$53689 ( \53664 , \53661 , \53663 );
xnor \U$53690 ( \53665 , RIc0dafa8_123, RIc0d7fd8_21);
buf \U$53691 ( \53666 , \53665 );
not \U$53692 ( \53667 , \53666 );
buf \U$53693 ( \53668 , \16692 );
nand \U$53694 ( \53669 , \53667 , \53668 );
buf \U$53695 ( \53670 , \53669 );
buf \U$53696 ( \53671 , \53670 );
nand \U$53697 ( \53672 , \53664 , \53671 );
buf \U$53698 ( \53673 , \53672 );
buf \U$53699 ( \53674 , \53673 );
xor \U$53700 ( \53675 , \53655 , \53674 );
buf \U$53701 ( \53676 , RIc0da288_95);
buf \U$53702 ( \53677 , RIc0d8d70_50);
xor \U$53703 ( \53678 , \53676 , \53677 );
buf \U$53704 ( \53679 , \53678 );
buf \U$53705 ( \53680 , \53679 );
not \U$53706 ( \53681 , \53680 );
buf \U$53707 ( \53682 , \330 );
not \U$53708 ( \53683 , \53682 );
or \U$53709 ( \53684 , \53681 , \53683 );
buf \U$53710 ( \53685 , \344 );
buf \U$53711 ( \53686 , RIc0da288_95);
buf \U$53712 ( \53687 , RIc0d8cf8_49);
and \U$53713 ( \53688 , \53686 , \53687 );
not \U$53714 ( \53689 , \53686 );
buf \U$53715 ( \53690 , \22504 );
and \U$53716 ( \53691 , \53689 , \53690 );
nor \U$53717 ( \53692 , \53688 , \53691 );
buf \U$53718 ( \53693 , \53692 );
buf \U$53719 ( \53694 , \53693 );
nand \U$53720 ( \53695 , \53685 , \53694 );
buf \U$53721 ( \53696 , \53695 );
buf \U$53722 ( \53697 , \53696 );
nand \U$53723 ( \53698 , \53684 , \53697 );
buf \U$53724 ( \53699 , \53698 );
buf \U$53725 ( \53700 , \53699 );
xor \U$53726 ( \53701 , \53675 , \53700 );
buf \U$53727 ( \53702 , \53701 );
buf \U$53728 ( \53703 , \53702 );
buf \U$53729 ( \53704 , RIc0da738_105);
buf \U$53730 ( \53705 , RIc0d88c0_40);
xor \U$53731 ( \53706 , \53704 , \53705 );
buf \U$53732 ( \53707 , \53706 );
buf \U$53733 ( \53708 , \53707 );
not \U$53734 ( \53709 , \53708 );
buf \U$53735 ( \53710 , \12736 );
not \U$53736 ( \53711 , \53710 );
or \U$53737 ( \53712 , \53709 , \53711 );
buf \U$53738 ( \53713 , \26301 );
xor \U$53739 ( \53714 , RIc0da738_105, RIc0d8848_39);
buf \U$53740 ( \53715 , \53714 );
nand \U$53741 ( \53716 , \53713 , \53715 );
buf \U$53742 ( \53717 , \53716 );
buf \U$53743 ( \53718 , \53717 );
nand \U$53744 ( \53719 , \53712 , \53718 );
buf \U$53745 ( \53720 , \53719 );
buf \U$53746 ( \53721 , RIc0d8aa0_44);
buf \U$53747 ( \53722 , RIc0da558_101);
xor \U$53748 ( \53723 , \53721 , \53722 );
buf \U$53749 ( \53724 , \53723 );
buf \U$53750 ( \53725 , \53724 );
not \U$53751 ( \53726 , \53725 );
buf \U$53752 ( \53727 , \4042 );
not \U$53753 ( \53728 , \53727 );
or \U$53754 ( \53729 , \53726 , \53728 );
buf \U$53755 ( \53730 , \3515 );
buf \U$53756 ( \53731 , RIc0d8a28_43);
buf \U$53757 ( \53732 , RIc0da558_101);
xor \U$53758 ( \53733 , \53731 , \53732 );
buf \U$53759 ( \53734 , \53733 );
buf \U$53760 ( \53735 , \53734 );
nand \U$53761 ( \53736 , \53730 , \53735 );
buf \U$53762 ( \53737 , \53736 );
buf \U$53763 ( \53738 , \53737 );
nand \U$53764 ( \53739 , \53729 , \53738 );
buf \U$53765 ( \53740 , \53739 );
xor \U$53766 ( \53741 , \53720 , \53740 );
buf \U$53767 ( \53742 , RIc0d8410_30);
buf \U$53768 ( \53743 , RIc0dabe8_115);
xor \U$53769 ( \53744 , \53742 , \53743 );
buf \U$53770 ( \53745 , \53744 );
buf \U$53771 ( \53746 , \53745 );
not \U$53772 ( \53747 , \53746 );
buf \U$53773 ( \53748 , \14186 );
not \U$53774 ( \53749 , \53748 );
or \U$53775 ( \53750 , \53747 , \53749 );
buf \U$53776 ( \53751 , \12303 );
xor \U$53777 ( \53752 , RIc0dabe8_115, RIc0d8398_29);
buf \U$53778 ( \53753 , \53752 );
nand \U$53779 ( \53754 , \53751 , \53753 );
buf \U$53780 ( \53755 , \53754 );
buf \U$53781 ( \53756 , \53755 );
nand \U$53782 ( \53757 , \53750 , \53756 );
buf \U$53783 ( \53758 , \53757 );
xnor \U$53784 ( \53759 , \53741 , \53758 );
buf \U$53785 ( \53760 , \53759 );
and \U$53786 ( \53761 , \53703 , \53760 );
not \U$53787 ( \53762 , \53703 );
buf \U$53788 ( \53763 , \53759 );
not \U$53789 ( \53764 , \53763 );
buf \U$53790 ( \53765 , \53764 );
buf \U$53791 ( \53766 , \53765 );
and \U$53792 ( \53767 , \53762 , \53766 );
nor \U$53793 ( \53768 , \53761 , \53767 );
buf \U$53794 ( \53769 , \53768 );
buf \U$53795 ( \53770 , RIc0d8b90_46);
buf \U$53796 ( \53771 , RIc0da468_99);
xor \U$53797 ( \53772 , \53770 , \53771 );
buf \U$53798 ( \53773 , \53772 );
buf \U$53799 ( \53774 , \53773 );
not \U$53800 ( \53775 , \53774 );
buf \U$53801 ( \53776 , \12578 );
not \U$53802 ( \53777 , \53776 );
or \U$53803 ( \53778 , \53775 , \53777 );
buf \U$53804 ( \53779 , \12584 );
buf \U$53805 ( \53780 , RIc0d8b18_45);
buf \U$53806 ( \53781 , RIc0da468_99);
xor \U$53807 ( \53782 , \53780 , \53781 );
buf \U$53808 ( \53783 , \53782 );
buf \U$53809 ( \53784 , \53783 );
nand \U$53810 ( \53785 , \53779 , \53784 );
buf \U$53811 ( \53786 , \53785 );
buf \U$53812 ( \53787 , \53786 );
nand \U$53813 ( \53788 , \53778 , \53787 );
buf \U$53814 ( \53789 , \53788 );
buf \U$53815 ( \53790 , \53789 );
not \U$53816 ( \53791 , \53790 );
xor \U$53817 ( \53792 , RIc0d9ec8_87, RIc0d9130_58);
buf \U$53818 ( \53793 , \53792 );
not \U$53819 ( \53794 , \53793 );
buf \U$53820 ( \53795 , \14325 );
not \U$53821 ( \53796 , \53795 );
or \U$53822 ( \53797 , \53794 , \53796 );
buf \U$53823 ( \53798 , \14331 );
buf \U$53824 ( \53799 , RIc0d90b8_57);
buf \U$53825 ( \53800 , RIc0d9ec8_87);
xor \U$53826 ( \53801 , \53799 , \53800 );
buf \U$53827 ( \53802 , \53801 );
buf \U$53828 ( \53803 , \53802 );
nand \U$53829 ( \53804 , \53798 , \53803 );
buf \U$53830 ( \53805 , \53804 );
buf \U$53831 ( \53806 , \53805 );
nand \U$53832 ( \53807 , \53797 , \53806 );
buf \U$53833 ( \53808 , \53807 );
buf \U$53834 ( \53809 , \53808 );
not \U$53835 ( \53810 , \53809 );
buf \U$53836 ( \53811 , \53810 );
buf \U$53837 ( \53812 , \53811 );
not \U$53838 ( \53813 , \53812 );
or \U$53839 ( \53814 , \53791 , \53813 );
buf \U$53840 ( \53815 , \53789 );
buf \U$53841 ( \53816 , \53811 );
or \U$53842 ( \53817 , \53815 , \53816 );
nand \U$53843 ( \53818 , \53814 , \53817 );
buf \U$53844 ( \53819 , \53818 );
buf \U$53845 ( \53820 , \53819 );
xor \U$53846 ( \53821 , RIc0d9dd8_85, RIc0d9220_60);
buf \U$53847 ( \53822 , \53821 );
not \U$53848 ( \53823 , \53822 );
buf \U$53849 ( \53824 , \5304 );
not \U$53850 ( \53825 , \53824 );
or \U$53851 ( \53826 , \53823 , \53825 );
buf \U$53852 ( \53827 , RIc0d91a8_59);
buf \U$53853 ( \53828 , RIc0d9dd8_85);
xnor \U$53854 ( \53829 , \53827 , \53828 );
buf \U$53855 ( \53830 , \53829 );
buf \U$53856 ( \53831 , \53830 );
not \U$53857 ( \53832 , \53831 );
buf \U$53858 ( \53833 , \1401 );
nand \U$53859 ( \53834 , \53832 , \53833 );
buf \U$53860 ( \53835 , \53834 );
buf \U$53861 ( \53836 , \53835 );
nand \U$53862 ( \53837 , \53826 , \53836 );
buf \U$53863 ( \53838 , \53837 );
buf \U$53864 ( \53839 , \53838 );
not \U$53865 ( \53840 , \53839 );
buf \U$53866 ( \53841 , \53840 );
buf \U$53867 ( \53842 , \53841 );
and \U$53868 ( \53843 , \53820 , \53842 );
not \U$53869 ( \53844 , \53820 );
buf \U$53870 ( \53845 , \53838 );
and \U$53871 ( \53846 , \53844 , \53845 );
nor \U$53872 ( \53847 , \53843 , \53846 );
buf \U$53873 ( \53848 , \53847 );
buf \U$53874 ( \53849 , \53848 );
not \U$53875 ( \53850 , \53849 );
buf \U$53876 ( \53851 , \53850 );
and \U$53877 ( \53852 , \53769 , \53851 );
not \U$53878 ( \53853 , \53769 );
and \U$53879 ( \53854 , \53853 , \53848 );
or \U$53880 ( \53855 , \53852 , \53854 );
buf \U$53881 ( \53856 , \53855 );
xor \U$53882 ( \53857 , \53634 , \53856 );
buf \U$53883 ( \53858 , RIc0d8b18_45);
buf \U$53884 ( \53859 , RIc0da558_101);
xor \U$53885 ( \53860 , \53858 , \53859 );
buf \U$53886 ( \53861 , \53860 );
buf \U$53887 ( \53862 , \53861 );
not \U$53888 ( \53863 , \53862 );
buf \U$53889 ( \53864 , \3535 );
not \U$53890 ( \53865 , \53864 );
or \U$53891 ( \53866 , \53863 , \53865 );
buf \U$53892 ( \53867 , \4049 );
buf \U$53893 ( \53868 , \53724 );
nand \U$53894 ( \53869 , \53867 , \53868 );
buf \U$53895 ( \53870 , \53869 );
buf \U$53896 ( \53871 , \53870 );
nand \U$53897 ( \53872 , \53866 , \53871 );
buf \U$53898 ( \53873 , \53872 );
xor \U$53899 ( \53874 , RIc0d9ec8_87, RIc0d91a8_59);
buf \U$53900 ( \53875 , \53874 );
not \U$53901 ( \53876 , \53875 );
buf \U$53902 ( \53877 , \618 );
not \U$53903 ( \53878 , \53877 );
or \U$53904 ( \53879 , \53876 , \53878 );
buf \U$53905 ( \53880 , \816 );
buf \U$53906 ( \53881 , \53792 );
nand \U$53907 ( \53882 , \53880 , \53881 );
buf \U$53908 ( \53883 , \53882 );
buf \U$53909 ( \53884 , \53883 );
nand \U$53910 ( \53885 , \53879 , \53884 );
buf \U$53911 ( \53886 , \53885 );
buf \U$53912 ( \53887 , RIc0d8848_39);
buf \U$53913 ( \53888 , RIc0da828_107);
xor \U$53914 ( \53889 , \53887 , \53888 );
buf \U$53915 ( \53890 , \53889 );
buf \U$53916 ( \53891 , \53890 );
not \U$53917 ( \53892 , \53891 );
buf \U$53918 ( \53893 , \21898 );
not \U$53919 ( \53894 , \53893 );
or \U$53920 ( \53895 , \53892 , \53894 );
buf \U$53921 ( \53896 , \12342 );
buf \U$53922 ( \53897 , \53537 );
nand \U$53923 ( \53898 , \53896 , \53897 );
buf \U$53924 ( \53899 , \53898 );
buf \U$53925 ( \53900 , \53899 );
nand \U$53926 ( \53901 , \53895 , \53900 );
buf \U$53927 ( \53902 , \53901 );
xnor \U$53928 ( \53903 , \53886 , \53902 );
not \U$53929 ( \53904 , \53903 );
xor \U$53930 ( \53905 , \53873 , \53904 );
buf \U$53931 ( \53906 , \53905 );
buf \U$53932 ( \53907 , \45089 );
buf \U$53933 ( \53908 , RIc0d8140_24);
buf \U$53934 ( \53909 , RIc0dafa8_123);
xor \U$53935 ( \53910 , \53908 , \53909 );
buf \U$53936 ( \53911 , \53910 );
buf \U$53937 ( \53912 , \53911 );
not \U$53938 ( \53913 , \53912 );
buf \U$53939 ( \53914 , \53913 );
buf \U$53940 ( \53915 , \53914 );
or \U$53941 ( \53916 , \53907 , \53915 );
buf \U$53942 ( \53917 , \16695 );
buf \U$53943 ( \53918 , RIc0dafa8_123);
buf \U$53944 ( \53919 , RIc0d80c8_23);
and \U$53945 ( \53920 , \53918 , \53919 );
not \U$53946 ( \53921 , \53918 );
buf \U$53947 ( \53922 , \7462 );
and \U$53948 ( \53923 , \53921 , \53922 );
nor \U$53949 ( \53924 , \53920 , \53923 );
buf \U$53950 ( \53925 , \53924 );
buf \U$53951 ( \53926 , \53925 );
not \U$53952 ( \53927 , \53926 );
buf \U$53953 ( \53928 , \53927 );
buf \U$53954 ( \53929 , \53928 );
or \U$53955 ( \53930 , \53917 , \53929 );
nand \U$53956 ( \53931 , \53916 , \53930 );
buf \U$53957 ( \53932 , \53931 );
buf \U$53958 ( \53933 , \53932 );
buf \U$53959 ( \53934 , RIc0d9dd8_85);
buf \U$53960 ( \53935 , RIc0d9310_62);
xor \U$53961 ( \53936 , \53934 , \53935 );
buf \U$53962 ( \53937 , \53936 );
buf \U$53963 ( \53938 , \53937 );
not \U$53964 ( \53939 , \53938 );
buf \U$53965 ( \53940 , \1389 );
not \U$53966 ( \53941 , \53940 );
or \U$53967 ( \53942 , \53939 , \53941 );
buf \U$53968 ( \53943 , \1401 );
buf \U$53969 ( \53944 , RIc0d9dd8_85);
buf \U$53970 ( \53945 , RIc0d9298_61);
xor \U$53971 ( \53946 , \53944 , \53945 );
buf \U$53972 ( \53947 , \53946 );
buf \U$53973 ( \53948 , \53947 );
nand \U$53974 ( \53949 , \53943 , \53948 );
buf \U$53975 ( \53950 , \53949 );
buf \U$53976 ( \53951 , \53950 );
nand \U$53977 ( \53952 , \53942 , \53951 );
buf \U$53978 ( \53953 , \53952 );
buf \U$53979 ( \53954 , \53953 );
buf \U$53980 ( \53955 , RIc0d9400_64);
buf \U$53981 ( \53956 , RIc0d9d60_84);
or \U$53982 ( \53957 , \53955 , \53956 );
buf \U$53983 ( \53958 , RIc0d9dd8_85);
nand \U$53984 ( \53959 , \53957 , \53958 );
buf \U$53985 ( \53960 , \53959 );
buf \U$53986 ( \53961 , \53960 );
buf \U$53987 ( \53962 , RIc0d9400_64);
buf \U$53988 ( \53963 , RIc0d9d60_84);
nand \U$53989 ( \53964 , \53962 , \53963 );
buf \U$53990 ( \53965 , \53964 );
buf \U$53991 ( \53966 , \53965 );
buf \U$53992 ( \53967 , RIc0d9ce8_83);
and \U$53993 ( \53968 , \53961 , \53966 , \53967 );
buf \U$53994 ( \53969 , \53968 );
buf \U$53995 ( \53970 , \53969 );
xor \U$53996 ( \53971 , \53954 , \53970 );
buf \U$53997 ( \53972 , \53971 );
buf \U$53998 ( \53973 , \53972 );
xor \U$53999 ( \53974 , \53933 , \53973 );
buf \U$54000 ( \53975 , \48214 );
not \U$54001 ( \53976 , \53975 );
buf \U$54002 ( \53977 , \27591 );
not \U$54003 ( \53978 , \53977 );
or \U$54004 ( \53979 , \53976 , \53978 );
buf \U$54005 ( \53980 , \344 );
buf \U$54006 ( \53981 , RIc0da288_95);
buf \U$54007 ( \53982 , RIc0d8e60_52);
xor \U$54008 ( \53983 , \53981 , \53982 );
buf \U$54009 ( \53984 , \53983 );
buf \U$54010 ( \53985 , \53984 );
nand \U$54011 ( \53986 , \53980 , \53985 );
buf \U$54012 ( \53987 , \53986 );
buf \U$54013 ( \53988 , \53987 );
nand \U$54014 ( \53989 , \53979 , \53988 );
buf \U$54015 ( \53990 , \53989 );
buf \U$54016 ( \53991 , \53990 );
buf \U$54017 ( \53992 , \48197 );
not \U$54018 ( \53993 , \53992 );
buf \U$54019 ( \53994 , \21959 );
not \U$54020 ( \53995 , \53994 );
or \U$54021 ( \53996 , \53993 , \53995 );
buf \U$54022 ( \53997 , \20211 );
buf \U$54023 ( \53998 , RIc0da918_109);
buf \U$54024 ( \53999 , RIc0d87d0_38);
xor \U$54025 ( \54000 , \53998 , \53999 );
buf \U$54026 ( \54001 , \54000 );
buf \U$54027 ( \54002 , \54001 );
nand \U$54028 ( \54003 , \53997 , \54002 );
buf \U$54029 ( \54004 , \54003 );
buf \U$54030 ( \54005 , \54004 );
nand \U$54031 ( \54006 , \53996 , \54005 );
buf \U$54032 ( \54007 , \54006 );
buf \U$54033 ( \54008 , \54007 );
nor \U$54034 ( \54009 , \53991 , \54008 );
buf \U$54035 ( \54010 , \54009 );
buf \U$54036 ( \54011 , \54010 );
buf \U$54037 ( \54012 , \48402 );
not \U$54038 ( \54013 , \54012 );
buf \U$54039 ( \54014 , \2066 );
not \U$54040 ( \54015 , \54014 );
or \U$54041 ( \54016 , \54013 , \54015 );
buf \U$54042 ( \54017 , \2070 );
buf \U$54043 ( \54018 , RIc0d8d70_50);
buf \U$54044 ( \54019 , RIc0da378_97);
xor \U$54045 ( \54020 , \54018 , \54019 );
buf \U$54046 ( \54021 , \54020 );
buf \U$54047 ( \54022 , \54021 );
nand \U$54048 ( \54023 , \54017 , \54022 );
buf \U$54049 ( \54024 , \54023 );
buf \U$54050 ( \54025 , \54024 );
nand \U$54051 ( \54026 , \54016 , \54025 );
buf \U$54052 ( \54027 , \54026 );
buf \U$54053 ( \54028 , \54027 );
not \U$54054 ( \54029 , \54028 );
buf \U$54055 ( \54030 , \54029 );
buf \U$54056 ( \54031 , \54030 );
or \U$54057 ( \54032 , \54011 , \54031 );
buf \U$54058 ( \54033 , \54007 );
buf \U$54059 ( \54034 , \53990 );
nand \U$54060 ( \54035 , \54033 , \54034 );
buf \U$54061 ( \54036 , \54035 );
buf \U$54062 ( \54037 , \54036 );
nand \U$54063 ( \54038 , \54032 , \54037 );
buf \U$54064 ( \54039 , \54038 );
buf \U$54065 ( \54040 , \54039 );
and \U$54066 ( \54041 , \53974 , \54040 );
and \U$54067 ( \54042 , \53933 , \53973 );
or \U$54068 ( \54043 , \54041 , \54042 );
buf \U$54069 ( \54044 , \54043 );
buf \U$54070 ( \54045 , \54044 );
xor \U$54071 ( \54046 , \53906 , \54045 );
buf \U$54072 ( \54047 , \816 );
buf \U$54073 ( \54048 , \606 );
buf \U$54074 ( \54049 , \48578 );
nand \U$54075 ( \54050 , \54048 , \54049 );
buf \U$54076 ( \54051 , \54050 );
buf \U$54077 ( \54052 , \54051 );
or \U$54078 ( \54053 , \54047 , \54052 );
buf \U$54079 ( \54054 , \634 );
not \U$54080 ( \54055 , \54054 );
xor \U$54081 ( \54056 , RIc0d9ec8_87, RIc0d9220_60);
buf \U$54082 ( \54057 , \54056 );
nand \U$54083 ( \54058 , \54055 , \54057 );
buf \U$54084 ( \54059 , \54058 );
buf \U$54085 ( \54060 , \54059 );
nand \U$54086 ( \54061 , \54053 , \54060 );
buf \U$54087 ( \54062 , \54061 );
buf \U$54088 ( \54063 , \54062 );
not \U$54089 ( \54064 , \54063 );
buf \U$54090 ( \54065 , \993 );
buf \U$54091 ( \54066 , RIc0d9400_64);
nand \U$54092 ( \54067 , \54065 , \54066 );
buf \U$54093 ( \54068 , \54067 );
buf \U$54094 ( \54069 , \54068 );
nand \U$54095 ( \54070 , \54064 , \54069 );
buf \U$54096 ( \54071 , \54070 );
buf \U$54097 ( \54072 , \54071 );
not \U$54098 ( \54073 , \54072 );
buf \U$54099 ( \54074 , \48145 );
not \U$54100 ( \54075 , \54074 );
buf \U$54101 ( \54076 , \12529 );
not \U$54102 ( \54077 , \54076 );
or \U$54103 ( \54078 , \54075 , \54077 );
buf \U$54104 ( \54079 , \18312 );
buf \U$54105 ( \54080 , RIc0daa08_111);
buf \U$54106 ( \54081 , RIc0d86e0_36);
xor \U$54107 ( \54082 , \54080 , \54081 );
buf \U$54108 ( \54083 , \54082 );
buf \U$54109 ( \54084 , \54083 );
nand \U$54110 ( \54085 , \54079 , \54084 );
buf \U$54111 ( \54086 , \54085 );
buf \U$54112 ( \54087 , \54086 );
nand \U$54113 ( \54088 , \54078 , \54087 );
buf \U$54114 ( \54089 , \54088 );
buf \U$54115 ( \54090 , \54089 );
not \U$54116 ( \54091 , \54090 );
or \U$54117 ( \54092 , \54073 , \54091 );
buf \U$54118 ( \54093 , \54068 );
not \U$54119 ( \54094 , \54093 );
buf \U$54120 ( \54095 , \54062 );
nand \U$54121 ( \54096 , \54094 , \54095 );
buf \U$54122 ( \54097 , \54096 );
buf \U$54123 ( \54098 , \54097 );
nand \U$54124 ( \54099 , \54092 , \54098 );
buf \U$54125 ( \54100 , \54099 );
buf \U$54126 ( \54101 , \54100 );
not \U$54127 ( \54102 , \54101 );
buf \U$54128 ( \54103 , \48247 );
not \U$54129 ( \54104 , \54103 );
buf \U$54130 ( \54105 , \15609 );
not \U$54131 ( \54106 , \54105 );
or \U$54132 ( \54107 , \54104 , \54106 );
buf \U$54133 ( \54108 , RIc0d7f60_20);
buf \U$54134 ( \54109 , RIc0db188_127);
xnor \U$54135 ( \54110 , \54108 , \54109 );
buf \U$54136 ( \54111 , \54110 );
buf \U$54137 ( \54112 , \54111 );
not \U$54138 ( \54113 , \54112 );
buf \U$54139 ( \54114 , RIc0db200_128);
nand \U$54140 ( \54115 , \54113 , \54114 );
buf \U$54141 ( \54116 , \54115 );
buf \U$54142 ( \54117 , \54116 );
nand \U$54143 ( \54118 , \54107 , \54117 );
buf \U$54144 ( \54119 , \54118 );
buf \U$54145 ( \54120 , \54119 );
buf \U$54146 ( \54121 , \48455 );
not \U$54147 ( \54122 , \54121 );
buf \U$54148 ( \54123 , \842 );
not \U$54149 ( \54124 , \54123 );
or \U$54150 ( \54125 , \54122 , \54124 );
buf \U$54151 ( \54126 , \442 );
buf \U$54152 ( \54127 , RIc0d9130_58);
buf \U$54153 ( \54128 , RIc0d9fb8_89);
xor \U$54154 ( \54129 , \54127 , \54128 );
buf \U$54155 ( \54130 , \54129 );
buf \U$54156 ( \54131 , \54130 );
nand \U$54157 ( \54132 , \54126 , \54131 );
buf \U$54158 ( \54133 , \54132 );
buf \U$54159 ( \54134 , \54133 );
nand \U$54160 ( \54135 , \54125 , \54134 );
buf \U$54161 ( \54136 , \54135 );
buf \U$54162 ( \54137 , \54136 );
xor \U$54163 ( \54138 , \54120 , \54137 );
buf \U$54164 ( \54139 , \48471 );
not \U$54165 ( \54140 , \54139 );
buf \U$54166 ( \54141 , \54140 );
buf \U$54167 ( \54142 , \54141 );
not \U$54168 ( \54143 , \54142 );
buf \U$54169 ( \54144 , \13042 );
not \U$54170 ( \54145 , \54144 );
or \U$54171 ( \54146 , \54143 , \54145 );
buf \U$54172 ( \54147 , \16584 );
buf \U$54173 ( \54148 , RIc0d8aa0_44);
buf \U$54174 ( \54149 , RIc0da648_103);
xor \U$54175 ( \54150 , \54148 , \54149 );
buf \U$54176 ( \54151 , \54150 );
buf \U$54177 ( \54152 , \54151 );
nand \U$54178 ( \54153 , \54147 , \54152 );
buf \U$54179 ( \54154 , \54153 );
buf \U$54180 ( \54155 , \54154 );
nand \U$54181 ( \54156 , \54146 , \54155 );
buf \U$54182 ( \54157 , \54156 );
buf \U$54183 ( \54158 , \54157 );
and \U$54184 ( \54159 , \54138 , \54158 );
and \U$54185 ( \54160 , \54120 , \54137 );
or \U$54186 ( \54161 , \54159 , \54160 );
buf \U$54187 ( \54162 , \54161 );
buf \U$54188 ( \54163 , \54162 );
not \U$54189 ( \54164 , \54163 );
or \U$54190 ( \54165 , \54102 , \54164 );
buf \U$54191 ( \54166 , \54162 );
buf \U$54192 ( \54167 , \54100 );
or \U$54193 ( \54168 , \54166 , \54167 );
buf \U$54194 ( \54169 , \48047 );
not \U$54195 ( \54170 , \54169 );
buf \U$54196 ( \54171 , \3415 );
not \U$54197 ( \54172 , \54171 );
or \U$54198 ( \54173 , \54170 , \54172 );
buf \U$54199 ( \54174 , \481 );
buf \U$54200 ( \54175 , RIc0d8f50_54);
buf \U$54201 ( \54176 , RIc0da198_93);
xor \U$54202 ( \54177 , \54175 , \54176 );
buf \U$54203 ( \54178 , \54177 );
buf \U$54204 ( \54179 , \54178 );
nand \U$54205 ( \54180 , \54174 , \54179 );
buf \U$54206 ( \54181 , \54180 );
buf \U$54207 ( \54182 , \54181 );
nand \U$54208 ( \54183 , \54173 , \54182 );
buf \U$54209 ( \54184 , \54183 );
buf \U$54210 ( \54185 , \54184 );
buf \U$54211 ( \54186 , \48181 );
not \U$54212 ( \54187 , \54186 );
buf \U$54213 ( \54188 , \25542 );
not \U$54214 ( \54189 , \54188 );
or \U$54215 ( \54190 , \54187 , \54189 );
buf \U$54216 ( \54191 , \13005 );
xor \U$54217 ( \54192 , RIc0dadc8_119, RIc0d8320_28);
buf \U$54218 ( \54193 , \54192 );
nand \U$54219 ( \54194 , \54191 , \54193 );
buf \U$54220 ( \54195 , \54194 );
buf \U$54221 ( \54196 , \54195 );
nand \U$54222 ( \54197 , \54190 , \54196 );
buf \U$54223 ( \54198 , \54197 );
buf \U$54224 ( \54199 , \54198 );
xor \U$54225 ( \54200 , \54185 , \54199 );
buf \U$54226 ( \54201 , \15789 );
not \U$54227 ( \54202 , \54201 );
buf \U$54228 ( \54203 , \54202 );
buf \U$54229 ( \54204 , \54203 );
buf \U$54230 ( \54205 , \48079 );
or \U$54231 ( \54206 , \54204 , \54205 );
buf \U$54232 ( \54207 , \22744 );
buf \U$54233 ( \54208 , RIc0db098_125);
buf \U$54234 ( \54209 , RIc0d8050_22);
xnor \U$54235 ( \54210 , \54208 , \54209 );
buf \U$54236 ( \54211 , \54210 );
buf \U$54237 ( \54212 , \54211 );
or \U$54238 ( \54213 , \54207 , \54212 );
nand \U$54239 ( \54214 , \54206 , \54213 );
buf \U$54240 ( \54215 , \54214 );
buf \U$54241 ( \54216 , \54215 );
and \U$54242 ( \54217 , \54200 , \54216 );
and \U$54243 ( \54218 , \54185 , \54199 );
or \U$54244 ( \54219 , \54217 , \54218 );
buf \U$54245 ( \54220 , \54219 );
buf \U$54246 ( \54221 , \54220 );
nand \U$54247 ( \54222 , \54168 , \54221 );
buf \U$54248 ( \54223 , \54222 );
buf \U$54249 ( \54224 , \54223 );
nand \U$54250 ( \54225 , \54165 , \54224 );
buf \U$54251 ( \54226 , \54225 );
buf \U$54252 ( \54227 , \54226 );
and \U$54253 ( \54228 , \54046 , \54227 );
and \U$54254 ( \54229 , \53906 , \54045 );
or \U$54255 ( \54230 , \54228 , \54229 );
buf \U$54256 ( \54231 , \54230 );
buf \U$54257 ( \54232 , \54231 );
xor \U$54258 ( \54233 , \53857 , \54232 );
buf \U$54259 ( \54234 , \54233 );
buf \U$54260 ( \54235 , \54234 );
buf \U$54261 ( \54236 , \48423 );
not \U$54262 ( \54237 , \54236 );
buf \U$54263 ( \54238 , \48395 );
not \U$54264 ( \54239 , \54238 );
or \U$54265 ( \54240 , \54237 , \54239 );
buf \U$54266 ( \54241 , \48395 );
buf \U$54267 ( \54242 , \48423 );
or \U$54268 ( \54243 , \54241 , \54242 );
buf \U$54269 ( \54244 , \48408 );
nand \U$54270 ( \54245 , \54243 , \54244 );
buf \U$54271 ( \54246 , \54245 );
buf \U$54272 ( \54247 , \54246 );
nand \U$54273 ( \54248 , \54240 , \54247 );
buf \U$54274 ( \54249 , \54248 );
buf \U$54275 ( \54250 , \54249 );
not \U$54276 ( \54251 , \54250 );
buf \U$54277 ( \54252 , \48203 );
buf \U$54278 ( \54253 , \48220 );
nor \U$54279 ( \54254 , \54252 , \54253 );
buf \U$54280 ( \54255 , \54254 );
buf \U$54281 ( \54256 , \54255 );
buf \U$54282 ( \54257 , \48190 );
or \U$54283 ( \54258 , \54256 , \54257 );
buf \U$54284 ( \54259 , \48203 );
buf \U$54285 ( \54260 , \48220 );
nand \U$54286 ( \54261 , \54259 , \54260 );
buf \U$54287 ( \54262 , \54261 );
buf \U$54288 ( \54263 , \54262 );
nand \U$54289 ( \54264 , \54258 , \54263 );
buf \U$54290 ( \54265 , \54264 );
buf \U$54291 ( \54266 , \54265 );
not \U$54292 ( \54267 , \54266 );
or \U$54293 ( \54268 , \54251 , \54267 );
buf \U$54294 ( \54269 , \54265 );
buf \U$54295 ( \54270 , \54249 );
or \U$54296 ( \54271 , \54269 , \54270 );
buf \U$54297 ( \54272 , \48526 );
not \U$54298 ( \54273 , \54272 );
buf \U$54299 ( \54274 , \54273 );
buf \U$54300 ( \54275 , \54274 );
not \U$54301 ( \54276 , \54275 );
buf \U$54302 ( \54277 , \48541 );
not \U$54303 ( \54278 , \54277 );
or \U$54304 ( \54279 , \54276 , \54278 );
buf \U$54305 ( \54280 , \48541 );
buf \U$54306 ( \54281 , \54274 );
or \U$54307 ( \54282 , \54280 , \54281 );
buf \U$54308 ( \54283 , \48509 );
nand \U$54309 ( \54284 , \54282 , \54283 );
buf \U$54310 ( \54285 , \54284 );
buf \U$54311 ( \54286 , \54285 );
nand \U$54312 ( \54287 , \54279 , \54286 );
buf \U$54313 ( \54288 , \54287 );
buf \U$54314 ( \54289 , \54288 );
nand \U$54315 ( \54290 , \54271 , \54289 );
buf \U$54316 ( \54291 , \54290 );
buf \U$54317 ( \54292 , \54291 );
nand \U$54318 ( \54293 , \54268 , \54292 );
buf \U$54319 ( \54294 , \54293 );
buf \U$54320 ( \54295 , \54294 );
not \U$54321 ( \54296 , \54295 );
buf \U$54322 ( \54297 , \54296 );
buf \U$54323 ( \54298 , \54297 );
not \U$54324 ( \54299 , \54298 );
xor \U$54325 ( \54300 , \54220 , \54100 );
xnor \U$54326 ( \54301 , \54300 , \54162 );
buf \U$54327 ( \54302 , \54301 );
not \U$54328 ( \54303 , \54302 );
or \U$54329 ( \54304 , \54299 , \54303 );
buf \U$54330 ( \54305 , \48135 );
not \U$54331 ( \54306 , \54305 );
buf \U$54332 ( \54307 , \48154 );
not \U$54333 ( \54308 , \54307 );
or \U$54334 ( \54309 , \54306 , \54308 );
buf \U$54335 ( \54310 , \48168 );
nand \U$54336 ( \54311 , \54309 , \54310 );
buf \U$54337 ( \54312 , \54311 );
buf \U$54338 ( \54313 , \54312 );
buf \U$54339 ( \54314 , \48135 );
not \U$54340 ( \54315 , \54314 );
buf \U$54341 ( \54316 , \48151 );
nand \U$54342 ( \54317 , \54315 , \54316 );
buf \U$54343 ( \54318 , \54317 );
buf \U$54344 ( \54319 , \54318 );
nand \U$54345 ( \54320 , \54313 , \54319 );
buf \U$54346 ( \54321 , \54320 );
buf \U$54347 ( \54322 , \54321 );
buf \U$54348 ( \54323 , \48272 );
buf \U$54349 ( \54324 , \48254 );
or \U$54350 ( \54325 , \54323 , \54324 );
buf \U$54351 ( \54326 , \48290 );
nand \U$54352 ( \54327 , \54325 , \54326 );
buf \U$54353 ( \54328 , \54327 );
buf \U$54354 ( \54329 , \54328 );
buf \U$54355 ( \54330 , \48272 );
buf \U$54356 ( \54331 , \48254 );
nand \U$54357 ( \54332 , \54330 , \54331 );
buf \U$54358 ( \54333 , \54332 );
buf \U$54359 ( \54334 , \54333 );
nand \U$54360 ( \54335 , \54329 , \54334 );
buf \U$54361 ( \54336 , \54335 );
buf \U$54362 ( \54337 , \54336 );
xor \U$54363 ( \54338 , \54322 , \54337 );
xor \U$54364 ( \54339 , \48445 , \48462 );
and \U$54365 ( \54340 , \54339 , \48476 );
and \U$54366 ( \54341 , \48445 , \48462 );
or \U$54367 ( \54342 , \54340 , \54341 );
buf \U$54368 ( \54343 , \54342 );
buf \U$54369 ( \54344 , \54343 );
and \U$54370 ( \54345 , \54338 , \54344 );
and \U$54371 ( \54346 , \54322 , \54337 );
or \U$54372 ( \54347 , \54345 , \54346 );
buf \U$54373 ( \54348 , \54347 );
buf \U$54374 ( \54349 , \54348 );
nand \U$54375 ( \54350 , \54304 , \54349 );
buf \U$54376 ( \54351 , \54350 );
buf \U$54377 ( \54352 , \54351 );
buf \U$54378 ( \54353 , \54301 );
not \U$54379 ( \54354 , \54353 );
buf \U$54380 ( \54355 , \54354 );
buf \U$54381 ( \54356 , \54355 );
buf \U$54382 ( \54357 , \54294 );
nand \U$54383 ( \54358 , \54356 , \54357 );
buf \U$54384 ( \54359 , \54358 );
buf \U$54385 ( \54360 , \54359 );
nand \U$54386 ( \54361 , \54352 , \54360 );
buf \U$54387 ( \54362 , \54361 );
buf \U$54388 ( \54363 , \54362 );
xor \U$54389 ( \54364 , \53906 , \54045 );
xor \U$54390 ( \54365 , \54364 , \54227 );
buf \U$54391 ( \54366 , \54365 );
buf \U$54392 ( \54367 , \54366 );
nor \U$54393 ( \54368 , \54363 , \54367 );
buf \U$54394 ( \54369 , \54368 );
buf \U$54395 ( \54370 , \54369 );
buf \U$54396 ( \54371 , \48053 );
not \U$54397 ( \54372 , \54371 );
buf \U$54398 ( \54373 , \48069 );
not \U$54399 ( \54374 , \54373 );
or \U$54400 ( \54375 , \54372 , \54374 );
buf \U$54401 ( \54376 , \48069 );
buf \U$54402 ( \54377 , \48053 );
or \U$54403 ( \54378 , \54376 , \54377 );
buf \U$54404 ( \54379 , \48087 );
nand \U$54405 ( \54380 , \54378 , \54379 );
buf \U$54406 ( \54381 , \54380 );
buf \U$54407 ( \54382 , \54381 );
nand \U$54408 ( \54383 , \54375 , \54382 );
buf \U$54409 ( \54384 , \54383 );
buf \U$54410 ( \54385 , \54384 );
buf \U$54411 ( \54386 , \54089 );
not \U$54412 ( \54387 , \54386 );
buf \U$54413 ( \54388 , \54062 );
not \U$54414 ( \54389 , \54388 );
buf \U$54415 ( \54390 , \54068 );
not \U$54416 ( \54391 , \54390 );
and \U$54417 ( \54392 , \54389 , \54391 );
buf \U$54418 ( \54393 , \54062 );
buf \U$54419 ( \54394 , \54068 );
and \U$54420 ( \54395 , \54393 , \54394 );
nor \U$54421 ( \54396 , \54392 , \54395 );
buf \U$54422 ( \54397 , \54396 );
buf \U$54423 ( \54398 , \54397 );
not \U$54424 ( \54399 , \54398 );
and \U$54425 ( \54400 , \54387 , \54399 );
buf \U$54426 ( \54401 , \54089 );
buf \U$54427 ( \54402 , \54397 );
and \U$54428 ( \54403 , \54401 , \54402 );
nor \U$54429 ( \54404 , \54400 , \54403 );
buf \U$54430 ( \54405 , \54404 );
buf \U$54431 ( \54406 , \54405 );
not \U$54432 ( \54407 , \54406 );
buf \U$54433 ( \54408 , \54407 );
buf \U$54434 ( \54409 , \54408 );
or \U$54435 ( \54410 , \54385 , \54409 );
buf \U$54436 ( \54411 , \48131 );
not \U$54437 ( \54412 , \54411 );
buf \U$54438 ( \54413 , \18767 );
not \U$54439 ( \54414 , \54413 );
or \U$54440 ( \54415 , \54412 , \54414 );
buf \U$54441 ( \54416 , \921 );
buf \U$54442 ( \54417 , \53937 );
nand \U$54443 ( \54418 , \54416 , \54417 );
buf \U$54444 ( \54419 , \54418 );
buf \U$54445 ( \54420 , \54419 );
nand \U$54446 ( \54421 , \54415 , \54420 );
buf \U$54447 ( \54422 , \54421 );
buf \U$54448 ( \54423 , \54422 );
buf \U$54449 ( \54424 , \48438 );
not \U$54450 ( \54425 , \54424 );
buf \U$54451 ( \54426 , \524 );
not \U$54452 ( \54427 , \54426 );
or \U$54453 ( \54428 , \54425 , \54427 );
buf \U$54454 ( \54429 , \1933 );
buf \U$54455 ( \54430 , RIc0da0a8_91);
buf \U$54456 ( \54431 , RIc0d9040_56);
xor \U$54457 ( \54432 , \54430 , \54431 );
buf \U$54458 ( \54433 , \54432 );
buf \U$54459 ( \54434 , \54433 );
nand \U$54460 ( \54435 , \54429 , \54434 );
buf \U$54461 ( \54436 , \54435 );
buf \U$54462 ( \54437 , \54436 );
nand \U$54463 ( \54438 , \54428 , \54437 );
buf \U$54464 ( \54439 , \54438 );
buf \U$54465 ( \54440 , \54439 );
xor \U$54466 ( \54441 , \54423 , \54440 );
buf \U$54467 ( \54442 , \48162 );
not \U$54468 ( \54443 , \54442 );
buf \U$54469 ( \54444 , \13146 );
not \U$54470 ( \54445 , \54444 );
or \U$54471 ( \54446 , \54443 , \54445 );
buf \U$54472 ( \54447 , RIc0dacd8_117);
buf \U$54473 ( \54448 , RIc0d8410_30);
xnor \U$54474 ( \54449 , \54447 , \54448 );
buf \U$54475 ( \54450 , \54449 );
buf \U$54476 ( \54451 , \54450 );
not \U$54477 ( \54452 , \54451 );
buf \U$54478 ( \54453 , \22356 );
nand \U$54479 ( \54454 , \54452 , \54453 );
buf \U$54480 ( \54455 , \54454 );
buf \U$54481 ( \54456 , \54455 );
nand \U$54482 ( \54457 , \54446 , \54456 );
buf \U$54483 ( \54458 , \54457 );
buf \U$54484 ( \54459 , \54458 );
xor \U$54485 ( \54460 , \54441 , \54459 );
buf \U$54486 ( \54461 , \54460 );
buf \U$54487 ( \54462 , \54461 );
nand \U$54488 ( \54463 , \54410 , \54462 );
buf \U$54489 ( \54464 , \54463 );
buf \U$54490 ( \54465 , \54464 );
buf \U$54491 ( \54466 , \54384 );
buf \U$54492 ( \54467 , \54408 );
nand \U$54493 ( \54468 , \54466 , \54467 );
buf \U$54494 ( \54469 , \54468 );
buf \U$54495 ( \54470 , \54469 );
nand \U$54496 ( \54471 , \54465 , \54470 );
buf \U$54497 ( \54472 , \54471 );
buf \U$54498 ( \54473 , \54472 );
xor \U$54499 ( \54474 , \54185 , \54199 );
xor \U$54500 ( \54475 , \54474 , \54216 );
buf \U$54501 ( \54476 , \54475 );
buf \U$54502 ( \54477 , \54476 );
not \U$54503 ( \54478 , \54477 );
buf \U$54504 ( \54479 , \48284 );
not \U$54505 ( \54480 , \54479 );
buf \U$54506 ( \54481 , \19695 );
not \U$54507 ( \54482 , \54481 );
or \U$54508 ( \54483 , \54480 , \54482 );
buf \U$54509 ( \54484 , \22006 );
xor \U$54510 ( \54485 , RIc0da468_99, RIc0d8c80_48);
buf \U$54511 ( \54486 , \54485 );
nand \U$54512 ( \54487 , \54484 , \54486 );
buf \U$54513 ( \54488 , \54487 );
buf \U$54514 ( \54489 , \54488 );
nand \U$54515 ( \54490 , \54483 , \54489 );
buf \U$54516 ( \54491 , \54490 );
buf \U$54517 ( \54492 , \54491 );
buf \U$54518 ( \54493 , \48063 );
not \U$54519 ( \54494 , \54493 );
buf \U$54520 ( \54495 , \15644 );
not \U$54521 ( \54496 , \54495 );
or \U$54522 ( \54497 , \54494 , \54496 );
buf \U$54523 ( \54498 , \12744 );
buf \U$54524 ( \54499 , RIc0da738_105);
buf \U$54525 ( \54500 , RIc0d89b0_42);
xor \U$54526 ( \54501 , \54499 , \54500 );
buf \U$54527 ( \54502 , \54501 );
buf \U$54528 ( \54503 , \54502 );
nand \U$54529 ( \54504 , \54498 , \54503 );
buf \U$54530 ( \54505 , \54504 );
buf \U$54531 ( \54506 , \54505 );
nand \U$54532 ( \54507 , \54497 , \54506 );
buf \U$54533 ( \54508 , \54507 );
buf \U$54534 ( \54509 , \54508 );
xor \U$54535 ( \54510 , \54492 , \54509 );
buf \U$54536 ( \54511 , \14888 );
buf \U$54537 ( \54512 , \48264 );
or \U$54538 ( \54513 , \54511 , \54512 );
buf \U$54539 ( \54514 , \34244 );
buf \U$54540 ( \54515 , RIc0daaf8_113);
buf \U$54541 ( \54516 , RIc0d85f0_34);
xor \U$54542 ( \54517 , \54515 , \54516 );
buf \U$54543 ( \54518 , \54517 );
buf \U$54544 ( \54519 , \54518 );
not \U$54545 ( \54520 , \54519 );
buf \U$54546 ( \54521 , \54520 );
buf \U$54547 ( \54522 , \54521 );
or \U$54548 ( \54523 , \54514 , \54522 );
nand \U$54549 ( \54524 , \54513 , \54523 );
buf \U$54550 ( \54525 , \54524 );
buf \U$54551 ( \54526 , \54525 );
xor \U$54552 ( \54527 , \54510 , \54526 );
buf \U$54553 ( \54528 , \54527 );
buf \U$54554 ( \54529 , \54528 );
not \U$54555 ( \54530 , \54529 );
or \U$54556 ( \54531 , \54478 , \54530 );
buf \U$54557 ( \54532 , \54528 );
buf \U$54558 ( \54533 , \54476 );
or \U$54559 ( \54534 , \54532 , \54533 );
xor \U$54560 ( \54535 , \54030 , \54007 );
not \U$54561 ( \54536 , \53990 );
xor \U$54562 ( \54537 , \54535 , \54536 );
buf \U$54563 ( \54538 , \54537 );
nand \U$54564 ( \54539 , \54534 , \54538 );
buf \U$54565 ( \54540 , \54539 );
buf \U$54566 ( \54541 , \54540 );
nand \U$54567 ( \54542 , \54531 , \54541 );
buf \U$54568 ( \54543 , \54542 );
buf \U$54569 ( \54544 , \54543 );
xor \U$54570 ( \54545 , \54473 , \54544 );
buf \U$54571 ( \54546 , \48389 );
not \U$54572 ( \54547 , \54546 );
buf \U$54573 ( \54548 , \17089 );
not \U$54574 ( \54549 , \54548 );
or \U$54575 ( \54550 , \54547 , \54549 );
buf \U$54576 ( \54551 , \13314 );
xor \U$54577 ( \54552 , RIc0daeb8_121, RIc0d8230_26);
buf \U$54578 ( \54553 , \54552 );
nand \U$54579 ( \54554 , \54551 , \54553 );
buf \U$54580 ( \54555 , \54554 );
buf \U$54581 ( \54556 , \54555 );
nand \U$54582 ( \54557 , \54550 , \54556 );
buf \U$54583 ( \54558 , \54557 );
buf \U$54584 ( \54559 , \54558 );
not \U$54585 ( \54560 , \54559 );
buf \U$54586 ( \54561 , \48417 );
not \U$54587 ( \54562 , \54561 );
buf \U$54588 ( \54563 , \22631 );
not \U$54589 ( \54564 , \54563 );
or \U$54590 ( \54565 , \54562 , \54564 );
buf \U$54591 ( \54566 , \15550 );
buf \U$54592 ( \54567 , RIc0da558_101);
buf \U$54593 ( \54568 , RIc0d8b90_46);
xor \U$54594 ( \54569 , \54567 , \54568 );
buf \U$54595 ( \54570 , \54569 );
buf \U$54596 ( \54571 , \54570 );
nand \U$54597 ( \54572 , \54566 , \54571 );
buf \U$54598 ( \54573 , \54572 );
buf \U$54599 ( \54574 , \54573 );
nand \U$54600 ( \54575 , \54565 , \54574 );
buf \U$54601 ( \54576 , \54575 );
buf \U$54602 ( \54577 , \54576 );
not \U$54603 ( \54578 , \54577 );
or \U$54604 ( \54579 , \54560 , \54578 );
buf \U$54605 ( \54580 , \54576 );
buf \U$54606 ( \54581 , \54558 );
or \U$54607 ( \54582 , \54580 , \54581 );
buf \U$54608 ( \54583 , \48520 );
not \U$54609 ( \54584 , \54583 );
buf \U$54610 ( \54585 , \54584 );
buf \U$54611 ( \54586 , \54585 );
not \U$54612 ( \54587 , \54586 );
buf \U$54613 ( \54588 , \27743 );
not \U$54614 ( \54589 , \54588 );
or \U$54615 ( \54590 , \54587 , \54589 );
buf \U$54616 ( \54591 , \12303 );
buf \U$54617 ( \54592 , RIc0dabe8_115);
buf \U$54618 ( \54593 , RIc0d8500_32);
xor \U$54619 ( \54594 , \54592 , \54593 );
buf \U$54620 ( \54595 , \54594 );
buf \U$54621 ( \54596 , \54595 );
nand \U$54622 ( \54597 , \54591 , \54596 );
buf \U$54623 ( \54598 , \54597 );
buf \U$54624 ( \54599 , \54598 );
nand \U$54625 ( \54600 , \54590 , \54599 );
buf \U$54626 ( \54601 , \54600 );
buf \U$54627 ( \54602 , \54601 );
nand \U$54628 ( \54603 , \54582 , \54602 );
buf \U$54629 ( \54604 , \54603 );
buf \U$54630 ( \54605 , \54604 );
nand \U$54631 ( \54606 , \54579 , \54605 );
buf \U$54632 ( \54607 , \54606 );
xor \U$54633 ( \54608 , \54492 , \54509 );
and \U$54634 ( \54609 , \54608 , \54526 );
and \U$54635 ( \54610 , \54492 , \54509 );
or \U$54636 ( \54611 , \54609 , \54610 );
buf \U$54637 ( \54612 , \54611 );
xor \U$54638 ( \54613 , \54607 , \54612 );
xor \U$54639 ( \54614 , \54423 , \54440 );
and \U$54640 ( \54615 , \54614 , \54459 );
and \U$54641 ( \54616 , \54423 , \54440 );
or \U$54642 ( \54617 , \54615 , \54616 );
buf \U$54643 ( \54618 , \54617 );
xor \U$54644 ( \54619 , \54613 , \54618 );
buf \U$54645 ( \54620 , \54619 );
and \U$54646 ( \54621 , \54545 , \54620 );
and \U$54647 ( \54622 , \54473 , \54544 );
or \U$54648 ( \54623 , \54621 , \54622 );
buf \U$54649 ( \54624 , \54623 );
buf \U$54650 ( \54625 , \54624 );
not \U$54651 ( \54626 , \54625 );
buf \U$54652 ( \54627 , \54626 );
buf \U$54653 ( \54628 , \54627 );
or \U$54654 ( \54629 , \54370 , \54628 );
buf \U$54655 ( \54630 , \54362 );
buf \U$54656 ( \54631 , \54366 );
nand \U$54657 ( \54632 , \54630 , \54631 );
buf \U$54658 ( \54633 , \54632 );
buf \U$54659 ( \54634 , \54633 );
nand \U$54660 ( \54635 , \54629 , \54634 );
buf \U$54661 ( \54636 , \54635 );
buf \U$54662 ( \54637 , \54636 );
xor \U$54663 ( \54638 , \54235 , \54637 );
buf \U$54664 ( \54639 , \54595 );
not \U$54665 ( \54640 , \54639 );
buf \U$54666 ( \54641 , \14186 );
not \U$54667 ( \54642 , \54641 );
or \U$54668 ( \54643 , \54640 , \54642 );
buf \U$54669 ( \54644 , \12303 );
buf \U$54670 ( \54645 , RIc0d8488_31);
buf \U$54671 ( \54646 , RIc0dabe8_115);
xor \U$54672 ( \54647 , \54645 , \54646 );
buf \U$54673 ( \54648 , \54647 );
buf \U$54674 ( \54649 , \54648 );
nand \U$54675 ( \54650 , \54644 , \54649 );
buf \U$54676 ( \54651 , \54650 );
buf \U$54677 ( \54652 , \54651 );
nand \U$54678 ( \54653 , \54643 , \54652 );
buf \U$54679 ( \54654 , \54653 );
buf \U$54680 ( \54655 , \54654 );
not \U$54681 ( \54656 , \54655 );
buf \U$54682 ( \54657 , \54656 );
buf \U$54683 ( \54658 , \54657 );
not \U$54684 ( \54659 , \54658 );
buf \U$54685 ( \54660 , \54001 );
not \U$54686 ( \54661 , \54660 );
buf \U$54687 ( \54662 , \20759 );
not \U$54688 ( \54663 , \54662 );
or \U$54689 ( \54664 , \54661 , \54663 );
buf \U$54690 ( \54665 , \20211 );
buf \U$54691 ( \54666 , RIc0da918_109);
buf \U$54692 ( \54667 , RIc0d8758_37);
xor \U$54693 ( \54668 , \54666 , \54667 );
buf \U$54694 ( \54669 , \54668 );
buf \U$54695 ( \54670 , \54669 );
nand \U$54696 ( \54671 , \54665 , \54670 );
buf \U$54697 ( \54672 , \54671 );
buf \U$54698 ( \54673 , \54672 );
nand \U$54699 ( \54674 , \54664 , \54673 );
buf \U$54700 ( \54675 , \54674 );
buf \U$54701 ( \54676 , \54675 );
not \U$54702 ( \54677 , \54676 );
buf \U$54703 ( \54678 , \54677 );
buf \U$54704 ( \54679 , \54678 );
not \U$54705 ( \54680 , \54679 );
or \U$54706 ( \54681 , \54659 , \54680 );
buf \U$54707 ( \54682 , RIc0d9ce8_83);
buf \U$54708 ( \54683 , RIc0d9400_64);
and \U$54709 ( \54684 , \54682 , \54683 );
not \U$54710 ( \54685 , \54682 );
buf \U$54711 ( \54686 , \43843 );
and \U$54712 ( \54687 , \54685 , \54686 );
nor \U$54713 ( \54688 , \54684 , \54687 );
buf \U$54714 ( \54689 , \54688 );
buf \U$54715 ( \54690 , \54689 );
not \U$54716 ( \54691 , \54690 );
buf \U$54717 ( \54692 , \2088 );
not \U$54718 ( \54693 , \54692 );
or \U$54719 ( \54694 , \54691 , \54693 );
buf \U$54720 ( \54695 , \993 );
buf \U$54721 ( \54696 , RIc0d9388_63);
buf \U$54722 ( \54697 , RIc0d9ce8_83);
xor \U$54723 ( \54698 , \54696 , \54697 );
buf \U$54724 ( \54699 , \54698 );
buf \U$54725 ( \54700 , \54699 );
nand \U$54726 ( \54701 , \54695 , \54700 );
buf \U$54727 ( \54702 , \54701 );
buf \U$54728 ( \54703 , \54702 );
nand \U$54729 ( \54704 , \54694 , \54703 );
buf \U$54730 ( \54705 , \54704 );
buf \U$54731 ( \54706 , \54705 );
nand \U$54732 ( \54707 , \54681 , \54706 );
buf \U$54733 ( \54708 , \54707 );
buf \U$54734 ( \54709 , \54708 );
buf \U$54735 ( \54710 , \54675 );
buf \U$54736 ( \54711 , \54654 );
nand \U$54737 ( \54712 , \54710 , \54711 );
buf \U$54738 ( \54713 , \54712 );
buf \U$54739 ( \54714 , \54713 );
nand \U$54740 ( \54715 , \54709 , \54714 );
buf \U$54741 ( \54716 , \54715 );
xor \U$54742 ( \54717 , RIc0da378_97, RIc0d8cf8_49);
buf \U$54743 ( \54718 , \54717 );
not \U$54744 ( \54719 , \54718 );
buf \U$54745 ( \54720 , \734 );
not \U$54746 ( \54721 , \54720 );
or \U$54747 ( \54722 , \54719 , \54721 );
buf \U$54748 ( \54723 , \737 );
buf \U$54749 ( \54724 , \54021 );
buf \U$54750 ( \54725 , \745 );
nand \U$54751 ( \54726 , \54723 , \54724 , \54725 );
buf \U$54752 ( \54727 , \54726 );
buf \U$54753 ( \54728 , \54727 );
nand \U$54754 ( \54729 , \54722 , \54728 );
buf \U$54755 ( \54730 , \54729 );
buf \U$54756 ( \54731 , \54730 );
not \U$54757 ( \54732 , \54731 );
buf \U$54758 ( \54733 , RIc0d88c0_40);
buf \U$54759 ( \54734 , RIc0da828_107);
xor \U$54760 ( \54735 , \54733 , \54734 );
buf \U$54761 ( \54736 , \54735 );
buf \U$54762 ( \54737 , \54736 );
not \U$54763 ( \54738 , \54737 );
buf \U$54764 ( \54739 , \12334 );
not \U$54765 ( \54740 , \54739 );
or \U$54766 ( \54741 , \54738 , \54740 );
buf \U$54767 ( \54742 , \16071 );
buf \U$54768 ( \54743 , \53890 );
nand \U$54769 ( \54744 , \54742 , \54743 );
buf \U$54770 ( \54745 , \54744 );
buf \U$54771 ( \54746 , \54745 );
nand \U$54772 ( \54747 , \54741 , \54746 );
buf \U$54773 ( \54748 , \54747 );
buf \U$54774 ( \54749 , \54748 );
not \U$54775 ( \54750 , \54749 );
or \U$54776 ( \54751 , \54732 , \54750 );
buf \U$54777 ( \54752 , \54748 );
buf \U$54778 ( \54753 , \54730 );
or \U$54779 ( \54754 , \54752 , \54753 );
buf \U$54780 ( \54755 , \54083 );
not \U$54781 ( \54756 , \54755 );
buf \U$54782 ( \54757 , \12529 );
not \U$54783 ( \54758 , \54757 );
or \U$54784 ( \54759 , \54756 , \54758 );
buf \U$54785 ( \54760 , RIc0d8668_35);
buf \U$54786 ( \54761 , RIc0daa08_111);
xnor \U$54787 ( \54762 , \54760 , \54761 );
buf \U$54788 ( \54763 , \54762 );
buf \U$54789 ( \54764 , \54763 );
not \U$54790 ( \54765 , \54764 );
buf \U$54791 ( \54766 , \15864 );
nand \U$54792 ( \54767 , \54765 , \54766 );
buf \U$54793 ( \54768 , \54767 );
buf \U$54794 ( \54769 , \54768 );
nand \U$54795 ( \54770 , \54759 , \54769 );
buf \U$54796 ( \54771 , \54770 );
buf \U$54797 ( \54772 , \54771 );
nand \U$54798 ( \54773 , \54754 , \54772 );
buf \U$54799 ( \54774 , \54773 );
buf \U$54800 ( \54775 , \54774 );
nand \U$54801 ( \54776 , \54751 , \54775 );
buf \U$54802 ( \54777 , \54776 );
buf \U$54803 ( \54778 , \54777 );
buf \U$54804 ( \54779 , \53953 );
buf \U$54805 ( \54780 , \53969 );
nand \U$54806 ( \54781 , \54779 , \54780 );
buf \U$54807 ( \54782 , \54781 );
buf \U$54808 ( \54783 , \54782 );
and \U$54809 ( \54784 , \54778 , \54783 );
not \U$54810 ( \54785 , \54778 );
buf \U$54811 ( \54786 , \54782 );
not \U$54812 ( \54787 , \54786 );
buf \U$54813 ( \54788 , \54787 );
buf \U$54814 ( \54789 , \54788 );
and \U$54815 ( \54790 , \54785 , \54789 );
nor \U$54816 ( \54791 , \54784 , \54790 );
buf \U$54817 ( \54792 , \54791 );
xnor \U$54818 ( \54793 , \54716 , \54792 );
buf \U$54819 ( \54794 , \54793 );
buf \U$54820 ( \54795 , \54518 );
not \U$54821 ( \54796 , \54795 );
buf \U$54822 ( \54797 , \14891 );
not \U$54823 ( \54798 , \54797 );
or \U$54824 ( \54799 , \54796 , \54798 );
buf \U$54825 ( \54800 , \12410 );
buf \U$54826 ( \54801 , RIc0d8578_33);
buf \U$54827 ( \54802 , RIc0daaf8_113);
xor \U$54828 ( \54803 , \54801 , \54802 );
buf \U$54829 ( \54804 , \54803 );
buf \U$54830 ( \54805 , \54804 );
nand \U$54831 ( \54806 , \54800 , \54805 );
buf \U$54832 ( \54807 , \54806 );
buf \U$54833 ( \54808 , \54807 );
nand \U$54834 ( \54809 , \54799 , \54808 );
buf \U$54835 ( \54810 , \54809 );
buf \U$54836 ( \54811 , \54810 );
buf \U$54837 ( \54812 , \54552 );
not \U$54838 ( \54813 , \54812 );
buf \U$54839 ( \54814 , \16382 );
not \U$54840 ( \54815 , \54814 );
or \U$54841 ( \54816 , \54813 , \54815 );
buf \U$54842 ( \54817 , \16386 );
buf \U$54843 ( \54818 , RIc0daeb8_121);
buf \U$54844 ( \54819 , RIc0d81b8_25);
xor \U$54845 ( \54820 , \54818 , \54819 );
buf \U$54846 ( \54821 , \54820 );
buf \U$54847 ( \54822 , \54821 );
nand \U$54848 ( \54823 , \54817 , \54822 );
buf \U$54849 ( \54824 , \54823 );
buf \U$54850 ( \54825 , \54824 );
nand \U$54851 ( \54826 , \54816 , \54825 );
buf \U$54852 ( \54827 , \54826 );
buf \U$54853 ( \54828 , \54827 );
xor \U$54854 ( \54829 , \54811 , \54828 );
buf \U$54855 ( \54830 , \2207 );
buf \U$54856 ( \54831 , \54485 );
not \U$54857 ( \54832 , \54831 );
buf \U$54858 ( \54833 , \54832 );
buf \U$54859 ( \54834 , \54833 );
or \U$54860 ( \54835 , \54830 , \54834 );
buf \U$54861 ( \54836 , \2199 );
xor \U$54862 ( \54837 , RIc0da468_99, RIc0d8c08_47);
buf \U$54863 ( \54838 , \54837 );
not \U$54864 ( \54839 , \54838 );
buf \U$54865 ( \54840 , \54839 );
buf \U$54866 ( \54841 , \54840 );
or \U$54867 ( \54842 , \54836 , \54841 );
nand \U$54868 ( \54843 , \54835 , \54842 );
buf \U$54869 ( \54844 , \54843 );
buf \U$54870 ( \54845 , \54844 );
xor \U$54871 ( \54846 , \54829 , \54845 );
buf \U$54872 ( \54847 , \54846 );
buf \U$54873 ( \54848 , \54847 );
not \U$54874 ( \54849 , \54848 );
buf \U$54875 ( \54850 , \54654 );
not \U$54876 ( \54851 , \54850 );
buf \U$54877 ( \54852 , \54678 );
not \U$54878 ( \54853 , \54852 );
or \U$54879 ( \54854 , \54851 , \54853 );
buf \U$54880 ( \54855 , \54657 );
buf \U$54881 ( \54856 , \54675 );
nand \U$54882 ( \54857 , \54855 , \54856 );
buf \U$54883 ( \54858 , \54857 );
buf \U$54884 ( \54859 , \54858 );
nand \U$54885 ( \54860 , \54854 , \54859 );
buf \U$54886 ( \54861 , \54860 );
buf \U$54887 ( \54862 , \54861 );
buf \U$54888 ( \54863 , \54705 );
not \U$54889 ( \54864 , \54863 );
buf \U$54890 ( \54865 , \54864 );
buf \U$54891 ( \54866 , \54865 );
and \U$54892 ( \54867 , \54862 , \54866 );
not \U$54893 ( \54868 , \54862 );
buf \U$54894 ( \54869 , \54705 );
and \U$54895 ( \54870 , \54868 , \54869 );
nor \U$54896 ( \54871 , \54867 , \54870 );
buf \U$54897 ( \54872 , \54871 );
buf \U$54898 ( \54873 , \54872 );
not \U$54899 ( \54874 , \54873 );
buf \U$54900 ( \54875 , \54874 );
buf \U$54901 ( \54876 , \54875 );
not \U$54902 ( \54877 , \54876 );
or \U$54903 ( \54878 , \54849 , \54877 );
buf \U$54904 ( \54879 , \54875 );
buf \U$54905 ( \54880 , \54847 );
or \U$54906 ( \54881 , \54879 , \54880 );
buf \U$54907 ( \54882 , \54433 );
not \U$54908 ( \54883 , \54882 );
buf \U$54909 ( \54884 , \704 );
not \U$54910 ( \54885 , \54884 );
or \U$54911 ( \54886 , \54883 , \54885 );
buf \U$54912 ( \54887 , \1933 );
buf \U$54913 ( \54888 , RIc0d8fc8_55);
buf \U$54914 ( \54889 , RIc0da0a8_91);
xor \U$54915 ( \54890 , \54888 , \54889 );
buf \U$54916 ( \54891 , \54890 );
buf \U$54917 ( \54892 , \54891 );
nand \U$54918 ( \54893 , \54887 , \54892 );
buf \U$54919 ( \54894 , \54893 );
buf \U$54920 ( \54895 , \54894 );
nand \U$54921 ( \54896 , \54886 , \54895 );
buf \U$54922 ( \54897 , \54896 );
buf \U$54923 ( \54898 , \54897 );
buf \U$54924 ( \54899 , \54502 );
not \U$54925 ( \54900 , \54899 );
buf \U$54926 ( \54901 , \15644 );
not \U$54927 ( \54902 , \54901 );
or \U$54928 ( \54903 , \54900 , \54902 );
buf \U$54929 ( \54904 , \12744 );
buf \U$54930 ( \54905 , RIc0da738_105);
buf \U$54931 ( \54906 , RIc0d8938_41);
xor \U$54932 ( \54907 , \54905 , \54906 );
buf \U$54933 ( \54908 , \54907 );
buf \U$54934 ( \54909 , \54908 );
nand \U$54935 ( \54910 , \54904 , \54909 );
buf \U$54936 ( \54911 , \54910 );
buf \U$54937 ( \54912 , \54911 );
nand \U$54938 ( \54913 , \54903 , \54912 );
buf \U$54939 ( \54914 , \54913 );
buf \U$54940 ( \54915 , \54914 );
xor \U$54941 ( \54916 , \54898 , \54915 );
buf \U$54942 ( \54917 , \54178 );
not \U$54943 ( \54918 , \54917 );
buf \U$54944 ( \54919 , \889 );
not \U$54945 ( \54920 , \54919 );
or \U$54946 ( \54921 , \54918 , \54920 );
buf \U$54947 ( \54922 , \4008 );
buf \U$54948 ( \54923 , RIc0da198_93);
buf \U$54949 ( \54924 , RIc0d8ed8_53);
xor \U$54950 ( \54925 , \54923 , \54924 );
buf \U$54951 ( \54926 , \54925 );
buf \U$54952 ( \54927 , \54926 );
nand \U$54953 ( \54928 , \54922 , \54927 );
buf \U$54954 ( \54929 , \54928 );
buf \U$54955 ( \54930 , \54929 );
nand \U$54956 ( \54931 , \54921 , \54930 );
buf \U$54957 ( \54932 , \54931 );
buf \U$54958 ( \54933 , \54932 );
xor \U$54959 ( \54934 , \54916 , \54933 );
buf \U$54960 ( \54935 , \54934 );
buf \U$54961 ( \54936 , \54935 );
nand \U$54962 ( \54937 , \54881 , \54936 );
buf \U$54963 ( \54938 , \54937 );
buf \U$54964 ( \54939 , \54938 );
nand \U$54965 ( \54940 , \54878 , \54939 );
buf \U$54966 ( \54941 , \54940 );
buf \U$54967 ( \54942 , \54941 );
xor \U$54968 ( \54943 , \54794 , \54942 );
xor \U$54969 ( \54944 , RIc0da648_103, RIc0d8a28_43);
buf \U$54970 ( \54945 , \54944 );
not \U$54971 ( \54946 , \54945 );
buf \U$54972 ( \54947 , \15403 );
not \U$54973 ( \54948 , \54947 );
or \U$54974 ( \54949 , \54946 , \54948 );
buf \U$54975 ( \54950 , \4475 );
buf \U$54976 ( \54951 , \54151 );
buf \U$54977 ( \54952 , \4479 );
nand \U$54978 ( \54953 , \54950 , \54951 , \54952 );
buf \U$54979 ( \54954 , \54953 );
buf \U$54980 ( \54955 , \54954 );
nand \U$54981 ( \54956 , \54949 , \54955 );
buf \U$54982 ( \54957 , \54956 );
buf \U$54983 ( \54958 , \54957 );
xor \U$54984 ( \54959 , RIc0db188_127, RIc0d7ee8_19);
not \U$54985 ( \54960 , \54959 );
not \U$54986 ( \54961 , RIc0db200_128);
or \U$54987 ( \54962 , \54960 , \54961 );
or \U$54988 ( \54963 , \18008 , \54111 );
nand \U$54989 ( \54964 , \54962 , \54963 );
buf \U$54990 ( \54965 , \54964 );
xor \U$54991 ( \54966 , \54958 , \54965 );
buf \U$54992 ( \54967 , \44882 );
buf \U$54993 ( \54968 , \54450 );
or \U$54994 ( \54969 , \54967 , \54968 );
buf \U$54995 ( \54970 , \44894 );
buf \U$54996 ( \54971 , RIc0d8398_29);
buf \U$54997 ( \54972 , RIc0dacd8_117);
xor \U$54998 ( \54973 , \54971 , \54972 );
buf \U$54999 ( \54974 , \54973 );
buf \U$55000 ( \54975 , \54974 );
not \U$55001 ( \54976 , \54975 );
buf \U$55002 ( \54977 , \54976 );
buf \U$55003 ( \54978 , \54977 );
or \U$55004 ( \54979 , \54970 , \54978 );
nand \U$55005 ( \54980 , \54969 , \54979 );
buf \U$55006 ( \54981 , \54980 );
buf \U$55007 ( \54982 , \54981 );
and \U$55008 ( \54983 , \54966 , \54982 );
and \U$55009 ( \54984 , \54958 , \54965 );
or \U$55010 ( \54985 , \54983 , \54984 );
buf \U$55011 ( \54986 , \54985 );
buf \U$55012 ( \54987 , \54986 );
buf \U$55013 ( \54988 , \53984 );
not \U$55014 ( \54989 , \54988 );
buf \U$55015 ( \54990 , \3714 );
not \U$55016 ( \54991 , \54990 );
or \U$55017 ( \54992 , \54989 , \54991 );
buf \U$55018 ( \54993 , \344 );
xor \U$55019 ( \54994 , RIc0da288_95, RIc0d8de8_51);
buf \U$55020 ( \54995 , \54994 );
nand \U$55021 ( \54996 , \54993 , \54995 );
buf \U$55022 ( \54997 , \54996 );
buf \U$55023 ( \54998 , \54997 );
nand \U$55024 ( \54999 , \54992 , \54998 );
buf \U$55025 ( \55000 , \54999 );
buf \U$55026 ( \55001 , \55000 );
not \U$55027 ( \55002 , \55001 );
buf \U$55028 ( \55003 , \54192 );
not \U$55029 ( \55004 , \55003 );
buf \U$55030 ( \55005 , \14569 );
not \U$55031 ( \55006 , \55005 );
or \U$55032 ( \55007 , \55004 , \55006 );
buf \U$55033 ( \55008 , \13005 );
buf \U$55034 ( \55009 , RIc0dadc8_119);
buf \U$55035 ( \55010 , RIc0d82a8_27);
xor \U$55036 ( \55011 , \55009 , \55010 );
buf \U$55037 ( \55012 , \55011 );
buf \U$55038 ( \55013 , \55012 );
nand \U$55039 ( \55014 , \55008 , \55013 );
buf \U$55040 ( \55015 , \55014 );
buf \U$55041 ( \55016 , \55015 );
nand \U$55042 ( \55017 , \55007 , \55016 );
buf \U$55043 ( \55018 , \55017 );
buf \U$55044 ( \55019 , \55018 );
not \U$55045 ( \55020 , \55019 );
or \U$55046 ( \55021 , \55002 , \55020 );
buf \U$55047 ( \55022 , \55000 );
buf \U$55048 ( \55023 , \55018 );
or \U$55049 ( \55024 , \55022 , \55023 );
buf \U$55050 ( \55025 , \17992 );
buf \U$55051 ( \55026 , \54211 );
or \U$55052 ( \55027 , \55025 , \55026 );
buf \U$55053 ( \55028 , \22744 );
buf \U$55054 ( \55029 , RIc0db098_125);
buf \U$55055 ( \55030 , RIc0d7fd8_21);
xnor \U$55056 ( \55031 , \55029 , \55030 );
buf \U$55057 ( \55032 , \55031 );
buf \U$55058 ( \55033 , \55032 );
or \U$55059 ( \55034 , \55028 , \55033 );
nand \U$55060 ( \55035 , \55027 , \55034 );
buf \U$55061 ( \55036 , \55035 );
buf \U$55062 ( \55037 , \55036 );
nand \U$55063 ( \55038 , \55024 , \55037 );
buf \U$55064 ( \55039 , \55038 );
buf \U$55065 ( \55040 , \55039 );
nand \U$55066 ( \55041 , \55021 , \55040 );
buf \U$55067 ( \55042 , \55041 );
buf \U$55068 ( \55043 , \55042 );
xor \U$55069 ( \55044 , \54987 , \55043 );
xor \U$55070 ( \55045 , \54811 , \54828 );
and \U$55071 ( \55046 , \55045 , \54845 );
and \U$55072 ( \55047 , \54811 , \54828 );
or \U$55073 ( \55048 , \55046 , \55047 );
buf \U$55074 ( \55049 , \55048 );
buf \U$55075 ( \55050 , \55049 );
xor \U$55076 ( \55051 , \55044 , \55050 );
buf \U$55077 ( \55052 , \55051 );
buf \U$55078 ( \55053 , \55052 );
xnor \U$55079 ( \55054 , \54943 , \55053 );
buf \U$55080 ( \55055 , \55054 );
buf \U$55081 ( \55056 , \55055 );
not \U$55082 ( \55057 , \55056 );
buf \U$55083 ( \55058 , \55057 );
buf \U$55084 ( \55059 , \55058 );
not \U$55085 ( \55060 , \55059 );
buf \U$55086 ( \55061 , \54607 );
buf \U$55087 ( \55062 , \54618 );
or \U$55088 ( \55063 , \55061 , \55062 );
buf \U$55089 ( \55064 , \54612 );
nand \U$55090 ( \55065 , \55063 , \55064 );
buf \U$55091 ( \55066 , \55065 );
buf \U$55092 ( \55067 , \55066 );
buf \U$55093 ( \55068 , \54607 );
buf \U$55094 ( \55069 , \54618 );
nand \U$55095 ( \55070 , \55068 , \55069 );
buf \U$55096 ( \55071 , \55070 );
buf \U$55097 ( \55072 , \55071 );
nand \U$55098 ( \55073 , \55067 , \55072 );
buf \U$55099 ( \55074 , \55073 );
buf \U$55100 ( \55075 , RIc0d8140_24);
buf \U$55101 ( \55076 , RIc0daeb8_121);
xor \U$55102 ( \55077 , \55075 , \55076 );
buf \U$55103 ( \55078 , \55077 );
buf \U$55104 ( \55079 , \55078 );
not \U$55105 ( \55080 , \55079 );
buf \U$55106 ( \55081 , \12975 );
not \U$55107 ( \55082 , \55081 );
or \U$55108 ( \55083 , \55080 , \55082 );
buf \U$55109 ( \55084 , \52081 );
buf \U$55110 ( \55085 , \54821 );
buf \U$55111 ( \55086 , \12964 );
nand \U$55112 ( \55087 , \55084 , \55085 , \55086 );
buf \U$55113 ( \55088 , \55087 );
buf \U$55114 ( \55089 , \55088 );
nand \U$55115 ( \55090 , \55083 , \55089 );
buf \U$55116 ( \55091 , \55090 );
buf \U$55117 ( \55092 , \55091 );
buf \U$55118 ( \55093 , \54804 );
not \U$55119 ( \55094 , \55093 );
buf \U$55120 ( \55095 , \12402 );
not \U$55121 ( \55096 , \55095 );
or \U$55122 ( \55097 , \55094 , \55096 );
buf \U$55123 ( \55098 , \12410 );
buf \U$55124 ( \55099 , \53515 );
nand \U$55125 ( \55100 , \55098 , \55099 );
buf \U$55126 ( \55101 , \55100 );
buf \U$55127 ( \55102 , \55101 );
nand \U$55128 ( \55103 , \55097 , \55102 );
buf \U$55129 ( \55104 , \55103 );
buf \U$55130 ( \55105 , \55104 );
xor \U$55131 ( \55106 , \55092 , \55105 );
buf \U$55132 ( \55107 , \53925 );
not \U$55133 ( \55108 , \55107 );
buf \U$55134 ( \55109 , \14982 );
not \U$55135 ( \55110 , \55109 );
or \U$55136 ( \55111 , \55108 , \55110 );
buf \U$55137 ( \55112 , \16692 );
buf \U$55138 ( \55113 , \53659 );
nand \U$55139 ( \55114 , \55112 , \55113 );
buf \U$55140 ( \55115 , \55114 );
buf \U$55141 ( \55116 , \55115 );
nand \U$55142 ( \55117 , \55111 , \55116 );
buf \U$55143 ( \55118 , \55117 );
buf \U$55144 ( \55119 , \55118 );
xor \U$55145 ( \55120 , \55106 , \55119 );
buf \U$55146 ( \55121 , \55120 );
buf \U$55147 ( \55122 , \55121 );
xor \U$55148 ( \55123 , \54898 , \54915 );
and \U$55149 ( \55124 , \55123 , \54933 );
and \U$55150 ( \55125 , \54898 , \54915 );
or \U$55151 ( \55126 , \55124 , \55125 );
buf \U$55152 ( \55127 , \55126 );
buf \U$55153 ( \55128 , \55127 );
xor \U$55154 ( \55129 , \55122 , \55128 );
buf \U$55155 ( \55130 , \54056 );
not \U$55156 ( \55131 , \55130 );
buf \U$55157 ( \55132 , \618 );
not \U$55158 ( \55133 , \55132 );
or \U$55159 ( \55134 , \55131 , \55133 );
buf \U$55160 ( \55135 , \816 );
buf \U$55161 ( \55136 , \53874 );
nand \U$55162 ( \55137 , \55135 , \55136 );
buf \U$55163 ( \55138 , \55137 );
buf \U$55164 ( \55139 , \55138 );
nand \U$55165 ( \55140 , \55134 , \55139 );
buf \U$55166 ( \55141 , \55140 );
buf \U$55167 ( \55142 , \55141 );
buf \U$55168 ( \55143 , \54130 );
not \U$55169 ( \55144 , \55143 );
buf \U$55170 ( \55145 , \437 );
not \U$55171 ( \55146 , \55145 );
or \U$55172 ( \55147 , \55144 , \55146 );
buf \U$55173 ( \55148 , \442 );
buf \U$55174 ( \55149 , RIc0d9fb8_89);
buf \U$55175 ( \55150 , RIc0d90b8_57);
xor \U$55176 ( \55151 , \55149 , \55150 );
buf \U$55177 ( \55152 , \55151 );
buf \U$55178 ( \55153 , \55152 );
nand \U$55179 ( \55154 , \55148 , \55153 );
buf \U$55180 ( \55155 , \55154 );
buf \U$55181 ( \55156 , \55155 );
nand \U$55182 ( \55157 , \55147 , \55156 );
buf \U$55183 ( \55158 , \55157 );
buf \U$55184 ( \55159 , \55158 );
or \U$55185 ( \55160 , \55142 , \55159 );
buf \U$55186 ( \55161 , \54570 );
not \U$55187 ( \55162 , \55161 );
buf \U$55188 ( \55163 , \3535 );
not \U$55189 ( \55164 , \55163 );
or \U$55190 ( \55165 , \55162 , \55164 );
buf \U$55191 ( \55166 , \16676 );
buf \U$55192 ( \55167 , \53861 );
nand \U$55193 ( \55168 , \55166 , \55167 );
buf \U$55194 ( \55169 , \55168 );
buf \U$55195 ( \55170 , \55169 );
nand \U$55196 ( \55171 , \55165 , \55170 );
buf \U$55197 ( \55172 , \55171 );
buf \U$55198 ( \55173 , \55172 );
nand \U$55199 ( \55174 , \55160 , \55173 );
buf \U$55200 ( \55175 , \55174 );
buf \U$55201 ( \55176 , \55175 );
buf \U$55202 ( \55177 , \55141 );
buf \U$55203 ( \55178 , \55158 );
nand \U$55204 ( \55179 , \55177 , \55178 );
buf \U$55205 ( \55180 , \55179 );
buf \U$55206 ( \55181 , \55180 );
nand \U$55207 ( \55182 , \55176 , \55181 );
buf \U$55208 ( \55183 , \55182 );
buf \U$55209 ( \55184 , \55183 );
xor \U$55210 ( \55185 , \55129 , \55184 );
buf \U$55211 ( \55186 , \55185 );
xor \U$55212 ( \55187 , \55074 , \55186 );
xor \U$55213 ( \55188 , \54748 , \54730 );
xor \U$55214 ( \55189 , \55188 , \54771 );
buf \U$55215 ( \55190 , \55189 );
not \U$55216 ( \55191 , \55190 );
xor \U$55217 ( \55192 , \54958 , \54965 );
xor \U$55218 ( \55193 , \55192 , \54982 );
buf \U$55219 ( \55194 , \55193 );
buf \U$55220 ( \55195 , \55194 );
not \U$55221 ( \55196 , \55195 );
or \U$55222 ( \55197 , \55191 , \55196 );
buf \U$55223 ( \55198 , \55194 );
buf \U$55224 ( \55199 , \55189 );
or \U$55225 ( \55200 , \55198 , \55199 );
xor \U$55226 ( \55201 , \55018 , \55000 );
xor \U$55227 ( \55202 , \55201 , \55036 );
buf \U$55228 ( \55203 , \55202 );
nand \U$55229 ( \55204 , \55200 , \55203 );
buf \U$55230 ( \55205 , \55204 );
buf \U$55231 ( \55206 , \55205 );
nand \U$55232 ( \55207 , \55197 , \55206 );
buf \U$55233 ( \55208 , \55207 );
xnor \U$55234 ( \55209 , \55187 , \55208 );
buf \U$55235 ( \55210 , \55209 );
not \U$55236 ( \55211 , \55210 );
buf \U$55237 ( \55212 , \55211 );
buf \U$55238 ( \55213 , \55212 );
not \U$55239 ( \55214 , \55213 );
or \U$55240 ( \55215 , \55060 , \55214 );
buf \U$55241 ( \55216 , \55055 );
not \U$55242 ( \55217 , \55216 );
buf \U$55243 ( \55218 , \55209 );
not \U$55244 ( \55219 , \55218 );
or \U$55245 ( \55220 , \55217 , \55219 );
buf \U$55246 ( \55221 , \54872 );
not \U$55247 ( \55222 , \55221 );
buf \U$55248 ( \55223 , \54935 );
not \U$55249 ( \55224 , \55223 );
or \U$55250 ( \55225 , \55222 , \55224 );
buf \U$55251 ( \55226 , \54935 );
buf \U$55252 ( \55227 , \54872 );
or \U$55253 ( \55228 , \55226 , \55227 );
nand \U$55254 ( \55229 , \55225 , \55228 );
buf \U$55255 ( \55230 , \55229 );
buf \U$55256 ( \55231 , \55230 );
buf \U$55257 ( \55232 , \54847 );
xor \U$55258 ( \55233 , \55231 , \55232 );
buf \U$55259 ( \55234 , \55233 );
buf \U$55260 ( \55235 , \55234 );
not \U$55261 ( \55236 , \55235 );
xor \U$55262 ( \55237 , \54120 , \54137 );
xor \U$55263 ( \55238 , \55237 , \54158 );
buf \U$55264 ( \55239 , \55238 );
buf \U$55265 ( \55240 , \55239 );
xor \U$55266 ( \55241 , \54558 , \54576 );
xor \U$55267 ( \55242 , \55241 , \54601 );
buf \U$55268 ( \55243 , \55242 );
xor \U$55269 ( \55244 , \55240 , \55243 );
buf \U$55270 ( \55245 , \48503 );
not \U$55271 ( \55246 , \55245 );
buf \U$55272 ( \55247 , \28794 );
not \U$55273 ( \55248 , \55247 );
or \U$55274 ( \55249 , \55246 , \55248 );
buf \U$55275 ( \55250 , \12342 );
buf \U$55276 ( \55251 , \54736 );
nand \U$55277 ( \55252 , \55250 , \55251 );
buf \U$55278 ( \55253 , \55252 );
buf \U$55279 ( \55254 , \55253 );
nand \U$55280 ( \55255 , \55249 , \55254 );
buf \U$55281 ( \55256 , \55255 );
buf \U$55282 ( \55257 , \55256 );
not \U$55283 ( \55258 , \55257 );
buf \U$55284 ( \55259 , \55258 );
buf \U$55285 ( \55260 , \48535 );
not \U$55286 ( \55261 , \55260 );
buf \U$55287 ( \55262 , \14982 );
not \U$55288 ( \55263 , \55262 );
or \U$55289 ( \55264 , \55261 , \55263 );
buf \U$55290 ( \55265 , \14278 );
buf \U$55291 ( \55266 , \53911 );
nand \U$55292 ( \55267 , \55265 , \55266 );
buf \U$55293 ( \55268 , \55267 );
buf \U$55294 ( \55269 , \55268 );
nand \U$55295 ( \55270 , \55264 , \55269 );
buf \U$55296 ( \55271 , \55270 );
xor \U$55297 ( \55272 , \55259 , \55271 );
buf \U$55298 ( \55273 , \48585 );
not \U$55299 ( \55274 , \55273 );
buf \U$55300 ( \55275 , \48600 );
nor \U$55301 ( \55276 , \55274 , \55275 );
buf \U$55302 ( \55277 , \55276 );
xnor \U$55303 ( \55278 , \55272 , \55277 );
buf \U$55304 ( \55279 , \55278 );
and \U$55305 ( \55280 , \55244 , \55279 );
and \U$55306 ( \55281 , \55240 , \55243 );
or \U$55307 ( \55282 , \55280 , \55281 );
buf \U$55308 ( \55283 , \55282 );
buf \U$55309 ( \55284 , \55283 );
not \U$55310 ( \55285 , \55284 );
or \U$55311 ( \55286 , \55236 , \55285 );
buf \U$55312 ( \55287 , \55234 );
buf \U$55313 ( \55288 , \55283 );
or \U$55314 ( \55289 , \55287 , \55288 );
xor \U$55315 ( \55290 , \55194 , \55202 );
xor \U$55316 ( \55291 , \55290 , \55189 );
buf \U$55317 ( \55292 , \55291 );
nand \U$55318 ( \55293 , \55289 , \55292 );
buf \U$55319 ( \55294 , \55293 );
buf \U$55320 ( \55295 , \55294 );
nand \U$55321 ( \55296 , \55286 , \55295 );
buf \U$55322 ( \55297 , \55296 );
buf \U$55323 ( \55298 , \55297 );
nand \U$55324 ( \55299 , \55220 , \55298 );
buf \U$55325 ( \55300 , \55299 );
buf \U$55326 ( \55301 , \55300 );
nand \U$55327 ( \55302 , \55215 , \55301 );
buf \U$55328 ( \55303 , \55302 );
buf \U$55329 ( \55304 , \55303 );
xor \U$55330 ( \55305 , \54638 , \55304 );
buf \U$55331 ( \55306 , \55305 );
buf \U$55332 ( \55307 , \55306 );
buf \U$55333 ( \55308 , \54788 );
not \U$55334 ( \55309 , \55308 );
buf \U$55335 ( \55310 , \54777 );
not \U$55336 ( \55311 , \55310 );
or \U$55337 ( \55312 , \55309 , \55311 );
buf \U$55338 ( \55313 , \54782 );
not \U$55339 ( \55314 , \55313 );
buf \U$55340 ( \55315 , \54777 );
not \U$55341 ( \55316 , \55315 );
buf \U$55342 ( \55317 , \55316 );
buf \U$55343 ( \55318 , \55317 );
not \U$55344 ( \55319 , \55318 );
or \U$55345 ( \55320 , \55314 , \55319 );
buf \U$55346 ( \55321 , \54716 );
nand \U$55347 ( \55322 , \55320 , \55321 );
buf \U$55348 ( \55323 , \55322 );
buf \U$55349 ( \55324 , \55323 );
nand \U$55350 ( \55325 , \55312 , \55324 );
buf \U$55351 ( \55326 , \55325 );
buf \U$55352 ( \55327 , \55326 );
buf \U$55353 ( \55328 , RIc0d9ce8_83);
buf \U$55354 ( \55329 , RIc0d9310_62);
xor \U$55355 ( \55330 , \55328 , \55329 );
buf \U$55356 ( \55331 , \55330 );
buf \U$55357 ( \55332 , \55331 );
not \U$55358 ( \55333 , \55332 );
buf \U$55359 ( \55334 , \1736 );
not \U$55360 ( \55335 , \55334 );
or \U$55361 ( \55336 , \55333 , \55335 );
buf \U$55362 ( \55337 , \584 );
buf \U$55363 ( \55338 , RIc0d9ce8_83);
buf \U$55364 ( \55339 , RIc0d9298_61);
xor \U$55365 ( \55340 , \55338 , \55339 );
buf \U$55366 ( \55341 , \55340 );
buf \U$55367 ( \55342 , \55341 );
nand \U$55368 ( \55343 , \55337 , \55342 );
buf \U$55369 ( \55344 , \55343 );
buf \U$55370 ( \55345 , \55344 );
nand \U$55371 ( \55346 , \55336 , \55345 );
buf \U$55372 ( \55347 , \55346 );
buf \U$55373 ( \55348 , \55347 );
buf \U$55374 ( \55349 , RIc0d9400_64);
buf \U$55375 ( \55350 , RIc0d9c70_82);
or \U$55376 ( \55351 , \55349 , \55350 );
buf \U$55377 ( \55352 , RIc0d9ce8_83);
nand \U$55378 ( \55353 , \55351 , \55352 );
buf \U$55379 ( \55354 , \55353 );
buf \U$55380 ( \55355 , \55354 );
buf \U$55381 ( \55356 , RIc0d9400_64);
buf \U$55382 ( \55357 , RIc0d9c70_82);
nand \U$55383 ( \55358 , \55356 , \55357 );
buf \U$55384 ( \55359 , \55358 );
buf \U$55385 ( \55360 , \55359 );
buf \U$55386 ( \55361 , RIc0d9bf8_81);
and \U$55387 ( \55362 , \55355 , \55360 , \55361 );
buf \U$55388 ( \55363 , \55362 );
buf \U$55389 ( \55364 , \55363 );
xor \U$55390 ( \55365 , \55348 , \55364 );
buf \U$55391 ( \55366 , \55365 );
buf \U$55392 ( \55367 , \55366 );
not \U$55393 ( \55368 , \55367 );
buf \U$55394 ( \55369 , \55368 );
buf \U$55395 ( \55370 , \55369 );
not \U$55396 ( \55371 , \55370 );
buf \U$55397 ( \55372 , \55078 );
not \U$55398 ( \55373 , \55372 );
buf \U$55399 ( \55374 , \24672 );
not \U$55400 ( \55375 , \55374 );
or \U$55401 ( \55376 , \55373 , \55375 );
buf \U$55402 ( \55377 , \13314 );
xor \U$55403 ( \55378 , RIc0daeb8_121, RIc0d80c8_23);
buf \U$55404 ( \55379 , \55378 );
nand \U$55405 ( \55380 , \55377 , \55379 );
buf \U$55406 ( \55381 , \55380 );
buf \U$55407 ( \55382 , \55381 );
nand \U$55408 ( \55383 , \55376 , \55382 );
buf \U$55409 ( \55384 , \55383 );
xor \U$55410 ( \55385 , RIc0db098_125, RIc0d7f60_20);
buf \U$55411 ( \55386 , \55385 );
not \U$55412 ( \55387 , \55386 );
buf \U$55413 ( \55388 , \44382 );
not \U$55414 ( \55389 , \55388 );
or \U$55415 ( \55390 , \55387 , \55389 );
buf \U$55416 ( \55391 , \15793 );
xor \U$55417 ( \55392 , RIc0db098_125, RIc0d7ee8_19);
buf \U$55418 ( \55393 , \55392 );
nand \U$55419 ( \55394 , \55391 , \55393 );
buf \U$55420 ( \55395 , \55394 );
buf \U$55421 ( \55396 , \55395 );
nand \U$55422 ( \55397 , \55390 , \55396 );
buf \U$55423 ( \55398 , \55397 );
xor \U$55424 ( \55399 , \55384 , \55398 );
buf \U$55425 ( \55400 , \55399 );
not \U$55426 ( \55401 , \55400 );
or \U$55427 ( \55402 , \55371 , \55401 );
buf \U$55428 ( \55403 , \55399 );
buf \U$55429 ( \55404 , \55369 );
or \U$55430 ( \55405 , \55403 , \55404 );
nand \U$55431 ( \55406 , \55402 , \55405 );
buf \U$55432 ( \55407 , \55406 );
buf \U$55433 ( \55408 , \55407 );
xor \U$55434 ( \55409 , \55327 , \55408 );
xor \U$55435 ( \55410 , \54987 , \55043 );
and \U$55436 ( \55411 , \55410 , \55050 );
and \U$55437 ( \55412 , \54987 , \55043 );
or \U$55438 ( \55413 , \55411 , \55412 );
buf \U$55439 ( \55414 , \55413 );
buf \U$55440 ( \55415 , \55414 );
xor \U$55441 ( \55416 , \55409 , \55415 );
buf \U$55442 ( \55417 , \55416 );
buf \U$55443 ( \55418 , \55417 );
buf \U$55444 ( \55419 , \55208 );
not \U$55445 ( \55420 , \55419 );
buf \U$55446 ( \55421 , \55074 );
not \U$55447 ( \55422 , \55421 );
or \U$55448 ( \55423 , \55420 , \55422 );
buf \U$55449 ( \55424 , \55074 );
buf \U$55450 ( \55425 , \55208 );
or \U$55451 ( \55426 , \55424 , \55425 );
buf \U$55452 ( \55427 , \55186 );
nand \U$55453 ( \55428 , \55426 , \55427 );
buf \U$55454 ( \55429 , \55428 );
buf \U$55455 ( \55430 , \55429 );
nand \U$55456 ( \55431 , \55423 , \55430 );
buf \U$55457 ( \55432 , \55431 );
buf \U$55458 ( \55433 , \55432 );
xor \U$55459 ( \55434 , \55418 , \55433 );
buf \U$55460 ( \55435 , \54793 );
not \U$55461 ( \55436 , \55435 );
buf \U$55462 ( \55437 , \55052 );
not \U$55463 ( \55438 , \55437 );
or \U$55464 ( \55439 , \55436 , \55438 );
buf \U$55465 ( \55440 , \55052 );
buf \U$55466 ( \55441 , \54793 );
or \U$55467 ( \55442 , \55440 , \55441 );
buf \U$55468 ( \55443 , \54941 );
nand \U$55469 ( \55444 , \55442 , \55443 );
buf \U$55470 ( \55445 , \55444 );
buf \U$55471 ( \55446 , \55445 );
nand \U$55472 ( \55447 , \55439 , \55446 );
buf \U$55473 ( \55448 , \55447 );
buf \U$55474 ( \55449 , \55448 );
xor \U$55475 ( \55450 , \55434 , \55449 );
buf \U$55476 ( \55451 , \55450 );
buf \U$55477 ( \55452 , \55451 );
buf \U$55478 ( \55453 , \1078 );
buf \U$55479 ( \55454 , RIc0d9400_64);
and \U$55480 ( \55455 , \55453 , \55454 );
buf \U$55481 ( \55456 , \55455 );
buf \U$55482 ( \55457 , \55456 );
buf \U$55483 ( \55458 , \53947 );
not \U$55484 ( \55459 , \55458 );
buf \U$55485 ( \55460 , \6029 );
not \U$55486 ( \55461 , \55460 );
or \U$55487 ( \55462 , \55459 , \55461 );
buf \U$55488 ( \55463 , \1401 );
buf \U$55489 ( \55464 , \53821 );
nand \U$55490 ( \55465 , \55463 , \55464 );
buf \U$55491 ( \55466 , \55465 );
buf \U$55492 ( \55467 , \55466 );
nand \U$55493 ( \55468 , \55462 , \55467 );
buf \U$55494 ( \55469 , \55468 );
buf \U$55495 ( \55470 , \55469 );
xor \U$55496 ( \55471 , \55457 , \55470 );
buf \U$55497 ( \55472 , \54669 );
not \U$55498 ( \55473 , \55472 );
buf \U$55499 ( \55474 , \14210 );
not \U$55500 ( \55475 , \55474 );
or \U$55501 ( \55476 , \55473 , \55475 );
buf \U$55502 ( \55477 , \15909 );
buf \U$55503 ( \55478 , \53638 );
nand \U$55504 ( \55479 , \55477 , \55478 );
buf \U$55505 ( \55480 , \55479 );
buf \U$55506 ( \55481 , \55480 );
nand \U$55507 ( \55482 , \55476 , \55481 );
buf \U$55508 ( \55483 , \55482 );
buf \U$55509 ( \55484 , \55483 );
xor \U$55510 ( \55485 , \55471 , \55484 );
buf \U$55511 ( \55486 , \55485 );
buf \U$55512 ( \55487 , \55486 );
buf \U$55513 ( \55488 , \54944 );
not \U$55514 ( \55489 , \55488 );
buf \U$55515 ( \55490 , \18220 );
not \U$55516 ( \55491 , \55490 );
or \U$55517 ( \55492 , \55489 , \55491 );
buf \U$55518 ( \55493 , \20243 );
buf \U$55519 ( \55494 , \53601 );
nand \U$55520 ( \55495 , \55493 , \55494 );
buf \U$55521 ( \55496 , \55495 );
buf \U$55522 ( \55497 , \55496 );
nand \U$55523 ( \55498 , \55492 , \55497 );
buf \U$55524 ( \55499 , \55498 );
buf \U$55525 ( \55500 , \54974 );
not \U$55526 ( \55501 , \55500 );
buf \U$55527 ( \55502 , \12923 );
not \U$55528 ( \55503 , \55502 );
or \U$55529 ( \55504 , \55501 , \55503 );
buf \U$55530 ( \55505 , \12937 );
buf \U$55531 ( \55506 , \53562 );
nand \U$55532 ( \55507 , \55505 , \55506 );
buf \U$55533 ( \55508 , \55507 );
buf \U$55534 ( \55509 , \55508 );
nand \U$55535 ( \55510 , \55504 , \55509 );
buf \U$55536 ( \55511 , \55510 );
xor \U$55537 ( \55512 , \55499 , \55511 );
buf \U$55538 ( \55513 , \55512 );
buf \U$55539 ( \55514 , \54891 );
not \U$55540 ( \55515 , \55514 );
buf \U$55541 ( \55516 , \2535 );
not \U$55542 ( \55517 , \55516 );
or \U$55543 ( \55518 , \55515 , \55517 );
buf \U$55544 ( \55519 , \714 );
buf \U$55545 ( \55520 , \53471 );
nand \U$55546 ( \55521 , \55519 , \55520 );
buf \U$55547 ( \55522 , \55521 );
buf \U$55548 ( \55523 , \55522 );
nand \U$55549 ( \55524 , \55518 , \55523 );
buf \U$55550 ( \55525 , \55524 );
buf \U$55551 ( \55526 , \55525 );
xor \U$55552 ( \55527 , \55513 , \55526 );
buf \U$55553 ( \55528 , \55527 );
buf \U$55554 ( \55529 , \55528 );
xor \U$55555 ( \55530 , \55487 , \55529 );
buf \U$55556 ( \55531 , \44640 );
buf \U$55557 ( \55532 , \54959 );
not \U$55558 ( \55533 , \55532 );
buf \U$55559 ( \55534 , \55533 );
buf \U$55560 ( \55535 , \55534 );
or \U$55561 ( \55536 , \55531 , \55535 );
buf \U$55562 ( \55537 , \12647 );
buf \U$55563 ( \55538 , \53428 );
not \U$55564 ( \55539 , \55538 );
buf \U$55565 ( \55540 , \55539 );
buf \U$55566 ( \55541 , \55540 );
or \U$55567 ( \55542 , \55537 , \55541 );
nand \U$55568 ( \55543 , \55536 , \55542 );
buf \U$55569 ( \55544 , \55543 );
buf \U$55570 ( \55545 , \55544 );
buf \U$55571 ( \55546 , \54717 );
not \U$55572 ( \55547 , \55546 );
buf \U$55573 ( \55548 , \2066 );
not \U$55574 ( \55549 , \55548 );
or \U$55575 ( \55550 , \55547 , \55549 );
buf \U$55576 ( \55551 , RIc0da378_97);
buf \U$55577 ( \55552 , RIc0d8c80_48);
xnor \U$55578 ( \55553 , \55551 , \55552 );
buf \U$55579 ( \55554 , \55553 );
buf \U$55580 ( \55555 , \55554 );
not \U$55581 ( \55556 , \55555 );
buf \U$55582 ( \55557 , \734 );
nand \U$55583 ( \55558 , \55556 , \55557 );
buf \U$55584 ( \55559 , \55558 );
buf \U$55585 ( \55560 , \55559 );
nand \U$55586 ( \55561 , \55550 , \55560 );
buf \U$55587 ( \55562 , \55561 );
buf \U$55588 ( \55563 , \55562 );
xor \U$55589 ( \55564 , \55545 , \55563 );
buf \U$55590 ( \55565 , \12532 );
buf \U$55591 ( \55566 , \54763 );
or \U$55592 ( \55567 , \55565 , \55566 );
buf \U$55593 ( \55568 , \49542 );
buf \U$55594 ( \55569 , RIc0daa08_111);
buf \U$55595 ( \55570 , RIc0d85f0_34);
xor \U$55596 ( \55571 , \55569 , \55570 );
buf \U$55597 ( \55572 , \55571 );
buf \U$55598 ( \55573 , \55572 );
not \U$55599 ( \55574 , \55573 );
buf \U$55600 ( \55575 , \55574 );
buf \U$55601 ( \55576 , \55575 );
or \U$55602 ( \55577 , \55568 , \55576 );
nand \U$55603 ( \55578 , \55567 , \55577 );
buf \U$55604 ( \55579 , \55578 );
buf \U$55605 ( \55580 , \55579 );
xor \U$55606 ( \55581 , \55564 , \55580 );
buf \U$55607 ( \55582 , \55581 );
buf \U$55608 ( \55583 , \55582 );
xor \U$55609 ( \55584 , \55530 , \55583 );
buf \U$55610 ( \55585 , \55584 );
buf \U$55611 ( \55586 , \55585 );
not \U$55612 ( \55587 , \55586 );
buf \U$55613 ( \55588 , \55587 );
buf \U$55614 ( \55589 , \55588 );
not \U$55615 ( \55590 , \55589 );
buf \U$55616 ( \55591 , \55271 );
not \U$55617 ( \55592 , \55591 );
buf \U$55618 ( \55593 , \55259 );
nand \U$55619 ( \55594 , \55592 , \55593 );
buf \U$55620 ( \55595 , \55594 );
buf \U$55621 ( \55596 , \55595 );
not \U$55622 ( \55597 , \55596 );
buf \U$55623 ( \55598 , \55277 );
not \U$55624 ( \55599 , \55598 );
or \U$55625 ( \55600 , \55597 , \55599 );
buf \U$55626 ( \55601 , \55256 );
buf \U$55627 ( \55602 , \55271 );
nand \U$55628 ( \55603 , \55601 , \55602 );
buf \U$55629 ( \55604 , \55603 );
buf \U$55630 ( \55605 , \55604 );
nand \U$55631 ( \55606 , \55600 , \55605 );
buf \U$55632 ( \55607 , \55606 );
buf \U$55633 ( \55608 , \55607 );
xor \U$55634 ( \55609 , \55172 , \55141 );
xor \U$55635 ( \55610 , \55609 , \55158 );
buf \U$55636 ( \55611 , \55610 );
xor \U$55637 ( \55612 , \55608 , \55611 );
xor \U$55638 ( \55613 , \53933 , \53973 );
xor \U$55639 ( \55614 , \55613 , \54040 );
buf \U$55640 ( \55615 , \55614 );
buf \U$55641 ( \55616 , \55615 );
and \U$55642 ( \55617 , \55612 , \55616 );
and \U$55643 ( \55618 , \55608 , \55611 );
or \U$55644 ( \55619 , \55617 , \55618 );
buf \U$55645 ( \55620 , \55619 );
buf \U$55646 ( \55621 , \55620 );
not \U$55647 ( \55622 , \55621 );
buf \U$55648 ( \55623 , \55622 );
buf \U$55649 ( \55624 , \55623 );
not \U$55650 ( \55625 , \55624 );
or \U$55651 ( \55626 , \55590 , \55625 );
buf \U$55652 ( \55627 , \54648 );
not \U$55653 ( \55628 , \55627 );
buf \U$55654 ( \55629 , \14684 );
not \U$55655 ( \55630 , \55629 );
or \U$55656 ( \55631 , \55628 , \55630 );
buf \U$55657 ( \55632 , \12303 );
buf \U$55658 ( \55633 , \53745 );
nand \U$55659 ( \55634 , \55632 , \55633 );
buf \U$55660 ( \55635 , \55634 );
buf \U$55661 ( \55636 , \55635 );
nand \U$55662 ( \55637 , \55631 , \55636 );
buf \U$55663 ( \55638 , \55637 );
buf \U$55664 ( \55639 , \55638 );
buf \U$55665 ( \55640 , \55152 );
not \U$55666 ( \55641 , \55640 );
buf \U$55667 ( \55642 , \18150 );
not \U$55668 ( \55643 , \55642 );
or \U$55669 ( \55644 , \55641 , \55643 );
buf \U$55670 ( \55645 , \846 );
buf \U$55671 ( \55646 , \53449 );
nand \U$55672 ( \55647 , \55645 , \55646 );
buf \U$55673 ( \55648 , \55647 );
buf \U$55674 ( \55649 , \55648 );
nand \U$55675 ( \55650 , \55644 , \55649 );
buf \U$55676 ( \55651 , \55650 );
buf \U$55677 ( \55652 , \55651 );
xor \U$55678 ( \55653 , \55639 , \55652 );
buf \U$55679 ( \55654 , \54699 );
not \U$55680 ( \55655 , \55654 );
buf \U$55681 ( \55656 , \1736 );
not \U$55682 ( \55657 , \55656 );
or \U$55683 ( \55658 , \55655 , \55657 );
buf \U$55684 ( \55659 , \584 );
buf \U$55685 ( \55660 , \55331 );
nand \U$55686 ( \55661 , \55659 , \55660 );
buf \U$55687 ( \55662 , \55661 );
buf \U$55688 ( \55663 , \55662 );
nand \U$55689 ( \55664 , \55658 , \55663 );
buf \U$55690 ( \55665 , \55664 );
buf \U$55691 ( \55666 , \55665 );
xor \U$55692 ( \55667 , \55653 , \55666 );
buf \U$55693 ( \55668 , \55667 );
buf \U$55694 ( \55669 , \55668 );
buf \U$55695 ( \55670 , \54837 );
not \U$55696 ( \55671 , \55670 );
buf \U$55697 ( \55672 , \2470 );
not \U$55698 ( \55673 , \55672 );
or \U$55699 ( \55674 , \55671 , \55673 );
buf \U$55700 ( \55675 , \2476 );
buf \U$55701 ( \55676 , \53773 );
nand \U$55702 ( \55677 , \55675 , \55676 );
buf \U$55703 ( \55678 , \55677 );
buf \U$55704 ( \55679 , \55678 );
nand \U$55705 ( \55680 , \55674 , \55679 );
buf \U$55706 ( \55681 , \55680 );
buf \U$55707 ( \55682 , \55681 );
buf \U$55708 ( \55683 , \55032 );
not \U$55709 ( \55684 , \55683 );
buf \U$55710 ( \55685 , \55684 );
buf \U$55711 ( \55686 , \55685 );
not \U$55712 ( \55687 , \55686 );
buf \U$55713 ( \55688 , \51095 );
not \U$55714 ( \55689 , \55688 );
or \U$55715 ( \55690 , \55687 , \55689 );
buf \U$55716 ( \55691 , \15793 );
buf \U$55717 ( \55692 , \55385 );
nand \U$55718 ( \55693 , \55691 , \55692 );
buf \U$55719 ( \55694 , \55693 );
buf \U$55720 ( \55695 , \55694 );
nand \U$55721 ( \55696 , \55690 , \55695 );
buf \U$55722 ( \55697 , \55696 );
buf \U$55723 ( \55698 , \55697 );
xor \U$55724 ( \55699 , \55682 , \55698 );
buf \U$55725 ( \55700 , \13949 );
not \U$55726 ( \55701 , \55700 );
buf \U$55727 ( \55702 , \55701 );
buf \U$55728 ( \55703 , \55702 );
buf \U$55729 ( \55704 , \55012 );
not \U$55730 ( \55705 , \55704 );
buf \U$55731 ( \55706 , \55705 );
buf \U$55732 ( \55707 , \55706 );
or \U$55733 ( \55708 , \55703 , \55707 );
buf \U$55734 ( \55709 , \45225 );
xor \U$55735 ( \55710 , RIc0dadc8_119, RIc0d8230_26);
buf \U$55736 ( \55711 , \55710 );
not \U$55737 ( \55712 , \55711 );
buf \U$55738 ( \55713 , \55712 );
buf \U$55739 ( \55714 , \55713 );
or \U$55740 ( \55715 , \55709 , \55714 );
nand \U$55741 ( \55716 , \55708 , \55715 );
buf \U$55742 ( \55717 , \55716 );
buf \U$55743 ( \55718 , \55717 );
xor \U$55744 ( \55719 , \55699 , \55718 );
buf \U$55745 ( \55720 , \55719 );
buf \U$55746 ( \55721 , \55720 );
xor \U$55747 ( \55722 , \55669 , \55721 );
buf \U$55748 ( \55723 , \54908 );
not \U$55749 ( \55724 , \55723 );
buf \U$55750 ( \55725 , \12736 );
not \U$55751 ( \55726 , \55725 );
or \U$55752 ( \55727 , \55724 , \55726 );
buf \U$55753 ( \55728 , \12744 );
buf \U$55754 ( \55729 , \53707 );
nand \U$55755 ( \55730 , \55728 , \55729 );
buf \U$55756 ( \55731 , \55730 );
buf \U$55757 ( \55732 , \55731 );
nand \U$55758 ( \55733 , \55727 , \55732 );
buf \U$55759 ( \55734 , \55733 );
buf \U$55760 ( \55735 , \54994 );
not \U$55761 ( \55736 , \55735 );
buf \U$55762 ( \55737 , \3714 );
not \U$55763 ( \55738 , \55737 );
or \U$55764 ( \55739 , \55736 , \55738 );
buf \U$55765 ( \55740 , \14707 );
buf \U$55766 ( \55741 , \53679 );
nand \U$55767 ( \55742 , \55740 , \55741 );
buf \U$55768 ( \55743 , \55742 );
buf \U$55769 ( \55744 , \55743 );
nand \U$55770 ( \55745 , \55739 , \55744 );
buf \U$55771 ( \55746 , \55745 );
xor \U$55772 ( \55747 , \55734 , \55746 );
buf \U$55773 ( \55748 , \54926 );
not \U$55774 ( \55749 , \55748 );
buf \U$55775 ( \55750 , \889 );
not \U$55776 ( \55751 , \55750 );
or \U$55777 ( \55752 , \55749 , \55751 );
buf \U$55778 ( \55753 , \4008 );
buf \U$55779 ( \55754 , \53582 );
nand \U$55780 ( \55755 , \55753 , \55754 );
buf \U$55781 ( \55756 , \55755 );
buf \U$55782 ( \55757 , \55756 );
nand \U$55783 ( \55758 , \55752 , \55757 );
buf \U$55784 ( \55759 , \55758 );
xor \U$55785 ( \55760 , \55747 , \55759 );
buf \U$55786 ( \55761 , \55760 );
xor \U$55787 ( \55762 , \55722 , \55761 );
buf \U$55788 ( \55763 , \55762 );
buf \U$55789 ( \55764 , \55763 );
nand \U$55790 ( \55765 , \55626 , \55764 );
buf \U$55791 ( \55766 , \55765 );
buf \U$55792 ( \55767 , \55766 );
buf \U$55793 ( \55768 , \55585 );
buf \U$55794 ( \55769 , \55620 );
nand \U$55795 ( \55770 , \55768 , \55769 );
buf \U$55796 ( \55771 , \55770 );
buf \U$55797 ( \55772 , \55771 );
nand \U$55798 ( \55773 , \55767 , \55772 );
buf \U$55799 ( \55774 , \55773 );
buf \U$55800 ( \55775 , \55774 );
xor \U$55801 ( \55776 , \55639 , \55652 );
and \U$55802 ( \55777 , \55776 , \55666 );
and \U$55803 ( \55778 , \55639 , \55652 );
or \U$55804 ( \55779 , \55777 , \55778 );
buf \U$55805 ( \55780 , \55779 );
buf \U$55806 ( \55781 , \55780 );
not \U$55807 ( \55782 , \55781 );
buf \U$55808 ( \55783 , \55511 );
buf \U$55809 ( \55784 , \55499 );
or \U$55810 ( \55785 , \55783 , \55784 );
buf \U$55811 ( \55786 , \55525 );
nand \U$55812 ( \55787 , \55785 , \55786 );
buf \U$55813 ( \55788 , \55787 );
buf \U$55814 ( \55789 , \55788 );
buf \U$55815 ( \55790 , \55511 );
buf \U$55816 ( \55791 , \55499 );
nand \U$55817 ( \55792 , \55790 , \55791 );
buf \U$55818 ( \55793 , \55792 );
buf \U$55819 ( \55794 , \55793 );
nand \U$55820 ( \55795 , \55789 , \55794 );
buf \U$55821 ( \55796 , \55795 );
buf \U$55822 ( \55797 , \55796 );
not \U$55823 ( \55798 , \55797 );
buf \U$55824 ( \55799 , \55798 );
buf \U$55825 ( \55800 , \55799 );
not \U$55826 ( \55801 , \55800 );
or \U$55827 ( \55802 , \55782 , \55801 );
not \U$55828 ( \55803 , \55780 );
buf \U$55829 ( \55804 , \55803 );
buf \U$55830 ( \55805 , \55796 );
nand \U$55831 ( \55806 , \55804 , \55805 );
buf \U$55832 ( \55807 , \55806 );
buf \U$55833 ( \55808 , \55807 );
nand \U$55834 ( \55809 , \55802 , \55808 );
buf \U$55835 ( \55810 , \55809 );
buf \U$55836 ( \55811 , \55810 );
buf \U$55837 ( \55812 , \55572 );
not \U$55838 ( \55813 , \55812 );
buf \U$55839 ( \55814 , \14346 );
not \U$55840 ( \55815 , \55814 );
or \U$55841 ( \55816 , \55813 , \55815 );
buf \U$55842 ( \55817 , \14353 );
buf \U$55843 ( \55818 , RIc0d8578_33);
buf \U$55844 ( \55819 , RIc0daa08_111);
xor \U$55845 ( \55820 , \55818 , \55819 );
buf \U$55846 ( \55821 , \55820 );
buf \U$55847 ( \55822 , \55821 );
nand \U$55848 ( \55823 , \55817 , \55822 );
buf \U$55849 ( \55824 , \55823 );
buf \U$55850 ( \55825 , \55824 );
nand \U$55851 ( \55826 , \55816 , \55825 );
buf \U$55852 ( \55827 , \55826 );
buf \U$55853 ( \55828 , \55827 );
buf \U$55854 ( \55829 , \55710 );
not \U$55855 ( \55830 , \55829 );
buf \U$55856 ( \55831 , \23985 );
not \U$55857 ( \55832 , \55831 );
or \U$55858 ( \55833 , \55830 , \55832 );
buf \U$55859 ( \55834 , \45225 );
not \U$55860 ( \55835 , \55834 );
buf \U$55861 ( \55836 , RIc0dadc8_119);
buf \U$55862 ( \55837 , RIc0d81b8_25);
xor \U$55863 ( \55838 , \55836 , \55837 );
buf \U$55864 ( \55839 , \55838 );
buf \U$55865 ( \55840 , \55839 );
nand \U$55866 ( \55841 , \55835 , \55840 );
buf \U$55867 ( \55842 , \55841 );
buf \U$55868 ( \55843 , \55842 );
nand \U$55869 ( \55844 , \55833 , \55843 );
buf \U$55870 ( \55845 , \55844 );
buf \U$55871 ( \55846 , \55845 );
xor \U$55872 ( \55847 , \55828 , \55846 );
buf \U$55873 ( \55848 , \2938 );
buf \U$55874 ( \55849 , \55554 );
or \U$55875 ( \55850 , \55848 , \55849 );
buf \U$55876 ( \55851 , \737 );
buf \U$55877 ( \55852 , RIc0da378_97);
buf \U$55878 ( \55853 , RIc0d8c08_47);
xor \U$55879 ( \55854 , \55852 , \55853 );
buf \U$55880 ( \55855 , \55854 );
buf \U$55881 ( \55856 , \55855 );
not \U$55882 ( \55857 , \55856 );
buf \U$55883 ( \55858 , \55857 );
buf \U$55884 ( \55859 , \55858 );
or \U$55885 ( \55860 , \55851 , \55859 );
nand \U$55886 ( \55861 , \55850 , \55860 );
buf \U$55887 ( \55862 , \55861 );
buf \U$55888 ( \55863 , \55862 );
xor \U$55889 ( \55864 , \55847 , \55863 );
buf \U$55890 ( \55865 , \55864 );
buf \U$55891 ( \55866 , \55865 );
xnor \U$55892 ( \55867 , \55811 , \55866 );
buf \U$55893 ( \55868 , \55867 );
buf \U$55894 ( \55869 , \55868 );
not \U$55895 ( \55870 , \55869 );
buf \U$55896 ( \55871 , \55870 );
buf \U$55897 ( \55872 , \55871 );
not \U$55898 ( \55873 , \55872 );
buf \U$55899 ( \55874 , \55873 );
buf \U$55900 ( \55875 , \55874 );
not \U$55901 ( \55876 , \55875 );
xor \U$55902 ( \55877 , \55669 , \55721 );
and \U$55903 ( \55878 , \55877 , \55761 );
and \U$55904 ( \55879 , \55669 , \55721 );
or \U$55905 ( \55880 , \55878 , \55879 );
buf \U$55906 ( \55881 , \55880 );
buf \U$55907 ( \55882 , \55881 );
not \U$55908 ( \55883 , \55882 );
xor \U$55909 ( \55884 , \55122 , \55128 );
and \U$55910 ( \55885 , \55884 , \55184 );
and \U$55911 ( \55886 , \55122 , \55128 );
or \U$55912 ( \55887 , \55885 , \55886 );
buf \U$55913 ( \55888 , \55887 );
buf \U$55914 ( \55889 , \55888 );
not \U$55915 ( \55890 , \55889 );
buf \U$55916 ( \55891 , \55890 );
buf \U$55917 ( \55892 , \55891 );
not \U$55918 ( \55893 , \55892 );
or \U$55919 ( \55894 , \55883 , \55893 );
buf \U$55920 ( \55895 , \55881 );
buf \U$55921 ( \55896 , \55891 );
or \U$55922 ( \55897 , \55895 , \55896 );
nand \U$55923 ( \55898 , \55894 , \55897 );
buf \U$55924 ( \55899 , \55898 );
buf \U$55925 ( \55900 , \55899 );
not \U$55926 ( \55901 , \55900 );
or \U$55927 ( \55902 , \55876 , \55901 );
buf \U$55928 ( \55903 , \55899 );
buf \U$55929 ( \55904 , \55874 );
or \U$55930 ( \55905 , \55903 , \55904 );
nand \U$55931 ( \55906 , \55902 , \55905 );
buf \U$55932 ( \55907 , \55906 );
buf \U$55933 ( \55908 , \55907 );
xor \U$55934 ( \55909 , \55775 , \55908 );
xor \U$55935 ( \55910 , \55487 , \55529 );
and \U$55936 ( \55911 , \55910 , \55583 );
and \U$55937 ( \55912 , \55487 , \55529 );
or \U$55938 ( \55913 , \55911 , \55912 );
buf \U$55939 ( \55914 , \55913 );
buf \U$55940 ( \55915 , \55914 );
xor \U$55941 ( \55916 , \55092 , \55105 );
and \U$55942 ( \55917 , \55916 , \55119 );
and \U$55943 ( \55918 , \55092 , \55105 );
or \U$55944 ( \55919 , \55917 , \55918 );
buf \U$55945 ( \55920 , \55919 );
buf \U$55946 ( \55921 , \55920 );
buf \U$55947 ( \55922 , \55746 );
buf \U$55948 ( \55923 , \55734 );
or \U$55949 ( \55924 , \55922 , \55923 );
buf \U$55950 ( \55925 , \55759 );
nand \U$55951 ( \55926 , \55924 , \55925 );
buf \U$55952 ( \55927 , \55926 );
buf \U$55953 ( \55928 , \55927 );
buf \U$55954 ( \55929 , \55746 );
buf \U$55955 ( \55930 , \55734 );
nand \U$55956 ( \55931 , \55929 , \55930 );
buf \U$55957 ( \55932 , \55931 );
buf \U$55958 ( \55933 , \55932 );
nand \U$55959 ( \55934 , \55928 , \55933 );
buf \U$55960 ( \55935 , \55934 );
buf \U$55961 ( \55936 , \55935 );
xor \U$55962 ( \55937 , \55921 , \55936 );
xor \U$55963 ( \55938 , \55682 , \55698 );
and \U$55964 ( \55939 , \55938 , \55718 );
and \U$55965 ( \55940 , \55682 , \55698 );
or \U$55966 ( \55941 , \55939 , \55940 );
buf \U$55967 ( \55942 , \55941 );
buf \U$55968 ( \55943 , \55942 );
xnor \U$55969 ( \55944 , \55937 , \55943 );
buf \U$55970 ( \55945 , \55944 );
buf \U$55971 ( \55946 , \55945 );
not \U$55972 ( \55947 , \55946 );
buf \U$55973 ( \55948 , \55947 );
buf \U$55974 ( \55949 , \55948 );
and \U$55975 ( \55950 , \55915 , \55949 );
not \U$55976 ( \55951 , \55915 );
buf \U$55977 ( \55952 , \55945 );
and \U$55978 ( \55953 , \55951 , \55952 );
nor \U$55979 ( \55954 , \55950 , \55953 );
buf \U$55980 ( \55955 , \55954 );
xor \U$55981 ( \55956 , \55457 , \55470 );
and \U$55982 ( \55957 , \55956 , \55484 );
and \U$55983 ( \55958 , \55457 , \55470 );
or \U$55984 ( \55959 , \55957 , \55958 );
buf \U$55985 ( \55960 , \55959 );
buf \U$55986 ( \55961 , \53886 );
buf \U$55987 ( \55962 , \53873 );
or \U$55988 ( \55963 , \55961 , \55962 );
buf \U$55989 ( \55964 , \53902 );
nand \U$55990 ( \55965 , \55963 , \55964 );
buf \U$55991 ( \55966 , \55965 );
buf \U$55992 ( \55967 , \55966 );
buf \U$55993 ( \55968 , \53886 );
buf \U$55994 ( \55969 , \53873 );
nand \U$55995 ( \55970 , \55968 , \55969 );
buf \U$55996 ( \55971 , \55970 );
buf \U$55997 ( \55972 , \55971 );
nand \U$55998 ( \55973 , \55967 , \55972 );
buf \U$55999 ( \55974 , \55973 );
xor \U$56000 ( \55975 , \55960 , \55974 );
xor \U$56001 ( \55976 , \55545 , \55563 );
and \U$56002 ( \55977 , \55976 , \55580 );
and \U$56003 ( \55978 , \55545 , \55563 );
or \U$56004 ( \55979 , \55977 , \55978 );
buf \U$56005 ( \55980 , \55979 );
xnor \U$56006 ( \55981 , \55975 , \55980 );
not \U$56007 ( \55982 , \55981 );
buf \U$56008 ( \55983 , \55982 );
xor \U$56009 ( \55984 , \55955 , \55983 );
buf \U$56010 ( \55985 , \55984 );
xor \U$56011 ( \55986 , \55909 , \55985 );
buf \U$56012 ( \55987 , \55986 );
buf \U$56013 ( \55988 , \55987 );
xor \U$56014 ( \55989 , \55452 , \55988 );
xor \U$56015 ( \55990 , \55585 , \55763 );
buf \U$56016 ( \55991 , \55990 );
buf \U$56017 ( \55992 , \55620 );
and \U$56018 ( \55993 , \55991 , \55992 );
not \U$56019 ( \55994 , \55991 );
buf \U$56020 ( \55995 , \55623 );
and \U$56021 ( \55996 , \55994 , \55995 );
nor \U$56022 ( \55997 , \55993 , \55996 );
buf \U$56023 ( \55998 , \55997 );
buf \U$56024 ( \55999 , \55998 );
buf \U$56025 ( \56000 , \48088 );
buf \U$56026 ( \56001 , \48033 );
buf \U$56027 ( \56002 , \48038 );
nor \U$56028 ( \56003 , \56001 , \56002 );
buf \U$56029 ( \56004 , \56003 );
buf \U$56030 ( \56005 , \56004 );
or \U$56031 ( \56006 , \56000 , \56005 );
buf \U$56032 ( \56007 , \48033 );
buf \U$56033 ( \56008 , \48038 );
nand \U$56034 ( \56009 , \56007 , \56008 );
buf \U$56035 ( \56010 , \56009 );
buf \U$56036 ( \56011 , \56010 );
nand \U$56037 ( \56012 , \56006 , \56011 );
buf \U$56038 ( \56013 , \56012 );
buf \U$56039 ( \56014 , \56013 );
buf \U$56040 ( \56015 , \48293 );
not \U$56041 ( \56016 , \56015 );
buf \U$56042 ( \56017 , \48221 );
not \U$56043 ( \56018 , \56017 );
or \U$56044 ( \56019 , \56016 , \56018 );
buf \U$56045 ( \56020 , \48169 );
nand \U$56046 ( \56021 , \56019 , \56020 );
buf \U$56047 ( \56022 , \56021 );
buf \U$56048 ( \56023 , \56022 );
buf \U$56049 ( \56024 , \48221 );
not \U$56050 ( \56025 , \56024 );
buf \U$56051 ( \56026 , \48296 );
nand \U$56052 ( \56027 , \56025 , \56026 );
buf \U$56053 ( \56028 , \56027 );
buf \U$56054 ( \56029 , \56028 );
nand \U$56055 ( \56030 , \56023 , \56029 );
buf \U$56056 ( \56031 , \56030 );
buf \U$56057 ( \56032 , \56031 );
xor \U$56058 ( \56033 , \56014 , \56032 );
buf \U$56059 ( \56034 , \48486 );
not \U$56060 ( \56035 , \56034 );
buf \U$56061 ( \56036 , \48555 );
not \U$56062 ( \56037 , \56036 );
or \U$56063 ( \56038 , \56035 , \56037 );
buf \U$56064 ( \56039 , \48426 );
not \U$56065 ( \56040 , \56039 );
buf \U$56066 ( \56041 , \48552 );
not \U$56067 ( \56042 , \56041 );
or \U$56068 ( \56043 , \56040 , \56042 );
buf \U$56069 ( \56044 , \48478 );
nand \U$56070 ( \56045 , \56043 , \56044 );
buf \U$56071 ( \56046 , \56045 );
buf \U$56072 ( \56047 , \56046 );
nand \U$56073 ( \56048 , \56038 , \56047 );
buf \U$56074 ( \56049 , \56048 );
buf \U$56075 ( \56050 , \56049 );
and \U$56076 ( \56051 , \56033 , \56050 );
and \U$56077 ( \56052 , \56014 , \56032 );
or \U$56078 ( \56053 , \56051 , \56052 );
buf \U$56079 ( \56054 , \56053 );
buf \U$56080 ( \56055 , \56054 );
not \U$56081 ( \56056 , \56055 );
xor \U$56082 ( \56057 , \54473 , \54544 );
xor \U$56083 ( \56058 , \56057 , \54620 );
buf \U$56084 ( \56059 , \56058 );
buf \U$56085 ( \56060 , \56059 );
not \U$56086 ( \56061 , \56060 );
or \U$56087 ( \56062 , \56056 , \56061 );
buf \U$56088 ( \56063 , \56059 );
buf \U$56089 ( \56064 , \56054 );
or \U$56090 ( \56065 , \56063 , \56064 );
xor \U$56091 ( \56066 , \54405 , \54384 );
xor \U$56092 ( \56067 , \56066 , \54461 );
buf \U$56093 ( \56068 , \56067 );
not \U$56094 ( \56069 , \56068 );
buf \U$56095 ( \56070 , \56069 );
not \U$56096 ( \56071 , \56070 );
xor \U$56097 ( \56072 , \54249 , \54265 );
xnor \U$56098 ( \56073 , \56072 , \54288 );
buf \U$56099 ( \56074 , \56073 );
not \U$56100 ( \56075 , \56074 );
buf \U$56101 ( \56076 , \56075 );
not \U$56102 ( \56077 , \56076 );
or \U$56103 ( \56078 , \56071 , \56077 );
not \U$56104 ( \56079 , \56067 );
not \U$56105 ( \56080 , \56073 );
or \U$56106 ( \56081 , \56079 , \56080 );
xor \U$56107 ( \56082 , \55240 , \55243 );
xor \U$56108 ( \56083 , \56082 , \55279 );
buf \U$56109 ( \56084 , \56083 );
nand \U$56110 ( \56085 , \56081 , \56084 );
nand \U$56111 ( \56086 , \56078 , \56085 );
buf \U$56112 ( \56087 , \56086 );
nand \U$56113 ( \56088 , \56065 , \56087 );
buf \U$56114 ( \56089 , \56088 );
buf \U$56115 ( \56090 , \56089 );
nand \U$56116 ( \56091 , \56062 , \56090 );
buf \U$56117 ( \56092 , \56091 );
buf \U$56118 ( \56093 , \56092 );
xor \U$56119 ( \56094 , \55999 , \56093 );
xor \U$56120 ( \56095 , \55608 , \55611 );
xor \U$56121 ( \56096 , \56095 , \55616 );
buf \U$56122 ( \56097 , \56096 );
buf \U$56123 ( \56098 , \56097 );
buf \U$56124 ( \56099 , \48656 );
not \U$56125 ( \56100 , \56099 );
buf \U$56126 ( \56101 , \48673 );
not \U$56127 ( \56102 , \56101 );
or \U$56128 ( \56103 , \56100 , \56102 );
buf \U$56129 ( \56104 , \48659 );
not \U$56130 ( \56105 , \56104 );
buf \U$56131 ( \56106 , \48679 );
not \U$56132 ( \56107 , \56106 );
or \U$56133 ( \56108 , \56105 , \56107 );
buf \U$56134 ( \56109 , \48640 );
nand \U$56135 ( \56110 , \56108 , \56109 );
buf \U$56136 ( \56111 , \56110 );
buf \U$56137 ( \56112 , \56111 );
nand \U$56138 ( \56113 , \56103 , \56112 );
buf \U$56139 ( \56114 , \56113 );
buf \U$56140 ( \56115 , \56114 );
buf \U$56141 ( \56116 , \48601 );
not \U$56142 ( \56117 , \56116 );
buf \U$56143 ( \56118 , \48625 );
not \U$56144 ( \56119 , \56118 );
or \U$56145 ( \56120 , \56117 , \56119 );
buf \U$56146 ( \56121 , \48607 );
nand \U$56147 ( \56122 , \56120 , \56121 );
buf \U$56148 ( \56123 , \56122 );
buf \U$56149 ( \56124 , \56123 );
buf \U$56150 ( \56125 , \48601 );
not \U$56151 ( \56126 , \56125 );
buf \U$56152 ( \56127 , \48622 );
nand \U$56153 ( \56128 , \56126 , \56127 );
buf \U$56154 ( \56129 , \56128 );
buf \U$56155 ( \56130 , \56129 );
nand \U$56156 ( \56131 , \56124 , \56130 );
buf \U$56157 ( \56132 , \56131 );
buf \U$56158 ( \56133 , \56132 );
xor \U$56159 ( \56134 , \56115 , \56133 );
xor \U$56160 ( \56135 , \54322 , \54337 );
xor \U$56161 ( \56136 , \56135 , \54344 );
buf \U$56162 ( \56137 , \56136 );
buf \U$56163 ( \56138 , \56137 );
and \U$56164 ( \56139 , \56134 , \56138 );
and \U$56165 ( \56140 , \56115 , \56133 );
or \U$56166 ( \56141 , \56139 , \56140 );
buf \U$56167 ( \56142 , \56141 );
buf \U$56168 ( \56143 , \56142 );
xor \U$56169 ( \56144 , \56098 , \56143 );
and \U$56170 ( \56145 , \54348 , \54297 );
not \U$56171 ( \56146 , \54348 );
and \U$56172 ( \56147 , \56146 , \54294 );
or \U$56173 ( \56148 , \56145 , \56147 );
buf \U$56174 ( \56149 , \56148 );
buf \U$56175 ( \56150 , \54301 );
and \U$56176 ( \56151 , \56149 , \56150 );
not \U$56177 ( \56152 , \56149 );
buf \U$56178 ( \56153 , \54355 );
and \U$56179 ( \56154 , \56152 , \56153 );
or \U$56180 ( \56155 , \56151 , \56154 );
buf \U$56181 ( \56156 , \56155 );
buf \U$56182 ( \56157 , \56156 );
and \U$56183 ( \56158 , \56144 , \56157 );
and \U$56184 ( \56159 , \56098 , \56143 );
or \U$56185 ( \56160 , \56158 , \56159 );
buf \U$56186 ( \56161 , \56160 );
buf \U$56187 ( \56162 , \56161 );
and \U$56188 ( \56163 , \56094 , \56162 );
and \U$56189 ( \56164 , \55999 , \56093 );
or \U$56190 ( \56165 , \56163 , \56164 );
buf \U$56191 ( \56166 , \56165 );
buf \U$56192 ( \56167 , \56166 );
xor \U$56193 ( \56168 , \55989 , \56167 );
buf \U$56194 ( \56169 , \56168 );
buf \U$56195 ( \56170 , \56169 );
xor \U$56196 ( \56171 , \55307 , \56170 );
buf \U$56197 ( \56172 , \55297 );
buf \U$56198 ( \56173 , \55055 );
and \U$56199 ( \56174 , \56172 , \56173 );
not \U$56200 ( \56175 , \56172 );
buf \U$56201 ( \56176 , \55058 );
and \U$56202 ( \56177 , \56175 , \56176 );
or \U$56203 ( \56178 , \56174 , \56177 );
buf \U$56204 ( \56179 , \56178 );
buf \U$56205 ( \56180 , \56179 );
buf \U$56206 ( \56181 , \55212 );
and \U$56207 ( \56182 , \56180 , \56181 );
not \U$56208 ( \56183 , \56180 );
buf \U$56209 ( \56184 , \55209 );
and \U$56210 ( \56185 , \56183 , \56184 );
nor \U$56211 ( \56186 , \56182 , \56185 );
buf \U$56212 ( \56187 , \56186 );
buf \U$56213 ( \56188 , \56187 );
xor \U$56214 ( \56189 , \54366 , \54362 );
buf \U$56215 ( \56190 , \56189 );
buf \U$56216 ( \56191 , \54624 );
and \U$56217 ( \56192 , \56190 , \56191 );
not \U$56218 ( \56193 , \56190 );
buf \U$56219 ( \56194 , \54627 );
and \U$56220 ( \56195 , \56193 , \56194 );
nor \U$56221 ( \56196 , \56192 , \56195 );
buf \U$56222 ( \56197 , \56196 );
buf \U$56223 ( \56198 , \56197 );
xor \U$56224 ( \56199 , \56188 , \56198 );
xor \U$56225 ( \56200 , \55999 , \56093 );
xor \U$56226 ( \56201 , \56200 , \56162 );
buf \U$56227 ( \56202 , \56201 );
buf \U$56228 ( \56203 , \56202 );
and \U$56229 ( \56204 , \56199 , \56203 );
and \U$56230 ( \56205 , \56188 , \56198 );
or \U$56231 ( \56206 , \56204 , \56205 );
buf \U$56232 ( \56207 , \56206 );
buf \U$56233 ( \56208 , \56207 );
xor \U$56234 ( \56209 , \56171 , \56208 );
buf \U$56235 ( \56210 , \56209 );
buf \U$56236 ( \56211 , \56210 );
buf \U$56237 ( \56212 , \56086 );
buf \U$56238 ( \56213 , \56054 );
xor \U$56239 ( \56214 , \56212 , \56213 );
buf \U$56240 ( \56215 , \56214 );
buf \U$56241 ( \56216 , \56215 );
buf \U$56242 ( \56217 , \56059 );
and \U$56243 ( \56218 , \56216 , \56217 );
not \U$56244 ( \56219 , \56216 );
buf \U$56245 ( \56220 , \56059 );
not \U$56246 ( \56221 , \56220 );
buf \U$56247 ( \56222 , \56221 );
buf \U$56248 ( \56223 , \56222 );
and \U$56249 ( \56224 , \56219 , \56223 );
nor \U$56250 ( \56225 , \56218 , \56224 );
buf \U$56251 ( \56226 , \56225 );
buf \U$56252 ( \56227 , \56226 );
buf \U$56253 ( \56228 , \48028 );
not \U$56254 ( \56229 , \56228 );
buf \U$56255 ( \56230 , \48098 );
not \U$56256 ( \56231 , \56230 );
or \U$56257 ( \56232 , \56229 , \56231 );
buf \U$56258 ( \56233 , \48098 );
buf \U$56259 ( \56234 , \48028 );
or \U$56260 ( \56235 , \56233 , \56234 );
buf \U$56261 ( \56236 , \48104 );
nand \U$56262 ( \56237 , \56235 , \56236 );
buf \U$56263 ( \56238 , \56237 );
buf \U$56264 ( \56239 , \56238 );
nand \U$56265 ( \56240 , \56232 , \56239 );
buf \U$56266 ( \56241 , \56240 );
buf \U$56267 ( \56242 , \56241 );
buf \U$56268 ( \56243 , \48633 );
not \U$56269 ( \56244 , \56243 );
buf \U$56270 ( \56245 , \48683 );
not \U$56271 ( \56246 , \56245 );
or \U$56272 ( \56247 , \56244 , \56246 );
buf \U$56273 ( \56248 , \48562 );
nand \U$56274 ( \56249 , \56247 , \56248 );
buf \U$56275 ( \56250 , \56249 );
buf \U$56276 ( \56251 , \56250 );
buf \U$56277 ( \56252 , \48633 );
not \U$56278 ( \56253 , \56252 );
buf \U$56279 ( \56254 , \48686 );
nand \U$56280 ( \56255 , \56253 , \56254 );
buf \U$56281 ( \56256 , \56255 );
buf \U$56282 ( \56257 , \56256 );
nand \U$56283 ( \56258 , \56251 , \56257 );
buf \U$56284 ( \56259 , \56258 );
buf \U$56285 ( \56260 , \56259 );
xor \U$56286 ( \56261 , \56242 , \56260 );
xor \U$56287 ( \56262 , \56014 , \56032 );
xor \U$56288 ( \56263 , \56262 , \56050 );
buf \U$56289 ( \56264 , \56263 );
buf \U$56290 ( \56265 , \56264 );
and \U$56291 ( \56266 , \56261 , \56265 );
and \U$56292 ( \56267 , \56242 , \56260 );
or \U$56293 ( \56268 , \56266 , \56267 );
buf \U$56294 ( \56269 , \56268 );
buf \U$56295 ( \56270 , \56269 );
xor \U$56296 ( \56271 , \56227 , \56270 );
not \U$56297 ( \56272 , \56070 );
not \U$56298 ( \56273 , \56073 );
or \U$56299 ( \56274 , \56272 , \56273 );
buf \U$56300 ( \56275 , \56076 );
buf \U$56301 ( \56276 , \56067 );
nand \U$56302 ( \56277 , \56275 , \56276 );
buf \U$56303 ( \56278 , \56277 );
nand \U$56304 ( \56279 , \56274 , \56278 );
buf \U$56305 ( \56280 , \56279 );
buf \U$56306 ( \56281 , \56084 );
xor \U$56307 ( \56282 , \56280 , \56281 );
buf \U$56308 ( \56283 , \56282 );
buf \U$56309 ( \56284 , \56283 );
xor \U$56310 ( \56285 , \48304 , \48310 );
and \U$56311 ( \56286 , \56285 , \48333 );
and \U$56312 ( \56287 , \48304 , \48310 );
or \U$56313 ( \56288 , \56286 , \56287 );
buf \U$56314 ( \56289 , \56288 );
buf \U$56315 ( \56290 , \56289 );
xor \U$56316 ( \56291 , \56284 , \56290 );
xor \U$56317 ( \56292 , \54537 , \54476 );
xor \U$56318 ( \56293 , \56292 , \54528 );
buf \U$56319 ( \56294 , \56293 );
xor \U$56320 ( \56295 , \48317 , \48323 );
and \U$56321 ( \56296 , \56295 , \48330 );
and \U$56322 ( \56297 , \48317 , \48323 );
or \U$56323 ( \56298 , \56296 , \56297 );
buf \U$56324 ( \56299 , \56298 );
buf \U$56325 ( \56300 , \56299 );
xor \U$56326 ( \56301 , \56294 , \56300 );
xor \U$56327 ( \56302 , \56115 , \56133 );
xor \U$56328 ( \56303 , \56302 , \56138 );
buf \U$56329 ( \56304 , \56303 );
buf \U$56330 ( \56305 , \56304 );
xor \U$56331 ( \56306 , \56301 , \56305 );
buf \U$56332 ( \56307 , \56306 );
buf \U$56333 ( \56308 , \56307 );
and \U$56334 ( \56309 , \56291 , \56308 );
and \U$56335 ( \56310 , \56284 , \56290 );
or \U$56336 ( \56311 , \56309 , \56310 );
buf \U$56337 ( \56312 , \56311 );
buf \U$56338 ( \56313 , \56312 );
and \U$56339 ( \56314 , \56271 , \56313 );
and \U$56340 ( \56315 , \56227 , \56270 );
or \U$56341 ( \56316 , \56314 , \56315 );
buf \U$56342 ( \56317 , \56316 );
buf \U$56343 ( \56318 , \56317 );
xor \U$56344 ( \56319 , \56188 , \56198 );
xor \U$56345 ( \56320 , \56319 , \56203 );
buf \U$56346 ( \56321 , \56320 );
buf \U$56347 ( \56322 , \56321 );
or \U$56348 ( \56323 , \56318 , \56322 );
xor \U$56349 ( \56324 , \55283 , \55234 );
xor \U$56350 ( \56325 , \56324 , \55291 );
buf \U$56351 ( \56326 , \56325 );
xor \U$56352 ( \56327 , \56294 , \56300 );
and \U$56353 ( \56328 , \56327 , \56305 );
and \U$56354 ( \56329 , \56294 , \56300 );
or \U$56355 ( \56330 , \56328 , \56329 );
buf \U$56356 ( \56331 , \56330 );
buf \U$56357 ( \56332 , \56331 );
xor \U$56358 ( \56333 , \56326 , \56332 );
xor \U$56359 ( \56334 , \56098 , \56143 );
xor \U$56360 ( \56335 , \56334 , \56157 );
buf \U$56361 ( \56336 , \56335 );
buf \U$56362 ( \56337 , \56336 );
and \U$56363 ( \56338 , \56333 , \56337 );
and \U$56364 ( \56339 , \56326 , \56332 );
or \U$56365 ( \56340 , \56338 , \56339 );
buf \U$56366 ( \56341 , \56340 );
buf \U$56367 ( \56342 , \56341 );
nand \U$56368 ( \56343 , \56323 , \56342 );
buf \U$56369 ( \56344 , \56343 );
buf \U$56370 ( \56345 , \56344 );
buf \U$56371 ( \56346 , \56321 );
buf \U$56372 ( \56347 , \56317 );
nand \U$56373 ( \56348 , \56346 , \56347 );
buf \U$56374 ( \56349 , \56348 );
buf \U$56375 ( \56350 , \56349 );
nand \U$56376 ( \56351 , \56345 , \56350 );
buf \U$56377 ( \56352 , \56351 );
buf \U$56378 ( \56353 , \56352 );
or \U$56379 ( \56354 , \56211 , \56353 );
buf \U$56380 ( \56355 , \56354 );
buf \U$56381 ( \56356 , \56355 );
xor \U$56382 ( \56357 , \56326 , \56332 );
xor \U$56383 ( \56358 , \56357 , \56337 );
buf \U$56384 ( \56359 , \56358 );
buf \U$56385 ( \56360 , \56359 );
xor \U$56386 ( \56361 , \48358 , \48375 );
and \U$56387 ( \56362 , \56361 , \48703 );
and \U$56388 ( \56363 , \48358 , \48375 );
or \U$56389 ( \56364 , \56362 , \56363 );
buf \U$56390 ( \56365 , \56364 );
buf \U$56391 ( \56366 , \56365 );
xor \U$56392 ( \56367 , \56242 , \56260 );
xor \U$56393 ( \56368 , \56367 , \56265 );
buf \U$56394 ( \56369 , \56368 );
buf \U$56395 ( \56370 , \56369 );
xor \U$56396 ( \56371 , \56366 , \56370 );
xor \U$56397 ( \56372 , \48106 , \48112 );
and \U$56398 ( \56373 , \56372 , \48336 );
and \U$56399 ( \56374 , \48106 , \48112 );
or \U$56400 ( \56375 , \56373 , \56374 );
buf \U$56401 ( \56376 , \56375 );
buf \U$56402 ( \56377 , \56376 );
and \U$56403 ( \56378 , \56371 , \56377 );
and \U$56404 ( \56379 , \56366 , \56370 );
or \U$56405 ( \56380 , \56378 , \56379 );
buf \U$56406 ( \56381 , \56380 );
buf \U$56407 ( \56382 , \56381 );
xor \U$56408 ( \56383 , \56360 , \56382 );
xor \U$56409 ( \56384 , \56227 , \56270 );
xor \U$56410 ( \56385 , \56384 , \56313 );
buf \U$56411 ( \56386 , \56385 );
buf \U$56412 ( \56387 , \56386 );
xor \U$56413 ( \56388 , \56383 , \56387 );
buf \U$56414 ( \56389 , \56388 );
buf \U$56415 ( \56390 , \56389 );
xor \U$56416 ( \56391 , \56284 , \56290 );
xor \U$56417 ( \56392 , \56391 , \56308 );
buf \U$56418 ( \56393 , \56392 );
buf \U$56419 ( \56394 , \56393 );
xor \U$56420 ( \56395 , \48352 , \48706 );
and \U$56421 ( \56396 , \56395 , \48713 );
and \U$56422 ( \56397 , \48352 , \48706 );
or \U$56423 ( \56398 , \56396 , \56397 );
buf \U$56424 ( \56399 , \56398 );
buf \U$56425 ( \56400 , \56399 );
xor \U$56426 ( \56401 , \56394 , \56400 );
xor \U$56427 ( \56402 , \56366 , \56370 );
xor \U$56428 ( \56403 , \56402 , \56377 );
buf \U$56429 ( \56404 , \56403 );
buf \U$56430 ( \56405 , \56404 );
and \U$56431 ( \56406 , \56401 , \56405 );
and \U$56432 ( \56407 , \56394 , \56400 );
or \U$56433 ( \56408 , \56406 , \56407 );
buf \U$56434 ( \56409 , \56408 );
buf \U$56435 ( \56410 , \56409 );
nor \U$56436 ( \56411 , \56390 , \56410 );
buf \U$56437 ( \56412 , \56411 );
not \U$56438 ( \56413 , \56412 );
buf \U$56439 ( \56414 , \56413 );
xor \U$56440 ( \56415 , \56360 , \56382 );
and \U$56441 ( \56416 , \56415 , \56387 );
and \U$56442 ( \56417 , \56360 , \56382 );
or \U$56443 ( \56418 , \56416 , \56417 );
buf \U$56444 ( \56419 , \56418 );
not \U$56445 ( \56420 , \56419 );
xor \U$56446 ( \56421 , \56341 , \56321 );
xnor \U$56447 ( \56422 , \56421 , \56317 );
nand \U$56448 ( \56423 , \56420 , \56422 );
buf \U$56449 ( \56424 , \56423 );
xor \U$56450 ( \56425 , \56394 , \56400 );
xor \U$56451 ( \56426 , \56425 , \56405 );
buf \U$56452 ( \56427 , \56426 );
buf \U$56453 ( \56428 , \56427 );
xor \U$56454 ( \56429 , \48339 , \48345 );
and \U$56455 ( \56430 , \56429 , \48716 );
and \U$56456 ( \56431 , \48339 , \48345 );
or \U$56457 ( \56432 , \56430 , \56431 );
buf \U$56458 ( \56433 , \56432 );
buf \U$56459 ( \56434 , \56433 );
or \U$56460 ( \56435 , \56428 , \56434 );
buf \U$56461 ( \56436 , \56435 );
buf \U$56462 ( \56437 , \56436 );
nand \U$56463 ( \56438 , \56356 , \56414 , \56424 , \56437 );
buf \U$56464 ( \56439 , \56438 );
buf \U$56465 ( \56440 , \56439 );
not \U$56466 ( \56441 , \56440 );
buf \U$56467 ( \56442 , \56441 );
buf \U$56468 ( \56443 , \56442 );
nand \U$56469 ( \56444 , \53424 , \56443 );
buf \U$56470 ( \56445 , \56444 );
buf \U$56471 ( \56446 , \56445 );
buf \U$56472 ( \56447 , \51433 );
buf \U$56473 ( \56448 , \53257 );
buf \U$56474 ( \56449 , \52871 );
not \U$56475 ( \56450 , \56449 );
buf \U$56476 ( \56451 , \56450 );
buf \U$56477 ( \56452 , \56451 );
buf \U$56478 ( \56453 , \53242 );
not \U$56479 ( \56454 , \56453 );
buf \U$56480 ( \56455 , \56454 );
buf \U$56481 ( \56456 , \56455 );
nand \U$56482 ( \56457 , \56452 , \56456 );
buf \U$56483 ( \56458 , \56457 );
buf \U$56484 ( \56459 , \56458 );
and \U$56485 ( \56460 , \56448 , \56459 );
buf \U$56486 ( \56461 , \56460 );
buf \U$56487 ( \56462 , \56461 );
buf \U$56488 ( \56463 , \53323 );
buf \U$56489 ( \56464 , \53290 );
and \U$56490 ( \56465 , \56462 , \56463 , \56464 );
buf \U$56491 ( \56466 , \56465 );
buf \U$56492 ( \56467 , \56466 );
buf \U$56493 ( \56468 , \51469 );
buf \U$56494 ( \56469 , \51489 );
and \U$56495 ( \56470 , \56447 , \56467 , \56468 , \56469 );
buf \U$56496 ( \56471 , \56470 );
not \U$56497 ( \56472 , \56471 );
nor \U$56498 ( \56473 , \56472 , \56439 );
buf \U$56499 ( \56474 , \56473 );
buf \U$56500 ( \56475 , \49374 );
buf \U$56501 ( \56476 , \52636 );
not \U$56502 ( \56477 , \56476 );
buf \U$56503 ( \56478 , \52645 );
buf \U$56504 ( \56479 , \52626 );
xnor \U$56505 ( \56480 , \56478 , \56479 );
buf \U$56506 ( \56481 , \56480 );
buf \U$56507 ( \56482 , \56481 );
not \U$56508 ( \56483 , \56482 );
or \U$56509 ( \56484 , \56477 , \56483 );
buf \U$56510 ( \56485 , \56481 );
buf \U$56511 ( \56486 , \52636 );
or \U$56512 ( \56487 , \56485 , \56486 );
nand \U$56513 ( \56488 , \56484 , \56487 );
buf \U$56514 ( \56489 , \56488 );
buf \U$56515 ( \56490 , \56489 );
xor \U$56516 ( \56491 , RIc0db188_127, RIc0d8848_39);
buf \U$56517 ( \56492 , \56491 );
not \U$56518 ( \56493 , \56492 );
buf \U$56519 ( \56494 , \46813 );
not \U$56520 ( \56495 , \56494 );
or \U$56521 ( \56496 , \56493 , \56495 );
buf \U$56522 ( \56497 , \52470 );
buf \U$56523 ( \56498 , RIc0db200_128);
nand \U$56524 ( \56499 , \56497 , \56498 );
buf \U$56525 ( \56500 , \56499 );
buf \U$56526 ( \56501 , \56500 );
nand \U$56527 ( \56502 , \56496 , \56501 );
buf \U$56528 ( \56503 , \56502 );
buf \U$56529 ( \56504 , \56503 );
not \U$56530 ( \56505 , \56504 );
buf \U$56531 ( \56506 , RIc0dadc8_119);
buf \U$56532 ( \56507 , RIc0d8c08_47);
xor \U$56533 ( \56508 , \56506 , \56507 );
buf \U$56534 ( \56509 , \56508 );
buf \U$56535 ( \56510 , \56509 );
not \U$56536 ( \56511 , \56510 );
buf \U$56537 ( \56512 , \25542 );
not \U$56538 ( \56513 , \56512 );
or \U$56539 ( \56514 , \56511 , \56513 );
buf \U$56540 ( \56515 , \13953 );
buf \U$56541 ( \56516 , \52732 );
nand \U$56542 ( \56517 , \56515 , \56516 );
buf \U$56543 ( \56518 , \56517 );
buf \U$56544 ( \56519 , \56518 );
nand \U$56545 ( \56520 , \56514 , \56519 );
buf \U$56546 ( \56521 , \56520 );
buf \U$56547 ( \56522 , \56521 );
not \U$56548 ( \56523 , \56522 );
or \U$56549 ( \56524 , \56505 , \56523 );
buf \U$56550 ( \56525 , RIc0d9310_62);
buf \U$56551 ( \56526 , RIc0da738_105);
xor \U$56552 ( \56527 , \56525 , \56526 );
buf \U$56553 ( \56528 , \56527 );
buf \U$56554 ( \56529 , \56528 );
not \U$56555 ( \56530 , \56529 );
buf \U$56556 ( \56531 , \12736 );
not \U$56557 ( \56532 , \56531 );
or \U$56558 ( \56533 , \56530 , \56532 );
buf \U$56559 ( \56534 , \12744 );
buf \U$56560 ( \56535 , \52925 );
nand \U$56561 ( \56536 , \56534 , \56535 );
buf \U$56562 ( \56537 , \56536 );
buf \U$56563 ( \56538 , \56537 );
nand \U$56564 ( \56539 , \56533 , \56538 );
buf \U$56565 ( \56540 , \56539 );
buf \U$56566 ( \56541 , \56540 );
buf \U$56567 ( \56542 , RIc0d9400_64);
buf \U$56568 ( \56543 , RIc0da6c0_104);
or \U$56569 ( \56544 , \56542 , \56543 );
buf \U$56570 ( \56545 , RIc0da738_105);
nand \U$56571 ( \56546 , \56544 , \56545 );
buf \U$56572 ( \56547 , \56546 );
buf \U$56573 ( \56548 , \56547 );
buf \U$56574 ( \56549 , RIc0d9400_64);
buf \U$56575 ( \56550 , RIc0da6c0_104);
nand \U$56576 ( \56551 , \56549 , \56550 );
buf \U$56577 ( \56552 , \56551 );
buf \U$56578 ( \56553 , \56552 );
buf \U$56579 ( \56554 , RIc0da648_103);
and \U$56580 ( \56555 , \56548 , \56553 , \56554 );
buf \U$56581 ( \56556 , \56555 );
buf \U$56582 ( \56557 , \56556 );
nand \U$56583 ( \56558 , \56541 , \56557 );
buf \U$56584 ( \56559 , \56558 );
buf \U$56585 ( \56560 , \56559 );
not \U$56586 ( \56561 , \56560 );
buf \U$56587 ( \56562 , \56561 );
buf \U$56588 ( \56563 , \56562 );
buf \U$56589 ( \56564 , \56521 );
not \U$56590 ( \56565 , \56564 );
buf \U$56591 ( \56566 , \56503 );
not \U$56592 ( \56567 , \56566 );
buf \U$56593 ( \56568 , \56567 );
buf \U$56594 ( \56569 , \56568 );
nand \U$56595 ( \56570 , \56565 , \56569 );
buf \U$56596 ( \56571 , \56570 );
buf \U$56597 ( \56572 , \56571 );
nand \U$56598 ( \56573 , \56563 , \56572 );
buf \U$56599 ( \56574 , \56573 );
buf \U$56600 ( \56575 , \56574 );
nand \U$56601 ( \56576 , \56524 , \56575 );
buf \U$56602 ( \56577 , \56576 );
buf \U$56603 ( \56578 , \56577 );
xor \U$56604 ( \56579 , \52722 , \52744 );
xor \U$56605 ( \56580 , \56579 , \52706 );
buf \U$56606 ( \56581 , \56580 );
xor \U$56607 ( \56582 , \56578 , \56581 );
xor \U$56608 ( \56583 , \52907 , \52918 );
xor \U$56609 ( \56584 , \56583 , \52962 );
buf \U$56610 ( \56585 , \56584 );
buf \U$56611 ( \56586 , \56585 );
and \U$56612 ( \56587 , \56582 , \56586 );
and \U$56613 ( \56588 , \56578 , \56581 );
or \U$56614 ( \56589 , \56587 , \56588 );
buf \U$56615 ( \56590 , \56589 );
buf \U$56616 ( \56591 , \56590 );
xor \U$56617 ( \56592 , \56490 , \56591 );
buf \U$56618 ( \56593 , RIc0d8d70_50);
buf \U$56619 ( \56594 , RIc0dacd8_117);
xor \U$56620 ( \56595 , \56593 , \56594 );
buf \U$56621 ( \56596 , \56595 );
buf \U$56622 ( \56597 , \56596 );
not \U$56623 ( \56598 , \56597 );
buf \U$56624 ( \56599 , \12929 );
not \U$56625 ( \56600 , \56599 );
or \U$56626 ( \56601 , \56598 , \56600 );
buf \U$56627 ( \56602 , \12937 );
buf \U$56628 ( \56603 , \53005 );
nand \U$56629 ( \56604 , \56602 , \56603 );
buf \U$56630 ( \56605 , \56604 );
buf \U$56631 ( \56606 , \56605 );
nand \U$56632 ( \56607 , \56601 , \56606 );
buf \U$56633 ( \56608 , \56607 );
buf \U$56634 ( \56609 , \56608 );
buf \U$56635 ( \56610 , RIc0d8c80_48);
buf \U$56636 ( \56611 , RIc0dadc8_119);
xor \U$56637 ( \56612 , \56610 , \56611 );
buf \U$56638 ( \56613 , \56612 );
buf \U$56639 ( \56614 , \56613 );
not \U$56640 ( \56615 , \56614 );
buf \U$56641 ( \56616 , \23985 );
not \U$56642 ( \56617 , \56616 );
or \U$56643 ( \56618 , \56615 , \56617 );
buf \U$56644 ( \56619 , \13953 );
buf \U$56645 ( \56620 , \56509 );
nand \U$56646 ( \56621 , \56619 , \56620 );
buf \U$56647 ( \56622 , \56621 );
buf \U$56648 ( \56623 , \56622 );
nand \U$56649 ( \56624 , \56618 , \56623 );
buf \U$56650 ( \56625 , \56624 );
buf \U$56651 ( \56626 , \56625 );
or \U$56652 ( \56627 , \56609 , \56626 );
buf \U$56653 ( \56628 , RIc0d9040_56);
buf \U$56654 ( \56629 , RIc0daa08_111);
xor \U$56655 ( \56630 , \56628 , \56629 );
buf \U$56656 ( \56631 , \56630 );
buf \U$56657 ( \56632 , \56631 );
not \U$56658 ( \56633 , \56632 );
buf \U$56659 ( \56634 , \18306 );
not \U$56660 ( \56635 , \56634 );
or \U$56661 ( \56636 , \56633 , \56635 );
buf \U$56662 ( \56637 , \52988 );
not \U$56663 ( \56638 , \56637 );
buf \U$56664 ( \56639 , \45728 );
nand \U$56665 ( \56640 , \56638 , \56639 );
buf \U$56666 ( \56641 , \56640 );
buf \U$56667 ( \56642 , \56641 );
nand \U$56668 ( \56643 , \56636 , \56642 );
buf \U$56669 ( \56644 , \56643 );
buf \U$56670 ( \56645 , \56644 );
nand \U$56671 ( \56646 , \56627 , \56645 );
buf \U$56672 ( \56647 , \56646 );
buf \U$56673 ( \56648 , \56647 );
buf \U$56674 ( \56649 , \56608 );
buf \U$56675 ( \56650 , \56625 );
nand \U$56676 ( \56651 , \56649 , \56650 );
buf \U$56677 ( \56652 , \56651 );
buf \U$56678 ( \56653 , \56652 );
nand \U$56679 ( \56654 , \56648 , \56653 );
buf \U$56680 ( \56655 , \56654 );
buf \U$56681 ( \56656 , \56655 );
not \U$56682 ( \56657 , \56656 );
buf \U$56683 ( \56658 , \56657 );
buf \U$56684 ( \56659 , \56658 );
not \U$56685 ( \56660 , \56659 );
buf \U$56686 ( \56661 , RIc0d8b90_46);
buf \U$56687 ( \56662 , RIc0daeb8_121);
xor \U$56688 ( \56663 , \56661 , \56662 );
buf \U$56689 ( \56664 , \56663 );
buf \U$56690 ( \56665 , \56664 );
not \U$56691 ( \56666 , \56665 );
buf \U$56692 ( \56667 , \13310 );
not \U$56693 ( \56668 , \56667 );
or \U$56694 ( \56669 , \56666 , \56668 );
buf \U$56695 ( \56670 , \53127 );
not \U$56696 ( \56671 , \56670 );
buf \U$56697 ( \56672 , \16386 );
nand \U$56698 ( \56673 , \56671 , \56672 );
buf \U$56699 ( \56674 , \56673 );
buf \U$56700 ( \56675 , \56674 );
nand \U$56701 ( \56676 , \56669 , \56675 );
buf \U$56702 ( \56677 , \56676 );
buf \U$56703 ( \56678 , \56677 );
not \U$56704 ( \56679 , \56678 );
buf \U$56705 ( \56680 , RIc0d9220_60);
buf \U$56706 ( \56681 , RIc0da828_107);
xor \U$56707 ( \56682 , \56680 , \56681 );
buf \U$56708 ( \56683 , \56682 );
buf \U$56709 ( \56684 , \56683 );
not \U$56710 ( \56685 , \56684 );
buf \U$56711 ( \56686 , \34202 );
not \U$56712 ( \56687 , \56686 );
or \U$56713 ( \56688 , \56685 , \56687 );
buf \U$56714 ( \56689 , \16071 );
buf \U$56715 ( \56690 , \53063 );
nand \U$56716 ( \56691 , \56689 , \56690 );
buf \U$56717 ( \56692 , \56691 );
buf \U$56718 ( \56693 , \56692 );
nand \U$56719 ( \56694 , \56688 , \56693 );
buf \U$56720 ( \56695 , \56694 );
buf \U$56721 ( \56696 , \56695 );
not \U$56722 ( \56697 , \56696 );
or \U$56723 ( \56698 , \56679 , \56697 );
buf \U$56724 ( \56699 , \56695 );
buf \U$56725 ( \56700 , \56677 );
or \U$56726 ( \56701 , \56699 , \56700 );
buf \U$56727 ( \56702 , RIc0d8aa0_44);
buf \U$56728 ( \56703 , RIc0dafa8_123);
xor \U$56729 ( \56704 , \56702 , \56703 );
buf \U$56730 ( \56705 , \56704 );
buf \U$56731 ( \56706 , \56705 );
not \U$56732 ( \56707 , \56706 );
buf \U$56733 ( \56708 , \47037 );
not \U$56734 ( \56709 , \56708 );
or \U$56735 ( \56710 , \56707 , \56709 );
buf \U$56736 ( \56711 , \16692 );
buf \U$56737 ( \56712 , \53090 );
nand \U$56738 ( \56713 , \56711 , \56712 );
buf \U$56739 ( \56714 , \56713 );
buf \U$56740 ( \56715 , \56714 );
nand \U$56741 ( \56716 , \56710 , \56715 );
buf \U$56742 ( \56717 , \56716 );
buf \U$56743 ( \56718 , \56717 );
nand \U$56744 ( \56719 , \56701 , \56718 );
buf \U$56745 ( \56720 , \56719 );
buf \U$56746 ( \56721 , \56720 );
nand \U$56747 ( \56722 , \56698 , \56721 );
buf \U$56748 ( \56723 , \56722 );
buf \U$56749 ( \56724 , \56723 );
not \U$56750 ( \56725 , \56724 );
buf \U$56751 ( \56726 , \56725 );
buf \U$56752 ( \56727 , \56726 );
not \U$56753 ( \56728 , \56727 );
or \U$56754 ( \56729 , \56660 , \56728 );
buf \U$56755 ( \56730 , RIc0d8e60_52);
buf \U$56756 ( \56731 , RIc0dabe8_115);
xor \U$56757 ( \56732 , \56730 , \56731 );
buf \U$56758 ( \56733 , \56732 );
buf \U$56759 ( \56734 , \56733 );
not \U$56760 ( \56735 , \56734 );
buf \U$56761 ( \56736 , \14186 );
not \U$56762 ( \56737 , \56736 );
or \U$56763 ( \56738 , \56735 , \56737 );
buf \U$56764 ( \56739 , \14690 );
buf \U$56765 ( \56740 , \52944 );
nand \U$56766 ( \56741 , \56739 , \56740 );
buf \U$56767 ( \56742 , \56741 );
buf \U$56768 ( \56743 , \56742 );
nand \U$56769 ( \56744 , \56738 , \56743 );
buf \U$56770 ( \56745 , \56744 );
buf \U$56771 ( \56746 , \56745 );
not \U$56772 ( \56747 , \56746 );
buf \U$56773 ( \56748 , RIc0d9130_58);
buf \U$56774 ( \56749 , RIc0da918_109);
xor \U$56775 ( \56750 , \56748 , \56749 );
buf \U$56776 ( \56751 , \56750 );
buf \U$56777 ( \56752 , \56751 );
not \U$56778 ( \56753 , \56752 );
buf \U$56779 ( \56754 , \20759 );
not \U$56780 ( \56755 , \56754 );
or \U$56781 ( \56756 , \56753 , \56755 );
buf \U$56782 ( \56757 , \16232 );
buf \U$56783 ( \56758 , \53028 );
nand \U$56784 ( \56759 , \56757 , \56758 );
buf \U$56785 ( \56760 , \56759 );
buf \U$56786 ( \56761 , \56760 );
nand \U$56787 ( \56762 , \56756 , \56761 );
buf \U$56788 ( \56763 , \56762 );
buf \U$56789 ( \56764 , \56763 );
not \U$56790 ( \56765 , \56764 );
or \U$56791 ( \56766 , \56747 , \56765 );
buf \U$56792 ( \56767 , \56763 );
buf \U$56793 ( \56768 , \56745 );
or \U$56794 ( \56769 , \56767 , \56768 );
buf \U$56795 ( \56770 , RIc0da648_103);
buf \U$56796 ( \56771 , RIc0d9400_64);
and \U$56797 ( \56772 , \56770 , \56771 );
not \U$56798 ( \56773 , \56770 );
buf \U$56799 ( \56774 , \43843 );
and \U$56800 ( \56775 , \56773 , \56774 );
nor \U$56801 ( \56776 , \56772 , \56775 );
buf \U$56802 ( \56777 , \56776 );
buf \U$56803 ( \56778 , \56777 );
not \U$56804 ( \56779 , \56778 );
buf \U$56805 ( \56780 , \17405 );
not \U$56806 ( \56781 , \56780 );
or \U$56807 ( \56782 , \56779 , \56781 );
buf \U$56808 ( \56783 , \13712 );
buf \U$56809 ( \56784 , \53045 );
nand \U$56810 ( \56785 , \56783 , \56784 );
buf \U$56811 ( \56786 , \56785 );
buf \U$56812 ( \56787 , \56786 );
nand \U$56813 ( \56788 , \56782 , \56787 );
buf \U$56814 ( \56789 , \56788 );
buf \U$56815 ( \56790 , \56789 );
nand \U$56816 ( \56791 , \56769 , \56790 );
buf \U$56817 ( \56792 , \56791 );
buf \U$56818 ( \56793 , \56792 );
nand \U$56819 ( \56794 , \56766 , \56793 );
buf \U$56820 ( \56795 , \56794 );
buf \U$56821 ( \56796 , \56795 );
nand \U$56822 ( \56797 , \56729 , \56796 );
buf \U$56823 ( \56798 , \56797 );
buf \U$56824 ( \56799 , \56798 );
buf \U$56825 ( \56800 , \56723 );
buf \U$56826 ( \56801 , \56655 );
nand \U$56827 ( \56802 , \56800 , \56801 );
buf \U$56828 ( \56803 , \56802 );
buf \U$56829 ( \56804 , \56803 );
nand \U$56830 ( \56805 , \56799 , \56804 );
buf \U$56831 ( \56806 , \56805 );
buf \U$56832 ( \56807 , \56806 );
not \U$56833 ( \56808 , \56807 );
buf \U$56834 ( \56809 , \56808 );
buf \U$56835 ( \56810 , \56809 );
not \U$56836 ( \56811 , \56810 );
buf \U$56837 ( \56812 , \53152 );
buf \U$56838 ( \56813 , \53080 );
xor \U$56839 ( \56814 , \56812 , \56813 );
buf \U$56840 ( \56815 , \56814 );
buf \U$56841 ( \56816 , \56815 );
buf \U$56842 ( \56817 , \53025 );
xnor \U$56843 ( \56818 , \56816 , \56817 );
buf \U$56844 ( \56819 , \56818 );
buf \U$56845 ( \56820 , \56819 );
not \U$56846 ( \56821 , \56820 );
or \U$56847 ( \56822 , \56811 , \56821 );
buf \U$56848 ( \56823 , RIc0daaf8_113);
buf \U$56849 ( \56824 , RIc0d8f50_54);
xor \U$56850 ( \56825 , \56823 , \56824 );
buf \U$56851 ( \56826 , \56825 );
buf \U$56852 ( \56827 , \56826 );
not \U$56853 ( \56828 , \56827 );
buf \U$56854 ( \56829 , \33224 );
not \U$56855 ( \56830 , \56829 );
or \U$56856 ( \56831 , \56828 , \56830 );
buf \U$56857 ( \56832 , \12410 );
buf \U$56858 ( \56833 , \53107 );
nand \U$56859 ( \56834 , \56832 , \56833 );
buf \U$56860 ( \56835 , \56834 );
buf \U$56861 ( \56836 , \56835 );
nand \U$56862 ( \56837 , \56831 , \56836 );
buf \U$56863 ( \56838 , \56837 );
buf \U$56864 ( \56839 , \56838 );
buf \U$56865 ( \56840 , \18008 );
not \U$56866 ( \56841 , \56840 );
buf \U$56867 ( \56842 , RIc0d88c0_40);
buf \U$56868 ( \56843 , RIc0db188_127);
xor \U$56869 ( \56844 , \56842 , \56843 );
buf \U$56870 ( \56845 , \56844 );
buf \U$56871 ( \56846 , \56845 );
not \U$56872 ( \56847 , \56846 );
buf \U$56873 ( \56848 , \56847 );
buf \U$56874 ( \56849 , \56848 );
not \U$56875 ( \56850 , \56849 );
and \U$56876 ( \56851 , \56841 , \56850 );
buf \U$56877 ( \56852 , \56491 );
buf \U$56878 ( \56853 , RIc0db200_128);
and \U$56879 ( \56854 , \56852 , \56853 );
nor \U$56880 ( \56855 , \56851 , \56854 );
buf \U$56881 ( \56856 , \56855 );
buf \U$56882 ( \56857 , \56856 );
not \U$56883 ( \56858 , \56857 );
buf \U$56884 ( \56859 , \56858 );
buf \U$56885 ( \56860 , \56859 );
nand \U$56886 ( \56861 , \56839 , \56860 );
buf \U$56887 ( \56862 , \56861 );
buf \U$56888 ( \56863 , \56862 );
buf \U$56889 ( \56864 , \56838 );
buf \U$56890 ( \56865 , \56859 );
or \U$56891 ( \56866 , \56864 , \56865 );
buf \U$56892 ( \56867 , RIc0d89b0_42);
buf \U$56893 ( \56868 , RIc0db098_125);
xnor \U$56894 ( \56869 , \56867 , \56868 );
buf \U$56895 ( \56870 , \56869 );
buf \U$56896 ( \56871 , \56870 );
not \U$56897 ( \56872 , \56871 );
buf \U$56898 ( \56873 , \56872 );
buf \U$56899 ( \56874 , \56873 );
not \U$56900 ( \56875 , \56874 );
buf \U$56901 ( \56876 , \17995 );
not \U$56902 ( \56877 , \56876 );
or \U$56903 ( \56878 , \56875 , \56877 );
buf \U$56904 ( \56879 , \13465 );
buf \U$56905 ( \56880 , \52969 );
nand \U$56906 ( \56881 , \56879 , \56880 );
buf \U$56907 ( \56882 , \56881 );
buf \U$56908 ( \56883 , \56882 );
nand \U$56909 ( \56884 , \56878 , \56883 );
buf \U$56910 ( \56885 , \56884 );
buf \U$56911 ( \56886 , \56885 );
nand \U$56912 ( \56887 , \56866 , \56886 );
buf \U$56913 ( \56888 , \56887 );
buf \U$56914 ( \56889 , \56888 );
nand \U$56915 ( \56890 , \56863 , \56889 );
buf \U$56916 ( \56891 , \56890 );
buf \U$56917 ( \56892 , \56891 );
xor \U$56918 ( \56893 , \52924 , \52939 );
xor \U$56919 ( \56894 , \56893 , \52957 );
buf \U$56920 ( \56895 , \56894 );
buf \U$56921 ( \56896 , \56895 );
xor \U$56922 ( \56897 , \56892 , \56896 );
buf \U$56923 ( \56898 , \53119 );
not \U$56924 ( \56899 , \56898 );
buf \U$56925 ( \56900 , \53138 );
not \U$56926 ( \56901 , \56900 );
or \U$56927 ( \56902 , \56899 , \56901 );
buf \U$56928 ( \56903 , \53119 );
buf \U$56929 ( \56904 , \53138 );
or \U$56930 ( \56905 , \56903 , \56904 );
nand \U$56931 ( \56906 , \56902 , \56905 );
buf \U$56932 ( \56907 , \56906 );
xor \U$56933 ( \56908 , \53102 , \56907 );
buf \U$56934 ( \56909 , \56908 );
and \U$56935 ( \56910 , \56897 , \56909 );
and \U$56936 ( \56911 , \56892 , \56896 );
or \U$56937 ( \56912 , \56910 , \56911 );
buf \U$56938 ( \56913 , \56912 );
buf \U$56939 ( \56914 , \56913 );
nand \U$56940 ( \56915 , \56822 , \56914 );
buf \U$56941 ( \56916 , \56915 );
buf \U$56942 ( \56917 , \56916 );
buf \U$56943 ( \56918 , \56819 );
not \U$56944 ( \56919 , \56918 );
buf \U$56945 ( \56920 , \56919 );
buf \U$56946 ( \56921 , \56920 );
buf \U$56947 ( \56922 , \56806 );
nand \U$56948 ( \56923 , \56921 , \56922 );
buf \U$56949 ( \56924 , \56923 );
buf \U$56950 ( \56925 , \56924 );
nand \U$56951 ( \56926 , \56917 , \56925 );
buf \U$56952 ( \56927 , \56926 );
buf \U$56953 ( \56928 , \56927 );
and \U$56954 ( \56929 , \56592 , \56928 );
and \U$56955 ( \56930 , \56490 , \56591 );
or \U$56956 ( \56931 , \56929 , \56930 );
buf \U$56957 ( \56932 , \56931 );
buf \U$56958 ( \56933 , \56932 );
not \U$56959 ( \56934 , \56933 );
xor \U$56960 ( \56935 , \52981 , \52999 );
xor \U$56961 ( \56936 , \56935 , \53017 );
buf \U$56962 ( \56937 , \56936 );
not \U$56963 ( \56938 , \56937 );
buf \U$56964 ( \56939 , \56568 );
not \U$56965 ( \56940 , \56939 );
buf \U$56966 ( \56941 , \56521 );
not \U$56967 ( \56942 , \56941 );
or \U$56968 ( \56943 , \56940 , \56942 );
buf \U$56969 ( \56944 , \56521 );
buf \U$56970 ( \56945 , \56568 );
or \U$56971 ( \56946 , \56944 , \56945 );
nand \U$56972 ( \56947 , \56943 , \56946 );
buf \U$56973 ( \56948 , \56947 );
buf \U$56974 ( \56949 , \56948 );
buf \U$56975 ( \56950 , \56559 );
and \U$56976 ( \56951 , \56949 , \56950 );
not \U$56977 ( \56952 , \56949 );
buf \U$56978 ( \56953 , \56562 );
and \U$56979 ( \56954 , \56952 , \56953 );
nor \U$56980 ( \56955 , \56951 , \56954 );
buf \U$56981 ( \56956 , \56955 );
buf \U$56982 ( \56957 , \56956 );
not \U$56983 ( \56958 , \56957 );
or \U$56984 ( \56959 , \56938 , \56958 );
xor \U$56985 ( \56960 , \53041 , \53058 );
xor \U$56986 ( \56961 , \56960 , \53076 );
buf \U$56987 ( \56962 , \56961 );
buf \U$56988 ( \56963 , \56962 );
nand \U$56989 ( \56964 , \56959 , \56963 );
buf \U$56990 ( \56965 , \56964 );
buf \U$56991 ( \56966 , \56965 );
buf \U$56992 ( \56967 , \56956 );
not \U$56993 ( \56968 , \56967 );
buf \U$56994 ( \56969 , \56936 );
not \U$56995 ( \56970 , \56969 );
buf \U$56996 ( \56971 , \56970 );
buf \U$56997 ( \56972 , \56971 );
nand \U$56998 ( \56973 , \56968 , \56972 );
buf \U$56999 ( \56974 , \56973 );
buf \U$57000 ( \56975 , \56974 );
nand \U$57001 ( \56976 , \56966 , \56975 );
buf \U$57002 ( \56977 , \56976 );
buf \U$57003 ( \56978 , \56977 );
xor \U$57004 ( \56979 , \53178 , \53199 );
xor \U$57005 ( \56980 , \56979 , \53203 );
buf \U$57006 ( \56981 , \56980 );
buf \U$57007 ( \56982 , \56981 );
xor \U$57008 ( \56983 , \56978 , \56982 );
xor \U$57009 ( \56984 , \56578 , \56581 );
xor \U$57010 ( \56985 , \56984 , \56586 );
buf \U$57011 ( \56986 , \56985 );
buf \U$57012 ( \56987 , \56986 );
and \U$57013 ( \56988 , \56983 , \56987 );
and \U$57014 ( \56989 , \56978 , \56982 );
or \U$57015 ( \56990 , \56988 , \56989 );
buf \U$57016 ( \56991 , \56990 );
buf \U$57017 ( \56992 , \56991 );
xor \U$57018 ( \56993 , \52888 , \52967 );
xor \U$57019 ( \56994 , \56993 , \53159 );
buf \U$57020 ( \56995 , \56994 );
buf \U$57021 ( \56996 , \56995 );
or \U$57022 ( \56997 , \56992 , \56996 );
xor \U$57023 ( \56998 , \53169 , \53173 );
xor \U$57024 ( \56999 , \56998 , \53208 );
buf \U$57025 ( \57000 , \56999 );
buf \U$57026 ( \57001 , \57000 );
nand \U$57027 ( \57002 , \56997 , \57001 );
buf \U$57028 ( \57003 , \57002 );
buf \U$57029 ( \57004 , \57003 );
buf \U$57030 ( \57005 , \56991 );
buf \U$57031 ( \57006 , \56995 );
nand \U$57032 ( \57007 , \57005 , \57006 );
buf \U$57033 ( \57008 , \57007 );
buf \U$57034 ( \57009 , \57008 );
nand \U$57035 ( \57010 , \57004 , \57009 );
buf \U$57036 ( \57011 , \57010 );
buf \U$57037 ( \57012 , \57011 );
not \U$57038 ( \57013 , \57012 );
buf \U$57039 ( \57014 , \57013 );
buf \U$57040 ( \57015 , \57014 );
not \U$57041 ( \57016 , \57015 );
or \U$57042 ( \57017 , \56934 , \57016 );
buf \U$57043 ( \57018 , \57014 );
buf \U$57044 ( \57019 , \56932 );
or \U$57045 ( \57020 , \57018 , \57019 );
nand \U$57046 ( \57021 , \57017 , \57020 );
buf \U$57047 ( \57022 , \57021 );
buf \U$57048 ( \57023 , \57022 );
not \U$57049 ( \57024 , \57023 );
buf \U$57050 ( \57025 , \52605 );
not \U$57051 ( \57026 , \57025 );
buf \U$57052 ( \57027 , \52439 );
not \U$57053 ( \57028 , \57027 );
buf \U$57054 ( \57029 , \52598 );
not \U$57055 ( \57030 , \57029 );
or \U$57056 ( \57031 , \57028 , \57030 );
buf \U$57057 ( \57032 , \52598 );
buf \U$57058 ( \57033 , \52439 );
or \U$57059 ( \57034 , \57032 , \57033 );
nand \U$57060 ( \57035 , \57031 , \57034 );
buf \U$57061 ( \57036 , \57035 );
buf \U$57062 ( \57037 , \57036 );
not \U$57063 ( \57038 , \57037 );
buf \U$57064 ( \57039 , \57038 );
buf \U$57065 ( \57040 , \57039 );
not \U$57066 ( \57041 , \57040 );
or \U$57067 ( \57042 , \57026 , \57041 );
buf \U$57068 ( \57043 , \52605 );
not \U$57069 ( \57044 , \57043 );
buf \U$57070 ( \57045 , \57036 );
nand \U$57071 ( \57046 , \57044 , \57045 );
buf \U$57072 ( \57047 , \57046 );
buf \U$57073 ( \57048 , \57047 );
nand \U$57074 ( \57049 , \57042 , \57048 );
buf \U$57075 ( \57050 , \57049 );
buf \U$57076 ( \57051 , \57050 );
xor \U$57077 ( \57052 , \52623 , \52652 );
xor \U$57078 ( \57053 , \57052 , \52820 );
buf \U$57079 ( \57054 , \57053 );
buf \U$57080 ( \57055 , \57054 );
not \U$57081 ( \57056 , \57055 );
buf \U$57082 ( \57057 , \57056 );
buf \U$57083 ( \57058 , \57057 );
and \U$57084 ( \57059 , \57051 , \57058 );
not \U$57085 ( \57060 , \57051 );
buf \U$57086 ( \57061 , \57054 );
and \U$57087 ( \57062 , \57060 , \57061 );
or \U$57088 ( \57063 , \57059 , \57062 );
buf \U$57089 ( \57064 , \57063 );
buf \U$57090 ( \57065 , \57064 );
xor \U$57091 ( \57066 , \52884 , \53164 );
xor \U$57092 ( \57067 , \57066 , \53213 );
buf \U$57093 ( \57068 , \57067 );
buf \U$57094 ( \57069 , \57068 );
xnor \U$57095 ( \57070 , \57065 , \57069 );
buf \U$57096 ( \57071 , \57070 );
buf \U$57097 ( \57072 , \57071 );
not \U$57098 ( \57073 , \57072 );
and \U$57099 ( \57074 , \57024 , \57073 );
buf \U$57100 ( \57075 , \57022 );
buf \U$57101 ( \57076 , \57071 );
and \U$57102 ( \57077 , \57075 , \57076 );
nor \U$57103 ( \57078 , \57074 , \57077 );
buf \U$57104 ( \57079 , \57078 );
buf \U$57105 ( \57080 , \57079 );
buf \U$57106 ( \57081 , \56809 );
not \U$57107 ( \57082 , \57081 );
buf \U$57108 ( \57083 , \56913 );
not \U$57109 ( \57084 , \57083 );
or \U$57110 ( \57085 , \57082 , \57084 );
buf \U$57111 ( \57086 , \56913 );
buf \U$57112 ( \57087 , \56809 );
or \U$57113 ( \57088 , \57086 , \57087 );
nand \U$57114 ( \57089 , \57085 , \57088 );
buf \U$57115 ( \57090 , \57089 );
buf \U$57116 ( \57091 , \57090 );
buf \U$57117 ( \57092 , \56819 );
and \U$57118 ( \57093 , \57091 , \57092 );
not \U$57119 ( \57094 , \57091 );
buf \U$57120 ( \57095 , \56920 );
and \U$57121 ( \57096 , \57094 , \57095 );
nor \U$57122 ( \57097 , \57093 , \57096 );
buf \U$57123 ( \57098 , \57097 );
buf \U$57124 ( \57099 , \57098 );
not \U$57125 ( \57100 , \57099 );
buf \U$57126 ( \57101 , \57100 );
not \U$57127 ( \57102 , \57101 );
buf \U$57128 ( \57103 , \56540 );
buf \U$57129 ( \57104 , \56556 );
xor \U$57130 ( \57105 , \57103 , \57104 );
buf \U$57131 ( \57106 , \57105 );
buf \U$57132 ( \57107 , \57106 );
buf \U$57133 ( \57108 , RIc0d8b18_45);
buf \U$57134 ( \57109 , RIc0dafa8_123);
xor \U$57135 ( \57110 , \57108 , \57109 );
buf \U$57136 ( \57111 , \57110 );
buf \U$57137 ( \57112 , \57111 );
not \U$57138 ( \57113 , \57112 );
buf \U$57139 ( \57114 , \14982 );
not \U$57140 ( \57115 , \57114 );
or \U$57141 ( \57116 , \57113 , \57115 );
buf \U$57142 ( \57117 , \16692 );
buf \U$57143 ( \57118 , \56705 );
nand \U$57144 ( \57119 , \57117 , \57118 );
buf \U$57145 ( \57120 , \57119 );
buf \U$57146 ( \57121 , \57120 );
nand \U$57147 ( \57122 , \57116 , \57121 );
buf \U$57148 ( \57123 , \57122 );
buf \U$57149 ( \57124 , \57123 );
not \U$57150 ( \57125 , \57124 );
xnor \U$57151 ( \57126 , RIc0dabe8_115, RIc0d8ed8_53);
buf \U$57152 ( \57127 , \57126 );
not \U$57153 ( \57128 , \57127 );
buf \U$57154 ( \57129 , \57128 );
buf \U$57155 ( \57130 , \57129 );
not \U$57156 ( \57131 , \57130 );
buf \U$57157 ( \57132 , \27743 );
not \U$57158 ( \57133 , \57132 );
or \U$57159 ( \57134 , \57131 , \57133 );
buf \U$57160 ( \57135 , \14690 );
buf \U$57161 ( \57136 , \56733 );
nand \U$57162 ( \57137 , \57135 , \57136 );
buf \U$57163 ( \57138 , \57137 );
buf \U$57164 ( \57139 , \57138 );
nand \U$57165 ( \57140 , \57134 , \57139 );
buf \U$57166 ( \57141 , \57140 );
buf \U$57167 ( \57142 , \57141 );
not \U$57168 ( \57143 , \57142 );
or \U$57169 ( \57144 , \57125 , \57143 );
buf \U$57170 ( \57145 , \57123 );
buf \U$57171 ( \57146 , \57141 );
or \U$57172 ( \57147 , \57145 , \57146 );
xor \U$57173 ( \57148 , RIc0dacd8_117, RIc0d8de8_51);
buf \U$57174 ( \57149 , \57148 );
not \U$57175 ( \57150 , \57149 );
buf \U$57176 ( \57151 , \13146 );
not \U$57177 ( \57152 , \57151 );
or \U$57178 ( \57153 , \57150 , \57152 );
buf \U$57179 ( \57154 , \12937 );
buf \U$57180 ( \57155 , \56596 );
nand \U$57181 ( \57156 , \57154 , \57155 );
buf \U$57182 ( \57157 , \57156 );
buf \U$57183 ( \57158 , \57157 );
nand \U$57184 ( \57159 , \57153 , \57158 );
buf \U$57185 ( \57160 , \57159 );
buf \U$57186 ( \57161 , \57160 );
nand \U$57187 ( \57162 , \57147 , \57161 );
buf \U$57188 ( \57163 , \57162 );
buf \U$57189 ( \57164 , \57163 );
nand \U$57190 ( \57165 , \57144 , \57164 );
buf \U$57191 ( \57166 , \57165 );
buf \U$57192 ( \57167 , \57166 );
xor \U$57193 ( \57168 , \57107 , \57167 );
xor \U$57194 ( \57169 , RIc0daa08_111, RIc0d90b8_57);
buf \U$57195 ( \57170 , \57169 );
not \U$57196 ( \57171 , \57170 );
buf \U$57197 ( \57172 , \14346 );
not \U$57198 ( \57173 , \57172 );
or \U$57199 ( \57174 , \57171 , \57173 );
buf \U$57200 ( \57175 , \14353 );
buf \U$57201 ( \57176 , \56631 );
nand \U$57202 ( \57177 , \57175 , \57176 );
buf \U$57203 ( \57178 , \57177 );
buf \U$57204 ( \57179 , \57178 );
nand \U$57205 ( \57180 , \57174 , \57179 );
buf \U$57206 ( \57181 , \57180 );
buf \U$57207 ( \57182 , \57181 );
buf \U$57208 ( \57183 , RIc0da738_105);
buf \U$57209 ( \57184 , RIc0d9388_63);
and \U$57210 ( \57185 , \57183 , \57184 );
not \U$57211 ( \57186 , \57183 );
buf \U$57212 ( \57187 , \43939 );
and \U$57213 ( \57188 , \57186 , \57187 );
nor \U$57214 ( \57189 , \57185 , \57188 );
buf \U$57215 ( \57190 , \57189 );
buf \U$57216 ( \57191 , \57190 );
not \U$57217 ( \57192 , \57191 );
buf \U$57218 ( \57193 , \12736 );
not \U$57219 ( \57194 , \57193 );
or \U$57220 ( \57195 , \57192 , \57194 );
buf \U$57221 ( \57196 , \21880 );
buf \U$57222 ( \57197 , \56528 );
nand \U$57223 ( \57198 , \57196 , \57197 );
buf \U$57224 ( \57199 , \57198 );
buf \U$57225 ( \57200 , \57199 );
nand \U$57226 ( \57201 , \57195 , \57200 );
buf \U$57227 ( \57202 , \57201 );
buf \U$57228 ( \57203 , \57202 );
xor \U$57229 ( \57204 , \57182 , \57203 );
buf \U$57230 ( \57205 , RIc0da918_109);
buf \U$57231 ( \57206 , RIc0d91a8_59);
xor \U$57232 ( \57207 , \57205 , \57206 );
buf \U$57233 ( \57208 , \57207 );
buf \U$57234 ( \57209 , \57208 );
not \U$57235 ( \57210 , \57209 );
buf \U$57236 ( \57211 , \14210 );
not \U$57237 ( \57212 , \57211 );
or \U$57238 ( \57213 , \57210 , \57212 );
buf \U$57239 ( \57214 , \20211 );
buf \U$57240 ( \57215 , \56751 );
nand \U$57241 ( \57216 , \57214 , \57215 );
buf \U$57242 ( \57217 , \57216 );
buf \U$57243 ( \57218 , \57217 );
nand \U$57244 ( \57219 , \57213 , \57218 );
buf \U$57245 ( \57220 , \57219 );
buf \U$57246 ( \57221 , \57220 );
and \U$57247 ( \57222 , \57204 , \57221 );
and \U$57248 ( \57223 , \57182 , \57203 );
or \U$57249 ( \57224 , \57222 , \57223 );
buf \U$57250 ( \57225 , \57224 );
buf \U$57251 ( \57226 , \57225 );
and \U$57252 ( \57227 , \57168 , \57226 );
and \U$57253 ( \57228 , \57107 , \57167 );
or \U$57254 ( \57229 , \57227 , \57228 );
buf \U$57255 ( \57230 , \57229 );
buf \U$57256 ( \57231 , \57230 );
not \U$57257 ( \57232 , \57231 );
buf \U$57258 ( \57233 , RIc0d8938_41);
buf \U$57259 ( \57234 , RIc0db188_127);
xor \U$57260 ( \57235 , \57233 , \57234 );
buf \U$57261 ( \57236 , \57235 );
buf \U$57262 ( \57237 , \57236 );
not \U$57263 ( \57238 , \57237 );
buf \U$57264 ( \57239 , \15609 );
not \U$57265 ( \57240 , \57239 );
or \U$57266 ( \57241 , \57238 , \57240 );
buf \U$57267 ( \57242 , \56845 );
buf \U$57268 ( \57243 , RIc0db200_128);
nand \U$57269 ( \57244 , \57242 , \57243 );
buf \U$57270 ( \57245 , \57244 );
buf \U$57271 ( \57246 , \57245 );
nand \U$57272 ( \57247 , \57241 , \57246 );
buf \U$57273 ( \57248 , \57247 );
buf \U$57274 ( \57249 , \57248 );
not \U$57275 ( \57250 , \57249 );
buf \U$57276 ( \57251 , RIc0daaf8_113);
buf \U$57277 ( \57252 , RIc0d8fc8_55);
xor \U$57278 ( \57253 , \57251 , \57252 );
buf \U$57279 ( \57254 , \57253 );
buf \U$57280 ( \57255 , \57254 );
not \U$57281 ( \57256 , \57255 );
buf \U$57282 ( \57257 , \28776 );
not \U$57283 ( \57258 , \57257 );
or \U$57284 ( \57259 , \57256 , \57258 );
buf \U$57285 ( \57260 , \12410 );
buf \U$57286 ( \57261 , \56826 );
nand \U$57287 ( \57262 , \57260 , \57261 );
buf \U$57288 ( \57263 , \57262 );
buf \U$57289 ( \57264 , \57263 );
nand \U$57290 ( \57265 , \57259 , \57264 );
buf \U$57291 ( \57266 , \57265 );
buf \U$57292 ( \57267 , \57266 );
not \U$57293 ( \57268 , \57267 );
or \U$57294 ( \57269 , \57250 , \57268 );
buf \U$57295 ( \57270 , \57266 );
buf \U$57296 ( \57271 , \57248 );
or \U$57297 ( \57272 , \57270 , \57271 );
buf \U$57298 ( \57273 , RIc0d8cf8_49);
buf \U$57299 ( \57274 , RIc0dadc8_119);
xor \U$57300 ( \57275 , \57273 , \57274 );
buf \U$57301 ( \57276 , \57275 );
buf \U$57302 ( \57277 , \57276 );
not \U$57303 ( \57278 , \57277 );
buf \U$57304 ( \57279 , \23985 );
not \U$57305 ( \57280 , \57279 );
or \U$57306 ( \57281 , \57278 , \57280 );
buf \U$57307 ( \57282 , \13953 );
buf \U$57308 ( \57283 , \56613 );
nand \U$57309 ( \57284 , \57282 , \57283 );
buf \U$57310 ( \57285 , \57284 );
buf \U$57311 ( \57286 , \57285 );
nand \U$57312 ( \57287 , \57281 , \57286 );
buf \U$57313 ( \57288 , \57287 );
buf \U$57314 ( \57289 , \57288 );
nand \U$57315 ( \57290 , \57272 , \57289 );
buf \U$57316 ( \57291 , \57290 );
buf \U$57317 ( \57292 , \57291 );
nand \U$57318 ( \57293 , \57269 , \57292 );
buf \U$57319 ( \57294 , \57293 );
buf \U$57320 ( \57295 , \57294 );
buf \U$57321 ( \57296 , \13048 );
buf \U$57322 ( \57297 , RIc0d9400_64);
and \U$57323 ( \57298 , \57296 , \57297 );
buf \U$57324 ( \57299 , \57298 );
buf \U$57325 ( \57300 , \57299 );
buf \U$57326 ( \57301 , RIc0d9298_61);
buf \U$57327 ( \57302 , RIc0da828_107);
xor \U$57328 ( \57303 , \57301 , \57302 );
buf \U$57329 ( \57304 , \57303 );
buf \U$57330 ( \57305 , \57304 );
not \U$57331 ( \57306 , \57305 );
buf \U$57332 ( \57307 , \28794 );
not \U$57333 ( \57308 , \57307 );
or \U$57334 ( \57309 , \57306 , \57308 );
buf \U$57335 ( \57310 , \12342 );
buf \U$57336 ( \57311 , \56683 );
nand \U$57337 ( \57312 , \57310 , \57311 );
buf \U$57338 ( \57313 , \57312 );
buf \U$57339 ( \57314 , \57313 );
nand \U$57340 ( \57315 , \57309 , \57314 );
buf \U$57341 ( \57316 , \57315 );
buf \U$57342 ( \57317 , \57316 );
xor \U$57343 ( \57318 , \57300 , \57317 );
buf \U$57344 ( \57319 , \46459 );
xnor \U$57345 ( \57320 , RIc0db098_125, RIc0d8a28_43);
buf \U$57346 ( \57321 , \57320 );
or \U$57347 ( \57322 , \57319 , \57321 );
buf \U$57348 ( \57323 , \22744 );
buf \U$57349 ( \57324 , \56870 );
or \U$57350 ( \57325 , \57323 , \57324 );
nand \U$57351 ( \57326 , \57322 , \57325 );
buf \U$57352 ( \57327 , \57326 );
buf \U$57353 ( \57328 , \57327 );
and \U$57354 ( \57329 , \57318 , \57328 );
and \U$57355 ( \57330 , \57300 , \57317 );
or \U$57356 ( \57331 , \57329 , \57330 );
buf \U$57357 ( \57332 , \57331 );
buf \U$57358 ( \57333 , \57332 );
xor \U$57359 ( \57334 , \57295 , \57333 );
xor \U$57360 ( \57335 , \56608 , \56625 );
xor \U$57361 ( \57336 , \57335 , \56644 );
buf \U$57362 ( \57337 , \57336 );
and \U$57363 ( \57338 , \57334 , \57337 );
and \U$57364 ( \57339 , \57295 , \57333 );
or \U$57365 ( \57340 , \57338 , \57339 );
buf \U$57366 ( \57341 , \57340 );
buf \U$57367 ( \57342 , \57341 );
not \U$57368 ( \57343 , \57342 );
or \U$57369 ( \57344 , \57232 , \57343 );
buf \U$57370 ( \57345 , \57341 );
buf \U$57371 ( \57346 , \57230 );
or \U$57372 ( \57347 , \57345 , \57346 );
buf \U$57373 ( \57348 , \56856 );
buf \U$57374 ( \57349 , \56838 );
xor \U$57375 ( \57350 , \57348 , \57349 );
buf \U$57376 ( \57351 , \56885 );
xnor \U$57377 ( \57352 , \57350 , \57351 );
buf \U$57378 ( \57353 , \57352 );
buf \U$57379 ( \57354 , \57353 );
xor \U$57380 ( \57355 , \56745 , \56789 );
xor \U$57381 ( \57356 , \57355 , \56763 );
buf \U$57382 ( \57357 , \57356 );
xor \U$57383 ( \57358 , \57354 , \57357 );
buf \U$57384 ( \57359 , \56695 );
buf \U$57385 ( \57360 , \56677 );
xor \U$57386 ( \57361 , \57359 , \57360 );
buf \U$57387 ( \57362 , \57361 );
buf \U$57388 ( \57363 , \57362 );
buf \U$57389 ( \57364 , \56717 );
xor \U$57390 ( \57365 , \57363 , \57364 );
buf \U$57391 ( \57366 , \57365 );
buf \U$57392 ( \57367 , \57366 );
and \U$57393 ( \57368 , \57358 , \57367 );
and \U$57394 ( \57369 , \57354 , \57357 );
or \U$57395 ( \57370 , \57368 , \57369 );
buf \U$57396 ( \57371 , \57370 );
buf \U$57397 ( \57372 , \57371 );
nand \U$57398 ( \57373 , \57347 , \57372 );
buf \U$57399 ( \57374 , \57373 );
buf \U$57400 ( \57375 , \57374 );
nand \U$57401 ( \57376 , \57344 , \57375 );
buf \U$57402 ( \57377 , \57376 );
not \U$57403 ( \57378 , \57377 );
or \U$57404 ( \57379 , \57102 , \57378 );
buf \U$57405 ( \57380 , \57377 );
not \U$57406 ( \57381 , \57380 );
buf \U$57407 ( \57382 , \57381 );
buf \U$57408 ( \57383 , \57382 );
not \U$57409 ( \57384 , \57383 );
buf \U$57410 ( \57385 , \57098 );
not \U$57411 ( \57386 , \57385 );
or \U$57412 ( \57387 , \57384 , \57386 );
buf \U$57413 ( \57388 , \56655 );
not \U$57414 ( \57389 , \57388 );
buf \U$57415 ( \57390 , \56795 );
buf \U$57416 ( \57391 , \56723 );
and \U$57417 ( \57392 , \57390 , \57391 );
not \U$57418 ( \57393 , \57390 );
buf \U$57419 ( \57394 , \56726 );
and \U$57420 ( \57395 , \57393 , \57394 );
nor \U$57421 ( \57396 , \57392 , \57395 );
buf \U$57422 ( \57397 , \57396 );
buf \U$57423 ( \57398 , \57397 );
not \U$57424 ( \57399 , \57398 );
buf \U$57425 ( \57400 , \57399 );
buf \U$57426 ( \57401 , \57400 );
not \U$57427 ( \57402 , \57401 );
or \U$57428 ( \57403 , \57389 , \57402 );
buf \U$57429 ( \57404 , \57397 );
buf \U$57430 ( \57405 , \56658 );
nand \U$57431 ( \57406 , \57404 , \57405 );
buf \U$57432 ( \57407 , \57406 );
buf \U$57433 ( \57408 , \57407 );
nand \U$57434 ( \57409 , \57403 , \57408 );
buf \U$57435 ( \57410 , \57409 );
buf \U$57436 ( \57411 , \57410 );
not \U$57437 ( \57412 , \57411 );
buf \U$57438 ( \57413 , \56962 );
not \U$57439 ( \57414 , \57413 );
buf \U$57440 ( \57415 , \56956 );
not \U$57441 ( \57416 , \57415 );
or \U$57442 ( \57417 , \57414 , \57416 );
buf \U$57443 ( \57418 , \56956 );
buf \U$57444 ( \57419 , \56962 );
or \U$57445 ( \57420 , \57418 , \57419 );
nand \U$57446 ( \57421 , \57417 , \57420 );
buf \U$57447 ( \57422 , \57421 );
buf \U$57448 ( \57423 , \57422 );
buf \U$57449 ( \57424 , \56971 );
and \U$57450 ( \57425 , \57423 , \57424 );
not \U$57451 ( \57426 , \57423 );
buf \U$57452 ( \57427 , \56936 );
and \U$57453 ( \57428 , \57426 , \57427 );
nor \U$57454 ( \57429 , \57425 , \57428 );
buf \U$57455 ( \57430 , \57429 );
buf \U$57456 ( \57431 , \57430 );
not \U$57457 ( \57432 , \57431 );
or \U$57458 ( \57433 , \57412 , \57432 );
buf \U$57459 ( \57434 , \57430 );
buf \U$57460 ( \57435 , \57410 );
or \U$57461 ( \57436 , \57434 , \57435 );
xor \U$57462 ( \57437 , \56892 , \56896 );
xor \U$57463 ( \57438 , \57437 , \56909 );
buf \U$57464 ( \57439 , \57438 );
buf \U$57465 ( \57440 , \57439 );
nand \U$57466 ( \57441 , \57436 , \57440 );
buf \U$57467 ( \57442 , \57441 );
buf \U$57468 ( \57443 , \57442 );
nand \U$57469 ( \57444 , \57433 , \57443 );
buf \U$57470 ( \57445 , \57444 );
buf \U$57471 ( \57446 , \57445 );
nand \U$57472 ( \57447 , \57387 , \57446 );
buf \U$57473 ( \57448 , \57447 );
nand \U$57474 ( \57449 , \57379 , \57448 );
buf \U$57475 ( \57450 , \57449 );
xor \U$57476 ( \57451 , \56490 , \56591 );
xor \U$57477 ( \57452 , \57451 , \56928 );
buf \U$57478 ( \57453 , \57452 );
buf \U$57479 ( \57454 , \57453 );
xor \U$57480 ( \57455 , \57450 , \57454 );
buf \U$57481 ( \57456 , \56995 );
buf \U$57482 ( \57457 , \57000 );
xor \U$57483 ( \57458 , \57456 , \57457 );
buf \U$57484 ( \57459 , \56991 );
xor \U$57485 ( \57460 , \57458 , \57459 );
buf \U$57486 ( \57461 , \57460 );
buf \U$57487 ( \57462 , \57461 );
and \U$57488 ( \57463 , \57455 , \57462 );
and \U$57489 ( \57464 , \57450 , \57454 );
or \U$57490 ( \57465 , \57463 , \57464 );
buf \U$57491 ( \57466 , \57465 );
buf \U$57492 ( \57467 , \57466 );
not \U$57493 ( \57468 , \57467 );
buf \U$57494 ( \57469 , \57468 );
buf \U$57495 ( \57470 , \57469 );
nand \U$57496 ( \57471 , \57080 , \57470 );
buf \U$57497 ( \57472 , \57471 );
buf \U$57498 ( \57473 , \57472 );
xor \U$57499 ( \57474 , \57450 , \57454 );
xor \U$57500 ( \57475 , \57474 , \57462 );
buf \U$57501 ( \57476 , \57475 );
buf \U$57502 ( \57477 , \57476 );
not \U$57503 ( \57478 , \57477 );
buf \U$57504 ( \57479 , \57478 );
buf \U$57505 ( \57480 , \57479 );
buf \U$57506 ( \57481 , \47570 );
buf \U$57507 ( \57482 , RIc0d8c08_47);
buf \U$57508 ( \57483 , RIc0daeb8_121);
xnor \U$57509 ( \57484 , \57482 , \57483 );
buf \U$57510 ( \57485 , \57484 );
buf \U$57511 ( \57486 , \57485 );
or \U$57512 ( \57487 , \57481 , \57486 );
buf \U$57513 ( \57488 , \45558 );
buf \U$57514 ( \57489 , \56664 );
not \U$57515 ( \57490 , \57489 );
buf \U$57516 ( \57491 , \57490 );
buf \U$57517 ( \57492 , \57491 );
or \U$57518 ( \57493 , \57488 , \57492 );
nand \U$57519 ( \57494 , \57487 , \57493 );
buf \U$57520 ( \57495 , \57494 );
buf \U$57521 ( \57496 , \57495 );
buf \U$57522 ( \57497 , RIc0da828_107);
buf \U$57523 ( \57498 , RIc0d9310_62);
xor \U$57524 ( \57499 , \57497 , \57498 );
buf \U$57525 ( \57500 , \57499 );
buf \U$57526 ( \57501 , \57500 );
not \U$57527 ( \57502 , \57501 );
buf \U$57528 ( \57503 , \19414 );
not \U$57529 ( \57504 , \57503 );
or \U$57530 ( \57505 , \57502 , \57504 );
buf \U$57531 ( \57506 , \12342 );
buf \U$57532 ( \57507 , \57304 );
nand \U$57533 ( \57508 , \57506 , \57507 );
buf \U$57534 ( \57509 , \57508 );
buf \U$57535 ( \57510 , \57509 );
nand \U$57536 ( \57511 , \57505 , \57510 );
buf \U$57537 ( \57512 , \57511 );
buf \U$57538 ( \57513 , \57512 );
not \U$57539 ( \57514 , \57513 );
buf \U$57540 ( \57515 , RIc0d9400_64);
buf \U$57541 ( \57516 , RIc0da7b0_106);
or \U$57542 ( \57517 , \57515 , \57516 );
buf \U$57543 ( \57518 , RIc0da828_107);
nand \U$57544 ( \57519 , \57517 , \57518 );
buf \U$57545 ( \57520 , \57519 );
buf \U$57546 ( \57521 , \57520 );
buf \U$57547 ( \57522 , RIc0d9400_64);
buf \U$57548 ( \57523 , RIc0da7b0_106);
nand \U$57549 ( \57524 , \57522 , \57523 );
buf \U$57550 ( \57525 , \57524 );
buf \U$57551 ( \57526 , \57525 );
buf \U$57552 ( \57527 , RIc0da738_105);
nand \U$57553 ( \57528 , \57521 , \57526 , \57527 );
buf \U$57554 ( \57529 , \57528 );
buf \U$57555 ( \57530 , \57529 );
nor \U$57556 ( \57531 , \57514 , \57530 );
buf \U$57557 ( \57532 , \57531 );
buf \U$57558 ( \57533 , \57532 );
xor \U$57559 ( \57534 , \57496 , \57533 );
buf \U$57560 ( \57535 , RIc0d89b0_42);
buf \U$57561 ( \57536 , RIc0db188_127);
xor \U$57562 ( \57537 , \57535 , \57536 );
buf \U$57563 ( \57538 , \57537 );
buf \U$57564 ( \57539 , \57538 );
not \U$57565 ( \57540 , \57539 );
buf \U$57566 ( \57541 , \15609 );
not \U$57567 ( \57542 , \57541 );
or \U$57568 ( \57543 , \57540 , \57542 );
buf \U$57569 ( \57544 , \57236 );
buf \U$57570 ( \57545 , RIc0db200_128);
nand \U$57571 ( \57546 , \57544 , \57545 );
buf \U$57572 ( \57547 , \57546 );
buf \U$57573 ( \57548 , \57547 );
nand \U$57574 ( \57549 , \57543 , \57548 );
buf \U$57575 ( \57550 , \57549 );
buf \U$57576 ( \57551 , \57550 );
not \U$57577 ( \57552 , \57551 );
buf \U$57578 ( \57553 , RIc0d9220_60);
buf \U$57579 ( \57554 , RIc0da918_109);
xor \U$57580 ( \57555 , \57553 , \57554 );
buf \U$57581 ( \57556 , \57555 );
buf \U$57582 ( \57557 , \57556 );
not \U$57583 ( \57558 , \57557 );
buf \U$57584 ( \57559 , \21959 );
not \U$57585 ( \57560 , \57559 );
or \U$57586 ( \57561 , \57558 , \57560 );
buf \U$57587 ( \57562 , \20211 );
buf \U$57588 ( \57563 , \57208 );
nand \U$57589 ( \57564 , \57562 , \57563 );
buf \U$57590 ( \57565 , \57564 );
buf \U$57591 ( \57566 , \57565 );
nand \U$57592 ( \57567 , \57561 , \57566 );
buf \U$57593 ( \57568 , \57567 );
buf \U$57594 ( \57569 , \57568 );
not \U$57595 ( \57570 , \57569 );
or \U$57596 ( \57571 , \57552 , \57570 );
buf \U$57597 ( \57572 , \57568 );
buf \U$57598 ( \57573 , \57550 );
or \U$57599 ( \57574 , \57572 , \57573 );
buf \U$57600 ( \57575 , RIc0d8b90_46);
buf \U$57601 ( \57576 , RIc0dafa8_123);
xnor \U$57602 ( \57577 , \57575 , \57576 );
buf \U$57603 ( \57578 , \57577 );
buf \U$57604 ( \57579 , \57578 );
not \U$57605 ( \57580 , \57579 );
buf \U$57606 ( \57581 , \57580 );
buf \U$57607 ( \57582 , \57581 );
not \U$57608 ( \57583 , \57582 );
buf \U$57609 ( \57584 , \47037 );
not \U$57610 ( \57585 , \57584 );
or \U$57611 ( \57586 , \57583 , \57585 );
buf \U$57612 ( \57587 , \14278 );
buf \U$57613 ( \57588 , \57111 );
nand \U$57614 ( \57589 , \57587 , \57588 );
buf \U$57615 ( \57590 , \57589 );
buf \U$57616 ( \57591 , \57590 );
nand \U$57617 ( \57592 , \57586 , \57591 );
buf \U$57618 ( \57593 , \57592 );
buf \U$57619 ( \57594 , \57593 );
nand \U$57620 ( \57595 , \57574 , \57594 );
buf \U$57621 ( \57596 , \57595 );
buf \U$57622 ( \57597 , \57596 );
nand \U$57623 ( \57598 , \57571 , \57597 );
buf \U$57624 ( \57599 , \57598 );
buf \U$57625 ( \57600 , \57599 );
and \U$57626 ( \57601 , \57534 , \57600 );
and \U$57627 ( \57602 , \57496 , \57533 );
or \U$57628 ( \57603 , \57601 , \57602 );
buf \U$57629 ( \57604 , \57603 );
buf \U$57630 ( \57605 , \57604 );
xor \U$57631 ( \57606 , \57266 , \57248 );
buf \U$57632 ( \57607 , \57606 );
buf \U$57633 ( \57608 , \57288 );
xnor \U$57634 ( \57609 , \57607 , \57608 );
buf \U$57635 ( \57610 , \57609 );
buf \U$57636 ( \57611 , \57610 );
not \U$57637 ( \57612 , \57611 );
buf \U$57638 ( \57613 , \14681 );
not \U$57639 ( \57614 , \57613 );
buf \U$57640 ( \57615 , RIc0dabe8_115);
buf \U$57641 ( \57616 , RIc0d8f50_54);
xnor \U$57642 ( \57617 , \57615 , \57616 );
buf \U$57643 ( \57618 , \57617 );
buf \U$57644 ( \57619 , \57618 );
not \U$57645 ( \57620 , \57619 );
and \U$57646 ( \57621 , \57614 , \57620 );
buf \U$57647 ( \57622 , \29865 );
buf \U$57648 ( \57623 , \57126 );
nor \U$57649 ( \57624 , \57622 , \57623 );
buf \U$57650 ( \57625 , \57624 );
buf \U$57651 ( \57626 , \57625 );
nor \U$57652 ( \57627 , \57621 , \57626 );
buf \U$57653 ( \57628 , \57627 );
buf \U$57654 ( \57629 , \57628 );
not \U$57655 ( \57630 , \57629 );
buf \U$57656 ( \57631 , RIc0d8e60_52);
buf \U$57657 ( \57632 , RIc0dacd8_117);
xor \U$57658 ( \57633 , \57631 , \57632 );
buf \U$57659 ( \57634 , \57633 );
buf \U$57660 ( \57635 , \57634 );
not \U$57661 ( \57636 , \57635 );
buf \U$57662 ( \57637 , \12929 );
not \U$57663 ( \57638 , \57637 );
or \U$57664 ( \57639 , \57636 , \57638 );
buf \U$57665 ( \57640 , \22356 );
buf \U$57666 ( \57641 , \57148 );
nand \U$57667 ( \57642 , \57640 , \57641 );
buf \U$57668 ( \57643 , \57642 );
buf \U$57669 ( \57644 , \57643 );
nand \U$57670 ( \57645 , \57639 , \57644 );
buf \U$57671 ( \57646 , \57645 );
buf \U$57672 ( \57647 , \57646 );
not \U$57673 ( \57648 , \57647 );
buf \U$57674 ( \57649 , \57648 );
buf \U$57675 ( \57650 , \57649 );
not \U$57676 ( \57651 , \57650 );
or \U$57677 ( \57652 , \57630 , \57651 );
buf \U$57678 ( \57653 , RIc0d8d70_50);
buf \U$57679 ( \57654 , RIc0dadc8_119);
xor \U$57680 ( \57655 , \57653 , \57654 );
buf \U$57681 ( \57656 , \57655 );
buf \U$57682 ( \57657 , \57656 );
not \U$57683 ( \57658 , \57657 );
buf \U$57684 ( \57659 , \13949 );
not \U$57685 ( \57660 , \57659 );
or \U$57686 ( \57661 , \57658 , \57660 );
buf \U$57687 ( \57662 , \13953 );
buf \U$57688 ( \57663 , \57276 );
nand \U$57689 ( \57664 , \57662 , \57663 );
buf \U$57690 ( \57665 , \57664 );
buf \U$57691 ( \57666 , \57665 );
nand \U$57692 ( \57667 , \57661 , \57666 );
buf \U$57693 ( \57668 , \57667 );
buf \U$57694 ( \57669 , \57668 );
nand \U$57695 ( \57670 , \57652 , \57669 );
buf \U$57696 ( \57671 , \57670 );
buf \U$57697 ( \57672 , \57671 );
buf \U$57698 ( \57673 , \57628 );
not \U$57699 ( \57674 , \57673 );
buf \U$57700 ( \57675 , \57646 );
nand \U$57701 ( \57676 , \57674 , \57675 );
buf \U$57702 ( \57677 , \57676 );
buf \U$57703 ( \57678 , \57677 );
nand \U$57704 ( \57679 , \57672 , \57678 );
buf \U$57705 ( \57680 , \57679 );
buf \U$57706 ( \57681 , \57680 );
not \U$57707 ( \57682 , \57681 );
buf \U$57708 ( \57683 , \57682 );
buf \U$57709 ( \57684 , \57683 );
not \U$57710 ( \57685 , \57684 );
or \U$57711 ( \57686 , \57612 , \57685 );
not \U$57712 ( \57687 , \14468 );
buf \U$57713 ( \57688 , RIc0d8aa0_44);
buf \U$57714 ( \57689 , RIc0db098_125);
xnor \U$57715 ( \57690 , \57688 , \57689 );
buf \U$57716 ( \57691 , \57690 );
not \U$57717 ( \57692 , \57691 );
and \U$57718 ( \57693 , \57687 , \57692 );
buf \U$57719 ( \57694 , \18699 );
buf \U$57720 ( \57695 , \57320 );
nor \U$57721 ( \57696 , \57694 , \57695 );
buf \U$57722 ( \57697 , \57696 );
nor \U$57723 ( \57698 , \57693 , \57697 );
buf \U$57724 ( \57699 , \57698 );
not \U$57725 ( \57700 , \57699 );
not \U$57726 ( \57701 , \33303 );
buf \U$57727 ( \57702 , RIc0d9130_58);
buf \U$57728 ( \57703 , RIc0daa08_111);
xnor \U$57729 ( \57704 , \57702 , \57703 );
buf \U$57730 ( \57705 , \57704 );
not \U$57731 ( \57706 , \57705 );
and \U$57732 ( \57707 , \57701 , \57706 );
and \U$57733 ( \57708 , \14106 , \57169 );
nor \U$57734 ( \57709 , \57707 , \57708 );
buf \U$57735 ( \57710 , \57709 );
not \U$57736 ( \57711 , \57710 );
or \U$57737 ( \57712 , \57700 , \57711 );
buf \U$57738 ( \57713 , RIc0d9400_64);
buf \U$57739 ( \57714 , RIc0da738_105);
xor \U$57740 ( \57715 , \57713 , \57714 );
buf \U$57741 ( \57716 , \57715 );
buf \U$57742 ( \57717 , \57716 );
not \U$57743 ( \57718 , \57717 );
buf \U$57744 ( \57719 , \12736 );
not \U$57745 ( \57720 , \57719 );
or \U$57746 ( \57721 , \57718 , \57720 );
buf \U$57747 ( \57722 , \15653 );
buf \U$57748 ( \57723 , \57190 );
nand \U$57749 ( \57724 , \57722 , \57723 );
buf \U$57750 ( \57725 , \57724 );
buf \U$57751 ( \57726 , \57725 );
nand \U$57752 ( \57727 , \57721 , \57726 );
buf \U$57753 ( \57728 , \57727 );
buf \U$57754 ( \57729 , \57728 );
nand \U$57755 ( \57730 , \57712 , \57729 );
buf \U$57756 ( \57731 , \57730 );
buf \U$57757 ( \57732 , \57731 );
buf \U$57758 ( \57733 , \57709 );
not \U$57759 ( \57734 , \57733 );
buf \U$57760 ( \57735 , \57734 );
buf \U$57761 ( \57736 , \57735 );
buf \U$57762 ( \57737 , \57698 );
not \U$57763 ( \57738 , \57737 );
buf \U$57764 ( \57739 , \57738 );
buf \U$57765 ( \57740 , \57739 );
nand \U$57766 ( \57741 , \57736 , \57740 );
buf \U$57767 ( \57742 , \57741 );
buf \U$57768 ( \57743 , \57742 );
and \U$57769 ( \57744 , \57732 , \57743 );
buf \U$57770 ( \57745 , \57744 );
buf \U$57771 ( \57746 , \57745 );
not \U$57772 ( \57747 , \57746 );
buf \U$57773 ( \57748 , \57747 );
buf \U$57774 ( \57749 , \57748 );
nand \U$57775 ( \57750 , \57686 , \57749 );
buf \U$57776 ( \57751 , \57750 );
buf \U$57777 ( \57752 , \57751 );
buf \U$57778 ( \57753 , \57610 );
not \U$57779 ( \57754 , \57753 );
buf \U$57780 ( \57755 , \57680 );
nand \U$57781 ( \57756 , \57754 , \57755 );
buf \U$57782 ( \57757 , \57756 );
buf \U$57783 ( \57758 , \57757 );
nand \U$57784 ( \57759 , \57752 , \57758 );
buf \U$57785 ( \57760 , \57759 );
buf \U$57786 ( \57761 , \57760 );
xor \U$57787 ( \57762 , \57605 , \57761 );
xor \U$57788 ( \57763 , \57295 , \57333 );
xor \U$57789 ( \57764 , \57763 , \57337 );
buf \U$57790 ( \57765 , \57764 );
buf \U$57791 ( \57766 , \57765 );
and \U$57792 ( \57767 , \57762 , \57766 );
and \U$57793 ( \57768 , \57605 , \57761 );
or \U$57794 ( \57769 , \57767 , \57768 );
buf \U$57795 ( \57770 , \57769 );
buf \U$57796 ( \57771 , \57770 );
xor \U$57797 ( \57772 , \57107 , \57167 );
xor \U$57798 ( \57773 , \57772 , \57226 );
buf \U$57799 ( \57774 , \57773 );
buf \U$57800 ( \57775 , \57774 );
xor \U$57801 ( \57776 , \57300 , \57317 );
xor \U$57802 ( \57777 , \57776 , \57328 );
buf \U$57803 ( \57778 , \57777 );
buf \U$57804 ( \57779 , \57778 );
xor \U$57805 ( \57780 , \57182 , \57203 );
xor \U$57806 ( \57781 , \57780 , \57221 );
buf \U$57807 ( \57782 , \57781 );
buf \U$57808 ( \57783 , \57782 );
xor \U$57809 ( \57784 , \57779 , \57783 );
xor \U$57810 ( \57785 , \57123 , \57160 );
xor \U$57811 ( \57786 , \57785 , \57141 );
buf \U$57812 ( \57787 , \57786 );
and \U$57813 ( \57788 , \57784 , \57787 );
and \U$57814 ( \57789 , \57779 , \57783 );
or \U$57815 ( \57790 , \57788 , \57789 );
buf \U$57816 ( \57791 , \57790 );
buf \U$57817 ( \57792 , \57791 );
xor \U$57818 ( \57793 , \57775 , \57792 );
xor \U$57819 ( \57794 , \57354 , \57357 );
xor \U$57820 ( \57795 , \57794 , \57367 );
buf \U$57821 ( \57796 , \57795 );
buf \U$57822 ( \57797 , \57796 );
and \U$57823 ( \57798 , \57793 , \57797 );
and \U$57824 ( \57799 , \57775 , \57792 );
or \U$57825 ( \57800 , \57798 , \57799 );
buf \U$57826 ( \57801 , \57800 );
buf \U$57827 ( \57802 , \57801 );
xor \U$57828 ( \57803 , \57771 , \57802 );
buf \U$57829 ( \57804 , \57371 );
not \U$57830 ( \57805 , \57804 );
xnor \U$57831 ( \57806 , \57341 , \57230 );
buf \U$57832 ( \57807 , \57806 );
not \U$57833 ( \57808 , \57807 );
or \U$57834 ( \57809 , \57805 , \57808 );
buf \U$57835 ( \57810 , \57806 );
buf \U$57836 ( \57811 , \57371 );
or \U$57837 ( \57812 , \57810 , \57811 );
nand \U$57838 ( \57813 , \57809 , \57812 );
buf \U$57839 ( \57814 , \57813 );
buf \U$57840 ( \57815 , \57814 );
and \U$57841 ( \57816 , \57803 , \57815 );
and \U$57842 ( \57817 , \57771 , \57802 );
or \U$57843 ( \57818 , \57816 , \57817 );
buf \U$57844 ( \57819 , \57818 );
buf \U$57845 ( \57820 , \57819 );
not \U$57846 ( \57821 , \57820 );
buf \U$57847 ( \57822 , \57821 );
buf \U$57848 ( \57823 , \57822 );
not \U$57849 ( \57824 , \57823 );
buf \U$57850 ( \57825 , \57377 );
buf \U$57851 ( \57826 , \57445 );
xor \U$57852 ( \57827 , \57825 , \57826 );
buf \U$57853 ( \57828 , \57101 );
xnor \U$57854 ( \57829 , \57827 , \57828 );
buf \U$57855 ( \57830 , \57829 );
buf \U$57856 ( \57831 , \57830 );
not \U$57857 ( \57832 , \57831 );
or \U$57858 ( \57833 , \57824 , \57832 );
xor \U$57859 ( \57834 , \56978 , \56982 );
xor \U$57860 ( \57835 , \57834 , \56987 );
buf \U$57861 ( \57836 , \57835 );
buf \U$57862 ( \57837 , \57836 );
nand \U$57863 ( \57838 , \57833 , \57837 );
buf \U$57864 ( \57839 , \57838 );
buf \U$57865 ( \57840 , \57839 );
buf \U$57866 ( \57841 , \57830 );
not \U$57867 ( \57842 , \57841 );
buf \U$57868 ( \57843 , \57842 );
buf \U$57869 ( \57844 , \57843 );
buf \U$57870 ( \57845 , \57819 );
nand \U$57871 ( \57846 , \57844 , \57845 );
buf \U$57872 ( \57847 , \57846 );
buf \U$57873 ( \57848 , \57847 );
nand \U$57874 ( \57849 , \57840 , \57848 );
buf \U$57875 ( \57850 , \57849 );
buf \U$57876 ( \57851 , \57850 );
not \U$57877 ( \57852 , \57851 );
buf \U$57878 ( \57853 , \57852 );
buf \U$57879 ( \57854 , \57853 );
nand \U$57880 ( \57855 , \57480 , \57854 );
buf \U$57881 ( \57856 , \57855 );
buf \U$57882 ( \57857 , \57856 );
and \U$57883 ( \57858 , \57473 , \57857 );
buf \U$57884 ( \57859 , \57858 );
buf \U$57885 ( \57860 , \57859 );
buf \U$57886 ( \57861 , \52824 );
buf \U$57887 ( \57862 , \52413 );
xor \U$57888 ( \57863 , \57861 , \57862 );
buf \U$57889 ( \57864 , \57863 );
xor \U$57890 ( \57865 , \52611 , \57864 );
buf \U$57891 ( \57866 , \57865 );
xor \U$57892 ( \57867 , \52876 , \52880 );
xor \U$57893 ( \57868 , \57867 , \53218 );
buf \U$57894 ( \57869 , \57868 );
buf \U$57895 ( \57870 , \57869 );
xor \U$57896 ( \57871 , \57866 , \57870 );
buf \U$57897 ( \57872 , \57050 );
not \U$57898 ( \57873 , \57872 );
buf \U$57899 ( \57874 , \57057 );
nand \U$57900 ( \57875 , \57873 , \57874 );
buf \U$57901 ( \57876 , \57875 );
buf \U$57902 ( \57877 , \57876 );
not \U$57903 ( \57878 , \57877 );
buf \U$57904 ( \57879 , \57068 );
not \U$57905 ( \57880 , \57879 );
or \U$57906 ( \57881 , \57878 , \57880 );
buf \U$57907 ( \57882 , \57050 );
buf \U$57908 ( \57883 , \57054 );
nand \U$57909 ( \57884 , \57882 , \57883 );
buf \U$57910 ( \57885 , \57884 );
buf \U$57911 ( \57886 , \57885 );
nand \U$57912 ( \57887 , \57881 , \57886 );
buf \U$57913 ( \57888 , \57887 );
buf \U$57914 ( \57889 , \57888 );
xnor \U$57915 ( \57890 , \57871 , \57889 );
buf \U$57916 ( \57891 , \57890 );
buf \U$57917 ( \57892 , \57891 );
buf \U$57918 ( \57893 , \56932 );
not \U$57919 ( \57894 , \57893 );
buf \U$57920 ( \57895 , \57014 );
nand \U$57921 ( \57896 , \57894 , \57895 );
buf \U$57922 ( \57897 , \57896 );
buf \U$57923 ( \57898 , \57897 );
not \U$57924 ( \57899 , \57898 );
buf \U$57925 ( \57900 , \57071 );
not \U$57926 ( \57901 , \57900 );
buf \U$57927 ( \57902 , \57901 );
buf \U$57928 ( \57903 , \57902 );
not \U$57929 ( \57904 , \57903 );
or \U$57930 ( \57905 , \57899 , \57904 );
buf \U$57931 ( \57906 , \57011 );
buf \U$57932 ( \57907 , \56932 );
nand \U$57933 ( \57908 , \57906 , \57907 );
buf \U$57934 ( \57909 , \57908 );
buf \U$57935 ( \57910 , \57909 );
nand \U$57936 ( \57911 , \57905 , \57910 );
buf \U$57937 ( \57912 , \57911 );
buf \U$57938 ( \57913 , \57912 );
not \U$57939 ( \57914 , \57913 );
buf \U$57940 ( \57915 , \57914 );
buf \U$57941 ( \57916 , \57915 );
nand \U$57942 ( \57917 , \57892 , \57916 );
buf \U$57943 ( \57918 , \57917 );
buf \U$57944 ( \57919 , \57918 );
buf \U$57945 ( \57920 , \57869 );
buf \U$57946 ( \57921 , \57888 );
or \U$57947 ( \57922 , \57920 , \57921 );
buf \U$57948 ( \57923 , \57865 );
nand \U$57949 ( \57924 , \57922 , \57923 );
buf \U$57950 ( \57925 , \57924 );
buf \U$57951 ( \57926 , \57925 );
buf \U$57952 ( \57927 , \57869 );
buf \U$57953 ( \57928 , \57888 );
nand \U$57954 ( \57929 , \57927 , \57928 );
buf \U$57955 ( \57930 , \57929 );
buf \U$57956 ( \57931 , \57930 );
and \U$57957 ( \57932 , \57926 , \57931 );
buf \U$57958 ( \57933 , \57932 );
buf \U$57959 ( \57934 , \57933 );
buf \U$57960 ( \57935 , \53226 );
buf \U$57961 ( \57936 , \53222 );
xor \U$57962 ( \57937 , \57935 , \57936 );
buf \U$57963 ( \57938 , \53231 );
xnor \U$57964 ( \57939 , \57937 , \57938 );
buf \U$57965 ( \57940 , \57939 );
buf \U$57966 ( \57941 , \57940 );
nand \U$57967 ( \57942 , \57934 , \57941 );
buf \U$57968 ( \57943 , \57942 );
buf \U$57969 ( \57944 , \57943 );
nand \U$57970 ( \57945 , \57860 , \57919 , \57944 );
buf \U$57971 ( \57946 , \57945 );
buf \U$57972 ( \57947 , \57946 );
xor \U$57973 ( \57948 , \57775 , \57792 );
xor \U$57974 ( \57949 , \57948 , \57797 );
buf \U$57975 ( \57950 , \57949 );
buf \U$57976 ( \57951 , \57950 );
not \U$57977 ( \57952 , \57951 );
buf \U$57978 ( \57953 , RIc0d9040_56);
buf \U$57979 ( \57954 , RIc0daaf8_113);
xor \U$57980 ( \57955 , \57953 , \57954 );
buf \U$57981 ( \57956 , \57955 );
buf \U$57982 ( \57957 , \57956 );
not \U$57983 ( \57958 , \57957 );
buf \U$57984 ( \57959 , \26484 );
not \U$57985 ( \57960 , \57959 );
or \U$57986 ( \57961 , \57958 , \57960 );
buf \U$57987 ( \57962 , \16995 );
buf \U$57988 ( \57963 , \57254 );
nand \U$57989 ( \57964 , \57962 , \57963 );
buf \U$57990 ( \57965 , \57964 );
buf \U$57991 ( \57966 , \57965 );
nand \U$57992 ( \57967 , \57961 , \57966 );
buf \U$57993 ( \57968 , \57967 );
buf \U$57994 ( \57969 , \57968 );
buf \U$57995 ( \57970 , \45548 );
buf \U$57996 ( \57971 , RIc0daeb8_121);
buf \U$57997 ( \57972 , RIc0d8c80_48);
xnor \U$57998 ( \57973 , \57971 , \57972 );
buf \U$57999 ( \57974 , \57973 );
buf \U$58000 ( \57975 , \57974 );
or \U$58001 ( \57976 , \57970 , \57975 );
buf \U$58002 ( \57977 , \26373 );
buf \U$58003 ( \57978 , \57485 );
or \U$58004 ( \57979 , \57977 , \57978 );
nand \U$58005 ( \57980 , \57976 , \57979 );
buf \U$58006 ( \57981 , \57980 );
buf \U$58007 ( \57982 , \57981 );
xor \U$58008 ( \57983 , \57969 , \57982 );
buf \U$58009 ( \57984 , \57529 );
not \U$58010 ( \57985 , \57984 );
buf \U$58011 ( \57986 , \57512 );
not \U$58012 ( \57987 , \57986 );
or \U$58013 ( \57988 , \57985 , \57987 );
buf \U$58014 ( \57989 , \57512 );
buf \U$58015 ( \57990 , \57529 );
or \U$58016 ( \57991 , \57989 , \57990 );
nand \U$58017 ( \57992 , \57988 , \57991 );
buf \U$58018 ( \57993 , \57992 );
buf \U$58019 ( \57994 , \57993 );
and \U$58020 ( \57995 , \57983 , \57994 );
and \U$58021 ( \57996 , \57969 , \57982 );
or \U$58022 ( \57997 , \57995 , \57996 );
buf \U$58023 ( \57998 , \57997 );
buf \U$58024 ( \57999 , \57998 );
xor \U$58025 ( \58000 , \57496 , \57533 );
xor \U$58026 ( \58001 , \58000 , \57600 );
buf \U$58027 ( \58002 , \58001 );
buf \U$58028 ( \58003 , \58002 );
xor \U$58029 ( \58004 , \57999 , \58003 );
buf \U$58030 ( \58005 , RIc0d90b8_57);
buf \U$58031 ( \58006 , RIc0daaf8_113);
xor \U$58032 ( \58007 , \58005 , \58006 );
buf \U$58033 ( \58008 , \58007 );
buf \U$58034 ( \58009 , \58008 );
not \U$58035 ( \58010 , \58009 );
buf \U$58036 ( \58011 , \16656 );
not \U$58037 ( \58012 , \58011 );
or \U$58038 ( \58013 , \58010 , \58012 );
buf \U$58039 ( \58014 , \14405 );
buf \U$58040 ( \58015 , \57956 );
nand \U$58041 ( \58016 , \58014 , \58015 );
buf \U$58042 ( \58017 , \58016 );
buf \U$58043 ( \58018 , \58017 );
nand \U$58044 ( \58019 , \58013 , \58018 );
buf \U$58045 ( \58020 , \58019 );
buf \U$58046 ( \58021 , \58020 );
not \U$58047 ( \58022 , \58021 );
buf \U$58048 ( \58023 , \58022 );
buf \U$58049 ( \58024 , \58023 );
not \U$58050 ( \58025 , \58024 );
buf \U$58051 ( \58026 , RIc0d9388_63);
buf \U$58052 ( \58027 , RIc0da828_107);
xor \U$58053 ( \58028 , \58026 , \58027 );
buf \U$58054 ( \58029 , \58028 );
buf \U$58055 ( \58030 , \58029 );
not \U$58056 ( \58031 , \58030 );
buf \U$58057 ( \58032 , \34202 );
not \U$58058 ( \58033 , \58032 );
or \U$58059 ( \58034 , \58031 , \58033 );
buf \U$58060 ( \58035 , \12342 );
buf \U$58061 ( \58036 , \57500 );
nand \U$58062 ( \58037 , \58035 , \58036 );
buf \U$58063 ( \58038 , \58037 );
buf \U$58064 ( \58039 , \58038 );
nand \U$58065 ( \58040 , \58034 , \58039 );
buf \U$58066 ( \58041 , \58040 );
buf \U$58067 ( \58042 , \58041 );
not \U$58068 ( \58043 , \58042 );
buf \U$58069 ( \58044 , \58043 );
buf \U$58070 ( \58045 , \58044 );
not \U$58071 ( \58046 , \58045 );
or \U$58072 ( \58047 , \58025 , \58046 );
buf \U$58073 ( \58048 , RIc0d91a8_59);
buf \U$58074 ( \58049 , RIc0daa08_111);
xor \U$58075 ( \58050 , \58048 , \58049 );
buf \U$58076 ( \58051 , \58050 );
buf \U$58077 ( \58052 , \58051 );
not \U$58078 ( \58053 , \58052 );
buf \U$58079 ( \58054 , \12529 );
not \U$58080 ( \58055 , \58054 );
or \U$58081 ( \58056 , \58053 , \58055 );
buf \U$58082 ( \58057 , \57705 );
not \U$58083 ( \58058 , \58057 );
buf \U$58084 ( \58059 , \14352 );
nand \U$58085 ( \58060 , \58058 , \58059 );
buf \U$58086 ( \58061 , \58060 );
buf \U$58087 ( \58062 , \58061 );
nand \U$58088 ( \58063 , \58056 , \58062 );
buf \U$58089 ( \58064 , \58063 );
buf \U$58090 ( \58065 , \58064 );
nand \U$58091 ( \58066 , \58047 , \58065 );
buf \U$58092 ( \58067 , \58066 );
buf \U$58093 ( \58068 , \58067 );
buf \U$58094 ( \58069 , \58041 );
buf \U$58095 ( \58070 , \58020 );
nand \U$58096 ( \58071 , \58069 , \58070 );
buf \U$58097 ( \58072 , \58071 );
buf \U$58098 ( \58073 , \58072 );
nand \U$58099 ( \58074 , \58068 , \58073 );
buf \U$58100 ( \58075 , \58074 );
buf \U$58101 ( \58076 , \58075 );
buf \U$58102 ( \58077 , \21880 );
buf \U$58103 ( \58078 , RIc0d9400_64);
and \U$58104 ( \58079 , \58077 , \58078 );
buf \U$58105 ( \58080 , \58079 );
buf \U$58106 ( \58081 , \58080 );
buf \U$58107 ( \58082 , RIc0da918_109);
buf \U$58108 ( \58083 , RIc0d9298_61);
xor \U$58109 ( \58084 , \58082 , \58083 );
buf \U$58110 ( \58085 , \58084 );
buf \U$58111 ( \58086 , \58085 );
not \U$58112 ( \58087 , \58086 );
buf \U$58113 ( \58088 , \14210 );
not \U$58114 ( \58089 , \58088 );
or \U$58115 ( \58090 , \58087 , \58089 );
buf \U$58116 ( \58091 , \16232 );
buf \U$58117 ( \58092 , \57556 );
nand \U$58118 ( \58093 , \58091 , \58092 );
buf \U$58119 ( \58094 , \58093 );
buf \U$58120 ( \58095 , \58094 );
nand \U$58121 ( \58096 , \58090 , \58095 );
buf \U$58122 ( \58097 , \58096 );
buf \U$58123 ( \58098 , \58097 );
xor \U$58124 ( \58099 , \58081 , \58098 );
buf \U$58125 ( \58100 , \46459 );
buf \U$58126 ( \58101 , RIc0d8b18_45);
buf \U$58127 ( \58102 , RIc0db098_125);
xnor \U$58128 ( \58103 , \58101 , \58102 );
buf \U$58129 ( \58104 , \58103 );
buf \U$58130 ( \58105 , \58104 );
or \U$58131 ( \58106 , \58100 , \58105 );
buf \U$58132 ( \58107 , \22744 );
buf \U$58133 ( \58108 , \57691 );
or \U$58134 ( \58109 , \58107 , \58108 );
nand \U$58135 ( \58110 , \58106 , \58109 );
buf \U$58136 ( \58111 , \58110 );
buf \U$58137 ( \58112 , \58111 );
and \U$58138 ( \58113 , \58099 , \58112 );
and \U$58139 ( \58114 , \58081 , \58098 );
or \U$58140 ( \58115 , \58113 , \58114 );
buf \U$58141 ( \58116 , \58115 );
buf \U$58142 ( \58117 , \58116 );
xor \U$58143 ( \58118 , \58076 , \58117 );
buf \U$58144 ( \58119 , RIc0d8cf8_49);
buf \U$58145 ( \58120 , RIc0daeb8_121);
xor \U$58146 ( \58121 , \58119 , \58120 );
buf \U$58147 ( \58122 , \58121 );
buf \U$58148 ( \58123 , \58122 );
not \U$58149 ( \58124 , \58123 );
buf \U$58150 ( \58125 , \19487 );
not \U$58151 ( \58126 , \58125 );
or \U$58152 ( \58127 , \58124 , \58126 );
buf \U$58153 ( \58128 , \57974 );
not \U$58154 ( \58129 , \58128 );
buf \U$58155 ( \58130 , \16386 );
nand \U$58156 ( \58131 , \58129 , \58130 );
buf \U$58157 ( \58132 , \58131 );
buf \U$58158 ( \58133 , \58132 );
nand \U$58159 ( \58134 , \58127 , \58133 );
buf \U$58160 ( \58135 , \58134 );
buf \U$58161 ( \58136 , \58135 );
buf \U$58162 ( \58137 , RIc0dabe8_115);
buf \U$58163 ( \58138 , RIc0d8fc8_55);
xor \U$58164 ( \58139 , \58137 , \58138 );
buf \U$58165 ( \58140 , \58139 );
buf \U$58166 ( \58141 , \58140 );
not \U$58167 ( \58142 , \58141 );
buf \U$58168 ( \58143 , \26466 );
not \U$58169 ( \58144 , \58143 );
or \U$58170 ( \58145 , \58142 , \58144 );
buf \U$58171 ( \58146 , \57618 );
not \U$58172 ( \58147 , \58146 );
buf \U$58173 ( \58148 , \12303 );
nand \U$58174 ( \58149 , \58147 , \58148 );
buf \U$58175 ( \58150 , \58149 );
buf \U$58176 ( \58151 , \58150 );
nand \U$58177 ( \58152 , \58145 , \58151 );
buf \U$58178 ( \58153 , \58152 );
buf \U$58179 ( \58154 , \58153 );
xor \U$58180 ( \58155 , \58136 , \58154 );
buf \U$58181 ( \58156 , \16688 );
buf \U$58182 ( \58157 , RIc0d8c08_47);
buf \U$58183 ( \58158 , RIc0dafa8_123);
xor \U$58184 ( \58159 , \58157 , \58158 );
buf \U$58185 ( \58160 , \58159 );
buf \U$58186 ( \58161 , \58160 );
not \U$58187 ( \58162 , \58161 );
buf \U$58188 ( \58163 , \58162 );
buf \U$58189 ( \58164 , \58163 );
or \U$58190 ( \58165 , \58156 , \58164 );
buf \U$58191 ( \58166 , \16695 );
buf \U$58192 ( \58167 , \57578 );
or \U$58193 ( \58168 , \58166 , \58167 );
nand \U$58194 ( \58169 , \58165 , \58168 );
buf \U$58195 ( \58170 , \58169 );
buf \U$58196 ( \58171 , \58170 );
and \U$58197 ( \58172 , \58155 , \58171 );
and \U$58198 ( \58173 , \58136 , \58154 );
or \U$58199 ( \58174 , \58172 , \58173 );
buf \U$58200 ( \58175 , \58174 );
buf \U$58201 ( \58176 , \58175 );
and \U$58202 ( \58177 , \58118 , \58176 );
and \U$58203 ( \58178 , \58076 , \58117 );
or \U$58204 ( \58179 , \58177 , \58178 );
buf \U$58205 ( \58180 , \58179 );
buf \U$58206 ( \58181 , \58180 );
and \U$58207 ( \58182 , \58004 , \58181 );
and \U$58208 ( \58183 , \57999 , \58003 );
or \U$58209 ( \58184 , \58182 , \58183 );
buf \U$58210 ( \58185 , \58184 );
buf \U$58211 ( \58186 , \58185 );
buf \U$58212 ( \58187 , \57550 );
buf \U$58213 ( \58188 , \57568 );
xor \U$58214 ( \58189 , \58187 , \58188 );
buf \U$58215 ( \58190 , \57593 );
xnor \U$58216 ( \58191 , \58189 , \58190 );
buf \U$58217 ( \58192 , \58191 );
buf \U$58218 ( \58193 , \58192 );
not \U$58219 ( \58194 , \58193 );
xor \U$58220 ( \58195 , \57668 , \57649 );
xnor \U$58221 ( \58196 , \58195 , \57628 );
buf \U$58222 ( \58197 , \58196 );
not \U$58223 ( \58198 , \58197 );
or \U$58224 ( \58199 , \58194 , \58198 );
not \U$58225 ( \58200 , \43781 );
buf \U$58226 ( \58201 , \58200 );
xor \U$58227 ( \58202 , RIc0db188_127, RIc0d8a28_43);
buf \U$58228 ( \58203 , \58202 );
not \U$58229 ( \58204 , \58203 );
buf \U$58230 ( \58205 , \58204 );
buf \U$58231 ( \58206 , \58205 );
or \U$58232 ( \58207 , \58201 , \58206 );
buf \U$58233 ( \58208 , \12647 );
buf \U$58234 ( \58209 , \57538 );
not \U$58235 ( \58210 , \58209 );
buf \U$58236 ( \58211 , \58210 );
buf \U$58237 ( \58212 , \58211 );
or \U$58238 ( \58213 , \58208 , \58212 );
nand \U$58239 ( \58214 , \58207 , \58213 );
buf \U$58240 ( \58215 , \58214 );
buf \U$58241 ( \58216 , \58215 );
buf \U$58242 ( \58217 , RIc0d8de8_51);
buf \U$58243 ( \58218 , RIc0dadc8_119);
xor \U$58244 ( \58219 , \58217 , \58218 );
buf \U$58245 ( \58220 , \58219 );
buf \U$58246 ( \58221 , \58220 );
not \U$58247 ( \58222 , \58221 );
buf \U$58248 ( \58223 , \14569 );
not \U$58249 ( \58224 , \58223 );
or \U$58250 ( \58225 , \58222 , \58224 );
buf \U$58251 ( \58226 , \13953 );
buf \U$58252 ( \58227 , \57656 );
nand \U$58253 ( \58228 , \58226 , \58227 );
buf \U$58254 ( \58229 , \58228 );
buf \U$58255 ( \58230 , \58229 );
nand \U$58256 ( \58231 , \58225 , \58230 );
buf \U$58257 ( \58232 , \58231 );
buf \U$58258 ( \58233 , \58232 );
xor \U$58259 ( \58234 , \58216 , \58233 );
buf \U$58260 ( \58235 , \12926 );
buf \U$58261 ( \58236 , RIc0d8ed8_53);
buf \U$58262 ( \58237 , RIc0dacd8_117);
xnor \U$58263 ( \58238 , \58236 , \58237 );
buf \U$58264 ( \58239 , \58238 );
buf \U$58265 ( \58240 , \58239 );
or \U$58266 ( \58241 , \58235 , \58240 );
buf \U$58267 ( \58242 , \44894 );
buf \U$58268 ( \58243 , \57634 );
not \U$58269 ( \58244 , \58243 );
buf \U$58270 ( \58245 , \58244 );
buf \U$58271 ( \58246 , \58245 );
or \U$58272 ( \58247 , \58242 , \58246 );
nand \U$58273 ( \58248 , \58241 , \58247 );
buf \U$58274 ( \58249 , \58248 );
buf \U$58275 ( \58250 , \58249 );
and \U$58276 ( \58251 , \58234 , \58250 );
and \U$58277 ( \58252 , \58216 , \58233 );
or \U$58278 ( \58253 , \58251 , \58252 );
buf \U$58279 ( \58254 , \58253 );
buf \U$58280 ( \58255 , \58254 );
nand \U$58281 ( \58256 , \58199 , \58255 );
buf \U$58282 ( \58257 , \58256 );
buf \U$58283 ( \58258 , \58257 );
buf \U$58284 ( \58259 , \58192 );
not \U$58285 ( \58260 , \58259 );
buf \U$58286 ( \58261 , \58196 );
not \U$58287 ( \58262 , \58261 );
buf \U$58288 ( \58263 , \58262 );
buf \U$58289 ( \58264 , \58263 );
nand \U$58290 ( \58265 , \58260 , \58264 );
buf \U$58291 ( \58266 , \58265 );
buf \U$58292 ( \58267 , \58266 );
nand \U$58293 ( \58268 , \58258 , \58267 );
buf \U$58294 ( \58269 , \58268 );
buf \U$58295 ( \58270 , \58269 );
not \U$58296 ( \58271 , \58270 );
buf \U$58297 ( \58272 , \57610 );
not \U$58298 ( \58273 , \58272 );
buf \U$58299 ( \58274 , \57680 );
not \U$58300 ( \58275 , \58274 );
buf \U$58301 ( \58276 , \57745 );
not \U$58302 ( \58277 , \58276 );
or \U$58303 ( \58278 , \58275 , \58277 );
buf \U$58304 ( \58279 , \57745 );
buf \U$58305 ( \58280 , \57680 );
or \U$58306 ( \58281 , \58279 , \58280 );
nand \U$58307 ( \58282 , \58278 , \58281 );
buf \U$58308 ( \58283 , \58282 );
buf \U$58309 ( \58284 , \58283 );
not \U$58310 ( \58285 , \58284 );
or \U$58311 ( \58286 , \58273 , \58285 );
buf \U$58312 ( \58287 , \58283 );
buf \U$58313 ( \58288 , \57610 );
or \U$58314 ( \58289 , \58287 , \58288 );
nand \U$58315 ( \58290 , \58286 , \58289 );
buf \U$58316 ( \58291 , \58290 );
buf \U$58317 ( \58292 , \58291 );
not \U$58318 ( \58293 , \58292 );
or \U$58319 ( \58294 , \58271 , \58293 );
buf \U$58320 ( \58295 , \58291 );
buf \U$58321 ( \58296 , \58269 );
or \U$58322 ( \58297 , \58295 , \58296 );
xor \U$58323 ( \58298 , \57779 , \57783 );
xor \U$58324 ( \58299 , \58298 , \57787 );
buf \U$58325 ( \58300 , \58299 );
buf \U$58326 ( \58301 , \58300 );
nand \U$58327 ( \58302 , \58297 , \58301 );
buf \U$58328 ( \58303 , \58302 );
buf \U$58329 ( \58304 , \58303 );
nand \U$58330 ( \58305 , \58294 , \58304 );
buf \U$58331 ( \58306 , \58305 );
buf \U$58332 ( \58307 , \58306 );
xor \U$58333 ( \58308 , \58186 , \58307 );
xor \U$58334 ( \58309 , \57605 , \57761 );
xor \U$58335 ( \58310 , \58309 , \57766 );
buf \U$58336 ( \58311 , \58310 );
buf \U$58337 ( \58312 , \58311 );
xnor \U$58338 ( \58313 , \58308 , \58312 );
buf \U$58339 ( \58314 , \58313 );
buf \U$58340 ( \58315 , \58314 );
not \U$58341 ( \58316 , \58315 );
buf \U$58342 ( \58317 , \58316 );
buf \U$58343 ( \58318 , \58317 );
not \U$58344 ( \58319 , \58318 );
or \U$58345 ( \58320 , \57952 , \58319 );
buf \U$58346 ( \58321 , \57950 );
not \U$58347 ( \58322 , \58321 );
buf \U$58348 ( \58323 , \58322 );
buf \U$58349 ( \58324 , \58323 );
not \U$58350 ( \58325 , \58324 );
buf \U$58351 ( \58326 , \58314 );
not \U$58352 ( \58327 , \58326 );
or \U$58353 ( \58328 , \58325 , \58327 );
and \U$58354 ( \58329 , \57728 , \57709 );
not \U$58355 ( \58330 , \57728 );
and \U$58356 ( \58331 , \58330 , \57735 );
or \U$58357 ( \58332 , \58329 , \58331 );
buf \U$58358 ( \58333 , \58332 );
buf \U$58359 ( \58334 , \57739 );
and \U$58360 ( \58335 , \58333 , \58334 );
not \U$58361 ( \58336 , \58333 );
buf \U$58362 ( \58337 , \57698 );
and \U$58363 ( \58338 , \58336 , \58337 );
nor \U$58364 ( \58339 , \58335 , \58338 );
buf \U$58365 ( \58340 , \58339 );
buf \U$58366 ( \58341 , \58340 );
xor \U$58367 ( \58342 , \57969 , \57982 );
xor \U$58368 ( \58343 , \58342 , \57994 );
buf \U$58369 ( \58344 , \58343 );
buf \U$58370 ( \58345 , \58344 );
xor \U$58371 ( \58346 , \58341 , \58345 );
buf \U$58372 ( \58347 , RIc0d9400_64);
buf \U$58373 ( \58348 , RIc0da8a0_108);
or \U$58374 ( \58349 , \58347 , \58348 );
buf \U$58375 ( \58350 , RIc0da918_109);
nand \U$58376 ( \58351 , \58349 , \58350 );
buf \U$58377 ( \58352 , \58351 );
buf \U$58378 ( \58353 , \58352 );
buf \U$58379 ( \58354 , RIc0d9400_64);
buf \U$58380 ( \58355 , RIc0da8a0_108);
nand \U$58381 ( \58356 , \58354 , \58355 );
buf \U$58382 ( \58357 , \58356 );
buf \U$58383 ( \58358 , \58357 );
buf \U$58384 ( \58359 , RIc0da828_107);
and \U$58385 ( \58360 , \58353 , \58358 , \58359 );
buf \U$58386 ( \58361 , \58360 );
buf \U$58387 ( \58362 , \58361 );
buf \U$58388 ( \58363 , RIc0da918_109);
buf \U$58389 ( \58364 , RIc0d9310_62);
xor \U$58390 ( \58365 , \58363 , \58364 );
buf \U$58391 ( \58366 , \58365 );
buf \U$58392 ( \58367 , \58366 );
not \U$58393 ( \58368 , \58367 );
buf \U$58394 ( \58369 , \20759 );
not \U$58395 ( \58370 , \58369 );
or \U$58396 ( \58371 , \58368 , \58370 );
buf \U$58397 ( \58372 , \20211 );
buf \U$58398 ( \58373 , \58085 );
nand \U$58399 ( \58374 , \58372 , \58373 );
buf \U$58400 ( \58375 , \58374 );
buf \U$58401 ( \58376 , \58375 );
nand \U$58402 ( \58377 , \58371 , \58376 );
buf \U$58403 ( \58378 , \58377 );
buf \U$58404 ( \58379 , \58378 );
and \U$58405 ( \58380 , \58362 , \58379 );
buf \U$58406 ( \58381 , \58380 );
buf \U$58407 ( \58382 , \58381 );
buf \U$58408 ( \58383 , RIc0daeb8_121);
buf \U$58409 ( \58384 , RIc0d8d70_50);
xor \U$58410 ( \58385 , \58383 , \58384 );
buf \U$58411 ( \58386 , \58385 );
buf \U$58412 ( \58387 , \58386 );
not \U$58413 ( \58388 , \58387 );
buf \U$58414 ( \58389 , \17089 );
not \U$58415 ( \58390 , \58389 );
or \U$58416 ( \58391 , \58388 , \58390 );
buf \U$58417 ( \58392 , \13314 );
buf \U$58418 ( \58393 , \58122 );
nand \U$58419 ( \58394 , \58392 , \58393 );
buf \U$58420 ( \58395 , \58394 );
buf \U$58421 ( \58396 , \58395 );
nand \U$58422 ( \58397 , \58391 , \58396 );
buf \U$58423 ( \58398 , \58397 );
buf \U$58424 ( \58399 , \58398 );
buf \U$58425 ( \58400 , RIc0dacd8_117);
buf \U$58426 ( \58401 , RIc0d8f50_54);
xor \U$58427 ( \58402 , \58400 , \58401 );
buf \U$58428 ( \58403 , \58402 );
buf \U$58429 ( \58404 , \58403 );
not \U$58430 ( \58405 , \58404 );
buf \U$58431 ( \58406 , \22350 );
not \U$58432 ( \58407 , \58406 );
or \U$58433 ( \58408 , \58405 , \58407 );
buf \U$58434 ( \58409 , \58239 );
not \U$58435 ( \58410 , \58409 );
buf \U$58436 ( \58411 , \12937 );
nand \U$58437 ( \58412 , \58410 , \58411 );
buf \U$58438 ( \58413 , \58412 );
buf \U$58439 ( \58414 , \58413 );
nand \U$58440 ( \58415 , \58408 , \58414 );
buf \U$58441 ( \58416 , \58415 );
buf \U$58442 ( \58417 , \58416 );
xor \U$58443 ( \58418 , \58399 , \58417 );
xnor \U$58444 ( \58419 , RIc0dabe8_115, RIc0d9040_56);
buf \U$58445 ( \58420 , \58419 );
not \U$58446 ( \58421 , \58420 );
buf \U$58447 ( \58422 , \58421 );
buf \U$58448 ( \58423 , \58422 );
not \U$58449 ( \58424 , \58423 );
buf \U$58450 ( \58425 , \46873 );
not \U$58451 ( \58426 , \58425 );
or \U$58452 ( \58427 , \58424 , \58426 );
buf \U$58453 ( \58428 , \12303 );
buf \U$58454 ( \58429 , \58140 );
nand \U$58455 ( \58430 , \58428 , \58429 );
buf \U$58456 ( \58431 , \58430 );
buf \U$58457 ( \58432 , \58431 );
nand \U$58458 ( \58433 , \58427 , \58432 );
buf \U$58459 ( \58434 , \58433 );
buf \U$58460 ( \58435 , \58434 );
and \U$58461 ( \58436 , \58418 , \58435 );
and \U$58462 ( \58437 , \58399 , \58417 );
or \U$58463 ( \58438 , \58436 , \58437 );
buf \U$58464 ( \58439 , \58438 );
buf \U$58465 ( \58440 , \58439 );
xor \U$58466 ( \58441 , \58382 , \58440 );
buf \U$58467 ( \58442 , RIc0daaf8_113);
buf \U$58468 ( \58443 , RIc0d9130_58);
xor \U$58469 ( \58444 , \58442 , \58443 );
buf \U$58470 ( \58445 , \58444 );
buf \U$58471 ( \58446 , \58445 );
not \U$58472 ( \58447 , \58446 );
buf \U$58473 ( \58448 , \28413 );
not \U$58474 ( \58449 , \58448 );
or \U$58475 ( \58450 , \58447 , \58449 );
buf \U$58476 ( \58451 , \16662 );
buf \U$58477 ( \58452 , \58008 );
nand \U$58478 ( \58453 , \58451 , \58452 );
buf \U$58479 ( \58454 , \58453 );
buf \U$58480 ( \58455 , \58454 );
nand \U$58481 ( \58456 , \58450 , \58455 );
buf \U$58482 ( \58457 , \58456 );
buf \U$58483 ( \58458 , \58457 );
not \U$58484 ( \58459 , \58458 );
buf \U$58485 ( \58460 , \54203 );
buf \U$58486 ( \58461 , RIc0db098_125);
buf \U$58487 ( \58462 , RIc0d8b90_46);
xnor \U$58488 ( \58463 , \58461 , \58462 );
buf \U$58489 ( \58464 , \58463 );
buf \U$58490 ( \58465 , \58464 );
or \U$58491 ( \58466 , \58460 , \58465 );
buf \U$58492 ( \58467 , \22744 );
buf \U$58493 ( \58468 , \58104 );
or \U$58494 ( \58469 , \58467 , \58468 );
nand \U$58495 ( \58470 , \58466 , \58469 );
buf \U$58496 ( \58471 , \58470 );
buf \U$58497 ( \58472 , \58471 );
not \U$58498 ( \58473 , \58472 );
or \U$58499 ( \58474 , \58459 , \58473 );
buf \U$58500 ( \58475 , \58471 );
buf \U$58501 ( \58476 , \58457 );
or \U$58502 ( \58477 , \58475 , \58476 );
buf \U$58503 ( \58478 , RIc0da828_107);
buf \U$58504 ( \58479 , RIc0d9400_64);
and \U$58505 ( \58480 , \58478 , \58479 );
not \U$58506 ( \58481 , \58478 );
buf \U$58507 ( \58482 , \43843 );
and \U$58508 ( \58483 , \58481 , \58482 );
nor \U$58509 ( \58484 , \58480 , \58483 );
buf \U$58510 ( \58485 , \58484 );
buf \U$58511 ( \58486 , \58485 );
not \U$58512 ( \58487 , \58486 );
buf \U$58513 ( \58488 , \37534 );
not \U$58514 ( \58489 , \58488 );
or \U$58515 ( \58490 , \58487 , \58489 );
buf \U$58516 ( \58491 , \12342 );
buf \U$58517 ( \58492 , \58029 );
nand \U$58518 ( \58493 , \58491 , \58492 );
buf \U$58519 ( \58494 , \58493 );
buf \U$58520 ( \58495 , \58494 );
nand \U$58521 ( \58496 , \58490 , \58495 );
buf \U$58522 ( \58497 , \58496 );
buf \U$58523 ( \58498 , \58497 );
nand \U$58524 ( \58499 , \58477 , \58498 );
buf \U$58525 ( \58500 , \58499 );
buf \U$58526 ( \58501 , \58500 );
nand \U$58527 ( \58502 , \58474 , \58501 );
buf \U$58528 ( \58503 , \58502 );
buf \U$58529 ( \58504 , \58503 );
and \U$58530 ( \58505 , \58441 , \58504 );
and \U$58531 ( \58506 , \58382 , \58440 );
or \U$58532 ( \58507 , \58505 , \58506 );
buf \U$58533 ( \58508 , \58507 );
buf \U$58534 ( \58509 , \58508 );
and \U$58535 ( \58510 , \58346 , \58509 );
and \U$58536 ( \58511 , \58341 , \58345 );
or \U$58537 ( \58512 , \58510 , \58511 );
buf \U$58538 ( \58513 , \58512 );
buf \U$58539 ( \58514 , \58513 );
buf \U$58540 ( \58515 , RIc0d8aa0_44);
buf \U$58541 ( \58516 , RIc0db188_127);
xor \U$58542 ( \58517 , \58515 , \58516 );
buf \U$58543 ( \58518 , \58517 );
buf \U$58544 ( \58519 , \58518 );
not \U$58545 ( \58520 , \58519 );
buf \U$58546 ( \58521 , \15609 );
buf \U$58547 ( \58522 , \58521 );
buf \U$58548 ( \58523 , \58522 );
not \U$58549 ( \58524 , \58523 );
or \U$58550 ( \58525 , \58520 , \58524 );
buf \U$58551 ( \58526 , \58202 );
buf \U$58552 ( \58527 , RIc0db200_128);
nand \U$58553 ( \58528 , \58526 , \58527 );
buf \U$58554 ( \58529 , \58528 );
buf \U$58555 ( \58530 , \58529 );
nand \U$58556 ( \58531 , \58525 , \58530 );
buf \U$58557 ( \58532 , \58531 );
buf \U$58558 ( \58533 , \58532 );
buf \U$58559 ( \58534 , RIc0d8e60_52);
buf \U$58560 ( \58535 , RIc0dadc8_119);
xor \U$58561 ( \58536 , \58534 , \58535 );
buf \U$58562 ( \58537 , \58536 );
buf \U$58563 ( \58538 , \58537 );
not \U$58564 ( \58539 , \58538 );
buf \U$58565 ( \58540 , \23985 );
not \U$58566 ( \58541 , \58540 );
or \U$58567 ( \58542 , \58539 , \58541 );
buf \U$58568 ( \58543 , \13953 );
buf \U$58569 ( \58544 , \58220 );
nand \U$58570 ( \58545 , \58543 , \58544 );
buf \U$58571 ( \58546 , \58545 );
buf \U$58572 ( \58547 , \58546 );
nand \U$58573 ( \58548 , \58542 , \58547 );
buf \U$58574 ( \58549 , \58548 );
buf \U$58575 ( \58550 , \58549 );
xor \U$58576 ( \58551 , \58533 , \58550 );
buf \U$58577 ( \58552 , \37704 );
buf \U$58578 ( \58553 , RIc0daa08_111);
buf \U$58579 ( \58554 , RIc0d9220_60);
xnor \U$58580 ( \58555 , \58553 , \58554 );
buf \U$58581 ( \58556 , \58555 );
buf \U$58582 ( \58557 , \58556 );
or \U$58583 ( \58558 , \58552 , \58557 );
buf \U$58584 ( \58559 , \45725 );
buf \U$58585 ( \58560 , \58051 );
not \U$58586 ( \58561 , \58560 );
buf \U$58587 ( \58562 , \58561 );
buf \U$58588 ( \58563 , \58562 );
or \U$58589 ( \58564 , \58559 , \58563 );
nand \U$58590 ( \58565 , \58558 , \58564 );
buf \U$58591 ( \58566 , \58565 );
buf \U$58592 ( \58567 , \58566 );
and \U$58593 ( \58568 , \58551 , \58567 );
and \U$58594 ( \58569 , \58533 , \58550 );
or \U$58595 ( \58570 , \58568 , \58569 );
buf \U$58596 ( \58571 , \58570 );
buf \U$58597 ( \58572 , \58571 );
not \U$58598 ( \58573 , \58572 );
buf \U$58599 ( \58574 , \58573 );
buf \U$58600 ( \58575 , \58574 );
not \U$58601 ( \58576 , \58575 );
xor \U$58602 ( \58577 , \58064 , \58044 );
xnor \U$58603 ( \58578 , \58577 , \58023 );
buf \U$58604 ( \58579 , \58578 );
not \U$58605 ( \58580 , \58579 );
or \U$58606 ( \58581 , \58576 , \58580 );
xor \U$58607 ( \58582 , \58136 , \58154 );
xor \U$58608 ( \58583 , \58582 , \58171 );
buf \U$58609 ( \58584 , \58583 );
buf \U$58610 ( \58585 , \58584 );
nand \U$58611 ( \58586 , \58581 , \58585 );
buf \U$58612 ( \58587 , \58586 );
buf \U$58613 ( \58588 , \58587 );
buf \U$58614 ( \58589 , \58578 );
not \U$58615 ( \58590 , \58589 );
buf \U$58616 ( \58591 , \58571 );
nand \U$58617 ( \58592 , \58590 , \58591 );
buf \U$58618 ( \58593 , \58592 );
buf \U$58619 ( \58594 , \58593 );
nand \U$58620 ( \58595 , \58588 , \58594 );
buf \U$58621 ( \58596 , \58595 );
buf \U$58622 ( \58597 , \58596 );
xor \U$58623 ( \58598 , \58076 , \58117 );
xor \U$58624 ( \58599 , \58598 , \58176 );
buf \U$58625 ( \58600 , \58599 );
buf \U$58626 ( \58601 , \58600 );
xor \U$58627 ( \58602 , \58597 , \58601 );
buf \U$58628 ( \58603 , \58254 );
not \U$58629 ( \58604 , \58603 );
buf \U$58630 ( \58605 , \58192 );
not \U$58631 ( \58606 , \58605 );
or \U$58632 ( \58607 , \58604 , \58606 );
buf \U$58633 ( \58608 , \58254 );
buf \U$58634 ( \58609 , \58192 );
or \U$58635 ( \58610 , \58608 , \58609 );
nand \U$58636 ( \58611 , \58607 , \58610 );
buf \U$58637 ( \58612 , \58611 );
buf \U$58638 ( \58613 , \58612 );
buf \U$58639 ( \58614 , \58263 );
and \U$58640 ( \58615 , \58613 , \58614 );
not \U$58641 ( \58616 , \58613 );
buf \U$58642 ( \58617 , \58196 );
and \U$58643 ( \58618 , \58616 , \58617 );
nor \U$58644 ( \58619 , \58615 , \58618 );
buf \U$58645 ( \58620 , \58619 );
buf \U$58646 ( \58621 , \58620 );
and \U$58647 ( \58622 , \58602 , \58621 );
and \U$58648 ( \58623 , \58597 , \58601 );
or \U$58649 ( \58624 , \58622 , \58623 );
buf \U$58650 ( \58625 , \58624 );
buf \U$58651 ( \58626 , \58625 );
xor \U$58652 ( \58627 , \58514 , \58626 );
xor \U$58653 ( \58628 , \57999 , \58003 );
xor \U$58654 ( \58629 , \58628 , \58181 );
buf \U$58655 ( \58630 , \58629 );
buf \U$58656 ( \58631 , \58630 );
and \U$58657 ( \58632 , \58627 , \58631 );
and \U$58658 ( \58633 , \58514 , \58626 );
or \U$58659 ( \58634 , \58632 , \58633 );
buf \U$58660 ( \58635 , \58634 );
buf \U$58661 ( \58636 , \58635 );
nand \U$58662 ( \58637 , \58328 , \58636 );
buf \U$58663 ( \58638 , \58637 );
buf \U$58664 ( \58639 , \58638 );
nand \U$58665 ( \58640 , \58320 , \58639 );
buf \U$58666 ( \58641 , \58640 );
buf \U$58667 ( \58642 , \58641 );
not \U$58668 ( \58643 , \58642 );
xor \U$58669 ( \58644 , \57410 , \57439 );
xor \U$58670 ( \58645 , \58644 , \57430 );
buf \U$58671 ( \58646 , \58645 );
not \U$58672 ( \58647 , \58646 );
buf \U$58673 ( \58648 , \58647 );
buf \U$58674 ( \58649 , \58648 );
not \U$58675 ( \58650 , \58649 );
buf \U$58676 ( \58651 , \58306 );
not \U$58677 ( \58652 , \58651 );
buf \U$58678 ( \58653 , \58311 );
not \U$58679 ( \58654 , \58653 );
or \U$58680 ( \58655 , \58652 , \58654 );
buf \U$58681 ( \58656 , \58306 );
buf \U$58682 ( \58657 , \58311 );
or \U$58683 ( \58658 , \58656 , \58657 );
buf \U$58684 ( \58659 , \58185 );
nand \U$58685 ( \58660 , \58658 , \58659 );
buf \U$58686 ( \58661 , \58660 );
buf \U$58687 ( \58662 , \58661 );
nand \U$58688 ( \58663 , \58655 , \58662 );
buf \U$58689 ( \58664 , \58663 );
buf \U$58690 ( \58665 , \58664 );
not \U$58691 ( \58666 , \58665 );
or \U$58692 ( \58667 , \58650 , \58666 );
buf \U$58693 ( \58668 , \58664 );
buf \U$58694 ( \58669 , \58648 );
or \U$58695 ( \58670 , \58668 , \58669 );
nand \U$58696 ( \58671 , \58667 , \58670 );
buf \U$58697 ( \58672 , \58671 );
buf \U$58698 ( \58673 , \58672 );
xor \U$58699 ( \58674 , \57771 , \57802 );
xor \U$58700 ( \58675 , \58674 , \57815 );
buf \U$58701 ( \58676 , \58675 );
buf \U$58702 ( \58677 , \58676 );
not \U$58703 ( \58678 , \58677 );
buf \U$58704 ( \58679 , \58678 );
buf \U$58705 ( \58680 , \58679 );
and \U$58706 ( \58681 , \58673 , \58680 );
not \U$58707 ( \58682 , \58673 );
buf \U$58708 ( \58683 , \58676 );
and \U$58709 ( \58684 , \58682 , \58683 );
nor \U$58710 ( \58685 , \58681 , \58684 );
buf \U$58711 ( \58686 , \58685 );
buf \U$58712 ( \58687 , \58686 );
nand \U$58713 ( \58688 , \58643 , \58687 );
buf \U$58714 ( \58689 , \58688 );
buf \U$58715 ( \58690 , \58689 );
buf \U$58716 ( \58691 , \58645 );
not \U$58717 ( \58692 , \58691 );
buf \U$58718 ( \58693 , \58664 );
not \U$58719 ( \58694 , \58693 );
or \U$58720 ( \58695 , \58692 , \58694 );
buf \U$58721 ( \58696 , \58676 );
buf \U$58722 ( \58697 , \58664 );
not \U$58723 ( \58698 , \58697 );
buf \U$58724 ( \58699 , \58648 );
nand \U$58725 ( \58700 , \58698 , \58699 );
buf \U$58726 ( \58701 , \58700 );
buf \U$58727 ( \58702 , \58701 );
nand \U$58728 ( \58703 , \58696 , \58702 );
buf \U$58729 ( \58704 , \58703 );
buf \U$58730 ( \58705 , \58704 );
nand \U$58731 ( \58706 , \58695 , \58705 );
buf \U$58732 ( \58707 , \58706 );
buf \U$58733 ( \58708 , \58707 );
not \U$58734 ( \58709 , \58708 );
buf \U$58735 ( \58710 , \57836 );
buf \U$58736 ( \58711 , \57819 );
xor \U$58737 ( \58712 , \58710 , \58711 );
buf \U$58738 ( \58713 , \57843 );
xnor \U$58739 ( \58714 , \58712 , \58713 );
buf \U$58740 ( \58715 , \58714 );
buf \U$58741 ( \58716 , \58715 );
nand \U$58742 ( \58717 , \58709 , \58716 );
buf \U$58743 ( \58718 , \58717 );
buf \U$58744 ( \58719 , \58718 );
and \U$58745 ( \58720 , \58690 , \58719 );
buf \U$58746 ( \58721 , \58720 );
buf \U$58747 ( \58722 , \58721 );
xor \U$58748 ( \58723 , \58291 , \58269 );
buf \U$58749 ( \58724 , \58723 );
buf \U$58750 ( \58725 , \58300 );
not \U$58751 ( \58726 , \58725 );
buf \U$58752 ( \58727 , \58726 );
buf \U$58753 ( \58728 , \58727 );
and \U$58754 ( \58729 , \58724 , \58728 );
not \U$58755 ( \58730 , \58724 );
buf \U$58756 ( \58731 , \58300 );
and \U$58757 ( \58732 , \58730 , \58731 );
or \U$58758 ( \58733 , \58729 , \58732 );
buf \U$58759 ( \58734 , \58733 );
buf \U$58760 ( \58735 , \58734 );
not \U$58761 ( \58736 , \58735 );
xor \U$58762 ( \58737 , \58081 , \58098 );
xor \U$58763 ( \58738 , \58737 , \58112 );
buf \U$58764 ( \58739 , \58738 );
buf \U$58765 ( \58740 , \58739 );
xor \U$58766 ( \58741 , \58216 , \58233 );
xor \U$58767 ( \58742 , \58741 , \58250 );
buf \U$58768 ( \58743 , \58742 );
buf \U$58769 ( \58744 , \58743 );
xor \U$58770 ( \58745 , \58740 , \58744 );
buf \U$58771 ( \58746 , RIc0d8c80_48);
buf \U$58772 ( \58747 , RIc0dafa8_123);
xor \U$58773 ( \58748 , \58746 , \58747 );
buf \U$58774 ( \58749 , \58748 );
buf \U$58775 ( \58750 , \58749 );
not \U$58776 ( \58751 , \58750 );
buf \U$58777 ( \58752 , \14982 );
not \U$58778 ( \58753 , \58752 );
or \U$58779 ( \58754 , \58751 , \58753 );
buf \U$58780 ( \58755 , \16692 );
buf \U$58781 ( \58756 , \58160 );
nand \U$58782 ( \58757 , \58755 , \58756 );
buf \U$58783 ( \58758 , \58757 );
buf \U$58784 ( \58759 , \58758 );
nand \U$58785 ( \58760 , \58754 , \58759 );
buf \U$58786 ( \58761 , \58760 );
buf \U$58787 ( \58762 , \58761 );
not \U$58788 ( \58763 , \58762 );
xor \U$58789 ( \58764 , \58362 , \58379 );
buf \U$58790 ( \58765 , \58764 );
buf \U$58791 ( \58766 , \58765 );
not \U$58792 ( \58767 , \58766 );
or \U$58793 ( \58768 , \58763 , \58767 );
buf \U$58794 ( \58769 , \58765 );
buf \U$58795 ( \58770 , \58761 );
or \U$58796 ( \58771 , \58769 , \58770 );
buf \U$58797 ( \58772 , \12342 );
buf \U$58798 ( \58773 , RIc0d9400_64);
and \U$58799 ( \58774 , \58772 , \58773 );
buf \U$58800 ( \58775 , \58774 );
buf \U$58801 ( \58776 , \58775 );
buf \U$58802 ( \58777 , RIc0d8de8_51);
buf \U$58803 ( \58778 , RIc0daeb8_121);
xor \U$58804 ( \58779 , \58777 , \58778 );
buf \U$58805 ( \58780 , \58779 );
buf \U$58806 ( \58781 , \58780 );
not \U$58807 ( \58782 , \58781 );
buf \U$58808 ( \58783 , \13310 );
not \U$58809 ( \58784 , \58783 );
or \U$58810 ( \58785 , \58782 , \58784 );
buf \U$58811 ( \58786 , \16386 );
buf \U$58812 ( \58787 , \58386 );
nand \U$58813 ( \58788 , \58786 , \58787 );
buf \U$58814 ( \58789 , \58788 );
buf \U$58815 ( \58790 , \58789 );
nand \U$58816 ( \58791 , \58785 , \58790 );
buf \U$58817 ( \58792 , \58791 );
buf \U$58818 ( \58793 , \58792 );
xor \U$58819 ( \58794 , \58776 , \58793 );
buf \U$58820 ( \58795 , RIc0daa08_111);
buf \U$58821 ( \58796 , RIc0d9298_61);
xor \U$58822 ( \58797 , \58795 , \58796 );
buf \U$58823 ( \58798 , \58797 );
buf \U$58824 ( \58799 , \58798 );
not \U$58825 ( \58800 , \58799 );
buf \U$58826 ( \58801 , \18306 );
not \U$58827 ( \58802 , \58801 );
or \U$58828 ( \58803 , \58800 , \58802 );
buf \U$58829 ( \58804 , \58556 );
not \U$58830 ( \58805 , \58804 );
buf \U$58831 ( \58806 , \18312 );
nand \U$58832 ( \58807 , \58805 , \58806 );
buf \U$58833 ( \58808 , \58807 );
buf \U$58834 ( \58809 , \58808 );
nand \U$58835 ( \58810 , \58803 , \58809 );
buf \U$58836 ( \58811 , \58810 );
buf \U$58837 ( \58812 , \58811 );
and \U$58838 ( \58813 , \58794 , \58812 );
and \U$58839 ( \58814 , \58776 , \58793 );
or \U$58840 ( \58815 , \58813 , \58814 );
buf \U$58841 ( \58816 , \58815 );
buf \U$58842 ( \58817 , \58816 );
nand \U$58843 ( \58818 , \58771 , \58817 );
buf \U$58844 ( \58819 , \58818 );
buf \U$58845 ( \58820 , \58819 );
nand \U$58846 ( \58821 , \58768 , \58820 );
buf \U$58847 ( \58822 , \58821 );
buf \U$58848 ( \58823 , \58822 );
and \U$58849 ( \58824 , \58745 , \58823 );
and \U$58850 ( \58825 , \58740 , \58744 );
or \U$58851 ( \58826 , \58824 , \58825 );
buf \U$58852 ( \58827 , \58826 );
buf \U$58853 ( \58828 , \58827 );
xor \U$58854 ( \58829 , \58341 , \58345 );
xor \U$58855 ( \58830 , \58829 , \58509 );
buf \U$58856 ( \58831 , \58830 );
buf \U$58857 ( \58832 , \58831 );
xor \U$58858 ( \58833 , \58828 , \58832 );
xor \U$58859 ( \58834 , \58597 , \58601 );
xor \U$58860 ( \58835 , \58834 , \58621 );
buf \U$58861 ( \58836 , \58835 );
buf \U$58862 ( \58837 , \58836 );
and \U$58863 ( \58838 , \58833 , \58837 );
and \U$58864 ( \58839 , \58828 , \58832 );
or \U$58865 ( \58840 , \58838 , \58839 );
buf \U$58866 ( \58841 , \58840 );
buf \U$58867 ( \58842 , \58841 );
not \U$58868 ( \58843 , \58842 );
or \U$58869 ( \58844 , \58736 , \58843 );
buf \U$58870 ( \58845 , \58841 );
buf \U$58871 ( \58846 , \58734 );
or \U$58872 ( \58847 , \58845 , \58846 );
xor \U$58873 ( \58848 , \58514 , \58626 );
xor \U$58874 ( \58849 , \58848 , \58631 );
buf \U$58875 ( \58850 , \58849 );
buf \U$58876 ( \58851 , \58850 );
nand \U$58877 ( \58852 , \58847 , \58851 );
buf \U$58878 ( \58853 , \58852 );
buf \U$58879 ( \58854 , \58853 );
nand \U$58880 ( \58855 , \58844 , \58854 );
buf \U$58881 ( \58856 , \58855 );
buf \U$58882 ( \58857 , \58856 );
not \U$58883 ( \58858 , \58857 );
buf \U$58884 ( \58859 , \57950 );
buf \U$58885 ( \58860 , \58635 );
xor \U$58886 ( \58861 , \58859 , \58860 );
buf \U$58887 ( \58862 , \58317 );
xnor \U$58888 ( \58863 , \58861 , \58862 );
buf \U$58889 ( \58864 , \58863 );
buf \U$58890 ( \58865 , \58864 );
nand \U$58891 ( \58866 , \58858 , \58865 );
buf \U$58892 ( \58867 , \58866 );
buf \U$58893 ( \58868 , \58867 );
buf \U$58894 ( \58869 , \58734 );
buf \U$58895 ( \58870 , \58841 );
xor \U$58896 ( \58871 , \58869 , \58870 );
buf \U$58897 ( \58872 , \58850 );
xnor \U$58898 ( \58873 , \58871 , \58872 );
buf \U$58899 ( \58874 , \58873 );
buf \U$58900 ( \58875 , \58874 );
buf \U$58901 ( \58876 , \58578 );
buf \U$58902 ( \58877 , \58574 );
and \U$58903 ( \58878 , \58876 , \58877 );
not \U$58904 ( \58879 , \58876 );
buf \U$58905 ( \58880 , \58571 );
and \U$58906 ( \58881 , \58879 , \58880 );
nor \U$58907 ( \58882 , \58878 , \58881 );
buf \U$58908 ( \58883 , \58882 );
buf \U$58909 ( \58884 , \58883 );
buf \U$58910 ( \58885 , \58584 );
and \U$58911 ( \58886 , \58884 , \58885 );
not \U$58912 ( \58887 , \58884 );
buf \U$58913 ( \58888 , \58584 );
not \U$58914 ( \58889 , \58888 );
buf \U$58915 ( \58890 , \58889 );
buf \U$58916 ( \58891 , \58890 );
and \U$58917 ( \58892 , \58887 , \58891 );
nor \U$58918 ( \58893 , \58886 , \58892 );
buf \U$58919 ( \58894 , \58893 );
buf \U$58920 ( \58895 , \58894 );
xor \U$58921 ( \58896 , \58740 , \58744 );
xor \U$58922 ( \58897 , \58896 , \58823 );
buf \U$58923 ( \58898 , \58897 );
buf \U$58924 ( \58899 , \58898 );
xor \U$58925 ( \58900 , \58895 , \58899 );
buf \U$58926 ( \58901 , RIc0d9130_58);
buf \U$58927 ( \58902 , RIc0dabe8_115);
xor \U$58928 ( \58903 , \58901 , \58902 );
buf \U$58929 ( \58904 , \58903 );
buf \U$58930 ( \58905 , \58904 );
not \U$58931 ( \58906 , \58905 );
buf \U$58932 ( \58907 , \14186 );
not \U$58933 ( \58908 , \58907 );
or \U$58934 ( \58909 , \58906 , \58908 );
buf \U$58935 ( \58910 , \12303 );
buf \U$58936 ( \58911 , RIc0d90b8_57);
buf \U$58937 ( \58912 , RIc0dabe8_115);
xor \U$58938 ( \58913 , \58911 , \58912 );
buf \U$58939 ( \58914 , \58913 );
buf \U$58940 ( \58915 , \58914 );
nand \U$58941 ( \58916 , \58910 , \58915 );
buf \U$58942 ( \58917 , \58916 );
buf \U$58943 ( \58918 , \58917 );
nand \U$58944 ( \58919 , \58909 , \58918 );
buf \U$58945 ( \58920 , \58919 );
buf \U$58946 ( \58921 , \58920 );
not \U$58947 ( \58922 , \58921 );
buf \U$58948 ( \58923 , RIc0d8e60_52);
buf \U$58949 ( \58924 , RIc0daeb8_121);
xor \U$58950 ( \58925 , \58923 , \58924 );
buf \U$58951 ( \58926 , \58925 );
buf \U$58952 ( \58927 , \58926 );
not \U$58953 ( \58928 , \58927 );
buf \U$58954 ( \58929 , \12971 );
not \U$58955 ( \58930 , \58929 );
or \U$58956 ( \58931 , \58928 , \58930 );
buf \U$58957 ( \58932 , \12975 );
buf \U$58958 ( \58933 , \58780 );
nand \U$58959 ( \58934 , \58932 , \58933 );
buf \U$58960 ( \58935 , \58934 );
buf \U$58961 ( \58936 , \58935 );
nand \U$58962 ( \58937 , \58931 , \58936 );
buf \U$58963 ( \58938 , \58937 );
buf \U$58964 ( \58939 , \58938 );
not \U$58965 ( \58940 , \58939 );
or \U$58966 ( \58941 , \58922 , \58940 );
buf \U$58967 ( \58942 , \58920 );
not \U$58968 ( \58943 , \58942 );
buf \U$58969 ( \58944 , \58938 );
not \U$58970 ( \58945 , \58944 );
buf \U$58971 ( \58946 , \58945 );
buf \U$58972 ( \58947 , \58946 );
nand \U$58973 ( \58948 , \58943 , \58947 );
buf \U$58974 ( \58949 , \58948 );
buf \U$58975 ( \58950 , \58949 );
buf \U$58976 ( \58951 , RIc0d9400_64);
buf \U$58977 ( \58952 , RIc0da918_109);
xor \U$58978 ( \58953 , \58951 , \58952 );
buf \U$58979 ( \58954 , \58953 );
buf \U$58980 ( \58955 , \58954 );
not \U$58981 ( \58956 , \58955 );
buf \U$58982 ( \58957 , \27660 );
not \U$58983 ( \58958 , \58957 );
or \U$58984 ( \58959 , \58956 , \58958 );
buf \U$58985 ( \58960 , \13426 );
buf \U$58986 ( \58961 , RIc0da918_109);
buf \U$58987 ( \58962 , RIc0d9388_63);
xor \U$58988 ( \58963 , \58961 , \58962 );
buf \U$58989 ( \58964 , \58963 );
buf \U$58990 ( \58965 , \58964 );
nand \U$58991 ( \58966 , \58960 , \58965 );
buf \U$58992 ( \58967 , \58966 );
buf \U$58993 ( \58968 , \58967 );
nand \U$58994 ( \58969 , \58959 , \58968 );
buf \U$58995 ( \58970 , \58969 );
buf \U$58996 ( \58971 , \58970 );
nand \U$58997 ( \58972 , \58950 , \58971 );
buf \U$58998 ( \58973 , \58972 );
buf \U$58999 ( \58974 , \58973 );
nand \U$59000 ( \58975 , \58941 , \58974 );
buf \U$59001 ( \58976 , \58975 );
buf \U$59002 ( \58977 , \58976 );
not \U$59003 ( \58978 , \58977 );
xor \U$59004 ( \58979 , RIc0db188_127, RIc0d8b90_46);
buf \U$59005 ( \58980 , \58979 );
not \U$59006 ( \58981 , \58980 );
buf \U$59007 ( \58982 , \58521 );
not \U$59008 ( \58983 , \58982 );
or \U$59009 ( \58984 , \58981 , \58983 );
buf \U$59010 ( \58985 , RIc0d8b18_45);
buf \U$59011 ( \58986 , RIc0db188_127);
xor \U$59012 ( \58987 , \58985 , \58986 );
buf \U$59013 ( \58988 , \58987 );
buf \U$59014 ( \58989 , \58988 );
buf \U$59015 ( \58990 , RIc0db200_128);
nand \U$59016 ( \58991 , \58989 , \58990 );
buf \U$59017 ( \58992 , \58991 );
buf \U$59018 ( \58993 , \58992 );
nand \U$59019 ( \58994 , \58984 , \58993 );
buf \U$59020 ( \58995 , \58994 );
buf \U$59021 ( \58996 , \58995 );
not \U$59022 ( \58997 , \58996 );
buf \U$59023 ( \58998 , RIc0daaf8_113);
buf \U$59024 ( \58999 , RIc0d9220_60);
xor \U$59025 ( \59000 , \58998 , \58999 );
buf \U$59026 ( \59001 , \59000 );
buf \U$59027 ( \59002 , \59001 );
not \U$59028 ( \59003 , \59002 );
buf \U$59029 ( \59004 , \16989 );
not \U$59030 ( \59005 , \59004 );
or \U$59031 ( \59006 , \59003 , \59005 );
buf \U$59032 ( \59007 , \16995 );
buf \U$59033 ( \59008 , RIc0daaf8_113);
buf \U$59034 ( \59009 , RIc0d91a8_59);
xor \U$59035 ( \59010 , \59008 , \59009 );
buf \U$59036 ( \59011 , \59010 );
buf \U$59037 ( \59012 , \59011 );
nand \U$59038 ( \59013 , \59007 , \59012 );
buf \U$59039 ( \59014 , \59013 );
buf \U$59040 ( \59015 , \59014 );
nand \U$59041 ( \59016 , \59006 , \59015 );
buf \U$59042 ( \59017 , \59016 );
buf \U$59043 ( \59018 , \59017 );
not \U$59044 ( \59019 , \59018 );
or \U$59045 ( \59020 , \58997 , \59019 );
buf \U$59046 ( \59021 , \59017 );
buf \U$59047 ( \59022 , \58995 );
or \U$59048 ( \59023 , \59021 , \59022 );
xor \U$59049 ( \59024 , RIc0dacd8_117, RIc0d9040_56);
buf \U$59050 ( \59025 , \59024 );
not \U$59051 ( \59026 , \59025 );
buf \U$59052 ( \59027 , \12929 );
not \U$59053 ( \59028 , \59027 );
or \U$59054 ( \59029 , \59026 , \59028 );
buf \U$59055 ( \59030 , \22356 );
buf \U$59056 ( \59031 , RIc0dacd8_117);
buf \U$59057 ( \59032 , RIc0d8fc8_55);
xor \U$59058 ( \59033 , \59031 , \59032 );
buf \U$59059 ( \59034 , \59033 );
buf \U$59060 ( \59035 , \59034 );
nand \U$59061 ( \59036 , \59030 , \59035 );
buf \U$59062 ( \59037 , \59036 );
buf \U$59063 ( \59038 , \59037 );
nand \U$59064 ( \59039 , \59029 , \59038 );
buf \U$59065 ( \59040 , \59039 );
buf \U$59066 ( \59041 , \59040 );
nand \U$59067 ( \59042 , \59023 , \59041 );
buf \U$59068 ( \59043 , \59042 );
buf \U$59069 ( \59044 , \59043 );
nand \U$59070 ( \59045 , \59020 , \59044 );
buf \U$59071 ( \59046 , \59045 );
buf \U$59072 ( \59047 , \59046 );
not \U$59073 ( \59048 , \59047 );
or \U$59074 ( \59049 , \58978 , \59048 );
or \U$59075 ( \59050 , \59046 , \58976 );
buf \U$59076 ( \59051 , RIc0db098_125);
buf \U$59077 ( \59052 , RIc0d8c80_48);
xor \U$59078 ( \59053 , \59051 , \59052 );
buf \U$59079 ( \59054 , \59053 );
buf \U$59080 ( \59055 , \59054 );
not \U$59081 ( \59056 , \59055 );
buf \U$59082 ( \59057 , \15789 );
not \U$59083 ( \59058 , \59057 );
or \U$59084 ( \59059 , \59056 , \59058 );
buf \U$59085 ( \59060 , \15793 );
xor \U$59086 ( \59061 , RIc0db098_125, RIc0d8c08_47);
buf \U$59087 ( \59062 , \59061 );
nand \U$59088 ( \59063 , \59060 , \59062 );
buf \U$59089 ( \59064 , \59063 );
buf \U$59090 ( \59065 , \59064 );
nand \U$59091 ( \59066 , \59059 , \59065 );
buf \U$59092 ( \59067 , \59066 );
buf \U$59093 ( \59068 , \59067 );
buf \U$59094 ( \59069 , RIc0d8d70_50);
buf \U$59095 ( \59070 , RIc0dafa8_123);
xor \U$59096 ( \59071 , \59069 , \59070 );
buf \U$59097 ( \59072 , \59071 );
buf \U$59098 ( \59073 , \59072 );
not \U$59099 ( \59074 , \59073 );
buf \U$59100 ( \59075 , \14982 );
not \U$59101 ( \59076 , \59075 );
or \U$59102 ( \59077 , \59074 , \59076 );
buf \U$59103 ( \59078 , \16692 );
xor \U$59104 ( \59079 , RIc0dafa8_123, RIc0d8cf8_49);
buf \U$59105 ( \59080 , \59079 );
nand \U$59106 ( \59081 , \59078 , \59080 );
buf \U$59107 ( \59082 , \59081 );
buf \U$59108 ( \59083 , \59082 );
nand \U$59109 ( \59084 , \59077 , \59083 );
buf \U$59110 ( \59085 , \59084 );
buf \U$59111 ( \59086 , \59085 );
xor \U$59112 ( \59087 , \59068 , \59086 );
buf \U$59113 ( \59088 , \55702 );
buf \U$59114 ( \59089 , RIc0dadc8_119);
buf \U$59115 ( \59090 , RIc0d8f50_54);
xnor \U$59116 ( \59091 , \59089 , \59090 );
buf \U$59117 ( \59092 , \59091 );
buf \U$59118 ( \59093 , \59092 );
or \U$59119 ( \59094 , \59088 , \59093 );
buf \U$59120 ( \59095 , \22798 );
buf \U$59121 ( \59096 , RIc0d8ed8_53);
buf \U$59122 ( \59097 , RIc0dadc8_119);
xor \U$59123 ( \59098 , \59096 , \59097 );
buf \U$59124 ( \59099 , \59098 );
buf \U$59125 ( \59100 , \59099 );
not \U$59126 ( \59101 , \59100 );
buf \U$59127 ( \59102 , \59101 );
buf \U$59128 ( \59103 , \59102 );
or \U$59129 ( \59104 , \59095 , \59103 );
nand \U$59130 ( \59105 , \59094 , \59104 );
buf \U$59131 ( \59106 , \59105 );
buf \U$59132 ( \59107 , \59106 );
and \U$59133 ( \59108 , \59087 , \59107 );
and \U$59134 ( \59109 , \59068 , \59086 );
or \U$59135 ( \59110 , \59108 , \59109 );
buf \U$59136 ( \59111 , \59110 );
nand \U$59137 ( \59112 , \59050 , \59111 );
buf \U$59138 ( \59113 , \59112 );
nand \U$59139 ( \59114 , \59049 , \59113 );
buf \U$59140 ( \59115 , \59114 );
buf \U$59141 ( \59116 , \59115 );
not \U$59142 ( \59117 , \59116 );
buf \U$59143 ( \59118 , \58761 );
not \U$59144 ( \59119 , \59118 );
buf \U$59145 ( \59120 , \59119 );
buf \U$59146 ( \59121 , \59120 );
not \U$59147 ( \59122 , \59121 );
buf \U$59148 ( \59123 , \58765 );
not \U$59149 ( \59124 , \59123 );
or \U$59150 ( \59125 , \59122 , \59124 );
buf \U$59151 ( \59126 , \58765 );
buf \U$59152 ( \59127 , \59120 );
or \U$59153 ( \59128 , \59126 , \59127 );
nand \U$59154 ( \59129 , \59125 , \59128 );
buf \U$59155 ( \59130 , \59129 );
buf \U$59156 ( \59131 , \59130 );
buf \U$59157 ( \59132 , \58816 );
xnor \U$59158 ( \59133 , \59131 , \59132 );
buf \U$59159 ( \59134 , \59133 );
buf \U$59160 ( \59135 , \59134 );
not \U$59161 ( \59136 , \59135 );
buf \U$59162 ( \59137 , \59136 );
buf \U$59163 ( \59138 , \59137 );
not \U$59164 ( \59139 , \59138 );
or \U$59165 ( \59140 , \59117 , \59139 );
buf \U$59166 ( \59141 , \58988 );
not \U$59167 ( \59142 , \59141 );
not \U$59168 ( \59143 , \43780 );
not \U$59169 ( \59144 , \59143 );
buf \U$59170 ( \59145 , \59144 );
not \U$59171 ( \59146 , \59145 );
or \U$59172 ( \59147 , \59142 , \59146 );
buf \U$59173 ( \59148 , \58518 );
buf \U$59174 ( \59149 , RIc0db200_128);
nand \U$59175 ( \59150 , \59148 , \59149 );
buf \U$59176 ( \59151 , \59150 );
buf \U$59177 ( \59152 , \59151 );
nand \U$59178 ( \59153 , \59147 , \59152 );
buf \U$59179 ( \59154 , \59153 );
buf \U$59180 ( \59155 , \59154 );
buf \U$59181 ( \59156 , \59034 );
not \U$59182 ( \59157 , \59156 );
buf \U$59183 ( \59158 , \22350 );
not \U$59184 ( \59159 , \59158 );
or \U$59185 ( \59160 , \59157 , \59159 );
buf \U$59186 ( \59161 , \16559 );
buf \U$59187 ( \59162 , \58403 );
nand \U$59188 ( \59163 , \59161 , \59162 );
buf \U$59189 ( \59164 , \59163 );
buf \U$59190 ( \59165 , \59164 );
nand \U$59191 ( \59166 , \59160 , \59165 );
buf \U$59192 ( \59167 , \59166 );
buf \U$59193 ( \59168 , \59167 );
xor \U$59194 ( \59169 , \59155 , \59168 );
buf \U$59195 ( \59170 , \51095 );
not \U$59196 ( \59171 , \59170 );
buf \U$59197 ( \59172 , \59061 );
not \U$59198 ( \59173 , \59172 );
or \U$59199 ( \59174 , \59171 , \59173 );
buf \U$59200 ( \59175 , \18699 );
buf \U$59201 ( \59176 , \58464 );
or \U$59202 ( \59177 , \59175 , \59176 );
nand \U$59203 ( \59178 , \59174 , \59177 );
buf \U$59204 ( \59179 , \59178 );
buf \U$59205 ( \59180 , \59179 );
and \U$59206 ( \59181 , \59169 , \59180 );
and \U$59207 ( \59182 , \59155 , \59168 );
or \U$59208 ( \59183 , \59181 , \59182 );
buf \U$59209 ( \59184 , \59183 );
buf \U$59210 ( \59185 , \59184 );
not \U$59211 ( \59186 , \59185 );
not \U$59212 ( \59187 , \58914 );
nor \U$59213 ( \59188 , \59187 , \22595 );
buf \U$59214 ( \59189 , \59188 );
buf \U$59215 ( \59190 , \29865 );
buf \U$59216 ( \59191 , \58419 );
nor \U$59217 ( \59192 , \59190 , \59191 );
buf \U$59218 ( \59193 , \59192 );
buf \U$59219 ( \59194 , \59193 );
nor \U$59220 ( \59195 , \59189 , \59194 );
buf \U$59221 ( \59196 , \59195 );
buf \U$59222 ( \59197 , \59196 );
not \U$59223 ( \59198 , \59197 );
buf \U$59224 ( \59199 , \59011 );
not \U$59225 ( \59200 , \59199 );
buf \U$59226 ( \59201 , \33224 );
not \U$59227 ( \59202 , \59201 );
or \U$59228 ( \59203 , \59200 , \59202 );
buf \U$59229 ( \59204 , \12410 );
buf \U$59230 ( \59205 , \58445 );
nand \U$59231 ( \59206 , \59204 , \59205 );
buf \U$59232 ( \59207 , \59206 );
buf \U$59233 ( \59208 , \59207 );
nand \U$59234 ( \59209 , \59203 , \59208 );
buf \U$59235 ( \59210 , \59209 );
buf \U$59236 ( \59211 , \59210 );
not \U$59237 ( \59212 , \59211 );
buf \U$59238 ( \59213 , \59212 );
buf \U$59239 ( \59214 , \59213 );
not \U$59240 ( \59215 , \59214 );
or \U$59241 ( \59216 , \59198 , \59215 );
buf \U$59242 ( \59217 , \58964 );
not \U$59243 ( \59218 , \59217 );
buf \U$59244 ( \59219 , \27660 );
not \U$59245 ( \59220 , \59219 );
or \U$59246 ( \59221 , \59218 , \59220 );
buf \U$59247 ( \59222 , \16232 );
buf \U$59248 ( \59223 , \58366 );
nand \U$59249 ( \59224 , \59222 , \59223 );
buf \U$59250 ( \59225 , \59224 );
buf \U$59251 ( \59226 , \59225 );
nand \U$59252 ( \59227 , \59221 , \59226 );
buf \U$59253 ( \59228 , \59227 );
buf \U$59254 ( \59229 , \59228 );
nand \U$59255 ( \59230 , \59216 , \59229 );
buf \U$59256 ( \59231 , \59230 );
buf \U$59257 ( \59232 , \59231 );
buf \U$59258 ( \59233 , \59210 );
buf \U$59259 ( \59234 , \59196 );
not \U$59260 ( \59235 , \59234 );
buf \U$59261 ( \59236 , \59235 );
buf \U$59262 ( \59237 , \59236 );
nand \U$59263 ( \59238 , \59233 , \59237 );
buf \U$59264 ( \59239 , \59238 );
buf \U$59265 ( \59240 , \59239 );
nand \U$59266 ( \59241 , \59232 , \59240 );
buf \U$59267 ( \59242 , \59241 );
buf \U$59268 ( \59243 , \59242 );
not \U$59269 ( \59244 , \59243 );
buf \U$59270 ( \59245 , \59244 );
buf \U$59271 ( \59246 , \59245 );
not \U$59272 ( \59247 , \59246 );
or \U$59273 ( \59248 , \59186 , \59247 );
buf \U$59274 ( \59249 , \59184 );
buf \U$59275 ( \59250 , \59245 );
or \U$59276 ( \59251 , \59249 , \59250 );
nand \U$59277 ( \59252 , \59248 , \59251 );
buf \U$59278 ( \59253 , \59252 );
buf \U$59279 ( \59254 , \59253 );
xor \U$59280 ( \59255 , \58399 , \58417 );
xor \U$59281 ( \59256 , \59255 , \58435 );
buf \U$59282 ( \59257 , \59256 );
buf \U$59283 ( \59258 , \59257 );
xnor \U$59284 ( \59259 , \59254 , \59258 );
buf \U$59285 ( \59260 , \59259 );
buf \U$59286 ( \59261 , \59260 );
not \U$59287 ( \59262 , \59261 );
buf \U$59288 ( \59263 , \59115 );
not \U$59289 ( \59264 , \59263 );
buf \U$59290 ( \59265 , \59134 );
nand \U$59291 ( \59266 , \59264 , \59265 );
buf \U$59292 ( \59267 , \59266 );
buf \U$59293 ( \59268 , \59267 );
nand \U$59294 ( \59269 , \59262 , \59268 );
buf \U$59295 ( \59270 , \59269 );
buf \U$59296 ( \59271 , \59270 );
nand \U$59297 ( \59272 , \59140 , \59271 );
buf \U$59298 ( \59273 , \59272 );
buf \U$59299 ( \59274 , \59273 );
and \U$59300 ( \59275 , \58900 , \59274 );
and \U$59301 ( \59276 , \58895 , \58899 );
or \U$59302 ( \59277 , \59275 , \59276 );
buf \U$59303 ( \59278 , \59277 );
buf \U$59304 ( \59279 , \59278 );
buf \U$59305 ( \59280 , \59099 );
not \U$59306 ( \59281 , \59280 );
buf \U$59307 ( \59282 , \14569 );
not \U$59308 ( \59283 , \59282 );
or \U$59309 ( \59284 , \59281 , \59283 );
buf \U$59310 ( \59285 , \13005 );
buf \U$59311 ( \59286 , \58537 );
nand \U$59312 ( \59287 , \59285 , \59286 );
buf \U$59313 ( \59288 , \59287 );
buf \U$59314 ( \59289 , \59288 );
nand \U$59315 ( \59290 , \59284 , \59289 );
buf \U$59316 ( \59291 , \59290 );
buf \U$59317 ( \59292 , \59291 );
not \U$59318 ( \59293 , \59292 );
buf \U$59319 ( \59294 , \59079 );
not \U$59320 ( \59295 , \59294 );
buf \U$59321 ( \59296 , \14982 );
not \U$59322 ( \59297 , \59296 );
or \U$59323 ( \59298 , \59295 , \59297 );
buf \U$59324 ( \59299 , \14278 );
buf \U$59325 ( \59300 , \58749 );
nand \U$59326 ( \59301 , \59299 , \59300 );
buf \U$59327 ( \59302 , \59301 );
buf \U$59328 ( \59303 , \59302 );
nand \U$59329 ( \59304 , \59298 , \59303 );
buf \U$59330 ( \59305 , \59304 );
buf \U$59331 ( \59306 , \59305 );
not \U$59332 ( \59307 , \59306 );
or \U$59333 ( \59308 , \59293 , \59307 );
buf \U$59334 ( \59309 , \59305 );
buf \U$59335 ( \59310 , \59291 );
or \U$59336 ( \59311 , \59309 , \59310 );
buf \U$59337 ( \59312 , RIc0daa08_111);
buf \U$59338 ( \59313 , RIc0d9310_62);
xor \U$59339 ( \59314 , \59312 , \59313 );
buf \U$59340 ( \59315 , \59314 );
buf \U$59341 ( \59316 , \59315 );
not \U$59342 ( \59317 , \59316 );
buf \U$59343 ( \59318 , \12529 );
not \U$59344 ( \59319 , \59318 );
or \U$59345 ( \59320 , \59317 , \59319 );
buf \U$59346 ( \59321 , \25649 );
buf \U$59347 ( \59322 , \58798 );
nand \U$59348 ( \59323 , \59321 , \59322 );
buf \U$59349 ( \59324 , \59323 );
buf \U$59350 ( \59325 , \59324 );
nand \U$59351 ( \59326 , \59320 , \59325 );
buf \U$59352 ( \59327 , \59326 );
buf \U$59353 ( \59328 , \59327 );
buf \U$59354 ( \59329 , RIc0d9400_64);
buf \U$59355 ( \59330 , RIc0da990_110);
or \U$59356 ( \59331 , \59329 , \59330 );
buf \U$59357 ( \59332 , RIc0daa08_111);
nand \U$59358 ( \59333 , \59331 , \59332 );
buf \U$59359 ( \59334 , \59333 );
buf \U$59360 ( \59335 , \59334 );
buf \U$59361 ( \59336 , RIc0d9400_64);
buf \U$59362 ( \59337 , RIc0da990_110);
nand \U$59363 ( \59338 , \59336 , \59337 );
buf \U$59364 ( \59339 , \59338 );
buf \U$59365 ( \59340 , \59339 );
buf \U$59366 ( \59341 , RIc0da918_109);
nand \U$59367 ( \59342 , \59335 , \59340 , \59341 );
buf \U$59368 ( \59343 , \59342 );
buf \U$59369 ( \59344 , \59343 );
not \U$59370 ( \59345 , \59344 );
buf \U$59371 ( \59346 , \59345 );
buf \U$59372 ( \59347 , \59346 );
and \U$59373 ( \59348 , \59328 , \59347 );
buf \U$59374 ( \59349 , \59348 );
buf \U$59375 ( \59350 , \59349 );
nand \U$59376 ( \59351 , \59311 , \59350 );
buf \U$59377 ( \59352 , \59351 );
buf \U$59378 ( \59353 , \59352 );
nand \U$59379 ( \59354 , \59308 , \59353 );
buf \U$59380 ( \59355 , \59354 );
buf \U$59381 ( \59356 , \59355 );
xor \U$59382 ( \59357 , \58533 , \58550 );
xor \U$59383 ( \59358 , \59357 , \58567 );
buf \U$59384 ( \59359 , \59358 );
buf \U$59385 ( \59360 , \59359 );
xor \U$59386 ( \59361 , \59356 , \59360 );
xor \U$59387 ( \59362 , \58457 , \58497 );
buf \U$59388 ( \59363 , \59362 );
buf \U$59389 ( \59364 , \58471 );
xor \U$59390 ( \59365 , \59363 , \59364 );
buf \U$59391 ( \59366 , \59365 );
buf \U$59392 ( \59367 , \59366 );
and \U$59393 ( \59368 , \59361 , \59367 );
and \U$59394 ( \59369 , \59356 , \59360 );
or \U$59395 ( \59370 , \59368 , \59369 );
buf \U$59396 ( \59371 , \59370 );
buf \U$59397 ( \59372 , \59371 );
xor \U$59398 ( \59373 , \58382 , \58440 );
xor \U$59399 ( \59374 , \59373 , \58504 );
buf \U$59400 ( \59375 , \59374 );
buf \U$59401 ( \59376 , \59375 );
xor \U$59402 ( \59377 , \59372 , \59376 );
buf \U$59403 ( \59378 , \59184 );
not \U$59404 ( \59379 , \59378 );
buf \U$59405 ( \59380 , \59257 );
not \U$59406 ( \59381 , \59380 );
or \U$59407 ( \59382 , \59379 , \59381 );
buf \U$59408 ( \59383 , \59257 );
buf \U$59409 ( \59384 , \59184 );
or \U$59410 ( \59385 , \59383 , \59384 );
buf \U$59411 ( \59386 , \59242 );
nand \U$59412 ( \59387 , \59385 , \59386 );
buf \U$59413 ( \59388 , \59387 );
buf \U$59414 ( \59389 , \59388 );
nand \U$59415 ( \59390 , \59382 , \59389 );
buf \U$59416 ( \59391 , \59390 );
buf \U$59417 ( \59392 , \59391 );
and \U$59418 ( \59393 , \59377 , \59392 );
and \U$59419 ( \59394 , \59372 , \59376 );
or \U$59420 ( \59395 , \59393 , \59394 );
buf \U$59421 ( \59396 , \59395 );
buf \U$59422 ( \59397 , \59396 );
or \U$59423 ( \59398 , \59279 , \59397 );
xor \U$59424 ( \59399 , \58828 , \58832 );
xor \U$59425 ( \59400 , \59399 , \58837 );
buf \U$59426 ( \59401 , \59400 );
buf \U$59427 ( \59402 , \59401 );
nand \U$59428 ( \59403 , \59398 , \59402 );
buf \U$59429 ( \59404 , \59403 );
buf \U$59430 ( \59405 , \59404 );
buf \U$59431 ( \59406 , \59278 );
buf \U$59432 ( \59407 , \59396 );
nand \U$59433 ( \59408 , \59406 , \59407 );
buf \U$59434 ( \59409 , \59408 );
buf \U$59435 ( \59410 , \59409 );
and \U$59436 ( \59411 , \59405 , \59410 );
buf \U$59437 ( \59412 , \59411 );
buf \U$59438 ( \59413 , \59412 );
nand \U$59439 ( \59414 , \58875 , \59413 );
buf \U$59440 ( \59415 , \59414 );
buf \U$59441 ( \59416 , \59415 );
and \U$59442 ( \59417 , \58868 , \59416 );
buf \U$59443 ( \59418 , \59417 );
buf \U$59444 ( \59419 , \59418 );
nand \U$59445 ( \59420 , \58722 , \59419 );
buf \U$59446 ( \59421 , \59420 );
buf \U$59447 ( \59422 , \59421 );
nor \U$59448 ( \59423 , \57947 , \59422 );
buf \U$59449 ( \59424 , \59423 );
buf \U$59450 ( \59425 , \59424 );
not \U$59451 ( \59426 , \59425 );
xor \U$59452 ( \59427 , \59372 , \59376 );
xor \U$59453 ( \59428 , \59427 , \59392 );
buf \U$59454 ( \59429 , \59428 );
buf \U$59455 ( \59430 , \59429 );
xor \U$59456 ( \59431 , \58776 , \58793 );
xor \U$59457 ( \59432 , \59431 , \58812 );
buf \U$59458 ( \59433 , \59432 );
buf \U$59459 ( \59434 , \59433 );
xor \U$59460 ( \59435 , \59155 , \59168 );
xor \U$59461 ( \59436 , \59435 , \59180 );
buf \U$59462 ( \59437 , \59436 );
buf \U$59463 ( \59438 , \59437 );
xor \U$59464 ( \59439 , \59434 , \59438 );
buf \U$59465 ( \59440 , \59228 );
not \U$59466 ( \59441 , \59440 );
buf \U$59467 ( \59442 , \59213 );
not \U$59468 ( \59443 , \59442 );
or \U$59469 ( \59444 , \59441 , \59443 );
buf \U$59470 ( \59445 , \59213 );
buf \U$59471 ( \59446 , \59228 );
or \U$59472 ( \59447 , \59445 , \59446 );
nand \U$59473 ( \59448 , \59444 , \59447 );
buf \U$59474 ( \59449 , \59448 );
buf \U$59475 ( \59450 , \59449 );
buf \U$59476 ( \59451 , \59236 );
and \U$59477 ( \59452 , \59450 , \59451 );
not \U$59478 ( \59453 , \59450 );
buf \U$59479 ( \59454 , \59196 );
and \U$59480 ( \59455 , \59453 , \59454 );
nor \U$59481 ( \59456 , \59452 , \59455 );
buf \U$59482 ( \59457 , \59456 );
buf \U$59483 ( \59458 , \59457 );
and \U$59484 ( \59459 , \59439 , \59458 );
and \U$59485 ( \59460 , \59434 , \59438 );
or \U$59486 ( \59461 , \59459 , \59460 );
buf \U$59487 ( \59462 , \59461 );
buf \U$59488 ( \59463 , \59462 );
xor \U$59489 ( \59464 , \59356 , \59360 );
xor \U$59490 ( \59465 , \59464 , \59367 );
buf \U$59491 ( \59466 , \59465 );
buf \U$59492 ( \59467 , \59466 );
xor \U$59493 ( \59468 , \59463 , \59467 );
buf \U$59494 ( \59469 , \59260 );
not \U$59495 ( \59470 , \59469 );
buf \U$59496 ( \59471 , \59115 );
not \U$59497 ( \59472 , \59471 );
buf \U$59498 ( \59473 , \59134 );
not \U$59499 ( \59474 , \59473 );
or \U$59500 ( \59475 , \59472 , \59474 );
buf \U$59501 ( \59476 , \59134 );
buf \U$59502 ( \59477 , \59115 );
or \U$59503 ( \59478 , \59476 , \59477 );
nand \U$59504 ( \59479 , \59475 , \59478 );
buf \U$59505 ( \59480 , \59479 );
buf \U$59506 ( \59481 , \59480 );
not \U$59507 ( \59482 , \59481 );
or \U$59508 ( \59483 , \59470 , \59482 );
buf \U$59509 ( \59484 , \59260 );
buf \U$59510 ( \59485 , \59480 );
or \U$59511 ( \59486 , \59484 , \59485 );
nand \U$59512 ( \59487 , \59483 , \59486 );
buf \U$59513 ( \59488 , \59487 );
buf \U$59514 ( \59489 , \59488 );
and \U$59515 ( \59490 , \59468 , \59489 );
and \U$59516 ( \59491 , \59463 , \59467 );
or \U$59517 ( \59492 , \59490 , \59491 );
buf \U$59518 ( \59493 , \59492 );
buf \U$59519 ( \59494 , \59493 );
xor \U$59520 ( \59495 , \59430 , \59494 );
xor \U$59521 ( \59496 , \58895 , \58899 );
xor \U$59522 ( \59497 , \59496 , \59274 );
buf \U$59523 ( \59498 , \59497 );
buf \U$59524 ( \59499 , \59498 );
xor \U$59525 ( \59500 , \59495 , \59499 );
buf \U$59526 ( \59501 , \59500 );
buf \U$59527 ( \59502 , \59501 );
xor \U$59528 ( \59503 , \59305 , \59291 );
xor \U$59529 ( \59504 , \59503 , \59349 );
buf \U$59530 ( \59505 , \59504 );
buf \U$59531 ( \59506 , \59343 );
not \U$59532 ( \59507 , \59506 );
buf \U$59533 ( \59508 , \59327 );
not \U$59534 ( \59509 , \59508 );
or \U$59535 ( \59510 , \59507 , \59509 );
buf \U$59536 ( \59511 , \59327 );
buf \U$59537 ( \59512 , \59343 );
or \U$59538 ( \59513 , \59511 , \59512 );
nand \U$59539 ( \59514 , \59510 , \59513 );
buf \U$59540 ( \59515 , \59514 );
buf \U$59541 ( \59516 , \59515 );
buf \U$59542 ( \59517 , RIc0d90b8_57);
buf \U$59543 ( \59518 , RIc0dacd8_117);
xor \U$59544 ( \59519 , \59517 , \59518 );
buf \U$59545 ( \59520 , \59519 );
buf \U$59546 ( \59521 , \59520 );
not \U$59547 ( \59522 , \59521 );
buf \U$59548 ( \59523 , \12929 );
not \U$59549 ( \59524 , \59523 );
or \U$59550 ( \59525 , \59522 , \59524 );
buf \U$59551 ( \59526 , \16559 );
buf \U$59552 ( \59527 , \59024 );
nand \U$59553 ( \59528 , \59526 , \59527 );
buf \U$59554 ( \59529 , \59528 );
buf \U$59555 ( \59530 , \59529 );
nand \U$59556 ( \59531 , \59525 , \59530 );
buf \U$59557 ( \59532 , \59531 );
buf \U$59558 ( \59533 , \59532 );
buf \U$59559 ( \59534 , RIc0d9388_63);
buf \U$59560 ( \59535 , RIc0daa08_111);
xor \U$59561 ( \59536 , \59534 , \59535 );
buf \U$59562 ( \59537 , \59536 );
buf \U$59563 ( \59538 , \59537 );
not \U$59564 ( \59539 , \59538 );
buf \U$59565 ( \59540 , \12529 );
not \U$59566 ( \59541 , \59540 );
or \U$59567 ( \59542 , \59539 , \59541 );
buf \U$59568 ( \59543 , \25649 );
buf \U$59569 ( \59544 , \59315 );
nand \U$59570 ( \59545 , \59543 , \59544 );
buf \U$59571 ( \59546 , \59545 );
buf \U$59572 ( \59547 , \59546 );
nand \U$59573 ( \59548 , \59542 , \59547 );
buf \U$59574 ( \59549 , \59548 );
buf \U$59575 ( \59550 , \59549 );
or \U$59576 ( \59551 , \59533 , \59550 );
buf \U$59577 ( \59552 , RIc0d91a8_59);
buf \U$59578 ( \59553 , RIc0dabe8_115);
xor \U$59579 ( \59554 , \59552 , \59553 );
buf \U$59580 ( \59555 , \59554 );
buf \U$59581 ( \59556 , \59555 );
not \U$59582 ( \59557 , \59556 );
buf \U$59583 ( \59558 , \46873 );
not \U$59584 ( \59559 , \59558 );
or \U$59585 ( \59560 , \59557 , \59559 );
buf \U$59586 ( \59561 , \12303 );
buf \U$59587 ( \59562 , \58904 );
nand \U$59588 ( \59563 , \59561 , \59562 );
buf \U$59589 ( \59564 , \59563 );
buf \U$59590 ( \59565 , \59564 );
nand \U$59591 ( \59566 , \59560 , \59565 );
buf \U$59592 ( \59567 , \59566 );
buf \U$59593 ( \59568 , \59567 );
nand \U$59594 ( \59569 , \59551 , \59568 );
buf \U$59595 ( \59570 , \59569 );
buf \U$59596 ( \59571 , \59570 );
buf \U$59597 ( \59572 , \59532 );
buf \U$59598 ( \59573 , \59549 );
nand \U$59599 ( \59574 , \59572 , \59573 );
buf \U$59600 ( \59575 , \59574 );
buf \U$59601 ( \59576 , \59575 );
nand \U$59602 ( \59577 , \59571 , \59576 );
buf \U$59603 ( \59578 , \59577 );
buf \U$59604 ( \59579 , \59578 );
xor \U$59605 ( \59580 , \59516 , \59579 );
buf \U$59606 ( \59581 , RIc0db200_128);
not \U$59607 ( \59582 , \59581 );
buf \U$59608 ( \59583 , \58979 );
not \U$59609 ( \59584 , \59583 );
or \U$59610 ( \59585 , \59582 , \59584 );
buf \U$59611 ( \59586 , \58200 );
buf \U$59612 ( \59587 , RIc0db188_127);
buf \U$59613 ( \59588 , RIc0d8c08_47);
xnor \U$59614 ( \59589 , \59587 , \59588 );
buf \U$59615 ( \59590 , \59589 );
buf \U$59616 ( \59591 , \59590 );
or \U$59617 ( \59592 , \59586 , \59591 );
nand \U$59618 ( \59593 , \59585 , \59592 );
buf \U$59619 ( \59594 , \59593 );
buf \U$59620 ( \59595 , \59594 );
buf \U$59621 ( \59596 , RIc0d8fc8_55);
buf \U$59622 ( \59597 , RIc0dadc8_119);
xor \U$59623 ( \59598 , \59596 , \59597 );
buf \U$59624 ( \59599 , \59598 );
buf \U$59625 ( \59600 , \59599 );
not \U$59626 ( \59601 , \59600 );
buf \U$59627 ( \59602 , \13949 );
not \U$59628 ( \59603 , \59602 );
or \U$59629 ( \59604 , \59601 , \59603 );
buf \U$59630 ( \59605 , \59092 );
not \U$59631 ( \59606 , \59605 );
buf \U$59632 ( \59607 , \13005 );
nand \U$59633 ( \59608 , \59606 , \59607 );
buf \U$59634 ( \59609 , \59608 );
buf \U$59635 ( \59610 , \59609 );
nand \U$59636 ( \59611 , \59604 , \59610 );
buf \U$59637 ( \59612 , \59611 );
buf \U$59638 ( \59613 , \59612 );
xor \U$59639 ( \59614 , \59595 , \59613 );
buf \U$59640 ( \59615 , \17992 );
buf \U$59641 ( \59616 , RIc0db098_125);
buf \U$59642 ( \59617 , \22504 );
and \U$59643 ( \59618 , \59616 , \59617 );
not \U$59644 ( \59619 , \59616 );
buf \U$59645 ( \59620 , RIc0d8cf8_49);
and \U$59646 ( \59621 , \59619 , \59620 );
nor \U$59647 ( \59622 , \59618 , \59621 );
buf \U$59648 ( \59623 , \59622 );
buf \U$59649 ( \59624 , \59623 );
or \U$59650 ( \59625 , \59615 , \59624 );
buf \U$59651 ( \59626 , \22744 );
buf \U$59652 ( \59627 , \59054 );
not \U$59653 ( \59628 , \59627 );
buf \U$59654 ( \59629 , \59628 );
buf \U$59655 ( \59630 , \59629 );
or \U$59656 ( \59631 , \59626 , \59630 );
nand \U$59657 ( \59632 , \59625 , \59631 );
buf \U$59658 ( \59633 , \59632 );
buf \U$59659 ( \59634 , \59633 );
and \U$59660 ( \59635 , \59614 , \59634 );
and \U$59661 ( \59636 , \59595 , \59613 );
or \U$59662 ( \59637 , \59635 , \59636 );
buf \U$59663 ( \59638 , \59637 );
buf \U$59664 ( \59639 , \59638 );
and \U$59665 ( \59640 , \59580 , \59639 );
and \U$59666 ( \59641 , \59516 , \59579 );
or \U$59667 ( \59642 , \59640 , \59641 );
buf \U$59668 ( \59643 , \59642 );
buf \U$59669 ( \59644 , \59643 );
xor \U$59670 ( \59645 , \59505 , \59644 );
buf \U$59671 ( \59646 , \15909 );
buf \U$59672 ( \59647 , RIc0d9400_64);
and \U$59673 ( \59648 , \59646 , \59647 );
buf \U$59674 ( \59649 , \59648 );
buf \U$59675 ( \59650 , \59649 );
buf \U$59676 ( \59651 , RIc0d9298_61);
buf \U$59677 ( \59652 , RIc0daaf8_113);
xor \U$59678 ( \59653 , \59651 , \59652 );
buf \U$59679 ( \59654 , \59653 );
buf \U$59680 ( \59655 , \59654 );
not \U$59681 ( \59656 , \59655 );
buf \U$59682 ( \59657 , \33224 );
not \U$59683 ( \59658 , \59657 );
or \U$59684 ( \59659 , \59656 , \59658 );
buf \U$59685 ( \59660 , \14405 );
buf \U$59686 ( \59661 , \59001 );
nand \U$59687 ( \59662 , \59660 , \59661 );
buf \U$59688 ( \59663 , \59662 );
buf \U$59689 ( \59664 , \59663 );
nand \U$59690 ( \59665 , \59659 , \59664 );
buf \U$59691 ( \59666 , \59665 );
buf \U$59692 ( \59667 , \59666 );
xor \U$59693 ( \59668 , \59650 , \59667 );
buf \U$59694 ( \59669 , \59072 );
not \U$59695 ( \59670 , \59669 );
buf \U$59696 ( \59671 , \16692 );
not \U$59697 ( \59672 , \59671 );
or \U$59698 ( \59673 , \59670 , \59672 );
buf \U$59699 ( \59674 , \45089 );
buf \U$59700 ( \59675 , RIc0d8de8_51);
buf \U$59701 ( \59676 , RIc0dafa8_123);
xnor \U$59702 ( \59677 , \59675 , \59676 );
buf \U$59703 ( \59678 , \59677 );
buf \U$59704 ( \59679 , \59678 );
or \U$59705 ( \59680 , \59674 , \59679 );
nand \U$59706 ( \59681 , \59673 , \59680 );
buf \U$59707 ( \59682 , \59681 );
buf \U$59708 ( \59683 , \59682 );
and \U$59709 ( \59684 , \59668 , \59683 );
and \U$59710 ( \59685 , \59650 , \59667 );
or \U$59711 ( \59686 , \59684 , \59685 );
buf \U$59712 ( \59687 , \59686 );
buf \U$59713 ( \59688 , \59687 );
xor \U$59714 ( \59689 , \59068 , \59086 );
xor \U$59715 ( \59690 , \59689 , \59107 );
buf \U$59716 ( \59691 , \59690 );
buf \U$59717 ( \59692 , \59691 );
xor \U$59718 ( \59693 , \59688 , \59692 );
xor \U$59719 ( \59694 , \58946 , \58970 );
xnor \U$59720 ( \59695 , \59694 , \58920 );
buf \U$59721 ( \59696 , \59695 );
and \U$59722 ( \59697 , \59693 , \59696 );
and \U$59723 ( \59698 , \59688 , \59692 );
or \U$59724 ( \59699 , \59697 , \59698 );
buf \U$59725 ( \59700 , \59699 );
buf \U$59726 ( \59701 , \59700 );
and \U$59727 ( \59702 , \59645 , \59701 );
and \U$59728 ( \59703 , \59505 , \59644 );
or \U$59729 ( \59704 , \59702 , \59703 );
buf \U$59730 ( \59705 , \59704 );
buf \U$59731 ( \59706 , \59705 );
not \U$59732 ( \59707 , \59706 );
xor \U$59733 ( \59708 , \59434 , \59438 );
xor \U$59734 ( \59709 , \59708 , \59458 );
buf \U$59735 ( \59710 , \59709 );
buf \U$59736 ( \59711 , \59710 );
buf \U$59737 ( \59712 , \58976 );
buf \U$59738 ( \59713 , \59046 );
xor \U$59739 ( \59714 , \59712 , \59713 );
buf \U$59740 ( \59715 , \59111 );
xor \U$59741 ( \59716 , \59714 , \59715 );
buf \U$59742 ( \59717 , \59716 );
buf \U$59743 ( \59718 , \59717 );
xor \U$59744 ( \59719 , \59711 , \59718 );
xor \U$59745 ( \59720 , \59505 , \59644 );
xor \U$59746 ( \59721 , \59720 , \59701 );
buf \U$59747 ( \59722 , \59721 );
buf \U$59748 ( \59723 , \59722 );
and \U$59749 ( \59724 , \59719 , \59723 );
and \U$59750 ( \59725 , \59711 , \59718 );
or \U$59751 ( \59726 , \59724 , \59725 );
buf \U$59752 ( \59727 , \59726 );
buf \U$59753 ( \59728 , \59727 );
not \U$59754 ( \59729 , \59728 );
or \U$59755 ( \59730 , \59707 , \59729 );
buf \U$59756 ( \59731 , \59727 );
buf \U$59757 ( \59732 , \59705 );
or \U$59758 ( \59733 , \59731 , \59732 );
xor \U$59759 ( \59734 , \59463 , \59467 );
xor \U$59760 ( \59735 , \59734 , \59489 );
buf \U$59761 ( \59736 , \59735 );
buf \U$59762 ( \59737 , \59736 );
nand \U$59763 ( \59738 , \59733 , \59737 );
buf \U$59764 ( \59739 , \59738 );
buf \U$59765 ( \59740 , \59739 );
nand \U$59766 ( \59741 , \59730 , \59740 );
buf \U$59767 ( \59742 , \59741 );
buf \U$59768 ( \59743 , \59742 );
or \U$59769 ( \59744 , \59502 , \59743 );
buf \U$59770 ( \59745 , \59744 );
buf \U$59771 ( \59746 , \59745 );
not \U$59772 ( \59747 , \59746 );
buf \U$59773 ( \59748 , \59040 );
not \U$59774 ( \59749 , \59748 );
buf \U$59775 ( \59750 , \59017 );
buf \U$59776 ( \59751 , \58995 );
xnor \U$59777 ( \59752 , \59750 , \59751 );
buf \U$59778 ( \59753 , \59752 );
buf \U$59779 ( \59754 , \59753 );
not \U$59780 ( \59755 , \59754 );
or \U$59781 ( \59756 , \59749 , \59755 );
buf \U$59782 ( \59757 , \59753 );
buf \U$59783 ( \59758 , \59040 );
or \U$59784 ( \59759 , \59757 , \59758 );
nand \U$59785 ( \59760 , \59756 , \59759 );
buf \U$59786 ( \59761 , \59760 );
buf \U$59787 ( \59762 , \59761 );
buf \U$59788 ( \59763 , \49672 );
buf \U$59789 ( \59764 , \13166 );
buf \U$59790 ( \59765 , RIc0d8ed8_53);
and \U$59791 ( \59766 , \59764 , \59765 );
buf \U$59792 ( \59767 , \23372 );
buf \U$59793 ( \59768 , RIc0daeb8_121);
and \U$59794 ( \59769 , \59767 , \59768 );
nor \U$59795 ( \59770 , \59766 , \59769 );
buf \U$59796 ( \59771 , \59770 );
buf \U$59797 ( \59772 , \59771 );
or \U$59798 ( \59773 , \59763 , \59772 );
buf \U$59799 ( \59774 , \26373 );
buf \U$59800 ( \59775 , \58926 );
not \U$59801 ( \59776 , \59775 );
buf \U$59802 ( \59777 , \59776 );
buf \U$59803 ( \59778 , \59777 );
or \U$59804 ( \59779 , \59774 , \59778 );
nand \U$59805 ( \59780 , \59773 , \59779 );
buf \U$59806 ( \59781 , \59780 );
buf \U$59807 ( \59782 , \59781 );
buf \U$59808 ( \59783 , RIc0d9400_64);
buf \U$59809 ( \59784 , RIc0daa80_112);
or \U$59810 ( \59785 , \59783 , \59784 );
buf \U$59811 ( \59786 , RIc0daaf8_113);
nand \U$59812 ( \59787 , \59785 , \59786 );
buf \U$59813 ( \59788 , \59787 );
buf \U$59814 ( \59789 , \59788 );
buf \U$59815 ( \59790 , RIc0d9400_64);
buf \U$59816 ( \59791 , RIc0daa80_112);
nand \U$59817 ( \59792 , \59790 , \59791 );
buf \U$59818 ( \59793 , \59792 );
buf \U$59819 ( \59794 , \59793 );
buf \U$59820 ( \59795 , RIc0daa08_111);
and \U$59821 ( \59796 , \59789 , \59794 , \59795 );
buf \U$59822 ( \59797 , \59796 );
buf \U$59823 ( \59798 , \59797 );
buf \U$59824 ( \59799 , \16989 );
not \U$59825 ( \59800 , \59799 );
buf \U$59826 ( \59801 , \59800 );
buf \U$59827 ( \59802 , \59801 );
buf \U$59828 ( \59803 , RIc0d9310_62);
buf \U$59829 ( \59804 , RIc0daaf8_113);
xnor \U$59830 ( \59805 , \59803 , \59804 );
buf \U$59831 ( \59806 , \59805 );
buf \U$59832 ( \59807 , \59806 );
or \U$59833 ( \59808 , \59802 , \59807 );
buf \U$59834 ( \59809 , \34244 );
buf \U$59835 ( \59810 , \59654 );
not \U$59836 ( \59811 , \59810 );
buf \U$59837 ( \59812 , \59811 );
buf \U$59838 ( \59813 , \59812 );
or \U$59839 ( \59814 , \59809 , \59813 );
nand \U$59840 ( \59815 , \59808 , \59814 );
buf \U$59841 ( \59816 , \59815 );
buf \U$59842 ( \59817 , \59816 );
and \U$59843 ( \59818 , \59798 , \59817 );
buf \U$59844 ( \59819 , \59818 );
buf \U$59845 ( \59820 , \59819 );
xor \U$59846 ( \59821 , \59782 , \59820 );
buf \U$59847 ( \59822 , RIc0d9130_58);
buf \U$59848 ( \59823 , RIc0dacd8_117);
xor \U$59849 ( \59824 , \59822 , \59823 );
buf \U$59850 ( \59825 , \59824 );
buf \U$59851 ( \59826 , \59825 );
not \U$59852 ( \59827 , \59826 );
buf \U$59853 ( \59828 , \13146 );
not \U$59854 ( \59829 , \59828 );
or \U$59855 ( \59830 , \59827 , \59829 );
buf \U$59856 ( \59831 , \22356 );
buf \U$59857 ( \59832 , \59520 );
nand \U$59858 ( \59833 , \59831 , \59832 );
buf \U$59859 ( \59834 , \59833 );
buf \U$59860 ( \59835 , \59834 );
nand \U$59861 ( \59836 , \59830 , \59835 );
buf \U$59862 ( \59837 , \59836 );
buf \U$59863 ( \59838 , \59837 );
buf \U$59864 ( \59839 , RIc0daa08_111);
buf \U$59865 ( \59840 , RIc0d9400_64);
and \U$59866 ( \59841 , \59839 , \59840 );
not \U$59867 ( \59842 , \59839 );
buf \U$59868 ( \59843 , \43843 );
and \U$59869 ( \59844 , \59842 , \59843 );
nor \U$59870 ( \59845 , \59841 , \59844 );
buf \U$59871 ( \59846 , \59845 );
buf \U$59872 ( \59847 , \59846 );
not \U$59873 ( \59848 , \59847 );
buf \U$59874 ( \59849 , \18306 );
not \U$59875 ( \59850 , \59849 );
or \U$59876 ( \59851 , \59848 , \59850 );
buf \U$59877 ( \59852 , \45728 );
buf \U$59878 ( \59853 , \59537 );
nand \U$59879 ( \59854 , \59852 , \59853 );
buf \U$59880 ( \59855 , \59854 );
buf \U$59881 ( \59856 , \59855 );
nand \U$59882 ( \59857 , \59851 , \59856 );
buf \U$59883 ( \59858 , \59857 );
buf \U$59884 ( \59859 , \59858 );
xor \U$59885 ( \59860 , \59838 , \59859 );
buf \U$59886 ( \59861 , \16688 );
buf \U$59887 ( \59862 , RIc0d8e60_52);
buf \U$59888 ( \59863 , RIc0dafa8_123);
xnor \U$59889 ( \59864 , \59862 , \59863 );
buf \U$59890 ( \59865 , \59864 );
buf \U$59891 ( \59866 , \59865 );
or \U$59892 ( \59867 , \59861 , \59866 );
buf \U$59893 ( \59868 , \16695 );
buf \U$59894 ( \59869 , \59678 );
or \U$59895 ( \59870 , \59868 , \59869 );
nand \U$59896 ( \59871 , \59867 , \59870 );
buf \U$59897 ( \59872 , \59871 );
buf \U$59898 ( \59873 , \59872 );
and \U$59899 ( \59874 , \59860 , \59873 );
and \U$59900 ( \59875 , \59838 , \59859 );
or \U$59901 ( \59876 , \59874 , \59875 );
buf \U$59902 ( \59877 , \59876 );
buf \U$59903 ( \59878 , \59877 );
and \U$59904 ( \59879 , \59821 , \59878 );
and \U$59905 ( \59880 , \59782 , \59820 );
or \U$59906 ( \59881 , \59879 , \59880 );
buf \U$59907 ( \59882 , \59881 );
buf \U$59908 ( \59883 , \59882 );
xor \U$59909 ( \59884 , \59762 , \59883 );
xor \U$59910 ( \59885 , \59516 , \59579 );
xor \U$59911 ( \59886 , \59885 , \59639 );
buf \U$59912 ( \59887 , \59886 );
buf \U$59913 ( \59888 , \59887 );
and \U$59914 ( \59889 , \59884 , \59888 );
and \U$59915 ( \59890 , \59762 , \59883 );
or \U$59916 ( \59891 , \59889 , \59890 );
buf \U$59917 ( \59892 , \59891 );
buf \U$59918 ( \59893 , \59892 );
buf \U$59919 ( \59894 , \58200 );
buf \U$59920 ( \59895 , RIc0db188_127);
buf \U$59921 ( \59896 , RIc0d8c80_48);
xnor \U$59922 ( \59897 , \59895 , \59896 );
buf \U$59923 ( \59898 , \59897 );
buf \U$59924 ( \59899 , \59898 );
or \U$59925 ( \59900 , \59894 , \59899 );
buf \U$59926 ( \59901 , \12647 );
buf \U$59927 ( \59902 , \59590 );
or \U$59928 ( \59903 , \59901 , \59902 );
nand \U$59929 ( \59904 , \59900 , \59903 );
buf \U$59930 ( \59905 , \59904 );
buf \U$59931 ( \59906 , \59905 );
buf \U$59932 ( \59907 , RIc0d9220_60);
buf \U$59933 ( \59908 , RIc0dabe8_115);
xor \U$59934 ( \59909 , \59907 , \59908 );
buf \U$59935 ( \59910 , \59909 );
buf \U$59936 ( \59911 , \59910 );
not \U$59937 ( \59912 , \59911 );
buf \U$59938 ( \59913 , \26466 );
not \U$59939 ( \59914 , \59913 );
or \U$59940 ( \59915 , \59912 , \59914 );
buf \U$59941 ( \59916 , \12303 );
buf \U$59942 ( \59917 , \59555 );
nand \U$59943 ( \59918 , \59916 , \59917 );
buf \U$59944 ( \59919 , \59918 );
buf \U$59945 ( \59920 , \59919 );
nand \U$59946 ( \59921 , \59915 , \59920 );
buf \U$59947 ( \59922 , \59921 );
buf \U$59948 ( \59923 , \59922 );
xor \U$59949 ( \59924 , \59906 , \59923 );
buf \U$59950 ( \59925 , \13178 );
buf \U$59951 ( \59926 , RIc0dadc8_119);
buf \U$59952 ( \59927 , RIc0d9040_56);
xnor \U$59953 ( \59928 , \59926 , \59927 );
buf \U$59954 ( \59929 , \59928 );
buf \U$59955 ( \59930 , \59929 );
or \U$59956 ( \59931 , \59925 , \59930 );
buf \U$59957 ( \59932 , \45225 );
buf \U$59958 ( \59933 , \59599 );
not \U$59959 ( \59934 , \59933 );
buf \U$59960 ( \59935 , \59934 );
buf \U$59961 ( \59936 , \59935 );
or \U$59962 ( \59937 , \59932 , \59936 );
nand \U$59963 ( \59938 , \59931 , \59937 );
buf \U$59964 ( \59939 , \59938 );
buf \U$59965 ( \59940 , \59939 );
and \U$59966 ( \59941 , \59924 , \59940 );
and \U$59967 ( \59942 , \59906 , \59923 );
or \U$59968 ( \59943 , \59941 , \59942 );
buf \U$59969 ( \59944 , \59943 );
buf \U$59970 ( \59945 , \59944 );
xor \U$59971 ( \59946 , \59595 , \59613 );
xor \U$59972 ( \59947 , \59946 , \59634 );
buf \U$59973 ( \59948 , \59947 );
buf \U$59974 ( \59949 , \59948 );
xor \U$59975 ( \59950 , \59945 , \59949 );
xor \U$59976 ( \59951 , \59650 , \59667 );
xor \U$59977 ( \59952 , \59951 , \59683 );
buf \U$59978 ( \59953 , \59952 );
buf \U$59979 ( \59954 , \59953 );
and \U$59980 ( \59955 , \59950 , \59954 );
and \U$59981 ( \59956 , \59945 , \59949 );
or \U$59982 ( \59957 , \59955 , \59956 );
buf \U$59983 ( \59958 , \59957 );
buf \U$59984 ( \59959 , \59958 );
xor \U$59985 ( \59960 , \59688 , \59692 );
xor \U$59986 ( \59961 , \59960 , \59696 );
buf \U$59987 ( \59962 , \59961 );
buf \U$59988 ( \59963 , \59962 );
xor \U$59989 ( \59964 , \59959 , \59963 );
xor \U$59990 ( \59965 , \59532 , \59549 );
xor \U$59991 ( \59966 , \59567 , \59965 );
buf \U$59992 ( \59967 , \59966 );
buf \U$59993 ( \59968 , \12968 );
buf \U$59994 ( \59969 , RIc0d8f50_54);
buf \U$59995 ( \59970 , RIc0daeb8_121);
xnor \U$59996 ( \59971 , \59969 , \59970 );
buf \U$59997 ( \59972 , \59971 );
buf \U$59998 ( \59973 , \59972 );
or \U$59999 ( \59974 , \59968 , \59973 );
buf \U$60000 ( \59975 , \26373 );
buf \U$60001 ( \59976 , \59771 );
or \U$60002 ( \59977 , \59975 , \59976 );
nand \U$60003 ( \59978 , \59974 , \59977 );
buf \U$60004 ( \59979 , \59978 );
buf \U$60005 ( \59980 , \59979 );
buf \U$60006 ( \59981 , \14468 );
buf \U$60007 ( \59982 , RIc0d8d70_50);
buf \U$60008 ( \59983 , RIc0db098_125);
xnor \U$60009 ( \59984 , \59982 , \59983 );
buf \U$60010 ( \59985 , \59984 );
buf \U$60011 ( \59986 , \59985 );
or \U$60012 ( \59987 , \59981 , \59986 );
buf \U$60013 ( \59988 , \22744 );
buf \U$60014 ( \59989 , \59623 );
or \U$60015 ( \59990 , \59988 , \59989 );
nand \U$60016 ( \59991 , \59987 , \59990 );
buf \U$60017 ( \59992 , \59991 );
buf \U$60018 ( \59993 , \59992 );
xor \U$60019 ( \59994 , \59980 , \59993 );
xor \U$60020 ( \59995 , \59798 , \59817 );
buf \U$60021 ( \59996 , \59995 );
buf \U$60022 ( \59997 , \59996 );
and \U$60023 ( \59998 , \59994 , \59997 );
and \U$60024 ( \59999 , \59980 , \59993 );
or \U$60025 ( \60000 , \59998 , \59999 );
buf \U$60026 ( \60001 , \60000 );
buf \U$60027 ( \60002 , \60001 );
xor \U$60028 ( \60003 , \59967 , \60002 );
xor \U$60029 ( \60004 , \59782 , \59820 );
xor \U$60030 ( \60005 , \60004 , \59878 );
buf \U$60031 ( \60006 , \60005 );
buf \U$60032 ( \60007 , \60006 );
and \U$60033 ( \60008 , \60003 , \60007 );
and \U$60034 ( \60009 , \59967 , \60002 );
or \U$60035 ( \60010 , \60008 , \60009 );
buf \U$60036 ( \60011 , \60010 );
buf \U$60037 ( \60012 , \60011 );
and \U$60038 ( \60013 , \59964 , \60012 );
and \U$60039 ( \60014 , \59959 , \59963 );
or \U$60040 ( \60015 , \60013 , \60014 );
buf \U$60041 ( \60016 , \60015 );
buf \U$60042 ( \60017 , \60016 );
xor \U$60043 ( \60018 , \59893 , \60017 );
xor \U$60044 ( \60019 , \59711 , \59718 );
xor \U$60045 ( \60020 , \60019 , \59723 );
buf \U$60046 ( \60021 , \60020 );
buf \U$60047 ( \60022 , \60021 );
xor \U$60048 ( \60023 , \60018 , \60022 );
buf \U$60049 ( \60024 , \60023 );
buf \U$60050 ( \60025 , \60024 );
xor \U$60051 ( \60026 , \59762 , \59883 );
xor \U$60052 ( \60027 , \60026 , \59888 );
buf \U$60053 ( \60028 , \60027 );
buf \U$60054 ( \60029 , \60028 );
not \U$60055 ( \60030 , \60029 );
buf \U$60056 ( \60031 , RIc0daaf8_113);
buf \U$60057 ( \60032 , RIc0d9388_63);
and \U$60058 ( \60033 , \60031 , \60032 );
not \U$60059 ( \60034 , \60031 );
buf \U$60060 ( \60035 , \43939 );
and \U$60061 ( \60036 , \60034 , \60035 );
nor \U$60062 ( \60037 , \60033 , \60036 );
buf \U$60063 ( \60038 , \60037 );
buf \U$60064 ( \60039 , \60038 );
not \U$60065 ( \60040 , \60039 );
buf \U$60066 ( \60041 , \25355 );
not \U$60067 ( \60042 , \60041 );
or \U$60068 ( \60043 , \60040 , \60042 );
buf \U$60069 ( \60044 , \59806 );
not \U$60070 ( \60045 , \60044 );
buf \U$60071 ( \60046 , \12410 );
nand \U$60072 ( \60047 , \60045 , \60046 );
buf \U$60073 ( \60048 , \60047 );
buf \U$60074 ( \60049 , \60048 );
nand \U$60075 ( \60050 , \60043 , \60049 );
buf \U$60076 ( \60051 , \60050 );
buf \U$60077 ( \60052 , \60051 );
buf \U$60078 ( \60053 , RIc0d8ed8_53);
buf \U$60079 ( \60054 , RIc0dafa8_123);
xor \U$60080 ( \60055 , \60053 , \60054 );
buf \U$60081 ( \60056 , \60055 );
buf \U$60082 ( \60057 , \60056 );
not \U$60083 ( \60058 , \60057 );
buf \U$60084 ( \60059 , \45570 );
not \U$60085 ( \60060 , \60059 );
or \U$60086 ( \60061 , \60058 , \60060 );
buf \U$60087 ( \60062 , \59865 );
not \U$60088 ( \60063 , \60062 );
buf \U$60089 ( \60064 , \16692 );
nand \U$60090 ( \60065 , \60063 , \60064 );
buf \U$60091 ( \60066 , \60065 );
buf \U$60092 ( \60067 , \60066 );
nand \U$60093 ( \60068 , \60061 , \60067 );
buf \U$60094 ( \60069 , \60068 );
buf \U$60095 ( \60070 , \60069 );
nor \U$60096 ( \60071 , \60052 , \60070 );
buf \U$60097 ( \60072 , \60071 );
buf \U$60098 ( \60073 , \60072 );
buf \U$60099 ( \60074 , RIc0d8fc8_55);
buf \U$60100 ( \60075 , RIc0daeb8_121);
xor \U$60101 ( \60076 , \60074 , \60075 );
buf \U$60102 ( \60077 , \60076 );
buf \U$60103 ( \60078 , \60077 );
not \U$60104 ( \60079 , \60078 );
buf \U$60105 ( \60080 , \24672 );
not \U$60106 ( \60081 , \60080 );
or \U$60107 ( \60082 , \60079 , \60081 );
buf \U$60108 ( \60083 , \59972 );
not \U$60109 ( \60084 , \60083 );
buf \U$60110 ( \60085 , \16386 );
nand \U$60111 ( \60086 , \60084 , \60085 );
buf \U$60112 ( \60087 , \60086 );
buf \U$60113 ( \60088 , \60087 );
nand \U$60114 ( \60089 , \60082 , \60088 );
buf \U$60115 ( \60090 , \60089 );
buf \U$60116 ( \60091 , \60090 );
not \U$60117 ( \60092 , \60091 );
buf \U$60118 ( \60093 , \60092 );
buf \U$60119 ( \60094 , \60093 );
or \U$60120 ( \60095 , \60073 , \60094 );
buf \U$60121 ( \60096 , \60051 );
buf \U$60122 ( \60097 , \60069 );
nand \U$60123 ( \60098 , \60096 , \60097 );
buf \U$60124 ( \60099 , \60098 );
buf \U$60125 ( \60100 , \60099 );
nand \U$60126 ( \60101 , \60095 , \60100 );
buf \U$60127 ( \60102 , \60101 );
buf \U$60128 ( \60103 , \60102 );
buf \U$60129 ( \60104 , \14106 );
buf \U$60130 ( \60105 , RIc0d9400_64);
and \U$60131 ( \60106 , \60104 , \60105 );
buf \U$60132 ( \60107 , \60106 );
buf \U$60133 ( \60108 , \60107 );
buf \U$60134 ( \60109 , RIc0d9298_61);
buf \U$60135 ( \60110 , RIc0dabe8_115);
xor \U$60136 ( \60111 , \60109 , \60110 );
buf \U$60137 ( \60112 , \60111 );
buf \U$60138 ( \60113 , \60112 );
not \U$60139 ( \60114 , \60113 );
buf \U$60140 ( \60115 , \26466 );
not \U$60141 ( \60116 , \60115 );
or \U$60142 ( \60117 , \60114 , \60116 );
buf \U$60143 ( \60118 , \12303 );
buf \U$60144 ( \60119 , \59910 );
nand \U$60145 ( \60120 , \60118 , \60119 );
buf \U$60146 ( \60121 , \60120 );
buf \U$60147 ( \60122 , \60121 );
nand \U$60148 ( \60123 , \60117 , \60122 );
buf \U$60149 ( \60124 , \60123 );
buf \U$60150 ( \60125 , \60124 );
xor \U$60151 ( \60126 , \60108 , \60125 );
buf \U$60152 ( \60127 , RIc0d8de8_51);
buf \U$60153 ( \60128 , RIc0db098_125);
xor \U$60154 ( \60129 , \60127 , \60128 );
buf \U$60155 ( \60130 , \60129 );
buf \U$60156 ( \60131 , \60130 );
not \U$60157 ( \60132 , \60131 );
buf \U$60158 ( \60133 , \14471 );
not \U$60159 ( \60134 , \60133 );
or \U$60160 ( \60135 , \60132 , \60134 );
buf \U$60161 ( \60136 , \59985 );
not \U$60162 ( \60137 , \60136 );
buf \U$60163 ( \60138 , \15793 );
nand \U$60164 ( \60139 , \60137 , \60138 );
buf \U$60165 ( \60140 , \60139 );
buf \U$60166 ( \60141 , \60140 );
nand \U$60167 ( \60142 , \60135 , \60141 );
buf \U$60168 ( \60143 , \60142 );
buf \U$60169 ( \60144 , \60143 );
and \U$60170 ( \60145 , \60126 , \60144 );
and \U$60171 ( \60146 , \60108 , \60125 );
or \U$60172 ( \60147 , \60145 , \60146 );
buf \U$60173 ( \60148 , \60147 );
buf \U$60174 ( \60149 , \60148 );
or \U$60175 ( \60150 , \60103 , \60149 );
not \U$60176 ( \60151 , \15609 );
buf \U$60177 ( \60152 , \60151 );
buf \U$60178 ( \60153 , RIc0db188_127);
buf \U$60179 ( \60154 , RIc0d8cf8_49);
xor \U$60180 ( \60155 , \60153 , \60154 );
buf \U$60181 ( \60156 , \60155 );
buf \U$60182 ( \60157 , \60156 );
not \U$60183 ( \60158 , \60157 );
buf \U$60184 ( \60159 , \60158 );
buf \U$60185 ( \60160 , \60159 );
or \U$60186 ( \60161 , \60152 , \60160 );
buf \U$60187 ( \60162 , \12647 );
buf \U$60188 ( \60163 , \59898 );
or \U$60189 ( \60164 , \60162 , \60163 );
nand \U$60190 ( \60165 , \60161 , \60164 );
buf \U$60191 ( \60166 , \60165 );
buf \U$60192 ( \60167 , \60166 );
buf \U$60193 ( \60168 , RIc0d90b8_57);
buf \U$60194 ( \60169 , RIc0dadc8_119);
xor \U$60195 ( \60170 , \60168 , \60169 );
buf \U$60196 ( \60171 , \60170 );
buf \U$60197 ( \60172 , \60171 );
not \U$60198 ( \60173 , \60172 );
buf \U$60199 ( \60174 , \14569 );
not \U$60200 ( \60175 , \60174 );
or \U$60201 ( \60176 , \60173 , \60175 );
buf \U$60202 ( \60177 , \59929 );
not \U$60203 ( \60178 , \60177 );
buf \U$60204 ( \60179 , \13005 );
nand \U$60205 ( \60180 , \60178 , \60179 );
buf \U$60206 ( \60181 , \60180 );
buf \U$60207 ( \60182 , \60181 );
nand \U$60208 ( \60183 , \60176 , \60182 );
buf \U$60209 ( \60184 , \60183 );
buf \U$60210 ( \60185 , \60184 );
xor \U$60211 ( \60186 , \60167 , \60185 );
buf \U$60212 ( \60187 , RIc0d91a8_59);
buf \U$60213 ( \60188 , RIc0dacd8_117);
xor \U$60214 ( \60189 , \60187 , \60188 );
buf \U$60215 ( \60190 , \60189 );
buf \U$60216 ( \60191 , \60190 );
not \U$60217 ( \60192 , \60191 );
buf \U$60218 ( \60193 , \12929 );
not \U$60219 ( \60194 , \60193 );
or \U$60220 ( \60195 , \60192 , \60194 );
buf \U$60221 ( \60196 , \12937 );
buf \U$60222 ( \60197 , \59825 );
nand \U$60223 ( \60198 , \60196 , \60197 );
buf \U$60224 ( \60199 , \60198 );
buf \U$60225 ( \60200 , \60199 );
nand \U$60226 ( \60201 , \60195 , \60200 );
buf \U$60227 ( \60202 , \60201 );
buf \U$60228 ( \60203 , \60202 );
and \U$60229 ( \60204 , \60186 , \60203 );
and \U$60230 ( \60205 , \60167 , \60185 );
or \U$60231 ( \60206 , \60204 , \60205 );
buf \U$60232 ( \60207 , \60206 );
buf \U$60233 ( \60208 , \60207 );
nand \U$60234 ( \60209 , \60150 , \60208 );
buf \U$60235 ( \60210 , \60209 );
buf \U$60236 ( \60211 , \60210 );
buf \U$60237 ( \60212 , \60102 );
buf \U$60238 ( \60213 , \60148 );
nand \U$60239 ( \60214 , \60212 , \60213 );
buf \U$60240 ( \60215 , \60214 );
buf \U$60241 ( \60216 , \60215 );
nand \U$60242 ( \60217 , \60211 , \60216 );
buf \U$60243 ( \60218 , \60217 );
buf \U$60244 ( \60219 , \60218 );
xor \U$60245 ( \60220 , \59945 , \59949 );
xor \U$60246 ( \60221 , \60220 , \59954 );
buf \U$60247 ( \60222 , \60221 );
buf \U$60248 ( \60223 , \60222 );
xor \U$60249 ( \60224 , \60219 , \60223 );
xor \U$60250 ( \60225 , \59906 , \59923 );
xor \U$60251 ( \60226 , \60225 , \59940 );
buf \U$60252 ( \60227 , \60226 );
buf \U$60253 ( \60228 , \60227 );
xor \U$60254 ( \60229 , \59838 , \59859 );
xor \U$60255 ( \60230 , \60229 , \59873 );
buf \U$60256 ( \60231 , \60230 );
buf \U$60257 ( \60232 , \60231 );
xor \U$60258 ( \60233 , \60228 , \60232 );
xor \U$60259 ( \60234 , \59980 , \59993 );
xor \U$60260 ( \60235 , \60234 , \59997 );
buf \U$60261 ( \60236 , \60235 );
buf \U$60262 ( \60237 , \60236 );
and \U$60263 ( \60238 , \60233 , \60237 );
and \U$60264 ( \60239 , \60228 , \60232 );
or \U$60265 ( \60240 , \60238 , \60239 );
buf \U$60266 ( \60241 , \60240 );
buf \U$60267 ( \60242 , \60241 );
and \U$60268 ( \60243 , \60224 , \60242 );
and \U$60269 ( \60244 , \60219 , \60223 );
or \U$60270 ( \60245 , \60243 , \60244 );
buf \U$60271 ( \60246 , \60245 );
buf \U$60272 ( \60247 , \60246 );
not \U$60273 ( \60248 , \60247 );
or \U$60274 ( \60249 , \60030 , \60248 );
buf \U$60275 ( \60250 , \60246 );
buf \U$60276 ( \60251 , \60028 );
or \U$60277 ( \60252 , \60250 , \60251 );
xor \U$60278 ( \60253 , \59959 , \59963 );
xor \U$60279 ( \60254 , \60253 , \60012 );
buf \U$60280 ( \60255 , \60254 );
buf \U$60281 ( \60256 , \60255 );
nand \U$60282 ( \60257 , \60252 , \60256 );
buf \U$60283 ( \60258 , \60257 );
buf \U$60284 ( \60259 , \60258 );
nand \U$60285 ( \60260 , \60249 , \60259 );
buf \U$60286 ( \60261 , \60260 );
buf \U$60287 ( \60262 , \60261 );
nand \U$60288 ( \60263 , \60025 , \60262 );
buf \U$60289 ( \60264 , \60263 );
buf \U$60290 ( \60265 , \60264 );
not \U$60291 ( \60266 , \60265 );
xor \U$60292 ( \60267 , \59893 , \60017 );
and \U$60293 ( \60268 , \60267 , \60022 );
and \U$60294 ( \60269 , \59893 , \60017 );
or \U$60295 ( \60270 , \60268 , \60269 );
buf \U$60296 ( \60271 , \60270 );
buf \U$60297 ( \60272 , \60271 );
not \U$60298 ( \60273 , \60272 );
buf \U$60299 ( \60274 , \59705 );
buf \U$60300 ( \60275 , \59736 );
xor \U$60301 ( \60276 , \60274 , \60275 );
buf \U$60302 ( \60277 , \59727 );
xnor \U$60303 ( \60278 , \60276 , \60277 );
buf \U$60304 ( \60279 , \60278 );
buf \U$60305 ( \60280 , \60279 );
nand \U$60306 ( \60281 , \60273 , \60280 );
buf \U$60307 ( \60282 , \60281 );
buf \U$60308 ( \60283 , \60282 );
nand \U$60309 ( \60284 , \60266 , \60283 );
buf \U$60310 ( \60285 , \60284 );
buf \U$60311 ( \60286 , \60285 );
buf \U$60312 ( \60287 , \60279 );
not \U$60313 ( \60288 , \60287 );
buf \U$60314 ( \60289 , \60271 );
nand \U$60315 ( \60290 , \60288 , \60289 );
buf \U$60316 ( \60291 , \60290 );
buf \U$60317 ( \60292 , \60291 );
nand \U$60318 ( \60293 , \60286 , \60292 );
buf \U$60319 ( \60294 , \60293 );
buf \U$60320 ( \60295 , \60294 );
not \U$60321 ( \60296 , \60295 );
or \U$60322 ( \60297 , \59747 , \60296 );
buf \U$60323 ( \60298 , \59501 );
buf \U$60324 ( \60299 , \59742 );
nand \U$60325 ( \60300 , \60298 , \60299 );
buf \U$60326 ( \60301 , \60300 );
buf \U$60327 ( \60302 , \60301 );
nand \U$60328 ( \60303 , \60297 , \60302 );
buf \U$60329 ( \60304 , \60303 );
buf \U$60330 ( \60305 , \60304 );
buf \U$60331 ( \60306 , \59396 );
not \U$60332 ( \60307 , \60306 );
buf \U$60333 ( \60308 , \60307 );
buf \U$60334 ( \60309 , \60308 );
not \U$60335 ( \60310 , \60309 );
buf \U$60336 ( \60311 , \59278 );
not \U$60337 ( \60312 , \60311 );
or \U$60338 ( \60313 , \60310 , \60312 );
buf \U$60339 ( \60314 , \59278 );
buf \U$60340 ( \60315 , \60308 );
or \U$60341 ( \60316 , \60314 , \60315 );
nand \U$60342 ( \60317 , \60313 , \60316 );
buf \U$60343 ( \60318 , \60317 );
buf \U$60344 ( \60319 , \60318 );
buf \U$60345 ( \60320 , \59401 );
xor \U$60346 ( \60321 , \60319 , \60320 );
buf \U$60347 ( \60322 , \60321 );
buf \U$60348 ( \60323 , \60322 );
xor \U$60349 ( \60324 , \59430 , \59494 );
and \U$60350 ( \60325 , \60324 , \59499 );
and \U$60351 ( \60326 , \59430 , \59494 );
or \U$60352 ( \60327 , \60325 , \60326 );
buf \U$60353 ( \60328 , \60327 );
buf \U$60354 ( \60329 , \60328 );
or \U$60355 ( \60330 , \60323 , \60329 );
buf \U$60356 ( \60331 , \60330 );
buf \U$60357 ( \60332 , \60331 );
nand \U$60358 ( \60333 , \60305 , \60332 );
buf \U$60359 ( \60334 , \60333 );
buf \U$60360 ( \60335 , \60334 );
xor \U$60361 ( \60336 , \59967 , \60002 );
xor \U$60362 ( \60337 , \60336 , \60007 );
buf \U$60363 ( \60338 , \60337 );
buf \U$60364 ( \60339 , \60338 );
buf \U$60365 ( \60340 , RIc0d9400_64);
buf \U$60366 ( \60341 , RIc0dab70_114);
or \U$60367 ( \60342 , \60340 , \60341 );
buf \U$60368 ( \60343 , RIc0dabe8_115);
nand \U$60369 ( \60344 , \60342 , \60343 );
buf \U$60370 ( \60345 , \60344 );
buf \U$60371 ( \60346 , \60345 );
buf \U$60372 ( \60347 , RIc0d9400_64);
buf \U$60373 ( \60348 , RIc0dab70_114);
nand \U$60374 ( \60349 , \60347 , \60348 );
buf \U$60375 ( \60350 , \60349 );
buf \U$60376 ( \60351 , \60350 );
buf \U$60377 ( \60352 , RIc0daaf8_113);
and \U$60378 ( \60353 , \60346 , \60351 , \60352 );
buf \U$60379 ( \60354 , \60353 );
buf \U$60380 ( \60355 , \60354 );
buf \U$60381 ( \60356 , RIc0dabe8_115);
buf \U$60382 ( \60357 , RIc0d9310_62);
and \U$60383 ( \60358 , \60356 , \60357 );
not \U$60384 ( \60359 , \60356 );
buf \U$60385 ( \60360 , RIc0d9310_62);
not \U$60386 ( \60361 , \60360 );
buf \U$60387 ( \60362 , \60361 );
buf \U$60388 ( \60363 , \60362 );
and \U$60389 ( \60364 , \60359 , \60363 );
nor \U$60390 ( \60365 , \60358 , \60364 );
buf \U$60391 ( \60366 , \60365 );
buf \U$60392 ( \60367 , \60366 );
not \U$60393 ( \60368 , \60367 );
buf \U$60394 ( \60369 , \27743 );
not \U$60395 ( \60370 , \60369 );
or \U$60396 ( \60371 , \60368 , \60370 );
buf \U$60397 ( \60372 , \12303 );
buf \U$60398 ( \60373 , \60112 );
nand \U$60399 ( \60374 , \60372 , \60373 );
buf \U$60400 ( \60375 , \60374 );
buf \U$60401 ( \60376 , \60375 );
nand \U$60402 ( \60377 , \60371 , \60376 );
buf \U$60403 ( \60378 , \60377 );
buf \U$60404 ( \60379 , \60378 );
and \U$60405 ( \60380 , \60355 , \60379 );
buf \U$60406 ( \60381 , \60380 );
buf \U$60407 ( \60382 , \60381 );
buf \U$60408 ( \60383 , \13178 );
buf \U$60409 ( \60384 , RIc0dadc8_119);
buf \U$60410 ( \60385 , RIc0d9130_58);
xnor \U$60411 ( \60386 , \60384 , \60385 );
buf \U$60412 ( \60387 , \60386 );
buf \U$60413 ( \60388 , \60387 );
or \U$60414 ( \60389 , \60383 , \60388 );
buf \U$60415 ( \60390 , \45225 );
buf \U$60416 ( \60391 , \60171 );
not \U$60417 ( \60392 , \60391 );
buf \U$60418 ( \60393 , \60392 );
buf \U$60419 ( \60394 , \60393 );
or \U$60420 ( \60395 , \60390 , \60394 );
nand \U$60421 ( \60396 , \60389 , \60395 );
buf \U$60422 ( \60397 , \60396 );
buf \U$60423 ( \60398 , \60397 );
buf \U$60424 ( \60399 , RIc0d8e60_52);
buf \U$60425 ( \60400 , RIc0db098_125);
xor \U$60426 ( \60401 , \60399 , \60400 );
buf \U$60427 ( \60402 , \60401 );
buf \U$60428 ( \60403 , \60402 );
not \U$60429 ( \60404 , \60403 );
buf \U$60430 ( \60405 , \44382 );
not \U$60431 ( \60406 , \60405 );
or \U$60432 ( \60407 , \60404 , \60406 );
buf \U$60433 ( \60408 , \13465 );
buf \U$60434 ( \60409 , \60130 );
nand \U$60435 ( \60410 , \60408 , \60409 );
buf \U$60436 ( \60411 , \60410 );
buf \U$60437 ( \60412 , \60411 );
nand \U$60438 ( \60413 , \60407 , \60412 );
buf \U$60439 ( \60414 , \60413 );
buf \U$60440 ( \60415 , \60414 );
xor \U$60441 ( \60416 , \60398 , \60415 );
buf \U$60442 ( \60417 , RIc0db188_127);
buf \U$60443 ( \60418 , RIc0d8d70_50);
xor \U$60444 ( \60419 , \60417 , \60418 );
buf \U$60445 ( \60420 , \60419 );
buf \U$60446 ( \60421 , \60420 );
not \U$60447 ( \60422 , \60421 );
buf \U$60448 ( \60423 , \59144 );
not \U$60449 ( \60424 , \60423 );
or \U$60450 ( \60425 , \60422 , \60424 );
buf \U$60451 ( \60426 , \60156 );
buf \U$60452 ( \60427 , RIc0db200_128);
nand \U$60453 ( \60428 , \60426 , \60427 );
buf \U$60454 ( \60429 , \60428 );
buf \U$60455 ( \60430 , \60429 );
nand \U$60456 ( \60431 , \60425 , \60430 );
buf \U$60457 ( \60432 , \60431 );
buf \U$60458 ( \60433 , \60432 );
and \U$60459 ( \60434 , \60416 , \60433 );
and \U$60460 ( \60435 , \60398 , \60415 );
or \U$60461 ( \60436 , \60434 , \60435 );
buf \U$60462 ( \60437 , \60436 );
buf \U$60463 ( \60438 , \60437 );
xor \U$60464 ( \60439 , \60382 , \60438 );
buf \U$60465 ( \60440 , RIc0d9040_56);
buf \U$60466 ( \60441 , RIc0daeb8_121);
xor \U$60467 ( \60442 , \60440 , \60441 );
buf \U$60468 ( \60443 , \60442 );
buf \U$60469 ( \60444 , \60443 );
not \U$60470 ( \60445 , \60444 );
buf \U$60471 ( \60446 , \16382 );
not \U$60472 ( \60447 , \60446 );
or \U$60473 ( \60448 , \60445 , \60447 );
buf \U$60474 ( \60449 , \13314 );
buf \U$60475 ( \60450 , \60077 );
nand \U$60476 ( \60451 , \60449 , \60450 );
buf \U$60477 ( \60452 , \60451 );
buf \U$60478 ( \60453 , \60452 );
nand \U$60479 ( \60454 , \60448 , \60453 );
buf \U$60480 ( \60455 , \60454 );
buf \U$60481 ( \60456 , \60455 );
buf \U$60482 ( \60457 , RIc0d9220_60);
buf \U$60483 ( \60458 , RIc0dacd8_117);
xor \U$60484 ( \60459 , \60457 , \60458 );
buf \U$60485 ( \60460 , \60459 );
buf \U$60486 ( \60461 , \60460 );
not \U$60487 ( \60462 , \60461 );
buf \U$60488 ( \60463 , \22350 );
not \U$60489 ( \60464 , \60463 );
or \U$60490 ( \60465 , \60462 , \60464 );
buf \U$60491 ( \60466 , \12937 );
buf \U$60492 ( \60467 , \60190 );
nand \U$60493 ( \60468 , \60466 , \60467 );
buf \U$60494 ( \60469 , \60468 );
buf \U$60495 ( \60470 , \60469 );
nand \U$60496 ( \60471 , \60465 , \60470 );
buf \U$60497 ( \60472 , \60471 );
buf \U$60498 ( \60473 , \60472 );
xor \U$60499 ( \60474 , \60456 , \60473 );
buf \U$60500 ( \60475 , RIc0d8f50_54);
buf \U$60501 ( \60476 , RIc0dafa8_123);
xnor \U$60502 ( \60477 , \60475 , \60476 );
buf \U$60503 ( \60478 , \60477 );
buf \U$60504 ( \60479 , \60478 );
not \U$60505 ( \60480 , \60479 );
buf \U$60506 ( \60481 , \60480 );
buf \U$60507 ( \60482 , \60481 );
not \U$60508 ( \60483 , \60482 );
buf \U$60509 ( \60484 , \47037 );
not \U$60510 ( \60485 , \60484 );
or \U$60511 ( \60486 , \60483 , \60485 );
buf \U$60512 ( \60487 , \14278 );
buf \U$60513 ( \60488 , \60056 );
nand \U$60514 ( \60489 , \60487 , \60488 );
buf \U$60515 ( \60490 , \60489 );
buf \U$60516 ( \60491 , \60490 );
nand \U$60517 ( \60492 , \60486 , \60491 );
buf \U$60518 ( \60493 , \60492 );
buf \U$60519 ( \60494 , \60493 );
and \U$60520 ( \60495 , \60474 , \60494 );
and \U$60521 ( \60496 , \60456 , \60473 );
or \U$60522 ( \60497 , \60495 , \60496 );
buf \U$60523 ( \60498 , \60497 );
buf \U$60524 ( \60499 , \60498 );
and \U$60525 ( \60500 , \60439 , \60499 );
and \U$60526 ( \60501 , \60382 , \60438 );
or \U$60527 ( \60502 , \60500 , \60501 );
buf \U$60528 ( \60503 , \60502 );
buf \U$60529 ( \60504 , \60503 );
xor \U$60530 ( \60505 , \60167 , \60185 );
xor \U$60531 ( \60506 , \60505 , \60203 );
buf \U$60532 ( \60507 , \60506 );
buf \U$60533 ( \60508 , \60507 );
not \U$60534 ( \60509 , \60508 );
xor \U$60535 ( \60510 , \60108 , \60125 );
xor \U$60536 ( \60511 , \60510 , \60144 );
buf \U$60537 ( \60512 , \60511 );
buf \U$60538 ( \60513 , \60512 );
not \U$60539 ( \60514 , \60513 );
or \U$60540 ( \60515 , \60509 , \60514 );
buf \U$60541 ( \60516 , \60507 );
buf \U$60542 ( \60517 , \60512 );
or \U$60543 ( \60518 , \60516 , \60517 );
buf \U$60544 ( \60519 , \60069 );
not \U$60545 ( \60520 , \60519 );
buf \U$60546 ( \60521 , \60520 );
buf \U$60547 ( \60522 , \60521 );
not \U$60548 ( \60523 , \60522 );
buf \U$60549 ( \60524 , \60051 );
not \U$60550 ( \60525 , \60524 );
buf \U$60551 ( \60526 , \60093 );
not \U$60552 ( \60527 , \60526 );
or \U$60553 ( \60528 , \60525 , \60527 );
buf \U$60554 ( \60529 , \60093 );
buf \U$60555 ( \60530 , \60051 );
or \U$60556 ( \60531 , \60529 , \60530 );
nand \U$60557 ( \60532 , \60528 , \60531 );
buf \U$60558 ( \60533 , \60532 );
buf \U$60559 ( \60534 , \60533 );
not \U$60560 ( \60535 , \60534 );
or \U$60561 ( \60536 , \60523 , \60535 );
buf \U$60562 ( \60537 , \60533 );
buf \U$60563 ( \60538 , \60521 );
or \U$60564 ( \60539 , \60537 , \60538 );
nand \U$60565 ( \60540 , \60536 , \60539 );
buf \U$60566 ( \60541 , \60540 );
buf \U$60567 ( \60542 , \60541 );
nand \U$60568 ( \60543 , \60518 , \60542 );
buf \U$60569 ( \60544 , \60543 );
buf \U$60570 ( \60545 , \60544 );
nand \U$60571 ( \60546 , \60515 , \60545 );
buf \U$60572 ( \60547 , \60546 );
buf \U$60573 ( \60548 , \60547 );
xor \U$60574 ( \60549 , \60504 , \60548 );
xor \U$60575 ( \60550 , \60207 , \60148 );
xor \U$60576 ( \60551 , \60550 , \60102 );
buf \U$60577 ( \60552 , \60551 );
and \U$60578 ( \60553 , \60549 , \60552 );
and \U$60579 ( \60554 , \60504 , \60548 );
or \U$60580 ( \60555 , \60553 , \60554 );
buf \U$60581 ( \60556 , \60555 );
buf \U$60582 ( \60557 , \60556 );
xor \U$60583 ( \60558 , \60339 , \60557 );
xor \U$60584 ( \60559 , \60219 , \60223 );
xor \U$60585 ( \60560 , \60559 , \60242 );
buf \U$60586 ( \60561 , \60560 );
buf \U$60587 ( \60562 , \60561 );
and \U$60588 ( \60563 , \60558 , \60562 );
and \U$60589 ( \60564 , \60339 , \60557 );
or \U$60590 ( \60565 , \60563 , \60564 );
buf \U$60591 ( \60566 , \60565 );
buf \U$60592 ( \60567 , \60566 );
not \U$60593 ( \60568 , \60567 );
buf \U$60594 ( \60569 , \60028 );
not \U$60595 ( \60570 , \60569 );
buf \U$60596 ( \60571 , \60570 );
buf \U$60597 ( \60572 , \60571 );
not \U$60598 ( \60573 , \60572 );
buf \U$60599 ( \60574 , \60246 );
not \U$60600 ( \60575 , \60574 );
or \U$60601 ( \60576 , \60573 , \60575 );
buf \U$60602 ( \60577 , \60246 );
buf \U$60603 ( \60578 , \60571 );
or \U$60604 ( \60579 , \60577 , \60578 );
nand \U$60605 ( \60580 , \60576 , \60579 );
buf \U$60606 ( \60581 , \60580 );
buf \U$60607 ( \60582 , \60581 );
buf \U$60608 ( \60583 , \60255 );
xnor \U$60609 ( \60584 , \60582 , \60583 );
buf \U$60610 ( \60585 , \60584 );
buf \U$60611 ( \60586 , \60585 );
nand \U$60612 ( \60587 , \60568 , \60586 );
buf \U$60613 ( \60588 , \60587 );
buf \U$60614 ( \60589 , \60588 );
xor \U$60615 ( \60590 , \60339 , \60557 );
xor \U$60616 ( \60591 , \60590 , \60562 );
buf \U$60617 ( \60592 , \60591 );
buf \U$60618 ( \60593 , \60592 );
xor \U$60619 ( \60594 , \60228 , \60232 );
xor \U$60620 ( \60595 , \60594 , \60237 );
buf \U$60621 ( \60596 , \60595 );
buf \U$60622 ( \60597 , \60596 );
buf \U$60623 ( \60598 , RIc0d9400_64);
buf \U$60624 ( \60599 , RIc0daaf8_113);
xor \U$60625 ( \60600 , \60598 , \60599 );
buf \U$60626 ( \60601 , \60600 );
buf \U$60627 ( \60602 , \60601 );
not \U$60628 ( \60603 , \60602 );
buf \U$60629 ( \60604 , \25355 );
not \U$60630 ( \60605 , \60604 );
or \U$60631 ( \60606 , \60603 , \60605 );
buf \U$60632 ( \60607 , \16995 );
buf \U$60633 ( \60608 , \60038 );
nand \U$60634 ( \60609 , \60607 , \60608 );
buf \U$60635 ( \60610 , \60609 );
buf \U$60636 ( \60611 , \60610 );
nand \U$60637 ( \60612 , \60606 , \60611 );
buf \U$60638 ( \60613 , \60612 );
buf \U$60639 ( \60614 , \60613 );
not \U$60640 ( \60615 , \60614 );
xor \U$60641 ( \60616 , \60355 , \60379 );
buf \U$60642 ( \60617 , \60616 );
buf \U$60643 ( \60618 , \60617 );
not \U$60644 ( \60619 , \60618 );
or \U$60645 ( \60620 , \60615 , \60619 );
buf \U$60646 ( \60621 , \60617 );
buf \U$60647 ( \60622 , \60613 );
or \U$60648 ( \60623 , \60621 , \60622 );
buf \U$60649 ( \60624 , \16662 );
buf \U$60650 ( \60625 , RIc0d9400_64);
and \U$60651 ( \60626 , \60624 , \60625 );
buf \U$60652 ( \60627 , \60626 );
buf \U$60653 ( \60628 , \60627 );
buf \U$60654 ( \60629 , RIc0d9298_61);
buf \U$60655 ( \60630 , RIc0dacd8_117);
xor \U$60656 ( \60631 , \60629 , \60630 );
buf \U$60657 ( \60632 , \60631 );
buf \U$60658 ( \60633 , \60632 );
not \U$60659 ( \60634 , \60633 );
buf \U$60660 ( \60635 , \22350 );
not \U$60661 ( \60636 , \60635 );
or \U$60662 ( \60637 , \60634 , \60636 );
buf \U$60663 ( \60638 , \12937 );
buf \U$60664 ( \60639 , \60460 );
nand \U$60665 ( \60640 , \60638 , \60639 );
buf \U$60666 ( \60641 , \60640 );
buf \U$60667 ( \60642 , \60641 );
nand \U$60668 ( \60643 , \60637 , \60642 );
buf \U$60669 ( \60644 , \60643 );
buf \U$60670 ( \60645 , \60644 );
xor \U$60671 ( \60646 , \60628 , \60645 );
buf \U$60672 ( \60647 , \16688 );
buf \U$60673 ( \60648 , RIc0d8fc8_55);
buf \U$60674 ( \60649 , RIc0dafa8_123);
xnor \U$60675 ( \60650 , \60648 , \60649 );
buf \U$60676 ( \60651 , \60650 );
buf \U$60677 ( \60652 , \60651 );
or \U$60678 ( \60653 , \60647 , \60652 );
buf \U$60679 ( \60654 , \16695 );
buf \U$60680 ( \60655 , \60478 );
or \U$60681 ( \60656 , \60654 , \60655 );
nand \U$60682 ( \60657 , \60653 , \60656 );
buf \U$60683 ( \60658 , \60657 );
buf \U$60684 ( \60659 , \60658 );
and \U$60685 ( \60660 , \60646 , \60659 );
and \U$60686 ( \60661 , \60628 , \60645 );
or \U$60687 ( \60662 , \60660 , \60661 );
buf \U$60688 ( \60663 , \60662 );
buf \U$60689 ( \60664 , \60663 );
nand \U$60690 ( \60665 , \60623 , \60664 );
buf \U$60691 ( \60666 , \60665 );
buf \U$60692 ( \60667 , \60666 );
nand \U$60693 ( \60668 , \60620 , \60667 );
buf \U$60694 ( \60669 , \60668 );
buf \U$60695 ( \60670 , \60669 );
buf \U$60696 ( \60671 , RIc0db200_128);
not \U$60697 ( \60672 , \60671 );
buf \U$60698 ( \60673 , \60420 );
not \U$60699 ( \60674 , \60673 );
or \U$60700 ( \60675 , \60672 , \60674 );
buf \U$60701 ( \60676 , \60151 );
xor \U$60702 ( \60677 , RIc0db188_127, RIc0d8de8_51);
buf \U$60703 ( \60678 , \60677 );
not \U$60704 ( \60679 , \60678 );
buf \U$60705 ( \60680 , \60679 );
buf \U$60706 ( \60681 , \60680 );
or \U$60707 ( \60682 , \60676 , \60681 );
nand \U$60708 ( \60683 , \60675 , \60682 );
buf \U$60709 ( \60684 , \60683 );
buf \U$60710 ( \60685 , \60684 );
buf \U$60711 ( \60686 , RIc0d91a8_59);
buf \U$60712 ( \60687 , RIc0dadc8_119);
xor \U$60713 ( \60688 , \60686 , \60687 );
buf \U$60714 ( \60689 , \60688 );
buf \U$60715 ( \60690 , \60689 );
not \U$60716 ( \60691 , \60690 );
buf \U$60717 ( \60692 , \14569 );
not \U$60718 ( \60693 , \60692 );
or \U$60719 ( \60694 , \60691 , \60693 );
buf \U$60720 ( \60695 , \60387 );
not \U$60721 ( \60696 , \60695 );
buf \U$60722 ( \60697 , \13953 );
nand \U$60723 ( \60698 , \60696 , \60697 );
buf \U$60724 ( \60699 , \60698 );
buf \U$60725 ( \60700 , \60699 );
nand \U$60726 ( \60701 , \60694 , \60700 );
buf \U$60727 ( \60702 , \60701 );
buf \U$60728 ( \60703 , \60702 );
xor \U$60729 ( \60704 , \60685 , \60703 );
buf \U$60730 ( \60705 , RIc0d8ed8_53);
buf \U$60731 ( \60706 , RIc0db098_125);
xor \U$60732 ( \60707 , \60705 , \60706 );
buf \U$60733 ( \60708 , \60707 );
buf \U$60734 ( \60709 , \60708 );
not \U$60735 ( \60710 , \60709 );
buf \U$60736 ( \60711 , \51095 );
not \U$60737 ( \60712 , \60711 );
or \U$60738 ( \60713 , \60710 , \60712 );
buf \U$60739 ( \60714 , \15793 );
buf \U$60740 ( \60715 , \60402 );
nand \U$60741 ( \60716 , \60714 , \60715 );
buf \U$60742 ( \60717 , \60716 );
buf \U$60743 ( \60718 , \60717 );
nand \U$60744 ( \60719 , \60713 , \60718 );
buf \U$60745 ( \60720 , \60719 );
buf \U$60746 ( \60721 , \60720 );
and \U$60747 ( \60722 , \60704 , \60721 );
and \U$60748 ( \60723 , \60685 , \60703 );
or \U$60749 ( \60724 , \60722 , \60723 );
buf \U$60750 ( \60725 , \60724 );
buf \U$60751 ( \60726 , \60725 );
not \U$60752 ( \60727 , \60726 );
xor \U$60753 ( \60728 , \60456 , \60473 );
xor \U$60754 ( \60729 , \60728 , \60494 );
buf \U$60755 ( \60730 , \60729 );
buf \U$60756 ( \60731 , \60730 );
not \U$60757 ( \60732 , \60731 );
or \U$60758 ( \60733 , \60727 , \60732 );
buf \U$60759 ( \60734 , \60730 );
buf \U$60760 ( \60735 , \60725 );
or \U$60761 ( \60736 , \60734 , \60735 );
xor \U$60762 ( \60737 , \60398 , \60415 );
xor \U$60763 ( \60738 , \60737 , \60433 );
buf \U$60764 ( \60739 , \60738 );
buf \U$60765 ( \60740 , \60739 );
nand \U$60766 ( \60741 , \60736 , \60740 );
buf \U$60767 ( \60742 , \60741 );
buf \U$60768 ( \60743 , \60742 );
nand \U$60769 ( \60744 , \60733 , \60743 );
buf \U$60770 ( \60745 , \60744 );
buf \U$60771 ( \60746 , \60745 );
xor \U$60772 ( \60747 , \60670 , \60746 );
xor \U$60773 ( \60748 , \60382 , \60438 );
xor \U$60774 ( \60749 , \60748 , \60499 );
buf \U$60775 ( \60750 , \60749 );
buf \U$60776 ( \60751 , \60750 );
and \U$60777 ( \60752 , \60747 , \60751 );
and \U$60778 ( \60753 , \60670 , \60746 );
or \U$60779 ( \60754 , \60752 , \60753 );
buf \U$60780 ( \60755 , \60754 );
buf \U$60781 ( \60756 , \60755 );
xor \U$60782 ( \60757 , \60597 , \60756 );
xor \U$60783 ( \60758 , \60504 , \60548 );
xor \U$60784 ( \60759 , \60758 , \60552 );
buf \U$60785 ( \60760 , \60759 );
buf \U$60786 ( \60761 , \60760 );
and \U$60787 ( \60762 , \60757 , \60761 );
and \U$60788 ( \60763 , \60597 , \60756 );
or \U$60789 ( \60764 , \60762 , \60763 );
buf \U$60790 ( \60765 , \60764 );
buf \U$60791 ( \60766 , \60765 );
or \U$60792 ( \60767 , \60593 , \60766 );
buf \U$60793 ( \60768 , \60767 );
buf \U$60794 ( \60769 , \60768 );
and \U$60795 ( \60770 , \60589 , \60769 );
buf \U$60796 ( \60771 , \60770 );
buf \U$60797 ( \60772 , \60771 );
buf \U$60798 ( \60773 , \54203 );
buf \U$60799 ( \60774 , RIc0d8fc8_55);
buf \U$60800 ( \60775 , RIc0db098_125);
xnor \U$60801 ( \60776 , \60774 , \60775 );
buf \U$60802 ( \60777 , \60776 );
buf \U$60803 ( \60778 , \60777 );
or \U$60804 ( \60779 , \60773 , \60778 );
buf \U$60805 ( \60780 , \22744 );
buf \U$60806 ( \60781 , RIc0d8f50_54);
buf \U$60807 ( \60782 , RIc0db098_125);
xor \U$60808 ( \60783 , \60781 , \60782 );
buf \U$60809 ( \60784 , \60783 );
buf \U$60810 ( \60785 , \60784 );
not \U$60811 ( \60786 , \60785 );
buf \U$60812 ( \60787 , \60786 );
buf \U$60813 ( \60788 , \60787 );
or \U$60814 ( \60789 , \60780 , \60788 );
nand \U$60815 ( \60790 , \60779 , \60789 );
buf \U$60816 ( \60791 , \60790 );
buf \U$60817 ( \60792 , \60791 );
buf \U$60818 ( \60793 , RIc0d9400_64);
buf \U$60819 ( \60794 , RIc0dad50_118);
or \U$60820 ( \60795 , \60793 , \60794 );
buf \U$60821 ( \60796 , RIc0dadc8_119);
nand \U$60822 ( \60797 , \60795 , \60796 );
buf \U$60823 ( \60798 , \60797 );
buf \U$60824 ( \60799 , \60798 );
buf \U$60825 ( \60800 , RIc0d9400_64);
buf \U$60826 ( \60801 , RIc0dad50_118);
nand \U$60827 ( \60802 , \60800 , \60801 );
buf \U$60828 ( \60803 , \60802 );
buf \U$60829 ( \60804 , \60803 );
buf \U$60830 ( \60805 , RIc0dacd8_117);
and \U$60831 ( \60806 , \60799 , \60804 , \60805 );
buf \U$60832 ( \60807 , \60806 );
buf \U$60833 ( \60808 , \60807 );
buf \U$60834 ( \60809 , RIc0d9310_62);
buf \U$60835 ( \60810 , RIc0dadc8_119);
xor \U$60836 ( \60811 , \60809 , \60810 );
buf \U$60837 ( \60812 , \60811 );
buf \U$60838 ( \60813 , \60812 );
not \U$60839 ( \60814 , \60813 );
buf \U$60840 ( \60815 , \13949 );
not \U$60841 ( \60816 , \60815 );
or \U$60842 ( \60817 , \60814 , \60816 );
buf \U$60843 ( \60818 , \13953 );
buf \U$60844 ( \60819 , RIc0dadc8_119);
buf \U$60845 ( \60820 , RIc0d9298_61);
xor \U$60846 ( \60821 , \60819 , \60820 );
buf \U$60847 ( \60822 , \60821 );
buf \U$60848 ( \60823 , \60822 );
nand \U$60849 ( \60824 , \60818 , \60823 );
buf \U$60850 ( \60825 , \60824 );
buf \U$60851 ( \60826 , \60825 );
nand \U$60852 ( \60827 , \60817 , \60826 );
buf \U$60853 ( \60828 , \60827 );
buf \U$60854 ( \60829 , \60828 );
and \U$60855 ( \60830 , \60808 , \60829 );
buf \U$60856 ( \60831 , \60830 );
buf \U$60857 ( \60832 , \60831 );
xor \U$60858 ( \60833 , \60792 , \60832 );
buf \U$60859 ( \60834 , RIc0daeb8_121);
buf \U$60860 ( \60835 , RIc0d9220_60);
xor \U$60861 ( \60836 , \60834 , \60835 );
buf \U$60862 ( \60837 , \60836 );
buf \U$60863 ( \60838 , \60837 );
not \U$60864 ( \60839 , \60838 );
buf \U$60865 ( \60840 , \13310 );
not \U$60866 ( \60841 , \60840 );
or \U$60867 ( \60842 , \60839 , \60841 );
buf \U$60868 ( \60843 , \16386 );
buf \U$60869 ( \60844 , RIc0daeb8_121);
buf \U$60870 ( \60845 , RIc0d91a8_59);
xor \U$60871 ( \60846 , \60844 , \60845 );
buf \U$60872 ( \60847 , \60846 );
buf \U$60873 ( \60848 , \60847 );
nand \U$60874 ( \60849 , \60843 , \60848 );
buf \U$60875 ( \60850 , \60849 );
buf \U$60876 ( \60851 , \60850 );
nand \U$60877 ( \60852 , \60842 , \60851 );
buf \U$60878 ( \60853 , \60852 );
buf \U$60879 ( \60854 , \60853 );
buf \U$60880 ( \60855 , RIc0dacd8_117);
buf \U$60881 ( \60856 , RIc0d9400_64);
and \U$60882 ( \60857 , \60855 , \60856 );
not \U$60883 ( \60858 , \60855 );
buf \U$60884 ( \60859 , \43843 );
and \U$60885 ( \60860 , \60858 , \60859 );
nor \U$60886 ( \60861 , \60857 , \60860 );
buf \U$60887 ( \60862 , \60861 );
buf \U$60888 ( \60863 , \60862 );
not \U$60889 ( \60864 , \60863 );
buf \U$60890 ( \60865 , \12929 );
not \U$60891 ( \60866 , \60865 );
or \U$60892 ( \60867 , \60864 , \60866 );
buf \U$60893 ( \60868 , \12937 );
buf \U$60894 ( \60869 , RIc0dacd8_117);
buf \U$60895 ( \60870 , RIc0d9388_63);
xor \U$60896 ( \60871 , \60869 , \60870 );
buf \U$60897 ( \60872 , \60871 );
buf \U$60898 ( \60873 , \60872 );
nand \U$60899 ( \60874 , \60868 , \60873 );
buf \U$60900 ( \60875 , \60874 );
buf \U$60901 ( \60876 , \60875 );
nand \U$60902 ( \60877 , \60867 , \60876 );
buf \U$60903 ( \60878 , \60877 );
buf \U$60904 ( \60879 , \60878 );
xor \U$60905 ( \60880 , \60854 , \60879 );
buf \U$60906 ( \60881 , \45089 );
xor \U$60907 ( \60882 , RIc0dafa8_123, RIc0d9130_58);
buf \U$60908 ( \60883 , \60882 );
not \U$60909 ( \60884 , \60883 );
buf \U$60910 ( \60885 , \60884 );
buf \U$60911 ( \60886 , \60885 );
or \U$60912 ( \60887 , \60881 , \60886 );
buf \U$60913 ( \60888 , \14275 );
buf \U$60914 ( \60889 , RIc0d90b8_57);
buf \U$60915 ( \60890 , RIc0dafa8_123);
xor \U$60916 ( \60891 , \60889 , \60890 );
buf \U$60917 ( \60892 , \60891 );
buf \U$60918 ( \60893 , \60892 );
not \U$60919 ( \60894 , \60893 );
buf \U$60920 ( \60895 , \60894 );
buf \U$60921 ( \60896 , \60895 );
or \U$60922 ( \60897 , \60888 , \60896 );
nand \U$60923 ( \60898 , \60887 , \60897 );
buf \U$60924 ( \60899 , \60898 );
buf \U$60925 ( \60900 , \60899 );
and \U$60926 ( \60901 , \60880 , \60900 );
and \U$60927 ( \60902 , \60854 , \60879 );
or \U$60928 ( \60903 , \60901 , \60902 );
buf \U$60929 ( \60904 , \60903 );
buf \U$60930 ( \60905 , \60904 );
xor \U$60931 ( \60906 , \60833 , \60905 );
buf \U$60932 ( \60907 , \60906 );
buf \U$60933 ( \60908 , \60907 );
not \U$60934 ( \60909 , \60908 );
not \U$60935 ( \60910 , \43781 );
not \U$60936 ( \60911 , \60910 );
not \U$60937 ( \60912 , \60911 );
buf \U$60938 ( \60913 , \60912 );
xor \U$60939 ( \60914 , RIc0db188_127, RIc0d8fc8_55);
buf \U$60940 ( \60915 , \60914 );
not \U$60941 ( \60916 , \60915 );
buf \U$60942 ( \60917 , \60916 );
buf \U$60943 ( \60918 , \60917 );
or \U$60944 ( \60919 , \60913 , \60918 );
buf \U$60945 ( \60920 , \12647 );
buf \U$60946 ( \60921 , RIc0db188_127);
buf \U$60947 ( \60922 , RIc0d8f50_54);
xnor \U$60948 ( \60923 , \60921 , \60922 );
buf \U$60949 ( \60924 , \60923 );
buf \U$60950 ( \60925 , \60924 );
or \U$60951 ( \60926 , \60920 , \60925 );
nand \U$60952 ( \60927 , \60919 , \60926 );
buf \U$60953 ( \60928 , \60927 );
buf \U$60954 ( \60929 , \60928 );
not \U$60955 ( \60930 , \60929 );
buf \U$60956 ( \60931 , RIc0d91a8_59);
buf \U$60957 ( \60932 , RIc0dafa8_123);
xor \U$60958 ( \60933 , \60931 , \60932 );
buf \U$60959 ( \60934 , \60933 );
buf \U$60960 ( \60935 , \60934 );
not \U$60961 ( \60936 , \60935 );
buf \U$60962 ( \60937 , \14982 );
not \U$60963 ( \60938 , \60937 );
or \U$60964 ( \60939 , \60936 , \60938 );
buf \U$60965 ( \60940 , \16692 );
buf \U$60966 ( \60941 , \60882 );
nand \U$60967 ( \60942 , \60940 , \60941 );
buf \U$60968 ( \60943 , \60942 );
buf \U$60969 ( \60944 , \60943 );
nand \U$60970 ( \60945 , \60939 , \60944 );
buf \U$60971 ( \60946 , \60945 );
buf \U$60972 ( \60947 , \60946 );
not \U$60973 ( \60948 , \60947 );
or \U$60974 ( \60949 , \60930 , \60948 );
buf \U$60975 ( \60950 , \60946 );
buf \U$60976 ( \60951 , \60928 );
or \U$60977 ( \60952 , \60950 , \60951 );
buf \U$60978 ( \60953 , RIc0db098_125);
buf \U$60979 ( \60954 , RIc0d90b8_57);
xor \U$60980 ( \60955 , \60953 , \60954 );
buf \U$60981 ( \60956 , \60955 );
buf \U$60982 ( \60957 , \60956 );
not \U$60983 ( \60958 , \60957 );
buf \U$60984 ( \60959 , \13461 );
not \U$60985 ( \60960 , \60959 );
or \U$60986 ( \60961 , \60958 , \60960 );
buf \U$60987 ( \60962 , \13465 );
buf \U$60988 ( \60963 , RIc0d9040_56);
buf \U$60989 ( \60964 , RIc0db098_125);
xor \U$60990 ( \60965 , \60963 , \60964 );
buf \U$60991 ( \60966 , \60965 );
buf \U$60992 ( \60967 , \60966 );
nand \U$60993 ( \60968 , \60962 , \60967 );
buf \U$60994 ( \60969 , \60968 );
buf \U$60995 ( \60970 , \60969 );
nand \U$60996 ( \60971 , \60961 , \60970 );
buf \U$60997 ( \60972 , \60971 );
buf \U$60998 ( \60973 , \60972 );
nand \U$60999 ( \60974 , \60952 , \60973 );
buf \U$61000 ( \60975 , \60974 );
buf \U$61001 ( \60976 , \60975 );
nand \U$61002 ( \60977 , \60949 , \60976 );
buf \U$61003 ( \60978 , \60977 );
buf \U$61004 ( \60979 , \60978 );
buf \U$61005 ( \60980 , \16556 );
buf \U$61006 ( \60981 , \43843 );
nor \U$61007 ( \60982 , \60980 , \60981 );
buf \U$61008 ( \60983 , \60982 );
buf \U$61009 ( \60984 , \60983 );
buf \U$61010 ( \60985 , RIc0d9298_61);
buf \U$61011 ( \60986 , RIc0daeb8_121);
xor \U$61012 ( \60987 , \60985 , \60986 );
buf \U$61013 ( \60988 , \60987 );
buf \U$61014 ( \60989 , \60988 );
not \U$61015 ( \60990 , \60989 );
buf \U$61016 ( \60991 , \16382 );
not \U$61017 ( \60992 , \60991 );
or \U$61018 ( \60993 , \60990 , \60992 );
buf \U$61019 ( \60994 , \12975 );
buf \U$61020 ( \60995 , \60837 );
nand \U$61021 ( \60996 , \60994 , \60995 );
buf \U$61022 ( \60997 , \60996 );
buf \U$61023 ( \60998 , \60997 );
nand \U$61024 ( \60999 , \60993 , \60998 );
buf \U$61025 ( \61000 , \60999 );
buf \U$61026 ( \61001 , \61000 );
xor \U$61027 ( \61002 , \60984 , \61001 );
buf \U$61028 ( \61003 , \13178 );
buf \U$61029 ( \61004 , RIc0dadc8_119);
buf \U$61030 ( \61005 , \43939 );
and \U$61031 ( \61006 , \61004 , \61005 );
not \U$61032 ( \61007 , \61004 );
buf \U$61033 ( \61008 , RIc0d9388_63);
and \U$61034 ( \61009 , \61007 , \61008 );
nor \U$61035 ( \61010 , \61006 , \61009 );
buf \U$61036 ( \61011 , \61010 );
buf \U$61037 ( \61012 , \61011 );
or \U$61038 ( \61013 , \61003 , \61012 );
buf \U$61039 ( \61014 , \45225 );
buf \U$61040 ( \61015 , \60812 );
not \U$61041 ( \61016 , \61015 );
buf \U$61042 ( \61017 , \61016 );
buf \U$61043 ( \61018 , \61017 );
or \U$61044 ( \61019 , \61014 , \61018 );
nand \U$61045 ( \61020 , \61013 , \61019 );
buf \U$61046 ( \61021 , \61020 );
buf \U$61047 ( \61022 , \61021 );
and \U$61048 ( \61023 , \61002 , \61022 );
and \U$61049 ( \61024 , \60984 , \61001 );
or \U$61050 ( \61025 , \61023 , \61024 );
buf \U$61051 ( \61026 , \61025 );
buf \U$61052 ( \61027 , \61026 );
xor \U$61053 ( \61028 , \60979 , \61027 );
xor \U$61054 ( \61029 , \60854 , \60879 );
xor \U$61055 ( \61030 , \61029 , \60900 );
buf \U$61056 ( \61031 , \61030 );
buf \U$61057 ( \61032 , \61031 );
and \U$61058 ( \61033 , \61028 , \61032 );
and \U$61059 ( \61034 , \60979 , \61027 );
or \U$61060 ( \61035 , \61033 , \61034 );
buf \U$61061 ( \61036 , \61035 );
buf \U$61062 ( \61037 , \61036 );
not \U$61063 ( \61038 , \61037 );
or \U$61064 ( \61039 , \60909 , \61038 );
buf \U$61065 ( \61040 , \61036 );
buf \U$61066 ( \61041 , \60907 );
or \U$61067 ( \61042 , \61040 , \61041 );
buf \U$61068 ( \61043 , \14690 );
buf \U$61069 ( \61044 , RIc0d9400_64);
and \U$61070 ( \61045 , \61043 , \61044 );
buf \U$61071 ( \61046 , \61045 );
buf \U$61072 ( \61047 , \61046 );
buf \U$61073 ( \61048 , \60847 );
not \U$61074 ( \61049 , \61048 );
buf \U$61075 ( \61050 , \19487 );
not \U$61076 ( \61051 , \61050 );
or \U$61077 ( \61052 , \61049 , \61051 );
buf \U$61078 ( \61053 , \13314 );
buf \U$61079 ( \61054 , RIc0daeb8_121);
buf \U$61080 ( \61055 , RIc0d9130_58);
xor \U$61081 ( \61056 , \61054 , \61055 );
buf \U$61082 ( \61057 , \61056 );
buf \U$61083 ( \61058 , \61057 );
nand \U$61084 ( \61059 , \61053 , \61058 );
buf \U$61085 ( \61060 , \61059 );
buf \U$61086 ( \61061 , \61060 );
nand \U$61087 ( \61062 , \61052 , \61061 );
buf \U$61088 ( \61063 , \61062 );
buf \U$61089 ( \61064 , \61063 );
xor \U$61090 ( \61065 , \61047 , \61064 );
buf \U$61091 ( \61066 , \60822 );
not \U$61092 ( \61067 , \61066 );
buf \U$61093 ( \61068 , \14569 );
not \U$61094 ( \61069 , \61068 );
or \U$61095 ( \61070 , \61067 , \61069 );
buf \U$61096 ( \61071 , \13953 );
buf \U$61097 ( \61072 , RIc0d9220_60);
buf \U$61098 ( \61073 , RIc0dadc8_119);
xor \U$61099 ( \61074 , \61072 , \61073 );
buf \U$61100 ( \61075 , \61074 );
buf \U$61101 ( \61076 , \61075 );
nand \U$61102 ( \61077 , \61071 , \61076 );
buf \U$61103 ( \61078 , \61077 );
buf \U$61104 ( \61079 , \61078 );
nand \U$61105 ( \61080 , \61070 , \61079 );
buf \U$61106 ( \61081 , \61080 );
buf \U$61107 ( \61082 , \61081 );
xor \U$61108 ( \61083 , \61065 , \61082 );
buf \U$61109 ( \61084 , \61083 );
buf \U$61110 ( \61085 , \61084 );
not \U$61111 ( \61086 , \61085 );
buf \U$61112 ( \61087 , \60872 );
not \U$61113 ( \61088 , \61087 );
buf \U$61114 ( \61089 , \12923 );
not \U$61115 ( \61090 , \61089 );
or \U$61116 ( \61091 , \61088 , \61090 );
buf \U$61117 ( \61092 , \16559 );
buf \U$61118 ( \61093 , RIc0dacd8_117);
buf \U$61119 ( \61094 , RIc0d9310_62);
xor \U$61120 ( \61095 , \61093 , \61094 );
buf \U$61121 ( \61096 , \61095 );
buf \U$61122 ( \61097 , \61096 );
nand \U$61123 ( \61098 , \61092 , \61097 );
buf \U$61124 ( \61099 , \61098 );
buf \U$61125 ( \61100 , \61099 );
nand \U$61126 ( \61101 , \61091 , \61100 );
buf \U$61127 ( \61102 , \61101 );
buf \U$61128 ( \61103 , \61102 );
not \U$61129 ( \61104 , \61103 );
buf \U$61130 ( \61105 , \61104 );
buf \U$61131 ( \61106 , \61105 );
buf \U$61132 ( \61107 , RIc0d8ed8_53);
buf \U$61133 ( \61108 , RIc0db188_127);
xor \U$61134 ( \61109 , \61107 , \61108 );
buf \U$61135 ( \61110 , \61109 );
buf \U$61136 ( \61111 , \61110 );
not \U$61137 ( \61112 , \61111 );
buf \U$61138 ( \61113 , \15609 );
not \U$61139 ( \61114 , \61113 );
or \U$61140 ( \61115 , \61112 , \61114 );
buf \U$61141 ( \61116 , RIc0d8e60_52);
buf \U$61142 ( \61117 , RIc0db188_127);
xor \U$61143 ( \61118 , \61116 , \61117 );
buf \U$61144 ( \61119 , \61118 );
buf \U$61145 ( \61120 , \61119 );
buf \U$61146 ( \61121 , RIc0db200_128);
nand \U$61147 ( \61122 , \61120 , \61121 );
buf \U$61148 ( \61123 , \61122 );
buf \U$61149 ( \61124 , \61123 );
nand \U$61150 ( \61125 , \61115 , \61124 );
buf \U$61151 ( \61126 , \61125 );
buf \U$61152 ( \61127 , \61126 );
not \U$61153 ( \61128 , \61127 );
buf \U$61154 ( \61129 , \61128 );
buf \U$61155 ( \61130 , \61129 );
and \U$61156 ( \61131 , \61106 , \61130 );
not \U$61157 ( \61132 , \61106 );
buf \U$61158 ( \61133 , \61126 );
and \U$61159 ( \61134 , \61132 , \61133 );
nor \U$61160 ( \61135 , \61131 , \61134 );
buf \U$61161 ( \61136 , \61135 );
buf \U$61162 ( \61137 , \61136 );
buf \U$61163 ( \61138 , \60892 );
not \U$61164 ( \61139 , \61138 );
buf \U$61165 ( \61140 , \14982 );
not \U$61166 ( \61141 , \61140 );
or \U$61167 ( \61142 , \61139 , \61141 );
buf \U$61168 ( \61143 , \14278 );
buf \U$61169 ( \61144 , RIc0d9040_56);
buf \U$61170 ( \61145 , RIc0dafa8_123);
xor \U$61171 ( \61146 , \61144 , \61145 );
buf \U$61172 ( \61147 , \61146 );
buf \U$61173 ( \61148 , \61147 );
nand \U$61174 ( \61149 , \61143 , \61148 );
buf \U$61175 ( \61150 , \61149 );
buf \U$61176 ( \61151 , \61150 );
nand \U$61177 ( \61152 , \61142 , \61151 );
buf \U$61178 ( \61153 , \61152 );
buf \U$61179 ( \61154 , \61153 );
not \U$61180 ( \61155 , \61154 );
buf \U$61181 ( \61156 , \61155 );
buf \U$61182 ( \61157 , \61156 );
and \U$61183 ( \61158 , \61137 , \61157 );
not \U$61184 ( \61159 , \61137 );
buf \U$61185 ( \61160 , \61153 );
and \U$61186 ( \61161 , \61159 , \61160 );
nor \U$61187 ( \61162 , \61158 , \61161 );
buf \U$61188 ( \61163 , \61162 );
buf \U$61189 ( \61164 , \61163 );
not \U$61190 ( \61165 , \61164 );
or \U$61191 ( \61166 , \61086 , \61165 );
buf \U$61192 ( \61167 , \61163 );
buf \U$61193 ( \61168 , \61084 );
or \U$61194 ( \61169 , \61167 , \61168 );
nand \U$61195 ( \61170 , \61166 , \61169 );
buf \U$61196 ( \61171 , \61170 );
buf \U$61197 ( \61172 , \61171 );
buf \U$61198 ( \61173 , \58200 );
buf \U$61199 ( \61174 , \60924 );
or \U$61200 ( \61175 , \61173 , \61174 );
buf \U$61201 ( \61176 , \12647 );
buf \U$61202 ( \61177 , \61110 );
not \U$61203 ( \61178 , \61177 );
buf \U$61204 ( \61179 , \61178 );
buf \U$61205 ( \61180 , \61179 );
or \U$61206 ( \61181 , \61176 , \61180 );
nand \U$61207 ( \61182 , \61175 , \61181 );
buf \U$61208 ( \61183 , \61182 );
buf \U$61209 ( \61184 , \61183 );
buf \U$61210 ( \61185 , \60966 );
not \U$61211 ( \61186 , \61185 );
buf \U$61212 ( \61187 , \14471 );
not \U$61213 ( \61188 , \61187 );
or \U$61214 ( \61189 , \61186 , \61188 );
buf \U$61215 ( \61190 , \60777 );
not \U$61216 ( \61191 , \61190 );
buf \U$61217 ( \61192 , \15793 );
nand \U$61218 ( \61193 , \61191 , \61192 );
buf \U$61219 ( \61194 , \61193 );
buf \U$61220 ( \61195 , \61194 );
nand \U$61221 ( \61196 , \61189 , \61195 );
buf \U$61222 ( \61197 , \61196 );
buf \U$61223 ( \61198 , \61197 );
xor \U$61224 ( \61199 , \61184 , \61198 );
xor \U$61225 ( \61200 , \60808 , \60829 );
buf \U$61226 ( \61201 , \61200 );
buf \U$61227 ( \61202 , \61201 );
and \U$61228 ( \61203 , \61199 , \61202 );
and \U$61229 ( \61204 , \61184 , \61198 );
or \U$61230 ( \61205 , \61203 , \61204 );
buf \U$61231 ( \61206 , \61205 );
buf \U$61232 ( \61207 , \61206 );
xor \U$61233 ( \61208 , \61172 , \61207 );
buf \U$61234 ( \61209 , \61208 );
buf \U$61235 ( \61210 , \61209 );
nand \U$61236 ( \61211 , \61042 , \61210 );
buf \U$61237 ( \61212 , \61211 );
buf \U$61238 ( \61213 , \61212 );
nand \U$61239 ( \61214 , \61039 , \61213 );
buf \U$61240 ( \61215 , \61214 );
buf \U$61241 ( \61216 , \61215 );
not \U$61242 ( \61217 , \61216 );
xor \U$61243 ( \61218 , \61047 , \61064 );
and \U$61244 ( \61219 , \61218 , \61082 );
and \U$61245 ( \61220 , \61047 , \61064 );
or \U$61246 ( \61221 , \61219 , \61220 );
buf \U$61247 ( \61222 , \61221 );
buf \U$61248 ( \61223 , \61222 );
not \U$61249 ( \61224 , \61223 );
buf \U$61250 ( \61225 , \61224 );
buf \U$61251 ( \61226 , \61225 );
not \U$61252 ( \61227 , \61226 );
buf \U$61253 ( \61228 , \61096 );
not \U$61254 ( \61229 , \61228 );
buf \U$61255 ( \61230 , \22350 );
not \U$61256 ( \61231 , \61230 );
or \U$61257 ( \61232 , \61229 , \61231 );
buf \U$61258 ( \61233 , \12937 );
buf \U$61259 ( \61234 , \60632 );
nand \U$61260 ( \61235 , \61233 , \61234 );
buf \U$61261 ( \61236 , \61235 );
buf \U$61262 ( \61237 , \61236 );
nand \U$61263 ( \61238 , \61232 , \61237 );
buf \U$61264 ( \61239 , \61238 );
buf \U$61265 ( \61240 , \61239 );
not \U$61266 ( \61241 , \61240 );
buf \U$61267 ( \61242 , RIc0d9400_64);
buf \U$61268 ( \61243 , RIc0dac60_116);
or \U$61269 ( \61244 , \61242 , \61243 );
buf \U$61270 ( \61245 , RIc0dacd8_117);
nand \U$61271 ( \61246 , \61244 , \61245 );
buf \U$61272 ( \61247 , \61246 );
buf \U$61273 ( \61248 , \61247 );
buf \U$61274 ( \61249 , RIc0d9400_64);
buf \U$61275 ( \61250 , RIc0dac60_116);
nand \U$61276 ( \61251 , \61249 , \61250 );
buf \U$61277 ( \61252 , \61251 );
buf \U$61278 ( \61253 , \61252 );
buf \U$61279 ( \61254 , RIc0dabe8_115);
nand \U$61280 ( \61255 , \61248 , \61253 , \61254 );
buf \U$61281 ( \61256 , \61255 );
buf \U$61282 ( \61257 , \61256 );
not \U$61283 ( \61258 , \61257 );
and \U$61284 ( \61259 , \61241 , \61258 );
buf \U$61285 ( \61260 , \61239 );
buf \U$61286 ( \61261 , \61256 );
and \U$61287 ( \61262 , \61260 , \61261 );
nor \U$61288 ( \61263 , \61259 , \61262 );
buf \U$61289 ( \61264 , \61263 );
buf \U$61290 ( \61265 , \61264 );
not \U$61291 ( \61266 , \61265 );
buf \U$61292 ( \61267 , \61266 );
buf \U$61293 ( \61268 , \61267 );
not \U$61294 ( \61269 , \61268 );
or \U$61295 ( \61270 , \61227 , \61269 );
buf \U$61296 ( \61271 , \61264 );
buf \U$61297 ( \61272 , \61222 );
nand \U$61298 ( \61273 , \61271 , \61272 );
buf \U$61299 ( \61274 , \61273 );
buf \U$61300 ( \61275 , \61274 );
nand \U$61301 ( \61276 , \61270 , \61275 );
buf \U$61302 ( \61277 , \61276 );
buf \U$61303 ( \61278 , \61277 );
buf \U$61304 ( \61279 , \61126 );
not \U$61305 ( \61280 , \61279 );
buf \U$61306 ( \61281 , \61102 );
not \U$61307 ( \61282 , \61281 );
or \U$61308 ( \61283 , \61280 , \61282 );
buf \U$61309 ( \61284 , \61129 );
not \U$61310 ( \61285 , \61284 );
buf \U$61311 ( \61286 , \61105 );
not \U$61312 ( \61287 , \61286 );
or \U$61313 ( \61288 , \61285 , \61287 );
buf \U$61314 ( \61289 , \61153 );
nand \U$61315 ( \61290 , \61288 , \61289 );
buf \U$61316 ( \61291 , \61290 );
buf \U$61317 ( \61292 , \61291 );
nand \U$61318 ( \61293 , \61283 , \61292 );
buf \U$61319 ( \61294 , \61293 );
buf \U$61320 ( \61295 , \61294 );
not \U$61321 ( \61296 , \61295 );
buf \U$61322 ( \61297 , \61296 );
buf \U$61323 ( \61298 , \61297 );
and \U$61324 ( \61299 , \61278 , \61298 );
not \U$61325 ( \61300 , \61278 );
buf \U$61326 ( \61301 , \61294 );
and \U$61327 ( \61302 , \61300 , \61301 );
nor \U$61328 ( \61303 , \61299 , \61302 );
buf \U$61329 ( \61304 , \61303 );
buf \U$61330 ( \61305 , \61304 );
buf \U$61331 ( \61306 , \61163 );
not \U$61332 ( \61307 , \61306 );
buf \U$61333 ( \61308 , \61307 );
buf \U$61334 ( \61309 , \61308 );
buf \U$61335 ( \61310 , \61084 );
or \U$61336 ( \61311 , \61309 , \61310 );
buf \U$61337 ( \61312 , \61206 );
nand \U$61338 ( \61313 , \61311 , \61312 );
buf \U$61339 ( \61314 , \61313 );
buf \U$61340 ( \61315 , \61314 );
buf \U$61341 ( \61316 , \61308 );
buf \U$61342 ( \61317 , \61084 );
nand \U$61343 ( \61318 , \61316 , \61317 );
buf \U$61344 ( \61319 , \61318 );
buf \U$61345 ( \61320 , \61319 );
nand \U$61346 ( \61321 , \61315 , \61320 );
buf \U$61347 ( \61322 , \61321 );
buf \U$61348 ( \61323 , \61322 );
not \U$61349 ( \61324 , \61323 );
buf \U$61350 ( \61325 , \61324 );
buf \U$61351 ( \61326 , \61325 );
xor \U$61352 ( \61327 , \61305 , \61326 );
buf \U$61353 ( \61328 , \61327 );
buf \U$61354 ( \61329 , \61328 );
not \U$61355 ( \61330 , \61329 );
buf \U$61356 ( \61331 , \61119 );
not \U$61357 ( \61332 , \61331 );
buf \U$61358 ( \61333 , \15609 );
not \U$61359 ( \61334 , \61333 );
or \U$61360 ( \61335 , \61332 , \61334 );
buf \U$61361 ( \61336 , \60677 );
buf \U$61362 ( \61337 , RIc0db200_128);
nand \U$61363 ( \61338 , \61336 , \61337 );
buf \U$61364 ( \61339 , \61338 );
buf \U$61365 ( \61340 , \61339 );
nand \U$61366 ( \61341 , \61335 , \61340 );
buf \U$61367 ( \61342 , \61341 );
buf \U$61368 ( \61343 , \61342 );
buf \U$61369 ( \61344 , \61075 );
not \U$61370 ( \61345 , \61344 );
buf \U$61371 ( \61346 , \13949 );
not \U$61372 ( \61347 , \61346 );
or \U$61373 ( \61348 , \61345 , \61347 );
buf \U$61374 ( \61349 , \13953 );
buf \U$61375 ( \61350 , \60689 );
nand \U$61376 ( \61351 , \61349 , \61350 );
buf \U$61377 ( \61352 , \61351 );
buf \U$61378 ( \61353 , \61352 );
nand \U$61379 ( \61354 , \61348 , \61353 );
buf \U$61380 ( \61355 , \61354 );
buf \U$61381 ( \61356 , \61355 );
xor \U$61382 ( \61357 , \61343 , \61356 );
buf \U$61383 ( \61358 , \61147 );
not \U$61384 ( \61359 , \61358 );
buf \U$61385 ( \61360 , \47037 );
not \U$61386 ( \61361 , \61360 );
or \U$61387 ( \61362 , \61359 , \61361 );
buf \U$61388 ( \61363 , \60651 );
not \U$61389 ( \61364 , \61363 );
buf \U$61390 ( \61365 , \16692 );
nand \U$61391 ( \61366 , \61364 , \61365 );
buf \U$61392 ( \61367 , \61366 );
buf \U$61393 ( \61368 , \61367 );
nand \U$61394 ( \61369 , \61362 , \61368 );
buf \U$61395 ( \61370 , \61369 );
buf \U$61396 ( \61371 , \61370 );
xnor \U$61397 ( \61372 , \61357 , \61371 );
buf \U$61398 ( \61373 , \61372 );
buf \U$61399 ( \61374 , \61373 );
not \U$61400 ( \61375 , \61374 );
buf \U$61401 ( \61376 , \61375 );
buf \U$61402 ( \61377 , \61376 );
not \U$61403 ( \61378 , \61377 );
buf \U$61404 ( \61379 , \60784 );
not \U$61405 ( \61380 , \61379 );
buf \U$61406 ( \61381 , \44382 );
not \U$61407 ( \61382 , \61381 );
or \U$61408 ( \61383 , \61380 , \61382 );
buf \U$61409 ( \61384 , \15793 );
buf \U$61410 ( \61385 , \60708 );
nand \U$61411 ( \61386 , \61384 , \61385 );
buf \U$61412 ( \61387 , \61386 );
buf \U$61413 ( \61388 , \61387 );
nand \U$61414 ( \61389 , \61383 , \61388 );
buf \U$61415 ( \61390 , \61389 );
buf \U$61416 ( \61391 , \61390 );
buf \U$61417 ( \61392 , \61057 );
not \U$61418 ( \61393 , \61392 );
buf \U$61419 ( \61394 , \19487 );
not \U$61420 ( \61395 , \61394 );
or \U$61421 ( \61396 , \61393 , \61395 );
buf \U$61422 ( \61397 , \13314 );
buf \U$61423 ( \61398 , RIc0d90b8_57);
buf \U$61424 ( \61399 , RIc0daeb8_121);
xor \U$61425 ( \61400 , \61398 , \61399 );
buf \U$61426 ( \61401 , \61400 );
buf \U$61427 ( \61402 , \61401 );
nand \U$61428 ( \61403 , \61397 , \61402 );
buf \U$61429 ( \61404 , \61403 );
buf \U$61430 ( \61405 , \61404 );
nand \U$61431 ( \61406 , \61396 , \61405 );
buf \U$61432 ( \61407 , \61406 );
buf \U$61433 ( \61408 , \61407 );
xor \U$61434 ( \61409 , \61391 , \61408 );
buf \U$61435 ( \61410 , \14681 );
buf \U$61436 ( \61411 , \12387 );
buf \U$61437 ( \61412 , RIc0d9400_64);
and \U$61438 ( \61413 , \61411 , \61412 );
buf \U$61439 ( \61414 , \43843 );
buf \U$61440 ( \61415 , RIc0dabe8_115);
and \U$61441 ( \61416 , \61414 , \61415 );
nor \U$61442 ( \61417 , \61413 , \61416 );
buf \U$61443 ( \61418 , \61417 );
buf \U$61444 ( \61419 , \61418 );
or \U$61445 ( \61420 , \61410 , \61419 );
buf \U$61446 ( \61421 , \29865 );
buf \U$61447 ( \61422 , RIc0d9388_63);
buf \U$61448 ( \61423 , RIc0dabe8_115);
xor \U$61449 ( \61424 , \61422 , \61423 );
buf \U$61450 ( \61425 , \61424 );
buf \U$61451 ( \61426 , \61425 );
not \U$61452 ( \61427 , \61426 );
buf \U$61453 ( \61428 , \61427 );
buf \U$61454 ( \61429 , \61428 );
or \U$61455 ( \61430 , \61421 , \61429 );
nand \U$61456 ( \61431 , \61420 , \61430 );
buf \U$61457 ( \61432 , \61431 );
buf \U$61458 ( \61433 , \61432 );
xor \U$61459 ( \61434 , \61409 , \61433 );
buf \U$61460 ( \61435 , \61434 );
buf \U$61461 ( \61436 , \61435 );
not \U$61462 ( \61437 , \61436 );
buf \U$61463 ( \61438 , \61437 );
buf \U$61464 ( \61439 , \61438 );
not \U$61465 ( \61440 , \61439 );
or \U$61466 ( \61441 , \61378 , \61440 );
buf \U$61467 ( \61442 , \61435 );
buf \U$61468 ( \61443 , \61373 );
nand \U$61469 ( \61444 , \61442 , \61443 );
buf \U$61470 ( \61445 , \61444 );
buf \U$61471 ( \61446 , \61445 );
nand \U$61472 ( \61447 , \61441 , \61446 );
buf \U$61473 ( \61448 , \61447 );
buf \U$61474 ( \61449 , \61448 );
xor \U$61475 ( \61450 , \60792 , \60832 );
and \U$61476 ( \61451 , \61450 , \60905 );
and \U$61477 ( \61452 , \60792 , \60832 );
or \U$61478 ( \61453 , \61451 , \61452 );
buf \U$61479 ( \61454 , \61453 );
buf \U$61480 ( \61455 , \61454 );
xnor \U$61481 ( \61456 , \61449 , \61455 );
buf \U$61482 ( \61457 , \61456 );
buf \U$61483 ( \61458 , \61457 );
not \U$61484 ( \61459 , \61458 );
and \U$61485 ( \61460 , \61330 , \61459 );
buf \U$61486 ( \61461 , \61328 );
buf \U$61487 ( \61462 , \61457 );
and \U$61488 ( \61463 , \61461 , \61462 );
nor \U$61489 ( \61464 , \61460 , \61463 );
buf \U$61490 ( \61465 , \61464 );
buf \U$61491 ( \61466 , \61465 );
nand \U$61492 ( \61467 , \61217 , \61466 );
buf \U$61493 ( \61468 , \61467 );
buf \U$61494 ( \61469 , \61468 );
xor \U$61495 ( \61470 , \61184 , \61198 );
xor \U$61496 ( \61471 , \61470 , \61202 );
buf \U$61497 ( \61472 , \61471 );
buf \U$61498 ( \61473 , \61472 );
xor \U$61499 ( \61474 , \60979 , \61027 );
xor \U$61500 ( \61475 , \61474 , \61032 );
buf \U$61501 ( \61476 , \61475 );
buf \U$61502 ( \61477 , \61476 );
or \U$61503 ( \61478 , \61473 , \61477 );
buf \U$61504 ( \61479 , RIc0d9400_64);
buf \U$61505 ( \61480 , RIc0dae40_120);
or \U$61506 ( \61481 , \61479 , \61480 );
buf \U$61507 ( \61482 , RIc0daeb8_121);
nand \U$61508 ( \61483 , \61481 , \61482 );
buf \U$61509 ( \61484 , \61483 );
buf \U$61510 ( \61485 , \61484 );
buf \U$61511 ( \61486 , RIc0d9400_64);
buf \U$61512 ( \61487 , RIc0dae40_120);
nand \U$61513 ( \61488 , \61486 , \61487 );
buf \U$61514 ( \61489 , \61488 );
buf \U$61515 ( \61490 , \61489 );
buf \U$61516 ( \61491 , RIc0dadc8_119);
and \U$61517 ( \61492 , \61485 , \61490 , \61491 );
buf \U$61518 ( \61493 , \61492 );
buf \U$61519 ( \61494 , \61493 );
buf \U$61520 ( \61495 , RIc0daeb8_121);
buf \U$61521 ( \61496 , RIc0d9310_62);
and \U$61522 ( \61497 , \61495 , \61496 );
not \U$61523 ( \61498 , \61495 );
buf \U$61524 ( \61499 , \60362 );
and \U$61525 ( \61500 , \61498 , \61499 );
nor \U$61526 ( \61501 , \61497 , \61500 );
buf \U$61527 ( \61502 , \61501 );
buf \U$61528 ( \61503 , \61502 );
not \U$61529 ( \61504 , \61503 );
buf \U$61530 ( \61505 , \13310 );
not \U$61531 ( \61506 , \61505 );
or \U$61532 ( \61507 , \61504 , \61506 );
buf \U$61533 ( \61508 , \12975 );
buf \U$61534 ( \61509 , \60988 );
nand \U$61535 ( \61510 , \61508 , \61509 );
buf \U$61536 ( \61511 , \61510 );
buf \U$61537 ( \61512 , \61511 );
nand \U$61538 ( \61513 , \61507 , \61512 );
buf \U$61539 ( \61514 , \61513 );
buf \U$61540 ( \61515 , \61514 );
and \U$61541 ( \61516 , \61494 , \61515 );
buf \U$61542 ( \61517 , \61516 );
buf \U$61543 ( \61518 , \61517 );
xor \U$61544 ( \61519 , \60984 , \61001 );
xor \U$61545 ( \61520 , \61519 , \61022 );
buf \U$61546 ( \61521 , \61520 );
buf \U$61547 ( \61522 , \61521 );
xor \U$61548 ( \61523 , \61518 , \61522 );
xor \U$61549 ( \61524 , RIc0db098_125, RIc0d9130_58);
buf \U$61550 ( \61525 , \61524 );
not \U$61551 ( \61526 , \61525 );
buf \U$61552 ( \61527 , \13461 );
not \U$61553 ( \61528 , \61527 );
or \U$61554 ( \61529 , \61526 , \61528 );
buf \U$61555 ( \61530 , \13465 );
buf \U$61556 ( \61531 , \60956 );
nand \U$61557 ( \61532 , \61530 , \61531 );
buf \U$61558 ( \61533 , \61532 );
buf \U$61559 ( \61534 , \61533 );
nand \U$61560 ( \61535 , \61529 , \61534 );
buf \U$61561 ( \61536 , \61535 );
buf \U$61562 ( \61537 , \61536 );
not \U$61563 ( \61538 , \61537 );
buf \U$61564 ( \61539 , RIc0d9040_56);
buf \U$61565 ( \61540 , RIc0db188_127);
xor \U$61566 ( \61541 , \61539 , \61540 );
buf \U$61567 ( \61542 , \61541 );
buf \U$61568 ( \61543 , \61542 );
not \U$61569 ( \61544 , \61543 );
buf \U$61570 ( \61545 , \46813 );
not \U$61571 ( \61546 , \61545 );
or \U$61572 ( \61547 , \61544 , \61546 );
buf \U$61573 ( \61548 , \60914 );
buf \U$61574 ( \61549 , RIc0db200_128);
nand \U$61575 ( \61550 , \61548 , \61549 );
buf \U$61576 ( \61551 , \61550 );
buf \U$61577 ( \61552 , \61551 );
nand \U$61578 ( \61553 , \61547 , \61552 );
buf \U$61579 ( \61554 , \61553 );
buf \U$61580 ( \61555 , \61554 );
not \U$61581 ( \61556 , \61555 );
or \U$61582 ( \61557 , \61538 , \61556 );
buf \U$61583 ( \61558 , \61554 );
buf \U$61584 ( \61559 , \61536 );
or \U$61585 ( \61560 , \61558 , \61559 );
buf \U$61586 ( \61561 , RIc0d9220_60);
buf \U$61587 ( \61562 , RIc0dafa8_123);
xor \U$61588 ( \61563 , \61561 , \61562 );
buf \U$61589 ( \61564 , \61563 );
buf \U$61590 ( \61565 , \61564 );
not \U$61591 ( \61566 , \61565 );
buf \U$61592 ( \61567 , \45570 );
not \U$61593 ( \61568 , \61567 );
or \U$61594 ( \61569 , \61566 , \61568 );
buf \U$61595 ( \61570 , \16692 );
buf \U$61596 ( \61571 , \60934 );
nand \U$61597 ( \61572 , \61570 , \61571 );
buf \U$61598 ( \61573 , \61572 );
buf \U$61599 ( \61574 , \61573 );
nand \U$61600 ( \61575 , \61569 , \61574 );
buf \U$61601 ( \61576 , \61575 );
buf \U$61602 ( \61577 , \61576 );
nand \U$61603 ( \61578 , \61560 , \61577 );
buf \U$61604 ( \61579 , \61578 );
buf \U$61605 ( \61580 , \61579 );
nand \U$61606 ( \61581 , \61557 , \61580 );
buf \U$61607 ( \61582 , \61581 );
buf \U$61608 ( \61583 , \61582 );
and \U$61609 ( \61584 , \61523 , \61583 );
and \U$61610 ( \61585 , \61518 , \61522 );
or \U$61611 ( \61586 , \61584 , \61585 );
buf \U$61612 ( \61587 , \61586 );
buf \U$61613 ( \61588 , \61587 );
nand \U$61614 ( \61589 , \61478 , \61588 );
buf \U$61615 ( \61590 , \61589 );
buf \U$61616 ( \61591 , \61590 );
buf \U$61617 ( \61592 , \61476 );
buf \U$61618 ( \61593 , \61472 );
nand \U$61619 ( \61594 , \61592 , \61593 );
buf \U$61620 ( \61595 , \61594 );
buf \U$61621 ( \61596 , \61595 );
nand \U$61622 ( \61597 , \61591 , \61596 );
buf \U$61623 ( \61598 , \61597 );
buf \U$61624 ( \61599 , \61598 );
not \U$61625 ( \61600 , \61599 );
buf \U$61626 ( \61601 , \60907 );
not \U$61627 ( \61602 , \61601 );
buf \U$61628 ( \61603 , \61036 );
not \U$61629 ( \61604 , \61603 );
buf \U$61630 ( \61605 , \61604 );
buf \U$61631 ( \61606 , \61605 );
not \U$61632 ( \61607 , \61606 );
or \U$61633 ( \61608 , \61602 , \61607 );
buf \U$61634 ( \61609 , \60907 );
not \U$61635 ( \61610 , \61609 );
buf \U$61636 ( \61611 , \61036 );
nand \U$61637 ( \61612 , \61610 , \61611 );
buf \U$61638 ( \61613 , \61612 );
buf \U$61639 ( \61614 , \61613 );
nand \U$61640 ( \61615 , \61608 , \61614 );
buf \U$61641 ( \61616 , \61615 );
buf \U$61642 ( \61617 , \61616 );
buf \U$61643 ( \61618 , \61209 );
xnor \U$61644 ( \61619 , \61617 , \61618 );
buf \U$61645 ( \61620 , \61619 );
buf \U$61646 ( \61621 , \61620 );
nor \U$61647 ( \61622 , \61600 , \61621 );
buf \U$61648 ( \61623 , \61622 );
buf \U$61649 ( \61624 , \61623 );
nand \U$61650 ( \61625 , \61469 , \61624 );
buf \U$61651 ( \61626 , \61625 );
buf \U$61652 ( \61627 , \61626 );
buf \U$61653 ( \61628 , \61465 );
not \U$61654 ( \61629 , \61628 );
buf \U$61655 ( \61630 , \61215 );
nand \U$61656 ( \61631 , \61629 , \61630 );
buf \U$61657 ( \61632 , \61631 );
buf \U$61658 ( \61633 , \61632 );
nand \U$61659 ( \61634 , \61627 , \61633 );
buf \U$61660 ( \61635 , \61634 );
buf \U$61661 ( \61636 , \61635 );
not \U$61662 ( \61637 , \61636 );
xor \U$61663 ( \61638 , \60628 , \60645 );
xor \U$61664 ( \61639 , \61638 , \60659 );
buf \U$61665 ( \61640 , \61639 );
buf \U$61666 ( \61641 , \61640 );
xor \U$61667 ( \61642 , \61391 , \61408 );
and \U$61668 ( \61643 , \61642 , \61433 );
and \U$61669 ( \61644 , \61391 , \61408 );
or \U$61670 ( \61645 , \61643 , \61644 );
buf \U$61671 ( \61646 , \61645 );
buf \U$61672 ( \61647 , \61646 );
xor \U$61673 ( \61648 , \61641 , \61647 );
buf \U$61674 ( \61649 , \61342 );
not \U$61675 ( \61650 , \61649 );
buf \U$61676 ( \61651 , \61370 );
not \U$61677 ( \61652 , \61651 );
or \U$61678 ( \61653 , \61650 , \61652 );
buf \U$61679 ( \61654 , \61370 );
buf \U$61680 ( \61655 , \61342 );
or \U$61681 ( \61656 , \61654 , \61655 );
buf \U$61682 ( \61657 , \61355 );
nand \U$61683 ( \61658 , \61656 , \61657 );
buf \U$61684 ( \61659 , \61658 );
buf \U$61685 ( \61660 , \61659 );
nand \U$61686 ( \61661 , \61653 , \61660 );
buf \U$61687 ( \61662 , \61661 );
buf \U$61688 ( \61663 , \61662 );
xor \U$61689 ( \61664 , \61648 , \61663 );
buf \U$61690 ( \61665 , \61664 );
xor \U$61691 ( \61666 , \60685 , \60703 );
xor \U$61692 ( \61667 , \61666 , \60721 );
buf \U$61693 ( \61668 , \61667 );
buf \U$61694 ( \61669 , \61668 );
buf \U$61695 ( \61670 , \61425 );
not \U$61696 ( \61671 , \61670 );
buf \U$61697 ( \61672 , \46873 );
not \U$61698 ( \61673 , \61672 );
or \U$61699 ( \61674 , \61671 , \61673 );
buf \U$61700 ( \61675 , \12303 );
buf \U$61701 ( \61676 , \60366 );
nand \U$61702 ( \61677 , \61675 , \61676 );
buf \U$61703 ( \61678 , \61677 );
buf \U$61704 ( \61679 , \61678 );
nand \U$61705 ( \61680 , \61674 , \61679 );
buf \U$61706 ( \61681 , \61680 );
buf \U$61707 ( \61682 , \61681 );
buf \U$61708 ( \61683 , \61401 );
not \U$61709 ( \61684 , \61683 );
buf \U$61710 ( \61685 , \16382 );
not \U$61711 ( \61686 , \61685 );
or \U$61712 ( \61687 , \61684 , \61686 );
buf \U$61713 ( \61688 , \13314 );
buf \U$61714 ( \61689 , \60443 );
nand \U$61715 ( \61690 , \61688 , \61689 );
buf \U$61716 ( \61691 , \61690 );
buf \U$61717 ( \61692 , \61691 );
nand \U$61718 ( \61693 , \61687 , \61692 );
buf \U$61719 ( \61694 , \61693 );
buf \U$61720 ( \61695 , \61694 );
xor \U$61721 ( \61696 , \61682 , \61695 );
buf \U$61722 ( \61697 , \61239 );
buf \U$61723 ( \61698 , \61256 );
not \U$61724 ( \61699 , \61698 );
buf \U$61725 ( \61700 , \61699 );
buf \U$61726 ( \61701 , \61700 );
and \U$61727 ( \61702 , \61697 , \61701 );
buf \U$61728 ( \61703 , \61702 );
buf \U$61729 ( \61704 , \61703 );
xor \U$61730 ( \61705 , \61696 , \61704 );
buf \U$61731 ( \61706 , \61705 );
buf \U$61732 ( \61707 , \61706 );
xor \U$61733 ( \61708 , \61669 , \61707 );
buf \U$61734 ( \61709 , \61267 );
not \U$61735 ( \61710 , \61709 );
buf \U$61736 ( \61711 , \61294 );
not \U$61737 ( \61712 , \61711 );
or \U$61738 ( \61713 , \61710 , \61712 );
buf \U$61739 ( \61714 , \61294 );
buf \U$61740 ( \61715 , \61267 );
or \U$61741 ( \61716 , \61714 , \61715 );
buf \U$61742 ( \61717 , \61222 );
nand \U$61743 ( \61718 , \61716 , \61717 );
buf \U$61744 ( \61719 , \61718 );
buf \U$61745 ( \61720 , \61719 );
nand \U$61746 ( \61721 , \61713 , \61720 );
buf \U$61747 ( \61722 , \61721 );
buf \U$61748 ( \61723 , \61722 );
xor \U$61749 ( \61724 , \61708 , \61723 );
buf \U$61750 ( \61725 , \61724 );
xor \U$61751 ( \61726 , \61665 , \61725 );
buf \U$61752 ( \61727 , \61726 );
buf \U$61753 ( \61728 , \61376 );
not \U$61754 ( \61729 , \61728 );
buf \U$61755 ( \61730 , \61435 );
not \U$61756 ( \61731 , \61730 );
or \U$61757 ( \61732 , \61729 , \61731 );
buf \U$61758 ( \61733 , \61454 );
buf \U$61759 ( \61734 , \61438 );
buf \U$61760 ( \61735 , \61373 );
nand \U$61761 ( \61736 , \61734 , \61735 );
buf \U$61762 ( \61737 , \61736 );
buf \U$61763 ( \61738 , \61737 );
nand \U$61764 ( \61739 , \61733 , \61738 );
buf \U$61765 ( \61740 , \61739 );
buf \U$61766 ( \61741 , \61740 );
nand \U$61767 ( \61742 , \61732 , \61741 );
buf \U$61768 ( \61743 , \61742 );
buf \U$61769 ( \61744 , \61743 );
xnor \U$61770 ( \61745 , \61727 , \61744 );
buf \U$61771 ( \61746 , \61745 );
buf \U$61772 ( \61747 , \61746 );
buf \U$61773 ( \61748 , \61322 );
not \U$61774 ( \61749 , \61748 );
buf \U$61775 ( \61750 , \61304 );
not \U$61776 ( \61751 , \61750 );
buf \U$61777 ( \61752 , \61751 );
buf \U$61778 ( \61753 , \61752 );
not \U$61779 ( \61754 , \61753 );
or \U$61780 ( \61755 , \61749 , \61754 );
and \U$61781 ( \61756 , \61305 , \61326 );
buf \U$61782 ( \61757 , \61756 );
or \U$61783 ( \61758 , \61757 , \61457 );
buf \U$61784 ( \61759 , \61758 );
nand \U$61785 ( \61760 , \61755 , \61759 );
buf \U$61786 ( \61761 , \61760 );
buf \U$61787 ( \61762 , \61761 );
not \U$61788 ( \61763 , \61762 );
buf \U$61789 ( \61764 , \61763 );
buf \U$61790 ( \61765 , \61764 );
nand \U$61791 ( \61766 , \61747 , \61765 );
buf \U$61792 ( \61767 , \61766 );
buf \U$61793 ( \61768 , \61767 );
not \U$61794 ( \61769 , \61768 );
or \U$61795 ( \61770 , \61637 , \61769 );
buf \U$61796 ( \61771 , \61746 );
not \U$61797 ( \61772 , \61771 );
buf \U$61798 ( \61773 , \61761 );
nand \U$61799 ( \61774 , \61772 , \61773 );
buf \U$61800 ( \61775 , \61774 );
buf \U$61801 ( \61776 , \61775 );
nand \U$61802 ( \61777 , \61770 , \61776 );
buf \U$61803 ( \61778 , \61777 );
buf \U$61804 ( \61779 , \61778 );
buf \U$61805 ( \61780 , \61665 );
not \U$61806 ( \61781 , \61780 );
buf \U$61807 ( \61782 , \61743 );
not \U$61808 ( \61783 , \61782 );
or \U$61809 ( \61784 , \61781 , \61783 );
buf \U$61810 ( \61785 , \61743 );
buf \U$61811 ( \61786 , \61665 );
or \U$61812 ( \61787 , \61785 , \61786 );
buf \U$61813 ( \61788 , \61725 );
nand \U$61814 ( \61789 , \61787 , \61788 );
buf \U$61815 ( \61790 , \61789 );
buf \U$61816 ( \61791 , \61790 );
nand \U$61817 ( \61792 , \61784 , \61791 );
buf \U$61818 ( \61793 , \61792 );
buf \U$61819 ( \61794 , \61793 );
not \U$61820 ( \61795 , \61794 );
xor \U$61821 ( \61796 , \61682 , \61695 );
and \U$61822 ( \61797 , \61796 , \61704 );
and \U$61823 ( \61798 , \61682 , \61695 );
or \U$61824 ( \61799 , \61797 , \61798 );
buf \U$61825 ( \61800 , \61799 );
buf \U$61826 ( \61801 , \60613 );
buf \U$61827 ( \61802 , \60617 );
xor \U$61828 ( \61803 , \61801 , \61802 );
buf \U$61829 ( \61804 , \60663 );
xnor \U$61830 ( \61805 , \61803 , \61804 );
buf \U$61831 ( \61806 , \61805 );
xor \U$61832 ( \61807 , \61800 , \61806 );
xor \U$61833 ( \61808 , \61641 , \61647 );
and \U$61834 ( \61809 , \61808 , \61663 );
and \U$61835 ( \61810 , \61641 , \61647 );
or \U$61836 ( \61811 , \61809 , \61810 );
buf \U$61837 ( \61812 , \61811 );
xor \U$61838 ( \61813 , \61807 , \61812 );
buf \U$61839 ( \61814 , \61813 );
not \U$61840 ( \61815 , \61814 );
xor \U$61841 ( \61816 , \60725 , \60730 );
xnor \U$61842 ( \61817 , \61816 , \60739 );
buf \U$61843 ( \61818 , \61817 );
not \U$61844 ( \61819 , \61818 );
xor \U$61845 ( \61820 , \61669 , \61707 );
and \U$61846 ( \61821 , \61820 , \61723 );
and \U$61847 ( \61822 , \61669 , \61707 );
or \U$61848 ( \61823 , \61821 , \61822 );
buf \U$61849 ( \61824 , \61823 );
buf \U$61850 ( \61825 , \61824 );
not \U$61851 ( \61826 , \61825 );
or \U$61852 ( \61827 , \61819 , \61826 );
buf \U$61853 ( \61828 , \61824 );
buf \U$61854 ( \61829 , \61817 );
or \U$61855 ( \61830 , \61828 , \61829 );
nand \U$61856 ( \61831 , \61827 , \61830 );
buf \U$61857 ( \61832 , \61831 );
buf \U$61858 ( \61833 , \61832 );
not \U$61859 ( \61834 , \61833 );
and \U$61860 ( \61835 , \61815 , \61834 );
buf \U$61861 ( \61836 , \61813 );
buf \U$61862 ( \61837 , \61832 );
and \U$61863 ( \61838 , \61836 , \61837 );
nor \U$61864 ( \61839 , \61835 , \61838 );
buf \U$61865 ( \61840 , \61839 );
buf \U$61866 ( \61841 , \61840 );
nand \U$61867 ( \61842 , \61795 , \61841 );
buf \U$61868 ( \61843 , \61842 );
buf \U$61869 ( \61844 , \61843 );
nand \U$61870 ( \61845 , \61779 , \61844 );
buf \U$61871 ( \61846 , \61845 );
buf \U$61872 ( \61847 , \61846 );
buf \U$61873 ( \61848 , \60910 );
xnor \U$61874 ( \61849 , RIc0db188_127, RIc0d90b8_57);
buf \U$61875 ( \61850 , \61849 );
or \U$61876 ( \61851 , \61848 , \61850 );
buf \U$61877 ( \61852 , \12647 );
buf \U$61878 ( \61853 , \61542 );
not \U$61879 ( \61854 , \61853 );
buf \U$61880 ( \61855 , \61854 );
buf \U$61881 ( \61856 , \61855 );
or \U$61882 ( \61857 , \61852 , \61856 );
nand \U$61883 ( \61858 , \61851 , \61857 );
buf \U$61884 ( \61859 , \61858 );
buf \U$61885 ( \61860 , \61859 );
buf \U$61886 ( \61861 , \13005 );
buf \U$61887 ( \61862 , RIc0d9400_64);
and \U$61888 ( \61863 , \61861 , \61862 );
buf \U$61889 ( \61864 , \61863 );
buf \U$61890 ( \61865 , \61864 );
xor \U$61891 ( \61866 , \61860 , \61865 );
buf \U$61892 ( \61867 , RIc0d9298_61);
buf \U$61893 ( \61868 , RIc0dafa8_123);
xor \U$61894 ( \61869 , \61867 , \61868 );
buf \U$61895 ( \61870 , \61869 );
buf \U$61896 ( \61871 , \61870 );
not \U$61897 ( \61872 , \61871 );
buf \U$61898 ( \61873 , \45570 );
not \U$61899 ( \61874 , \61873 );
or \U$61900 ( \61875 , \61872 , \61874 );
buf \U$61901 ( \61876 , \14278 );
buf \U$61902 ( \61877 , \61564 );
nand \U$61903 ( \61878 , \61876 , \61877 );
buf \U$61904 ( \61879 , \61878 );
buf \U$61905 ( \61880 , \61879 );
nand \U$61906 ( \61881 , \61875 , \61880 );
buf \U$61907 ( \61882 , \61881 );
buf \U$61908 ( \61883 , \61882 );
xor \U$61909 ( \61884 , \61866 , \61883 );
buf \U$61910 ( \61885 , \61884 );
buf \U$61911 ( \61886 , \61885 );
not \U$61912 ( \61887 , \58522 );
buf \U$61913 ( \61888 , \61887 );
buf \U$61914 ( \61889 , RIc0db188_127);
buf \U$61915 ( \61890 , RIc0d9130_58);
xnor \U$61916 ( \61891 , \61889 , \61890 );
buf \U$61917 ( \61892 , \61891 );
buf \U$61918 ( \61893 , \61892 );
or \U$61919 ( \61894 , \61888 , \61893 );
buf \U$61920 ( \61895 , \61849 );
buf \U$61921 ( \61896 , \12647 );
or \U$61922 ( \61897 , \61895 , \61896 );
nand \U$61923 ( \61898 , \61894 , \61897 );
buf \U$61924 ( \61899 , \61898 );
buf \U$61925 ( \61900 , \61899 );
buf \U$61926 ( \61901 , RIc0d9220_60);
buf \U$61927 ( \61902 , RIc0db098_125);
xor \U$61928 ( \61903 , \61901 , \61902 );
buf \U$61929 ( \61904 , \61903 );
buf \U$61930 ( \61905 , \61904 );
not \U$61931 ( \61906 , \61905 );
buf \U$61932 ( \61907 , \13461 );
not \U$61933 ( \61908 , \61907 );
or \U$61934 ( \61909 , \61906 , \61908 );
buf \U$61935 ( \61910 , RIc0d91a8_59);
buf \U$61936 ( \61911 , RIc0db098_125);
xnor \U$61937 ( \61912 , \61910 , \61911 );
buf \U$61938 ( \61913 , \61912 );
buf \U$61939 ( \61914 , \61913 );
not \U$61940 ( \61915 , \61914 );
buf \U$61941 ( \61916 , \15793 );
nand \U$61942 ( \61917 , \61915 , \61916 );
buf \U$61943 ( \61918 , \61917 );
buf \U$61944 ( \61919 , \61918 );
nand \U$61945 ( \61920 , \61909 , \61919 );
buf \U$61946 ( \61921 , \61920 );
buf \U$61947 ( \61922 , \61921 );
xor \U$61948 ( \61923 , \61900 , \61922 );
buf \U$61949 ( \61924 , \49672 );
buf \U$61950 ( \61925 , \13166 );
buf \U$61951 ( \61926 , RIc0d9400_64);
and \U$61952 ( \61927 , \61925 , \61926 );
buf \U$61953 ( \61928 , \43843 );
buf \U$61954 ( \61929 , RIc0daeb8_121);
and \U$61955 ( \61930 , \61928 , \61929 );
nor \U$61956 ( \61931 , \61927 , \61930 );
buf \U$61957 ( \61932 , \61931 );
buf \U$61958 ( \61933 , \61932 );
or \U$61959 ( \61934 , \61924 , \61933 );
buf \U$61960 ( \61935 , \27558 );
buf \U$61961 ( \61936 , RIc0d9388_63);
buf \U$61962 ( \61937 , RIc0daeb8_121);
xor \U$61963 ( \61938 , \61936 , \61937 );
buf \U$61964 ( \61939 , \61938 );
buf \U$61965 ( \61940 , \61939 );
not \U$61966 ( \61941 , \61940 );
buf \U$61967 ( \61942 , \61941 );
buf \U$61968 ( \61943 , \61942 );
or \U$61969 ( \61944 , \61935 , \61943 );
nand \U$61970 ( \61945 , \61934 , \61944 );
buf \U$61971 ( \61946 , \61945 );
buf \U$61972 ( \61947 , \61946 );
and \U$61973 ( \61948 , \61923 , \61947 );
and \U$61974 ( \61949 , \61900 , \61922 );
or \U$61975 ( \61950 , \61948 , \61949 );
buf \U$61976 ( \61951 , \61950 );
buf \U$61977 ( \61952 , \61951 );
xor \U$61978 ( \61953 , \61886 , \61952 );
buf \U$61979 ( \61954 , \61939 );
not \U$61980 ( \61955 , \61954 );
buf \U$61981 ( \61956 , \13310 );
not \U$61982 ( \61957 , \61956 );
or \U$61983 ( \61958 , \61955 , \61957 );
buf \U$61984 ( \61959 , \16386 );
buf \U$61985 ( \61960 , \61502 );
nand \U$61986 ( \61961 , \61959 , \61960 );
buf \U$61987 ( \61962 , \61961 );
buf \U$61988 ( \61963 , \61962 );
nand \U$61989 ( \61964 , \61958 , \61963 );
buf \U$61990 ( \61965 , \61964 );
buf \U$61991 ( \61966 , \61965 );
not \U$61992 ( \61967 , \61966 );
not \U$61993 ( \61968 , \14468 );
not \U$61994 ( \61969 , \61913 );
and \U$61995 ( \61970 , \61968 , \61969 );
and \U$61996 ( \61971 , \13465 , \61524 );
nor \U$61997 ( \61972 , \61970 , \61971 );
buf \U$61998 ( \61973 , \61972 );
not \U$61999 ( \61974 , \61973 );
or \U$62000 ( \61975 , \61967 , \61974 );
buf \U$62001 ( \61976 , \61972 );
buf \U$62002 ( \61977 , \61965 );
or \U$62003 ( \61978 , \61976 , \61977 );
nand \U$62004 ( \61979 , \61975 , \61978 );
buf \U$62005 ( \61980 , \61979 );
buf \U$62006 ( \61981 , \61980 );
buf \U$62007 ( \61982 , RIc0d9310_62);
buf \U$62008 ( \61983 , RIc0dafa8_123);
xor \U$62009 ( \61984 , \61982 , \61983 );
buf \U$62010 ( \61985 , \61984 );
buf \U$62011 ( \61986 , \61985 );
not \U$62012 ( \61987 , \61986 );
buf \U$62013 ( \61988 , \47037 );
not \U$62014 ( \61989 , \61988 );
or \U$62015 ( \61990 , \61987 , \61989 );
buf \U$62016 ( \61991 , \16692 );
buf \U$62017 ( \61992 , \61870 );
nand \U$62018 ( \61993 , \61991 , \61992 );
buf \U$62019 ( \61994 , \61993 );
buf \U$62020 ( \61995 , \61994 );
nand \U$62021 ( \61996 , \61990 , \61995 );
buf \U$62022 ( \61997 , \61996 );
buf \U$62023 ( \61998 , \61997 );
buf \U$62024 ( \61999 , RIc0d9400_64);
buf \U$62025 ( \62000 , RIc0daf30_122);
or \U$62026 ( \62001 , \61999 , \62000 );
buf \U$62027 ( \62002 , RIc0dafa8_123);
nand \U$62028 ( \62003 , \62001 , \62002 );
buf \U$62029 ( \62004 , \62003 );
buf \U$62030 ( \62005 , \62004 );
buf \U$62031 ( \62006 , RIc0d9400_64);
buf \U$62032 ( \62007 , RIc0daf30_122);
nand \U$62033 ( \62008 , \62006 , \62007 );
buf \U$62034 ( \62009 , \62008 );
buf \U$62035 ( \62010 , \62009 );
buf \U$62036 ( \62011 , RIc0daeb8_121);
and \U$62037 ( \62012 , \62005 , \62010 , \62011 );
buf \U$62038 ( \62013 , \62012 );
buf \U$62039 ( \62014 , \62013 );
nand \U$62040 ( \62015 , \61998 , \62014 );
buf \U$62041 ( \62016 , \62015 );
buf \U$62042 ( \62017 , \62016 );
xnor \U$62043 ( \62018 , \61981 , \62017 );
buf \U$62044 ( \62019 , \62018 );
buf \U$62045 ( \62020 , \62019 );
and \U$62046 ( \62021 , \61953 , \62020 );
and \U$62047 ( \62022 , \61886 , \61952 );
or \U$62048 ( \62023 , \62021 , \62022 );
buf \U$62049 ( \62024 , \62023 );
buf \U$62050 ( \62025 , \62024 );
not \U$62051 ( \62026 , \62025 );
buf \U$62052 ( \62027 , \61965 );
buf \U$62053 ( \62028 , \61972 );
not \U$62054 ( \62029 , \62028 );
buf \U$62055 ( \62030 , \62029 );
buf \U$62056 ( \62031 , \62030 );
nor \U$62057 ( \62032 , \62027 , \62031 );
buf \U$62058 ( \62033 , \62032 );
buf \U$62059 ( \62034 , \62033 );
buf \U$62060 ( \62035 , \62016 );
or \U$62061 ( \62036 , \62034 , \62035 );
buf \U$62062 ( \62037 , \61965 );
buf \U$62063 ( \62038 , \62030 );
nand \U$62064 ( \62039 , \62037 , \62038 );
buf \U$62065 ( \62040 , \62039 );
buf \U$62066 ( \62041 , \62040 );
nand \U$62067 ( \62042 , \62036 , \62041 );
buf \U$62068 ( \62043 , \62042 );
buf \U$62069 ( \62044 , \61554 );
buf \U$62070 ( \62045 , \61536 );
xor \U$62071 ( \62046 , \62044 , \62045 );
buf \U$62072 ( \62047 , \61576 );
xnor \U$62073 ( \62048 , \62046 , \62047 );
buf \U$62074 ( \62049 , \62048 );
xnor \U$62075 ( \62050 , \62043 , \62049 );
buf \U$62076 ( \62051 , \62050 );
not \U$62077 ( \62052 , \62051 );
buf \U$62078 ( \62053 , \13178 );
buf \U$62079 ( \62054 , \12911 );
buf \U$62080 ( \62055 , RIc0d9400_64);
and \U$62081 ( \62056 , \62054 , \62055 );
buf \U$62082 ( \62057 , \43843 );
buf \U$62083 ( \62058 , RIc0dadc8_119);
and \U$62084 ( \62059 , \62057 , \62058 );
nor \U$62085 ( \62060 , \62056 , \62059 );
buf \U$62086 ( \62061 , \62060 );
buf \U$62087 ( \62062 , \62061 );
nor \U$62088 ( \62063 , \62053 , \62062 );
buf \U$62089 ( \62064 , \62063 );
buf \U$62090 ( \62065 , \62064 );
buf \U$62091 ( \62066 , \45225 );
buf \U$62092 ( \62067 , \61011 );
nor \U$62093 ( \62068 , \62066 , \62067 );
buf \U$62094 ( \62069 , \62068 );
buf \U$62095 ( \62070 , \62069 );
nor \U$62096 ( \62071 , \62065 , \62070 );
buf \U$62097 ( \62072 , \62071 );
xor \U$62098 ( \62073 , \61494 , \61515 );
buf \U$62099 ( \62074 , \62073 );
xnor \U$62100 ( \62075 , \62072 , \62074 );
xor \U$62101 ( \62076 , \61860 , \61865 );
and \U$62102 ( \62077 , \62076 , \61883 );
and \U$62103 ( \62078 , \61860 , \61865 );
or \U$62104 ( \62079 , \62077 , \62078 );
buf \U$62105 ( \62080 , \62079 );
xnor \U$62106 ( \62081 , \62075 , \62080 );
buf \U$62107 ( \62082 , \62081 );
not \U$62108 ( \62083 , \62082 );
and \U$62109 ( \62084 , \62052 , \62083 );
buf \U$62110 ( \62085 , \62081 );
buf \U$62111 ( \62086 , \62050 );
and \U$62112 ( \62087 , \62085 , \62086 );
nor \U$62113 ( \62088 , \62084 , \62087 );
buf \U$62114 ( \62089 , \62088 );
buf \U$62115 ( \62090 , \62089 );
nand \U$62116 ( \62091 , \62026 , \62090 );
buf \U$62117 ( \62092 , \62091 );
buf \U$62118 ( \62093 , \62092 );
not \U$62119 ( \62094 , \62093 );
xor \U$62120 ( \62095 , \61886 , \61952 );
xor \U$62121 ( \62096 , \62095 , \62020 );
buf \U$62122 ( \62097 , \62096 );
buf \U$62123 ( \62098 , \62097 );
buf \U$62124 ( \62099 , \61997 );
buf \U$62125 ( \62100 , \62013 );
xor \U$62126 ( \62101 , \62099 , \62100 );
buf \U$62127 ( \62102 , \62101 );
buf \U$62128 ( \62103 , \62102 );
buf \U$62129 ( \62104 , \13314 );
buf \U$62130 ( \62105 , RIc0d9400_64);
and \U$62131 ( \62106 , \62104 , \62105 );
buf \U$62132 ( \62107 , \62106 );
buf \U$62133 ( \62108 , \62107 );
buf \U$62134 ( \62109 , RIc0dafa8_123);
buf \U$62135 ( \62110 , RIc0d9388_63);
and \U$62136 ( \62111 , \62109 , \62110 );
not \U$62137 ( \62112 , \62109 );
buf \U$62138 ( \62113 , \43939 );
and \U$62139 ( \62114 , \62112 , \62113 );
nor \U$62140 ( \62115 , \62111 , \62114 );
buf \U$62141 ( \62116 , \62115 );
buf \U$62142 ( \62117 , \62116 );
not \U$62143 ( \62118 , \62117 );
buf \U$62144 ( \62119 , \14982 );
not \U$62145 ( \62120 , \62119 );
or \U$62146 ( \62121 , \62118 , \62120 );
buf \U$62147 ( \62122 , \16692 );
buf \U$62148 ( \62123 , \61985 );
nand \U$62149 ( \62124 , \62122 , \62123 );
buf \U$62150 ( \62125 , \62124 );
buf \U$62151 ( \62126 , \62125 );
nand \U$62152 ( \62127 , \62121 , \62126 );
buf \U$62153 ( \62128 , \62127 );
buf \U$62154 ( \62129 , \62128 );
xor \U$62155 ( \62130 , \62108 , \62129 );
buf \U$62156 ( \62131 , RIc0d9298_61);
buf \U$62157 ( \62132 , RIc0db098_125);
xor \U$62158 ( \62133 , \62131 , \62132 );
buf \U$62159 ( \62134 , \62133 );
buf \U$62160 ( \62135 , \62134 );
not \U$62161 ( \62136 , \62135 );
buf \U$62162 ( \62137 , \13461 );
not \U$62163 ( \62138 , \62137 );
or \U$62164 ( \62139 , \62136 , \62138 );
buf \U$62165 ( \62140 , \15793 );
buf \U$62166 ( \62141 , \61904 );
nand \U$62167 ( \62142 , \62140 , \62141 );
buf \U$62168 ( \62143 , \62142 );
buf \U$62169 ( \62144 , \62143 );
nand \U$62170 ( \62145 , \62139 , \62144 );
buf \U$62171 ( \62146 , \62145 );
buf \U$62172 ( \62147 , \62146 );
and \U$62173 ( \62148 , \62130 , \62147 );
and \U$62174 ( \62149 , \62108 , \62129 );
or \U$62175 ( \62150 , \62148 , \62149 );
buf \U$62176 ( \62151 , \62150 );
buf \U$62177 ( \62152 , \62151 );
xor \U$62178 ( \62153 , \62103 , \62152 );
xor \U$62179 ( \62154 , \61900 , \61922 );
xor \U$62180 ( \62155 , \62154 , \61947 );
buf \U$62181 ( \62156 , \62155 );
buf \U$62182 ( \62157 , \62156 );
and \U$62183 ( \62158 , \62153 , \62157 );
and \U$62184 ( \62159 , \62103 , \62152 );
or \U$62185 ( \62160 , \62158 , \62159 );
buf \U$62186 ( \62161 , \62160 );
buf \U$62187 ( \62162 , \62161 );
nor \U$62188 ( \62163 , \62098 , \62162 );
buf \U$62189 ( \62164 , \62163 );
buf \U$62190 ( \62165 , \62164 );
nor \U$62191 ( \62166 , \62094 , \62165 );
buf \U$62192 ( \62167 , \62166 );
buf \U$62193 ( \62168 , \62167 );
buf \U$62194 ( \62169 , RIc0d9220_60);
buf \U$62195 ( \62170 , RIc0db188_127);
xor \U$62196 ( \62171 , \62169 , \62170 );
buf \U$62197 ( \62172 , \62171 );
buf \U$62198 ( \62173 , \62172 );
not \U$62199 ( \62174 , \62173 );
buf \U$62200 ( \62175 , \15609 );
not \U$62201 ( \62176 , \62175 );
or \U$62202 ( \62177 , \62174 , \62176 );
buf \U$62203 ( \62178 , RIc0db188_127);
not \U$62204 ( \62179 , \62178 );
buf \U$62205 ( \62180 , \16956 );
not \U$62206 ( \62181 , \62180 );
or \U$62207 ( \62182 , \62179 , \62181 );
buf \U$62208 ( \62183 , RIc0db188_127);
not \U$62209 ( \62184 , \62183 );
buf \U$62210 ( \62185 , RIc0d91a8_59);
nand \U$62211 ( \62186 , \62184 , \62185 );
buf \U$62212 ( \62187 , \62186 );
buf \U$62213 ( \62188 , \62187 );
nand \U$62214 ( \62189 , \62182 , \62188 );
buf \U$62215 ( \62190 , \62189 );
buf \U$62216 ( \62191 , \62190 );
buf \U$62217 ( \62192 , RIc0db200_128);
nand \U$62218 ( \62193 , \62191 , \62192 );
buf \U$62219 ( \62194 , \62193 );
buf \U$62220 ( \62195 , \62194 );
nand \U$62221 ( \62196 , \62177 , \62195 );
buf \U$62222 ( \62197 , \62196 );
buf \U$62223 ( \62198 , \62197 );
not \U$62224 ( \62199 , \62198 );
buf \U$62225 ( \62200 , RIc0d9400_64);
buf \U$62226 ( \62201 , RIc0db020_124);
or \U$62227 ( \62202 , \62200 , \62201 );
buf \U$62228 ( \62203 , RIc0db098_125);
nand \U$62229 ( \62204 , \62202 , \62203 );
buf \U$62230 ( \62205 , \62204 );
buf \U$62231 ( \62206 , \62205 );
buf \U$62232 ( \62207 , RIc0d9400_64);
buf \U$62233 ( \62208 , RIc0db020_124);
nand \U$62234 ( \62209 , \62207 , \62208 );
buf \U$62235 ( \62210 , \62209 );
buf \U$62236 ( \62211 , \62210 );
buf \U$62237 ( \62212 , RIc0dafa8_123);
nand \U$62238 ( \62213 , \62206 , \62211 , \62212 );
buf \U$62239 ( \62214 , \62213 );
buf \U$62240 ( \62215 , \62214 );
nor \U$62241 ( \62216 , \62199 , \62215 );
buf \U$62242 ( \62217 , \62216 );
buf \U$62243 ( \62218 , \62217 );
not \U$62244 ( \62219 , \62218 );
buf \U$62245 ( \62220 , \62190 );
not \U$62246 ( \62221 , \62220 );
buf \U$62247 ( \62222 , \60911 );
not \U$62248 ( \62223 , \62222 );
or \U$62249 ( \62224 , \62221 , \62223 );
buf \U$62250 ( \62225 , \61892 );
not \U$62251 ( \62226 , \62225 );
buf \U$62252 ( \62227 , RIc0db200_128);
nand \U$62253 ( \62228 , \62226 , \62227 );
buf \U$62254 ( \62229 , \62228 );
buf \U$62255 ( \62230 , \62229 );
nand \U$62256 ( \62231 , \62224 , \62230 );
buf \U$62257 ( \62232 , \62231 );
buf \U$62258 ( \62233 , \62232 );
not \U$62259 ( \62234 , \62233 );
or \U$62260 ( \62235 , \62219 , \62234 );
buf \U$62261 ( \62236 , \62217 );
buf \U$62262 ( \62237 , \62232 );
or \U$62263 ( \62238 , \62236 , \62237 );
xor \U$62264 ( \62239 , \62108 , \62129 );
xor \U$62265 ( \62240 , \62239 , \62147 );
buf \U$62266 ( \62241 , \62240 );
buf \U$62267 ( \62242 , \62241 );
nand \U$62268 ( \62243 , \62238 , \62242 );
buf \U$62269 ( \62244 , \62243 );
buf \U$62270 ( \62245 , \62244 );
nand \U$62271 ( \62246 , \62235 , \62245 );
buf \U$62272 ( \62247 , \62246 );
buf \U$62273 ( \62248 , \62247 );
xor \U$62274 ( \62249 , \62103 , \62152 );
xor \U$62275 ( \62250 , \62249 , \62157 );
buf \U$62276 ( \62251 , \62250 );
buf \U$62277 ( \62252 , \62251 );
xor \U$62278 ( \62253 , \62248 , \62252 );
buf \U$62279 ( \62254 , RIc0d9310_62);
buf \U$62280 ( \62255 , RIc0db098_125);
xor \U$62281 ( \62256 , \62254 , \62255 );
buf \U$62282 ( \62257 , \62256 );
buf \U$62283 ( \62258 , \62257 );
not \U$62284 ( \62259 , \62258 );
buf \U$62285 ( \62260 , \51095 );
not \U$62286 ( \62261 , \62260 );
or \U$62287 ( \62262 , \62259 , \62261 );
buf \U$62288 ( \62263 , \15793 );
buf \U$62289 ( \62264 , \62134 );
nand \U$62290 ( \62265 , \62263 , \62264 );
buf \U$62291 ( \62266 , \62265 );
buf \U$62292 ( \62267 , \62266 );
nand \U$62293 ( \62268 , \62262 , \62267 );
buf \U$62294 ( \62269 , \62268 );
buf \U$62295 ( \62270 , \62269 );
not \U$62296 ( \62271 , \62270 );
buf \U$62297 ( \62272 , \62197 );
not \U$62298 ( \62273 , \62272 );
buf \U$62299 ( \62274 , \62214 );
not \U$62300 ( \62275 , \62274 );
and \U$62301 ( \62276 , \62273 , \62275 );
buf \U$62302 ( \62277 , \62197 );
buf \U$62303 ( \62278 , \62214 );
and \U$62304 ( \62279 , \62277 , \62278 );
nor \U$62305 ( \62280 , \62276 , \62279 );
buf \U$62306 ( \62281 , \62280 );
buf \U$62307 ( \62282 , \62281 );
not \U$62308 ( \62283 , \62282 );
buf \U$62309 ( \62284 , \62283 );
buf \U$62310 ( \62285 , \62284 );
not \U$62311 ( \62286 , \62285 );
or \U$62312 ( \62287 , \62271 , \62286 );
buf \U$62313 ( \62288 , \62284 );
buf \U$62314 ( \62289 , \62269 );
or \U$62315 ( \62290 , \62288 , \62289 );
buf \U$62316 ( \62291 , \62116 );
not \U$62317 ( \62292 , \62291 );
buf \U$62318 ( \62293 , \16692 );
not \U$62319 ( \62294 , \62293 );
or \U$62320 ( \62295 , \62292 , \62294 );
buf \U$62321 ( \62296 , \45089 );
buf \U$62322 ( \62297 , RIc0dafa8_123);
buf \U$62323 ( \62298 , \43843 );
and \U$62324 ( \62299 , \62297 , \62298 );
not \U$62325 ( \62300 , \62297 );
buf \U$62326 ( \62301 , RIc0d9400_64);
and \U$62327 ( \62302 , \62300 , \62301 );
nor \U$62328 ( \62303 , \62299 , \62302 );
buf \U$62329 ( \62304 , \62303 );
buf \U$62330 ( \62305 , \62304 );
or \U$62331 ( \62306 , \62296 , \62305 );
nand \U$62332 ( \62307 , \62295 , \62306 );
buf \U$62333 ( \62308 , \62307 );
buf \U$62334 ( \62309 , \62308 );
nand \U$62335 ( \62310 , \62290 , \62309 );
buf \U$62336 ( \62311 , \62310 );
buf \U$62337 ( \62312 , \62311 );
nand \U$62338 ( \62313 , \62287 , \62312 );
buf \U$62339 ( \62314 , \62313 );
buf \U$62340 ( \62315 , \62314 );
not \U$62341 ( \62316 , \62315 );
buf \U$62342 ( \62317 , \62241 );
buf \U$62343 ( \62318 , \62217 );
buf \U$62344 ( \62319 , \62232 );
xor \U$62345 ( \62320 , \62318 , \62319 );
buf \U$62346 ( \62321 , \62320 );
buf \U$62347 ( \62322 , \62321 );
xnor \U$62348 ( \62323 , \62317 , \62322 );
buf \U$62349 ( \62324 , \62323 );
buf \U$62350 ( \62325 , \62324 );
nand \U$62351 ( \62326 , \62316 , \62325 );
buf \U$62352 ( \62327 , \62326 );
not \U$62353 ( \62328 , \62327 );
buf \U$62354 ( \62329 , RIc0d9400_64);
buf \U$62355 ( \62330 , RIc0db110_126);
or \U$62356 ( \62331 , \62329 , \62330 );
buf \U$62357 ( \62332 , RIc0db188_127);
nand \U$62358 ( \62333 , \62331 , \62332 );
buf \U$62359 ( \62334 , \62333 );
buf \U$62360 ( \62335 , \62334 );
buf \U$62361 ( \62336 , RIc0d9400_64);
buf \U$62362 ( \62337 , RIc0db110_126);
nand \U$62363 ( \62338 , \62336 , \62337 );
buf \U$62364 ( \62339 , \62338 );
buf \U$62365 ( \62340 , \62339 );
buf \U$62366 ( \62341 , RIc0db098_125);
and \U$62367 ( \62342 , \62335 , \62340 , \62341 );
buf \U$62368 ( \62343 , \62342 );
buf \U$62369 ( \62344 , \62343 );
buf \U$62370 ( \62345 , RIc0db200_128);
not \U$62371 ( \62346 , \62345 );
buf \U$62372 ( \62347 , RIc0d9298_61);
buf \U$62373 ( \62348 , RIc0db188_127);
xor \U$62374 ( \62349 , \62347 , \62348 );
buf \U$62375 ( \62350 , \62349 );
buf \U$62376 ( \62351 , \62350 );
not \U$62377 ( \62352 , \62351 );
or \U$62378 ( \62353 , \62346 , \62352 );
buf \U$62379 ( \62354 , \47878 );
buf \U$62380 ( \62355 , RIc0d9310_62);
buf \U$62381 ( \62356 , RIc0db188_127);
xor \U$62382 ( \62357 , \62355 , \62356 );
buf \U$62383 ( \62358 , \62357 );
buf \U$62384 ( \62359 , \62358 );
not \U$62385 ( \62360 , \62359 );
buf \U$62386 ( \62361 , \62360 );
buf \U$62387 ( \62362 , \62361 );
or \U$62388 ( \62363 , \62354 , \62362 );
nand \U$62389 ( \62364 , \62353 , \62363 );
buf \U$62390 ( \62365 , \62364 );
buf \U$62391 ( \62366 , \62365 );
and \U$62392 ( \62367 , \62344 , \62366 );
buf \U$62393 ( \62368 , \62367 );
buf \U$62394 ( \62369 , \62368 );
not \U$62395 ( \62370 , \62369 );
buf \U$62396 ( \62371 , \16692 );
buf \U$62397 ( \62372 , RIc0d9400_64);
and \U$62398 ( \62373 , \62371 , \62372 );
buf \U$62399 ( \62374 , \62373 );
buf \U$62400 ( \62375 , \43781 );
buf \U$62401 ( \62376 , \62350 );
and \U$62402 ( \62377 , \62375 , \62376 );
buf \U$62403 ( \62378 , \62172 );
not \U$62404 ( \62379 , \62378 );
buf \U$62405 ( \62380 , \12647 );
nor \U$62406 ( \62381 , \62379 , \62380 );
buf \U$62407 ( \62382 , \62381 );
buf \U$62408 ( \62383 , \62382 );
nor \U$62409 ( \62384 , \62377 , \62383 );
buf \U$62410 ( \62385 , \62384 );
xor \U$62411 ( \62386 , \62374 , \62385 );
xnor \U$62412 ( \62387 , RIc0db098_125, RIc0d9388_63);
buf \U$62413 ( \62388 , \62387 );
not \U$62414 ( \62389 , \62388 );
buf \U$62415 ( \62390 , \62389 );
buf \U$62416 ( \62391 , \62390 );
not \U$62417 ( \62392 , \62391 );
buf \U$62418 ( \62393 , \44382 );
not \U$62419 ( \62394 , \62393 );
or \U$62420 ( \62395 , \62392 , \62394 );
buf \U$62421 ( \62396 , \13465 );
buf \U$62422 ( \62397 , \62257 );
nand \U$62423 ( \62398 , \62396 , \62397 );
buf \U$62424 ( \62399 , \62398 );
buf \U$62425 ( \62400 , \62399 );
nand \U$62426 ( \62401 , \62395 , \62400 );
buf \U$62427 ( \62402 , \62401 );
xor \U$62428 ( \62403 , \62386 , \62402 );
buf \U$62429 ( \62404 , \62403 );
nand \U$62430 ( \62405 , \62370 , \62404 );
buf \U$62431 ( \62406 , \62405 );
not \U$62432 ( \62407 , \62406 );
buf \U$62433 ( \62408 , \15609 );
not \U$62434 ( \62409 , \62408 );
buf \U$62435 ( \62410 , RIc0db188_127);
buf \U$62436 ( \62411 , RIc0d9388_63);
and \U$62437 ( \62412 , \62410 , \62411 );
not \U$62438 ( \62413 , \62410 );
buf \U$62439 ( \62414 , \43939 );
and \U$62440 ( \62415 , \62413 , \62414 );
nor \U$62441 ( \62416 , \62412 , \62415 );
buf \U$62442 ( \62417 , \62416 );
buf \U$62443 ( \62418 , \62417 );
not \U$62444 ( \62419 , \62418 );
or \U$62445 ( \62420 , \62409 , \62419 );
buf \U$62446 ( \62421 , \62358 );
buf \U$62447 ( \62422 , RIc0db200_128);
nand \U$62448 ( \62423 , \62421 , \62422 );
buf \U$62449 ( \62424 , \62423 );
buf \U$62450 ( \62425 , \62424 );
nand \U$62451 ( \62426 , \62420 , \62425 );
buf \U$62452 ( \62427 , \62426 );
buf \U$62453 ( \62428 , \62427 );
not \U$62454 ( \62429 , \62428 );
buf \U$62455 ( \62430 , \15793 );
buf \U$62456 ( \62431 , RIc0d9400_64);
nand \U$62457 ( \62432 , \62430 , \62431 );
buf \U$62458 ( \62433 , \62432 );
buf \U$62459 ( \62434 , \62433 );
nand \U$62460 ( \62435 , \62429 , \62434 );
buf \U$62461 ( \62436 , \62435 );
buf \U$62462 ( \62437 , \62436 );
buf \U$62463 ( \62438 , \43843 );
not \U$62464 ( \62439 , \62438 );
buf \U$62465 ( \62440 , \15609 );
not \U$62466 ( \62441 , \62440 );
or \U$62467 ( \62442 , \62439 , \62441 );
buf \U$62468 ( \62443 , RIc0db200_128);
buf \U$62469 ( \62444 , \62417 );
nand \U$62470 ( \62445 , \62443 , \62444 );
buf \U$62471 ( \62446 , \62445 );
buf \U$62472 ( \62447 , \62446 );
nand \U$62473 ( \62448 , \62442 , \62447 );
buf \U$62474 ( \62449 , \62448 );
buf \U$62475 ( \62450 , \62449 );
buf \U$62476 ( \62451 , RIc0d9400_64);
buf \U$62477 ( \62452 , RIc0db200_128);
nand \U$62478 ( \62453 , \62451 , \62452 );
buf \U$62479 ( \62454 , \62453 );
and \U$62480 ( \62455 , \62454 , RIc0db188_127);
buf \U$62481 ( \62456 , \62455 );
and \U$62482 ( \62457 , \62450 , \62456 );
buf \U$62483 ( \62458 , \62457 );
buf \U$62484 ( \62459 , \62458 );
nand \U$62485 ( \62460 , \62437 , \62459 );
buf \U$62486 ( \62461 , \62460 );
buf \U$62487 ( \62462 , \62461 );
buf \U$62488 ( \62463 , \62433 );
not \U$62489 ( \62464 , \62463 );
buf \U$62490 ( \62465 , \62427 );
nand \U$62491 ( \62466 , \62464 , \62465 );
buf \U$62492 ( \62467 , \62466 );
buf \U$62493 ( \62468 , \62467 );
and \U$62494 ( \62469 , \62462 , \62468 );
buf \U$62495 ( \62470 , \62469 );
buf \U$62496 ( \62471 , \62470 );
xor \U$62497 ( \62472 , \62344 , \62366 );
buf \U$62498 ( \62473 , \62472 );
buf \U$62499 ( \62474 , \62473 );
buf \U$62500 ( \62475 , \46459 );
buf \U$62501 ( \62476 , RIc0db098_125);
buf \U$62502 ( \62477 , \43843 );
and \U$62503 ( \62478 , \62476 , \62477 );
not \U$62504 ( \62479 , \62476 );
buf \U$62505 ( \62480 , RIc0d9400_64);
and \U$62506 ( \62481 , \62479 , \62480 );
nor \U$62507 ( \62482 , \62478 , \62481 );
buf \U$62508 ( \62483 , \62482 );
buf \U$62509 ( \62484 , \62483 );
or \U$62510 ( \62485 , \62475 , \62484 );
buf \U$62511 ( \62486 , \18699 );
buf \U$62512 ( \62487 , \62387 );
or \U$62513 ( \62488 , \62486 , \62487 );
nand \U$62514 ( \62489 , \62485 , \62488 );
buf \U$62515 ( \62490 , \62489 );
buf \U$62516 ( \62491 , \62490 );
nor \U$62517 ( \62492 , \62474 , \62491 );
buf \U$62518 ( \62493 , \62492 );
buf \U$62519 ( \62494 , \62493 );
or \U$62520 ( \62495 , \62471 , \62494 );
buf \U$62521 ( \62496 , \62473 );
buf \U$62522 ( \62497 , \62490 );
nand \U$62523 ( \62498 , \62496 , \62497 );
buf \U$62524 ( \62499 , \62498 );
buf \U$62525 ( \62500 , \62499 );
nand \U$62526 ( \62501 , \62495 , \62500 );
buf \U$62527 ( \62502 , \62501 );
not \U$62528 ( \62503 , \62502 );
or \U$62529 ( \62504 , \62407 , \62503 );
buf \U$62530 ( \62505 , \62403 );
not \U$62531 ( \62506 , \62505 );
buf \U$62532 ( \62507 , \62368 );
nand \U$62533 ( \62508 , \62506 , \62507 );
buf \U$62534 ( \62509 , \62508 );
nand \U$62535 ( \62510 , \62504 , \62509 );
buf \U$62536 ( \62511 , \62510 );
buf \U$62537 ( \62512 , \62385 );
not \U$62538 ( \62513 , \62512 );
buf \U$62539 ( \62514 , \62513 );
buf \U$62540 ( \62515 , \62514 );
not \U$62541 ( \62516 , \62515 );
buf \U$62542 ( \62517 , \62374 );
not \U$62543 ( \62518 , \62517 );
or \U$62544 ( \62519 , \62516 , \62518 );
buf \U$62545 ( \62520 , \62374 );
buf \U$62546 ( \62521 , \62514 );
or \U$62547 ( \62522 , \62520 , \62521 );
buf \U$62548 ( \62523 , \62402 );
nand \U$62549 ( \62524 , \62522 , \62523 );
buf \U$62550 ( \62525 , \62524 );
buf \U$62551 ( \62526 , \62525 );
nand \U$62552 ( \62527 , \62519 , \62526 );
buf \U$62553 ( \62528 , \62527 );
buf \U$62554 ( \62529 , \62528 );
not \U$62555 ( \62530 , \62529 );
xor \U$62556 ( \62531 , \62269 , \62281 );
xor \U$62557 ( \62532 , \62531 , \62308 );
buf \U$62558 ( \62533 , \62532 );
nand \U$62559 ( \62534 , \62530 , \62533 );
buf \U$62560 ( \62535 , \62534 );
buf \U$62561 ( \62536 , \62535 );
nand \U$62562 ( \62537 , \62511 , \62536 );
buf \U$62563 ( \62538 , \62537 );
buf \U$62564 ( \62539 , \62538 );
buf \U$62565 ( \62540 , \62532 );
not \U$62566 ( \62541 , \62540 );
buf \U$62567 ( \62542 , \62541 );
buf \U$62568 ( \62543 , \62542 );
buf \U$62569 ( \62544 , \62528 );
nand \U$62570 ( \62545 , \62543 , \62544 );
buf \U$62571 ( \62546 , \62545 );
buf \U$62572 ( \62547 , \62546 );
nand \U$62573 ( \62548 , \62539 , \62547 );
buf \U$62574 ( \62549 , \62548 );
not \U$62575 ( \62550 , \62549 );
or \U$62576 ( \62551 , \62328 , \62550 );
buf \U$62577 ( \62552 , \62324 );
not \U$62578 ( \62553 , \62552 );
buf \U$62579 ( \62554 , \62314 );
nand \U$62580 ( \62555 , \62553 , \62554 );
buf \U$62581 ( \62556 , \62555 );
nand \U$62582 ( \62557 , \62551 , \62556 );
buf \U$62583 ( \62558 , \62557 );
and \U$62584 ( \62559 , \62253 , \62558 );
and \U$62585 ( \62560 , \62248 , \62252 );
or \U$62586 ( \62561 , \62559 , \62560 );
buf \U$62587 ( \62562 , \62561 );
buf \U$62588 ( \62563 , \62562 );
nand \U$62589 ( \62564 , \62168 , \62563 );
buf \U$62590 ( \62565 , \62564 );
buf \U$62591 ( \62566 , \62565 );
not \U$62592 ( \62567 , \62566 );
buf \U$62593 ( \62568 , \62097 );
buf \U$62594 ( \62569 , \62161 );
nand \U$62595 ( \62570 , \62568 , \62569 );
buf \U$62596 ( \62571 , \62570 );
buf \U$62597 ( \62572 , \62571 );
not \U$62598 ( \62573 , \62572 );
buf \U$62599 ( \62574 , \62092 );
nand \U$62600 ( \62575 , \62573 , \62574 );
buf \U$62601 ( \62576 , \62575 );
buf \U$62602 ( \62577 , \62576 );
buf \U$62603 ( \62578 , \62089 );
not \U$62604 ( \62579 , \62578 );
buf \U$62605 ( \62580 , \62024 );
nand \U$62606 ( \62581 , \62579 , \62580 );
buf \U$62607 ( \62582 , \62581 );
buf \U$62608 ( \62583 , \62582 );
nand \U$62609 ( \62584 , \62577 , \62583 );
buf \U$62610 ( \62585 , \62584 );
buf \U$62611 ( \62586 , \62585 );
buf \U$62612 ( \62587 , \62081 );
not \U$62613 ( \62588 , \62587 );
buf \U$62614 ( \62589 , \62043 );
not \U$62615 ( \62590 , \62589 );
buf \U$62616 ( \62591 , \62049 );
nand \U$62617 ( \62592 , \62590 , \62591 );
buf \U$62618 ( \62593 , \62592 );
buf \U$62619 ( \62594 , \62593 );
nand \U$62620 ( \62595 , \62588 , \62594 );
buf \U$62621 ( \62596 , \62595 );
buf \U$62622 ( \62597 , \62596 );
buf \U$62623 ( \62598 , \62049 );
not \U$62624 ( \62599 , \62598 );
buf \U$62625 ( \62600 , \62043 );
nand \U$62626 ( \62601 , \62599 , \62600 );
buf \U$62627 ( \62602 , \62601 );
buf \U$62628 ( \62603 , \62602 );
nand \U$62629 ( \62604 , \62597 , \62603 );
buf \U$62630 ( \62605 , \62604 );
buf \U$62631 ( \62606 , \62605 );
not \U$62632 ( \62607 , \62606 );
buf \U$62633 ( \62608 , \62072 );
not \U$62634 ( \62609 , \62608 );
buf \U$62635 ( \62610 , \62609 );
buf \U$62636 ( \62611 , \62610 );
not \U$62637 ( \62612 , \62611 );
buf \U$62638 ( \62613 , \62074 );
not \U$62639 ( \62614 , \62613 );
or \U$62640 ( \62615 , \62612 , \62614 );
buf \U$62641 ( \62616 , \62072 );
not \U$62642 ( \62617 , \62616 );
buf \U$62643 ( \62618 , \62074 );
not \U$62644 ( \62619 , \62618 );
buf \U$62645 ( \62620 , \62619 );
buf \U$62646 ( \62621 , \62620 );
not \U$62647 ( \62622 , \62621 );
or \U$62648 ( \62623 , \62617 , \62622 );
buf \U$62649 ( \62624 , \62080 );
nand \U$62650 ( \62625 , \62623 , \62624 );
buf \U$62651 ( \62626 , \62625 );
buf \U$62652 ( \62627 , \62626 );
nand \U$62653 ( \62628 , \62615 , \62627 );
buf \U$62654 ( \62629 , \62628 );
buf \U$62655 ( \62630 , \62629 );
not \U$62656 ( \62631 , \62630 );
xor \U$62657 ( \62632 , \60972 , \60946 );
xor \U$62658 ( \62633 , \62632 , \60928 );
buf \U$62659 ( \62634 , \62633 );
not \U$62660 ( \62635 , \62634 );
buf \U$62661 ( \62636 , \62635 );
buf \U$62662 ( \62637 , \62636 );
not \U$62663 ( \62638 , \62637 );
and \U$62664 ( \62639 , \62631 , \62638 );
buf \U$62665 ( \62640 , \62629 );
buf \U$62666 ( \62641 , \62636 );
and \U$62667 ( \62642 , \62640 , \62641 );
nor \U$62668 ( \62643 , \62639 , \62642 );
buf \U$62669 ( \62644 , \62643 );
xor \U$62670 ( \62645 , \61518 , \61522 );
xor \U$62671 ( \62646 , \62645 , \61583 );
buf \U$62672 ( \62647 , \62646 );
xor \U$62673 ( \62648 , \62644 , \62647 );
buf \U$62674 ( \62649 , \62648 );
nor \U$62675 ( \62650 , \62607 , \62649 );
buf \U$62676 ( \62651 , \62650 );
buf \U$62677 ( \62652 , \62651 );
nor \U$62678 ( \62653 , \62586 , \62652 );
buf \U$62679 ( \62654 , \62653 );
buf \U$62680 ( \62655 , \62654 );
not \U$62681 ( \62656 , \62655 );
or \U$62682 ( \62657 , \62567 , \62656 );
buf \U$62683 ( \62658 , \62633 );
not \U$62684 ( \62659 , \62658 );
buf \U$62685 ( \62660 , \62647 );
not \U$62686 ( \62661 , \62660 );
or \U$62687 ( \62662 , \62659 , \62661 );
buf \U$62688 ( \62663 , \62647 );
buf \U$62689 ( \62664 , \62633 );
or \U$62690 ( \62665 , \62663 , \62664 );
buf \U$62691 ( \62666 , \62629 );
nand \U$62692 ( \62667 , \62665 , \62666 );
buf \U$62693 ( \62668 , \62667 );
buf \U$62694 ( \62669 , \62668 );
nand \U$62695 ( \62670 , \62662 , \62669 );
buf \U$62696 ( \62671 , \62670 );
buf \U$62697 ( \62672 , \62671 );
not \U$62698 ( \62673 , \62672 );
buf \U$62699 ( \62674 , \61472 );
buf \U$62700 ( \62675 , \61587 );
xor \U$62701 ( \62676 , \62674 , \62675 );
buf \U$62702 ( \62677 , \61476 );
xnor \U$62703 ( \62678 , \62676 , \62677 );
buf \U$62704 ( \62679 , \62678 );
buf \U$62705 ( \62680 , \62679 );
nand \U$62706 ( \62681 , \62673 , \62680 );
buf \U$62707 ( \62682 , \62681 );
buf \U$62708 ( \62683 , \62682 );
buf \U$62709 ( \62684 , \62605 );
not \U$62710 ( \62685 , \62684 );
buf \U$62711 ( \62686 , \62648 );
nand \U$62712 ( \62687 , \62685 , \62686 );
buf \U$62713 ( \62688 , \62687 );
buf \U$62714 ( \62689 , \62688 );
and \U$62715 ( \62690 , \62683 , \62689 );
buf \U$62716 ( \62691 , \62690 );
buf \U$62717 ( \62692 , \62691 );
nand \U$62718 ( \62693 , \62657 , \62692 );
buf \U$62719 ( \62694 , \62693 );
buf \U$62720 ( \62695 , \62694 );
buf \U$62721 ( \62696 , \62679 );
not \U$62722 ( \62697 , \62696 );
buf \U$62723 ( \62698 , \62671 );
nand \U$62724 ( \62699 , \62697 , \62698 );
buf \U$62725 ( \62700 , \62699 );
buf \U$62726 ( \62701 , \62700 );
nand \U$62727 ( \62702 , \62695 , \62701 );
buf \U$62728 ( \62703 , \62702 );
buf \U$62729 ( \62704 , \62703 );
buf \U$62730 ( \62705 , \61767 );
not \U$62731 ( \62706 , \62705 );
buf \U$62732 ( \62707 , \61468 );
buf \U$62733 ( \62708 , \61598 );
not \U$62734 ( \62709 , \62708 );
buf \U$62735 ( \62710 , \61620 );
nand \U$62736 ( \62711 , \62709 , \62710 );
buf \U$62737 ( \62712 , \62711 );
buf \U$62738 ( \62713 , \62712 );
nand \U$62739 ( \62714 , \62707 , \62713 );
buf \U$62740 ( \62715 , \62714 );
buf \U$62741 ( \62716 , \62715 );
nor \U$62742 ( \62717 , \62706 , \62716 );
buf \U$62743 ( \62718 , \62717 );
buf \U$62744 ( \62719 , \62718 );
buf \U$62745 ( \62720 , \61843 );
nand \U$62746 ( \62721 , \62704 , \62719 , \62720 );
buf \U$62747 ( \62722 , \62721 );
buf \U$62748 ( \62723 , \62722 );
buf \U$62749 ( \62724 , \61840 );
not \U$62750 ( \62725 , \62724 );
buf \U$62751 ( \62726 , \61793 );
nand \U$62752 ( \62727 , \62725 , \62726 );
buf \U$62753 ( \62728 , \62727 );
buf \U$62754 ( \62729 , \62728 );
nand \U$62755 ( \62730 , \61847 , \62723 , \62729 );
buf \U$62756 ( \62731 , \62730 );
buf \U$62757 ( \62732 , \62731 );
xor \U$62758 ( \62733 , \60597 , \60756 );
xor \U$62759 ( \62734 , \62733 , \60761 );
buf \U$62760 ( \62735 , \62734 );
buf \U$62761 ( \62736 , \62735 );
buf \U$62762 ( \62737 , \60507 );
buf \U$62763 ( \62738 , \60512 );
xor \U$62764 ( \62739 , \62737 , \62738 );
buf \U$62765 ( \62740 , \60541 );
xor \U$62766 ( \62741 , \62739 , \62740 );
buf \U$62767 ( \62742 , \62741 );
buf \U$62768 ( \62743 , \62742 );
buf \U$62769 ( \62744 , \61800 );
not \U$62770 ( \62745 , \62744 );
buf \U$62771 ( \62746 , \61806 );
not \U$62772 ( \62747 , \62746 );
buf \U$62773 ( \62748 , \62747 );
buf \U$62774 ( \62749 , \62748 );
not \U$62775 ( \62750 , \62749 );
or \U$62776 ( \62751 , \62745 , \62750 );
buf \U$62777 ( \62752 , \62748 );
buf \U$62778 ( \62753 , \61800 );
or \U$62779 ( \62754 , \62752 , \62753 );
buf \U$62780 ( \62755 , \61812 );
nand \U$62781 ( \62756 , \62754 , \62755 );
buf \U$62782 ( \62757 , \62756 );
buf \U$62783 ( \62758 , \62757 );
nand \U$62784 ( \62759 , \62751 , \62758 );
buf \U$62785 ( \62760 , \62759 );
buf \U$62786 ( \62761 , \62760 );
xor \U$62787 ( \62762 , \62743 , \62761 );
xor \U$62788 ( \62763 , \60670 , \60746 );
xor \U$62789 ( \62764 , \62763 , \60751 );
buf \U$62790 ( \62765 , \62764 );
buf \U$62791 ( \62766 , \62765 );
and \U$62792 ( \62767 , \62762 , \62766 );
and \U$62793 ( \62768 , \62743 , \62761 );
or \U$62794 ( \62769 , \62767 , \62768 );
buf \U$62795 ( \62770 , \62769 );
buf \U$62796 ( \62771 , \62770 );
or \U$62797 ( \62772 , \62736 , \62771 );
buf \U$62798 ( \62773 , \62772 );
buf \U$62799 ( \62774 , \62773 );
buf \U$62800 ( \62775 , \61824 );
not \U$62801 ( \62776 , \62775 );
buf \U$62802 ( \62777 , \61813 );
not \U$62803 ( \62778 , \62777 );
buf \U$62804 ( \62779 , \62778 );
buf \U$62805 ( \62780 , \62779 );
not \U$62806 ( \62781 , \62780 );
or \U$62807 ( \62782 , \62776 , \62781 );
buf \U$62808 ( \62783 , \61817 );
not \U$62809 ( \62784 , \62783 );
buf \U$62810 ( \62785 , \61824 );
not \U$62811 ( \62786 , \62785 );
buf \U$62812 ( \62787 , \61813 );
nand \U$62813 ( \62788 , \62786 , \62787 );
buf \U$62814 ( \62789 , \62788 );
buf \U$62815 ( \62790 , \62789 );
nand \U$62816 ( \62791 , \62784 , \62790 );
buf \U$62817 ( \62792 , \62791 );
buf \U$62818 ( \62793 , \62792 );
nand \U$62819 ( \62794 , \62782 , \62793 );
buf \U$62820 ( \62795 , \62794 );
buf \U$62821 ( \62796 , \62795 );
xor \U$62822 ( \62797 , \62743 , \62761 );
xor \U$62823 ( \62798 , \62797 , \62766 );
buf \U$62824 ( \62799 , \62798 );
buf \U$62825 ( \62800 , \62799 );
or \U$62826 ( \62801 , \62796 , \62800 );
buf \U$62827 ( \62802 , \62801 );
buf \U$62828 ( \62803 , \62802 );
and \U$62829 ( \62804 , \62774 , \62803 );
buf \U$62830 ( \62805 , \62804 );
buf \U$62831 ( \62806 , \62805 );
nand \U$62832 ( \62807 , \60772 , \62732 , \62806 );
buf \U$62833 ( \62808 , \62807 );
buf \U$62834 ( \62809 , \62808 );
buf \U$62835 ( \62810 , \60771 );
buf \U$62836 ( \62811 , \62799 );
buf \U$62837 ( \62812 , \62795 );
nand \U$62838 ( \62813 , \62811 , \62812 );
buf \U$62839 ( \62814 , \62813 );
buf \U$62840 ( \62815 , \62814 );
not \U$62841 ( \62816 , \62815 );
buf \U$62842 ( \62817 , \62773 );
nand \U$62843 ( \62818 , \62816 , \62817 );
buf \U$62844 ( \62819 , \62818 );
buf \U$62845 ( \62820 , \62819 );
buf \U$62846 ( \62821 , \62735 );
buf \U$62847 ( \62822 , \62770 );
nand \U$62848 ( \62823 , \62821 , \62822 );
buf \U$62849 ( \62824 , \62823 );
buf \U$62850 ( \62825 , \62824 );
nand \U$62851 ( \62826 , \62820 , \62825 );
buf \U$62852 ( \62827 , \62826 );
buf \U$62853 ( \62828 , \62827 );
nand \U$62854 ( \62829 , \62810 , \62828 );
buf \U$62855 ( \62830 , \62829 );
buf \U$62856 ( \62831 , \62830 );
buf \U$62857 ( \62832 , \60592 );
buf \U$62858 ( \62833 , \60765 );
nand \U$62859 ( \62834 , \62832 , \62833 );
buf \U$62860 ( \62835 , \62834 );
buf \U$62861 ( \62836 , \62835 );
not \U$62862 ( \62837 , \62836 );
buf \U$62863 ( \62838 , \60588 );
nand \U$62864 ( \62839 , \62837 , \62838 );
buf \U$62865 ( \62840 , \62839 );
buf \U$62866 ( \62841 , \62840 );
buf \U$62867 ( \62842 , \60585 );
not \U$62868 ( \62843 , \62842 );
buf \U$62869 ( \62844 , \60566 );
nand \U$62870 ( \62845 , \62843 , \62844 );
buf \U$62871 ( \62846 , \62845 );
buf \U$62872 ( \62847 , \62846 );
and \U$62873 ( \62848 , \62841 , \62847 );
buf \U$62874 ( \62849 , \62848 );
buf \U$62875 ( \62850 , \62849 );
nand \U$62876 ( \62851 , \62809 , \62831 , \62850 );
buf \U$62877 ( \62852 , \62851 );
buf \U$62878 ( \62853 , \62852 );
buf \U$62879 ( \62854 , \60024 );
buf \U$62880 ( \62855 , \60261 );
or \U$62881 ( \62856 , \62854 , \62855 );
buf \U$62882 ( \62857 , \62856 );
buf \U$62883 ( \62858 , \62857 );
buf \U$62884 ( \62859 , \60282 );
nand \U$62885 ( \62860 , \62858 , \62859 );
buf \U$62886 ( \62861 , \62860 );
buf \U$62887 ( \62862 , \62861 );
buf \U$62888 ( \62863 , \60331 );
buf \U$62889 ( \62864 , \59745 );
nand \U$62890 ( \62865 , \62863 , \62864 );
buf \U$62891 ( \62866 , \62865 );
buf \U$62892 ( \62867 , \62866 );
nor \U$62893 ( \62868 , \62862 , \62867 );
buf \U$62894 ( \62869 , \62868 );
buf \U$62895 ( \62870 , \62869 );
nand \U$62896 ( \62871 , \62853 , \62870 );
buf \U$62897 ( \62872 , \62871 );
buf \U$62898 ( \62873 , \62872 );
buf \U$62899 ( \62874 , \60322 );
buf \U$62900 ( \62875 , \60328 );
nand \U$62901 ( \62876 , \62874 , \62875 );
buf \U$62902 ( \62877 , \62876 );
buf \U$62903 ( \62878 , \62877 );
nand \U$62904 ( \62879 , \60335 , \62873 , \62878 );
buf \U$62905 ( \62880 , \62879 );
buf \U$62906 ( \62881 , \62880 );
not \U$62907 ( \62882 , \62881 );
or \U$62908 ( \62883 , \59426 , \62882 );
buf \U$62909 ( \62884 , \57946 );
not \U$62910 ( \62885 , \62884 );
buf \U$62911 ( \62886 , \62885 );
buf \U$62912 ( \62887 , \62886 );
buf \U$62913 ( \62888 , \58721 );
not \U$62914 ( \62889 , \62888 );
buf \U$62915 ( \62890 , \58867 );
buf \U$62916 ( \62891 , \58874 );
buf \U$62917 ( \62892 , \59412 );
nor \U$62918 ( \62893 , \62891 , \62892 );
buf \U$62919 ( \62894 , \62893 );
buf \U$62920 ( \62895 , \62894 );
nand \U$62921 ( \62896 , \62890 , \62895 );
buf \U$62922 ( \62897 , \62896 );
buf \U$62923 ( \62898 , \62897 );
buf \U$62924 ( \62899 , \58686 );
not \U$62925 ( \62900 , \62899 );
buf \U$62926 ( \62901 , \58641 );
nand \U$62927 ( \62902 , \62900 , \62901 );
buf \U$62928 ( \62903 , \62902 );
buf \U$62929 ( \62904 , \62903 );
buf \U$62930 ( \62905 , \58864 );
not \U$62931 ( \62906 , \62905 );
buf \U$62932 ( \62907 , \58856 );
nand \U$62933 ( \62908 , \62906 , \62907 );
buf \U$62934 ( \62909 , \62908 );
buf \U$62935 ( \62910 , \62909 );
nand \U$62936 ( \62911 , \62898 , \62904 , \62910 );
buf \U$62937 ( \62912 , \62911 );
buf \U$62938 ( \62913 , \62912 );
not \U$62939 ( \62914 , \62913 );
or \U$62940 ( \62915 , \62889 , \62914 );
buf \U$62941 ( \62916 , \58715 );
not \U$62942 ( \62917 , \62916 );
buf \U$62943 ( \62918 , \58707 );
nand \U$62944 ( \62919 , \62917 , \62918 );
buf \U$62945 ( \62920 , \62919 );
buf \U$62946 ( \62921 , \62920 );
nand \U$62947 ( \62922 , \62915 , \62921 );
buf \U$62948 ( \62923 , \62922 );
buf \U$62949 ( \62924 , \62923 );
and \U$62950 ( \62925 , \62887 , \62924 );
buf \U$62951 ( \62926 , \57476 );
buf \U$62952 ( \62927 , \57850 );
nand \U$62953 ( \62928 , \62926 , \62927 );
buf \U$62954 ( \62929 , \62928 );
buf \U$62955 ( \62930 , \62929 );
not \U$62956 ( \62931 , \62930 );
buf \U$62957 ( \62932 , \57472 );
nand \U$62958 ( \62933 , \62931 , \62932 );
buf \U$62959 ( \62934 , \62933 );
buf \U$62960 ( \62935 , \62934 );
buf \U$62961 ( \62936 , \57079 );
not \U$62962 ( \62937 , \62936 );
buf \U$62963 ( \62938 , \57466 );
nand \U$62964 ( \62939 , \62937 , \62938 );
buf \U$62965 ( \62940 , \62939 );
buf \U$62966 ( \62941 , \62940 );
nand \U$62967 ( \62942 , \62935 , \62941 );
buf \U$62968 ( \62943 , \62942 );
buf \U$62969 ( \62944 , \62943 );
buf \U$62970 ( \62945 , \57943 );
buf \U$62971 ( \62946 , \57918 );
nand \U$62972 ( \62947 , \62944 , \62945 , \62946 );
buf \U$62973 ( \62948 , \62947 );
buf \U$62974 ( \62949 , \62948 );
buf \U$62975 ( \62950 , \57943 );
buf \U$62976 ( \62951 , \57915 );
buf \U$62977 ( \62952 , \57891 );
nor \U$62978 ( \62953 , \62951 , \62952 );
buf \U$62979 ( \62954 , \62953 );
buf \U$62980 ( \62955 , \62954 );
and \U$62981 ( \62956 , \62950 , \62955 );
buf \U$62982 ( \62957 , \57933 );
buf \U$62983 ( \62958 , \57940 );
nor \U$62984 ( \62959 , \62957 , \62958 );
buf \U$62985 ( \62960 , \62959 );
buf \U$62986 ( \62961 , \62960 );
nor \U$62987 ( \62962 , \62956 , \62961 );
buf \U$62988 ( \62963 , \62962 );
buf \U$62989 ( \62964 , \62963 );
nand \U$62990 ( \62965 , \62949 , \62964 );
buf \U$62991 ( \62966 , \62965 );
buf \U$62992 ( \62967 , \62966 );
nor \U$62993 ( \62968 , \62925 , \62967 );
buf \U$62994 ( \62969 , \62968 );
buf \U$62995 ( \62970 , \62969 );
nand \U$62996 ( \62971 , \62883 , \62970 );
buf \U$62997 ( \62972 , \62971 );
buf \U$62998 ( \62973 , \62972 );
and \U$62999 ( \62974 , \56474 , \56475 , \62973 );
buf \U$63000 ( \62975 , \56355 );
not \U$63001 ( \62976 , \62975 );
buf \U$63002 ( \62977 , \56423 );
not \U$63003 ( \62978 , \62977 );
buf \U$63004 ( \62979 , \56412 );
buf \U$63005 ( \62980 , \56427 );
buf \U$63006 ( \62981 , \56433 );
nand \U$63007 ( \62982 , \62980 , \62981 );
buf \U$63008 ( \62983 , \62982 );
buf \U$63009 ( \62984 , \62983 );
or \U$63010 ( \62985 , \62979 , \62984 );
buf \U$63011 ( \62986 , \56389 );
buf \U$63012 ( \62987 , \56409 );
nand \U$63013 ( \62988 , \62986 , \62987 );
buf \U$63014 ( \62989 , \62988 );
buf \U$63015 ( \62990 , \62989 );
nand \U$63016 ( \62991 , \62985 , \62990 );
buf \U$63017 ( \62992 , \62991 );
buf \U$63018 ( \62993 , \62992 );
not \U$63019 ( \62994 , \62993 );
or \U$63020 ( \62995 , \62978 , \62994 );
buf \U$63021 ( \62996 , \56422 );
not \U$63022 ( \62997 , \62996 );
buf \U$63023 ( \62998 , \56419 );
nand \U$63024 ( \62999 , \62997 , \62998 );
buf \U$63025 ( \63000 , \62999 );
buf \U$63026 ( \63001 , \63000 );
nand \U$63027 ( \63002 , \62995 , \63001 );
buf \U$63028 ( \63003 , \63002 );
buf \U$63029 ( \63004 , \63003 );
not \U$63030 ( \63005 , \63004 );
or \U$63031 ( \63006 , \62976 , \63005 );
buf \U$63032 ( \63007 , \56210 );
buf \U$63033 ( \63008 , \56352 );
nand \U$63034 ( \63009 , \63007 , \63008 );
buf \U$63035 ( \63010 , \63009 );
buf \U$63036 ( \63011 , \63010 );
nand \U$63037 ( \63012 , \63006 , \63011 );
buf \U$63038 ( \63013 , \63012 );
buf \U$63039 ( \63014 , \63013 );
nor \U$63040 ( \63015 , \62974 , \63014 );
buf \U$63041 ( \63016 , \63015 );
buf \U$63042 ( \63017 , \63016 );
nand \U$63043 ( \63018 , \56446 , \63017 );
buf \U$63044 ( \63019 , \63018 );
buf \U$63045 ( \63020 , \63019 );
not \U$63046 ( \63021 , \63020 );
buf \U$63047 ( \63022 , \6141 );
buf \U$63048 ( \63023 , RIc0d9400_64);
and \U$63049 ( \63024 , \63022 , \63023 );
buf \U$63050 ( \63025 , \63024 );
buf \U$63051 ( \63026 , \63025 );
buf \U$63052 ( \63027 , RIc0d9bf8_81);
buf \U$63053 ( \63028 , RIc0d9298_61);
xor \U$63054 ( \63029 , \63027 , \63028 );
buf \U$63055 ( \63030 , \63029 );
buf \U$63056 ( \63031 , \63030 );
not \U$63057 ( \63032 , \63031 );
buf \U$63058 ( \63033 , \17141 );
not \U$63059 ( \63034 , \63033 );
or \U$63060 ( \63035 , \63032 , \63034 );
buf \U$63061 ( \63036 , \1078 );
buf \U$63062 ( \63037 , RIc0d9bf8_81);
buf \U$63063 ( \63038 , RIc0d9220_60);
xor \U$63064 ( \63039 , \63037 , \63038 );
buf \U$63065 ( \63040 , \63039 );
buf \U$63066 ( \63041 , \63040 );
nand \U$63067 ( \63042 , \63036 , \63041 );
buf \U$63068 ( \63043 , \63042 );
buf \U$63069 ( \63044 , \63043 );
nand \U$63070 ( \63045 , \63035 , \63044 );
buf \U$63071 ( \63046 , \63045 );
buf \U$63072 ( \63047 , \63046 );
xor \U$63073 ( \63048 , \63026 , \63047 );
buf \U$63074 ( \63049 , RIc0dadc8_119);
buf \U$63075 ( \63050 , RIc0d80c8_23);
xor \U$63076 ( \63051 , \63049 , \63050 );
buf \U$63077 ( \63052 , \63051 );
buf \U$63078 ( \63053 , \63052 );
not \U$63079 ( \63054 , \63053 );
buf \U$63080 ( \63055 , \23985 );
not \U$63081 ( \63056 , \63055 );
or \U$63082 ( \63057 , \63054 , \63056 );
buf \U$63083 ( \63058 , \13005 );
xor \U$63084 ( \63059 , RIc0dadc8_119, RIc0d8050_22);
buf \U$63085 ( \63060 , \63059 );
nand \U$63086 ( \63061 , \63058 , \63060 );
buf \U$63087 ( \63062 , \63061 );
buf \U$63088 ( \63063 , \63062 );
nand \U$63089 ( \63064 , \63057 , \63063 );
buf \U$63090 ( \63065 , \63064 );
buf \U$63091 ( \63066 , \63065 );
xor \U$63092 ( \63067 , \63048 , \63066 );
buf \U$63093 ( \63068 , \63067 );
buf \U$63094 ( \63069 , \63068 );
buf \U$63095 ( \63070 , RIc0d7d08_15);
buf \U$63096 ( \63071 , RIc0db188_127);
xor \U$63097 ( \63072 , \63070 , \63071 );
buf \U$63098 ( \63073 , \63072 );
buf \U$63099 ( \63074 , \63073 );
not \U$63100 ( \63075 , \63074 );
buf \U$63101 ( \63076 , \15609 );
not \U$63102 ( \63077 , \63076 );
or \U$63103 ( \63078 , \63075 , \63077 );
buf \U$63104 ( \63079 , RIc0d7c90_14);
buf \U$63105 ( \63080 , RIc0db188_127);
xor \U$63106 ( \63081 , \63079 , \63080 );
buf \U$63107 ( \63082 , \63081 );
buf \U$63108 ( \63083 , \63082 );
buf \U$63109 ( \63084 , RIc0db200_128);
nand \U$63110 ( \63085 , \63083 , \63084 );
buf \U$63111 ( \63086 , \63085 );
buf \U$63112 ( \63087 , \63086 );
nand \U$63113 ( \63088 , \63078 , \63087 );
buf \U$63114 ( \63089 , \63088 );
buf \U$63115 ( \63090 , \63089 );
buf \U$63116 ( \63091 , RIc0d9fb8_89);
buf \U$63117 ( \63092 , RIc0d8ed8_53);
xor \U$63118 ( \63093 , \63091 , \63092 );
buf \U$63119 ( \63094 , \63093 );
buf \U$63120 ( \63095 , \63094 );
not \U$63121 ( \63096 , \63095 );
buf \U$63122 ( \63097 , \18150 );
not \U$63123 ( \63098 , \63097 );
or \U$63124 ( \63099 , \63096 , \63098 );
buf \U$63125 ( \63100 , \846 );
buf \U$63126 ( \63101 , RIc0d9fb8_89);
buf \U$63127 ( \63102 , RIc0d8e60_52);
xor \U$63128 ( \63103 , \63101 , \63102 );
buf \U$63129 ( \63104 , \63103 );
buf \U$63130 ( \63105 , \63104 );
nand \U$63131 ( \63106 , \63100 , \63105 );
buf \U$63132 ( \63107 , \63106 );
buf \U$63133 ( \63108 , \63107 );
nand \U$63134 ( \63109 , \63099 , \63108 );
buf \U$63135 ( \63110 , \63109 );
buf \U$63136 ( \63111 , \63110 );
xor \U$63137 ( \63112 , \63090 , \63111 );
xor \U$63138 ( \63113 , RIc0da0a8_91, RIc0d8de8_51);
buf \U$63139 ( \63114 , \63113 );
not \U$63140 ( \63115 , \63114 );
buf \U$63141 ( \63116 , \524 );
not \U$63142 ( \63117 , \63116 );
or \U$63143 ( \63118 , \63115 , \63117 );
buf \U$63144 ( \63119 , \13293 );
buf \U$63145 ( \63120 , RIc0d8d70_50);
buf \U$63146 ( \63121 , RIc0da0a8_91);
xor \U$63147 ( \63122 , \63120 , \63121 );
buf \U$63148 ( \63123 , \63122 );
buf \U$63149 ( \63124 , \63123 );
nand \U$63150 ( \63125 , \63119 , \63124 );
buf \U$63151 ( \63126 , \63125 );
buf \U$63152 ( \63127 , \63126 );
nand \U$63153 ( \63128 , \63118 , \63127 );
buf \U$63154 ( \63129 , \63128 );
buf \U$63155 ( \63130 , \63129 );
xor \U$63156 ( \63131 , \63112 , \63130 );
buf \U$63157 ( \63132 , \63131 );
buf \U$63158 ( \63133 , \63132 );
nor \U$63159 ( \63134 , \63069 , \63133 );
buf \U$63160 ( \63135 , \63134 );
buf \U$63161 ( \63136 , \63135 );
buf \U$63162 ( \63137 , RIc0dabe8_115);
buf \U$63163 ( \63138 , RIc0d82a8_27);
xor \U$63164 ( \63139 , \63137 , \63138 );
buf \U$63165 ( \63140 , \63139 );
buf \U$63166 ( \63141 , \63140 );
not \U$63167 ( \63142 , \63141 );
buf \U$63168 ( \63143 , \14186 );
not \U$63169 ( \63144 , \63143 );
or \U$63170 ( \63145 , \63142 , \63144 );
buf \U$63171 ( \63146 , \14690 );
buf \U$63172 ( \63147 , RIc0dabe8_115);
buf \U$63173 ( \63148 , RIc0d8230_26);
xor \U$63174 ( \63149 , \63147 , \63148 );
buf \U$63175 ( \63150 , \63149 );
buf \U$63176 ( \63151 , \63150 );
nand \U$63177 ( \63152 , \63146 , \63151 );
buf \U$63178 ( \63153 , \63152 );
buf \U$63179 ( \63154 , \63153 );
nand \U$63180 ( \63155 , \63145 , \63154 );
buf \U$63181 ( \63156 , \63155 );
buf \U$63182 ( \63157 , RIc0da558_101);
buf \U$63183 ( \63158 , RIc0d8938_41);
xor \U$63184 ( \63159 , \63157 , \63158 );
buf \U$63185 ( \63160 , \63159 );
buf \U$63186 ( \63161 , \63160 );
not \U$63187 ( \63162 , \63161 );
buf \U$63188 ( \63163 , \22631 );
not \U$63189 ( \63164 , \63163 );
or \U$63190 ( \63165 , \63162 , \63164 );
buf \U$63191 ( \63166 , \26354 );
xor \U$63192 ( \63167 , RIc0da558_101, RIc0d88c0_40);
buf \U$63193 ( \63168 , \63167 );
nand \U$63194 ( \63169 , \63166 , \63168 );
buf \U$63195 ( \63170 , \63169 );
buf \U$63196 ( \63171 , \63170 );
nand \U$63197 ( \63172 , \63165 , \63171 );
buf \U$63198 ( \63173 , \63172 );
xor \U$63199 ( \63174 , \63156 , \63173 );
xor \U$63200 ( \63175 , RIc0d9ec8_87, RIc0d8fc8_55);
buf \U$63201 ( \63176 , \63175 );
not \U$63202 ( \63177 , \63176 );
buf \U$63203 ( \63178 , \4527 );
not \U$63204 ( \63179 , \63178 );
or \U$63205 ( \63180 , \63177 , \63179 );
buf \U$63206 ( \63181 , \816 );
buf \U$63207 ( \63182 , RIc0d8f50_54);
buf \U$63208 ( \63183 , RIc0d9ec8_87);
xor \U$63209 ( \63184 , \63182 , \63183 );
buf \U$63210 ( \63185 , \63184 );
buf \U$63211 ( \63186 , \63185 );
nand \U$63212 ( \63187 , \63181 , \63186 );
buf \U$63213 ( \63188 , \63187 );
buf \U$63214 ( \63189 , \63188 );
nand \U$63215 ( \63190 , \63180 , \63189 );
buf \U$63216 ( \63191 , \63190 );
xnor \U$63217 ( \63192 , \63174 , \63191 );
buf \U$63218 ( \63193 , \63192 );
or \U$63219 ( \63194 , \63136 , \63193 );
buf \U$63220 ( \63195 , \63068 );
buf \U$63221 ( \63196 , \63132 );
nand \U$63222 ( \63197 , \63195 , \63196 );
buf \U$63223 ( \63198 , \63197 );
buf \U$63224 ( \63199 , \63198 );
nand \U$63225 ( \63200 , \63194 , \63199 );
buf \U$63226 ( \63201 , \63200 );
buf \U$63227 ( \63202 , \63201 );
buf \U$63228 ( \63203 , RIc0d8b18_45);
buf \U$63229 ( \63204 , RIc0da378_97);
xor \U$63230 ( \63205 , \63203 , \63204 );
buf \U$63231 ( \63206 , \63205 );
buf \U$63232 ( \63207 , \63206 );
not \U$63233 ( \63208 , \63207 );
buf \U$63234 ( \63209 , \2066 );
not \U$63235 ( \63210 , \63209 );
or \U$63236 ( \63211 , \63208 , \63210 );
buf \U$63237 ( \63212 , \2070 );
buf \U$63238 ( \63213 , RIc0da378_97);
buf \U$63239 ( \63214 , RIc0d8aa0_44);
xor \U$63240 ( \63215 , \63213 , \63214 );
buf \U$63241 ( \63216 , \63215 );
buf \U$63242 ( \63217 , \63216 );
nand \U$63243 ( \63218 , \63212 , \63217 );
buf \U$63244 ( \63219 , \63218 );
buf \U$63245 ( \63220 , \63219 );
nand \U$63246 ( \63221 , \63211 , \63220 );
buf \U$63247 ( \63222 , \63221 );
buf \U$63248 ( \63223 , \63222 );
buf \U$63249 ( \63224 , RIc0d9ce8_83);
buf \U$63250 ( \63225 , RIc0d91a8_59);
xor \U$63251 ( \63226 , \63224 , \63225 );
buf \U$63252 ( \63227 , \63226 );
buf \U$63253 ( \63228 , \63227 );
not \U$63254 ( \63229 , \63228 );
buf \U$63255 ( \63230 , \1736 );
not \U$63256 ( \63231 , \63230 );
or \U$63257 ( \63232 , \63229 , \63231 );
buf \U$63258 ( \63233 , \993 );
buf \U$63259 ( \63234 , RIc0d9ce8_83);
buf \U$63260 ( \63235 , RIc0d9130_58);
xor \U$63261 ( \63236 , \63234 , \63235 );
buf \U$63262 ( \63237 , \63236 );
buf \U$63263 ( \63238 , \63237 );
nand \U$63264 ( \63239 , \63233 , \63238 );
buf \U$63265 ( \63240 , \63239 );
buf \U$63266 ( \63241 , \63240 );
nand \U$63267 ( \63242 , \63232 , \63241 );
buf \U$63268 ( \63243 , \63242 );
buf \U$63269 ( \63244 , \63243 );
or \U$63270 ( \63245 , \63223 , \63244 );
buf \U$63271 ( \63246 , RIc0daeb8_121);
buf \U$63272 ( \63247 , RIc0d7fd8_21);
xor \U$63273 ( \63248 , \63246 , \63247 );
buf \U$63274 ( \63249 , \63248 );
buf \U$63275 ( \63250 , \63249 );
not \U$63276 ( \63251 , \63250 );
buf \U$63277 ( \63252 , \24672 );
not \U$63278 ( \63253 , \63252 );
or \U$63279 ( \63254 , \63251 , \63253 );
buf \U$63280 ( \63255 , \16386 );
xor \U$63281 ( \63256 , RIc0daeb8_121, RIc0d7f60_20);
buf \U$63282 ( \63257 , \63256 );
nand \U$63283 ( \63258 , \63255 , \63257 );
buf \U$63284 ( \63259 , \63258 );
buf \U$63285 ( \63260 , \63259 );
nand \U$63286 ( \63261 , \63254 , \63260 );
buf \U$63287 ( \63262 , \63261 );
buf \U$63288 ( \63263 , \63262 );
nand \U$63289 ( \63264 , \63245 , \63263 );
buf \U$63290 ( \63265 , \63264 );
buf \U$63291 ( \63266 , \63265 );
buf \U$63292 ( \63267 , \63222 );
buf \U$63293 ( \63268 , \63243 );
nand \U$63294 ( \63269 , \63267 , \63268 );
buf \U$63295 ( \63270 , \63269 );
buf \U$63296 ( \63271 , \63270 );
nand \U$63297 ( \63272 , \63266 , \63271 );
buf \U$63298 ( \63273 , \63272 );
buf \U$63299 ( \63274 , \63273 );
xor \U$63300 ( \63275 , \63026 , \63047 );
and \U$63301 ( \63276 , \63275 , \63066 );
and \U$63302 ( \63277 , \63026 , \63047 );
or \U$63303 ( \63278 , \63276 , \63277 );
buf \U$63304 ( \63279 , \63278 );
buf \U$63305 ( \63280 , \63279 );
xor \U$63306 ( \63281 , \63274 , \63280 );
buf \U$63307 ( \63282 , \63191 );
not \U$63308 ( \63283 , \63282 );
buf \U$63309 ( \63284 , \63173 );
not \U$63310 ( \63285 , \63284 );
or \U$63311 ( \63286 , \63283 , \63285 );
buf \U$63312 ( \63287 , \63173 );
buf \U$63313 ( \63288 , \63191 );
or \U$63314 ( \63289 , \63287 , \63288 );
buf \U$63315 ( \63290 , \63156 );
nand \U$63316 ( \63291 , \63289 , \63290 );
buf \U$63317 ( \63292 , \63291 );
buf \U$63318 ( \63293 , \63292 );
nand \U$63319 ( \63294 , \63286 , \63293 );
buf \U$63320 ( \63295 , \63294 );
buf \U$63321 ( \63296 , \63295 );
xor \U$63322 ( \63297 , \63281 , \63296 );
buf \U$63323 ( \63298 , \63297 );
buf \U$63324 ( \63299 , \63298 );
xor \U$63325 ( \63300 , \63202 , \63299 );
xor \U$63326 ( \63301 , RIc0da738_105, RIc0d8758_37);
buf \U$63327 ( \63302 , \63301 );
not \U$63328 ( \63303 , \63302 );
buf \U$63329 ( \63304 , \12736 );
not \U$63330 ( \63305 , \63304 );
or \U$63331 ( \63306 , \63303 , \63305 );
buf \U$63332 ( \63307 , \12744 );
buf \U$63333 ( \63308 , RIc0da738_105);
buf \U$63334 ( \63309 , RIc0d86e0_36);
xor \U$63335 ( \63310 , \63308 , \63309 );
buf \U$63336 ( \63311 , \63310 );
buf \U$63337 ( \63312 , \63311 );
nand \U$63338 ( \63313 , \63307 , \63312 );
buf \U$63339 ( \63314 , \63313 );
buf \U$63340 ( \63315 , \63314 );
nand \U$63341 ( \63316 , \63306 , \63315 );
buf \U$63342 ( \63317 , \63316 );
buf \U$63343 ( \63318 , \63317 );
not \U$63344 ( \63319 , \63318 );
buf \U$63345 ( \63320 , RIc0d8398_29);
buf \U$63346 ( \63321 , RIc0daaf8_113);
xor \U$63347 ( \63322 , \63320 , \63321 );
buf \U$63348 ( \63323 , \63322 );
buf \U$63349 ( \63324 , \63323 );
not \U$63350 ( \63325 , \63324 );
buf \U$63351 ( \63326 , \25355 );
not \U$63352 ( \63327 , \63326 );
or \U$63353 ( \63328 , \63325 , \63327 );
buf \U$63354 ( \63329 , \16995 );
buf \U$63355 ( \63330 , RIc0daaf8_113);
buf \U$63356 ( \63331 , RIc0d8320_28);
xor \U$63357 ( \63332 , \63330 , \63331 );
buf \U$63358 ( \63333 , \63332 );
buf \U$63359 ( \63334 , \63333 );
nand \U$63360 ( \63335 , \63329 , \63334 );
buf \U$63361 ( \63336 , \63335 );
buf \U$63362 ( \63337 , \63336 );
nand \U$63363 ( \63338 , \63328 , \63337 );
buf \U$63364 ( \63339 , \63338 );
buf \U$63365 ( \63340 , \63339 );
not \U$63366 ( \63341 , \63340 );
or \U$63367 ( \63342 , \63319 , \63341 );
buf \U$63368 ( \63343 , \63339 );
buf \U$63369 ( \63344 , \63317 );
or \U$63370 ( \63345 , \63343 , \63344 );
xor \U$63371 ( \63346 , RIc0da468_99, RIc0d8a28_43);
buf \U$63372 ( \63347 , \63346 );
not \U$63373 ( \63348 , \63347 );
buf \U$63374 ( \63349 , \19695 );
not \U$63375 ( \63350 , \63349 );
or \U$63376 ( \63351 , \63348 , \63350 );
buf \U$63377 ( \63352 , \16750 );
buf \U$63378 ( \63353 , RIc0da468_99);
buf \U$63379 ( \63354 , RIc0d89b0_42);
xor \U$63380 ( \63355 , \63353 , \63354 );
buf \U$63381 ( \63356 , \63355 );
buf \U$63382 ( \63357 , \63356 );
nand \U$63383 ( \63358 , \63352 , \63357 );
buf \U$63384 ( \63359 , \63358 );
buf \U$63385 ( \63360 , \63359 );
nand \U$63386 ( \63361 , \63351 , \63360 );
buf \U$63387 ( \63362 , \63361 );
buf \U$63388 ( \63363 , \63362 );
nand \U$63389 ( \63364 , \63345 , \63363 );
buf \U$63390 ( \63365 , \63364 );
buf \U$63391 ( \63366 , \63365 );
nand \U$63392 ( \63367 , \63342 , \63366 );
buf \U$63393 ( \63368 , \63367 );
buf \U$63394 ( \63369 , \63368 );
buf \U$63395 ( \63370 , RIc0d9b08_79);
buf \U$63396 ( \63371 , RIc0d9388_63);
xor \U$63397 ( \63372 , \63370 , \63371 );
buf \U$63398 ( \63373 , \63372 );
buf \U$63399 ( \63374 , \63373 );
not \U$63400 ( \63375 , \63374 );
buf \U$63401 ( \63376 , \14940 );
not \U$63402 ( \63377 , \63376 );
or \U$63403 ( \63378 , \63375 , \63377 );
buf \U$63404 ( \63379 , \1025 );
xor \U$63405 ( \63380 , RIc0d9b08_79, RIc0d9310_62);
buf \U$63406 ( \63381 , \63380 );
nand \U$63407 ( \63382 , \63379 , \63381 );
buf \U$63408 ( \63383 , \63382 );
buf \U$63409 ( \63384 , \63383 );
nand \U$63410 ( \63385 , \63378 , \63384 );
buf \U$63411 ( \63386 , \63385 );
not \U$63412 ( \63387 , \63386 );
buf \U$63413 ( \63388 , RIc0d9dd8_85);
buf \U$63414 ( \63389 , RIc0d90b8_57);
xor \U$63415 ( \63390 , \63388 , \63389 );
buf \U$63416 ( \63391 , \63390 );
buf \U$63417 ( \63392 , \63391 );
not \U$63418 ( \63393 , \63392 );
buf \U$63419 ( \63394 , \5304 );
not \U$63420 ( \63395 , \63394 );
or \U$63421 ( \63396 , \63393 , \63395 );
buf \U$63422 ( \63397 , \1401 );
xor \U$63423 ( \63398 , RIc0d9dd8_85, RIc0d9040_56);
buf \U$63424 ( \63399 , \63398 );
nand \U$63425 ( \63400 , \63397 , \63399 );
buf \U$63426 ( \63401 , \63400 );
buf \U$63427 ( \63402 , \63401 );
nand \U$63428 ( \63403 , \63396 , \63402 );
buf \U$63429 ( \63404 , \63403 );
not \U$63430 ( \63405 , \63404 );
or \U$63431 ( \63406 , \63387 , \63405 );
buf \U$63432 ( \63407 , \63386 );
buf \U$63433 ( \63408 , \63404 );
or \U$63434 ( \63409 , \63407 , \63408 );
buf \U$63435 ( \63410 , RIc0daa08_111);
buf \U$63436 ( \63411 , RIc0d8488_31);
xor \U$63437 ( \63412 , \63410 , \63411 );
buf \U$63438 ( \63413 , \63412 );
buf \U$63439 ( \63414 , \63413 );
not \U$63440 ( \63415 , \63414 );
buf \U$63441 ( \63416 , \14346 );
not \U$63442 ( \63417 , \63416 );
or \U$63443 ( \63418 , \63415 , \63417 );
buf \U$63444 ( \63419 , \15864 );
xor \U$63445 ( \63420 , RIc0daa08_111, RIc0d8410_30);
buf \U$63446 ( \63421 , \63420 );
nand \U$63447 ( \63422 , \63419 , \63421 );
buf \U$63448 ( \63423 , \63422 );
buf \U$63449 ( \63424 , \63423 );
nand \U$63450 ( \63425 , \63418 , \63424 );
buf \U$63451 ( \63426 , \63425 );
buf \U$63452 ( \63427 , \63426 );
nand \U$63453 ( \63428 , \63409 , \63427 );
buf \U$63454 ( \63429 , \63428 );
nand \U$63455 ( \63430 , \63406 , \63429 );
buf \U$63456 ( \63431 , \63430 );
xor \U$63457 ( \63432 , \63369 , \63431 );
xor \U$63458 ( \63433 , RIc0da828_107, RIc0d8668_35);
buf \U$63459 ( \63434 , \63433 );
not \U$63460 ( \63435 , \63434 );
buf \U$63461 ( \63436 , \12334 );
not \U$63462 ( \63437 , \63436 );
or \U$63463 ( \63438 , \63435 , \63437 );
buf \U$63464 ( \63439 , \12342 );
buf \U$63465 ( \63440 , RIc0da828_107);
buf \U$63466 ( \63441 , RIc0d85f0_34);
xor \U$63467 ( \63442 , \63440 , \63441 );
buf \U$63468 ( \63443 , \63442 );
buf \U$63469 ( \63444 , \63443 );
nand \U$63470 ( \63445 , \63439 , \63444 );
buf \U$63471 ( \63446 , \63445 );
buf \U$63472 ( \63447 , \63446 );
nand \U$63473 ( \63448 , \63438 , \63447 );
buf \U$63474 ( \63449 , \63448 );
buf \U$63475 ( \63450 , \63449 );
buf \U$63476 ( \63451 , RIc0da198_93);
buf \U$63477 ( \63452 , RIc0d8cf8_49);
xor \U$63478 ( \63453 , \63451 , \63452 );
buf \U$63479 ( \63454 , \63453 );
buf \U$63480 ( \63455 , \63454 );
not \U$63481 ( \63456 , \63455 );
buf \U$63482 ( \63457 , \476 );
not \U$63483 ( \63458 , \63457 );
or \U$63484 ( \63459 , \63456 , \63458 );
buf \U$63485 ( \63460 , \4008 );
xor \U$63486 ( \63461 , RIc0da198_93, RIc0d8c80_48);
buf \U$63487 ( \63462 , \63461 );
nand \U$63488 ( \63463 , \63460 , \63462 );
buf \U$63489 ( \63464 , \63463 );
buf \U$63490 ( \63465 , \63464 );
nand \U$63491 ( \63466 , \63459 , \63465 );
buf \U$63492 ( \63467 , \63466 );
buf \U$63493 ( \63468 , \63467 );
or \U$63494 ( \63469 , \63450 , \63468 );
xor \U$63495 ( \63470 , RIc0dafa8_123, RIc0d7ee8_19);
buf \U$63496 ( \63471 , \63470 );
not \U$63497 ( \63472 , \63471 );
buf \U$63498 ( \63473 , \14982 );
not \U$63499 ( \63474 , \63473 );
or \U$63500 ( \63475 , \63472 , \63474 );
buf \U$63501 ( \63476 , \16692 );
buf \U$63502 ( \63477 , RIc0dafa8_123);
buf \U$63503 ( \63478 , RIc0d7e70_18);
xor \U$63504 ( \63479 , \63477 , \63478 );
buf \U$63505 ( \63480 , \63479 );
buf \U$63506 ( \63481 , \63480 );
nand \U$63507 ( \63482 , \63476 , \63481 );
buf \U$63508 ( \63483 , \63482 );
buf \U$63509 ( \63484 , \63483 );
nand \U$63510 ( \63485 , \63475 , \63484 );
buf \U$63511 ( \63486 , \63485 );
buf \U$63512 ( \63487 , \63486 );
nand \U$63513 ( \63488 , \63469 , \63487 );
buf \U$63514 ( \63489 , \63488 );
buf \U$63515 ( \63490 , \63489 );
buf \U$63516 ( \63491 , \63449 );
buf \U$63517 ( \63492 , \63467 );
nand \U$63518 ( \63493 , \63491 , \63492 );
buf \U$63519 ( \63494 , \63493 );
buf \U$63520 ( \63495 , \63494 );
nand \U$63521 ( \63496 , \63490 , \63495 );
buf \U$63522 ( \63497 , \63496 );
buf \U$63523 ( \63498 , \63497 );
xor \U$63524 ( \63499 , \63432 , \63498 );
buf \U$63525 ( \63500 , \63499 );
buf \U$63526 ( \63501 , \63500 );
xor \U$63527 ( \63502 , \63300 , \63501 );
buf \U$63528 ( \63503 , \63502 );
buf \U$63529 ( \63504 , \63503 );
xor \U$63530 ( \63505 , RIc0da0a8_91, RIc0d8e60_52);
buf \U$63531 ( \63506 , \63505 );
not \U$63532 ( \63507 , \63506 );
buf \U$63533 ( \63508 , \704 );
not \U$63534 ( \63509 , \63508 );
or \U$63535 ( \63510 , \63507 , \63509 );
buf \U$63536 ( \63511 , \533 );
buf \U$63537 ( \63512 , \63113 );
nand \U$63538 ( \63513 , \63511 , \63512 );
buf \U$63539 ( \63514 , \63513 );
buf \U$63540 ( \63515 , \63514 );
nand \U$63541 ( \63516 , \63510 , \63515 );
buf \U$63542 ( \63517 , \63516 );
buf \U$63543 ( \63518 , \63517 );
buf \U$63544 ( \63519 , RIc0d9ec8_87);
buf \U$63545 ( \63520 , RIc0d9040_56);
xor \U$63546 ( \63521 , \63519 , \63520 );
buf \U$63547 ( \63522 , \63521 );
buf \U$63548 ( \63523 , \63522 );
not \U$63549 ( \63524 , \63523 );
buf \U$63550 ( \63525 , \2607 );
not \U$63551 ( \63526 , \63525 );
or \U$63552 ( \63527 , \63524 , \63526 );
buf \U$63553 ( \63528 , \3631 );
buf \U$63554 ( \63529 , \63175 );
nand \U$63555 ( \63530 , \63528 , \63529 );
buf \U$63556 ( \63531 , \63530 );
buf \U$63557 ( \63532 , \63531 );
nand \U$63558 ( \63533 , \63527 , \63532 );
buf \U$63559 ( \63534 , \63533 );
buf \U$63560 ( \63535 , \63534 );
xor \U$63561 ( \63536 , \63518 , \63535 );
buf \U$63562 ( \63537 , RIc0dabe8_115);
buf \U$63563 ( \63538 , RIc0d8320_28);
xor \U$63564 ( \63539 , \63537 , \63538 );
buf \U$63565 ( \63540 , \63539 );
buf \U$63566 ( \63541 , \63540 );
not \U$63567 ( \63542 , \63541 );
buf \U$63568 ( \63543 , \26466 );
not \U$63569 ( \63544 , \63543 );
or \U$63570 ( \63545 , \63542 , \63544 );
buf \U$63571 ( \63546 , \12303 );
buf \U$63572 ( \63547 , \63140 );
nand \U$63573 ( \63548 , \63546 , \63547 );
buf \U$63574 ( \63549 , \63548 );
buf \U$63575 ( \63550 , \63549 );
nand \U$63576 ( \63551 , \63545 , \63550 );
buf \U$63577 ( \63552 , \63551 );
buf \U$63578 ( \63553 , \63552 );
and \U$63579 ( \63554 , \63536 , \63553 );
and \U$63580 ( \63555 , \63518 , \63535 );
or \U$63581 ( \63556 , \63554 , \63555 );
buf \U$63582 ( \63557 , \63556 );
buf \U$63583 ( \63558 , \63557 );
buf \U$63584 ( \63559 , RIc0d7d80_16);
buf \U$63585 ( \63560 , RIc0db188_127);
xor \U$63586 ( \63561 , \63559 , \63560 );
buf \U$63587 ( \63562 , \63561 );
buf \U$63588 ( \63563 , \63562 );
not \U$63589 ( \63564 , \63563 );
buf \U$63590 ( \63565 , \43780 );
not \U$63591 ( \63566 , \63565 );
or \U$63592 ( \63567 , \63564 , \63566 );
buf \U$63593 ( \63568 , \63073 );
buf \U$63594 ( \63569 , RIc0db200_128);
nand \U$63595 ( \63570 , \63568 , \63569 );
buf \U$63596 ( \63571 , \63570 );
buf \U$63597 ( \63572 , \63571 );
nand \U$63598 ( \63573 , \63567 , \63572 );
buf \U$63599 ( \63574 , \63573 );
buf \U$63600 ( \63575 , \63574 );
buf \U$63601 ( \63576 , RIc0d9fb8_89);
buf \U$63602 ( \63577 , RIc0d8f50_54);
xor \U$63603 ( \63578 , \63576 , \63577 );
buf \U$63604 ( \63579 , \63578 );
buf \U$63605 ( \63580 , \63579 );
not \U$63606 ( \63581 , \63580 );
buf \U$63607 ( \63582 , \437 );
not \U$63608 ( \63583 , \63582 );
or \U$63609 ( \63584 , \63581 , \63583 );
buf \U$63610 ( \63585 , \846 );
buf \U$63611 ( \63586 , \63094 );
nand \U$63612 ( \63587 , \63585 , \63586 );
buf \U$63613 ( \63588 , \63587 );
buf \U$63614 ( \63589 , \63588 );
nand \U$63615 ( \63590 , \63584 , \63589 );
buf \U$63616 ( \63591 , \63590 );
buf \U$63617 ( \63592 , \63591 );
or \U$63618 ( \63593 , \63575 , \63592 );
buf \U$63619 ( \63594 , RIc0da738_105);
buf \U$63620 ( \63595 , RIc0d87d0_38);
xor \U$63621 ( \63596 , \63594 , \63595 );
buf \U$63622 ( \63597 , \63596 );
buf \U$63623 ( \63598 , \63597 );
not \U$63624 ( \63599 , \63598 );
buf \U$63625 ( \63600 , \12736 );
not \U$63626 ( \63601 , \63600 );
or \U$63627 ( \63602 , \63599 , \63601 );
buf \U$63628 ( \63603 , \26301 );
buf \U$63629 ( \63604 , \63301 );
nand \U$63630 ( \63605 , \63603 , \63604 );
buf \U$63631 ( \63606 , \63605 );
buf \U$63632 ( \63607 , \63606 );
nand \U$63633 ( \63608 , \63602 , \63607 );
buf \U$63634 ( \63609 , \63608 );
buf \U$63635 ( \63610 , \63609 );
nand \U$63636 ( \63611 , \63593 , \63610 );
buf \U$63637 ( \63612 , \63611 );
buf \U$63638 ( \63613 , \63612 );
buf \U$63639 ( \63614 , \63591 );
buf \U$63640 ( \63615 , \63574 );
nand \U$63641 ( \63616 , \63614 , \63615 );
buf \U$63642 ( \63617 , \63616 );
buf \U$63643 ( \63618 , \63617 );
nand \U$63644 ( \63619 , \63613 , \63618 );
buf \U$63645 ( \63620 , \63619 );
buf \U$63646 ( \63621 , \63620 );
or \U$63647 ( \63622 , \63558 , \63621 );
buf \U$63648 ( \63623 , \63386 );
buf \U$63649 ( \63624 , \63404 );
xor \U$63650 ( \63625 , \63623 , \63624 );
buf \U$63651 ( \63626 , \63426 );
xor \U$63652 ( \63627 , \63625 , \63626 );
buf \U$63653 ( \63628 , \63627 );
buf \U$63654 ( \63629 , \63628 );
nand \U$63655 ( \63630 , \63622 , \63629 );
buf \U$63656 ( \63631 , \63630 );
buf \U$63657 ( \63632 , \63631 );
buf \U$63658 ( \63633 , \63557 );
buf \U$63659 ( \63634 , \63620 );
nand \U$63660 ( \63635 , \63633 , \63634 );
buf \U$63661 ( \63636 , \63635 );
buf \U$63662 ( \63637 , \63636 );
nand \U$63663 ( \63638 , \63632 , \63637 );
buf \U$63664 ( \63639 , \63638 );
buf \U$63665 ( \63640 , \63639 );
xor \U$63666 ( \63641 , RIc0da198_93, RIc0d8d70_50);
buf \U$63667 ( \63642 , \63641 );
not \U$63668 ( \63643 , \63642 );
buf \U$63669 ( \63644 , \3415 );
not \U$63670 ( \63645 , \63644 );
or \U$63671 ( \63646 , \63643 , \63645 );
buf \U$63672 ( \63647 , \4008 );
buf \U$63673 ( \63648 , \63454 );
nand \U$63674 ( \63649 , \63647 , \63648 );
buf \U$63675 ( \63650 , \63649 );
buf \U$63676 ( \63651 , \63650 );
nand \U$63677 ( \63652 , \63646 , \63651 );
buf \U$63678 ( \63653 , \63652 );
buf \U$63679 ( \63654 , \63653 );
buf \U$63680 ( \63655 , RIc0da828_107);
buf \U$63681 ( \63656 , RIc0d86e0_36);
xor \U$63682 ( \63657 , \63655 , \63656 );
buf \U$63683 ( \63658 , \63657 );
buf \U$63684 ( \63659 , \63658 );
not \U$63685 ( \63660 , \63659 );
buf \U$63686 ( \63661 , \17595 );
not \U$63687 ( \63662 , \63661 );
or \U$63688 ( \63663 , \63660 , \63662 );
buf \U$63689 ( \63664 , \12342 );
buf \U$63690 ( \63665 , \63433 );
nand \U$63691 ( \63666 , \63664 , \63665 );
buf \U$63692 ( \63667 , \63666 );
buf \U$63693 ( \63668 , \63667 );
nand \U$63694 ( \63669 , \63663 , \63668 );
buf \U$63695 ( \63670 , \63669 );
buf \U$63696 ( \63671 , \63670 );
nor \U$63697 ( \63672 , \63654 , \63671 );
buf \U$63698 ( \63673 , \63672 );
buf \U$63699 ( \63674 , \63673 );
buf \U$63700 ( \63675 , RIc0daeb8_121);
buf \U$63701 ( \63676 , RIc0d8050_22);
xor \U$63702 ( \63677 , \63675 , \63676 );
buf \U$63703 ( \63678 , \63677 );
buf \U$63704 ( \63679 , \63678 );
not \U$63705 ( \63680 , \63679 );
buf \U$63706 ( \63681 , \16382 );
not \U$63707 ( \63682 , \63681 );
or \U$63708 ( \63683 , \63680 , \63682 );
buf \U$63709 ( \63684 , \13314 );
buf \U$63710 ( \63685 , \63249 );
nand \U$63711 ( \63686 , \63684 , \63685 );
buf \U$63712 ( \63687 , \63686 );
buf \U$63713 ( \63688 , \63687 );
nand \U$63714 ( \63689 , \63683 , \63688 );
buf \U$63715 ( \63690 , \63689 );
buf \U$63716 ( \63691 , \63690 );
not \U$63717 ( \63692 , \63691 );
buf \U$63718 ( \63693 , \63692 );
buf \U$63719 ( \63694 , \63693 );
or \U$63720 ( \63695 , \63674 , \63694 );
buf \U$63721 ( \63696 , \63653 );
buf \U$63722 ( \63697 , \63670 );
nand \U$63723 ( \63698 , \63696 , \63697 );
buf \U$63724 ( \63699 , \63698 );
buf \U$63725 ( \63700 , \63699 );
nand \U$63726 ( \63701 , \63695 , \63700 );
buf \U$63727 ( \63702 , \63701 );
buf \U$63728 ( \63703 , \63702 );
buf \U$63729 ( \63704 , RIc0d8aa0_44);
buf \U$63730 ( \63705 , RIc0da468_99);
xor \U$63731 ( \63706 , \63704 , \63705 );
buf \U$63732 ( \63707 , \63706 );
buf \U$63733 ( \63708 , \63707 );
not \U$63734 ( \63709 , \63708 );
buf \U$63735 ( \63710 , \21461 );
not \U$63736 ( \63711 , \63710 );
or \U$63737 ( \63712 , \63709 , \63711 );
buf \U$63738 ( \63713 , \16750 );
buf \U$63739 ( \63714 , \63346 );
nand \U$63740 ( \63715 , \63713 , \63714 );
buf \U$63741 ( \63716 , \63715 );
buf \U$63742 ( \63717 , \63716 );
nand \U$63743 ( \63718 , \63712 , \63717 );
buf \U$63744 ( \63719 , \63718 );
buf \U$63745 ( \63720 , \63719 );
xnor \U$63746 ( \63721 , RIc0dafa8_123, RIc0d7f60_20);
buf \U$63747 ( \63722 , \63721 );
not \U$63748 ( \63723 , \63722 );
buf \U$63749 ( \63724 , \63723 );
buf \U$63750 ( \63725 , \63724 );
not \U$63751 ( \63726 , \63725 );
buf \U$63752 ( \63727 , \14982 );
not \U$63753 ( \63728 , \63727 );
or \U$63754 ( \63729 , \63726 , \63728 );
buf \U$63755 ( \63730 , \16692 );
buf \U$63756 ( \63731 , \63470 );
nand \U$63757 ( \63732 , \63730 , \63731 );
buf \U$63758 ( \63733 , \63732 );
buf \U$63759 ( \63734 , \63733 );
nand \U$63760 ( \63735 , \63729 , \63734 );
buf \U$63761 ( \63736 , \63735 );
buf \U$63763 ( \63737 , \63736 );
xor \U$63764 ( \63738 , \63720 , \63737 );
buf \U$63765 ( \63739 , RIc0daaf8_113);
buf \U$63766 ( \63740 , RIc0d8410_30);
xor \U$63767 ( \63741 , \63739 , \63740 );
buf \U$63768 ( \63742 , \63741 );
buf \U$63769 ( \63743 , \63742 );
not \U$63770 ( \63744 , \63743 );
buf \U$63771 ( \63745 , \16989 );
not \U$63772 ( \63746 , \63745 );
or \U$63773 ( \63747 , \63744 , \63746 );
buf \U$63774 ( \63748 , \12410 );
buf \U$63775 ( \63749 , \63323 );
nand \U$63776 ( \63750 , \63748 , \63749 );
buf \U$63777 ( \63751 , \63750 );
buf \U$63778 ( \63752 , \63751 );
nand \U$63779 ( \63753 , \63747 , \63752 );
buf \U$63780 ( \63754 , \63753 );
buf \U$63781 ( \63755 , \63754 );
and \U$63782 ( \63756 , \63738 , \63755 );
and \U$63783 ( \63757 , \63720 , \63737 );
or \U$63784 ( \63758 , \63756 , \63757 );
buf \U$63785 ( \63759 , \63758 );
buf \U$63786 ( \63760 , \63759 );
xor \U$63787 ( \63761 , \63703 , \63760 );
buf \U$63788 ( \63762 , RIc0d8500_32);
buf \U$63789 ( \63763 , RIc0daa08_111);
xor \U$63790 ( \63764 , \63762 , \63763 );
buf \U$63791 ( \63765 , \63764 );
buf \U$63792 ( \63766 , \63765 );
not \U$63793 ( \63767 , \63766 );
buf \U$63794 ( \63768 , \14346 );
not \U$63795 ( \63769 , \63768 );
or \U$63796 ( \63770 , \63767 , \63769 );
buf \U$63797 ( \63771 , \25649 );
buf \U$63798 ( \63772 , \63413 );
nand \U$63799 ( \63773 , \63771 , \63772 );
buf \U$63800 ( \63774 , \63773 );
buf \U$63801 ( \63775 , \63774 );
nand \U$63802 ( \63776 , \63770 , \63775 );
buf \U$63803 ( \63777 , \63776 );
buf \U$63804 ( \63778 , \63777 );
buf \U$63805 ( \63779 , RIc0dadc8_119);
buf \U$63806 ( \63780 , RIc0d8140_24);
xor \U$63807 ( \63781 , \63779 , \63780 );
buf \U$63808 ( \63782 , \63781 );
buf \U$63809 ( \63783 , \63782 );
not \U$63810 ( \63784 , \63783 );
buf \U$63811 ( \63785 , \25542 );
not \U$63812 ( \63786 , \63785 );
or \U$63813 ( \63787 , \63784 , \63786 );
buf \U$63814 ( \63788 , \13005 );
buf \U$63815 ( \63789 , \63052 );
nand \U$63816 ( \63790 , \63788 , \63789 );
buf \U$63817 ( \63791 , \63790 );
buf \U$63818 ( \63792 , \63791 );
nand \U$63819 ( \63793 , \63787 , \63792 );
buf \U$63820 ( \63794 , \63793 );
buf \U$63821 ( \63795 , \63794 );
xor \U$63822 ( \63796 , \63778 , \63795 );
buf \U$63823 ( \63797 , RIc0d9b08_79);
buf \U$63824 ( \63798 , RIc0d9400_64);
and \U$63825 ( \63799 , \63797 , \63798 );
not \U$63826 ( \63800 , \63797 );
buf \U$63827 ( \63801 , \43843 );
and \U$63828 ( \63802 , \63800 , \63801 );
nor \U$63829 ( \63803 , \63799 , \63802 );
buf \U$63830 ( \63804 , \63803 );
buf \U$63831 ( \63805 , \63804 );
not \U$63832 ( \63806 , \63805 );
buf \U$63833 ( \63807 , \1021 );
not \U$63834 ( \63808 , \63807 );
or \U$63835 ( \63809 , \63806 , \63808 );
buf \U$63836 ( \63810 , \1026 );
buf \U$63837 ( \63811 , \63373 );
nand \U$63838 ( \63812 , \63810 , \63811 );
buf \U$63839 ( \63813 , \63812 );
buf \U$63840 ( \63814 , \63813 );
nand \U$63841 ( \63815 , \63809 , \63814 );
buf \U$63842 ( \63816 , \63815 );
buf \U$63843 ( \63817 , \63816 );
and \U$63844 ( \63818 , \63796 , \63817 );
and \U$63845 ( \63819 , \63778 , \63795 );
or \U$63846 ( \63820 , \63818 , \63819 );
buf \U$63847 ( \63821 , \63820 );
buf \U$63848 ( \63822 , \63821 );
and \U$63849 ( \63823 , \63761 , \63822 );
and \U$63850 ( \63824 , \63703 , \63760 );
or \U$63851 ( \63825 , \63823 , \63824 );
buf \U$63852 ( \63826 , \63825 );
buf \U$63853 ( \63827 , \63826 );
xor \U$63854 ( \63828 , \63640 , \63827 );
xor \U$63855 ( \63829 , \63362 , \63339 );
xor \U$63856 ( \63830 , \63829 , \63317 );
buf \U$63857 ( \63831 , \63830 );
not \U$63858 ( \63832 , \63831 );
xor \U$63859 ( \63833 , \63449 , \63467 );
xor \U$63860 ( \63834 , \63833 , \63486 );
buf \U$63861 ( \63835 , \63834 );
not \U$63862 ( \63836 , \63835 );
or \U$63863 ( \63837 , \63832 , \63836 );
buf \U$63864 ( \63838 , \63834 );
buf \U$63865 ( \63839 , \63830 );
or \U$63866 ( \63840 , \63838 , \63839 );
xor \U$63867 ( \63841 , \63222 , \63262 );
xor \U$63868 ( \63842 , \63841 , \63243 );
buf \U$63869 ( \63843 , \63842 );
nand \U$63870 ( \63844 , \63840 , \63843 );
buf \U$63871 ( \63845 , \63844 );
buf \U$63872 ( \63846 , \63845 );
nand \U$63873 ( \63847 , \63837 , \63846 );
buf \U$63874 ( \63848 , \63847 );
buf \U$63875 ( \63849 , \63848 );
xor \U$63876 ( \63850 , \63828 , \63849 );
buf \U$63877 ( \63851 , \63850 );
buf \U$63878 ( \63852 , \63851 );
or \U$63879 ( \63853 , \63504 , \63852 );
buf \U$63880 ( \63854 , RIc0dacd8_117);
buf \U$63881 ( \63855 , RIc0d81b8_25);
xor \U$63882 ( \63856 , \63854 , \63855 );
buf \U$63883 ( \63857 , \63856 );
buf \U$63884 ( \63858 , \63857 );
not \U$63885 ( \63859 , \63858 );
buf \U$63886 ( \63860 , \22350 );
not \U$63887 ( \63861 , \63860 );
or \U$63888 ( \63862 , \63859 , \63861 );
buf \U$63889 ( \63863 , \12937 );
buf \U$63890 ( \63864 , RIc0d8140_24);
buf \U$63891 ( \63865 , RIc0dacd8_117);
xor \U$63892 ( \63866 , \63864 , \63865 );
buf \U$63893 ( \63867 , \63866 );
buf \U$63894 ( \63868 , \63867 );
nand \U$63895 ( \63869 , \63863 , \63868 );
buf \U$63896 ( \63870 , \63869 );
buf \U$63897 ( \63871 , \63870 );
nand \U$63898 ( \63872 , \63862 , \63871 );
buf \U$63899 ( \63873 , \63872 );
buf \U$63900 ( \63874 , \63873 );
buf \U$63901 ( \63875 , RIc0d7df8_17);
buf \U$63902 ( \63876 , RIc0db098_125);
xor \U$63903 ( \63877 , \63875 , \63876 );
buf \U$63904 ( \63878 , \63877 );
buf \U$63905 ( \63879 , \63878 );
not \U$63906 ( \63880 , \63879 );
buf \U$63907 ( \63881 , \13461 );
not \U$63908 ( \63882 , \63881 );
or \U$63909 ( \63883 , \63880 , \63882 );
buf \U$63910 ( \63884 , RIc0d7d80_16);
buf \U$63911 ( \63885 , RIc0db098_125);
xnor \U$63912 ( \63886 , \63884 , \63885 );
buf \U$63913 ( \63887 , \63886 );
buf \U$63914 ( \63888 , \63887 );
buf \U$63915 ( \63889 , \22744 );
or \U$63916 ( \63890 , \63888 , \63889 );
buf \U$63917 ( \63891 , \63890 );
buf \U$63918 ( \63892 , \63891 );
nand \U$63919 ( \63893 , \63883 , \63892 );
buf \U$63920 ( \63894 , \63893 );
buf \U$63921 ( \63895 , \63894 );
xor \U$63922 ( \63896 , \63874 , \63895 );
buf \U$63923 ( \63897 , RIc0d9bf8_81);
buf \U$63924 ( \63898 , RIc0d9310_62);
xor \U$63925 ( \63899 , \63897 , \63898 );
buf \U$63926 ( \63900 , \63899 );
buf \U$63927 ( \63901 , \63900 );
not \U$63928 ( \63902 , \63901 );
buf \U$63929 ( \63903 , \17141 );
not \U$63930 ( \63904 , \63903 );
or \U$63931 ( \63905 , \63902 , \63904 );
buf \U$63932 ( \63906 , \1078 );
buf \U$63933 ( \63907 , \63030 );
nand \U$63934 ( \63908 , \63906 , \63907 );
buf \U$63935 ( \63909 , \63908 );
buf \U$63936 ( \63910 , \63909 );
nand \U$63937 ( \63911 , \63905 , \63910 );
buf \U$63938 ( \63912 , \63911 );
buf \U$63939 ( \63913 , \63912 );
not \U$63940 ( \63914 , \63913 );
buf \U$63941 ( \63915 , RIc0d9400_64);
buf \U$63942 ( \63916 , RIc0d9b80_80);
or \U$63943 ( \63917 , \63915 , \63916 );
buf \U$63944 ( \63918 , RIc0d9bf8_81);
nand \U$63945 ( \63919 , \63917 , \63918 );
buf \U$63946 ( \63920 , \63919 );
buf \U$63947 ( \63921 , \63920 );
buf \U$63948 ( \63922 , RIc0d9400_64);
buf \U$63949 ( \63923 , RIc0d9b80_80);
nand \U$63950 ( \63924 , \63922 , \63923 );
buf \U$63951 ( \63925 , \63924 );
buf \U$63952 ( \63926 , \63925 );
buf \U$63953 ( \63927 , RIc0d9b08_79);
nand \U$63954 ( \63928 , \63921 , \63926 , \63927 );
buf \U$63955 ( \63929 , \63928 );
buf \U$63956 ( \63930 , \63929 );
nor \U$63957 ( \63931 , \63914 , \63930 );
buf \U$63958 ( \63932 , \63931 );
buf \U$63959 ( \63933 , \63932 );
and \U$63960 ( \63934 , \63896 , \63933 );
and \U$63961 ( \63935 , \63874 , \63895 );
or \U$63962 ( \63936 , \63934 , \63935 );
buf \U$63963 ( \63937 , \63936 );
buf \U$63964 ( \63938 , \63937 );
buf \U$63965 ( \63939 , RIc0da918_109);
buf \U$63966 ( \63940 , RIc0d85f0_34);
xor \U$63967 ( \63941 , \63939 , \63940 );
buf \U$63968 ( \63942 , \63941 );
buf \U$63969 ( \63943 , \63942 );
not \U$63970 ( \63944 , \63943 );
buf \U$63971 ( \63945 , \20759 );
not \U$63972 ( \63946 , \63945 );
or \U$63973 ( \63947 , \63944 , \63946 );
buf \U$63974 ( \63948 , \15909 );
buf \U$63975 ( \63949 , RIc0da918_109);
buf \U$63976 ( \63950 , RIc0d8578_33);
xor \U$63977 ( \63951 , \63949 , \63950 );
buf \U$63978 ( \63952 , \63951 );
buf \U$63979 ( \63953 , \63952 );
nand \U$63980 ( \63954 , \63948 , \63953 );
buf \U$63981 ( \63955 , \63954 );
buf \U$63982 ( \63956 , \63955 );
nand \U$63983 ( \63957 , \63947 , \63956 );
buf \U$63984 ( \63958 , \63957 );
buf \U$63985 ( \63959 , \63958 );
not \U$63986 ( \63960 , \63959 );
buf \U$63987 ( \63961 , RIc0dacd8_117);
buf \U$63988 ( \63962 , RIc0d8230_26);
xor \U$63989 ( \63963 , \63961 , \63962 );
buf \U$63990 ( \63964 , \63963 );
buf \U$63991 ( \63965 , \63964 );
not \U$63992 ( \63966 , \63965 );
buf \U$63993 ( \63967 , \13146 );
not \U$63994 ( \63968 , \63967 );
or \U$63995 ( \63969 , \63966 , \63968 );
buf \U$63996 ( \63970 , \12937 );
buf \U$63997 ( \63971 , \63857 );
nand \U$63998 ( \63972 , \63970 , \63971 );
buf \U$63999 ( \63973 , \63972 );
buf \U$64000 ( \63974 , \63973 );
nand \U$64001 ( \63975 , \63969 , \63974 );
buf \U$64002 ( \63976 , \63975 );
buf \U$64003 ( \63977 , \63976 );
not \U$64004 ( \63978 , \63977 );
or \U$64005 ( \63979 , \63960 , \63978 );
buf \U$64006 ( \63980 , \63976 );
buf \U$64007 ( \63981 , \63958 );
or \U$64008 ( \63982 , \63980 , \63981 );
buf \U$64009 ( \63983 , RIc0d7e70_18);
buf \U$64010 ( \63984 , RIc0db098_125);
xor \U$64011 ( \63985 , \63983 , \63984 );
buf \U$64012 ( \63986 , \63985 );
buf \U$64013 ( \63987 , \63986 );
not \U$64014 ( \63988 , \63987 );
buf \U$64015 ( \63989 , \13461 );
not \U$64016 ( \63990 , \63989 );
or \U$64017 ( \63991 , \63988 , \63990 );
buf \U$64018 ( \63992 , \15793 );
buf \U$64019 ( \63993 , \63878 );
nand \U$64020 ( \63994 , \63992 , \63993 );
buf \U$64021 ( \63995 , \63994 );
buf \U$64022 ( \63996 , \63995 );
nand \U$64023 ( \63997 , \63991 , \63996 );
buf \U$64024 ( \63998 , \63997 );
buf \U$64025 ( \63999 , \63998 );
nand \U$64026 ( \64000 , \63982 , \63999 );
buf \U$64027 ( \64001 , \64000 );
buf \U$64028 ( \64002 , \64001 );
nand \U$64029 ( \64003 , \63979 , \64002 );
buf \U$64030 ( \64004 , \64003 );
buf \U$64031 ( \64005 , \64004 );
not \U$64032 ( \64006 , \64005 );
buf \U$64033 ( \64007 , \64006 );
buf \U$64034 ( \64008 , \64007 );
not \U$64035 ( \64009 , \64008 );
xor \U$64036 ( \64010 , RIc0da558_101, RIc0d89b0_42);
buf \U$64037 ( \64011 , \64010 );
not \U$64038 ( \64012 , \64011 );
buf \U$64039 ( \64013 , \22631 );
not \U$64040 ( \64014 , \64013 );
or \U$64041 ( \64015 , \64012 , \64014 );
buf \U$64042 ( \64016 , \16676 );
buf \U$64043 ( \64017 , \63160 );
nand \U$64044 ( \64018 , \64016 , \64017 );
buf \U$64045 ( \64019 , \64018 );
buf \U$64046 ( \64020 , \64019 );
nand \U$64047 ( \64021 , \64015 , \64020 );
buf \U$64048 ( \64022 , \64021 );
buf \U$64049 ( \64023 , \64022 );
not \U$64050 ( \64024 , \64023 );
xor \U$64051 ( \64025 , RIc0da288_95, RIc0d8c80_48);
buf \U$64052 ( \64026 , \64025 );
not \U$64053 ( \64027 , \64026 );
buf \U$64054 ( \64028 , \330 );
not \U$64055 ( \64029 , \64028 );
or \U$64056 ( \64030 , \64027 , \64029 );
buf \U$64057 ( \64031 , \14707 );
buf \U$64058 ( \64032 , RIc0da288_95);
buf \U$64059 ( \64033 , RIc0d8c08_47);
xor \U$64060 ( \64034 , \64032 , \64033 );
buf \U$64061 ( \64035 , \64034 );
buf \U$64062 ( \64036 , \64035 );
nand \U$64063 ( \64037 , \64031 , \64036 );
buf \U$64064 ( \64038 , \64037 );
buf \U$64065 ( \64039 , \64038 );
nand \U$64066 ( \64040 , \64030 , \64039 );
buf \U$64067 ( \64041 , \64040 );
buf \U$64068 ( \64042 , \64041 );
not \U$64069 ( \64043 , \64042 );
or \U$64070 ( \64044 , \64024 , \64043 );
buf \U$64071 ( \64045 , \64041 );
buf \U$64072 ( \64046 , \64022 );
or \U$64073 ( \64047 , \64045 , \64046 );
buf \U$64074 ( \64048 , RIc0d88c0_40);
buf \U$64075 ( \64049 , RIc0da648_103);
xor \U$64076 ( \64050 , \64048 , \64049 );
buf \U$64077 ( \64051 , \64050 );
buf \U$64078 ( \64052 , \64051 );
not \U$64079 ( \64053 , \64052 );
buf \U$64080 ( \64054 , \13706 );
not \U$64081 ( \64055 , \64054 );
or \U$64082 ( \64056 , \64053 , \64055 );
buf \U$64083 ( \64057 , \18416 );
buf \U$64084 ( \64058 , RIc0d8848_39);
buf \U$64085 ( \64059 , RIc0da648_103);
xor \U$64086 ( \64060 , \64058 , \64059 );
buf \U$64087 ( \64061 , \64060 );
buf \U$64088 ( \64062 , \64061 );
nand \U$64089 ( \64063 , \64057 , \64062 );
buf \U$64090 ( \64064 , \64063 );
buf \U$64091 ( \64065 , \64064 );
nand \U$64092 ( \64066 , \64056 , \64065 );
buf \U$64093 ( \64067 , \64066 );
buf \U$64094 ( \64068 , \64067 );
nand \U$64095 ( \64069 , \64047 , \64068 );
buf \U$64096 ( \64070 , \64069 );
buf \U$64097 ( \64071 , \64070 );
nand \U$64098 ( \64072 , \64044 , \64071 );
buf \U$64099 ( \64073 , \64072 );
buf \U$64100 ( \64074 , \64073 );
not \U$64101 ( \64075 , \64074 );
buf \U$64102 ( \64076 , \64075 );
buf \U$64103 ( \64077 , \64076 );
not \U$64104 ( \64078 , \64077 );
or \U$64105 ( \64079 , \64009 , \64078 );
xor \U$64106 ( \64080 , RIc0d9ce8_83, RIc0d9220_60);
buf \U$64107 ( \64081 , \64080 );
not \U$64108 ( \64082 , \64081 );
buf \U$64109 ( \64083 , \2088 );
not \U$64110 ( \64084 , \64083 );
or \U$64111 ( \64085 , \64082 , \64084 );
buf \U$64112 ( \64086 , \993 );
buf \U$64113 ( \64087 , \63227 );
nand \U$64114 ( \64088 , \64086 , \64087 );
buf \U$64115 ( \64089 , \64088 );
buf \U$64116 ( \64090 , \64089 );
nand \U$64117 ( \64091 , \64085 , \64090 );
buf \U$64118 ( \64092 , \64091 );
buf \U$64119 ( \64093 , \64092 );
xor \U$64120 ( \64094 , RIc0d9dd8_85, RIc0d9130_58);
buf \U$64121 ( \64095 , \64094 );
not \U$64122 ( \64096 , \64095 );
buf \U$64123 ( \64097 , \1389 );
not \U$64124 ( \64098 , \64097 );
or \U$64125 ( \64099 , \64096 , \64098 );
buf \U$64126 ( \64100 , \921 );
buf \U$64127 ( \64101 , \63391 );
nand \U$64128 ( \64102 , \64100 , \64101 );
buf \U$64129 ( \64103 , \64102 );
buf \U$64130 ( \64104 , \64103 );
nand \U$64131 ( \64105 , \64099 , \64104 );
buf \U$64132 ( \64106 , \64105 );
buf \U$64133 ( \64107 , \64106 );
xor \U$64134 ( \64108 , \64093 , \64107 );
xor \U$64135 ( \64109 , RIc0da378_97, RIc0d8b90_46);
buf \U$64136 ( \64110 , \64109 );
not \U$64137 ( \64111 , \64110 );
buf \U$64138 ( \64112 , \26572 );
not \U$64139 ( \64113 , \64112 );
or \U$64140 ( \64114 , \64111 , \64113 );
buf \U$64141 ( \64115 , \734 );
buf \U$64142 ( \64116 , \63206 );
nand \U$64143 ( \64117 , \64115 , \64116 );
buf \U$64144 ( \64118 , \64117 );
buf \U$64145 ( \64119 , \64118 );
nand \U$64146 ( \64120 , \64114 , \64119 );
buf \U$64147 ( \64121 , \64120 );
buf \U$64148 ( \64122 , \64121 );
and \U$64149 ( \64123 , \64108 , \64122 );
and \U$64150 ( \64124 , \64093 , \64107 );
or \U$64151 ( \64125 , \64123 , \64124 );
buf \U$64152 ( \64126 , \64125 );
buf \U$64153 ( \64127 , \64126 );
nand \U$64154 ( \64128 , \64079 , \64127 );
buf \U$64155 ( \64129 , \64128 );
buf \U$64156 ( \64130 , \64129 );
buf \U$64157 ( \64131 , \64073 );
buf \U$64158 ( \64132 , \64004 );
nand \U$64159 ( \64133 , \64131 , \64132 );
buf \U$64160 ( \64134 , \64133 );
buf \U$64161 ( \64135 , \64134 );
nand \U$64162 ( \64136 , \64130 , \64135 );
buf \U$64163 ( \64137 , \64136 );
buf \U$64164 ( \64138 , \64137 );
xor \U$64165 ( \64139 , \63938 , \64138 );
buf \U$64166 ( \64140 , \44382 );
not \U$64167 ( \64141 , \64140 );
buf \U$64168 ( \64142 , \64141 );
buf \U$64169 ( \64143 , \64142 );
not \U$64170 ( \64144 , \64143 );
buf \U$64171 ( \64145 , \63887 );
not \U$64172 ( \64146 , \64145 );
and \U$64173 ( \64147 , \64144 , \64146 );
buf \U$64174 ( \64148 , RIc0db098_125);
buf \U$64175 ( \64149 , RIc0d7d08_15);
xor \U$64176 ( \64150 , \64148 , \64149 );
buf \U$64177 ( \64151 , \64150 );
buf \U$64178 ( \64152 , \64151 );
not \U$64179 ( \64153 , \64152 );
buf \U$64180 ( \64154 , \18699 );
nor \U$64181 ( \64155 , \64153 , \64154 );
buf \U$64182 ( \64156 , \64155 );
buf \U$64183 ( \64157 , \64156 );
nor \U$64184 ( \64158 , \64147 , \64157 );
buf \U$64185 ( \64159 , \64158 );
buf \U$64186 ( \64160 , \64159 );
buf \U$64187 ( \64161 , \63380 );
not \U$64188 ( \64162 , \64161 );
buf \U$64189 ( \64163 , \396 );
not \U$64190 ( \64164 , \64163 );
or \U$64191 ( \64165 , \64162 , \64164 );
buf \U$64192 ( \64166 , \402 );
buf \U$64193 ( \64167 , RIc0d9298_61);
buf \U$64194 ( \64168 , RIc0d9b08_79);
xor \U$64195 ( \64169 , \64167 , \64168 );
buf \U$64196 ( \64170 , \64169 );
buf \U$64197 ( \64171 , \64170 );
nand \U$64198 ( \64172 , \64166 , \64171 );
buf \U$64199 ( \64173 , \64172 );
buf \U$64200 ( \64174 , \64173 );
nand \U$64201 ( \64175 , \64165 , \64174 );
buf \U$64202 ( \64176 , \64175 );
buf \U$64203 ( \64177 , \64176 );
not \U$64204 ( \64178 , \64177 );
buf \U$64205 ( \64179 , RIc0d9400_64);
buf \U$64206 ( \64180 , RIc0d9a90_78);
or \U$64207 ( \64181 , \64179 , \64180 );
buf \U$64208 ( \64182 , RIc0d9b08_79);
nand \U$64209 ( \64183 , \64181 , \64182 );
buf \U$64210 ( \64184 , \64183 );
buf \U$64211 ( \64185 , \64184 );
buf \U$64212 ( \64186 , RIc0d9400_64);
buf \U$64213 ( \64187 , RIc0d9a90_78);
nand \U$64214 ( \64188 , \64186 , \64187 );
buf \U$64215 ( \64189 , \64188 );
buf \U$64216 ( \64190 , \64189 );
buf \U$64217 ( \64191 , RIc0d9a18_77);
and \U$64218 ( \64192 , \64185 , \64190 , \64191 );
buf \U$64219 ( \64193 , \64192 );
buf \U$64220 ( \64194 , \64193 );
not \U$64221 ( \64195 , \64194 );
buf \U$64222 ( \64196 , \64195 );
buf \U$64223 ( \64197 , \64196 );
not \U$64224 ( \64198 , \64197 );
and \U$64225 ( \64199 , \64178 , \64198 );
buf \U$64226 ( \64200 , \64176 );
buf \U$64227 ( \64201 , \64196 );
and \U$64228 ( \64202 , \64200 , \64201 );
nor \U$64229 ( \64203 , \64199 , \64202 );
buf \U$64230 ( \64204 , \64203 );
buf \U$64231 ( \64205 , \64204 );
not \U$64232 ( \64206 , \64205 );
buf \U$64233 ( \64207 , \64206 );
buf \U$64234 ( \64208 , \64207 );
xor \U$64235 ( \64209 , \64160 , \64208 );
buf \U$64236 ( \64210 , \64035 );
not \U$64237 ( \64211 , \64210 );
buf \U$64238 ( \64212 , \3714 );
not \U$64239 ( \64213 , \64212 );
or \U$64240 ( \64214 , \64211 , \64213 );
buf \U$64241 ( \64215 , \343 );
buf \U$64242 ( \64216 , RIc0da288_95);
buf \U$64243 ( \64217 , RIc0d8b90_46);
xor \U$64244 ( \64218 , \64216 , \64217 );
buf \U$64245 ( \64219 , \64218 );
buf \U$64246 ( \64220 , \64219 );
nand \U$64247 ( \64221 , \64215 , \64220 );
buf \U$64248 ( \64222 , \64221 );
buf \U$64249 ( \64223 , \64222 );
nand \U$64250 ( \64224 , \64214 , \64223 );
buf \U$64251 ( \64225 , \64224 );
buf \U$64252 ( \64226 , \64225 );
buf \U$64253 ( \64227 , \63952 );
not \U$64254 ( \64228 , \64227 );
buf \U$64255 ( \64229 , \21959 );
not \U$64256 ( \64230 , \64229 );
or \U$64257 ( \64231 , \64228 , \64230 );
buf \U$64258 ( \64232 , \20211 );
buf \U$64259 ( \64233 , RIc0da918_109);
buf \U$64260 ( \64234 , RIc0d8500_32);
xor \U$64261 ( \64235 , \64233 , \64234 );
buf \U$64262 ( \64236 , \64235 );
buf \U$64263 ( \64237 , \64236 );
nand \U$64264 ( \64238 , \64232 , \64237 );
buf \U$64265 ( \64239 , \64238 );
buf \U$64266 ( \64240 , \64239 );
nand \U$64267 ( \64241 , \64231 , \64240 );
buf \U$64268 ( \64242 , \64241 );
buf \U$64269 ( \64243 , \64242 );
or \U$64270 ( \64244 , \64226 , \64243 );
buf \U$64271 ( \64245 , \64061 );
not \U$64272 ( \64246 , \64245 );
buf \U$64273 ( \64247 , \13042 );
not \U$64274 ( \64248 , \64247 );
or \U$64275 ( \64249 , \64246 , \64248 );
buf \U$64276 ( \64250 , \16584 );
buf \U$64277 ( \64251 , RIc0d87d0_38);
buf \U$64278 ( \64252 , RIc0da648_103);
xor \U$64279 ( \64253 , \64251 , \64252 );
buf \U$64280 ( \64254 , \64253 );
buf \U$64281 ( \64255 , \64254 );
nand \U$64282 ( \64256 , \64250 , \64255 );
buf \U$64283 ( \64257 , \64256 );
buf \U$64284 ( \64258 , \64257 );
nand \U$64285 ( \64259 , \64249 , \64258 );
buf \U$64286 ( \64260 , \64259 );
buf \U$64287 ( \64261 , \64260 );
nand \U$64288 ( \64262 , \64244 , \64261 );
buf \U$64289 ( \64263 , \64262 );
buf \U$64290 ( \64264 , \64263 );
buf \U$64291 ( \64265 , \64225 );
buf \U$64292 ( \64266 , \64242 );
nand \U$64293 ( \64267 , \64265 , \64266 );
buf \U$64294 ( \64268 , \64267 );
buf \U$64295 ( \64269 , \64268 );
nand \U$64296 ( \64270 , \64264 , \64269 );
buf \U$64297 ( \64271 , \64270 );
buf \U$64298 ( \64272 , \64271 );
xnor \U$64299 ( \64273 , \64209 , \64272 );
buf \U$64300 ( \64274 , \64273 );
buf \U$64301 ( \64275 , \64274 );
xor \U$64302 ( \64276 , \64139 , \64275 );
buf \U$64303 ( \64277 , \64276 );
buf \U$64304 ( \64278 , \64277 );
nand \U$64305 ( \64279 , \63853 , \64278 );
buf \U$64306 ( \64280 , \64279 );
buf \U$64307 ( \64281 , \64280 );
buf \U$64308 ( \64282 , \63503 );
buf \U$64309 ( \64283 , \63851 );
nand \U$64310 ( \64284 , \64282 , \64283 );
buf \U$64311 ( \64285 , \64284 );
buf \U$64312 ( \64286 , \64285 );
nand \U$64313 ( \64287 , \64281 , \64286 );
buf \U$64314 ( \64288 , \64287 );
buf \U$64315 ( \64289 , \64288 );
xor \U$64316 ( \64290 , \63938 , \64138 );
and \U$64317 ( \64291 , \64290 , \64275 );
and \U$64318 ( \64292 , \63938 , \64138 );
or \U$64319 ( \64293 , \64291 , \64292 );
buf \U$64320 ( \64294 , \64293 );
buf \U$64321 ( \64295 , \64294 );
xor \U$64322 ( \64296 , \63202 , \63299 );
and \U$64323 ( \64297 , \64296 , \63501 );
and \U$64324 ( \64298 , \63202 , \63299 );
or \U$64325 ( \64299 , \64297 , \64298 );
buf \U$64326 ( \64300 , \64299 );
buf \U$64327 ( \64301 , \64300 );
xor \U$64328 ( \64302 , \64295 , \64301 );
buf \U$64329 ( \64303 , \64204 );
buf \U$64330 ( \64304 , \64159 );
nand \U$64331 ( \64305 , \64303 , \64304 );
buf \U$64332 ( \64306 , \64305 );
not \U$64333 ( \64307 , \64306 );
not \U$64334 ( \64308 , \64271 );
or \U$64335 ( \64309 , \64307 , \64308 );
buf \U$64336 ( \64310 , \64159 );
not \U$64337 ( \64311 , \64310 );
buf \U$64338 ( \64312 , \64207 );
nand \U$64339 ( \64313 , \64311 , \64312 );
buf \U$64340 ( \64314 , \64313 );
nand \U$64341 ( \64315 , \64309 , \64314 );
buf \U$64342 ( \64316 , \64315 );
buf \U$64343 ( \64317 , \63430 );
buf \U$64344 ( \64318 , \63497 );
or \U$64345 ( \64319 , \64317 , \64318 );
buf \U$64346 ( \64320 , \63368 );
nand \U$64347 ( \64321 , \64319 , \64320 );
buf \U$64348 ( \64322 , \64321 );
buf \U$64349 ( \64323 , \64322 );
buf \U$64350 ( \64324 , \63497 );
buf \U$64351 ( \64325 , \63430 );
nand \U$64352 ( \64326 , \64324 , \64325 );
buf \U$64353 ( \64327 , \64326 );
buf \U$64354 ( \64328 , \64327 );
nand \U$64355 ( \64329 , \64323 , \64328 );
buf \U$64356 ( \64330 , \64329 );
buf \U$64357 ( \64331 , \64330 );
xor \U$64358 ( \64332 , \64316 , \64331 );
xor \U$64359 ( \64333 , \63274 , \63280 );
and \U$64360 ( \64334 , \64333 , \63296 );
and \U$64361 ( \64335 , \63274 , \63280 );
or \U$64362 ( \64336 , \64334 , \64335 );
buf \U$64363 ( \64337 , \64336 );
buf \U$64364 ( \64338 , \64337 );
xor \U$64365 ( \64339 , \64332 , \64338 );
buf \U$64366 ( \64340 , \64339 );
buf \U$64367 ( \64341 , \64340 );
xor \U$64368 ( \64342 , \64302 , \64341 );
buf \U$64369 ( \64343 , \64342 );
buf \U$64370 ( \64344 , \64343 );
xor \U$64371 ( \64345 , \64289 , \64344 );
xor \U$64372 ( \64346 , \63640 , \63827 );
and \U$64373 ( \64347 , \64346 , \63849 );
and \U$64374 ( \64348 , \63640 , \63827 );
or \U$64375 ( \64349 , \64347 , \64348 );
buf \U$64376 ( \64350 , \64349 );
buf \U$64377 ( \64351 , \64350 );
xor \U$64378 ( \64352 , \63090 , \63111 );
and \U$64379 ( \64353 , \64352 , \63130 );
and \U$64380 ( \64354 , \63090 , \63111 );
or \U$64381 ( \64355 , \64353 , \64354 );
buf \U$64382 ( \64356 , \64355 );
buf \U$64383 ( \64357 , \64356 );
buf \U$64384 ( \64358 , \63167 );
not \U$64385 ( \64359 , \64358 );
buf \U$64386 ( \64360 , \4042 );
not \U$64387 ( \64361 , \64360 );
or \U$64388 ( \64362 , \64359 , \64361 );
buf \U$64389 ( \64363 , \12839 );
xor \U$64390 ( \64364 , RIc0da558_101, RIc0d8848_39);
buf \U$64391 ( \64365 , \64364 );
nand \U$64392 ( \64366 , \64363 , \64365 );
buf \U$64393 ( \64367 , \64366 );
buf \U$64394 ( \64368 , \64367 );
nand \U$64395 ( \64369 , \64362 , \64368 );
buf \U$64396 ( \64370 , \64369 );
buf \U$64397 ( \64371 , \64370 );
buf \U$64398 ( \64372 , \63150 );
not \U$64399 ( \64373 , \64372 );
buf \U$64400 ( \64374 , \14186 );
not \U$64401 ( \64375 , \64374 );
or \U$64402 ( \64376 , \64373 , \64375 );
buf \U$64403 ( \64377 , \12303 );
buf \U$64404 ( \64378 , RIc0d81b8_25);
buf \U$64405 ( \64379 , RIc0dabe8_115);
xor \U$64406 ( \64380 , \64378 , \64379 );
buf \U$64407 ( \64381 , \64380 );
buf \U$64408 ( \64382 , \64381 );
nand \U$64409 ( \64383 , \64377 , \64382 );
buf \U$64410 ( \64384 , \64383 );
buf \U$64411 ( \64385 , \64384 );
nand \U$64412 ( \64386 , \64376 , \64385 );
buf \U$64413 ( \64387 , \64386 );
buf \U$64414 ( \64388 , \64387 );
xor \U$64415 ( \64389 , \64371 , \64388 );
buf \U$64416 ( \64390 , \63443 );
not \U$64417 ( \64391 , \64390 );
buf \U$64418 ( \64392 , \17595 );
not \U$64419 ( \64393 , \64392 );
or \U$64420 ( \64394 , \64391 , \64393 );
buf \U$64421 ( \64395 , \12342 );
xor \U$64422 ( \64396 , RIc0da828_107, RIc0d8578_33);
buf \U$64423 ( \64397 , \64396 );
nand \U$64424 ( \64398 , \64395 , \64397 );
buf \U$64425 ( \64399 , \64398 );
buf \U$64426 ( \64400 , \64399 );
nand \U$64427 ( \64401 , \64394 , \64400 );
buf \U$64428 ( \64402 , \64401 );
buf \U$64429 ( \64403 , \64402 );
xor \U$64430 ( \64404 , \64389 , \64403 );
buf \U$64431 ( \64405 , \64404 );
buf \U$64432 ( \64406 , \64405 );
xor \U$64433 ( \64407 , \64357 , \64406 );
buf \U$64434 ( \64408 , \63867 );
not \U$64435 ( \64409 , \64408 );
buf \U$64436 ( \64410 , \22350 );
not \U$64437 ( \64411 , \64410 );
or \U$64438 ( \64412 , \64409 , \64411 );
buf \U$64439 ( \64413 , \12937 );
buf \U$64440 ( \64414 , RIc0dacd8_117);
buf \U$64441 ( \64415 , RIc0d80c8_23);
xor \U$64442 ( \64416 , \64414 , \64415 );
buf \U$64443 ( \64417 , \64416 );
buf \U$64444 ( \64418 , \64417 );
nand \U$64445 ( \64419 , \64413 , \64418 );
buf \U$64446 ( \64420 , \64419 );
buf \U$64447 ( \64421 , \64420 );
nand \U$64448 ( \64422 , \64412 , \64421 );
buf \U$64449 ( \64423 , \64422 );
buf \U$64450 ( \64424 , \64236 );
not \U$64451 ( \64425 , \64424 );
buf \U$64452 ( \64426 , \14210 );
not \U$64453 ( \64427 , \64426 );
or \U$64454 ( \64428 , \64425 , \64427 );
buf \U$64455 ( \64429 , \20211 );
buf \U$64456 ( \64430 , RIc0d8488_31);
buf \U$64457 ( \64431 , RIc0da918_109);
xor \U$64458 ( \64432 , \64430 , \64431 );
buf \U$64459 ( \64433 , \64432 );
buf \U$64460 ( \64434 , \64433 );
nand \U$64461 ( \64435 , \64429 , \64434 );
buf \U$64462 ( \64436 , \64435 );
buf \U$64463 ( \64437 , \64436 );
nand \U$64464 ( \64438 , \64428 , \64437 );
buf \U$64465 ( \64439 , \64438 );
xor \U$64466 ( \64440 , \64423 , \64439 );
buf \U$64467 ( \64441 , \43843 );
buf \U$64468 ( \64442 , RIc0d9a18_77);
or \U$64469 ( \64443 , \64441 , \64442 );
buf \U$64470 ( \64444 , \1113 );
buf \U$64471 ( \64445 , RIc0d9400_64);
or \U$64472 ( \64446 , \64444 , \64445 );
nand \U$64473 ( \64447 , \64443 , \64446 );
buf \U$64474 ( \64448 , \64447 );
buf \U$64475 ( \64449 , \64448 );
not \U$64476 ( \64450 , \64449 );
buf \U$64477 ( \64451 , \1183 );
not \U$64478 ( \64452 , \64451 );
or \U$64479 ( \64453 , \64450 , \64452 );
buf \U$64480 ( \64454 , \14374 );
buf \U$64481 ( \64455 , RIc0d9a18_77);
buf \U$64482 ( \64456 , RIc0d9388_63);
xor \U$64483 ( \64457 , \64455 , \64456 );
buf \U$64484 ( \64458 , \64457 );
buf \U$64485 ( \64459 , \64458 );
nand \U$64486 ( \64460 , \64454 , \64459 );
buf \U$64487 ( \64461 , \64460 );
buf \U$64488 ( \64462 , \64461 );
nand \U$64489 ( \64463 , \64453 , \64462 );
buf \U$64490 ( \64464 , \64463 );
xor \U$64491 ( \64465 , \64440 , \64464 );
buf \U$64492 ( \64466 , \64465 );
xnor \U$64493 ( \64467 , \64407 , \64466 );
buf \U$64494 ( \64468 , \64467 );
buf \U$64495 ( \64469 , \64468 );
not \U$64496 ( \64470 , \64469 );
buf \U$64497 ( \64471 , \63082 );
not \U$64498 ( \64472 , \64471 );
buf \U$64499 ( \64473 , \15609 );
not \U$64500 ( \64474 , \64473 );
or \U$64501 ( \64475 , \64472 , \64474 );
buf \U$64502 ( \64476 , RIc0d7c18_13);
buf \U$64503 ( \64477 , RIc0db188_127);
xor \U$64504 ( \64478 , \64476 , \64477 );
buf \U$64505 ( \64479 , \64478 );
buf \U$64506 ( \64480 , \64479 );
buf \U$64507 ( \64481 , RIc0db200_128);
nand \U$64508 ( \64482 , \64480 , \64481 );
buf \U$64509 ( \64483 , \64482 );
buf \U$64510 ( \64484 , \64483 );
nand \U$64511 ( \64485 , \64475 , \64484 );
buf \U$64512 ( \64486 , \64485 );
buf \U$64513 ( \64487 , \64486 );
buf \U$64514 ( \64488 , \63356 );
not \U$64515 ( \64489 , \64488 );
buf \U$64516 ( \64490 , \25371 );
not \U$64517 ( \64491 , \64490 );
or \U$64518 ( \64492 , \64489 , \64491 );
buf \U$64519 ( \64493 , \2476 );
xor \U$64520 ( \64494 , RIc0da468_99, RIc0d8938_41);
buf \U$64521 ( \64495 , \64494 );
nand \U$64522 ( \64496 , \64493 , \64495 );
buf \U$64523 ( \64497 , \64496 );
buf \U$64524 ( \64498 , \64497 );
nand \U$64525 ( \64499 , \64492 , \64498 );
buf \U$64526 ( \64500 , \64499 );
buf \U$64527 ( \64501 , \64500 );
xor \U$64528 ( \64502 , \64487 , \64501 );
buf \U$64529 ( \64503 , \63461 );
not \U$64530 ( \64504 , \64503 );
buf \U$64531 ( \64505 , \64504 );
buf \U$64532 ( \64506 , \64505 );
buf \U$64533 ( \64507 , \473 );
or \U$64534 ( \64508 , \64506 , \64507 );
buf \U$64535 ( \64509 , \40339 );
buf \U$64536 ( \64510 , RIc0d8c08_47);
buf \U$64537 ( \64511 , RIc0da198_93);
xor \U$64538 ( \64512 , \64510 , \64511 );
buf \U$64539 ( \64513 , \64512 );
buf \U$64540 ( \64514 , \64513 );
not \U$64541 ( \64515 , \64514 );
buf \U$64542 ( \64516 , \64515 );
buf \U$64543 ( \64517 , \64516 );
or \U$64544 ( \64518 , \64509 , \64517 );
nand \U$64545 ( \64519 , \64508 , \64518 );
buf \U$64546 ( \64520 , \64519 );
buf \U$64547 ( \64521 , \64520 );
xor \U$64548 ( \64522 , \64502 , \64521 );
buf \U$64549 ( \64523 , \64522 );
buf \U$64550 ( \64524 , \64219 );
not \U$64551 ( \64525 , \64524 );
buf \U$64552 ( \64526 , \330 );
not \U$64553 ( \64527 , \64526 );
or \U$64554 ( \64528 , \64525 , \64527 );
buf \U$64555 ( \64529 , \14707 );
buf \U$64556 ( \64530 , RIc0d8b18_45);
buf \U$64557 ( \64531 , RIc0da288_95);
xor \U$64558 ( \64532 , \64530 , \64531 );
buf \U$64559 ( \64533 , \64532 );
buf \U$64560 ( \64534 , \64533 );
nand \U$64561 ( \64535 , \64529 , \64534 );
buf \U$64562 ( \64536 , \64535 );
buf \U$64563 ( \64537 , \64536 );
nand \U$64564 ( \64538 , \64528 , \64537 );
buf \U$64565 ( \64539 , \64538 );
buf \U$64566 ( \64540 , \64539 );
not \U$64567 ( \64541 , \64540 );
buf \U$64568 ( \64542 , \63237 );
not \U$64569 ( \64543 , \64542 );
buf \U$64570 ( \64544 , \2088 );
not \U$64571 ( \64545 , \64544 );
or \U$64572 ( \64546 , \64543 , \64545 );
buf \U$64573 ( \64547 , \993 );
buf \U$64574 ( \64548 , RIc0d9ce8_83);
buf \U$64575 ( \64549 , RIc0d90b8_57);
xor \U$64576 ( \64550 , \64548 , \64549 );
buf \U$64577 ( \64551 , \64550 );
buf \U$64578 ( \64552 , \64551 );
nand \U$64579 ( \64553 , \64547 , \64552 );
buf \U$64580 ( \64554 , \64553 );
buf \U$64581 ( \64555 , \64554 );
nand \U$64582 ( \64556 , \64546 , \64555 );
buf \U$64583 ( \64557 , \64556 );
buf \U$64584 ( \64558 , \64557 );
not \U$64585 ( \64559 , \64558 );
buf \U$64586 ( \64560 , \64559 );
buf \U$64587 ( \64561 , \64560 );
not \U$64588 ( \64562 , \64561 );
or \U$64589 ( \64563 , \64541 , \64562 );
buf \U$64590 ( \64564 , \64539 );
buf \U$64591 ( \64565 , \64560 );
or \U$64592 ( \64566 , \64564 , \64565 );
nand \U$64593 ( \64567 , \64563 , \64566 );
buf \U$64594 ( \64568 , \64567 );
buf \U$64595 ( \64569 , \64568 );
buf \U$64596 ( \64570 , \63040 );
not \U$64597 ( \64571 , \64570 );
buf \U$64598 ( \64572 , \1063 );
not \U$64599 ( \64573 , \64572 );
or \U$64600 ( \64574 , \64571 , \64573 );
buf \U$64601 ( \64575 , \1078 );
xor \U$64602 ( \64576 , RIc0d9bf8_81, RIc0d91a8_59);
buf \U$64603 ( \64577 , \64576 );
nand \U$64604 ( \64578 , \64575 , \64577 );
buf \U$64605 ( \64579 , \64578 );
buf \U$64606 ( \64580 , \64579 );
nand \U$64607 ( \64581 , \64574 , \64580 );
buf \U$64608 ( \64582 , \64581 );
buf \U$64609 ( \64583 , \64582 );
not \U$64610 ( \64584 , \64583 );
buf \U$64611 ( \64585 , \64584 );
buf \U$64612 ( \64586 , \64585 );
and \U$64613 ( \64587 , \64569 , \64586 );
not \U$64614 ( \64588 , \64569 );
buf \U$64615 ( \64589 , \64582 );
and \U$64616 ( \64590 , \64588 , \64589 );
nor \U$64617 ( \64591 , \64587 , \64590 );
buf \U$64618 ( \64592 , \64591 );
and \U$64619 ( \64593 , \64523 , \64592 );
not \U$64620 ( \64594 , \64523 );
buf \U$64621 ( \64595 , \64592 );
not \U$64622 ( \64596 , \64595 );
buf \U$64623 ( \64597 , \64596 );
and \U$64624 ( \64598 , \64594 , \64597 );
or \U$64625 ( \64599 , \64593 , \64598 );
buf \U$64626 ( \64600 , \64599 );
buf \U$64627 ( \64601 , \63333 );
not \U$64628 ( \64602 , \64601 );
buf \U$64629 ( \64603 , \28776 );
not \U$64630 ( \64604 , \64603 );
or \U$64631 ( \64605 , \64602 , \64604 );
buf \U$64632 ( \64606 , \14405 );
buf \U$64633 ( \64607 , RIc0d82a8_27);
buf \U$64634 ( \64608 , RIc0daaf8_113);
xor \U$64635 ( \64609 , \64607 , \64608 );
buf \U$64636 ( \64610 , \64609 );
buf \U$64637 ( \64611 , \64610 );
nand \U$64638 ( \64612 , \64606 , \64611 );
buf \U$64639 ( \64613 , \64612 );
buf \U$64640 ( \64614 , \64613 );
nand \U$64641 ( \64615 , \64605 , \64614 );
buf \U$64642 ( \64616 , \64615 );
buf \U$64643 ( \64617 , \64616 );
not \U$64644 ( \64618 , \64617 );
buf \U$64645 ( \64619 , \64618 );
buf \U$64646 ( \64620 , \64619 );
buf \U$64647 ( \64621 , \63104 );
not \U$64648 ( \64622 , \64621 );
buf \U$64649 ( \64623 , \3384 );
not \U$64650 ( \64624 , \64623 );
or \U$64651 ( \64625 , \64622 , \64624 );
buf \U$64652 ( \64626 , \13494 );
not \U$64653 ( \64627 , \64626 );
buf \U$64654 ( \64628 , RIc0d8de8_51);
buf \U$64655 ( \64629 , RIc0d9fb8_89);
xor \U$64656 ( \64630 , \64628 , \64629 );
buf \U$64657 ( \64631 , \64630 );
buf \U$64658 ( \64632 , \64631 );
nand \U$64659 ( \64633 , \64627 , \64632 );
buf \U$64660 ( \64634 , \64633 );
buf \U$64661 ( \64635 , \64634 );
nand \U$64662 ( \64636 , \64625 , \64635 );
buf \U$64663 ( \64637 , \64636 );
buf \U$64664 ( \64638 , \64637 );
not \U$64665 ( \64639 , \64638 );
buf \U$64666 ( \64640 , \64639 );
buf \U$64667 ( \64641 , \64640 );
and \U$64668 ( \64642 , \64620 , \64641 );
not \U$64669 ( \64643 , \64620 );
buf \U$64670 ( \64644 , \64637 );
and \U$64671 ( \64645 , \64643 , \64644 );
nor \U$64672 ( \64646 , \64642 , \64645 );
buf \U$64673 ( \64647 , \64646 );
buf \U$64674 ( \64648 , \64647 );
buf \U$64675 ( \64649 , \63398 );
not \U$64676 ( \64650 , \64649 );
buf \U$64677 ( \64651 , \5305 );
not \U$64678 ( \64652 , \64651 );
or \U$64679 ( \64653 , \64650 , \64652 );
buf \U$64680 ( \64654 , \921 );
xor \U$64681 ( \64655 , RIc0d9dd8_85, RIc0d8fc8_55);
buf \U$64682 ( \64656 , \64655 );
nand \U$64683 ( \64657 , \64654 , \64656 );
buf \U$64684 ( \64658 , \64657 );
buf \U$64685 ( \64659 , \64658 );
nand \U$64686 ( \64660 , \64653 , \64659 );
buf \U$64687 ( \64661 , \64660 );
buf \U$64688 ( \64662 , \64661 );
xor \U$64689 ( \64663 , \64648 , \64662 );
buf \U$64690 ( \64664 , \64663 );
buf \U$64691 ( \64665 , \64664 );
xnor \U$64692 ( \64666 , \64600 , \64665 );
buf \U$64693 ( \64667 , \64666 );
buf \U$64694 ( \64668 , \64667 );
not \U$64695 ( \64669 , \64668 );
or \U$64696 ( \64670 , \64470 , \64669 );
buf \U$64697 ( \64671 , \63059 );
not \U$64698 ( \64672 , \64671 );
buf \U$64699 ( \64673 , \13949 );
not \U$64700 ( \64674 , \64673 );
or \U$64701 ( \64675 , \64672 , \64674 );
buf \U$64702 ( \64676 , \13005 );
buf \U$64703 ( \64677 , RIc0d7fd8_21);
buf \U$64704 ( \64678 , RIc0dadc8_119);
xor \U$64705 ( \64679 , \64677 , \64678 );
buf \U$64706 ( \64680 , \64679 );
buf \U$64707 ( \64681 , \64680 );
nand \U$64708 ( \64682 , \64676 , \64681 );
buf \U$64709 ( \64683 , \64682 );
buf \U$64710 ( \64684 , \64683 );
nand \U$64711 ( \64685 , \64675 , \64684 );
buf \U$64712 ( \64686 , \64685 );
buf \U$64713 ( \64687 , \64686 );
not \U$64714 ( \64688 , \64687 );
buf \U$64715 ( \64689 , \63311 );
not \U$64716 ( \64690 , \64689 );
buf \U$64717 ( \64691 , \12736 );
not \U$64718 ( \64692 , \64691 );
or \U$64719 ( \64693 , \64690 , \64692 );
buf \U$64720 ( \64694 , \12744 );
buf \U$64721 ( \64695 , RIc0da738_105);
buf \U$64722 ( \64696 , RIc0d8668_35);
xor \U$64723 ( \64697 , \64695 , \64696 );
buf \U$64724 ( \64698 , \64697 );
buf \U$64725 ( \64699 , \64698 );
nand \U$64726 ( \64700 , \64694 , \64699 );
buf \U$64727 ( \64701 , \64700 );
buf \U$64728 ( \64702 , \64701 );
nand \U$64729 ( \64703 , \64693 , \64702 );
buf \U$64730 ( \64704 , \64703 );
buf \U$64731 ( \64705 , \64704 );
not \U$64732 ( \64706 , \64705 );
buf \U$64733 ( \64707 , \64706 );
buf \U$64734 ( \64708 , \64707 );
not \U$64735 ( \64709 , \64708 );
or \U$64736 ( \64710 , \64688 , \64709 );
buf \U$64737 ( \64711 , \64704 );
buf \U$64738 ( \64712 , \64686 );
not \U$64739 ( \64713 , \64712 );
buf \U$64740 ( \64714 , \64713 );
buf \U$64741 ( \64715 , \64714 );
nand \U$64742 ( \64716 , \64711 , \64715 );
buf \U$64743 ( \64717 , \64716 );
buf \U$64744 ( \64718 , \64717 );
nand \U$64745 ( \64719 , \64710 , \64718 );
buf \U$64746 ( \64720 , \64719 );
buf \U$64747 ( \64721 , \64720 );
buf \U$64748 ( \64722 , \63123 );
not \U$64749 ( \64723 , \64722 );
buf \U$64750 ( \64724 , \704 );
not \U$64751 ( \64725 , \64724 );
or \U$64752 ( \64726 , \64723 , \64725 );
buf \U$64753 ( \64727 , \13293 );
xor \U$64754 ( \64728 , RIc0da0a8_91, RIc0d8cf8_49);
buf \U$64755 ( \64729 , \64728 );
nand \U$64756 ( \64730 , \64727 , \64729 );
buf \U$64757 ( \64731 , \64730 );
buf \U$64758 ( \64732 , \64731 );
nand \U$64759 ( \64733 , \64726 , \64732 );
buf \U$64760 ( \64734 , \64733 );
buf \U$64761 ( \64735 , \64734 );
xor \U$64762 ( \64736 , \64721 , \64735 );
buf \U$64763 ( \64737 , \64736 );
buf \U$64764 ( \64738 , \64737 );
buf \U$64765 ( \64739 , \63480 );
not \U$64766 ( \64740 , \64739 );
buf \U$64767 ( \64741 , \14982 );
not \U$64768 ( \64742 , \64741 );
or \U$64769 ( \64743 , \64740 , \64742 );
buf \U$64770 ( \64744 , \16692 );
buf \U$64771 ( \64745 , RIc0dafa8_123);
buf \U$64772 ( \64746 , RIc0d7df8_17);
xor \U$64773 ( \64747 , \64745 , \64746 );
buf \U$64774 ( \64748 , \64747 );
buf \U$64775 ( \64749 , \64748 );
nand \U$64776 ( \64750 , \64744 , \64749 );
buf \U$64777 ( \64751 , \64750 );
buf \U$64778 ( \64752 , \64751 );
nand \U$64779 ( \64753 , \64743 , \64752 );
buf \U$64780 ( \64754 , \64753 );
buf \U$64781 ( \64755 , \64754 );
buf \U$64782 ( \64756 , \64254 );
not \U$64783 ( \64757 , \64756 );
buf \U$64784 ( \64758 , \16578 );
not \U$64785 ( \64759 , \64758 );
or \U$64786 ( \64760 , \64757 , \64759 );
buf \U$64787 ( \64761 , \13048 );
buf \U$64788 ( \64762 , RIc0da648_103);
buf \U$64789 ( \64763 , RIc0d8758_37);
xor \U$64790 ( \64764 , \64762 , \64763 );
buf \U$64791 ( \64765 , \64764 );
buf \U$64792 ( \64766 , \64765 );
nand \U$64793 ( \64767 , \64761 , \64766 );
buf \U$64794 ( \64768 , \64767 );
buf \U$64795 ( \64769 , \64768 );
nand \U$64796 ( \64770 , \64760 , \64769 );
buf \U$64797 ( \64771 , \64770 );
buf \U$64798 ( \64772 , \64771 );
xor \U$64799 ( \64773 , \64755 , \64772 );
buf \U$64800 ( \64774 , \63185 );
not \U$64801 ( \64775 , \64774 );
buf \U$64802 ( \64776 , \4527 );
not \U$64803 ( \64777 , \64776 );
or \U$64804 ( \64778 , \64775 , \64777 );
buf \U$64805 ( \64779 , \3631 );
xor \U$64806 ( \64780 , RIc0d9ec8_87, RIc0d8ed8_53);
buf \U$64807 ( \64781 , \64780 );
nand \U$64808 ( \64782 , \64779 , \64781 );
buf \U$64809 ( \64783 , \64782 );
buf \U$64810 ( \64784 , \64783 );
nand \U$64811 ( \64785 , \64778 , \64784 );
buf \U$64812 ( \64786 , \64785 );
buf \U$64813 ( \64787 , \64786 );
xor \U$64814 ( \64788 , \64773 , \64787 );
buf \U$64815 ( \64789 , \64788 );
buf \U$64816 ( \64790 , \64789 );
xor \U$64817 ( \64791 , \64738 , \64790 );
buf \U$64818 ( \64792 , \63216 );
not \U$64819 ( \64793 , \64792 );
buf \U$64820 ( \64794 , \16358 );
not \U$64821 ( \64795 , \64794 );
or \U$64822 ( \64796 , \64793 , \64795 );
buf \U$64823 ( \64797 , \734 );
buf \U$64824 ( \64798 , RIc0d8a28_43);
buf \U$64825 ( \64799 , RIc0da378_97);
xor \U$64826 ( \64800 , \64798 , \64799 );
buf \U$64827 ( \64801 , \64800 );
buf \U$64828 ( \64802 , \64801 );
nand \U$64829 ( \64803 , \64797 , \64802 );
buf \U$64830 ( \64804 , \64803 );
buf \U$64831 ( \64805 , \64804 );
nand \U$64832 ( \64806 , \64796 , \64805 );
buf \U$64833 ( \64807 , \64806 );
buf \U$64834 ( \64808 , \64807 );
not \U$64835 ( \64809 , \64808 );
buf \U$64836 ( \64810 , \64809 );
buf \U$64837 ( \64811 , \64810 );
buf \U$64838 ( \64812 , \63256 );
not \U$64839 ( \64813 , \64812 );
buf \U$64840 ( \64814 , \16382 );
not \U$64841 ( \64815 , \64814 );
or \U$64842 ( \64816 , \64813 , \64815 );
buf \U$64843 ( \64817 , \12975 );
xor \U$64844 ( \64818 , RIc0daeb8_121, RIc0d7ee8_19);
buf \U$64845 ( \64819 , \64818 );
nand \U$64846 ( \64820 , \64817 , \64819 );
buf \U$64847 ( \64821 , \64820 );
buf \U$64848 ( \64822 , \64821 );
nand \U$64849 ( \64823 , \64816 , \64822 );
buf \U$64850 ( \64824 , \64823 );
buf \U$64851 ( \64825 , \64824 );
not \U$64852 ( \64826 , \64825 );
buf \U$64853 ( \64827 , \64826 );
buf \U$64854 ( \64828 , \64827 );
and \U$64855 ( \64829 , \64811 , \64828 );
not \U$64856 ( \64830 , \64811 );
buf \U$64857 ( \64831 , \64824 );
and \U$64858 ( \64832 , \64830 , \64831 );
nor \U$64859 ( \64833 , \64829 , \64832 );
buf \U$64860 ( \64834 , \64833 );
buf \U$64861 ( \64835 , \64834 );
buf \U$64862 ( \64836 , \63420 );
not \U$64863 ( \64837 , \64836 );
buf \U$64864 ( \64838 , \12529 );
not \U$64865 ( \64839 , \64838 );
or \U$64866 ( \64840 , \64837 , \64839 );
buf \U$64867 ( \64841 , \45728 );
buf \U$64868 ( \64842 , RIc0d8398_29);
buf \U$64869 ( \64843 , RIc0daa08_111);
xor \U$64870 ( \64844 , \64842 , \64843 );
buf \U$64871 ( \64845 , \64844 );
buf \U$64872 ( \64846 , \64845 );
nand \U$64873 ( \64847 , \64841 , \64846 );
buf \U$64874 ( \64848 , \64847 );
buf \U$64875 ( \64849 , \64848 );
nand \U$64876 ( \64850 , \64840 , \64849 );
buf \U$64877 ( \64851 , \64850 );
buf \U$64878 ( \64852 , \64851 );
xor \U$64879 ( \64853 , \64835 , \64852 );
buf \U$64880 ( \64854 , \64853 );
buf \U$64881 ( \64855 , \64854 );
xor \U$64882 ( \64856 , \64791 , \64855 );
buf \U$64883 ( \64857 , \64856 );
buf \U$64884 ( \64858 , \64857 );
nand \U$64885 ( \64859 , \64670 , \64858 );
buf \U$64886 ( \64860 , \64859 );
buf \U$64887 ( \64861 , \64860 );
buf \U$64888 ( \64862 , \64468 );
not \U$64889 ( \64863 , \64862 );
buf \U$64890 ( \64864 , \64667 );
not \U$64891 ( \64865 , \64864 );
buf \U$64892 ( \64866 , \64865 );
buf \U$64893 ( \64867 , \64866 );
nand \U$64894 ( \64868 , \64863 , \64867 );
buf \U$64895 ( \64869 , \64868 );
buf \U$64896 ( \64870 , \64869 );
nand \U$64897 ( \64871 , \64861 , \64870 );
buf \U$64898 ( \64872 , \64871 );
buf \U$64899 ( \64873 , \64872 );
xor \U$64900 ( \64874 , \64351 , \64873 );
xor \U$64901 ( \64875 , \64371 , \64388 );
and \U$64902 ( \64876 , \64875 , \64403 );
and \U$64903 ( \64877 , \64371 , \64388 );
or \U$64904 ( \64878 , \64876 , \64877 );
buf \U$64905 ( \64879 , \64878 );
buf \U$64906 ( \64880 , \64464 );
not \U$64907 ( \64881 , \64880 );
buf \U$64908 ( \64882 , \64423 );
not \U$64909 ( \64883 , \64882 );
or \U$64910 ( \64884 , \64881 , \64883 );
buf \U$64911 ( \64885 , \64464 );
buf \U$64912 ( \64886 , \64423 );
or \U$64913 ( \64887 , \64885 , \64886 );
buf \U$64914 ( \64888 , \64439 );
nand \U$64915 ( \64889 , \64887 , \64888 );
buf \U$64916 ( \64890 , \64889 );
buf \U$64917 ( \64891 , \64890 );
nand \U$64918 ( \64892 , \64884 , \64891 );
buf \U$64919 ( \64893 , \64892 );
xor \U$64920 ( \64894 , \64879 , \64893 );
buf \U$64921 ( \64895 , \64582 );
not \U$64922 ( \64896 , \64895 );
buf \U$64923 ( \64897 , \64539 );
not \U$64924 ( \64898 , \64897 );
or \U$64925 ( \64899 , \64896 , \64898 );
buf \U$64926 ( \64900 , \64539 );
buf \U$64927 ( \64901 , \64582 );
or \U$64928 ( \64902 , \64900 , \64901 );
buf \U$64929 ( \64903 , \64557 );
nand \U$64930 ( \64904 , \64902 , \64903 );
buf \U$64931 ( \64905 , \64904 );
buf \U$64932 ( \64906 , \64905 );
nand \U$64933 ( \64907 , \64899 , \64906 );
buf \U$64934 ( \64908 , \64907 );
xor \U$64935 ( \64909 , \64894 , \64908 );
buf \U$64936 ( \64910 , \64909 );
xor \U$64937 ( \64911 , \64738 , \64790 );
and \U$64938 ( \64912 , \64911 , \64855 );
and \U$64939 ( \64913 , \64738 , \64790 );
or \U$64940 ( \64914 , \64912 , \64913 );
buf \U$64941 ( \64915 , \64914 );
buf \U$64942 ( \64916 , \64915 );
xor \U$64943 ( \64917 , \64910 , \64916 );
xor \U$64944 ( \64918 , \64755 , \64772 );
and \U$64945 ( \64919 , \64918 , \64787 );
and \U$64946 ( \64920 , \64755 , \64772 );
or \U$64947 ( \64921 , \64919 , \64920 );
buf \U$64948 ( \64922 , \64921 );
buf \U$64949 ( \64923 , \64714 );
not \U$64950 ( \64924 , \64923 );
buf \U$64951 ( \64925 , \64707 );
not \U$64952 ( \64926 , \64925 );
or \U$64953 ( \64927 , \64924 , \64926 );
buf \U$64954 ( \64928 , \64734 );
nand \U$64955 ( \64929 , \64927 , \64928 );
buf \U$64956 ( \64930 , \64929 );
buf \U$64957 ( \64931 , \64930 );
buf \U$64958 ( \64932 , \64704 );
buf \U$64959 ( \64933 , \64686 );
nand \U$64960 ( \64934 , \64932 , \64933 );
buf \U$64961 ( \64935 , \64934 );
buf \U$64962 ( \64936 , \64935 );
nand \U$64963 ( \64937 , \64931 , \64936 );
buf \U$64964 ( \64938 , \64937 );
xor \U$64965 ( \64939 , \64922 , \64938 );
buf \U$64966 ( \64940 , \64827 );
not \U$64967 ( \64941 , \64940 );
buf \U$64968 ( \64942 , \64810 );
not \U$64969 ( \64943 , \64942 );
or \U$64970 ( \64944 , \64941 , \64943 );
buf \U$64971 ( \64945 , \64851 );
nand \U$64972 ( \64946 , \64944 , \64945 );
buf \U$64973 ( \64947 , \64946 );
buf \U$64974 ( \64948 , \64947 );
buf \U$64975 ( \64949 , \64807 );
buf \U$64976 ( \64950 , \64824 );
nand \U$64977 ( \64951 , \64949 , \64950 );
buf \U$64978 ( \64952 , \64951 );
buf \U$64979 ( \64953 , \64952 );
nand \U$64980 ( \64954 , \64948 , \64953 );
buf \U$64981 ( \64955 , \64954 );
xor \U$64982 ( \64956 , \64939 , \64955 );
buf \U$64983 ( \64957 , \64956 );
xor \U$64984 ( \64958 , \64917 , \64957 );
buf \U$64985 ( \64959 , \64958 );
buf \U$64986 ( \64960 , \64959 );
xor \U$64987 ( \64961 , \64874 , \64960 );
buf \U$64988 ( \64962 , \64961 );
buf \U$64989 ( \64963 , \64962 );
xor \U$64990 ( \64964 , \64345 , \64963 );
buf \U$64991 ( \64965 , \64964 );
buf \U$64992 ( \64966 , \64965 );
buf \U$64993 ( \64967 , \64277 );
buf \U$64994 ( \64968 , \63503 );
xor \U$64995 ( \64969 , \64967 , \64968 );
buf \U$64996 ( \64970 , \63851 );
xor \U$64997 ( \64971 , \64969 , \64970 );
buf \U$64998 ( \64972 , \64971 );
buf \U$64999 ( \64973 , \64972 );
xor \U$65000 ( \64974 , \63703 , \63760 );
xor \U$65001 ( \64975 , \64974 , \63822 );
buf \U$65002 ( \64976 , \64975 );
buf \U$65003 ( \64977 , \64976 );
buf \U$65004 ( \64978 , \63068 );
buf \U$65005 ( \64979 , \63132 );
xor \U$65006 ( \64980 , \64978 , \64979 );
buf \U$65007 ( \64981 , \63192 );
xnor \U$65008 ( \64982 , \64980 , \64981 );
buf \U$65009 ( \64983 , \64982 );
buf \U$65010 ( \64984 , \64983 );
xor \U$65011 ( \64985 , \64977 , \64984 );
xor \U$65012 ( \64986 , \63834 , \63842 );
xor \U$65013 ( \64987 , \64986 , \63830 );
buf \U$65014 ( \64988 , \64987 );
and \U$65015 ( \64989 , \64985 , \64988 );
and \U$65016 ( \64990 , \64977 , \64984 );
or \U$65017 ( \64991 , \64989 , \64990 );
buf \U$65018 ( \64992 , \64991 );
buf \U$65019 ( \64993 , \64992 );
buf \U$65020 ( \64994 , \64468 );
not \U$65021 ( \64995 , \64994 );
buf \U$65022 ( \64996 , \64857 );
not \U$65023 ( \64997 , \64996 );
or \U$65024 ( \64998 , \64995 , \64997 );
buf \U$65025 ( \64999 , \64468 );
buf \U$65026 ( \65000 , \64857 );
or \U$65027 ( \65001 , \64999 , \65000 );
nand \U$65028 ( \65002 , \64998 , \65001 );
buf \U$65029 ( \65003 , \65002 );
buf \U$65030 ( \65004 , \65003 );
buf \U$65031 ( \65005 , \64866 );
and \U$65032 ( \65006 , \65004 , \65005 );
not \U$65033 ( \65007 , \65004 );
buf \U$65034 ( \65008 , \64667 );
and \U$65035 ( \65009 , \65007 , \65008 );
nor \U$65036 ( \65010 , \65006 , \65009 );
buf \U$65037 ( \65011 , \65010 );
buf \U$65038 ( \65012 , \65011 );
xor \U$65039 ( \65013 , \64993 , \65012 );
xor \U$65040 ( \65014 , \63720 , \63737 );
xor \U$65041 ( \65015 , \65014 , \63755 );
buf \U$65042 ( \65016 , \65015 );
buf \U$65043 ( \65017 , \65016 );
xor \U$65044 ( \65018 , \64022 , \64041 );
xor \U$65045 ( \65019 , \65018 , \64067 );
buf \U$65046 ( \65020 , \65019 );
xor \U$65047 ( \65021 , \65017 , \65020 );
xor \U$65048 ( \65022 , \53511 , \53532 );
and \U$65049 ( \65023 , \65022 , \53554 );
and \U$65050 ( \65024 , \53511 , \53532 );
or \U$65051 ( \65025 , \65023 , \65024 );
buf \U$65052 ( \65026 , \65025 );
buf \U$65053 ( \65027 , \65026 );
buf \U$65054 ( \65028 , \53465 );
buf \U$65055 ( \65029 , \53444 );
or \U$65056 ( \65030 , \65028 , \65029 );
buf \U$65057 ( \65031 , \53487 );
nand \U$65058 ( \65032 , \65030 , \65031 );
buf \U$65059 ( \65033 , \65032 );
buf \U$65060 ( \65034 , \65033 );
buf \U$65061 ( \65035 , \53465 );
buf \U$65062 ( \65036 , \53444 );
nand \U$65063 ( \65037 , \65035 , \65036 );
buf \U$65064 ( \65038 , \65037 );
buf \U$65065 ( \65039 , \65038 );
nand \U$65066 ( \65040 , \65034 , \65039 );
buf \U$65067 ( \65041 , \65040 );
buf \U$65068 ( \65042 , \65041 );
or \U$65069 ( \65043 , \65027 , \65042 );
xor \U$65070 ( \65044 , \53655 , \53674 );
and \U$65071 ( \65045 , \65044 , \53700 );
and \U$65072 ( \65046 , \53655 , \53674 );
or \U$65073 ( \65047 , \65045 , \65046 );
buf \U$65074 ( \65048 , \65047 );
buf \U$65075 ( \65049 , \65048 );
nand \U$65076 ( \65050 , \65043 , \65049 );
buf \U$65077 ( \65051 , \65050 );
buf \U$65078 ( \65052 , \65051 );
buf \U$65079 ( \65053 , \65026 );
buf \U$65080 ( \65054 , \65041 );
nand \U$65081 ( \65055 , \65053 , \65054 );
buf \U$65082 ( \65056 , \65055 );
buf \U$65083 ( \65057 , \65056 );
nand \U$65084 ( \65058 , \65052 , \65057 );
buf \U$65085 ( \65059 , \65058 );
buf \U$65086 ( \65060 , \65059 );
and \U$65087 ( \65061 , \65021 , \65060 );
and \U$65088 ( \65062 , \65017 , \65020 );
or \U$65089 ( \65063 , \65061 , \65062 );
buf \U$65090 ( \65064 , \65063 );
buf \U$65091 ( \65065 , \65064 );
xor \U$65092 ( \65066 , \64242 , \64225 );
xor \U$65093 ( \65067 , \64260 , \65066 );
buf \U$65094 ( \65068 , \65067 );
xor \U$65095 ( \65069 , \63874 , \63895 );
xor \U$65096 ( \65070 , \65069 , \63933 );
buf \U$65097 ( \65071 , \65070 );
buf \U$65098 ( \65072 , \65071 );
xor \U$65099 ( \65073 , \65068 , \65072 );
buf \U$65100 ( \65074 , \2037 );
not \U$65101 ( \65075 , \65074 );
buf \U$65102 ( \65076 , \65075 );
buf \U$65103 ( \65077 , \65076 );
buf \U$65104 ( \65078 , \53459 );
not \U$65105 ( \65079 , \65078 );
buf \U$65106 ( \65080 , \65079 );
buf \U$65107 ( \65081 , \65080 );
or \U$65108 ( \65082 , \65077 , \65081 );
buf \U$65109 ( \65083 , \13494 );
buf \U$65110 ( \65084 , \63579 );
not \U$65111 ( \65085 , \65084 );
buf \U$65112 ( \65086 , \65085 );
buf \U$65113 ( \65087 , \65086 );
or \U$65114 ( \65088 , \65083 , \65087 );
nand \U$65115 ( \65089 , \65082 , \65088 );
buf \U$65116 ( \65090 , \65089 );
buf \U$65117 ( \65091 , \53481 );
not \U$65118 ( \65092 , \65091 );
buf \U$65119 ( \65093 , \524 );
not \U$65120 ( \65094 , \65093 );
or \U$65121 ( \65095 , \65092 , \65094 );
buf \U$65122 ( \65096 , \13293 );
buf \U$65123 ( \65097 , \63505 );
nand \U$65124 ( \65098 , \65096 , \65097 );
buf \U$65125 ( \65099 , \65098 );
buf \U$65126 ( \65100 , \65099 );
nand \U$65127 ( \65101 , \65095 , \65100 );
buf \U$65128 ( \65102 , \65101 );
or \U$65129 ( \65103 , \65090 , \65102 );
buf \U$65130 ( \65104 , \53592 );
not \U$65131 ( \65105 , \65104 );
buf \U$65132 ( \65106 , \13569 );
not \U$65133 ( \65107 , \65106 );
or \U$65134 ( \65108 , \65105 , \65107 );
buf \U$65135 ( \65109 , \4008 );
buf \U$65136 ( \65110 , \63641 );
nand \U$65137 ( \65111 , \65109 , \65110 );
buf \U$65138 ( \65112 , \65111 );
buf \U$65139 ( \65113 , \65112 );
nand \U$65140 ( \65114 , \65108 , \65113 );
buf \U$65141 ( \65115 , \65114 );
nand \U$65142 ( \65116 , \65103 , \65115 );
buf \U$65143 ( \65117 , \65090 );
buf \U$65144 ( \65118 , \65102 );
nand \U$65145 ( \65119 , \65117 , \65118 );
buf \U$65146 ( \65120 , \65119 );
nand \U$65147 ( \65121 , \65116 , \65120 );
buf \U$65148 ( \65122 , \65121 );
buf \U$65149 ( \65123 , \55821 );
not \U$65150 ( \65124 , \65123 );
buf \U$65151 ( \65125 , \14100 );
not \U$65152 ( \65126 , \65125 );
or \U$65153 ( \65127 , \65124 , \65126 );
buf \U$65154 ( \65128 , \14353 );
buf \U$65155 ( \65129 , \63765 );
nand \U$65156 ( \65130 , \65128 , \65129 );
buf \U$65157 ( \65131 , \65130 );
buf \U$65158 ( \65132 , \65131 );
nand \U$65159 ( \65133 , \65127 , \65132 );
buf \U$65160 ( \65134 , \65133 );
not \U$65161 ( \65135 , \65134 );
buf \U$65162 ( \65136 , \55855 );
not \U$65163 ( \65137 , \65136 );
buf \U$65164 ( \65138 , \26572 );
not \U$65165 ( \65139 , \65138 );
or \U$65166 ( \65140 , \65137 , \65139 );
buf \U$65167 ( \65141 , \734 );
buf \U$65168 ( \65142 , \64109 );
nand \U$65169 ( \65143 , \65141 , \65142 );
buf \U$65170 ( \65144 , \65143 );
buf \U$65171 ( \65145 , \65144 );
nand \U$65172 ( \65146 , \65140 , \65145 );
buf \U$65173 ( \65147 , \65146 );
buf \U$65174 ( \65148 , \65147 );
not \U$65175 ( \65149 , \65148 );
buf \U$65176 ( \65150 , \65149 );
nand \U$65177 ( \65151 , \65135 , \65150 );
not \U$65178 ( \65152 , \65151 );
buf \U$65179 ( \65153 , \55392 );
not \U$65180 ( \65154 , \65153 );
buf \U$65181 ( \65155 , \44382 );
not \U$65182 ( \65156 , \65155 );
or \U$65183 ( \65157 , \65154 , \65156 );
buf \U$65184 ( \65158 , \15793 );
buf \U$65185 ( \65159 , \63986 );
nand \U$65186 ( \65160 , \65158 , \65159 );
buf \U$65187 ( \65161 , \65160 );
buf \U$65188 ( \65162 , \65161 );
nand \U$65189 ( \65163 , \65157 , \65162 );
buf \U$65190 ( \65164 , \65163 );
not \U$65191 ( \65165 , \65164 );
or \U$65192 ( \65166 , \65152 , \65165 );
buf \U$65193 ( \65167 , \65147 );
buf \U$65194 ( \65168 , \65134 );
nand \U$65195 ( \65169 , \65167 , \65168 );
buf \U$65196 ( \65170 , \65169 );
nand \U$65197 ( \65171 , \65166 , \65170 );
buf \U$65198 ( \65172 , \65171 );
or \U$65199 ( \65173 , \65122 , \65172 );
buf \U$65200 ( \65174 , \53572 );
not \U$65201 ( \65175 , \65174 );
buf \U$65202 ( \65176 , \13146 );
not \U$65203 ( \65177 , \65176 );
or \U$65204 ( \65178 , \65175 , \65177 );
buf \U$65205 ( \65179 , \12937 );
buf \U$65206 ( \65180 , \63964 );
nand \U$65207 ( \65181 , \65179 , \65180 );
buf \U$65208 ( \65182 , \65181 );
buf \U$65209 ( \65183 , \65182 );
nand \U$65210 ( \65184 , \65178 , \65183 );
buf \U$65211 ( \65185 , \65184 );
buf \U$65212 ( \65186 , \65185 );
not \U$65213 ( \65187 , \65186 );
buf \U$65214 ( \65188 , \65187 );
buf \U$65215 ( \65189 , \65188 );
not \U$65216 ( \65190 , \65189 );
buf \U$65217 ( \65191 , \55839 );
not \U$65218 ( \65192 , \65191 );
buf \U$65219 ( \65193 , \14569 );
not \U$65220 ( \65194 , \65193 );
or \U$65221 ( \65195 , \65192 , \65194 );
buf \U$65222 ( \65196 , \13005 );
buf \U$65223 ( \65197 , \63782 );
nand \U$65224 ( \65198 , \65196 , \65197 );
buf \U$65225 ( \65199 , \65198 );
buf \U$65226 ( \65200 , \65199 );
nand \U$65227 ( \65201 , \65195 , \65200 );
buf \U$65228 ( \65202 , \65201 );
buf \U$65229 ( \65203 , \65202 );
not \U$65230 ( \65204 , \65203 );
buf \U$65231 ( \65205 , \65204 );
buf \U$65232 ( \65206 , \65205 );
not \U$65233 ( \65207 , \65206 );
or \U$65234 ( \65208 , \65190 , \65207 );
buf \U$65235 ( \65209 , \53608 );
not \U$65236 ( \65210 , \65209 );
buf \U$65237 ( \65211 , \13706 );
not \U$65238 ( \65212 , \65211 );
or \U$65239 ( \65213 , \65210 , \65212 );
buf \U$65240 ( \65214 , \16584 );
buf \U$65241 ( \65215 , \64051 );
nand \U$65242 ( \65216 , \65214 , \65215 );
buf \U$65243 ( \65217 , \65216 );
buf \U$65244 ( \65218 , \65217 );
nand \U$65245 ( \65219 , \65213 , \65218 );
buf \U$65246 ( \65220 , \65219 );
buf \U$65247 ( \65221 , \65220 );
nand \U$65248 ( \65222 , \65208 , \65221 );
buf \U$65249 ( \65223 , \65222 );
buf \U$65250 ( \65224 , \65223 );
buf \U$65251 ( \65225 , \65202 );
buf \U$65252 ( \65226 , \65185 );
nand \U$65253 ( \65227 , \65225 , \65226 );
buf \U$65254 ( \65228 , \65227 );
buf \U$65255 ( \65229 , \65228 );
nand \U$65256 ( \65230 , \65224 , \65229 );
buf \U$65257 ( \65231 , \65230 );
buf \U$65258 ( \65232 , \65231 );
nand \U$65259 ( \65233 , \65173 , \65232 );
buf \U$65260 ( \65234 , \65233 );
buf \U$65261 ( \65235 , \65234 );
buf \U$65262 ( \65236 , \65121 );
buf \U$65263 ( \65237 , \65171 );
nand \U$65264 ( \65238 , \65236 , \65237 );
buf \U$65265 ( \65239 , \65238 );
buf \U$65266 ( \65240 , \65239 );
nand \U$65267 ( \65241 , \65235 , \65240 );
buf \U$65268 ( \65242 , \65241 );
buf \U$65269 ( \65243 , \65242 );
xor \U$65270 ( \65244 , \65073 , \65243 );
buf \U$65271 ( \65245 , \65244 );
buf \U$65272 ( \65246 , \65245 );
xor \U$65273 ( \65247 , \65065 , \65246 );
buf \U$65274 ( \65248 , \2396 );
not \U$65275 ( \65249 , \65248 );
buf \U$65276 ( \65250 , \53830 );
not \U$65277 ( \65251 , \65250 );
and \U$65278 ( \65252 , \65249 , \65251 );
buf \U$65279 ( \65253 , \2960 );
buf \U$65280 ( \65254 , \64094 );
and \U$65281 ( \65255 , \65253 , \65254 );
nor \U$65282 ( \65256 , \65252 , \65255 );
buf \U$65283 ( \65257 , \65256 );
buf \U$65284 ( \65258 , \65257 );
not \U$65285 ( \65259 , \65258 );
buf \U$65286 ( \65260 , \65259 );
buf \U$65287 ( \65261 , \65260 );
not \U$65288 ( \65262 , \65261 );
buf \U$65289 ( \65263 , \53783 );
not \U$65290 ( \65264 , \65263 );
buf \U$65291 ( \65265 , \12578 );
not \U$65292 ( \65266 , \65265 );
or \U$65293 ( \65267 , \65264 , \65266 );
buf \U$65294 ( \65268 , \12584 );
buf \U$65295 ( \65269 , \63707 );
nand \U$65296 ( \65270 , \65268 , \65269 );
buf \U$65297 ( \65271 , \65270 );
buf \U$65298 ( \65272 , \65271 );
nand \U$65299 ( \65273 , \65267 , \65272 );
buf \U$65300 ( \65274 , \65273 );
buf \U$65301 ( \65275 , \65274 );
not \U$65302 ( \65276 , \65275 );
or \U$65303 ( \65277 , \65262 , \65276 );
buf \U$65304 ( \65278 , \65274 );
not \U$65305 ( \65279 , \65278 );
buf \U$65306 ( \65280 , \65257 );
nand \U$65307 ( \65281 , \65279 , \65280 );
buf \U$65308 ( \65282 , \65281 );
buf \U$65309 ( \65283 , \65282 );
buf \U$65310 ( \65284 , \45089 );
buf \U$65311 ( \65285 , \53665 );
or \U$65312 ( \65286 , \65284 , \65285 );
buf \U$65313 ( \65287 , \14275 );
buf \U$65314 ( \65288 , \63721 );
or \U$65315 ( \65289 , \65287 , \65288 );
nand \U$65316 ( \65290 , \65286 , \65289 );
buf \U$65317 ( \65291 , \65290 );
buf \U$65318 ( \65292 , \65291 );
nand \U$65319 ( \65293 , \65283 , \65292 );
buf \U$65320 ( \65294 , \65293 );
buf \U$65321 ( \65295 , \65294 );
nand \U$65322 ( \65296 , \65277 , \65295 );
buf \U$65323 ( \65297 , \65296 );
buf \U$65324 ( \65298 , \65297 );
not \U$65325 ( \65299 , \65298 );
buf \U$65326 ( \65300 , \63912 );
not \U$65327 ( \65301 , \65300 );
buf \U$65328 ( \65302 , \63929 );
not \U$65329 ( \65303 , \65302 );
and \U$65330 ( \65304 , \65301 , \65303 );
buf \U$65331 ( \65305 , \63912 );
buf \U$65332 ( \65306 , \63929 );
and \U$65333 ( \65307 , \65305 , \65306 );
nor \U$65334 ( \65308 , \65304 , \65307 );
buf \U$65335 ( \65309 , \65308 );
buf \U$65336 ( \65310 , \65309 );
not \U$65337 ( \65311 , \65310 );
or \U$65338 ( \65312 , \65299 , \65311 );
buf \U$65339 ( \65313 , \65297 );
buf \U$65340 ( \65314 , \65309 );
or \U$65341 ( \65315 , \65313 , \65314 );
nand \U$65342 ( \65316 , \65312 , \65315 );
buf \U$65343 ( \65317 , \65316 );
buf \U$65344 ( \65318 , \65317 );
buf \U$65345 ( \65319 , \53802 );
not \U$65346 ( \65320 , \65319 );
buf \U$65347 ( \65321 , \2607 );
not \U$65348 ( \65322 , \65321 );
or \U$65349 ( \65323 , \65320 , \65322 );
buf \U$65350 ( \65324 , \816 );
buf \U$65351 ( \65325 , \63522 );
nand \U$65352 ( \65326 , \65324 , \65325 );
buf \U$65353 ( \65327 , \65326 );
buf \U$65354 ( \65328 , \65327 );
nand \U$65355 ( \65329 , \65323 , \65328 );
buf \U$65356 ( \65330 , \65329 );
buf \U$65357 ( \65331 , \65330 );
not \U$65358 ( \65332 , \65331 );
buf \U$65359 ( \65333 , \53525 );
not \U$65360 ( \65334 , \65333 );
buf \U$65361 ( \65335 , \16989 );
not \U$65362 ( \65336 , \65335 );
or \U$65363 ( \65337 , \65334 , \65336 );
buf \U$65364 ( \65338 , \12410 );
buf \U$65365 ( \65339 , \63742 );
nand \U$65366 ( \65340 , \65338 , \65339 );
buf \U$65367 ( \65341 , \65340 );
buf \U$65368 ( \65342 , \65341 );
nand \U$65369 ( \65343 , \65337 , \65342 );
buf \U$65370 ( \65344 , \65343 );
buf \U$65371 ( \65345 , \65344 );
not \U$65372 ( \65346 , \65345 );
or \U$65373 ( \65347 , \65332 , \65346 );
buf \U$65374 ( \65348 , \65344 );
buf \U$65375 ( \65349 , \65330 );
or \U$65376 ( \65350 , \65348 , \65349 );
buf \U$65377 ( \65351 , \53504 );
not \U$65378 ( \65352 , \65351 );
buf \U$65379 ( \65353 , \2766 );
not \U$65380 ( \65354 , \65353 );
or \U$65381 ( \65355 , \65352 , \65354 );
buf \U$65382 ( \65356 , \1078 );
buf \U$65383 ( \65357 , \63900 );
nand \U$65384 ( \65358 , \65356 , \65357 );
buf \U$65385 ( \65359 , \65358 );
buf \U$65386 ( \65360 , \65359 );
nand \U$65387 ( \65361 , \65355 , \65360 );
buf \U$65388 ( \65362 , \65361 );
buf \U$65389 ( \65363 , \65362 );
nand \U$65390 ( \65364 , \65350 , \65363 );
buf \U$65391 ( \65365 , \65364 );
buf \U$65392 ( \65366 , \65365 );
nand \U$65393 ( \65367 , \65347 , \65366 );
buf \U$65394 ( \65368 , \65367 );
buf \U$65395 ( \65369 , \65368 );
not \U$65396 ( \65370 , \65369 );
buf \U$65397 ( \65371 , \65370 );
buf \U$65398 ( \65372 , \65371 );
and \U$65399 ( \65373 , \65318 , \65372 );
not \U$65400 ( \65374 , \65318 );
buf \U$65401 ( \65375 , \65368 );
and \U$65402 ( \65376 , \65374 , \65375 );
nor \U$65403 ( \65377 , \65373 , \65376 );
buf \U$65404 ( \65378 , \65377 );
buf \U$65405 ( \65379 , \65378 );
not \U$65406 ( \65380 , \65379 );
buf \U$65407 ( \65381 , \65380 );
buf \U$65408 ( \65382 , \65381 );
not \U$65409 ( \65383 , \65382 );
buf \U$65410 ( \65384 , \65185 );
not \U$65411 ( \65385 , \65384 );
buf \U$65412 ( \65386 , \65205 );
not \U$65413 ( \65387 , \65386 );
or \U$65414 ( \65388 , \65385 , \65387 );
buf \U$65415 ( \65389 , \65202 );
buf \U$65416 ( \65390 , \65188 );
nand \U$65417 ( \65391 , \65389 , \65390 );
buf \U$65418 ( \65392 , \65391 );
buf \U$65419 ( \65393 , \65392 );
nand \U$65420 ( \65394 , \65388 , \65393 );
buf \U$65421 ( \65395 , \65394 );
buf \U$65422 ( \65396 , \65395 );
buf \U$65423 ( \65397 , \65220 );
xnor \U$65424 ( \65398 , \65396 , \65397 );
buf \U$65425 ( \65399 , \65398 );
buf \U$65426 ( \65400 , \65399 );
not \U$65427 ( \65401 , \65400 );
xor \U$65428 ( \65402 , \65134 , \65150 );
xor \U$65429 ( \65403 , \65402 , \65164 );
buf \U$65430 ( \65404 , \65403 );
not \U$65431 ( \65405 , \65404 );
or \U$65432 ( \65406 , \65401 , \65405 );
xor \U$65433 ( \65407 , \65344 , \65330 );
xor \U$65434 ( \65408 , \65407 , \65362 );
buf \U$65435 ( \65409 , \65408 );
nand \U$65436 ( \65410 , \65406 , \65409 );
buf \U$65437 ( \65411 , \65410 );
buf \U$65438 ( \65412 , \65411 );
buf \U$65439 ( \65413 , \65403 );
not \U$65440 ( \65414 , \65413 );
buf \U$65441 ( \65415 , \65414 );
buf \U$65442 ( \65416 , \65415 );
buf \U$65443 ( \65417 , \65399 );
not \U$65444 ( \65418 , \65417 );
buf \U$65445 ( \65419 , \65418 );
buf \U$65446 ( \65420 , \65419 );
nand \U$65447 ( \65421 , \65416 , \65420 );
buf \U$65448 ( \65422 , \65421 );
buf \U$65449 ( \65423 , \65422 );
nand \U$65450 ( \65424 , \65412 , \65423 );
buf \U$65451 ( \65425 , \65424 );
buf \U$65452 ( \65426 , \65425 );
not \U$65453 ( \65427 , \65426 );
or \U$65454 ( \65428 , \65383 , \65427 );
buf \U$65455 ( \65429 , \65425 );
buf \U$65456 ( \65430 , \65381 );
or \U$65457 ( \65431 , \65429 , \65430 );
buf \U$65458 ( \65432 , \55341 );
not \U$65459 ( \65433 , \65432 );
buf \U$65460 ( \65434 , \573 );
not \U$65461 ( \65435 , \65434 );
or \U$65462 ( \65436 , \65433 , \65435 );
buf \U$65463 ( \65437 , \584 );
buf \U$65464 ( \65438 , \64080 );
nand \U$65465 ( \65439 , \65437 , \65438 );
buf \U$65466 ( \65440 , \65439 );
buf \U$65467 ( \65441 , \65440 );
nand \U$65468 ( \65442 , \65436 , \65441 );
buf \U$65469 ( \65443 , \65442 );
buf \U$65470 ( \65444 , \3985 );
buf \U$65471 ( \65445 , RIc0d9400_64);
nand \U$65472 ( \65446 , \65444 , \65445 );
buf \U$65473 ( \65447 , \65446 );
xor \U$65474 ( \65448 , \65443 , \65447 );
buf \U$65475 ( \65449 , \53547 );
not \U$65476 ( \65450 , \65449 );
buf \U$65477 ( \65451 , \21898 );
not \U$65478 ( \65452 , \65451 );
or \U$65479 ( \65453 , \65450 , \65452 );
buf \U$65480 ( \65454 , \12342 );
buf \U$65481 ( \65455 , \63658 );
nand \U$65482 ( \65456 , \65454 , \65455 );
buf \U$65483 ( \65457 , \65456 );
buf \U$65484 ( \65458 , \65457 );
nand \U$65485 ( \65459 , \65453 , \65458 );
buf \U$65486 ( \65460 , \65459 );
xor \U$65487 ( \65461 , \65448 , \65460 );
buf \U$65488 ( \65462 , \65461 );
not \U$65489 ( \65463 , \65462 );
buf \U$65490 ( \65464 , \65463 );
buf \U$65491 ( \65465 , \65464 );
not \U$65492 ( \65466 , \65465 );
buf \U$65493 ( \65467 , \53734 );
not \U$65494 ( \65468 , \65467 );
buf \U$65495 ( \65469 , \3534 );
not \U$65496 ( \65470 , \65469 );
or \U$65497 ( \65471 , \65468 , \65470 );
buf \U$65498 ( \65472 , \16676 );
buf \U$65499 ( \65473 , \64010 );
nand \U$65500 ( \65474 , \65472 , \65473 );
buf \U$65501 ( \65475 , \65474 );
buf \U$65502 ( \65476 , \65475 );
nand \U$65503 ( \65477 , \65471 , \65476 );
buf \U$65504 ( \65478 , \65477 );
buf \U$65505 ( \65479 , \65478 );
buf \U$65506 ( \65480 , \53437 );
not \U$65507 ( \65481 , \65480 );
not \U$65508 ( \65482 , \18008 );
buf \U$65509 ( \65483 , \65482 );
not \U$65510 ( \65484 , \65483 );
or \U$65511 ( \65485 , \65481 , \65484 );
buf \U$65512 ( \65486 , \63562 );
buf \U$65513 ( \65487 , RIc0db200_128);
nand \U$65514 ( \65488 , \65486 , \65487 );
buf \U$65515 ( \65489 , \65488 );
buf \U$65516 ( \65490 , \65489 );
nand \U$65517 ( \65491 , \65485 , \65490 );
buf \U$65518 ( \65492 , \65491 );
buf \U$65519 ( \65493 , \65492 );
xor \U$65520 ( \65494 , \65479 , \65493 );
buf \U$65521 ( \65495 , \53752 );
not \U$65522 ( \65496 , \65495 );
buf \U$65523 ( \65497 , \26466 );
not \U$65524 ( \65498 , \65497 );
or \U$65525 ( \65499 , \65496 , \65498 );
buf \U$65526 ( \65500 , \12303 );
buf \U$65527 ( \65501 , \63540 );
nand \U$65528 ( \65502 , \65500 , \65501 );
buf \U$65529 ( \65503 , \65502 );
buf \U$65530 ( \65504 , \65503 );
nand \U$65531 ( \65505 , \65499 , \65504 );
buf \U$65532 ( \65506 , \65505 );
buf \U$65533 ( \65507 , \65506 );
xnor \U$65534 ( \65508 , \65494 , \65507 );
buf \U$65535 ( \65509 , \65508 );
buf \U$65536 ( \65510 , \65509 );
not \U$65537 ( \65511 , \65510 );
buf \U$65538 ( \65512 , \65511 );
buf \U$65539 ( \65513 , \65512 );
not \U$65540 ( \65514 , \65513 );
or \U$65541 ( \65515 , \65466 , \65514 );
buf \U$65542 ( \65516 , \65461 );
not \U$65543 ( \65517 , \65516 );
buf \U$65544 ( \65518 , \65509 );
not \U$65545 ( \65519 , \65518 );
or \U$65546 ( \65520 , \65517 , \65519 );
xor \U$65547 ( \65521 , \65090 , \65115 );
xor \U$65548 ( \65522 , \65521 , \65102 );
buf \U$65549 ( \65523 , \65522 );
nand \U$65550 ( \65524 , \65520 , \65523 );
buf \U$65551 ( \65525 , \65524 );
buf \U$65552 ( \65526 , \65525 );
nand \U$65553 ( \65527 , \65515 , \65526 );
buf \U$65554 ( \65528 , \65527 );
buf \U$65555 ( \65529 , \65528 );
nand \U$65556 ( \65530 , \65431 , \65529 );
buf \U$65557 ( \65531 , \65530 );
buf \U$65558 ( \65532 , \65531 );
nand \U$65559 ( \65533 , \65428 , \65532 );
buf \U$65560 ( \65534 , \65533 );
buf \U$65561 ( \65535 , \65534 );
and \U$65562 ( \65536 , \65247 , \65535 );
and \U$65563 ( \65537 , \65065 , \65246 );
or \U$65564 ( \65538 , \65536 , \65537 );
buf \U$65565 ( \65539 , \65538 );
buf \U$65566 ( \65540 , \65539 );
xor \U$65567 ( \65541 , \65013 , \65540 );
buf \U$65568 ( \65542 , \65541 );
buf \U$65569 ( \65543 , \65542 );
xor \U$65570 ( \65544 , \64973 , \65543 );
xor \U$65571 ( \65545 , \65065 , \65246 );
xor \U$65572 ( \65546 , \65545 , \65535 );
buf \U$65573 ( \65547 , \65546 );
buf \U$65574 ( \65548 , \65547 );
buf \U$65575 ( \65549 , \53851 );
not \U$65576 ( \65550 , \65549 );
buf \U$65577 ( \65551 , \53765 );
not \U$65578 ( \65552 , \65551 );
or \U$65579 ( \65553 , \65550 , \65552 );
buf \U$65580 ( \65554 , \53848 );
not \U$65581 ( \65555 , \65554 );
buf \U$65582 ( \65556 , \53759 );
not \U$65583 ( \65557 , \65556 );
or \U$65584 ( \65558 , \65555 , \65557 );
buf \U$65585 ( \65559 , \53702 );
nand \U$65586 ( \65560 , \65558 , \65559 );
buf \U$65587 ( \65561 , \65560 );
buf \U$65588 ( \65562 , \65561 );
nand \U$65589 ( \65563 , \65553 , \65562 );
buf \U$65590 ( \65564 , \65563 );
not \U$65591 ( \65565 , \65564 );
buf \U$65592 ( \65566 , \53624 );
buf \U$65593 ( \65567 , \53490 );
nand \U$65594 ( \65568 , \65566 , \65567 );
buf \U$65595 ( \65569 , \65568 );
buf \U$65596 ( \65570 , \65569 );
buf \U$65597 ( \65571 , \53556 );
and \U$65598 ( \65572 , \65570 , \65571 );
buf \U$65599 ( \65573 , \53624 );
buf \U$65600 ( \65574 , \53490 );
nor \U$65601 ( \65575 , \65573 , \65574 );
buf \U$65602 ( \65576 , \65575 );
buf \U$65603 ( \65577 , \65576 );
nor \U$65604 ( \65578 , \65572 , \65577 );
buf \U$65605 ( \65579 , \65578 );
nand \U$65606 ( \65580 , \65565 , \65579 );
not \U$65607 ( \65581 , \65580 );
not \U$65608 ( \65582 , \55803 );
buf \U$65609 ( \65583 , \65582 );
not \U$65610 ( \65584 , \65583 );
buf \U$65611 ( \65585 , \55796 );
not \U$65612 ( \65586 , \65585 );
or \U$65613 ( \65587 , \65584 , \65586 );
buf \U$65614 ( \65588 , \55803 );
not \U$65615 ( \65589 , \65588 );
buf \U$65616 ( \65590 , \55799 );
not \U$65617 ( \65591 , \65590 );
or \U$65618 ( \65592 , \65589 , \65591 );
buf \U$65619 ( \65593 , \55865 );
nand \U$65620 ( \65594 , \65592 , \65593 );
buf \U$65621 ( \65595 , \65594 );
buf \U$65622 ( \65596 , \65595 );
nand \U$65623 ( \65597 , \65587 , \65596 );
buf \U$65624 ( \65598 , \65597 );
not \U$65625 ( \65599 , \65598 );
or \U$65626 ( \65600 , \65581 , \65599 );
buf \U$65627 ( \65601 , \65564 );
buf \U$65628 ( \65602 , \65579 );
not \U$65629 ( \65603 , \65602 );
buf \U$65630 ( \65604 , \65603 );
buf \U$65631 ( \65605 , \65604 );
nand \U$65632 ( \65606 , \65601 , \65605 );
buf \U$65633 ( \65607 , \65606 );
nand \U$65634 ( \65608 , \65600 , \65607 );
buf \U$65635 ( \65609 , \65608 );
buf \U$65636 ( \65610 , \55378 );
not \U$65637 ( \65611 , \65610 );
buf \U$65638 ( \65612 , \16382 );
not \U$65639 ( \65613 , \65612 );
or \U$65640 ( \65614 , \65611 , \65613 );
buf \U$65641 ( \65615 , \13314 );
buf \U$65642 ( \65616 , \63678 );
nand \U$65643 ( \65617 , \65615 , \65616 );
buf \U$65644 ( \65618 , \65617 );
buf \U$65645 ( \65619 , \65618 );
nand \U$65646 ( \65620 , \65614 , \65619 );
buf \U$65647 ( \65621 , \65620 );
buf \U$65648 ( \65622 , \65621 );
not \U$65649 ( \65623 , \65622 );
buf \U$65650 ( \65624 , \55347 );
buf \U$65651 ( \65625 , \55363 );
nand \U$65652 ( \65626 , \65624 , \65625 );
buf \U$65653 ( \65627 , \65626 );
buf \U$65654 ( \65628 , \65627 );
nand \U$65655 ( \65629 , \65623 , \65628 );
buf \U$65656 ( \65630 , \65629 );
buf \U$65657 ( \65631 , \65630 );
not \U$65658 ( \65632 , \65631 );
buf \U$65659 ( \65633 , \53740 );
not \U$65660 ( \65634 , \65633 );
buf \U$65661 ( \65635 , \53758 );
not \U$65662 ( \65636 , \65635 );
or \U$65663 ( \65637 , \65634 , \65636 );
buf \U$65664 ( \65638 , \53758 );
buf \U$65665 ( \65639 , \53740 );
or \U$65666 ( \65640 , \65638 , \65639 );
buf \U$65667 ( \65641 , \53720 );
nand \U$65668 ( \65642 , \65640 , \65641 );
buf \U$65669 ( \65643 , \65642 );
buf \U$65670 ( \65644 , \65643 );
nand \U$65671 ( \65645 , \65637 , \65644 );
buf \U$65672 ( \65646 , \65645 );
buf \U$65673 ( \65647 , \65646 );
not \U$65674 ( \65648 , \65647 );
or \U$65675 ( \65649 , \65632 , \65648 );
buf \U$65676 ( \65650 , \65627 );
not \U$65677 ( \65651 , \65650 );
buf \U$65678 ( \65652 , \65621 );
nand \U$65679 ( \65653 , \65651 , \65652 );
buf \U$65680 ( \65654 , \65653 );
buf \U$65681 ( \65655 , \65654 );
nand \U$65682 ( \65656 , \65649 , \65655 );
buf \U$65683 ( \65657 , \65656 );
buf \U$65684 ( \65658 , \65657 );
not \U$65685 ( \65659 , \53808 );
not \U$65686 ( \65660 , \53838 );
or \U$65687 ( \65661 , \65659 , \65660 );
not \U$65688 ( \65662 , \53811 );
not \U$65689 ( \65663 , \53841 );
or \U$65690 ( \65664 , \65662 , \65663 );
nand \U$65691 ( \65665 , \65664 , \53789 );
nand \U$65692 ( \65666 , \65661 , \65665 );
buf \U$65693 ( \65667 , \65666 );
xor \U$65694 ( \65668 , \55828 , \55846 );
and \U$65695 ( \65669 , \65668 , \55863 );
and \U$65696 ( \65670 , \55828 , \55846 );
or \U$65697 ( \65671 , \65669 , \65670 );
buf \U$65698 ( \65672 , \65671 );
buf \U$65699 ( \65673 , \65672 );
xor \U$65700 ( \65674 , \65667 , \65673 );
buf \U$65701 ( \65675 , \53578 );
not \U$65702 ( \65676 , \65675 );
buf \U$65703 ( \65677 , \53598 );
not \U$65704 ( \65678 , \65677 );
or \U$65705 ( \65679 , \65676 , \65678 );
buf \U$65706 ( \65680 , \53598 );
buf \U$65707 ( \65681 , \53578 );
or \U$65708 ( \65682 , \65680 , \65681 );
buf \U$65709 ( \65683 , \53614 );
nand \U$65710 ( \65684 , \65682 , \65683 );
buf \U$65711 ( \65685 , \65684 );
buf \U$65712 ( \65686 , \65685 );
nand \U$65713 ( \65687 , \65679 , \65686 );
buf \U$65714 ( \65688 , \65687 );
buf \U$65715 ( \65689 , \65688 );
and \U$65716 ( \65690 , \65674 , \65689 );
and \U$65717 ( \65691 , \65667 , \65673 );
or \U$65718 ( \65692 , \65690 , \65691 );
buf \U$65719 ( \65693 , \65692 );
buf \U$65720 ( \65694 , \65693 );
xor \U$65721 ( \65695 , \65658 , \65694 );
xor \U$65722 ( \65696 , \65171 , \65231 );
xor \U$65723 ( \65697 , \65696 , \65121 );
buf \U$65724 ( \65698 , \65697 );
xor \U$65725 ( \65699 , \65695 , \65698 );
buf \U$65726 ( \65700 , \65699 );
buf \U$65727 ( \65701 , \65700 );
xor \U$65728 ( \65702 , \65609 , \65701 );
buf \U$65729 ( \65703 , \65425 );
not \U$65730 ( \65704 , \65703 );
buf \U$65731 ( \65705 , \65704 );
buf \U$65732 ( \65706 , \65705 );
not \U$65733 ( \65707 , \65706 );
buf \U$65734 ( \65708 , \65378 );
not \U$65735 ( \65709 , \65708 );
buf \U$65736 ( \65710 , \65528 );
not \U$65737 ( \65711 , \65710 );
or \U$65738 ( \65712 , \65709 , \65711 );
buf \U$65739 ( \65713 , \65528 );
buf \U$65740 ( \65714 , \65378 );
or \U$65741 ( \65715 , \65713 , \65714 );
nand \U$65742 ( \65716 , \65712 , \65715 );
buf \U$65743 ( \65717 , \65716 );
buf \U$65744 ( \65718 , \65717 );
not \U$65745 ( \65719 , \65718 );
or \U$65746 ( \65720 , \65707 , \65719 );
buf \U$65747 ( \65721 , \65717 );
buf \U$65748 ( \65722 , \65705 );
or \U$65749 ( \65723 , \65721 , \65722 );
nand \U$65750 ( \65724 , \65720 , \65723 );
buf \U$65751 ( \65725 , \65724 );
buf \U$65752 ( \65726 , \65725 );
and \U$65753 ( \65727 , \65702 , \65726 );
and \U$65754 ( \65728 , \65609 , \65701 );
or \U$65755 ( \65729 , \65727 , \65728 );
buf \U$65756 ( \65730 , \65729 );
buf \U$65757 ( \65731 , \65730 );
xor \U$65758 ( \65732 , \65548 , \65731 );
xor \U$65759 ( \65733 , \65658 , \65694 );
and \U$65760 ( \65734 , \65733 , \65698 );
and \U$65761 ( \65735 , \65658 , \65694 );
or \U$65762 ( \65736 , \65734 , \65735 );
buf \U$65763 ( \65737 , \65736 );
buf \U$65764 ( \65738 , \65737 );
buf \U$65765 ( \65739 , \65309 );
not \U$65766 ( \65740 , \65739 );
buf \U$65767 ( \65741 , \65371 );
not \U$65768 ( \65742 , \65741 );
or \U$65769 ( \65743 , \65740 , \65742 );
buf \U$65770 ( \65744 , \65297 );
nand \U$65771 ( \65745 , \65743 , \65744 );
buf \U$65772 ( \65746 , \65745 );
buf \U$65773 ( \65747 , \65746 );
buf \U$65774 ( \65748 , \65309 );
not \U$65775 ( \65749 , \65748 );
buf \U$65776 ( \65750 , \65368 );
nand \U$65777 ( \65751 , \65749 , \65750 );
buf \U$65778 ( \65752 , \65751 );
buf \U$65779 ( \65753 , \65752 );
nand \U$65780 ( \65754 , \65747 , \65753 );
buf \U$65781 ( \65755 , \65754 );
buf \U$65782 ( \65756 , \65755 );
buf \U$65783 ( \65757 , \65447 );
not \U$65784 ( \65758 , \65757 );
buf \U$65785 ( \65759 , \65443 );
not \U$65786 ( \65760 , \65759 );
buf \U$65787 ( \65761 , \65760 );
buf \U$65788 ( \65762 , \65761 );
not \U$65789 ( \65763 , \65762 );
or \U$65790 ( \65764 , \65758 , \65763 );
buf \U$65791 ( \65765 , \65460 );
nand \U$65792 ( \65766 , \65764 , \65765 );
buf \U$65793 ( \65767 , \65766 );
buf \U$65794 ( \65768 , \65767 );
buf \U$65795 ( \65769 , \65447 );
not \U$65796 ( \65770 , \65769 );
buf \U$65797 ( \65771 , \65443 );
nand \U$65798 ( \65772 , \65770 , \65771 );
buf \U$65799 ( \65773 , \65772 );
buf \U$65800 ( \65774 , \65773 );
nand \U$65801 ( \65775 , \65768 , \65774 );
buf \U$65802 ( \65776 , \65775 );
buf \U$65803 ( \65777 , \65776 );
buf \U$65804 ( \65778 , \65492 );
buf \U$65805 ( \65779 , \65478 );
or \U$65806 ( \65780 , \65778 , \65779 );
buf \U$65807 ( \65781 , \65506 );
nand \U$65808 ( \65782 , \65780 , \65781 );
buf \U$65809 ( \65783 , \65782 );
buf \U$65810 ( \65784 , \65783 );
buf \U$65811 ( \65785 , \65478 );
buf \U$65812 ( \65786 , \65492 );
nand \U$65813 ( \65787 , \65785 , \65786 );
buf \U$65814 ( \65788 , \65787 );
buf \U$65815 ( \65789 , \65788 );
nand \U$65816 ( \65790 , \65784 , \65789 );
buf \U$65817 ( \65791 , \65790 );
buf \U$65818 ( \65792 , \65791 );
xor \U$65819 ( \65793 , \65777 , \65792 );
buf \U$65820 ( \65794 , \53648 );
not \U$65821 ( \65795 , \65794 );
buf \U$65822 ( \65796 , \14210 );
not \U$65823 ( \65797 , \65796 );
or \U$65824 ( \65798 , \65795 , \65797 );
buf \U$65825 ( \65799 , \20211 );
buf \U$65826 ( \65800 , \63942 );
nand \U$65827 ( \65801 , \65799 , \65800 );
buf \U$65828 ( \65802 , \65801 );
buf \U$65829 ( \65803 , \65802 );
nand \U$65830 ( \65804 , \65798 , \65803 );
buf \U$65831 ( \65805 , \65804 );
buf \U$65832 ( \65806 , \65805 );
not \U$65833 ( \65807 , \65806 );
buf \U$65834 ( \65808 , \53693 );
not \U$65835 ( \65809 , \65808 );
buf \U$65836 ( \65810 , \330 );
not \U$65837 ( \65811 , \65810 );
or \U$65838 ( \65812 , \65809 , \65811 );
buf \U$65839 ( \65813 , \344 );
buf \U$65840 ( \65814 , \64025 );
nand \U$65841 ( \65815 , \65813 , \65814 );
buf \U$65842 ( \65816 , \65815 );
buf \U$65843 ( \65817 , \65816 );
nand \U$65844 ( \65818 , \65812 , \65817 );
buf \U$65845 ( \65819 , \65818 );
buf \U$65846 ( \65820 , \65819 );
not \U$65847 ( \65821 , \65820 );
or \U$65848 ( \65822 , \65807 , \65821 );
buf \U$65849 ( \65823 , \65819 );
buf \U$65850 ( \65824 , \65805 );
or \U$65851 ( \65825 , \65823 , \65824 );
buf \U$65852 ( \65826 , \53714 );
not \U$65853 ( \65827 , \65826 );
buf \U$65854 ( \65828 , \25475 );
not \U$65855 ( \65829 , \65828 );
or \U$65856 ( \65830 , \65827 , \65829 );
buf \U$65857 ( \65831 , \12744 );
buf \U$65858 ( \65832 , \63597 );
nand \U$65859 ( \65833 , \65831 , \65832 );
buf \U$65860 ( \65834 , \65833 );
buf \U$65861 ( \65835 , \65834 );
nand \U$65862 ( \65836 , \65830 , \65835 );
buf \U$65863 ( \65837 , \65836 );
buf \U$65864 ( \65838 , \65837 );
nand \U$65865 ( \65839 , \65825 , \65838 );
buf \U$65866 ( \65840 , \65839 );
buf \U$65867 ( \65841 , \65840 );
nand \U$65868 ( \65842 , \65822 , \65841 );
buf \U$65869 ( \65843 , \65842 );
buf \U$65870 ( \65844 , \65843 );
and \U$65871 ( \65845 , \65793 , \65844 );
and \U$65872 ( \65846 , \65777 , \65792 );
or \U$65873 ( \65847 , \65845 , \65846 );
buf \U$65874 ( \65848 , \65847 );
buf \U$65875 ( \65849 , \65848 );
xor \U$65876 ( \65850 , \65756 , \65849 );
xor \U$65877 ( \65851 , \63557 , \63620 );
xor \U$65878 ( \65852 , \65851 , \63628 );
buf \U$65879 ( \65853 , \65852 );
xor \U$65880 ( \65854 , \65850 , \65853 );
buf \U$65881 ( \65855 , \65854 );
buf \U$65882 ( \65856 , \65855 );
xor \U$65883 ( \65857 , \65738 , \65856 );
xor \U$65884 ( \65858 , \65777 , \65792 );
xor \U$65885 ( \65859 , \65858 , \65844 );
buf \U$65886 ( \65860 , \65859 );
buf \U$65887 ( \65861 , \65860 );
buf \U$65888 ( \65862 , \55398 );
not \U$65889 ( \65863 , \65862 );
buf \U$65890 ( \65864 , \55384 );
not \U$65891 ( \65865 , \65864 );
or \U$65892 ( \65866 , \65863 , \65865 );
buf \U$65893 ( \65867 , \55384 );
buf \U$65894 ( \65868 , \55398 );
or \U$65895 ( \65869 , \65867 , \65868 );
buf \U$65896 ( \65870 , \55366 );
nand \U$65897 ( \65871 , \65869 , \65870 );
buf \U$65898 ( \65872 , \65871 );
buf \U$65899 ( \65873 , \65872 );
nand \U$65900 ( \65874 , \65866 , \65873 );
buf \U$65901 ( \65875 , \65874 );
buf \U$65902 ( \65876 , \65875 );
buf \U$65903 ( \65877 , \65260 );
buf \U$65904 ( \65878 , \65274 );
xor \U$65905 ( \65879 , \65877 , \65878 );
buf \U$65906 ( \65880 , \65291 );
xor \U$65907 ( \65881 , \65879 , \65880 );
buf \U$65908 ( \65882 , \65881 );
buf \U$65909 ( \65883 , \65882 );
xor \U$65910 ( \65884 , \65876 , \65883 );
xor \U$65911 ( \65885 , \65805 , \65819 );
xor \U$65912 ( \65886 , \65885 , \65837 );
buf \U$65913 ( \65887 , \65886 );
and \U$65914 ( \65888 , \65884 , \65887 );
and \U$65915 ( \65889 , \65876 , \65883 );
or \U$65916 ( \65890 , \65888 , \65889 );
buf \U$65917 ( \65891 , \65890 );
buf \U$65918 ( \65892 , \65891 );
xor \U$65919 ( \65893 , \65861 , \65892 );
xor \U$65920 ( \65894 , \63958 , \63976 );
xnor \U$65921 ( \65895 , \65894 , \63998 );
xor \U$65922 ( \65896 , \63778 , \63795 );
xor \U$65923 ( \65897 , \65896 , \63817 );
buf \U$65924 ( \65898 , \65897 );
xor \U$65925 ( \65899 , \65895 , \65898 );
xor \U$65926 ( \65900 , \63518 , \63535 );
xor \U$65927 ( \65901 , \65900 , \63553 );
buf \U$65928 ( \65902 , \65901 );
xnor \U$65929 ( \65903 , \65899 , \65902 );
buf \U$65930 ( \65904 , \65903 );
and \U$65931 ( \65905 , \65893 , \65904 );
and \U$65932 ( \65906 , \65861 , \65892 );
or \U$65933 ( \65907 , \65905 , \65906 );
buf \U$65934 ( \65908 , \65907 );
buf \U$65935 ( \65909 , \65908 );
xor \U$65936 ( \65910 , \65857 , \65909 );
buf \U$65937 ( \65911 , \65910 );
buf \U$65938 ( \65912 , \65911 );
and \U$65939 ( \65913 , \65732 , \65912 );
and \U$65940 ( \65914 , \65548 , \65731 );
or \U$65941 ( \65915 , \65913 , \65914 );
buf \U$65942 ( \65916 , \65915 );
buf \U$65943 ( \65917 , \65916 );
and \U$65944 ( \65918 , \65544 , \65917 );
and \U$65945 ( \65919 , \64973 , \65543 );
or \U$65946 ( \65920 , \65918 , \65919 );
buf \U$65947 ( \65921 , \65920 );
buf \U$65948 ( \65922 , \65921 );
xor \U$65949 ( \65923 , \64966 , \65922 );
buf \U$65950 ( \65924 , \64356 );
not \U$65951 ( \65925 , \65924 );
buf \U$65952 ( \65926 , \64405 );
not \U$65953 ( \65927 , \65926 );
or \U$65954 ( \65928 , \65925 , \65927 );
buf \U$65955 ( \65929 , \64405 );
buf \U$65956 ( \65930 , \64356 );
or \U$65957 ( \65931 , \65929 , \65930 );
buf \U$65958 ( \65932 , \64465 );
nand \U$65959 ( \65933 , \65931 , \65932 );
buf \U$65960 ( \65934 , \65933 );
buf \U$65961 ( \65935 , \65934 );
nand \U$65962 ( \65936 , \65928 , \65935 );
buf \U$65963 ( \65937 , \65936 );
buf \U$65964 ( \65938 , \64176 );
buf \U$65965 ( \65939 , \64193 );
and \U$65966 ( \65940 , \65938 , \65939 );
buf \U$65967 ( \65941 , \65940 );
buf \U$65968 ( \65942 , \65941 );
xor \U$65969 ( \65943 , \64487 , \64501 );
and \U$65970 ( \65944 , \65943 , \64521 );
and \U$65971 ( \65945 , \64487 , \64501 );
or \U$65972 ( \65946 , \65944 , \65945 );
buf \U$65973 ( \65947 , \65946 );
buf \U$65974 ( \65948 , \65947 );
xor \U$65975 ( \65949 , \65942 , \65948 );
buf \U$65976 ( \65950 , \64637 );
not \U$65977 ( \65951 , \65950 );
buf \U$65978 ( \65952 , \64616 );
not \U$65979 ( \65953 , \65952 );
or \U$65980 ( \65954 , \65951 , \65953 );
buf \U$65981 ( \65955 , \64640 );
not \U$65982 ( \65956 , \65955 );
buf \U$65983 ( \65957 , \64619 );
not \U$65984 ( \65958 , \65957 );
or \U$65985 ( \65959 , \65956 , \65958 );
buf \U$65986 ( \65960 , \64661 );
nand \U$65987 ( \65961 , \65959 , \65960 );
buf \U$65988 ( \65962 , \65961 );
buf \U$65989 ( \65963 , \65962 );
nand \U$65990 ( \65964 , \65954 , \65963 );
buf \U$65991 ( \65965 , \65964 );
buf \U$65992 ( \65966 , \65965 );
xor \U$65993 ( \65967 , \65949 , \65966 );
buf \U$65994 ( \65968 , \65967 );
xor \U$65995 ( \65969 , \65937 , \65968 );
buf \U$65996 ( \65970 , \64664 );
buf \U$65997 ( \65971 , \64523 );
or \U$65998 ( \65972 , \65970 , \65971 );
buf \U$65999 ( \65973 , \64597 );
nand \U$66000 ( \65974 , \65972 , \65973 );
buf \U$66001 ( \65975 , \65974 );
buf \U$66002 ( \65976 , \65975 );
buf \U$66003 ( \65977 , \64664 );
buf \U$66004 ( \65978 , \64523 );
nand \U$66005 ( \65979 , \65977 , \65978 );
buf \U$66006 ( \65980 , \65979 );
buf \U$66007 ( \65981 , \65980 );
nand \U$66008 ( \65982 , \65976 , \65981 );
buf \U$66009 ( \65983 , \65982 );
xor \U$66010 ( \65984 , \65969 , \65983 );
buf \U$66011 ( \65985 , \65984 );
buf \U$66012 ( \65986 , \64610 );
not \U$66013 ( \65987 , \65986 );
buf \U$66014 ( \65988 , \12402 );
not \U$66015 ( \65989 , \65988 );
or \U$66016 ( \65990 , \65987 , \65989 );
buf \U$66017 ( \65991 , \16662 );
buf \U$66018 ( \65992 , RIc0d8230_26);
buf \U$66019 ( \65993 , RIc0daaf8_113);
xor \U$66020 ( \65994 , \65992 , \65993 );
buf \U$66021 ( \65995 , \65994 );
buf \U$66022 ( \65996 , \65995 );
nand \U$66023 ( \65997 , \65991 , \65996 );
buf \U$66024 ( \65998 , \65997 );
buf \U$66025 ( \65999 , \65998 );
nand \U$66026 ( \66000 , \65990 , \65999 );
buf \U$66027 ( \66001 , \66000 );
buf \U$66028 ( \66002 , \66001 );
buf \U$66029 ( \66003 , \64494 );
not \U$66030 ( \66004 , \66003 );
buf \U$66031 ( \66005 , \14419 );
not \U$66032 ( \66006 , \66005 );
or \U$66033 ( \66007 , \66004 , \66006 );
buf \U$66034 ( \66008 , \22006 );
buf \U$66035 ( \66009 , RIc0d88c0_40);
buf \U$66036 ( \66010 , RIc0da468_99);
xor \U$66037 ( \66011 , \66009 , \66010 );
buf \U$66038 ( \66012 , \66011 );
buf \U$66039 ( \66013 , \66012 );
nand \U$66040 ( \66014 , \66008 , \66013 );
buf \U$66041 ( \66015 , \66014 );
buf \U$66042 ( \66016 , \66015 );
nand \U$66043 ( \66017 , \66007 , \66016 );
buf \U$66044 ( \66018 , \66017 );
buf \U$66045 ( \66019 , \66018 );
xor \U$66046 ( \66020 , \66002 , \66019 );
buf \U$66047 ( \66021 , \64655 );
not \U$66048 ( \66022 , \66021 );
buf \U$66049 ( \66023 , \18767 );
not \U$66050 ( \66024 , \66023 );
or \U$66051 ( \66025 , \66022 , \66024 );
buf \U$66052 ( \66026 , \2960 );
buf \U$66053 ( \66027 , RIc0d9dd8_85);
buf \U$66054 ( \66028 , RIc0d8f50_54);
xor \U$66055 ( \66029 , \66027 , \66028 );
buf \U$66056 ( \66030 , \66029 );
buf \U$66057 ( \66031 , \66030 );
nand \U$66058 ( \66032 , \66026 , \66031 );
buf \U$66059 ( \66033 , \66032 );
buf \U$66060 ( \66034 , \66033 );
nand \U$66061 ( \66035 , \66025 , \66034 );
buf \U$66062 ( \66036 , \66035 );
buf \U$66063 ( \66037 , \66036 );
xor \U$66064 ( \66038 , \66020 , \66037 );
buf \U$66065 ( \66039 , \66038 );
buf \U$66066 ( \66040 , \64533 );
not \U$66067 ( \66041 , \66040 );
buf \U$66068 ( \66042 , \13860 );
not \U$66069 ( \66043 , \66042 );
or \U$66070 ( \66044 , \66041 , \66043 );
buf \U$66071 ( \66045 , \13873 );
buf \U$66072 ( \66046 , RIc0d8aa0_44);
buf \U$66073 ( \66047 , RIc0da288_95);
xor \U$66074 ( \66048 , \66046 , \66047 );
buf \U$66075 ( \66049 , \66048 );
buf \U$66076 ( \66050 , \66049 );
nand \U$66077 ( \66051 , \66045 , \66050 );
buf \U$66078 ( \66052 , \66051 );
buf \U$66079 ( \66053 , \66052 );
nand \U$66080 ( \66054 , \66044 , \66053 );
buf \U$66081 ( \66055 , \66054 );
buf \U$66082 ( \66056 , \66055 );
buf \U$66083 ( \66057 , \64680 );
not \U$66084 ( \66058 , \66057 );
buf \U$66085 ( \66059 , \13001 );
not \U$66086 ( \66060 , \66059 );
or \U$66087 ( \66061 , \66058 , \66060 );
buf \U$66088 ( \66062 , \13005 );
buf \U$66089 ( \66063 , RIc0d7f60_20);
buf \U$66090 ( \66064 , RIc0dadc8_119);
xor \U$66091 ( \66065 , \66063 , \66064 );
buf \U$66092 ( \66066 , \66065 );
buf \U$66093 ( \66067 , \66066 );
nand \U$66094 ( \66068 , \66062 , \66067 );
buf \U$66095 ( \66069 , \66068 );
buf \U$66096 ( \66070 , \66069 );
nand \U$66097 ( \66071 , \66061 , \66070 );
buf \U$66098 ( \66072 , \66071 );
buf \U$66099 ( \66073 , \66072 );
xor \U$66100 ( \66074 , \66056 , \66073 );
buf \U$66101 ( \66075 , \64576 );
not \U$66102 ( \66076 , \66075 );
buf \U$66103 ( \66077 , \17141 );
not \U$66104 ( \66078 , \66077 );
or \U$66105 ( \66079 , \66076 , \66078 );
buf \U$66106 ( \66080 , \1078 );
xor \U$66107 ( \66081 , RIc0d9bf8_81, RIc0d9130_58);
buf \U$66108 ( \66082 , \66081 );
nand \U$66109 ( \66083 , \66080 , \66082 );
buf \U$66110 ( \66084 , \66083 );
buf \U$66111 ( \66085 , \66084 );
nand \U$66112 ( \66086 , \66079 , \66085 );
buf \U$66113 ( \66087 , \66086 );
buf \U$66114 ( \66088 , \66087 );
xor \U$66115 ( \66089 , \66074 , \66088 );
buf \U$66116 ( \66090 , \66089 );
xor \U$66117 ( \66091 , \66039 , \66090 );
buf \U$66118 ( \66092 , \64845 );
not \U$66119 ( \66093 , \66092 );
buf \U$66120 ( \66094 , \14100 );
not \U$66121 ( \66095 , \66094 );
or \U$66122 ( \66096 , \66093 , \66095 );
buf \U$66123 ( \66097 , \18312 );
buf \U$66124 ( \66098 , RIc0d8320_28);
buf \U$66125 ( \66099 , RIc0daa08_111);
xor \U$66126 ( \66100 , \66098 , \66099 );
buf \U$66127 ( \66101 , \66100 );
buf \U$66128 ( \66102 , \66101 );
nand \U$66129 ( \66103 , \66097 , \66102 );
buf \U$66130 ( \66104 , \66103 );
buf \U$66131 ( \66105 , \66104 );
nand \U$66132 ( \66106 , \66096 , \66105 );
buf \U$66133 ( \66107 , \66106 );
buf \U$66134 ( \66108 , \66107 );
buf \U$66135 ( \66109 , \64801 );
not \U$66136 ( \66110 , \66109 );
buf \U$66137 ( \66111 , \15329 );
not \U$66138 ( \66112 , \66111 );
or \U$66139 ( \66113 , \66110 , \66112 );
buf \U$66140 ( \66114 , \734 );
buf \U$66141 ( \66115 , RIc0d89b0_42);
buf \U$66142 ( \66116 , RIc0da378_97);
xor \U$66143 ( \66117 , \66115 , \66116 );
buf \U$66144 ( \66118 , \66117 );
buf \U$66145 ( \66119 , \66118 );
nand \U$66146 ( \66120 , \66114 , \66119 );
buf \U$66147 ( \66121 , \66120 );
buf \U$66148 ( \66122 , \66121 );
nand \U$66149 ( \66123 , \66113 , \66122 );
buf \U$66150 ( \66124 , \66123 );
buf \U$66151 ( \66125 , \66124 );
xor \U$66152 ( \66126 , \66108 , \66125 );
buf \U$66153 ( \66127 , \64748 );
not \U$66154 ( \66128 , \66127 );
buf \U$66155 ( \66129 , \14982 );
not \U$66156 ( \66130 , \66129 );
or \U$66157 ( \66131 , \66128 , \66130 );
buf \U$66158 ( \66132 , \16692 );
buf \U$66159 ( \66133 , RIc0dafa8_123);
buf \U$66160 ( \66134 , RIc0d7d80_16);
xor \U$66161 ( \66135 , \66133 , \66134 );
buf \U$66162 ( \66136 , \66135 );
buf \U$66163 ( \66137 , \66136 );
nand \U$66164 ( \66138 , \66132 , \66137 );
buf \U$66165 ( \66139 , \66138 );
buf \U$66166 ( \66140 , \66139 );
nand \U$66167 ( \66141 , \66131 , \66140 );
buf \U$66168 ( \66142 , \66141 );
buf \U$66169 ( \66143 , \66142 );
xor \U$66170 ( \66144 , \66126 , \66143 );
buf \U$66171 ( \66145 , \66144 );
xor \U$66172 ( \66146 , \66091 , \66145 );
buf \U$66173 ( \66147 , \66146 );
buf \U$66174 ( \66148 , \64458 );
not \U$66175 ( \66149 , \66148 );
buf \U$66176 ( \66150 , \1183 );
not \U$66177 ( \66151 , \66150 );
or \U$66178 ( \66152 , \66149 , \66151 );
buf \U$66179 ( \66153 , \14374 );
buf \U$66180 ( \66154 , RIc0d9a18_77);
buf \U$66181 ( \66155 , RIc0d9310_62);
xor \U$66182 ( \66156 , \66154 , \66155 );
buf \U$66183 ( \66157 , \66156 );
buf \U$66184 ( \66158 , \66157 );
nand \U$66185 ( \66159 , \66153 , \66158 );
buf \U$66186 ( \66160 , \66159 );
buf \U$66187 ( \66161 , \66160 );
nand \U$66188 ( \66162 , \66152 , \66161 );
buf \U$66189 ( \66163 , \66162 );
buf \U$66190 ( \66164 , \66163 );
buf \U$66191 ( \66165 , \64551 );
not \U$66192 ( \66166 , \66165 );
buf \U$66193 ( \66167 , \1736 );
not \U$66194 ( \66168 , \66167 );
or \U$66195 ( \66169 , \66166 , \66168 );
buf \U$66196 ( \66170 , \993 );
buf \U$66197 ( \66171 , RIc0d9ce8_83);
buf \U$66198 ( \66172 , RIc0d9040_56);
xor \U$66199 ( \66173 , \66171 , \66172 );
buf \U$66200 ( \66174 , \66173 );
buf \U$66201 ( \66175 , \66174 );
nand \U$66202 ( \66176 , \66170 , \66175 );
buf \U$66203 ( \66177 , \66176 );
buf \U$66204 ( \66178 , \66177 );
nand \U$66205 ( \66179 , \66169 , \66178 );
buf \U$66206 ( \66180 , \66179 );
buf \U$66207 ( \66181 , \66180 );
xor \U$66208 ( \66182 , \66164 , \66181 );
buf \U$66209 ( \66183 , \64433 );
not \U$66210 ( \66184 , \66183 );
buf \U$66211 ( \66185 , \27660 );
not \U$66212 ( \66186 , \66185 );
or \U$66213 ( \66187 , \66184 , \66186 );
buf \U$66214 ( \66188 , \16232 );
buf \U$66215 ( \66189 , RIc0da918_109);
buf \U$66216 ( \66190 , RIc0d8410_30);
xor \U$66217 ( \66191 , \66189 , \66190 );
buf \U$66218 ( \66192 , \66191 );
buf \U$66219 ( \66193 , \66192 );
nand \U$66220 ( \66194 , \66188 , \66193 );
buf \U$66221 ( \66195 , \66194 );
buf \U$66222 ( \66196 , \66195 );
nand \U$66223 ( \66197 , \66187 , \66196 );
buf \U$66224 ( \66198 , \66197 );
buf \U$66225 ( \66199 , \66198 );
xor \U$66226 ( \66200 , \66182 , \66199 );
buf \U$66227 ( \66201 , \66200 );
buf \U$66228 ( \66202 , \66201 );
buf \U$66229 ( \66203 , \64396 );
not \U$66230 ( \66204 , \66203 );
buf \U$66231 ( \66205 , \16065 );
not \U$66232 ( \66206 , \66205 );
or \U$66233 ( \66207 , \66204 , \66206 );
buf \U$66234 ( \66208 , \16071 );
xor \U$66235 ( \66209 , RIc0da828_107, RIc0d8500_32);
buf \U$66236 ( \66210 , \66209 );
nand \U$66237 ( \66211 , \66208 , \66210 );
buf \U$66238 ( \66212 , \66211 );
buf \U$66239 ( \66213 , \66212 );
nand \U$66240 ( \66214 , \66207 , \66213 );
buf \U$66241 ( \66215 , \66214 );
buf \U$66242 ( \66216 , \64381 );
not \U$66243 ( \66217 , \66216 );
buf \U$66244 ( \66218 , \12299 );
not \U$66245 ( \66219 , \66218 );
or \U$66246 ( \66220 , \66217 , \66219 );
buf \U$66247 ( \66221 , \12303 );
buf \U$66248 ( \66222 , RIc0d8140_24);
buf \U$66249 ( \66223 , RIc0dabe8_115);
xor \U$66250 ( \66224 , \66222 , \66223 );
buf \U$66251 ( \66225 , \66224 );
buf \U$66252 ( \66226 , \66225 );
nand \U$66253 ( \66227 , \66221 , \66226 );
buf \U$66254 ( \66228 , \66227 );
buf \U$66255 ( \66229 , \66228 );
nand \U$66256 ( \66230 , \66220 , \66229 );
buf \U$66257 ( \66231 , \66230 );
xor \U$66258 ( \66232 , \66215 , \66231 );
buf \U$66259 ( \66233 , \64151 );
not \U$66260 ( \66234 , \66233 );
buf \U$66261 ( \66235 , \17995 );
not \U$66262 ( \66236 , \66235 );
or \U$66263 ( \66237 , \66234 , \66236 );
buf \U$66264 ( \66238 , \13465 );
xor \U$66265 ( \66239 , RIc0db098_125, RIc0d7c90_14);
buf \U$66266 ( \66240 , \66239 );
nand \U$66267 ( \66241 , \66238 , \66240 );
buf \U$66268 ( \66242 , \66241 );
buf \U$66269 ( \66243 , \66242 );
nand \U$66270 ( \66244 , \66237 , \66243 );
buf \U$66271 ( \66245 , \66244 );
not \U$66272 ( \66246 , \66245 );
xor \U$66273 ( \66247 , \66232 , \66246 );
buf \U$66274 ( \66248 , \66247 );
not \U$66275 ( \66249 , \66248 );
buf \U$66276 ( \66250 , \66249 );
buf \U$66277 ( \66251 , \66250 );
and \U$66278 ( \66252 , \66202 , \66251 );
not \U$66279 ( \66253 , \66202 );
buf \U$66280 ( \66254 , \66247 );
and \U$66281 ( \66255 , \66253 , \66254 );
nor \U$66282 ( \66256 , \66252 , \66255 );
buf \U$66283 ( \66257 , \66256 );
buf \U$66284 ( \66258 , \66257 );
buf \U$66285 ( \66259 , \13389 );
buf \U$66286 ( \66260 , RIc0d9400_64);
nand \U$66287 ( \66261 , \66259 , \66260 );
buf \U$66288 ( \66262 , \66261 );
buf \U$66289 ( \66263 , \66262 );
buf \U$66290 ( \66264 , \64170 );
not \U$66291 ( \66265 , \66264 );
buf \U$66292 ( \66266 , \14940 );
not \U$66293 ( \66267 , \66266 );
or \U$66294 ( \66268 , \66265 , \66267 );
buf \U$66295 ( \66269 , \1025 );
buf \U$66296 ( \66270 , RIc0d9220_60);
buf \U$66297 ( \66271 , RIc0d9b08_79);
xor \U$66298 ( \66272 , \66270 , \66271 );
buf \U$66299 ( \66273 , \66272 );
buf \U$66300 ( \66274 , \66273 );
nand \U$66301 ( \66275 , \66269 , \66274 );
buf \U$66302 ( \66276 , \66275 );
buf \U$66303 ( \66277 , \66276 );
nand \U$66304 ( \66278 , \66268 , \66277 );
buf \U$66305 ( \66279 , \66278 );
buf \U$66306 ( \66280 , \66279 );
xor \U$66307 ( \66281 , \66263 , \66280 );
buf \U$66308 ( \66282 , \64417 );
not \U$66309 ( \66283 , \66282 );
buf \U$66310 ( \66284 , \22350 );
not \U$66311 ( \66285 , \66284 );
or \U$66312 ( \66286 , \66283 , \66285 );
buf \U$66313 ( \66287 , \22356 );
buf \U$66314 ( \66288 , RIc0dacd8_117);
buf \U$66315 ( \66289 , RIc0d8050_22);
xor \U$66316 ( \66290 , \66288 , \66289 );
buf \U$66317 ( \66291 , \66290 );
buf \U$66318 ( \66292 , \66291 );
nand \U$66319 ( \66293 , \66287 , \66292 );
buf \U$66320 ( \66294 , \66293 );
buf \U$66321 ( \66295 , \66294 );
nand \U$66322 ( \66296 , \66286 , \66295 );
buf \U$66323 ( \66297 , \66296 );
buf \U$66324 ( \66298 , \66297 );
xor \U$66325 ( \66299 , \66281 , \66298 );
buf \U$66326 ( \66300 , \66299 );
buf \U$66327 ( \66301 , \66300 );
not \U$66328 ( \66302 , \66301 );
buf \U$66329 ( \66303 , \66302 );
buf \U$66330 ( \66304 , \66303 );
and \U$66331 ( \66305 , \66258 , \66304 );
not \U$66332 ( \66306 , \66258 );
buf \U$66333 ( \66307 , \66300 );
and \U$66334 ( \66308 , \66306 , \66307 );
nor \U$66335 ( \66309 , \66305 , \66308 );
buf \U$66336 ( \66310 , \66309 );
buf \U$66337 ( \66311 , \66310 );
xor \U$66338 ( \66312 , \66147 , \66311 );
buf \U$66339 ( \66313 , \64479 );
not \U$66340 ( \66314 , \66313 );
buf \U$66341 ( \66315 , \44639 );
not \U$66342 ( \66316 , \66315 );
or \U$66343 ( \66317 , \66314 , \66316 );
buf \U$66344 ( \66318 , RIc0d7ba0_12);
buf \U$66345 ( \66319 , RIc0db188_127);
xor \U$66346 ( \66320 , \66318 , \66319 );
buf \U$66347 ( \66321 , \66320 );
buf \U$66348 ( \66322 , \66321 );
buf \U$66349 ( \66323 , RIc0db200_128);
nand \U$66350 ( \66324 , \66322 , \66323 );
buf \U$66351 ( \66325 , \66324 );
buf \U$66352 ( \66326 , \66325 );
nand \U$66353 ( \66327 , \66317 , \66326 );
buf \U$66354 ( \66328 , \66327 );
buf \U$66355 ( \66329 , \66328 );
buf \U$66356 ( \66330 , \64513 );
not \U$66357 ( \66331 , \66330 );
buf \U$66358 ( \66332 , \15995 );
not \U$66359 ( \66333 , \66332 );
or \U$66360 ( \66334 , \66331 , \66333 );
buf \U$66361 ( \66335 , \481 );
buf \U$66362 ( \66336 , RIc0d8b90_46);
buf \U$66363 ( \66337 , RIc0da198_93);
xor \U$66364 ( \66338 , \66336 , \66337 );
buf \U$66365 ( \66339 , \66338 );
buf \U$66366 ( \66340 , \66339 );
nand \U$66367 ( \66341 , \66335 , \66340 );
buf \U$66368 ( \66342 , \66341 );
buf \U$66369 ( \66343 , \66342 );
nand \U$66370 ( \66344 , \66334 , \66343 );
buf \U$66371 ( \66345 , \66344 );
buf \U$66372 ( \66346 , \66345 );
xor \U$66373 ( \66347 , \66329 , \66346 );
buf \U$66374 ( \66348 , \64364 );
not \U$66375 ( \66349 , \66348 );
buf \U$66376 ( \66350 , \3534 );
not \U$66377 ( \66351 , \66350 );
or \U$66378 ( \66352 , \66349 , \66351 );
buf \U$66379 ( \66353 , \16676 );
buf \U$66380 ( \66354 , RIc0da558_101);
buf \U$66381 ( \66355 , RIc0d87d0_38);
xor \U$66382 ( \66356 , \66354 , \66355 );
buf \U$66383 ( \66357 , \66356 );
buf \U$66384 ( \66358 , \66357 );
nand \U$66385 ( \66359 , \66353 , \66358 );
buf \U$66386 ( \66360 , \66359 );
buf \U$66387 ( \66361 , \66360 );
nand \U$66388 ( \66362 , \66352 , \66361 );
buf \U$66389 ( \66363 , \66362 );
buf \U$66390 ( \66364 , \66363 );
xor \U$66391 ( \66365 , \66347 , \66364 );
buf \U$66392 ( \66366 , \66365 );
buf \U$66393 ( \66367 , \66366 );
buf \U$66394 ( \66368 , \64631 );
not \U$66395 ( \66369 , \66368 );
buf \U$66396 ( \66370 , \16942 );
not \U$66397 ( \66371 , \66370 );
or \U$66398 ( \66372 , \66369 , \66371 );
buf \U$66399 ( \66373 , \13618 );
buf \U$66400 ( \66374 , RIc0d8d70_50);
buf \U$66401 ( \66375 , RIc0d9fb8_89);
xor \U$66402 ( \66376 , \66374 , \66375 );
buf \U$66403 ( \66377 , \66376 );
buf \U$66404 ( \66378 , \66377 );
nand \U$66405 ( \66379 , \66373 , \66378 );
buf \U$66406 ( \66380 , \66379 );
buf \U$66407 ( \66381 , \66380 );
nand \U$66408 ( \66382 , \66372 , \66381 );
buf \U$66409 ( \66383 , \66382 );
buf \U$66410 ( \66384 , \66383 );
buf \U$66411 ( \66385 , \64780 );
not \U$66412 ( \66386 , \66385 );
buf \U$66413 ( \66387 , \14325 );
not \U$66414 ( \66388 , \66387 );
or \U$66415 ( \66389 , \66386 , \66388 );
buf \U$66416 ( \66390 , \816 );
buf \U$66417 ( \66391 , RIc0d8e60_52);
buf \U$66418 ( \66392 , RIc0d9ec8_87);
xor \U$66419 ( \66393 , \66391 , \66392 );
buf \U$66420 ( \66394 , \66393 );
buf \U$66421 ( \66395 , \66394 );
nand \U$66422 ( \66396 , \66390 , \66395 );
buf \U$66423 ( \66397 , \66396 );
buf \U$66424 ( \66398 , \66397 );
nand \U$66425 ( \66399 , \66389 , \66398 );
buf \U$66426 ( \66400 , \66399 );
buf \U$66427 ( \66401 , \66400 );
xor \U$66428 ( \66402 , \66384 , \66401 );
buf \U$66429 ( \66403 , \64765 );
not \U$66430 ( \66404 , \66403 );
buf \U$66431 ( \66405 , \16578 );
not \U$66432 ( \66406 , \66405 );
or \U$66433 ( \66407 , \66404 , \66406 );
buf \U$66434 ( \66408 , \13048 );
xor \U$66435 ( \66409 , RIc0da648_103, RIc0d86e0_36);
buf \U$66436 ( \66410 , \66409 );
nand \U$66437 ( \66411 , \66408 , \66410 );
buf \U$66438 ( \66412 , \66411 );
buf \U$66439 ( \66413 , \66412 );
nand \U$66440 ( \66414 , \66407 , \66413 );
buf \U$66441 ( \66415 , \66414 );
buf \U$66442 ( \66416 , \66415 );
xor \U$66443 ( \66417 , \66402 , \66416 );
buf \U$66444 ( \66418 , \66417 );
buf \U$66445 ( \66419 , \66418 );
xor \U$66446 ( \66420 , \66367 , \66419 );
buf \U$66447 ( \66421 , \64728 );
not \U$66448 ( \66422 , \66421 );
buf \U$66449 ( \66423 , \16402 );
not \U$66450 ( \66424 , \66423 );
or \U$66451 ( \66425 , \66422 , \66424 );
buf \U$66452 ( \66426 , \533 );
buf \U$66453 ( \66427 , RIc0d8c80_48);
buf \U$66454 ( \66428 , RIc0da0a8_91);
xor \U$66455 ( \66429 , \66427 , \66428 );
buf \U$66456 ( \66430 , \66429 );
buf \U$66457 ( \66431 , \66430 );
nand \U$66458 ( \66432 , \66426 , \66431 );
buf \U$66459 ( \66433 , \66432 );
buf \U$66460 ( \66434 , \66433 );
nand \U$66461 ( \66435 , \66425 , \66434 );
buf \U$66462 ( \66436 , \66435 );
buf \U$66463 ( \66437 , \66436 );
buf \U$66464 ( \66438 , \64698 );
not \U$66465 ( \66439 , \66438 );
buf \U$66466 ( \66440 , \25475 );
not \U$66467 ( \66441 , \66440 );
or \U$66468 ( \66442 , \66439 , \66441 );
buf \U$66469 ( \66443 , \15653 );
buf \U$66470 ( \66444 , RIc0da738_105);
buf \U$66471 ( \66445 , RIc0d85f0_34);
xor \U$66472 ( \66446 , \66444 , \66445 );
buf \U$66473 ( \66447 , \66446 );
buf \U$66474 ( \66448 , \66447 );
nand \U$66475 ( \66449 , \66443 , \66448 );
buf \U$66476 ( \66450 , \66449 );
buf \U$66477 ( \66451 , \66450 );
nand \U$66478 ( \66452 , \66442 , \66451 );
buf \U$66479 ( \66453 , \66452 );
buf \U$66480 ( \66454 , \66453 );
xor \U$66481 ( \66455 , \66437 , \66454 );
buf \U$66482 ( \66456 , \64818 );
not \U$66483 ( \66457 , \66456 );
buf \U$66484 ( \66458 , \13310 );
not \U$66485 ( \66459 , \66458 );
or \U$66486 ( \66460 , \66457 , \66459 );
buf \U$66487 ( \66461 , \13314 );
xor \U$66488 ( \66462 , RIc0daeb8_121, RIc0d7e70_18);
buf \U$66489 ( \66463 , \66462 );
nand \U$66490 ( \66464 , \66461 , \66463 );
buf \U$66491 ( \66465 , \66464 );
buf \U$66492 ( \66466 , \66465 );
nand \U$66493 ( \66467 , \66460 , \66466 );
buf \U$66494 ( \66468 , \66467 );
buf \U$66495 ( \66469 , \66468 );
xor \U$66496 ( \66470 , \66455 , \66469 );
buf \U$66497 ( \66471 , \66470 );
buf \U$66498 ( \66472 , \66471 );
xor \U$66499 ( \66473 , \66420 , \66472 );
buf \U$66500 ( \66474 , \66473 );
buf \U$66501 ( \66475 , \66474 );
xor \U$66502 ( \66476 , \66312 , \66475 );
buf \U$66503 ( \66477 , \66476 );
buf \U$66504 ( \66478 , \66477 );
xor \U$66505 ( \66479 , \65985 , \66478 );
xor \U$66506 ( \66480 , \65068 , \65072 );
and \U$66507 ( \66481 , \66480 , \65243 );
and \U$66508 ( \66482 , \65068 , \65072 );
or \U$66509 ( \66483 , \66481 , \66482 );
buf \U$66510 ( \66484 , \66483 );
buf \U$66511 ( \66485 , \66484 );
buf \U$66512 ( \66486 , \64004 );
not \U$66513 ( \66487 , \66486 );
buf \U$66514 ( \66488 , \64076 );
not \U$66515 ( \66489 , \66488 );
or \U$66516 ( \66490 , \66487 , \66489 );
buf \U$66517 ( \66491 , \64073 );
buf \U$66518 ( \66492 , \64007 );
nand \U$66519 ( \66493 , \66491 , \66492 );
buf \U$66520 ( \66494 , \66493 );
buf \U$66521 ( \66495 , \66494 );
nand \U$66522 ( \66496 , \66490 , \66495 );
buf \U$66523 ( \66497 , \66496 );
buf \U$66524 ( \66498 , \66497 );
buf \U$66525 ( \66499 , \64126 );
xnor \U$66526 ( \66500 , \66498 , \66499 );
buf \U$66527 ( \66501 , \66500 );
buf \U$66528 ( \66502 , \66501 );
not \U$66529 ( \66503 , \66502 );
buf \U$66530 ( \66504 , \65902 );
not \U$66531 ( \66505 , \66504 );
buf \U$66532 ( \66506 , \65898 );
not \U$66533 ( \66507 , \66506 );
or \U$66534 ( \66508 , \66505 , \66507 );
buf \U$66535 ( \66509 , \65898 );
buf \U$66536 ( \66510 , \65902 );
or \U$66537 ( \66511 , \66509 , \66510 );
buf \U$66538 ( \66512 , \65895 );
not \U$66539 ( \66513 , \66512 );
buf \U$66540 ( \66514 , \66513 );
buf \U$66541 ( \66515 , \66514 );
nand \U$66542 ( \66516 , \66511 , \66515 );
buf \U$66543 ( \66517 , \66516 );
buf \U$66544 ( \66518 , \66517 );
nand \U$66545 ( \66519 , \66508 , \66518 );
buf \U$66546 ( \66520 , \66519 );
buf \U$66547 ( \66521 , \66520 );
not \U$66548 ( \66522 , \66521 );
buf \U$66549 ( \66523 , \66522 );
buf \U$66550 ( \66524 , \66523 );
not \U$66551 ( \66525 , \66524 );
or \U$66552 ( \66526 , \66503 , \66525 );
xor \U$66553 ( \66527 , \63670 , \63693 );
xor \U$66554 ( \66528 , \66527 , \63653 );
buf \U$66555 ( \66529 , \66528 );
not \U$66556 ( \66530 , \66529 );
buf \U$66557 ( \66531 , \63574 );
buf \U$66558 ( \66532 , \63609 );
xor \U$66559 ( \66533 , \66531 , \66532 );
buf \U$66560 ( \66534 , \63591 );
xnor \U$66561 ( \66535 , \66533 , \66534 );
buf \U$66562 ( \66536 , \66535 );
buf \U$66563 ( \66537 , \66536 );
not \U$66564 ( \66538 , \66537 );
or \U$66565 ( \66539 , \66530 , \66538 );
xor \U$66566 ( \66540 , \64093 , \64107 );
xor \U$66567 ( \66541 , \66540 , \64122 );
buf \U$66568 ( \66542 , \66541 );
buf \U$66569 ( \66543 , \66542 );
nand \U$66570 ( \66544 , \66539 , \66543 );
buf \U$66571 ( \66545 , \66544 );
buf \U$66572 ( \66546 , \66545 );
buf \U$66573 ( \66547 , \66536 );
not \U$66574 ( \66548 , \66547 );
buf \U$66575 ( \66549 , \66528 );
not \U$66576 ( \66550 , \66549 );
buf \U$66577 ( \66551 , \66550 );
buf \U$66578 ( \66552 , \66551 );
nand \U$66579 ( \66553 , \66548 , \66552 );
buf \U$66580 ( \66554 , \66553 );
buf \U$66581 ( \66555 , \66554 );
nand \U$66582 ( \66556 , \66546 , \66555 );
buf \U$66583 ( \66557 , \66556 );
buf \U$66584 ( \66558 , \66557 );
nand \U$66585 ( \66559 , \66526 , \66558 );
buf \U$66586 ( \66560 , \66559 );
buf \U$66587 ( \66561 , \66560 );
buf \U$66588 ( \66562 , \66501 );
not \U$66589 ( \66563 , \66562 );
buf \U$66590 ( \66564 , \66563 );
buf \U$66591 ( \66565 , \66564 );
buf \U$66592 ( \66566 , \66520 );
nand \U$66593 ( \66567 , \66565 , \66566 );
buf \U$66594 ( \66568 , \66567 );
buf \U$66595 ( \66569 , \66568 );
nand \U$66596 ( \66570 , \66561 , \66569 );
buf \U$66597 ( \66571 , \66570 );
buf \U$66598 ( \66572 , \66571 );
xor \U$66599 ( \66573 , \66485 , \66572 );
xor \U$66600 ( \66574 , \65756 , \65849 );
and \U$66601 ( \66575 , \66574 , \65853 );
and \U$66602 ( \66576 , \65756 , \65849 );
or \U$66603 ( \66577 , \66575 , \66576 );
buf \U$66604 ( \66578 , \66577 );
buf \U$66605 ( \66579 , \66578 );
and \U$66606 ( \66580 , \66573 , \66579 );
and \U$66607 ( \66581 , \66485 , \66572 );
or \U$66608 ( \66582 , \66580 , \66581 );
buf \U$66609 ( \66583 , \66582 );
buf \U$66610 ( \66584 , \66583 );
xor \U$66611 ( \66585 , \66479 , \66584 );
buf \U$66612 ( \66586 , \66585 );
buf \U$66613 ( \66587 , \66586 );
xor \U$66614 ( \66588 , \64993 , \65012 );
and \U$66615 ( \66589 , \66588 , \65540 );
and \U$66616 ( \66590 , \64993 , \65012 );
or \U$66617 ( \66591 , \66589 , \66590 );
buf \U$66618 ( \66592 , \66591 );
buf \U$66619 ( \66593 , \66592 );
xor \U$66620 ( \66594 , \66587 , \66593 );
xor \U$66621 ( \66595 , \66485 , \66572 );
xor \U$66622 ( \66596 , \66595 , \66579 );
buf \U$66623 ( \66597 , \66596 );
buf \U$66624 ( \66598 , \66597 );
xor \U$66625 ( \66599 , \65738 , \65856 );
and \U$66626 ( \66600 , \66599 , \65909 );
and \U$66627 ( \66601 , \65738 , \65856 );
or \U$66628 ( \66602 , \66600 , \66601 );
buf \U$66629 ( \66603 , \66602 );
buf \U$66630 ( \66604 , \66603 );
xor \U$66631 ( \66605 , \66598 , \66604 );
buf \U$66632 ( \66606 , \66520 );
not \U$66633 ( \66607 , \66606 );
buf \U$66634 ( \66608 , \66557 );
not \U$66635 ( \66609 , \66608 );
buf \U$66636 ( \66610 , \66609 );
buf \U$66637 ( \66611 , \66610 );
not \U$66638 ( \66612 , \66611 );
or \U$66639 ( \66613 , \66607 , \66612 );
buf \U$66640 ( \66614 , \66610 );
buf \U$66641 ( \66615 , \66520 );
or \U$66642 ( \66616 , \66614 , \66615 );
nand \U$66643 ( \66617 , \66613 , \66616 );
buf \U$66644 ( \66618 , \66617 );
buf \U$66645 ( \66619 , \66618 );
buf \U$66646 ( \66620 , \66564 );
and \U$66647 ( \66621 , \66619 , \66620 );
not \U$66648 ( \66622 , \66619 );
buf \U$66649 ( \66623 , \66501 );
and \U$66650 ( \66624 , \66622 , \66623 );
nor \U$66651 ( \66625 , \66621 , \66624 );
buf \U$66652 ( \66626 , \66625 );
buf \U$66653 ( \66627 , \66626 );
buf \U$66654 ( \66628 , \66528 );
not \U$66655 ( \66629 , \66628 );
xnor \U$66656 ( \66630 , \66536 , \66542 );
buf \U$66657 ( \66631 , \66630 );
not \U$66658 ( \66632 , \66631 );
or \U$66659 ( \66633 , \66629 , \66632 );
buf \U$66660 ( \66634 , \66630 );
buf \U$66661 ( \66635 , \66528 );
or \U$66662 ( \66636 , \66634 , \66635 );
nand \U$66663 ( \66637 , \66633 , \66636 );
buf \U$66664 ( \66638 , \66637 );
buf \U$66665 ( \66639 , \66638 );
xor \U$66666 ( \66640 , \65017 , \65020 );
xor \U$66667 ( \66641 , \66640 , \65060 );
buf \U$66668 ( \66642 , \66641 );
buf \U$66669 ( \66643 , \66642 );
xor \U$66670 ( \66644 , \66639 , \66643 );
buf \U$66671 ( \66645 , \55920 );
not \U$66672 ( \66646 , \66645 );
buf \U$66673 ( \66647 , \55935 );
not \U$66674 ( \66648 , \66647 );
or \U$66675 ( \66649 , \66646 , \66648 );
buf \U$66676 ( \66650 , \55920 );
buf \U$66677 ( \66651 , \55935 );
or \U$66678 ( \66652 , \66650 , \66651 );
buf \U$66679 ( \66653 , \55942 );
nand \U$66680 ( \66654 , \66652 , \66653 );
buf \U$66681 ( \66655 , \66654 );
buf \U$66682 ( \66656 , \66655 );
nand \U$66683 ( \66657 , \66649 , \66656 );
buf \U$66684 ( \66658 , \66657 );
buf \U$66685 ( \66659 , \66658 );
not \U$66686 ( \66660 , \66659 );
buf \U$66687 ( \66661 , \65646 );
not \U$66688 ( \66662 , \66661 );
buf \U$66689 ( \66663 , \65627 );
not \U$66690 ( \66664 , \66663 );
buf \U$66691 ( \66665 , \65621 );
not \U$66692 ( \66666 , \66665 );
and \U$66693 ( \66667 , \66664 , \66666 );
buf \U$66694 ( \66668 , \65627 );
buf \U$66695 ( \66669 , \65621 );
and \U$66696 ( \66670 , \66668 , \66669 );
nor \U$66697 ( \66671 , \66667 , \66670 );
buf \U$66698 ( \66672 , \66671 );
buf \U$66699 ( \66673 , \66672 );
not \U$66700 ( \66674 , \66673 );
and \U$66701 ( \66675 , \66662 , \66674 );
buf \U$66702 ( \66676 , \65646 );
buf \U$66703 ( \66677 , \66672 );
and \U$66704 ( \66678 , \66676 , \66677 );
nor \U$66705 ( \66679 , \66675 , \66678 );
buf \U$66706 ( \66680 , \66679 );
buf \U$66707 ( \66681 , \66680 );
not \U$66708 ( \66682 , \66681 );
buf \U$66709 ( \66683 , \66682 );
buf \U$66710 ( \66684 , \66683 );
not \U$66711 ( \66685 , \66684 );
or \U$66712 ( \66686 , \66660 , \66685 );
buf \U$66713 ( \66687 , \66683 );
buf \U$66714 ( \66688 , \66658 );
or \U$66715 ( \66689 , \66687 , \66688 );
buf \U$66716 ( \66690 , \55974 );
not \U$66717 ( \66691 , \66690 );
buf \U$66718 ( \66692 , \55960 );
not \U$66719 ( \66693 , \66692 );
or \U$66720 ( \66694 , \66691 , \66693 );
buf \U$66721 ( \66695 , \55960 );
buf \U$66722 ( \66696 , \55974 );
or \U$66723 ( \66697 , \66695 , \66696 );
buf \U$66724 ( \66698 , \55980 );
nand \U$66725 ( \66699 , \66697 , \66698 );
buf \U$66726 ( \66700 , \66699 );
buf \U$66727 ( \66701 , \66700 );
nand \U$66728 ( \66702 , \66694 , \66701 );
buf \U$66729 ( \66703 , \66702 );
buf \U$66730 ( \66704 , \66703 );
nand \U$66731 ( \66705 , \66689 , \66704 );
buf \U$66732 ( \66706 , \66705 );
buf \U$66733 ( \66707 , \66706 );
nand \U$66734 ( \66708 , \66686 , \66707 );
buf \U$66735 ( \66709 , \66708 );
buf \U$66736 ( \66710 , \66709 );
and \U$66737 ( \66711 , \66644 , \66710 );
and \U$66738 ( \66712 , \66639 , \66643 );
or \U$66739 ( \66713 , \66711 , \66712 );
buf \U$66740 ( \66714 , \66713 );
buf \U$66741 ( \66715 , \66714 );
xor \U$66742 ( \66716 , \66627 , \66715 );
xor \U$66743 ( \66717 , \64977 , \64984 );
xor \U$66744 ( \66718 , \66717 , \64988 );
buf \U$66745 ( \66719 , \66718 );
buf \U$66746 ( \66720 , \66719 );
and \U$66747 ( \66721 , \66716 , \66720 );
and \U$66748 ( \66722 , \66627 , \66715 );
or \U$66749 ( \66723 , \66721 , \66722 );
buf \U$66750 ( \66724 , \66723 );
buf \U$66751 ( \66725 , \66724 );
and \U$66752 ( \66726 , \66605 , \66725 );
and \U$66753 ( \66727 , \66598 , \66604 );
or \U$66754 ( \66728 , \66726 , \66727 );
buf \U$66755 ( \66729 , \66728 );
buf \U$66756 ( \66730 , \66729 );
xor \U$66757 ( \66731 , \66594 , \66730 );
buf \U$66758 ( \66732 , \66731 );
buf \U$66759 ( \66733 , \66732 );
and \U$66760 ( \66734 , \65923 , \66733 );
and \U$66761 ( \66735 , \64966 , \65922 );
or \U$66762 ( \66736 , \66734 , \66735 );
buf \U$66763 ( \66737 , \66736 );
buf \U$66764 ( \66738 , \66737 );
not \U$66765 ( \66739 , \66738 );
buf \U$66766 ( \66740 , \65968 );
not \U$66767 ( \66741 , \66740 );
buf \U$66768 ( \66742 , \65937 );
not \U$66769 ( \66743 , \66742 );
or \U$66770 ( \66744 , \66741 , \66743 );
buf \U$66771 ( \66745 , \65937 );
buf \U$66772 ( \66746 , \65968 );
or \U$66773 ( \66747 , \66745 , \66746 );
buf \U$66774 ( \66748 , \65983 );
nand \U$66775 ( \66749 , \66747 , \66748 );
buf \U$66776 ( \66750 , \66749 );
buf \U$66777 ( \66751 , \66750 );
nand \U$66778 ( \66752 , \66744 , \66751 );
buf \U$66779 ( \66753 , \66752 );
xor \U$66780 ( \66754 , \64316 , \64331 );
and \U$66781 ( \66755 , \66754 , \64338 );
and \U$66782 ( \66756 , \64316 , \64331 );
or \U$66783 ( \66757 , \66755 , \66756 );
buf \U$66784 ( \66758 , \66757 );
buf \U$66785 ( \66759 , \66758 );
not \U$66786 ( \66760 , \66759 );
buf \U$66787 ( \66761 , \66760 );
xor \U$66788 ( \66762 , \66753 , \66761 );
buf \U$66789 ( \66763 , \64938 );
not \U$66790 ( \66764 , \66763 );
buf \U$66791 ( \66765 , \64955 );
not \U$66792 ( \66766 , \66765 );
or \U$66793 ( \66767 , \66764 , \66766 );
buf \U$66794 ( \66768 , \64955 );
buf \U$66795 ( \66769 , \64938 );
or \U$66796 ( \66770 , \66768 , \66769 );
buf \U$66797 ( \66771 , \64922 );
nand \U$66798 ( \66772 , \66770 , \66771 );
buf \U$66799 ( \66773 , \66772 );
buf \U$66800 ( \66774 , \66773 );
nand \U$66801 ( \66775 , \66767 , \66774 );
buf \U$66802 ( \66776 , \66775 );
buf \U$66803 ( \66777 , \65965 );
buf \U$66804 ( \66778 , \65941 );
or \U$66805 ( \66779 , \66777 , \66778 );
buf \U$66806 ( \66780 , \65947 );
nand \U$66807 ( \66781 , \66779 , \66780 );
buf \U$66808 ( \66782 , \66781 );
buf \U$66809 ( \66783 , \66782 );
buf \U$66810 ( \66784 , \65965 );
buf \U$66811 ( \66785 , \65941 );
nand \U$66812 ( \66786 , \66784 , \66785 );
buf \U$66813 ( \66787 , \66786 );
buf \U$66814 ( \66788 , \66787 );
nand \U$66815 ( \66789 , \66783 , \66788 );
buf \U$66816 ( \66790 , \66789 );
buf \U$66817 ( \66791 , \66790 );
not \U$66818 ( \66792 , \66791 );
buf \U$66819 ( \66793 , \66792 );
xor \U$66820 ( \66794 , \66776 , \66793 );
buf \U$66821 ( \66795 , \64908 );
not \U$66822 ( \66796 , \66795 );
buf \U$66823 ( \66797 , \64879 );
not \U$66824 ( \66798 , \66797 );
or \U$66825 ( \66799 , \66796 , \66798 );
buf \U$66826 ( \66800 , \64879 );
buf \U$66827 ( \66801 , \64908 );
or \U$66828 ( \66802 , \66800 , \66801 );
buf \U$66829 ( \66803 , \64893 );
nand \U$66830 ( \66804 , \66802 , \66803 );
buf \U$66831 ( \66805 , \66804 );
buf \U$66832 ( \66806 , \66805 );
nand \U$66833 ( \66807 , \66799 , \66806 );
buf \U$66834 ( \66808 , \66807 );
buf \U$66835 ( \66809 , \66808 );
not \U$66836 ( \66810 , \66809 );
buf \U$66837 ( \66811 , \66810 );
xnor \U$66838 ( \66812 , \66794 , \66811 );
buf \U$66839 ( \66813 , \66812 );
not \U$66840 ( \66814 , \66813 );
buf \U$66841 ( \66815 , \66814 );
xnor \U$66842 ( \66816 , \66762 , \66815 );
xor \U$66843 ( \66817 , \64351 , \64873 );
and \U$66844 ( \66818 , \66817 , \64960 );
and \U$66845 ( \66819 , \64351 , \64873 );
or \U$66846 ( \66820 , \66818 , \66819 );
buf \U$66847 ( \66821 , \66820 );
xor \U$66848 ( \66822 , \66816 , \66821 );
xor \U$66849 ( \66823 , \66384 , \66401 );
and \U$66850 ( \66824 , \66823 , \66416 );
and \U$66851 ( \66825 , \66384 , \66401 );
or \U$66852 ( \66826 , \66824 , \66825 );
buf \U$66853 ( \66827 , \66826 );
buf \U$66854 ( \66828 , \66827 );
buf \U$66855 ( \66829 , \66231 );
not \U$66856 ( \66830 , \66829 );
buf \U$66857 ( \66831 , \66215 );
not \U$66858 ( \66832 , \66831 );
or \U$66859 ( \66833 , \66830 , \66832 );
buf \U$66860 ( \66834 , \66215 );
buf \U$66861 ( \66835 , \66231 );
or \U$66862 ( \66836 , \66834 , \66835 );
buf \U$66863 ( \66837 , \66245 );
nand \U$66864 ( \66838 , \66836 , \66837 );
buf \U$66865 ( \66839 , \66838 );
buf \U$66866 ( \66840 , \66839 );
nand \U$66867 ( \66841 , \66833 , \66840 );
buf \U$66868 ( \66842 , \66841 );
buf \U$66869 ( \66843 , \66842 );
xor \U$66870 ( \66844 , \66828 , \66843 );
xor \U$66871 ( \66845 , \66002 , \66019 );
and \U$66872 ( \66846 , \66845 , \66037 );
and \U$66873 ( \66847 , \66002 , \66019 );
or \U$66874 ( \66848 , \66846 , \66847 );
buf \U$66875 ( \66849 , \66848 );
buf \U$66876 ( \66850 , \66849 );
xor \U$66877 ( \66851 , \66844 , \66850 );
buf \U$66878 ( \66852 , \66851 );
buf \U$66879 ( \66853 , \66852 );
not \U$66880 ( \66854 , \66853 );
buf \U$66881 ( \66855 , \66039 );
not \U$66882 ( \66856 , \66855 );
buf \U$66883 ( \66857 , \66090 );
not \U$66884 ( \66858 , \66857 );
or \U$66885 ( \66859 , \66856 , \66858 );
buf \U$66886 ( \66860 , \66039 );
buf \U$66887 ( \66861 , \66090 );
or \U$66888 ( \66862 , \66860 , \66861 );
buf \U$66889 ( \66863 , \66145 );
nand \U$66890 ( \66864 , \66862 , \66863 );
buf \U$66891 ( \66865 , \66864 );
buf \U$66892 ( \66866 , \66865 );
nand \U$66893 ( \66867 , \66859 , \66866 );
buf \U$66894 ( \66868 , \66867 );
buf \U$66895 ( \66869 , \66868 );
buf \U$66896 ( \66870 , \66418 );
not \U$66897 ( \66871 , \66870 );
buf \U$66898 ( \66872 , \66366 );
not \U$66899 ( \66873 , \66872 );
or \U$66900 ( \66874 , \66871 , \66873 );
buf \U$66901 ( \66875 , \66366 );
buf \U$66902 ( \66876 , \66418 );
or \U$66903 ( \66877 , \66875 , \66876 );
buf \U$66904 ( \66878 , \66471 );
nand \U$66905 ( \66879 , \66877 , \66878 );
buf \U$66906 ( \66880 , \66879 );
buf \U$66907 ( \66881 , \66880 );
nand \U$66908 ( \66882 , \66874 , \66881 );
buf \U$66909 ( \66883 , \66882 );
buf \U$66910 ( \66884 , \66883 );
xnor \U$66911 ( \66885 , \66869 , \66884 );
buf \U$66912 ( \66886 , \66885 );
buf \U$66913 ( \66887 , \66886 );
not \U$66914 ( \66888 , \66887 );
or \U$66915 ( \66889 , \66854 , \66888 );
buf \U$66916 ( \66890 , \66886 );
buf \U$66917 ( \66891 , \66852 );
or \U$66918 ( \66892 , \66890 , \66891 );
nand \U$66919 ( \66893 , \66889 , \66892 );
buf \U$66920 ( \66894 , \66893 );
buf \U$66921 ( \66895 , \66894 );
buf \U$66922 ( \66896 , \66300 );
not \U$66923 ( \66897 , \66896 );
buf \U$66924 ( \66898 , \66247 );
not \U$66925 ( \66899 , \66898 );
or \U$66926 ( \66900 , \66897 , \66899 );
buf \U$66927 ( \66901 , \66201 );
nand \U$66928 ( \66902 , \66900 , \66901 );
buf \U$66929 ( \66903 , \66902 );
buf \U$66930 ( \66904 , \66903 );
buf \U$66931 ( \66905 , \66250 );
buf \U$66932 ( \66906 , \66303 );
nand \U$66933 ( \66907 , \66905 , \66906 );
buf \U$66934 ( \66908 , \66907 );
buf \U$66935 ( \66909 , \66908 );
nand \U$66936 ( \66910 , \66904 , \66909 );
buf \U$66937 ( \66911 , \66910 );
xor \U$66938 ( \66912 , \66108 , \66125 );
and \U$66939 ( \66913 , \66912 , \66143 );
and \U$66940 ( \66914 , \66108 , \66125 );
or \U$66941 ( \66915 , \66913 , \66914 );
buf \U$66942 ( \66916 , \66915 );
buf \U$66943 ( \66917 , \66916 );
xor \U$66944 ( \66918 , \66056 , \66073 );
and \U$66945 ( \66919 , \66918 , \66088 );
and \U$66946 ( \66920 , \66056 , \66073 );
or \U$66947 ( \66921 , \66919 , \66920 );
buf \U$66948 ( \66922 , \66921 );
buf \U$66949 ( \66923 , \66922 );
xor \U$66950 ( \66924 , \66917 , \66923 );
xor \U$66951 ( \66925 , \66437 , \66454 );
and \U$66952 ( \66926 , \66925 , \66469 );
and \U$66953 ( \66927 , \66437 , \66454 );
or \U$66954 ( \66928 , \66926 , \66927 );
buf \U$66955 ( \66929 , \66928 );
buf \U$66956 ( \66930 , \66929 );
xor \U$66957 ( \66931 , \66924 , \66930 );
buf \U$66958 ( \66932 , \66931 );
xor \U$66959 ( \66933 , \66911 , \66932 );
buf \U$66960 ( \66934 , \66279 );
buf \U$66961 ( \66935 , \66262 );
not \U$66962 ( \66936 , \66935 );
buf \U$66963 ( \66937 , \66936 );
buf \U$66964 ( \66938 , \66937 );
or \U$66965 ( \66939 , \66934 , \66938 );
buf \U$66966 ( \66940 , \66297 );
nand \U$66967 ( \66941 , \66939 , \66940 );
buf \U$66968 ( \66942 , \66941 );
buf \U$66969 ( \66943 , \66942 );
buf \U$66970 ( \66944 , \66279 );
buf \U$66971 ( \66945 , \66937 );
nand \U$66972 ( \66946 , \66944 , \66945 );
buf \U$66973 ( \66947 , \66946 );
buf \U$66974 ( \66948 , \66947 );
nand \U$66975 ( \66949 , \66943 , \66948 );
buf \U$66976 ( \66950 , \66949 );
buf \U$66977 ( \66951 , \66950 );
xor \U$66978 ( \66952 , \66329 , \66346 );
and \U$66979 ( \66953 , \66952 , \66364 );
and \U$66980 ( \66954 , \66329 , \66346 );
or \U$66981 ( \66955 , \66953 , \66954 );
buf \U$66982 ( \66956 , \66955 );
buf \U$66983 ( \66957 , \66956 );
xor \U$66984 ( \66958 , \66951 , \66957 );
xor \U$66985 ( \66959 , \66164 , \66181 );
and \U$66986 ( \66960 , \66959 , \66199 );
and \U$66987 ( \66961 , \66164 , \66181 );
or \U$66988 ( \66962 , \66960 , \66961 );
buf \U$66989 ( \66963 , \66962 );
buf \U$66990 ( \66964 , \66963 );
xor \U$66991 ( \66965 , \66958 , \66964 );
buf \U$66992 ( \66966 , \66965 );
xor \U$66993 ( \66967 , \66933 , \66966 );
buf \U$66994 ( \66968 , \66967 );
xor \U$66995 ( \66969 , \66895 , \66968 );
xor \U$66996 ( \66970 , \64910 , \64916 );
and \U$66997 ( \66971 , \66970 , \64957 );
and \U$66998 ( \66972 , \64910 , \64916 );
or \U$66999 ( \66973 , \66971 , \66972 );
buf \U$67000 ( \66974 , \66973 );
buf \U$67001 ( \66975 , \66974 );
xor \U$67002 ( \66976 , \66969 , \66975 );
buf \U$67003 ( \66977 , \66976 );
xor \U$67004 ( \66978 , \66822 , \66977 );
buf \U$67005 ( \66979 , \66978 );
xor \U$67006 ( \66980 , \66587 , \66593 );
and \U$67007 ( \66981 , \66980 , \66730 );
and \U$67008 ( \66982 , \66587 , \66593 );
or \U$67009 ( \66983 , \66981 , \66982 );
buf \U$67010 ( \66984 , \66983 );
buf \U$67011 ( \66985 , \66984 );
xor \U$67012 ( \66986 , \66979 , \66985 );
xor \U$67013 ( \66987 , \65985 , \66478 );
and \U$67014 ( \66988 , \66987 , \66584 );
and \U$67015 ( \66989 , \65985 , \66478 );
or \U$67016 ( \66990 , \66988 , \66989 );
buf \U$67017 ( \66991 , \66990 );
buf \U$67018 ( \66992 , \66991 );
xor \U$67019 ( \66993 , \66147 , \66311 );
and \U$67020 ( \66994 , \66993 , \66475 );
and \U$67021 ( \66995 , \66147 , \66311 );
or \U$67022 ( \66996 , \66994 , \66995 );
buf \U$67023 ( \66997 , \66996 );
buf \U$67024 ( \66998 , \66997 );
buf \U$67025 ( \66999 , \59143 );
buf \U$67026 ( \67000 , \66321 );
not \U$67027 ( \67001 , \67000 );
buf \U$67028 ( \67002 , \67001 );
buf \U$67029 ( \67003 , \67002 );
or \U$67030 ( \67004 , \66999 , \67003 );
buf \U$67031 ( \67005 , RIc0d7b28_11);
buf \U$67032 ( \67006 , RIc0db188_127);
xor \U$67033 ( \67007 , \67005 , \67006 );
buf \U$67034 ( \67008 , \67007 );
buf \U$67035 ( \67009 , \67008 );
buf \U$67036 ( \67010 , RIc0db200_128);
nand \U$67037 ( \67011 , \67009 , \67010 );
buf \U$67038 ( \67012 , \67011 );
buf \U$67039 ( \67013 , \67012 );
nand \U$67040 ( \67014 , \67004 , \67013 );
buf \U$67041 ( \67015 , \67014 );
buf \U$67042 ( \67016 , \67015 );
buf \U$67043 ( \67017 , \65995 );
not \U$67044 ( \67018 , \67017 );
buf \U$67045 ( \67019 , \28413 );
not \U$67046 ( \67020 , \67019 );
or \U$67047 ( \67021 , \67018 , \67020 );
buf \U$67048 ( \67022 , \12410 );
xor \U$67049 ( \67023 , RIc0daaf8_113, RIc0d81b8_25);
buf \U$67050 ( \67024 , \67023 );
nand \U$67051 ( \67025 , \67022 , \67024 );
buf \U$67052 ( \67026 , \67025 );
buf \U$67053 ( \67027 , \67026 );
nand \U$67054 ( \67028 , \67021 , \67027 );
buf \U$67055 ( \67029 , \67028 );
buf \U$67056 ( \67030 , \67029 );
xor \U$67057 ( \67031 , \67016 , \67030 );
buf \U$67058 ( \67032 , \66447 );
not \U$67059 ( \67033 , \67032 );
buf \U$67060 ( \67034 , \12736 );
not \U$67061 ( \67035 , \67034 );
or \U$67062 ( \67036 , \67033 , \67035 );
buf \U$67063 ( \67037 , RIc0d8578_33);
buf \U$67064 ( \67038 , RIc0da738_105);
xnor \U$67065 ( \67039 , \67037 , \67038 );
buf \U$67066 ( \67040 , \67039 );
buf \U$67067 ( \67041 , \67040 );
not \U$67068 ( \67042 , \67041 );
buf \U$67069 ( \67043 , \12744 );
nand \U$67070 ( \67044 , \67042 , \67043 );
buf \U$67071 ( \67045 , \67044 );
buf \U$67072 ( \67046 , \67045 );
nand \U$67073 ( \67047 , \67036 , \67046 );
buf \U$67074 ( \67048 , \67047 );
buf \U$67075 ( \67049 , \67048 );
xor \U$67076 ( \67050 , \67031 , \67049 );
buf \U$67077 ( \67051 , \67050 );
buf \U$67078 ( \67052 , \67051 );
buf \U$67079 ( \67053 , \66273 );
not \U$67080 ( \67054 , \67053 );
buf \U$67081 ( \67055 , \14940 );
not \U$67082 ( \67056 , \67055 );
or \U$67083 ( \67057 , \67054 , \67056 );
buf \U$67084 ( \67058 , \1025 );
xor \U$67085 ( \67059 , RIc0d9b08_79, RIc0d91a8_59);
buf \U$67086 ( \67060 , \67059 );
nand \U$67087 ( \67061 , \67058 , \67060 );
buf \U$67088 ( \67062 , \67061 );
buf \U$67089 ( \67063 , \67062 );
nand \U$67090 ( \67064 , \67057 , \67063 );
buf \U$67091 ( \67065 , \67064 );
buf \U$67092 ( \67066 , \66081 );
not \U$67093 ( \67067 , \67066 );
buf \U$67094 ( \67068 , \17141 );
not \U$67095 ( \67069 , \67068 );
or \U$67096 ( \67070 , \67067 , \67069 );
buf \U$67097 ( \67071 , \1078 );
buf \U$67098 ( \67072 , RIc0d9bf8_81);
buf \U$67099 ( \67073 , RIc0d90b8_57);
xor \U$67100 ( \67074 , \67072 , \67073 );
buf \U$67101 ( \67075 , \67074 );
buf \U$67102 ( \67076 , \67075 );
nand \U$67103 ( \67077 , \67071 , \67076 );
buf \U$67104 ( \67078 , \67077 );
buf \U$67105 ( \67079 , \67078 );
nand \U$67106 ( \67080 , \67070 , \67079 );
buf \U$67107 ( \67081 , \67080 );
xor \U$67108 ( \67082 , \67065 , \67081 );
buf \U$67109 ( \67083 , \66339 );
not \U$67110 ( \67084 , \67083 );
buf \U$67111 ( \67085 , \476 );
not \U$67112 ( \67086 , \67085 );
or \U$67113 ( \67087 , \67084 , \67086 );
buf \U$67114 ( \67088 , \4008 );
buf \U$67115 ( \67089 , RIc0d8b18_45);
buf \U$67116 ( \67090 , RIc0da198_93);
xor \U$67117 ( \67091 , \67089 , \67090 );
buf \U$67118 ( \67092 , \67091 );
buf \U$67119 ( \67093 , \67092 );
nand \U$67120 ( \67094 , \67088 , \67093 );
buf \U$67121 ( \67095 , \67094 );
buf \U$67122 ( \67096 , \67095 );
nand \U$67123 ( \67097 , \67087 , \67096 );
buf \U$67124 ( \67098 , \67097 );
xor \U$67125 ( \67099 , \67082 , \67098 );
buf \U$67126 ( \67100 , \67099 );
xor \U$67127 ( \67101 , \67052 , \67100 );
buf \U$67128 ( \67102 , \66430 );
not \U$67129 ( \67103 , \67102 );
buf \U$67130 ( \67104 , \1927 );
not \U$67131 ( \67105 , \67104 );
or \U$67132 ( \67106 , \67103 , \67105 );
buf \U$67133 ( \67107 , \714 );
xor \U$67134 ( \67108 , RIc0da0a8_91, RIc0d8c08_47);
buf \U$67135 ( \67109 , \67108 );
nand \U$67136 ( \67110 , \67107 , \67109 );
buf \U$67137 ( \67111 , \67110 );
buf \U$67138 ( \67112 , \67111 );
nand \U$67139 ( \67113 , \67106 , \67112 );
buf \U$67140 ( \67114 , \67113 );
buf \U$67141 ( \67115 , \67114 );
buf \U$67142 ( \67116 , \66118 );
not \U$67143 ( \67117 , \67116 );
buf \U$67144 ( \67118 , \16358 );
not \U$67145 ( \67119 , \67118 );
or \U$67146 ( \67120 , \67117 , \67119 );
buf \U$67147 ( \67121 , \734 );
buf \U$67148 ( \67122 , RIc0d8938_41);
buf \U$67149 ( \67123 , RIc0da378_97);
xor \U$67150 ( \67124 , \67122 , \67123 );
buf \U$67151 ( \67125 , \67124 );
buf \U$67152 ( \67126 , \67125 );
nand \U$67153 ( \67127 , \67121 , \67126 );
buf \U$67154 ( \67128 , \67127 );
buf \U$67155 ( \67129 , \67128 );
nand \U$67156 ( \67130 , \67120 , \67129 );
buf \U$67157 ( \67131 , \67130 );
buf \U$67158 ( \67132 , \67131 );
xor \U$67159 ( \67133 , \67115 , \67132 );
buf \U$67160 ( \67134 , \66409 );
not \U$67161 ( \67135 , \67134 );
buf \U$67162 ( \67136 , \13042 );
not \U$67163 ( \67137 , \67136 );
or \U$67164 ( \67138 , \67135 , \67137 );
buf \U$67165 ( \67139 , RIc0d8668_35);
buf \U$67166 ( \67140 , RIc0da648_103);
xnor \U$67167 ( \67141 , \67139 , \67140 );
buf \U$67168 ( \67142 , \67141 );
buf \U$67169 ( \67143 , \67142 );
not \U$67170 ( \67144 , \67143 );
buf \U$67171 ( \67145 , \16584 );
nand \U$67172 ( \67146 , \67144 , \67145 );
buf \U$67173 ( \67147 , \67146 );
buf \U$67174 ( \67148 , \67147 );
nand \U$67175 ( \67149 , \67138 , \67148 );
buf \U$67176 ( \67150 , \67149 );
buf \U$67177 ( \67151 , \67150 );
xor \U$67178 ( \67152 , \67133 , \67151 );
buf \U$67179 ( \67153 , \67152 );
buf \U$67180 ( \67154 , \67153 );
xor \U$67181 ( \67155 , \67101 , \67154 );
buf \U$67182 ( \67156 , \67155 );
buf \U$67183 ( \67157 , \67156 );
not \U$67184 ( \67158 , \67157 );
buf \U$67185 ( \67159 , \66462 );
not \U$67186 ( \67160 , \67159 );
buf \U$67187 ( \67161 , \15420 );
not \U$67188 ( \67162 , \67161 );
or \U$67189 ( \67163 , \67160 , \67162 );
buf \U$67190 ( \67164 , \12975 );
xor \U$67191 ( \67165 , RIc0daeb8_121, RIc0d7df8_17);
buf \U$67192 ( \67166 , \67165 );
nand \U$67193 ( \67167 , \67164 , \67166 );
buf \U$67194 ( \67168 , \67167 );
buf \U$67195 ( \67169 , \67168 );
nand \U$67196 ( \67170 , \67163 , \67169 );
buf \U$67197 ( \67171 , \67170 );
buf \U$67198 ( \67172 , \67171 );
buf \U$67199 ( \67173 , \66030 );
not \U$67200 ( \67174 , \67173 );
buf \U$67201 ( \67175 , \1389 );
not \U$67202 ( \67176 , \67175 );
or \U$67203 ( \67177 , \67174 , \67176 );
buf \U$67204 ( \67178 , \1401 );
buf \U$67205 ( \67179 , RIc0d8ed8_53);
buf \U$67206 ( \67180 , RIc0d9dd8_85);
xor \U$67207 ( \67181 , \67179 , \67180 );
buf \U$67208 ( \67182 , \67181 );
buf \U$67209 ( \67183 , \67182 );
nand \U$67210 ( \67184 , \67178 , \67183 );
buf \U$67211 ( \67185 , \67184 );
buf \U$67212 ( \67186 , \67185 );
nand \U$67213 ( \67187 , \67177 , \67186 );
buf \U$67214 ( \67188 , \67187 );
buf \U$67215 ( \67189 , \67188 );
xor \U$67216 ( \67190 , \67172 , \67189 );
buf \U$67217 ( \67191 , \66136 );
not \U$67218 ( \67192 , \67191 );
buf \U$67219 ( \67193 , \14982 );
not \U$67220 ( \67194 , \67193 );
or \U$67221 ( \67195 , \67192 , \67194 );
buf \U$67222 ( \67196 , RIc0dafa8_123);
buf \U$67223 ( \67197 , RIc0d7d08_15);
xnor \U$67224 ( \67198 , \67196 , \67197 );
buf \U$67225 ( \67199 , \67198 );
buf \U$67226 ( \67200 , \67199 );
not \U$67227 ( \67201 , \67200 );
buf \U$67228 ( \67202 , \14278 );
nand \U$67229 ( \67203 , \67201 , \67202 );
buf \U$67230 ( \67204 , \67203 );
buf \U$67231 ( \67205 , \67204 );
nand \U$67232 ( \67206 , \67195 , \67205 );
buf \U$67233 ( \67207 , \67206 );
buf \U$67234 ( \67208 , \67207 );
xor \U$67235 ( \67209 , \67190 , \67208 );
buf \U$67236 ( \67210 , \67209 );
buf \U$67237 ( \67211 , \67210 );
not \U$67238 ( \67212 , \67211 );
buf \U$67239 ( \67213 , \67212 );
buf \U$67240 ( \67214 , \67213 );
not \U$67241 ( \67215 , \67214 );
buf \U$67242 ( \67216 , \66291 );
not \U$67243 ( \67217 , \67216 );
buf \U$67244 ( \67218 , \22350 );
not \U$67245 ( \67219 , \67218 );
or \U$67246 ( \67220 , \67217 , \67219 );
buf \U$67247 ( \67221 , \16559 );
buf \U$67248 ( \67222 , RIc0d7fd8_21);
buf \U$67249 ( \67223 , RIc0dacd8_117);
xor \U$67250 ( \67224 , \67222 , \67223 );
buf \U$67251 ( \67225 , \67224 );
buf \U$67252 ( \67226 , \67225 );
nand \U$67253 ( \67227 , \67221 , \67226 );
buf \U$67254 ( \67228 , \67227 );
buf \U$67255 ( \67229 , \67228 );
nand \U$67256 ( \67230 , \67220 , \67229 );
buf \U$67257 ( \67231 , \67230 );
buf \U$67258 ( \67232 , \66239 );
not \U$67259 ( \67233 , \67232 );
buf \U$67260 ( \67234 , \15789 );
not \U$67261 ( \67235 , \67234 );
or \U$67262 ( \67236 , \67233 , \67235 );
buf \U$67263 ( \67237 , \15793 );
buf \U$67264 ( \67238 , RIc0d7c18_13);
buf \U$67265 ( \67239 , RIc0db098_125);
xor \U$67266 ( \67240 , \67238 , \67239 );
buf \U$67267 ( \67241 , \67240 );
buf \U$67268 ( \67242 , \67241 );
nand \U$67269 ( \67243 , \67237 , \67242 );
buf \U$67270 ( \67244 , \67243 );
buf \U$67271 ( \67245 , \67244 );
nand \U$67272 ( \67246 , \67236 , \67245 );
buf \U$67273 ( \67247 , \67246 );
buf \U$67274 ( \67248 , \67247 );
not \U$67275 ( \67249 , \67248 );
buf \U$67276 ( \67250 , \67249 );
xor \U$67277 ( \67251 , \67231 , \67250 );
buf \U$67278 ( \67252 , \66377 );
not \U$67279 ( \67253 , \67252 );
buf \U$67280 ( \67254 , \18150 );
not \U$67281 ( \67255 , \67254 );
or \U$67282 ( \67256 , \67253 , \67255 );
buf \U$67283 ( \67257 , \846 );
xor \U$67284 ( \67258 , RIc0d9fb8_89, RIc0d8cf8_49);
buf \U$67285 ( \67259 , \67258 );
nand \U$67286 ( \67260 , \67257 , \67259 );
buf \U$67287 ( \67261 , \67260 );
buf \U$67288 ( \67262 , \67261 );
nand \U$67289 ( \67263 , \67256 , \67262 );
buf \U$67290 ( \67264 , \67263 );
xor \U$67291 ( \67265 , \67251 , \67264 );
buf \U$67292 ( \67266 , \67265 );
not \U$67293 ( \67267 , \67266 );
buf \U$67294 ( \67268 , \67267 );
buf \U$67295 ( \67269 , \67268 );
not \U$67296 ( \67270 , \67269 );
or \U$67297 ( \67271 , \67215 , \67270 );
buf \U$67298 ( \67272 , \67265 );
buf \U$67299 ( \67273 , \67210 );
nand \U$67300 ( \67274 , \67272 , \67273 );
buf \U$67301 ( \67275 , \67274 );
buf \U$67302 ( \67276 , \67275 );
nand \U$67303 ( \67277 , \67271 , \67276 );
buf \U$67304 ( \67278 , \67277 );
buf \U$67305 ( \67279 , \67278 );
buf \U$67306 ( \67280 , \66174 );
not \U$67307 ( \67281 , \67280 );
buf \U$67308 ( \67282 , \1736 );
not \U$67309 ( \67283 , \67282 );
or \U$67310 ( \67284 , \67281 , \67283 );
buf \U$67311 ( \67285 , \584 );
buf \U$67312 ( \67286 , RIc0d8fc8_55);
buf \U$67313 ( \67287 , RIc0d9ce8_83);
xor \U$67314 ( \67288 , \67286 , \67287 );
buf \U$67315 ( \67289 , \67288 );
buf \U$67316 ( \67290 , \67289 );
nand \U$67317 ( \67291 , \67285 , \67290 );
buf \U$67318 ( \67292 , \67291 );
buf \U$67319 ( \67293 , \67292 );
nand \U$67320 ( \67294 , \67284 , \67293 );
buf \U$67321 ( \67295 , \67294 );
buf \U$67322 ( \67296 , \66101 );
not \U$67323 ( \67297 , \67296 );
buf \U$67324 ( \67298 , \12529 );
not \U$67325 ( \67299 , \67298 );
or \U$67326 ( \67300 , \67297 , \67299 );
buf \U$67327 ( \67301 , \14106 );
xor \U$67328 ( \67302 , RIc0daa08_111, RIc0d82a8_27);
buf \U$67329 ( \67303 , \67302 );
nand \U$67330 ( \67304 , \67301 , \67303 );
buf \U$67331 ( \67305 , \67304 );
buf \U$67332 ( \67306 , \67305 );
nand \U$67333 ( \67307 , \67300 , \67306 );
buf \U$67334 ( \67308 , \67307 );
xor \U$67335 ( \67309 , \67295 , \67308 );
buf \U$67336 ( \67310 , \66394 );
not \U$67337 ( \67311 , \67310 );
buf \U$67338 ( \67312 , \1765 );
not \U$67339 ( \67313 , \67312 );
or \U$67340 ( \67314 , \67311 , \67313 );
buf \U$67341 ( \67315 , \816 );
buf \U$67342 ( \67316 , RIc0d8de8_51);
buf \U$67343 ( \67317 , RIc0d9ec8_87);
xor \U$67344 ( \67318 , \67316 , \67317 );
buf \U$67345 ( \67319 , \67318 );
buf \U$67346 ( \67320 , \67319 );
nand \U$67347 ( \67321 , \67315 , \67320 );
buf \U$67348 ( \67322 , \67321 );
buf \U$67349 ( \67323 , \67322 );
nand \U$67350 ( \67324 , \67314 , \67323 );
buf \U$67351 ( \67325 , \67324 );
xnor \U$67352 ( \67326 , \67309 , \67325 );
buf \U$67353 ( \67327 , \67326 );
and \U$67354 ( \67328 , \67279 , \67327 );
not \U$67355 ( \67329 , \67279 );
buf \U$67356 ( \67330 , \67326 );
not \U$67357 ( \67331 , \67330 );
buf \U$67358 ( \67332 , \67331 );
buf \U$67359 ( \67333 , \67332 );
and \U$67360 ( \67334 , \67329 , \67333 );
nor \U$67361 ( \67335 , \67328 , \67334 );
buf \U$67362 ( \67336 , \67335 );
buf \U$67363 ( \67337 , \67336 );
not \U$67364 ( \67338 , \67337 );
or \U$67365 ( \67339 , \67158 , \67338 );
buf \U$67366 ( \67340 , \67156 );
buf \U$67367 ( \67341 , \67336 );
or \U$67368 ( \67342 , \67340 , \67341 );
nand \U$67369 ( \67343 , \67339 , \67342 );
buf \U$67370 ( \67344 , \67343 );
buf \U$67371 ( \67345 , \67344 );
buf \U$67372 ( \67346 , RIc0d9400_64);
buf \U$67373 ( \67347 , RIc0d9928_75);
xor \U$67374 ( \67348 , \67346 , \67347 );
buf \U$67375 ( \67349 , \67348 );
buf \U$67376 ( \67350 , \67349 );
not \U$67377 ( \67351 , \67350 );
buf \U$67378 ( \67352 , \2358 );
not \U$67379 ( \67353 , \67352 );
or \U$67380 ( \67354 , \67351 , \67353 );
buf \U$67381 ( \67355 , \13389 );
buf \U$67382 ( \67356 , RIc0d9388_63);
buf \U$67383 ( \67357 , RIc0d9928_75);
xor \U$67384 ( \67358 , \67356 , \67357 );
buf \U$67385 ( \67359 , \67358 );
buf \U$67386 ( \67360 , \67359 );
nand \U$67387 ( \67361 , \67355 , \67360 );
buf \U$67388 ( \67362 , \67361 );
buf \U$67389 ( \67363 , \67362 );
nand \U$67390 ( \67364 , \67354 , \67363 );
buf \U$67391 ( \67365 , \67364 );
buf \U$67392 ( \67366 , \67365 );
buf \U$67393 ( \67367 , \66357 );
not \U$67394 ( \67368 , \67367 );
buf \U$67395 ( \67369 , \22631 );
not \U$67396 ( \67370 , \67369 );
or \U$67397 ( \67371 , \67368 , \67370 );
buf \U$67398 ( \67372 , \26354 );
xor \U$67399 ( \67373 , RIc0da558_101, RIc0d8758_37);
buf \U$67400 ( \67374 , \67373 );
nand \U$67401 ( \67375 , \67372 , \67374 );
buf \U$67402 ( \67376 , \67375 );
buf \U$67403 ( \67377 , \67376 );
nand \U$67404 ( \67378 , \67371 , \67377 );
buf \U$67405 ( \67379 , \67378 );
buf \U$67406 ( \67380 , \67379 );
xor \U$67407 ( \67381 , \67366 , \67380 );
buf \U$67408 ( \67382 , \66209 );
not \U$67409 ( \67383 , \67382 );
buf \U$67410 ( \67384 , \17595 );
not \U$67411 ( \67385 , \67384 );
or \U$67412 ( \67386 , \67383 , \67385 );
buf \U$67413 ( \67387 , \12342 );
buf \U$67414 ( \67388 , RIc0d8488_31);
buf \U$67415 ( \67389 , RIc0da828_107);
xor \U$67416 ( \67390 , \67388 , \67389 );
buf \U$67417 ( \67391 , \67390 );
buf \U$67418 ( \67392 , \67391 );
nand \U$67419 ( \67393 , \67387 , \67392 );
buf \U$67420 ( \67394 , \67393 );
buf \U$67421 ( \67395 , \67394 );
nand \U$67422 ( \67396 , \67386 , \67395 );
buf \U$67423 ( \67397 , \67396 );
buf \U$67424 ( \67398 , \67397 );
xor \U$67425 ( \67399 , \67381 , \67398 );
buf \U$67426 ( \67400 , \67399 );
buf \U$67427 ( \67401 , \67400 );
not \U$67428 ( \67402 , \67401 );
buf \U$67429 ( \67403 , \67402 );
buf \U$67430 ( \67404 , \67403 );
not \U$67431 ( \67405 , \67404 );
buf \U$67432 ( \67406 , \66049 );
not \U$67433 ( \67407 , \67406 );
buf \U$67434 ( \67408 , \330 );
not \U$67435 ( \67409 , \67408 );
or \U$67436 ( \67410 , \67407 , \67409 );
buf \U$67437 ( \67411 , \343 );
buf \U$67438 ( \67412 , RIc0da288_95);
buf \U$67439 ( \67413 , RIc0d8a28_43);
xor \U$67440 ( \67414 , \67412 , \67413 );
buf \U$67441 ( \67415 , \67414 );
buf \U$67442 ( \67416 , \67415 );
nand \U$67443 ( \67417 , \67411 , \67416 );
buf \U$67444 ( \67418 , \67417 );
buf \U$67445 ( \67419 , \67418 );
nand \U$67446 ( \67420 , \67410 , \67419 );
buf \U$67447 ( \67421 , \67420 );
buf \U$67448 ( \67422 , \67421 );
not \U$67449 ( \67423 , \67422 );
buf \U$67450 ( \67424 , \66066 );
not \U$67451 ( \67425 , \67424 );
buf \U$67452 ( \67426 , \13949 );
not \U$67453 ( \67427 , \67426 );
or \U$67454 ( \67428 , \67425 , \67427 );
buf \U$67455 ( \67429 , \13953 );
buf \U$67456 ( \67430 , RIc0d7ee8_19);
buf \U$67457 ( \67431 , RIc0dadc8_119);
xor \U$67458 ( \67432 , \67430 , \67431 );
buf \U$67459 ( \67433 , \67432 );
buf \U$67460 ( \67434 , \67433 );
nand \U$67461 ( \67435 , \67429 , \67434 );
buf \U$67462 ( \67436 , \67435 );
buf \U$67463 ( \67437 , \67436 );
nand \U$67464 ( \67438 , \67428 , \67437 );
buf \U$67465 ( \67439 , \67438 );
buf \U$67466 ( \67440 , \67439 );
not \U$67467 ( \67441 , \67440 );
buf \U$67468 ( \67442 , \67441 );
buf \U$67469 ( \67443 , \67442 );
not \U$67470 ( \67444 , \67443 );
or \U$67471 ( \67445 , \67423 , \67444 );
buf \U$67472 ( \67446 , \67421 );
not \U$67473 ( \67447 , \67446 );
buf \U$67474 ( \67448 , \67439 );
nand \U$67475 ( \67449 , \67447 , \67448 );
buf \U$67476 ( \67450 , \67449 );
buf \U$67477 ( \67451 , \67450 );
nand \U$67478 ( \67452 , \67445 , \67451 );
buf \U$67479 ( \67453 , \67452 );
buf \U$67480 ( \67454 , \67453 );
buf \U$67481 ( \67455 , \66192 );
not \U$67482 ( \67456 , \67455 );
buf \U$67483 ( \67457 , \21959 );
not \U$67484 ( \67458 , \67457 );
or \U$67485 ( \67459 , \67456 , \67458 );
buf \U$67486 ( \67460 , \15909 );
buf \U$67487 ( \67461 , RIc0d8398_29);
buf \U$67488 ( \67462 , RIc0da918_109);
xor \U$67489 ( \67463 , \67461 , \67462 );
buf \U$67490 ( \67464 , \67463 );
buf \U$67491 ( \67465 , \67464 );
nand \U$67492 ( \67466 , \67460 , \67465 );
buf \U$67493 ( \67467 , \67466 );
buf \U$67494 ( \67468 , \67467 );
nand \U$67495 ( \67469 , \67459 , \67468 );
buf \U$67496 ( \67470 , \67469 );
buf \U$67497 ( \67471 , \67470 );
not \U$67498 ( \67472 , \67471 );
buf \U$67499 ( \67473 , \67472 );
buf \U$67500 ( \67474 , \67473 );
and \U$67501 ( \67475 , \67454 , \67474 );
not \U$67502 ( \67476 , \67454 );
buf \U$67503 ( \67477 , \67470 );
and \U$67504 ( \67478 , \67476 , \67477 );
nor \U$67505 ( \67479 , \67475 , \67478 );
buf \U$67506 ( \67480 , \67479 );
buf \U$67507 ( \67481 , \67480 );
not \U$67508 ( \67482 , \67481 );
buf \U$67509 ( \67483 , \67482 );
buf \U$67510 ( \67484 , \67483 );
not \U$67511 ( \67485 , \67484 );
or \U$67512 ( \67486 , \67405 , \67485 );
buf \U$67513 ( \67487 , \67480 );
buf \U$67514 ( \67488 , \67400 );
nand \U$67515 ( \67489 , \67487 , \67488 );
buf \U$67516 ( \67490 , \67489 );
buf \U$67517 ( \67491 , \67490 );
nand \U$67518 ( \67492 , \67486 , \67491 );
buf \U$67519 ( \67493 , \67492 );
buf \U$67520 ( \67494 , \67493 );
buf \U$67521 ( \67495 , \66157 );
not \U$67522 ( \67496 , \67495 );
buf \U$67523 ( \67497 , \1183 );
not \U$67524 ( \67498 , \67497 );
or \U$67525 ( \67499 , \67496 , \67498 );
buf \U$67526 ( \67500 , \3742 );
xor \U$67527 ( \67501 , RIc0d9a18_77, RIc0d9298_61);
buf \U$67528 ( \67502 , \67501 );
nand \U$67529 ( \67503 , \67500 , \67502 );
buf \U$67530 ( \67504 , \67503 );
buf \U$67531 ( \67505 , \67504 );
nand \U$67532 ( \67506 , \67499 , \67505 );
buf \U$67533 ( \67507 , \67506 );
buf \U$67534 ( \67508 , RIc0d9400_64);
buf \U$67535 ( \67509 , RIc0d99a0_76);
nand \U$67536 ( \67510 , \67508 , \67509 );
buf \U$67537 ( \67511 , \67510 );
buf \U$67538 ( \67512 , RIc0d9400_64);
buf \U$67539 ( \67513 , RIc0d99a0_76);
or \U$67540 ( \67514 , \67512 , \67513 );
buf \U$67541 ( \67515 , RIc0d9a18_77);
nand \U$67542 ( \67516 , \67514 , \67515 );
buf \U$67543 ( \67517 , \67516 );
nand \U$67544 ( \67518 , \67511 , RIc0d9928_75, \67517 );
xor \U$67545 ( \67519 , \67507 , \67518 );
buf \U$67546 ( \67520 , \67519 );
not \U$67547 ( \67521 , \67520 );
buf \U$67548 ( \67522 , \66012 );
not \U$67549 ( \67523 , \67522 );
buf \U$67550 ( \67524 , \21461 );
not \U$67551 ( \67525 , \67524 );
or \U$67552 ( \67526 , \67523 , \67525 );
buf \U$67553 ( \67527 , \22006 );
xor \U$67554 ( \67528 , RIc0da468_99, RIc0d8848_39);
buf \U$67555 ( \67529 , \67528 );
nand \U$67556 ( \67530 , \67527 , \67529 );
buf \U$67557 ( \67531 , \67530 );
buf \U$67558 ( \67532 , \67531 );
nand \U$67559 ( \67533 , \67526 , \67532 );
buf \U$67560 ( \67534 , \67533 );
buf \U$67561 ( \67535 , \67534 );
buf \U$67562 ( \67536 , \66225 );
not \U$67563 ( \67537 , \67536 );
buf \U$67564 ( \67538 , \26466 );
not \U$67565 ( \67539 , \67538 );
or \U$67566 ( \67540 , \67537 , \67539 );
buf \U$67567 ( \67541 , \12303 );
buf \U$67568 ( \67542 , RIc0dabe8_115);
buf \U$67569 ( \67543 , RIc0d80c8_23);
xor \U$67570 ( \67544 , \67542 , \67543 );
buf \U$67571 ( \67545 , \67544 );
buf \U$67572 ( \67546 , \67545 );
nand \U$67573 ( \67547 , \67541 , \67546 );
buf \U$67574 ( \67548 , \67547 );
buf \U$67575 ( \67549 , \67548 );
nand \U$67576 ( \67550 , \67540 , \67549 );
buf \U$67577 ( \67551 , \67550 );
buf \U$67578 ( \67552 , \67551 );
xor \U$67579 ( \67553 , \67535 , \67552 );
buf \U$67580 ( \67554 , \67553 );
buf \U$67581 ( \67555 , \67554 );
not \U$67582 ( \67556 , \67555 );
or \U$67583 ( \67557 , \67521 , \67556 );
buf \U$67584 ( \67558 , \67519 );
buf \U$67585 ( \67559 , \67554 );
or \U$67586 ( \67560 , \67558 , \67559 );
nand \U$67587 ( \67561 , \67557 , \67560 );
buf \U$67588 ( \67562 , \67561 );
buf \U$67589 ( \67563 , \67562 );
xor \U$67590 ( \67564 , \67494 , \67563 );
buf \U$67591 ( \67565 , \67564 );
buf \U$67592 ( \67566 , \67565 );
xor \U$67593 ( \67567 , \67345 , \67566 );
buf \U$67594 ( \67568 , \67567 );
buf \U$67595 ( \67569 , \67568 );
xor \U$67596 ( \67570 , \66998 , \67569 );
xor \U$67597 ( \67571 , \64295 , \64301 );
and \U$67598 ( \67572 , \67571 , \64341 );
and \U$67599 ( \67573 , \64295 , \64301 );
or \U$67600 ( \67574 , \67572 , \67573 );
buf \U$67601 ( \67575 , \67574 );
buf \U$67602 ( \67576 , \67575 );
xor \U$67603 ( \67577 , \67570 , \67576 );
buf \U$67604 ( \67578 , \67577 );
buf \U$67605 ( \67579 , \67578 );
xor \U$67606 ( \67580 , \66992 , \67579 );
xor \U$67607 ( \67581 , \64289 , \64344 );
and \U$67608 ( \67582 , \67581 , \64963 );
and \U$67609 ( \67583 , \64289 , \64344 );
or \U$67610 ( \67584 , \67582 , \67583 );
buf \U$67611 ( \67585 , \67584 );
buf \U$67612 ( \67586 , \67585 );
xor \U$67613 ( \67587 , \67580 , \67586 );
buf \U$67614 ( \67588 , \67587 );
buf \U$67615 ( \67589 , \67588 );
xor \U$67616 ( \67590 , \66986 , \67589 );
buf \U$67617 ( \67591 , \67590 );
buf \U$67618 ( \67592 , \67591 );
not \U$67619 ( \67593 , \67592 );
buf \U$67620 ( \67594 , \67593 );
buf \U$67621 ( \67595 , \67594 );
nand \U$67622 ( \67596 , \66739 , \67595 );
buf \U$67623 ( \67597 , \67596 );
buf \U$67624 ( \67598 , \67597 );
xor \U$67625 ( \67599 , \64966 , \65922 );
xor \U$67626 ( \67600 , \67599 , \66733 );
buf \U$67627 ( \67601 , \67600 );
buf \U$67628 ( \67602 , \67601 );
xor \U$67629 ( \67603 , \65667 , \65673 );
xor \U$67630 ( \67604 , \67603 , \65689 );
buf \U$67631 ( \67605 , \67604 );
buf \U$67632 ( \67606 , \67605 );
buf \U$67633 ( \67607 , \65041 );
not \U$67634 ( \67608 , \67607 );
buf \U$67635 ( \67609 , \67608 );
buf \U$67636 ( \67610 , \67609 );
not \U$67637 ( \67611 , \67610 );
xor \U$67638 ( \67612 , \65026 , \65048 );
buf \U$67639 ( \67613 , \67612 );
not \U$67640 ( \67614 , \67613 );
or \U$67641 ( \67615 , \67611 , \67614 );
buf \U$67642 ( \67616 , \67612 );
buf \U$67643 ( \67617 , \67609 );
or \U$67644 ( \67618 , \67616 , \67617 );
nand \U$67645 ( \67619 , \67615 , \67618 );
buf \U$67646 ( \67620 , \67619 );
buf \U$67647 ( \67621 , \67620 );
xor \U$67648 ( \67622 , \67606 , \67621 );
and \U$67649 ( \67623 , \65408 , \65403 );
not \U$67650 ( \67624 , \65408 );
and \U$67651 ( \67625 , \67624 , \65415 );
or \U$67652 ( \67626 , \67623 , \67625 );
buf \U$67653 ( \67627 , \67626 );
buf \U$67654 ( \67628 , \65419 );
and \U$67655 ( \67629 , \67627 , \67628 );
not \U$67656 ( \67630 , \67627 );
buf \U$67657 ( \67631 , \65399 );
and \U$67658 ( \67632 , \67630 , \67631 );
nor \U$67659 ( \67633 , \67629 , \67632 );
buf \U$67660 ( \67634 , \67633 );
buf \U$67661 ( \67635 , \67634 );
and \U$67662 ( \67636 , \67622 , \67635 );
and \U$67663 ( \67637 , \67606 , \67621 );
or \U$67664 ( \67638 , \67636 , \67637 );
buf \U$67665 ( \67639 , \67638 );
buf \U$67666 ( \67640 , \67639 );
xor \U$67667 ( \67641 , \55327 , \55408 );
and \U$67668 ( \67642 , \67641 , \55415 );
and \U$67669 ( \67643 , \55327 , \55408 );
or \U$67670 ( \67644 , \67642 , \67643 );
buf \U$67671 ( \67645 , \67644 );
buf \U$67672 ( \67646 , \67645 );
not \U$67673 ( \67647 , \67646 );
buf \U$67674 ( \67648 , \65461 );
not \U$67675 ( \67649 , \67648 );
buf \U$67676 ( \67650 , \65512 );
not \U$67677 ( \67651 , \67650 );
or \U$67678 ( \67652 , \67649 , \67651 );
buf \U$67679 ( \67653 , \65509 );
buf \U$67680 ( \67654 , \65464 );
nand \U$67681 ( \67655 , \67653 , \67654 );
buf \U$67682 ( \67656 , \67655 );
buf \U$67683 ( \67657 , \67656 );
nand \U$67684 ( \67658 , \67652 , \67657 );
buf \U$67685 ( \67659 , \67658 );
buf \U$67686 ( \67660 , \67659 );
buf \U$67687 ( \67661 , \65522 );
xnor \U$67688 ( \67662 , \67660 , \67661 );
buf \U$67689 ( \67663 , \67662 );
buf \U$67690 ( \67664 , \67663 );
not \U$67691 ( \67665 , \67664 );
buf \U$67692 ( \67666 , \67665 );
buf \U$67693 ( \67667 , \67666 );
not \U$67694 ( \67668 , \67667 );
or \U$67695 ( \67669 , \67647 , \67668 );
not \U$67696 ( \67670 , \67663 );
buf \U$67697 ( \67671 , \67645 );
not \U$67698 ( \67672 , \67671 );
buf \U$67699 ( \67673 , \67672 );
not \U$67700 ( \67674 , \67673 );
or \U$67701 ( \67675 , \67670 , \67674 );
xor \U$67702 ( \67676 , \65876 , \65883 );
xor \U$67703 ( \67677 , \67676 , \65887 );
buf \U$67704 ( \67678 , \67677 );
nand \U$67705 ( \67679 , \67675 , \67678 );
buf \U$67706 ( \67680 , \67679 );
nand \U$67707 ( \67681 , \67669 , \67680 );
buf \U$67708 ( \67682 , \67681 );
buf \U$67709 ( \67683 , \67682 );
xor \U$67710 ( \67684 , \67640 , \67683 );
xor \U$67711 ( \67685 , \65861 , \65892 );
xor \U$67712 ( \67686 , \67685 , \65904 );
buf \U$67713 ( \67687 , \67686 );
buf \U$67714 ( \67688 , \67687 );
and \U$67715 ( \67689 , \67684 , \67688 );
and \U$67716 ( \67690 , \67640 , \67683 );
or \U$67717 ( \67691 , \67689 , \67690 );
buf \U$67718 ( \67692 , \67691 );
buf \U$67719 ( \67693 , \67692 );
xor \U$67720 ( \67694 , \66627 , \66715 );
xor \U$67721 ( \67695 , \67694 , \66720 );
buf \U$67722 ( \67696 , \67695 );
buf \U$67723 ( \67697 , \67696 );
xor \U$67724 ( \67698 , \67693 , \67697 );
xor \U$67725 ( \67699 , \66639 , \66643 );
xor \U$67726 ( \67700 , \67699 , \66710 );
buf \U$67727 ( \67701 , \67700 );
buf \U$67728 ( \67702 , \67701 );
buf \U$67729 ( \67703 , \66658 );
not \U$67730 ( \67704 , \67703 );
buf \U$67731 ( \67705 , \66680 );
not \U$67732 ( \67706 , \67705 );
or \U$67733 ( \67707 , \67704 , \67706 );
buf \U$67734 ( \67708 , \66658 );
buf \U$67735 ( \67709 , \66680 );
or \U$67736 ( \67710 , \67708 , \67709 );
nand \U$67737 ( \67711 , \67707 , \67710 );
buf \U$67738 ( \67712 , \67711 );
buf \U$67739 ( \67713 , \67712 );
buf \U$67740 ( \67714 , \66703 );
not \U$67741 ( \67715 , \67714 );
buf \U$67742 ( \67716 , \67715 );
buf \U$67743 ( \67717 , \67716 );
and \U$67744 ( \67718 , \67713 , \67717 );
not \U$67745 ( \67719 , \67713 );
buf \U$67746 ( \67720 , \66703 );
and \U$67747 ( \67721 , \67719 , \67720 );
nor \U$67748 ( \67722 , \67718 , \67721 );
buf \U$67749 ( \67723 , \67722 );
buf \U$67750 ( \67724 , \67723 );
not \U$67751 ( \67725 , \67724 );
buf \U$67752 ( \67726 , \67725 );
buf \U$67753 ( \67727 , \67726 );
not \U$67754 ( \67728 , \67727 );
not \U$67755 ( \67729 , \55982 );
not \U$67756 ( \67730 , \55948 );
or \U$67757 ( \67731 , \67729 , \67730 );
not \U$67758 ( \67732 , \55945 );
not \U$67759 ( \67733 , \55981 );
or \U$67760 ( \67734 , \67732 , \67733 );
nand \U$67761 ( \67735 , \67734 , \55914 );
nand \U$67762 ( \67736 , \67731 , \67735 );
buf \U$67763 ( \67737 , \67736 );
not \U$67764 ( \67738 , \67737 );
or \U$67765 ( \67739 , \67728 , \67738 );
buf \U$67766 ( \67740 , \67736 );
buf \U$67767 ( \67741 , \67726 );
or \U$67768 ( \67742 , \67740 , \67741 );
buf \U$67769 ( \67743 , \55888 );
not \U$67770 ( \67744 , \67743 );
buf \U$67771 ( \67745 , \55871 );
not \U$67772 ( \67746 , \67745 );
or \U$67773 ( \67747 , \67744 , \67746 );
buf \U$67774 ( \67748 , \55891 );
not \U$67775 ( \67749 , \67748 );
buf \U$67776 ( \67750 , \55868 );
not \U$67777 ( \67751 , \67750 );
or \U$67778 ( \67752 , \67749 , \67751 );
buf \U$67779 ( \67753 , \55881 );
nand \U$67780 ( \67754 , \67752 , \67753 );
buf \U$67781 ( \67755 , \67754 );
buf \U$67782 ( \67756 , \67755 );
nand \U$67783 ( \67757 , \67747 , \67756 );
buf \U$67784 ( \67758 , \67757 );
buf \U$67785 ( \67759 , \67758 );
nand \U$67786 ( \67760 , \67742 , \67759 );
buf \U$67787 ( \67761 , \67760 );
buf \U$67788 ( \67762 , \67761 );
nand \U$67789 ( \67763 , \67739 , \67762 );
buf \U$67790 ( \67764 , \67763 );
buf \U$67791 ( \67765 , \67764 );
xor \U$67792 ( \67766 , \67702 , \67765 );
xor \U$67793 ( \67767 , \65609 , \65701 );
xor \U$67794 ( \67768 , \67767 , \65726 );
buf \U$67795 ( \67769 , \67768 );
buf \U$67796 ( \67770 , \67769 );
and \U$67797 ( \67771 , \67766 , \67770 );
and \U$67798 ( \67772 , \67702 , \67765 );
or \U$67799 ( \67773 , \67771 , \67772 );
buf \U$67800 ( \67774 , \67773 );
buf \U$67801 ( \67775 , \67774 );
and \U$67802 ( \67776 , \67698 , \67775 );
and \U$67803 ( \67777 , \67693 , \67697 );
or \U$67804 ( \67778 , \67776 , \67777 );
buf \U$67805 ( \67779 , \67778 );
not \U$67806 ( \67780 , \67779 );
xor \U$67807 ( \67781 , \66598 , \66604 );
xor \U$67808 ( \67782 , \67781 , \66725 );
buf \U$67809 ( \67783 , \67782 );
not \U$67810 ( \67784 , \67783 );
or \U$67811 ( \67785 , \67780 , \67784 );
buf \U$67812 ( \67786 , \67783 );
not \U$67813 ( \67787 , \67786 );
buf \U$67814 ( \67788 , \67787 );
not \U$67815 ( \67789 , \67788 );
buf \U$67816 ( \67790 , \67779 );
not \U$67817 ( \67791 , \67790 );
buf \U$67818 ( \67792 , \67791 );
not \U$67819 ( \67793 , \67792 );
or \U$67820 ( \67794 , \67789 , \67793 );
xor \U$67821 ( \67795 , \64973 , \65543 );
xor \U$67822 ( \67796 , \67795 , \65917 );
buf \U$67823 ( \67797 , \67796 );
nand \U$67824 ( \67798 , \67794 , \67797 );
nand \U$67825 ( \67799 , \67785 , \67798 );
buf \U$67826 ( \67800 , \67799 );
or \U$67827 ( \67801 , \67602 , \67800 );
buf \U$67828 ( \67802 , \67801 );
buf \U$67829 ( \67803 , \67802 );
and \U$67830 ( \67804 , \67598 , \67803 );
buf \U$67831 ( \67805 , \67804 );
buf \U$67832 ( \67806 , \67805 );
xor \U$67833 ( \67807 , \66828 , \66843 );
and \U$67834 ( \67808 , \67807 , \66850 );
and \U$67835 ( \67809 , \66828 , \66843 );
or \U$67836 ( \67810 , \67808 , \67809 );
buf \U$67837 ( \67811 , \67810 );
buf \U$67838 ( \67812 , \67811 );
xor \U$67839 ( \67813 , \66917 , \66923 );
and \U$67840 ( \67814 , \67813 , \66930 );
and \U$67841 ( \67815 , \66917 , \66923 );
or \U$67842 ( \67816 , \67814 , \67815 );
buf \U$67843 ( \67817 , \67816 );
buf \U$67844 ( \67818 , \67817 );
xor \U$67845 ( \67819 , \67812 , \67818 );
xor \U$67846 ( \67820 , \66951 , \66957 );
and \U$67847 ( \67821 , \67820 , \66964 );
and \U$67848 ( \67822 , \66951 , \66957 );
or \U$67849 ( \67823 , \67821 , \67822 );
buf \U$67850 ( \67824 , \67823 );
buf \U$67851 ( \67825 , \67824 );
xor \U$67852 ( \67826 , \67819 , \67825 );
buf \U$67853 ( \67827 , \67826 );
buf \U$67854 ( \67828 , \67827 );
buf \U$67855 ( \67829 , \67156 );
buf \U$67856 ( \67830 , \67565 );
or \U$67857 ( \67831 , \67829 , \67830 );
buf \U$67858 ( \67832 , \67336 );
not \U$67859 ( \67833 , \67832 );
buf \U$67860 ( \67834 , \67833 );
buf \U$67861 ( \67835 , \67834 );
nand \U$67862 ( \67836 , \67831 , \67835 );
buf \U$67863 ( \67837 , \67836 );
buf \U$67864 ( \67838 , \67837 );
buf \U$67865 ( \67839 , \67565 );
buf \U$67866 ( \67840 , \67156 );
nand \U$67867 ( \67841 , \67839 , \67840 );
buf \U$67868 ( \67842 , \67841 );
buf \U$67869 ( \67843 , \67842 );
nand \U$67870 ( \67844 , \67838 , \67843 );
buf \U$67871 ( \67845 , \67844 );
buf \U$67872 ( \67846 , \67845 );
xor \U$67873 ( \67847 , \67828 , \67846 );
buf \U$67874 ( \67848 , \67065 );
not \U$67875 ( \67849 , \67848 );
buf \U$67876 ( \67850 , \67081 );
not \U$67877 ( \67851 , \67850 );
or \U$67878 ( \67852 , \67849 , \67851 );
buf \U$67879 ( \67853 , \67081 );
buf \U$67880 ( \67854 , \67065 );
or \U$67881 ( \67855 , \67853 , \67854 );
buf \U$67882 ( \67856 , \67098 );
nand \U$67883 ( \67857 , \67855 , \67856 );
buf \U$67884 ( \67858 , \67857 );
buf \U$67885 ( \67859 , \67858 );
nand \U$67886 ( \67860 , \67852 , \67859 );
buf \U$67887 ( \67861 , \67860 );
buf \U$67888 ( \67862 , \67861 );
xor \U$67889 ( \67863 , \67016 , \67030 );
and \U$67890 ( \67864 , \67863 , \67049 );
and \U$67891 ( \67865 , \67016 , \67030 );
or \U$67892 ( \67866 , \67864 , \67865 );
buf \U$67893 ( \67867 , \67866 );
buf \U$67894 ( \67868 , \67867 );
xor \U$67895 ( \67869 , \67862 , \67868 );
xor \U$67896 ( \67870 , \67366 , \67380 );
and \U$67897 ( \67871 , \67870 , \67398 );
and \U$67898 ( \67872 , \67366 , \67380 );
or \U$67899 ( \67873 , \67871 , \67872 );
buf \U$67900 ( \67874 , \67873 );
buf \U$67901 ( \67875 , \67874 );
xor \U$67902 ( \67876 , \67869 , \67875 );
buf \U$67903 ( \67877 , \67876 );
xor \U$67904 ( \67878 , \67172 , \67189 );
and \U$67905 ( \67879 , \67878 , \67208 );
and \U$67906 ( \67880 , \67172 , \67189 );
or \U$67907 ( \67881 , \67879 , \67880 );
buf \U$67908 ( \67882 , \67881 );
buf \U$67909 ( \67883 , \67882 );
xor \U$67910 ( \67884 , \67115 , \67132 );
and \U$67911 ( \67885 , \67884 , \67151 );
and \U$67912 ( \67886 , \67115 , \67132 );
or \U$67913 ( \67887 , \67885 , \67886 );
buf \U$67914 ( \67888 , \67887 );
buf \U$67915 ( \67889 , \67888 );
xor \U$67916 ( \67890 , \67883 , \67889 );
buf \U$67917 ( \67891 , \67325 );
not \U$67918 ( \67892 , \67891 );
buf \U$67919 ( \67893 , \67308 );
not \U$67920 ( \67894 , \67893 );
or \U$67921 ( \67895 , \67892 , \67894 );
buf \U$67922 ( \67896 , \67308 );
buf \U$67923 ( \67897 , \67325 );
or \U$67924 ( \67898 , \67896 , \67897 );
buf \U$67925 ( \67899 , \67295 );
nand \U$67926 ( \67900 , \67898 , \67899 );
buf \U$67927 ( \67901 , \67900 );
buf \U$67928 ( \67902 , \67901 );
nand \U$67929 ( \67903 , \67895 , \67902 );
buf \U$67930 ( \67904 , \67903 );
buf \U$67931 ( \67905 , \67904 );
xor \U$67932 ( \67906 , \67890 , \67905 );
buf \U$67933 ( \67907 , \67906 );
xor \U$67934 ( \67908 , \67877 , \67907 );
xor \U$67935 ( \67909 , \67052 , \67100 );
and \U$67936 ( \67910 , \67909 , \67154 );
and \U$67937 ( \67911 , \67052 , \67100 );
or \U$67938 ( \67912 , \67910 , \67911 );
buf \U$67939 ( \67913 , \67912 );
xor \U$67940 ( \67914 , \67908 , \67913 );
buf \U$67941 ( \67915 , \67914 );
and \U$67942 ( \67916 , \67847 , \67915 );
and \U$67943 ( \67917 , \67828 , \67846 );
or \U$67944 ( \67918 , \67916 , \67917 );
buf \U$67945 ( \67919 , \67918 );
buf \U$67946 ( \67920 , RIc0d8500_32);
buf \U$67947 ( \67921 , RIc0da738_105);
xnor \U$67948 ( \67922 , \67920 , \67921 );
buf \U$67949 ( \67923 , \67922 );
buf \U$67950 ( \67924 , \67923 );
not \U$67951 ( \67925 , \67924 );
buf \U$67952 ( \67926 , \67925 );
buf \U$67953 ( \67927 , \67926 );
not \U$67954 ( \67928 , \67927 );
buf \U$67955 ( \67929 , \25475 );
not \U$67956 ( \67930 , \67929 );
or \U$67957 ( \67931 , \67928 , \67930 );
buf \U$67958 ( \67932 , \12744 );
buf \U$67959 ( \67933 , RIc0d8488_31);
buf \U$67960 ( \67934 , RIc0da738_105);
xor \U$67961 ( \67935 , \67933 , \67934 );
buf \U$67962 ( \67936 , \67935 );
buf \U$67963 ( \67937 , \67936 );
nand \U$67964 ( \67938 , \67932 , \67937 );
buf \U$67965 ( \67939 , \67938 );
buf \U$67966 ( \67940 , \67939 );
nand \U$67967 ( \67941 , \67931 , \67940 );
buf \U$67968 ( \67942 , \67941 );
xor \U$67969 ( \67943 , RIc0da468_99, RIc0d87d0_38);
buf \U$67970 ( \67944 , \67943 );
not \U$67971 ( \67945 , \67944 );
buf \U$67972 ( \67946 , \19695 );
not \U$67973 ( \67947 , \67946 );
or \U$67974 ( \67948 , \67945 , \67947 );
buf \U$67975 ( \67949 , \12584 );
xor \U$67976 ( \67950 , RIc0da468_99, RIc0d8758_37);
buf \U$67977 ( \67951 , \67950 );
nand \U$67978 ( \67952 , \67949 , \67951 );
buf \U$67979 ( \67953 , \67952 );
buf \U$67980 ( \67954 , \67953 );
nand \U$67981 ( \67955 , \67948 , \67954 );
buf \U$67982 ( \67956 , \67955 );
xor \U$67983 ( \67957 , \67942 , \67956 );
buf \U$67984 ( \67958 , \67957 );
buf \U$67985 ( \67959 , RIc0d9400_64);
buf \U$67986 ( \67960 , RIc0d9838_73);
xor \U$67987 ( \67961 , \67959 , \67960 );
buf \U$67988 ( \67962 , \67961 );
buf \U$67989 ( \67963 , \67962 );
not \U$67990 ( \67964 , \67963 );
buf \U$67991 ( \67965 , \2871 );
not \U$67992 ( \67966 , \67965 );
or \U$67993 ( \67967 , \67964 , \67966 );
buf \U$67994 ( \67968 , \1856 );
buf \U$67995 ( \67969 , RIc0d9388_63);
buf \U$67996 ( \67970 , RIc0d9838_73);
xor \U$67997 ( \67971 , \67969 , \67970 );
buf \U$67998 ( \67972 , \67971 );
buf \U$67999 ( \67973 , \67972 );
nand \U$68000 ( \67974 , \67968 , \67973 );
buf \U$68001 ( \67975 , \67974 );
buf \U$68002 ( \67976 , \67975 );
nand \U$68003 ( \67977 , \67967 , \67976 );
buf \U$68004 ( \67978 , \67977 );
buf \U$68005 ( \67979 , \67978 );
xor \U$68006 ( \67980 , \67958 , \67979 );
buf \U$68007 ( \67981 , \67980 );
buf \U$68008 ( \67982 , \67981 );
buf \U$68009 ( \67983 , \67507 );
not \U$68010 ( \67984 , \67983 );
buf \U$68011 ( \67985 , \67518 );
nor \U$68012 ( \67986 , \67984 , \67985 );
buf \U$68013 ( \67987 , \67986 );
buf \U$68014 ( \67988 , \67987 );
buf \U$68015 ( \67989 , \67545 );
not \U$68016 ( \67990 , \67989 );
buf \U$68017 ( \67991 , \27743 );
not \U$68018 ( \67992 , \67991 );
or \U$68019 ( \67993 , \67990 , \67992 );
buf \U$68020 ( \67994 , \12303 );
buf \U$68021 ( \67995 , RIc0d8050_22);
buf \U$68022 ( \67996 , RIc0dabe8_115);
xor \U$68023 ( \67997 , \67995 , \67996 );
buf \U$68024 ( \67998 , \67997 );
buf \U$68025 ( \67999 , \67998 );
nand \U$68026 ( \68000 , \67994 , \67999 );
buf \U$68027 ( \68001 , \68000 );
buf \U$68028 ( \68002 , \68001 );
nand \U$68029 ( \68003 , \67993 , \68002 );
buf \U$68030 ( \68004 , \68003 );
buf \U$68031 ( \68005 , \68004 );
or \U$68032 ( \68006 , \67988 , \68005 );
buf \U$68033 ( \68007 , \68006 );
buf \U$68034 ( \68008 , \68007 );
not \U$68035 ( \68009 , \68008 );
buf \U$68036 ( \68010 , \67439 );
not \U$68037 ( \68011 , \68010 );
buf \U$68038 ( \68012 , \67421 );
not \U$68039 ( \68013 , \68012 );
or \U$68040 ( \68014 , \68011 , \68013 );
buf \U$68041 ( \68015 , \67439 );
buf \U$68042 ( \68016 , \67421 );
or \U$68043 ( \68017 , \68015 , \68016 );
buf \U$68044 ( \68018 , \67470 );
nand \U$68045 ( \68019 , \68017 , \68018 );
buf \U$68046 ( \68020 , \68019 );
buf \U$68047 ( \68021 , \68020 );
nand \U$68048 ( \68022 , \68014 , \68021 );
buf \U$68049 ( \68023 , \68022 );
buf \U$68050 ( \68024 , \68023 );
not \U$68051 ( \68025 , \68024 );
or \U$68052 ( \68026 , \68009 , \68025 );
buf \U$68053 ( \68027 , \67987 );
buf \U$68054 ( \68028 , \68004 );
nand \U$68055 ( \68029 , \68027 , \68028 );
buf \U$68056 ( \68030 , \68029 );
buf \U$68057 ( \68031 , \68030 );
nand \U$68058 ( \68032 , \68026 , \68031 );
buf \U$68059 ( \68033 , \68032 );
buf \U$68060 ( \68034 , \68033 );
xor \U$68061 ( \68035 , \67982 , \68034 );
xor \U$68062 ( \68036 , \67883 , \67889 );
and \U$68063 ( \68037 , \68036 , \67905 );
and \U$68064 ( \68038 , \67883 , \67889 );
or \U$68065 ( \68039 , \68037 , \68038 );
buf \U$68066 ( \68040 , \68039 );
buf \U$68067 ( \68041 , \68040 );
xnor \U$68068 ( \68042 , \68035 , \68041 );
buf \U$68069 ( \68043 , \68042 );
buf \U$68070 ( \68044 , \67907 );
not \U$68071 ( \68045 , \68044 );
buf \U$68072 ( \68046 , \67877 );
not \U$68073 ( \68047 , \68046 );
or \U$68074 ( \68048 , \68045 , \68047 );
buf \U$68075 ( \68049 , \67877 );
buf \U$68076 ( \68050 , \67907 );
or \U$68077 ( \68051 , \68049 , \68050 );
buf \U$68078 ( \68052 , \67913 );
nand \U$68079 ( \68053 , \68051 , \68052 );
buf \U$68080 ( \68054 , \68053 );
buf \U$68081 ( \68055 , \68054 );
nand \U$68082 ( \68056 , \68048 , \68055 );
buf \U$68083 ( \68057 , \68056 );
xor \U$68084 ( \68058 , \68043 , \68057 );
buf \U$68085 ( \68059 , \67289 );
not \U$68086 ( \68060 , \68059 );
buf \U$68087 ( \68061 , \12254 );
not \U$68088 ( \68062 , \68061 );
or \U$68089 ( \68063 , \68060 , \68062 );
buf \U$68090 ( \68064 , \993 );
buf \U$68091 ( \68065 , RIc0d8f50_54);
buf \U$68092 ( \68066 , RIc0d9ce8_83);
xor \U$68093 ( \68067 , \68065 , \68066 );
buf \U$68094 ( \68068 , \68067 );
buf \U$68095 ( \68069 , \68068 );
nand \U$68096 ( \68070 , \68064 , \68069 );
buf \U$68097 ( \68071 , \68070 );
buf \U$68098 ( \68072 , \68071 );
nand \U$68099 ( \68073 , \68063 , \68072 );
buf \U$68100 ( \68074 , \68073 );
buf \U$68101 ( \68075 , \68074 );
buf \U$68102 ( \68076 , \67302 );
not \U$68103 ( \68077 , \68076 );
buf \U$68104 ( \68078 , \14346 );
not \U$68105 ( \68079 , \68078 );
or \U$68106 ( \68080 , \68077 , \68079 );
buf \U$68107 ( \68081 , \25649 );
buf \U$68108 ( \68082 , RIc0d8230_26);
buf \U$68109 ( \68083 , RIc0daa08_111);
xor \U$68110 ( \68084 , \68082 , \68083 );
buf \U$68111 ( \68085 , \68084 );
buf \U$68112 ( \68086 , \68085 );
nand \U$68113 ( \68087 , \68081 , \68086 );
buf \U$68114 ( \68088 , \68087 );
buf \U$68115 ( \68089 , \68088 );
nand \U$68116 ( \68090 , \68080 , \68089 );
buf \U$68117 ( \68091 , \68090 );
buf \U$68118 ( \68092 , \68091 );
xor \U$68119 ( \68093 , \68075 , \68092 );
buf \U$68120 ( \68094 , \67125 );
not \U$68121 ( \68095 , \68094 );
buf \U$68122 ( \68096 , \13092 );
not \U$68123 ( \68097 , \68096 );
or \U$68124 ( \68098 , \68095 , \68097 );
buf \U$68125 ( \68099 , \734 );
buf \U$68126 ( \68100 , RIc0da378_97);
buf \U$68127 ( \68101 , RIc0d88c0_40);
xor \U$68128 ( \68102 , \68100 , \68101 );
buf \U$68129 ( \68103 , \68102 );
buf \U$68130 ( \68104 , \68103 );
nand \U$68131 ( \68105 , \68099 , \68104 );
buf \U$68132 ( \68106 , \68105 );
buf \U$68133 ( \68107 , \68106 );
nand \U$68134 ( \68108 , \68098 , \68107 );
buf \U$68135 ( \68109 , \68108 );
buf \U$68136 ( \68110 , \68109 );
xor \U$68137 ( \68111 , \68093 , \68110 );
buf \U$68138 ( \68112 , \68111 );
buf \U$68139 ( \68113 , \68112 );
buf \U$68140 ( \68114 , \1351 );
buf \U$68141 ( \68115 , \67059 );
and \U$68142 ( \68116 , \68114 , \68115 );
buf \U$68143 ( \68117 , \1026 );
buf \U$68144 ( \68118 , RIc0d9130_58);
buf \U$68145 ( \68119 , RIc0d9b08_79);
xor \U$68146 ( \68120 , \68118 , \68119 );
buf \U$68147 ( \68121 , \68120 );
buf \U$68148 ( \68122 , \68121 );
and \U$68149 ( \68123 , \68117 , \68122 );
nor \U$68150 ( \68124 , \68116 , \68123 );
buf \U$68151 ( \68125 , \68124 );
buf \U$68152 ( \68126 , \68125 );
not \U$68153 ( \68127 , \68126 );
buf \U$68154 ( \68128 , \67241 );
not \U$68155 ( \68129 , \68128 );
buf \U$68156 ( \68130 , \13460 );
not \U$68157 ( \68131 , \68130 );
or \U$68158 ( \68132 , \68129 , \68131 );
buf \U$68159 ( \68133 , \15793 );
xor \U$68160 ( \68134 , RIc0db098_125, RIc0d7ba0_12);
buf \U$68161 ( \68135 , \68134 );
nand \U$68162 ( \68136 , \68133 , \68135 );
buf \U$68163 ( \68137 , \68136 );
buf \U$68164 ( \68138 , \68137 );
nand \U$68165 ( \68139 , \68132 , \68138 );
buf \U$68166 ( \68140 , \68139 );
buf \U$68167 ( \68141 , \68140 );
not \U$68168 ( \68142 , \68141 );
buf \U$68169 ( \68143 , \67092 );
not \U$68170 ( \68144 , \68143 );
buf \U$68171 ( \68145 , \15995 );
not \U$68172 ( \68146 , \68145 );
or \U$68173 ( \68147 , \68144 , \68146 );
buf \U$68174 ( \68148 , \481 );
xor \U$68175 ( \68149 , RIc0da198_93, RIc0d8aa0_44);
buf \U$68176 ( \68150 , \68149 );
nand \U$68177 ( \68151 , \68148 , \68150 );
buf \U$68178 ( \68152 , \68151 );
buf \U$68179 ( \68153 , \68152 );
nand \U$68180 ( \68154 , \68147 , \68153 );
buf \U$68181 ( \68155 , \68154 );
buf \U$68182 ( \68156 , \68155 );
not \U$68183 ( \68157 , \68156 );
buf \U$68184 ( \68158 , \68157 );
buf \U$68185 ( \68159 , \68158 );
not \U$68186 ( \68160 , \68159 );
or \U$68187 ( \68161 , \68142 , \68160 );
buf \U$68188 ( \68162 , \68158 );
buf \U$68189 ( \68163 , \68140 );
or \U$68190 ( \68164 , \68162 , \68163 );
nand \U$68191 ( \68165 , \68161 , \68164 );
buf \U$68192 ( \68166 , \68165 );
buf \U$68193 ( \68167 , \68166 );
not \U$68194 ( \68168 , \68167 );
or \U$68195 ( \68169 , \68127 , \68168 );
buf \U$68196 ( \68170 , \68166 );
buf \U$68197 ( \68171 , \68125 );
or \U$68198 ( \68172 , \68170 , \68171 );
nand \U$68199 ( \68173 , \68169 , \68172 );
buf \U$68200 ( \68174 , \68173 );
buf \U$68201 ( \68175 , \68174 );
xor \U$68202 ( \68176 , \68113 , \68175 );
not \U$68203 ( \68177 , \921 );
buf \U$68204 ( \68178 , RIc0d8e60_52);
buf \U$68205 ( \68179 , RIc0d9dd8_85);
xor \U$68206 ( \68180 , \68178 , \68179 );
buf \U$68207 ( \68181 , \68180 );
not \U$68208 ( \68182 , \68181 );
or \U$68209 ( \68183 , \68177 , \68182 );
buf \U$68210 ( \68184 , \67182 );
not \U$68211 ( \68185 , \68184 );
buf \U$68212 ( \68186 , \68185 );
or \U$68213 ( \68187 , \954 , \68186 );
nand \U$68214 ( \68188 , \68183 , \68187 );
buf \U$68215 ( \68189 , \68188 );
buf \U$68216 ( \68190 , \67319 );
not \U$68217 ( \68191 , \68190 );
buf \U$68218 ( \68192 , \618 );
not \U$68219 ( \68193 , \68192 );
or \U$68220 ( \68194 , \68191 , \68193 );
buf \U$68221 ( \68195 , \816 );
xor \U$68222 ( \68196 , RIc0d9ec8_87, RIc0d8d70_50);
buf \U$68223 ( \68197 , \68196 );
nand \U$68224 ( \68198 , \68195 , \68197 );
buf \U$68225 ( \68199 , \68198 );
buf \U$68226 ( \68200 , \68199 );
nand \U$68227 ( \68201 , \68194 , \68200 );
buf \U$68228 ( \68202 , \68201 );
buf \U$68229 ( \68203 , \68202 );
xor \U$68230 ( \68204 , \68189 , \68203 );
buf \U$68231 ( \68205 , RIc0d7c90_14);
buf \U$68232 ( \68206 , RIc0dafa8_123);
xor \U$68233 ( \68207 , \68205 , \68206 );
buf \U$68234 ( \68208 , \68207 );
buf \U$68235 ( \68209 , \68208 );
not \U$68236 ( \68210 , \68209 );
buf \U$68237 ( \68211 , \14278 );
not \U$68238 ( \68212 , \68211 );
or \U$68239 ( \68213 , \68210 , \68212 );
buf \U$68240 ( \68214 , \46183 );
buf \U$68241 ( \68215 , \67199 );
or \U$68242 ( \68216 , \68214 , \68215 );
nand \U$68243 ( \68217 , \68213 , \68216 );
buf \U$68244 ( \68218 , \68217 );
buf \U$68245 ( \68219 , \68218 );
xor \U$68246 ( \68220 , \68204 , \68219 );
buf \U$68247 ( \68221 , \68220 );
buf \U$68248 ( \68222 , \68221 );
and \U$68249 ( \68223 , \68176 , \68222 );
and \U$68250 ( \68224 , \68113 , \68175 );
or \U$68251 ( \68225 , \68223 , \68224 );
buf \U$68252 ( \68226 , \68225 );
buf \U$68253 ( \68227 , \68226 );
not \U$68254 ( \68228 , \68227 );
buf \U$68255 ( \68229 , \68228 );
buf \U$68256 ( \68230 , \68229 );
buf \U$68257 ( \68231 , \67247 );
not \U$68258 ( \68232 , \68231 );
buf \U$68259 ( \68233 , \67264 );
not \U$68260 ( \68234 , \68233 );
or \U$68261 ( \68235 , \68232 , \68234 );
buf \U$68262 ( \68236 , \67250 );
not \U$68263 ( \68237 , \68236 );
buf \U$68264 ( \68238 , \67264 );
not \U$68265 ( \68239 , \68238 );
buf \U$68266 ( \68240 , \68239 );
buf \U$68267 ( \68241 , \68240 );
not \U$68268 ( \68242 , \68241 );
or \U$68269 ( \68243 , \68237 , \68242 );
buf \U$68270 ( \68244 , \67231 );
nand \U$68271 ( \68245 , \68243 , \68244 );
buf \U$68272 ( \68246 , \68245 );
buf \U$68273 ( \68247 , \68246 );
nand \U$68274 ( \68248 , \68235 , \68247 );
buf \U$68275 ( \68249 , \68248 );
buf \U$68276 ( \68250 , \68249 );
not \U$68277 ( \68251 , \68250 );
buf \U$68278 ( \68252 , \68251 );
buf \U$68279 ( \68253 , \68252 );
not \U$68280 ( \68254 , \68253 );
buf \U$68281 ( \68255 , \67391 );
not \U$68282 ( \68256 , \68255 );
buf \U$68283 ( \68257 , \16065 );
not \U$68284 ( \68258 , \68257 );
or \U$68285 ( \68259 , \68256 , \68258 );
buf \U$68286 ( \68260 , \12342 );
buf \U$68287 ( \68261 , RIc0d8410_30);
buf \U$68288 ( \68262 , RIc0da828_107);
xor \U$68289 ( \68263 , \68261 , \68262 );
buf \U$68290 ( \68264 , \68263 );
buf \U$68291 ( \68265 , \68264 );
nand \U$68292 ( \68266 , \68260 , \68265 );
buf \U$68293 ( \68267 , \68266 );
buf \U$68294 ( \68268 , \68267 );
nand \U$68295 ( \68269 , \68259 , \68268 );
buf \U$68296 ( \68270 , \68269 );
buf \U$68297 ( \68271 , \67359 );
not \U$68298 ( \68272 , \68271 );
buf \U$68299 ( \68273 , \13991 );
not \U$68300 ( \68274 , \68273 );
or \U$68301 ( \68275 , \68272 , \68274 );
buf \U$68302 ( \68276 , \13998 );
buf \U$68303 ( \68277 , RIc0d9310_62);
buf \U$68304 ( \68278 , RIc0d9928_75);
xor \U$68305 ( \68279 , \68277 , \68278 );
buf \U$68306 ( \68280 , \68279 );
buf \U$68307 ( \68281 , \68280 );
nand \U$68308 ( \68282 , \68276 , \68281 );
buf \U$68309 ( \68283 , \68282 );
buf \U$68310 ( \68284 , \68283 );
nand \U$68311 ( \68285 , \68275 , \68284 );
buf \U$68312 ( \68286 , \68285 );
xor \U$68313 ( \68287 , \68270 , \68286 );
buf \U$68314 ( \68288 , \67075 );
not \U$68315 ( \68289 , \68288 );
buf \U$68316 ( \68290 , \14532 );
not \U$68317 ( \68291 , \68290 );
or \U$68318 ( \68292 , \68289 , \68291 );
buf \U$68319 ( \68293 , RIc0d9040_56);
buf \U$68320 ( \68294 , RIc0d9bf8_81);
xnor \U$68321 ( \68295 , \68293 , \68294 );
buf \U$68322 ( \68296 , \68295 );
buf \U$68323 ( \68297 , \68296 );
not \U$68324 ( \68298 , \68297 );
buf \U$68325 ( \68299 , \1078 );
nand \U$68326 ( \68300 , \68298 , \68299 );
buf \U$68327 ( \68301 , \68300 );
buf \U$68328 ( \68302 , \68301 );
nand \U$68329 ( \68303 , \68292 , \68302 );
buf \U$68330 ( \68304 , \68303 );
xnor \U$68331 ( \68305 , \68287 , \68304 );
buf \U$68332 ( \68306 , \68305 );
not \U$68333 ( \68307 , \68306 );
or \U$68334 ( \68308 , \68254 , \68307 );
buf \U$68335 ( \68309 , \67008 );
not \U$68336 ( \68310 , \68309 );
buf \U$68337 ( \68311 , \15609 );
not \U$68338 ( \68312 , \68311 );
or \U$68339 ( \68313 , \68310 , \68312 );
buf \U$68340 ( \68314 , RIc0d7ab0_10);
buf \U$68341 ( \68315 , RIc0db188_127);
xor \U$68342 ( \68316 , \68314 , \68315 );
buf \U$68343 ( \68317 , \68316 );
buf \U$68344 ( \68318 , \68317 );
buf \U$68345 ( \68319 , RIc0db200_128);
nand \U$68346 ( \68320 , \68318 , \68319 );
buf \U$68347 ( \68321 , \68320 );
buf \U$68348 ( \68322 , \68321 );
nand \U$68349 ( \68323 , \68313 , \68322 );
buf \U$68350 ( \68324 , \68323 );
buf \U$68351 ( \68325 , \68324 );
buf \U$68352 ( \68326 , \67108 );
not \U$68353 ( \68327 , \68326 );
buf \U$68354 ( \68328 , \2535 );
not \U$68355 ( \68329 , \68328 );
or \U$68356 ( \68330 , \68327 , \68329 );
buf \U$68357 ( \68331 , \714 );
xor \U$68358 ( \68332 , RIc0da0a8_91, RIc0d8b90_46);
buf \U$68359 ( \68333 , \68332 );
nand \U$68360 ( \68334 , \68331 , \68333 );
buf \U$68361 ( \68335 , \68334 );
buf \U$68362 ( \68336 , \68335 );
nand \U$68363 ( \68337 , \68330 , \68336 );
buf \U$68364 ( \68338 , \68337 );
buf \U$68365 ( \68339 , \68338 );
xor \U$68366 ( \68340 , \68325 , \68339 );
buf \U$68367 ( \68341 , \20243 );
not \U$68368 ( \68342 , \68341 );
buf \U$68369 ( \68343 , RIc0d85f0_34);
buf \U$68370 ( \68344 , RIc0da648_103);
xor \U$68371 ( \68345 , \68343 , \68344 );
buf \U$68372 ( \68346 , \68345 );
buf \U$68373 ( \68347 , \68346 );
not \U$68374 ( \68348 , \68347 );
or \U$68375 ( \68349 , \68342 , \68348 );
buf \U$68376 ( \68350 , \4483 );
buf \U$68377 ( \68351 , \67142 );
or \U$68378 ( \68352 , \68350 , \68351 );
nand \U$68379 ( \68353 , \68349 , \68352 );
buf \U$68380 ( \68354 , \68353 );
buf \U$68381 ( \68355 , \68354 );
xor \U$68382 ( \68356 , \68340 , \68355 );
buf \U$68383 ( \68357 , \68356 );
buf \U$68384 ( \68358 , \68357 );
nand \U$68385 ( \68359 , \68308 , \68358 );
buf \U$68386 ( \68360 , \68359 );
buf \U$68387 ( \68361 , \68360 );
buf \U$68388 ( \68362 , \68305 );
not \U$68389 ( \68363 , \68362 );
buf \U$68390 ( \68364 , \68249 );
nand \U$68391 ( \68365 , \68363 , \68364 );
buf \U$68392 ( \68366 , \68365 );
buf \U$68393 ( \68367 , \68366 );
nand \U$68394 ( \68368 , \68361 , \68367 );
buf \U$68395 ( \68369 , \68368 );
buf \U$68396 ( \68370 , \68369 );
not \U$68397 ( \68371 , \68370 );
buf \U$68398 ( \68372 , \68371 );
buf \U$68399 ( \68373 , \68372 );
and \U$68400 ( \68374 , \68230 , \68373 );
not \U$68401 ( \68375 , \68230 );
buf \U$68402 ( \68376 , \68369 );
and \U$68403 ( \68377 , \68375 , \68376 );
nor \U$68404 ( \68378 , \68374 , \68377 );
buf \U$68405 ( \68379 , \68378 );
buf \U$68406 ( \68380 , \68379 );
buf \U$68407 ( \68381 , \791 );
buf \U$68408 ( \68382 , RIc0d9400_64);
and \U$68409 ( \68383 , \68381 , \68382 );
buf \U$68410 ( \68384 , \68383 );
buf \U$68411 ( \68385 , \68384 );
buf \U$68412 ( \68386 , \67501 );
not \U$68413 ( \68387 , \68386 );
buf \U$68414 ( \68388 , \1431 );
not \U$68415 ( \68389 , \68388 );
or \U$68416 ( \68390 , \68387 , \68389 );
buf \U$68417 ( \68391 , \1196 );
buf \U$68418 ( \68392 , RIc0d9220_60);
buf \U$68419 ( \68393 , RIc0d9a18_77);
xor \U$68420 ( \68394 , \68392 , \68393 );
buf \U$68421 ( \68395 , \68394 );
buf \U$68422 ( \68396 , \68395 );
nand \U$68423 ( \68397 , \68391 , \68396 );
buf \U$68424 ( \68398 , \68397 );
buf \U$68425 ( \68399 , \68398 );
nand \U$68426 ( \68400 , \68390 , \68399 );
buf \U$68427 ( \68401 , \68400 );
buf \U$68428 ( \68402 , \68401 );
xor \U$68429 ( \68403 , \68385 , \68402 );
buf \U$68430 ( \68404 , \67373 );
not \U$68431 ( \68405 , \68404 );
buf \U$68432 ( \68406 , \3535 );
not \U$68433 ( \68407 , \68406 );
or \U$68434 ( \68408 , \68405 , \68407 );
buf \U$68435 ( \68409 , \15550 );
xor \U$68436 ( \68410 , RIc0da558_101, RIc0d86e0_36);
buf \U$68437 ( \68411 , \68410 );
nand \U$68438 ( \68412 , \68409 , \68411 );
buf \U$68439 ( \68413 , \68412 );
buf \U$68440 ( \68414 , \68413 );
nand \U$68441 ( \68415 , \68408 , \68414 );
buf \U$68442 ( \68416 , \68415 );
buf \U$68443 ( \68417 , \68416 );
xnor \U$68444 ( \68418 , \68403 , \68417 );
buf \U$68445 ( \68419 , \68418 );
buf \U$68446 ( \68420 , \68419 );
not \U$68447 ( \68421 , \68420 );
buf \U$68448 ( \68422 , \67225 );
not \U$68449 ( \68423 , \68422 );
buf \U$68450 ( \68424 , \13684 );
not \U$68451 ( \68425 , \68424 );
or \U$68452 ( \68426 , \68423 , \68425 );
buf \U$68453 ( \68427 , \12937 );
buf \U$68454 ( \68428 , RIc0d7f60_20);
buf \U$68455 ( \68429 , RIc0dacd8_117);
xor \U$68456 ( \68430 , \68428 , \68429 );
buf \U$68457 ( \68431 , \68430 );
buf \U$68458 ( \68432 , \68431 );
nand \U$68459 ( \68433 , \68427 , \68432 );
buf \U$68460 ( \68434 , \68433 );
buf \U$68461 ( \68435 , \68434 );
nand \U$68462 ( \68436 , \68426 , \68435 );
buf \U$68463 ( \68437 , \68436 );
buf \U$68464 ( \68438 , \67433 );
not \U$68465 ( \68439 , \68438 );
buf \U$68466 ( \68440 , \13001 );
not \U$68467 ( \68441 , \68440 );
or \U$68468 ( \68442 , \68439 , \68441 );
buf \U$68469 ( \68443 , \13005 );
buf \U$68470 ( \68444 , RIc0d7e70_18);
buf \U$68471 ( \68445 , RIc0dadc8_119);
xor \U$68472 ( \68446 , \68444 , \68445 );
buf \U$68473 ( \68447 , \68446 );
buf \U$68474 ( \68448 , \68447 );
nand \U$68475 ( \68449 , \68443 , \68448 );
buf \U$68476 ( \68450 , \68449 );
buf \U$68477 ( \68451 , \68450 );
nand \U$68478 ( \68452 , \68442 , \68451 );
buf \U$68479 ( \68453 , \68452 );
xor \U$68480 ( \68454 , \68437 , \68453 );
buf \U$68481 ( \68455 , \67258 );
not \U$68482 ( \68456 , \68455 );
buf \U$68483 ( \68457 , \436 );
not \U$68484 ( \68458 , \68457 );
or \U$68485 ( \68459 , \68456 , \68458 );
buf \U$68486 ( \68460 , \441 );
xor \U$68487 ( \68461 , RIc0d9fb8_89, RIc0d8c80_48);
buf \U$68488 ( \68462 , \68461 );
nand \U$68489 ( \68463 , \68460 , \68462 );
buf \U$68490 ( \68464 , \68463 );
buf \U$68491 ( \68465 , \68464 );
nand \U$68492 ( \68466 , \68459 , \68465 );
buf \U$68493 ( \68467 , \68466 );
not \U$68494 ( \68468 , \68467 );
xor \U$68495 ( \68469 , \68454 , \68468 );
buf \U$68496 ( \68470 , \68469 );
not \U$68497 ( \68471 , \68470 );
or \U$68498 ( \68472 , \68421 , \68471 );
buf \U$68499 ( \68473 , \67165 );
not \U$68500 ( \68474 , \68473 );
buf \U$68501 ( \68475 , \19487 );
not \U$68502 ( \68476 , \68475 );
or \U$68503 ( \68477 , \68474 , \68476 );
buf \U$68504 ( \68478 , \13314 );
buf \U$68505 ( \68479 , RIc0d7d80_16);
buf \U$68506 ( \68480 , RIc0daeb8_121);
xor \U$68507 ( \68481 , \68479 , \68480 );
buf \U$68508 ( \68482 , \68481 );
buf \U$68509 ( \68483 , \68482 );
nand \U$68510 ( \68484 , \68478 , \68483 );
buf \U$68511 ( \68485 , \68484 );
buf \U$68512 ( \68486 , \68485 );
nand \U$68513 ( \68487 , \68477 , \68486 );
buf \U$68514 ( \68488 , \68487 );
buf \U$68515 ( \68489 , \67464 );
not \U$68516 ( \68490 , \68489 );
buf \U$68517 ( \68491 , \13419 );
not \U$68518 ( \68492 , \68491 );
or \U$68519 ( \68493 , \68490 , \68492 );
buf \U$68520 ( \68494 , \20211 );
buf \U$68521 ( \68495 , RIc0d8320_28);
buf \U$68522 ( \68496 , RIc0da918_109);
xor \U$68523 ( \68497 , \68495 , \68496 );
buf \U$68524 ( \68498 , \68497 );
buf \U$68525 ( \68499 , \68498 );
nand \U$68526 ( \68500 , \68494 , \68499 );
buf \U$68527 ( \68501 , \68500 );
buf \U$68528 ( \68502 , \68501 );
nand \U$68529 ( \68503 , \68493 , \68502 );
buf \U$68530 ( \68504 , \68503 );
xor \U$68531 ( \68505 , \68488 , \68504 );
buf \U$68532 ( \68506 , \67415 );
not \U$68533 ( \68507 , \68506 );
buf \U$68534 ( \68508 , \330 );
not \U$68535 ( \68509 , \68508 );
or \U$68536 ( \68510 , \68507 , \68509 );
buf \U$68537 ( \68511 , \344 );
xor \U$68538 ( \68512 , RIc0da288_95, RIc0d89b0_42);
buf \U$68539 ( \68513 , \68512 );
nand \U$68540 ( \68514 , \68511 , \68513 );
buf \U$68541 ( \68515 , \68514 );
buf \U$68542 ( \68516 , \68515 );
nand \U$68543 ( \68517 , \68510 , \68516 );
buf \U$68544 ( \68518 , \68517 );
xor \U$68545 ( \68519 , \68505 , \68518 );
buf \U$68546 ( \68520 , \68519 );
nand \U$68547 ( \68521 , \68472 , \68520 );
buf \U$68548 ( \68522 , \68521 );
buf \U$68549 ( \68523 , \68522 );
buf \U$68550 ( \68524 , \68469 );
not \U$68551 ( \68525 , \68524 );
buf \U$68552 ( \68526 , \68419 );
not \U$68553 ( \68527 , \68526 );
buf \U$68554 ( \68528 , \68527 );
buf \U$68555 ( \68529 , \68528 );
nand \U$68556 ( \68530 , \68525 , \68529 );
buf \U$68557 ( \68531 , \68530 );
buf \U$68558 ( \68532 , \68531 );
nand \U$68559 ( \68533 , \68523 , \68532 );
buf \U$68560 ( \68534 , \68533 );
buf \U$68561 ( \68535 , \68534 );
and \U$68562 ( \68536 , \68380 , \68535 );
not \U$68563 ( \68537 , \68380 );
buf \U$68564 ( \68538 , \68534 );
not \U$68565 ( \68539 , \68538 );
buf \U$68566 ( \68540 , \68539 );
buf \U$68567 ( \68541 , \68540 );
and \U$68568 ( \68542 , \68537 , \68541 );
nor \U$68569 ( \68543 , \68536 , \68542 );
buf \U$68570 ( \68544 , \68543 );
xor \U$68571 ( \68545 , \68058 , \68544 );
xor \U$68572 ( \68546 , \67919 , \68545 );
buf \U$68573 ( \68547 , \67400 );
buf \U$68574 ( \68548 , \67562 );
or \U$68575 ( \68549 , \68547 , \68548 );
buf \U$68576 ( \68550 , \67483 );
nand \U$68577 ( \68551 , \68549 , \68550 );
buf \U$68578 ( \68552 , \68551 );
buf \U$68579 ( \68553 , \68552 );
buf \U$68580 ( \68554 , \67562 );
buf \U$68581 ( \68555 , \67400 );
nand \U$68582 ( \68556 , \68554 , \68555 );
buf \U$68583 ( \68557 , \68556 );
buf \U$68584 ( \68558 , \68557 );
nand \U$68585 ( \68559 , \68553 , \68558 );
buf \U$68586 ( \68560 , \68559 );
buf \U$68587 ( \68561 , \68560 );
xor \U$68588 ( \68562 , \68469 , \68519 );
xnor \U$68589 ( \68563 , \68562 , \68528 );
buf \U$68590 ( \68564 , \68563 );
xor \U$68591 ( \68565 , \68561 , \68564 );
buf \U$68592 ( \68566 , \66811 );
not \U$68593 ( \68567 , \68566 );
buf \U$68594 ( \68568 , \66793 );
not \U$68595 ( \68569 , \68568 );
or \U$68596 ( \68570 , \68567 , \68569 );
buf \U$68597 ( \68571 , \66776 );
nand \U$68598 ( \68572 , \68570 , \68571 );
buf \U$68599 ( \68573 , \68572 );
buf \U$68600 ( \68574 , \68573 );
buf \U$68601 ( \68575 , \66790 );
buf \U$68602 ( \68576 , \66808 );
nand \U$68603 ( \68577 , \68575 , \68576 );
buf \U$68604 ( \68578 , \68577 );
buf \U$68605 ( \68579 , \68578 );
nand \U$68606 ( \68580 , \68574 , \68579 );
buf \U$68607 ( \68581 , \68580 );
buf \U$68608 ( \68582 , \68581 );
and \U$68609 ( \68583 , \68565 , \68582 );
and \U$68610 ( \68584 , \68561 , \68564 );
or \U$68611 ( \68585 , \68583 , \68584 );
buf \U$68612 ( \68586 , \68585 );
buf \U$68613 ( \68587 , \68586 );
not \U$68614 ( \68588 , \68587 );
buf \U$68615 ( \68589 , \68588 );
buf \U$68616 ( \68590 , \68589 );
not \U$68617 ( \68591 , \68590 );
buf \U$68618 ( \68592 , \68249 );
not \U$68619 ( \68593 , \68592 );
buf \U$68620 ( \68594 , \68305 );
not \U$68621 ( \68595 , \68594 );
or \U$68622 ( \68596 , \68593 , \68595 );
buf \U$68623 ( \68597 , \68249 );
buf \U$68624 ( \68598 , \68305 );
or \U$68625 ( \68599 , \68597 , \68598 );
nand \U$68626 ( \68600 , \68596 , \68599 );
buf \U$68627 ( \68601 , \68600 );
buf \U$68628 ( \68602 , \68601 );
buf \U$68629 ( \68603 , \68357 );
not \U$68630 ( \68604 , \68603 );
buf \U$68631 ( \68605 , \68604 );
buf \U$68632 ( \68606 , \68605 );
and \U$68633 ( \68607 , \68602 , \68606 );
not \U$68634 ( \68608 , \68602 );
buf \U$68635 ( \68609 , \68357 );
and \U$68636 ( \68610 , \68608 , \68609 );
nor \U$68637 ( \68611 , \68607 , \68610 );
buf \U$68638 ( \68612 , \68611 );
buf \U$68639 ( \68613 , \68612 );
not \U$68640 ( \68614 , \68613 );
buf \U$68641 ( \68615 , \67210 );
not \U$68642 ( \68616 , \68615 );
buf \U$68643 ( \68617 , \67332 );
not \U$68644 ( \68618 , \68617 );
or \U$68645 ( \68619 , \68616 , \68618 );
buf \U$68646 ( \68620 , \67213 );
not \U$68647 ( \68621 , \68620 );
buf \U$68648 ( \68622 , \67326 );
not \U$68649 ( \68623 , \68622 );
or \U$68650 ( \68624 , \68621 , \68623 );
buf \U$68651 ( \68625 , \67268 );
nand \U$68652 ( \68626 , \68624 , \68625 );
buf \U$68653 ( \68627 , \68626 );
buf \U$68654 ( \68628 , \68627 );
nand \U$68655 ( \68629 , \68619 , \68628 );
buf \U$68656 ( \68630 , \68629 );
buf \U$68657 ( \68631 , \68630 );
not \U$68658 ( \68632 , \68631 );
buf \U$68659 ( \68633 , \68632 );
buf \U$68660 ( \68634 , \68633 );
not \U$68661 ( \68635 , \68634 );
or \U$68662 ( \68636 , \68614 , \68635 );
xor \U$68663 ( \68637 , \68113 , \68175 );
xor \U$68664 ( \68638 , \68637 , \68222 );
buf \U$68665 ( \68639 , \68638 );
buf \U$68666 ( \68640 , \68639 );
nand \U$68667 ( \68641 , \68636 , \68640 );
buf \U$68668 ( \68642 , \68641 );
buf \U$68669 ( \68643 , \68642 );
buf \U$68670 ( \68644 , \68630 );
buf \U$68671 ( \68645 , \68612 );
not \U$68672 ( \68646 , \68645 );
buf \U$68673 ( \68647 , \68646 );
buf \U$68674 ( \68648 , \68647 );
nand \U$68675 ( \68649 , \68644 , \68648 );
buf \U$68676 ( \68650 , \68649 );
buf \U$68677 ( \68651 , \68650 );
nand \U$68678 ( \68652 , \68643 , \68651 );
buf \U$68679 ( \68653 , \68652 );
buf \U$68680 ( \68654 , \68653 );
not \U$68681 ( \68655 , \68654 );
buf \U$68682 ( \68656 , \67861 );
not \U$68683 ( \68657 , \68656 );
buf \U$68684 ( \68658 , \67867 );
not \U$68685 ( \68659 , \68658 );
or \U$68686 ( \68660 , \68657 , \68659 );
buf \U$68687 ( \68661 , \67867 );
buf \U$68688 ( \68662 , \67861 );
or \U$68689 ( \68663 , \68661 , \68662 );
buf \U$68690 ( \68664 , \67874 );
nand \U$68691 ( \68665 , \68663 , \68664 );
buf \U$68692 ( \68666 , \68665 );
buf \U$68693 ( \68667 , \68666 );
nand \U$68694 ( \68668 , \68660 , \68667 );
buf \U$68695 ( \68669 , \68668 );
buf \U$68696 ( \68670 , \68280 );
not \U$68697 ( \68671 , \68670 );
buf \U$68698 ( \68672 , \1556 );
not \U$68699 ( \68673 , \68672 );
or \U$68700 ( \68674 , \68671 , \68673 );
buf \U$68701 ( \68675 , \1143 );
xor \U$68702 ( \68676 , RIc0d9928_75, RIc0d9298_61);
buf \U$68703 ( \68677 , \68676 );
nand \U$68704 ( \68678 , \68675 , \68677 );
buf \U$68705 ( \68679 , \68678 );
buf \U$68706 ( \68680 , \68679 );
nand \U$68707 ( \68681 , \68674 , \68680 );
buf \U$68708 ( \68682 , \68681 );
buf \U$68709 ( \68683 , \68682 );
not \U$68710 ( \68684 , \68683 );
buf \U$68711 ( \68685 , RIc0d9400_64);
buf \U$68712 ( \68686 , RIc0d98b0_74);
or \U$68713 ( \68687 , \68685 , \68686 );
buf \U$68714 ( \68688 , RIc0d9928_75);
nand \U$68715 ( \68689 , \68687 , \68688 );
buf \U$68716 ( \68690 , \68689 );
buf \U$68717 ( \68691 , \68690 );
buf \U$68718 ( \68692 , RIc0d9400_64);
buf \U$68719 ( \68693 , RIc0d98b0_74);
nand \U$68720 ( \68694 , \68692 , \68693 );
buf \U$68721 ( \68695 , \68694 );
buf \U$68722 ( \68696 , \68695 );
buf \U$68723 ( \68697 , RIc0d9838_73);
nand \U$68724 ( \68698 , \68691 , \68696 , \68697 );
buf \U$68725 ( \68699 , \68698 );
buf \U$68726 ( \68700 , \68699 );
not \U$68727 ( \68701 , \68700 );
and \U$68728 ( \68702 , \68684 , \68701 );
buf \U$68729 ( \68703 , \68682 );
buf \U$68730 ( \68704 , \68699 );
and \U$68731 ( \68705 , \68703 , \68704 );
nor \U$68732 ( \68706 , \68702 , \68705 );
buf \U$68733 ( \68707 , \68706 );
buf \U$68734 ( \68708 , \68707 );
not \U$68735 ( \68709 , \68708 );
buf \U$68736 ( \68710 , \68467 );
not \U$68737 ( \68711 , \68710 );
buf \U$68738 ( \68712 , \68453 );
not \U$68739 ( \68713 , \68712 );
or \U$68740 ( \68714 , \68711 , \68713 );
buf \U$68741 ( \68715 , \68453 );
buf \U$68742 ( \68716 , \68467 );
or \U$68743 ( \68717 , \68715 , \68716 );
buf \U$68744 ( \68718 , \68437 );
nand \U$68745 ( \68719 , \68717 , \68718 );
buf \U$68746 ( \68720 , \68719 );
buf \U$68747 ( \68721 , \68720 );
nand \U$68748 ( \68722 , \68714 , \68721 );
buf \U$68749 ( \68723 , \68722 );
buf \U$68750 ( \68724 , \68723 );
not \U$68751 ( \68725 , \68724 );
or \U$68752 ( \68726 , \68709 , \68725 );
buf \U$68753 ( \68727 , \68723 );
buf \U$68754 ( \68728 , \68707 );
or \U$68755 ( \68729 , \68727 , \68728 );
nand \U$68756 ( \68730 , \68726 , \68729 );
buf \U$68757 ( \68731 , \68730 );
buf \U$68758 ( \68732 , \68731 );
not \U$68759 ( \68733 , \68732 );
buf \U$68760 ( \68734 , \68504 );
not \U$68761 ( \68735 , \68734 );
buf \U$68762 ( \68736 , \68518 );
not \U$68763 ( \68737 , \68736 );
or \U$68764 ( \68738 , \68735 , \68737 );
buf \U$68765 ( \68739 , \68518 );
buf \U$68766 ( \68740 , \68504 );
or \U$68767 ( \68741 , \68739 , \68740 );
buf \U$68768 ( \68742 , \68488 );
nand \U$68769 ( \68743 , \68741 , \68742 );
buf \U$68770 ( \68744 , \68743 );
buf \U$68771 ( \68745 , \68744 );
nand \U$68772 ( \68746 , \68738 , \68745 );
buf \U$68773 ( \68747 , \68746 );
buf \U$68774 ( \68748 , \68747 );
not \U$68775 ( \68749 , \68748 );
buf \U$68776 ( \68750 , \68749 );
buf \U$68777 ( \68751 , \68750 );
not \U$68778 ( \68752 , \68751 );
and \U$68779 ( \68753 , \68733 , \68752 );
buf \U$68780 ( \68754 , \68731 );
buf \U$68781 ( \68755 , \68750 );
and \U$68782 ( \68756 , \68754 , \68755 );
nor \U$68783 ( \68757 , \68753 , \68756 );
buf \U$68784 ( \68758 , \68757 );
xor \U$68785 ( \68759 , \68669 , \68758 );
xor \U$68786 ( \68760 , \68325 , \68339 );
and \U$68787 ( \68761 , \68760 , \68355 );
and \U$68788 ( \68762 , \68325 , \68339 );
or \U$68789 ( \68763 , \68761 , \68762 );
buf \U$68790 ( \68764 , \68763 );
buf \U$68791 ( \68765 , \68764 );
xor \U$68792 ( \68766 , \68189 , \68203 );
and \U$68793 ( \68767 , \68766 , \68219 );
and \U$68794 ( \68768 , \68189 , \68203 );
or \U$68795 ( \68769 , \68767 , \68768 );
buf \U$68796 ( \68770 , \68769 );
buf \U$68797 ( \68771 , \68770 );
xor \U$68798 ( \68772 , \68765 , \68771 );
xor \U$68799 ( \68773 , \68075 , \68092 );
and \U$68800 ( \68774 , \68773 , \68110 );
and \U$68801 ( \68775 , \68075 , \68092 );
or \U$68802 ( \68776 , \68774 , \68775 );
buf \U$68803 ( \68777 , \68776 );
buf \U$68804 ( \68778 , \68777 );
xor \U$68805 ( \68779 , \68772 , \68778 );
buf \U$68806 ( \68780 , \68779 );
xor \U$68807 ( \68781 , \68759 , \68780 );
buf \U$68808 ( \68782 , \68781 );
not \U$68809 ( \68783 , \68782 );
or \U$68810 ( \68784 , \68655 , \68783 );
buf \U$68811 ( \68785 , \68653 );
buf \U$68812 ( \68786 , \68781 );
or \U$68813 ( \68787 , \68785 , \68786 );
nand \U$68814 ( \68788 , \68784 , \68787 );
buf \U$68815 ( \68789 , \68788 );
buf \U$68816 ( \68790 , \68789 );
not \U$68817 ( \68791 , \68790 );
and \U$68818 ( \68792 , \68591 , \68791 );
buf \U$68819 ( \68793 , \68589 );
buf \U$68820 ( \68794 , \68789 );
and \U$68821 ( \68795 , \68793 , \68794 );
nor \U$68822 ( \68796 , \68792 , \68795 );
buf \U$68823 ( \68797 , \68796 );
and \U$68824 ( \68798 , \68546 , \68797 );
not \U$68825 ( \68799 , \68546 );
buf \U$68826 ( \68800 , \68797 );
not \U$68827 ( \68801 , \68800 );
buf \U$68828 ( \68802 , \68801 );
and \U$68829 ( \68803 , \68799 , \68802 );
nor \U$68830 ( \68804 , \68798 , \68803 );
buf \U$68831 ( \68805 , \68804 );
xor \U$68832 ( \68806 , \66998 , \67569 );
and \U$68833 ( \68807 , \68806 , \67576 );
and \U$68834 ( \68808 , \66998 , \67569 );
or \U$68835 ( \68809 , \68807 , \68808 );
buf \U$68836 ( \68810 , \68809 );
buf \U$68837 ( \68811 , \68810 );
buf \U$68838 ( \68812 , \68633 );
not \U$68839 ( \68813 , \68812 );
buf \U$68840 ( \68814 , \68639 );
not \U$68841 ( \68815 , \68814 );
or \U$68842 ( \68816 , \68813 , \68815 );
buf \U$68843 ( \68817 , \68639 );
buf \U$68844 ( \68818 , \68633 );
or \U$68845 ( \68819 , \68817 , \68818 );
nand \U$68846 ( \68820 , \68816 , \68819 );
buf \U$68847 ( \68821 , \68820 );
buf \U$68848 ( \68822 , \68821 );
buf \U$68849 ( \68823 , \68612 );
and \U$68850 ( \68824 , \68822 , \68823 );
not \U$68851 ( \68825 , \68822 );
buf \U$68852 ( \68826 , \68647 );
and \U$68853 ( \68827 , \68825 , \68826 );
nor \U$68854 ( \68828 , \68824 , \68827 );
buf \U$68855 ( \68829 , \68828 );
buf \U$68856 ( \68830 , \68829 );
not \U$68857 ( \68831 , \68830 );
xor \U$68858 ( \68832 , \68561 , \68564 );
xor \U$68859 ( \68833 , \68832 , \68582 );
buf \U$68860 ( \68834 , \68833 );
buf \U$68861 ( \68835 , \68834 );
not \U$68862 ( \68836 , \68835 );
or \U$68863 ( \68837 , \68831 , \68836 );
buf \U$68864 ( \68838 , \68834 );
buf \U$68865 ( \68839 , \68829 );
or \U$68866 ( \68840 , \68838 , \68839 );
nand \U$68867 ( \68841 , \68837 , \68840 );
buf \U$68868 ( \68842 , \68841 );
buf \U$68869 ( \68843 , \68842 );
buf \U$68870 ( \68844 , \66761 );
not \U$68871 ( \68845 , \68844 );
buf \U$68872 ( \68846 , \66812 );
not \U$68873 ( \68847 , \68846 );
or \U$68874 ( \68848 , \68845 , \68847 );
buf \U$68875 ( \68849 , \66753 );
nand \U$68876 ( \68850 , \68848 , \68849 );
buf \U$68877 ( \68851 , \68850 );
buf \U$68878 ( \68852 , \68851 );
buf \U$68879 ( \68853 , \66815 );
buf \U$68880 ( \68854 , \66758 );
nand \U$68881 ( \68855 , \68853 , \68854 );
buf \U$68882 ( \68856 , \68855 );
buf \U$68883 ( \68857 , \68856 );
nand \U$68884 ( \68858 , \68852 , \68857 );
buf \U$68885 ( \68859 , \68858 );
buf \U$68886 ( \68860 , \68859 );
and \U$68887 ( \68861 , \68843 , \68860 );
not \U$68888 ( \68862 , \68843 );
buf \U$68889 ( \68863 , \68859 );
not \U$68890 ( \68864 , \68863 );
buf \U$68891 ( \68865 , \68864 );
buf \U$68892 ( \68866 , \68865 );
and \U$68893 ( \68867 , \68862 , \68866 );
nor \U$68894 ( \68868 , \68861 , \68867 );
buf \U$68895 ( \68869 , \68868 );
buf \U$68896 ( \68870 , \68869 );
xor \U$68897 ( \68871 , \68811 , \68870 );
buf \U$68898 ( \68872 , \66816 );
not \U$68899 ( \68873 , \68872 );
buf \U$68900 ( \68874 , \66977 );
not \U$68901 ( \68875 , \68874 );
or \U$68902 ( \68876 , \68873 , \68875 );
buf \U$68903 ( \68877 , \66977 );
buf \U$68904 ( \68878 , \66816 );
or \U$68905 ( \68879 , \68877 , \68878 );
buf \U$68906 ( \68880 , \66821 );
nand \U$68907 ( \68881 , \68879 , \68880 );
buf \U$68908 ( \68882 , \68881 );
buf \U$68909 ( \68883 , \68882 );
nand \U$68910 ( \68884 , \68876 , \68883 );
buf \U$68911 ( \68885 , \68884 );
buf \U$68912 ( \68886 , \68885 );
and \U$68913 ( \68887 , \68871 , \68886 );
and \U$68914 ( \68888 , \68811 , \68870 );
or \U$68915 ( \68889 , \68887 , \68888 );
buf \U$68916 ( \68890 , \68889 );
buf \U$68917 ( \68891 , \68890 );
xor \U$68918 ( \68892 , \68805 , \68891 );
buf \U$68919 ( \68893 , \68834 );
not \U$68920 ( \68894 , \68893 );
buf \U$68921 ( \68895 , \68865 );
nand \U$68922 ( \68896 , \68894 , \68895 );
buf \U$68923 ( \68897 , \68896 );
buf \U$68924 ( \68898 , \68897 );
buf \U$68925 ( \68899 , \68829 );
not \U$68926 ( \68900 , \68899 );
buf \U$68927 ( \68901 , \68900 );
buf \U$68928 ( \68902 , \68901 );
and \U$68929 ( \68903 , \68898 , \68902 );
buf \U$68930 ( \68904 , \68834 );
not \U$68931 ( \68905 , \68904 );
buf \U$68932 ( \68906 , \68865 );
nor \U$68933 ( \68907 , \68905 , \68906 );
buf \U$68934 ( \68908 , \68907 );
buf \U$68935 ( \68909 , \68908 );
nor \U$68936 ( \68910 , \68903 , \68909 );
buf \U$68937 ( \68911 , \68910 );
buf \U$68938 ( \68912 , \68911 );
buf \U$68939 ( \68913 , \68158 );
not \U$68940 ( \68914 , \68913 );
buf \U$68941 ( \68915 , \68125 );
not \U$68942 ( \68916 , \68915 );
or \U$68943 ( \68917 , \68914 , \68916 );
buf \U$68944 ( \68918 , \68140 );
nand \U$68945 ( \68919 , \68917 , \68918 );
buf \U$68946 ( \68920 , \68919 );
buf \U$68947 ( \68921 , \68920 );
buf \U$68948 ( \68922 , \68125 );
not \U$68949 ( \68923 , \68922 );
buf \U$68950 ( \68924 , \68155 );
nand \U$68951 ( \68925 , \68923 , \68924 );
buf \U$68952 ( \68926 , \68925 );
buf \U$68953 ( \68927 , \68926 );
nand \U$68954 ( \68928 , \68921 , \68927 );
buf \U$68955 ( \68929 , \68928 );
buf \U$68956 ( \68930 , \68929 );
not \U$68957 ( \68931 , \68930 );
buf \U$68958 ( \68932 , \68931 );
buf \U$68959 ( \68933 , \68932 );
not \U$68960 ( \68934 , \68933 );
buf \U$68961 ( \68935 , \68317 );
not \U$68962 ( \68936 , \68935 );
buf \U$68963 ( \68937 , \43780 );
not \U$68964 ( \68938 , \68937 );
or \U$68965 ( \68939 , \68936 , \68938 );
buf \U$68966 ( \68940 , RIc0d7a38_9);
buf \U$68967 ( \68941 , RIc0db188_127);
xor \U$68968 ( \68942 , \68940 , \68941 );
buf \U$68969 ( \68943 , \68942 );
buf \U$68970 ( \68944 , \68943 );
buf \U$68971 ( \68945 , RIc0db200_128);
nand \U$68972 ( \68946 , \68944 , \68945 );
buf \U$68973 ( \68947 , \68946 );
buf \U$68974 ( \68948 , \68947 );
nand \U$68975 ( \68949 , \68939 , \68948 );
buf \U$68976 ( \68950 , \68949 );
buf \U$68977 ( \68951 , \68950 );
xor \U$68978 ( \68952 , RIc0daaf8_113, RIc0d8140_24);
buf \U$68979 ( \68953 , \68952 );
not \U$68980 ( \68954 , \68953 );
buf \U$68981 ( \68955 , \28776 );
not \U$68982 ( \68956 , \68955 );
or \U$68983 ( \68957 , \68954 , \68956 );
buf \U$68984 ( \68958 , \16995 );
xor \U$68985 ( \68959 , RIc0daaf8_113, RIc0d80c8_23);
buf \U$68986 ( \68960 , \68959 );
nand \U$68987 ( \68961 , \68958 , \68960 );
buf \U$68988 ( \68962 , \68961 );
buf \U$68989 ( \68963 , \68962 );
nand \U$68990 ( \68964 , \68957 , \68963 );
buf \U$68991 ( \68965 , \68964 );
buf \U$68992 ( \68966 , \68965 );
xor \U$68993 ( \68967 , \68951 , \68966 );
buf \U$68994 ( \68968 , \68103 );
not \U$68995 ( \68969 , \68968 );
buf \U$68996 ( \68970 , \13092 );
not \U$68997 ( \68971 , \68970 );
or \U$68998 ( \68972 , \68969 , \68971 );
buf \U$68999 ( \68973 , \734 );
buf \U$69000 ( \68974 , \20273 );
nand \U$69001 ( \68975 , \68973 , \68974 );
buf \U$69002 ( \68976 , \68975 );
buf \U$69003 ( \68977 , \68976 );
nand \U$69004 ( \68978 , \68972 , \68977 );
buf \U$69005 ( \68979 , \68978 );
buf \U$69006 ( \68980 , \68979 );
xor \U$69007 ( \68981 , \68967 , \68980 );
buf \U$69008 ( \68982 , \68981 );
buf \U$69009 ( \68983 , \68982 );
not \U$69010 ( \68984 , \68983 );
or \U$69011 ( \68985 , \68934 , \68984 );
buf \U$69012 ( \68986 , \68982 );
buf \U$69013 ( \68987 , \68932 );
or \U$69014 ( \68988 , \68986 , \68987 );
nand \U$69015 ( \68989 , \68985 , \68988 );
buf \U$69016 ( \68990 , \68989 );
buf \U$69017 ( \68991 , \68990 );
buf \U$69018 ( \68992 , \68121 );
not \U$69019 ( \68993 , \68992 );
buf \U$69020 ( \68994 , \12361 );
not \U$69021 ( \68995 , \68994 );
or \U$69022 ( \68996 , \68993 , \68995 );
buf \U$69023 ( \68997 , \402 );
buf \U$69024 ( \68998 , RIc0d90b8_57);
buf \U$69025 ( \68999 , RIc0d9b08_79);
xor \U$69026 ( \69000 , \68998 , \68999 );
buf \U$69027 ( \69001 , \69000 );
buf \U$69028 ( \69002 , \69001 );
nand \U$69029 ( \69003 , \68997 , \69002 );
buf \U$69030 ( \69004 , \69003 );
buf \U$69031 ( \69005 , \69004 );
nand \U$69032 ( \69006 , \68996 , \69005 );
buf \U$69033 ( \69007 , \69006 );
not \U$69034 ( \69008 , \69007 );
buf \U$69035 ( \69009 , \68395 );
not \U$69036 ( \69010 , \69009 );
buf \U$69037 ( \69011 , \14825 );
not \U$69038 ( \69012 , \69011 );
or \U$69039 ( \69013 , \69010 , \69012 );
buf \U$69040 ( \69014 , \3742 );
buf \U$69041 ( \69015 , RIc0d91a8_59);
buf \U$69042 ( \69016 , RIc0d9a18_77);
xor \U$69043 ( \69017 , \69015 , \69016 );
buf \U$69044 ( \69018 , \69017 );
buf \U$69045 ( \69019 , \69018 );
nand \U$69046 ( \69020 , \69014 , \69019 );
buf \U$69047 ( \69021 , \69020 );
buf \U$69048 ( \69022 , \69021 );
nand \U$69049 ( \69023 , \69013 , \69022 );
buf \U$69050 ( \69024 , \69023 );
buf \U$69051 ( \69025 , \69024 );
not \U$69052 ( \69026 , \69025 );
buf \U$69053 ( \69027 , \69026 );
not \U$69054 ( \69028 , \69027 );
or \U$69055 ( \69029 , \69008 , \69028 );
buf \U$69056 ( \69030 , \69024 );
buf \U$69057 ( \69031 , \69007 );
not \U$69058 ( \69032 , \69031 );
buf \U$69059 ( \69033 , \69032 );
buf \U$69060 ( \69034 , \69033 );
nand \U$69061 ( \69035 , \69030 , \69034 );
buf \U$69062 ( \69036 , \69035 );
nand \U$69063 ( \69037 , \69029 , \69036 );
buf \U$69064 ( \69038 , \68332 );
not \U$69065 ( \69039 , \69038 );
buf \U$69066 ( \69040 , \704 );
not \U$69067 ( \69041 , \69040 );
or \U$69068 ( \69042 , \69039 , \69041 );
buf \U$69069 ( \69043 , \714 );
buf \U$69070 ( \69044 , RIc0d8b18_45);
buf \U$69071 ( \69045 , RIc0da0a8_91);
xor \U$69072 ( \69046 , \69044 , \69045 );
buf \U$69073 ( \69047 , \69046 );
buf \U$69074 ( \69048 , \69047 );
nand \U$69075 ( \69049 , \69043 , \69048 );
buf \U$69076 ( \69050 , \69049 );
buf \U$69077 ( \69051 , \69050 );
nand \U$69078 ( \69052 , \69042 , \69051 );
buf \U$69079 ( \69053 , \69052 );
xnor \U$69080 ( \69054 , \69037 , \69053 );
buf \U$69081 ( \69055 , \69054 );
not \U$69082 ( \69056 , \69055 );
buf \U$69083 ( \69057 , \69056 );
buf \U$69084 ( \69058 , \69057 );
and \U$69085 ( \69059 , \68991 , \69058 );
not \U$69086 ( \69060 , \68991 );
buf \U$69087 ( \69061 , \69054 );
and \U$69088 ( \69062 , \69060 , \69061 );
nor \U$69089 ( \69063 , \69059 , \69062 );
buf \U$69090 ( \69064 , \69063 );
buf \U$69091 ( \69065 , \69064 );
not \U$69092 ( \69066 , \69065 );
buf \U$69093 ( \69067 , \68384 );
not \U$69094 ( \69068 , \69067 );
buf \U$69095 ( \69069 , \68401 );
not \U$69096 ( \69070 , \69069 );
or \U$69097 ( \69071 , \69068 , \69070 );
buf \U$69098 ( \69072 , \68401 );
buf \U$69099 ( \69073 , \68384 );
or \U$69100 ( \69074 , \69072 , \69073 );
buf \U$69101 ( \69075 , \68416 );
nand \U$69102 ( \69076 , \69074 , \69075 );
buf \U$69103 ( \69077 , \69076 );
buf \U$69104 ( \69078 , \69077 );
nand \U$69105 ( \69079 , \69071 , \69078 );
buf \U$69106 ( \69080 , \69079 );
buf \U$69107 ( \69081 , \15644 );
not \U$69108 ( \69082 , \69081 );
buf \U$69109 ( \69083 , \67040 );
nor \U$69110 ( \69084 , \69082 , \69083 );
buf \U$69111 ( \69085 , \69084 );
buf \U$69112 ( \69086 , \69085 );
buf \U$69113 ( \69087 , \26301 );
not \U$69114 ( \69088 , \69087 );
buf \U$69115 ( \69089 , \67923 );
nor \U$69116 ( \69090 , \69088 , \69089 );
buf \U$69117 ( \69091 , \69090 );
buf \U$69118 ( \69092 , \69091 );
nor \U$69119 ( \69093 , \69086 , \69092 );
buf \U$69120 ( \69094 , \69093 );
buf \U$69121 ( \69095 , \69094 );
not \U$69122 ( \69096 , \69095 );
buf \U$69123 ( \69097 , \67023 );
not \U$69124 ( \69098 , \69097 );
buf \U$69125 ( \69099 , \16656 );
not \U$69126 ( \69100 , \69099 );
or \U$69127 ( \69101 , \69098 , \69100 );
buf \U$69128 ( \69102 , \12410 );
buf \U$69129 ( \69103 , \68952 );
nand \U$69130 ( \69104 , \69102 , \69103 );
buf \U$69131 ( \69105 , \69104 );
buf \U$69132 ( \69106 , \69105 );
nand \U$69133 ( \69107 , \69101 , \69106 );
buf \U$69134 ( \69108 , \69107 );
buf \U$69135 ( \69109 , \69108 );
not \U$69136 ( \69110 , \69109 );
buf \U$69137 ( \69111 , \69110 );
buf \U$69138 ( \69112 , \69111 );
not \U$69139 ( \69113 , \69112 );
or \U$69140 ( \69114 , \69096 , \69113 );
buf \U$69141 ( \69115 , \67528 );
not \U$69142 ( \69116 , \69115 );
buf \U$69143 ( \69117 , \19695 );
not \U$69144 ( \69118 , \69117 );
or \U$69145 ( \69119 , \69116 , \69118 );
buf \U$69146 ( \69120 , \12584 );
buf \U$69147 ( \69121 , \67943 );
nand \U$69148 ( \69122 , \69120 , \69121 );
buf \U$69149 ( \69123 , \69122 );
buf \U$69150 ( \69124 , \69123 );
nand \U$69151 ( \69125 , \69119 , \69124 );
buf \U$69152 ( \69126 , \69125 );
buf \U$69153 ( \69127 , \69126 );
nand \U$69154 ( \69128 , \69114 , \69127 );
buf \U$69155 ( \69129 , \69128 );
buf \U$69156 ( \69130 , \69129 );
buf \U$69157 ( \69131 , \69094 );
not \U$69158 ( \69132 , \69131 );
buf \U$69159 ( \69133 , \69108 );
nand \U$69160 ( \69134 , \69132 , \69133 );
buf \U$69161 ( \69135 , \69134 );
buf \U$69162 ( \69136 , \69135 );
nand \U$69163 ( \69137 , \69130 , \69136 );
buf \U$69164 ( \69138 , \69137 );
xor \U$69165 ( \69139 , \69080 , \69138 );
buf \U$69166 ( \69140 , \68286 );
not \U$69167 ( \69141 , \69140 );
buf \U$69168 ( \69142 , \68304 );
not \U$69169 ( \69143 , \69142 );
or \U$69170 ( \69144 , \69141 , \69143 );
buf \U$69171 ( \69145 , \68304 );
buf \U$69172 ( \69146 , \68286 );
or \U$69173 ( \69147 , \69145 , \69146 );
buf \U$69174 ( \69148 , \68270 );
nand \U$69175 ( \69149 , \69147 , \69148 );
buf \U$69176 ( \69150 , \69149 );
buf \U$69177 ( \69151 , \69150 );
nand \U$69178 ( \69152 , \69144 , \69151 );
buf \U$69179 ( \69153 , \69152 );
xnor \U$69180 ( \69154 , \69139 , \69153 );
buf \U$69181 ( \69155 , \69154 );
not \U$69182 ( \69156 , \69155 );
or \U$69183 ( \69157 , \69066 , \69156 );
buf \U$69184 ( \69158 , \69154 );
buf \U$69185 ( \69159 , \69064 );
or \U$69186 ( \69160 , \69158 , \69159 );
nand \U$69187 ( \69161 , \69157 , \69160 );
buf \U$69188 ( \69162 , \69161 );
buf \U$69189 ( \69163 , \69162 );
buf \U$69190 ( \69164 , \68498 );
not \U$69191 ( \69165 , \69164 );
buf \U$69192 ( \69166 , \27660 );
not \U$69193 ( \69167 , \69166 );
or \U$69194 ( \69168 , \69165 , \69167 );
buf \U$69195 ( \69169 , \16232 );
buf \U$69196 ( \69170 , \20205 );
nand \U$69197 ( \69171 , \69169 , \69170 );
buf \U$69198 ( \69172 , \69171 );
buf \U$69199 ( \69173 , \69172 );
nand \U$69200 ( \69174 , \69168 , \69173 );
buf \U$69201 ( \69175 , \69174 );
buf \U$69202 ( \69176 , \69175 );
not \U$69203 ( \69177 , \69176 );
buf \U$69204 ( \69178 , \68181 );
not \U$69205 ( \69179 , \69178 );
buf \U$69206 ( \69180 , \13737 );
not \U$69207 ( \69181 , \69180 );
or \U$69208 ( \69182 , \69179 , \69181 );
buf \U$69209 ( \69183 , \2960 );
buf \U$69210 ( \69184 , \20113 );
nand \U$69211 ( \69185 , \69183 , \69184 );
buf \U$69212 ( \69186 , \69185 );
buf \U$69213 ( \69187 , \69186 );
nand \U$69214 ( \69188 , \69182 , \69187 );
buf \U$69215 ( \69189 , \69188 );
buf \U$69216 ( \69190 , \69189 );
not \U$69217 ( \69191 , \69190 );
buf \U$69218 ( \69192 , \69191 );
buf \U$69219 ( \69193 , \69192 );
not \U$69220 ( \69194 , \69193 );
or \U$69221 ( \69195 , \69177 , \69194 );
buf \U$69222 ( \69196 , \69175 );
buf \U$69223 ( \69197 , \69192 );
or \U$69224 ( \69198 , \69196 , \69197 );
nand \U$69225 ( \69199 , \69195 , \69198 );
buf \U$69226 ( \69200 , \69199 );
buf \U$69227 ( \69201 , \69200 );
not \U$69228 ( \69202 , \69201 );
buf \U$69229 ( \69203 , \1078 );
buf \U$69230 ( \69204 , \20159 );
and \U$69231 ( \69205 , \69203 , \69204 );
buf \U$69232 ( \69206 , \69205 );
buf \U$69233 ( \69207 , \69206 );
buf \U$69234 ( \69208 , \1060 );
buf \U$69235 ( \69209 , \68296 );
nor \U$69236 ( \69210 , \69208 , \69209 );
buf \U$69237 ( \69211 , \69210 );
buf \U$69238 ( \69212 , \69211 );
nor \U$69239 ( \69213 , \69207 , \69212 );
buf \U$69240 ( \69214 , \69213 );
buf \U$69241 ( \69215 , \69214 );
not \U$69242 ( \69216 , \69215 );
and \U$69243 ( \69217 , \69202 , \69216 );
buf \U$69244 ( \69218 , \69200 );
buf \U$69245 ( \69219 , \69214 );
and \U$69246 ( \69220 , \69218 , \69219 );
nor \U$69247 ( \69221 , \69217 , \69220 );
buf \U$69248 ( \69222 , \69221 );
buf \U$69249 ( \69223 , \69222 );
not \U$69250 ( \69224 , \69223 );
buf \U$69251 ( \69225 , \68512 );
not \U$69252 ( \69226 , \69225 );
buf \U$69253 ( \69227 , \13860 );
not \U$69254 ( \69228 , \69227 );
or \U$69255 ( \69229 , \69226 , \69228 );
buf \U$69256 ( \69230 , \13873 );
buf \U$69257 ( \69231 , \20184 );
nand \U$69258 ( \69232 , \69230 , \69231 );
buf \U$69259 ( \69233 , \69232 );
buf \U$69260 ( \69234 , \69233 );
nand \U$69261 ( \69235 , \69229 , \69234 );
buf \U$69262 ( \69236 , \69235 );
buf \U$69263 ( \69237 , \69236 );
not \U$69264 ( \69238 , \69237 );
buf \U$69265 ( \69239 , \68208 );
not \U$69266 ( \69240 , \69239 );
buf \U$69267 ( \69241 , \14982 );
not \U$69268 ( \69242 , \69241 );
or \U$69269 ( \69243 , \69240 , \69242 );
buf \U$69270 ( \69244 , \16692 );
buf \U$69271 ( \69245 , RIc0d7c18_13);
buf \U$69272 ( \69246 , RIc0dafa8_123);
xor \U$69273 ( \69247 , \69245 , \69246 );
buf \U$69274 ( \69248 , \69247 );
buf \U$69275 ( \69249 , \69248 );
nand \U$69276 ( \69250 , \69244 , \69249 );
buf \U$69277 ( \69251 , \69250 );
buf \U$69278 ( \69252 , \69251 );
nand \U$69279 ( \69253 , \69243 , \69252 );
buf \U$69280 ( \69254 , \69253 );
buf \U$69281 ( \69255 , \69254 );
not \U$69282 ( \69256 , \69255 );
buf \U$69283 ( \69257 , \69256 );
buf \U$69284 ( \69258 , \69257 );
not \U$69285 ( \69259 , \69258 );
or \U$69286 ( \69260 , \69238 , \69259 );
buf \U$69287 ( \69261 , \69236 );
not \U$69288 ( \69262 , \69261 );
buf \U$69289 ( \69263 , \69254 );
nand \U$69290 ( \69264 , \69262 , \69263 );
buf \U$69291 ( \69265 , \69264 );
buf \U$69292 ( \69266 , \69265 );
nand \U$69293 ( \69267 , \69260 , \69266 );
buf \U$69294 ( \69268 , \69267 );
buf \U$69295 ( \69269 , \69268 );
buf \U$69296 ( \69270 , \68461 );
not \U$69297 ( \69271 , \69270 );
buf \U$69298 ( \69272 , \436 );
not \U$69299 ( \69273 , \69272 );
or \U$69300 ( \69274 , \69271 , \69273 );
buf \U$69301 ( \69275 , \442 );
xor \U$69302 ( \69276 , RIc0d9fb8_89, RIc0d8c08_47);
buf \U$69303 ( \69277 , \69276 );
nand \U$69304 ( \69278 , \69275 , \69277 );
buf \U$69305 ( \69279 , \69278 );
buf \U$69306 ( \69280 , \69279 );
nand \U$69307 ( \69281 , \69274 , \69280 );
buf \U$69308 ( \69282 , \69281 );
buf \U$69309 ( \69283 , \69282 );
xor \U$69310 ( \69284 , \69269 , \69283 );
buf \U$69311 ( \69285 , \69284 );
buf \U$69312 ( \69286 , \69285 );
not \U$69313 ( \69287 , \69286 );
or \U$69314 ( \69288 , \69224 , \69287 );
buf \U$69315 ( \69289 , \69222 );
buf \U$69316 ( \69290 , \69285 );
or \U$69317 ( \69291 , \69289 , \69290 );
nand \U$69318 ( \69292 , \69288 , \69291 );
buf \U$69319 ( \69293 , \69292 );
buf \U$69320 ( \69294 , \69293 );
buf \U$69321 ( \69295 , \67998 );
not \U$69322 ( \69296 , \69295 );
buf \U$69323 ( \69297 , \27743 );
not \U$69324 ( \69298 , \69297 );
or \U$69325 ( \69299 , \69296 , \69298 );
buf \U$69326 ( \69300 , \12303 );
buf \U$69327 ( \69301 , RIc0d7fd8_21);
buf \U$69328 ( \69302 , RIc0dabe8_115);
xor \U$69329 ( \69303 , \69301 , \69302 );
buf \U$69330 ( \69304 , \69303 );
buf \U$69331 ( \69305 , \69304 );
nand \U$69332 ( \69306 , \69300 , \69305 );
buf \U$69333 ( \69307 , \69306 );
buf \U$69334 ( \69308 , \69307 );
nand \U$69335 ( \69309 , \69299 , \69308 );
buf \U$69336 ( \69310 , \69309 );
buf \U$69337 ( \69311 , \69310 );
not \U$69338 ( \69312 , \69311 );
buf \U$69339 ( \69313 , \68431 );
not \U$69340 ( \69314 , \69313 );
buf \U$69341 ( \69315 , \13684 );
not \U$69342 ( \69316 , \69315 );
or \U$69343 ( \69317 , \69314 , \69316 );
buf \U$69344 ( \69318 , \12936 );
xor \U$69345 ( \69319 , RIc0dacd8_117, RIc0d7ee8_19);
buf \U$69346 ( \69320 , \69319 );
nand \U$69347 ( \69321 , \69318 , \69320 );
buf \U$69348 ( \69322 , \69321 );
buf \U$69349 ( \69323 , \69322 );
nand \U$69350 ( \69324 , \69317 , \69323 );
buf \U$69351 ( \69325 , \69324 );
buf \U$69352 ( \69326 , \69325 );
not \U$69353 ( \69327 , \69326 );
buf \U$69354 ( \69328 , \69327 );
buf \U$69355 ( \69329 , \69328 );
not \U$69356 ( \69330 , \69329 );
or \U$69357 ( \69331 , \69312 , \69330 );
buf \U$69358 ( \69332 , \69310 );
buf \U$69359 ( \69333 , \69328 );
or \U$69360 ( \69334 , \69332 , \69333 );
nand \U$69361 ( \69335 , \69331 , \69334 );
buf \U$69362 ( \69336 , \69335 );
buf \U$69363 ( \69337 , \69336 );
buf \U$69364 ( \69338 , \68196 );
not \U$69365 ( \69339 , \69338 );
buf \U$69366 ( \69340 , \4527 );
not \U$69367 ( \69341 , \69340 );
or \U$69368 ( \69342 , \69339 , \69341 );
buf \U$69369 ( \69343 , \14331 );
buf \U$69370 ( \69344 , RIc0d8cf8_49);
buf \U$69371 ( \69345 , RIc0d9ec8_87);
xor \U$69372 ( \69346 , \69344 , \69345 );
buf \U$69373 ( \69347 , \69346 );
buf \U$69374 ( \69348 , \69347 );
nand \U$69375 ( \69349 , \69343 , \69348 );
buf \U$69376 ( \69350 , \69349 );
buf \U$69377 ( \69351 , \69350 );
nand \U$69378 ( \69352 , \69342 , \69351 );
buf \U$69379 ( \69353 , \69352 );
buf \U$69380 ( \69354 , \69353 );
xor \U$69381 ( \69355 , \69337 , \69354 );
buf \U$69382 ( \69356 , \69355 );
buf \U$69383 ( \69357 , \69356 );
not \U$69384 ( \69358 , \69357 );
buf \U$69385 ( \69359 , \69358 );
buf \U$69386 ( \69360 , \69359 );
and \U$69387 ( \69361 , \69294 , \69360 );
not \U$69388 ( \69362 , \69294 );
buf \U$69389 ( \69363 , \69356 );
and \U$69390 ( \69364 , \69362 , \69363 );
nor \U$69391 ( \69365 , \69361 , \69364 );
buf \U$69392 ( \69366 , \69365 );
buf \U$69395 ( \69367 , \69366 );
buf \U$69396 ( \69368 , \69367 );
and \U$69397 ( \69369 , \69163 , \69368 );
not \U$69398 ( \69370 , \69163 );
buf \U$69399 ( \69371 , \69367 );
not \U$69400 ( \69372 , \69371 );
buf \U$69401 ( \69373 , \69372 );
buf \U$69402 ( \69374 , \69373 );
and \U$69403 ( \69375 , \69370 , \69374 );
nor \U$69404 ( \69376 , \69369 , \69375 );
buf \U$69405 ( \69377 , \69376 );
buf \U$69406 ( \69378 , \69377 );
not \U$69407 ( \69379 , \69378 );
buf \U$69408 ( \69380 , \69379 );
buf \U$69409 ( \69381 , \69380 );
not \U$69410 ( \69382 , \69381 );
buf \U$69411 ( \69383 , \66868 );
not \U$69412 ( \69384 , \69383 );
buf \U$69413 ( \69385 , \66852 );
not \U$69414 ( \69386 , \69385 );
or \U$69415 ( \69387 , \69384 , \69386 );
buf \U$69416 ( \69388 , \66852 );
buf \U$69417 ( \69389 , \66868 );
or \U$69418 ( \69390 , \69388 , \69389 );
buf \U$69419 ( \69391 , \66883 );
nand \U$69420 ( \69392 , \69390 , \69391 );
buf \U$69421 ( \69393 , \69392 );
buf \U$69422 ( \69394 , \69393 );
nand \U$69423 ( \69395 , \69387 , \69394 );
buf \U$69424 ( \69396 , \69395 );
buf \U$69425 ( \69397 , \69396 );
not \U$69426 ( \69398 , \69397 );
buf \U$69427 ( \69399 , \66966 );
not \U$69428 ( \69400 , \69399 );
buf \U$69429 ( \69401 , \66911 );
not \U$69430 ( \69402 , \69401 );
or \U$69431 ( \69403 , \69400 , \69402 );
buf \U$69432 ( \69404 , \66911 );
buf \U$69433 ( \69405 , \66966 );
or \U$69434 ( \69406 , \69404 , \69405 );
buf \U$69435 ( \69407 , \66932 );
nand \U$69436 ( \69408 , \69406 , \69407 );
buf \U$69437 ( \69409 , \69408 );
buf \U$69438 ( \69410 , \69409 );
nand \U$69439 ( \69411 , \69403 , \69410 );
buf \U$69440 ( \69412 , \69411 );
buf \U$69441 ( \69413 , \69412 );
not \U$69442 ( \69414 , \69413 );
or \U$69443 ( \69415 , \69398 , \69414 );
buf \U$69444 ( \69416 , \69412 );
buf \U$69445 ( \69417 , \69396 );
or \U$69446 ( \69418 , \69416 , \69417 );
buf \U$69447 ( \69419 , \68004 );
buf \U$69448 ( \69420 , \67987 );
xor \U$69449 ( \69421 , \69419 , \69420 );
buf \U$69450 ( \69422 , \68023 );
xnor \U$69451 ( \69423 , \69421 , \69422 );
buf \U$69452 ( \69424 , \69423 );
buf \U$69453 ( \69425 , \69424 );
not \U$69454 ( \69426 , \69425 );
buf \U$69455 ( \69427 , \67519 );
buf \U$69456 ( \69428 , \67551 );
buf \U$69457 ( \69429 , \67534 );
nor \U$69458 ( \69430 , \69428 , \69429 );
buf \U$69459 ( \69431 , \69430 );
buf \U$69460 ( \69432 , \69431 );
or \U$69461 ( \69433 , \69427 , \69432 );
buf \U$69462 ( \69434 , \67551 );
buf \U$69463 ( \69435 , \67534 );
nand \U$69464 ( \69436 , \69434 , \69435 );
buf \U$69465 ( \69437 , \69436 );
buf \U$69466 ( \69438 , \69437 );
nand \U$69467 ( \69439 , \69433 , \69438 );
buf \U$69468 ( \69440 , \69439 );
buf \U$69469 ( \69441 , \69440 );
not \U$69470 ( \69442 , \69441 );
buf \U$69471 ( \69443 , \69126 );
not \U$69472 ( \69444 , \69443 );
buf \U$69473 ( \69445 , \69111 );
not \U$69474 ( \69446 , \69445 );
or \U$69475 ( \69447 , \69444 , \69446 );
buf \U$69476 ( \69448 , \69126 );
buf \U$69477 ( \69449 , \69111 );
or \U$69478 ( \69450 , \69448 , \69449 );
nand \U$69479 ( \69451 , \69447 , \69450 );
buf \U$69480 ( \69452 , \69451 );
buf \U$69481 ( \69453 , \69452 );
not \U$69482 ( \69454 , \69453 );
buf \U$69483 ( \69455 , \69094 );
not \U$69484 ( \69456 , \69455 );
and \U$69485 ( \69457 , \69454 , \69456 );
buf \U$69486 ( \69458 , \69452 );
buf \U$69487 ( \69459 , \69094 );
and \U$69488 ( \69460 , \69458 , \69459 );
nor \U$69489 ( \69461 , \69457 , \69460 );
buf \U$69490 ( \69462 , \69461 );
buf \U$69491 ( \69463 , \69462 );
not \U$69492 ( \69464 , \69463 );
or \U$69493 ( \69465 , \69442 , \69464 );
buf \U$69494 ( \69466 , \69440 );
buf \U$69495 ( \69467 , \69462 );
or \U$69496 ( \69468 , \69466 , \69467 );
nand \U$69497 ( \69469 , \69465 , \69468 );
buf \U$69498 ( \69470 , \69469 );
buf \U$69499 ( \69471 , \69470 );
not \U$69500 ( \69472 , \69471 );
and \U$69501 ( \69473 , \69426 , \69472 );
buf \U$69502 ( \69474 , \69424 );
buf \U$69503 ( \69475 , \69470 );
and \U$69504 ( \69476 , \69474 , \69475 );
nor \U$69505 ( \69477 , \69473 , \69476 );
buf \U$69506 ( \69478 , \69477 );
buf \U$69507 ( \69479 , \69478 );
not \U$69508 ( \69480 , \69479 );
buf \U$69509 ( \69481 , \69480 );
buf \U$69510 ( \69482 , \69481 );
nand \U$69511 ( \69483 , \69418 , \69482 );
buf \U$69512 ( \69484 , \69483 );
buf \U$69513 ( \69485 , \69484 );
nand \U$69514 ( \69486 , \69415 , \69485 );
buf \U$69515 ( \69487 , \69486 );
buf \U$69516 ( \69488 , \69487 );
not \U$69517 ( \69489 , \69488 );
buf \U$69518 ( \69490 , \69489 );
buf \U$69519 ( \69491 , \69490 );
not \U$69520 ( \69492 , \69491 );
or \U$69521 ( \69493 , \69382 , \69492 );
buf \U$69522 ( \69494 , \69487 );
buf \U$69523 ( \69495 , \69377 );
nand \U$69524 ( \69496 , \69494 , \69495 );
buf \U$69525 ( \69497 , \69496 );
buf \U$69526 ( \69498 , \69497 );
nand \U$69527 ( \69499 , \69493 , \69498 );
buf \U$69528 ( \69500 , \69499 );
buf \U$69529 ( \69501 , \69500 );
buf \U$69530 ( \69502 , \68149 );
not \U$69531 ( \69503 , \69502 );
buf \U$69532 ( \69504 , \3415 );
not \U$69533 ( \69505 , \69504 );
or \U$69534 ( \69506 , \69503 , \69505 );
buf \U$69535 ( \69507 , \4008 );
buf \U$69536 ( \69508 , RIc0d8a28_43);
buf \U$69537 ( \69509 , RIc0da198_93);
xor \U$69538 ( \69510 , \69508 , \69509 );
buf \U$69539 ( \69511 , \69510 );
buf \U$69540 ( \69512 , \69511 );
nand \U$69541 ( \69513 , \69507 , \69512 );
buf \U$69542 ( \69514 , \69513 );
buf \U$69543 ( \69515 , \69514 );
nand \U$69544 ( \69516 , \69506 , \69515 );
buf \U$69545 ( \69517 , \69516 );
buf \U$69546 ( \69518 , \69517 );
buf \U$69547 ( \69519 , \68264 );
not \U$69548 ( \69520 , \69519 );
buf \U$69549 ( \69521 , \21898 );
not \U$69550 ( \69522 , \69521 );
or \U$69551 ( \69523 , \69520 , \69522 );
buf \U$69552 ( \69524 , \12342 );
buf \U$69553 ( \69525 , RIc0d8398_29);
buf \U$69554 ( \69526 , RIc0da828_107);
xor \U$69555 ( \69527 , \69525 , \69526 );
buf \U$69556 ( \69528 , \69527 );
buf \U$69557 ( \69529 , \69528 );
nand \U$69558 ( \69530 , \69524 , \69529 );
buf \U$69559 ( \69531 , \69530 );
buf \U$69560 ( \69532 , \69531 );
nand \U$69561 ( \69533 , \69523 , \69532 );
buf \U$69562 ( \69534 , \69533 );
buf \U$69563 ( \69535 , \69534 );
xor \U$69564 ( \69536 , \69518 , \69535 );
buf \U$69565 ( \69537 , \68134 );
not \U$69566 ( \69538 , \69537 );
buf \U$69567 ( \69539 , \13461 );
not \U$69568 ( \69540 , \69539 );
or \U$69569 ( \69541 , \69538 , \69540 );
buf \U$69570 ( \69542 , \13465 );
buf \U$69571 ( \69543 , RIc0d7b28_11);
buf \U$69572 ( \69544 , RIc0db098_125);
xor \U$69573 ( \69545 , \69543 , \69544 );
buf \U$69574 ( \69546 , \69545 );
buf \U$69575 ( \69547 , \69546 );
nand \U$69576 ( \69548 , \69542 , \69547 );
buf \U$69577 ( \69549 , \69548 );
buf \U$69578 ( \69550 , \69549 );
nand \U$69579 ( \69551 , \69541 , \69550 );
buf \U$69580 ( \69552 , \69551 );
buf \U$69581 ( \69553 , \69552 );
xor \U$69582 ( \69554 , \69536 , \69553 );
buf \U$69583 ( \69555 , \69554 );
buf \U$69584 ( \69556 , \68085 );
not \U$69585 ( \69557 , \69556 );
buf \U$69586 ( \69558 , \14100 );
not \U$69587 ( \69559 , \69558 );
or \U$69588 ( \69560 , \69557 , \69559 );
buf \U$69589 ( \69561 , \14352 );
buf \U$69590 ( \69562 , \20255 );
nand \U$69591 ( \69563 , \69561 , \69562 );
buf \U$69592 ( \69564 , \69563 );
buf \U$69593 ( \69565 , \69564 );
nand \U$69594 ( \69566 , \69560 , \69565 );
buf \U$69595 ( \69567 , \69566 );
buf \U$69596 ( \69568 , \69567 );
buf \U$69597 ( \69569 , \68410 );
not \U$69598 ( \69570 , \69569 );
buf \U$69599 ( \69571 , \4042 );
not \U$69600 ( \69572 , \69571 );
or \U$69601 ( \69573 , \69570 , \69572 );
buf \U$69602 ( \69574 , \3515 );
buf \U$69603 ( \69575 , RIc0d8668_35);
buf \U$69604 ( \69576 , RIc0da558_101);
xor \U$69605 ( \69577 , \69575 , \69576 );
buf \U$69606 ( \69578 , \69577 );
buf \U$69607 ( \69579 , \69578 );
nand \U$69608 ( \69580 , \69574 , \69579 );
buf \U$69609 ( \69581 , \69580 );
buf \U$69610 ( \69582 , \69581 );
nand \U$69611 ( \69583 , \69573 , \69582 );
buf \U$69612 ( \69584 , \69583 );
buf \U$69613 ( \69585 , \69584 );
xor \U$69614 ( \69586 , \69568 , \69585 );
buf \U$69615 ( \69587 , \68346 );
not \U$69616 ( \69588 , \69587 );
buf \U$69617 ( \69589 , \17405 );
not \U$69618 ( \69590 , \69589 );
or \U$69619 ( \69591 , \69588 , \69590 );
buf \U$69620 ( \69592 , \18416 );
buf \U$69621 ( \69593 , \20235 );
nand \U$69622 ( \69594 , \69592 , \69593 );
buf \U$69623 ( \69595 , \69594 );
buf \U$69624 ( \69596 , \69595 );
nand \U$69625 ( \69597 , \69591 , \69596 );
buf \U$69626 ( \69598 , \69597 );
buf \U$69627 ( \69599 , \69598 );
xor \U$69628 ( \69600 , \69586 , \69599 );
buf \U$69629 ( \69601 , \69600 );
xor \U$69630 ( \69602 , \69555 , \69601 );
buf \U$69631 ( \69603 , \68068 );
not \U$69632 ( \69604 , \69603 );
buf \U$69633 ( \69605 , \2088 );
not \U$69634 ( \69606 , \69605 );
or \U$69635 ( \69607 , \69604 , \69606 );
buf \U$69636 ( \69608 , \993 );
buf \U$69637 ( \69609 , \20131 );
nand \U$69638 ( \69610 , \69608 , \69609 );
buf \U$69639 ( \69611 , \69610 );
buf \U$69640 ( \69612 , \69611 );
nand \U$69641 ( \69613 , \69607 , \69612 );
buf \U$69642 ( \69614 , \69613 );
buf \U$69643 ( \69615 , \69614 );
not \U$69644 ( \69616 , \69615 );
buf \U$69645 ( \69617 , \69616 );
buf \U$69646 ( \69618 , \69617 );
not \U$69647 ( \69619 , \69618 );
buf \U$69648 ( \69620 , \68482 );
not \U$69649 ( \69621 , \69620 );
buf \U$69650 ( \69622 , \20098 );
not \U$69651 ( \69623 , \69622 );
or \U$69652 ( \69624 , \69621 , \69623 );
buf \U$69653 ( \69625 , \12975 );
buf \U$69654 ( \69626 , \20092 );
nand \U$69655 ( \69627 , \69625 , \69626 );
buf \U$69656 ( \69628 , \69627 );
buf \U$69657 ( \69629 , \69628 );
nand \U$69658 ( \69630 , \69624 , \69629 );
buf \U$69659 ( \69631 , \69630 );
buf \U$69660 ( \69632 , \69631 );
not \U$69661 ( \69633 , \69632 );
buf \U$69662 ( \69634 , \68447 );
not \U$69663 ( \69635 , \69634 );
buf \U$69664 ( \69636 , \13001 );
not \U$69665 ( \69637 , \69636 );
or \U$69666 ( \69638 , \69635 , \69637 );
buf \U$69667 ( \69639 , \13005 );
buf \U$69668 ( \69640 , RIc0d7df8_17);
buf \U$69669 ( \69641 , RIc0dadc8_119);
xor \U$69670 ( \69642 , \69640 , \69641 );
buf \U$69671 ( \69643 , \69642 );
buf \U$69672 ( \69644 , \69643 );
nand \U$69673 ( \69645 , \69639 , \69644 );
buf \U$69674 ( \69646 , \69645 );
buf \U$69675 ( \69647 , \69646 );
nand \U$69676 ( \69648 , \69638 , \69647 );
buf \U$69677 ( \69649 , \69648 );
buf \U$69678 ( \69650 , \69649 );
not \U$69679 ( \69651 , \69650 );
buf \U$69680 ( \69652 , \69651 );
buf \U$69681 ( \69653 , \69652 );
not \U$69682 ( \69654 , \69653 );
or \U$69683 ( \69655 , \69633 , \69654 );
buf \U$69684 ( \69656 , \69652 );
buf \U$69685 ( \69657 , \69631 );
or \U$69686 ( \69658 , \69656 , \69657 );
nand \U$69687 ( \69659 , \69655 , \69658 );
buf \U$69688 ( \69660 , \69659 );
buf \U$69689 ( \69661 , \69660 );
not \U$69690 ( \69662 , \69661 );
or \U$69691 ( \69663 , \69619 , \69662 );
buf \U$69692 ( \69664 , \69660 );
buf \U$69693 ( \69665 , \69617 );
or \U$69694 ( \69666 , \69664 , \69665 );
nand \U$69695 ( \69667 , \69663 , \69666 );
buf \U$69696 ( \69668 , \69667 );
xor \U$69697 ( \69669 , \69602 , \69668 );
buf \U$69698 ( \69670 , \69669 );
buf \U$69699 ( \69671 , \69440 );
not \U$69700 ( \69672 , \69671 );
buf \U$69701 ( \69673 , \69462 );
nand \U$69702 ( \69674 , \69672 , \69673 );
buf \U$69703 ( \69675 , \69674 );
buf \U$69704 ( \69676 , \69675 );
not \U$69705 ( \69677 , \69676 );
buf \U$69706 ( \69678 , \69424 );
not \U$69707 ( \69679 , \69678 );
buf \U$69708 ( \69680 , \69679 );
buf \U$69709 ( \69681 , \69680 );
not \U$69710 ( \69682 , \69681 );
or \U$69711 ( \69683 , \69677 , \69682 );
buf \U$69712 ( \69684 , \69462 );
not \U$69713 ( \69685 , \69684 );
buf \U$69714 ( \69686 , \69440 );
nand \U$69715 ( \69687 , \69685 , \69686 );
buf \U$69716 ( \69688 , \69687 );
buf \U$69717 ( \69689 , \69688 );
nand \U$69718 ( \69690 , \69683 , \69689 );
buf \U$69719 ( \69691 , \69690 );
buf \U$69720 ( \69692 , \69691 );
xor \U$69721 ( \69693 , \69670 , \69692 );
xor \U$69722 ( \69694 , \67812 , \67818 );
and \U$69723 ( \69695 , \69694 , \67825 );
and \U$69724 ( \69696 , \67812 , \67818 );
or \U$69725 ( \69697 , \69695 , \69696 );
buf \U$69726 ( \69698 , \69697 );
buf \U$69727 ( \69699 , \69698 );
xor \U$69728 ( \69700 , \69693 , \69699 );
buf \U$69729 ( \69701 , \69700 );
buf \U$69730 ( \69702 , \69701 );
not \U$69731 ( \69703 , \69702 );
buf \U$69732 ( \69704 , \69703 );
buf \U$69733 ( \69705 , \69704 );
and \U$69734 ( \69706 , \69501 , \69705 );
not \U$69735 ( \69707 , \69501 );
buf \U$69736 ( \69708 , \69701 );
and \U$69737 ( \69709 , \69707 , \69708 );
nor \U$69738 ( \69710 , \69706 , \69709 );
buf \U$69739 ( \69711 , \69710 );
buf \U$69740 ( \69712 , \69711 );
and \U$69741 ( \69713 , \68912 , \69712 );
not \U$69742 ( \69714 , \68912 );
buf \U$69743 ( \69715 , \69711 );
not \U$69744 ( \69716 , \69715 );
buf \U$69745 ( \69717 , \69716 );
buf \U$69746 ( \69718 , \69717 );
and \U$69747 ( \69719 , \69714 , \69718 );
nor \U$69748 ( \69720 , \69713 , \69719 );
buf \U$69749 ( \69721 , \69720 );
buf \U$69750 ( \69722 , \69721 );
buf \U$69753 ( \69723 , \69412 );
buf \U$69754 ( \69724 , \69723 );
not \U$69755 ( \69725 , \69724 );
buf \U$69756 ( \69726 , \69396 );
not \U$69757 ( \69727 , \69726 );
buf \U$69758 ( \69728 , \69478 );
not \U$69759 ( \69729 , \69728 );
and \U$69760 ( \69730 , \69727 , \69729 );
buf \U$69761 ( \69731 , \69396 );
buf \U$69762 ( \69732 , \69478 );
and \U$69763 ( \69733 , \69731 , \69732 );
nor \U$69764 ( \69734 , \69730 , \69733 );
buf \U$69765 ( \69735 , \69734 );
buf \U$69766 ( \69736 , \69735 );
not \U$69767 ( \69737 , \69736 );
or \U$69768 ( \69738 , \69725 , \69737 );
buf \U$69769 ( \69739 , \69735 );
buf \U$69770 ( \69740 , \69723 );
or \U$69771 ( \69741 , \69739 , \69740 );
nand \U$69772 ( \69742 , \69738 , \69741 );
buf \U$69773 ( \69743 , \69742 );
buf \U$69774 ( \69744 , \69743 );
xor \U$69775 ( \69745 , \66895 , \66968 );
and \U$69776 ( \69746 , \69745 , \66975 );
and \U$69777 ( \69747 , \66895 , \66968 );
or \U$69778 ( \69748 , \69746 , \69747 );
buf \U$69779 ( \69749 , \69748 );
buf \U$69780 ( \69750 , \69749 );
xor \U$69781 ( \69751 , \69744 , \69750 );
xor \U$69782 ( \69752 , \67828 , \67846 );
xor \U$69783 ( \69753 , \69752 , \67915 );
buf \U$69784 ( \69754 , \69753 );
buf \U$69785 ( \69755 , \69754 );
and \U$69786 ( \69756 , \69751 , \69755 );
and \U$69787 ( \69757 , \69744 , \69750 );
or \U$69788 ( \69758 , \69756 , \69757 );
buf \U$69789 ( \69759 , \69758 );
buf \U$69790 ( \69760 , \69759 );
and \U$69791 ( \69761 , \69722 , \69760 );
not \U$69792 ( \69762 , \69722 );
buf \U$69793 ( \69763 , \69759 );
not \U$69794 ( \69764 , \69763 );
buf \U$69795 ( \69765 , \69764 );
buf \U$69796 ( \69766 , \69765 );
and \U$69797 ( \69767 , \69762 , \69766 );
nor \U$69798 ( \69768 , \69761 , \69767 );
buf \U$69799 ( \69769 , \69768 );
buf \U$69800 ( \69770 , \69769 );
xor \U$69801 ( \69771 , \68892 , \69770 );
buf \U$69802 ( \69772 , \69771 );
buf \U$69803 ( \69773 , \69772 );
xor \U$69804 ( \69774 , \69744 , \69750 );
xor \U$69805 ( \69775 , \69774 , \69755 );
buf \U$69806 ( \69776 , \69775 );
buf \U$69807 ( \69777 , \69776 );
xor \U$69808 ( \69778 , \68811 , \68870 );
xor \U$69809 ( \69779 , \69778 , \68886 );
buf \U$69810 ( \69780 , \69779 );
buf \U$69811 ( \69781 , \69780 );
xor \U$69812 ( \69782 , \69777 , \69781 );
xor \U$69813 ( \69783 , \66992 , \67579 );
and \U$69814 ( \69784 , \69783 , \67586 );
and \U$69815 ( \69785 , \66992 , \67579 );
or \U$69816 ( \69786 , \69784 , \69785 );
buf \U$69817 ( \69787 , \69786 );
buf \U$69818 ( \69788 , \69787 );
and \U$69819 ( \69789 , \69782 , \69788 );
and \U$69820 ( \69790 , \69777 , \69781 );
or \U$69821 ( \69791 , \69789 , \69790 );
buf \U$69822 ( \69792 , \69791 );
buf \U$69823 ( \69793 , \69792 );
or \U$69824 ( \69794 , \69773 , \69793 );
buf \U$69825 ( \69795 , \69794 );
buf \U$69826 ( \69796 , \69795 );
xor \U$69827 ( \69797 , \69777 , \69781 );
xor \U$69828 ( \69798 , \69797 , \69788 );
buf \U$69829 ( \69799 , \69798 );
buf \U$69830 ( \69800 , \69799 );
not \U$69831 ( \69801 , \69800 );
buf \U$69832 ( \69802 , \69801 );
buf \U$69833 ( \69803 , \69802 );
xor \U$69834 ( \69804 , \66979 , \66985 );
and \U$69835 ( \69805 , \69804 , \67589 );
and \U$69836 ( \69806 , \66979 , \66985 );
or \U$69837 ( \69807 , \69805 , \69806 );
buf \U$69838 ( \69808 , \69807 );
buf \U$69839 ( \69809 , \69808 );
not \U$69840 ( \69810 , \69809 );
buf \U$69841 ( \69811 , \69810 );
buf \U$69842 ( \69812 , \69811 );
nand \U$69843 ( \69813 , \69803 , \69812 );
buf \U$69844 ( \69814 , \69813 );
buf \U$69845 ( \69815 , \69814 );
and \U$69846 ( \69816 , \69796 , \69815 );
buf \U$69847 ( \69817 , \69816 );
buf \U$69848 ( \69818 , \69817 );
buf \U$69849 ( \69819 , \67783 );
not \U$69850 ( \69820 , \69819 );
buf \U$69851 ( \69821 , \67797 );
not \U$69852 ( \69822 , \69821 );
buf \U$69853 ( \69823 , \69822 );
buf \U$69854 ( \69824 , \69823 );
not \U$69855 ( \69825 , \69824 );
or \U$69856 ( \69826 , \69820 , \69825 );
buf \U$69857 ( \69827 , \67783 );
not \U$69858 ( \69828 , \69827 );
buf \U$69859 ( \69829 , \67797 );
nand \U$69860 ( \69830 , \69828 , \69829 );
buf \U$69861 ( \69831 , \69830 );
buf \U$69862 ( \69832 , \69831 );
nand \U$69863 ( \69833 , \69826 , \69832 );
buf \U$69864 ( \69834 , \69833 );
buf \U$69865 ( \69835 , \69834 );
buf \U$69866 ( \69836 , \67792 );
and \U$69867 ( \69837 , \69835 , \69836 );
not \U$69868 ( \69838 , \69835 );
buf \U$69869 ( \69839 , \67779 );
and \U$69870 ( \69840 , \69838 , \69839 );
nor \U$69871 ( \69841 , \69837 , \69840 );
buf \U$69872 ( \69842 , \69841 );
buf \U$69873 ( \69843 , \69842 );
buf \U$69874 ( \69844 , \65564 );
buf \U$69875 ( \69845 , \65598 );
xnor \U$69876 ( \69846 , \69844 , \69845 );
buf \U$69877 ( \69847 , \69846 );
buf \U$69878 ( \69848 , \69847 );
buf \U$69879 ( \69849 , \65579 );
and \U$69880 ( \69850 , \69848 , \69849 );
not \U$69881 ( \69851 , \69848 );
buf \U$69882 ( \69852 , \65604 );
and \U$69883 ( \69853 , \69851 , \69852 );
nor \U$69884 ( \69854 , \69850 , \69853 );
buf \U$69885 ( \69855 , \69854 );
buf \U$69886 ( \69856 , \69855 );
xor \U$69887 ( \69857 , \67606 , \67621 );
xor \U$69888 ( \69858 , \69857 , \67635 );
buf \U$69889 ( \69859 , \69858 );
buf \U$69890 ( \69860 , \69859 );
xor \U$69891 ( \69861 , \69856 , \69860 );
buf \U$69892 ( \69862 , \67645 );
not \U$69893 ( \69863 , \69862 );
buf \U$69894 ( \69864 , \67678 );
not \U$69895 ( \69865 , \69864 );
buf \U$69896 ( \69866 , \67663 );
not \U$69897 ( \69867 , \69866 );
and \U$69898 ( \69868 , \69865 , \69867 );
buf \U$69899 ( \69869 , \67678 );
buf \U$69900 ( \69870 , \67663 );
and \U$69901 ( \69871 , \69869 , \69870 );
nor \U$69902 ( \69872 , \69868 , \69871 );
buf \U$69903 ( \69873 , \69872 );
buf \U$69904 ( \69874 , \69873 );
not \U$69905 ( \69875 , \69874 );
or \U$69906 ( \69876 , \69863 , \69875 );
buf \U$69907 ( \69877 , \69873 );
buf \U$69908 ( \69878 , \67645 );
or \U$69909 ( \69879 , \69877 , \69878 );
nand \U$69910 ( \69880 , \69876 , \69879 );
buf \U$69911 ( \69881 , \69880 );
buf \U$69912 ( \69882 , \69881 );
and \U$69913 ( \69883 , \69861 , \69882 );
and \U$69914 ( \69884 , \69856 , \69860 );
or \U$69915 ( \69885 , \69883 , \69884 );
buf \U$69916 ( \69886 , \69885 );
buf \U$69917 ( \69887 , \69886 );
xor \U$69918 ( \69888 , \67640 , \67683 );
xor \U$69919 ( \69889 , \69888 , \67688 );
buf \U$69920 ( \69890 , \69889 );
buf \U$69921 ( \69891 , \69890 );
xor \U$69922 ( \69892 , \69887 , \69891 );
xor \U$69923 ( \69893 , \53634 , \53856 );
and \U$69924 ( \69894 , \69893 , \54232 );
and \U$69925 ( \69895 , \53634 , \53856 );
or \U$69926 ( \69896 , \69894 , \69895 );
buf \U$69927 ( \69897 , \69896 );
buf \U$69928 ( \69898 , \69897 );
xor \U$69929 ( \69899 , \55418 , \55433 );
and \U$69930 ( \69900 , \69899 , \55449 );
and \U$69931 ( \69901 , \55418 , \55433 );
or \U$69932 ( \69902 , \69900 , \69901 );
buf \U$69933 ( \69903 , \69902 );
buf \U$69934 ( \69904 , \69903 );
xor \U$69935 ( \69905 , \69898 , \69904 );
buf \U$69936 ( \69906 , \67736 );
not \U$69937 ( \69907 , \69906 );
buf \U$69938 ( \69908 , \69907 );
buf \U$69939 ( \69909 , \69908 );
not \U$69940 ( \69910 , \69909 );
buf \U$69941 ( \69911 , \67723 );
not \U$69942 ( \69912 , \69911 );
buf \U$69943 ( \69913 , \67758 );
not \U$69944 ( \69914 , \69913 );
or \U$69945 ( \69915 , \69912 , \69914 );
buf \U$69946 ( \69916 , \67758 );
buf \U$69947 ( \69917 , \67723 );
or \U$69948 ( \69918 , \69916 , \69917 );
nand \U$69949 ( \69919 , \69915 , \69918 );
buf \U$69950 ( \69920 , \69919 );
buf \U$69951 ( \69921 , \69920 );
not \U$69952 ( \69922 , \69921 );
or \U$69953 ( \69923 , \69910 , \69922 );
buf \U$69954 ( \69924 , \69920 );
buf \U$69955 ( \69925 , \69908 );
or \U$69956 ( \69926 , \69924 , \69925 );
nand \U$69957 ( \69927 , \69923 , \69926 );
buf \U$69958 ( \69928 , \69927 );
buf \U$69959 ( \69929 , \69928 );
and \U$69960 ( \69930 , \69905 , \69929 );
and \U$69961 ( \69931 , \69898 , \69904 );
or \U$69962 ( \69932 , \69930 , \69931 );
buf \U$69963 ( \69933 , \69932 );
buf \U$69964 ( \69934 , \69933 );
and \U$69965 ( \69935 , \69892 , \69934 );
and \U$69966 ( \69936 , \69887 , \69891 );
or \U$69967 ( \69937 , \69935 , \69936 );
buf \U$69968 ( \69938 , \69937 );
buf \U$69969 ( \69939 , \69938 );
xor \U$69970 ( \69940 , \65548 , \65731 );
xor \U$69971 ( \69941 , \69940 , \65912 );
buf \U$69972 ( \69942 , \69941 );
buf \U$69973 ( \69943 , \69942 );
or \U$69974 ( \69944 , \69939 , \69943 );
xor \U$69975 ( \69945 , \67693 , \67697 );
xor \U$69976 ( \69946 , \69945 , \67775 );
buf \U$69977 ( \69947 , \69946 );
buf \U$69978 ( \69948 , \69947 );
nand \U$69979 ( \69949 , \69944 , \69948 );
buf \U$69980 ( \69950 , \69949 );
buf \U$69981 ( \69951 , \69950 );
buf \U$69982 ( \69952 , \69938 );
buf \U$69983 ( \69953 , \69942 );
nand \U$69984 ( \69954 , \69952 , \69953 );
buf \U$69985 ( \69955 , \69954 );
buf \U$69986 ( \69956 , \69955 );
and \U$69987 ( \69957 , \69951 , \69956 );
buf \U$69988 ( \69958 , \69957 );
buf \U$69989 ( \69959 , \69958 );
nand \U$69990 ( \69960 , \69843 , \69959 );
buf \U$69991 ( \69961 , \69960 );
buf \U$69992 ( \69962 , \69961 );
buf \U$69993 ( \69963 , \69942 );
buf \U$69994 ( \69964 , \69947 );
xor \U$69995 ( \69965 , \69963 , \69964 );
buf \U$69996 ( \69966 , \69938 );
xnor \U$69997 ( \69967 , \69965 , \69966 );
buf \U$69998 ( \69968 , \69967 );
buf \U$69999 ( \69969 , \69968 );
xor \U$70000 ( \69970 , \67702 , \67765 );
xor \U$70001 ( \69971 , \69970 , \67770 );
buf \U$70002 ( \69972 , \69971 );
buf \U$70003 ( \69973 , \69972 );
xor \U$70004 ( \69974 , \55775 , \55908 );
and \U$70005 ( \69975 , \69974 , \55985 );
and \U$70006 ( \69976 , \55775 , \55908 );
or \U$70007 ( \69977 , \69975 , \69976 );
buf \U$70008 ( \69978 , \69977 );
buf \U$70009 ( \69979 , \69978 );
xor \U$70010 ( \69980 , \54235 , \54637 );
and \U$70011 ( \69981 , \69980 , \55304 );
and \U$70012 ( \69982 , \54235 , \54637 );
or \U$70013 ( \69983 , \69981 , \69982 );
buf \U$70014 ( \69984 , \69983 );
buf \U$70015 ( \69985 , \69984 );
xor \U$70016 ( \69986 , \69979 , \69985 );
xor \U$70017 ( \69987 , \69856 , \69860 );
xor \U$70018 ( \69988 , \69987 , \69882 );
buf \U$70019 ( \69989 , \69988 );
buf \U$70020 ( \69990 , \69989 );
and \U$70021 ( \69991 , \69986 , \69990 );
and \U$70022 ( \69992 , \69979 , \69985 );
or \U$70023 ( \69993 , \69991 , \69992 );
buf \U$70024 ( \69994 , \69993 );
buf \U$70025 ( \69995 , \69994 );
xor \U$70026 ( \69996 , \69973 , \69995 );
xor \U$70027 ( \69997 , \69887 , \69891 );
xor \U$70028 ( \69998 , \69997 , \69934 );
buf \U$70029 ( \69999 , \69998 );
buf \U$70030 ( \70000 , \69999 );
and \U$70031 ( \70001 , \69996 , \70000 );
and \U$70032 ( \70002 , \69973 , \69995 );
or \U$70033 ( \70003 , \70001 , \70002 );
buf \U$70034 ( \70004 , \70003 );
buf \U$70035 ( \70005 , \70004 );
not \U$70036 ( \70006 , \70005 );
buf \U$70037 ( \70007 , \70006 );
buf \U$70038 ( \70008 , \70007 );
nand \U$70039 ( \70009 , \69969 , \70008 );
buf \U$70040 ( \70010 , \70009 );
buf \U$70041 ( \70011 , \70010 );
nand \U$70042 ( \70012 , \69962 , \70011 );
buf \U$70043 ( \70013 , \70012 );
buf \U$70044 ( \70014 , \70013 );
xor \U$70045 ( \70015 , \69898 , \69904 );
xor \U$70046 ( \70016 , \70015 , \69929 );
buf \U$70047 ( \70017 , \70016 );
buf \U$70048 ( \70018 , \70017 );
xor \U$70049 ( \70019 , \55452 , \55988 );
and \U$70050 ( \70020 , \70019 , \56167 );
and \U$70051 ( \70021 , \55452 , \55988 );
or \U$70052 ( \70022 , \70020 , \70021 );
buf \U$70053 ( \70023 , \70022 );
buf \U$70054 ( \70024 , \70023 );
xor \U$70055 ( \70025 , \70018 , \70024 );
xor \U$70056 ( \70026 , \69979 , \69985 );
xor \U$70057 ( \70027 , \70026 , \69990 );
buf \U$70058 ( \70028 , \70027 );
buf \U$70059 ( \70029 , \70028 );
and \U$70060 ( \70030 , \70025 , \70029 );
and \U$70061 ( \70031 , \70018 , \70024 );
or \U$70062 ( \70032 , \70030 , \70031 );
buf \U$70063 ( \70033 , \70032 );
buf \U$70064 ( \70034 , \70033 );
not \U$70065 ( \70035 , \70034 );
xor \U$70066 ( \70036 , \69973 , \69995 );
xor \U$70067 ( \70037 , \70036 , \70000 );
buf \U$70068 ( \70038 , \70037 );
buf \U$70069 ( \70039 , \70038 );
not \U$70070 ( \70040 , \70039 );
buf \U$70071 ( \70041 , \70040 );
buf \U$70072 ( \70042 , \70041 );
nand \U$70073 ( \70043 , \70035 , \70042 );
buf \U$70074 ( \70044 , \70043 );
buf \U$70075 ( \70045 , \70044 );
xor \U$70076 ( \70046 , \70018 , \70024 );
xor \U$70077 ( \70047 , \70046 , \70029 );
buf \U$70078 ( \70048 , \70047 );
buf \U$70079 ( \70049 , \70048 );
xor \U$70080 ( \70050 , \55307 , \56170 );
and \U$70081 ( \70051 , \70050 , \56208 );
and \U$70082 ( \70052 , \55307 , \56170 );
or \U$70083 ( \70053 , \70051 , \70052 );
buf \U$70084 ( \70054 , \70053 );
buf \U$70085 ( \70055 , \70054 );
or \U$70086 ( \70056 , \70049 , \70055 );
buf \U$70087 ( \70057 , \70056 );
buf \U$70088 ( \70058 , \70057 );
nand \U$70089 ( \70059 , \70045 , \70058 );
buf \U$70090 ( \70060 , \70059 );
buf \U$70091 ( \70061 , \70060 );
nor \U$70092 ( \70062 , \70014 , \70061 );
buf \U$70093 ( \70063 , \70062 );
buf \U$70094 ( \70064 , \70063 );
and \U$70095 ( \70065 , \67806 , \69818 , \70064 );
buf \U$70096 ( \70066 , \70065 );
buf \U$70097 ( \70067 , \70066 );
buf \U$70098 ( \70068 , \20171 );
buf \U$70099 ( \70069 , \20218 );
xor \U$70100 ( \70070 , \70068 , \70069 );
buf \U$70101 ( \70071 , \20198 );
xor \U$70102 ( \70072 , \70070 , \70071 );
buf \U$70103 ( \70073 , \70072 );
buf \U$70104 ( \70074 , \70073 );
not \U$70105 ( \70075 , \70074 );
buf \U$70106 ( \70076 , \69578 );
not \U$70107 ( \70077 , \70076 );
buf \U$70108 ( \70078 , \20798 );
not \U$70109 ( \70079 , \70078 );
or \U$70110 ( \70080 , \70077 , \70079 );
buf \U$70111 ( \70081 , \15550 );
buf \U$70112 ( \70082 , \19935 );
nand \U$70113 ( \70083 , \70081 , \70082 );
buf \U$70114 ( \70084 , \70083 );
buf \U$70115 ( \70085 , \70084 );
nand \U$70116 ( \70086 , \70080 , \70085 );
buf \U$70117 ( \70087 , \70086 );
buf \U$70118 ( \70088 , \69248 );
not \U$70119 ( \70089 , \70088 );
buf \U$70120 ( \70090 , \12870 );
not \U$70121 ( \70091 , \70090 );
or \U$70122 ( \70092 , \70089 , \70091 );
buf \U$70123 ( \70093 , \12877 );
buf \U$70124 ( \70094 , \19353 );
nand \U$70125 ( \70095 , \70093 , \70094 );
buf \U$70126 ( \70096 , \70095 );
buf \U$70127 ( \70097 , \70096 );
nand \U$70128 ( \70098 , \70092 , \70097 );
buf \U$70129 ( \70099 , \70098 );
xnor \U$70130 ( \70100 , \70087 , \70099 );
buf \U$70131 ( \70101 , \69276 );
not \U$70132 ( \70102 , \70101 );
buf \U$70133 ( \70103 , \436 );
not \U$70134 ( \70104 , \70103 );
or \U$70135 ( \70105 , \70102 , \70104 );
buf \U$70136 ( \70106 , \442 );
buf \U$70137 ( \70107 , \18145 );
nand \U$70138 ( \70108 , \70106 , \70107 );
buf \U$70139 ( \70109 , \70108 );
buf \U$70140 ( \70110 , \70109 );
nand \U$70141 ( \70111 , \70105 , \70110 );
buf \U$70142 ( \70112 , \70111 );
and \U$70143 ( \70113 , \70100 , \70112 );
not \U$70144 ( \70114 , \70100 );
buf \U$70145 ( \70115 , \70112 );
not \U$70146 ( \70116 , \70115 );
buf \U$70147 ( \70117 , \70116 );
and \U$70148 ( \70118 , \70114 , \70117 );
nor \U$70149 ( \70119 , \70113 , \70118 );
buf \U$70150 ( \70120 , \70119 );
not \U$70151 ( \70121 , \70120 );
buf \U$70152 ( \70122 , \70121 );
buf \U$70153 ( \70123 , \70122 );
not \U$70154 ( \70124 , \70123 );
or \U$70155 ( \70125 , \70075 , \70124 );
buf \U$70156 ( \70126 , \70073 );
not \U$70157 ( \70127 , \70126 );
buf \U$70158 ( \70128 , \70127 );
buf \U$70159 ( \70129 , \70128 );
buf \U$70160 ( \70130 , \70119 );
nand \U$70161 ( \70131 , \70129 , \70130 );
buf \U$70162 ( \70132 , \70131 );
buf \U$70163 ( \70133 , \70132 );
nand \U$70164 ( \70134 , \70125 , \70133 );
buf \U$70165 ( \70135 , \70134 );
buf \U$70166 ( \70136 , \70135 );
buf \U$70167 ( \70137 , \69347 );
not \U$70168 ( \70138 , \70137 );
buf \U$70169 ( \70139 , \2607 );
not \U$70170 ( \70140 , \70139 );
or \U$70171 ( \70141 , \70138 , \70140 );
buf \U$70172 ( \70142 , \816 );
buf \U$70173 ( \70143 , \19439 );
nand \U$70174 ( \70144 , \70142 , \70143 );
buf \U$70175 ( \70145 , \70144 );
buf \U$70176 ( \70146 , \70145 );
nand \U$70177 ( \70147 , \70141 , \70146 );
buf \U$70178 ( \70148 , \70147 );
buf \U$70179 ( \70149 , \70148 );
not \U$70180 ( \70150 , \70149 );
buf \U$70181 ( \70151 , \70150 );
buf \U$70182 ( \70152 , \70151 );
not \U$70183 ( \70153 , \70152 );
buf \U$70184 ( \70154 , \69319 );
not \U$70185 ( \70155 , \70154 );
buf \U$70186 ( \70156 , \13684 );
not \U$70187 ( \70157 , \70156 );
or \U$70188 ( \70158 , \70155 , \70157 );
buf \U$70189 ( \70159 , \12937 );
buf \U$70190 ( \70160 , \19331 );
nand \U$70191 ( \70161 , \70159 , \70160 );
buf \U$70192 ( \70162 , \70161 );
buf \U$70193 ( \70163 , \70162 );
nand \U$70194 ( \70164 , \70158 , \70163 );
buf \U$70195 ( \70165 , \70164 );
buf \U$70196 ( \70166 , \70165 );
not \U$70197 ( \70167 , \70166 );
buf \U$70198 ( \70168 , \69546 );
not \U$70199 ( \70169 , \70168 );
buf \U$70200 ( \70170 , \16914 );
not \U$70201 ( \70171 , \70170 );
or \U$70202 ( \70172 , \70169 , \70171 );
buf \U$70203 ( \70173 , \15793 );
buf \U$70204 ( \70174 , \19523 );
nand \U$70205 ( \70175 , \70173 , \70174 );
buf \U$70206 ( \70176 , \70175 );
buf \U$70207 ( \70177 , \70176 );
nand \U$70208 ( \70178 , \70172 , \70177 );
buf \U$70209 ( \70179 , \70178 );
buf \U$70210 ( \70180 , \70179 );
not \U$70211 ( \70181 , \70180 );
buf \U$70212 ( \70182 , \70181 );
buf \U$70213 ( \70183 , \70182 );
not \U$70214 ( \70184 , \70183 );
or \U$70215 ( \70185 , \70167 , \70184 );
buf \U$70216 ( \70186 , \70165 );
buf \U$70217 ( \70187 , \70182 );
or \U$70218 ( \70188 , \70186 , \70187 );
nand \U$70219 ( \70189 , \70185 , \70188 );
buf \U$70220 ( \70190 , \70189 );
buf \U$70221 ( \70191 , \70190 );
not \U$70222 ( \70192 , \70191 );
or \U$70223 ( \70193 , \70153 , \70192 );
buf \U$70224 ( \70194 , \70190 );
buf \U$70225 ( \70195 , \70151 );
or \U$70226 ( \70196 , \70194 , \70195 );
nand \U$70227 ( \70197 , \70193 , \70196 );
buf \U$70228 ( \70198 , \70197 );
buf \U$70229 ( \70199 , \70198 );
xnor \U$70230 ( \70200 , \70136 , \70199 );
buf \U$70231 ( \70201 , \70200 );
buf \U$70232 ( \70202 , \70201 );
not \U$70233 ( \70203 , \70202 );
buf \U$70234 ( \70204 , \20125 );
buf \U$70235 ( \70205 , \20108 );
xor \U$70236 ( \70206 , \70204 , \70205 );
buf \U$70237 ( \70207 , \20143 );
xor \U$70238 ( \70208 , \70206 , \70207 );
buf \U$70239 ( \70209 , \70208 );
buf \U$70240 ( \70210 , \69528 );
not \U$70241 ( \70211 , \70210 );
buf \U$70242 ( \70212 , \16065 );
not \U$70243 ( \70213 , \70212 );
or \U$70244 ( \70214 , \70211 , \70213 );
buf \U$70245 ( \70215 , \16071 );
buf \U$70246 ( \70216 , \19409 );
nand \U$70247 ( \70217 , \70215 , \70216 );
buf \U$70248 ( \70218 , \70217 );
buf \U$70249 ( \70219 , \70218 );
nand \U$70250 ( \70220 , \70214 , \70219 );
buf \U$70251 ( \70221 , \70220 );
buf \U$70252 ( \70222 , \70221 );
not \U$70253 ( \70223 , \70222 );
buf \U$70254 ( \70224 , \69511 );
not \U$70255 ( \70225 , \70224 );
buf \U$70256 ( \70226 , \15995 );
not \U$70257 ( \70227 , \70226 );
or \U$70258 ( \70228 , \70225 , \70227 );
buf \U$70259 ( \70229 , \481 );
buf \U$70260 ( \70230 , \19460 );
nand \U$70261 ( \70231 , \70229 , \70230 );
buf \U$70262 ( \70232 , \70231 );
buf \U$70263 ( \70233 , \70232 );
nand \U$70264 ( \70234 , \70228 , \70233 );
buf \U$70265 ( \70235 , \70234 );
buf \U$70266 ( \70236 , \70235 );
not \U$70267 ( \70237 , \70236 );
buf \U$70268 ( \70238 , \70237 );
buf \U$70269 ( \70239 , \70238 );
not \U$70270 ( \70240 , \70239 );
or \U$70271 ( \70241 , \70223 , \70240 );
buf \U$70272 ( \70242 , \70235 );
buf \U$70273 ( \70243 , \70221 );
not \U$70274 ( \70244 , \70243 );
buf \U$70275 ( \70245 , \70244 );
buf \U$70276 ( \70246 , \70245 );
nand \U$70277 ( \70247 , \70242 , \70246 );
buf \U$70278 ( \70248 , \70247 );
buf \U$70279 ( \70249 , \70248 );
nand \U$70280 ( \70250 , \70241 , \70249 );
buf \U$70281 ( \70251 , \70250 );
buf \U$70282 ( \70252 , \70251 );
buf \U$70283 ( \70253 , \69643 );
not \U$70284 ( \70254 , \70253 );
buf \U$70285 ( \70255 , \13949 );
not \U$70286 ( \70256 , \70255 );
or \U$70287 ( \70257 , \70254 , \70256 );
buf \U$70288 ( \70258 , \13005 );
buf \U$70289 ( \70259 , \19560 );
nand \U$70290 ( \70260 , \70258 , \70259 );
buf \U$70291 ( \70261 , \70260 );
buf \U$70292 ( \70262 , \70261 );
nand \U$70293 ( \70263 , \70257 , \70262 );
buf \U$70294 ( \70264 , \70263 );
buf \U$70295 ( \70265 , \70264 );
not \U$70296 ( \70266 , \70265 );
buf \U$70297 ( \70267 , \70266 );
buf \U$70298 ( \70268 , \70267 );
and \U$70299 ( \70269 , \70252 , \70268 );
not \U$70300 ( \70270 , \70252 );
buf \U$70301 ( \70271 , \70264 );
and \U$70302 ( \70272 , \70270 , \70271 );
nor \U$70303 ( \70273 , \70269 , \70272 );
buf \U$70304 ( \70274 , \70273 );
xor \U$70305 ( \70275 , \70209 , \70274 );
xor \U$70306 ( \70276 , \20251 , \20268 );
xor \U$70307 ( \70277 , \70276 , \20286 );
buf \U$70308 ( \70278 , \70277 );
xor \U$70309 ( \70279 , \70275 , \70278 );
buf \U$70310 ( \70280 , \70279 );
not \U$70311 ( \70281 , \70280 );
or \U$70312 ( \70282 , \70203 , \70281 );
buf \U$70313 ( \70283 , \67978 );
not \U$70314 ( \70284 , \70283 );
buf \U$70315 ( \70285 , \67956 );
not \U$70316 ( \70286 , \70285 );
or \U$70317 ( \70287 , \70284 , \70286 );
buf \U$70318 ( \70288 , \67956 );
buf \U$70319 ( \70289 , \67978 );
or \U$70320 ( \70290 , \70288 , \70289 );
buf \U$70321 ( \70291 , \67942 );
nand \U$70322 ( \70292 , \70290 , \70291 );
buf \U$70323 ( \70293 , \70292 );
buf \U$70324 ( \70294 , \70293 );
nand \U$70325 ( \70295 , \70287 , \70294 );
buf \U$70326 ( \70296 , \70295 );
buf \U$70327 ( \70297 , \70296 );
not \U$70328 ( \70298 , \70297 );
xor \U$70329 ( \70299 , \69568 , \69585 );
and \U$70330 ( \70300 , \70299 , \69599 );
and \U$70331 ( \70301 , \69568 , \69585 );
or \U$70332 ( \70302 , \70300 , \70301 );
buf \U$70333 ( \70303 , \70302 );
buf \U$70334 ( \70304 , \70303 );
not \U$70335 ( \70305 , \70304 );
buf \U$70336 ( \70306 , \70305 );
buf \U$70337 ( \70307 , \70306 );
not \U$70338 ( \70308 , \70307 );
or \U$70339 ( \70309 , \70298 , \70308 );
buf \U$70340 ( \70310 , \70306 );
buf \U$70341 ( \70311 , \70296 );
or \U$70342 ( \70312 , \70310 , \70311 );
nand \U$70343 ( \70313 , \70309 , \70312 );
buf \U$70344 ( \70314 , \70313 );
buf \U$70345 ( \70315 , \70314 );
xor \U$70346 ( \70316 , \68951 , \68966 );
and \U$70347 ( \70317 , \70316 , \68980 );
and \U$70348 ( \70318 , \68951 , \68966 );
or \U$70349 ( \70319 , \70317 , \70318 );
buf \U$70350 ( \70320 , \70319 );
buf \U$70351 ( \70321 , \70320 );
and \U$70352 ( \70322 , \70315 , \70321 );
not \U$70353 ( \70323 , \70315 );
buf \U$70354 ( \70324 , \70320 );
not \U$70355 ( \70325 , \70324 );
buf \U$70356 ( \70326 , \70325 );
buf \U$70357 ( \70327 , \70326 );
and \U$70358 ( \70328 , \70323 , \70327 );
nor \U$70359 ( \70329 , \70322 , \70328 );
buf \U$70360 ( \70330 , \70329 );
buf \U$70361 ( \70331 , \70330 );
nand \U$70362 ( \70332 , \70282 , \70331 );
buf \U$70363 ( \70333 , \70332 );
buf \U$70364 ( \70334 , \70333 );
buf \U$70365 ( \70335 , \70201 );
not \U$70366 ( \70336 , \70335 );
buf \U$70367 ( \70337 , \70279 );
not \U$70368 ( \70338 , \70337 );
buf \U$70369 ( \70339 , \70338 );
buf \U$70370 ( \70340 , \70339 );
nand \U$70371 ( \70341 , \70336 , \70340 );
buf \U$70372 ( \70342 , \70341 );
buf \U$70373 ( \70343 , \70342 );
nand \U$70374 ( \70344 , \70334 , \70343 );
buf \U$70375 ( \70345 , \70344 );
buf \U$70376 ( \70346 , \70345 );
buf \U$70377 ( \70347 , \69033 );
not \U$70378 ( \70348 , \70347 );
buf \U$70379 ( \70349 , \69027 );
not \U$70380 ( \70350 , \70349 );
or \U$70381 ( \70351 , \70348 , \70350 );
buf \U$70382 ( \70352 , \69053 );
nand \U$70383 ( \70353 , \70351 , \70352 );
buf \U$70384 ( \70354 , \70353 );
buf \U$70385 ( \70355 , \70354 );
buf \U$70386 ( \70356 , \69024 );
buf \U$70387 ( \70357 , \69007 );
nand \U$70388 ( \70358 , \70356 , \70357 );
buf \U$70389 ( \70359 , \70358 );
buf \U$70390 ( \70360 , \70359 );
nand \U$70391 ( \70361 , \70355 , \70360 );
buf \U$70392 ( \70362 , \70361 );
buf \U$70393 ( \70363 , \70362 );
buf \U$70394 ( \70364 , \69353 );
not \U$70395 ( \70365 , \70364 );
buf \U$70396 ( \70366 , \70365 );
buf \U$70397 ( \70367 , \70366 );
not \U$70398 ( \70368 , \70367 );
buf \U$70399 ( \70369 , \69328 );
not \U$70400 ( \70370 , \70369 );
or \U$70401 ( \70371 , \70368 , \70370 );
buf \U$70402 ( \70372 , \69310 );
nand \U$70403 ( \70373 , \70371 , \70372 );
buf \U$70404 ( \70374 , \70373 );
buf \U$70405 ( \70375 , \70374 );
buf \U$70406 ( \70376 , \69325 );
buf \U$70407 ( \70377 , \69353 );
nand \U$70408 ( \70378 , \70376 , \70377 );
buf \U$70409 ( \70379 , \70378 );
buf \U$70410 ( \70380 , \70379 );
nand \U$70411 ( \70381 , \70375 , \70380 );
buf \U$70412 ( \70382 , \70381 );
buf \U$70413 ( \70383 , \70382 );
xor \U$70414 ( \70384 , \70363 , \70383 );
xor \U$70415 ( \70385 , \69518 , \69535 );
and \U$70416 ( \70386 , \70385 , \69553 );
and \U$70417 ( \70387 , \69518 , \69535 );
or \U$70418 ( \70388 , \70386 , \70387 );
buf \U$70419 ( \70389 , \70388 );
buf \U$70420 ( \70390 , \70389 );
and \U$70421 ( \70391 , \70384 , \70390 );
and \U$70422 ( \70392 , \70363 , \70383 );
or \U$70423 ( \70393 , \70391 , \70392 );
buf \U$70424 ( \70394 , \70393 );
buf \U$70425 ( \70395 , \70394 );
xor \U$70426 ( \70396 , \20155 , \20230 );
xor \U$70427 ( \70397 , \70396 , \20291 );
buf \U$70428 ( \70398 , \70397 );
buf \U$70429 ( \70399 , \70398 );
xor \U$70430 ( \70400 , \70395 , \70399 );
not \U$70431 ( \70401 , \70235 );
not \U$70432 ( \70402 , \70221 );
or \U$70433 ( \70403 , \70401 , \70402 );
not \U$70434 ( \70404 , \70245 );
not \U$70435 ( \70405 , \70238 );
or \U$70436 ( \70406 , \70404 , \70405 );
nand \U$70437 ( \70407 , \70406 , \70264 );
nand \U$70438 ( \70408 , \70403 , \70407 );
buf \U$70439 ( \70409 , \70408 );
buf \U$70440 ( \70410 , \70165 );
buf \U$70441 ( \70411 , \70148 );
nor \U$70442 ( \70412 , \70410 , \70411 );
buf \U$70443 ( \70413 , \70412 );
buf \U$70444 ( \70414 , \70413 );
buf \U$70445 ( \70415 , \70182 );
or \U$70446 ( \70416 , \70414 , \70415 );
buf \U$70447 ( \70417 , \70165 );
buf \U$70448 ( \70418 , \70148 );
nand \U$70449 ( \70419 , \70417 , \70418 );
buf \U$70450 ( \70420 , \70419 );
buf \U$70451 ( \70421 , \70420 );
nand \U$70452 ( \70422 , \70416 , \70421 );
buf \U$70453 ( \70423 , \70422 );
buf \U$70454 ( \70424 , \70423 );
xor \U$70455 ( \70425 , \70409 , \70424 );
buf \U$70456 ( \70426 , \69047 );
not \U$70457 ( \70427 , \70426 );
buf \U$70458 ( \70428 , \16402 );
not \U$70459 ( \70429 , \70428 );
or \U$70460 ( \70430 , \70427 , \70429 );
buf \U$70461 ( \70431 , \1933 );
buf \U$70462 ( \70432 , \19599 );
nand \U$70463 ( \70433 , \70431 , \70432 );
buf \U$70464 ( \70434 , \70433 );
buf \U$70465 ( \70435 , \70434 );
nand \U$70466 ( \70436 , \70430 , \70435 );
buf \U$70467 ( \70437 , \70436 );
buf \U$70468 ( \70438 , \70437 );
not \U$70469 ( \70439 , \70438 );
buf \U$70470 ( \70440 , \70439 );
buf \U$70471 ( \70441 , \70440 );
not \U$70472 ( \70442 , \70441 );
buf \U$70473 ( \70443 , \69018 );
not \U$70474 ( \70444 , \70443 );
buf \U$70475 ( \70445 , \1183 );
not \U$70476 ( \70446 , \70445 );
or \U$70477 ( \70447 , \70444 , \70446 );
buf \U$70478 ( \70448 , \27267 );
buf \U$70479 ( \70449 , \18095 );
nand \U$70480 ( \70450 , \70448 , \70449 );
buf \U$70481 ( \70451 , \70450 );
buf \U$70482 ( \70452 , \70451 );
nand \U$70483 ( \70453 , \70447 , \70452 );
buf \U$70484 ( \70454 , \70453 );
buf \U$70485 ( \70455 , \70454 );
not \U$70486 ( \70456 , \70455 );
buf \U$70487 ( \70457 , \70456 );
buf \U$70488 ( \70458 , \70457 );
not \U$70489 ( \70459 , \70458 );
or \U$70490 ( \70460 , \70442 , \70459 );
buf \U$70491 ( \70461 , \69304 );
not \U$70492 ( \70462 , \70461 );
buf \U$70493 ( \70463 , \12299 );
not \U$70494 ( \70464 , \70463 );
or \U$70495 ( \70465 , \70462 , \70464 );
buf \U$70496 ( \70466 , \12303 );
buf \U$70497 ( \70467 , \19581 );
nand \U$70498 ( \70468 , \70466 , \70467 );
buf \U$70499 ( \70469 , \70468 );
buf \U$70500 ( \70470 , \70469 );
nand \U$70501 ( \70471 , \70465 , \70470 );
buf \U$70502 ( \70472 , \70471 );
buf \U$70503 ( \70473 , \70472 );
nand \U$70504 ( \70474 , \70460 , \70473 );
buf \U$70505 ( \70475 , \70474 );
buf \U$70506 ( \70476 , \70475 );
buf \U$70507 ( \70477 , \70440 );
not \U$70508 ( \70478 , \70477 );
buf \U$70509 ( \70479 , \70454 );
nand \U$70510 ( \70480 , \70478 , \70479 );
buf \U$70511 ( \70481 , \70480 );
buf \U$70512 ( \70482 , \70481 );
nand \U$70513 ( \70483 , \70476 , \70482 );
buf \U$70514 ( \70484 , \70483 );
buf \U$70515 ( \70485 , \70484 );
xor \U$70516 ( \70486 , \70425 , \70485 );
buf \U$70517 ( \70487 , \70486 );
buf \U$70518 ( \70488 , \70487 );
xor \U$70519 ( \70489 , \70400 , \70488 );
buf \U$70520 ( \70490 , \70489 );
buf \U$70521 ( \70491 , \70490 );
xor \U$70522 ( \70492 , \70346 , \70491 );
buf \U$70523 ( \70493 , \70274 );
not \U$70524 ( \70494 , \70493 );
buf \U$70525 ( \70495 , \70494 );
buf \U$70526 ( \70496 , \70495 );
buf \U$70527 ( \70497 , \70209 );
or \U$70528 ( \70498 , \70496 , \70497 );
buf \U$70529 ( \70499 , \70278 );
nand \U$70530 ( \70500 , \70498 , \70499 );
buf \U$70531 ( \70501 , \70500 );
buf \U$70532 ( \70502 , \70501 );
buf \U$70533 ( \70503 , \70209 );
buf \U$70534 ( \70504 , \70495 );
nand \U$70535 ( \70505 , \70503 , \70504 );
buf \U$70536 ( \70506 , \70505 );
buf \U$70537 ( \70507 , \70506 );
nand \U$70538 ( \70508 , \70502 , \70507 );
buf \U$70539 ( \70509 , \70508 );
buf \U$70540 ( \70510 , \70509 );
xor \U$70541 ( \70511 , \19536 , \19555 );
xor \U$70542 ( \70512 , \70511 , \19573 );
buf \U$70543 ( \70513 , \70512 );
buf \U$70544 ( \70514 , \70513 );
buf \U$70545 ( \70515 , \68682 );
not \U$70546 ( \70516 , \70515 );
buf \U$70547 ( \70517 , \68699 );
nor \U$70548 ( \70518 , \70516 , \70517 );
buf \U$70549 ( \70519 , \70518 );
buf \U$70550 ( \70520 , \70519 );
not \U$70551 ( \70521 , \70520 );
buf \U$70552 ( \70522 , \14888 );
not \U$70553 ( \70523 , \70522 );
buf \U$70554 ( \70524 , \68959 );
not \U$70555 ( \70525 , \70524 );
buf \U$70556 ( \70526 , \70525 );
buf \U$70557 ( \70527 , \70526 );
not \U$70558 ( \70528 , \70527 );
and \U$70559 ( \70529 , \70523 , \70528 );
buf \U$70560 ( \70530 , \19671 );
not \U$70561 ( \70531 , \70530 );
buf \U$70562 ( \70532 , \34244 );
nor \U$70563 ( \70533 , \70531 , \70532 );
buf \U$70564 ( \70534 , \70533 );
buf \U$70565 ( \70535 , \70534 );
nor \U$70566 ( \70536 , \70529 , \70535 );
buf \U$70567 ( \70537 , \70536 );
buf \U$70568 ( \70538 , \70537 );
buf \U$70569 ( \70539 , \18008 );
not \U$70570 ( \70540 , \70539 );
buf \U$70571 ( \70541 , \68943 );
not \U$70572 ( \70542 , \70541 );
buf \U$70573 ( \70543 , \70542 );
buf \U$70574 ( \70544 , \70543 );
not \U$70575 ( \70545 , \70544 );
and \U$70576 ( \70546 , \70540 , \70545 );
buf \U$70577 ( \70547 , RIc0d79c0_8);
buf \U$70578 ( \70548 , RIc0db188_127);
xor \U$70579 ( \70549 , \70547 , \70548 );
buf \U$70580 ( \70550 , \70549 );
buf \U$70581 ( \70551 , \70550 );
buf \U$70582 ( \70552 , RIc0db200_128);
and \U$70583 ( \70553 , \70551 , \70552 );
nor \U$70584 ( \70554 , \70546 , \70553 );
buf \U$70585 ( \70555 , \70554 );
buf \U$70586 ( \70556 , \70555 );
nand \U$70587 ( \70557 , \70538 , \70556 );
buf \U$70588 ( \70558 , \70557 );
buf \U$70589 ( \70559 , \70558 );
not \U$70590 ( \70560 , \70559 );
or \U$70591 ( \70561 , \70521 , \70560 );
buf \U$70592 ( \70562 , \70537 );
not \U$70593 ( \70563 , \70562 );
buf \U$70594 ( \70564 , \70563 );
buf \U$70595 ( \70565 , \70564 );
buf \U$70596 ( \70566 , \70555 );
not \U$70597 ( \70567 , \70566 );
buf \U$70598 ( \70568 , \70567 );
buf \U$70599 ( \70569 , \70568 );
nand \U$70600 ( \70570 , \70565 , \70569 );
buf \U$70601 ( \70571 , \70570 );
buf \U$70602 ( \70572 , \70571 );
nand \U$70603 ( \70573 , \70561 , \70572 );
buf \U$70604 ( \70574 , \70573 );
buf \U$70605 ( \70575 , \70574 );
xor \U$70606 ( \70576 , \70514 , \70575 );
xor \U$70607 ( \70577 , \19390 , \19404 );
xor \U$70608 ( \70578 , \70577 , \19425 );
buf \U$70609 ( \70579 , \70578 );
buf \U$70610 ( \70580 , \70579 );
xor \U$70611 ( \70581 , \70576 , \70580 );
buf \U$70612 ( \70582 , \70581 );
buf \U$70613 ( \70583 , \70582 );
xor \U$70614 ( \70584 , \70510 , \70583 );
xor \U$70615 ( \70585 , \19343 , \19325 );
xor \U$70616 ( \70586 , \70585 , \19365 );
buf \U$70617 ( \70587 , \70586 );
and \U$70618 ( \70588 , \19705 , \19686 );
not \U$70619 ( \70589 , \19705 );
and \U$70620 ( \70590 , \70589 , \19683 );
or \U$70621 ( \70591 , \70588 , \70590 );
and \U$70622 ( \70592 , \70591 , \19665 );
not \U$70623 ( \70593 , \70591 );
and \U$70624 ( \70594 , \70593 , \19668 );
nor \U$70625 ( \70595 , \70592 , \70594 );
buf \U$70626 ( \70596 , \70595 );
xor \U$70627 ( \70597 , \70587 , \70596 );
buf \U$70628 ( \70598 , \19475 );
not \U$70629 ( \70599 , \70598 );
buf \U$70630 ( \70600 , \19497 );
not \U$70631 ( \70601 , \70600 );
or \U$70632 ( \70602 , \70599 , \70601 );
buf \U$70633 ( \70603 , \19497 );
buf \U$70634 ( \70604 , \19475 );
or \U$70635 ( \70605 , \70603 , \70604 );
nand \U$70636 ( \70606 , \70602 , \70605 );
buf \U$70637 ( \70607 , \70606 );
buf \U$70638 ( \70608 , \70607 );
buf \U$70639 ( \70609 , \19451 );
xor \U$70640 ( \70610 , \70608 , \70609 );
buf \U$70641 ( \70611 , \70610 );
buf \U$70642 ( \70612 , \70611 );
xor \U$70643 ( \70613 , \70597 , \70612 );
buf \U$70644 ( \70614 , \70613 );
buf \U$70645 ( \70615 , \70614 );
xor \U$70646 ( \70616 , \70584 , \70615 );
buf \U$70647 ( \70617 , \70616 );
buf \U$70648 ( \70618 , \70617 );
xor \U$70649 ( \70619 , \70492 , \70618 );
buf \U$70650 ( \70620 , \70619 );
buf \U$70651 ( \70621 , \70620 );
not \U$70652 ( \70622 , \70621 );
xor \U$70653 ( \70623 , \70363 , \70383 );
xor \U$70654 ( \70624 , \70623 , \70390 );
buf \U$70655 ( \70625 , \70624 );
buf \U$70656 ( \70626 , \70625 );
not \U$70657 ( \70627 , \70626 );
buf \U$70658 ( \70628 , \68707 );
not \U$70659 ( \70629 , \70628 );
buf \U$70660 ( \70630 , \68750 );
not \U$70661 ( \70631 , \70630 );
or \U$70662 ( \70632 , \70629 , \70631 );
buf \U$70663 ( \70633 , \68723 );
nand \U$70664 ( \70634 , \70632 , \70633 );
buf \U$70665 ( \70635 , \70634 );
buf \U$70666 ( \70636 , \70635 );
buf \U$70667 ( \70637 , \68707 );
not \U$70668 ( \70638 , \70637 );
buf \U$70669 ( \70639 , \68747 );
nand \U$70670 ( \70640 , \70638 , \70639 );
buf \U$70671 ( \70641 , \70640 );
buf \U$70672 ( \70642 , \70641 );
nand \U$70673 ( \70643 , \70636 , \70642 );
buf \U$70674 ( \70644 , \70643 );
buf \U$70675 ( \70645 , \69631 );
not \U$70676 ( \70646 , \70645 );
buf \U$70677 ( \70647 , \70646 );
buf \U$70678 ( \70648 , \70647 );
not \U$70679 ( \70649 , \70648 );
buf \U$70680 ( \70650 , \69652 );
not \U$70681 ( \70651 , \70650 );
or \U$70682 ( \70652 , \70649 , \70651 );
buf \U$70683 ( \70653 , \69614 );
nand \U$70684 ( \70654 , \70652 , \70653 );
buf \U$70685 ( \70655 , \70654 );
buf \U$70686 ( \70656 , \70655 );
buf \U$70687 ( \70657 , \69649 );
buf \U$70688 ( \70658 , \69631 );
nand \U$70689 ( \70659 , \70657 , \70658 );
buf \U$70690 ( \70660 , \70659 );
buf \U$70691 ( \70661 , \70660 );
nand \U$70692 ( \70662 , \70656 , \70661 );
buf \U$70693 ( \70663 , \70662 );
buf \U$70694 ( \70664 , \70663 );
buf \U$70695 ( \70665 , \69282 );
not \U$70696 ( \70666 , \70665 );
buf \U$70697 ( \70667 , \69236 );
not \U$70698 ( \70668 , \70667 );
or \U$70699 ( \70669 , \70666 , \70668 );
buf \U$70700 ( \70670 , \69282 );
buf \U$70701 ( \70671 , \69236 );
or \U$70702 ( \70672 , \70670 , \70671 );
buf \U$70703 ( \70673 , \69254 );
nand \U$70704 ( \70674 , \70672 , \70673 );
buf \U$70705 ( \70675 , \70674 );
buf \U$70706 ( \70676 , \70675 );
nand \U$70707 ( \70677 , \70669 , \70676 );
buf \U$70708 ( \70678 , \70677 );
buf \U$70709 ( \70679 , \70678 );
xor \U$70710 ( \70680 , \70664 , \70679 );
buf \U$70711 ( \70681 , \69214 );
not \U$70712 ( \70682 , \70681 );
buf \U$70713 ( \70683 , \69192 );
not \U$70714 ( \70684 , \70683 );
or \U$70715 ( \70685 , \70682 , \70684 );
buf \U$70716 ( \70686 , \69175 );
nand \U$70717 ( \70687 , \70685 , \70686 );
buf \U$70718 ( \70688 , \70687 );
buf \U$70719 ( \70689 , \70688 );
buf \U$70720 ( \70690 , \69214 );
not \U$70721 ( \70691 , \70690 );
buf \U$70722 ( \70692 , \69189 );
nand \U$70723 ( \70693 , \70691 , \70692 );
buf \U$70724 ( \70694 , \70693 );
buf \U$70725 ( \70695 , \70694 );
nand \U$70726 ( \70696 , \70689 , \70695 );
buf \U$70727 ( \70697 , \70696 );
buf \U$70728 ( \70698 , \70697 );
xor \U$70729 ( \70699 , \70680 , \70698 );
buf \U$70730 ( \70700 , \70699 );
xnor \U$70731 ( \70701 , \70644 , \70700 );
buf \U$70732 ( \70702 , \70701 );
not \U$70733 ( \70703 , \70702 );
or \U$70734 ( \70704 , \70627 , \70703 );
buf \U$70735 ( \70705 , \70701 );
buf \U$70736 ( \70706 , \70625 );
or \U$70737 ( \70707 , \70705 , \70706 );
nand \U$70738 ( \70708 , \70704 , \70707 );
buf \U$70739 ( \70709 , \70708 );
buf \U$70740 ( \70710 , \70709 );
buf \U$70741 ( \70711 , \69154 );
not \U$70742 ( \70712 , \70711 );
buf \U$70743 ( \70713 , \69366 );
not \U$70744 ( \70714 , \70713 );
or \U$70745 ( \70715 , \70712 , \70714 );
buf \U$70746 ( \70716 , \69064 );
nand \U$70747 ( \70717 , \70715 , \70716 );
buf \U$70748 ( \70718 , \70717 );
buf \U$70749 ( \70719 , \70718 );
buf \U$70750 ( \70720 , \69366 );
not \U$70751 ( \70721 , \70720 );
buf \U$70752 ( \70722 , \70721 );
buf \U$70753 ( \70723 , \70722 );
buf \U$70754 ( \70724 , \69154 );
not \U$70755 ( \70725 , \70724 );
buf \U$70756 ( \70726 , \70725 );
buf \U$70757 ( \70727 , \70726 );
nand \U$70758 ( \70728 , \70723 , \70727 );
buf \U$70759 ( \70729 , \70728 );
buf \U$70760 ( \70730 , \70729 );
nand \U$70761 ( \70731 , \70719 , \70730 );
buf \U$70762 ( \70732 , \70731 );
buf \U$70763 ( \70733 , \70732 );
xor \U$70764 ( \70734 , \70710 , \70733 );
buf \U$70765 ( \70735 , \70339 );
not \U$70766 ( \70736 , \70735 );
buf \U$70767 ( \70737 , \70201 );
not \U$70768 ( \70738 , \70737 );
buf \U$70769 ( \70739 , \70330 );
not \U$70770 ( \70740 , \70739 );
and \U$70771 ( \70741 , \70738 , \70740 );
buf \U$70772 ( \70742 , \70201 );
buf \U$70773 ( \70743 , \70330 );
and \U$70774 ( \70744 , \70742 , \70743 );
nor \U$70775 ( \70745 , \70741 , \70744 );
buf \U$70776 ( \70746 , \70745 );
buf \U$70777 ( \70747 , \70746 );
not \U$70778 ( \70748 , \70747 );
or \U$70779 ( \70749 , \70736 , \70748 );
buf \U$70780 ( \70750 , \70746 );
buf \U$70781 ( \70751 , \70339 );
or \U$70782 ( \70752 , \70750 , \70751 );
nand \U$70783 ( \70753 , \70749 , \70752 );
buf \U$70784 ( \70754 , \70753 );
buf \U$70785 ( \70755 , \70754 );
and \U$70786 ( \70756 , \70734 , \70755 );
and \U$70787 ( \70757 , \70710 , \70733 );
or \U$70788 ( \70758 , \70756 , \70757 );
buf \U$70789 ( \70759 , \70758 );
buf \U$70790 ( \70760 , \70759 );
buf \U$70791 ( \70761 , \70644 );
not \U$70792 ( \70762 , \70761 );
buf \U$70793 ( \70763 , \70625 );
not \U$70794 ( \70764 , \70763 );
or \U$70795 ( \70765 , \70762 , \70764 );
buf \U$70796 ( \70766 , \70625 );
buf \U$70797 ( \70767 , \70644 );
or \U$70798 ( \70768 , \70766 , \70767 );
buf \U$70799 ( \70769 , \70700 );
nand \U$70800 ( \70770 , \70768 , \70769 );
buf \U$70801 ( \70771 , \70770 );
buf \U$70802 ( \70772 , \70771 );
nand \U$70803 ( \70773 , \70765 , \70772 );
buf \U$70804 ( \70774 , \70773 );
buf \U$70805 ( \70775 , \70774 );
not \U$70806 ( \70776 , \70775 );
buf \U$70807 ( \70777 , \69668 );
buf \U$70808 ( \70778 , \69601 );
or \U$70809 ( \70779 , \70777 , \70778 );
buf \U$70810 ( \70780 , \69555 );
nand \U$70811 ( \70781 , \70779 , \70780 );
buf \U$70812 ( \70782 , \70781 );
buf \U$70813 ( \70783 , \70782 );
buf \U$70814 ( \70784 , \69668 );
buf \U$70815 ( \70785 , \69601 );
nand \U$70816 ( \70786 , \70784 , \70785 );
buf \U$70817 ( \70787 , \70786 );
buf \U$70818 ( \70788 , \70787 );
nand \U$70819 ( \70789 , \70783 , \70788 );
buf \U$70820 ( \70790 , \70789 );
buf \U$70821 ( \70791 , \70790 );
not \U$70822 ( \70792 , \70791 );
buf \U$70823 ( \70793 , \69054 );
not \U$70824 ( \70794 , \70793 );
buf \U$70825 ( \70795 , \68932 );
not \U$70826 ( \70796 , \70795 );
or \U$70827 ( \70797 , \70794 , \70796 );
buf \U$70828 ( \70798 , \68982 );
nand \U$70829 ( \70799 , \70797 , \70798 );
buf \U$70830 ( \70800 , \70799 );
buf \U$70831 ( \70801 , \70800 );
buf \U$70832 ( \70802 , \68929 );
buf \U$70833 ( \70803 , \69057 );
nand \U$70834 ( \70804 , \70802 , \70803 );
buf \U$70835 ( \70805 , \70804 );
buf \U$70836 ( \70806 , \70805 );
nand \U$70837 ( \70807 , \70801 , \70806 );
buf \U$70838 ( \70808 , \70807 );
buf \U$70839 ( \70809 , \70808 );
not \U$70840 ( \70810 , \70809 );
or \U$70841 ( \70811 , \70792 , \70810 );
buf \U$70842 ( \70812 , \69356 );
buf \U$70843 ( \70813 , \69285 );
or \U$70844 ( \70814 , \70812 , \70813 );
buf \U$70845 ( \70815 , \69222 );
not \U$70846 ( \70816 , \70815 );
buf \U$70847 ( \70817 , \70816 );
buf \U$70848 ( \70818 , \70817 );
nand \U$70849 ( \70819 , \70814 , \70818 );
buf \U$70850 ( \70820 , \70819 );
buf \U$70851 ( \70821 , \70820 );
buf \U$70852 ( \70822 , \69285 );
buf \U$70853 ( \70823 , \69356 );
nand \U$70854 ( \70824 , \70822 , \70823 );
buf \U$70855 ( \70825 , \70824 );
buf \U$70856 ( \70826 , \70825 );
nand \U$70857 ( \70827 , \70821 , \70826 );
buf \U$70858 ( \70828 , \70827 );
buf \U$70859 ( \70829 , \70828 );
buf \U$70860 ( \70830 , \70808 );
not \U$70861 ( \70831 , \70830 );
buf \U$70862 ( \70832 , \70790 );
not \U$70863 ( \70833 , \70832 );
buf \U$70864 ( \70834 , \70833 );
buf \U$70865 ( \70835 , \70834 );
nand \U$70866 ( \70836 , \70831 , \70835 );
buf \U$70867 ( \70837 , \70836 );
buf \U$70868 ( \70838 , \70837 );
nand \U$70869 ( \70839 , \70829 , \70838 );
buf \U$70870 ( \70840 , \70839 );
buf \U$70871 ( \70841 , \70840 );
nand \U$70872 ( \70842 , \70811 , \70841 );
buf \U$70873 ( \70843 , \70842 );
buf \U$70874 ( \70844 , \70843 );
not \U$70875 ( \70845 , \70844 );
buf \U$70876 ( \70846 , \70845 );
buf \U$70877 ( \70847 , \70846 );
not \U$70878 ( \70848 , \70847 );
or \U$70879 ( \70849 , \70776 , \70848 );
buf \U$70880 ( \70850 , \70774 );
not \U$70881 ( \70851 , \70850 );
buf \U$70882 ( \70852 , \70851 );
buf \U$70883 ( \70853 , \70852 );
buf \U$70884 ( \70854 , \70843 );
nand \U$70885 ( \70855 , \70853 , \70854 );
buf \U$70886 ( \70856 , \70855 );
buf \U$70887 ( \70857 , \70856 );
nand \U$70888 ( \70858 , \70849 , \70857 );
buf \U$70889 ( \70859 , \70858 );
buf \U$70890 ( \70860 , \70859 );
buf \U$70891 ( \70861 , \70472 );
buf \U$70892 ( \70862 , \70437 );
and \U$70893 ( \70863 , \70861 , \70862 );
not \U$70894 ( \70864 , \70861 );
buf \U$70895 ( \70865 , \70440 );
and \U$70896 ( \70866 , \70864 , \70865 );
nor \U$70897 ( \70867 , \70863 , \70866 );
buf \U$70898 ( \70868 , \70867 );
buf \U$70899 ( \70869 , \70868 );
not \U$70900 ( \70870 , \70869 );
buf \U$70901 ( \70871 , \70457 );
not \U$70902 ( \70872 , \70871 );
and \U$70903 ( \70873 , \70870 , \70872 );
buf \U$70904 ( \70874 , \70868 );
buf \U$70905 ( \70875 , \70457 );
and \U$70906 ( \70876 , \70874 , \70875 );
nor \U$70907 ( \70877 , \70873 , \70876 );
buf \U$70908 ( \70878 , \70877 );
buf \U$70909 ( \70879 , \70878 );
not \U$70910 ( \70880 , \70879 );
buf \U$70911 ( \70881 , \70880 );
buf \U$70912 ( \70882 , \70881 );
not \U$70913 ( \70883 , \70882 );
buf \U$70914 ( \70884 , \67972 );
not \U$70915 ( \70885 , \70884 );
buf \U$70916 ( \70886 , \14608 );
not \U$70917 ( \70887 , \70886 );
or \U$70918 ( \70888 , \70885 , \70887 );
buf \U$70919 ( \70889 , \791 );
buf \U$70920 ( \70890 , \18052 );
nand \U$70921 ( \70891 , \70889 , \70890 );
buf \U$70922 ( \70892 , \70891 );
buf \U$70923 ( \70893 , \70892 );
nand \U$70924 ( \70894 , \70888 , \70893 );
buf \U$70925 ( \70895 , \70894 );
buf \U$70926 ( \70896 , \70895 );
not \U$70927 ( \70897 , \70896 );
buf \U$70928 ( \70898 , \70897 );
buf \U$70929 ( \70899 , \70898 );
not \U$70930 ( \70900 , \70899 );
buf \U$70931 ( \70901 , \67936 );
not \U$70932 ( \70902 , \70901 );
buf \U$70933 ( \70903 , \16014 );
not \U$70934 ( \70904 , \70903 );
or \U$70935 ( \70905 , \70902 , \70904 );
buf \U$70936 ( \70906 , \26301 );
buf \U$70937 ( \70907 , \19629 );
nand \U$70938 ( \70908 , \70906 , \70907 );
buf \U$70939 ( \70909 , \70908 );
buf \U$70940 ( \70910 , \70909 );
nand \U$70941 ( \70911 , \70905 , \70910 );
buf \U$70942 ( \70912 , \70911 );
buf \U$70943 ( \70913 , \70912 );
not \U$70944 ( \70914 , \70913 );
or \U$70945 ( \70915 , \70900 , \70914 );
buf \U$70946 ( \70916 , \70912 );
buf \U$70947 ( \70917 , \70898 );
or \U$70948 ( \70918 , \70916 , \70917 );
nand \U$70949 ( \70919 , \70915 , \70918 );
buf \U$70950 ( \70920 , \70919 );
buf \U$70951 ( \70921 , \70920 );
buf \U$70952 ( \70922 , \69001 );
not \U$70953 ( \70923 , \70922 );
buf \U$70954 ( \70924 , \396 );
not \U$70955 ( \70925 , \70924 );
or \U$70956 ( \70926 , \70923 , \70925 );
buf \U$70957 ( \70927 , \1025 );
buf \U$70958 ( \70928 , \19391 );
nand \U$70959 ( \70929 , \70927 , \70928 );
buf \U$70960 ( \70930 , \70929 );
buf \U$70961 ( \70931 , \70930 );
nand \U$70962 ( \70932 , \70926 , \70931 );
buf \U$70963 ( \70933 , \70932 );
buf \U$70964 ( \70934 , \70933 );
not \U$70965 ( \70935 , \70934 );
buf \U$70966 ( \70936 , \70935 );
buf \U$70967 ( \70937 , \70936 );
and \U$70968 ( \70938 , \70921 , \70937 );
not \U$70969 ( \70939 , \70921 );
buf \U$70970 ( \70940 , \70933 );
and \U$70971 ( \70941 , \70939 , \70940 );
nor \U$70972 ( \70942 , \70938 , \70941 );
buf \U$70973 ( \70943 , \70942 );
buf \U$70974 ( \70944 , \70943 );
not \U$70975 ( \70945 , \70944 );
buf \U$70976 ( \70946 , \70945 );
buf \U$70977 ( \70947 , \70946 );
not \U$70978 ( \70948 , \70947 );
or \U$70979 ( \70949 , \70883 , \70948 );
buf \U$70980 ( \70950 , \70878 );
not \U$70981 ( \70951 , \70950 );
buf \U$70982 ( \70952 , \70943 );
not \U$70983 ( \70953 , \70952 );
or \U$70984 ( \70954 , \70951 , \70953 );
buf \U$70985 ( \70955 , \12683 );
buf \U$70986 ( \70956 , RIc0d9400_64);
and \U$70987 ( \70957 , \70955 , \70956 );
buf \U$70988 ( \70958 , \70957 );
buf \U$70989 ( \70959 , \70958 );
buf \U$70990 ( \70960 , \68676 );
not \U$70991 ( \70961 , \70960 );
buf \U$70992 ( \70962 , \2358 );
not \U$70993 ( \70963 , \70962 );
or \U$70994 ( \70964 , \70961 , \70963 );
buf \U$70995 ( \70965 , \13998 );
buf \U$70996 ( \70966 , \18117 );
nand \U$70997 ( \70967 , \70965 , \70966 );
buf \U$70998 ( \70968 , \70967 );
buf \U$70999 ( \70969 , \70968 );
nand \U$71000 ( \70970 , \70964 , \70969 );
buf \U$71001 ( \70971 , \70970 );
buf \U$71002 ( \70972 , \70971 );
xor \U$71003 ( \70973 , \70959 , \70972 );
buf \U$71004 ( \70974 , \67950 );
not \U$71005 ( \70975 , \70974 );
buf \U$71006 ( \70976 , \14419 );
not \U$71007 ( \70977 , \70976 );
or \U$71008 ( \70978 , \70975 , \70977 );
buf \U$71009 ( \70979 , \14648 );
buf \U$71010 ( \70980 , \19690 );
nand \U$71011 ( \70981 , \70979 , \70980 );
buf \U$71012 ( \70982 , \70981 );
buf \U$71013 ( \70983 , \70982 );
nand \U$71014 ( \70984 , \70978 , \70983 );
buf \U$71015 ( \70985 , \70984 );
buf \U$71016 ( \70986 , \70985 );
xor \U$71017 ( \70987 , \70973 , \70986 );
buf \U$71018 ( \70988 , \70987 );
buf \U$71019 ( \70989 , \70988 );
nand \U$71020 ( \70990 , \70954 , \70989 );
buf \U$71021 ( \70991 , \70990 );
buf \U$71022 ( \70992 , \70991 );
nand \U$71023 ( \70993 , \70949 , \70992 );
buf \U$71024 ( \70994 , \70993 );
buf \U$71025 ( \70995 , \70128 );
not \U$71026 ( \70996 , \70995 );
buf \U$71027 ( \70997 , \70122 );
not \U$71028 ( \70998 , \70997 );
or \U$71029 ( \70999 , \70996 , \70998 );
not \U$71030 ( \71000 , \70119 );
not \U$71031 ( \71001 , \70073 );
or \U$71032 ( \71002 , \71000 , \71001 );
nand \U$71033 ( \71003 , \71002 , \70198 );
buf \U$71034 ( \71004 , \71003 );
nand \U$71035 ( \71005 , \70999 , \71004 );
buf \U$71036 ( \71006 , \71005 );
xor \U$71037 ( \71007 , \70994 , \71006 );
xor \U$71038 ( \71008 , \70959 , \70972 );
and \U$71039 ( \71009 , \71008 , \70986 );
and \U$71040 ( \71010 , \70959 , \70972 );
or \U$71041 ( \71011 , \71009 , \71010 );
buf \U$71042 ( \71012 , \71011 );
buf \U$71043 ( \71013 , \71012 );
buf \U$71044 ( \71014 , \70087 );
not \U$71045 ( \71015 , \71014 );
buf \U$71046 ( \71016 , \70112 );
not \U$71047 ( \71017 , \71016 );
or \U$71048 ( \71018 , \71015 , \71017 );
buf \U$71049 ( \71019 , \70087 );
buf \U$71050 ( \71020 , \70112 );
or \U$71051 ( \71021 , \71019 , \71020 );
buf \U$71052 ( \71022 , \70099 );
nand \U$71053 ( \71023 , \71021 , \71022 );
buf \U$71054 ( \71024 , \71023 );
buf \U$71055 ( \71025 , \71024 );
nand \U$71056 ( \71026 , \71018 , \71025 );
buf \U$71057 ( \71027 , \71026 );
buf \U$71058 ( \71028 , \71027 );
xor \U$71059 ( \71029 , \71013 , \71028 );
buf \U$71060 ( \71030 , \19593 );
not \U$71061 ( \71031 , \71030 );
buf \U$71062 ( \71032 , \19622 );
not \U$71063 ( \71033 , \71032 );
or \U$71064 ( \71034 , \71031 , \71033 );
buf \U$71065 ( \71035 , \19617 );
buf \U$71066 ( \71036 , \19611 );
nand \U$71067 ( \71037 , \71035 , \71036 );
buf \U$71068 ( \71038 , \71037 );
buf \U$71069 ( \71039 , \71038 );
nand \U$71070 ( \71040 , \71034 , \71039 );
buf \U$71071 ( \71041 , \71040 );
buf \U$71072 ( \71042 , \71041 );
buf \U$71073 ( \71043 , \19641 );
xor \U$71074 ( \71044 , \71042 , \71043 );
buf \U$71075 ( \71045 , \71044 );
buf \U$71076 ( \71046 , \71045 );
xor \U$71077 ( \71047 , \71029 , \71046 );
buf \U$71078 ( \71048 , \71047 );
buf \U$71081 ( \71049 , \71048 );
xor \U$71082 ( \71050 , \71007 , \71049 );
buf \U$71083 ( \71051 , \71050 );
and \U$71084 ( \71052 , \70860 , \71051 );
not \U$71085 ( \71053 , \70860 );
buf \U$71086 ( \71054 , \71050 );
not \U$71087 ( \71055 , \71054 );
buf \U$71088 ( \71056 , \71055 );
buf \U$71089 ( \71057 , \71056 );
and \U$71090 ( \71058 , \71053 , \71057 );
nor \U$71091 ( \71059 , \71052 , \71058 );
buf \U$71092 ( \71060 , \71059 );
buf \U$71093 ( \71061 , \71060 );
xor \U$71094 ( \71062 , \70760 , \71061 );
buf \U$71095 ( \71063 , \71062 );
buf \U$71096 ( \71064 , \71063 );
not \U$71097 ( \71065 , \71064 );
buf \U$71098 ( \71066 , \71065 );
buf \U$71099 ( \71067 , \71066 );
not \U$71100 ( \71068 , \71067 );
or \U$71101 ( \71069 , \70622 , \71068 );
buf \U$71102 ( \71070 , \70620 );
not \U$71103 ( \71071 , \71070 );
buf \U$71104 ( \71072 , \71063 );
nand \U$71105 ( \71073 , \71071 , \71072 );
buf \U$71106 ( \71074 , \71073 );
buf \U$71107 ( \71075 , \71074 );
nand \U$71108 ( \71076 , \71069 , \71075 );
buf \U$71109 ( \71077 , \71076 );
buf \U$71110 ( \71078 , \71077 );
buf \U$71111 ( \71079 , \69490 );
not \U$71112 ( \71080 , \71079 );
buf \U$71113 ( \71081 , \69377 );
not \U$71114 ( \71082 , \71081 );
or \U$71115 ( \71083 , \71080 , \71082 );
buf \U$71116 ( \71084 , \69701 );
nand \U$71117 ( \71085 , \71083 , \71084 );
buf \U$71118 ( \71086 , \71085 );
buf \U$71119 ( \71087 , \71086 );
buf \U$71120 ( \71088 , \69487 );
buf \U$71121 ( \71089 , \69380 );
nand \U$71122 ( \71090 , \71088 , \71089 );
buf \U$71123 ( \71091 , \71090 );
buf \U$71124 ( \71092 , \71091 );
nand \U$71125 ( \71093 , \71087 , \71092 );
buf \U$71126 ( \71094 , \71093 );
buf \U$71127 ( \71095 , \71094 );
xor \U$71128 ( \71096 , \69670 , \69692 );
and \U$71129 ( \71097 , \71096 , \69699 );
and \U$71130 ( \71098 , \69670 , \69692 );
or \U$71131 ( \71099 , \71097 , \71098 );
buf \U$71132 ( \71100 , \71099 );
buf \U$71133 ( \71101 , \71100 );
buf \U$71134 ( \71102 , \70881 );
not \U$71135 ( \71103 , \71102 );
buf \U$71136 ( \71104 , \70988 );
buf \U$71137 ( \71105 , \70943 );
and \U$71138 ( \71106 , \71104 , \71105 );
not \U$71139 ( \71107 , \71104 );
buf \U$71140 ( \71108 , \70946 );
and \U$71141 ( \71109 , \71107 , \71108 );
nor \U$71142 ( \71110 , \71106 , \71109 );
buf \U$71143 ( \71111 , \71110 );
buf \U$71144 ( \71112 , \71111 );
not \U$71145 ( \71113 , \71112 );
or \U$71146 ( \71114 , \71103 , \71113 );
buf \U$71147 ( \71115 , \71111 );
buf \U$71148 ( \71116 , \70881 );
or \U$71149 ( \71117 , \71115 , \71116 );
nand \U$71150 ( \71118 , \71114 , \71117 );
buf \U$71151 ( \71119 , \71118 );
buf \U$71152 ( \71120 , \71119 );
buf \U$71153 ( \71121 , \67981 );
not \U$71154 ( \71122 , \71121 );
buf \U$71155 ( \71123 , \68033 );
not \U$71156 ( \71124 , \71123 );
or \U$71157 ( \71125 , \71122 , \71124 );
buf \U$71158 ( \71126 , \67981 );
buf \U$71159 ( \71127 , \68033 );
or \U$71160 ( \71128 , \71126 , \71127 );
buf \U$71161 ( \71129 , \68040 );
nand \U$71162 ( \71130 , \71128 , \71129 );
buf \U$71163 ( \71131 , \71130 );
buf \U$71164 ( \71132 , \71131 );
nand \U$71165 ( \71133 , \71125 , \71132 );
buf \U$71166 ( \71134 , \71133 );
buf \U$71167 ( \71135 , \71134 );
xor \U$71168 ( \71136 , \71120 , \71135 );
buf \U$71169 ( \71137 , \70564 );
buf \U$71170 ( \71138 , \70568 );
and \U$71171 ( \71139 , \71137 , \71138 );
not \U$71172 ( \71140 , \71137 );
buf \U$71173 ( \71141 , \70555 );
and \U$71174 ( \71142 , \71140 , \71141 );
nor \U$71175 ( \71143 , \71139 , \71142 );
buf \U$71176 ( \71144 , \71143 );
buf \U$71177 ( \71145 , \71144 );
buf \U$71178 ( \71146 , \70519 );
xor \U$71179 ( \71147 , \71145 , \71146 );
buf \U$71180 ( \71148 , \71147 );
buf \U$71181 ( \71149 , \71148 );
xor \U$71182 ( \71150 , \68765 , \68771 );
and \U$71183 ( \71151 , \71150 , \68778 );
and \U$71184 ( \71152 , \68765 , \68771 );
or \U$71185 ( \71153 , \71151 , \71152 );
buf \U$71186 ( \71154 , \71153 );
buf \U$71187 ( \71155 , \71154 );
xor \U$71188 ( \71156 , \71149 , \71155 );
buf \U$71189 ( \71157 , \69080 );
not \U$71190 ( \71158 , \71157 );
buf \U$71191 ( \71159 , \69138 );
not \U$71192 ( \71160 , \71159 );
or \U$71193 ( \71161 , \71158 , \71160 );
buf \U$71194 ( \71162 , \69138 );
buf \U$71195 ( \71163 , \69080 );
or \U$71196 ( \71164 , \71162 , \71163 );
buf \U$71197 ( \71165 , \69153 );
nand \U$71198 ( \71166 , \71164 , \71165 );
buf \U$71199 ( \71167 , \71166 );
buf \U$71200 ( \71168 , \71167 );
nand \U$71201 ( \71169 , \71161 , \71168 );
buf \U$71202 ( \71170 , \71169 );
buf \U$71203 ( \71171 , \71170 );
xor \U$71204 ( \71172 , \71156 , \71171 );
buf \U$71205 ( \71173 , \71172 );
buf \U$71206 ( \71174 , \71173 );
xor \U$71207 ( \71175 , \71136 , \71174 );
buf \U$71208 ( \71176 , \71175 );
buf \U$71209 ( \71177 , \71176 );
xor \U$71210 ( \71178 , \71101 , \71177 );
buf \U$71211 ( \71179 , \68043 );
not \U$71212 ( \71180 , \71179 );
buf \U$71213 ( \71181 , \71180 );
buf \U$71214 ( \71182 , \71181 );
not \U$71215 ( \71183 , \71182 );
buf \U$71216 ( \71184 , \68057 );
not \U$71217 ( \71185 , \71184 );
or \U$71218 ( \71186 , \71183 , \71185 );
buf \U$71219 ( \71187 , \68057 );
buf \U$71220 ( \71188 , \71181 );
or \U$71221 ( \71189 , \71187 , \71188 );
buf \U$71222 ( \71190 , \68544 );
nand \U$71223 ( \71191 , \71189 , \71190 );
buf \U$71224 ( \71192 , \71191 );
buf \U$71225 ( \71193 , \71192 );
nand \U$71226 ( \71194 , \71186 , \71193 );
buf \U$71227 ( \71195 , \71194 );
buf \U$71228 ( \71196 , \71195 );
xor \U$71229 ( \71197 , \71178 , \71196 );
buf \U$71230 ( \71198 , \71197 );
buf \U$71231 ( \71199 , \71198 );
xor \U$71232 ( \71200 , \71095 , \71199 );
buf \U$71233 ( \71201 , \68545 );
not \U$71234 ( \71202 , \71201 );
buf \U$71235 ( \71203 , \68797 );
not \U$71236 ( \71204 , \71203 );
or \U$71237 ( \71205 , \71202 , \71204 );
buf \U$71238 ( \71206 , \67919 );
nand \U$71239 ( \71207 , \71205 , \71206 );
buf \U$71240 ( \71208 , \71207 );
buf \U$71241 ( \71209 , \71208 );
buf \U$71242 ( \71210 , \68545 );
not \U$71243 ( \71211 , \71210 );
buf \U$71244 ( \71212 , \68802 );
nand \U$71245 ( \71213 , \71211 , \71212 );
buf \U$71246 ( \71214 , \71213 );
buf \U$71247 ( \71215 , \71214 );
nand \U$71248 ( \71216 , \71209 , \71215 );
buf \U$71249 ( \71217 , \71216 );
buf \U$71250 ( \71218 , \71217 );
and \U$71251 ( \71219 , \71200 , \71218 );
and \U$71252 ( \71220 , \71095 , \71199 );
or \U$71253 ( \71221 , \71219 , \71220 );
buf \U$71254 ( \71222 , \71221 );
buf \U$71255 ( \71223 , \71222 );
xor \U$71256 ( \71224 , \71078 , \71223 );
xor \U$71257 ( \71225 , \71101 , \71177 );
and \U$71258 ( \71226 , \71225 , \71196 );
and \U$71259 ( \71227 , \71101 , \71177 );
or \U$71260 ( \71228 , \71226 , \71227 );
buf \U$71261 ( \71229 , \71228 );
buf \U$71262 ( \71230 , \71229 );
xor \U$71263 ( \71231 , \71120 , \71135 );
and \U$71264 ( \71232 , \71231 , \71174 );
and \U$71265 ( \71233 , \71120 , \71135 );
or \U$71266 ( \71234 , \71232 , \71233 );
buf \U$71267 ( \71235 , \71234 );
buf \U$71268 ( \71236 , \71235 );
buf \U$71269 ( \71237 , \68229 );
buf \U$71270 ( \71238 , \68369 );
buf \U$71271 ( \71239 , \68534 );
nor \U$71272 ( \71240 , \71238 , \71239 );
buf \U$71273 ( \71241 , \71240 );
buf \U$71274 ( \71242 , \71241 );
or \U$71275 ( \71243 , \71237 , \71242 );
buf \U$71276 ( \71244 , \68534 );
buf \U$71277 ( \71245 , \68369 );
nand \U$71278 ( \71246 , \71244 , \71245 );
buf \U$71279 ( \71247 , \71246 );
buf \U$71280 ( \71248 , \71247 );
nand \U$71281 ( \71249 , \71243 , \71248 );
buf \U$71282 ( \71250 , \71249 );
buf \U$71283 ( \71251 , \71250 );
not \U$71284 ( \71252 , \68669 );
nand \U$71285 ( \71253 , \71252 , \68758 );
not \U$71286 ( \71254 , \71253 );
not \U$71287 ( \71255 , \68780 );
or \U$71288 ( \71256 , \71254 , \71255 );
buf \U$71289 ( \71257 , \68758 );
not \U$71290 ( \71258 , \71257 );
buf \U$71291 ( \71259 , \68669 );
nand \U$71292 ( \71260 , \71258 , \71259 );
buf \U$71293 ( \71261 , \71260 );
nand \U$71294 ( \71262 , \71256 , \71261 );
buf \U$71295 ( \71263 , \71262 );
xor \U$71296 ( \71264 , \71251 , \71263 );
buf \U$71297 ( \71265 , \70808 );
buf \U$71298 ( \71266 , \70790 );
xor \U$71299 ( \71267 , \71265 , \71266 );
buf \U$71300 ( \71268 , \70828 );
xor \U$71301 ( \71269 , \71267 , \71268 );
buf \U$71302 ( \71270 , \71269 );
buf \U$71303 ( \71271 , \71270 );
and \U$71304 ( \71272 , \71264 , \71271 );
and \U$71305 ( \71273 , \71251 , \71263 );
or \U$71306 ( \71274 , \71272 , \71273 );
buf \U$71307 ( \71275 , \71274 );
buf \U$71308 ( \71276 , \71275 );
xor \U$71309 ( \71277 , \71236 , \71276 );
buf \U$71310 ( \71278 , \18188 );
buf \U$71311 ( \71279 , \18209 );
xor \U$71312 ( \71280 , \71278 , \71279 );
buf \U$71313 ( \71281 , \18231 );
xor \U$71314 ( \71282 , \71280 , \71281 );
buf \U$71315 ( \71283 , \71282 );
xor \U$71316 ( \71284 , \19948 , \19963 );
xor \U$71317 ( \71285 , \71284 , \19981 );
buf \U$71318 ( \71286 , \71285 );
xor \U$71319 ( \71287 , \71283 , \71286 );
buf \U$71320 ( \71288 , \18111 );
not \U$71321 ( \71289 , \71288 );
buf \U$71322 ( \71290 , \18130 );
not \U$71323 ( \71291 , \71290 );
or \U$71324 ( \71292 , \71289 , \71291 );
buf \U$71325 ( \71293 , \18133 );
buf \U$71326 ( \71294 , \18139 );
nand \U$71327 ( \71295 , \71293 , \71294 );
buf \U$71328 ( \71296 , \71295 );
buf \U$71329 ( \71297 , \71296 );
nand \U$71330 ( \71298 , \71292 , \71297 );
buf \U$71331 ( \71299 , \71298 );
buf \U$71332 ( \71300 , \71299 );
buf \U$71333 ( \71301 , \18160 );
xor \U$71334 ( \71302 , \71300 , \71301 );
buf \U$71335 ( \71303 , \71302 );
xor \U$71336 ( \71304 , \71287 , \71303 );
buf \U$71337 ( \71305 , \71304 );
xor \U$71338 ( \71306 , \71149 , \71155 );
and \U$71339 ( \71307 , \71306 , \71171 );
and \U$71340 ( \71308 , \71149 , \71155 );
or \U$71341 ( \71309 , \71307 , \71308 );
buf \U$71342 ( \71310 , \71309 );
buf \U$71343 ( \71311 , \71310 );
xor \U$71344 ( \71312 , \71305 , \71311 );
buf \U$71345 ( \71313 , \61887 );
buf \U$71346 ( \71314 , \70550 );
not \U$71347 ( \71315 , \71314 );
buf \U$71348 ( \71316 , \71315 );
buf \U$71349 ( \71317 , \71316 );
or \U$71350 ( \71318 , \71313 , \71317 );
buf \U$71351 ( \71319 , \12647 );
buf \U$71352 ( \71320 , \17203 );
not \U$71353 ( \71321 , \71320 );
buf \U$71354 ( \71322 , \71321 );
buf \U$71355 ( \71323 , \71322 );
or \U$71356 ( \71324 , \71319 , \71323 );
nand \U$71357 ( \71325 , \71318 , \71324 );
buf \U$71358 ( \71326 , \71325 );
buf \U$71359 ( \71327 , \71326 );
buf \U$71360 ( \71328 , \18071 );
buf \U$71361 ( \71329 , \18087 );
xor \U$71362 ( \71330 , \71328 , \71329 );
buf \U$71363 ( \71331 , \71330 );
buf \U$71364 ( \71332 , \71331 );
xor \U$71365 ( \71333 , \71327 , \71332 );
buf \U$71366 ( \71334 , \70898 );
not \U$71367 ( \71335 , \71334 );
buf \U$71368 ( \71336 , \70936 );
not \U$71369 ( \71337 , \71336 );
or \U$71370 ( \71338 , \71335 , \71337 );
buf \U$71371 ( \71339 , \70912 );
nand \U$71372 ( \71340 , \71338 , \71339 );
buf \U$71373 ( \71341 , \71340 );
buf \U$71374 ( \71342 , \71341 );
buf \U$71375 ( \71343 , \70933 );
buf \U$71376 ( \71344 , \70895 );
nand \U$71377 ( \71345 , \71343 , \71344 );
buf \U$71378 ( \71346 , \71345 );
buf \U$71379 ( \71347 , \71346 );
nand \U$71380 ( \71348 , \71342 , \71347 );
buf \U$71381 ( \71349 , \71348 );
buf \U$71382 ( \71350 , \71349 );
xor \U$71383 ( \71351 , \71333 , \71350 );
buf \U$71384 ( \71352 , \71351 );
buf \U$71385 ( \71353 , \71352 );
not \U$71386 ( \71354 , \71353 );
xor \U$71387 ( \71355 , \70664 , \70679 );
and \U$71388 ( \71356 , \71355 , \70698 );
and \U$71389 ( \71357 , \70664 , \70679 );
or \U$71390 ( \71358 , \71356 , \71357 );
buf \U$71391 ( \71359 , \71358 );
buf \U$71392 ( \71360 , \70326 );
not \U$71393 ( \71361 , \71360 );
buf \U$71394 ( \71362 , \70306 );
not \U$71395 ( \71363 , \71362 );
or \U$71396 ( \71364 , \71361 , \71363 );
buf \U$71397 ( \71365 , \70296 );
nand \U$71398 ( \71366 , \71364 , \71365 );
buf \U$71399 ( \71367 , \71366 );
buf \U$71400 ( \71368 , \71367 );
buf \U$71401 ( \71369 , \70303 );
buf \U$71402 ( \71370 , \70320 );
nand \U$71403 ( \71371 , \71369 , \71370 );
buf \U$71404 ( \71372 , \71371 );
buf \U$71405 ( \71373 , \71372 );
nand \U$71406 ( \71374 , \71368 , \71373 );
buf \U$71407 ( \71375 , \71374 );
xnor \U$71408 ( \71376 , \71359 , \71375 );
buf \U$71409 ( \71377 , \71376 );
not \U$71410 ( \71378 , \71377 );
or \U$71411 ( \71379 , \71354 , \71378 );
buf \U$71412 ( \71380 , \71376 );
buf \U$71413 ( \71381 , \71352 );
or \U$71414 ( \71382 , \71380 , \71381 );
nand \U$71415 ( \71383 , \71379 , \71382 );
buf \U$71416 ( \71384 , \71383 );
buf \U$71417 ( \71385 , \71384 );
xor \U$71418 ( \71386 , \71312 , \71385 );
buf \U$71419 ( \71387 , \71386 );
buf \U$71420 ( \71388 , \71387 );
xor \U$71421 ( \71389 , \71277 , \71388 );
buf \U$71422 ( \71390 , \71389 );
buf \U$71423 ( \71391 , \71390 );
xor \U$71424 ( \71392 , \71230 , \71391 );
xor \U$71425 ( \71393 , \71251 , \71263 );
xor \U$71426 ( \71394 , \71393 , \71271 );
buf \U$71427 ( \71395 , \71394 );
buf \U$71428 ( \71396 , \71395 );
xor \U$71429 ( \71397 , \70710 , \70733 );
xor \U$71430 ( \71398 , \71397 , \70755 );
buf \U$71431 ( \71399 , \71398 );
buf \U$71432 ( \71400 , \71399 );
xor \U$71433 ( \71401 , \71396 , \71400 );
buf \U$71434 ( \71402 , \68586 );
buf \U$71435 ( \71403 , \68781 );
not \U$71436 ( \71404 , \71403 );
buf \U$71437 ( \71405 , \71404 );
buf \U$71438 ( \71406 , \71405 );
or \U$71439 ( \71407 , \71402 , \71406 );
buf \U$71440 ( \71408 , \68653 );
nand \U$71441 ( \71409 , \71407 , \71408 );
buf \U$71442 ( \71410 , \71409 );
buf \U$71443 ( \71411 , \71410 );
buf \U$71444 ( \71412 , \68586 );
buf \U$71445 ( \71413 , \71405 );
nand \U$71446 ( \71414 , \71412 , \71413 );
buf \U$71447 ( \71415 , \71414 );
buf \U$71448 ( \71416 , \71415 );
nand \U$71449 ( \71417 , \71411 , \71416 );
buf \U$71450 ( \71418 , \71417 );
buf \U$71451 ( \71419 , \71418 );
and \U$71452 ( \71420 , \71401 , \71419 );
and \U$71453 ( \71421 , \71396 , \71400 );
or \U$71454 ( \71422 , \71420 , \71421 );
buf \U$71455 ( \71423 , \71422 );
buf \U$71456 ( \71424 , \71423 );
xor \U$71457 ( \71425 , \71392 , \71424 );
buf \U$71458 ( \71426 , \71425 );
buf \U$71459 ( \71427 , \71426 );
xor \U$71460 ( \71428 , \71224 , \71427 );
buf \U$71461 ( \71429 , \71428 );
buf \U$71462 ( \71430 , \71429 );
not \U$71463 ( \71431 , \71430 );
buf \U$71464 ( \71432 , \71431 );
buf \U$71465 ( \71433 , \71432 );
xor \U$71466 ( \71434 , \71396 , \71400 );
xor \U$71467 ( \71435 , \71434 , \71419 );
buf \U$71468 ( \71436 , \71435 );
buf \U$71469 ( \71437 , \71436 );
not \U$71470 ( \71438 , \71437 );
buf \U$71471 ( \71439 , \69717 );
not \U$71472 ( \71440 , \71439 );
buf \U$71473 ( \71441 , \68911 );
not \U$71474 ( \71442 , \71441 );
buf \U$71475 ( \71443 , \71442 );
buf \U$71476 ( \71444 , \71443 );
not \U$71477 ( \71445 , \71444 );
or \U$71478 ( \71446 , \71440 , \71445 );
buf \U$71479 ( \71447 , \69711 );
not \U$71480 ( \71448 , \71447 );
buf \U$71481 ( \71449 , \68911 );
not \U$71482 ( \71450 , \71449 );
or \U$71483 ( \71451 , \71448 , \71450 );
buf \U$71484 ( \71452 , \69759 );
nand \U$71485 ( \71453 , \71451 , \71452 );
buf \U$71486 ( \71454 , \71453 );
buf \U$71487 ( \71455 , \71454 );
nand \U$71488 ( \71456 , \71446 , \71455 );
buf \U$71489 ( \71457 , \71456 );
buf \U$71490 ( \71458 , \71457 );
not \U$71491 ( \71459 , \71458 );
or \U$71492 ( \71460 , \71438 , \71459 );
or \U$71493 ( \71461 , \71457 , \71436 );
xor \U$71494 ( \71462 , \71095 , \71199 );
xor \U$71495 ( \71463 , \71462 , \71218 );
buf \U$71496 ( \71464 , \71463 );
nand \U$71497 ( \71465 , \71461 , \71464 );
buf \U$71498 ( \71466 , \71465 );
nand \U$71499 ( \71467 , \71460 , \71466 );
buf \U$71500 ( \71468 , \71467 );
buf \U$71501 ( \71469 , \71468 );
not \U$71502 ( \71470 , \71469 );
buf \U$71503 ( \71471 , \71470 );
buf \U$71504 ( \71472 , \71471 );
nand \U$71505 ( \71473 , \71433 , \71472 );
buf \U$71506 ( \71474 , \71473 );
buf \U$71507 ( \71475 , \71474 );
buf \U$71508 ( \71476 , \71060 );
not \U$71509 ( \71477 , \71476 );
buf \U$71510 ( \71478 , \70759 );
not \U$71511 ( \71479 , \71478 );
or \U$71512 ( \71480 , \71477 , \71479 );
buf \U$71513 ( \71481 , \70759 );
buf \U$71514 ( \71482 , \71060 );
or \U$71515 ( \71483 , \71481 , \71482 );
buf \U$71516 ( \71484 , \70620 );
nand \U$71517 ( \71485 , \71483 , \71484 );
buf \U$71518 ( \71486 , \71485 );
buf \U$71519 ( \71487 , \71486 );
nand \U$71520 ( \71488 , \71480 , \71487 );
buf \U$71521 ( \71489 , \71488 );
buf \U$71522 ( \71490 , \71489 );
buf \U$71523 ( \71491 , \71048 );
not \U$71524 ( \71492 , \71491 );
buf \U$71525 ( \71493 , \71006 );
not \U$71526 ( \71494 , \71493 );
or \U$71527 ( \71495 , \71492 , \71494 );
buf \U$71528 ( \71496 , \71048 );
buf \U$71529 ( \71497 , \71006 );
or \U$71530 ( \71498 , \71496 , \71497 );
buf \U$71531 ( \71499 , \70994 );
nand \U$71532 ( \71500 , \71498 , \71499 );
buf \U$71533 ( \71501 , \71500 );
buf \U$71534 ( \71502 , \71501 );
nand \U$71535 ( \71503 , \71495 , \71502 );
buf \U$71536 ( \71504 , \71503 );
buf \U$71537 ( \71505 , \71504 );
buf \U$71538 ( \71506 , \70394 );
not \U$71539 ( \71507 , \71506 );
buf \U$71540 ( \71508 , \70398 );
not \U$71541 ( \71509 , \71508 );
or \U$71542 ( \71510 , \71507 , \71509 );
buf \U$71543 ( \71511 , \70398 );
buf \U$71544 ( \71512 , \70394 );
or \U$71545 ( \71513 , \71511 , \71512 );
buf \U$71546 ( \71514 , \70487 );
nand \U$71547 ( \71515 , \71513 , \71514 );
buf \U$71548 ( \71516 , \71515 );
buf \U$71549 ( \71517 , \71516 );
nand \U$71550 ( \71518 , \71510 , \71517 );
buf \U$71551 ( \71519 , \71518 );
buf \U$71552 ( \71520 , \71519 );
xor \U$71553 ( \71521 , \71505 , \71520 );
buf \U$71554 ( \71522 , \71521 );
buf \U$71555 ( \71523 , \71522 );
xor \U$71556 ( \71524 , \70510 , \70583 );
and \U$71557 ( \71525 , \71524 , \70615 );
and \U$71558 ( \71526 , \70510 , \70583 );
or \U$71559 ( \71527 , \71525 , \71526 );
buf \U$71560 ( \71528 , \71527 );
buf \U$71561 ( \71529 , \71528 );
xor \U$71562 ( \71530 , \71523 , \71529 );
buf \U$71563 ( \71531 , \71530 );
buf \U$71564 ( \71532 , \71531 );
xor \U$71565 ( \71533 , \70346 , \70491 );
and \U$71566 ( \71534 , \71533 , \70618 );
and \U$71567 ( \71535 , \70346 , \70491 );
or \U$71568 ( \71536 , \71534 , \71535 );
buf \U$71569 ( \71537 , \71536 );
buf \U$71570 ( \71538 , \71537 );
xor \U$71571 ( \71539 , \71532 , \71538 );
xor \U$71572 ( \71540 , \71013 , \71028 );
and \U$71573 ( \71541 , \71540 , \71046 );
and \U$71574 ( \71542 , \71013 , \71028 );
or \U$71575 ( \71543 , \71541 , \71542 );
buf \U$71576 ( \71544 , \71543 );
buf \U$71577 ( \71545 , \71544 );
xor \U$71578 ( \71546 , \19931 , \19986 );
xor \U$71579 ( \71547 , \71546 , \19997 );
buf \U$71580 ( \71548 , \71547 );
buf \U$71581 ( \71549 , \71548 );
xor \U$71582 ( \71550 , \71545 , \71549 );
xor \U$71583 ( \71551 , \70587 , \70596 );
and \U$71584 ( \71552 , \71551 , \70612 );
and \U$71585 ( \71553 , \70587 , \70596 );
or \U$71586 ( \71554 , \71552 , \71553 );
buf \U$71587 ( \71555 , \71554 );
buf \U$71588 ( \71556 , \71555 );
xor \U$71589 ( \71557 , \71550 , \71556 );
buf \U$71590 ( \71558 , \71557 );
buf \U$71591 ( \71559 , \71558 );
not \U$71592 ( \71560 , \71559 );
xor \U$71593 ( \71561 , \18091 , \18167 );
xor \U$71594 ( \71562 , \71561 , \18243 );
buf \U$71595 ( \71563 , \71562 );
buf \U$71596 ( \71564 , \71563 );
buf \U$71597 ( \71565 , \71303 );
not \U$71598 ( \71566 , \71565 );
buf \U$71599 ( \71567 , \71286 );
not \U$71600 ( \71568 , \71567 );
or \U$71601 ( \71569 , \71566 , \71568 );
buf \U$71602 ( \71570 , \71286 );
buf \U$71603 ( \71571 , \71303 );
or \U$71604 ( \71572 , \71570 , \71571 );
buf \U$71605 ( \71573 , \71283 );
nand \U$71606 ( \71574 , \71572 , \71573 );
buf \U$71607 ( \71575 , \71574 );
buf \U$71608 ( \71576 , \71575 );
nand \U$71609 ( \71577 , \71569 , \71576 );
buf \U$71610 ( \71578 , \71577 );
buf \U$71611 ( \71579 , \71578 );
xor \U$71612 ( \71580 , \71564 , \71579 );
buf \U$71613 ( \71581 , \19429 );
not \U$71614 ( \71582 , \71581 );
buf \U$71615 ( \71583 , \71582 );
buf \U$71616 ( \71584 , \71583 );
not \U$71617 ( \71585 , \71584 );
xor \U$71618 ( \71586 , \19508 , \19371 );
buf \U$71619 ( \71587 , \71586 );
not \U$71620 ( \71588 , \71587 );
or \U$71621 ( \71589 , \71585 , \71588 );
buf \U$71622 ( \71590 , \71586 );
buf \U$71623 ( \71591 , \71583 );
or \U$71624 ( \71592 , \71590 , \71591 );
nand \U$71625 ( \71593 , \71589 , \71592 );
buf \U$71626 ( \71594 , \71593 );
buf \U$71627 ( \71595 , \71594 );
xor \U$71628 ( \71596 , \71580 , \71595 );
buf \U$71629 ( \71597 , \71596 );
buf \U$71630 ( \71598 , \71597 );
not \U$71631 ( \71599 , \71598 );
buf \U$71632 ( \71600 , \71599 );
buf \U$71633 ( \71601 , \71600 );
not \U$71634 ( \71602 , \71601 );
or \U$71635 ( \71603 , \71560 , \71602 );
buf \U$71636 ( \71604 , \71558 );
not \U$71637 ( \71605 , \71604 );
buf \U$71638 ( \71606 , \71605 );
buf \U$71639 ( \71607 , \71606 );
buf \U$71640 ( \71608 , \71597 );
nand \U$71641 ( \71609 , \71607 , \71608 );
buf \U$71642 ( \71610 , \71609 );
buf \U$71643 ( \71611 , \71610 );
nand \U$71644 ( \71612 , \71603 , \71611 );
buf \U$71645 ( \71613 , \71612 );
buf \U$71646 ( \71614 , \71613 );
buf \U$71647 ( \71615 , \19788 );
not \U$71648 ( \71616 , \71615 );
buf \U$71649 ( \71617 , \19796 );
not \U$71650 ( \71618 , \71617 );
or \U$71651 ( \71619 , \71616 , \71618 );
buf \U$71652 ( \71620 , \19796 );
buf \U$71653 ( \71621 , \19788 );
or \U$71654 ( \71622 , \71620 , \71621 );
nand \U$71655 ( \71623 , \71619 , \71622 );
buf \U$71656 ( \71624 , \71623 );
buf \U$71657 ( \71625 , \71624 );
buf \U$71658 ( \71626 , \19771 );
not \U$71659 ( \71627 , \71626 );
buf \U$71660 ( \71628 , \71627 );
buf \U$71661 ( \71629 , \71628 );
and \U$71662 ( \71630 , \71625 , \71629 );
not \U$71663 ( \71631 , \71625 );
buf \U$71664 ( \71632 , \19771 );
and \U$71665 ( \71633 , \71631 , \71632 );
nor \U$71666 ( \71634 , \71630 , \71633 );
buf \U$71667 ( \71635 , \71634 );
xor \U$71668 ( \71636 , \70514 , \70575 );
and \U$71669 ( \71637 , \71636 , \70580 );
and \U$71670 ( \71638 , \70514 , \70575 );
or \U$71671 ( \71639 , \71637 , \71638 );
buf \U$71672 ( \71640 , \71639 );
and \U$71673 ( \71641 , \71635 , \71640 );
not \U$71674 ( \71642 , \71635 );
buf \U$71675 ( \71643 , \71640 );
not \U$71676 ( \71644 , \71643 );
buf \U$71677 ( \71645 , \71644 );
and \U$71678 ( \71646 , \71642 , \71645 );
nor \U$71679 ( \71647 , \71641 , \71646 );
buf \U$71680 ( \71648 , \20047 );
not \U$71681 ( \71649 , \71648 );
buf \U$71682 ( \71650 , \20012 );
not \U$71683 ( \71651 , \71650 );
buf \U$71684 ( \71652 , \71651 );
buf \U$71685 ( \71653 , \71652 );
not \U$71686 ( \71654 , \71653 );
or \U$71687 ( \71655 , \71649 , \71654 );
buf \U$71688 ( \71656 , \20012 );
buf \U$71689 ( \71657 , \20044 );
nand \U$71690 ( \71658 , \71656 , \71657 );
buf \U$71691 ( \71659 , \71658 );
buf \U$71692 ( \71660 , \71659 );
nand \U$71693 ( \71661 , \71655 , \71660 );
buf \U$71694 ( \71662 , \71661 );
buf \U$71695 ( \71663 , \71662 );
buf \U$71696 ( \71664 , \20016 );
xor \U$71697 ( \71665 , \71663 , \71664 );
buf \U$71698 ( \71666 , \71665 );
xor \U$71699 ( \71667 , \71647 , \71666 );
buf \U$71700 ( \71668 , \71667 );
not \U$71701 ( \71669 , \71668 );
buf \U$71702 ( \71670 , \71669 );
buf \U$71703 ( \71671 , \71670 );
and \U$71704 ( \71672 , \71614 , \71671 );
not \U$71705 ( \71673 , \71614 );
buf \U$71706 ( \71674 , \71667 );
and \U$71707 ( \71675 , \71673 , \71674 );
nor \U$71708 ( \71676 , \71672 , \71675 );
buf \U$71709 ( \71677 , \71676 );
buf \U$71710 ( \71678 , \71677 );
xor \U$71711 ( \71679 , \71539 , \71678 );
buf \U$71712 ( \71680 , \71679 );
buf \U$71713 ( \71681 , \71680 );
xor \U$71714 ( \71682 , \71490 , \71681 );
xor \U$71715 ( \71683 , \71236 , \71276 );
and \U$71716 ( \71684 , \71683 , \71388 );
and \U$71717 ( \71685 , \71236 , \71276 );
or \U$71718 ( \71686 , \71684 , \71685 );
buf \U$71719 ( \71687 , \71686 );
buf \U$71720 ( \71688 , \71687 );
not \U$71721 ( \71689 , \71688 );
buf \U$71722 ( \71690 , \71689 );
buf \U$71723 ( \71691 , \71690 );
not \U$71724 ( \71692 , \71691 );
xor \U$71725 ( \71693 , \20084 , \20087 );
xor \U$71726 ( \71694 , \71693 , \20296 );
buf \U$71727 ( \71695 , \71694 );
buf \U$71728 ( \71696 , \71695 );
buf \U$71729 ( \71697 , \71375 );
not \U$71730 ( \71698 , \71697 );
buf \U$71731 ( \71699 , \71352 );
not \U$71732 ( \71700 , \71699 );
or \U$71733 ( \71701 , \71698 , \71700 );
buf \U$71734 ( \71702 , \71352 );
buf \U$71735 ( \71703 , \71375 );
or \U$71736 ( \71704 , \71702 , \71703 );
buf \U$71737 ( \71705 , \71359 );
nand \U$71738 ( \71706 , \71704 , \71705 );
buf \U$71739 ( \71707 , \71706 );
buf \U$71740 ( \71708 , \71707 );
nand \U$71741 ( \71709 , \71701 , \71708 );
buf \U$71742 ( \71710 , \71709 );
buf \U$71743 ( \71711 , \71710 );
xor \U$71744 ( \71712 , \71696 , \71711 );
xor \U$71745 ( \71713 , \71327 , \71332 );
and \U$71746 ( \71714 , \71713 , \71350 );
and \U$71747 ( \71715 , \71327 , \71332 );
or \U$71748 ( \71716 , \71714 , \71715 );
buf \U$71749 ( \71717 , \71716 );
buf \U$71750 ( \71718 , \71717 );
xor \U$71751 ( \71719 , \70409 , \70424 );
and \U$71752 ( \71720 , \71719 , \70485 );
and \U$71753 ( \71721 , \70409 , \70424 );
or \U$71754 ( \71722 , \71720 , \71721 );
buf \U$71755 ( \71723 , \71722 );
buf \U$71756 ( \71724 , \71723 );
xor \U$71757 ( \71725 , \71718 , \71724 );
xor \U$71758 ( \71726 , \19577 , \19647 );
xor \U$71759 ( \71727 , \71726 , \19716 );
buf \U$71760 ( \71728 , \71727 );
xor \U$71761 ( \71729 , \71725 , \71728 );
buf \U$71762 ( \71730 , \71729 );
buf \U$71763 ( \71731 , \71730 );
xor \U$71764 ( \71732 , \71712 , \71731 );
buf \U$71765 ( \71733 , \71732 );
buf \U$71766 ( \71734 , \70843 );
not \U$71767 ( \71735 , \71734 );
buf \U$71768 ( \71736 , \70774 );
not \U$71769 ( \71737 , \71736 );
or \U$71770 ( \71738 , \71735 , \71737 );
buf \U$71771 ( \71739 , \70774 );
buf \U$71772 ( \71740 , \70843 );
or \U$71773 ( \71741 , \71739 , \71740 );
buf \U$71774 ( \71742 , \71050 );
nand \U$71775 ( \71743 , \71741 , \71742 );
buf \U$71776 ( \71744 , \71743 );
buf \U$71777 ( \71745 , \71744 );
nand \U$71778 ( \71746 , \71738 , \71745 );
buf \U$71779 ( \71747 , \71746 );
xor \U$71780 ( \71748 , \71733 , \71747 );
buf \U$71781 ( \71749 , \71748 );
xor \U$71782 ( \71750 , \71305 , \71311 );
and \U$71783 ( \71751 , \71750 , \71385 );
and \U$71784 ( \71752 , \71305 , \71311 );
or \U$71785 ( \71753 , \71751 , \71752 );
buf \U$71786 ( \71754 , \71753 );
buf \U$71787 ( \71755 , \71754 );
not \U$71788 ( \71756 , \71755 );
buf \U$71789 ( \71757 , \71756 );
buf \U$71790 ( \71758 , \71757 );
and \U$71791 ( \71759 , \71749 , \71758 );
not \U$71792 ( \71760 , \71749 );
buf \U$71793 ( \71761 , \71754 );
and \U$71794 ( \71762 , \71760 , \71761 );
nor \U$71795 ( \71763 , \71759 , \71762 );
buf \U$71796 ( \71764 , \71763 );
not \U$71797 ( \71765 , \71764 );
buf \U$71798 ( \71766 , \71765 );
not \U$71799 ( \71767 , \71766 );
or \U$71800 ( \71768 , \71692 , \71767 );
buf \U$71801 ( \71769 , \71764 );
buf \U$71802 ( \71770 , \71687 );
nand \U$71803 ( \71771 , \71769 , \71770 );
buf \U$71804 ( \71772 , \71771 );
buf \U$71805 ( \71773 , \71772 );
nand \U$71806 ( \71774 , \71768 , \71773 );
buf \U$71807 ( \71775 , \71774 );
buf \U$71808 ( \71776 , \71775 );
xor \U$71809 ( \71777 , \71682 , \71776 );
buf \U$71810 ( \71778 , \71777 );
buf \U$71811 ( \71779 , \71778 );
xor \U$71812 ( \71780 , \71230 , \71391 );
and \U$71813 ( \71781 , \71780 , \71424 );
and \U$71814 ( \71782 , \71230 , \71391 );
or \U$71815 ( \71783 , \71781 , \71782 );
buf \U$71816 ( \71784 , \71783 );
buf \U$71817 ( \71785 , \71784 );
xnor \U$71818 ( \71786 , \71779 , \71785 );
buf \U$71819 ( \71787 , \71786 );
buf \U$71820 ( \71788 , \71787 );
buf \U$71821 ( \71789 , \71222 );
buf \U$71822 ( \71790 , \71077 );
or \U$71823 ( \71791 , \71789 , \71790 );
buf \U$71824 ( \71792 , \71791 );
buf \U$71825 ( \71793 , \71792 );
buf \U$71826 ( \71794 , \71426 );
and \U$71827 ( \71795 , \71793 , \71794 );
buf \U$71828 ( \71796 , \71222 );
buf \U$71829 ( \71797 , \71077 );
and \U$71830 ( \71798 , \71796 , \71797 );
buf \U$71831 ( \71799 , \71798 );
buf \U$71832 ( \71800 , \71799 );
nor \U$71833 ( \71801 , \71795 , \71800 );
buf \U$71834 ( \71802 , \71801 );
buf \U$71835 ( \71803 , \71802 );
nand \U$71836 ( \71804 , \71788 , \71803 );
buf \U$71837 ( \71805 , \71804 );
buf \U$71838 ( \71806 , \71805 );
xor \U$71839 ( \71807 , \71545 , \71549 );
and \U$71840 ( \71808 , \71807 , \71556 );
and \U$71841 ( \71809 , \71545 , \71549 );
or \U$71842 ( \71810 , \71808 , \71809 );
buf \U$71843 ( \71811 , \71810 );
buf \U$71844 ( \71812 , \71811 );
xor \U$71845 ( \71813 , \19761 , \19768 );
xor \U$71846 ( \71814 , \71813 , \19808 );
buf \U$71847 ( \71815 , \71814 );
buf \U$71848 ( \71816 , \71815 );
xor \U$71849 ( \71817 , \71812 , \71816 );
xor \U$71850 ( \71818 , \20061 , \20080 );
xor \U$71851 ( \71819 , \71818 , \20301 );
buf \U$71852 ( \71820 , \71819 );
buf \U$71853 ( \71821 , \71820 );
xor \U$71854 ( \71822 , \71817 , \71821 );
buf \U$71855 ( \71823 , \71822 );
buf \U$71856 ( \71824 , \71823 );
buf \U$71857 ( \71825 , \71597 );
not \U$71858 ( \71826 , \71825 );
buf \U$71859 ( \71827 , \71670 );
not \U$71860 ( \71828 , \71827 );
or \U$71861 ( \71829 , \71826 , \71828 );
buf \U$71862 ( \71830 , \71600 );
not \U$71863 ( \71831 , \71830 );
buf \U$71864 ( \71832 , \71667 );
not \U$71865 ( \71833 , \71832 );
or \U$71866 ( \71834 , \71831 , \71833 );
buf \U$71867 ( \71835 , \71558 );
nand \U$71868 ( \71836 , \71834 , \71835 );
buf \U$71869 ( \71837 , \71836 );
buf \U$71870 ( \71838 , \71837 );
nand \U$71871 ( \71839 , \71829 , \71838 );
buf \U$71872 ( \71840 , \71839 );
buf \U$71873 ( \71841 , \71840 );
and \U$71874 ( \71842 , \71824 , \71841 );
not \U$71875 ( \71843 , \71824 );
buf \U$71876 ( \71844 , \71840 );
not \U$71877 ( \71845 , \71844 );
buf \U$71878 ( \71846 , \71845 );
buf \U$71879 ( \71847 , \71846 );
and \U$71880 ( \71848 , \71843 , \71847 );
nor \U$71881 ( \71849 , \71842 , \71848 );
buf \U$71882 ( \71850 , \71849 );
buf \U$71883 ( \71851 , \71850 );
xor \U$71884 ( \71852 , \71718 , \71724 );
and \U$71885 ( \71853 , \71852 , \71728 );
and \U$71886 ( \71854 , \71718 , \71724 );
or \U$71887 ( \71855 , \71853 , \71854 );
buf \U$71888 ( \71856 , \71855 );
buf \U$71889 ( \71857 , \71856 );
not \U$71890 ( \71858 , \71857 );
buf \U$71891 ( \71859 , \71858 );
buf \U$71892 ( \71860 , \71859 );
not \U$71893 ( \71861 , \71860 );
buf \U$71894 ( \71862 , \71645 );
not \U$71895 ( \71863 , \71862 );
buf \U$71896 ( \71864 , \71863 );
buf \U$71897 ( \71865 , \71864 );
not \U$71898 ( \71866 , \71865 );
buf \U$71899 ( \71867 , \71635 );
not \U$71900 ( \71868 , \71867 );
buf \U$71901 ( \71869 , \71868 );
buf \U$71902 ( \71870 , \71869 );
not \U$71903 ( \71871 , \71870 );
or \U$71904 ( \71872 , \71866 , \71871 );
buf \U$71905 ( \71873 , \71864 );
buf \U$71906 ( \71874 , \71869 );
or \U$71907 ( \71875 , \71873 , \71874 );
buf \U$71908 ( \71876 , \71666 );
nand \U$71909 ( \71877 , \71875 , \71876 );
buf \U$71910 ( \71878 , \71877 );
buf \U$71911 ( \71879 , \71878 );
nand \U$71912 ( \71880 , \71872 , \71879 );
buf \U$71913 ( \71881 , \71880 );
buf \U$71914 ( \71882 , \71881 );
not \U$71915 ( \71883 , \71882 );
or \U$71916 ( \71884 , \71861 , \71883 );
buf \U$71917 ( \71885 , \71881 );
buf \U$71918 ( \71886 , \71859 );
or \U$71919 ( \71887 , \71885 , \71886 );
nand \U$71920 ( \71888 , \71884 , \71887 );
buf \U$71921 ( \71889 , \71888 );
buf \U$71922 ( \71890 , \71889 );
buf \U$71923 ( \71891 , \20006 );
not \U$71924 ( \71892 , \71891 );
buf \U$71925 ( \71893 , \20053 );
not \U$71926 ( \71894 , \71893 );
or \U$71927 ( \71895 , \71892 , \71894 );
buf \U$71928 ( \71896 , \20053 );
buf \U$71929 ( \71897 , \20006 );
or \U$71930 ( \71898 , \71896 , \71897 );
nand \U$71931 ( \71899 , \71895 , \71898 );
buf \U$71932 ( \71900 , \71899 );
buf \U$71933 ( \71901 , \71900 );
buf \U$71934 ( \71902 , \19923 );
and \U$71935 ( \71903 , \71901 , \71902 );
not \U$71936 ( \71904 , \71901 );
buf \U$71937 ( \71905 , \19926 );
and \U$71938 ( \71906 , \71904 , \71905 );
nor \U$71939 ( \71907 , \71903 , \71906 );
buf \U$71940 ( \71908 , \71907 );
buf \U$71941 ( \71909 , \71908 );
and \U$71942 ( \71910 , \71890 , \71909 );
not \U$71943 ( \71911 , \71890 );
buf \U$71944 ( \71912 , \71908 );
not \U$71945 ( \71913 , \71912 );
buf \U$71946 ( \71914 , \71913 );
buf \U$71947 ( \71915 , \71914 );
and \U$71948 ( \71916 , \71911 , \71915 );
nor \U$71949 ( \71917 , \71910 , \71916 );
buf \U$71950 ( \71918 , \71917 );
buf \U$71951 ( \71919 , \71918 );
not \U$71952 ( \71920 , \71919 );
buf \U$71953 ( \71921 , \71920 );
buf \U$71957 ( \71922 , \71921 );
xor \U$71958 ( \71923 , \71851 , \71922 );
buf \U$71959 ( \71924 , \71923 );
buf \U$71960 ( \71925 , \71924 );
buf \U$71961 ( \71926 , \71489 );
not \U$71962 ( \71927 , \71926 );
not \U$71963 ( \71928 , \71764 );
buf \U$71964 ( \71929 , \71928 );
not \U$71965 ( \71930 , \71929 );
or \U$71966 ( \71931 , \71927 , \71930 );
buf \U$71967 ( \71932 , \71489 );
buf \U$71968 ( \71933 , \71928 );
or \U$71969 ( \71934 , \71932 , \71933 );
buf \U$71970 ( \71935 , \71687 );
nand \U$71971 ( \71936 , \71934 , \71935 );
buf \U$71972 ( \71937 , \71936 );
buf \U$71973 ( \71938 , \71937 );
nand \U$71974 ( \71939 , \71931 , \71938 );
buf \U$71975 ( \71940 , \71939 );
buf \U$71976 ( \71941 , \71940 );
xor \U$71977 ( \71942 , \71925 , \71941 );
buf \U$71978 ( \71943 , \71747 );
buf \U$71979 ( \71944 , \71733 );
or \U$71980 ( \71945 , \71943 , \71944 );
buf \U$71981 ( \71946 , \71754 );
nand \U$71982 ( \71947 , \71945 , \71946 );
buf \U$71983 ( \71948 , \71947 );
buf \U$71984 ( \71949 , \71948 );
buf \U$71985 ( \71950 , \71733 );
buf \U$71986 ( \71951 , \71747 );
nand \U$71987 ( \71952 , \71950 , \71951 );
buf \U$71988 ( \71953 , \71952 );
buf \U$71989 ( \71954 , \71953 );
and \U$71990 ( \71955 , \71949 , \71954 );
buf \U$71991 ( \71956 , \71955 );
buf \U$71992 ( \71957 , \71956 );
buf \U$71993 ( \71958 , \71519 );
buf \U$71994 ( \71959 , \71504 );
or \U$71995 ( \71960 , \71958 , \71959 );
buf \U$71996 ( \71961 , \71528 );
nand \U$71997 ( \71962 , \71960 , \71961 );
buf \U$71998 ( \71963 , \71962 );
buf \U$71999 ( \71964 , \71963 );
buf \U$72000 ( \71965 , \71504 );
buf \U$72001 ( \71966 , \71519 );
nand \U$72002 ( \71967 , \71965 , \71966 );
buf \U$72003 ( \71968 , \71967 );
buf \U$72004 ( \71969 , \71968 );
nand \U$72005 ( \71970 , \71964 , \71969 );
buf \U$72006 ( \71971 , \71970 );
buf \U$72007 ( \71972 , \71971 );
xor \U$72008 ( \71973 , \71696 , \71711 );
and \U$72009 ( \71974 , \71973 , \71731 );
and \U$72010 ( \71975 , \71696 , \71711 );
or \U$72011 ( \71976 , \71974 , \71975 );
buf \U$72012 ( \71977 , \71976 );
buf \U$72013 ( \71978 , \71977 );
xor \U$72014 ( \71979 , \71972 , \71978 );
xor \U$72015 ( \71980 , \18038 , \18047 );
xor \U$72016 ( \71981 , \71980 , \18248 );
buf \U$72017 ( \71982 , \71981 );
buf \U$72018 ( \71983 , \71982 );
buf \U$72019 ( \71984 , \71563 );
not \U$72020 ( \71985 , \71984 );
buf \U$72021 ( \71986 , \71594 );
not \U$72022 ( \71987 , \71986 );
or \U$72023 ( \71988 , \71985 , \71987 );
buf \U$72024 ( \71989 , \71594 );
buf \U$72025 ( \71990 , \71563 );
or \U$72026 ( \71991 , \71989 , \71990 );
buf \U$72027 ( \71992 , \71578 );
nand \U$72028 ( \71993 , \71991 , \71992 );
buf \U$72029 ( \71994 , \71993 );
buf \U$72030 ( \71995 , \71994 );
nand \U$72031 ( \71996 , \71988 , \71995 );
buf \U$72032 ( \71997 , \71996 );
buf \U$72033 ( \71998 , \71997 );
xor \U$72034 ( \71999 , \71983 , \71998 );
buf \U$72035 ( \72000 , \19514 );
not \U$72036 ( \72001 , \72000 );
buf \U$72037 ( \72002 , \19722 );
not \U$72038 ( \72003 , \72002 );
or \U$72039 ( \72004 , \72001 , \72003 );
buf \U$72040 ( \72005 , \19719 );
buf \U$72041 ( \72006 , \19517 );
nand \U$72042 ( \72007 , \72005 , \72006 );
buf \U$72043 ( \72008 , \72007 );
buf \U$72044 ( \72009 , \72008 );
nand \U$72045 ( \72010 , \72004 , \72009 );
buf \U$72046 ( \72011 , \72010 );
buf \U$72047 ( \72012 , \72011 );
buf \U$72048 ( \72013 , \19727 );
xor \U$72049 ( \72014 , \72012 , \72013 );
buf \U$72050 ( \72015 , \72014 );
buf \U$72051 ( \72016 , \72015 );
xnor \U$72052 ( \72017 , \71999 , \72016 );
buf \U$72053 ( \72018 , \72017 );
buf \U$72054 ( \72019 , \72018 );
not \U$72055 ( \72020 , \72019 );
buf \U$72056 ( \72021 , \72020 );
buf \U$72057 ( \72022 , \72021 );
xnor \U$72058 ( \72023 , \71979 , \72022 );
buf \U$72059 ( \72024 , \72023 );
buf \U$72060 ( \72025 , \72024 );
xor \U$72061 ( \72026 , \71957 , \72025 );
xor \U$72062 ( \72027 , \71532 , \71538 );
and \U$72063 ( \72028 , \72027 , \71678 );
and \U$72064 ( \72029 , \71532 , \71538 );
or \U$72065 ( \72030 , \72028 , \72029 );
buf \U$72066 ( \72031 , \72030 );
buf \U$72067 ( \72032 , \72031 );
not \U$72068 ( \72033 , \72032 );
buf \U$72069 ( \72034 , \72033 );
buf \U$72070 ( \72035 , \72034 );
xor \U$72071 ( \72036 , \72026 , \72035 );
buf \U$72072 ( \72037 , \72036 );
buf \U$72073 ( \72038 , \72037 );
not \U$72074 ( \72039 , \72038 );
buf \U$72075 ( \72040 , \72039 );
buf \U$72076 ( \72041 , \72040 );
xnor \U$72077 ( \72042 , \71942 , \72041 );
buf \U$72078 ( \72043 , \72042 );
buf \U$72079 ( \72044 , \72043 );
buf \U$72080 ( \72045 , \71784 );
buf \U$72081 ( \72046 , \71680 );
not \U$72082 ( \72047 , \72046 );
buf \U$72083 ( \72048 , \71775 );
buf \U$72084 ( \72049 , \71489 );
xnor \U$72085 ( \72050 , \72048 , \72049 );
buf \U$72086 ( \72051 , \72050 );
buf \U$72087 ( \72052 , \72051 );
nand \U$72088 ( \72053 , \72047 , \72052 );
buf \U$72089 ( \72054 , \72053 );
buf \U$72090 ( \72055 , \72054 );
nand \U$72091 ( \72056 , \72045 , \72055 );
buf \U$72092 ( \72057 , \72056 );
buf \U$72093 ( \72058 , \72057 );
buf \U$72094 ( \72059 , \72051 );
not \U$72095 ( \72060 , \72059 );
buf \U$72096 ( \72061 , \71680 );
nand \U$72097 ( \72062 , \72060 , \72061 );
buf \U$72098 ( \72063 , \72062 );
buf \U$72099 ( \72064 , \72063 );
nand \U$72100 ( \72065 , \72044 , \72058 , \72064 );
buf \U$72101 ( \72066 , \72065 );
buf \U$72102 ( \72067 , \72066 );
xor \U$72103 ( \72068 , \68805 , \68891 );
and \U$72104 ( \72069 , \72068 , \69770 );
and \U$72105 ( \72070 , \68805 , \68891 );
or \U$72106 ( \72071 , \72069 , \72070 );
buf \U$72107 ( \72072 , \72071 );
buf \U$72108 ( \72073 , \72072 );
not \U$72109 ( \72074 , \72073 );
buf \U$72110 ( \72075 , \71436 );
buf \U$72111 ( \72076 , \71457 );
xor \U$72112 ( \72077 , \72075 , \72076 );
buf \U$72113 ( \72078 , \71464 );
xnor \U$72114 ( \72079 , \72077 , \72078 );
buf \U$72115 ( \72080 , \72079 );
buf \U$72116 ( \72081 , \72080 );
nand \U$72117 ( \72082 , \72074 , \72081 );
buf \U$72118 ( \72083 , \72082 );
buf \U$72119 ( \72084 , \72083 );
and \U$72120 ( \72085 , \71475 , \71806 , \72067 , \72084 );
buf \U$72121 ( \72086 , \72085 );
buf \U$72124 ( \72087 , \72086 );
buf \U$72125 ( \72088 , \72087 );
buf \U$72126 ( \72089 , \19824 );
not \U$72127 ( \72090 , \72089 );
buf \U$72128 ( \72091 , \19853 );
not \U$72129 ( \72092 , \72091 );
or \U$72130 ( \72093 , \72090 , \72092 );
buf \U$72131 ( \72094 , \19853 );
not \U$72132 ( \72095 , \72094 );
buf \U$72133 ( \72096 , \19862 );
nand \U$72134 ( \72097 , \72095 , \72096 );
buf \U$72135 ( \72098 , \72097 );
buf \U$72136 ( \72099 , \72098 );
nand \U$72137 ( \72100 , \72093 , \72099 );
buf \U$72138 ( \72101 , \72100 );
buf \U$72139 ( \72102 , \72101 );
buf \U$72143 ( \72103 , \19847 );
xor \U$72144 ( \72104 , \72102 , \72103 );
buf \U$72145 ( \72105 , \72104 );
buf \U$72146 ( \72106 , \72105 );
not \U$72147 ( \72107 , \72106 );
xor \U$72148 ( \72108 , \71812 , \71816 );
and \U$72149 ( \72109 , \72108 , \71821 );
and \U$72150 ( \72110 , \71812 , \71816 );
or \U$72151 ( \72111 , \72109 , \72110 );
buf \U$72152 ( \72112 , \72111 );
buf \U$72153 ( \72113 , \72112 );
not \U$72154 ( \72114 , \72113 );
or \U$72155 ( \72115 , \72107 , \72114 );
buf \U$72156 ( \72116 , \72112 );
buf \U$72157 ( \72117 , \72105 );
or \U$72158 ( \72118 , \72116 , \72117 );
nand \U$72159 ( \72119 , \72115 , \72118 );
buf \U$72160 ( \72120 , \72119 );
buf \U$72161 ( \72121 , \72120 );
not \U$72162 ( \72122 , \72121 );
xor \U$72163 ( \72123 , \19902 , \20056 );
xor \U$72164 ( \72124 , \72123 , \20306 );
buf \U$72165 ( \72125 , \72124 );
buf \U$72166 ( \72126 , \72125 );
not \U$72167 ( \72127 , \72126 );
buf \U$72168 ( \72128 , \72127 );
buf \U$72169 ( \72129 , \72128 );
not \U$72170 ( \72130 , \72129 );
and \U$72171 ( \72131 , \72122 , \72130 );
buf \U$72172 ( \72132 , \72120 );
buf \U$72173 ( \72133 , \72128 );
and \U$72174 ( \72134 , \72132 , \72133 );
nor \U$72175 ( \72135 , \72131 , \72134 );
buf \U$72176 ( \72136 , \72135 );
buf \U$72177 ( \72137 , \72136 );
xor \U$72178 ( \72138 , \71957 , \72025 );
and \U$72179 ( \72139 , \72138 , \72035 );
and \U$72180 ( \72140 , \71957 , \72025 );
or \U$72181 ( \72141 , \72139 , \72140 );
buf \U$72182 ( \72142 , \72141 );
buf \U$72183 ( \72143 , \72142 );
and \U$72184 ( \72144 , \72137 , \72143 );
buf \U$72185 ( \72145 , \72144 );
buf \U$72186 ( \72146 , \72145 );
buf \U$72187 ( \72147 , \71971 );
not \U$72188 ( \72148 , \72147 );
buf \U$72189 ( \72149 , \72148 );
buf \U$72190 ( \72150 , \72149 );
not \U$72191 ( \72151 , \72150 );
buf \U$72192 ( \72152 , \72018 );
not \U$72193 ( \72153 , \72152 );
or \U$72194 ( \72154 , \72151 , \72153 );
buf \U$72195 ( \72155 , \71977 );
nand \U$72196 ( \72156 , \72154 , \72155 );
buf \U$72197 ( \72157 , \72156 );
buf \U$72198 ( \72158 , \72157 );
buf \U$72199 ( \72159 , \72149 );
not \U$72200 ( \72160 , \72159 );
buf \U$72201 ( \72161 , \72021 );
nand \U$72202 ( \72162 , \72160 , \72161 );
buf \U$72203 ( \72163 , \72162 );
buf \U$72204 ( \72164 , \72163 );
nand \U$72205 ( \72165 , \72158 , \72164 );
buf \U$72206 ( \72166 , \72165 );
buf \U$72207 ( \72167 , \72166 );
not \U$72208 ( \72168 , \71921 );
not \U$72209 ( \72169 , \71840 );
or \U$72210 ( \72170 , \72168 , \72169 );
not \U$72211 ( \72171 , \71918 );
not \U$72212 ( \72172 , \71846 );
or \U$72213 ( \72173 , \72171 , \72172 );
nand \U$72214 ( \72174 , \72173 , \71823 );
nand \U$72215 ( \72175 , \72170 , \72174 );
buf \U$72216 ( \72176 , \72175 );
xor \U$72217 ( \72177 , \72167 , \72176 );
buf \U$72218 ( \72178 , \71997 );
buf \U$72219 ( \72179 , \71982 );
or \U$72220 ( \72180 , \72178 , \72179 );
buf \U$72221 ( \72181 , \72015 );
nand \U$72222 ( \72182 , \72180 , \72181 );
buf \U$72223 ( \72183 , \72182 );
buf \U$72224 ( \72184 , \72183 );
buf \U$72225 ( \72185 , \71997 );
buf \U$72226 ( \72186 , \71982 );
nand \U$72227 ( \72187 , \72185 , \72186 );
buf \U$72228 ( \72188 , \72187 );
buf \U$72229 ( \72189 , \72188 );
nand \U$72230 ( \72190 , \72184 , \72189 );
buf \U$72231 ( \72191 , \72190 );
buf \U$72232 ( \72192 , \72191 );
buf \U$72233 ( \72193 , \71856 );
not \U$72234 ( \72194 , \72193 );
buf \U$72235 ( \72195 , \71914 );
not \U$72236 ( \72196 , \72195 );
or \U$72237 ( \72197 , \72194 , \72196 );
buf \U$72238 ( \72198 , \71859 );
not \U$72239 ( \72199 , \72198 );
buf \U$72240 ( \72200 , \71908 );
not \U$72241 ( \72201 , \72200 );
or \U$72242 ( \72202 , \72199 , \72201 );
buf \U$72243 ( \72203 , \71881 );
nand \U$72244 ( \72204 , \72202 , \72203 );
buf \U$72245 ( \72205 , \72204 );
buf \U$72246 ( \72206 , \72205 );
nand \U$72247 ( \72207 , \72197 , \72206 );
buf \U$72248 ( \72208 , \72207 );
buf \U$72249 ( \72209 , \72208 );
xor \U$72250 ( \72210 , \72192 , \72209 );
xor \U$72251 ( \72211 , \19739 , \19756 );
xor \U$72252 ( \72212 , \72211 , \19813 );
buf \U$72253 ( \72213 , \72212 );
buf \U$72254 ( \72214 , \72213 );
xor \U$72255 ( \72215 , \72210 , \72214 );
buf \U$72256 ( \72216 , \72215 );
buf \U$72257 ( \72217 , \72216 );
xor \U$72258 ( \72218 , \72177 , \72217 );
buf \U$72259 ( \72219 , \72218 );
buf \U$72260 ( \72220 , \72219 );
not \U$72261 ( \72221 , \72220 );
buf \U$72262 ( \72222 , \72221 );
buf \U$72263 ( \72223 , \72222 );
or \U$72264 ( \72224 , \72146 , \72223 );
buf \U$72265 ( \72225 , \72142 );
buf \U$72266 ( \72226 , \72136 );
or \U$72267 ( \72227 , \72225 , \72226 );
buf \U$72268 ( \72228 , \72227 );
buf \U$72269 ( \72229 , \72228 );
nand \U$72270 ( \72230 , \72224 , \72229 );
buf \U$72271 ( \72231 , \72230 );
buf \U$72272 ( \72232 , \72231 );
not \U$72273 ( \72233 , \72232 );
xor \U$72274 ( \72234 , \20310 , \20323 );
xnor \U$72275 ( \72235 , \72234 , \20315 );
buf \U$72276 ( \72236 , \72235 );
xor \U$72277 ( \72237 , \72167 , \72176 );
and \U$72278 ( \72238 , \72237 , \72217 );
and \U$72279 ( \72239 , \72167 , \72176 );
or \U$72280 ( \72240 , \72238 , \72239 );
buf \U$72281 ( \72241 , \72240 );
buf \U$72282 ( \72242 , \72241 );
not \U$72283 ( \72243 , \72242 );
buf \U$72284 ( \72244 , \72243 );
buf \U$72285 ( \72245 , \72244 );
xor \U$72286 ( \72246 , \72236 , \72245 );
buf \U$72287 ( \72247 , \72246 );
buf \U$72288 ( \72248 , \72247 );
xor \U$72289 ( \72249 , \72192 , \72209 );
and \U$72290 ( \72250 , \72249 , \72214 );
and \U$72291 ( \72251 , \72192 , \72209 );
or \U$72292 ( \72252 , \72250 , \72251 );
buf \U$72293 ( \72253 , \72252 );
buf \U$72294 ( \72254 , \72253 );
not \U$72295 ( \72255 , \72254 );
buf \U$72296 ( \72256 , \72255 );
buf \U$72297 ( \72257 , \72256 );
not \U$72298 ( \72258 , \72257 );
xor \U$72299 ( \72259 , \19868 , \19817 );
buf \U$72300 ( \72260 , \72259 );
buf \U$72301 ( \72261 , \19873 );
not \U$72302 ( \72262 , \72261 );
buf \U$72303 ( \72263 , \72262 );
buf \U$72304 ( \72264 , \72263 );
and \U$72305 ( \72265 , \72260 , \72264 );
not \U$72306 ( \72266 , \72260 );
buf \U$72307 ( \72267 , \19873 );
and \U$72308 ( \72268 , \72266 , \72267 );
nor \U$72309 ( \72269 , \72265 , \72268 );
buf \U$72310 ( \72270 , \72269 );
buf \U$72311 ( \72271 , \72270 );
not \U$72312 ( \72272 , \72271 );
buf \U$72313 ( \72273 , \72272 );
buf \U$72314 ( \72274 , \72273 );
not \U$72315 ( \72275 , \72274 );
or \U$72316 ( \72276 , \72258 , \72275 );
buf \U$72317 ( \72277 , \72270 );
buf \U$72318 ( \72278 , \72253 );
nand \U$72319 ( \72279 , \72277 , \72278 );
buf \U$72320 ( \72280 , \72279 );
buf \U$72321 ( \72281 , \72280 );
nand \U$72322 ( \72282 , \72276 , \72281 );
buf \U$72323 ( \72283 , \72282 );
buf \U$72324 ( \72284 , \72283 );
buf \U$72325 ( \72285 , \72105 );
not \U$72326 ( \72286 , \72285 );
buf \U$72327 ( \72287 , \72286 );
buf \U$72328 ( \72288 , \72287 );
not \U$72329 ( \72289 , \72288 );
buf \U$72330 ( \72290 , \72112 );
not \U$72331 ( \72291 , \72290 );
or \U$72332 ( \72292 , \72289 , \72291 );
buf \U$72333 ( \72293 , \72287 );
buf \U$72334 ( \72294 , \72112 );
or \U$72335 ( \72295 , \72293 , \72294 );
buf \U$72336 ( \72296 , \72125 );
nand \U$72337 ( \72297 , \72295 , \72296 );
buf \U$72338 ( \72298 , \72297 );
buf \U$72339 ( \72299 , \72298 );
nand \U$72340 ( \72300 , \72292 , \72299 );
buf \U$72341 ( \72301 , \72300 );
buf \U$72342 ( \72302 , \72301 );
not \U$72343 ( \72303 , \72302 );
buf \U$72344 ( \72304 , \72303 );
buf \U$72345 ( \72305 , \72304 );
and \U$72346 ( \72306 , \72284 , \72305 );
not \U$72347 ( \72307 , \72284 );
buf \U$72348 ( \72308 , \72301 );
and \U$72349 ( \72309 , \72307 , \72308 );
nor \U$72350 ( \72310 , \72306 , \72309 );
buf \U$72351 ( \72311 , \72310 );
buf \U$72352 ( \72312 , \72311 );
xor \U$72353 ( \72313 , \72248 , \72312 );
buf \U$72354 ( \72314 , \72313 );
buf \U$72355 ( \72315 , \72314 );
nand \U$72356 ( \72316 , \72233 , \72315 );
buf \U$72357 ( \72317 , \72316 );
buf \U$72358 ( \72318 , \72317 );
buf \U$72359 ( \72319 , \71924 );
not \U$72360 ( \72320 , \72319 );
buf \U$72361 ( \72321 , \72320 );
buf \U$72362 ( \72322 , \72321 );
not \U$72363 ( \72323 , \72322 );
buf \U$72364 ( \72324 , \72037 );
not \U$72365 ( \72325 , \72324 );
or \U$72366 ( \72326 , \72323 , \72325 );
buf \U$72367 ( \72327 , \71940 );
nand \U$72368 ( \72328 , \72326 , \72327 );
buf \U$72369 ( \72329 , \72328 );
buf \U$72370 ( \72330 , \72329 );
buf \U$72371 ( \72331 , \72040 );
buf \U$72372 ( \72332 , \71924 );
nand \U$72373 ( \72333 , \72331 , \72332 );
buf \U$72374 ( \72334 , \72333 );
buf \U$72375 ( \72335 , \72334 );
nand \U$72376 ( \72336 , \72330 , \72335 );
buf \U$72377 ( \72337 , \72336 );
buf \U$72378 ( \72338 , \72337 );
not \U$72379 ( \72339 , \72338 );
xor \U$72380 ( \72340 , \72137 , \72143 );
buf \U$72381 ( \72341 , \72340 );
buf \U$72382 ( \72342 , \72341 );
buf \U$72383 ( \72343 , \72222 );
and \U$72384 ( \72344 , \72342 , \72343 );
not \U$72385 ( \72345 , \72342 );
buf \U$72386 ( \72346 , \72219 );
and \U$72387 ( \72347 , \72345 , \72346 );
nor \U$72388 ( \72348 , \72344 , \72347 );
buf \U$72389 ( \72349 , \72348 );
buf \U$72390 ( \72350 , \72349 );
nand \U$72391 ( \72351 , \72339 , \72350 );
buf \U$72392 ( \72352 , \72351 );
buf \U$72393 ( \72353 , \72352 );
and \U$72394 ( \72354 , \72318 , \72353 );
buf \U$72395 ( \72355 , \72354 );
buf \U$72398 ( \72356 , \72355 );
buf \U$72399 ( \72357 , \72356 );
and \U$72400 ( \72358 , \72236 , \72245 );
buf \U$72401 ( \72359 , \72358 );
buf \U$72402 ( \72360 , \72359 );
buf \U$72403 ( \72361 , \72311 );
or \U$72404 ( \72362 , \72360 , \72361 );
buf \U$72405 ( \72363 , \72235 );
not \U$72406 ( \72364 , \72363 );
buf \U$72407 ( \72365 , \72241 );
nand \U$72408 ( \72366 , \72364 , \72365 );
buf \U$72409 ( \72367 , \72366 );
buf \U$72410 ( \72368 , \72367 );
nand \U$72411 ( \72369 , \72362 , \72368 );
buf \U$72412 ( \72370 , \72369 );
buf \U$72413 ( \72371 , \72370 );
not \U$72414 ( \72372 , \72371 );
xor \U$72415 ( \72373 , \17945 , \18571 );
xor \U$72416 ( \72374 , \72373 , \18830 );
buf \U$72417 ( \72375 , \72374 );
buf \U$72418 ( \72376 , \19887 );
not \U$72419 ( \72377 , \72376 );
buf \U$72420 ( \72378 , \19892 );
not \U$72421 ( \72379 , \72378 );
or \U$72422 ( \72380 , \72377 , \72379 );
buf \U$72423 ( \72381 , \19887 );
buf \U$72424 ( \72382 , \19892 );
or \U$72425 ( \72383 , \72381 , \72382 );
nand \U$72426 ( \72384 , \72380 , \72383 );
buf \U$72427 ( \72385 , \72384 );
buf \U$72428 ( \72386 , \72385 );
buf \U$72429 ( \72387 , \20329 );
not \U$72430 ( \72388 , \72387 );
buf \U$72431 ( \72389 , \72388 );
buf \U$72432 ( \72390 , \72389 );
and \U$72433 ( \72391 , \72386 , \72390 );
not \U$72434 ( \72392 , \72386 );
buf \U$72435 ( \72393 , \20329 );
and \U$72436 ( \72394 , \72392 , \72393 );
nor \U$72437 ( \72395 , \72391 , \72394 );
buf \U$72438 ( \72396 , \72395 );
xor \U$72439 ( \72397 , \72375 , \72396 );
buf \U$72440 ( \72398 , \72253 );
not \U$72441 ( \72399 , \72398 );
buf \U$72442 ( \72400 , \72301 );
not \U$72443 ( \72401 , \72400 );
or \U$72444 ( \72402 , \72399 , \72401 );
buf \U$72445 ( \72403 , \72256 );
not \U$72446 ( \72404 , \72403 );
buf \U$72447 ( \72405 , \72304 );
not \U$72448 ( \72406 , \72405 );
or \U$72449 ( \72407 , \72404 , \72406 );
buf \U$72450 ( \72408 , \72270 );
not \U$72451 ( \72409 , \72408 );
buf \U$72452 ( \72410 , \72409 );
buf \U$72453 ( \72411 , \72410 );
nand \U$72454 ( \72412 , \72407 , \72411 );
buf \U$72455 ( \72413 , \72412 );
buf \U$72456 ( \72414 , \72413 );
nand \U$72457 ( \72415 , \72402 , \72414 );
buf \U$72458 ( \72416 , \72415 );
xor \U$72459 ( \72417 , \72397 , \72416 );
buf \U$72460 ( \72418 , \72417 );
nand \U$72461 ( \72419 , \72372 , \72418 );
buf \U$72462 ( \72420 , \72419 );
buf \U$72463 ( \72421 , \72420 );
not \U$72464 ( \72422 , \72375 );
nand \U$72465 ( \72423 , \72422 , \72396 );
not \U$72466 ( \72424 , \72423 );
not \U$72467 ( \72425 , \72416 );
or \U$72468 ( \72426 , \72424 , \72425 );
buf \U$72469 ( \72427 , \72396 );
not \U$72470 ( \72428 , \72427 );
buf \U$72471 ( \72429 , \72375 );
nand \U$72472 ( \72430 , \72428 , \72429 );
buf \U$72473 ( \72431 , \72430 );
nand \U$72474 ( \72432 , \72426 , \72431 );
buf \U$72475 ( \72433 , \72432 );
not \U$72476 ( \72434 , \72433 );
buf \U$72477 ( \72435 , \19307 );
buf \U$72478 ( \72436 , \20352 );
xor \U$72479 ( \72437 , \72435 , \72436 );
buf \U$72480 ( \72438 , \20346 );
xor \U$72481 ( \72439 , \72437 , \72438 );
buf \U$72482 ( \72440 , \72439 );
buf \U$72483 ( \72441 , \72440 );
nand \U$72484 ( \72442 , \72434 , \72441 );
buf \U$72485 ( \72443 , \72442 );
buf \U$72486 ( \72444 , \72443 );
nand \U$72487 ( \72445 , \72421 , \72444 );
buf \U$72488 ( \72446 , \72445 );
buf \U$72489 ( \72447 , \72446 );
not \U$72490 ( \72448 , \72447 );
buf \U$72491 ( \72449 , \72448 );
buf \U$72492 ( \72450 , \72449 );
and \U$72493 ( \72451 , \70067 , \72088 , \72357 , \72450 );
buf \U$72494 ( \72452 , \72451 );
buf \U$72495 ( \72453 , \72452 );
not \U$72496 ( \72454 , \72453 );
or \U$72497 ( \72455 , \63021 , \72454 );
buf \U$72498 ( \72456 , \72086 );
buf \U$72499 ( \72457 , \72355 );
buf \U$72500 ( \72458 , \72449 );
and \U$72501 ( \72459 , \72456 , \72457 , \72458 );
buf \U$72502 ( \72460 , \72459 );
buf \U$72503 ( \72461 , \72460 );
not \U$72504 ( \72462 , \72461 );
buf \U$72505 ( \72463 , \67805 );
buf \U$72506 ( \72464 , \69817 );
nand \U$72507 ( \72465 , \72463 , \72464 );
buf \U$72508 ( \72466 , \72465 );
buf \U$72509 ( \72467 , \72466 );
buf \U$72510 ( \72468 , \69968 );
buf \U$72511 ( \72469 , \70007 );
nor \U$72512 ( \72470 , \72468 , \72469 );
buf \U$72513 ( \72471 , \72470 );
buf \U$72514 ( \72472 , \72471 );
buf \U$72515 ( \72473 , \69842 );
buf \U$72516 ( \72474 , \69958 );
nor \U$72517 ( \72475 , \72473 , \72474 );
buf \U$72518 ( \72476 , \72475 );
buf \U$72519 ( \72477 , \72476 );
nor \U$72520 ( \72478 , \72472 , \72477 );
buf \U$72521 ( \72479 , \72478 );
buf \U$72522 ( \72480 , \72479 );
not \U$72523 ( \72481 , \72480 );
buf \U$72524 ( \72482 , \70038 );
buf \U$72525 ( \72483 , \70033 );
nand \U$72526 ( \72484 , \72482 , \72483 );
buf \U$72527 ( \72485 , \72484 );
buf \U$72528 ( \72486 , \72485 );
buf \U$72529 ( \72487 , \70048 );
buf \U$72530 ( \72488 , \70054 );
nand \U$72531 ( \72489 , \72487 , \72488 );
buf \U$72532 ( \72490 , \72489 );
buf \U$72533 ( \72491 , \72490 );
nand \U$72534 ( \72492 , \72486 , \72491 );
buf \U$72535 ( \72493 , \72492 );
buf \U$72536 ( \72494 , \72493 );
buf \U$72537 ( \72495 , \70010 );
buf \U$72538 ( \72496 , \70044 );
nand \U$72539 ( \72497 , \72494 , \72495 , \72496 );
buf \U$72540 ( \72498 , \72497 );
buf \U$72541 ( \72499 , \72498 );
not \U$72542 ( \72500 , \72499 );
or \U$72543 ( \72501 , \72481 , \72500 );
buf \U$72544 ( \72502 , \69961 );
nand \U$72545 ( \72503 , \72501 , \72502 );
buf \U$72546 ( \72504 , \72503 );
buf \U$72547 ( \72505 , \72504 );
or \U$72548 ( \72506 , \72467 , \72505 );
buf \U$72549 ( \72507 , \67601 );
buf \U$72550 ( \72508 , \67799 );
nand \U$72551 ( \72509 , \72507 , \72508 );
buf \U$72552 ( \72510 , \72509 );
buf \U$72553 ( \72511 , \72510 );
buf \U$72554 ( \72512 , \66737 );
buf \U$72555 ( \72513 , \67591 );
nand \U$72556 ( \72514 , \72512 , \72513 );
buf \U$72557 ( \72515 , \72514 );
buf \U$72558 ( \72516 , \72515 );
and \U$72559 ( \72517 , \72511 , \72516 );
buf \U$72560 ( \72518 , \72517 );
buf \U$72561 ( \72519 , \72518 );
buf \U$72562 ( \72520 , \67597 );
buf \U$72563 ( \72521 , \69814 );
nand \U$72564 ( \72522 , \72520 , \72521 );
buf \U$72565 ( \72523 , \72522 );
buf \U$72566 ( \72524 , \72523 );
or \U$72567 ( \72525 , \72519 , \72524 );
buf \U$72568 ( \72526 , \69772 );
buf \U$72569 ( \72527 , \69792 );
nand \U$72570 ( \72528 , \72526 , \72527 );
buf \U$72571 ( \72529 , \72528 );
buf \U$72572 ( \72530 , \72529 );
buf \U$72573 ( \72531 , \69799 );
buf \U$72574 ( \72532 , \69808 );
nand \U$72575 ( \72533 , \72531 , \72532 );
buf \U$72576 ( \72534 , \72533 );
buf \U$72577 ( \72535 , \72534 );
and \U$72578 ( \72536 , \72530 , \72535 );
buf \U$72579 ( \72537 , \72536 );
buf \U$72580 ( \72538 , \72537 );
nand \U$72581 ( \72539 , \72525 , \72538 );
buf \U$72582 ( \72540 , \72539 );
buf \U$72583 ( \72541 , \72540 );
buf \U$72584 ( \72542 , \69795 );
buf \U$72585 ( \72543 , \72542 );
nand \U$72586 ( \72544 , \72541 , \72543 );
buf \U$72587 ( \72545 , \72544 );
buf \U$72588 ( \72546 , \72545 );
nand \U$72589 ( \72547 , \72506 , \72546 );
buf \U$72590 ( \72548 , \72547 );
buf \U$72591 ( \72549 , \72548 );
not \U$72592 ( \72550 , \72549 );
or \U$72593 ( \72551 , \72462 , \72550 );
not \U$72594 ( \72552 , \72314 );
buf \U$72595 ( \72553 , \72552 );
buf \U$72597 ( \72554 , \72231 );
nand \U$72598 ( \72555 , \72553 , \72554 );
buf \U$72599 ( \72556 , \72555 );
not \U$72600 ( \72557 , \72556 );
buf \U$72601 ( \72558 , \72349 );
not \U$72602 ( \72559 , \72558 );
buf \U$72603 ( \72560 , \72559 );
buf \U$72604 ( \72561 , \72560 );
buf \U$72605 ( \72562 , \72337 );
nand \U$72606 ( \72563 , \72561 , \72562 );
buf \U$72607 ( \72564 , \72563 );
not \U$72608 ( \72565 , \72564 );
or \U$72609 ( \72566 , \72557 , \72565 );
nand \U$72610 ( \72567 , \72566 , \72317 );
buf \U$72611 ( \72568 , \72567 );
buf \U$72612 ( \72569 , \72420 );
not \U$72613 ( \72570 , \72569 );
buf \U$72614 ( \72571 , \72570 );
buf \U$72615 ( \72572 , \72571 );
or \U$72616 ( \72573 , \72568 , \72572 );
buf \U$72617 ( \72574 , \72417 );
not \U$72618 ( \72575 , \72574 );
buf \U$72619 ( \72576 , \72370 );
nand \U$72620 ( \72577 , \72575 , \72576 );
buf \U$72621 ( \72578 , \72577 );
buf \U$72622 ( \72579 , \72578 );
nand \U$72623 ( \72580 , \72573 , \72579 );
buf \U$72624 ( \72581 , \72580 );
buf \U$72625 ( \72582 , \72581 );
buf \U$72628 ( \72583 , \72443 );
buf \U$72629 ( \72584 , \72583 );
and \U$72630 ( \72585 , \72582 , \72584 );
buf \U$72631 ( \72586 , \72355 );
buf \U$72632 ( \72587 , \72446 );
not \U$72633 ( \72588 , \72587 );
buf \U$72634 ( \72589 , \72588 );
buf \U$72635 ( \72590 , \72589 );
and \U$72636 ( \72591 , \72057 , \72063 );
nor \U$72637 ( \72592 , \72591 , \72043 );
buf \U$72638 ( \72593 , \72592 );
nand \U$72639 ( \72594 , \72586 , \72590 , \72593 );
buf \U$72640 ( \72595 , \72594 );
buf \U$72641 ( \72596 , \72595 );
buf \U$72642 ( \72597 , \72440 );
not \U$72643 ( \72598 , \72597 );
buf \U$72644 ( \72599 , \72432 );
nand \U$72645 ( \72600 , \72598 , \72599 );
buf \U$72646 ( \72601 , \72600 );
buf \U$72647 ( \72602 , \72601 );
nand \U$72648 ( \72603 , \72596 , \72602 );
buf \U$72649 ( \72604 , \72603 );
buf \U$72650 ( \72605 , \72604 );
nor \U$72651 ( \72606 , \72585 , \72605 );
buf \U$72652 ( \72607 , \72606 );
buf \U$72653 ( \72608 , \72607 );
nand \U$72654 ( \72609 , \72551 , \72608 );
buf \U$72655 ( \72610 , \72609 );
buf \U$72656 ( \72611 , \72610 );
buf \U$72657 ( \72612 , \72356 );
buf \U$72658 ( \72613 , \72449 );
nand \U$72659 ( \72614 , \72612 , \72613 );
buf \U$72660 ( \72615 , \72614 );
buf \U$72661 ( \72616 , \72615 );
buf \U$72662 ( \72617 , \71474 );
buf \U$72663 ( \72618 , \71468 );
buf \U$72664 ( \72619 , \71429 );
nand \U$72665 ( \72620 , \72618 , \72619 );
buf \U$72666 ( \72621 , \72620 );
buf \U$72667 ( \72622 , \72621 );
buf \U$72668 ( \72623 , \72080 );
not \U$72669 ( \72624 , \72623 );
buf \U$72670 ( \72625 , \72072 );
nand \U$72671 ( \72626 , \72624 , \72625 );
buf \U$72672 ( \72627 , \72626 );
buf \U$72673 ( \72628 , \72627 );
nand \U$72674 ( \72629 , \72622 , \72628 );
buf \U$72675 ( \72630 , \72629 );
buf \U$72676 ( \72631 , \72630 );
nand \U$72677 ( \72632 , \72617 , \72631 );
buf \U$72678 ( \72633 , \72632 );
buf \U$72679 ( \72634 , \72633 );
buf \U$72680 ( \72635 , \71805 );
not \U$72681 ( \72636 , \72635 );
buf \U$72682 ( \72637 , \72636 );
buf \U$72683 ( \72638 , \72637 );
or \U$72684 ( \72639 , \72634 , \72638 );
buf \U$72685 ( \72640 , \71787 );
buf \U$72686 ( \72641 , \71802 );
or \U$72687 ( \72642 , \72640 , \72641 );
buf \U$72688 ( \72643 , \72642 );
buf \U$72689 ( \72644 , \72643 );
nand \U$72690 ( \72645 , \72639 , \72644 );
buf \U$72691 ( \72646 , \72645 );
buf \U$72692 ( \72647 , \72646 );
buf \U$72695 ( \72648 , \72066 );
buf \U$72696 ( \72649 , \72648 );
nand \U$72697 ( \72650 , \72647 , \72649 );
buf \U$72698 ( \72651 , \72650 );
buf \U$72699 ( \72652 , \72651 );
nor \U$72700 ( \72653 , \72616 , \72652 );
buf \U$72701 ( \72654 , \72653 );
buf \U$72702 ( \72655 , \72654 );
nor \U$72703 ( \72656 , \72611 , \72655 );
buf \U$72704 ( \72657 , \72656 );
buf \U$72705 ( \72658 , \72657 );
nand \U$72706 ( \72659 , \72455 , \72658 );
buf \U$72707 ( \72660 , \72659 );
buf \U$72708 ( \72661 , \72660 );
nand \U$72709 ( \72662 , \43778 , \72661 );
buf \U$72710 ( \72663 , \72662 );
buf \U$72711 ( \72664 , \72663 );
nand \U$72712 ( \72665 , \43747 , \72664 );
buf \U$72713 ( \72666 , \72665 );
buf \U$72714 ( \72667 , \72666 );
buf \U$72715 ( \72668 , \72667 );
not \U$72716 ( \72669 , \72668 );
or \U$72717 ( \72670 , \12244 , \72669 );
buf \U$72718 ( \72671 , \11697 );
not \U$72719 ( \72672 , \72671 );
buf \U$72720 ( \72673 , \8741 );
not \U$72721 ( \72674 , \72673 );
buf \U$72722 ( \72675 , \8748 );
buf \U$72723 ( \72676 , \8754 );
and \U$72724 ( \72677 , \72675 , \72676 );
buf \U$72725 ( \72678 , \72677 );
not \U$72726 ( \72679 , \72678 );
not \U$72727 ( \72680 , \8410 );
or \U$72728 ( \72681 , \72679 , \72680 );
buf \U$72729 ( \72682 , \8387 );
buf \U$72730 ( \72683 , \8407 );
nand \U$72731 ( \72684 , \72682 , \72683 );
buf \U$72732 ( \72685 , \72684 );
nand \U$72733 ( \72686 , \72681 , \72685 );
buf \U$72734 ( \72687 , \72686 );
nand \U$72735 ( \72688 , \72674 , \72687 );
buf \U$72736 ( \72689 , \72688 );
buf \U$72737 ( \72690 , \72689 );
buf \U$72738 ( \72691 , \8732 );
buf \U$72739 ( \72692 , \8738 );
nand \U$72740 ( \72693 , \72691 , \72692 );
buf \U$72741 ( \72694 , \72693 );
buf \U$72742 ( \72695 , \72694 );
nand \U$72743 ( \72696 , \72690 , \72695 );
buf \U$72744 ( \72697 , \72696 );
not \U$72745 ( \72698 , \72697 );
not \U$72746 ( \72699 , \9026 );
or \U$72747 ( \72700 , \72698 , \72699 );
buf \U$72748 ( \72701 , \9023 );
buf \U$72749 ( \72702 , \8763 );
nand \U$72750 ( \72703 , \72701 , \72702 );
buf \U$72751 ( \72704 , \72703 );
nand \U$72752 ( \72705 , \72700 , \72704 );
buf \U$72753 ( \72706 , \72705 );
not \U$72754 ( \72707 , \72706 );
buf \U$72755 ( \72708 , \5615 );
not \U$72756 ( \72709 , \72708 );
buf \U$72757 ( \72710 , \5131 );
not \U$72758 ( \72711 , \72710 );
buf \U$72759 ( \72712 , \72711 );
buf \U$72760 ( \72713 , \72712 );
buf \U$72761 ( \72714 , \3944 );
buf \U$72762 ( \72715 , \4614 );
nand \U$72763 ( \72716 , \72714 , \72715 );
buf \U$72764 ( \72717 , \72716 );
buf \U$72765 ( \72718 , \72717 );
or \U$72766 ( \72719 , \72713 , \72718 );
buf \U$72767 ( \72720 , \5116 );
buf \U$72768 ( \72721 , \5125 );
nand \U$72769 ( \72722 , \72720 , \72721 );
buf \U$72770 ( \72723 , \72722 );
buf \U$72771 ( \72724 , \72723 );
nand \U$72772 ( \72725 , \72719 , \72724 );
buf \U$72773 ( \72726 , \72725 );
buf \U$72774 ( \72727 , \72726 );
not \U$72775 ( \72728 , \72727 );
or \U$72776 ( \72729 , \72709 , \72728 );
buf \U$72777 ( \72730 , \5606 );
buf \U$72778 ( \72731 , \5612 );
nand \U$72779 ( \72732 , \72730 , \72731 );
buf \U$72780 ( \72733 , \72732 );
buf \U$72781 ( \72734 , \72733 );
nand \U$72782 ( \72735 , \72729 , \72734 );
buf \U$72783 ( \72736 , \72735 );
not \U$72784 ( \72737 , \72736 );
buf \U$72785 ( \72738 , \6091 );
buf \U$72786 ( \72739 , \6097 );
nand \U$72787 ( \72740 , \72738 , \72739 );
buf \U$72788 ( \72741 , \72740 );
buf \U$72789 ( \72742 , \72741 );
not \U$72790 ( \72743 , \72742 );
buf \U$72791 ( \72744 , \72743 );
not \U$72792 ( \72745 , \72744 );
and \U$72793 ( \72746 , \72737 , \72745 );
not \U$72794 ( \72747 , \6100 );
nand \U$72795 ( \72748 , \72747 , \7718 );
nor \U$72796 ( \72749 , \72746 , \72748 );
buf \U$72797 ( \72750 , \72749 );
buf \U$72798 ( \72751 , \7715 );
not \U$72799 ( \72752 , \72751 );
buf \U$72800 ( \72753 , \7337 );
not \U$72801 ( \72754 , \72753 );
buf \U$72802 ( \72755 , \6937 );
not \U$72803 ( \72756 , \72755 );
buf \U$72804 ( \72757 , \6944 );
nor \U$72805 ( \72758 , \72756 , \72757 );
buf \U$72806 ( \72759 , \72758 );
not \U$72807 ( \72760 , \72759 );
not \U$72808 ( \72761 , \6931 );
or \U$72809 ( \72762 , \72760 , \72761 );
buf \U$72810 ( \72763 , \6930 );
buf \U$72811 ( \72764 , \6529 );
nand \U$72812 ( \72765 , \72763 , \72764 );
buf \U$72813 ( \72766 , \72765 );
nand \U$72814 ( \72767 , \72762 , \72766 );
buf \U$72815 ( \72768 , \72767 );
not \U$72816 ( \72769 , \72768 );
or \U$72817 ( \72770 , \72754 , \72769 );
buf \U$72818 ( \72771 , \7328 );
buf \U$72819 ( \72772 , \7334 );
nand \U$72820 ( \72773 , \72771 , \72772 );
buf \U$72821 ( \72774 , \72773 );
buf \U$72822 ( \72775 , \72774 );
nand \U$72823 ( \72776 , \72770 , \72775 );
buf \U$72824 ( \72777 , \72776 );
buf \U$72825 ( \72778 , \72777 );
not \U$72826 ( \72779 , \72778 );
or \U$72827 ( \72780 , \72752 , \72779 );
buf \U$72828 ( \72781 , \7706 );
buf \U$72829 ( \72782 , \7712 );
nand \U$72830 ( \72783 , \72781 , \72782 );
buf \U$72831 ( \72784 , \72783 );
buf \U$72832 ( \72785 , \72784 );
nand \U$72833 ( \72786 , \72780 , \72785 );
buf \U$72834 ( \72787 , \72786 );
buf \U$72835 ( \72788 , \72787 );
or \U$72836 ( \72789 , \72750 , \72788 );
buf \U$72837 ( \72790 , \9029 );
nand \U$72838 ( \72791 , \72789 , \72790 );
buf \U$72839 ( \72792 , \72791 );
buf \U$72840 ( \72793 , \72792 );
nand \U$72841 ( \72794 , \72707 , \72793 );
buf \U$72842 ( \72795 , \72794 );
buf \U$72843 ( \72796 , \72795 );
buf \U$72844 ( \72797 , \10108 );
nand \U$72845 ( \72798 , \72796 , \72797 );
buf \U$72846 ( \72799 , \72798 );
buf \U$72847 ( \72800 , \72799 );
buf \U$72848 ( \72801 , \9855 );
not \U$72849 ( \72802 , \72801 );
buf \U$72850 ( \72803 , \9586 );
buf \U$72851 ( \72804 , \9590 );
buf \U$72852 ( \72805 , \9596 );
nand \U$72853 ( \72806 , \72804 , \72805 );
buf \U$72854 ( \72807 , \72806 );
buf \U$72855 ( \72808 , \72807 );
or \U$72856 ( \72809 , \72803 , \72808 );
buf \U$72857 ( \72810 , \9583 );
buf \U$72858 ( \72811 , \9318 );
nand \U$72859 ( \72812 , \72810 , \72811 );
buf \U$72860 ( \72813 , \72812 );
buf \U$72861 ( \72814 , \72813 );
nand \U$72862 ( \72815 , \72809 , \72814 );
buf \U$72863 ( \72816 , \72815 );
buf \U$72864 ( \72817 , \72816 );
not \U$72865 ( \72818 , \72817 );
or \U$72866 ( \72819 , \72802 , \72818 );
buf \U$72867 ( \72820 , \9843 );
buf \U$72868 ( \72821 , \9852 );
nand \U$72869 ( \72822 , \72820 , \72821 );
buf \U$72870 ( \72823 , \72822 );
buf \U$72871 ( \72824 , \72823 );
nand \U$72872 ( \72825 , \72819 , \72824 );
buf \U$72873 ( \72826 , \72825 );
buf \U$72874 ( \72827 , \72826 );
buf \U$72875 ( \72828 , \10105 );
and \U$72876 ( \72829 , \72827 , \72828 );
buf \U$72877 ( \72830 , \10102 );
buf \U$72878 ( \72831 , \9867 );
and \U$72879 ( \72832 , \72830 , \72831 );
buf \U$72880 ( \72833 , \72832 );
buf \U$72881 ( \72834 , \72833 );
nor \U$72882 ( \72835 , \72829 , \72834 );
buf \U$72883 ( \72836 , \72835 );
buf \U$72884 ( \72837 , \72836 );
nand \U$72885 ( \72838 , \72800 , \72837 );
buf \U$72886 ( \72839 , \72838 );
buf \U$72887 ( \72840 , \72839 );
not \U$72888 ( \72841 , \72840 );
or \U$72889 ( \72842 , \72672 , \72841 );
buf \U$72890 ( \72843 , \10577 );
buf \U$72891 ( \72844 , \10340 );
buf \U$72892 ( \72845 , \10346 );
nand \U$72893 ( \72846 , \72844 , \72845 );
buf \U$72894 ( \72847 , \72846 );
buf \U$72895 ( \72848 , \72847 );
or \U$72896 ( \72849 , \72843 , \72848 );
buf \U$72897 ( \72850 , \10568 );
buf \U$72898 ( \72851 , \10574 );
nand \U$72899 ( \72852 , \72850 , \72851 );
buf \U$72900 ( \72853 , \72852 );
buf \U$72901 ( \72854 , \72853 );
nand \U$72902 ( \72855 , \72849 , \72854 );
buf \U$72903 ( \72856 , \72855 );
buf \U$72904 ( \72857 , \72856 );
buf \U$72905 ( \72858 , \10825 );
and \U$72906 ( \72859 , \72857 , \72858 );
buf \U$72907 ( \72860 , \10816 );
buf \U$72908 ( \72861 , \10822 );
nand \U$72909 ( \72862 , \72860 , \72861 );
buf \U$72910 ( \72863 , \72862 );
buf \U$72911 ( \72864 , \72863 );
not \U$72912 ( \72865 , \72864 );
buf \U$72913 ( \72866 , \72865 );
buf \U$72914 ( \72867 , \72866 );
nor \U$72915 ( \72868 , \72859 , \72867 );
buf \U$72916 ( \72869 , \72868 );
buf \U$72917 ( \72870 , \72869 );
buf \U$72918 ( \72871 , \11054 );
or \U$72919 ( \72872 , \72870 , \72871 );
buf \U$72920 ( \72873 , \10834 );
buf \U$72921 ( \72874 , \11051 );
nand \U$72922 ( \72875 , \72873 , \72874 );
buf \U$72923 ( \72876 , \72875 );
buf \U$72924 ( \72877 , \72876 );
nand \U$72925 ( \72878 , \72872 , \72877 );
buf \U$72926 ( \72879 , \72878 );
buf \U$72927 ( \72880 , \72879 );
buf \U$72928 ( \72881 , \11691 );
and \U$72929 ( \72882 , \72880 , \72881 );
buf \U$72930 ( \72883 , \11553 );
not \U$72931 ( \72884 , \72883 );
buf \U$72932 ( \72885 , \11531 );
buf \U$72933 ( \72886 , \11537 );
nand \U$72934 ( \72887 , \72885 , \72886 );
buf \U$72935 ( \72888 , \72887 );
buf \U$72936 ( \72889 , \72888 );
not \U$72937 ( \72890 , \72889 );
and \U$72938 ( \72891 , \72884 , \72890 );
buf \U$72939 ( \72892 , \11544 );
buf \U$72940 ( \72893 , \11550 );
and \U$72941 ( \72894 , \72892 , \72893 );
buf \U$72942 ( \72895 , \72894 );
buf \U$72943 ( \72896 , \72895 );
nor \U$72944 ( \72897 , \72891 , \72896 );
buf \U$72945 ( \72898 , \72897 );
buf \U$72946 ( \72899 , \72898 );
buf \U$72947 ( \72900 , \11510 );
or \U$72948 ( \72901 , \72899 , \72900 );
buf \U$72949 ( \72902 , \11472 );
buf \U$72950 ( \72903 , \11507 );
nand \U$72951 ( \72904 , \72902 , \72903 );
buf \U$72952 ( \72905 , \72904 );
buf \U$72953 ( \72906 , \72905 );
nand \U$72954 ( \72907 , \72901 , \72906 );
buf \U$72955 ( \72908 , \72907 );
buf \U$72956 ( \72909 , \72908 );
not \U$72957 ( \72910 , \72909 );
buf \U$72958 ( \72911 , \72910 );
buf \U$72959 ( \72912 , \72911 );
buf \U$72960 ( \72913 , \11688 );
or \U$72961 ( \72914 , \72912 , \72913 );
buf \U$72962 ( \72915 , \11565 );
buf \U$72963 ( \72916 , \11685 );
nand \U$72964 ( \72917 , \72915 , \72916 );
buf \U$72965 ( \72918 , \72917 );
buf \U$72966 ( \72919 , \72918 );
nand \U$72967 ( \72920 , \72914 , \72919 );
buf \U$72968 ( \72921 , \72920 );
buf \U$72969 ( \72922 , \72921 );
nor \U$72970 ( \72923 , \72882 , \72922 );
buf \U$72971 ( \72924 , \72923 );
buf \U$72972 ( \72925 , \72924 );
nand \U$72973 ( \72926 , \72842 , \72925 );
buf \U$72974 ( \72927 , \72926 );
buf \U$72975 ( \72928 , \72927 );
buf \U$72976 ( \72929 , \12239 );
and \U$72977 ( \72930 , \72928 , \72929 );
buf \U$72978 ( \72931 , \12082 );
buf \U$72979 ( \72932 , \12088 );
nand \U$72980 ( \72933 , \72931 , \72932 );
buf \U$72981 ( \72934 , \72933 );
buf \U$72982 ( \72935 , \72934 );
buf \U$72983 ( \72936 , \12148 );
or \U$72984 ( \72937 , \72935 , \72936 );
buf \U$72985 ( \72938 , \12136 );
buf \U$72986 ( \72939 , \12145 );
nand \U$72987 ( \72940 , \72938 , \72939 );
buf \U$72988 ( \72941 , \72940 );
buf \U$72989 ( \72942 , \72941 );
nand \U$72990 ( \72943 , \72937 , \72942 );
buf \U$72991 ( \72944 , \72943 );
buf \U$72992 ( \72945 , \72944 );
buf \U$72993 ( \72946 , \12177 );
and \U$72994 ( \72947 , \72945 , \72946 );
buf \U$72995 ( \72948 , \12165 );
buf \U$72996 ( \72949 , \12174 );
and \U$72997 ( \72950 , \72948 , \72949 );
buf \U$72998 ( \72951 , \72950 );
buf \U$72999 ( \72952 , \72951 );
nor \U$73000 ( \72953 , \72947 , \72952 );
buf \U$73001 ( \72954 , \72953 );
buf \U$73002 ( \72955 , \72954 );
buf \U$73003 ( \72956 , \12197 );
or \U$73004 ( \72957 , \72955 , \72956 );
buf \U$73005 ( \72958 , \12189 );
buf \U$73006 ( \72959 , \12194 );
nand \U$73007 ( \72960 , \72958 , \72959 );
buf \U$73008 ( \72961 , \72960 );
buf \U$73009 ( \72962 , \72961 );
nand \U$73010 ( \72963 , \72957 , \72962 );
buf \U$73011 ( \72964 , \72963 );
buf \U$73012 ( \72965 , \72964 );
buf \U$73013 ( \72966 , \11995 );
and \U$73014 ( \72967 , \72965 , \72966 );
buf \U$73015 ( \72968 , \11889 );
buf \U$73016 ( \72969 , \11931 );
nand \U$73017 ( \72970 , \72968 , \72969 );
buf \U$73018 ( \72971 , \72970 );
buf \U$73019 ( \72972 , \72971 );
buf \U$73020 ( \72973 , \11992 );
or \U$73021 ( \72974 , \72972 , \72973 );
buf \U$73022 ( \72975 , \11943 );
buf \U$73023 ( \72976 , \11989 );
nand \U$73024 ( \72977 , \72975 , \72976 );
buf \U$73025 ( \72978 , \72977 );
buf \U$73026 ( \72979 , \72978 );
nand \U$73027 ( \72980 , \72974 , \72979 );
buf \U$73028 ( \72981 , \72980 );
buf \U$73029 ( \72982 , \72981 );
nor \U$73030 ( \72983 , \72967 , \72982 );
buf \U$73031 ( \72984 , \72983 );
buf \U$73032 ( \72985 , \72984 );
buf \U$73033 ( \72986 , \12236 );
or \U$73034 ( \72987 , \72985 , \72986 );
buf \U$73035 ( \72988 , \12207 );
buf \U$73036 ( \72989 , \12233 );
nand \U$73037 ( \72990 , \72988 , \72989 );
buf \U$73038 ( \72991 , \72990 );
buf \U$73039 ( \72992 , \72991 );
nand \U$73040 ( \72993 , \72987 , \72992 );
buf \U$73041 ( \72994 , \72993 );
buf \U$73042 ( \72995 , \72994 );
nor \U$73043 ( \72996 , \72930 , \72995 );
buf \U$73044 ( \72997 , \72996 );
buf \U$73045 ( \72998 , \72997 );
nand \U$73046 ( \72999 , \72670 , \72998 );
buf \U$73047 ( \73000 , \72999 );
buf \U$73048 ( \73001 , \73000 );
buf \U$73049 ( \73002 , \12223 );
not \U$73050 ( \73003 , \73002 );
buf \U$73051 ( \73004 , RIc0d7678_1);
buf \U$73052 ( \73005 , RIc0d9478_65);
nand \U$73053 ( \73006 , \73004 , \73005 );
buf \U$73054 ( \73007 , \73006 );
buf \U$73055 ( \73008 , \73007 );
not \U$73056 ( \73009 , \73008 );
or \U$73057 ( \73010 , \1235 , \3781 );
nand \U$73058 ( \73011 , \73010 , RIc0d9478_65);
buf \U$73059 ( \73012 , \73011 );
not \U$73060 ( \73013 , \73012 );
or \U$73061 ( \73014 , \73009 , \73013 );
buf \U$73062 ( \73015 , \73011 );
buf \U$73063 ( \73016 , \73007 );
or \U$73064 ( \73017 , \73015 , \73016 );
nand \U$73065 ( \73018 , \73014 , \73017 );
buf \U$73066 ( \73019 , \73018 );
buf \U$73067 ( \73020 , \73019 );
not \U$73068 ( \73021 , \73020 );
or \U$73069 ( \73022 , \73003 , \73021 );
buf \U$73070 ( \73023 , \73019 );
buf \U$73071 ( \73024 , \12223 );
or \U$73072 ( \73025 , \73023 , \73024 );
nand \U$73073 ( \73026 , \73022 , \73025 );
buf \U$73074 ( \73027 , \73026 );
buf \U$73075 ( \73028 , \73027 );
not \U$73076 ( \73029 , \73028 );
xor \U$73077 ( \73030 , \12219 , \12224 );
and \U$73078 ( \73031 , \73030 , \12231 );
and \U$73079 ( \73032 , \12219 , \12224 );
or \U$73080 ( \73033 , \73031 , \73032 );
buf \U$73081 ( \73034 , \73033 );
buf \U$73082 ( \73035 , \73034 );
not \U$73083 ( \73036 , \73035 );
or \U$73084 ( \73037 , \73029 , \73036 );
buf \U$73085 ( \73038 , \73034 );
buf \U$73086 ( \73039 , \73027 );
or \U$73087 ( \73040 , \73038 , \73039 );
nand \U$73088 ( \73041 , \73037 , \73040 );
buf \U$73089 ( \73042 , \73041 );
buf \U$73090 ( \73043 , \73042 );
not \U$73091 ( \73044 , \73043 );
buf \U$73092 ( \73045 , \73044 );
buf \U$73093 ( \73046 , \73045 );
and \U$73094 ( \73047 , \73001 , \73046 );
not \U$73095 ( \73048 , \73001 );
buf \U$73096 ( \73049 , \73042 );
and \U$73097 ( \73050 , \73048 , \73049 );
nor \U$73098 ( \73051 , \73047 , \73050 );
buf \U$73099 ( \73052 , \73051 );
buf \U$73100 ( \73053 , \73052 );
buf \U$73101 ( \73054 , \12200 );
buf \U$73102 ( \73055 , \11697 );
buf \U$73103 ( \73056 , \11995 );
and \U$73104 ( \73057 , \73054 , \73055 , \73056 );
buf \U$73105 ( \73058 , \73057 );
buf \U$73106 ( \73059 , \73058 );
not \U$73107 ( \73060 , \73059 );
buf \U$73108 ( \73061 , \43525 );
buf \U$73109 ( \73062 , \43737 );
not \U$73110 ( \73063 , \73062 );
buf \U$73111 ( \73064 , \73063 );
buf \U$73112 ( \73065 , \73064 );
and \U$73113 ( \73066 , \73061 , \73065 );
buf \U$73114 ( \73067 , \73066 );
buf \U$73115 ( \73068 , \73067 );
buf \U$73116 ( \73069 , \72663 );
buf \U$73119 ( \73070 , \43691 );
buf \U$73120 ( \73071 , \73070 );
buf \U$73121 ( \73072 , \43516 );
nand \U$73122 ( \73073 , \73071 , \73072 );
buf \U$73123 ( \73074 , \73073 );
buf \U$73124 ( \73075 , \73074 );
nand \U$73125 ( \73076 , \73068 , \73069 , \73075 );
buf \U$73126 ( \73077 , \73076 );
buf \U$73127 ( \73078 , \73077 );
buf \U$73130 ( \73079 , \10111 );
buf \U$73131 ( \73080 , \73079 );
and \U$73132 ( \73081 , \73078 , \73080 );
buf \U$73133 ( \73082 , \73081 );
buf \U$73134 ( \73083 , \73082 );
not \U$73135 ( \73084 , \73083 );
or \U$73136 ( \73085 , \73060 , \73084 );
buf \U$73137 ( \73086 , \72839 );
buf \U$73138 ( \73087 , \73058 );
and \U$73139 ( \73088 , \73086 , \73087 );
buf \U$73140 ( \73089 , \72924 );
not \U$73141 ( \73090 , \73089 );
buf \U$73142 ( \73091 , \73090 );
buf \U$73143 ( \73092 , \73091 );
buf \U$73144 ( \73093 , \12200 );
and \U$73145 ( \73094 , \73092 , \73093 );
buf \U$73146 ( \73095 , \72964 );
nor \U$73147 ( \73096 , \73094 , \73095 );
buf \U$73148 ( \73097 , \73096 );
buf \U$73149 ( \73098 , \73097 );
not \U$73150 ( \73099 , \73098 );
buf \U$73151 ( \73100 , \73099 );
buf \U$73152 ( \73101 , \73100 );
buf \U$73153 ( \73102 , \11995 );
and \U$73154 ( \73103 , \73101 , \73102 );
buf \U$73155 ( \73104 , \72981 );
nor \U$73156 ( \73105 , \73088 , \73103 , \73104 );
buf \U$73157 ( \73106 , \73105 );
buf \U$73158 ( \73107 , \73106 );
nand \U$73159 ( \73108 , \73085 , \73107 );
buf \U$73160 ( \73109 , \73108 );
buf \U$73161 ( \73110 , \73109 );
buf \U$73162 ( \73111 , \12236 );
not \U$73163 ( \73112 , \73111 );
buf \U$73164 ( \73113 , \72991 );
nand \U$73165 ( \73114 , \73112 , \73113 );
buf \U$73166 ( \73115 , \73114 );
buf \U$73167 ( \73116 , \73115 );
not \U$73168 ( \73117 , \73116 );
buf \U$73169 ( \73118 , \73117 );
buf \U$73170 ( \73119 , \73118 );
and \U$73171 ( \73120 , \73110 , \73119 );
not \U$73172 ( \73121 , \73110 );
buf \U$73173 ( \73122 , \73115 );
and \U$73174 ( \73123 , \73121 , \73122 );
nor \U$73175 ( \73124 , \73120 , \73123 );
buf \U$73176 ( \73125 , \73124 );
buf \U$73177 ( \73126 , \73125 );
buf \U$73178 ( \73127 , \11694 );
buf \U$73179 ( \73128 , \12201 );
buf \U$73180 ( \73129 , \11934 );
nor \U$73181 ( \73130 , \73127 , \73128 , \73129 );
buf \U$73182 ( \73131 , \73130 );
buf \U$73183 ( \73132 , \73131 );
not \U$73184 ( \73133 , \73132 );
buf \U$73185 ( \73134 , \73082 );
not \U$73186 ( \73135 , \73134 );
or \U$73187 ( \73136 , \73133 , \73135 );
buf \U$73190 ( \73137 , \72839 );
buf \U$73191 ( \73138 , \73137 );
buf \U$73192 ( \73139 , \73131 );
and \U$73193 ( \73140 , \73138 , \73139 );
buf \U$73194 ( \73141 , \11934 );
buf \U$73195 ( \73142 , \73097 );
or \U$73196 ( \73143 , \73141 , \73142 );
buf \U$73197 ( \73144 , \72971 );
nand \U$73198 ( \73145 , \73143 , \73144 );
buf \U$73199 ( \73146 , \73145 );
buf \U$73200 ( \73147 , \73146 );
nor \U$73201 ( \73148 , \73140 , \73147 );
buf \U$73202 ( \73149 , \73148 );
buf \U$73203 ( \73150 , \73149 );
nand \U$73204 ( \73151 , \73136 , \73150 );
buf \U$73205 ( \73152 , \73151 );
buf \U$73206 ( \73153 , \73152 );
buf \U$73207 ( \73154 , \11992 );
not \U$73208 ( \73155 , \73154 );
buf \U$73209 ( \73156 , \72978 );
nand \U$73210 ( \73157 , \73155 , \73156 );
buf \U$73211 ( \73158 , \73157 );
buf \U$73212 ( \73159 , \73158 );
not \U$73213 ( \73160 , \73159 );
buf \U$73214 ( \73161 , \73160 );
buf \U$73215 ( \73162 , \73161 );
and \U$73216 ( \73163 , \73153 , \73162 );
not \U$73217 ( \73164 , \73153 );
buf \U$73218 ( \73165 , \73158 );
and \U$73219 ( \73166 , \73164 , \73165 );
nor \U$73220 ( \73167 , \73163 , \73166 );
buf \U$73221 ( \73168 , \73167 );
buf \U$73222 ( \73169 , \73168 );
buf \U$73223 ( \73170 , \12200 );
buf \U$73224 ( \73171 , \11700 );
and \U$73225 ( \73172 , \73170 , \73171 );
buf \U$73226 ( \73173 , \73172 );
buf \U$73227 ( \73174 , \73173 );
not \U$73228 ( \73175 , \73174 );
buf \U$73229 ( \73176 , \72667 );
not \U$73230 ( \73177 , \73176 );
or \U$73231 ( \73178 , \73175 , \73177 );
buf \U$73232 ( \73179 , \72927 );
buf \U$73233 ( \73180 , \12200 );
and \U$73234 ( \73181 , \73179 , \73180 );
buf \U$73235 ( \73182 , \72964 );
nor \U$73236 ( \73183 , \73181 , \73182 );
buf \U$73237 ( \73184 , \73183 );
buf \U$73238 ( \73185 , \73184 );
nand \U$73239 ( \73186 , \73178 , \73185 );
buf \U$73240 ( \73187 , \73186 );
buf \U$73241 ( \73188 , \73187 );
buf \U$73242 ( \73189 , \11934 );
not \U$73243 ( \73190 , \73189 );
buf \U$73244 ( \73191 , \72971 );
nand \U$73245 ( \73192 , \73190 , \73191 );
buf \U$73246 ( \73193 , \73192 );
buf \U$73247 ( \73194 , \73193 );
not \U$73248 ( \73195 , \73194 );
buf \U$73249 ( \73196 , \73195 );
buf \U$73250 ( \73197 , \73196 );
and \U$73251 ( \73198 , \73188 , \73197 );
not \U$73252 ( \73199 , \73188 );
buf \U$73253 ( \73200 , \73193 );
and \U$73254 ( \73201 , \73199 , \73200 );
nor \U$73255 ( \73202 , \73198 , \73201 );
buf \U$73256 ( \73203 , \73202 );
buf \U$73257 ( \73204 , \73203 );
buf \U$73258 ( \73205 , \11694 );
buf \U$73259 ( \73206 , \12180 );
nor \U$73260 ( \73207 , \73205 , \73206 );
buf \U$73261 ( \73208 , \73207 );
buf \U$73262 ( \73209 , \73208 );
not \U$73263 ( \73210 , \73209 );
buf \U$73264 ( \73211 , \73082 );
not \U$73265 ( \73212 , \73211 );
or \U$73266 ( \73213 , \73210 , \73212 );
buf \U$73267 ( \73214 , \73137 );
buf \U$73268 ( \73215 , \73208 );
and \U$73269 ( \73216 , \73214 , \73215 );
buf \U$73270 ( \73217 , \72924 );
buf \U$73271 ( \73218 , \12180 );
or \U$73272 ( \73219 , \73217 , \73218 );
buf \U$73273 ( \73220 , \72954 );
nand \U$73274 ( \73221 , \73219 , \73220 );
buf \U$73275 ( \73222 , \73221 );
buf \U$73276 ( \73223 , \73222 );
nor \U$73277 ( \73224 , \73216 , \73223 );
buf \U$73278 ( \73225 , \73224 );
buf \U$73279 ( \73226 , \73225 );
nand \U$73280 ( \73227 , \73213 , \73226 );
buf \U$73281 ( \73228 , \73227 );
buf \U$73282 ( \73229 , \73228 );
buf \U$73283 ( \73230 , \12197 );
not \U$73284 ( \73231 , \73230 );
buf \U$73285 ( \73232 , \72961 );
nand \U$73286 ( \73233 , \73231 , \73232 );
buf \U$73287 ( \73234 , \73233 );
buf \U$73288 ( \73235 , \73234 );
not \U$73289 ( \73236 , \73235 );
buf \U$73290 ( \73237 , \73236 );
buf \U$73291 ( \73238 , \73237 );
and \U$73292 ( \73239 , \73229 , \73238 );
not \U$73293 ( \73240 , \73229 );
buf \U$73294 ( \73241 , \73234 );
and \U$73295 ( \73242 , \73240 , \73241 );
nor \U$73296 ( \73243 , \73239 , \73242 );
buf \U$73297 ( \73244 , \73243 );
buf \U$73298 ( \73245 , \73244 );
buf \U$73299 ( \73246 , \12151 );
buf \U$73300 ( \73247 , \11700 );
and \U$73301 ( \73248 , \73246 , \73247 );
buf \U$73302 ( \73249 , \73248 );
buf \U$73303 ( \73250 , \73249 );
not \U$73304 ( \73251 , \73250 );
buf \U$73305 ( \73252 , \72667 );
not \U$73306 ( \73253 , \73252 );
or \U$73307 ( \73254 , \73251 , \73253 );
buf \U$73308 ( \73255 , \72927 );
buf \U$73309 ( \73256 , \12151 );
and \U$73310 ( \73257 , \73255 , \73256 );
buf \U$73311 ( \73258 , \72944 );
nor \U$73312 ( \73259 , \73257 , \73258 );
buf \U$73313 ( \73260 , \73259 );
buf \U$73314 ( \73261 , \73260 );
nand \U$73315 ( \73262 , \73254 , \73261 );
buf \U$73316 ( \73263 , \73262 );
buf \U$73317 ( \73264 , \73263 );
buf \U$73318 ( \73265 , \72951 );
not \U$73319 ( \73266 , \73265 );
buf \U$73320 ( \73267 , \12177 );
nand \U$73321 ( \73268 , \73266 , \73267 );
buf \U$73322 ( \73269 , \73268 );
buf \U$73323 ( \73270 , \73269 );
not \U$73324 ( \73271 , \73270 );
buf \U$73325 ( \73272 , \73271 );
buf \U$73326 ( \73273 , \73272 );
and \U$73327 ( \73274 , \73264 , \73273 );
not \U$73328 ( \73275 , \73264 );
buf \U$73329 ( \73276 , \73269 );
and \U$73330 ( \73277 , \73275 , \73276 );
nor \U$73331 ( \73278 , \73274 , \73277 );
buf \U$73332 ( \73279 , \73278 );
buf \U$73333 ( \73280 , \73279 );
buf \U$73334 ( \73281 , \11700 );
buf \U$73335 ( \73282 , \12091 );
and \U$73336 ( \73283 , \73281 , \73282 );
buf \U$73337 ( \73284 , \73283 );
buf \U$73338 ( \73285 , \73284 );
not \U$73339 ( \73286 , \73285 );
buf \U$73340 ( \73287 , \72667 );
not \U$73341 ( \73288 , \73287 );
or \U$73342 ( \73289 , \73286 , \73288 );
buf \U$73343 ( \73290 , \72927 );
buf \U$73344 ( \73291 , \12091 );
and \U$73345 ( \73292 , \73290 , \73291 );
buf \U$73346 ( \73293 , \72934 );
not \U$73347 ( \73294 , \73293 );
buf \U$73348 ( \73295 , \73294 );
buf \U$73349 ( \73296 , \73295 );
nor \U$73350 ( \73297 , \73292 , \73296 );
buf \U$73351 ( \73298 , \73297 );
buf \U$73352 ( \73299 , \73298 );
nand \U$73353 ( \73300 , \73289 , \73299 );
buf \U$73354 ( \73301 , \73300 );
buf \U$73355 ( \73302 , \73301 );
buf \U$73356 ( \73303 , \12148 );
not \U$73357 ( \73304 , \73303 );
buf \U$73358 ( \73305 , \72941 );
nand \U$73359 ( \73306 , \73304 , \73305 );
buf \U$73360 ( \73307 , \73306 );
buf \U$73361 ( \73308 , \73307 );
not \U$73362 ( \73309 , \73308 );
buf \U$73363 ( \73310 , \73309 );
buf \U$73364 ( \73311 , \73310 );
and \U$73365 ( \73312 , \73302 , \73311 );
not \U$73366 ( \73313 , \73302 );
buf \U$73367 ( \73314 , \73307 );
and \U$73368 ( \73315 , \73313 , \73314 );
nor \U$73369 ( \73316 , \73312 , \73315 );
buf \U$73370 ( \73317 , \73316 );
buf \U$73371 ( \73318 , \73317 );
buf \U$73372 ( \73319 , \11700 );
not \U$73373 ( \73320 , \73319 );
buf \U$73374 ( \73321 , \72667 );
not \U$73375 ( \73322 , \73321 );
or \U$73376 ( \73323 , \73320 , \73322 );
buf \U$73377 ( \73324 , \72927 );
not \U$73378 ( \73325 , \73324 );
buf \U$73379 ( \73326 , \73325 );
buf \U$73380 ( \73327 , \73326 );
nand \U$73381 ( \73328 , \73323 , \73327 );
buf \U$73382 ( \73329 , \73328 );
buf \U$73383 ( \73330 , \73329 );
buf \U$73384 ( \73331 , \72934 );
buf \U$73385 ( \73332 , \12091 );
nand \U$73386 ( \73333 , \73331 , \73332 );
buf \U$73387 ( \73334 , \73333 );
buf \U$73388 ( \73335 , \73334 );
not \U$73389 ( \73336 , \73335 );
buf \U$73390 ( \73337 , \73336 );
buf \U$73391 ( \73338 , \73337 );
and \U$73392 ( \73339 , \73330 , \73338 );
not \U$73393 ( \73340 , \73330 );
buf \U$73394 ( \73341 , \73334 );
and \U$73395 ( \73342 , \73340 , \73341 );
nor \U$73396 ( \73343 , \73339 , \73342 );
buf \U$73397 ( \73344 , \73343 );
buf \U$73398 ( \73345 , \73344 );
buf \U$73399 ( \73346 , \11057 );
buf \U$73400 ( \73347 , \11559 );
not \U$73401 ( \73348 , \73347 );
buf \U$73402 ( \73349 , \73348 );
buf \U$73403 ( \73350 , \73349 );
and \U$73404 ( \73351 , \73346 , \73350 );
buf \U$73405 ( \73352 , \73351 );
buf \U$73406 ( \73353 , \73352 );
not \U$73407 ( \73354 , \73353 );
buf \U$73408 ( \73355 , \73082 );
not \U$73409 ( \73356 , \73355 );
or \U$73410 ( \73357 , \73354 , \73356 );
buf \U$73411 ( \73358 , \72839 );
buf \U$73412 ( \73359 , \73352 );
and \U$73413 ( \73360 , \73358 , \73359 );
buf \U$73414 ( \73361 , \72879 );
buf \U$73415 ( \73362 , \73349 );
and \U$73416 ( \73363 , \73361 , \73362 );
buf \U$73417 ( \73364 , \72908 );
nor \U$73418 ( \73365 , \73360 , \73363 , \73364 );
buf \U$73419 ( \73366 , \73365 );
buf \U$73420 ( \73367 , \73366 );
nand \U$73421 ( \73368 , \73357 , \73367 );
buf \U$73422 ( \73369 , \73368 );
buf \U$73423 ( \73370 , \73369 );
buf \U$73424 ( \73371 , \11688 );
not \U$73425 ( \73372 , \73371 );
buf \U$73426 ( \73373 , \72918 );
nand \U$73427 ( \73374 , \73372 , \73373 );
buf \U$73428 ( \73375 , \73374 );
buf \U$73429 ( \73376 , \73375 );
not \U$73430 ( \73377 , \73376 );
buf \U$73431 ( \73378 , \73377 );
buf \U$73432 ( \73379 , \73378 );
and \U$73433 ( \73380 , \73370 , \73379 );
not \U$73434 ( \73381 , \73370 );
buf \U$73435 ( \73382 , \73375 );
and \U$73436 ( \73383 , \73381 , \73382 );
nor \U$73437 ( \73384 , \73380 , \73383 );
buf \U$73438 ( \73385 , \73384 );
buf \U$73439 ( \73386 , \73385 );
buf \U$73440 ( \73387 , \11556 );
not \U$73441 ( \73388 , \73387 );
buf \U$73442 ( \73389 , \43740 );
not \U$73443 ( \73390 , \73389 );
buf \U$73444 ( \73391 , \73390 );
buf \U$73445 ( \73392 , \73391 );
not \U$73446 ( \73393 , \73392 );
buf \U$73447 ( \73394 , \10111 );
buf \U$73448 ( \73395 , \11057 );
and \U$73449 ( \73396 , \73394 , \73395 );
buf \U$73450 ( \73397 , \73396 );
buf \U$73451 ( \73398 , \73397 );
not \U$73452 ( \73399 , \73398 );
or \U$73453 ( \73400 , \73393 , \73399 );
buf \U$73454 ( \73401 , \11057 );
buf \U$73455 ( \73402 , \72839 );
and \U$73456 ( \73403 , \73401 , \73402 );
buf \U$73457 ( \73404 , \72879 );
nor \U$73458 ( \73405 , \73403 , \73404 );
buf \U$73459 ( \73406 , \73405 );
buf \U$73460 ( \73407 , \73406 );
nand \U$73461 ( \73408 , \73400 , \73407 );
buf \U$73462 ( \73409 , \73408 );
buf \U$73463 ( \73410 , \73409 );
not \U$73464 ( \73411 , \73410 );
buf \U$73465 ( \73412 , \73411 );
buf \U$73466 ( \73413 , \73412 );
buf \U$73467 ( \73414 , \72663 );
not \U$73468 ( \73415 , \73414 );
buf \U$73469 ( \73416 , \43525 );
not \U$73470 ( \73417 , \73416 );
or \U$73471 ( \73418 , \73415 , \73417 );
buf \U$73472 ( \73419 , \73397 );
nand \U$73473 ( \73420 , \73418 , \73419 );
buf \U$73474 ( \73421 , \73420 );
buf \U$73475 ( \73422 , \73421 );
nand \U$73476 ( \73423 , \73413 , \73422 );
buf \U$73477 ( \73424 , \73423 );
buf \U$73478 ( \73425 , \73424 );
not \U$73479 ( \73426 , \73425 );
or \U$73480 ( \73427 , \73388 , \73426 );
buf \U$73481 ( \73428 , \72898 );
nand \U$73482 ( \73429 , \73427 , \73428 );
buf \U$73483 ( \73430 , \73429 );
buf \U$73484 ( \73431 , \73430 );
buf \U$73485 ( \73432 , \11510 );
not \U$73486 ( \73433 , \73432 );
buf \U$73487 ( \73434 , \72905 );
nand \U$73488 ( \73435 , \73433 , \73434 );
buf \U$73489 ( \73436 , \73435 );
buf \U$73490 ( \73437 , \73436 );
not \U$73491 ( \73438 , \73437 );
buf \U$73492 ( \73439 , \73438 );
buf \U$73493 ( \73440 , \73439 );
and \U$73494 ( \73441 , \73431 , \73440 );
not \U$73495 ( \73442 , \73431 );
buf \U$73496 ( \73443 , \73436 );
and \U$73497 ( \73444 , \73442 , \73443 );
nor \U$73498 ( \73445 , \73441 , \73444 );
buf \U$73499 ( \73446 , \73445 );
buf \U$73500 ( \73447 , \73446 );
buf \U$73501 ( \73448 , \11540 );
not \U$73502 ( \73449 , \73448 );
buf \U$73503 ( \73450 , \73449 );
buf \U$73504 ( \73451 , \73450 );
not \U$73505 ( \73452 , \73451 );
buf \U$73506 ( \73453 , \73424 );
not \U$73507 ( \73454 , \73453 );
or \U$73508 ( \73455 , \73452 , \73454 );
buf \U$73509 ( \73456 , \72888 );
nand \U$73510 ( \73457 , \73455 , \73456 );
buf \U$73511 ( \73458 , \73457 );
buf \U$73512 ( \73459 , \73458 );
buf \U$73513 ( \73460 , \72895 );
buf \U$73514 ( \73461 , \11553 );
nor \U$73515 ( \73462 , \73460 , \73461 );
buf \U$73516 ( \73463 , \73462 );
buf \U$73517 ( \73464 , \73463 );
and \U$73518 ( \73465 , \73459 , \73464 );
not \U$73519 ( \73466 , \73459 );
buf \U$73520 ( \73467 , \73463 );
not \U$73521 ( \73468 , \73467 );
buf \U$73522 ( \73469 , \73468 );
buf \U$73523 ( \73470 , \73469 );
and \U$73524 ( \73471 , \73466 , \73470 );
nor \U$73525 ( \73472 , \73465 , \73471 );
buf \U$73526 ( \73473 , \73472 );
buf \U$73527 ( \73474 , \73473 );
buf \U$73528 ( \73475 , \73424 );
buf \U$73529 ( \73476 , \73450 );
buf \U$73530 ( \73477 , \72888 );
nand \U$73531 ( \73478 , \73476 , \73477 );
buf \U$73532 ( \73479 , \73478 );
buf \U$73533 ( \73480 , \73479 );
not \U$73534 ( \73481 , \73480 );
buf \U$73535 ( \73482 , \73481 );
buf \U$73536 ( \73483 , \73482 );
and \U$73537 ( \73484 , \73475 , \73483 );
not \U$73538 ( \73485 , \73475 );
buf \U$73539 ( \73486 , \73479 );
and \U$73540 ( \73487 , \73485 , \73486 );
nor \U$73541 ( \73488 , \73484 , \73487 );
buf \U$73542 ( \73489 , \73488 );
buf \U$73543 ( \73490 , \73489 );
buf \U$73544 ( \73491 , \73079 );
not \U$73545 ( \73492 , \73491 );
buf \U$73546 ( \73493 , \10828 );
nor \U$73547 ( \73494 , \73492 , \73493 );
buf \U$73548 ( \73495 , \73494 );
buf \U$73549 ( \73496 , \73495 );
not \U$73550 ( \73497 , \73496 );
buf \U$73551 ( \73498 , \72667 );
not \U$73552 ( \73499 , \73498 );
or \U$73553 ( \73500 , \73497 , \73499 );
buf \U$73554 ( \73501 , \10825 );
not \U$73555 ( \73502 , \73501 );
buf \U$73556 ( \73503 , \10580 );
not \U$73557 ( \73504 , \73503 );
buf \U$73558 ( \73505 , \72839 );
not \U$73559 ( \73506 , \73505 );
or \U$73560 ( \73507 , \73504 , \73506 );
buf \U$73561 ( \73508 , \72856 );
not \U$73562 ( \73509 , \73508 );
buf \U$73563 ( \73510 , \73509 );
buf \U$73564 ( \73511 , \73510 );
nand \U$73565 ( \73512 , \73507 , \73511 );
buf \U$73566 ( \73513 , \73512 );
buf \U$73567 ( \73514 , \73513 );
not \U$73568 ( \73515 , \73514 );
or \U$73569 ( \73516 , \73502 , \73515 );
buf \U$73570 ( \73517 , \72863 );
nand \U$73571 ( \73518 , \73516 , \73517 );
buf \U$73572 ( \73519 , \73518 );
buf \U$73573 ( \73520 , \73519 );
not \U$73574 ( \73521 , \73520 );
buf \U$73575 ( \73522 , \73521 );
buf \U$73576 ( \73523 , \73522 );
nand \U$73577 ( \73524 , \73500 , \73523 );
buf \U$73578 ( \73525 , \73524 );
buf \U$73579 ( \73526 , \73525 );
buf \U$73580 ( \73527 , \11054 );
not \U$73581 ( \73528 , \73527 );
buf \U$73582 ( \73529 , \72876 );
nand \U$73583 ( \73530 , \73528 , \73529 );
buf \U$73584 ( \73531 , \73530 );
buf \U$73585 ( \73532 , \73531 );
not \U$73586 ( \73533 , \73532 );
buf \U$73587 ( \73534 , \73533 );
buf \U$73588 ( \73535 , \73534 );
and \U$73589 ( \73536 , \73526 , \73535 );
not \U$73590 ( \73537 , \73526 );
buf \U$73591 ( \73538 , \73531 );
and \U$73592 ( \73539 , \73537 , \73538 );
nor \U$73593 ( \73540 , \73536 , \73539 );
buf \U$73594 ( \73541 , \73540 );
buf \U$73595 ( \73542 , \73541 );
not \U$73596 ( \73543 , \10340 );
not \U$73597 ( \73544 , \10346 );
and \U$73598 ( \73545 , \73543 , \73544 );
nor \U$73599 ( \73546 , \73545 , \10577 );
not \U$73600 ( \73547 , \73546 );
not \U$73601 ( \73548 , \73082 );
or \U$73602 ( \73549 , \73547 , \73548 );
buf \U$73603 ( \73550 , \73513 );
not \U$73604 ( \73551 , \73550 );
buf \U$73605 ( \73552 , \73551 );
nand \U$73606 ( \73553 , \73549 , \73552 );
buf \U$73607 ( \73554 , \73553 );
buf \U$73608 ( \73555 , \72863 );
buf \U$73609 ( \73556 , \10825 );
nand \U$73610 ( \73557 , \73555 , \73556 );
buf \U$73611 ( \73558 , \73557 );
buf \U$73612 ( \73559 , \73558 );
not \U$73613 ( \73560 , \73559 );
buf \U$73614 ( \73561 , \73560 );
buf \U$73615 ( \73562 , \73561 );
and \U$73616 ( \73563 , \73554 , \73562 );
not \U$73617 ( \73564 , \73554 );
buf \U$73618 ( \73565 , \73558 );
and \U$73619 ( \73566 , \73564 , \73565 );
nor \U$73620 ( \73567 , \73563 , \73566 );
buf \U$73621 ( \73568 , \73567 );
buf \U$73622 ( \73569 , \73568 );
buf \U$73623 ( \73570 , \73079 );
buf \U$73624 ( \73571 , \10349 );
not \U$73625 ( \73572 , \73571 );
buf \U$73626 ( \73573 , \73572 );
buf \U$73627 ( \73574 , \73573 );
and \U$73628 ( \73575 , \73570 , \73574 );
buf \U$73629 ( \73576 , \73575 );
buf \U$73630 ( \73577 , \73576 );
not \U$73631 ( \73578 , \73577 );
buf \U$73632 ( \73579 , \72667 );
not \U$73633 ( \73580 , \73579 );
or \U$73634 ( \73581 , \73578 , \73580 );
buf \U$73635 ( \73582 , \73137 );
buf \U$73636 ( \73583 , \73573 );
and \U$73637 ( \73584 , \73582 , \73583 );
buf \U$73638 ( \73585 , \72847 );
not \U$73639 ( \73586 , \73585 );
buf \U$73640 ( \73587 , \73586 );
buf \U$73641 ( \73588 , \73587 );
nor \U$73642 ( \73589 , \73584 , \73588 );
buf \U$73643 ( \73590 , \73589 );
buf \U$73644 ( \73591 , \73590 );
nand \U$73645 ( \73592 , \73581 , \73591 );
buf \U$73646 ( \73593 , \73592 );
buf \U$73647 ( \73594 , \73593 );
buf \U$73648 ( \73595 , \10577 );
not \U$73649 ( \73596 , \73595 );
buf \U$73650 ( \73597 , \72853 );
nand \U$73651 ( \73598 , \73596 , \73597 );
buf \U$73652 ( \73599 , \73598 );
buf \U$73653 ( \73600 , \73599 );
not \U$73654 ( \73601 , \73600 );
buf \U$73655 ( \73602 , \73601 );
buf \U$73656 ( \73603 , \73602 );
and \U$73657 ( \73604 , \73594 , \73603 );
not \U$73658 ( \73605 , \73594 );
buf \U$73659 ( \73606 , \73599 );
and \U$73660 ( \73607 , \73605 , \73606 );
nor \U$73661 ( \73608 , \73604 , \73607 );
buf \U$73662 ( \73609 , \73608 );
buf \U$73663 ( \73610 , \73609 );
not \U$73664 ( \73611 , \73082 );
buf \U$73665 ( \73612 , \73611 );
buf \U$73666 ( \73613 , \73137 );
not \U$73667 ( \73614 , \73613 );
buf \U$73668 ( \73615 , \73614 );
buf \U$73669 ( \73616 , \73615 );
nand \U$73670 ( \73617 , \73612 , \73616 );
buf \U$73671 ( \73618 , \73617 );
buf \U$73672 ( \73619 , \73618 );
buf \U$73673 ( \73620 , \73573 );
buf \U$73674 ( \73621 , \72847 );
nand \U$73675 ( \73622 , \73620 , \73621 );
buf \U$73676 ( \73623 , \73622 );
buf \U$73677 ( \73624 , \73623 );
not \U$73678 ( \73625 , \73624 );
buf \U$73679 ( \73626 , \73625 );
buf \U$73680 ( \73627 , \73626 );
and \U$73681 ( \73628 , \73619 , \73627 );
not \U$73682 ( \73629 , \73619 );
buf \U$73683 ( \73630 , \73623 );
and \U$73684 ( \73631 , \73629 , \73630 );
nor \U$73685 ( \73632 , \73628 , \73631 );
buf \U$73686 ( \73633 , \73632 );
buf \U$73687 ( \73634 , \73633 );
buf \U$73688 ( \73635 , \7721 );
buf \U$73689 ( \73636 , \73635 );
not \U$73690 ( \73637 , \73636 );
buf \U$73691 ( \73638 , \9029 );
buf \U$73692 ( \73639 , \9858 );
nand \U$73693 ( \73640 , \73638 , \73639 );
buf \U$73694 ( \73641 , \73640 );
buf \U$73695 ( \73642 , \73641 );
nor \U$73696 ( \73643 , \73637 , \73642 );
buf \U$73697 ( \73644 , \73643 );
buf \U$73698 ( \73645 , \73644 );
not \U$73699 ( \73646 , \73645 );
buf \U$73700 ( \73647 , \72667 );
not \U$73701 ( \73648 , \73647 );
or \U$73702 ( \73649 , \73646 , \73648 );
buf \U$73703 ( \73650 , \72705 );
buf \U$73704 ( \73651 , \73650 );
buf \U$73705 ( \73652 , \9858 );
and \U$73706 ( \73653 , \73651 , \73652 );
buf \U$73707 ( \73654 , \7718 );
not \U$73708 ( \73655 , \73654 );
not \U$73709 ( \73656 , \72736 );
buf \U$73710 ( \73657 , \6100 );
not \U$73711 ( \73658 , \73657 );
buf \U$73712 ( \73659 , \73658 );
not \U$73713 ( \73660 , \73659 );
or \U$73714 ( \73661 , \73656 , \73660 );
nand \U$73715 ( \73662 , \73661 , \72741 );
buf \U$73716 ( \73663 , \73662 );
not \U$73717 ( \73664 , \73663 );
or \U$73718 ( \73665 , \73655 , \73664 );
buf \U$73719 ( \73666 , \72787 );
not \U$73720 ( \73667 , \73666 );
buf \U$73721 ( \73668 , \73667 );
buf \U$73722 ( \73669 , \73668 );
nand \U$73723 ( \73670 , \73665 , \73669 );
buf \U$73724 ( \73671 , \73670 );
buf \U$73725 ( \73672 , \73671 );
not \U$73726 ( \73673 , \73672 );
buf \U$73727 ( \73674 , \73673 );
buf \U$73728 ( \73675 , \73674 );
buf \U$73729 ( \73676 , \73641 );
nor \U$73730 ( \73677 , \73675 , \73676 );
buf \U$73731 ( \73678 , \73677 );
buf \U$73732 ( \73679 , \73678 );
buf \U$73733 ( \73680 , \72826 );
nor \U$73734 ( \73681 , \73653 , \73679 , \73680 );
buf \U$73735 ( \73682 , \73681 );
buf \U$73736 ( \73683 , \73682 );
nand \U$73737 ( \73684 , \73649 , \73683 );
buf \U$73738 ( \73685 , \73684 );
buf \U$73739 ( \73686 , \73685 );
buf \U$73740 ( \73687 , \72833 );
not \U$73741 ( \73688 , \73687 );
buf \U$73742 ( \73689 , \10105 );
nand \U$73743 ( \73690 , \73688 , \73689 );
buf \U$73744 ( \73691 , \73690 );
buf \U$73745 ( \73692 , \73691 );
not \U$73746 ( \73693 , \73692 );
buf \U$73747 ( \73694 , \73693 );
buf \U$73748 ( \73695 , \73694 );
and \U$73749 ( \73696 , \73686 , \73695 );
not \U$73750 ( \73697 , \73686 );
buf \U$73751 ( \73698 , \73691 );
and \U$73752 ( \73699 , \73697 , \73698 );
nor \U$73753 ( \73700 , \73696 , \73699 );
buf \U$73754 ( \73701 , \73700 );
buf \U$73755 ( \73702 , \73701 );
buf \U$73756 ( \73703 , \9602 );
not \U$73757 ( \73704 , \73703 );
buf \U$73758 ( \73705 , \72666 );
buf \U$73759 ( \73706 , \9032 );
and \U$73760 ( \73707 , \73705 , \73706 );
buf \U$73761 ( \73708 , \73707 );
buf \U$73762 ( \73709 , \73708 );
not \U$73763 ( \73710 , \73709 );
or \U$73764 ( \73711 , \73704 , \73710 );
buf \U$73765 ( \73712 , \73650 );
not \U$73766 ( \73713 , \73712 );
buf \U$73767 ( \73714 , \73671 );
buf \U$73768 ( \73715 , \9029 );
nand \U$73769 ( \73716 , \73714 , \73715 );
buf \U$73770 ( \73717 , \73716 );
buf \U$73771 ( \73718 , \73717 );
nand \U$73772 ( \73719 , \73713 , \73718 );
buf \U$73773 ( \73720 , \73719 );
buf \U$73774 ( \73721 , \73720 );
buf \U$73775 ( \73722 , \9602 );
and \U$73776 ( \73723 , \73721 , \73722 );
buf \U$73777 ( \73724 , \72816 );
nor \U$73778 ( \73725 , \73723 , \73724 );
buf \U$73779 ( \73726 , \73725 );
buf \U$73780 ( \73727 , \73726 );
nand \U$73781 ( \73728 , \73711 , \73727 );
buf \U$73782 ( \73729 , \73728 );
buf \U$73783 ( \73730 , \73729 );
buf \U$73784 ( \73731 , \9855 );
buf \U$73785 ( \73732 , \72823 );
nand \U$73786 ( \73733 , \73731 , \73732 );
buf \U$73787 ( \73734 , \73733 );
buf \U$73788 ( \73735 , \73734 );
not \U$73789 ( \73736 , \73735 );
buf \U$73790 ( \73737 , \73736 );
buf \U$73791 ( \73738 , \73737 );
and \U$73792 ( \73739 , \73730 , \73738 );
not \U$73793 ( \73740 , \73730 );
buf \U$73794 ( \73741 , \73734 );
and \U$73795 ( \73742 , \73740 , \73741 );
nor \U$73796 ( \73743 , \73739 , \73742 );
buf \U$73797 ( \73744 , \73743 );
buf \U$73798 ( \73745 , \73744 );
buf \U$73799 ( \73746 , \9599 );
not \U$73800 ( \73747 , \73746 );
buf \U$73801 ( \73748 , \73747 );
buf \U$73802 ( \73749 , \73748 );
not \U$73803 ( \73750 , \73749 );
buf \U$73804 ( \73751 , \73708 );
not \U$73805 ( \73752 , \73751 );
or \U$73806 ( \73753 , \73750 , \73752 );
buf \U$73807 ( \73754 , \73720 );
buf \U$73808 ( \73755 , \73748 );
and \U$73809 ( \73756 , \73754 , \73755 );
buf \U$73810 ( \73757 , \72807 );
not \U$73811 ( \73758 , \73757 );
buf \U$73812 ( \73759 , \73758 );
buf \U$73813 ( \73760 , \73759 );
nor \U$73814 ( \73761 , \73756 , \73760 );
buf \U$73815 ( \73762 , \73761 );
buf \U$73816 ( \73763 , \73762 );
nand \U$73817 ( \73764 , \73753 , \73763 );
buf \U$73818 ( \73765 , \73764 );
buf \U$73819 ( \73766 , \73765 );
buf \U$73820 ( \73767 , \9586 );
not \U$73821 ( \73768 , \73767 );
buf \U$73822 ( \73769 , \72813 );
nand \U$73823 ( \73770 , \73768 , \73769 );
buf \U$73824 ( \73771 , \73770 );
buf \U$73825 ( \73772 , \73771 );
not \U$73826 ( \73773 , \73772 );
buf \U$73827 ( \73774 , \73773 );
buf \U$73828 ( \73775 , \73774 );
and \U$73829 ( \73776 , \73766 , \73775 );
not \U$73830 ( \73777 , \73766 );
buf \U$73831 ( \73778 , \73771 );
and \U$73832 ( \73779 , \73777 , \73778 );
nor \U$73833 ( \73780 , \73776 , \73779 );
buf \U$73834 ( \73781 , \73780 );
buf \U$73835 ( \73782 , \73781 );
buf \U$73836 ( \73783 , \9032 );
not \U$73837 ( \73784 , \73783 );
buf \U$73838 ( \73785 , \72667 );
not \U$73839 ( \73786 , \73785 );
or \U$73840 ( \73787 , \73784 , \73786 );
buf \U$73841 ( \73788 , \73720 );
not \U$73842 ( \73789 , \73788 );
buf \U$73843 ( \73790 , \73789 );
buf \U$73844 ( \73791 , \73790 );
nand \U$73845 ( \73792 , \73787 , \73791 );
buf \U$73846 ( \73793 , \73792 );
buf \U$73847 ( \73794 , \73793 );
buf \U$73848 ( \73795 , \73748 );
buf \U$73849 ( \73796 , \72807 );
nand \U$73850 ( \73797 , \73795 , \73796 );
buf \U$73851 ( \73798 , \73797 );
buf \U$73852 ( \73799 , \73798 );
not \U$73853 ( \73800 , \73799 );
buf \U$73854 ( \73801 , \73800 );
buf \U$73855 ( \73802 , \73801 );
and \U$73856 ( \73803 , \73794 , \73802 );
not \U$73857 ( \73804 , \73794 );
buf \U$73858 ( \73805 , \73798 );
and \U$73859 ( \73806 , \73804 , \73805 );
nor \U$73860 ( \73807 , \73803 , \73806 );
buf \U$73861 ( \73808 , \73807 );
buf \U$73862 ( \73809 , \73808 );
buf \U$73863 ( \73810 , \8744 );
not \U$73864 ( \73811 , \73810 );
buf \U$73865 ( \73812 , \72666 );
buf \U$73866 ( \73813 , \73635 );
buf \U$73867 ( \73814 , \8757 );
and \U$73868 ( \73815 , \73813 , \73814 );
buf \U$73869 ( \73816 , \73815 );
buf \U$73870 ( \73817 , \73816 );
and \U$73871 ( \73818 , \73812 , \73817 );
buf \U$73872 ( \73819 , \73818 );
buf \U$73873 ( \73820 , \73819 );
not \U$73874 ( \73821 , \73820 );
or \U$73875 ( \73822 , \73811 , \73821 );
buf \U$73876 ( \73823 , \73671 );
buf \U$73877 ( \73824 , \8757 );
and \U$73878 ( \73825 , \73823 , \73824 );
buf \U$73879 ( \73826 , \73825 );
buf \U$73880 ( \73827 , \73826 );
buf \U$73881 ( \73828 , \8410 );
and \U$73882 ( \73829 , \73827 , \73828 );
buf \U$73883 ( \73830 , \72686 );
nor \U$73884 ( \73831 , \73829 , \73830 );
buf \U$73885 ( \73832 , \73831 );
not \U$73886 ( \73833 , \73832 );
not \U$73887 ( \73834 , \8741 );
and \U$73888 ( \73835 , \73833 , \73834 );
buf \U$73889 ( \73836 , \72694 );
not \U$73890 ( \73837 , \73836 );
buf \U$73891 ( \73838 , \73837 );
nor \U$73892 ( \73839 , \73835 , \73838 );
buf \U$73893 ( \73840 , \73839 );
nand \U$73894 ( \73841 , \73822 , \73840 );
buf \U$73895 ( \73842 , \73841 );
buf \U$73896 ( \73843 , \73842 );
buf \U$73897 ( \73844 , \9026 );
buf \U$73898 ( \73845 , \72704 );
nand \U$73899 ( \73846 , \73844 , \73845 );
buf \U$73900 ( \73847 , \73846 );
buf \U$73901 ( \73848 , \73847 );
not \U$73902 ( \73849 , \73848 );
buf \U$73903 ( \73850 , \73849 );
buf \U$73904 ( \73851 , \73850 );
and \U$73905 ( \73852 , \73843 , \73851 );
not \U$73906 ( \73853 , \73843 );
buf \U$73907 ( \73854 , \73847 );
and \U$73908 ( \73855 , \73853 , \73854 );
nor \U$73909 ( \73856 , \73852 , \73855 );
buf \U$73910 ( \73857 , \73856 );
buf \U$73911 ( \73858 , \73857 );
buf \U$73912 ( \73859 , \8410 );
not \U$73913 ( \73860 , \73859 );
buf \U$73914 ( \73861 , \73819 );
not \U$73915 ( \73862 , \73861 );
or \U$73916 ( \73863 , \73860 , \73862 );
buf \U$73917 ( \73864 , \73832 );
nand \U$73918 ( \73865 , \73863 , \73864 );
buf \U$73919 ( \73866 , \73865 );
buf \U$73920 ( \73867 , \73866 );
buf \U$73921 ( \73868 , \73838 );
buf \U$73922 ( \73869 , \8741 );
nor \U$73923 ( \73870 , \73868 , \73869 );
buf \U$73924 ( \73871 , \73870 );
buf \U$73925 ( \73872 , \73871 );
and \U$73926 ( \73873 , \73867 , \73872 );
not \U$73927 ( \73874 , \73867 );
buf \U$73928 ( \73875 , \73871 );
not \U$73929 ( \73876 , \73875 );
buf \U$73930 ( \73877 , \73876 );
buf \U$73931 ( \73878 , \73877 );
and \U$73932 ( \73879 , \73874 , \73878 );
nor \U$73933 ( \73880 , \73873 , \73879 );
buf \U$73934 ( \73881 , \73880 );
buf \U$73935 ( \73882 , \73881 );
buf \U$73936 ( \73883 , \73816 );
not \U$73937 ( \73884 , \73883 );
buf \U$73938 ( \73885 , \72667 );
not \U$73939 ( \73886 , \73885 );
or \U$73940 ( \73887 , \73884 , \73886 );
buf \U$73941 ( \73888 , \73826 );
buf \U$73942 ( \73889 , \72678 );
nor \U$73943 ( \73890 , \73888 , \73889 );
buf \U$73944 ( \73891 , \73890 );
buf \U$73945 ( \73892 , \73891 );
nand \U$73946 ( \73893 , \73887 , \73892 );
buf \U$73947 ( \73894 , \73893 );
buf \U$73948 ( \73895 , \73894 );
buf \U$73949 ( \73896 , \72685 );
buf \U$73950 ( \73897 , \8410 );
nand \U$73951 ( \73898 , \73896 , \73897 );
buf \U$73952 ( \73899 , \73898 );
buf \U$73953 ( \73900 , \73899 );
not \U$73954 ( \73901 , \73900 );
buf \U$73955 ( \73902 , \73901 );
buf \U$73956 ( \73903 , \73902 );
and \U$73957 ( \73904 , \73895 , \73903 );
not \U$73958 ( \73905 , \73895 );
buf \U$73959 ( \73906 , \73899 );
and \U$73960 ( \73907 , \73905 , \73906 );
nor \U$73961 ( \73908 , \73904 , \73907 );
buf \U$73962 ( \73909 , \73908 );
buf \U$73963 ( \73910 , \73909 );
buf \U$73964 ( \73911 , \73635 );
not \U$73965 ( \73912 , \73911 );
buf \U$73966 ( \73913 , \72667 );
not \U$73967 ( \73914 , \73913 );
or \U$73968 ( \73915 , \73912 , \73914 );
buf \U$73969 ( \73916 , \73674 );
nand \U$73970 ( \73917 , \73915 , \73916 );
buf \U$73971 ( \73918 , \73917 );
buf \U$73972 ( \73919 , \73918 );
buf \U$73973 ( \73920 , \72678 );
not \U$73974 ( \73921 , \73920 );
buf \U$73975 ( \73922 , \8757 );
nand \U$73976 ( \73923 , \73921 , \73922 );
buf \U$73977 ( \73924 , \73923 );
buf \U$73978 ( \73925 , \73924 );
not \U$73979 ( \73926 , \73925 );
buf \U$73980 ( \73927 , \73926 );
buf \U$73981 ( \73928 , \73927 );
and \U$73982 ( \73929 , \73919 , \73928 );
not \U$73983 ( \73930 , \73919 );
buf \U$73984 ( \73931 , \73924 );
and \U$73985 ( \73932 , \73930 , \73931 );
nor \U$73986 ( \73933 , \73929 , \73932 );
buf \U$73987 ( \73934 , \73933 );
buf \U$73988 ( \73935 , \73934 );
buf \U$73991 ( \73936 , \6103 );
buf \U$73992 ( \73937 , \73936 );
buf \U$73993 ( \73938 , \6950 );
and \U$73994 ( \73939 , \73937 , \73938 );
buf \U$73995 ( \73940 , \73939 );
buf \U$73996 ( \73941 , \73940 );
buf \U$73997 ( \73942 , \7337 );
and \U$73998 ( \73943 , \73941 , \73942 );
buf \U$73999 ( \73944 , \73943 );
buf \U$74000 ( \73945 , \73944 );
not \U$74001 ( \73946 , \73945 );
buf \U$74002 ( \73947 , \72667 );
not \U$74003 ( \73948 , \73947 );
or \U$74004 ( \73949 , \73946 , \73948 );
buf \U$74005 ( \73950 , \73662 );
buf \U$74006 ( \73951 , \6950 );
and \U$74007 ( \73952 , \73950 , \73951 );
buf \U$74008 ( \73953 , \72767 );
nor \U$74009 ( \73954 , \73952 , \73953 );
buf \U$74010 ( \73955 , \73954 );
buf \U$74011 ( \73956 , \73955 );
not \U$74012 ( \73957 , \73956 );
buf \U$74013 ( \73958 , \73957 );
buf \U$74014 ( \73959 , \73958 );
buf \U$74015 ( \73960 , \7337 );
and \U$74016 ( \73961 , \73959 , \73960 );
buf \U$74017 ( \73962 , \72774 );
not \U$74018 ( \73963 , \73962 );
buf \U$74019 ( \73964 , \73963 );
buf \U$74020 ( \73965 , \73964 );
nor \U$74021 ( \73966 , \73961 , \73965 );
buf \U$74022 ( \73967 , \73966 );
buf \U$74023 ( \73968 , \73967 );
nand \U$74024 ( \73969 , \73949 , \73968 );
buf \U$74025 ( \73970 , \73969 );
buf \U$74026 ( \73971 , \73970 );
buf \U$74027 ( \73972 , \72784 );
buf \U$74028 ( \73973 , \7715 );
nand \U$74029 ( \73974 , \73972 , \73973 );
buf \U$74030 ( \73975 , \73974 );
buf \U$74031 ( \73976 , \73975 );
not \U$74032 ( \73977 , \73976 );
buf \U$74033 ( \73978 , \73977 );
buf \U$74034 ( \73979 , \73978 );
and \U$74035 ( \73980 , \73971 , \73979 );
not \U$74036 ( \73981 , \73971 );
buf \U$74037 ( \73982 , \73975 );
and \U$74038 ( \73983 , \73981 , \73982 );
nor \U$74039 ( \73984 , \73980 , \73983 );
buf \U$74040 ( \73985 , \73984 );
buf \U$74041 ( \73986 , \73985 );
buf \U$74042 ( \73987 , \73940 );
not \U$74043 ( \73988 , \73987 );
buf \U$74044 ( \73989 , \72667 );
not \U$74045 ( \73990 , \73989 );
or \U$74046 ( \73991 , \73988 , \73990 );
buf \U$74047 ( \73992 , \73955 );
nand \U$74048 ( \73993 , \73991 , \73992 );
buf \U$74049 ( \73994 , \73993 );
buf \U$74050 ( \73995 , \73994 );
buf \U$74051 ( \73996 , \7337 );
buf \U$74052 ( \73997 , \72774 );
nand \U$74053 ( \73998 , \73996 , \73997 );
buf \U$74054 ( \73999 , \73998 );
buf \U$74055 ( \74000 , \73999 );
not \U$74056 ( \74001 , \74000 );
buf \U$74057 ( \74002 , \74001 );
buf \U$74058 ( \74003 , \74002 );
and \U$74059 ( \74004 , \73995 , \74003 );
not \U$74060 ( \74005 , \73995 );
buf \U$74061 ( \74006 , \73999 );
and \U$74062 ( \74007 , \74005 , \74006 );
nor \U$74063 ( \74008 , \74004 , \74007 );
buf \U$74064 ( \74009 , \74008 );
buf \U$74065 ( \74010 , \74009 );
buf \U$74066 ( \74011 , \73936 );
buf \U$74067 ( \74012 , \6947 );
and \U$74068 ( \74013 , \74011 , \74012 );
buf \U$74069 ( \74014 , \74013 );
buf \U$74070 ( \74015 , \74014 );
not \U$74071 ( \74016 , \74015 );
buf \U$74072 ( \74017 , \72667 );
not \U$74073 ( \74018 , \74017 );
or \U$74074 ( \74019 , \74016 , \74018 );
buf \U$74075 ( \74020 , \73662 );
buf \U$74076 ( \74021 , \6947 );
and \U$74077 ( \74022 , \74020 , \74021 );
buf \U$74078 ( \74023 , \72759 );
nor \U$74079 ( \74024 , \74022 , \74023 );
buf \U$74080 ( \74025 , \74024 );
buf \U$74081 ( \74026 , \74025 );
nand \U$74082 ( \74027 , \74019 , \74026 );
buf \U$74083 ( \74028 , \74027 );
buf \U$74084 ( \74029 , \74028 );
buf \U$74085 ( \74030 , \6931 );
buf \U$74086 ( \74031 , \72766 );
nand \U$74087 ( \74032 , \74030 , \74031 );
buf \U$74088 ( \74033 , \74032 );
buf \U$74089 ( \74034 , \74033 );
not \U$74090 ( \74035 , \74034 );
buf \U$74091 ( \74036 , \74035 );
buf \U$74092 ( \74037 , \74036 );
and \U$74093 ( \74038 , \74029 , \74037 );
not \U$74094 ( \74039 , \74029 );
buf \U$74095 ( \74040 , \74033 );
and \U$74096 ( \74041 , \74039 , \74040 );
nor \U$74097 ( \74042 , \74038 , \74041 );
buf \U$74098 ( \74043 , \74042 );
buf \U$74099 ( \74044 , \74043 );
buf \U$74100 ( \74045 , \73936 );
not \U$74101 ( \74046 , \74045 );
buf \U$74102 ( \74047 , \72667 );
not \U$74103 ( \74048 , \74047 );
or \U$74104 ( \74049 , \74046 , \74048 );
buf \U$74105 ( \74050 , \73662 );
not \U$74106 ( \74051 , \74050 );
buf \U$74107 ( \74052 , \74051 );
buf \U$74108 ( \74053 , \74052 );
nand \U$74109 ( \74054 , \74049 , \74053 );
buf \U$74110 ( \74055 , \74054 );
buf \U$74111 ( \74056 , \74055 );
buf \U$74112 ( \74057 , \72759 );
not \U$74113 ( \74058 , \74057 );
buf \U$74114 ( \74059 , \6947 );
nand \U$74115 ( \74060 , \74058 , \74059 );
buf \U$74116 ( \74061 , \74060 );
buf \U$74117 ( \74062 , \74061 );
not \U$74118 ( \74063 , \74062 );
buf \U$74119 ( \74064 , \74063 );
buf \U$74120 ( \74065 , \74064 );
and \U$74121 ( \74066 , \74056 , \74065 );
not \U$74122 ( \74067 , \74056 );
buf \U$74123 ( \74068 , \74061 );
and \U$74124 ( \74069 , \74067 , \74068 );
nor \U$74125 ( \74070 , \74066 , \74069 );
buf \U$74126 ( \74071 , \74070 );
buf \U$74127 ( \74072 , \74071 );
buf \U$74128 ( \74073 , \5618 );
not \U$74129 ( \74074 , \74073 );
buf \U$74130 ( \74075 , \74074 );
buf \U$74131 ( \74076 , \74075 );
not \U$74132 ( \74077 , \74076 );
buf \U$74133 ( \74078 , \72667 );
not \U$74134 ( \74079 , \74078 );
or \U$74135 ( \74080 , \74077 , \74079 );
buf \U$74136 ( \74081 , \72736 );
not \U$74137 ( \74082 , \74081 );
buf \U$74138 ( \74083 , \74082 );
buf \U$74139 ( \74084 , \74083 );
nand \U$74140 ( \74085 , \74080 , \74084 );
buf \U$74141 ( \74086 , \74085 );
buf \U$74142 ( \74087 , \74086 );
buf \U$74143 ( \74088 , \73659 );
buf \U$74144 ( \74089 , \72741 );
nand \U$74145 ( \74090 , \74088 , \74089 );
buf \U$74146 ( \74091 , \74090 );
buf \U$74147 ( \74092 , \74091 );
not \U$74148 ( \74093 , \74092 );
buf \U$74149 ( \74094 , \74093 );
buf \U$74150 ( \74095 , \74094 );
and \U$74151 ( \74096 , \74087 , \74095 );
not \U$74152 ( \74097 , \74087 );
buf \U$74153 ( \74098 , \74091 );
and \U$74154 ( \74099 , \74097 , \74098 );
nor \U$74155 ( \74100 , \74096 , \74099 );
buf \U$74156 ( \74101 , \74100 );
buf \U$74157 ( \74102 , \74101 );
buf \U$74158 ( \74103 , \5134 );
not \U$74159 ( \74104 , \74103 );
buf \U$74160 ( \74105 , \74104 );
buf \U$74161 ( \74106 , \74105 );
not \U$74162 ( \74107 , \74106 );
buf \U$74163 ( \74108 , \72667 );
not \U$74164 ( \74109 , \74108 );
or \U$74165 ( \74110 , \74107 , \74109 );
buf \U$74166 ( \74111 , \72726 );
not \U$74167 ( \74112 , \74111 );
buf \U$74168 ( \74113 , \74112 );
buf \U$74169 ( \74114 , \74113 );
nand \U$74170 ( \74115 , \74110 , \74114 );
buf \U$74171 ( \74116 , \74115 );
buf \U$74172 ( \74117 , \74116 );
buf \U$74173 ( \74118 , \72733 );
buf \U$74174 ( \74119 , \5615 );
nand \U$74175 ( \74120 , \74118 , \74119 );
buf \U$74176 ( \74121 , \74120 );
buf \U$74177 ( \74122 , \74121 );
not \U$74178 ( \74123 , \74122 );
buf \U$74179 ( \74124 , \74123 );
buf \U$74180 ( \74125 , \74124 );
and \U$74181 ( \74126 , \74117 , \74125 );
not \U$74182 ( \74127 , \74117 );
buf \U$74183 ( \74128 , \74121 );
and \U$74184 ( \74129 , \74127 , \74128 );
nor \U$74185 ( \74130 , \74126 , \74129 );
buf \U$74186 ( \74131 , \74130 );
buf \U$74187 ( \74132 , \74131 );
buf \U$74188 ( \74133 , \4617 );
not \U$74189 ( \74134 , \74133 );
buf \U$74190 ( \74135 , \72667 );
not \U$74191 ( \74136 , \74135 );
or \U$74192 ( \74137 , \74134 , \74136 );
buf \U$74193 ( \74138 , \72717 );
nand \U$74194 ( \74139 , \74137 , \74138 );
buf \U$74195 ( \74140 , \74139 );
buf \U$74196 ( \74141 , \74140 );
buf \U$74197 ( \74142 , \5131 );
buf \U$74198 ( \74143 , \72723 );
nand \U$74199 ( \74144 , \74142 , \74143 );
buf \U$74200 ( \74145 , \74144 );
buf \U$74201 ( \74146 , \74145 );
not \U$74202 ( \74147 , \74146 );
buf \U$74203 ( \74148 , \74147 );
buf \U$74204 ( \74149 , \74148 );
and \U$74205 ( \74150 , \74141 , \74149 );
not \U$74206 ( \74151 , \74141 );
buf \U$74207 ( \74152 , \74145 );
and \U$74208 ( \74153 , \74151 , \74152 );
nor \U$74209 ( \74154 , \74150 , \74153 );
buf \U$74210 ( \74155 , \74154 );
buf \U$74211 ( \74156 , \74155 );
buf \U$74212 ( \74157 , \72717 );
buf \U$74213 ( \74158 , \4617 );
and \U$74214 ( \74159 , \74157 , \74158 );
buf \U$74215 ( \74160 , \74159 );
buf \U$74216 ( \74161 , \74160 );
not \U$74217 ( \74162 , \74161 );
not \U$74218 ( \74163 , \72667 );
buf \U$74219 ( \74164 , \74163 );
not \U$74220 ( \74165 , \74164 );
or \U$74221 ( \74166 , \74162 , \74165 );
buf \U$74222 ( \74167 , \74160 );
buf \U$74223 ( \74168 , \74163 );
or \U$74224 ( \74169 , \74167 , \74168 );
nand \U$74225 ( \74170 , \74166 , \74169 );
buf \U$74226 ( \74171 , \74170 );
buf \U$74227 ( \74172 , \74171 );
buf \U$74228 ( \74173 , \43336 );
buf \U$74229 ( \74174 , \43500 );
and \U$74230 ( \74175 , \74173 , \74174 );
buf \U$74231 ( \74176 , \74175 );
buf \U$74232 ( \74177 , \74176 );
not \U$74233 ( \74178 , \74177 );
not \U$74234 ( \74179 , \35570 );
buf \U$74235 ( \74180 , \43772 );
buf \U$74236 ( \74181 , \72452 );
buf \U$74237 ( \74182 , \63013 );
not \U$74238 ( \74183 , \74182 );
buf \U$74239 ( \74184 , \56473 );
buf \U$74240 ( \74185 , \49374 );
buf \U$74241 ( \74186 , \62972 );
nand \U$74242 ( \74187 , \74184 , \74185 , \74186 );
buf \U$74243 ( \74188 , \74187 );
buf \U$74244 ( \74189 , \74188 );
buf \U$74245 ( \74190 , \56445 );
nand \U$74246 ( \74191 , \74183 , \74189 , \74190 );
buf \U$74247 ( \74192 , \74191 );
buf \U$74248 ( \74193 , \74192 );
nand \U$74249 ( \74194 , \74180 , \74181 , \74193 );
buf \U$74250 ( \74195 , \74194 );
buf \U$74251 ( \74196 , \72657 );
not \U$74252 ( \74197 , \74196 );
buf \U$74253 ( \74198 , \43772 );
nand \U$74254 ( \74199 , \74197 , \74198 );
buf \U$74255 ( \74200 , \74199 );
nand \U$74256 ( \74201 , \74179 , \74195 , \74200 );
buf \U$74257 ( \74202 , \74201 );
buf \U$74258 ( \74203 , \41971 );
buf \U$74259 ( \74204 , \74203 );
and \U$74260 ( \74205 , \74202 , \74204 );
buf \U$74261 ( \74206 , \74205 );
buf \U$74262 ( \74207 , \74206 );
not \U$74263 ( \74208 , \74207 );
or \U$74264 ( \74209 , \74178 , \74208 );
buf \U$74265 ( \74210 , \74176 );
buf \U$74266 ( \74211 , \41637 );
not \U$74267 ( \74212 , \74211 );
buf \U$74268 ( \74213 , \41945 );
not \U$74269 ( \74214 , \74213 );
buf \U$74270 ( \74215 , \41968 );
not \U$74271 ( \74216 , \74215 );
buf \U$74272 ( \74217 , \43608 );
not \U$74273 ( \74218 , \74217 );
or \U$74274 ( \74219 , \74216 , \74218 );
buf \U$74277 ( \74220 , \43624 );
buf \U$74278 ( \74221 , \74220 );
nand \U$74279 ( \74222 , \74219 , \74221 );
buf \U$74280 ( \74223 , \74222 );
buf \U$74281 ( \74224 , \74223 );
not \U$74282 ( \74225 , \74224 );
or \U$74283 ( \74226 , \74214 , \74225 );
buf \U$74284 ( \74227 , \43635 );
nand \U$74285 ( \74228 , \74226 , \74227 );
buf \U$74286 ( \74229 , \74228 );
buf \U$74287 ( \74230 , \74229 );
not \U$74288 ( \74231 , \74230 );
or \U$74289 ( \74232 , \74212 , \74231 );
buf \U$74290 ( \74233 , \43684 );
not \U$74291 ( \74234 , \74233 );
buf \U$74292 ( \74235 , \74234 );
buf \U$74293 ( \74236 , \74235 );
nand \U$74294 ( \74237 , \74232 , \74236 );
buf \U$74295 ( \74238 , \74237 );
buf \U$74296 ( \74239 , \74238 );
and \U$74297 ( \74240 , \74210 , \74239 );
buf \U$74298 ( \74241 , \43500 );
not \U$74299 ( \74242 , \74241 );
buf \U$74300 ( \74243 , \43570 );
not \U$74301 ( \74244 , \74243 );
or \U$74302 ( \74245 , \74242 , \74244 );
buf \U$74303 ( \74246 , \43727 );
not \U$74304 ( \74247 , \74246 );
buf \U$74305 ( \74248 , \74247 );
buf \U$74306 ( \74249 , \74248 );
nand \U$74307 ( \74250 , \74245 , \74249 );
buf \U$74308 ( \74251 , \74250 );
buf \U$74309 ( \74252 , \74251 );
nor \U$74310 ( \74253 , \74240 , \74252 );
buf \U$74311 ( \74254 , \74253 );
buf \U$74312 ( \74255 , \74254 );
nand \U$74313 ( \74256 , \74209 , \74255 );
buf \U$74314 ( \74257 , \74256 );
buf \U$74315 ( \74258 , \74257 );
buf \U$74316 ( \74259 , \43513 );
buf \U$74317 ( \74260 , \43734 );
nand \U$74318 ( \74261 , \74259 , \74260 );
buf \U$74319 ( \74262 , \74261 );
buf \U$74320 ( \74263 , \74262 );
not \U$74321 ( \74264 , \74263 );
buf \U$74322 ( \74265 , \74264 );
buf \U$74323 ( \74266 , \74265 );
and \U$74324 ( \74267 , \74258 , \74266 );
not \U$74325 ( \74268 , \74258 );
buf \U$74326 ( \74269 , \74262 );
and \U$74327 ( \74270 , \74268 , \74269 );
nor \U$74328 ( \74271 , \74267 , \74270 );
buf \U$74329 ( \74272 , \74271 );
buf \U$74330 ( \74273 , \74272 );
buf \U$74331 ( \74274 , \43339 );
not \U$74332 ( \74275 , \74274 );
buf \U$74333 ( \74276 , \74275 );
buf \U$74334 ( \74277 , \74276 );
buf \U$74335 ( \74278 , \43462 );
nor \U$74336 ( \74279 , \74277 , \74278 );
buf \U$74337 ( \74280 , \74279 );
buf \U$74338 ( \74281 , \74280 );
not \U$74339 ( \74282 , \74281 );
buf \U$74340 ( \74283 , \74201 );
buf \U$74342 ( \74284 , \74283 );
buf \U$74343 ( \74285 , \74284 );
not \U$74344 ( \74286 , \74285 );
or \U$74345 ( \74287 , \74282 , \74286 );
buf \U$74346 ( \74288 , \73070 );
buf \U$74347 ( \74289 , \43462 );
not \U$74348 ( \74290 , \74289 );
buf \U$74349 ( \74291 , \74290 );
buf \U$74350 ( \74292 , \74291 );
and \U$74351 ( \74293 , \74288 , \74292 );
buf \U$74352 ( \74294 , \43717 );
nor \U$74353 ( \74295 , \74293 , \74294 );
buf \U$74354 ( \74296 , \74295 );
buf \U$74355 ( \74297 , \74296 );
nand \U$74356 ( \74298 , \74287 , \74297 );
buf \U$74357 ( \74299 , \74298 );
buf \U$74358 ( \74300 , \74299 );
buf \U$74359 ( \74301 , \43699 );
buf \U$74360 ( \74302 , \43724 );
nand \U$74361 ( \74303 , \74301 , \74302 );
buf \U$74362 ( \74304 , \74303 );
buf \U$74363 ( \74305 , \74304 );
not \U$74364 ( \74306 , \74305 );
buf \U$74365 ( \74307 , \74306 );
buf \U$74366 ( \74308 , \74307 );
and \U$74367 ( \74309 , \74300 , \74308 );
not \U$74368 ( \74310 , \74300 );
buf \U$74369 ( \74311 , \74304 );
and \U$74370 ( \74312 , \74310 , \74311 );
nor \U$74371 ( \74313 , \74309 , \74312 );
buf \U$74372 ( \74314 , \74313 );
buf \U$74373 ( \74315 , \74314 );
buf \U$74374 ( \74316 , \74276 );
buf \U$74375 ( \74317 , \43417 );
not \U$74376 ( \74318 , \74317 );
buf \U$74377 ( \74319 , \74318 );
nor \U$74378 ( \74320 , \74316 , \74319 );
buf \U$74379 ( \74321 , \74320 );
buf \U$74380 ( \74322 , \74321 );
not \U$74381 ( \74323 , \74322 );
buf \U$74382 ( \74324 , \74284 );
not \U$74383 ( \74325 , \74324 );
or \U$74384 ( \74326 , \74323 , \74325 );
buf \U$74385 ( \74327 , \73070 );
buf \U$74386 ( \74328 , \74317 );
and \U$74387 ( \74329 , \74327 , \74328 );
buf \U$74388 ( \74330 , \43707 );
buf \U$74389 ( \74331 , \74330 );
nor \U$74390 ( \74332 , \74329 , \74331 );
buf \U$74391 ( \74333 , \74332 );
buf \U$74392 ( \74334 , \74333 );
nand \U$74393 ( \74335 , \74326 , \74334 );
buf \U$74394 ( \74336 , \74335 );
buf \U$74395 ( \74337 , \74336 );
buf \U$74396 ( \74338 , \43459 );
buf \U$74397 ( \74339 , \43714 );
nand \U$74398 ( \74340 , \74338 , \74339 );
buf \U$74399 ( \74341 , \74340 );
buf \U$74400 ( \74342 , \74341 );
not \U$74401 ( \74343 , \74342 );
buf \U$74402 ( \74344 , \74343 );
buf \U$74403 ( \74345 , \74344 );
and \U$74404 ( \74346 , \74337 , \74345 );
not \U$74405 ( \74347 , \74337 );
buf \U$74406 ( \74348 , \74341 );
and \U$74407 ( \74349 , \74347 , \74348 );
nor \U$74408 ( \74350 , \74346 , \74349 );
buf \U$74409 ( \74351 , \74350 );
buf \U$74410 ( \74352 , \74351 );
buf \U$74411 ( \74353 , \43339 );
not \U$74412 ( \74354 , \74353 );
buf \U$74413 ( \74355 , \74284 );
not \U$74414 ( \74356 , \74355 );
or \U$74415 ( \74357 , \74354 , \74356 );
buf \U$74416 ( \74358 , \73070 );
not \U$74417 ( \74359 , \74358 );
buf \U$74418 ( \74360 , \74359 );
buf \U$74419 ( \74361 , \74360 );
nand \U$74420 ( \74362 , \74357 , \74361 );
buf \U$74421 ( \74363 , \74362 );
buf \U$74422 ( \74364 , \74363 );
buf \U$74423 ( \74365 , \74330 );
buf \U$74424 ( \74366 , \74318 );
nor \U$74425 ( \74367 , \74365 , \74366 );
buf \U$74426 ( \74368 , \74367 );
buf \U$74427 ( \74369 , \74368 );
and \U$74428 ( \74370 , \74364 , \74369 );
not \U$74429 ( \74371 , \74364 );
buf \U$74430 ( \74372 , \74368 );
not \U$74431 ( \74373 , \74372 );
buf \U$74432 ( \74374 , \74373 );
buf \U$74433 ( \74375 , \74374 );
and \U$74434 ( \74376 , \74371 , \74375 );
nor \U$74435 ( \74377 , \74370 , \74376 );
buf \U$74436 ( \74378 , \74377 );
buf \U$74437 ( \74379 , \74378 );
buf \U$74438 ( \74380 , \74203 );
buf \U$74439 ( \74381 , \42892 );
buf \U$74440 ( \74382 , \43139 );
and \U$74441 ( \74383 , \74380 , \74381 , \74382 );
buf \U$74442 ( \74384 , \74383 );
buf \U$74443 ( \74385 , \74384 );
not \U$74444 ( \74386 , \74385 );
buf \U$74445 ( \74387 , \74284 );
not \U$74446 ( \74388 , \74387 );
or \U$74447 ( \74389 , \74386 , \74388 );
buf \U$74448 ( \74390 , \43139 );
not \U$74449 ( \74391 , \74390 );
buf \U$74450 ( \74392 , \42892 );
not \U$74451 ( \74393 , \74392 );
buf \U$74452 ( \74394 , \74238 );
not \U$74453 ( \74395 , \74394 );
or \U$74454 ( \74396 , \74393 , \74395 );
buf \U$74455 ( \74397 , \43546 );
not \U$74456 ( \74398 , \74397 );
buf \U$74457 ( \74399 , \74398 );
buf \U$74458 ( \74400 , \74399 );
nand \U$74459 ( \74401 , \74396 , \74400 );
buf \U$74460 ( \74402 , \74401 );
buf \U$74461 ( \74403 , \74402 );
not \U$74462 ( \74404 , \74403 );
or \U$74463 ( \74405 , \74391 , \74404 );
buf \U$74464 ( \74406 , \43553 );
nand \U$74465 ( \74407 , \74405 , \74406 );
buf \U$74466 ( \74408 , \74407 );
buf \U$74467 ( \74409 , \74408 );
not \U$74468 ( \74410 , \74409 );
buf \U$74469 ( \74411 , \74410 );
buf \U$74470 ( \74412 , \74411 );
nand \U$74471 ( \74413 , \74389 , \74412 );
buf \U$74472 ( \74414 , \74413 );
buf \U$74473 ( \74415 , \74414 );
buf \U$74474 ( \74416 , \43567 );
buf \U$74475 ( \74417 , \43558 );
nand \U$74476 ( \74418 , \74416 , \74417 );
buf \U$74477 ( \74419 , \74418 );
buf \U$74478 ( \74420 , \74419 );
not \U$74479 ( \74421 , \74420 );
buf \U$74480 ( \74422 , \74421 );
buf \U$74481 ( \74423 , \74422 );
and \U$74482 ( \74424 , \74415 , \74423 );
not \U$74483 ( \74425 , \74415 );
buf \U$74484 ( \74426 , \74419 );
and \U$74485 ( \74427 , \74425 , \74426 );
nor \U$74486 ( \74428 , \74424 , \74427 );
buf \U$74487 ( \74429 , \74428 );
buf \U$74488 ( \74430 , \74429 );
buf \U$74489 ( \74431 , \42892 );
not \U$74490 ( \74432 , \74431 );
buf \U$74491 ( \74433 , \74206 );
not \U$74492 ( \74434 , \74433 );
or \U$74493 ( \74435 , \74432 , \74434 );
buf \U$74494 ( \74436 , \74402 );
not \U$74495 ( \74437 , \74436 );
buf \U$74496 ( \74438 , \74437 );
buf \U$74497 ( \74439 , \74438 );
nand \U$74498 ( \74440 , \74435 , \74439 );
buf \U$74499 ( \74441 , \74440 );
buf \U$74500 ( \74442 , \74441 );
buf \U$74501 ( \74443 , \43139 );
buf \U$74502 ( \74444 , \43553 );
nand \U$74503 ( \74445 , \74443 , \74444 );
buf \U$74504 ( \74446 , \74445 );
buf \U$74505 ( \74447 , \74446 );
not \U$74506 ( \74448 , \74447 );
buf \U$74507 ( \74449 , \74448 );
buf \U$74508 ( \74450 , \74449 );
and \U$74509 ( \74451 , \74442 , \74450 );
not \U$74510 ( \74452 , \74442 );
buf \U$74511 ( \74453 , \74446 );
and \U$74512 ( \74454 , \74452 , \74453 );
nor \U$74513 ( \74455 , \74451 , \74454 );
buf \U$74514 ( \74456 , \74455 );
buf \U$74515 ( \74457 , \74456 );
buf \U$74516 ( \74458 , \42525 );
not \U$74517 ( \74459 , \74458 );
buf \U$74518 ( \74460 , \74206 );
not \U$74519 ( \74461 , \74460 );
or \U$74520 ( \74462 , \74459 , \74461 );
buf \U$74521 ( \74463 , \42525 );
buf \U$74522 ( \74464 , \74238 );
and \U$74523 ( \74465 , \74463 , \74464 );
buf \U$74524 ( \74466 , \43536 );
not \U$74525 ( \74467 , \74466 );
buf \U$74526 ( \74468 , \74467 );
buf \U$74527 ( \74469 , \74468 );
nor \U$74528 ( \74470 , \74465 , \74469 );
buf \U$74529 ( \74471 , \74470 );
buf \U$74530 ( \74472 , \74471 );
nand \U$74531 ( \74473 , \74462 , \74472 );
buf \U$74532 ( \74474 , \74473 );
buf \U$74533 ( \74475 , \74474 );
buf \U$74534 ( \74476 , \43531 );
not \U$74535 ( \74477 , \74476 );
buf \U$74536 ( \74478 , \43543 );
nand \U$74537 ( \74479 , \74477 , \74478 );
buf \U$74538 ( \74480 , \74479 );
buf \U$74539 ( \74481 , \74480 );
not \U$74540 ( \74482 , \74481 );
buf \U$74541 ( \74483 , \74482 );
buf \U$74542 ( \74484 , \74483 );
and \U$74543 ( \74485 , \74475 , \74484 );
not \U$74544 ( \74486 , \74475 );
buf \U$74545 ( \74487 , \74480 );
and \U$74546 ( \74488 , \74486 , \74487 );
nor \U$74547 ( \74489 , \74485 , \74488 );
buf \U$74548 ( \74490 , \74489 );
buf \U$74549 ( \74491 , \74490 );
buf \U$74550 ( \74492 , \74203 );
not \U$74551 ( \74493 , \74492 );
buf \U$74552 ( \74494 , \74284 );
not \U$74553 ( \74495 , \74494 );
or \U$74554 ( \74496 , \74493 , \74495 );
buf \U$74555 ( \74497 , \74238 );
not \U$74556 ( \74498 , \74497 );
buf \U$74557 ( \74499 , \74498 );
buf \U$74558 ( \74500 , \74499 );
nand \U$74559 ( \74501 , \74496 , \74500 );
buf \U$74560 ( \74502 , \74501 );
buf \U$74561 ( \74503 , \74502 );
buf \U$74562 ( \74504 , \43536 );
buf \U$74563 ( \74505 , \42525 );
nand \U$74564 ( \74506 , \74504 , \74505 );
buf \U$74565 ( \74507 , \74506 );
buf \U$74566 ( \74508 , \74507 );
not \U$74567 ( \74509 , \74508 );
buf \U$74568 ( \74510 , \74509 );
buf \U$74569 ( \74511 , \74510 );
and \U$74570 ( \74512 , \74503 , \74511 );
not \U$74571 ( \74513 , \74503 );
buf \U$74572 ( \74514 , \74507 );
and \U$74573 ( \74515 , \74513 , \74514 );
nor \U$74574 ( \74516 , \74512 , \74515 );
buf \U$74575 ( \74517 , \74516 );
buf \U$74576 ( \74518 , \74517 );
buf \U$74579 ( \74519 , \41631 );
buf \U$74580 ( \74520 , \74519 );
not \U$74581 ( \74521 , \74520 );
buf \U$74582 ( \74522 , \41895 );
buf \U$74583 ( \74523 , \41968 );
and \U$74584 ( \74524 , \74522 , \74523 );
buf \U$74585 ( \74525 , \74524 );
buf \U$74586 ( \74526 , \74525 );
buf \U$74587 ( \74527 , \41945 );
and \U$74588 ( \74528 , \74526 , \74527 );
buf \U$74589 ( \74529 , \74528 );
buf \U$74590 ( \74530 , \74529 );
buf \U$74591 ( \74531 , \40147 );
not \U$74592 ( \74532 , \74531 );
buf \U$74593 ( \74533 , \74532 );
buf \U$74594 ( \74534 , \74533 );
and \U$74595 ( \74535 , \74530 , \74534 );
buf \U$74596 ( \74536 , \74535 );
buf \U$74597 ( \74537 , \74536 );
not \U$74598 ( \74538 , \74537 );
buf \U$74599 ( \74539 , \74201 );
not \U$74600 ( \74540 , \74539 );
or \U$74601 ( \74541 , \74538 , \74540 );
buf \U$74602 ( \74542 , \74229 );
buf \U$74603 ( \74543 , \74533 );
nand \U$74604 ( \74544 , \74542 , \74543 );
buf \U$74605 ( \74545 , \74544 );
buf \U$74606 ( \74546 , \74545 );
nand \U$74607 ( \74547 , \74541 , \74546 );
buf \U$74608 ( \74548 , \74547 );
buf \U$74609 ( \74549 , \74548 );
not \U$74610 ( \74550 , \74549 );
or \U$74611 ( \74551 , \74521 , \74550 );
buf \U$74612 ( \74552 , \43665 );
buf \U$74613 ( \74553 , \74519 );
and \U$74614 ( \74554 , \74552 , \74553 );
buf \U$74615 ( \74555 , \43674 );
not \U$74616 ( \74556 , \74555 );
buf \U$74617 ( \74557 , \74556 );
buf \U$74618 ( \74558 , \74557 );
nor \U$74619 ( \74559 , \74554 , \74558 );
buf \U$74620 ( \74560 , \74559 );
buf \U$74621 ( \74561 , \74560 );
nand \U$74622 ( \74562 , \74551 , \74561 );
buf \U$74623 ( \74563 , \74562 );
buf \U$74624 ( \74564 , \74563 );
buf \U$74625 ( \74565 , \43680 );
buf \U$74626 ( \74566 , \41605 );
nor \U$74627 ( \74567 , \74565 , \74566 );
buf \U$74628 ( \74568 , \74567 );
buf \U$74629 ( \74569 , \74568 );
and \U$74630 ( \74570 , \74564 , \74569 );
not \U$74631 ( \74571 , \74564 );
buf \U$74632 ( \74572 , \74568 );
not \U$74633 ( \74573 , \74572 );
buf \U$74634 ( \74574 , \74573 );
buf \U$74635 ( \74575 , \74574 );
and \U$74636 ( \74576 , \74571 , \74575 );
nor \U$74637 ( \74577 , \74570 , \74576 );
buf \U$74638 ( \74578 , \74577 );
buf \U$74639 ( \74579 , \74578 );
buf \U$74640 ( \74580 , \74548 );
buf \U$74641 ( \74581 , \43665 );
nor \U$74642 ( \74582 , \74580 , \74581 );
buf \U$74643 ( \74583 , \74582 );
buf \U$74644 ( \74584 , \74583 );
buf \U$74645 ( \74585 , \74557 );
not \U$74646 ( \74586 , \74585 );
buf \U$74647 ( \74587 , \74519 );
nand \U$74648 ( \74588 , \74586 , \74587 );
buf \U$74649 ( \74589 , \74588 );
buf \U$74650 ( \74590 , \74589 );
and \U$74651 ( \74591 , \74584 , \74590 );
not \U$74652 ( \74592 , \74584 );
buf \U$74653 ( \74593 , \74589 );
not \U$74654 ( \74594 , \74593 );
buf \U$74655 ( \74595 , \74594 );
buf \U$74656 ( \74596 , \74595 );
and \U$74657 ( \74597 , \74592 , \74596 );
nor \U$74658 ( \74598 , \74591 , \74597 );
buf \U$74659 ( \74599 , \74598 );
buf \U$74660 ( \74600 , \74599 );
buf \U$74661 ( \74601 , \40144 );
not \U$74662 ( \74602 , \74601 );
buf \U$74663 ( \74603 , \74529 );
not \U$74664 ( \74604 , \74603 );
buf \U$74665 ( \74605 , \74201 );
not \U$74666 ( \74606 , \74605 );
or \U$74667 ( \74607 , \74604 , \74606 );
buf \U$74668 ( \74608 , \74229 );
not \U$74669 ( \74609 , \74608 );
buf \U$74670 ( \74610 , \74609 );
buf \U$74671 ( \74611 , \74610 );
nand \U$74672 ( \74612 , \74607 , \74611 );
buf \U$74673 ( \74613 , \74612 );
buf \U$74674 ( \74614 , \74613 );
not \U$74675 ( \74615 , \74614 );
or \U$74676 ( \74616 , \74602 , \74615 );
buf \U$74677 ( \74617 , \43655 );
nand \U$74678 ( \74618 , \74616 , \74617 );
buf \U$74679 ( \74619 , \74618 );
buf \U$74680 ( \74620 , \74619 );
buf \U$74681 ( \74621 , \43647 );
not \U$74682 ( \74622 , \74621 );
buf \U$74683 ( \74623 , \43662 );
nand \U$74684 ( \74624 , \74622 , \74623 );
buf \U$74685 ( \74625 , \74624 );
buf \U$74686 ( \74626 , \74625 );
not \U$74687 ( \74627 , \74626 );
buf \U$74688 ( \74628 , \74627 );
buf \U$74689 ( \74629 , \74628 );
and \U$74690 ( \74630 , \74620 , \74629 );
not \U$74691 ( \74631 , \74620 );
buf \U$74692 ( \74632 , \74625 );
and \U$74693 ( \74633 , \74631 , \74632 );
nor \U$74694 ( \74634 , \74630 , \74633 );
buf \U$74695 ( \74635 , \74634 );
buf \U$74696 ( \74636 , \74635 );
buf \U$74697 ( \74637 , \43655 );
buf \U$74698 ( \74638 , \40144 );
nand \U$74699 ( \74639 , \74637 , \74638 );
buf \U$74700 ( \74640 , \74639 );
buf \U$74701 ( \74641 , \74640 );
not \U$74702 ( \74642 , \74641 );
buf \U$74703 ( \74643 , \74613 );
not \U$74704 ( \74644 , \74643 );
or \U$74705 ( \74645 , \74642 , \74644 );
buf \U$74706 ( \74646 , \74640 );
buf \U$74707 ( \74647 , \74613 );
or \U$74708 ( \74648 , \74646 , \74647 );
nand \U$74709 ( \74649 , \74645 , \74648 );
buf \U$74710 ( \74650 , \74649 );
buf \U$74711 ( \74651 , \74650 );
buf \U$74712 ( \74652 , \74525 );
not \U$74713 ( \74653 , \74652 );
buf \U$74714 ( \74654 , \74284 );
not \U$74715 ( \74655 , \74654 );
or \U$74716 ( \74656 , \74653 , \74655 );
buf \U$74717 ( \74657 , \74223 );
not \U$74718 ( \74658 , \74657 );
buf \U$74719 ( \74659 , \74658 );
buf \U$74720 ( \74660 , \74659 );
nand \U$74721 ( \74661 , \74656 , \74660 );
buf \U$74722 ( \74662 , \74661 );
buf \U$74723 ( \74663 , \74662 );
buf \U$74724 ( \74664 , \41945 );
buf \U$74725 ( \74665 , \43635 );
nand \U$74726 ( \74666 , \74664 , \74665 );
buf \U$74727 ( \74667 , \74666 );
buf \U$74728 ( \74668 , \74667 );
not \U$74729 ( \74669 , \74668 );
buf \U$74730 ( \74670 , \74669 );
buf \U$74731 ( \74671 , \74670 );
and \U$74732 ( \74672 , \74663 , \74671 );
not \U$74733 ( \74673 , \74663 );
buf \U$74734 ( \74674 , \74667 );
and \U$74735 ( \74675 , \74673 , \74674 );
nor \U$74736 ( \74676 , \74672 , \74675 );
buf \U$74737 ( \74677 , \74676 );
buf \U$74738 ( \74678 , \74677 );
buf \U$74739 ( \74679 , \41895 );
not \U$74740 ( \74680 , \74679 );
buf \U$74741 ( \74681 , \74284 );
not \U$74742 ( \74682 , \74681 );
or \U$74743 ( \74683 , \74680 , \74682 );
buf \U$74744 ( \74684 , \43608 );
not \U$74745 ( \74685 , \74684 );
buf \U$74746 ( \74686 , \74685 );
buf \U$74747 ( \74687 , \74686 );
nand \U$74748 ( \74688 , \74683 , \74687 );
buf \U$74749 ( \74689 , \74688 );
buf \U$74750 ( \74690 , \74689 );
buf \U$74751 ( \74691 , \41968 );
buf \U$74752 ( \74692 , \74220 );
nand \U$74753 ( \74693 , \74691 , \74692 );
buf \U$74754 ( \74694 , \74693 );
buf \U$74755 ( \74695 , \74694 );
not \U$74756 ( \74696 , \74695 );
buf \U$74757 ( \74697 , \74696 );
buf \U$74758 ( \74698 , \74697 );
and \U$74759 ( \74699 , \74690 , \74698 );
not \U$74760 ( \74700 , \74690 );
buf \U$74761 ( \74701 , \74694 );
and \U$74762 ( \74702 , \74700 , \74701 );
nor \U$74763 ( \74703 , \74699 , \74702 );
buf \U$74764 ( \74704 , \74703 );
buf \U$74765 ( \74705 , \74704 );
buf \U$74766 ( \74706 , \41892 );
not \U$74767 ( \74707 , \74706 );
buf \U$74768 ( \74708 , \74284 );
not \U$74769 ( \74709 , \74708 );
or \U$74770 ( \74710 , \74707 , \74709 );
buf \U$74771 ( \74711 , \43594 );
nand \U$74772 ( \74712 , \74710 , \74711 );
buf \U$74773 ( \74713 , \74712 );
buf \U$74774 ( \74714 , \74713 );
buf \U$74775 ( \74715 , \43605 );
buf \U$74776 ( \74716 , \43597 );
nand \U$74777 ( \74717 , \74715 , \74716 );
buf \U$74778 ( \74718 , \74717 );
buf \U$74779 ( \74719 , \74718 );
not \U$74780 ( \74720 , \74719 );
buf \U$74781 ( \74721 , \74720 );
buf \U$74782 ( \74722 , \74721 );
and \U$74783 ( \74723 , \74714 , \74722 );
not \U$74784 ( \74724 , \74714 );
buf \U$74785 ( \74725 , \74718 );
and \U$74786 ( \74726 , \74724 , \74725 );
nor \U$74787 ( \74727 , \74723 , \74726 );
buf \U$74788 ( \74728 , \74727 );
buf \U$74789 ( \74729 , \74728 );
buf \U$74790 ( \74730 , \74201 );
not \U$74791 ( \74731 , \74730 );
buf \U$74792 ( \74732 , \74731 );
buf \U$74793 ( \74733 , \74732 );
not \U$74794 ( \74734 , \74733 );
buf \U$74795 ( \74735 , \41892 );
buf \U$74796 ( \74736 , \43594 );
and \U$74797 ( \74737 , \74735 , \74736 );
buf \U$74798 ( \74738 , \74737 );
buf \U$74799 ( \74739 , \74738 );
not \U$74800 ( \74740 , \74739 );
or \U$74801 ( \74741 , \74734 , \74740 );
buf \U$74802 ( \74742 , \74738 );
buf \U$74803 ( \74743 , \74732 );
or \U$74804 ( \74744 , \74742 , \74743 );
nand \U$74805 ( \74745 , \74741 , \74744 );
buf \U$74806 ( \74746 , \74745 );
buf \U$74807 ( \74747 , \74746 );
buf \U$74808 ( \74748 , \43767 );
not \U$74809 ( \74749 , \74748 );
buf \U$74810 ( \74750 , \72660 );
not \U$74811 ( \74751 , \74750 );
or \U$74812 ( \74752 , \74749 , \74751 );
buf \U$74813 ( \74753 , \27849 );
buf \U$74814 ( \74754 , \35325 );
and \U$74815 ( \74755 , \74753 , \74754 );
buf \U$74816 ( \74756 , \74755 );
buf \U$74817 ( \74757 , \74756 );
nand \U$74818 ( \74758 , \74752 , \74757 );
buf \U$74819 ( \74759 , \74758 );
buf \U$74820 ( \74760 , \74759 );
buf \U$74821 ( \74761 , \35415 );
buf \U$74822 ( \74762 , \74761 );
buf \U$74823 ( \74763 , \35464 );
buf \U$74824 ( \74764 , \35497 );
and \U$74825 ( \74765 , \74762 , \74763 , \74764 );
buf \U$74826 ( \74766 , \74765 );
buf \U$74827 ( \74767 , \74766 );
buf \U$74828 ( \74768 , \35513 );
and \U$74829 ( \74769 , \74767 , \74768 );
buf \U$74830 ( \74770 , \74769 );
buf \U$74831 ( \74771 , \74770 );
buf \U$74832 ( \74772 , \35338 );
not \U$74833 ( \74773 , \74772 );
buf \U$74834 ( \74774 , \74773 );
buf \U$74835 ( \74775 , \74774 );
buf \U$74838 ( \74776 , \33620 );
buf \U$74839 ( \74777 , \74776 );
nand \U$74840 ( \74778 , \74760 , \74771 , \74775 , \74777 );
buf \U$74841 ( \74779 , \74778 );
buf \U$74842 ( \74780 , \74779 );
buf \U$74843 ( \74781 , \74776 );
not \U$74844 ( \74782 , \74781 );
buf \U$74845 ( \74783 , \74774 );
not \U$74846 ( \74784 , \74783 );
buf \U$74849 ( \74785 , \35563 );
buf \U$74850 ( \74786 , \74785 );
not \U$74851 ( \74787 , \74786 );
or \U$74852 ( \74788 , \74784 , \74787 );
buf \U$74853 ( \74789 , \35255 );
not \U$74854 ( \74790 , \74789 );
buf \U$74855 ( \74791 , \74790 );
buf \U$74856 ( \74792 , \74791 );
nand \U$74857 ( \74793 , \74788 , \74792 );
buf \U$74858 ( \74794 , \74793 );
buf \U$74859 ( \74795 , \74794 );
not \U$74860 ( \74796 , \74795 );
or \U$74861 ( \74797 , \74782 , \74796 );
buf \U$74862 ( \74798 , \35264 );
not \U$74863 ( \74799 , \74798 );
buf \U$74864 ( \74800 , \74799 );
buf \U$74865 ( \74801 , \74800 );
nand \U$74866 ( \74802 , \74797 , \74801 );
buf \U$74867 ( \74803 , \74802 );
buf \U$74868 ( \74804 , \74803 );
not \U$74869 ( \74805 , \74804 );
buf \U$74870 ( \74806 , \74805 );
buf \U$74871 ( \74807 , \74806 );
nand \U$74872 ( \74808 , \74780 , \74807 );
buf \U$74873 ( \74809 , \74808 );
buf \U$74874 ( \74810 , \74809 );
buf \U$74875 ( \74811 , \34578 );
not \U$74876 ( \74812 , \74811 );
buf \U$74877 ( \74813 , \35276 );
nor \U$74878 ( \74814 , \74812 , \74813 );
buf \U$74879 ( \74815 , \74814 );
buf \U$74880 ( \74816 , \74815 );
and \U$74881 ( \74817 , \74810 , \74816 );
not \U$74882 ( \74818 , \74810 );
buf \U$74883 ( \74819 , \74815 );
not \U$74884 ( \74820 , \74819 );
buf \U$74885 ( \74821 , \74820 );
buf \U$74886 ( \74822 , \74821 );
and \U$74887 ( \74823 , \74818 , \74822 );
nor \U$74888 ( \74824 , \74817 , \74823 );
buf \U$74889 ( \74825 , \74824 );
buf \U$74890 ( \74826 , \74825 );
buf \U$74891 ( \74827 , \74774 );
not \U$74892 ( \74828 , \74827 );
buf \U$74893 ( \74829 , \74759 );
buf \U$74894 ( \74830 , \74770 );
and \U$74895 ( \74831 , \74829 , \74830 );
buf \U$74896 ( \74832 , \74831 );
buf \U$74897 ( \74833 , \74832 );
not \U$74898 ( \74834 , \74833 );
or \U$74899 ( \74835 , \74828 , \74834 );
buf \U$74900 ( \74836 , \74794 );
not \U$74901 ( \74837 , \74836 );
buf \U$74902 ( \74838 , \74837 );
buf \U$74903 ( \74839 , \74838 );
nand \U$74904 ( \74840 , \74835 , \74839 );
buf \U$74905 ( \74841 , \74840 );
buf \U$74906 ( \74842 , \74841 );
buf \U$74907 ( \74843 , \74800 );
buf \U$74908 ( \74844 , \74776 );
nand \U$74909 ( \74845 , \74843 , \74844 );
buf \U$74910 ( \74846 , \74845 );
buf \U$74911 ( \74847 , \74846 );
not \U$74912 ( \74848 , \74847 );
buf \U$74913 ( \74849 , \74848 );
buf \U$74914 ( \74850 , \74849 );
and \U$74915 ( \74851 , \74842 , \74850 );
not \U$74916 ( \74852 , \74842 );
buf \U$74917 ( \74853 , \74846 );
and \U$74918 ( \74854 , \74852 , \74853 );
nor \U$74919 ( \74855 , \74851 , \74854 );
buf \U$74920 ( \74856 , \74855 );
buf \U$74921 ( \74857 , \74856 );
buf \U$74922 ( \74858 , \35335 );
not \U$74923 ( \74859 , \74858 );
buf \U$74924 ( \74860 , \74832 );
not \U$74925 ( \74861 , \74860 );
or \U$74926 ( \74862 , \74859 , \74861 );
buf \U$74927 ( \74863 , \74785 );
buf \U$74928 ( \74864 , \35335 );
and \U$74929 ( \74865 , \74863 , \74864 );
buf \U$74930 ( \74866 , \35181 );
nor \U$74931 ( \74867 , \74865 , \74866 );
buf \U$74932 ( \74868 , \74867 );
buf \U$74933 ( \74869 , \74868 );
nand \U$74934 ( \74870 , \74862 , \74869 );
buf \U$74935 ( \74871 , \74870 );
buf \U$74936 ( \74872 , \74871 );
buf \U$74937 ( \74873 , \35252 );
buf \U$74938 ( \74874 , \35243 );
nand \U$74939 ( \74875 , \74873 , \74874 );
buf \U$74940 ( \74876 , \74875 );
buf \U$74941 ( \74877 , \74876 );
not \U$74942 ( \74878 , \74877 );
buf \U$74943 ( \74879 , \74878 );
buf \U$74944 ( \74880 , \74879 );
and \U$74945 ( \74881 , \74872 , \74880 );
not \U$74946 ( \74882 , \74872 );
buf \U$74947 ( \74883 , \74876 );
and \U$74948 ( \74884 , \74882 , \74883 );
nor \U$74949 ( \74885 , \74881 , \74884 );
buf \U$74950 ( \74886 , \74885 );
buf \U$74951 ( \74887 , \74886 );
buf \U$74952 ( \74888 , \74770 );
not \U$74953 ( \74889 , \74888 );
buf \U$74954 ( \74890 , \74759 );
not \U$74955 ( \74891 , \74890 );
or \U$74956 ( \74892 , \74889 , \74891 );
buf \U$74957 ( \74893 , \74785 );
not \U$74958 ( \74894 , \74893 );
buf \U$74959 ( \74895 , \74894 );
buf \U$74960 ( \74896 , \74895 );
nand \U$74961 ( \74897 , \74892 , \74896 );
buf \U$74962 ( \74898 , \74897 );
buf \U$74963 ( \74899 , \74898 );
buf \U$74964 ( \74900 , \35181 );
not \U$74965 ( \74901 , \74900 );
buf \U$74966 ( \74902 , \35335 );
nand \U$74967 ( \74903 , \74901 , \74902 );
buf \U$74968 ( \74904 , \74903 );
buf \U$74969 ( \74905 , \74904 );
not \U$74970 ( \74906 , \74905 );
buf \U$74971 ( \74907 , \74906 );
buf \U$74972 ( \74908 , \74907 );
and \U$74973 ( \74909 , \74899 , \74908 );
not \U$74974 ( \74910 , \74899 );
buf \U$74975 ( \74911 , \74904 );
and \U$74976 ( \74912 , \74910 , \74911 );
nor \U$74977 ( \74913 , \74909 , \74912 );
buf \U$74978 ( \74914 , \74913 );
buf \U$74979 ( \74915 , \74914 );
buf \U$74980 ( \74916 , \74766 );
not \U$74981 ( \74917 , \74916 );
buf \U$74982 ( \74918 , \74759 );
not \U$74983 ( \74919 , \74918 );
or \U$74984 ( \74920 , \74917 , \74919 );
buf \U$74985 ( \74921 , \35552 );
not \U$74986 ( \74922 , \74921 );
buf \U$74987 ( \74923 , \74922 );
buf \U$74988 ( \74924 , \74923 );
nand \U$74989 ( \74925 , \74920 , \74924 );
buf \U$74990 ( \74926 , \74925 );
buf \U$74991 ( \74927 , \74926 );
buf \U$74992 ( \74928 , \35513 );
buf \U$74993 ( \74929 , \35560 );
nand \U$74994 ( \74930 , \74928 , \74929 );
buf \U$74995 ( \74931 , \74930 );
buf \U$74996 ( \74932 , \74931 );
not \U$74997 ( \74933 , \74932 );
buf \U$74998 ( \74934 , \74933 );
buf \U$74999 ( \74935 , \74934 );
and \U$75000 ( \74936 , \74927 , \74935 );
not \U$75001 ( \74937 , \74927 );
buf \U$75002 ( \74938 , \74931 );
and \U$75003 ( \74939 , \74937 , \74938 );
nor \U$75004 ( \74940 , \74936 , \74939 );
buf \U$75005 ( \74941 , \74940 );
buf \U$75006 ( \74942 , \74941 );
buf \U$75007 ( \74943 , \35467 );
not \U$75008 ( \74944 , \74943 );
buf \U$75009 ( \74945 , \74759 );
not \U$75010 ( \74946 , \74945 );
or \U$75011 ( \74947 , \74944 , \74946 );
buf \U$75012 ( \74948 , \35530 );
not \U$75013 ( \74949 , \74948 );
buf \U$75014 ( \74950 , \74949 );
buf \U$75015 ( \74951 , \74950 );
not \U$75016 ( \74952 , \74951 );
buf \U$75017 ( \74953 , \35539 );
not \U$75018 ( \74954 , \74953 );
or \U$75019 ( \74955 , \74952 , \74954 );
buf \U$75020 ( \74956 , \35464 );
nand \U$75021 ( \74957 , \74955 , \74956 );
buf \U$75022 ( \74958 , \74957 );
buf \U$75023 ( \74959 , \74958 );
nand \U$75024 ( \74960 , \74947 , \74959 );
buf \U$75025 ( \74961 , \74960 );
buf \U$75026 ( \74962 , \74961 );
buf \U$75027 ( \74963 , \35497 );
buf \U$75028 ( \74964 , \35549 );
nand \U$75029 ( \74965 , \74963 , \74964 );
buf \U$75030 ( \74966 , \74965 );
buf \U$75031 ( \74967 , \74966 );
not \U$75032 ( \74968 , \74967 );
buf \U$75033 ( \74969 , \74968 );
buf \U$75034 ( \74970 , \74969 );
and \U$75035 ( \74971 , \74962 , \74970 );
not \U$75036 ( \74972 , \74962 );
buf \U$75037 ( \74973 , \74966 );
and \U$75038 ( \74974 , \74972 , \74973 );
nor \U$75039 ( \74975 , \74971 , \74974 );
buf \U$75040 ( \74976 , \74975 );
buf \U$75041 ( \74977 , \74976 );
buf \U$75042 ( \74978 , \74761 );
not \U$75043 ( \74979 , \74978 );
buf \U$75044 ( \74980 , \74759 );
not \U$75045 ( \74981 , \74980 );
or \U$75046 ( \74982 , \74979 , \74981 );
buf \U$75047 ( \74983 , \74950 );
nand \U$75048 ( \74984 , \74982 , \74983 );
buf \U$75049 ( \74985 , \74984 );
buf \U$75050 ( \74986 , \74985 );
buf \U$75051 ( \74987 , \35464 );
buf \U$75052 ( \74988 , \35539 );
nand \U$75053 ( \74989 , \74987 , \74988 );
buf \U$75054 ( \74990 , \74989 );
buf \U$75055 ( \74991 , \74990 );
not \U$75056 ( \74992 , \74991 );
buf \U$75057 ( \74993 , \74992 );
buf \U$75058 ( \74994 , \74993 );
and \U$75059 ( \74995 , \74986 , \74994 );
not \U$75060 ( \74996 , \74986 );
buf \U$75061 ( \74997 , \74990 );
and \U$75062 ( \74998 , \74996 , \74997 );
nor \U$75063 ( \74999 , \74995 , \74998 );
buf \U$75064 ( \75000 , \74999 );
buf \U$75065 ( \75001 , \75000 );
buf \U$75066 ( \75002 , \74950 );
buf \U$75067 ( \75003 , \74761 );
nand \U$75068 ( \75004 , \75002 , \75003 );
buf \U$75069 ( \75005 , \75004 );
buf \U$75070 ( \75006 , \75005 );
not \U$75071 ( \75007 , \75006 );
buf \U$75072 ( \75008 , \74759 );
not \U$75073 ( \75009 , \75008 );
or \U$75074 ( \75010 , \75007 , \75009 );
buf \U$75075 ( \75011 , \74759 );
buf \U$75076 ( \75012 , \75005 );
or \U$75077 ( \75013 , \75011 , \75012 );
nand \U$75078 ( \75014 , \75010 , \75013 );
buf \U$75079 ( \75015 , \75014 );
buf \U$75080 ( \75016 , \75015 );
buf \U$75081 ( \75017 , \43750 );
buf \U$75082 ( \75018 , \26954 );
and \U$75083 ( \75019 , \75017 , \75018 );
buf \U$75084 ( \75020 , \75019 );
buf \U$75085 ( \75021 , \75020 );
not \U$75086 ( \75022 , \75021 );
buf \U$75087 ( \75023 , \23729 );
buf \U$75088 ( \75024 , \43764 );
buf \U$75089 ( \75025 , \75024 );
and \U$75090 ( \75026 , \75023 , \75025 );
buf \U$75091 ( \75027 , \75026 );
buf \U$75092 ( \75028 , \75027 );
not \U$75093 ( \75029 , \75028 );
buf \U$75094 ( \75030 , \72660 );
buf \U$75095 ( \75031 , \75030 );
not \U$75096 ( \75032 , \75031 );
or \U$75097 ( \75033 , \75029 , \75032 );
buf \U$75098 ( \75034 , \23756 );
not \U$75099 ( \75035 , \75034 );
buf \U$75100 ( \75036 , \75035 );
buf \U$75101 ( \75037 , \75036 );
nand \U$75102 ( \75038 , \75033 , \75037 );
buf \U$75103 ( \75039 , \75038 );
buf \U$75104 ( \75040 , \75039 );
not \U$75105 ( \75041 , \75040 );
or \U$75106 ( \75042 , \75022 , \75041 );
buf \U$75107 ( \75043 , \35311 );
buf \U$75108 ( \75044 , \35293 );
buf \U$75109 ( \75045 , \75044 );
nand \U$75110 ( \75046 , \75043 , \75045 );
buf \U$75111 ( \75047 , \75046 );
buf \U$75112 ( \75048 , \75047 );
buf \U$75113 ( \75049 , \26954 );
and \U$75114 ( \75050 , \75048 , \75049 );
buf \U$75115 ( \75051 , \35285 );
not \U$75116 ( \75052 , \75051 );
buf \U$75117 ( \75053 , \75052 );
buf \U$75118 ( \75054 , \75053 );
nor \U$75119 ( \75055 , \75050 , \75054 );
buf \U$75120 ( \75056 , \75055 );
buf \U$75121 ( \75057 , \75056 );
nand \U$75122 ( \75058 , \75042 , \75057 );
buf \U$75123 ( \75059 , \75058 );
buf \U$75124 ( \75060 , \75059 );
buf \U$75125 ( \75061 , \27840 );
buf \U$75126 ( \75062 , \35298 );
nand \U$75127 ( \75063 , \75061 , \75062 );
buf \U$75128 ( \75064 , \75063 );
buf \U$75129 ( \75065 , \75064 );
not \U$75130 ( \75066 , \75065 );
buf \U$75131 ( \75067 , \75066 );
buf \U$75132 ( \75068 , \75067 );
and \U$75133 ( \75069 , \75060 , \75068 );
not \U$75134 ( \75070 , \75060 );
buf \U$75135 ( \75071 , \75064 );
and \U$75136 ( \75072 , \75070 , \75071 );
nor \U$75137 ( \75073 , \75069 , \75072 );
buf \U$75138 ( \75074 , \75073 );
buf \U$75139 ( \75075 , \75074 );
buf \U$75140 ( \75076 , \43750 );
not \U$75141 ( \75077 , \75076 );
buf \U$75142 ( \75078 , \75039 );
not \U$75143 ( \75079 , \75078 );
or \U$75144 ( \75080 , \75077 , \75079 );
buf \U$75145 ( \75081 , \75047 );
not \U$75146 ( \75082 , \75081 );
buf \U$75147 ( \75083 , \75082 );
buf \U$75148 ( \75084 , \75083 );
nand \U$75149 ( \75085 , \75080 , \75084 );
buf \U$75150 ( \75086 , \75085 );
buf \U$75151 ( \75087 , \75086 );
buf \U$75152 ( \75088 , \26954 );
buf \U$75153 ( \75089 , \35285 );
nand \U$75154 ( \75090 , \75088 , \75089 );
buf \U$75155 ( \75091 , \75090 );
buf \U$75156 ( \75092 , \75091 );
not \U$75157 ( \75093 , \75092 );
buf \U$75158 ( \75094 , \75093 );
buf \U$75159 ( \75095 , \75094 );
and \U$75160 ( \75096 , \75087 , \75095 );
not \U$75161 ( \75097 , \75087 );
buf \U$75162 ( \75098 , \75091 );
and \U$75163 ( \75099 , \75097 , \75098 );
nor \U$75164 ( \75100 , \75096 , \75099 );
buf \U$75165 ( \75101 , \75100 );
buf \U$75166 ( \75102 , \75101 );
buf \U$75167 ( \75103 , \24891 );
not \U$75168 ( \75104 , \75103 );
buf \U$75169 ( \75105 , \75039 );
not \U$75170 ( \75106 , \75105 );
or \U$75171 ( \75107 , \75104 , \75106 );
buf \U$75172 ( \75108 , \35308 );
not \U$75173 ( \75109 , \75108 );
buf \U$75174 ( \75110 , \75109 );
buf \U$75175 ( \75111 , \75110 );
nand \U$75176 ( \75112 , \75107 , \75111 );
buf \U$75177 ( \75113 , \75112 );
buf \U$75178 ( \75114 , \75113 );
buf \U$75179 ( \75115 , \75044 );
buf \U$75180 ( \75116 , \25929 );
nand \U$75181 ( \75117 , \75115 , \75116 );
buf \U$75182 ( \75118 , \75117 );
buf \U$75183 ( \75119 , \75118 );
not \U$75184 ( \75120 , \75119 );
buf \U$75185 ( \75121 , \75120 );
buf \U$75186 ( \75122 , \75121 );
and \U$75187 ( \75123 , \75114 , \75122 );
not \U$75188 ( \75124 , \75114 );
buf \U$75189 ( \75125 , \75118 );
and \U$75190 ( \75126 , \75124 , \75125 );
nor \U$75191 ( \75127 , \75123 , \75126 );
buf \U$75192 ( \75128 , \75127 );
buf \U$75193 ( \75129 , \75128 );
buf \U$75194 ( \75130 , \75110 );
buf \U$75195 ( \75131 , \24891 );
nand \U$75196 ( \75132 , \75130 , \75131 );
buf \U$75197 ( \75133 , \75132 );
buf \U$75198 ( \75134 , \75133 );
not \U$75199 ( \75135 , \75134 );
buf \U$75200 ( \75136 , \75039 );
not \U$75201 ( \75137 , \75136 );
or \U$75202 ( \75138 , \75135 , \75137 );
buf \U$75203 ( \75139 , \75133 );
buf \U$75204 ( \75140 , \75039 );
or \U$75205 ( \75141 , \75139 , \75140 );
nand \U$75206 ( \75142 , \75138 , \75141 );
buf \U$75207 ( \75143 , \75142 );
buf \U$75208 ( \75144 , \75143 );
buf \U$75209 ( \75145 , \23726 );
not \U$75210 ( \75146 , \75145 );
buf \U$75211 ( \75147 , \75024 );
not \U$75212 ( \75148 , \75147 );
buf \U$75213 ( \75149 , \75030 );
not \U$75214 ( \75150 , \75149 );
or \U$75215 ( \75151 , \75148 , \75150 );
buf \U$75216 ( \75152 , \21571 );
not \U$75217 ( \75153 , \75152 );
buf \U$75218 ( \75154 , \20364 );
not \U$75219 ( \75155 , \75154 );
and \U$75220 ( \75156 , \75153 , \75155 );
buf \U$75221 ( \75157 , \21561 );
not \U$75222 ( \75158 , \75157 );
buf \U$75223 ( \75159 , \75158 );
buf \U$75224 ( \75160 , \75159 );
nor \U$75225 ( \75161 , \75156 , \75160 );
buf \U$75226 ( \75162 , \75161 );
buf \U$75227 ( \75163 , \75162 );
nand \U$75228 ( \75164 , \75151 , \75163 );
buf \U$75229 ( \75165 , \75164 );
buf \U$75230 ( \75166 , \75165 );
not \U$75231 ( \75167 , \75166 );
or \U$75232 ( \75168 , \75146 , \75167 );
buf \U$75233 ( \75169 , \23737 );
not \U$75234 ( \75170 , \75169 );
buf \U$75235 ( \75171 , \75170 );
buf \U$75236 ( \75172 , \75171 );
nand \U$75237 ( \75173 , \75168 , \75172 );
buf \U$75238 ( \75174 , \75173 );
buf \U$75239 ( \75175 , \75174 );
buf \U$75240 ( \75176 , \23713 );
buf \U$75241 ( \75177 , \23749 );
nand \U$75242 ( \75178 , \75176 , \75177 );
buf \U$75243 ( \75179 , \75178 );
buf \U$75244 ( \75180 , \75179 );
not \U$75245 ( \75181 , \75180 );
buf \U$75246 ( \75182 , \75181 );
buf \U$75247 ( \75183 , \75182 );
and \U$75248 ( \75184 , \75175 , \75183 );
not \U$75249 ( \75185 , \75175 );
buf \U$75250 ( \75186 , \75179 );
and \U$75251 ( \75187 , \75185 , \75186 );
nor \U$75252 ( \75188 , \75184 , \75187 );
buf \U$75253 ( \75189 , \75188 );
buf \U$75254 ( \75190 , \75189 );
buf \U$75255 ( \75191 , \75171 );
buf \U$75256 ( \75192 , \23726 );
nand \U$75257 ( \75193 , \75191 , \75192 );
buf \U$75258 ( \75194 , \75193 );
buf \U$75259 ( \75195 , \75194 );
not \U$75260 ( \75196 , \75195 );
buf \U$75261 ( \75197 , \75165 );
not \U$75262 ( \75198 , \75197 );
or \U$75263 ( \75199 , \75196 , \75198 );
buf \U$75264 ( \75200 , \75194 );
buf \U$75265 ( \75201 , \75165 );
or \U$75266 ( \75202 , \75200 , \75201 );
nand \U$75267 ( \75203 , \75199 , \75202 );
buf \U$75268 ( \75204 , \75203 );
buf \U$75269 ( \75205 , \75204 );
buf \U$75270 ( \75206 , \43761 );
not \U$75271 ( \75207 , \75206 );
buf \U$75272 ( \75208 , \75030 );
not \U$75273 ( \75209 , \75208 );
or \U$75274 ( \75210 , \75207 , \75209 );
buf \U$75275 ( \75211 , \20364 );
nand \U$75276 ( \75212 , \75210 , \75211 );
buf \U$75277 ( \75213 , \75212 );
buf \U$75278 ( \75214 , \75213 );
buf \U$75279 ( \75215 , \21568 );
buf \U$75280 ( \75216 , \21561 );
nand \U$75281 ( \75217 , \75215 , \75216 );
buf \U$75282 ( \75218 , \75217 );
buf \U$75283 ( \75219 , \75218 );
not \U$75284 ( \75220 , \75219 );
buf \U$75285 ( \75221 , \75220 );
buf \U$75286 ( \75222 , \75221 );
and \U$75287 ( \75223 , \75214 , \75222 );
not \U$75288 ( \75224 , \75214 );
buf \U$75289 ( \75225 , \75218 );
and \U$75290 ( \75226 , \75224 , \75225 );
nor \U$75291 ( \75227 , \75223 , \75226 );
buf \U$75292 ( \75228 , \75227 );
buf \U$75293 ( \75229 , \75228 );
buf \U$75294 ( \75230 , \20364 );
buf \U$75295 ( \75231 , \43761 );
nand \U$75296 ( \75232 , \75230 , \75231 );
buf \U$75297 ( \75233 , \75232 );
buf \U$75298 ( \75234 , \75233 );
buf \U$75299 ( \75235 , \75030 );
not \U$75300 ( \75236 , \75235 );
xor \U$75301 ( \75237 , \75234 , \75236 );
buf \U$75302 ( \75238 , \75237 );
buf \U$75303 ( \75239 , \75238 );
buf \U$75304 ( \75240 , \72356 );
buf \U$75305 ( \75241 , \72420 );
and \U$75306 ( \75242 , \75240 , \75241 );
buf \U$75307 ( \75243 , \75242 );
buf \U$75308 ( \75244 , \75243 );
buf \U$75309 ( \75245 , \72087 );
and \U$75310 ( \75246 , \75244 , \75245 );
buf \U$75311 ( \75247 , \75246 );
buf \U$75312 ( \75248 , \75247 );
not \U$75313 ( \75249 , \75248 );
buf \U$75314 ( \75250 , \70066 );
not \U$75315 ( \75251 , \75250 );
buf \U$75316 ( \75252 , \63019 );
not \U$75317 ( \75253 , \75252 );
or \U$75318 ( \75254 , \75251 , \75253 );
buf \U$75319 ( \75255 , \72548 );
not \U$75320 ( \75256 , \75255 );
buf \U$75321 ( \75257 , \75256 );
buf \U$75322 ( \75258 , \75257 );
nand \U$75323 ( \75259 , \75254 , \75258 );
buf \U$75324 ( \75260 , \75259 );
buf \U$75325 ( \75261 , \75260 );
not \U$75326 ( \75262 , \75261 );
or \U$75327 ( \75263 , \75249 , \75262 );
buf \U$75328 ( \75264 , \72651 );
not \U$75329 ( \75265 , \72592 );
buf \U$75330 ( \75266 , \75265 );
and \U$75331 ( \75267 , \75264 , \75266 );
buf \U$75332 ( \75268 , \75267 );
buf \U$75333 ( \75269 , \75268 );
not \U$75334 ( \75270 , \75269 );
buf \U$75335 ( \75271 , \75270 );
buf \U$75336 ( \75272 , \75271 );
buf \U$75337 ( \75273 , \75243 );
and \U$75338 ( \75274 , \75272 , \75273 );
buf \U$75339 ( \75275 , \72581 );
nor \U$75340 ( \75276 , \75274 , \75275 );
buf \U$75341 ( \75277 , \75276 );
buf \U$75342 ( \75278 , \75277 );
nand \U$75343 ( \75279 , \75263 , \75278 );
buf \U$75344 ( \75280 , \75279 );
buf \U$75345 ( \75281 , \75280 );
buf \U$75346 ( \75282 , \72601 );
buf \U$75347 ( \75283 , \72583 );
nand \U$75348 ( \75284 , \75282 , \75283 );
buf \U$75349 ( \75285 , \75284 );
buf \U$75350 ( \75286 , \75285 );
not \U$75351 ( \75287 , \75286 );
buf \U$75352 ( \75288 , \75287 );
buf \U$75353 ( \75289 , \75288 );
and \U$75354 ( \75290 , \75281 , \75289 );
not \U$75355 ( \75291 , \75281 );
buf \U$75356 ( \75292 , \75285 );
and \U$75357 ( \75293 , \75291 , \75292 );
nor \U$75358 ( \75294 , \75290 , \75293 );
buf \U$75359 ( \75295 , \75294 );
buf \U$75360 ( \75296 , \75295 );
buf \U$75361 ( \75297 , \72356 );
not \U$75362 ( \75298 , \75297 );
buf \U$75363 ( \75299 , \72087 );
not \U$75364 ( \75300 , \75299 );
buf \U$75365 ( \75301 , \75260 );
not \U$75366 ( \75302 , \75301 );
or \U$75367 ( \75303 , \75300 , \75302 );
buf \U$75368 ( \75304 , \75268 );
nand \U$75369 ( \75305 , \75303 , \75304 );
buf \U$75370 ( \75306 , \75305 );
buf \U$75371 ( \75307 , \75306 );
not \U$75372 ( \75308 , \75307 );
or \U$75373 ( \75309 , \75298 , \75308 );
buf \U$75374 ( \75310 , \72567 );
nand \U$75375 ( \75311 , \75309 , \75310 );
buf \U$75376 ( \75312 , \75311 );
buf \U$75377 ( \75313 , \75312 );
buf \U$75378 ( \75314 , \72578 );
buf \U$75379 ( \75315 , \72420 );
nand \U$75380 ( \75316 , \75314 , \75315 );
buf \U$75381 ( \75317 , \75316 );
buf \U$75382 ( \75318 , \75317 );
not \U$75383 ( \75319 , \75318 );
buf \U$75384 ( \75320 , \75319 );
buf \U$75385 ( \75321 , \75320 );
and \U$75386 ( \75322 , \75313 , \75321 );
not \U$75387 ( \75323 , \75313 );
buf \U$75388 ( \75324 , \75317 );
and \U$75389 ( \75325 , \75323 , \75324 );
nor \U$75390 ( \75326 , \75322 , \75325 );
buf \U$75391 ( \75327 , \75326 );
buf \U$75392 ( \75328 , \75327 );
buf \U$75393 ( \75329 , \72352 );
not \U$75394 ( \75330 , \75329 );
buf \U$75395 ( \75331 , \75306 );
not \U$75396 ( \75332 , \75331 );
or \U$75397 ( \75333 , \75330 , \75332 );
buf \U$75398 ( \75334 , \72564 );
nand \U$75399 ( \75335 , \75333 , \75334 );
buf \U$75400 ( \75336 , \75335 );
buf \U$75401 ( \75337 , \75336 );
buf \U$75402 ( \75338 , \72317 );
buf \U$75403 ( \75339 , \72556 );
nand \U$75404 ( \75340 , \75338 , \75339 );
buf \U$75405 ( \75341 , \75340 );
buf \U$75406 ( \75342 , \75341 );
not \U$75407 ( \75343 , \75342 );
buf \U$75408 ( \75344 , \75343 );
buf \U$75409 ( \75345 , \75344 );
and \U$75410 ( \75346 , \75337 , \75345 );
not \U$75411 ( \75347 , \75337 );
buf \U$75412 ( \75348 , \75341 );
and \U$75413 ( \75349 , \75347 , \75348 );
nor \U$75414 ( \75350 , \75346 , \75349 );
buf \U$75415 ( \75351 , \75350 );
buf \U$75416 ( \75352 , \75351 );
buf \U$75417 ( \75353 , \72564 );
buf \U$75418 ( \75354 , \72352 );
nand \U$75419 ( \75355 , \75353 , \75354 );
buf \U$75420 ( \75356 , \75355 );
buf \U$75421 ( \75357 , \75356 );
not \U$75422 ( \75358 , \75357 );
buf \U$75423 ( \75359 , \75306 );
not \U$75424 ( \75360 , \75359 );
or \U$75425 ( \75361 , \75358 , \75360 );
buf \U$75426 ( \75362 , \75356 );
buf \U$75427 ( \75363 , \75306 );
or \U$75428 ( \75364 , \75362 , \75363 );
nand \U$75429 ( \75365 , \75361 , \75364 );
buf \U$75430 ( \75366 , \75365 );
buf \U$75431 ( \75367 , \75366 );
buf \U$75432 ( \75368 , \72637 );
not \U$75433 ( \75369 , \75368 );
buf \U$75434 ( \75370 , \75369 );
buf \U$75435 ( \75371 , \75370 );
not \U$75436 ( \75372 , \75371 );
buf \U$75437 ( \75373 , \71474 );
buf \U$75438 ( \75374 , \75373 );
buf \U$75439 ( \75375 , \72083 );
and \U$75440 ( \75376 , \75374 , \75375 );
buf \U$75441 ( \75377 , \75376 );
buf \U$75442 ( \75378 , \75377 );
not \U$75443 ( \75379 , \75378 );
buf \U$75444 ( \75380 , \75260 );
not \U$75445 ( \75381 , \75380 );
or \U$75446 ( \75382 , \75379 , \75381 );
buf \U$75448 ( \75383 , \72633 );
nand \U$75449 ( \75384 , \75382 , \75383 );
buf \U$75450 ( \75385 , \75384 );
buf \U$75451 ( \75386 , \75385 );
not \U$75452 ( \75387 , \75386 );
or \U$75453 ( \75388 , \75372 , \75387 );
buf \U$75454 ( \75389 , \72643 );
nand \U$75455 ( \75390 , \75388 , \75389 );
buf \U$75456 ( \75391 , \75390 );
buf \U$75457 ( \75392 , \75391 );
buf \U$75458 ( \75393 , \72648 );
buf \U$75459 ( \75394 , \75265 );
nand \U$75460 ( \75395 , \75393 , \75394 );
buf \U$75461 ( \75396 , \75395 );
buf \U$75462 ( \75397 , \75396 );
not \U$75463 ( \75398 , \75397 );
buf \U$75464 ( \75399 , \75398 );
buf \U$75465 ( \75400 , \75399 );
and \U$75466 ( \75401 , \75392 , \75400 );
not \U$75467 ( \75402 , \75392 );
buf \U$75468 ( \75403 , \75396 );
and \U$75469 ( \75404 , \75402 , \75403 );
nor \U$75470 ( \75405 , \75401 , \75404 );
buf \U$75471 ( \75406 , \75405 );
buf \U$75472 ( \75407 , \75406 );
buf \U$75473 ( \75408 , \75370 );
buf \U$75474 ( \75409 , \72643 );
nand \U$75475 ( \75410 , \75408 , \75409 );
buf \U$75476 ( \75411 , \75410 );
buf \U$75477 ( \75412 , \75411 );
not \U$75478 ( \75413 , \75412 );
buf \U$75479 ( \75414 , \75385 );
not \U$75480 ( \75415 , \75414 );
or \U$75481 ( \75416 , \75413 , \75415 );
buf \U$75482 ( \75417 , \75411 );
buf \U$75483 ( \75418 , \75385 );
or \U$75484 ( \75419 , \75417 , \75418 );
nand \U$75485 ( \75420 , \75416 , \75419 );
buf \U$75486 ( \75421 , \75420 );
buf \U$75487 ( \75422 , \75421 );
buf \U$75488 ( \75423 , \72083 );
not \U$75489 ( \75424 , \75423 );
buf \U$75490 ( \75425 , \75260 );
not \U$75491 ( \75426 , \75425 );
or \U$75492 ( \75427 , \75424 , \75426 );
buf \U$75493 ( \75428 , \72627 );
nand \U$75494 ( \75429 , \75427 , \75428 );
buf \U$75495 ( \75430 , \75429 );
buf \U$75496 ( \75431 , \75430 );
buf \U$75497 ( \75432 , \72621 );
buf \U$75498 ( \75433 , \75373 );
nand \U$75499 ( \75434 , \75432 , \75433 );
buf \U$75500 ( \75435 , \75434 );
buf \U$75501 ( \75436 , \75435 );
not \U$75502 ( \75437 , \75436 );
buf \U$75503 ( \75438 , \75437 );
buf \U$75504 ( \75439 , \75438 );
and \U$75505 ( \75440 , \75431 , \75439 );
not \U$75506 ( \75441 , \75431 );
buf \U$75507 ( \75442 , \75435 );
and \U$75508 ( \75443 , \75441 , \75442 );
nor \U$75509 ( \75444 , \75440 , \75443 );
buf \U$75510 ( \75445 , \75444 );
buf \U$75511 ( \75446 , \75445 );
buf \U$75512 ( \75447 , \72627 );
buf \U$75513 ( \75448 , \72083 );
nand \U$75514 ( \75449 , \75447 , \75448 );
buf \U$75515 ( \75450 , \75449 );
buf \U$75516 ( \75451 , \75450 );
not \U$75517 ( \75452 , \75451 );
buf \U$75518 ( \75453 , \75260 );
not \U$75519 ( \75454 , \75453 );
or \U$75520 ( \75455 , \75452 , \75454 );
buf \U$75521 ( \75456 , \75450 );
buf \U$75522 ( \75457 , \75260 );
or \U$75523 ( \75458 , \75456 , \75457 );
nand \U$75524 ( \75459 , \75455 , \75458 );
buf \U$75525 ( \75460 , \75459 );
buf \U$75526 ( \75461 , \75460 );
buf \U$75527 ( \75462 , \69814 );
not \U$75528 ( \75463 , \75462 );
buf \U$75529 ( \75464 , \67805 );
not \U$75530 ( \75465 , \75464 );
buf \U$75531 ( \75466 , \70063 );
not \U$75532 ( \75467 , \75466 );
buf \U$75533 ( \75468 , \63019 );
not \U$75534 ( \75469 , \75468 );
or \U$75535 ( \75470 , \75467 , \75469 );
buf \U$75536 ( \75471 , \72504 );
nand \U$75537 ( \75472 , \75470 , \75471 );
buf \U$75538 ( \75473 , \75472 );
buf \U$75539 ( \75474 , \75473 );
not \U$75540 ( \75475 , \75474 );
or \U$75541 ( \75476 , \75465 , \75475 );
buf \U$75542 ( \75477 , \72518 );
not \U$75543 ( \75478 , \75477 );
buf \U$75544 ( \75479 , \67597 );
nand \U$75545 ( \75480 , \75478 , \75479 );
buf \U$75546 ( \75481 , \75480 );
buf \U$75547 ( \75482 , \75481 );
nand \U$75548 ( \75483 , \75476 , \75482 );
buf \U$75549 ( \75484 , \75483 );
buf \U$75550 ( \75485 , \75484 );
not \U$75551 ( \75486 , \75485 );
or \U$75552 ( \75487 , \75463 , \75486 );
buf \U$75553 ( \75488 , \72534 );
nand \U$75554 ( \75489 , \75487 , \75488 );
buf \U$75555 ( \75490 , \75489 );
buf \U$75556 ( \75491 , \75490 );
buf \U$75557 ( \75492 , \72529 );
buf \U$75558 ( \75493 , \72542 );
nand \U$75559 ( \75494 , \75492 , \75493 );
buf \U$75560 ( \75495 , \75494 );
buf \U$75561 ( \75496 , \75495 );
not \U$75562 ( \75497 , \75496 );
buf \U$75563 ( \75498 , \75497 );
buf \U$75564 ( \75499 , \75498 );
and \U$75565 ( \75500 , \75491 , \75499 );
not \U$75566 ( \75501 , \75491 );
buf \U$75567 ( \75502 , \75495 );
and \U$75568 ( \75503 , \75501 , \75502 );
nor \U$75569 ( \75504 , \75500 , \75503 );
buf \U$75570 ( \75505 , \75504 );
buf \U$75571 ( \75506 , \75505 );
buf \U$75572 ( \75507 , \72534 );
buf \U$75573 ( \75508 , \69814 );
nand \U$75574 ( \75509 , \75507 , \75508 );
buf \U$75575 ( \75510 , \75509 );
buf \U$75576 ( \75511 , \75510 );
not \U$75577 ( \75512 , \75511 );
buf \U$75578 ( \75513 , \75484 );
not \U$75579 ( \75514 , \75513 );
or \U$75580 ( \75515 , \75512 , \75514 );
buf \U$75581 ( \75516 , \75510 );
buf \U$75582 ( \75517 , \75484 );
or \U$75583 ( \75518 , \75516 , \75517 );
nand \U$75584 ( \75519 , \75515 , \75518 );
buf \U$75585 ( \75520 , \75519 );
buf \U$75586 ( \75521 , \75520 );
buf \U$75587 ( \75522 , \67802 );
not \U$75588 ( \75523 , \75522 );
buf \U$75589 ( \75524 , \75473 );
not \U$75590 ( \75525 , \75524 );
or \U$75591 ( \75526 , \75523 , \75525 );
buf \U$75592 ( \75527 , \72510 );
nand \U$75593 ( \75528 , \75526 , \75527 );
buf \U$75594 ( \75529 , \75528 );
buf \U$75595 ( \75530 , \75529 );
buf \U$75596 ( \75531 , \67597 );
buf \U$75597 ( \75532 , \72515 );
nand \U$75598 ( \75533 , \75531 , \75532 );
buf \U$75599 ( \75534 , \75533 );
buf \U$75600 ( \75535 , \75534 );
not \U$75601 ( \75536 , \75535 );
buf \U$75602 ( \75537 , \75536 );
buf \U$75603 ( \75538 , \75537 );
and \U$75604 ( \75539 , \75530 , \75538 );
not \U$75605 ( \75540 , \75530 );
buf \U$75606 ( \75541 , \75534 );
and \U$75607 ( \75542 , \75540 , \75541 );
nor \U$75608 ( \75543 , \75539 , \75542 );
buf \U$75609 ( \75544 , \75543 );
buf \U$75610 ( \75545 , \75544 );
buf \U$75611 ( \75546 , \72510 );
buf \U$75612 ( \75547 , \67802 );
nand \U$75613 ( \75548 , \75546 , \75547 );
buf \U$75614 ( \75549 , \75548 );
buf \U$75615 ( \75550 , \75549 );
not \U$75616 ( \75551 , \75550 );
buf \U$75617 ( \75552 , \75473 );
not \U$75618 ( \75553 , \75552 );
or \U$75619 ( \75554 , \75551 , \75553 );
buf \U$75620 ( \75555 , \75549 );
buf \U$75621 ( \75556 , \75473 );
or \U$75622 ( \75557 , \75555 , \75556 );
nand \U$75623 ( \75558 , \75554 , \75557 );
buf \U$75624 ( \75559 , \75558 );
buf \U$75625 ( \75560 , \75559 );
buf \U$75626 ( \75561 , \70010 );
not \U$75627 ( \75562 , \75561 );
buf \U$75628 ( \75563 , \70060 );
not \U$75629 ( \75564 , \75563 );
buf \U$75630 ( \75565 , \75564 );
buf \U$75631 ( \75566 , \75565 );
not \U$75632 ( \75567 , \75566 );
buf \U$75633 ( \75568 , \74192 );
not \U$75634 ( \75569 , \75568 );
or \U$75635 ( \75570 , \75567 , \75569 );
buf \U$75636 ( \75571 , \72493 );
buf \U$75637 ( \75572 , \70044 );
nand \U$75638 ( \75573 , \75571 , \75572 );
buf \U$75639 ( \75574 , \75573 );
buf \U$75640 ( \75575 , \75574 );
nand \U$75641 ( \75576 , \75570 , \75575 );
buf \U$75642 ( \75577 , \75576 );
buf \U$75643 ( \75578 , \75577 );
not \U$75644 ( \75579 , \75578 );
or \U$75645 ( \75580 , \75562 , \75579 );
buf \U$75646 ( \75581 , \72471 );
not \U$75647 ( \75582 , \75581 );
buf \U$75648 ( \75583 , \75582 );
buf \U$75649 ( \75584 , \75583 );
nand \U$75650 ( \75585 , \75580 , \75584 );
buf \U$75651 ( \75586 , \75585 );
buf \U$75652 ( \75587 , \75586 );
buf \U$75653 ( \75588 , \72476 );
not \U$75654 ( \75589 , \75588 );
buf \U$75655 ( \75590 , \69961 );
nand \U$75656 ( \75591 , \75589 , \75590 );
buf \U$75657 ( \75592 , \75591 );
buf \U$75658 ( \75593 , \75592 );
not \U$75659 ( \75594 , \75593 );
buf \U$75660 ( \75595 , \75594 );
buf \U$75661 ( \75596 , \75595 );
and \U$75662 ( \75597 , \75587 , \75596 );
not \U$75663 ( \75598 , \75587 );
buf \U$75664 ( \75599 , \75592 );
and \U$75665 ( \75600 , \75598 , \75599 );
nor \U$75666 ( \75601 , \75597 , \75600 );
buf \U$75667 ( \75602 , \75601 );
buf \U$75668 ( \75603 , \75602 );
buf \U$75669 ( \75604 , \75583 );
buf \U$75670 ( \75605 , \70010 );
nand \U$75671 ( \75606 , \75604 , \75605 );
buf \U$75672 ( \75607 , \75606 );
buf \U$75673 ( \75608 , \75607 );
not \U$75674 ( \75609 , \75608 );
buf \U$75675 ( \75610 , \75577 );
not \U$75676 ( \75611 , \75610 );
or \U$75677 ( \75612 , \75609 , \75611 );
buf \U$75678 ( \75613 , \75607 );
buf \U$75679 ( \75614 , \75577 );
or \U$75680 ( \75615 , \75613 , \75614 );
nand \U$75681 ( \75616 , \75612 , \75615 );
buf \U$75682 ( \75617 , \75616 );
buf \U$75683 ( \75618 , \75617 );
buf \U$75684 ( \75619 , \70057 );
not \U$75685 ( \75620 , \75619 );
buf \U$75686 ( \75621 , \74192 );
not \U$75687 ( \75622 , \75621 );
or \U$75688 ( \75623 , \75620 , \75622 );
buf \U$75689 ( \75624 , \72490 );
nand \U$75690 ( \75625 , \75623 , \75624 );
buf \U$75691 ( \75626 , \75625 );
buf \U$75692 ( \75627 , \75626 );
buf \U$75693 ( \75628 , \70044 );
buf \U$75694 ( \75629 , \72485 );
nand \U$75695 ( \75630 , \75628 , \75629 );
buf \U$75696 ( \75631 , \75630 );
buf \U$75697 ( \75632 , \75631 );
not \U$75698 ( \75633 , \75632 );
buf \U$75699 ( \75634 , \75633 );
buf \U$75700 ( \75635 , \75634 );
and \U$75701 ( \75636 , \75627 , \75635 );
not \U$75702 ( \75637 , \75627 );
buf \U$75703 ( \75638 , \75631 );
and \U$75704 ( \75639 , \75637 , \75638 );
nor \U$75705 ( \75640 , \75636 , \75639 );
buf \U$75706 ( \75641 , \75640 );
buf \U$75707 ( \75642 , \75641 );
buf \U$75708 ( \75643 , \72490 );
buf \U$75709 ( \75644 , \70057 );
nand \U$75710 ( \75645 , \75643 , \75644 );
buf \U$75711 ( \75646 , \75645 );
buf \U$75712 ( \75647 , \75646 );
not \U$75713 ( \75648 , \75647 );
buf \U$75714 ( \75649 , \74192 );
not \U$75715 ( \75650 , \75649 );
or \U$75716 ( \75651 , \75648 , \75650 );
buf \U$75717 ( \75652 , \75646 );
buf \U$75718 ( \75653 , \74192 );
or \U$75719 ( \75654 , \75652 , \75653 );
nand \U$75720 ( \75655 , \75651 , \75654 );
buf \U$75721 ( \75656 , \75655 );
buf \U$75722 ( \75657 , \75656 );
buf \U$75723 ( \75658 , \56423 );
not \U$75724 ( \75659 , \75658 );
and \U$75725 ( \75660 , \56436 , \56413 );
buf \U$75726 ( \75661 , \75660 );
not \U$75727 ( \75662 , \75661 );
buf \U$75728 ( \75663 , \49374 );
not \U$75729 ( \75664 , \75663 );
buf \U$75730 ( \75665 , \62972 );
not \U$75731 ( \75666 , \75665 );
buf \U$75732 ( \75667 , \56471 );
not \U$75733 ( \75668 , \75667 );
or \U$75734 ( \75669 , \75666 , \75668 );
buf \U$75735 ( \75670 , \53378 );
nand \U$75736 ( \75671 , \75669 , \75670 );
buf \U$75737 ( \75672 , \75671 );
buf \U$75738 ( \75673 , \75672 );
not \U$75739 ( \75674 , \75673 );
or \U$75740 ( \75675 , \75664 , \75674 );
buf \U$75741 ( \75676 , \53420 );
nand \U$75742 ( \75677 , \75675 , \75676 );
buf \U$75743 ( \75678 , \75677 );
buf \U$75744 ( \75679 , \75678 );
not \U$75745 ( \75680 , \75679 );
or \U$75746 ( \75681 , \75662 , \75680 );
buf \U$75747 ( \75682 , \62992 );
not \U$75748 ( \75683 , \75682 );
buf \U$75749 ( \75684 , \75683 );
buf \U$75750 ( \75685 , \75684 );
nand \U$75751 ( \75686 , \75681 , \75685 );
buf \U$75752 ( \75687 , \75686 );
buf \U$75753 ( \75688 , \75687 );
not \U$75754 ( \75689 , \75688 );
or \U$75755 ( \75690 , \75659 , \75689 );
buf \U$75756 ( \75691 , \63000 );
nand \U$75757 ( \75692 , \75690 , \75691 );
buf \U$75758 ( \75693 , \75692 );
buf \U$75759 ( \75694 , \75693 );
buf \U$75760 ( \75695 , \56355 );
buf \U$75761 ( \75696 , \63010 );
nand \U$75762 ( \75697 , \75695 , \75696 );
buf \U$75763 ( \75698 , \75697 );
buf \U$75764 ( \75699 , \75698 );
not \U$75765 ( \75700 , \75699 );
buf \U$75766 ( \75701 , \75700 );
buf \U$75767 ( \75702 , \75701 );
and \U$75768 ( \75703 , \75694 , \75702 );
not \U$75769 ( \75704 , \75694 );
buf \U$75770 ( \75705 , \75698 );
and \U$75771 ( \75706 , \75704 , \75705 );
nor \U$75772 ( \75707 , \75703 , \75706 );
buf \U$75773 ( \75708 , \75707 );
buf \U$75774 ( \75709 , \75708 );
buf \U$75775 ( \75710 , \75687 );
not \U$75776 ( \75711 , \75710 );
buf \U$75777 ( \75712 , \63000 );
buf \U$75778 ( \75713 , \56423 );
nand \U$75779 ( \75714 , \75712 , \75713 );
buf \U$75780 ( \75715 , \75714 );
buf \U$75781 ( \75716 , \75715 );
not \U$75782 ( \75717 , \75716 );
or \U$75783 ( \75718 , \75711 , \75717 );
buf \U$75784 ( \75719 , \75715 );
buf \U$75785 ( \75720 , \75687 );
or \U$75786 ( \75721 , \75719 , \75720 );
nand \U$75787 ( \75722 , \75718 , \75721 );
buf \U$75788 ( \75723 , \75722 );
buf \U$75789 ( \75724 , \75723 );
buf \U$75790 ( \75725 , \56436 );
not \U$75791 ( \75726 , \75725 );
buf \U$75792 ( \75727 , \75678 );
not \U$75793 ( \75728 , \75727 );
or \U$75794 ( \75729 , \75726 , \75728 );
buf \U$75795 ( \75730 , \62983 );
buf \U$75796 ( \75731 , \75730 );
nand \U$75797 ( \75732 , \75729 , \75731 );
buf \U$75798 ( \75733 , \75732 );
buf \U$75799 ( \75734 , \75733 );
buf \U$75800 ( \75735 , \56413 );
buf \U$75801 ( \75736 , \62989 );
nand \U$75802 ( \75737 , \75735 , \75736 );
buf \U$75803 ( \75738 , \75737 );
buf \U$75804 ( \75739 , \75738 );
not \U$75805 ( \75740 , \75739 );
buf \U$75806 ( \75741 , \75740 );
buf \U$75807 ( \75742 , \75741 );
and \U$75808 ( \75743 , \75734 , \75742 );
not \U$75809 ( \75744 , \75734 );
buf \U$75810 ( \75745 , \75738 );
and \U$75811 ( \75746 , \75744 , \75745 );
nor \U$75812 ( \75747 , \75743 , \75746 );
buf \U$75813 ( \75748 , \75747 );
buf \U$75814 ( \75749 , \75748 );
buf \U$75815 ( \75750 , \56436 );
buf \U$75816 ( \75751 , \75730 );
nand \U$75817 ( \75752 , \75750 , \75751 );
buf \U$75818 ( \75753 , \75752 );
buf \U$75819 ( \75754 , \75753 );
not \U$75820 ( \75755 , \75754 );
buf \U$75821 ( \75756 , \75678 );
not \U$75822 ( \75757 , \75756 );
or \U$75823 ( \75758 , \75755 , \75757 );
buf \U$75824 ( \75759 , \75753 );
buf \U$75825 ( \75760 , \75678 );
or \U$75826 ( \75761 , \75759 , \75760 );
nand \U$75827 ( \75762 , \75758 , \75761 );
buf \U$75828 ( \75763 , \75762 );
buf \U$75829 ( \75764 , \75763 );
buf \U$75830 ( \75765 , \47442 );
not \U$75831 ( \75766 , \75765 );
buf \U$75832 ( \75767 , \48013 );
buf \U$75833 ( \75768 , \49371 );
and \U$75834 ( \75769 , \75767 , \75768 );
buf \U$75835 ( \75770 , \75769 );
buf \U$75836 ( \75771 , \75770 );
not \U$75837 ( \75772 , \75771 );
buf \U$75838 ( \75773 , \75672 );
not \U$75839 ( \75774 , \75773 );
or \U$75840 ( \75775 , \75772 , \75774 );
buf \U$75841 ( \75776 , \53408 );
buf \U$75842 ( \75777 , \53414 );
and \U$75843 ( \75778 , \75776 , \75777 );
buf \U$75844 ( \75779 , \75778 );
buf \U$75845 ( \75780 , \75779 );
nand \U$75846 ( \75781 , \75775 , \75780 );
buf \U$75847 ( \75782 , \75781 );
buf \U$75848 ( \75783 , \75782 );
not \U$75849 ( \75784 , \75783 );
or \U$75850 ( \75785 , \75766 , \75784 );
buf \U$75851 ( \75786 , \53396 );
nand \U$75852 ( \75787 , \75785 , \75786 );
buf \U$75853 ( \75788 , \75787 );
buf \U$75854 ( \75789 , \75788 );
buf \U$75855 ( \75790 , \53387 );
buf \U$75856 ( \75791 , \48727 );
nand \U$75857 ( \75792 , \75790 , \75791 );
buf \U$75858 ( \75793 , \75792 );
buf \U$75859 ( \75794 , \75793 );
not \U$75860 ( \75795 , \75794 );
buf \U$75861 ( \75796 , \75795 );
buf \U$75862 ( \75797 , \75796 );
and \U$75863 ( \75798 , \75789 , \75797 );
not \U$75864 ( \75799 , \75789 );
buf \U$75865 ( \75800 , \75793 );
and \U$75866 ( \75801 , \75799 , \75800 );
nor \U$75867 ( \75802 , \75798 , \75801 );
buf \U$75868 ( \75803 , \75802 );
buf \U$75869 ( \75804 , \75803 );
buf \U$75870 ( \75805 , \47442 );
buf \U$75871 ( \75806 , \53396 );
nand \U$75872 ( \75807 , \75805 , \75806 );
buf \U$75873 ( \75808 , \75807 );
buf \U$75874 ( \75809 , \75808 );
not \U$75875 ( \75810 , \75809 );
buf \U$75876 ( \75811 , \75782 );
not \U$75877 ( \75812 , \75811 );
or \U$75878 ( \75813 , \75810 , \75812 );
buf \U$75879 ( \75814 , \75808 );
buf \U$75880 ( \75815 , \75782 );
or \U$75881 ( \75816 , \75814 , \75815 );
nand \U$75882 ( \75817 , \75813 , \75816 );
buf \U$75883 ( \75818 , \75817 );
buf \U$75884 ( \75819 , \75818 );
buf \U$75885 ( \75820 , \49371 );
not \U$75886 ( \75821 , \75820 );
buf \U$75887 ( \75822 , \75672 );
not \U$75888 ( \75823 , \75822 );
or \U$75889 ( \75824 , \75821 , \75823 );
buf \U$75890 ( \75825 , \53405 );
not \U$75891 ( \75826 , \75825 );
buf \U$75892 ( \75827 , \75826 );
buf \U$75893 ( \75828 , \75827 );
nand \U$75894 ( \75829 , \75824 , \75828 );
buf \U$75895 ( \75830 , \75829 );
buf \U$75896 ( \75831 , \75830 );
buf \U$75897 ( \75832 , \48013 );
buf \U$75898 ( \75833 , \53414 );
nand \U$75899 ( \75834 , \75832 , \75833 );
buf \U$75900 ( \75835 , \75834 );
buf \U$75901 ( \75836 , \75835 );
not \U$75902 ( \75837 , \75836 );
buf \U$75903 ( \75838 , \75837 );
buf \U$75904 ( \75839 , \75838 );
and \U$75905 ( \75840 , \75831 , \75839 );
not \U$75906 ( \75841 , \75831 );
buf \U$75907 ( \75842 , \75835 );
and \U$75908 ( \75843 , \75841 , \75842 );
nor \U$75909 ( \75844 , \75840 , \75843 );
buf \U$75910 ( \75845 , \75844 );
buf \U$75911 ( \75846 , \75845 );
buf \U$75912 ( \75847 , \75827 );
buf \U$75913 ( \75848 , \49371 );
nand \U$75914 ( \75849 , \75847 , \75848 );
buf \U$75915 ( \75850 , \75849 );
buf \U$75916 ( \75851 , \75850 );
not \U$75917 ( \75852 , \75851 );
buf \U$75918 ( \75853 , \75672 );
not \U$75919 ( \75854 , \75853 );
or \U$75920 ( \75855 , \75852 , \75854 );
buf \U$75921 ( \75856 , \75850 );
buf \U$75922 ( \75857 , \75672 );
or \U$75923 ( \75858 , \75856 , \75857 );
nand \U$75924 ( \75859 , \75855 , \75858 );
buf \U$75925 ( \75860 , \75859 );
buf \U$75926 ( \75861 , \75860 );
buf \U$75927 ( \75862 , \51469 );
not \U$75928 ( \75863 , \75862 );
buf \U$75929 ( \75864 , \51433 );
not \U$75930 ( \75865 , \75864 );
buf \U$75931 ( \75866 , \56466 );
not \U$75932 ( \75867 , \75866 );
buf \U$75933 ( \75868 , \62972 );
not \U$75934 ( \75869 , \75868 );
or \U$75935 ( \75870 , \75867 , \75869 );
buf \U$75936 ( \75871 , \53326 );
nand \U$75937 ( \75872 , \75870 , \75871 );
buf \U$75938 ( \75873 , \75872 );
buf \U$75939 ( \75874 , \75873 );
not \U$75940 ( \75875 , \75874 );
or \U$75941 ( \75876 , \75865 , \75875 );
buf \U$75942 ( \75877 , \53355 );
not \U$75943 ( \75878 , \75877 );
buf \U$75944 ( \75879 , \75878 );
buf \U$75945 ( \75880 , \75879 );
nand \U$75946 ( \75881 , \75876 , \75880 );
buf \U$75947 ( \75882 , \75881 );
buf \U$75948 ( \75883 , \75882 );
not \U$75949 ( \75884 , \75883 );
or \U$75950 ( \75885 , \75863 , \75884 );
buf \U$75951 ( \75886 , \53367 );
nand \U$75952 ( \75887 , \75885 , \75886 );
buf \U$75953 ( \75888 , \75887 );
buf \U$75954 ( \75889 , \75888 );
buf \U$75955 ( \75890 , \53333 );
buf \U$75956 ( \75891 , \51489 );
nand \U$75957 ( \75892 , \75890 , \75891 );
buf \U$75958 ( \75893 , \75892 );
buf \U$75959 ( \75894 , \75893 );
not \U$75960 ( \75895 , \75894 );
buf \U$75961 ( \75896 , \75895 );
buf \U$75962 ( \75897 , \75896 );
and \U$75963 ( \75898 , \75889 , \75897 );
not \U$75964 ( \75899 , \75889 );
buf \U$75965 ( \75900 , \75893 );
and \U$75966 ( \75901 , \75899 , \75900 );
nor \U$75967 ( \75902 , \75898 , \75901 );
buf \U$75968 ( \75903 , \75902 );
buf \U$75969 ( \75904 , \75903 );
buf \U$75970 ( \75905 , \75882 );
not \U$75971 ( \75906 , \75905 );
buf \U$75972 ( \75907 , \51469 );
buf \U$75973 ( \75908 , \53367 );
nand \U$75974 ( \75909 , \75907 , \75908 );
buf \U$75975 ( \75910 , \75909 );
buf \U$75976 ( \75911 , \75910 );
not \U$75977 ( \75912 , \75911 );
or \U$75978 ( \75913 , \75906 , \75912 );
buf \U$75979 ( \75914 , \75910 );
buf \U$75980 ( \75915 , \75882 );
or \U$75981 ( \75916 , \75914 , \75915 );
nand \U$75982 ( \75917 , \75913 , \75916 );
buf \U$75983 ( \75918 , \75917 );
buf \U$75984 ( \75919 , \75918 );
buf \U$75985 ( \75920 , \51430 );
not \U$75986 ( \75921 , \75920 );
buf \U$75987 ( \75922 , \75873 );
not \U$75988 ( \75923 , \75922 );
or \U$75989 ( \75924 , \75921 , \75923 );
buf \U$75990 ( \75925 , \53343 );
not \U$75991 ( \75926 , \75925 );
buf \U$75992 ( \75927 , \75926 );
buf \U$75993 ( \75928 , \75927 );
nand \U$75994 ( \75929 , \75924 , \75928 );
buf \U$75995 ( \75930 , \75929 );
buf \U$75996 ( \75931 , \75930 );
buf \U$75997 ( \75932 , \50976 );
buf \U$75998 ( \75933 , \53352 );
nand \U$75999 ( \75934 , \75932 , \75933 );
buf \U$76000 ( \75935 , \75934 );
buf \U$76001 ( \75936 , \75935 );
not \U$76002 ( \75937 , \75936 );
buf \U$76003 ( \75938 , \75937 );
buf \U$76004 ( \75939 , \75938 );
and \U$76005 ( \75940 , \75931 , \75939 );
not \U$76006 ( \75941 , \75931 );
buf \U$76007 ( \75942 , \75935 );
and \U$76008 ( \75943 , \75941 , \75942 );
nor \U$76009 ( \75944 , \75940 , \75943 );
buf \U$76010 ( \75945 , \75944 );
buf \U$76011 ( \75946 , \75945 );
buf \U$76012 ( \75947 , \75927 );
buf \U$76013 ( \75948 , \51430 );
nand \U$76014 ( \75949 , \75947 , \75948 );
buf \U$76015 ( \75950 , \75949 );
buf \U$76016 ( \75951 , \75950 );
not \U$76017 ( \75952 , \75951 );
buf \U$76018 ( \75953 , \75873 );
not \U$76019 ( \75954 , \75953 );
or \U$76020 ( \75955 , \75952 , \75954 );
buf \U$76021 ( \75956 , \75950 );
buf \U$76022 ( \75957 , \75873 );
or \U$76023 ( \75958 , \75956 , \75957 );
nand \U$76024 ( \75959 , \75955 , \75958 );
buf \U$76025 ( \75960 , \75959 );
buf \U$76026 ( \75961 , \75960 );
buf \U$76027 ( \75962 , \53290 );
not \U$76028 ( \75963 , \75962 );
buf \U$76029 ( \75964 , \56461 );
not \U$76030 ( \75965 , \75964 );
buf \U$76031 ( \75966 , \62972 );
not \U$76032 ( \75967 , \75966 );
or \U$76033 ( \75968 , \75965 , \75967 );
buf \U$76034 ( \75969 , \53258 );
nand \U$76035 ( \75970 , \75968 , \75969 );
buf \U$76036 ( \75971 , \75970 );
buf \U$76037 ( \75972 , \75971 );
not \U$76038 ( \75973 , \75972 );
or \U$76039 ( \75974 , \75963 , \75973 );
buf \U$76040 ( \75975 , \53312 );
nand \U$76041 ( \75976 , \75974 , \75975 );
buf \U$76042 ( \75977 , \75976 );
buf \U$76043 ( \75978 , \75977 );
buf \U$76044 ( \75979 , \53323 );
buf \U$76045 ( \75980 , \53307 );
nand \U$76046 ( \75981 , \75979 , \75980 );
buf \U$76047 ( \75982 , \75981 );
buf \U$76048 ( \75983 , \75982 );
not \U$76049 ( \75984 , \75983 );
buf \U$76050 ( \75985 , \75984 );
buf \U$76051 ( \75986 , \75985 );
and \U$76052 ( \75987 , \75978 , \75986 );
not \U$76053 ( \75988 , \75978 );
buf \U$76054 ( \75989 , \75982 );
and \U$76055 ( \75990 , \75988 , \75989 );
nor \U$76056 ( \75991 , \75987 , \75990 );
buf \U$76057 ( \75992 , \75991 );
buf \U$76058 ( \75993 , \75992 );
buf \U$76059 ( \75994 , \53312 );
buf \U$76060 ( \75995 , \53290 );
nand \U$76061 ( \75996 , \75994 , \75995 );
buf \U$76062 ( \75997 , \75996 );
buf \U$76063 ( \75998 , \75997 );
not \U$76064 ( \75999 , \75998 );
buf \U$76065 ( \76000 , \75971 );
not \U$76066 ( \76001 , \76000 );
or \U$76067 ( \76002 , \75999 , \76001 );
buf \U$76068 ( \76003 , \75997 );
buf \U$76069 ( \76004 , \75971 );
or \U$76070 ( \76005 , \76003 , \76004 );
nand \U$76071 ( \76006 , \76002 , \76005 );
buf \U$76072 ( \76007 , \76006 );
buf \U$76073 ( \76008 , \76007 );
buf \U$76074 ( \76009 , \56458 );
not \U$76075 ( \76010 , \76009 );
buf \U$76076 ( \76011 , \62972 );
not \U$76077 ( \76012 , \76011 );
or \U$76078 ( \76013 , \76010 , \76012 );
buf \U$76079 ( \76014 , \53245 );
nand \U$76080 ( \76015 , \76013 , \76014 );
buf \U$76081 ( \76016 , \76015 );
buf \U$76082 ( \76017 , \76016 );
buf \U$76083 ( \76018 , \52867 );
buf \U$76084 ( \76019 , \53257 );
nand \U$76085 ( \76020 , \76018 , \76019 );
buf \U$76086 ( \76021 , \76020 );
buf \U$76087 ( \76022 , \76021 );
not \U$76088 ( \76023 , \76022 );
buf \U$76089 ( \76024 , \76023 );
buf \U$76090 ( \76025 , \76024 );
and \U$76091 ( \76026 , \76017 , \76025 );
not \U$76092 ( \76027 , \76017 );
buf \U$76093 ( \76028 , \76021 );
and \U$76094 ( \76029 , \76027 , \76028 );
nor \U$76095 ( \76030 , \76026 , \76029 );
buf \U$76096 ( \76031 , \76030 );
buf \U$76097 ( \76032 , \76031 );
buf \U$76098 ( \76033 , \62972 );
buf \U$76099 ( \76034 , \56458 );
buf \U$76100 ( \76035 , \53245 );
nand \U$76101 ( \76036 , \76034 , \76035 );
buf \U$76102 ( \76037 , \76036 );
buf \U$76103 ( \76038 , \76037 );
not \U$76104 ( \76039 , \76038 );
buf \U$76105 ( \76040 , \76039 );
buf \U$76106 ( \76041 , \76040 );
and \U$76107 ( \76042 , \76033 , \76041 );
not \U$76108 ( \76043 , \76033 );
buf \U$76109 ( \76044 , \76037 );
and \U$76110 ( \76045 , \76043 , \76044 );
nor \U$76111 ( \76046 , \76042 , \76045 );
buf \U$76112 ( \76047 , \76046 );
buf \U$76113 ( \76048 , \76047 );
buf \U$76114 ( \76049 , \57918 );
not \U$76115 ( \76050 , \76049 );
buf \U$76116 ( \76051 , \57859 );
not \U$76117 ( \76052 , \76051 );
buf \U$76118 ( \76053 , \59421 );
not \U$76119 ( \76054 , \76053 );
buf \U$76120 ( \76055 , \76054 );
buf \U$76121 ( \76056 , \76055 );
not \U$76122 ( \76057 , \76056 );
buf \U$76123 ( \76058 , \62880 );
not \U$76124 ( \76059 , \76058 );
or \U$76125 ( \76060 , \76057 , \76059 );
buf \U$76126 ( \76061 , \62923 );
not \U$76127 ( \76062 , \76061 );
buf \U$76128 ( \76063 , \76062 );
buf \U$76129 ( \76064 , \76063 );
nand \U$76130 ( \76065 , \76060 , \76064 );
buf \U$76131 ( \76066 , \76065 );
buf \U$76132 ( \76067 , \76066 );
not \U$76133 ( \76068 , \76067 );
or \U$76134 ( \76069 , \76052 , \76068 );
buf \U$76135 ( \76070 , \62943 );
not \U$76136 ( \76071 , \76070 );
buf \U$76137 ( \76072 , \76071 );
buf \U$76138 ( \76073 , \76072 );
nand \U$76139 ( \76074 , \76069 , \76073 );
buf \U$76140 ( \76075 , \76074 );
buf \U$76141 ( \76076 , \76075 );
not \U$76142 ( \76077 , \76076 );
or \U$76143 ( \76078 , \76050 , \76077 );
buf \U$76144 ( \76079 , \62954 );
not \U$76145 ( \76080 , \76079 );
buf \U$76146 ( \76081 , \76080 );
buf \U$76147 ( \76082 , \76081 );
nand \U$76148 ( \76083 , \76078 , \76082 );
buf \U$76149 ( \76084 , \76083 );
buf \U$76150 ( \76085 , \76084 );
buf \U$76151 ( \76086 , \62960 );
not \U$76152 ( \76087 , \76086 );
buf \U$76153 ( \76088 , \57943 );
nand \U$76154 ( \76089 , \76087 , \76088 );
buf \U$76155 ( \76090 , \76089 );
buf \U$76156 ( \76091 , \76090 );
not \U$76157 ( \76092 , \76091 );
buf \U$76158 ( \76093 , \76092 );
buf \U$76159 ( \76094 , \76093 );
and \U$76160 ( \76095 , \76085 , \76094 );
not \U$76161 ( \76096 , \76085 );
buf \U$76162 ( \76097 , \76090 );
and \U$76163 ( \76098 , \76096 , \76097 );
nor \U$76164 ( \76099 , \76095 , \76098 );
buf \U$76165 ( \76100 , \76099 );
buf \U$76166 ( \76101 , \76100 );
buf \U$76167 ( \76102 , \57918 );
buf \U$76168 ( \76103 , \76081 );
nand \U$76169 ( \76104 , \76102 , \76103 );
buf \U$76170 ( \76105 , \76104 );
buf \U$76171 ( \76106 , \76105 );
not \U$76172 ( \76107 , \76106 );
buf \U$76173 ( \76108 , \76075 );
not \U$76174 ( \76109 , \76108 );
or \U$76175 ( \76110 , \76107 , \76109 );
buf \U$76176 ( \76111 , \76105 );
buf \U$76177 ( \76112 , \76075 );
or \U$76178 ( \76113 , \76111 , \76112 );
nand \U$76179 ( \76114 , \76110 , \76113 );
buf \U$76180 ( \76115 , \76114 );
buf \U$76181 ( \76116 , \76115 );
buf \U$76182 ( \76117 , \57856 );
not \U$76183 ( \76118 , \76117 );
buf \U$76184 ( \76119 , \76066 );
not \U$76185 ( \76120 , \76119 );
or \U$76186 ( \76121 , \76118 , \76120 );
buf \U$76187 ( \76122 , \62929 );
nand \U$76188 ( \76123 , \76121 , \76122 );
buf \U$76189 ( \76124 , \76123 );
buf \U$76190 ( \76125 , \76124 );
buf \U$76191 ( \76126 , \57472 );
buf \U$76192 ( \76127 , \62940 );
nand \U$76193 ( \76128 , \76126 , \76127 );
buf \U$76194 ( \76129 , \76128 );
buf \U$76195 ( \76130 , \76129 );
not \U$76196 ( \76131 , \76130 );
buf \U$76197 ( \76132 , \76131 );
buf \U$76198 ( \76133 , \76132 );
and \U$76199 ( \76134 , \76125 , \76133 );
not \U$76200 ( \76135 , \76125 );
buf \U$76201 ( \76136 , \76129 );
and \U$76202 ( \76137 , \76135 , \76136 );
nor \U$76203 ( \76138 , \76134 , \76137 );
buf \U$76204 ( \76139 , \76138 );
buf \U$76205 ( \76140 , \76139 );
buf \U$76206 ( \76141 , \62929 );
buf \U$76207 ( \76142 , \57856 );
nand \U$76208 ( \76143 , \76141 , \76142 );
buf \U$76209 ( \76144 , \76143 );
buf \U$76210 ( \76145 , \76144 );
not \U$76211 ( \76146 , \76145 );
buf \U$76212 ( \76147 , \76066 );
not \U$76213 ( \76148 , \76147 );
or \U$76214 ( \76149 , \76146 , \76148 );
buf \U$76215 ( \76150 , \76144 );
buf \U$76216 ( \76151 , \76066 );
or \U$76217 ( \76152 , \76150 , \76151 );
nand \U$76218 ( \76153 , \76149 , \76152 );
buf \U$76219 ( \76154 , \76153 );
buf \U$76220 ( \76155 , \76154 );
buf \U$76221 ( \76156 , \58689 );
not \U$76222 ( \76157 , \76156 );
buf \U$76223 ( \76158 , \59418 );
not \U$76224 ( \76159 , \76158 );
buf \U$76225 ( \76160 , \62880 );
not \U$76226 ( \76161 , \76160 );
or \U$76227 ( \76162 , \76159 , \76161 );
buf \U$76228 ( \76163 , \62897 );
not \U$76229 ( \76164 , \76163 );
buf \U$76230 ( \76165 , \62909 );
not \U$76231 ( \76166 , \76165 );
buf \U$76232 ( \76167 , \76166 );
buf \U$76233 ( \76168 , \76167 );
nor \U$76234 ( \76169 , \76164 , \76168 );
buf \U$76235 ( \76170 , \76169 );
buf \U$76236 ( \76171 , \76170 );
nand \U$76237 ( \76172 , \76162 , \76171 );
buf \U$76238 ( \76173 , \76172 );
buf \U$76239 ( \76174 , \76173 );
not \U$76240 ( \76175 , \76174 );
or \U$76241 ( \76176 , \76157 , \76175 );
buf \U$76242 ( \76177 , \62903 );
nand \U$76243 ( \76178 , \76176 , \76177 );
buf \U$76244 ( \76179 , \76178 );
buf \U$76245 ( \76180 , \76179 );
buf \U$76246 ( \76181 , \62920 );
buf \U$76247 ( \76182 , \58718 );
nand \U$76248 ( \76183 , \76181 , \76182 );
buf \U$76249 ( \76184 , \76183 );
buf \U$76250 ( \76185 , \76184 );
not \U$76251 ( \76186 , \76185 );
buf \U$76252 ( \76187 , \76186 );
buf \U$76253 ( \76188 , \76187 );
and \U$76254 ( \76189 , \76180 , \76188 );
not \U$76255 ( \76190 , \76180 );
buf \U$76256 ( \76191 , \76184 );
and \U$76257 ( \76192 , \76190 , \76191 );
nor \U$76258 ( \76193 , \76189 , \76192 );
buf \U$76259 ( \76194 , \76193 );
buf \U$76260 ( \76195 , \76194 );
buf \U$76261 ( \76196 , \58689 );
buf \U$76262 ( \76197 , \62903 );
nand \U$76263 ( \76198 , \76196 , \76197 );
buf \U$76264 ( \76199 , \76198 );
buf \U$76265 ( \76200 , \76199 );
not \U$76266 ( \76201 , \76200 );
buf \U$76267 ( \76202 , \76173 );
not \U$76268 ( \76203 , \76202 );
or \U$76269 ( \76204 , \76201 , \76203 );
buf \U$76270 ( \76205 , \76199 );
buf \U$76271 ( \76206 , \76173 );
or \U$76272 ( \76207 , \76205 , \76206 );
nand \U$76273 ( \76208 , \76204 , \76207 );
buf \U$76274 ( \76209 , \76208 );
buf \U$76275 ( \76210 , \76209 );
buf \U$76276 ( \76211 , \59415 );
not \U$76277 ( \76212 , \76211 );
buf \U$76278 ( \76213 , \62880 );
not \U$76279 ( \76214 , \76213 );
or \U$76280 ( \76215 , \76212 , \76214 );
buf \U$76281 ( \76216 , \62894 );
not \U$76282 ( \76217 , \76216 );
buf \U$76283 ( \76218 , \76217 );
buf \U$76284 ( \76219 , \76218 );
nand \U$76285 ( \76220 , \76215 , \76219 );
buf \U$76286 ( \76221 , \76220 );
buf \U$76287 ( \76222 , \76221 );
buf \U$76288 ( \76223 , \58867 );
not \U$76289 ( \76224 , \76223 );
buf \U$76290 ( \76225 , \76167 );
nor \U$76291 ( \76226 , \76224 , \76225 );
buf \U$76292 ( \76227 , \76226 );
buf \U$76293 ( \76228 , \76227 );
and \U$76294 ( \76229 , \76222 , \76228 );
not \U$76295 ( \76230 , \76222 );
buf \U$76296 ( \76231 , \76227 );
not \U$76297 ( \76232 , \76231 );
buf \U$76298 ( \76233 , \76232 );
buf \U$76299 ( \76234 , \76233 );
and \U$76300 ( \76235 , \76230 , \76234 );
nor \U$76301 ( \76236 , \76229 , \76235 );
buf \U$76302 ( \76237 , \76236 );
buf \U$76303 ( \76238 , \76237 );
buf \U$76304 ( \76239 , \62880 );
buf \U$76305 ( \76240 , \76218 );
buf \U$76306 ( \76241 , \59415 );
nand \U$76307 ( \76242 , \76240 , \76241 );
buf \U$76308 ( \76243 , \76242 );
buf \U$76309 ( \76244 , \76243 );
not \U$76310 ( \76245 , \76244 );
buf \U$76311 ( \76246 , \76245 );
buf \U$76312 ( \76247 , \76246 );
and \U$76313 ( \76248 , \76239 , \76247 );
not \U$76314 ( \76249 , \76239 );
buf \U$76315 ( \76250 , \76243 );
and \U$76316 ( \76251 , \76249 , \76250 );
nor \U$76317 ( \76252 , \76248 , \76251 );
buf \U$76318 ( \76253 , \76252 );
buf \U$76319 ( \76254 , \76253 );
buf \U$76320 ( \76255 , \59745 );
not \U$76321 ( \76256 , \76255 );
buf \U$76322 ( \76257 , \62861 );
not \U$76323 ( \76258 , \76257 );
buf \U$76324 ( \76259 , \76258 );
buf \U$76325 ( \76260 , \76259 );
not \U$76326 ( \76261 , \76260 );
buf \U$76327 ( \76262 , \62852 );
not \U$76328 ( \76263 , \76262 );
or \U$76329 ( \76264 , \76261 , \76263 );
buf \U$76330 ( \76265 , \60294 );
not \U$76331 ( \76266 , \76265 );
buf \U$76332 ( \76267 , \76266 );
buf \U$76333 ( \76268 , \76267 );
nand \U$76334 ( \76269 , \76264 , \76268 );
buf \U$76335 ( \76270 , \76269 );
buf \U$76336 ( \76271 , \76270 );
not \U$76337 ( \76272 , \76271 );
or \U$76338 ( \76273 , \76256 , \76272 );
buf \U$76339 ( \76274 , \60301 );
nand \U$76340 ( \76275 , \76273 , \76274 );
buf \U$76341 ( \76276 , \76275 );
buf \U$76342 ( \76277 , \76276 );
buf \U$76343 ( \76278 , \62877 );
buf \U$76344 ( \76279 , \60331 );
nand \U$76345 ( \76280 , \76278 , \76279 );
buf \U$76346 ( \76281 , \76280 );
buf \U$76347 ( \76282 , \76281 );
xnor \U$76348 ( \76283 , \76277 , \76282 );
buf \U$76349 ( \76284 , \76283 );
buf \U$76350 ( \76285 , \76284 );
buf \U$76351 ( \76286 , \60301 );
buf \U$76352 ( \76287 , \59745 );
nand \U$76353 ( \76288 , \76286 , \76287 );
buf \U$76354 ( \76289 , \76288 );
buf \U$76355 ( \76290 , \76289 );
not \U$76356 ( \76291 , \76290 );
buf \U$76357 ( \76292 , \76270 );
not \U$76358 ( \76293 , \76292 );
or \U$76359 ( \76294 , \76291 , \76293 );
buf \U$76360 ( \76295 , \76289 );
buf \U$76361 ( \76296 , \76270 );
or \U$76362 ( \76297 , \76295 , \76296 );
nand \U$76363 ( \76298 , \76294 , \76297 );
buf \U$76364 ( \76299 , \76298 );
buf \U$76365 ( \76300 , \76299 );
buf \U$76366 ( \76301 , \62857 );
not \U$76367 ( \76302 , \76301 );
buf \U$76368 ( \76303 , \62852 );
not \U$76369 ( \76304 , \76303 );
or \U$76370 ( \76305 , \76302 , \76304 );
buf \U$76371 ( \76306 , \60264 );
nand \U$76372 ( \76307 , \76305 , \76306 );
buf \U$76373 ( \76308 , \76307 );
buf \U$76374 ( \76309 , \76308 );
buf \U$76375 ( \76310 , \60291 );
buf \U$76376 ( \76311 , \60282 );
nand \U$76377 ( \76312 , \76310 , \76311 );
buf \U$76378 ( \76313 , \76312 );
buf \U$76379 ( \76314 , \76313 );
xnor \U$76380 ( \76315 , \76309 , \76314 );
buf \U$76381 ( \76316 , \76315 );
buf \U$76382 ( \76317 , \76316 );
buf \U$76383 ( \76318 , \62852 );
buf \U$76384 ( \76319 , \62857 );
buf \U$76385 ( \76320 , \60264 );
nand \U$76386 ( \76321 , \76319 , \76320 );
buf \U$76387 ( \76322 , \76321 );
buf \U$76388 ( \76323 , \76322 );
xnor \U$76389 ( \76324 , \76318 , \76323 );
buf \U$76390 ( \76325 , \76324 );
buf \U$76391 ( \76326 , \76325 );
buf \U$76392 ( \76327 , \60768 );
buf \U$76393 ( \76328 , \62805 );
not \U$76394 ( \76329 , \76328 );
buf \U$76395 ( \76330 , \62731 );
not \U$76396 ( \76331 , \76330 );
or \U$76397 ( \76332 , \76329 , \76331 );
buf \U$76398 ( \76333 , \62827 );
not \U$76399 ( \76334 , \76333 );
buf \U$76400 ( \76335 , \76334 );
buf \U$76401 ( \76336 , \76335 );
nand \U$76402 ( \76337 , \76332 , \76336 );
buf \U$76403 ( \76338 , \76337 );
buf \U$76404 ( \76339 , \76338 );
nand \U$76405 ( \76340 , \76327 , \76339 );
buf \U$76406 ( \76341 , \76340 );
buf \U$76407 ( \76342 , \76341 );
buf \U$76408 ( \76343 , \62835 );
nand \U$76409 ( \76344 , \76342 , \76343 );
buf \U$76410 ( \76345 , \76344 );
buf \U$76411 ( \76346 , \76345 );
buf \U$76412 ( \76347 , \60588 );
buf \U$76413 ( \76348 , \62846 );
nand \U$76414 ( \76349 , \76347 , \76348 );
buf \U$76415 ( \76350 , \76349 );
buf \U$76416 ( \76351 , \76350 );
xnor \U$76417 ( \76352 , \76346 , \76351 );
buf \U$76418 ( \76353 , \76352 );
buf \U$76419 ( \76354 , \76353 );
buf \U$76420 ( \76355 , \62835 );
buf \U$76421 ( \76356 , \60768 );
nand \U$76422 ( \76357 , \76355 , \76356 );
buf \U$76423 ( \76358 , \76357 );
buf \U$76424 ( \76359 , \76358 );
not \U$76425 ( \76360 , \76359 );
buf \U$76426 ( \76361 , \76338 );
not \U$76427 ( \76362 , \76361 );
or \U$76428 ( \76363 , \76360 , \76362 );
buf \U$76429 ( \76364 , \76358 );
buf \U$76430 ( \76365 , \76338 );
or \U$76431 ( \76366 , \76364 , \76365 );
nand \U$76432 ( \76367 , \76363 , \76366 );
buf \U$76433 ( \76368 , \76367 );
buf \U$76434 ( \76369 , \76368 );
buf \U$76435 ( \76370 , \62773 );
buf \U$76436 ( \76371 , \62824 );
nand \U$76437 ( \76372 , \76370 , \76371 );
buf \U$76438 ( \76373 , \76372 );
buf \U$76439 ( \76374 , \76373 );
not \U$76440 ( \76375 , \76374 );
buf \U$76441 ( \76376 , \62802 );
not \U$76442 ( \76377 , \76376 );
buf \U$76443 ( \76378 , \62731 );
not \U$76444 ( \76379 , \76378 );
or \U$76445 ( \76380 , \76377 , \76379 );
buf \U$76446 ( \76381 , \62814 );
nand \U$76447 ( \76382 , \76380 , \76381 );
buf \U$76448 ( \76383 , \76382 );
buf \U$76449 ( \76384 , \76383 );
not \U$76450 ( \76385 , \76384 );
or \U$76451 ( \76386 , \76375 , \76385 );
buf \U$76452 ( \76387 , \76373 );
buf \U$76453 ( \76388 , \76383 );
or \U$76454 ( \76389 , \76387 , \76388 );
nand \U$76455 ( \76390 , \76386 , \76389 );
buf \U$76456 ( \76391 , \76390 );
buf \U$76457 ( \76392 , \76391 );
buf \U$76458 ( \76393 , \62814 );
buf \U$76459 ( \76394 , \62802 );
nand \U$76460 ( \76395 , \76393 , \76394 );
buf \U$76461 ( \76396 , \76395 );
buf \U$76462 ( \76397 , \76396 );
not \U$76463 ( \76398 , \76397 );
buf \U$76464 ( \76399 , \62731 );
not \U$76465 ( \76400 , \76399 );
or \U$76466 ( \76401 , \76398 , \76400 );
buf \U$76467 ( \76402 , \76396 );
buf \U$76468 ( \76403 , \62731 );
or \U$76469 ( \76404 , \76402 , \76403 );
nand \U$76470 ( \76405 , \76401 , \76404 );
buf \U$76471 ( \76406 , \76405 );
buf \U$76472 ( \76407 , \76406 );
buf \U$76473 ( \76408 , \61843 );
buf \U$76474 ( \76409 , \62728 );
nand \U$76475 ( \76410 , \76408 , \76409 );
buf \U$76476 ( \76411 , \76410 );
buf \U$76477 ( \76412 , \76411 );
not \U$76478 ( \76413 , \76412 );
buf \U$76481 ( \76414 , \62703 );
buf \U$76482 ( \76415 , \76414 );
buf \U$76483 ( \76416 , \62715 );
not \U$76484 ( \76417 , \76416 );
buf \U$76485 ( \76418 , \76417 );
buf \U$76486 ( \76419 , \76418 );
and \U$76487 ( \76420 , \76415 , \76419 );
buf \U$76488 ( \76421 , \61635 );
nor \U$76489 ( \76422 , \76420 , \76421 );
buf \U$76490 ( \76423 , \76422 );
buf \U$76491 ( \76424 , \76423 );
not \U$76492 ( \76425 , \76424 );
buf \U$76493 ( \76426 , \61767 );
nand \U$76494 ( \76427 , \76425 , \76426 );
buf \U$76495 ( \76428 , \76427 );
buf \U$76496 ( \76429 , \76428 );
buf \U$76497 ( \76430 , \61775 );
nand \U$76498 ( \76431 , \76429 , \76430 );
buf \U$76499 ( \76432 , \76431 );
buf \U$76500 ( \76433 , \76432 );
not \U$76501 ( \76434 , \76433 );
or \U$76502 ( \76435 , \76413 , \76434 );
buf \U$76503 ( \76436 , \76411 );
buf \U$76504 ( \76437 , \76432 );
or \U$76505 ( \76438 , \76436 , \76437 );
nand \U$76506 ( \76439 , \76435 , \76438 );
buf \U$76507 ( \76440 , \76439 );
buf \U$76508 ( \76441 , \76440 );
buf \U$76509 ( \76442 , \61775 );
buf \U$76510 ( \76443 , \61767 );
and \U$76511 ( \76444 , \76442 , \76443 );
buf \U$76512 ( \76445 , \76444 );
buf \U$76513 ( \76446 , \76445 );
not \U$76514 ( \76447 , \76446 );
buf \U$76515 ( \76448 , \76423 );
not \U$76516 ( \76449 , \76448 );
or \U$76517 ( \76450 , \76447 , \76449 );
buf \U$76518 ( \76451 , \76445 );
buf \U$76519 ( \76452 , \76423 );
or \U$76520 ( \76453 , \76451 , \76452 );
nand \U$76521 ( \76454 , \76450 , \76453 );
buf \U$76522 ( \76455 , \76454 );
buf \U$76523 ( \76456 , \76455 );
buf \U$76524 ( \76457 , \61632 );
buf \U$76525 ( \76458 , \61468 );
nand \U$76526 ( \76459 , \76457 , \76458 );
buf \U$76527 ( \76460 , \76459 );
buf \U$76528 ( \76461 , \76460 );
not \U$76529 ( \76462 , \76461 );
buf \U$76530 ( \76463 , \62712 );
not \U$76531 ( \76464 , \76463 );
buf \U$76532 ( \76465 , \76414 );
not \U$76533 ( \76466 , \76465 );
or \U$76534 ( \76467 , \76464 , \76466 );
buf \U$76535 ( \76468 , \61623 );
not \U$76536 ( \76469 , \76468 );
buf \U$76537 ( \76470 , \76469 );
buf \U$76538 ( \76471 , \76470 );
nand \U$76539 ( \76472 , \76467 , \76471 );
buf \U$76540 ( \76473 , \76472 );
buf \U$76541 ( \76474 , \76473 );
not \U$76542 ( \76475 , \76474 );
or \U$76543 ( \76476 , \76462 , \76475 );
buf \U$76544 ( \76477 , \76460 );
buf \U$76545 ( \76478 , \76473 );
or \U$76546 ( \76479 , \76477 , \76478 );
nand \U$76547 ( \76480 , \76476 , \76479 );
buf \U$76548 ( \76481 , \76480 );
buf \U$76549 ( \76482 , \76481 );
endmodule

